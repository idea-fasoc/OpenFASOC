* NGSPICE file created from diff_pair_sample_0104.ext - technology: sky130A

.subckt diff_pair_sample_0104 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1097 pd=37.24 as=7.1097 ps=37.24 w=18.23 l=3.89
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1097 pd=37.24 as=0 ps=0 w=18.23 l=3.89
X2 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.1097 pd=37.24 as=7.1097 ps=37.24 w=18.23 l=3.89
X3 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1097 pd=37.24 as=7.1097 ps=37.24 w=18.23 l=3.89
X4 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.1097 pd=37.24 as=0 ps=0 w=18.23 l=3.89
X5 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=7.1097 pd=37.24 as=7.1097 ps=37.24 w=18.23 l=3.89
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.1097 pd=37.24 as=0 ps=0 w=18.23 l=3.89
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1097 pd=37.24 as=0 ps=0 w=18.23 l=3.89
R0 VN VN.t1 200.589
R1 VN VN.t0 148.6
R2 VTAIL.n402 VTAIL.n306 289.615
R3 VTAIL.n96 VTAIL.n0 289.615
R4 VTAIL.n300 VTAIL.n204 289.615
R5 VTAIL.n198 VTAIL.n102 289.615
R6 VTAIL.n338 VTAIL.n337 185
R7 VTAIL.n343 VTAIL.n342 185
R8 VTAIL.n345 VTAIL.n344 185
R9 VTAIL.n334 VTAIL.n333 185
R10 VTAIL.n351 VTAIL.n350 185
R11 VTAIL.n353 VTAIL.n352 185
R12 VTAIL.n330 VTAIL.n329 185
R13 VTAIL.n359 VTAIL.n358 185
R14 VTAIL.n361 VTAIL.n360 185
R15 VTAIL.n326 VTAIL.n325 185
R16 VTAIL.n367 VTAIL.n366 185
R17 VTAIL.n369 VTAIL.n368 185
R18 VTAIL.n322 VTAIL.n321 185
R19 VTAIL.n375 VTAIL.n374 185
R20 VTAIL.n377 VTAIL.n376 185
R21 VTAIL.n318 VTAIL.n317 185
R22 VTAIL.n384 VTAIL.n383 185
R23 VTAIL.n385 VTAIL.n316 185
R24 VTAIL.n387 VTAIL.n386 185
R25 VTAIL.n314 VTAIL.n313 185
R26 VTAIL.n393 VTAIL.n392 185
R27 VTAIL.n395 VTAIL.n394 185
R28 VTAIL.n310 VTAIL.n309 185
R29 VTAIL.n401 VTAIL.n400 185
R30 VTAIL.n403 VTAIL.n402 185
R31 VTAIL.n32 VTAIL.n31 185
R32 VTAIL.n37 VTAIL.n36 185
R33 VTAIL.n39 VTAIL.n38 185
R34 VTAIL.n28 VTAIL.n27 185
R35 VTAIL.n45 VTAIL.n44 185
R36 VTAIL.n47 VTAIL.n46 185
R37 VTAIL.n24 VTAIL.n23 185
R38 VTAIL.n53 VTAIL.n52 185
R39 VTAIL.n55 VTAIL.n54 185
R40 VTAIL.n20 VTAIL.n19 185
R41 VTAIL.n61 VTAIL.n60 185
R42 VTAIL.n63 VTAIL.n62 185
R43 VTAIL.n16 VTAIL.n15 185
R44 VTAIL.n69 VTAIL.n68 185
R45 VTAIL.n71 VTAIL.n70 185
R46 VTAIL.n12 VTAIL.n11 185
R47 VTAIL.n78 VTAIL.n77 185
R48 VTAIL.n79 VTAIL.n10 185
R49 VTAIL.n81 VTAIL.n80 185
R50 VTAIL.n8 VTAIL.n7 185
R51 VTAIL.n87 VTAIL.n86 185
R52 VTAIL.n89 VTAIL.n88 185
R53 VTAIL.n4 VTAIL.n3 185
R54 VTAIL.n95 VTAIL.n94 185
R55 VTAIL.n97 VTAIL.n96 185
R56 VTAIL.n301 VTAIL.n300 185
R57 VTAIL.n299 VTAIL.n298 185
R58 VTAIL.n208 VTAIL.n207 185
R59 VTAIL.n293 VTAIL.n292 185
R60 VTAIL.n291 VTAIL.n290 185
R61 VTAIL.n212 VTAIL.n211 185
R62 VTAIL.n285 VTAIL.n284 185
R63 VTAIL.n283 VTAIL.n214 185
R64 VTAIL.n282 VTAIL.n281 185
R65 VTAIL.n217 VTAIL.n215 185
R66 VTAIL.n276 VTAIL.n275 185
R67 VTAIL.n274 VTAIL.n273 185
R68 VTAIL.n221 VTAIL.n220 185
R69 VTAIL.n268 VTAIL.n267 185
R70 VTAIL.n266 VTAIL.n265 185
R71 VTAIL.n225 VTAIL.n224 185
R72 VTAIL.n260 VTAIL.n259 185
R73 VTAIL.n258 VTAIL.n257 185
R74 VTAIL.n229 VTAIL.n228 185
R75 VTAIL.n252 VTAIL.n251 185
R76 VTAIL.n250 VTAIL.n249 185
R77 VTAIL.n233 VTAIL.n232 185
R78 VTAIL.n244 VTAIL.n243 185
R79 VTAIL.n242 VTAIL.n241 185
R80 VTAIL.n237 VTAIL.n236 185
R81 VTAIL.n199 VTAIL.n198 185
R82 VTAIL.n197 VTAIL.n196 185
R83 VTAIL.n106 VTAIL.n105 185
R84 VTAIL.n191 VTAIL.n190 185
R85 VTAIL.n189 VTAIL.n188 185
R86 VTAIL.n110 VTAIL.n109 185
R87 VTAIL.n183 VTAIL.n182 185
R88 VTAIL.n181 VTAIL.n112 185
R89 VTAIL.n180 VTAIL.n179 185
R90 VTAIL.n115 VTAIL.n113 185
R91 VTAIL.n174 VTAIL.n173 185
R92 VTAIL.n172 VTAIL.n171 185
R93 VTAIL.n119 VTAIL.n118 185
R94 VTAIL.n166 VTAIL.n165 185
R95 VTAIL.n164 VTAIL.n163 185
R96 VTAIL.n123 VTAIL.n122 185
R97 VTAIL.n158 VTAIL.n157 185
R98 VTAIL.n156 VTAIL.n155 185
R99 VTAIL.n127 VTAIL.n126 185
R100 VTAIL.n150 VTAIL.n149 185
R101 VTAIL.n148 VTAIL.n147 185
R102 VTAIL.n131 VTAIL.n130 185
R103 VTAIL.n142 VTAIL.n141 185
R104 VTAIL.n140 VTAIL.n139 185
R105 VTAIL.n135 VTAIL.n134 185
R106 VTAIL.n339 VTAIL.t3 147.659
R107 VTAIL.n33 VTAIL.t0 147.659
R108 VTAIL.n238 VTAIL.t1 147.659
R109 VTAIL.n136 VTAIL.t2 147.659
R110 VTAIL.n343 VTAIL.n337 104.615
R111 VTAIL.n344 VTAIL.n343 104.615
R112 VTAIL.n344 VTAIL.n333 104.615
R113 VTAIL.n351 VTAIL.n333 104.615
R114 VTAIL.n352 VTAIL.n351 104.615
R115 VTAIL.n352 VTAIL.n329 104.615
R116 VTAIL.n359 VTAIL.n329 104.615
R117 VTAIL.n360 VTAIL.n359 104.615
R118 VTAIL.n360 VTAIL.n325 104.615
R119 VTAIL.n367 VTAIL.n325 104.615
R120 VTAIL.n368 VTAIL.n367 104.615
R121 VTAIL.n368 VTAIL.n321 104.615
R122 VTAIL.n375 VTAIL.n321 104.615
R123 VTAIL.n376 VTAIL.n375 104.615
R124 VTAIL.n376 VTAIL.n317 104.615
R125 VTAIL.n384 VTAIL.n317 104.615
R126 VTAIL.n385 VTAIL.n384 104.615
R127 VTAIL.n386 VTAIL.n385 104.615
R128 VTAIL.n386 VTAIL.n313 104.615
R129 VTAIL.n393 VTAIL.n313 104.615
R130 VTAIL.n394 VTAIL.n393 104.615
R131 VTAIL.n394 VTAIL.n309 104.615
R132 VTAIL.n401 VTAIL.n309 104.615
R133 VTAIL.n402 VTAIL.n401 104.615
R134 VTAIL.n37 VTAIL.n31 104.615
R135 VTAIL.n38 VTAIL.n37 104.615
R136 VTAIL.n38 VTAIL.n27 104.615
R137 VTAIL.n45 VTAIL.n27 104.615
R138 VTAIL.n46 VTAIL.n45 104.615
R139 VTAIL.n46 VTAIL.n23 104.615
R140 VTAIL.n53 VTAIL.n23 104.615
R141 VTAIL.n54 VTAIL.n53 104.615
R142 VTAIL.n54 VTAIL.n19 104.615
R143 VTAIL.n61 VTAIL.n19 104.615
R144 VTAIL.n62 VTAIL.n61 104.615
R145 VTAIL.n62 VTAIL.n15 104.615
R146 VTAIL.n69 VTAIL.n15 104.615
R147 VTAIL.n70 VTAIL.n69 104.615
R148 VTAIL.n70 VTAIL.n11 104.615
R149 VTAIL.n78 VTAIL.n11 104.615
R150 VTAIL.n79 VTAIL.n78 104.615
R151 VTAIL.n80 VTAIL.n79 104.615
R152 VTAIL.n80 VTAIL.n7 104.615
R153 VTAIL.n87 VTAIL.n7 104.615
R154 VTAIL.n88 VTAIL.n87 104.615
R155 VTAIL.n88 VTAIL.n3 104.615
R156 VTAIL.n95 VTAIL.n3 104.615
R157 VTAIL.n96 VTAIL.n95 104.615
R158 VTAIL.n300 VTAIL.n299 104.615
R159 VTAIL.n299 VTAIL.n207 104.615
R160 VTAIL.n292 VTAIL.n207 104.615
R161 VTAIL.n292 VTAIL.n291 104.615
R162 VTAIL.n291 VTAIL.n211 104.615
R163 VTAIL.n284 VTAIL.n211 104.615
R164 VTAIL.n284 VTAIL.n283 104.615
R165 VTAIL.n283 VTAIL.n282 104.615
R166 VTAIL.n282 VTAIL.n215 104.615
R167 VTAIL.n275 VTAIL.n215 104.615
R168 VTAIL.n275 VTAIL.n274 104.615
R169 VTAIL.n274 VTAIL.n220 104.615
R170 VTAIL.n267 VTAIL.n220 104.615
R171 VTAIL.n267 VTAIL.n266 104.615
R172 VTAIL.n266 VTAIL.n224 104.615
R173 VTAIL.n259 VTAIL.n224 104.615
R174 VTAIL.n259 VTAIL.n258 104.615
R175 VTAIL.n258 VTAIL.n228 104.615
R176 VTAIL.n251 VTAIL.n228 104.615
R177 VTAIL.n251 VTAIL.n250 104.615
R178 VTAIL.n250 VTAIL.n232 104.615
R179 VTAIL.n243 VTAIL.n232 104.615
R180 VTAIL.n243 VTAIL.n242 104.615
R181 VTAIL.n242 VTAIL.n236 104.615
R182 VTAIL.n198 VTAIL.n197 104.615
R183 VTAIL.n197 VTAIL.n105 104.615
R184 VTAIL.n190 VTAIL.n105 104.615
R185 VTAIL.n190 VTAIL.n189 104.615
R186 VTAIL.n189 VTAIL.n109 104.615
R187 VTAIL.n182 VTAIL.n109 104.615
R188 VTAIL.n182 VTAIL.n181 104.615
R189 VTAIL.n181 VTAIL.n180 104.615
R190 VTAIL.n180 VTAIL.n113 104.615
R191 VTAIL.n173 VTAIL.n113 104.615
R192 VTAIL.n173 VTAIL.n172 104.615
R193 VTAIL.n172 VTAIL.n118 104.615
R194 VTAIL.n165 VTAIL.n118 104.615
R195 VTAIL.n165 VTAIL.n164 104.615
R196 VTAIL.n164 VTAIL.n122 104.615
R197 VTAIL.n157 VTAIL.n122 104.615
R198 VTAIL.n157 VTAIL.n156 104.615
R199 VTAIL.n156 VTAIL.n126 104.615
R200 VTAIL.n149 VTAIL.n126 104.615
R201 VTAIL.n149 VTAIL.n148 104.615
R202 VTAIL.n148 VTAIL.n130 104.615
R203 VTAIL.n141 VTAIL.n130 104.615
R204 VTAIL.n141 VTAIL.n140 104.615
R205 VTAIL.n140 VTAIL.n134 104.615
R206 VTAIL.t3 VTAIL.n337 52.3082
R207 VTAIL.t0 VTAIL.n31 52.3082
R208 VTAIL.t1 VTAIL.n236 52.3082
R209 VTAIL.t2 VTAIL.n134 52.3082
R210 VTAIL.n203 VTAIL.n101 35.3583
R211 VTAIL.n407 VTAIL.n406 31.9914
R212 VTAIL.n101 VTAIL.n100 31.9914
R213 VTAIL.n305 VTAIL.n304 31.9914
R214 VTAIL.n203 VTAIL.n202 31.9914
R215 VTAIL.n407 VTAIL.n305 31.7203
R216 VTAIL.n339 VTAIL.n338 15.6677
R217 VTAIL.n33 VTAIL.n32 15.6677
R218 VTAIL.n238 VTAIL.n237 15.6677
R219 VTAIL.n136 VTAIL.n135 15.6677
R220 VTAIL.n387 VTAIL.n316 13.1884
R221 VTAIL.n81 VTAIL.n10 13.1884
R222 VTAIL.n285 VTAIL.n214 13.1884
R223 VTAIL.n183 VTAIL.n112 13.1884
R224 VTAIL.n342 VTAIL.n341 12.8005
R225 VTAIL.n383 VTAIL.n382 12.8005
R226 VTAIL.n388 VTAIL.n314 12.8005
R227 VTAIL.n36 VTAIL.n35 12.8005
R228 VTAIL.n77 VTAIL.n76 12.8005
R229 VTAIL.n82 VTAIL.n8 12.8005
R230 VTAIL.n286 VTAIL.n212 12.8005
R231 VTAIL.n281 VTAIL.n216 12.8005
R232 VTAIL.n241 VTAIL.n240 12.8005
R233 VTAIL.n184 VTAIL.n110 12.8005
R234 VTAIL.n179 VTAIL.n114 12.8005
R235 VTAIL.n139 VTAIL.n138 12.8005
R236 VTAIL.n345 VTAIL.n336 12.0247
R237 VTAIL.n381 VTAIL.n318 12.0247
R238 VTAIL.n392 VTAIL.n391 12.0247
R239 VTAIL.n39 VTAIL.n30 12.0247
R240 VTAIL.n75 VTAIL.n12 12.0247
R241 VTAIL.n86 VTAIL.n85 12.0247
R242 VTAIL.n290 VTAIL.n289 12.0247
R243 VTAIL.n280 VTAIL.n217 12.0247
R244 VTAIL.n244 VTAIL.n235 12.0247
R245 VTAIL.n188 VTAIL.n187 12.0247
R246 VTAIL.n178 VTAIL.n115 12.0247
R247 VTAIL.n142 VTAIL.n133 12.0247
R248 VTAIL.n346 VTAIL.n334 11.249
R249 VTAIL.n378 VTAIL.n377 11.249
R250 VTAIL.n395 VTAIL.n312 11.249
R251 VTAIL.n40 VTAIL.n28 11.249
R252 VTAIL.n72 VTAIL.n71 11.249
R253 VTAIL.n89 VTAIL.n6 11.249
R254 VTAIL.n293 VTAIL.n210 11.249
R255 VTAIL.n277 VTAIL.n276 11.249
R256 VTAIL.n245 VTAIL.n233 11.249
R257 VTAIL.n191 VTAIL.n108 11.249
R258 VTAIL.n175 VTAIL.n174 11.249
R259 VTAIL.n143 VTAIL.n131 11.249
R260 VTAIL.n350 VTAIL.n349 10.4732
R261 VTAIL.n374 VTAIL.n320 10.4732
R262 VTAIL.n396 VTAIL.n310 10.4732
R263 VTAIL.n44 VTAIL.n43 10.4732
R264 VTAIL.n68 VTAIL.n14 10.4732
R265 VTAIL.n90 VTAIL.n4 10.4732
R266 VTAIL.n294 VTAIL.n208 10.4732
R267 VTAIL.n273 VTAIL.n219 10.4732
R268 VTAIL.n249 VTAIL.n248 10.4732
R269 VTAIL.n192 VTAIL.n106 10.4732
R270 VTAIL.n171 VTAIL.n117 10.4732
R271 VTAIL.n147 VTAIL.n146 10.4732
R272 VTAIL.n353 VTAIL.n332 9.69747
R273 VTAIL.n373 VTAIL.n322 9.69747
R274 VTAIL.n400 VTAIL.n399 9.69747
R275 VTAIL.n47 VTAIL.n26 9.69747
R276 VTAIL.n67 VTAIL.n16 9.69747
R277 VTAIL.n94 VTAIL.n93 9.69747
R278 VTAIL.n298 VTAIL.n297 9.69747
R279 VTAIL.n272 VTAIL.n221 9.69747
R280 VTAIL.n252 VTAIL.n231 9.69747
R281 VTAIL.n196 VTAIL.n195 9.69747
R282 VTAIL.n170 VTAIL.n119 9.69747
R283 VTAIL.n150 VTAIL.n129 9.69747
R284 VTAIL.n406 VTAIL.n405 9.45567
R285 VTAIL.n100 VTAIL.n99 9.45567
R286 VTAIL.n304 VTAIL.n303 9.45567
R287 VTAIL.n202 VTAIL.n201 9.45567
R288 VTAIL.n405 VTAIL.n404 9.3005
R289 VTAIL.n308 VTAIL.n307 9.3005
R290 VTAIL.n399 VTAIL.n398 9.3005
R291 VTAIL.n397 VTAIL.n396 9.3005
R292 VTAIL.n312 VTAIL.n311 9.3005
R293 VTAIL.n391 VTAIL.n390 9.3005
R294 VTAIL.n389 VTAIL.n388 9.3005
R295 VTAIL.n328 VTAIL.n327 9.3005
R296 VTAIL.n357 VTAIL.n356 9.3005
R297 VTAIL.n355 VTAIL.n354 9.3005
R298 VTAIL.n332 VTAIL.n331 9.3005
R299 VTAIL.n349 VTAIL.n348 9.3005
R300 VTAIL.n347 VTAIL.n346 9.3005
R301 VTAIL.n336 VTAIL.n335 9.3005
R302 VTAIL.n341 VTAIL.n340 9.3005
R303 VTAIL.n363 VTAIL.n362 9.3005
R304 VTAIL.n365 VTAIL.n364 9.3005
R305 VTAIL.n324 VTAIL.n323 9.3005
R306 VTAIL.n371 VTAIL.n370 9.3005
R307 VTAIL.n373 VTAIL.n372 9.3005
R308 VTAIL.n320 VTAIL.n319 9.3005
R309 VTAIL.n379 VTAIL.n378 9.3005
R310 VTAIL.n381 VTAIL.n380 9.3005
R311 VTAIL.n382 VTAIL.n315 9.3005
R312 VTAIL.n99 VTAIL.n98 9.3005
R313 VTAIL.n2 VTAIL.n1 9.3005
R314 VTAIL.n93 VTAIL.n92 9.3005
R315 VTAIL.n91 VTAIL.n90 9.3005
R316 VTAIL.n6 VTAIL.n5 9.3005
R317 VTAIL.n85 VTAIL.n84 9.3005
R318 VTAIL.n83 VTAIL.n82 9.3005
R319 VTAIL.n22 VTAIL.n21 9.3005
R320 VTAIL.n51 VTAIL.n50 9.3005
R321 VTAIL.n49 VTAIL.n48 9.3005
R322 VTAIL.n26 VTAIL.n25 9.3005
R323 VTAIL.n43 VTAIL.n42 9.3005
R324 VTAIL.n41 VTAIL.n40 9.3005
R325 VTAIL.n30 VTAIL.n29 9.3005
R326 VTAIL.n35 VTAIL.n34 9.3005
R327 VTAIL.n57 VTAIL.n56 9.3005
R328 VTAIL.n59 VTAIL.n58 9.3005
R329 VTAIL.n18 VTAIL.n17 9.3005
R330 VTAIL.n65 VTAIL.n64 9.3005
R331 VTAIL.n67 VTAIL.n66 9.3005
R332 VTAIL.n14 VTAIL.n13 9.3005
R333 VTAIL.n73 VTAIL.n72 9.3005
R334 VTAIL.n75 VTAIL.n74 9.3005
R335 VTAIL.n76 VTAIL.n9 9.3005
R336 VTAIL.n264 VTAIL.n263 9.3005
R337 VTAIL.n223 VTAIL.n222 9.3005
R338 VTAIL.n270 VTAIL.n269 9.3005
R339 VTAIL.n272 VTAIL.n271 9.3005
R340 VTAIL.n219 VTAIL.n218 9.3005
R341 VTAIL.n278 VTAIL.n277 9.3005
R342 VTAIL.n280 VTAIL.n279 9.3005
R343 VTAIL.n216 VTAIL.n213 9.3005
R344 VTAIL.n303 VTAIL.n302 9.3005
R345 VTAIL.n206 VTAIL.n205 9.3005
R346 VTAIL.n297 VTAIL.n296 9.3005
R347 VTAIL.n295 VTAIL.n294 9.3005
R348 VTAIL.n210 VTAIL.n209 9.3005
R349 VTAIL.n289 VTAIL.n288 9.3005
R350 VTAIL.n287 VTAIL.n286 9.3005
R351 VTAIL.n262 VTAIL.n261 9.3005
R352 VTAIL.n227 VTAIL.n226 9.3005
R353 VTAIL.n256 VTAIL.n255 9.3005
R354 VTAIL.n254 VTAIL.n253 9.3005
R355 VTAIL.n231 VTAIL.n230 9.3005
R356 VTAIL.n248 VTAIL.n247 9.3005
R357 VTAIL.n246 VTAIL.n245 9.3005
R358 VTAIL.n235 VTAIL.n234 9.3005
R359 VTAIL.n240 VTAIL.n239 9.3005
R360 VTAIL.n162 VTAIL.n161 9.3005
R361 VTAIL.n121 VTAIL.n120 9.3005
R362 VTAIL.n168 VTAIL.n167 9.3005
R363 VTAIL.n170 VTAIL.n169 9.3005
R364 VTAIL.n117 VTAIL.n116 9.3005
R365 VTAIL.n176 VTAIL.n175 9.3005
R366 VTAIL.n178 VTAIL.n177 9.3005
R367 VTAIL.n114 VTAIL.n111 9.3005
R368 VTAIL.n201 VTAIL.n200 9.3005
R369 VTAIL.n104 VTAIL.n103 9.3005
R370 VTAIL.n195 VTAIL.n194 9.3005
R371 VTAIL.n193 VTAIL.n192 9.3005
R372 VTAIL.n108 VTAIL.n107 9.3005
R373 VTAIL.n187 VTAIL.n186 9.3005
R374 VTAIL.n185 VTAIL.n184 9.3005
R375 VTAIL.n160 VTAIL.n159 9.3005
R376 VTAIL.n125 VTAIL.n124 9.3005
R377 VTAIL.n154 VTAIL.n153 9.3005
R378 VTAIL.n152 VTAIL.n151 9.3005
R379 VTAIL.n129 VTAIL.n128 9.3005
R380 VTAIL.n146 VTAIL.n145 9.3005
R381 VTAIL.n144 VTAIL.n143 9.3005
R382 VTAIL.n133 VTAIL.n132 9.3005
R383 VTAIL.n138 VTAIL.n137 9.3005
R384 VTAIL.n354 VTAIL.n330 8.92171
R385 VTAIL.n370 VTAIL.n369 8.92171
R386 VTAIL.n403 VTAIL.n308 8.92171
R387 VTAIL.n48 VTAIL.n24 8.92171
R388 VTAIL.n64 VTAIL.n63 8.92171
R389 VTAIL.n97 VTAIL.n2 8.92171
R390 VTAIL.n301 VTAIL.n206 8.92171
R391 VTAIL.n269 VTAIL.n268 8.92171
R392 VTAIL.n253 VTAIL.n229 8.92171
R393 VTAIL.n199 VTAIL.n104 8.92171
R394 VTAIL.n167 VTAIL.n166 8.92171
R395 VTAIL.n151 VTAIL.n127 8.92171
R396 VTAIL.n358 VTAIL.n357 8.14595
R397 VTAIL.n366 VTAIL.n324 8.14595
R398 VTAIL.n404 VTAIL.n306 8.14595
R399 VTAIL.n52 VTAIL.n51 8.14595
R400 VTAIL.n60 VTAIL.n18 8.14595
R401 VTAIL.n98 VTAIL.n0 8.14595
R402 VTAIL.n302 VTAIL.n204 8.14595
R403 VTAIL.n265 VTAIL.n223 8.14595
R404 VTAIL.n257 VTAIL.n256 8.14595
R405 VTAIL.n200 VTAIL.n102 8.14595
R406 VTAIL.n163 VTAIL.n121 8.14595
R407 VTAIL.n155 VTAIL.n154 8.14595
R408 VTAIL.n361 VTAIL.n328 7.3702
R409 VTAIL.n365 VTAIL.n326 7.3702
R410 VTAIL.n55 VTAIL.n22 7.3702
R411 VTAIL.n59 VTAIL.n20 7.3702
R412 VTAIL.n264 VTAIL.n225 7.3702
R413 VTAIL.n260 VTAIL.n227 7.3702
R414 VTAIL.n162 VTAIL.n123 7.3702
R415 VTAIL.n158 VTAIL.n125 7.3702
R416 VTAIL.n362 VTAIL.n361 6.59444
R417 VTAIL.n362 VTAIL.n326 6.59444
R418 VTAIL.n56 VTAIL.n55 6.59444
R419 VTAIL.n56 VTAIL.n20 6.59444
R420 VTAIL.n261 VTAIL.n225 6.59444
R421 VTAIL.n261 VTAIL.n260 6.59444
R422 VTAIL.n159 VTAIL.n123 6.59444
R423 VTAIL.n159 VTAIL.n158 6.59444
R424 VTAIL.n358 VTAIL.n328 5.81868
R425 VTAIL.n366 VTAIL.n365 5.81868
R426 VTAIL.n406 VTAIL.n306 5.81868
R427 VTAIL.n52 VTAIL.n22 5.81868
R428 VTAIL.n60 VTAIL.n59 5.81868
R429 VTAIL.n100 VTAIL.n0 5.81868
R430 VTAIL.n304 VTAIL.n204 5.81868
R431 VTAIL.n265 VTAIL.n264 5.81868
R432 VTAIL.n257 VTAIL.n227 5.81868
R433 VTAIL.n202 VTAIL.n102 5.81868
R434 VTAIL.n163 VTAIL.n162 5.81868
R435 VTAIL.n155 VTAIL.n125 5.81868
R436 VTAIL.n357 VTAIL.n330 5.04292
R437 VTAIL.n369 VTAIL.n324 5.04292
R438 VTAIL.n404 VTAIL.n403 5.04292
R439 VTAIL.n51 VTAIL.n24 5.04292
R440 VTAIL.n63 VTAIL.n18 5.04292
R441 VTAIL.n98 VTAIL.n97 5.04292
R442 VTAIL.n302 VTAIL.n301 5.04292
R443 VTAIL.n268 VTAIL.n223 5.04292
R444 VTAIL.n256 VTAIL.n229 5.04292
R445 VTAIL.n200 VTAIL.n199 5.04292
R446 VTAIL.n166 VTAIL.n121 5.04292
R447 VTAIL.n154 VTAIL.n127 5.04292
R448 VTAIL.n340 VTAIL.n339 4.38563
R449 VTAIL.n34 VTAIL.n33 4.38563
R450 VTAIL.n239 VTAIL.n238 4.38563
R451 VTAIL.n137 VTAIL.n136 4.38563
R452 VTAIL.n354 VTAIL.n353 4.26717
R453 VTAIL.n370 VTAIL.n322 4.26717
R454 VTAIL.n400 VTAIL.n308 4.26717
R455 VTAIL.n48 VTAIL.n47 4.26717
R456 VTAIL.n64 VTAIL.n16 4.26717
R457 VTAIL.n94 VTAIL.n2 4.26717
R458 VTAIL.n298 VTAIL.n206 4.26717
R459 VTAIL.n269 VTAIL.n221 4.26717
R460 VTAIL.n253 VTAIL.n252 4.26717
R461 VTAIL.n196 VTAIL.n104 4.26717
R462 VTAIL.n167 VTAIL.n119 4.26717
R463 VTAIL.n151 VTAIL.n150 4.26717
R464 VTAIL.n350 VTAIL.n332 3.49141
R465 VTAIL.n374 VTAIL.n373 3.49141
R466 VTAIL.n399 VTAIL.n310 3.49141
R467 VTAIL.n44 VTAIL.n26 3.49141
R468 VTAIL.n68 VTAIL.n67 3.49141
R469 VTAIL.n93 VTAIL.n4 3.49141
R470 VTAIL.n297 VTAIL.n208 3.49141
R471 VTAIL.n273 VTAIL.n272 3.49141
R472 VTAIL.n249 VTAIL.n231 3.49141
R473 VTAIL.n195 VTAIL.n106 3.49141
R474 VTAIL.n171 VTAIL.n170 3.49141
R475 VTAIL.n147 VTAIL.n129 3.49141
R476 VTAIL.n349 VTAIL.n334 2.71565
R477 VTAIL.n377 VTAIL.n320 2.71565
R478 VTAIL.n396 VTAIL.n395 2.71565
R479 VTAIL.n43 VTAIL.n28 2.71565
R480 VTAIL.n71 VTAIL.n14 2.71565
R481 VTAIL.n90 VTAIL.n89 2.71565
R482 VTAIL.n294 VTAIL.n293 2.71565
R483 VTAIL.n276 VTAIL.n219 2.71565
R484 VTAIL.n248 VTAIL.n233 2.71565
R485 VTAIL.n192 VTAIL.n191 2.71565
R486 VTAIL.n174 VTAIL.n117 2.71565
R487 VTAIL.n146 VTAIL.n131 2.71565
R488 VTAIL.n305 VTAIL.n203 2.28929
R489 VTAIL.n346 VTAIL.n345 1.93989
R490 VTAIL.n378 VTAIL.n318 1.93989
R491 VTAIL.n392 VTAIL.n312 1.93989
R492 VTAIL.n40 VTAIL.n39 1.93989
R493 VTAIL.n72 VTAIL.n12 1.93989
R494 VTAIL.n86 VTAIL.n6 1.93989
R495 VTAIL.n290 VTAIL.n210 1.93989
R496 VTAIL.n277 VTAIL.n217 1.93989
R497 VTAIL.n245 VTAIL.n244 1.93989
R498 VTAIL.n188 VTAIL.n108 1.93989
R499 VTAIL.n175 VTAIL.n115 1.93989
R500 VTAIL.n143 VTAIL.n142 1.93989
R501 VTAIL VTAIL.n101 1.438
R502 VTAIL.n342 VTAIL.n336 1.16414
R503 VTAIL.n383 VTAIL.n381 1.16414
R504 VTAIL.n391 VTAIL.n314 1.16414
R505 VTAIL.n36 VTAIL.n30 1.16414
R506 VTAIL.n77 VTAIL.n75 1.16414
R507 VTAIL.n85 VTAIL.n8 1.16414
R508 VTAIL.n289 VTAIL.n212 1.16414
R509 VTAIL.n281 VTAIL.n280 1.16414
R510 VTAIL.n241 VTAIL.n235 1.16414
R511 VTAIL.n187 VTAIL.n110 1.16414
R512 VTAIL.n179 VTAIL.n178 1.16414
R513 VTAIL.n139 VTAIL.n133 1.16414
R514 VTAIL VTAIL.n407 0.851793
R515 VTAIL.n341 VTAIL.n338 0.388379
R516 VTAIL.n382 VTAIL.n316 0.388379
R517 VTAIL.n388 VTAIL.n387 0.388379
R518 VTAIL.n35 VTAIL.n32 0.388379
R519 VTAIL.n76 VTAIL.n10 0.388379
R520 VTAIL.n82 VTAIL.n81 0.388379
R521 VTAIL.n286 VTAIL.n285 0.388379
R522 VTAIL.n216 VTAIL.n214 0.388379
R523 VTAIL.n240 VTAIL.n237 0.388379
R524 VTAIL.n184 VTAIL.n183 0.388379
R525 VTAIL.n114 VTAIL.n112 0.388379
R526 VTAIL.n138 VTAIL.n135 0.388379
R527 VTAIL.n340 VTAIL.n335 0.155672
R528 VTAIL.n347 VTAIL.n335 0.155672
R529 VTAIL.n348 VTAIL.n347 0.155672
R530 VTAIL.n348 VTAIL.n331 0.155672
R531 VTAIL.n355 VTAIL.n331 0.155672
R532 VTAIL.n356 VTAIL.n355 0.155672
R533 VTAIL.n356 VTAIL.n327 0.155672
R534 VTAIL.n363 VTAIL.n327 0.155672
R535 VTAIL.n364 VTAIL.n363 0.155672
R536 VTAIL.n364 VTAIL.n323 0.155672
R537 VTAIL.n371 VTAIL.n323 0.155672
R538 VTAIL.n372 VTAIL.n371 0.155672
R539 VTAIL.n372 VTAIL.n319 0.155672
R540 VTAIL.n379 VTAIL.n319 0.155672
R541 VTAIL.n380 VTAIL.n379 0.155672
R542 VTAIL.n380 VTAIL.n315 0.155672
R543 VTAIL.n389 VTAIL.n315 0.155672
R544 VTAIL.n390 VTAIL.n389 0.155672
R545 VTAIL.n390 VTAIL.n311 0.155672
R546 VTAIL.n397 VTAIL.n311 0.155672
R547 VTAIL.n398 VTAIL.n397 0.155672
R548 VTAIL.n398 VTAIL.n307 0.155672
R549 VTAIL.n405 VTAIL.n307 0.155672
R550 VTAIL.n34 VTAIL.n29 0.155672
R551 VTAIL.n41 VTAIL.n29 0.155672
R552 VTAIL.n42 VTAIL.n41 0.155672
R553 VTAIL.n42 VTAIL.n25 0.155672
R554 VTAIL.n49 VTAIL.n25 0.155672
R555 VTAIL.n50 VTAIL.n49 0.155672
R556 VTAIL.n50 VTAIL.n21 0.155672
R557 VTAIL.n57 VTAIL.n21 0.155672
R558 VTAIL.n58 VTAIL.n57 0.155672
R559 VTAIL.n58 VTAIL.n17 0.155672
R560 VTAIL.n65 VTAIL.n17 0.155672
R561 VTAIL.n66 VTAIL.n65 0.155672
R562 VTAIL.n66 VTAIL.n13 0.155672
R563 VTAIL.n73 VTAIL.n13 0.155672
R564 VTAIL.n74 VTAIL.n73 0.155672
R565 VTAIL.n74 VTAIL.n9 0.155672
R566 VTAIL.n83 VTAIL.n9 0.155672
R567 VTAIL.n84 VTAIL.n83 0.155672
R568 VTAIL.n84 VTAIL.n5 0.155672
R569 VTAIL.n91 VTAIL.n5 0.155672
R570 VTAIL.n92 VTAIL.n91 0.155672
R571 VTAIL.n92 VTAIL.n1 0.155672
R572 VTAIL.n99 VTAIL.n1 0.155672
R573 VTAIL.n303 VTAIL.n205 0.155672
R574 VTAIL.n296 VTAIL.n205 0.155672
R575 VTAIL.n296 VTAIL.n295 0.155672
R576 VTAIL.n295 VTAIL.n209 0.155672
R577 VTAIL.n288 VTAIL.n209 0.155672
R578 VTAIL.n288 VTAIL.n287 0.155672
R579 VTAIL.n287 VTAIL.n213 0.155672
R580 VTAIL.n279 VTAIL.n213 0.155672
R581 VTAIL.n279 VTAIL.n278 0.155672
R582 VTAIL.n278 VTAIL.n218 0.155672
R583 VTAIL.n271 VTAIL.n218 0.155672
R584 VTAIL.n271 VTAIL.n270 0.155672
R585 VTAIL.n270 VTAIL.n222 0.155672
R586 VTAIL.n263 VTAIL.n222 0.155672
R587 VTAIL.n263 VTAIL.n262 0.155672
R588 VTAIL.n262 VTAIL.n226 0.155672
R589 VTAIL.n255 VTAIL.n226 0.155672
R590 VTAIL.n255 VTAIL.n254 0.155672
R591 VTAIL.n254 VTAIL.n230 0.155672
R592 VTAIL.n247 VTAIL.n230 0.155672
R593 VTAIL.n247 VTAIL.n246 0.155672
R594 VTAIL.n246 VTAIL.n234 0.155672
R595 VTAIL.n239 VTAIL.n234 0.155672
R596 VTAIL.n201 VTAIL.n103 0.155672
R597 VTAIL.n194 VTAIL.n103 0.155672
R598 VTAIL.n194 VTAIL.n193 0.155672
R599 VTAIL.n193 VTAIL.n107 0.155672
R600 VTAIL.n186 VTAIL.n107 0.155672
R601 VTAIL.n186 VTAIL.n185 0.155672
R602 VTAIL.n185 VTAIL.n111 0.155672
R603 VTAIL.n177 VTAIL.n111 0.155672
R604 VTAIL.n177 VTAIL.n176 0.155672
R605 VTAIL.n176 VTAIL.n116 0.155672
R606 VTAIL.n169 VTAIL.n116 0.155672
R607 VTAIL.n169 VTAIL.n168 0.155672
R608 VTAIL.n168 VTAIL.n120 0.155672
R609 VTAIL.n161 VTAIL.n120 0.155672
R610 VTAIL.n161 VTAIL.n160 0.155672
R611 VTAIL.n160 VTAIL.n124 0.155672
R612 VTAIL.n153 VTAIL.n124 0.155672
R613 VTAIL.n153 VTAIL.n152 0.155672
R614 VTAIL.n152 VTAIL.n128 0.155672
R615 VTAIL.n145 VTAIL.n128 0.155672
R616 VTAIL.n145 VTAIL.n144 0.155672
R617 VTAIL.n144 VTAIL.n132 0.155672
R618 VTAIL.n137 VTAIL.n132 0.155672
R619 VDD2.n197 VDD2.n101 289.615
R620 VDD2.n96 VDD2.n0 289.615
R621 VDD2.n198 VDD2.n197 185
R622 VDD2.n196 VDD2.n195 185
R623 VDD2.n105 VDD2.n104 185
R624 VDD2.n190 VDD2.n189 185
R625 VDD2.n188 VDD2.n187 185
R626 VDD2.n109 VDD2.n108 185
R627 VDD2.n182 VDD2.n181 185
R628 VDD2.n180 VDD2.n111 185
R629 VDD2.n179 VDD2.n178 185
R630 VDD2.n114 VDD2.n112 185
R631 VDD2.n173 VDD2.n172 185
R632 VDD2.n171 VDD2.n170 185
R633 VDD2.n118 VDD2.n117 185
R634 VDD2.n165 VDD2.n164 185
R635 VDD2.n163 VDD2.n162 185
R636 VDD2.n122 VDD2.n121 185
R637 VDD2.n157 VDD2.n156 185
R638 VDD2.n155 VDD2.n154 185
R639 VDD2.n126 VDD2.n125 185
R640 VDD2.n149 VDD2.n148 185
R641 VDD2.n147 VDD2.n146 185
R642 VDD2.n130 VDD2.n129 185
R643 VDD2.n141 VDD2.n140 185
R644 VDD2.n139 VDD2.n138 185
R645 VDD2.n134 VDD2.n133 185
R646 VDD2.n32 VDD2.n31 185
R647 VDD2.n37 VDD2.n36 185
R648 VDD2.n39 VDD2.n38 185
R649 VDD2.n28 VDD2.n27 185
R650 VDD2.n45 VDD2.n44 185
R651 VDD2.n47 VDD2.n46 185
R652 VDD2.n24 VDD2.n23 185
R653 VDD2.n53 VDD2.n52 185
R654 VDD2.n55 VDD2.n54 185
R655 VDD2.n20 VDD2.n19 185
R656 VDD2.n61 VDD2.n60 185
R657 VDD2.n63 VDD2.n62 185
R658 VDD2.n16 VDD2.n15 185
R659 VDD2.n69 VDD2.n68 185
R660 VDD2.n71 VDD2.n70 185
R661 VDD2.n12 VDD2.n11 185
R662 VDD2.n78 VDD2.n77 185
R663 VDD2.n79 VDD2.n10 185
R664 VDD2.n81 VDD2.n80 185
R665 VDD2.n8 VDD2.n7 185
R666 VDD2.n87 VDD2.n86 185
R667 VDD2.n89 VDD2.n88 185
R668 VDD2.n4 VDD2.n3 185
R669 VDD2.n95 VDD2.n94 185
R670 VDD2.n97 VDD2.n96 185
R671 VDD2.n135 VDD2.t0 147.659
R672 VDD2.n33 VDD2.t1 147.659
R673 VDD2.n197 VDD2.n196 104.615
R674 VDD2.n196 VDD2.n104 104.615
R675 VDD2.n189 VDD2.n104 104.615
R676 VDD2.n189 VDD2.n188 104.615
R677 VDD2.n188 VDD2.n108 104.615
R678 VDD2.n181 VDD2.n108 104.615
R679 VDD2.n181 VDD2.n180 104.615
R680 VDD2.n180 VDD2.n179 104.615
R681 VDD2.n179 VDD2.n112 104.615
R682 VDD2.n172 VDD2.n112 104.615
R683 VDD2.n172 VDD2.n171 104.615
R684 VDD2.n171 VDD2.n117 104.615
R685 VDD2.n164 VDD2.n117 104.615
R686 VDD2.n164 VDD2.n163 104.615
R687 VDD2.n163 VDD2.n121 104.615
R688 VDD2.n156 VDD2.n121 104.615
R689 VDD2.n156 VDD2.n155 104.615
R690 VDD2.n155 VDD2.n125 104.615
R691 VDD2.n148 VDD2.n125 104.615
R692 VDD2.n148 VDD2.n147 104.615
R693 VDD2.n147 VDD2.n129 104.615
R694 VDD2.n140 VDD2.n129 104.615
R695 VDD2.n140 VDD2.n139 104.615
R696 VDD2.n139 VDD2.n133 104.615
R697 VDD2.n37 VDD2.n31 104.615
R698 VDD2.n38 VDD2.n37 104.615
R699 VDD2.n38 VDD2.n27 104.615
R700 VDD2.n45 VDD2.n27 104.615
R701 VDD2.n46 VDD2.n45 104.615
R702 VDD2.n46 VDD2.n23 104.615
R703 VDD2.n53 VDD2.n23 104.615
R704 VDD2.n54 VDD2.n53 104.615
R705 VDD2.n54 VDD2.n19 104.615
R706 VDD2.n61 VDD2.n19 104.615
R707 VDD2.n62 VDD2.n61 104.615
R708 VDD2.n62 VDD2.n15 104.615
R709 VDD2.n69 VDD2.n15 104.615
R710 VDD2.n70 VDD2.n69 104.615
R711 VDD2.n70 VDD2.n11 104.615
R712 VDD2.n78 VDD2.n11 104.615
R713 VDD2.n79 VDD2.n78 104.615
R714 VDD2.n80 VDD2.n79 104.615
R715 VDD2.n80 VDD2.n7 104.615
R716 VDD2.n87 VDD2.n7 104.615
R717 VDD2.n88 VDD2.n87 104.615
R718 VDD2.n88 VDD2.n3 104.615
R719 VDD2.n95 VDD2.n3 104.615
R720 VDD2.n96 VDD2.n95 104.615
R721 VDD2.n202 VDD2.n100 95.321
R722 VDD2.t0 VDD2.n133 52.3082
R723 VDD2.t1 VDD2.n31 52.3082
R724 VDD2.n202 VDD2.n201 48.6702
R725 VDD2.n135 VDD2.n134 15.6677
R726 VDD2.n33 VDD2.n32 15.6677
R727 VDD2.n182 VDD2.n111 13.1884
R728 VDD2.n81 VDD2.n10 13.1884
R729 VDD2.n183 VDD2.n109 12.8005
R730 VDD2.n178 VDD2.n113 12.8005
R731 VDD2.n138 VDD2.n137 12.8005
R732 VDD2.n36 VDD2.n35 12.8005
R733 VDD2.n77 VDD2.n76 12.8005
R734 VDD2.n82 VDD2.n8 12.8005
R735 VDD2.n187 VDD2.n186 12.0247
R736 VDD2.n177 VDD2.n114 12.0247
R737 VDD2.n141 VDD2.n132 12.0247
R738 VDD2.n39 VDD2.n30 12.0247
R739 VDD2.n75 VDD2.n12 12.0247
R740 VDD2.n86 VDD2.n85 12.0247
R741 VDD2.n190 VDD2.n107 11.249
R742 VDD2.n174 VDD2.n173 11.249
R743 VDD2.n142 VDD2.n130 11.249
R744 VDD2.n40 VDD2.n28 11.249
R745 VDD2.n72 VDD2.n71 11.249
R746 VDD2.n89 VDD2.n6 11.249
R747 VDD2.n191 VDD2.n105 10.4732
R748 VDD2.n170 VDD2.n116 10.4732
R749 VDD2.n146 VDD2.n145 10.4732
R750 VDD2.n44 VDD2.n43 10.4732
R751 VDD2.n68 VDD2.n14 10.4732
R752 VDD2.n90 VDD2.n4 10.4732
R753 VDD2.n195 VDD2.n194 9.69747
R754 VDD2.n169 VDD2.n118 9.69747
R755 VDD2.n149 VDD2.n128 9.69747
R756 VDD2.n47 VDD2.n26 9.69747
R757 VDD2.n67 VDD2.n16 9.69747
R758 VDD2.n94 VDD2.n93 9.69747
R759 VDD2.n201 VDD2.n200 9.45567
R760 VDD2.n100 VDD2.n99 9.45567
R761 VDD2.n161 VDD2.n160 9.3005
R762 VDD2.n120 VDD2.n119 9.3005
R763 VDD2.n167 VDD2.n166 9.3005
R764 VDD2.n169 VDD2.n168 9.3005
R765 VDD2.n116 VDD2.n115 9.3005
R766 VDD2.n175 VDD2.n174 9.3005
R767 VDD2.n177 VDD2.n176 9.3005
R768 VDD2.n113 VDD2.n110 9.3005
R769 VDD2.n200 VDD2.n199 9.3005
R770 VDD2.n103 VDD2.n102 9.3005
R771 VDD2.n194 VDD2.n193 9.3005
R772 VDD2.n192 VDD2.n191 9.3005
R773 VDD2.n107 VDD2.n106 9.3005
R774 VDD2.n186 VDD2.n185 9.3005
R775 VDD2.n184 VDD2.n183 9.3005
R776 VDD2.n159 VDD2.n158 9.3005
R777 VDD2.n124 VDD2.n123 9.3005
R778 VDD2.n153 VDD2.n152 9.3005
R779 VDD2.n151 VDD2.n150 9.3005
R780 VDD2.n128 VDD2.n127 9.3005
R781 VDD2.n145 VDD2.n144 9.3005
R782 VDD2.n143 VDD2.n142 9.3005
R783 VDD2.n132 VDD2.n131 9.3005
R784 VDD2.n137 VDD2.n136 9.3005
R785 VDD2.n99 VDD2.n98 9.3005
R786 VDD2.n2 VDD2.n1 9.3005
R787 VDD2.n93 VDD2.n92 9.3005
R788 VDD2.n91 VDD2.n90 9.3005
R789 VDD2.n6 VDD2.n5 9.3005
R790 VDD2.n85 VDD2.n84 9.3005
R791 VDD2.n83 VDD2.n82 9.3005
R792 VDD2.n22 VDD2.n21 9.3005
R793 VDD2.n51 VDD2.n50 9.3005
R794 VDD2.n49 VDD2.n48 9.3005
R795 VDD2.n26 VDD2.n25 9.3005
R796 VDD2.n43 VDD2.n42 9.3005
R797 VDD2.n41 VDD2.n40 9.3005
R798 VDD2.n30 VDD2.n29 9.3005
R799 VDD2.n35 VDD2.n34 9.3005
R800 VDD2.n57 VDD2.n56 9.3005
R801 VDD2.n59 VDD2.n58 9.3005
R802 VDD2.n18 VDD2.n17 9.3005
R803 VDD2.n65 VDD2.n64 9.3005
R804 VDD2.n67 VDD2.n66 9.3005
R805 VDD2.n14 VDD2.n13 9.3005
R806 VDD2.n73 VDD2.n72 9.3005
R807 VDD2.n75 VDD2.n74 9.3005
R808 VDD2.n76 VDD2.n9 9.3005
R809 VDD2.n198 VDD2.n103 8.92171
R810 VDD2.n166 VDD2.n165 8.92171
R811 VDD2.n150 VDD2.n126 8.92171
R812 VDD2.n48 VDD2.n24 8.92171
R813 VDD2.n64 VDD2.n63 8.92171
R814 VDD2.n97 VDD2.n2 8.92171
R815 VDD2.n199 VDD2.n101 8.14595
R816 VDD2.n162 VDD2.n120 8.14595
R817 VDD2.n154 VDD2.n153 8.14595
R818 VDD2.n52 VDD2.n51 8.14595
R819 VDD2.n60 VDD2.n18 8.14595
R820 VDD2.n98 VDD2.n0 8.14595
R821 VDD2.n161 VDD2.n122 7.3702
R822 VDD2.n157 VDD2.n124 7.3702
R823 VDD2.n55 VDD2.n22 7.3702
R824 VDD2.n59 VDD2.n20 7.3702
R825 VDD2.n158 VDD2.n122 6.59444
R826 VDD2.n158 VDD2.n157 6.59444
R827 VDD2.n56 VDD2.n55 6.59444
R828 VDD2.n56 VDD2.n20 6.59444
R829 VDD2.n201 VDD2.n101 5.81868
R830 VDD2.n162 VDD2.n161 5.81868
R831 VDD2.n154 VDD2.n124 5.81868
R832 VDD2.n52 VDD2.n22 5.81868
R833 VDD2.n60 VDD2.n59 5.81868
R834 VDD2.n100 VDD2.n0 5.81868
R835 VDD2.n199 VDD2.n198 5.04292
R836 VDD2.n165 VDD2.n120 5.04292
R837 VDD2.n153 VDD2.n126 5.04292
R838 VDD2.n51 VDD2.n24 5.04292
R839 VDD2.n63 VDD2.n18 5.04292
R840 VDD2.n98 VDD2.n97 5.04292
R841 VDD2.n136 VDD2.n135 4.38563
R842 VDD2.n34 VDD2.n33 4.38563
R843 VDD2.n195 VDD2.n103 4.26717
R844 VDD2.n166 VDD2.n118 4.26717
R845 VDD2.n150 VDD2.n149 4.26717
R846 VDD2.n48 VDD2.n47 4.26717
R847 VDD2.n64 VDD2.n16 4.26717
R848 VDD2.n94 VDD2.n2 4.26717
R849 VDD2.n194 VDD2.n105 3.49141
R850 VDD2.n170 VDD2.n169 3.49141
R851 VDD2.n146 VDD2.n128 3.49141
R852 VDD2.n44 VDD2.n26 3.49141
R853 VDD2.n68 VDD2.n67 3.49141
R854 VDD2.n93 VDD2.n4 3.49141
R855 VDD2.n191 VDD2.n190 2.71565
R856 VDD2.n173 VDD2.n116 2.71565
R857 VDD2.n145 VDD2.n130 2.71565
R858 VDD2.n43 VDD2.n28 2.71565
R859 VDD2.n71 VDD2.n14 2.71565
R860 VDD2.n90 VDD2.n89 2.71565
R861 VDD2.n187 VDD2.n107 1.93989
R862 VDD2.n174 VDD2.n114 1.93989
R863 VDD2.n142 VDD2.n141 1.93989
R864 VDD2.n40 VDD2.n39 1.93989
R865 VDD2.n72 VDD2.n12 1.93989
R866 VDD2.n86 VDD2.n6 1.93989
R867 VDD2.n186 VDD2.n109 1.16414
R868 VDD2.n178 VDD2.n177 1.16414
R869 VDD2.n138 VDD2.n132 1.16414
R870 VDD2.n36 VDD2.n30 1.16414
R871 VDD2.n77 VDD2.n75 1.16414
R872 VDD2.n85 VDD2.n8 1.16414
R873 VDD2 VDD2.n202 0.968172
R874 VDD2.n183 VDD2.n182 0.388379
R875 VDD2.n113 VDD2.n111 0.388379
R876 VDD2.n137 VDD2.n134 0.388379
R877 VDD2.n35 VDD2.n32 0.388379
R878 VDD2.n76 VDD2.n10 0.388379
R879 VDD2.n82 VDD2.n81 0.388379
R880 VDD2.n200 VDD2.n102 0.155672
R881 VDD2.n193 VDD2.n102 0.155672
R882 VDD2.n193 VDD2.n192 0.155672
R883 VDD2.n192 VDD2.n106 0.155672
R884 VDD2.n185 VDD2.n106 0.155672
R885 VDD2.n185 VDD2.n184 0.155672
R886 VDD2.n184 VDD2.n110 0.155672
R887 VDD2.n176 VDD2.n110 0.155672
R888 VDD2.n176 VDD2.n175 0.155672
R889 VDD2.n175 VDD2.n115 0.155672
R890 VDD2.n168 VDD2.n115 0.155672
R891 VDD2.n168 VDD2.n167 0.155672
R892 VDD2.n167 VDD2.n119 0.155672
R893 VDD2.n160 VDD2.n119 0.155672
R894 VDD2.n160 VDD2.n159 0.155672
R895 VDD2.n159 VDD2.n123 0.155672
R896 VDD2.n152 VDD2.n123 0.155672
R897 VDD2.n152 VDD2.n151 0.155672
R898 VDD2.n151 VDD2.n127 0.155672
R899 VDD2.n144 VDD2.n127 0.155672
R900 VDD2.n144 VDD2.n143 0.155672
R901 VDD2.n143 VDD2.n131 0.155672
R902 VDD2.n136 VDD2.n131 0.155672
R903 VDD2.n34 VDD2.n29 0.155672
R904 VDD2.n41 VDD2.n29 0.155672
R905 VDD2.n42 VDD2.n41 0.155672
R906 VDD2.n42 VDD2.n25 0.155672
R907 VDD2.n49 VDD2.n25 0.155672
R908 VDD2.n50 VDD2.n49 0.155672
R909 VDD2.n50 VDD2.n21 0.155672
R910 VDD2.n57 VDD2.n21 0.155672
R911 VDD2.n58 VDD2.n57 0.155672
R912 VDD2.n58 VDD2.n17 0.155672
R913 VDD2.n65 VDD2.n17 0.155672
R914 VDD2.n66 VDD2.n65 0.155672
R915 VDD2.n66 VDD2.n13 0.155672
R916 VDD2.n73 VDD2.n13 0.155672
R917 VDD2.n74 VDD2.n73 0.155672
R918 VDD2.n74 VDD2.n9 0.155672
R919 VDD2.n83 VDD2.n9 0.155672
R920 VDD2.n84 VDD2.n83 0.155672
R921 VDD2.n84 VDD2.n5 0.155672
R922 VDD2.n91 VDD2.n5 0.155672
R923 VDD2.n92 VDD2.n91 0.155672
R924 VDD2.n92 VDD2.n1 0.155672
R925 VDD2.n99 VDD2.n1 0.155672
R926 B.n923 B.n922 585
R927 B.n924 B.n923 585
R928 B.n388 B.n127 585
R929 B.n387 B.n386 585
R930 B.n385 B.n384 585
R931 B.n383 B.n382 585
R932 B.n381 B.n380 585
R933 B.n379 B.n378 585
R934 B.n377 B.n376 585
R935 B.n375 B.n374 585
R936 B.n373 B.n372 585
R937 B.n371 B.n370 585
R938 B.n369 B.n368 585
R939 B.n367 B.n366 585
R940 B.n365 B.n364 585
R941 B.n363 B.n362 585
R942 B.n361 B.n360 585
R943 B.n359 B.n358 585
R944 B.n357 B.n356 585
R945 B.n355 B.n354 585
R946 B.n353 B.n352 585
R947 B.n351 B.n350 585
R948 B.n349 B.n348 585
R949 B.n347 B.n346 585
R950 B.n345 B.n344 585
R951 B.n343 B.n342 585
R952 B.n341 B.n340 585
R953 B.n339 B.n338 585
R954 B.n337 B.n336 585
R955 B.n335 B.n334 585
R956 B.n333 B.n332 585
R957 B.n331 B.n330 585
R958 B.n329 B.n328 585
R959 B.n327 B.n326 585
R960 B.n325 B.n324 585
R961 B.n323 B.n322 585
R962 B.n321 B.n320 585
R963 B.n319 B.n318 585
R964 B.n317 B.n316 585
R965 B.n315 B.n314 585
R966 B.n313 B.n312 585
R967 B.n311 B.n310 585
R968 B.n309 B.n308 585
R969 B.n307 B.n306 585
R970 B.n305 B.n304 585
R971 B.n303 B.n302 585
R972 B.n301 B.n300 585
R973 B.n299 B.n298 585
R974 B.n297 B.n296 585
R975 B.n295 B.n294 585
R976 B.n293 B.n292 585
R977 B.n291 B.n290 585
R978 B.n289 B.n288 585
R979 B.n287 B.n286 585
R980 B.n285 B.n284 585
R981 B.n283 B.n282 585
R982 B.n281 B.n280 585
R983 B.n279 B.n278 585
R984 B.n277 B.n276 585
R985 B.n275 B.n274 585
R986 B.n273 B.n272 585
R987 B.n270 B.n269 585
R988 B.n268 B.n267 585
R989 B.n266 B.n265 585
R990 B.n264 B.n263 585
R991 B.n262 B.n261 585
R992 B.n260 B.n259 585
R993 B.n258 B.n257 585
R994 B.n256 B.n255 585
R995 B.n254 B.n253 585
R996 B.n252 B.n251 585
R997 B.n250 B.n249 585
R998 B.n248 B.n247 585
R999 B.n246 B.n245 585
R1000 B.n244 B.n243 585
R1001 B.n242 B.n241 585
R1002 B.n240 B.n239 585
R1003 B.n238 B.n237 585
R1004 B.n236 B.n235 585
R1005 B.n234 B.n233 585
R1006 B.n232 B.n231 585
R1007 B.n230 B.n229 585
R1008 B.n228 B.n227 585
R1009 B.n226 B.n225 585
R1010 B.n224 B.n223 585
R1011 B.n222 B.n221 585
R1012 B.n220 B.n219 585
R1013 B.n218 B.n217 585
R1014 B.n216 B.n215 585
R1015 B.n214 B.n213 585
R1016 B.n212 B.n211 585
R1017 B.n210 B.n209 585
R1018 B.n208 B.n207 585
R1019 B.n206 B.n205 585
R1020 B.n204 B.n203 585
R1021 B.n202 B.n201 585
R1022 B.n200 B.n199 585
R1023 B.n198 B.n197 585
R1024 B.n196 B.n195 585
R1025 B.n194 B.n193 585
R1026 B.n192 B.n191 585
R1027 B.n190 B.n189 585
R1028 B.n188 B.n187 585
R1029 B.n186 B.n185 585
R1030 B.n184 B.n183 585
R1031 B.n182 B.n181 585
R1032 B.n180 B.n179 585
R1033 B.n178 B.n177 585
R1034 B.n176 B.n175 585
R1035 B.n174 B.n173 585
R1036 B.n172 B.n171 585
R1037 B.n170 B.n169 585
R1038 B.n168 B.n167 585
R1039 B.n166 B.n165 585
R1040 B.n164 B.n163 585
R1041 B.n162 B.n161 585
R1042 B.n160 B.n159 585
R1043 B.n158 B.n157 585
R1044 B.n156 B.n155 585
R1045 B.n154 B.n153 585
R1046 B.n152 B.n151 585
R1047 B.n150 B.n149 585
R1048 B.n148 B.n147 585
R1049 B.n146 B.n145 585
R1050 B.n144 B.n143 585
R1051 B.n142 B.n141 585
R1052 B.n140 B.n139 585
R1053 B.n138 B.n137 585
R1054 B.n136 B.n135 585
R1055 B.n134 B.n133 585
R1056 B.n921 B.n62 585
R1057 B.n925 B.n62 585
R1058 B.n920 B.n61 585
R1059 B.n926 B.n61 585
R1060 B.n919 B.n918 585
R1061 B.n918 B.n57 585
R1062 B.n917 B.n56 585
R1063 B.n932 B.n56 585
R1064 B.n916 B.n55 585
R1065 B.n933 B.n55 585
R1066 B.n915 B.n54 585
R1067 B.n934 B.n54 585
R1068 B.n914 B.n913 585
R1069 B.n913 B.n50 585
R1070 B.n912 B.n49 585
R1071 B.n940 B.n49 585
R1072 B.n911 B.n48 585
R1073 B.n941 B.n48 585
R1074 B.n910 B.n47 585
R1075 B.n942 B.n47 585
R1076 B.n909 B.n908 585
R1077 B.n908 B.n43 585
R1078 B.n907 B.n42 585
R1079 B.n948 B.n42 585
R1080 B.n906 B.n41 585
R1081 B.n949 B.n41 585
R1082 B.n905 B.n40 585
R1083 B.n950 B.n40 585
R1084 B.n904 B.n903 585
R1085 B.n903 B.n36 585
R1086 B.n902 B.n35 585
R1087 B.n956 B.n35 585
R1088 B.n901 B.n34 585
R1089 B.n957 B.n34 585
R1090 B.n900 B.n33 585
R1091 B.n958 B.n33 585
R1092 B.n899 B.n898 585
R1093 B.n898 B.n29 585
R1094 B.n897 B.n28 585
R1095 B.n964 B.n28 585
R1096 B.n896 B.n27 585
R1097 B.n965 B.n27 585
R1098 B.n895 B.n26 585
R1099 B.n966 B.n26 585
R1100 B.n894 B.n893 585
R1101 B.n893 B.n22 585
R1102 B.n892 B.n21 585
R1103 B.n972 B.n21 585
R1104 B.n891 B.n20 585
R1105 B.n973 B.n20 585
R1106 B.n890 B.n19 585
R1107 B.n974 B.n19 585
R1108 B.n889 B.n888 585
R1109 B.n888 B.n15 585
R1110 B.n887 B.n14 585
R1111 B.n980 B.n14 585
R1112 B.n886 B.n13 585
R1113 B.n981 B.n13 585
R1114 B.n885 B.n12 585
R1115 B.n982 B.n12 585
R1116 B.n884 B.n883 585
R1117 B.n883 B.n8 585
R1118 B.n882 B.n7 585
R1119 B.n988 B.n7 585
R1120 B.n881 B.n6 585
R1121 B.n989 B.n6 585
R1122 B.n880 B.n5 585
R1123 B.n990 B.n5 585
R1124 B.n879 B.n878 585
R1125 B.n878 B.n4 585
R1126 B.n877 B.n389 585
R1127 B.n877 B.n876 585
R1128 B.n867 B.n390 585
R1129 B.n391 B.n390 585
R1130 B.n869 B.n868 585
R1131 B.n870 B.n869 585
R1132 B.n866 B.n396 585
R1133 B.n396 B.n395 585
R1134 B.n865 B.n864 585
R1135 B.n864 B.n863 585
R1136 B.n398 B.n397 585
R1137 B.n399 B.n398 585
R1138 B.n856 B.n855 585
R1139 B.n857 B.n856 585
R1140 B.n854 B.n404 585
R1141 B.n404 B.n403 585
R1142 B.n853 B.n852 585
R1143 B.n852 B.n851 585
R1144 B.n406 B.n405 585
R1145 B.n407 B.n406 585
R1146 B.n844 B.n843 585
R1147 B.n845 B.n844 585
R1148 B.n842 B.n412 585
R1149 B.n412 B.n411 585
R1150 B.n841 B.n840 585
R1151 B.n840 B.n839 585
R1152 B.n414 B.n413 585
R1153 B.n415 B.n414 585
R1154 B.n832 B.n831 585
R1155 B.n833 B.n832 585
R1156 B.n830 B.n420 585
R1157 B.n420 B.n419 585
R1158 B.n829 B.n828 585
R1159 B.n828 B.n827 585
R1160 B.n422 B.n421 585
R1161 B.n423 B.n422 585
R1162 B.n820 B.n819 585
R1163 B.n821 B.n820 585
R1164 B.n818 B.n428 585
R1165 B.n428 B.n427 585
R1166 B.n817 B.n816 585
R1167 B.n816 B.n815 585
R1168 B.n430 B.n429 585
R1169 B.n431 B.n430 585
R1170 B.n808 B.n807 585
R1171 B.n809 B.n808 585
R1172 B.n806 B.n436 585
R1173 B.n436 B.n435 585
R1174 B.n805 B.n804 585
R1175 B.n804 B.n803 585
R1176 B.n438 B.n437 585
R1177 B.n439 B.n438 585
R1178 B.n796 B.n795 585
R1179 B.n797 B.n796 585
R1180 B.n794 B.n444 585
R1181 B.n444 B.n443 585
R1182 B.n793 B.n792 585
R1183 B.n792 B.n791 585
R1184 B.n446 B.n445 585
R1185 B.n447 B.n446 585
R1186 B.n784 B.n783 585
R1187 B.n785 B.n784 585
R1188 B.n782 B.n452 585
R1189 B.n452 B.n451 585
R1190 B.n776 B.n775 585
R1191 B.n774 B.n518 585
R1192 B.n773 B.n517 585
R1193 B.n778 B.n517 585
R1194 B.n772 B.n771 585
R1195 B.n770 B.n769 585
R1196 B.n768 B.n767 585
R1197 B.n766 B.n765 585
R1198 B.n764 B.n763 585
R1199 B.n762 B.n761 585
R1200 B.n760 B.n759 585
R1201 B.n758 B.n757 585
R1202 B.n756 B.n755 585
R1203 B.n754 B.n753 585
R1204 B.n752 B.n751 585
R1205 B.n750 B.n749 585
R1206 B.n748 B.n747 585
R1207 B.n746 B.n745 585
R1208 B.n744 B.n743 585
R1209 B.n742 B.n741 585
R1210 B.n740 B.n739 585
R1211 B.n738 B.n737 585
R1212 B.n736 B.n735 585
R1213 B.n734 B.n733 585
R1214 B.n732 B.n731 585
R1215 B.n730 B.n729 585
R1216 B.n728 B.n727 585
R1217 B.n726 B.n725 585
R1218 B.n724 B.n723 585
R1219 B.n722 B.n721 585
R1220 B.n720 B.n719 585
R1221 B.n718 B.n717 585
R1222 B.n716 B.n715 585
R1223 B.n714 B.n713 585
R1224 B.n712 B.n711 585
R1225 B.n710 B.n709 585
R1226 B.n708 B.n707 585
R1227 B.n706 B.n705 585
R1228 B.n704 B.n703 585
R1229 B.n702 B.n701 585
R1230 B.n700 B.n699 585
R1231 B.n698 B.n697 585
R1232 B.n696 B.n695 585
R1233 B.n694 B.n693 585
R1234 B.n692 B.n691 585
R1235 B.n690 B.n689 585
R1236 B.n688 B.n687 585
R1237 B.n686 B.n685 585
R1238 B.n684 B.n683 585
R1239 B.n682 B.n681 585
R1240 B.n680 B.n679 585
R1241 B.n678 B.n677 585
R1242 B.n676 B.n675 585
R1243 B.n674 B.n673 585
R1244 B.n672 B.n671 585
R1245 B.n670 B.n669 585
R1246 B.n668 B.n667 585
R1247 B.n666 B.n665 585
R1248 B.n664 B.n663 585
R1249 B.n662 B.n661 585
R1250 B.n660 B.n659 585
R1251 B.n657 B.n656 585
R1252 B.n655 B.n654 585
R1253 B.n653 B.n652 585
R1254 B.n651 B.n650 585
R1255 B.n649 B.n648 585
R1256 B.n647 B.n646 585
R1257 B.n645 B.n644 585
R1258 B.n643 B.n642 585
R1259 B.n641 B.n640 585
R1260 B.n639 B.n638 585
R1261 B.n637 B.n636 585
R1262 B.n635 B.n634 585
R1263 B.n633 B.n632 585
R1264 B.n631 B.n630 585
R1265 B.n629 B.n628 585
R1266 B.n627 B.n626 585
R1267 B.n625 B.n624 585
R1268 B.n623 B.n622 585
R1269 B.n621 B.n620 585
R1270 B.n619 B.n618 585
R1271 B.n617 B.n616 585
R1272 B.n615 B.n614 585
R1273 B.n613 B.n612 585
R1274 B.n611 B.n610 585
R1275 B.n609 B.n608 585
R1276 B.n607 B.n606 585
R1277 B.n605 B.n604 585
R1278 B.n603 B.n602 585
R1279 B.n601 B.n600 585
R1280 B.n599 B.n598 585
R1281 B.n597 B.n596 585
R1282 B.n595 B.n594 585
R1283 B.n593 B.n592 585
R1284 B.n591 B.n590 585
R1285 B.n589 B.n588 585
R1286 B.n587 B.n586 585
R1287 B.n585 B.n584 585
R1288 B.n583 B.n582 585
R1289 B.n581 B.n580 585
R1290 B.n579 B.n578 585
R1291 B.n577 B.n576 585
R1292 B.n575 B.n574 585
R1293 B.n573 B.n572 585
R1294 B.n571 B.n570 585
R1295 B.n569 B.n568 585
R1296 B.n567 B.n566 585
R1297 B.n565 B.n564 585
R1298 B.n563 B.n562 585
R1299 B.n561 B.n560 585
R1300 B.n559 B.n558 585
R1301 B.n557 B.n556 585
R1302 B.n555 B.n554 585
R1303 B.n553 B.n552 585
R1304 B.n551 B.n550 585
R1305 B.n549 B.n548 585
R1306 B.n547 B.n546 585
R1307 B.n545 B.n544 585
R1308 B.n543 B.n542 585
R1309 B.n541 B.n540 585
R1310 B.n539 B.n538 585
R1311 B.n537 B.n536 585
R1312 B.n535 B.n534 585
R1313 B.n533 B.n532 585
R1314 B.n531 B.n530 585
R1315 B.n529 B.n528 585
R1316 B.n527 B.n526 585
R1317 B.n525 B.n524 585
R1318 B.n454 B.n453 585
R1319 B.n781 B.n780 585
R1320 B.n450 B.n449 585
R1321 B.n451 B.n450 585
R1322 B.n787 B.n786 585
R1323 B.n786 B.n785 585
R1324 B.n788 B.n448 585
R1325 B.n448 B.n447 585
R1326 B.n790 B.n789 585
R1327 B.n791 B.n790 585
R1328 B.n442 B.n441 585
R1329 B.n443 B.n442 585
R1330 B.n799 B.n798 585
R1331 B.n798 B.n797 585
R1332 B.n800 B.n440 585
R1333 B.n440 B.n439 585
R1334 B.n802 B.n801 585
R1335 B.n803 B.n802 585
R1336 B.n434 B.n433 585
R1337 B.n435 B.n434 585
R1338 B.n811 B.n810 585
R1339 B.n810 B.n809 585
R1340 B.n812 B.n432 585
R1341 B.n432 B.n431 585
R1342 B.n814 B.n813 585
R1343 B.n815 B.n814 585
R1344 B.n426 B.n425 585
R1345 B.n427 B.n426 585
R1346 B.n823 B.n822 585
R1347 B.n822 B.n821 585
R1348 B.n824 B.n424 585
R1349 B.n424 B.n423 585
R1350 B.n826 B.n825 585
R1351 B.n827 B.n826 585
R1352 B.n418 B.n417 585
R1353 B.n419 B.n418 585
R1354 B.n835 B.n834 585
R1355 B.n834 B.n833 585
R1356 B.n836 B.n416 585
R1357 B.n416 B.n415 585
R1358 B.n838 B.n837 585
R1359 B.n839 B.n838 585
R1360 B.n410 B.n409 585
R1361 B.n411 B.n410 585
R1362 B.n847 B.n846 585
R1363 B.n846 B.n845 585
R1364 B.n848 B.n408 585
R1365 B.n408 B.n407 585
R1366 B.n850 B.n849 585
R1367 B.n851 B.n850 585
R1368 B.n402 B.n401 585
R1369 B.n403 B.n402 585
R1370 B.n859 B.n858 585
R1371 B.n858 B.n857 585
R1372 B.n860 B.n400 585
R1373 B.n400 B.n399 585
R1374 B.n862 B.n861 585
R1375 B.n863 B.n862 585
R1376 B.n394 B.n393 585
R1377 B.n395 B.n394 585
R1378 B.n872 B.n871 585
R1379 B.n871 B.n870 585
R1380 B.n873 B.n392 585
R1381 B.n392 B.n391 585
R1382 B.n875 B.n874 585
R1383 B.n876 B.n875 585
R1384 B.n2 B.n0 585
R1385 B.n4 B.n2 585
R1386 B.n3 B.n1 585
R1387 B.n989 B.n3 585
R1388 B.n987 B.n986 585
R1389 B.n988 B.n987 585
R1390 B.n985 B.n9 585
R1391 B.n9 B.n8 585
R1392 B.n984 B.n983 585
R1393 B.n983 B.n982 585
R1394 B.n11 B.n10 585
R1395 B.n981 B.n11 585
R1396 B.n979 B.n978 585
R1397 B.n980 B.n979 585
R1398 B.n977 B.n16 585
R1399 B.n16 B.n15 585
R1400 B.n976 B.n975 585
R1401 B.n975 B.n974 585
R1402 B.n18 B.n17 585
R1403 B.n973 B.n18 585
R1404 B.n971 B.n970 585
R1405 B.n972 B.n971 585
R1406 B.n969 B.n23 585
R1407 B.n23 B.n22 585
R1408 B.n968 B.n967 585
R1409 B.n967 B.n966 585
R1410 B.n25 B.n24 585
R1411 B.n965 B.n25 585
R1412 B.n963 B.n962 585
R1413 B.n964 B.n963 585
R1414 B.n961 B.n30 585
R1415 B.n30 B.n29 585
R1416 B.n960 B.n959 585
R1417 B.n959 B.n958 585
R1418 B.n32 B.n31 585
R1419 B.n957 B.n32 585
R1420 B.n955 B.n954 585
R1421 B.n956 B.n955 585
R1422 B.n953 B.n37 585
R1423 B.n37 B.n36 585
R1424 B.n952 B.n951 585
R1425 B.n951 B.n950 585
R1426 B.n39 B.n38 585
R1427 B.n949 B.n39 585
R1428 B.n947 B.n946 585
R1429 B.n948 B.n947 585
R1430 B.n945 B.n44 585
R1431 B.n44 B.n43 585
R1432 B.n944 B.n943 585
R1433 B.n943 B.n942 585
R1434 B.n46 B.n45 585
R1435 B.n941 B.n46 585
R1436 B.n939 B.n938 585
R1437 B.n940 B.n939 585
R1438 B.n937 B.n51 585
R1439 B.n51 B.n50 585
R1440 B.n936 B.n935 585
R1441 B.n935 B.n934 585
R1442 B.n53 B.n52 585
R1443 B.n933 B.n53 585
R1444 B.n931 B.n930 585
R1445 B.n932 B.n931 585
R1446 B.n929 B.n58 585
R1447 B.n58 B.n57 585
R1448 B.n928 B.n927 585
R1449 B.n927 B.n926 585
R1450 B.n60 B.n59 585
R1451 B.n925 B.n60 585
R1452 B.n992 B.n991 585
R1453 B.n991 B.n990 585
R1454 B.n776 B.n450 526.135
R1455 B.n133 B.n60 526.135
R1456 B.n780 B.n452 526.135
R1457 B.n923 B.n62 526.135
R1458 B.n521 B.t12 471.396
R1459 B.n128 B.t4 471.396
R1460 B.n519 B.t9 471.396
R1461 B.n130 B.t14 471.396
R1462 B.n522 B.t11 389.553
R1463 B.n129 B.t5 389.553
R1464 B.n520 B.t8 389.553
R1465 B.n131 B.t15 389.553
R1466 B.n521 B.t10 322.353
R1467 B.n519 B.t6 322.353
R1468 B.n130 B.t13 322.353
R1469 B.n128 B.t2 322.353
R1470 B.n924 B.n126 256.663
R1471 B.n924 B.n125 256.663
R1472 B.n924 B.n124 256.663
R1473 B.n924 B.n123 256.663
R1474 B.n924 B.n122 256.663
R1475 B.n924 B.n121 256.663
R1476 B.n924 B.n120 256.663
R1477 B.n924 B.n119 256.663
R1478 B.n924 B.n118 256.663
R1479 B.n924 B.n117 256.663
R1480 B.n924 B.n116 256.663
R1481 B.n924 B.n115 256.663
R1482 B.n924 B.n114 256.663
R1483 B.n924 B.n113 256.663
R1484 B.n924 B.n112 256.663
R1485 B.n924 B.n111 256.663
R1486 B.n924 B.n110 256.663
R1487 B.n924 B.n109 256.663
R1488 B.n924 B.n108 256.663
R1489 B.n924 B.n107 256.663
R1490 B.n924 B.n106 256.663
R1491 B.n924 B.n105 256.663
R1492 B.n924 B.n104 256.663
R1493 B.n924 B.n103 256.663
R1494 B.n924 B.n102 256.663
R1495 B.n924 B.n101 256.663
R1496 B.n924 B.n100 256.663
R1497 B.n924 B.n99 256.663
R1498 B.n924 B.n98 256.663
R1499 B.n924 B.n97 256.663
R1500 B.n924 B.n96 256.663
R1501 B.n924 B.n95 256.663
R1502 B.n924 B.n94 256.663
R1503 B.n924 B.n93 256.663
R1504 B.n924 B.n92 256.663
R1505 B.n924 B.n91 256.663
R1506 B.n924 B.n90 256.663
R1507 B.n924 B.n89 256.663
R1508 B.n924 B.n88 256.663
R1509 B.n924 B.n87 256.663
R1510 B.n924 B.n86 256.663
R1511 B.n924 B.n85 256.663
R1512 B.n924 B.n84 256.663
R1513 B.n924 B.n83 256.663
R1514 B.n924 B.n82 256.663
R1515 B.n924 B.n81 256.663
R1516 B.n924 B.n80 256.663
R1517 B.n924 B.n79 256.663
R1518 B.n924 B.n78 256.663
R1519 B.n924 B.n77 256.663
R1520 B.n924 B.n76 256.663
R1521 B.n924 B.n75 256.663
R1522 B.n924 B.n74 256.663
R1523 B.n924 B.n73 256.663
R1524 B.n924 B.n72 256.663
R1525 B.n924 B.n71 256.663
R1526 B.n924 B.n70 256.663
R1527 B.n924 B.n69 256.663
R1528 B.n924 B.n68 256.663
R1529 B.n924 B.n67 256.663
R1530 B.n924 B.n66 256.663
R1531 B.n924 B.n65 256.663
R1532 B.n924 B.n64 256.663
R1533 B.n924 B.n63 256.663
R1534 B.n778 B.n777 256.663
R1535 B.n778 B.n455 256.663
R1536 B.n778 B.n456 256.663
R1537 B.n778 B.n457 256.663
R1538 B.n778 B.n458 256.663
R1539 B.n778 B.n459 256.663
R1540 B.n778 B.n460 256.663
R1541 B.n778 B.n461 256.663
R1542 B.n778 B.n462 256.663
R1543 B.n778 B.n463 256.663
R1544 B.n778 B.n464 256.663
R1545 B.n778 B.n465 256.663
R1546 B.n778 B.n466 256.663
R1547 B.n778 B.n467 256.663
R1548 B.n778 B.n468 256.663
R1549 B.n778 B.n469 256.663
R1550 B.n778 B.n470 256.663
R1551 B.n778 B.n471 256.663
R1552 B.n778 B.n472 256.663
R1553 B.n778 B.n473 256.663
R1554 B.n778 B.n474 256.663
R1555 B.n778 B.n475 256.663
R1556 B.n778 B.n476 256.663
R1557 B.n778 B.n477 256.663
R1558 B.n778 B.n478 256.663
R1559 B.n778 B.n479 256.663
R1560 B.n778 B.n480 256.663
R1561 B.n778 B.n481 256.663
R1562 B.n778 B.n482 256.663
R1563 B.n778 B.n483 256.663
R1564 B.n778 B.n484 256.663
R1565 B.n778 B.n485 256.663
R1566 B.n778 B.n486 256.663
R1567 B.n778 B.n487 256.663
R1568 B.n778 B.n488 256.663
R1569 B.n778 B.n489 256.663
R1570 B.n778 B.n490 256.663
R1571 B.n778 B.n491 256.663
R1572 B.n778 B.n492 256.663
R1573 B.n778 B.n493 256.663
R1574 B.n778 B.n494 256.663
R1575 B.n778 B.n495 256.663
R1576 B.n778 B.n496 256.663
R1577 B.n778 B.n497 256.663
R1578 B.n778 B.n498 256.663
R1579 B.n778 B.n499 256.663
R1580 B.n778 B.n500 256.663
R1581 B.n778 B.n501 256.663
R1582 B.n778 B.n502 256.663
R1583 B.n778 B.n503 256.663
R1584 B.n778 B.n504 256.663
R1585 B.n778 B.n505 256.663
R1586 B.n778 B.n506 256.663
R1587 B.n778 B.n507 256.663
R1588 B.n778 B.n508 256.663
R1589 B.n778 B.n509 256.663
R1590 B.n778 B.n510 256.663
R1591 B.n778 B.n511 256.663
R1592 B.n778 B.n512 256.663
R1593 B.n778 B.n513 256.663
R1594 B.n778 B.n514 256.663
R1595 B.n778 B.n515 256.663
R1596 B.n778 B.n516 256.663
R1597 B.n779 B.n778 256.663
R1598 B.n786 B.n450 163.367
R1599 B.n786 B.n448 163.367
R1600 B.n790 B.n448 163.367
R1601 B.n790 B.n442 163.367
R1602 B.n798 B.n442 163.367
R1603 B.n798 B.n440 163.367
R1604 B.n802 B.n440 163.367
R1605 B.n802 B.n434 163.367
R1606 B.n810 B.n434 163.367
R1607 B.n810 B.n432 163.367
R1608 B.n814 B.n432 163.367
R1609 B.n814 B.n426 163.367
R1610 B.n822 B.n426 163.367
R1611 B.n822 B.n424 163.367
R1612 B.n826 B.n424 163.367
R1613 B.n826 B.n418 163.367
R1614 B.n834 B.n418 163.367
R1615 B.n834 B.n416 163.367
R1616 B.n838 B.n416 163.367
R1617 B.n838 B.n410 163.367
R1618 B.n846 B.n410 163.367
R1619 B.n846 B.n408 163.367
R1620 B.n850 B.n408 163.367
R1621 B.n850 B.n402 163.367
R1622 B.n858 B.n402 163.367
R1623 B.n858 B.n400 163.367
R1624 B.n862 B.n400 163.367
R1625 B.n862 B.n394 163.367
R1626 B.n871 B.n394 163.367
R1627 B.n871 B.n392 163.367
R1628 B.n875 B.n392 163.367
R1629 B.n875 B.n2 163.367
R1630 B.n991 B.n2 163.367
R1631 B.n991 B.n3 163.367
R1632 B.n987 B.n3 163.367
R1633 B.n987 B.n9 163.367
R1634 B.n983 B.n9 163.367
R1635 B.n983 B.n11 163.367
R1636 B.n979 B.n11 163.367
R1637 B.n979 B.n16 163.367
R1638 B.n975 B.n16 163.367
R1639 B.n975 B.n18 163.367
R1640 B.n971 B.n18 163.367
R1641 B.n971 B.n23 163.367
R1642 B.n967 B.n23 163.367
R1643 B.n967 B.n25 163.367
R1644 B.n963 B.n25 163.367
R1645 B.n963 B.n30 163.367
R1646 B.n959 B.n30 163.367
R1647 B.n959 B.n32 163.367
R1648 B.n955 B.n32 163.367
R1649 B.n955 B.n37 163.367
R1650 B.n951 B.n37 163.367
R1651 B.n951 B.n39 163.367
R1652 B.n947 B.n39 163.367
R1653 B.n947 B.n44 163.367
R1654 B.n943 B.n44 163.367
R1655 B.n943 B.n46 163.367
R1656 B.n939 B.n46 163.367
R1657 B.n939 B.n51 163.367
R1658 B.n935 B.n51 163.367
R1659 B.n935 B.n53 163.367
R1660 B.n931 B.n53 163.367
R1661 B.n931 B.n58 163.367
R1662 B.n927 B.n58 163.367
R1663 B.n927 B.n60 163.367
R1664 B.n518 B.n517 163.367
R1665 B.n771 B.n517 163.367
R1666 B.n769 B.n768 163.367
R1667 B.n765 B.n764 163.367
R1668 B.n761 B.n760 163.367
R1669 B.n757 B.n756 163.367
R1670 B.n753 B.n752 163.367
R1671 B.n749 B.n748 163.367
R1672 B.n745 B.n744 163.367
R1673 B.n741 B.n740 163.367
R1674 B.n737 B.n736 163.367
R1675 B.n733 B.n732 163.367
R1676 B.n729 B.n728 163.367
R1677 B.n725 B.n724 163.367
R1678 B.n721 B.n720 163.367
R1679 B.n717 B.n716 163.367
R1680 B.n713 B.n712 163.367
R1681 B.n709 B.n708 163.367
R1682 B.n705 B.n704 163.367
R1683 B.n701 B.n700 163.367
R1684 B.n697 B.n696 163.367
R1685 B.n693 B.n692 163.367
R1686 B.n689 B.n688 163.367
R1687 B.n685 B.n684 163.367
R1688 B.n681 B.n680 163.367
R1689 B.n677 B.n676 163.367
R1690 B.n673 B.n672 163.367
R1691 B.n669 B.n668 163.367
R1692 B.n665 B.n664 163.367
R1693 B.n661 B.n660 163.367
R1694 B.n656 B.n655 163.367
R1695 B.n652 B.n651 163.367
R1696 B.n648 B.n647 163.367
R1697 B.n644 B.n643 163.367
R1698 B.n640 B.n639 163.367
R1699 B.n636 B.n635 163.367
R1700 B.n632 B.n631 163.367
R1701 B.n628 B.n627 163.367
R1702 B.n624 B.n623 163.367
R1703 B.n620 B.n619 163.367
R1704 B.n616 B.n615 163.367
R1705 B.n612 B.n611 163.367
R1706 B.n608 B.n607 163.367
R1707 B.n604 B.n603 163.367
R1708 B.n600 B.n599 163.367
R1709 B.n596 B.n595 163.367
R1710 B.n592 B.n591 163.367
R1711 B.n588 B.n587 163.367
R1712 B.n584 B.n583 163.367
R1713 B.n580 B.n579 163.367
R1714 B.n576 B.n575 163.367
R1715 B.n572 B.n571 163.367
R1716 B.n568 B.n567 163.367
R1717 B.n564 B.n563 163.367
R1718 B.n560 B.n559 163.367
R1719 B.n556 B.n555 163.367
R1720 B.n552 B.n551 163.367
R1721 B.n548 B.n547 163.367
R1722 B.n544 B.n543 163.367
R1723 B.n540 B.n539 163.367
R1724 B.n536 B.n535 163.367
R1725 B.n532 B.n531 163.367
R1726 B.n528 B.n527 163.367
R1727 B.n524 B.n454 163.367
R1728 B.n784 B.n452 163.367
R1729 B.n784 B.n446 163.367
R1730 B.n792 B.n446 163.367
R1731 B.n792 B.n444 163.367
R1732 B.n796 B.n444 163.367
R1733 B.n796 B.n438 163.367
R1734 B.n804 B.n438 163.367
R1735 B.n804 B.n436 163.367
R1736 B.n808 B.n436 163.367
R1737 B.n808 B.n430 163.367
R1738 B.n816 B.n430 163.367
R1739 B.n816 B.n428 163.367
R1740 B.n820 B.n428 163.367
R1741 B.n820 B.n422 163.367
R1742 B.n828 B.n422 163.367
R1743 B.n828 B.n420 163.367
R1744 B.n832 B.n420 163.367
R1745 B.n832 B.n414 163.367
R1746 B.n840 B.n414 163.367
R1747 B.n840 B.n412 163.367
R1748 B.n844 B.n412 163.367
R1749 B.n844 B.n406 163.367
R1750 B.n852 B.n406 163.367
R1751 B.n852 B.n404 163.367
R1752 B.n856 B.n404 163.367
R1753 B.n856 B.n398 163.367
R1754 B.n864 B.n398 163.367
R1755 B.n864 B.n396 163.367
R1756 B.n869 B.n396 163.367
R1757 B.n869 B.n390 163.367
R1758 B.n877 B.n390 163.367
R1759 B.n878 B.n877 163.367
R1760 B.n878 B.n5 163.367
R1761 B.n6 B.n5 163.367
R1762 B.n7 B.n6 163.367
R1763 B.n883 B.n7 163.367
R1764 B.n883 B.n12 163.367
R1765 B.n13 B.n12 163.367
R1766 B.n14 B.n13 163.367
R1767 B.n888 B.n14 163.367
R1768 B.n888 B.n19 163.367
R1769 B.n20 B.n19 163.367
R1770 B.n21 B.n20 163.367
R1771 B.n893 B.n21 163.367
R1772 B.n893 B.n26 163.367
R1773 B.n27 B.n26 163.367
R1774 B.n28 B.n27 163.367
R1775 B.n898 B.n28 163.367
R1776 B.n898 B.n33 163.367
R1777 B.n34 B.n33 163.367
R1778 B.n35 B.n34 163.367
R1779 B.n903 B.n35 163.367
R1780 B.n903 B.n40 163.367
R1781 B.n41 B.n40 163.367
R1782 B.n42 B.n41 163.367
R1783 B.n908 B.n42 163.367
R1784 B.n908 B.n47 163.367
R1785 B.n48 B.n47 163.367
R1786 B.n49 B.n48 163.367
R1787 B.n913 B.n49 163.367
R1788 B.n913 B.n54 163.367
R1789 B.n55 B.n54 163.367
R1790 B.n56 B.n55 163.367
R1791 B.n918 B.n56 163.367
R1792 B.n918 B.n61 163.367
R1793 B.n62 B.n61 163.367
R1794 B.n137 B.n136 163.367
R1795 B.n141 B.n140 163.367
R1796 B.n145 B.n144 163.367
R1797 B.n149 B.n148 163.367
R1798 B.n153 B.n152 163.367
R1799 B.n157 B.n156 163.367
R1800 B.n161 B.n160 163.367
R1801 B.n165 B.n164 163.367
R1802 B.n169 B.n168 163.367
R1803 B.n173 B.n172 163.367
R1804 B.n177 B.n176 163.367
R1805 B.n181 B.n180 163.367
R1806 B.n185 B.n184 163.367
R1807 B.n189 B.n188 163.367
R1808 B.n193 B.n192 163.367
R1809 B.n197 B.n196 163.367
R1810 B.n201 B.n200 163.367
R1811 B.n205 B.n204 163.367
R1812 B.n209 B.n208 163.367
R1813 B.n213 B.n212 163.367
R1814 B.n217 B.n216 163.367
R1815 B.n221 B.n220 163.367
R1816 B.n225 B.n224 163.367
R1817 B.n229 B.n228 163.367
R1818 B.n233 B.n232 163.367
R1819 B.n237 B.n236 163.367
R1820 B.n241 B.n240 163.367
R1821 B.n245 B.n244 163.367
R1822 B.n249 B.n248 163.367
R1823 B.n253 B.n252 163.367
R1824 B.n257 B.n256 163.367
R1825 B.n261 B.n260 163.367
R1826 B.n265 B.n264 163.367
R1827 B.n269 B.n268 163.367
R1828 B.n274 B.n273 163.367
R1829 B.n278 B.n277 163.367
R1830 B.n282 B.n281 163.367
R1831 B.n286 B.n285 163.367
R1832 B.n290 B.n289 163.367
R1833 B.n294 B.n293 163.367
R1834 B.n298 B.n297 163.367
R1835 B.n302 B.n301 163.367
R1836 B.n306 B.n305 163.367
R1837 B.n310 B.n309 163.367
R1838 B.n314 B.n313 163.367
R1839 B.n318 B.n317 163.367
R1840 B.n322 B.n321 163.367
R1841 B.n326 B.n325 163.367
R1842 B.n330 B.n329 163.367
R1843 B.n334 B.n333 163.367
R1844 B.n338 B.n337 163.367
R1845 B.n342 B.n341 163.367
R1846 B.n346 B.n345 163.367
R1847 B.n350 B.n349 163.367
R1848 B.n354 B.n353 163.367
R1849 B.n358 B.n357 163.367
R1850 B.n362 B.n361 163.367
R1851 B.n366 B.n365 163.367
R1852 B.n370 B.n369 163.367
R1853 B.n374 B.n373 163.367
R1854 B.n378 B.n377 163.367
R1855 B.n382 B.n381 163.367
R1856 B.n386 B.n385 163.367
R1857 B.n923 B.n127 163.367
R1858 B.n522 B.n521 81.8429
R1859 B.n520 B.n519 81.8429
R1860 B.n131 B.n130 81.8429
R1861 B.n129 B.n128 81.8429
R1862 B.n777 B.n776 71.676
R1863 B.n771 B.n455 71.676
R1864 B.n768 B.n456 71.676
R1865 B.n764 B.n457 71.676
R1866 B.n760 B.n458 71.676
R1867 B.n756 B.n459 71.676
R1868 B.n752 B.n460 71.676
R1869 B.n748 B.n461 71.676
R1870 B.n744 B.n462 71.676
R1871 B.n740 B.n463 71.676
R1872 B.n736 B.n464 71.676
R1873 B.n732 B.n465 71.676
R1874 B.n728 B.n466 71.676
R1875 B.n724 B.n467 71.676
R1876 B.n720 B.n468 71.676
R1877 B.n716 B.n469 71.676
R1878 B.n712 B.n470 71.676
R1879 B.n708 B.n471 71.676
R1880 B.n704 B.n472 71.676
R1881 B.n700 B.n473 71.676
R1882 B.n696 B.n474 71.676
R1883 B.n692 B.n475 71.676
R1884 B.n688 B.n476 71.676
R1885 B.n684 B.n477 71.676
R1886 B.n680 B.n478 71.676
R1887 B.n676 B.n479 71.676
R1888 B.n672 B.n480 71.676
R1889 B.n668 B.n481 71.676
R1890 B.n664 B.n482 71.676
R1891 B.n660 B.n483 71.676
R1892 B.n655 B.n484 71.676
R1893 B.n651 B.n485 71.676
R1894 B.n647 B.n486 71.676
R1895 B.n643 B.n487 71.676
R1896 B.n639 B.n488 71.676
R1897 B.n635 B.n489 71.676
R1898 B.n631 B.n490 71.676
R1899 B.n627 B.n491 71.676
R1900 B.n623 B.n492 71.676
R1901 B.n619 B.n493 71.676
R1902 B.n615 B.n494 71.676
R1903 B.n611 B.n495 71.676
R1904 B.n607 B.n496 71.676
R1905 B.n603 B.n497 71.676
R1906 B.n599 B.n498 71.676
R1907 B.n595 B.n499 71.676
R1908 B.n591 B.n500 71.676
R1909 B.n587 B.n501 71.676
R1910 B.n583 B.n502 71.676
R1911 B.n579 B.n503 71.676
R1912 B.n575 B.n504 71.676
R1913 B.n571 B.n505 71.676
R1914 B.n567 B.n506 71.676
R1915 B.n563 B.n507 71.676
R1916 B.n559 B.n508 71.676
R1917 B.n555 B.n509 71.676
R1918 B.n551 B.n510 71.676
R1919 B.n547 B.n511 71.676
R1920 B.n543 B.n512 71.676
R1921 B.n539 B.n513 71.676
R1922 B.n535 B.n514 71.676
R1923 B.n531 B.n515 71.676
R1924 B.n527 B.n516 71.676
R1925 B.n779 B.n454 71.676
R1926 B.n133 B.n63 71.676
R1927 B.n137 B.n64 71.676
R1928 B.n141 B.n65 71.676
R1929 B.n145 B.n66 71.676
R1930 B.n149 B.n67 71.676
R1931 B.n153 B.n68 71.676
R1932 B.n157 B.n69 71.676
R1933 B.n161 B.n70 71.676
R1934 B.n165 B.n71 71.676
R1935 B.n169 B.n72 71.676
R1936 B.n173 B.n73 71.676
R1937 B.n177 B.n74 71.676
R1938 B.n181 B.n75 71.676
R1939 B.n185 B.n76 71.676
R1940 B.n189 B.n77 71.676
R1941 B.n193 B.n78 71.676
R1942 B.n197 B.n79 71.676
R1943 B.n201 B.n80 71.676
R1944 B.n205 B.n81 71.676
R1945 B.n209 B.n82 71.676
R1946 B.n213 B.n83 71.676
R1947 B.n217 B.n84 71.676
R1948 B.n221 B.n85 71.676
R1949 B.n225 B.n86 71.676
R1950 B.n229 B.n87 71.676
R1951 B.n233 B.n88 71.676
R1952 B.n237 B.n89 71.676
R1953 B.n241 B.n90 71.676
R1954 B.n245 B.n91 71.676
R1955 B.n249 B.n92 71.676
R1956 B.n253 B.n93 71.676
R1957 B.n257 B.n94 71.676
R1958 B.n261 B.n95 71.676
R1959 B.n265 B.n96 71.676
R1960 B.n269 B.n97 71.676
R1961 B.n274 B.n98 71.676
R1962 B.n278 B.n99 71.676
R1963 B.n282 B.n100 71.676
R1964 B.n286 B.n101 71.676
R1965 B.n290 B.n102 71.676
R1966 B.n294 B.n103 71.676
R1967 B.n298 B.n104 71.676
R1968 B.n302 B.n105 71.676
R1969 B.n306 B.n106 71.676
R1970 B.n310 B.n107 71.676
R1971 B.n314 B.n108 71.676
R1972 B.n318 B.n109 71.676
R1973 B.n322 B.n110 71.676
R1974 B.n326 B.n111 71.676
R1975 B.n330 B.n112 71.676
R1976 B.n334 B.n113 71.676
R1977 B.n338 B.n114 71.676
R1978 B.n342 B.n115 71.676
R1979 B.n346 B.n116 71.676
R1980 B.n350 B.n117 71.676
R1981 B.n354 B.n118 71.676
R1982 B.n358 B.n119 71.676
R1983 B.n362 B.n120 71.676
R1984 B.n366 B.n121 71.676
R1985 B.n370 B.n122 71.676
R1986 B.n374 B.n123 71.676
R1987 B.n378 B.n124 71.676
R1988 B.n382 B.n125 71.676
R1989 B.n386 B.n126 71.676
R1990 B.n127 B.n126 71.676
R1991 B.n385 B.n125 71.676
R1992 B.n381 B.n124 71.676
R1993 B.n377 B.n123 71.676
R1994 B.n373 B.n122 71.676
R1995 B.n369 B.n121 71.676
R1996 B.n365 B.n120 71.676
R1997 B.n361 B.n119 71.676
R1998 B.n357 B.n118 71.676
R1999 B.n353 B.n117 71.676
R2000 B.n349 B.n116 71.676
R2001 B.n345 B.n115 71.676
R2002 B.n341 B.n114 71.676
R2003 B.n337 B.n113 71.676
R2004 B.n333 B.n112 71.676
R2005 B.n329 B.n111 71.676
R2006 B.n325 B.n110 71.676
R2007 B.n321 B.n109 71.676
R2008 B.n317 B.n108 71.676
R2009 B.n313 B.n107 71.676
R2010 B.n309 B.n106 71.676
R2011 B.n305 B.n105 71.676
R2012 B.n301 B.n104 71.676
R2013 B.n297 B.n103 71.676
R2014 B.n293 B.n102 71.676
R2015 B.n289 B.n101 71.676
R2016 B.n285 B.n100 71.676
R2017 B.n281 B.n99 71.676
R2018 B.n277 B.n98 71.676
R2019 B.n273 B.n97 71.676
R2020 B.n268 B.n96 71.676
R2021 B.n264 B.n95 71.676
R2022 B.n260 B.n94 71.676
R2023 B.n256 B.n93 71.676
R2024 B.n252 B.n92 71.676
R2025 B.n248 B.n91 71.676
R2026 B.n244 B.n90 71.676
R2027 B.n240 B.n89 71.676
R2028 B.n236 B.n88 71.676
R2029 B.n232 B.n87 71.676
R2030 B.n228 B.n86 71.676
R2031 B.n224 B.n85 71.676
R2032 B.n220 B.n84 71.676
R2033 B.n216 B.n83 71.676
R2034 B.n212 B.n82 71.676
R2035 B.n208 B.n81 71.676
R2036 B.n204 B.n80 71.676
R2037 B.n200 B.n79 71.676
R2038 B.n196 B.n78 71.676
R2039 B.n192 B.n77 71.676
R2040 B.n188 B.n76 71.676
R2041 B.n184 B.n75 71.676
R2042 B.n180 B.n74 71.676
R2043 B.n176 B.n73 71.676
R2044 B.n172 B.n72 71.676
R2045 B.n168 B.n71 71.676
R2046 B.n164 B.n70 71.676
R2047 B.n160 B.n69 71.676
R2048 B.n156 B.n68 71.676
R2049 B.n152 B.n67 71.676
R2050 B.n148 B.n66 71.676
R2051 B.n144 B.n65 71.676
R2052 B.n140 B.n64 71.676
R2053 B.n136 B.n63 71.676
R2054 B.n777 B.n518 71.676
R2055 B.n769 B.n455 71.676
R2056 B.n765 B.n456 71.676
R2057 B.n761 B.n457 71.676
R2058 B.n757 B.n458 71.676
R2059 B.n753 B.n459 71.676
R2060 B.n749 B.n460 71.676
R2061 B.n745 B.n461 71.676
R2062 B.n741 B.n462 71.676
R2063 B.n737 B.n463 71.676
R2064 B.n733 B.n464 71.676
R2065 B.n729 B.n465 71.676
R2066 B.n725 B.n466 71.676
R2067 B.n721 B.n467 71.676
R2068 B.n717 B.n468 71.676
R2069 B.n713 B.n469 71.676
R2070 B.n709 B.n470 71.676
R2071 B.n705 B.n471 71.676
R2072 B.n701 B.n472 71.676
R2073 B.n697 B.n473 71.676
R2074 B.n693 B.n474 71.676
R2075 B.n689 B.n475 71.676
R2076 B.n685 B.n476 71.676
R2077 B.n681 B.n477 71.676
R2078 B.n677 B.n478 71.676
R2079 B.n673 B.n479 71.676
R2080 B.n669 B.n480 71.676
R2081 B.n665 B.n481 71.676
R2082 B.n661 B.n482 71.676
R2083 B.n656 B.n483 71.676
R2084 B.n652 B.n484 71.676
R2085 B.n648 B.n485 71.676
R2086 B.n644 B.n486 71.676
R2087 B.n640 B.n487 71.676
R2088 B.n636 B.n488 71.676
R2089 B.n632 B.n489 71.676
R2090 B.n628 B.n490 71.676
R2091 B.n624 B.n491 71.676
R2092 B.n620 B.n492 71.676
R2093 B.n616 B.n493 71.676
R2094 B.n612 B.n494 71.676
R2095 B.n608 B.n495 71.676
R2096 B.n604 B.n496 71.676
R2097 B.n600 B.n497 71.676
R2098 B.n596 B.n498 71.676
R2099 B.n592 B.n499 71.676
R2100 B.n588 B.n500 71.676
R2101 B.n584 B.n501 71.676
R2102 B.n580 B.n502 71.676
R2103 B.n576 B.n503 71.676
R2104 B.n572 B.n504 71.676
R2105 B.n568 B.n505 71.676
R2106 B.n564 B.n506 71.676
R2107 B.n560 B.n507 71.676
R2108 B.n556 B.n508 71.676
R2109 B.n552 B.n509 71.676
R2110 B.n548 B.n510 71.676
R2111 B.n544 B.n511 71.676
R2112 B.n540 B.n512 71.676
R2113 B.n536 B.n513 71.676
R2114 B.n532 B.n514 71.676
R2115 B.n528 B.n515 71.676
R2116 B.n524 B.n516 71.676
R2117 B.n780 B.n779 71.676
R2118 B.n523 B.n522 59.5399
R2119 B.n658 B.n520 59.5399
R2120 B.n132 B.n131 59.5399
R2121 B.n271 B.n129 59.5399
R2122 B.n778 B.n451 55.6908
R2123 B.n925 B.n924 55.6908
R2124 B.n134 B.n59 34.1859
R2125 B.n922 B.n921 34.1859
R2126 B.n782 B.n781 34.1859
R2127 B.n775 B.n449 34.1859
R2128 B.n785 B.n451 31.8235
R2129 B.n785 B.n447 31.8235
R2130 B.n791 B.n447 31.8235
R2131 B.n791 B.n443 31.8235
R2132 B.n797 B.n443 31.8235
R2133 B.n797 B.n439 31.8235
R2134 B.n803 B.n439 31.8235
R2135 B.n803 B.n435 31.8235
R2136 B.n809 B.n435 31.8235
R2137 B.n815 B.n431 31.8235
R2138 B.n815 B.n427 31.8235
R2139 B.n821 B.n427 31.8235
R2140 B.n821 B.n423 31.8235
R2141 B.n827 B.n423 31.8235
R2142 B.n827 B.n419 31.8235
R2143 B.n833 B.n419 31.8235
R2144 B.n833 B.n415 31.8235
R2145 B.n839 B.n415 31.8235
R2146 B.n839 B.n411 31.8235
R2147 B.n845 B.n411 31.8235
R2148 B.n845 B.n407 31.8235
R2149 B.n851 B.n407 31.8235
R2150 B.n851 B.n403 31.8235
R2151 B.n857 B.n403 31.8235
R2152 B.n863 B.n399 31.8235
R2153 B.n863 B.n395 31.8235
R2154 B.n870 B.n395 31.8235
R2155 B.n870 B.n391 31.8235
R2156 B.n876 B.n391 31.8235
R2157 B.n876 B.n4 31.8235
R2158 B.n990 B.n4 31.8235
R2159 B.n990 B.n989 31.8235
R2160 B.n989 B.n988 31.8235
R2161 B.n988 B.n8 31.8235
R2162 B.n982 B.n8 31.8235
R2163 B.n982 B.n981 31.8235
R2164 B.n981 B.n980 31.8235
R2165 B.n980 B.n15 31.8235
R2166 B.n974 B.n973 31.8235
R2167 B.n973 B.n972 31.8235
R2168 B.n972 B.n22 31.8235
R2169 B.n966 B.n22 31.8235
R2170 B.n966 B.n965 31.8235
R2171 B.n965 B.n964 31.8235
R2172 B.n964 B.n29 31.8235
R2173 B.n958 B.n29 31.8235
R2174 B.n958 B.n957 31.8235
R2175 B.n957 B.n956 31.8235
R2176 B.n956 B.n36 31.8235
R2177 B.n950 B.n36 31.8235
R2178 B.n950 B.n949 31.8235
R2179 B.n949 B.n948 31.8235
R2180 B.n948 B.n43 31.8235
R2181 B.n942 B.n941 31.8235
R2182 B.n941 B.n940 31.8235
R2183 B.n940 B.n50 31.8235
R2184 B.n934 B.n50 31.8235
R2185 B.n934 B.n933 31.8235
R2186 B.n933 B.n932 31.8235
R2187 B.n932 B.n57 31.8235
R2188 B.n926 B.n57 31.8235
R2189 B.n926 B.n925 31.8235
R2190 B.t0 B.n399 25.7397
R2191 B.t1 B.n15 25.7397
R2192 B.n809 B.t7 18.2519
R2193 B.n942 B.t3 18.2519
R2194 B B.n992 18.0485
R2195 B.t7 B.n431 13.5721
R2196 B.t3 B.n43 13.5721
R2197 B.n135 B.n134 10.6151
R2198 B.n138 B.n135 10.6151
R2199 B.n139 B.n138 10.6151
R2200 B.n142 B.n139 10.6151
R2201 B.n143 B.n142 10.6151
R2202 B.n146 B.n143 10.6151
R2203 B.n147 B.n146 10.6151
R2204 B.n150 B.n147 10.6151
R2205 B.n151 B.n150 10.6151
R2206 B.n154 B.n151 10.6151
R2207 B.n155 B.n154 10.6151
R2208 B.n158 B.n155 10.6151
R2209 B.n159 B.n158 10.6151
R2210 B.n162 B.n159 10.6151
R2211 B.n163 B.n162 10.6151
R2212 B.n166 B.n163 10.6151
R2213 B.n167 B.n166 10.6151
R2214 B.n170 B.n167 10.6151
R2215 B.n171 B.n170 10.6151
R2216 B.n174 B.n171 10.6151
R2217 B.n175 B.n174 10.6151
R2218 B.n178 B.n175 10.6151
R2219 B.n179 B.n178 10.6151
R2220 B.n182 B.n179 10.6151
R2221 B.n183 B.n182 10.6151
R2222 B.n186 B.n183 10.6151
R2223 B.n187 B.n186 10.6151
R2224 B.n190 B.n187 10.6151
R2225 B.n191 B.n190 10.6151
R2226 B.n194 B.n191 10.6151
R2227 B.n195 B.n194 10.6151
R2228 B.n198 B.n195 10.6151
R2229 B.n199 B.n198 10.6151
R2230 B.n202 B.n199 10.6151
R2231 B.n203 B.n202 10.6151
R2232 B.n206 B.n203 10.6151
R2233 B.n207 B.n206 10.6151
R2234 B.n210 B.n207 10.6151
R2235 B.n211 B.n210 10.6151
R2236 B.n214 B.n211 10.6151
R2237 B.n215 B.n214 10.6151
R2238 B.n218 B.n215 10.6151
R2239 B.n219 B.n218 10.6151
R2240 B.n222 B.n219 10.6151
R2241 B.n223 B.n222 10.6151
R2242 B.n226 B.n223 10.6151
R2243 B.n227 B.n226 10.6151
R2244 B.n230 B.n227 10.6151
R2245 B.n231 B.n230 10.6151
R2246 B.n234 B.n231 10.6151
R2247 B.n235 B.n234 10.6151
R2248 B.n238 B.n235 10.6151
R2249 B.n239 B.n238 10.6151
R2250 B.n242 B.n239 10.6151
R2251 B.n243 B.n242 10.6151
R2252 B.n246 B.n243 10.6151
R2253 B.n247 B.n246 10.6151
R2254 B.n250 B.n247 10.6151
R2255 B.n251 B.n250 10.6151
R2256 B.n255 B.n254 10.6151
R2257 B.n258 B.n255 10.6151
R2258 B.n259 B.n258 10.6151
R2259 B.n262 B.n259 10.6151
R2260 B.n263 B.n262 10.6151
R2261 B.n266 B.n263 10.6151
R2262 B.n267 B.n266 10.6151
R2263 B.n270 B.n267 10.6151
R2264 B.n275 B.n272 10.6151
R2265 B.n276 B.n275 10.6151
R2266 B.n279 B.n276 10.6151
R2267 B.n280 B.n279 10.6151
R2268 B.n283 B.n280 10.6151
R2269 B.n284 B.n283 10.6151
R2270 B.n287 B.n284 10.6151
R2271 B.n288 B.n287 10.6151
R2272 B.n291 B.n288 10.6151
R2273 B.n292 B.n291 10.6151
R2274 B.n295 B.n292 10.6151
R2275 B.n296 B.n295 10.6151
R2276 B.n299 B.n296 10.6151
R2277 B.n300 B.n299 10.6151
R2278 B.n303 B.n300 10.6151
R2279 B.n304 B.n303 10.6151
R2280 B.n307 B.n304 10.6151
R2281 B.n308 B.n307 10.6151
R2282 B.n311 B.n308 10.6151
R2283 B.n312 B.n311 10.6151
R2284 B.n315 B.n312 10.6151
R2285 B.n316 B.n315 10.6151
R2286 B.n319 B.n316 10.6151
R2287 B.n320 B.n319 10.6151
R2288 B.n323 B.n320 10.6151
R2289 B.n324 B.n323 10.6151
R2290 B.n327 B.n324 10.6151
R2291 B.n328 B.n327 10.6151
R2292 B.n331 B.n328 10.6151
R2293 B.n332 B.n331 10.6151
R2294 B.n335 B.n332 10.6151
R2295 B.n336 B.n335 10.6151
R2296 B.n339 B.n336 10.6151
R2297 B.n340 B.n339 10.6151
R2298 B.n343 B.n340 10.6151
R2299 B.n344 B.n343 10.6151
R2300 B.n347 B.n344 10.6151
R2301 B.n348 B.n347 10.6151
R2302 B.n351 B.n348 10.6151
R2303 B.n352 B.n351 10.6151
R2304 B.n355 B.n352 10.6151
R2305 B.n356 B.n355 10.6151
R2306 B.n359 B.n356 10.6151
R2307 B.n360 B.n359 10.6151
R2308 B.n363 B.n360 10.6151
R2309 B.n364 B.n363 10.6151
R2310 B.n367 B.n364 10.6151
R2311 B.n368 B.n367 10.6151
R2312 B.n371 B.n368 10.6151
R2313 B.n372 B.n371 10.6151
R2314 B.n375 B.n372 10.6151
R2315 B.n376 B.n375 10.6151
R2316 B.n379 B.n376 10.6151
R2317 B.n380 B.n379 10.6151
R2318 B.n383 B.n380 10.6151
R2319 B.n384 B.n383 10.6151
R2320 B.n387 B.n384 10.6151
R2321 B.n388 B.n387 10.6151
R2322 B.n922 B.n388 10.6151
R2323 B.n783 B.n782 10.6151
R2324 B.n783 B.n445 10.6151
R2325 B.n793 B.n445 10.6151
R2326 B.n794 B.n793 10.6151
R2327 B.n795 B.n794 10.6151
R2328 B.n795 B.n437 10.6151
R2329 B.n805 B.n437 10.6151
R2330 B.n806 B.n805 10.6151
R2331 B.n807 B.n806 10.6151
R2332 B.n807 B.n429 10.6151
R2333 B.n817 B.n429 10.6151
R2334 B.n818 B.n817 10.6151
R2335 B.n819 B.n818 10.6151
R2336 B.n819 B.n421 10.6151
R2337 B.n829 B.n421 10.6151
R2338 B.n830 B.n829 10.6151
R2339 B.n831 B.n830 10.6151
R2340 B.n831 B.n413 10.6151
R2341 B.n841 B.n413 10.6151
R2342 B.n842 B.n841 10.6151
R2343 B.n843 B.n842 10.6151
R2344 B.n843 B.n405 10.6151
R2345 B.n853 B.n405 10.6151
R2346 B.n854 B.n853 10.6151
R2347 B.n855 B.n854 10.6151
R2348 B.n855 B.n397 10.6151
R2349 B.n865 B.n397 10.6151
R2350 B.n866 B.n865 10.6151
R2351 B.n868 B.n866 10.6151
R2352 B.n868 B.n867 10.6151
R2353 B.n867 B.n389 10.6151
R2354 B.n879 B.n389 10.6151
R2355 B.n880 B.n879 10.6151
R2356 B.n881 B.n880 10.6151
R2357 B.n882 B.n881 10.6151
R2358 B.n884 B.n882 10.6151
R2359 B.n885 B.n884 10.6151
R2360 B.n886 B.n885 10.6151
R2361 B.n887 B.n886 10.6151
R2362 B.n889 B.n887 10.6151
R2363 B.n890 B.n889 10.6151
R2364 B.n891 B.n890 10.6151
R2365 B.n892 B.n891 10.6151
R2366 B.n894 B.n892 10.6151
R2367 B.n895 B.n894 10.6151
R2368 B.n896 B.n895 10.6151
R2369 B.n897 B.n896 10.6151
R2370 B.n899 B.n897 10.6151
R2371 B.n900 B.n899 10.6151
R2372 B.n901 B.n900 10.6151
R2373 B.n902 B.n901 10.6151
R2374 B.n904 B.n902 10.6151
R2375 B.n905 B.n904 10.6151
R2376 B.n906 B.n905 10.6151
R2377 B.n907 B.n906 10.6151
R2378 B.n909 B.n907 10.6151
R2379 B.n910 B.n909 10.6151
R2380 B.n911 B.n910 10.6151
R2381 B.n912 B.n911 10.6151
R2382 B.n914 B.n912 10.6151
R2383 B.n915 B.n914 10.6151
R2384 B.n916 B.n915 10.6151
R2385 B.n917 B.n916 10.6151
R2386 B.n919 B.n917 10.6151
R2387 B.n920 B.n919 10.6151
R2388 B.n921 B.n920 10.6151
R2389 B.n775 B.n774 10.6151
R2390 B.n774 B.n773 10.6151
R2391 B.n773 B.n772 10.6151
R2392 B.n772 B.n770 10.6151
R2393 B.n770 B.n767 10.6151
R2394 B.n767 B.n766 10.6151
R2395 B.n766 B.n763 10.6151
R2396 B.n763 B.n762 10.6151
R2397 B.n762 B.n759 10.6151
R2398 B.n759 B.n758 10.6151
R2399 B.n758 B.n755 10.6151
R2400 B.n755 B.n754 10.6151
R2401 B.n754 B.n751 10.6151
R2402 B.n751 B.n750 10.6151
R2403 B.n750 B.n747 10.6151
R2404 B.n747 B.n746 10.6151
R2405 B.n746 B.n743 10.6151
R2406 B.n743 B.n742 10.6151
R2407 B.n742 B.n739 10.6151
R2408 B.n739 B.n738 10.6151
R2409 B.n738 B.n735 10.6151
R2410 B.n735 B.n734 10.6151
R2411 B.n734 B.n731 10.6151
R2412 B.n731 B.n730 10.6151
R2413 B.n730 B.n727 10.6151
R2414 B.n727 B.n726 10.6151
R2415 B.n726 B.n723 10.6151
R2416 B.n723 B.n722 10.6151
R2417 B.n722 B.n719 10.6151
R2418 B.n719 B.n718 10.6151
R2419 B.n718 B.n715 10.6151
R2420 B.n715 B.n714 10.6151
R2421 B.n714 B.n711 10.6151
R2422 B.n711 B.n710 10.6151
R2423 B.n710 B.n707 10.6151
R2424 B.n707 B.n706 10.6151
R2425 B.n706 B.n703 10.6151
R2426 B.n703 B.n702 10.6151
R2427 B.n702 B.n699 10.6151
R2428 B.n699 B.n698 10.6151
R2429 B.n698 B.n695 10.6151
R2430 B.n695 B.n694 10.6151
R2431 B.n694 B.n691 10.6151
R2432 B.n691 B.n690 10.6151
R2433 B.n690 B.n687 10.6151
R2434 B.n687 B.n686 10.6151
R2435 B.n686 B.n683 10.6151
R2436 B.n683 B.n682 10.6151
R2437 B.n682 B.n679 10.6151
R2438 B.n679 B.n678 10.6151
R2439 B.n678 B.n675 10.6151
R2440 B.n675 B.n674 10.6151
R2441 B.n674 B.n671 10.6151
R2442 B.n671 B.n670 10.6151
R2443 B.n670 B.n667 10.6151
R2444 B.n667 B.n666 10.6151
R2445 B.n666 B.n663 10.6151
R2446 B.n663 B.n662 10.6151
R2447 B.n662 B.n659 10.6151
R2448 B.n657 B.n654 10.6151
R2449 B.n654 B.n653 10.6151
R2450 B.n653 B.n650 10.6151
R2451 B.n650 B.n649 10.6151
R2452 B.n649 B.n646 10.6151
R2453 B.n646 B.n645 10.6151
R2454 B.n645 B.n642 10.6151
R2455 B.n642 B.n641 10.6151
R2456 B.n638 B.n637 10.6151
R2457 B.n637 B.n634 10.6151
R2458 B.n634 B.n633 10.6151
R2459 B.n633 B.n630 10.6151
R2460 B.n630 B.n629 10.6151
R2461 B.n629 B.n626 10.6151
R2462 B.n626 B.n625 10.6151
R2463 B.n625 B.n622 10.6151
R2464 B.n622 B.n621 10.6151
R2465 B.n621 B.n618 10.6151
R2466 B.n618 B.n617 10.6151
R2467 B.n617 B.n614 10.6151
R2468 B.n614 B.n613 10.6151
R2469 B.n613 B.n610 10.6151
R2470 B.n610 B.n609 10.6151
R2471 B.n609 B.n606 10.6151
R2472 B.n606 B.n605 10.6151
R2473 B.n605 B.n602 10.6151
R2474 B.n602 B.n601 10.6151
R2475 B.n601 B.n598 10.6151
R2476 B.n598 B.n597 10.6151
R2477 B.n597 B.n594 10.6151
R2478 B.n594 B.n593 10.6151
R2479 B.n593 B.n590 10.6151
R2480 B.n590 B.n589 10.6151
R2481 B.n589 B.n586 10.6151
R2482 B.n586 B.n585 10.6151
R2483 B.n585 B.n582 10.6151
R2484 B.n582 B.n581 10.6151
R2485 B.n581 B.n578 10.6151
R2486 B.n578 B.n577 10.6151
R2487 B.n577 B.n574 10.6151
R2488 B.n574 B.n573 10.6151
R2489 B.n573 B.n570 10.6151
R2490 B.n570 B.n569 10.6151
R2491 B.n569 B.n566 10.6151
R2492 B.n566 B.n565 10.6151
R2493 B.n565 B.n562 10.6151
R2494 B.n562 B.n561 10.6151
R2495 B.n561 B.n558 10.6151
R2496 B.n558 B.n557 10.6151
R2497 B.n557 B.n554 10.6151
R2498 B.n554 B.n553 10.6151
R2499 B.n553 B.n550 10.6151
R2500 B.n550 B.n549 10.6151
R2501 B.n549 B.n546 10.6151
R2502 B.n546 B.n545 10.6151
R2503 B.n545 B.n542 10.6151
R2504 B.n542 B.n541 10.6151
R2505 B.n541 B.n538 10.6151
R2506 B.n538 B.n537 10.6151
R2507 B.n537 B.n534 10.6151
R2508 B.n534 B.n533 10.6151
R2509 B.n533 B.n530 10.6151
R2510 B.n530 B.n529 10.6151
R2511 B.n529 B.n526 10.6151
R2512 B.n526 B.n525 10.6151
R2513 B.n525 B.n453 10.6151
R2514 B.n781 B.n453 10.6151
R2515 B.n787 B.n449 10.6151
R2516 B.n788 B.n787 10.6151
R2517 B.n789 B.n788 10.6151
R2518 B.n789 B.n441 10.6151
R2519 B.n799 B.n441 10.6151
R2520 B.n800 B.n799 10.6151
R2521 B.n801 B.n800 10.6151
R2522 B.n801 B.n433 10.6151
R2523 B.n811 B.n433 10.6151
R2524 B.n812 B.n811 10.6151
R2525 B.n813 B.n812 10.6151
R2526 B.n813 B.n425 10.6151
R2527 B.n823 B.n425 10.6151
R2528 B.n824 B.n823 10.6151
R2529 B.n825 B.n824 10.6151
R2530 B.n825 B.n417 10.6151
R2531 B.n835 B.n417 10.6151
R2532 B.n836 B.n835 10.6151
R2533 B.n837 B.n836 10.6151
R2534 B.n837 B.n409 10.6151
R2535 B.n847 B.n409 10.6151
R2536 B.n848 B.n847 10.6151
R2537 B.n849 B.n848 10.6151
R2538 B.n849 B.n401 10.6151
R2539 B.n859 B.n401 10.6151
R2540 B.n860 B.n859 10.6151
R2541 B.n861 B.n860 10.6151
R2542 B.n861 B.n393 10.6151
R2543 B.n872 B.n393 10.6151
R2544 B.n873 B.n872 10.6151
R2545 B.n874 B.n873 10.6151
R2546 B.n874 B.n0 10.6151
R2547 B.n986 B.n1 10.6151
R2548 B.n986 B.n985 10.6151
R2549 B.n985 B.n984 10.6151
R2550 B.n984 B.n10 10.6151
R2551 B.n978 B.n10 10.6151
R2552 B.n978 B.n977 10.6151
R2553 B.n977 B.n976 10.6151
R2554 B.n976 B.n17 10.6151
R2555 B.n970 B.n17 10.6151
R2556 B.n970 B.n969 10.6151
R2557 B.n969 B.n968 10.6151
R2558 B.n968 B.n24 10.6151
R2559 B.n962 B.n24 10.6151
R2560 B.n962 B.n961 10.6151
R2561 B.n961 B.n960 10.6151
R2562 B.n960 B.n31 10.6151
R2563 B.n954 B.n31 10.6151
R2564 B.n954 B.n953 10.6151
R2565 B.n953 B.n952 10.6151
R2566 B.n952 B.n38 10.6151
R2567 B.n946 B.n38 10.6151
R2568 B.n946 B.n945 10.6151
R2569 B.n945 B.n944 10.6151
R2570 B.n944 B.n45 10.6151
R2571 B.n938 B.n45 10.6151
R2572 B.n938 B.n937 10.6151
R2573 B.n937 B.n936 10.6151
R2574 B.n936 B.n52 10.6151
R2575 B.n930 B.n52 10.6151
R2576 B.n930 B.n929 10.6151
R2577 B.n929 B.n928 10.6151
R2578 B.n928 B.n59 10.6151
R2579 B.n254 B.n132 6.5566
R2580 B.n271 B.n270 6.5566
R2581 B.n658 B.n657 6.5566
R2582 B.n641 B.n523 6.5566
R2583 B.n857 B.t0 6.08431
R2584 B.n974 B.t1 6.08431
R2585 B.n251 B.n132 4.05904
R2586 B.n272 B.n271 4.05904
R2587 B.n659 B.n658 4.05904
R2588 B.n638 B.n523 4.05904
R2589 B.n992 B.n0 2.81026
R2590 B.n992 B.n1 2.81026
R2591 VP.n0 VP.t1 200.776
R2592 VP.n0 VP.t0 147.98
R2593 VP VP.n0 0.621237
R2594 VDD1.n96 VDD1.n0 289.615
R2595 VDD1.n197 VDD1.n101 289.615
R2596 VDD1.n97 VDD1.n96 185
R2597 VDD1.n95 VDD1.n94 185
R2598 VDD1.n4 VDD1.n3 185
R2599 VDD1.n89 VDD1.n88 185
R2600 VDD1.n87 VDD1.n86 185
R2601 VDD1.n8 VDD1.n7 185
R2602 VDD1.n81 VDD1.n80 185
R2603 VDD1.n79 VDD1.n10 185
R2604 VDD1.n78 VDD1.n77 185
R2605 VDD1.n13 VDD1.n11 185
R2606 VDD1.n72 VDD1.n71 185
R2607 VDD1.n70 VDD1.n69 185
R2608 VDD1.n17 VDD1.n16 185
R2609 VDD1.n64 VDD1.n63 185
R2610 VDD1.n62 VDD1.n61 185
R2611 VDD1.n21 VDD1.n20 185
R2612 VDD1.n56 VDD1.n55 185
R2613 VDD1.n54 VDD1.n53 185
R2614 VDD1.n25 VDD1.n24 185
R2615 VDD1.n48 VDD1.n47 185
R2616 VDD1.n46 VDD1.n45 185
R2617 VDD1.n29 VDD1.n28 185
R2618 VDD1.n40 VDD1.n39 185
R2619 VDD1.n38 VDD1.n37 185
R2620 VDD1.n33 VDD1.n32 185
R2621 VDD1.n133 VDD1.n132 185
R2622 VDD1.n138 VDD1.n137 185
R2623 VDD1.n140 VDD1.n139 185
R2624 VDD1.n129 VDD1.n128 185
R2625 VDD1.n146 VDD1.n145 185
R2626 VDD1.n148 VDD1.n147 185
R2627 VDD1.n125 VDD1.n124 185
R2628 VDD1.n154 VDD1.n153 185
R2629 VDD1.n156 VDD1.n155 185
R2630 VDD1.n121 VDD1.n120 185
R2631 VDD1.n162 VDD1.n161 185
R2632 VDD1.n164 VDD1.n163 185
R2633 VDD1.n117 VDD1.n116 185
R2634 VDD1.n170 VDD1.n169 185
R2635 VDD1.n172 VDD1.n171 185
R2636 VDD1.n113 VDD1.n112 185
R2637 VDD1.n179 VDD1.n178 185
R2638 VDD1.n180 VDD1.n111 185
R2639 VDD1.n182 VDD1.n181 185
R2640 VDD1.n109 VDD1.n108 185
R2641 VDD1.n188 VDD1.n187 185
R2642 VDD1.n190 VDD1.n189 185
R2643 VDD1.n105 VDD1.n104 185
R2644 VDD1.n196 VDD1.n195 185
R2645 VDD1.n198 VDD1.n197 185
R2646 VDD1.n34 VDD1.t0 147.659
R2647 VDD1.n134 VDD1.t1 147.659
R2648 VDD1.n96 VDD1.n95 104.615
R2649 VDD1.n95 VDD1.n3 104.615
R2650 VDD1.n88 VDD1.n3 104.615
R2651 VDD1.n88 VDD1.n87 104.615
R2652 VDD1.n87 VDD1.n7 104.615
R2653 VDD1.n80 VDD1.n7 104.615
R2654 VDD1.n80 VDD1.n79 104.615
R2655 VDD1.n79 VDD1.n78 104.615
R2656 VDD1.n78 VDD1.n11 104.615
R2657 VDD1.n71 VDD1.n11 104.615
R2658 VDD1.n71 VDD1.n70 104.615
R2659 VDD1.n70 VDD1.n16 104.615
R2660 VDD1.n63 VDD1.n16 104.615
R2661 VDD1.n63 VDD1.n62 104.615
R2662 VDD1.n62 VDD1.n20 104.615
R2663 VDD1.n55 VDD1.n20 104.615
R2664 VDD1.n55 VDD1.n54 104.615
R2665 VDD1.n54 VDD1.n24 104.615
R2666 VDD1.n47 VDD1.n24 104.615
R2667 VDD1.n47 VDD1.n46 104.615
R2668 VDD1.n46 VDD1.n28 104.615
R2669 VDD1.n39 VDD1.n28 104.615
R2670 VDD1.n39 VDD1.n38 104.615
R2671 VDD1.n38 VDD1.n32 104.615
R2672 VDD1.n138 VDD1.n132 104.615
R2673 VDD1.n139 VDD1.n138 104.615
R2674 VDD1.n139 VDD1.n128 104.615
R2675 VDD1.n146 VDD1.n128 104.615
R2676 VDD1.n147 VDD1.n146 104.615
R2677 VDD1.n147 VDD1.n124 104.615
R2678 VDD1.n154 VDD1.n124 104.615
R2679 VDD1.n155 VDD1.n154 104.615
R2680 VDD1.n155 VDD1.n120 104.615
R2681 VDD1.n162 VDD1.n120 104.615
R2682 VDD1.n163 VDD1.n162 104.615
R2683 VDD1.n163 VDD1.n116 104.615
R2684 VDD1.n170 VDD1.n116 104.615
R2685 VDD1.n171 VDD1.n170 104.615
R2686 VDD1.n171 VDD1.n112 104.615
R2687 VDD1.n179 VDD1.n112 104.615
R2688 VDD1.n180 VDD1.n179 104.615
R2689 VDD1.n181 VDD1.n180 104.615
R2690 VDD1.n181 VDD1.n108 104.615
R2691 VDD1.n188 VDD1.n108 104.615
R2692 VDD1.n189 VDD1.n188 104.615
R2693 VDD1.n189 VDD1.n104 104.615
R2694 VDD1.n196 VDD1.n104 104.615
R2695 VDD1.n197 VDD1.n196 104.615
R2696 VDD1 VDD1.n201 96.7553
R2697 VDD1.t0 VDD1.n32 52.3082
R2698 VDD1.t1 VDD1.n132 52.3082
R2699 VDD1 VDD1.n100 49.6379
R2700 VDD1.n34 VDD1.n33 15.6677
R2701 VDD1.n134 VDD1.n133 15.6677
R2702 VDD1.n81 VDD1.n10 13.1884
R2703 VDD1.n182 VDD1.n111 13.1884
R2704 VDD1.n82 VDD1.n8 12.8005
R2705 VDD1.n77 VDD1.n12 12.8005
R2706 VDD1.n37 VDD1.n36 12.8005
R2707 VDD1.n137 VDD1.n136 12.8005
R2708 VDD1.n178 VDD1.n177 12.8005
R2709 VDD1.n183 VDD1.n109 12.8005
R2710 VDD1.n86 VDD1.n85 12.0247
R2711 VDD1.n76 VDD1.n13 12.0247
R2712 VDD1.n40 VDD1.n31 12.0247
R2713 VDD1.n140 VDD1.n131 12.0247
R2714 VDD1.n176 VDD1.n113 12.0247
R2715 VDD1.n187 VDD1.n186 12.0247
R2716 VDD1.n89 VDD1.n6 11.249
R2717 VDD1.n73 VDD1.n72 11.249
R2718 VDD1.n41 VDD1.n29 11.249
R2719 VDD1.n141 VDD1.n129 11.249
R2720 VDD1.n173 VDD1.n172 11.249
R2721 VDD1.n190 VDD1.n107 11.249
R2722 VDD1.n90 VDD1.n4 10.4732
R2723 VDD1.n69 VDD1.n15 10.4732
R2724 VDD1.n45 VDD1.n44 10.4732
R2725 VDD1.n145 VDD1.n144 10.4732
R2726 VDD1.n169 VDD1.n115 10.4732
R2727 VDD1.n191 VDD1.n105 10.4732
R2728 VDD1.n94 VDD1.n93 9.69747
R2729 VDD1.n68 VDD1.n17 9.69747
R2730 VDD1.n48 VDD1.n27 9.69747
R2731 VDD1.n148 VDD1.n127 9.69747
R2732 VDD1.n168 VDD1.n117 9.69747
R2733 VDD1.n195 VDD1.n194 9.69747
R2734 VDD1.n100 VDD1.n99 9.45567
R2735 VDD1.n201 VDD1.n200 9.45567
R2736 VDD1.n60 VDD1.n59 9.3005
R2737 VDD1.n19 VDD1.n18 9.3005
R2738 VDD1.n66 VDD1.n65 9.3005
R2739 VDD1.n68 VDD1.n67 9.3005
R2740 VDD1.n15 VDD1.n14 9.3005
R2741 VDD1.n74 VDD1.n73 9.3005
R2742 VDD1.n76 VDD1.n75 9.3005
R2743 VDD1.n12 VDD1.n9 9.3005
R2744 VDD1.n99 VDD1.n98 9.3005
R2745 VDD1.n2 VDD1.n1 9.3005
R2746 VDD1.n93 VDD1.n92 9.3005
R2747 VDD1.n91 VDD1.n90 9.3005
R2748 VDD1.n6 VDD1.n5 9.3005
R2749 VDD1.n85 VDD1.n84 9.3005
R2750 VDD1.n83 VDD1.n82 9.3005
R2751 VDD1.n58 VDD1.n57 9.3005
R2752 VDD1.n23 VDD1.n22 9.3005
R2753 VDD1.n52 VDD1.n51 9.3005
R2754 VDD1.n50 VDD1.n49 9.3005
R2755 VDD1.n27 VDD1.n26 9.3005
R2756 VDD1.n44 VDD1.n43 9.3005
R2757 VDD1.n42 VDD1.n41 9.3005
R2758 VDD1.n31 VDD1.n30 9.3005
R2759 VDD1.n36 VDD1.n35 9.3005
R2760 VDD1.n200 VDD1.n199 9.3005
R2761 VDD1.n103 VDD1.n102 9.3005
R2762 VDD1.n194 VDD1.n193 9.3005
R2763 VDD1.n192 VDD1.n191 9.3005
R2764 VDD1.n107 VDD1.n106 9.3005
R2765 VDD1.n186 VDD1.n185 9.3005
R2766 VDD1.n184 VDD1.n183 9.3005
R2767 VDD1.n123 VDD1.n122 9.3005
R2768 VDD1.n152 VDD1.n151 9.3005
R2769 VDD1.n150 VDD1.n149 9.3005
R2770 VDD1.n127 VDD1.n126 9.3005
R2771 VDD1.n144 VDD1.n143 9.3005
R2772 VDD1.n142 VDD1.n141 9.3005
R2773 VDD1.n131 VDD1.n130 9.3005
R2774 VDD1.n136 VDD1.n135 9.3005
R2775 VDD1.n158 VDD1.n157 9.3005
R2776 VDD1.n160 VDD1.n159 9.3005
R2777 VDD1.n119 VDD1.n118 9.3005
R2778 VDD1.n166 VDD1.n165 9.3005
R2779 VDD1.n168 VDD1.n167 9.3005
R2780 VDD1.n115 VDD1.n114 9.3005
R2781 VDD1.n174 VDD1.n173 9.3005
R2782 VDD1.n176 VDD1.n175 9.3005
R2783 VDD1.n177 VDD1.n110 9.3005
R2784 VDD1.n97 VDD1.n2 8.92171
R2785 VDD1.n65 VDD1.n64 8.92171
R2786 VDD1.n49 VDD1.n25 8.92171
R2787 VDD1.n149 VDD1.n125 8.92171
R2788 VDD1.n165 VDD1.n164 8.92171
R2789 VDD1.n198 VDD1.n103 8.92171
R2790 VDD1.n98 VDD1.n0 8.14595
R2791 VDD1.n61 VDD1.n19 8.14595
R2792 VDD1.n53 VDD1.n52 8.14595
R2793 VDD1.n153 VDD1.n152 8.14595
R2794 VDD1.n161 VDD1.n119 8.14595
R2795 VDD1.n199 VDD1.n101 8.14595
R2796 VDD1.n60 VDD1.n21 7.3702
R2797 VDD1.n56 VDD1.n23 7.3702
R2798 VDD1.n156 VDD1.n123 7.3702
R2799 VDD1.n160 VDD1.n121 7.3702
R2800 VDD1.n57 VDD1.n21 6.59444
R2801 VDD1.n57 VDD1.n56 6.59444
R2802 VDD1.n157 VDD1.n156 6.59444
R2803 VDD1.n157 VDD1.n121 6.59444
R2804 VDD1.n100 VDD1.n0 5.81868
R2805 VDD1.n61 VDD1.n60 5.81868
R2806 VDD1.n53 VDD1.n23 5.81868
R2807 VDD1.n153 VDD1.n123 5.81868
R2808 VDD1.n161 VDD1.n160 5.81868
R2809 VDD1.n201 VDD1.n101 5.81868
R2810 VDD1.n98 VDD1.n97 5.04292
R2811 VDD1.n64 VDD1.n19 5.04292
R2812 VDD1.n52 VDD1.n25 5.04292
R2813 VDD1.n152 VDD1.n125 5.04292
R2814 VDD1.n164 VDD1.n119 5.04292
R2815 VDD1.n199 VDD1.n198 5.04292
R2816 VDD1.n35 VDD1.n34 4.38563
R2817 VDD1.n135 VDD1.n134 4.38563
R2818 VDD1.n94 VDD1.n2 4.26717
R2819 VDD1.n65 VDD1.n17 4.26717
R2820 VDD1.n49 VDD1.n48 4.26717
R2821 VDD1.n149 VDD1.n148 4.26717
R2822 VDD1.n165 VDD1.n117 4.26717
R2823 VDD1.n195 VDD1.n103 4.26717
R2824 VDD1.n93 VDD1.n4 3.49141
R2825 VDD1.n69 VDD1.n68 3.49141
R2826 VDD1.n45 VDD1.n27 3.49141
R2827 VDD1.n145 VDD1.n127 3.49141
R2828 VDD1.n169 VDD1.n168 3.49141
R2829 VDD1.n194 VDD1.n105 3.49141
R2830 VDD1.n90 VDD1.n89 2.71565
R2831 VDD1.n72 VDD1.n15 2.71565
R2832 VDD1.n44 VDD1.n29 2.71565
R2833 VDD1.n144 VDD1.n129 2.71565
R2834 VDD1.n172 VDD1.n115 2.71565
R2835 VDD1.n191 VDD1.n190 2.71565
R2836 VDD1.n86 VDD1.n6 1.93989
R2837 VDD1.n73 VDD1.n13 1.93989
R2838 VDD1.n41 VDD1.n40 1.93989
R2839 VDD1.n141 VDD1.n140 1.93989
R2840 VDD1.n173 VDD1.n113 1.93989
R2841 VDD1.n187 VDD1.n107 1.93989
R2842 VDD1.n85 VDD1.n8 1.16414
R2843 VDD1.n77 VDD1.n76 1.16414
R2844 VDD1.n37 VDD1.n31 1.16414
R2845 VDD1.n137 VDD1.n131 1.16414
R2846 VDD1.n178 VDD1.n176 1.16414
R2847 VDD1.n186 VDD1.n109 1.16414
R2848 VDD1.n82 VDD1.n81 0.388379
R2849 VDD1.n12 VDD1.n10 0.388379
R2850 VDD1.n36 VDD1.n33 0.388379
R2851 VDD1.n136 VDD1.n133 0.388379
R2852 VDD1.n177 VDD1.n111 0.388379
R2853 VDD1.n183 VDD1.n182 0.388379
R2854 VDD1.n99 VDD1.n1 0.155672
R2855 VDD1.n92 VDD1.n1 0.155672
R2856 VDD1.n92 VDD1.n91 0.155672
R2857 VDD1.n91 VDD1.n5 0.155672
R2858 VDD1.n84 VDD1.n5 0.155672
R2859 VDD1.n84 VDD1.n83 0.155672
R2860 VDD1.n83 VDD1.n9 0.155672
R2861 VDD1.n75 VDD1.n9 0.155672
R2862 VDD1.n75 VDD1.n74 0.155672
R2863 VDD1.n74 VDD1.n14 0.155672
R2864 VDD1.n67 VDD1.n14 0.155672
R2865 VDD1.n67 VDD1.n66 0.155672
R2866 VDD1.n66 VDD1.n18 0.155672
R2867 VDD1.n59 VDD1.n18 0.155672
R2868 VDD1.n59 VDD1.n58 0.155672
R2869 VDD1.n58 VDD1.n22 0.155672
R2870 VDD1.n51 VDD1.n22 0.155672
R2871 VDD1.n51 VDD1.n50 0.155672
R2872 VDD1.n50 VDD1.n26 0.155672
R2873 VDD1.n43 VDD1.n26 0.155672
R2874 VDD1.n43 VDD1.n42 0.155672
R2875 VDD1.n42 VDD1.n30 0.155672
R2876 VDD1.n35 VDD1.n30 0.155672
R2877 VDD1.n135 VDD1.n130 0.155672
R2878 VDD1.n142 VDD1.n130 0.155672
R2879 VDD1.n143 VDD1.n142 0.155672
R2880 VDD1.n143 VDD1.n126 0.155672
R2881 VDD1.n150 VDD1.n126 0.155672
R2882 VDD1.n151 VDD1.n150 0.155672
R2883 VDD1.n151 VDD1.n122 0.155672
R2884 VDD1.n158 VDD1.n122 0.155672
R2885 VDD1.n159 VDD1.n158 0.155672
R2886 VDD1.n159 VDD1.n118 0.155672
R2887 VDD1.n166 VDD1.n118 0.155672
R2888 VDD1.n167 VDD1.n166 0.155672
R2889 VDD1.n167 VDD1.n114 0.155672
R2890 VDD1.n174 VDD1.n114 0.155672
R2891 VDD1.n175 VDD1.n174 0.155672
R2892 VDD1.n175 VDD1.n110 0.155672
R2893 VDD1.n184 VDD1.n110 0.155672
R2894 VDD1.n185 VDD1.n184 0.155672
R2895 VDD1.n185 VDD1.n106 0.155672
R2896 VDD1.n192 VDD1.n106 0.155672
R2897 VDD1.n193 VDD1.n192 0.155672
R2898 VDD1.n193 VDD1.n102 0.155672
R2899 VDD1.n200 VDD1.n102 0.155672
C0 VN VDD2 4.3157f
C1 VTAIL VDD2 6.94237f
C2 VN VP 7.215569f
C3 VN VDD1 0.148715f
C4 VTAIL VP 3.77564f
C5 VTAIL VDD1 6.88303f
C6 VDD2 VP 0.386611f
C7 VDD1 VDD2 0.819859f
C8 VDD1 VP 4.5518f
C9 VN VTAIL 3.76035f
C10 VDD2 B 6.010192f
C11 VDD1 B 9.4691f
C12 VTAIL B 10.543526f
C13 VN B 13.42495f
C14 VP B 8.416918f
C15 VDD1.n0 B 0.028482f
C16 VDD1.n1 B 0.020361f
C17 VDD1.n2 B 0.010941f
C18 VDD1.n3 B 0.025861f
C19 VDD1.n4 B 0.011585f
C20 VDD1.n5 B 0.020361f
C21 VDD1.n6 B 0.010941f
C22 VDD1.n7 B 0.025861f
C23 VDD1.n8 B 0.011585f
C24 VDD1.n9 B 0.020361f
C25 VDD1.n10 B 0.011263f
C26 VDD1.n11 B 0.025861f
C27 VDD1.n12 B 0.010941f
C28 VDD1.n13 B 0.011585f
C29 VDD1.n14 B 0.020361f
C30 VDD1.n15 B 0.010941f
C31 VDD1.n16 B 0.025861f
C32 VDD1.n17 B 0.011585f
C33 VDD1.n18 B 0.020361f
C34 VDD1.n19 B 0.010941f
C35 VDD1.n20 B 0.025861f
C36 VDD1.n21 B 0.011585f
C37 VDD1.n22 B 0.020361f
C38 VDD1.n23 B 0.010941f
C39 VDD1.n24 B 0.025861f
C40 VDD1.n25 B 0.011585f
C41 VDD1.n26 B 0.020361f
C42 VDD1.n27 B 0.010941f
C43 VDD1.n28 B 0.025861f
C44 VDD1.n29 B 0.011585f
C45 VDD1.n30 B 0.020361f
C46 VDD1.n31 B 0.010941f
C47 VDD1.n32 B 0.019396f
C48 VDD1.n33 B 0.015277f
C49 VDD1.t0 B 0.042867f
C50 VDD1.n34 B 0.149288f
C51 VDD1.n35 B 1.62612f
C52 VDD1.n36 B 0.010941f
C53 VDD1.n37 B 0.011585f
C54 VDD1.n38 B 0.025861f
C55 VDD1.n39 B 0.025861f
C56 VDD1.n40 B 0.011585f
C57 VDD1.n41 B 0.010941f
C58 VDD1.n42 B 0.020361f
C59 VDD1.n43 B 0.020361f
C60 VDD1.n44 B 0.010941f
C61 VDD1.n45 B 0.011585f
C62 VDD1.n46 B 0.025861f
C63 VDD1.n47 B 0.025861f
C64 VDD1.n48 B 0.011585f
C65 VDD1.n49 B 0.010941f
C66 VDD1.n50 B 0.020361f
C67 VDD1.n51 B 0.020361f
C68 VDD1.n52 B 0.010941f
C69 VDD1.n53 B 0.011585f
C70 VDD1.n54 B 0.025861f
C71 VDD1.n55 B 0.025861f
C72 VDD1.n56 B 0.011585f
C73 VDD1.n57 B 0.010941f
C74 VDD1.n58 B 0.020361f
C75 VDD1.n59 B 0.020361f
C76 VDD1.n60 B 0.010941f
C77 VDD1.n61 B 0.011585f
C78 VDD1.n62 B 0.025861f
C79 VDD1.n63 B 0.025861f
C80 VDD1.n64 B 0.011585f
C81 VDD1.n65 B 0.010941f
C82 VDD1.n66 B 0.020361f
C83 VDD1.n67 B 0.020361f
C84 VDD1.n68 B 0.010941f
C85 VDD1.n69 B 0.011585f
C86 VDD1.n70 B 0.025861f
C87 VDD1.n71 B 0.025861f
C88 VDD1.n72 B 0.011585f
C89 VDD1.n73 B 0.010941f
C90 VDD1.n74 B 0.020361f
C91 VDD1.n75 B 0.020361f
C92 VDD1.n76 B 0.010941f
C93 VDD1.n77 B 0.011585f
C94 VDD1.n78 B 0.025861f
C95 VDD1.n79 B 0.025861f
C96 VDD1.n80 B 0.025861f
C97 VDD1.n81 B 0.011263f
C98 VDD1.n82 B 0.010941f
C99 VDD1.n83 B 0.020361f
C100 VDD1.n84 B 0.020361f
C101 VDD1.n85 B 0.010941f
C102 VDD1.n86 B 0.011585f
C103 VDD1.n87 B 0.025861f
C104 VDD1.n88 B 0.025861f
C105 VDD1.n89 B 0.011585f
C106 VDD1.n90 B 0.010941f
C107 VDD1.n91 B 0.020361f
C108 VDD1.n92 B 0.020361f
C109 VDD1.n93 B 0.010941f
C110 VDD1.n94 B 0.011585f
C111 VDD1.n95 B 0.025861f
C112 VDD1.n96 B 0.055741f
C113 VDD1.n97 B 0.011585f
C114 VDD1.n98 B 0.010941f
C115 VDD1.n99 B 0.046785f
C116 VDD1.n100 B 0.047216f
C117 VDD1.n101 B 0.028482f
C118 VDD1.n102 B 0.020361f
C119 VDD1.n103 B 0.010941f
C120 VDD1.n104 B 0.025861f
C121 VDD1.n105 B 0.011585f
C122 VDD1.n106 B 0.020361f
C123 VDD1.n107 B 0.010941f
C124 VDD1.n108 B 0.025861f
C125 VDD1.n109 B 0.011585f
C126 VDD1.n110 B 0.020361f
C127 VDD1.n111 B 0.011263f
C128 VDD1.n112 B 0.025861f
C129 VDD1.n113 B 0.011585f
C130 VDD1.n114 B 0.020361f
C131 VDD1.n115 B 0.010941f
C132 VDD1.n116 B 0.025861f
C133 VDD1.n117 B 0.011585f
C134 VDD1.n118 B 0.020361f
C135 VDD1.n119 B 0.010941f
C136 VDD1.n120 B 0.025861f
C137 VDD1.n121 B 0.011585f
C138 VDD1.n122 B 0.020361f
C139 VDD1.n123 B 0.010941f
C140 VDD1.n124 B 0.025861f
C141 VDD1.n125 B 0.011585f
C142 VDD1.n126 B 0.020361f
C143 VDD1.n127 B 0.010941f
C144 VDD1.n128 B 0.025861f
C145 VDD1.n129 B 0.011585f
C146 VDD1.n130 B 0.020361f
C147 VDD1.n131 B 0.010941f
C148 VDD1.n132 B 0.019396f
C149 VDD1.n133 B 0.015277f
C150 VDD1.t1 B 0.042867f
C151 VDD1.n134 B 0.149288f
C152 VDD1.n135 B 1.62612f
C153 VDD1.n136 B 0.010941f
C154 VDD1.n137 B 0.011585f
C155 VDD1.n138 B 0.025861f
C156 VDD1.n139 B 0.025861f
C157 VDD1.n140 B 0.011585f
C158 VDD1.n141 B 0.010941f
C159 VDD1.n142 B 0.020361f
C160 VDD1.n143 B 0.020361f
C161 VDD1.n144 B 0.010941f
C162 VDD1.n145 B 0.011585f
C163 VDD1.n146 B 0.025861f
C164 VDD1.n147 B 0.025861f
C165 VDD1.n148 B 0.011585f
C166 VDD1.n149 B 0.010941f
C167 VDD1.n150 B 0.020361f
C168 VDD1.n151 B 0.020361f
C169 VDD1.n152 B 0.010941f
C170 VDD1.n153 B 0.011585f
C171 VDD1.n154 B 0.025861f
C172 VDD1.n155 B 0.025861f
C173 VDD1.n156 B 0.011585f
C174 VDD1.n157 B 0.010941f
C175 VDD1.n158 B 0.020361f
C176 VDD1.n159 B 0.020361f
C177 VDD1.n160 B 0.010941f
C178 VDD1.n161 B 0.011585f
C179 VDD1.n162 B 0.025861f
C180 VDD1.n163 B 0.025861f
C181 VDD1.n164 B 0.011585f
C182 VDD1.n165 B 0.010941f
C183 VDD1.n166 B 0.020361f
C184 VDD1.n167 B 0.020361f
C185 VDD1.n168 B 0.010941f
C186 VDD1.n169 B 0.011585f
C187 VDD1.n170 B 0.025861f
C188 VDD1.n171 B 0.025861f
C189 VDD1.n172 B 0.011585f
C190 VDD1.n173 B 0.010941f
C191 VDD1.n174 B 0.020361f
C192 VDD1.n175 B 0.020361f
C193 VDD1.n176 B 0.010941f
C194 VDD1.n177 B 0.010941f
C195 VDD1.n178 B 0.011585f
C196 VDD1.n179 B 0.025861f
C197 VDD1.n180 B 0.025861f
C198 VDD1.n181 B 0.025861f
C199 VDD1.n182 B 0.011263f
C200 VDD1.n183 B 0.010941f
C201 VDD1.n184 B 0.020361f
C202 VDD1.n185 B 0.020361f
C203 VDD1.n186 B 0.010941f
C204 VDD1.n187 B 0.011585f
C205 VDD1.n188 B 0.025861f
C206 VDD1.n189 B 0.025861f
C207 VDD1.n190 B 0.011585f
C208 VDD1.n191 B 0.010941f
C209 VDD1.n192 B 0.020361f
C210 VDD1.n193 B 0.020361f
C211 VDD1.n194 B 0.010941f
C212 VDD1.n195 B 0.011585f
C213 VDD1.n196 B 0.025861f
C214 VDD1.n197 B 0.055741f
C215 VDD1.n198 B 0.011585f
C216 VDD1.n199 B 0.010941f
C217 VDD1.n200 B 0.046785f
C218 VDD1.n201 B 0.920243f
C219 VP.t1 B 5.65547f
C220 VP.t0 B 4.89312f
C221 VP.n0 B 4.95104f
C222 VDD2.n0 B 0.027921f
C223 VDD2.n1 B 0.01996f
C224 VDD2.n2 B 0.010726f
C225 VDD2.n3 B 0.025352f
C226 VDD2.n4 B 0.011357f
C227 VDD2.n5 B 0.01996f
C228 VDD2.n6 B 0.010726f
C229 VDD2.n7 B 0.025352f
C230 VDD2.n8 B 0.011357f
C231 VDD2.n9 B 0.01996f
C232 VDD2.n10 B 0.011041f
C233 VDD2.n11 B 0.025352f
C234 VDD2.n12 B 0.011357f
C235 VDD2.n13 B 0.01996f
C236 VDD2.n14 B 0.010726f
C237 VDD2.n15 B 0.025352f
C238 VDD2.n16 B 0.011357f
C239 VDD2.n17 B 0.01996f
C240 VDD2.n18 B 0.010726f
C241 VDD2.n19 B 0.025352f
C242 VDD2.n20 B 0.011357f
C243 VDD2.n21 B 0.01996f
C244 VDD2.n22 B 0.010726f
C245 VDD2.n23 B 0.025352f
C246 VDD2.n24 B 0.011357f
C247 VDD2.n25 B 0.01996f
C248 VDD2.n26 B 0.010726f
C249 VDD2.n27 B 0.025352f
C250 VDD2.n28 B 0.011357f
C251 VDD2.n29 B 0.01996f
C252 VDD2.n30 B 0.010726f
C253 VDD2.n31 B 0.019014f
C254 VDD2.n32 B 0.014976f
C255 VDD2.t1 B 0.042024f
C256 VDD2.n33 B 0.146351f
C257 VDD2.n34 B 1.59413f
C258 VDD2.n35 B 0.010726f
C259 VDD2.n36 B 0.011357f
C260 VDD2.n37 B 0.025352f
C261 VDD2.n38 B 0.025352f
C262 VDD2.n39 B 0.011357f
C263 VDD2.n40 B 0.010726f
C264 VDD2.n41 B 0.01996f
C265 VDD2.n42 B 0.01996f
C266 VDD2.n43 B 0.010726f
C267 VDD2.n44 B 0.011357f
C268 VDD2.n45 B 0.025352f
C269 VDD2.n46 B 0.025352f
C270 VDD2.n47 B 0.011357f
C271 VDD2.n48 B 0.010726f
C272 VDD2.n49 B 0.01996f
C273 VDD2.n50 B 0.01996f
C274 VDD2.n51 B 0.010726f
C275 VDD2.n52 B 0.011357f
C276 VDD2.n53 B 0.025352f
C277 VDD2.n54 B 0.025352f
C278 VDD2.n55 B 0.011357f
C279 VDD2.n56 B 0.010726f
C280 VDD2.n57 B 0.01996f
C281 VDD2.n58 B 0.01996f
C282 VDD2.n59 B 0.010726f
C283 VDD2.n60 B 0.011357f
C284 VDD2.n61 B 0.025352f
C285 VDD2.n62 B 0.025352f
C286 VDD2.n63 B 0.011357f
C287 VDD2.n64 B 0.010726f
C288 VDD2.n65 B 0.01996f
C289 VDD2.n66 B 0.01996f
C290 VDD2.n67 B 0.010726f
C291 VDD2.n68 B 0.011357f
C292 VDD2.n69 B 0.025352f
C293 VDD2.n70 B 0.025352f
C294 VDD2.n71 B 0.011357f
C295 VDD2.n72 B 0.010726f
C296 VDD2.n73 B 0.01996f
C297 VDD2.n74 B 0.01996f
C298 VDD2.n75 B 0.010726f
C299 VDD2.n76 B 0.010726f
C300 VDD2.n77 B 0.011357f
C301 VDD2.n78 B 0.025352f
C302 VDD2.n79 B 0.025352f
C303 VDD2.n80 B 0.025352f
C304 VDD2.n81 B 0.011041f
C305 VDD2.n82 B 0.010726f
C306 VDD2.n83 B 0.01996f
C307 VDD2.n84 B 0.01996f
C308 VDD2.n85 B 0.010726f
C309 VDD2.n86 B 0.011357f
C310 VDD2.n87 B 0.025352f
C311 VDD2.n88 B 0.025352f
C312 VDD2.n89 B 0.011357f
C313 VDD2.n90 B 0.010726f
C314 VDD2.n91 B 0.01996f
C315 VDD2.n92 B 0.01996f
C316 VDD2.n93 B 0.010726f
C317 VDD2.n94 B 0.011357f
C318 VDD2.n95 B 0.025352f
C319 VDD2.n96 B 0.054645f
C320 VDD2.n97 B 0.011357f
C321 VDD2.n98 B 0.010726f
C322 VDD2.n99 B 0.045865f
C323 VDD2.n100 B 0.848843f
C324 VDD2.n101 B 0.027921f
C325 VDD2.n102 B 0.01996f
C326 VDD2.n103 B 0.010726f
C327 VDD2.n104 B 0.025352f
C328 VDD2.n105 B 0.011357f
C329 VDD2.n106 B 0.01996f
C330 VDD2.n107 B 0.010726f
C331 VDD2.n108 B 0.025352f
C332 VDD2.n109 B 0.011357f
C333 VDD2.n110 B 0.01996f
C334 VDD2.n111 B 0.011041f
C335 VDD2.n112 B 0.025352f
C336 VDD2.n113 B 0.010726f
C337 VDD2.n114 B 0.011357f
C338 VDD2.n115 B 0.01996f
C339 VDD2.n116 B 0.010726f
C340 VDD2.n117 B 0.025352f
C341 VDD2.n118 B 0.011357f
C342 VDD2.n119 B 0.01996f
C343 VDD2.n120 B 0.010726f
C344 VDD2.n121 B 0.025352f
C345 VDD2.n122 B 0.011357f
C346 VDD2.n123 B 0.01996f
C347 VDD2.n124 B 0.010726f
C348 VDD2.n125 B 0.025352f
C349 VDD2.n126 B 0.011357f
C350 VDD2.n127 B 0.01996f
C351 VDD2.n128 B 0.010726f
C352 VDD2.n129 B 0.025352f
C353 VDD2.n130 B 0.011357f
C354 VDD2.n131 B 0.01996f
C355 VDD2.n132 B 0.010726f
C356 VDD2.n133 B 0.019014f
C357 VDD2.n134 B 0.014976f
C358 VDD2.t0 B 0.042024f
C359 VDD2.n135 B 0.146351f
C360 VDD2.n136 B 1.59413f
C361 VDD2.n137 B 0.010726f
C362 VDD2.n138 B 0.011357f
C363 VDD2.n139 B 0.025352f
C364 VDD2.n140 B 0.025352f
C365 VDD2.n141 B 0.011357f
C366 VDD2.n142 B 0.010726f
C367 VDD2.n143 B 0.01996f
C368 VDD2.n144 B 0.01996f
C369 VDD2.n145 B 0.010726f
C370 VDD2.n146 B 0.011357f
C371 VDD2.n147 B 0.025352f
C372 VDD2.n148 B 0.025352f
C373 VDD2.n149 B 0.011357f
C374 VDD2.n150 B 0.010726f
C375 VDD2.n151 B 0.01996f
C376 VDD2.n152 B 0.01996f
C377 VDD2.n153 B 0.010726f
C378 VDD2.n154 B 0.011357f
C379 VDD2.n155 B 0.025352f
C380 VDD2.n156 B 0.025352f
C381 VDD2.n157 B 0.011357f
C382 VDD2.n158 B 0.010726f
C383 VDD2.n159 B 0.01996f
C384 VDD2.n160 B 0.01996f
C385 VDD2.n161 B 0.010726f
C386 VDD2.n162 B 0.011357f
C387 VDD2.n163 B 0.025352f
C388 VDD2.n164 B 0.025352f
C389 VDD2.n165 B 0.011357f
C390 VDD2.n166 B 0.010726f
C391 VDD2.n167 B 0.01996f
C392 VDD2.n168 B 0.01996f
C393 VDD2.n169 B 0.010726f
C394 VDD2.n170 B 0.011357f
C395 VDD2.n171 B 0.025352f
C396 VDD2.n172 B 0.025352f
C397 VDD2.n173 B 0.011357f
C398 VDD2.n174 B 0.010726f
C399 VDD2.n175 B 0.01996f
C400 VDD2.n176 B 0.01996f
C401 VDD2.n177 B 0.010726f
C402 VDD2.n178 B 0.011357f
C403 VDD2.n179 B 0.025352f
C404 VDD2.n180 B 0.025352f
C405 VDD2.n181 B 0.025352f
C406 VDD2.n182 B 0.011041f
C407 VDD2.n183 B 0.010726f
C408 VDD2.n184 B 0.01996f
C409 VDD2.n185 B 0.01996f
C410 VDD2.n186 B 0.010726f
C411 VDD2.n187 B 0.011357f
C412 VDD2.n188 B 0.025352f
C413 VDD2.n189 B 0.025352f
C414 VDD2.n190 B 0.011357f
C415 VDD2.n191 B 0.010726f
C416 VDD2.n192 B 0.01996f
C417 VDD2.n193 B 0.01996f
C418 VDD2.n194 B 0.010726f
C419 VDD2.n195 B 0.011357f
C420 VDD2.n196 B 0.025352f
C421 VDD2.n197 B 0.054645f
C422 VDD2.n198 B 0.011357f
C423 VDD2.n199 B 0.010726f
C424 VDD2.n200 B 0.045865f
C425 VDD2.n201 B 0.044327f
C426 VDD2.n202 B 3.13405f
C427 VTAIL.n0 B 0.028058f
C428 VTAIL.n1 B 0.020058f
C429 VTAIL.n2 B 0.010778f
C430 VTAIL.n3 B 0.025476f
C431 VTAIL.n4 B 0.011412f
C432 VTAIL.n5 B 0.020058f
C433 VTAIL.n6 B 0.010778f
C434 VTAIL.n7 B 0.025476f
C435 VTAIL.n8 B 0.011412f
C436 VTAIL.n9 B 0.020058f
C437 VTAIL.n10 B 0.011095f
C438 VTAIL.n11 B 0.025476f
C439 VTAIL.n12 B 0.011412f
C440 VTAIL.n13 B 0.020058f
C441 VTAIL.n14 B 0.010778f
C442 VTAIL.n15 B 0.025476f
C443 VTAIL.n16 B 0.011412f
C444 VTAIL.n17 B 0.020058f
C445 VTAIL.n18 B 0.010778f
C446 VTAIL.n19 B 0.025476f
C447 VTAIL.n20 B 0.011412f
C448 VTAIL.n21 B 0.020058f
C449 VTAIL.n22 B 0.010778f
C450 VTAIL.n23 B 0.025476f
C451 VTAIL.n24 B 0.011412f
C452 VTAIL.n25 B 0.020058f
C453 VTAIL.n26 B 0.010778f
C454 VTAIL.n27 B 0.025476f
C455 VTAIL.n28 B 0.011412f
C456 VTAIL.n29 B 0.020058f
C457 VTAIL.n30 B 0.010778f
C458 VTAIL.n31 B 0.019107f
C459 VTAIL.n32 B 0.015049f
C460 VTAIL.t0 B 0.042229f
C461 VTAIL.n33 B 0.147065f
C462 VTAIL.n34 B 1.6019f
C463 VTAIL.n35 B 0.010778f
C464 VTAIL.n36 B 0.011412f
C465 VTAIL.n37 B 0.025476f
C466 VTAIL.n38 B 0.025476f
C467 VTAIL.n39 B 0.011412f
C468 VTAIL.n40 B 0.010778f
C469 VTAIL.n41 B 0.020058f
C470 VTAIL.n42 B 0.020058f
C471 VTAIL.n43 B 0.010778f
C472 VTAIL.n44 B 0.011412f
C473 VTAIL.n45 B 0.025476f
C474 VTAIL.n46 B 0.025476f
C475 VTAIL.n47 B 0.011412f
C476 VTAIL.n48 B 0.010778f
C477 VTAIL.n49 B 0.020058f
C478 VTAIL.n50 B 0.020058f
C479 VTAIL.n51 B 0.010778f
C480 VTAIL.n52 B 0.011412f
C481 VTAIL.n53 B 0.025476f
C482 VTAIL.n54 B 0.025476f
C483 VTAIL.n55 B 0.011412f
C484 VTAIL.n56 B 0.010778f
C485 VTAIL.n57 B 0.020058f
C486 VTAIL.n58 B 0.020058f
C487 VTAIL.n59 B 0.010778f
C488 VTAIL.n60 B 0.011412f
C489 VTAIL.n61 B 0.025476f
C490 VTAIL.n62 B 0.025476f
C491 VTAIL.n63 B 0.011412f
C492 VTAIL.n64 B 0.010778f
C493 VTAIL.n65 B 0.020058f
C494 VTAIL.n66 B 0.020058f
C495 VTAIL.n67 B 0.010778f
C496 VTAIL.n68 B 0.011412f
C497 VTAIL.n69 B 0.025476f
C498 VTAIL.n70 B 0.025476f
C499 VTAIL.n71 B 0.011412f
C500 VTAIL.n72 B 0.010778f
C501 VTAIL.n73 B 0.020058f
C502 VTAIL.n74 B 0.020058f
C503 VTAIL.n75 B 0.010778f
C504 VTAIL.n76 B 0.010778f
C505 VTAIL.n77 B 0.011412f
C506 VTAIL.n78 B 0.025476f
C507 VTAIL.n79 B 0.025476f
C508 VTAIL.n80 B 0.025476f
C509 VTAIL.n81 B 0.011095f
C510 VTAIL.n82 B 0.010778f
C511 VTAIL.n83 B 0.020058f
C512 VTAIL.n84 B 0.020058f
C513 VTAIL.n85 B 0.010778f
C514 VTAIL.n86 B 0.011412f
C515 VTAIL.n87 B 0.025476f
C516 VTAIL.n88 B 0.025476f
C517 VTAIL.n89 B 0.011412f
C518 VTAIL.n90 B 0.010778f
C519 VTAIL.n91 B 0.020058f
C520 VTAIL.n92 B 0.020058f
C521 VTAIL.n93 B 0.010778f
C522 VTAIL.n94 B 0.011412f
C523 VTAIL.n95 B 0.025476f
C524 VTAIL.n96 B 0.054911f
C525 VTAIL.n97 B 0.011412f
C526 VTAIL.n98 B 0.010778f
C527 VTAIL.n99 B 0.046089f
C528 VTAIL.n100 B 0.030692f
C529 VTAIL.n101 B 1.86829f
C530 VTAIL.n102 B 0.028058f
C531 VTAIL.n103 B 0.020058f
C532 VTAIL.n104 B 0.010778f
C533 VTAIL.n105 B 0.025476f
C534 VTAIL.n106 B 0.011412f
C535 VTAIL.n107 B 0.020058f
C536 VTAIL.n108 B 0.010778f
C537 VTAIL.n109 B 0.025476f
C538 VTAIL.n110 B 0.011412f
C539 VTAIL.n111 B 0.020058f
C540 VTAIL.n112 B 0.011095f
C541 VTAIL.n113 B 0.025476f
C542 VTAIL.n114 B 0.010778f
C543 VTAIL.n115 B 0.011412f
C544 VTAIL.n116 B 0.020058f
C545 VTAIL.n117 B 0.010778f
C546 VTAIL.n118 B 0.025476f
C547 VTAIL.n119 B 0.011412f
C548 VTAIL.n120 B 0.020058f
C549 VTAIL.n121 B 0.010778f
C550 VTAIL.n122 B 0.025476f
C551 VTAIL.n123 B 0.011412f
C552 VTAIL.n124 B 0.020058f
C553 VTAIL.n125 B 0.010778f
C554 VTAIL.n126 B 0.025476f
C555 VTAIL.n127 B 0.011412f
C556 VTAIL.n128 B 0.020058f
C557 VTAIL.n129 B 0.010778f
C558 VTAIL.n130 B 0.025476f
C559 VTAIL.n131 B 0.011412f
C560 VTAIL.n132 B 0.020058f
C561 VTAIL.n133 B 0.010778f
C562 VTAIL.n134 B 0.019107f
C563 VTAIL.n135 B 0.015049f
C564 VTAIL.t2 B 0.042229f
C565 VTAIL.n136 B 0.147065f
C566 VTAIL.n137 B 1.6019f
C567 VTAIL.n138 B 0.010778f
C568 VTAIL.n139 B 0.011412f
C569 VTAIL.n140 B 0.025476f
C570 VTAIL.n141 B 0.025476f
C571 VTAIL.n142 B 0.011412f
C572 VTAIL.n143 B 0.010778f
C573 VTAIL.n144 B 0.020058f
C574 VTAIL.n145 B 0.020058f
C575 VTAIL.n146 B 0.010778f
C576 VTAIL.n147 B 0.011412f
C577 VTAIL.n148 B 0.025476f
C578 VTAIL.n149 B 0.025476f
C579 VTAIL.n150 B 0.011412f
C580 VTAIL.n151 B 0.010778f
C581 VTAIL.n152 B 0.020058f
C582 VTAIL.n153 B 0.020058f
C583 VTAIL.n154 B 0.010778f
C584 VTAIL.n155 B 0.011412f
C585 VTAIL.n156 B 0.025476f
C586 VTAIL.n157 B 0.025476f
C587 VTAIL.n158 B 0.011412f
C588 VTAIL.n159 B 0.010778f
C589 VTAIL.n160 B 0.020058f
C590 VTAIL.n161 B 0.020058f
C591 VTAIL.n162 B 0.010778f
C592 VTAIL.n163 B 0.011412f
C593 VTAIL.n164 B 0.025476f
C594 VTAIL.n165 B 0.025476f
C595 VTAIL.n166 B 0.011412f
C596 VTAIL.n167 B 0.010778f
C597 VTAIL.n168 B 0.020058f
C598 VTAIL.n169 B 0.020058f
C599 VTAIL.n170 B 0.010778f
C600 VTAIL.n171 B 0.011412f
C601 VTAIL.n172 B 0.025476f
C602 VTAIL.n173 B 0.025476f
C603 VTAIL.n174 B 0.011412f
C604 VTAIL.n175 B 0.010778f
C605 VTAIL.n176 B 0.020058f
C606 VTAIL.n177 B 0.020058f
C607 VTAIL.n178 B 0.010778f
C608 VTAIL.n179 B 0.011412f
C609 VTAIL.n180 B 0.025476f
C610 VTAIL.n181 B 0.025476f
C611 VTAIL.n182 B 0.025476f
C612 VTAIL.n183 B 0.011095f
C613 VTAIL.n184 B 0.010778f
C614 VTAIL.n185 B 0.020058f
C615 VTAIL.n186 B 0.020058f
C616 VTAIL.n187 B 0.010778f
C617 VTAIL.n188 B 0.011412f
C618 VTAIL.n189 B 0.025476f
C619 VTAIL.n190 B 0.025476f
C620 VTAIL.n191 B 0.011412f
C621 VTAIL.n192 B 0.010778f
C622 VTAIL.n193 B 0.020058f
C623 VTAIL.n194 B 0.020058f
C624 VTAIL.n195 B 0.010778f
C625 VTAIL.n196 B 0.011412f
C626 VTAIL.n197 B 0.025476f
C627 VTAIL.n198 B 0.054911f
C628 VTAIL.n199 B 0.011412f
C629 VTAIL.n200 B 0.010778f
C630 VTAIL.n201 B 0.046089f
C631 VTAIL.n202 B 0.030692f
C632 VTAIL.n203 B 1.92331f
C633 VTAIL.n204 B 0.028058f
C634 VTAIL.n205 B 0.020058f
C635 VTAIL.n206 B 0.010778f
C636 VTAIL.n207 B 0.025476f
C637 VTAIL.n208 B 0.011412f
C638 VTAIL.n209 B 0.020058f
C639 VTAIL.n210 B 0.010778f
C640 VTAIL.n211 B 0.025476f
C641 VTAIL.n212 B 0.011412f
C642 VTAIL.n213 B 0.020058f
C643 VTAIL.n214 B 0.011095f
C644 VTAIL.n215 B 0.025476f
C645 VTAIL.n216 B 0.010778f
C646 VTAIL.n217 B 0.011412f
C647 VTAIL.n218 B 0.020058f
C648 VTAIL.n219 B 0.010778f
C649 VTAIL.n220 B 0.025476f
C650 VTAIL.n221 B 0.011412f
C651 VTAIL.n222 B 0.020058f
C652 VTAIL.n223 B 0.010778f
C653 VTAIL.n224 B 0.025476f
C654 VTAIL.n225 B 0.011412f
C655 VTAIL.n226 B 0.020058f
C656 VTAIL.n227 B 0.010778f
C657 VTAIL.n228 B 0.025476f
C658 VTAIL.n229 B 0.011412f
C659 VTAIL.n230 B 0.020058f
C660 VTAIL.n231 B 0.010778f
C661 VTAIL.n232 B 0.025476f
C662 VTAIL.n233 B 0.011412f
C663 VTAIL.n234 B 0.020058f
C664 VTAIL.n235 B 0.010778f
C665 VTAIL.n236 B 0.019107f
C666 VTAIL.n237 B 0.015049f
C667 VTAIL.t1 B 0.042229f
C668 VTAIL.n238 B 0.147065f
C669 VTAIL.n239 B 1.6019f
C670 VTAIL.n240 B 0.010778f
C671 VTAIL.n241 B 0.011412f
C672 VTAIL.n242 B 0.025476f
C673 VTAIL.n243 B 0.025476f
C674 VTAIL.n244 B 0.011412f
C675 VTAIL.n245 B 0.010778f
C676 VTAIL.n246 B 0.020058f
C677 VTAIL.n247 B 0.020058f
C678 VTAIL.n248 B 0.010778f
C679 VTAIL.n249 B 0.011412f
C680 VTAIL.n250 B 0.025476f
C681 VTAIL.n251 B 0.025476f
C682 VTAIL.n252 B 0.011412f
C683 VTAIL.n253 B 0.010778f
C684 VTAIL.n254 B 0.020058f
C685 VTAIL.n255 B 0.020058f
C686 VTAIL.n256 B 0.010778f
C687 VTAIL.n257 B 0.011412f
C688 VTAIL.n258 B 0.025476f
C689 VTAIL.n259 B 0.025476f
C690 VTAIL.n260 B 0.011412f
C691 VTAIL.n261 B 0.010778f
C692 VTAIL.n262 B 0.020058f
C693 VTAIL.n263 B 0.020058f
C694 VTAIL.n264 B 0.010778f
C695 VTAIL.n265 B 0.011412f
C696 VTAIL.n266 B 0.025476f
C697 VTAIL.n267 B 0.025476f
C698 VTAIL.n268 B 0.011412f
C699 VTAIL.n269 B 0.010778f
C700 VTAIL.n270 B 0.020058f
C701 VTAIL.n271 B 0.020058f
C702 VTAIL.n272 B 0.010778f
C703 VTAIL.n273 B 0.011412f
C704 VTAIL.n274 B 0.025476f
C705 VTAIL.n275 B 0.025476f
C706 VTAIL.n276 B 0.011412f
C707 VTAIL.n277 B 0.010778f
C708 VTAIL.n278 B 0.020058f
C709 VTAIL.n279 B 0.020058f
C710 VTAIL.n280 B 0.010778f
C711 VTAIL.n281 B 0.011412f
C712 VTAIL.n282 B 0.025476f
C713 VTAIL.n283 B 0.025476f
C714 VTAIL.n284 B 0.025476f
C715 VTAIL.n285 B 0.011095f
C716 VTAIL.n286 B 0.010778f
C717 VTAIL.n287 B 0.020058f
C718 VTAIL.n288 B 0.020058f
C719 VTAIL.n289 B 0.010778f
C720 VTAIL.n290 B 0.011412f
C721 VTAIL.n291 B 0.025476f
C722 VTAIL.n292 B 0.025476f
C723 VTAIL.n293 B 0.011412f
C724 VTAIL.n294 B 0.010778f
C725 VTAIL.n295 B 0.020058f
C726 VTAIL.n296 B 0.020058f
C727 VTAIL.n297 B 0.010778f
C728 VTAIL.n298 B 0.011412f
C729 VTAIL.n299 B 0.025476f
C730 VTAIL.n300 B 0.054911f
C731 VTAIL.n301 B 0.011412f
C732 VTAIL.n302 B 0.010778f
C733 VTAIL.n303 B 0.046089f
C734 VTAIL.n304 B 0.030692f
C735 VTAIL.n305 B 1.68819f
C736 VTAIL.n306 B 0.028058f
C737 VTAIL.n307 B 0.020058f
C738 VTAIL.n308 B 0.010778f
C739 VTAIL.n309 B 0.025476f
C740 VTAIL.n310 B 0.011412f
C741 VTAIL.n311 B 0.020058f
C742 VTAIL.n312 B 0.010778f
C743 VTAIL.n313 B 0.025476f
C744 VTAIL.n314 B 0.011412f
C745 VTAIL.n315 B 0.020058f
C746 VTAIL.n316 B 0.011095f
C747 VTAIL.n317 B 0.025476f
C748 VTAIL.n318 B 0.011412f
C749 VTAIL.n319 B 0.020058f
C750 VTAIL.n320 B 0.010778f
C751 VTAIL.n321 B 0.025476f
C752 VTAIL.n322 B 0.011412f
C753 VTAIL.n323 B 0.020058f
C754 VTAIL.n324 B 0.010778f
C755 VTAIL.n325 B 0.025476f
C756 VTAIL.n326 B 0.011412f
C757 VTAIL.n327 B 0.020058f
C758 VTAIL.n328 B 0.010778f
C759 VTAIL.n329 B 0.025476f
C760 VTAIL.n330 B 0.011412f
C761 VTAIL.n331 B 0.020058f
C762 VTAIL.n332 B 0.010778f
C763 VTAIL.n333 B 0.025476f
C764 VTAIL.n334 B 0.011412f
C765 VTAIL.n335 B 0.020058f
C766 VTAIL.n336 B 0.010778f
C767 VTAIL.n337 B 0.019107f
C768 VTAIL.n338 B 0.015049f
C769 VTAIL.t3 B 0.042229f
C770 VTAIL.n339 B 0.147065f
C771 VTAIL.n340 B 1.6019f
C772 VTAIL.n341 B 0.010778f
C773 VTAIL.n342 B 0.011412f
C774 VTAIL.n343 B 0.025476f
C775 VTAIL.n344 B 0.025476f
C776 VTAIL.n345 B 0.011412f
C777 VTAIL.n346 B 0.010778f
C778 VTAIL.n347 B 0.020058f
C779 VTAIL.n348 B 0.020058f
C780 VTAIL.n349 B 0.010778f
C781 VTAIL.n350 B 0.011412f
C782 VTAIL.n351 B 0.025476f
C783 VTAIL.n352 B 0.025476f
C784 VTAIL.n353 B 0.011412f
C785 VTAIL.n354 B 0.010778f
C786 VTAIL.n355 B 0.020058f
C787 VTAIL.n356 B 0.020058f
C788 VTAIL.n357 B 0.010778f
C789 VTAIL.n358 B 0.011412f
C790 VTAIL.n359 B 0.025476f
C791 VTAIL.n360 B 0.025476f
C792 VTAIL.n361 B 0.011412f
C793 VTAIL.n362 B 0.010778f
C794 VTAIL.n363 B 0.020058f
C795 VTAIL.n364 B 0.020058f
C796 VTAIL.n365 B 0.010778f
C797 VTAIL.n366 B 0.011412f
C798 VTAIL.n367 B 0.025476f
C799 VTAIL.n368 B 0.025476f
C800 VTAIL.n369 B 0.011412f
C801 VTAIL.n370 B 0.010778f
C802 VTAIL.n371 B 0.020058f
C803 VTAIL.n372 B 0.020058f
C804 VTAIL.n373 B 0.010778f
C805 VTAIL.n374 B 0.011412f
C806 VTAIL.n375 B 0.025476f
C807 VTAIL.n376 B 0.025476f
C808 VTAIL.n377 B 0.011412f
C809 VTAIL.n378 B 0.010778f
C810 VTAIL.n379 B 0.020058f
C811 VTAIL.n380 B 0.020058f
C812 VTAIL.n381 B 0.010778f
C813 VTAIL.n382 B 0.010778f
C814 VTAIL.n383 B 0.011412f
C815 VTAIL.n384 B 0.025476f
C816 VTAIL.n385 B 0.025476f
C817 VTAIL.n386 B 0.025476f
C818 VTAIL.n387 B 0.011095f
C819 VTAIL.n388 B 0.010778f
C820 VTAIL.n389 B 0.020058f
C821 VTAIL.n390 B 0.020058f
C822 VTAIL.n391 B 0.010778f
C823 VTAIL.n392 B 0.011412f
C824 VTAIL.n393 B 0.025476f
C825 VTAIL.n394 B 0.025476f
C826 VTAIL.n395 B 0.011412f
C827 VTAIL.n396 B 0.010778f
C828 VTAIL.n397 B 0.020058f
C829 VTAIL.n398 B 0.020058f
C830 VTAIL.n399 B 0.010778f
C831 VTAIL.n400 B 0.011412f
C832 VTAIL.n401 B 0.025476f
C833 VTAIL.n402 B 0.054911f
C834 VTAIL.n403 B 0.011412f
C835 VTAIL.n404 B 0.010778f
C836 VTAIL.n405 B 0.046089f
C837 VTAIL.n406 B 0.030692f
C838 VTAIL.n407 B 1.59528f
C839 VN.t0 B 4.7953f
C840 VN.t1 B 5.53317f
.ends

