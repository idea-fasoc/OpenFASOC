* NGSPICE file created from diff_pair_sample_1636.ext - technology: sky130A

.subckt diff_pair_sample_1636 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=6.6924 pd=35.1 as=0 ps=0 w=17.16 l=0.71
X1 VTAIL.t11 VN.t0 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8314 pd=17.49 as=2.8314 ps=17.49 w=17.16 l=0.71
X2 VDD1.t5 VP.t0 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8314 pd=17.49 as=6.6924 ps=35.1 w=17.16 l=0.71
X3 VDD2.t1 VN.t1 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6924 pd=35.1 as=2.8314 ps=17.49 w=17.16 l=0.71
X4 VTAIL.t5 VP.t1 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8314 pd=17.49 as=2.8314 ps=17.49 w=17.16 l=0.71
X5 VDD1.t3 VP.t2 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8314 pd=17.49 as=6.6924 ps=35.1 w=17.16 l=0.71
X6 VTAIL.t9 VN.t2 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8314 pd=17.49 as=2.8314 ps=17.49 w=17.16 l=0.71
X7 VTAIL.t3 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8314 pd=17.49 as=2.8314 ps=17.49 w=17.16 l=0.71
X8 VDD1.t1 VP.t4 VTAIL.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6924 pd=35.1 as=2.8314 ps=17.49 w=17.16 l=0.71
X9 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=6.6924 pd=35.1 as=0 ps=0 w=17.16 l=0.71
X10 VDD2.t3 VN.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8314 pd=17.49 as=6.6924 ps=35.1 w=17.16 l=0.71
X11 VDD2.t5 VN.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8314 pd=17.49 as=6.6924 ps=35.1 w=17.16 l=0.71
X12 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6924 pd=35.1 as=0 ps=0 w=17.16 l=0.71
X13 VDD1.t0 VP.t5 VTAIL.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6924 pd=35.1 as=2.8314 ps=17.49 w=17.16 l=0.71
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.6924 pd=35.1 as=0 ps=0 w=17.16 l=0.71
X15 VDD2.t2 VN.t5 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6924 pd=35.1 as=2.8314 ps=17.49 w=17.16 l=0.71
R0 B.n107 B.t10 785.317
R1 B.n104 B.t6 785.317
R2 B.n418 B.t17 785.317
R3 B.n424 B.t13 785.317
R4 B.n791 B.n790 585
R5 B.n792 B.n791 585
R6 B.n350 B.n103 585
R7 B.n349 B.n348 585
R8 B.n347 B.n346 585
R9 B.n345 B.n344 585
R10 B.n343 B.n342 585
R11 B.n341 B.n340 585
R12 B.n339 B.n338 585
R13 B.n337 B.n336 585
R14 B.n335 B.n334 585
R15 B.n333 B.n332 585
R16 B.n331 B.n330 585
R17 B.n329 B.n328 585
R18 B.n327 B.n326 585
R19 B.n325 B.n324 585
R20 B.n323 B.n322 585
R21 B.n321 B.n320 585
R22 B.n319 B.n318 585
R23 B.n317 B.n316 585
R24 B.n315 B.n314 585
R25 B.n313 B.n312 585
R26 B.n311 B.n310 585
R27 B.n309 B.n308 585
R28 B.n307 B.n306 585
R29 B.n305 B.n304 585
R30 B.n303 B.n302 585
R31 B.n301 B.n300 585
R32 B.n299 B.n298 585
R33 B.n297 B.n296 585
R34 B.n295 B.n294 585
R35 B.n293 B.n292 585
R36 B.n291 B.n290 585
R37 B.n289 B.n288 585
R38 B.n287 B.n286 585
R39 B.n285 B.n284 585
R40 B.n283 B.n282 585
R41 B.n281 B.n280 585
R42 B.n279 B.n278 585
R43 B.n277 B.n276 585
R44 B.n275 B.n274 585
R45 B.n273 B.n272 585
R46 B.n271 B.n270 585
R47 B.n269 B.n268 585
R48 B.n267 B.n266 585
R49 B.n265 B.n264 585
R50 B.n263 B.n262 585
R51 B.n261 B.n260 585
R52 B.n259 B.n258 585
R53 B.n257 B.n256 585
R54 B.n255 B.n254 585
R55 B.n253 B.n252 585
R56 B.n251 B.n250 585
R57 B.n249 B.n248 585
R58 B.n247 B.n246 585
R59 B.n245 B.n244 585
R60 B.n243 B.n242 585
R61 B.n241 B.n240 585
R62 B.n239 B.n238 585
R63 B.n237 B.n236 585
R64 B.n235 B.n234 585
R65 B.n233 B.n232 585
R66 B.n231 B.n230 585
R67 B.n229 B.n228 585
R68 B.n227 B.n226 585
R69 B.n225 B.n224 585
R70 B.n223 B.n222 585
R71 B.n220 B.n219 585
R72 B.n218 B.n217 585
R73 B.n216 B.n215 585
R74 B.n214 B.n213 585
R75 B.n212 B.n211 585
R76 B.n210 B.n209 585
R77 B.n208 B.n207 585
R78 B.n206 B.n205 585
R79 B.n204 B.n203 585
R80 B.n202 B.n201 585
R81 B.n200 B.n199 585
R82 B.n198 B.n197 585
R83 B.n196 B.n195 585
R84 B.n194 B.n193 585
R85 B.n192 B.n191 585
R86 B.n190 B.n189 585
R87 B.n188 B.n187 585
R88 B.n186 B.n185 585
R89 B.n184 B.n183 585
R90 B.n182 B.n181 585
R91 B.n180 B.n179 585
R92 B.n178 B.n177 585
R93 B.n176 B.n175 585
R94 B.n174 B.n173 585
R95 B.n172 B.n171 585
R96 B.n170 B.n169 585
R97 B.n168 B.n167 585
R98 B.n166 B.n165 585
R99 B.n164 B.n163 585
R100 B.n162 B.n161 585
R101 B.n160 B.n159 585
R102 B.n158 B.n157 585
R103 B.n156 B.n155 585
R104 B.n154 B.n153 585
R105 B.n152 B.n151 585
R106 B.n150 B.n149 585
R107 B.n148 B.n147 585
R108 B.n146 B.n145 585
R109 B.n144 B.n143 585
R110 B.n142 B.n141 585
R111 B.n140 B.n139 585
R112 B.n138 B.n137 585
R113 B.n136 B.n135 585
R114 B.n134 B.n133 585
R115 B.n132 B.n131 585
R116 B.n130 B.n129 585
R117 B.n128 B.n127 585
R118 B.n126 B.n125 585
R119 B.n124 B.n123 585
R120 B.n122 B.n121 585
R121 B.n120 B.n119 585
R122 B.n118 B.n117 585
R123 B.n116 B.n115 585
R124 B.n114 B.n113 585
R125 B.n112 B.n111 585
R126 B.n110 B.n109 585
R127 B.n40 B.n39 585
R128 B.n789 B.n41 585
R129 B.n793 B.n41 585
R130 B.n788 B.n787 585
R131 B.n787 B.n37 585
R132 B.n786 B.n36 585
R133 B.n799 B.n36 585
R134 B.n785 B.n35 585
R135 B.n800 B.n35 585
R136 B.n784 B.n34 585
R137 B.n801 B.n34 585
R138 B.n783 B.n782 585
R139 B.n782 B.n30 585
R140 B.n781 B.n29 585
R141 B.n807 B.n29 585
R142 B.n780 B.n28 585
R143 B.n808 B.n28 585
R144 B.n779 B.n27 585
R145 B.n809 B.n27 585
R146 B.n778 B.n777 585
R147 B.n777 B.n23 585
R148 B.n776 B.n22 585
R149 B.n815 B.n22 585
R150 B.n775 B.n21 585
R151 B.n816 B.n21 585
R152 B.n774 B.n20 585
R153 B.n817 B.n20 585
R154 B.n773 B.n772 585
R155 B.n772 B.n16 585
R156 B.n771 B.n15 585
R157 B.n823 B.n15 585
R158 B.n770 B.n14 585
R159 B.n824 B.n14 585
R160 B.n769 B.n13 585
R161 B.n825 B.n13 585
R162 B.n768 B.n767 585
R163 B.n767 B.n12 585
R164 B.n766 B.n765 585
R165 B.n766 B.n8 585
R166 B.n764 B.n7 585
R167 B.n832 B.n7 585
R168 B.n763 B.n6 585
R169 B.n833 B.n6 585
R170 B.n762 B.n5 585
R171 B.n834 B.n5 585
R172 B.n761 B.n760 585
R173 B.n760 B.n4 585
R174 B.n759 B.n351 585
R175 B.n759 B.n758 585
R176 B.n748 B.n352 585
R177 B.n751 B.n352 585
R178 B.n750 B.n749 585
R179 B.n752 B.n750 585
R180 B.n747 B.n357 585
R181 B.n357 B.n356 585
R182 B.n746 B.n745 585
R183 B.n745 B.n744 585
R184 B.n359 B.n358 585
R185 B.n360 B.n359 585
R186 B.n737 B.n736 585
R187 B.n738 B.n737 585
R188 B.n735 B.n364 585
R189 B.n368 B.n364 585
R190 B.n734 B.n733 585
R191 B.n733 B.n732 585
R192 B.n366 B.n365 585
R193 B.n367 B.n366 585
R194 B.n725 B.n724 585
R195 B.n726 B.n725 585
R196 B.n723 B.n373 585
R197 B.n373 B.n372 585
R198 B.n722 B.n721 585
R199 B.n721 B.n720 585
R200 B.n375 B.n374 585
R201 B.n376 B.n375 585
R202 B.n713 B.n712 585
R203 B.n714 B.n713 585
R204 B.n711 B.n381 585
R205 B.n381 B.n380 585
R206 B.n710 B.n709 585
R207 B.n709 B.n708 585
R208 B.n383 B.n382 585
R209 B.n384 B.n383 585
R210 B.n701 B.n700 585
R211 B.n702 B.n701 585
R212 B.n387 B.n386 585
R213 B.n457 B.n456 585
R214 B.n458 B.n454 585
R215 B.n454 B.n388 585
R216 B.n460 B.n459 585
R217 B.n462 B.n453 585
R218 B.n465 B.n464 585
R219 B.n466 B.n452 585
R220 B.n468 B.n467 585
R221 B.n470 B.n451 585
R222 B.n473 B.n472 585
R223 B.n474 B.n450 585
R224 B.n476 B.n475 585
R225 B.n478 B.n449 585
R226 B.n481 B.n480 585
R227 B.n482 B.n448 585
R228 B.n484 B.n483 585
R229 B.n486 B.n447 585
R230 B.n489 B.n488 585
R231 B.n490 B.n446 585
R232 B.n492 B.n491 585
R233 B.n494 B.n445 585
R234 B.n497 B.n496 585
R235 B.n498 B.n444 585
R236 B.n500 B.n499 585
R237 B.n502 B.n443 585
R238 B.n505 B.n504 585
R239 B.n506 B.n442 585
R240 B.n508 B.n507 585
R241 B.n510 B.n441 585
R242 B.n513 B.n512 585
R243 B.n514 B.n440 585
R244 B.n516 B.n515 585
R245 B.n518 B.n439 585
R246 B.n521 B.n520 585
R247 B.n522 B.n438 585
R248 B.n524 B.n523 585
R249 B.n526 B.n437 585
R250 B.n529 B.n528 585
R251 B.n530 B.n436 585
R252 B.n532 B.n531 585
R253 B.n534 B.n435 585
R254 B.n537 B.n536 585
R255 B.n538 B.n434 585
R256 B.n540 B.n539 585
R257 B.n542 B.n433 585
R258 B.n545 B.n544 585
R259 B.n546 B.n432 585
R260 B.n548 B.n547 585
R261 B.n550 B.n431 585
R262 B.n553 B.n552 585
R263 B.n554 B.n430 585
R264 B.n556 B.n555 585
R265 B.n558 B.n429 585
R266 B.n561 B.n560 585
R267 B.n562 B.n428 585
R268 B.n564 B.n563 585
R269 B.n566 B.n427 585
R270 B.n569 B.n568 585
R271 B.n570 B.n423 585
R272 B.n572 B.n571 585
R273 B.n574 B.n422 585
R274 B.n577 B.n576 585
R275 B.n578 B.n421 585
R276 B.n580 B.n579 585
R277 B.n582 B.n420 585
R278 B.n585 B.n584 585
R279 B.n587 B.n417 585
R280 B.n589 B.n588 585
R281 B.n591 B.n416 585
R282 B.n594 B.n593 585
R283 B.n595 B.n415 585
R284 B.n597 B.n596 585
R285 B.n599 B.n414 585
R286 B.n602 B.n601 585
R287 B.n603 B.n413 585
R288 B.n605 B.n604 585
R289 B.n607 B.n412 585
R290 B.n610 B.n609 585
R291 B.n611 B.n411 585
R292 B.n613 B.n612 585
R293 B.n615 B.n410 585
R294 B.n618 B.n617 585
R295 B.n619 B.n409 585
R296 B.n621 B.n620 585
R297 B.n623 B.n408 585
R298 B.n626 B.n625 585
R299 B.n627 B.n407 585
R300 B.n629 B.n628 585
R301 B.n631 B.n406 585
R302 B.n634 B.n633 585
R303 B.n635 B.n405 585
R304 B.n637 B.n636 585
R305 B.n639 B.n404 585
R306 B.n642 B.n641 585
R307 B.n643 B.n403 585
R308 B.n645 B.n644 585
R309 B.n647 B.n402 585
R310 B.n650 B.n649 585
R311 B.n651 B.n401 585
R312 B.n653 B.n652 585
R313 B.n655 B.n400 585
R314 B.n658 B.n657 585
R315 B.n659 B.n399 585
R316 B.n661 B.n660 585
R317 B.n663 B.n398 585
R318 B.n666 B.n665 585
R319 B.n667 B.n397 585
R320 B.n669 B.n668 585
R321 B.n671 B.n396 585
R322 B.n674 B.n673 585
R323 B.n675 B.n395 585
R324 B.n677 B.n676 585
R325 B.n679 B.n394 585
R326 B.n682 B.n681 585
R327 B.n683 B.n393 585
R328 B.n685 B.n684 585
R329 B.n687 B.n392 585
R330 B.n690 B.n689 585
R331 B.n691 B.n391 585
R332 B.n693 B.n692 585
R333 B.n695 B.n390 585
R334 B.n698 B.n697 585
R335 B.n699 B.n389 585
R336 B.n704 B.n703 585
R337 B.n703 B.n702 585
R338 B.n705 B.n385 585
R339 B.n385 B.n384 585
R340 B.n707 B.n706 585
R341 B.n708 B.n707 585
R342 B.n379 B.n378 585
R343 B.n380 B.n379 585
R344 B.n716 B.n715 585
R345 B.n715 B.n714 585
R346 B.n717 B.n377 585
R347 B.n377 B.n376 585
R348 B.n719 B.n718 585
R349 B.n720 B.n719 585
R350 B.n371 B.n370 585
R351 B.n372 B.n371 585
R352 B.n728 B.n727 585
R353 B.n727 B.n726 585
R354 B.n729 B.n369 585
R355 B.n369 B.n367 585
R356 B.n731 B.n730 585
R357 B.n732 B.n731 585
R358 B.n363 B.n362 585
R359 B.n368 B.n363 585
R360 B.n740 B.n739 585
R361 B.n739 B.n738 585
R362 B.n741 B.n361 585
R363 B.n361 B.n360 585
R364 B.n743 B.n742 585
R365 B.n744 B.n743 585
R366 B.n355 B.n354 585
R367 B.n356 B.n355 585
R368 B.n754 B.n753 585
R369 B.n753 B.n752 585
R370 B.n755 B.n353 585
R371 B.n751 B.n353 585
R372 B.n757 B.n756 585
R373 B.n758 B.n757 585
R374 B.n3 B.n0 585
R375 B.n4 B.n3 585
R376 B.n831 B.n1 585
R377 B.n832 B.n831 585
R378 B.n830 B.n829 585
R379 B.n830 B.n8 585
R380 B.n828 B.n9 585
R381 B.n12 B.n9 585
R382 B.n827 B.n826 585
R383 B.n826 B.n825 585
R384 B.n11 B.n10 585
R385 B.n824 B.n11 585
R386 B.n822 B.n821 585
R387 B.n823 B.n822 585
R388 B.n820 B.n17 585
R389 B.n17 B.n16 585
R390 B.n819 B.n818 585
R391 B.n818 B.n817 585
R392 B.n19 B.n18 585
R393 B.n816 B.n19 585
R394 B.n814 B.n813 585
R395 B.n815 B.n814 585
R396 B.n812 B.n24 585
R397 B.n24 B.n23 585
R398 B.n811 B.n810 585
R399 B.n810 B.n809 585
R400 B.n26 B.n25 585
R401 B.n808 B.n26 585
R402 B.n806 B.n805 585
R403 B.n807 B.n806 585
R404 B.n804 B.n31 585
R405 B.n31 B.n30 585
R406 B.n803 B.n802 585
R407 B.n802 B.n801 585
R408 B.n33 B.n32 585
R409 B.n800 B.n33 585
R410 B.n798 B.n797 585
R411 B.n799 B.n798 585
R412 B.n796 B.n38 585
R413 B.n38 B.n37 585
R414 B.n795 B.n794 585
R415 B.n794 B.n793 585
R416 B.n835 B.n834 585
R417 B.n833 B.n2 585
R418 B.n794 B.n40 487.695
R419 B.n791 B.n41 487.695
R420 B.n701 B.n389 487.695
R421 B.n703 B.n387 487.695
R422 B.n792 B.n102 256.663
R423 B.n792 B.n101 256.663
R424 B.n792 B.n100 256.663
R425 B.n792 B.n99 256.663
R426 B.n792 B.n98 256.663
R427 B.n792 B.n97 256.663
R428 B.n792 B.n96 256.663
R429 B.n792 B.n95 256.663
R430 B.n792 B.n94 256.663
R431 B.n792 B.n93 256.663
R432 B.n792 B.n92 256.663
R433 B.n792 B.n91 256.663
R434 B.n792 B.n90 256.663
R435 B.n792 B.n89 256.663
R436 B.n792 B.n88 256.663
R437 B.n792 B.n87 256.663
R438 B.n792 B.n86 256.663
R439 B.n792 B.n85 256.663
R440 B.n792 B.n84 256.663
R441 B.n792 B.n83 256.663
R442 B.n792 B.n82 256.663
R443 B.n792 B.n81 256.663
R444 B.n792 B.n80 256.663
R445 B.n792 B.n79 256.663
R446 B.n792 B.n78 256.663
R447 B.n792 B.n77 256.663
R448 B.n792 B.n76 256.663
R449 B.n792 B.n75 256.663
R450 B.n792 B.n74 256.663
R451 B.n792 B.n73 256.663
R452 B.n792 B.n72 256.663
R453 B.n792 B.n71 256.663
R454 B.n792 B.n70 256.663
R455 B.n792 B.n69 256.663
R456 B.n792 B.n68 256.663
R457 B.n792 B.n67 256.663
R458 B.n792 B.n66 256.663
R459 B.n792 B.n65 256.663
R460 B.n792 B.n64 256.663
R461 B.n792 B.n63 256.663
R462 B.n792 B.n62 256.663
R463 B.n792 B.n61 256.663
R464 B.n792 B.n60 256.663
R465 B.n792 B.n59 256.663
R466 B.n792 B.n58 256.663
R467 B.n792 B.n57 256.663
R468 B.n792 B.n56 256.663
R469 B.n792 B.n55 256.663
R470 B.n792 B.n54 256.663
R471 B.n792 B.n53 256.663
R472 B.n792 B.n52 256.663
R473 B.n792 B.n51 256.663
R474 B.n792 B.n50 256.663
R475 B.n792 B.n49 256.663
R476 B.n792 B.n48 256.663
R477 B.n792 B.n47 256.663
R478 B.n792 B.n46 256.663
R479 B.n792 B.n45 256.663
R480 B.n792 B.n44 256.663
R481 B.n792 B.n43 256.663
R482 B.n792 B.n42 256.663
R483 B.n455 B.n388 256.663
R484 B.n461 B.n388 256.663
R485 B.n463 B.n388 256.663
R486 B.n469 B.n388 256.663
R487 B.n471 B.n388 256.663
R488 B.n477 B.n388 256.663
R489 B.n479 B.n388 256.663
R490 B.n485 B.n388 256.663
R491 B.n487 B.n388 256.663
R492 B.n493 B.n388 256.663
R493 B.n495 B.n388 256.663
R494 B.n501 B.n388 256.663
R495 B.n503 B.n388 256.663
R496 B.n509 B.n388 256.663
R497 B.n511 B.n388 256.663
R498 B.n517 B.n388 256.663
R499 B.n519 B.n388 256.663
R500 B.n525 B.n388 256.663
R501 B.n527 B.n388 256.663
R502 B.n533 B.n388 256.663
R503 B.n535 B.n388 256.663
R504 B.n541 B.n388 256.663
R505 B.n543 B.n388 256.663
R506 B.n549 B.n388 256.663
R507 B.n551 B.n388 256.663
R508 B.n557 B.n388 256.663
R509 B.n559 B.n388 256.663
R510 B.n565 B.n388 256.663
R511 B.n567 B.n388 256.663
R512 B.n573 B.n388 256.663
R513 B.n575 B.n388 256.663
R514 B.n581 B.n388 256.663
R515 B.n583 B.n388 256.663
R516 B.n590 B.n388 256.663
R517 B.n592 B.n388 256.663
R518 B.n598 B.n388 256.663
R519 B.n600 B.n388 256.663
R520 B.n606 B.n388 256.663
R521 B.n608 B.n388 256.663
R522 B.n614 B.n388 256.663
R523 B.n616 B.n388 256.663
R524 B.n622 B.n388 256.663
R525 B.n624 B.n388 256.663
R526 B.n630 B.n388 256.663
R527 B.n632 B.n388 256.663
R528 B.n638 B.n388 256.663
R529 B.n640 B.n388 256.663
R530 B.n646 B.n388 256.663
R531 B.n648 B.n388 256.663
R532 B.n654 B.n388 256.663
R533 B.n656 B.n388 256.663
R534 B.n662 B.n388 256.663
R535 B.n664 B.n388 256.663
R536 B.n670 B.n388 256.663
R537 B.n672 B.n388 256.663
R538 B.n678 B.n388 256.663
R539 B.n680 B.n388 256.663
R540 B.n686 B.n388 256.663
R541 B.n688 B.n388 256.663
R542 B.n694 B.n388 256.663
R543 B.n696 B.n388 256.663
R544 B.n837 B.n836 256.663
R545 B.n111 B.n110 163.367
R546 B.n115 B.n114 163.367
R547 B.n119 B.n118 163.367
R548 B.n123 B.n122 163.367
R549 B.n127 B.n126 163.367
R550 B.n131 B.n130 163.367
R551 B.n135 B.n134 163.367
R552 B.n139 B.n138 163.367
R553 B.n143 B.n142 163.367
R554 B.n147 B.n146 163.367
R555 B.n151 B.n150 163.367
R556 B.n155 B.n154 163.367
R557 B.n159 B.n158 163.367
R558 B.n163 B.n162 163.367
R559 B.n167 B.n166 163.367
R560 B.n171 B.n170 163.367
R561 B.n175 B.n174 163.367
R562 B.n179 B.n178 163.367
R563 B.n183 B.n182 163.367
R564 B.n187 B.n186 163.367
R565 B.n191 B.n190 163.367
R566 B.n195 B.n194 163.367
R567 B.n199 B.n198 163.367
R568 B.n203 B.n202 163.367
R569 B.n207 B.n206 163.367
R570 B.n211 B.n210 163.367
R571 B.n215 B.n214 163.367
R572 B.n219 B.n218 163.367
R573 B.n224 B.n223 163.367
R574 B.n228 B.n227 163.367
R575 B.n232 B.n231 163.367
R576 B.n236 B.n235 163.367
R577 B.n240 B.n239 163.367
R578 B.n244 B.n243 163.367
R579 B.n248 B.n247 163.367
R580 B.n252 B.n251 163.367
R581 B.n256 B.n255 163.367
R582 B.n260 B.n259 163.367
R583 B.n264 B.n263 163.367
R584 B.n268 B.n267 163.367
R585 B.n272 B.n271 163.367
R586 B.n276 B.n275 163.367
R587 B.n280 B.n279 163.367
R588 B.n284 B.n283 163.367
R589 B.n288 B.n287 163.367
R590 B.n292 B.n291 163.367
R591 B.n296 B.n295 163.367
R592 B.n300 B.n299 163.367
R593 B.n304 B.n303 163.367
R594 B.n308 B.n307 163.367
R595 B.n312 B.n311 163.367
R596 B.n316 B.n315 163.367
R597 B.n320 B.n319 163.367
R598 B.n324 B.n323 163.367
R599 B.n328 B.n327 163.367
R600 B.n332 B.n331 163.367
R601 B.n336 B.n335 163.367
R602 B.n340 B.n339 163.367
R603 B.n344 B.n343 163.367
R604 B.n348 B.n347 163.367
R605 B.n791 B.n103 163.367
R606 B.n701 B.n383 163.367
R607 B.n709 B.n383 163.367
R608 B.n709 B.n381 163.367
R609 B.n713 B.n381 163.367
R610 B.n713 B.n375 163.367
R611 B.n721 B.n375 163.367
R612 B.n721 B.n373 163.367
R613 B.n725 B.n373 163.367
R614 B.n725 B.n366 163.367
R615 B.n733 B.n366 163.367
R616 B.n733 B.n364 163.367
R617 B.n737 B.n364 163.367
R618 B.n737 B.n359 163.367
R619 B.n745 B.n359 163.367
R620 B.n745 B.n357 163.367
R621 B.n750 B.n357 163.367
R622 B.n750 B.n352 163.367
R623 B.n759 B.n352 163.367
R624 B.n760 B.n759 163.367
R625 B.n760 B.n5 163.367
R626 B.n6 B.n5 163.367
R627 B.n7 B.n6 163.367
R628 B.n766 B.n7 163.367
R629 B.n767 B.n766 163.367
R630 B.n767 B.n13 163.367
R631 B.n14 B.n13 163.367
R632 B.n15 B.n14 163.367
R633 B.n772 B.n15 163.367
R634 B.n772 B.n20 163.367
R635 B.n21 B.n20 163.367
R636 B.n22 B.n21 163.367
R637 B.n777 B.n22 163.367
R638 B.n777 B.n27 163.367
R639 B.n28 B.n27 163.367
R640 B.n29 B.n28 163.367
R641 B.n782 B.n29 163.367
R642 B.n782 B.n34 163.367
R643 B.n35 B.n34 163.367
R644 B.n36 B.n35 163.367
R645 B.n787 B.n36 163.367
R646 B.n787 B.n41 163.367
R647 B.n456 B.n454 163.367
R648 B.n460 B.n454 163.367
R649 B.n464 B.n462 163.367
R650 B.n468 B.n452 163.367
R651 B.n472 B.n470 163.367
R652 B.n476 B.n450 163.367
R653 B.n480 B.n478 163.367
R654 B.n484 B.n448 163.367
R655 B.n488 B.n486 163.367
R656 B.n492 B.n446 163.367
R657 B.n496 B.n494 163.367
R658 B.n500 B.n444 163.367
R659 B.n504 B.n502 163.367
R660 B.n508 B.n442 163.367
R661 B.n512 B.n510 163.367
R662 B.n516 B.n440 163.367
R663 B.n520 B.n518 163.367
R664 B.n524 B.n438 163.367
R665 B.n528 B.n526 163.367
R666 B.n532 B.n436 163.367
R667 B.n536 B.n534 163.367
R668 B.n540 B.n434 163.367
R669 B.n544 B.n542 163.367
R670 B.n548 B.n432 163.367
R671 B.n552 B.n550 163.367
R672 B.n556 B.n430 163.367
R673 B.n560 B.n558 163.367
R674 B.n564 B.n428 163.367
R675 B.n568 B.n566 163.367
R676 B.n572 B.n423 163.367
R677 B.n576 B.n574 163.367
R678 B.n580 B.n421 163.367
R679 B.n584 B.n582 163.367
R680 B.n589 B.n417 163.367
R681 B.n593 B.n591 163.367
R682 B.n597 B.n415 163.367
R683 B.n601 B.n599 163.367
R684 B.n605 B.n413 163.367
R685 B.n609 B.n607 163.367
R686 B.n613 B.n411 163.367
R687 B.n617 B.n615 163.367
R688 B.n621 B.n409 163.367
R689 B.n625 B.n623 163.367
R690 B.n629 B.n407 163.367
R691 B.n633 B.n631 163.367
R692 B.n637 B.n405 163.367
R693 B.n641 B.n639 163.367
R694 B.n645 B.n403 163.367
R695 B.n649 B.n647 163.367
R696 B.n653 B.n401 163.367
R697 B.n657 B.n655 163.367
R698 B.n661 B.n399 163.367
R699 B.n665 B.n663 163.367
R700 B.n669 B.n397 163.367
R701 B.n673 B.n671 163.367
R702 B.n677 B.n395 163.367
R703 B.n681 B.n679 163.367
R704 B.n685 B.n393 163.367
R705 B.n689 B.n687 163.367
R706 B.n693 B.n391 163.367
R707 B.n697 B.n695 163.367
R708 B.n703 B.n385 163.367
R709 B.n707 B.n385 163.367
R710 B.n707 B.n379 163.367
R711 B.n715 B.n379 163.367
R712 B.n715 B.n377 163.367
R713 B.n719 B.n377 163.367
R714 B.n719 B.n371 163.367
R715 B.n727 B.n371 163.367
R716 B.n727 B.n369 163.367
R717 B.n731 B.n369 163.367
R718 B.n731 B.n363 163.367
R719 B.n739 B.n363 163.367
R720 B.n739 B.n361 163.367
R721 B.n743 B.n361 163.367
R722 B.n743 B.n355 163.367
R723 B.n753 B.n355 163.367
R724 B.n753 B.n353 163.367
R725 B.n757 B.n353 163.367
R726 B.n757 B.n3 163.367
R727 B.n835 B.n3 163.367
R728 B.n831 B.n2 163.367
R729 B.n831 B.n830 163.367
R730 B.n830 B.n9 163.367
R731 B.n826 B.n9 163.367
R732 B.n826 B.n11 163.367
R733 B.n822 B.n11 163.367
R734 B.n822 B.n17 163.367
R735 B.n818 B.n17 163.367
R736 B.n818 B.n19 163.367
R737 B.n814 B.n19 163.367
R738 B.n814 B.n24 163.367
R739 B.n810 B.n24 163.367
R740 B.n810 B.n26 163.367
R741 B.n806 B.n26 163.367
R742 B.n806 B.n31 163.367
R743 B.n802 B.n31 163.367
R744 B.n802 B.n33 163.367
R745 B.n798 B.n33 163.367
R746 B.n798 B.n38 163.367
R747 B.n794 B.n38 163.367
R748 B.n104 B.t8 90.574
R749 B.n418 B.t19 90.574
R750 B.n107 B.t11 90.5512
R751 B.n424 B.t16 90.5512
R752 B.n42 B.n40 71.676
R753 B.n111 B.n43 71.676
R754 B.n115 B.n44 71.676
R755 B.n119 B.n45 71.676
R756 B.n123 B.n46 71.676
R757 B.n127 B.n47 71.676
R758 B.n131 B.n48 71.676
R759 B.n135 B.n49 71.676
R760 B.n139 B.n50 71.676
R761 B.n143 B.n51 71.676
R762 B.n147 B.n52 71.676
R763 B.n151 B.n53 71.676
R764 B.n155 B.n54 71.676
R765 B.n159 B.n55 71.676
R766 B.n163 B.n56 71.676
R767 B.n167 B.n57 71.676
R768 B.n171 B.n58 71.676
R769 B.n175 B.n59 71.676
R770 B.n179 B.n60 71.676
R771 B.n183 B.n61 71.676
R772 B.n187 B.n62 71.676
R773 B.n191 B.n63 71.676
R774 B.n195 B.n64 71.676
R775 B.n199 B.n65 71.676
R776 B.n203 B.n66 71.676
R777 B.n207 B.n67 71.676
R778 B.n211 B.n68 71.676
R779 B.n215 B.n69 71.676
R780 B.n219 B.n70 71.676
R781 B.n224 B.n71 71.676
R782 B.n228 B.n72 71.676
R783 B.n232 B.n73 71.676
R784 B.n236 B.n74 71.676
R785 B.n240 B.n75 71.676
R786 B.n244 B.n76 71.676
R787 B.n248 B.n77 71.676
R788 B.n252 B.n78 71.676
R789 B.n256 B.n79 71.676
R790 B.n260 B.n80 71.676
R791 B.n264 B.n81 71.676
R792 B.n268 B.n82 71.676
R793 B.n272 B.n83 71.676
R794 B.n276 B.n84 71.676
R795 B.n280 B.n85 71.676
R796 B.n284 B.n86 71.676
R797 B.n288 B.n87 71.676
R798 B.n292 B.n88 71.676
R799 B.n296 B.n89 71.676
R800 B.n300 B.n90 71.676
R801 B.n304 B.n91 71.676
R802 B.n308 B.n92 71.676
R803 B.n312 B.n93 71.676
R804 B.n316 B.n94 71.676
R805 B.n320 B.n95 71.676
R806 B.n324 B.n96 71.676
R807 B.n328 B.n97 71.676
R808 B.n332 B.n98 71.676
R809 B.n336 B.n99 71.676
R810 B.n340 B.n100 71.676
R811 B.n344 B.n101 71.676
R812 B.n348 B.n102 71.676
R813 B.n103 B.n102 71.676
R814 B.n347 B.n101 71.676
R815 B.n343 B.n100 71.676
R816 B.n339 B.n99 71.676
R817 B.n335 B.n98 71.676
R818 B.n331 B.n97 71.676
R819 B.n327 B.n96 71.676
R820 B.n323 B.n95 71.676
R821 B.n319 B.n94 71.676
R822 B.n315 B.n93 71.676
R823 B.n311 B.n92 71.676
R824 B.n307 B.n91 71.676
R825 B.n303 B.n90 71.676
R826 B.n299 B.n89 71.676
R827 B.n295 B.n88 71.676
R828 B.n291 B.n87 71.676
R829 B.n287 B.n86 71.676
R830 B.n283 B.n85 71.676
R831 B.n279 B.n84 71.676
R832 B.n275 B.n83 71.676
R833 B.n271 B.n82 71.676
R834 B.n267 B.n81 71.676
R835 B.n263 B.n80 71.676
R836 B.n259 B.n79 71.676
R837 B.n255 B.n78 71.676
R838 B.n251 B.n77 71.676
R839 B.n247 B.n76 71.676
R840 B.n243 B.n75 71.676
R841 B.n239 B.n74 71.676
R842 B.n235 B.n73 71.676
R843 B.n231 B.n72 71.676
R844 B.n227 B.n71 71.676
R845 B.n223 B.n70 71.676
R846 B.n218 B.n69 71.676
R847 B.n214 B.n68 71.676
R848 B.n210 B.n67 71.676
R849 B.n206 B.n66 71.676
R850 B.n202 B.n65 71.676
R851 B.n198 B.n64 71.676
R852 B.n194 B.n63 71.676
R853 B.n190 B.n62 71.676
R854 B.n186 B.n61 71.676
R855 B.n182 B.n60 71.676
R856 B.n178 B.n59 71.676
R857 B.n174 B.n58 71.676
R858 B.n170 B.n57 71.676
R859 B.n166 B.n56 71.676
R860 B.n162 B.n55 71.676
R861 B.n158 B.n54 71.676
R862 B.n154 B.n53 71.676
R863 B.n150 B.n52 71.676
R864 B.n146 B.n51 71.676
R865 B.n142 B.n50 71.676
R866 B.n138 B.n49 71.676
R867 B.n134 B.n48 71.676
R868 B.n130 B.n47 71.676
R869 B.n126 B.n46 71.676
R870 B.n122 B.n45 71.676
R871 B.n118 B.n44 71.676
R872 B.n114 B.n43 71.676
R873 B.n110 B.n42 71.676
R874 B.n455 B.n387 71.676
R875 B.n461 B.n460 71.676
R876 B.n464 B.n463 71.676
R877 B.n469 B.n468 71.676
R878 B.n472 B.n471 71.676
R879 B.n477 B.n476 71.676
R880 B.n480 B.n479 71.676
R881 B.n485 B.n484 71.676
R882 B.n488 B.n487 71.676
R883 B.n493 B.n492 71.676
R884 B.n496 B.n495 71.676
R885 B.n501 B.n500 71.676
R886 B.n504 B.n503 71.676
R887 B.n509 B.n508 71.676
R888 B.n512 B.n511 71.676
R889 B.n517 B.n516 71.676
R890 B.n520 B.n519 71.676
R891 B.n525 B.n524 71.676
R892 B.n528 B.n527 71.676
R893 B.n533 B.n532 71.676
R894 B.n536 B.n535 71.676
R895 B.n541 B.n540 71.676
R896 B.n544 B.n543 71.676
R897 B.n549 B.n548 71.676
R898 B.n552 B.n551 71.676
R899 B.n557 B.n556 71.676
R900 B.n560 B.n559 71.676
R901 B.n565 B.n564 71.676
R902 B.n568 B.n567 71.676
R903 B.n573 B.n572 71.676
R904 B.n576 B.n575 71.676
R905 B.n581 B.n580 71.676
R906 B.n584 B.n583 71.676
R907 B.n590 B.n589 71.676
R908 B.n593 B.n592 71.676
R909 B.n598 B.n597 71.676
R910 B.n601 B.n600 71.676
R911 B.n606 B.n605 71.676
R912 B.n609 B.n608 71.676
R913 B.n614 B.n613 71.676
R914 B.n617 B.n616 71.676
R915 B.n622 B.n621 71.676
R916 B.n625 B.n624 71.676
R917 B.n630 B.n629 71.676
R918 B.n633 B.n632 71.676
R919 B.n638 B.n637 71.676
R920 B.n641 B.n640 71.676
R921 B.n646 B.n645 71.676
R922 B.n649 B.n648 71.676
R923 B.n654 B.n653 71.676
R924 B.n657 B.n656 71.676
R925 B.n662 B.n661 71.676
R926 B.n665 B.n664 71.676
R927 B.n670 B.n669 71.676
R928 B.n673 B.n672 71.676
R929 B.n678 B.n677 71.676
R930 B.n681 B.n680 71.676
R931 B.n686 B.n685 71.676
R932 B.n689 B.n688 71.676
R933 B.n694 B.n693 71.676
R934 B.n697 B.n696 71.676
R935 B.n456 B.n455 71.676
R936 B.n462 B.n461 71.676
R937 B.n463 B.n452 71.676
R938 B.n470 B.n469 71.676
R939 B.n471 B.n450 71.676
R940 B.n478 B.n477 71.676
R941 B.n479 B.n448 71.676
R942 B.n486 B.n485 71.676
R943 B.n487 B.n446 71.676
R944 B.n494 B.n493 71.676
R945 B.n495 B.n444 71.676
R946 B.n502 B.n501 71.676
R947 B.n503 B.n442 71.676
R948 B.n510 B.n509 71.676
R949 B.n511 B.n440 71.676
R950 B.n518 B.n517 71.676
R951 B.n519 B.n438 71.676
R952 B.n526 B.n525 71.676
R953 B.n527 B.n436 71.676
R954 B.n534 B.n533 71.676
R955 B.n535 B.n434 71.676
R956 B.n542 B.n541 71.676
R957 B.n543 B.n432 71.676
R958 B.n550 B.n549 71.676
R959 B.n551 B.n430 71.676
R960 B.n558 B.n557 71.676
R961 B.n559 B.n428 71.676
R962 B.n566 B.n565 71.676
R963 B.n567 B.n423 71.676
R964 B.n574 B.n573 71.676
R965 B.n575 B.n421 71.676
R966 B.n582 B.n581 71.676
R967 B.n583 B.n417 71.676
R968 B.n591 B.n590 71.676
R969 B.n592 B.n415 71.676
R970 B.n599 B.n598 71.676
R971 B.n600 B.n413 71.676
R972 B.n607 B.n606 71.676
R973 B.n608 B.n411 71.676
R974 B.n615 B.n614 71.676
R975 B.n616 B.n409 71.676
R976 B.n623 B.n622 71.676
R977 B.n624 B.n407 71.676
R978 B.n631 B.n630 71.676
R979 B.n632 B.n405 71.676
R980 B.n639 B.n638 71.676
R981 B.n640 B.n403 71.676
R982 B.n647 B.n646 71.676
R983 B.n648 B.n401 71.676
R984 B.n655 B.n654 71.676
R985 B.n656 B.n399 71.676
R986 B.n663 B.n662 71.676
R987 B.n664 B.n397 71.676
R988 B.n671 B.n670 71.676
R989 B.n672 B.n395 71.676
R990 B.n679 B.n678 71.676
R991 B.n680 B.n393 71.676
R992 B.n687 B.n686 71.676
R993 B.n688 B.n391 71.676
R994 B.n695 B.n694 71.676
R995 B.n696 B.n389 71.676
R996 B.n836 B.n835 71.676
R997 B.n836 B.n2 71.676
R998 B.n105 B.t9 70.4043
R999 B.n419 B.t18 70.4043
R1000 B.n108 B.t12 70.3815
R1001 B.n425 B.t15 70.3815
R1002 B.n221 B.n108 59.5399
R1003 B.n106 B.n105 59.5399
R1004 B.n586 B.n419 59.5399
R1005 B.n426 B.n425 59.5399
R1006 B.n702 B.n388 55.405
R1007 B.n793 B.n792 55.405
R1008 B.n702 B.n384 33.3413
R1009 B.n708 B.n384 33.3413
R1010 B.n708 B.n380 33.3413
R1011 B.n714 B.n380 33.3413
R1012 B.n720 B.n376 33.3413
R1013 B.n720 B.n372 33.3413
R1014 B.n726 B.n372 33.3413
R1015 B.n726 B.n367 33.3413
R1016 B.n732 B.n367 33.3413
R1017 B.n732 B.n368 33.3413
R1018 B.n738 B.n360 33.3413
R1019 B.n744 B.n360 33.3413
R1020 B.n752 B.n356 33.3413
R1021 B.n752 B.n751 33.3413
R1022 B.n758 B.n4 33.3413
R1023 B.n834 B.n4 33.3413
R1024 B.n834 B.n833 33.3413
R1025 B.n833 B.n832 33.3413
R1026 B.n832 B.n8 33.3413
R1027 B.n825 B.n12 33.3413
R1028 B.n825 B.n824 33.3413
R1029 B.n823 B.n16 33.3413
R1030 B.n817 B.n16 33.3413
R1031 B.n816 B.n815 33.3413
R1032 B.n815 B.n23 33.3413
R1033 B.n809 B.n23 33.3413
R1034 B.n809 B.n808 33.3413
R1035 B.n808 B.n807 33.3413
R1036 B.n807 B.n30 33.3413
R1037 B.n801 B.n800 33.3413
R1038 B.n800 B.n799 33.3413
R1039 B.n799 B.n37 33.3413
R1040 B.n793 B.n37 33.3413
R1041 B.n714 B.t14 32.851
R1042 B.n801 B.t7 32.851
R1043 B.n704 B.n386 31.6883
R1044 B.n700 B.n699 31.6883
R1045 B.n790 B.n789 31.6883
R1046 B.n795 B.n39 31.6883
R1047 B.n738 B.t5 25.0061
R1048 B.n817 B.t2 25.0061
R1049 B.t0 B.n356 23.0448
R1050 B.n824 B.t3 23.0448
R1051 B.n758 B.t1 21.0836
R1052 B.t4 B.n8 21.0836
R1053 B.n108 B.n107 20.1702
R1054 B.n105 B.n104 20.1702
R1055 B.n419 B.n418 20.1702
R1056 B.n425 B.n424 20.1702
R1057 B B.n837 18.0485
R1058 B.n751 B.t1 12.2581
R1059 B.n12 B.t4 12.2581
R1060 B.n705 B.n704 10.6151
R1061 B.n706 B.n705 10.6151
R1062 B.n706 B.n378 10.6151
R1063 B.n716 B.n378 10.6151
R1064 B.n717 B.n716 10.6151
R1065 B.n718 B.n717 10.6151
R1066 B.n718 B.n370 10.6151
R1067 B.n728 B.n370 10.6151
R1068 B.n729 B.n728 10.6151
R1069 B.n730 B.n729 10.6151
R1070 B.n730 B.n362 10.6151
R1071 B.n740 B.n362 10.6151
R1072 B.n741 B.n740 10.6151
R1073 B.n742 B.n741 10.6151
R1074 B.n742 B.n354 10.6151
R1075 B.n754 B.n354 10.6151
R1076 B.n755 B.n754 10.6151
R1077 B.n756 B.n755 10.6151
R1078 B.n756 B.n0 10.6151
R1079 B.n457 B.n386 10.6151
R1080 B.n458 B.n457 10.6151
R1081 B.n459 B.n458 10.6151
R1082 B.n459 B.n453 10.6151
R1083 B.n465 B.n453 10.6151
R1084 B.n466 B.n465 10.6151
R1085 B.n467 B.n466 10.6151
R1086 B.n467 B.n451 10.6151
R1087 B.n473 B.n451 10.6151
R1088 B.n474 B.n473 10.6151
R1089 B.n475 B.n474 10.6151
R1090 B.n475 B.n449 10.6151
R1091 B.n481 B.n449 10.6151
R1092 B.n482 B.n481 10.6151
R1093 B.n483 B.n482 10.6151
R1094 B.n483 B.n447 10.6151
R1095 B.n489 B.n447 10.6151
R1096 B.n490 B.n489 10.6151
R1097 B.n491 B.n490 10.6151
R1098 B.n491 B.n445 10.6151
R1099 B.n497 B.n445 10.6151
R1100 B.n498 B.n497 10.6151
R1101 B.n499 B.n498 10.6151
R1102 B.n499 B.n443 10.6151
R1103 B.n505 B.n443 10.6151
R1104 B.n506 B.n505 10.6151
R1105 B.n507 B.n506 10.6151
R1106 B.n507 B.n441 10.6151
R1107 B.n513 B.n441 10.6151
R1108 B.n514 B.n513 10.6151
R1109 B.n515 B.n514 10.6151
R1110 B.n515 B.n439 10.6151
R1111 B.n521 B.n439 10.6151
R1112 B.n522 B.n521 10.6151
R1113 B.n523 B.n522 10.6151
R1114 B.n523 B.n437 10.6151
R1115 B.n529 B.n437 10.6151
R1116 B.n530 B.n529 10.6151
R1117 B.n531 B.n530 10.6151
R1118 B.n531 B.n435 10.6151
R1119 B.n537 B.n435 10.6151
R1120 B.n538 B.n537 10.6151
R1121 B.n539 B.n538 10.6151
R1122 B.n539 B.n433 10.6151
R1123 B.n545 B.n433 10.6151
R1124 B.n546 B.n545 10.6151
R1125 B.n547 B.n546 10.6151
R1126 B.n547 B.n431 10.6151
R1127 B.n553 B.n431 10.6151
R1128 B.n554 B.n553 10.6151
R1129 B.n555 B.n554 10.6151
R1130 B.n555 B.n429 10.6151
R1131 B.n561 B.n429 10.6151
R1132 B.n562 B.n561 10.6151
R1133 B.n563 B.n562 10.6151
R1134 B.n563 B.n427 10.6151
R1135 B.n570 B.n569 10.6151
R1136 B.n571 B.n570 10.6151
R1137 B.n571 B.n422 10.6151
R1138 B.n577 B.n422 10.6151
R1139 B.n578 B.n577 10.6151
R1140 B.n579 B.n578 10.6151
R1141 B.n579 B.n420 10.6151
R1142 B.n585 B.n420 10.6151
R1143 B.n588 B.n587 10.6151
R1144 B.n588 B.n416 10.6151
R1145 B.n594 B.n416 10.6151
R1146 B.n595 B.n594 10.6151
R1147 B.n596 B.n595 10.6151
R1148 B.n596 B.n414 10.6151
R1149 B.n602 B.n414 10.6151
R1150 B.n603 B.n602 10.6151
R1151 B.n604 B.n603 10.6151
R1152 B.n604 B.n412 10.6151
R1153 B.n610 B.n412 10.6151
R1154 B.n611 B.n610 10.6151
R1155 B.n612 B.n611 10.6151
R1156 B.n612 B.n410 10.6151
R1157 B.n618 B.n410 10.6151
R1158 B.n619 B.n618 10.6151
R1159 B.n620 B.n619 10.6151
R1160 B.n620 B.n408 10.6151
R1161 B.n626 B.n408 10.6151
R1162 B.n627 B.n626 10.6151
R1163 B.n628 B.n627 10.6151
R1164 B.n628 B.n406 10.6151
R1165 B.n634 B.n406 10.6151
R1166 B.n635 B.n634 10.6151
R1167 B.n636 B.n635 10.6151
R1168 B.n636 B.n404 10.6151
R1169 B.n642 B.n404 10.6151
R1170 B.n643 B.n642 10.6151
R1171 B.n644 B.n643 10.6151
R1172 B.n644 B.n402 10.6151
R1173 B.n650 B.n402 10.6151
R1174 B.n651 B.n650 10.6151
R1175 B.n652 B.n651 10.6151
R1176 B.n652 B.n400 10.6151
R1177 B.n658 B.n400 10.6151
R1178 B.n659 B.n658 10.6151
R1179 B.n660 B.n659 10.6151
R1180 B.n660 B.n398 10.6151
R1181 B.n666 B.n398 10.6151
R1182 B.n667 B.n666 10.6151
R1183 B.n668 B.n667 10.6151
R1184 B.n668 B.n396 10.6151
R1185 B.n674 B.n396 10.6151
R1186 B.n675 B.n674 10.6151
R1187 B.n676 B.n675 10.6151
R1188 B.n676 B.n394 10.6151
R1189 B.n682 B.n394 10.6151
R1190 B.n683 B.n682 10.6151
R1191 B.n684 B.n683 10.6151
R1192 B.n684 B.n392 10.6151
R1193 B.n690 B.n392 10.6151
R1194 B.n691 B.n690 10.6151
R1195 B.n692 B.n691 10.6151
R1196 B.n692 B.n390 10.6151
R1197 B.n698 B.n390 10.6151
R1198 B.n699 B.n698 10.6151
R1199 B.n700 B.n382 10.6151
R1200 B.n710 B.n382 10.6151
R1201 B.n711 B.n710 10.6151
R1202 B.n712 B.n711 10.6151
R1203 B.n712 B.n374 10.6151
R1204 B.n722 B.n374 10.6151
R1205 B.n723 B.n722 10.6151
R1206 B.n724 B.n723 10.6151
R1207 B.n724 B.n365 10.6151
R1208 B.n734 B.n365 10.6151
R1209 B.n735 B.n734 10.6151
R1210 B.n736 B.n735 10.6151
R1211 B.n736 B.n358 10.6151
R1212 B.n746 B.n358 10.6151
R1213 B.n747 B.n746 10.6151
R1214 B.n749 B.n747 10.6151
R1215 B.n749 B.n748 10.6151
R1216 B.n748 B.n351 10.6151
R1217 B.n761 B.n351 10.6151
R1218 B.n762 B.n761 10.6151
R1219 B.n763 B.n762 10.6151
R1220 B.n764 B.n763 10.6151
R1221 B.n765 B.n764 10.6151
R1222 B.n768 B.n765 10.6151
R1223 B.n769 B.n768 10.6151
R1224 B.n770 B.n769 10.6151
R1225 B.n771 B.n770 10.6151
R1226 B.n773 B.n771 10.6151
R1227 B.n774 B.n773 10.6151
R1228 B.n775 B.n774 10.6151
R1229 B.n776 B.n775 10.6151
R1230 B.n778 B.n776 10.6151
R1231 B.n779 B.n778 10.6151
R1232 B.n780 B.n779 10.6151
R1233 B.n781 B.n780 10.6151
R1234 B.n783 B.n781 10.6151
R1235 B.n784 B.n783 10.6151
R1236 B.n785 B.n784 10.6151
R1237 B.n786 B.n785 10.6151
R1238 B.n788 B.n786 10.6151
R1239 B.n789 B.n788 10.6151
R1240 B.n829 B.n1 10.6151
R1241 B.n829 B.n828 10.6151
R1242 B.n828 B.n827 10.6151
R1243 B.n827 B.n10 10.6151
R1244 B.n821 B.n10 10.6151
R1245 B.n821 B.n820 10.6151
R1246 B.n820 B.n819 10.6151
R1247 B.n819 B.n18 10.6151
R1248 B.n813 B.n18 10.6151
R1249 B.n813 B.n812 10.6151
R1250 B.n812 B.n811 10.6151
R1251 B.n811 B.n25 10.6151
R1252 B.n805 B.n25 10.6151
R1253 B.n805 B.n804 10.6151
R1254 B.n804 B.n803 10.6151
R1255 B.n803 B.n32 10.6151
R1256 B.n797 B.n32 10.6151
R1257 B.n797 B.n796 10.6151
R1258 B.n796 B.n795 10.6151
R1259 B.n109 B.n39 10.6151
R1260 B.n112 B.n109 10.6151
R1261 B.n113 B.n112 10.6151
R1262 B.n116 B.n113 10.6151
R1263 B.n117 B.n116 10.6151
R1264 B.n120 B.n117 10.6151
R1265 B.n121 B.n120 10.6151
R1266 B.n124 B.n121 10.6151
R1267 B.n125 B.n124 10.6151
R1268 B.n128 B.n125 10.6151
R1269 B.n129 B.n128 10.6151
R1270 B.n132 B.n129 10.6151
R1271 B.n133 B.n132 10.6151
R1272 B.n136 B.n133 10.6151
R1273 B.n137 B.n136 10.6151
R1274 B.n140 B.n137 10.6151
R1275 B.n141 B.n140 10.6151
R1276 B.n144 B.n141 10.6151
R1277 B.n145 B.n144 10.6151
R1278 B.n148 B.n145 10.6151
R1279 B.n149 B.n148 10.6151
R1280 B.n152 B.n149 10.6151
R1281 B.n153 B.n152 10.6151
R1282 B.n156 B.n153 10.6151
R1283 B.n157 B.n156 10.6151
R1284 B.n160 B.n157 10.6151
R1285 B.n161 B.n160 10.6151
R1286 B.n164 B.n161 10.6151
R1287 B.n165 B.n164 10.6151
R1288 B.n168 B.n165 10.6151
R1289 B.n169 B.n168 10.6151
R1290 B.n172 B.n169 10.6151
R1291 B.n173 B.n172 10.6151
R1292 B.n176 B.n173 10.6151
R1293 B.n177 B.n176 10.6151
R1294 B.n180 B.n177 10.6151
R1295 B.n181 B.n180 10.6151
R1296 B.n184 B.n181 10.6151
R1297 B.n185 B.n184 10.6151
R1298 B.n188 B.n185 10.6151
R1299 B.n189 B.n188 10.6151
R1300 B.n192 B.n189 10.6151
R1301 B.n193 B.n192 10.6151
R1302 B.n196 B.n193 10.6151
R1303 B.n197 B.n196 10.6151
R1304 B.n200 B.n197 10.6151
R1305 B.n201 B.n200 10.6151
R1306 B.n204 B.n201 10.6151
R1307 B.n205 B.n204 10.6151
R1308 B.n208 B.n205 10.6151
R1309 B.n209 B.n208 10.6151
R1310 B.n212 B.n209 10.6151
R1311 B.n213 B.n212 10.6151
R1312 B.n216 B.n213 10.6151
R1313 B.n217 B.n216 10.6151
R1314 B.n220 B.n217 10.6151
R1315 B.n225 B.n222 10.6151
R1316 B.n226 B.n225 10.6151
R1317 B.n229 B.n226 10.6151
R1318 B.n230 B.n229 10.6151
R1319 B.n233 B.n230 10.6151
R1320 B.n234 B.n233 10.6151
R1321 B.n237 B.n234 10.6151
R1322 B.n238 B.n237 10.6151
R1323 B.n242 B.n241 10.6151
R1324 B.n245 B.n242 10.6151
R1325 B.n246 B.n245 10.6151
R1326 B.n249 B.n246 10.6151
R1327 B.n250 B.n249 10.6151
R1328 B.n253 B.n250 10.6151
R1329 B.n254 B.n253 10.6151
R1330 B.n257 B.n254 10.6151
R1331 B.n258 B.n257 10.6151
R1332 B.n261 B.n258 10.6151
R1333 B.n262 B.n261 10.6151
R1334 B.n265 B.n262 10.6151
R1335 B.n266 B.n265 10.6151
R1336 B.n269 B.n266 10.6151
R1337 B.n270 B.n269 10.6151
R1338 B.n273 B.n270 10.6151
R1339 B.n274 B.n273 10.6151
R1340 B.n277 B.n274 10.6151
R1341 B.n278 B.n277 10.6151
R1342 B.n281 B.n278 10.6151
R1343 B.n282 B.n281 10.6151
R1344 B.n285 B.n282 10.6151
R1345 B.n286 B.n285 10.6151
R1346 B.n289 B.n286 10.6151
R1347 B.n290 B.n289 10.6151
R1348 B.n293 B.n290 10.6151
R1349 B.n294 B.n293 10.6151
R1350 B.n297 B.n294 10.6151
R1351 B.n298 B.n297 10.6151
R1352 B.n301 B.n298 10.6151
R1353 B.n302 B.n301 10.6151
R1354 B.n305 B.n302 10.6151
R1355 B.n306 B.n305 10.6151
R1356 B.n309 B.n306 10.6151
R1357 B.n310 B.n309 10.6151
R1358 B.n313 B.n310 10.6151
R1359 B.n314 B.n313 10.6151
R1360 B.n317 B.n314 10.6151
R1361 B.n318 B.n317 10.6151
R1362 B.n321 B.n318 10.6151
R1363 B.n322 B.n321 10.6151
R1364 B.n325 B.n322 10.6151
R1365 B.n326 B.n325 10.6151
R1366 B.n329 B.n326 10.6151
R1367 B.n330 B.n329 10.6151
R1368 B.n333 B.n330 10.6151
R1369 B.n334 B.n333 10.6151
R1370 B.n337 B.n334 10.6151
R1371 B.n338 B.n337 10.6151
R1372 B.n341 B.n338 10.6151
R1373 B.n342 B.n341 10.6151
R1374 B.n345 B.n342 10.6151
R1375 B.n346 B.n345 10.6151
R1376 B.n349 B.n346 10.6151
R1377 B.n350 B.n349 10.6151
R1378 B.n790 B.n350 10.6151
R1379 B.n744 B.t0 10.2969
R1380 B.t3 B.n823 10.2969
R1381 B.n368 B.t5 8.33569
R1382 B.t2 B.n816 8.33569
R1383 B.n837 B.n0 8.11757
R1384 B.n837 B.n1 8.11757
R1385 B.n569 B.n426 6.5566
R1386 B.n586 B.n585 6.5566
R1387 B.n222 B.n221 6.5566
R1388 B.n238 B.n106 6.5566
R1389 B.n427 B.n426 4.05904
R1390 B.n587 B.n586 4.05904
R1391 B.n221 B.n220 4.05904
R1392 B.n241 B.n106 4.05904
R1393 B.t14 B.n376 0.490805
R1394 B.t7 B.n30 0.490805
R1395 VN.n1 VN.t5 659.592
R1396 VN.n7 VN.t4 659.592
R1397 VN.n2 VN.t0 637.802
R1398 VN.n4 VN.t3 637.802
R1399 VN.n8 VN.t2 637.802
R1400 VN.n10 VN.t1 637.802
R1401 VN.n5 VN.n4 161.3
R1402 VN.n11 VN.n10 161.3
R1403 VN.n9 VN.n6 161.3
R1404 VN.n3 VN.n0 161.3
R1405 VN VN.n11 45.5403
R1406 VN.n7 VN.n6 44.8565
R1407 VN.n1 VN.n0 44.8565
R1408 VN.n4 VN.n3 27.0217
R1409 VN.n10 VN.n9 27.0217
R1410 VN.n3 VN.n2 21.1793
R1411 VN.n9 VN.n8 21.1793
R1412 VN.n2 VN.n1 20.1275
R1413 VN.n8 VN.n7 20.1275
R1414 VN.n11 VN.n6 0.189894
R1415 VN.n5 VN.n0 0.189894
R1416 VN VN.n5 0.0516364
R1417 VDD2.n1 VDD2.t2 62.4728
R1418 VDD2.n2 VDD2.t1 61.8558
R1419 VDD2.n1 VDD2.n0 60.8706
R1420 VDD2 VDD2.n3 60.8678
R1421 VDD2.n2 VDD2.n1 41.4222
R1422 VDD2.n3 VDD2.t4 1.15435
R1423 VDD2.n3 VDD2.t5 1.15435
R1424 VDD2.n0 VDD2.t0 1.15435
R1425 VDD2.n0 VDD2.t3 1.15435
R1426 VDD2 VDD2.n2 0.731103
R1427 VTAIL.n7 VTAIL.t7 45.1771
R1428 VTAIL.n11 VTAIL.t8 45.1769
R1429 VTAIL.n2 VTAIL.t4 45.1769
R1430 VTAIL.n10 VTAIL.t0 45.1769
R1431 VTAIL.n9 VTAIL.n8 44.0233
R1432 VTAIL.n6 VTAIL.n5 44.0233
R1433 VTAIL.n1 VTAIL.n0 44.023
R1434 VTAIL.n4 VTAIL.n3 44.023
R1435 VTAIL.n6 VTAIL.n4 28.9531
R1436 VTAIL.n11 VTAIL.n10 28.0565
R1437 VTAIL.n0 VTAIL.t6 1.15435
R1438 VTAIL.n0 VTAIL.t11 1.15435
R1439 VTAIL.n3 VTAIL.t2 1.15435
R1440 VTAIL.n3 VTAIL.t3 1.15435
R1441 VTAIL.n8 VTAIL.t1 1.15435
R1442 VTAIL.n8 VTAIL.t5 1.15435
R1443 VTAIL.n5 VTAIL.t10 1.15435
R1444 VTAIL.n5 VTAIL.t9 1.15435
R1445 VTAIL.n9 VTAIL.n7 0.918603
R1446 VTAIL.n2 VTAIL.n1 0.918603
R1447 VTAIL.n7 VTAIL.n6 0.897052
R1448 VTAIL.n10 VTAIL.n9 0.897052
R1449 VTAIL.n4 VTAIL.n2 0.897052
R1450 VTAIL VTAIL.n11 0.614724
R1451 VTAIL VTAIL.n1 0.282828
R1452 VP.n3 VP.t4 659.592
R1453 VP.n8 VP.t5 637.802
R1454 VP.n12 VP.t3 637.802
R1455 VP.n14 VP.t2 637.802
R1456 VP.n6 VP.t0 637.802
R1457 VP.n4 VP.t1 637.802
R1458 VP.n15 VP.n14 161.3
R1459 VP.n5 VP.n2 161.3
R1460 VP.n7 VP.n6 161.3
R1461 VP.n13 VP.n0 161.3
R1462 VP.n12 VP.n11 161.3
R1463 VP.n10 VP.n1 161.3
R1464 VP.n9 VP.n8 161.3
R1465 VP.n9 VP.n7 45.1596
R1466 VP.n3 VP.n2 44.8565
R1467 VP.n8 VP.n1 27.0217
R1468 VP.n14 VP.n13 27.0217
R1469 VP.n6 VP.n5 27.0217
R1470 VP.n12 VP.n1 21.1793
R1471 VP.n13 VP.n12 21.1793
R1472 VP.n5 VP.n4 21.1793
R1473 VP.n4 VP.n3 20.1275
R1474 VP.n7 VP.n2 0.189894
R1475 VP.n10 VP.n9 0.189894
R1476 VP.n11 VP.n10 0.189894
R1477 VP.n11 VP.n0 0.189894
R1478 VP.n15 VP.n0 0.189894
R1479 VP VP.n15 0.0516364
R1480 VDD1 VDD1.t1 62.5865
R1481 VDD1.n1 VDD1.t0 62.4728
R1482 VDD1.n1 VDD1.n0 60.8706
R1483 VDD1.n3 VDD1.n2 60.7019
R1484 VDD1.n3 VDD1.n1 42.4535
R1485 VDD1.n2 VDD1.t4 1.15435
R1486 VDD1.n2 VDD1.t5 1.15435
R1487 VDD1.n0 VDD1.t2 1.15435
R1488 VDD1.n0 VDD1.t3 1.15435
R1489 VDD1 VDD1.n3 0.166448
C0 VDD1 VTAIL 13.3213f
C1 VDD2 VTAIL 13.3527f
C2 VTAIL VN 5.5892f
C3 VDD1 VP 6.25171f
C4 VDD2 VP 0.299377f
C5 VP VN 6.04401f
C6 VDD2 VDD1 0.714428f
C7 VDD1 VN 0.148281f
C8 VDD2 VN 6.1069f
C9 VP VTAIL 5.60402f
C10 VDD2 B 5.423726f
C11 VDD1 B 5.660459f
C12 VTAIL B 8.289088f
C13 VN B 8.38039f
C14 VP B 6.145907f
C15 VDD1.t1 B 3.68605f
C16 VDD1.t0 B 3.68538f
C17 VDD1.t2 B 0.316968f
C18 VDD1.t3 B 0.316968f
C19 VDD1.n0 B 2.88259f
C20 VDD1.n1 B 2.32864f
C21 VDD1.t4 B 0.316968f
C22 VDD1.t5 B 0.316968f
C23 VDD1.n2 B 2.88179f
C24 VDD1.n3 B 2.48184f
C25 VP.n0 B 0.046052f
C26 VP.n1 B 0.01045f
C27 VP.n2 B 0.191508f
C28 VP.t0 B 1.59166f
C29 VP.t1 B 1.59166f
C30 VP.t4 B 1.61159f
C31 VP.n3 B 0.587998f
C32 VP.n4 B 0.607271f
C33 VP.n5 B 0.01045f
C34 VP.n6 B 0.600418f
C35 VP.n7 B 2.13906f
C36 VP.t5 B 1.59166f
C37 VP.n8 B 0.600418f
C38 VP.n9 B 2.17582f
C39 VP.n10 B 0.046052f
C40 VP.n11 B 0.046052f
C41 VP.t3 B 1.59166f
C42 VP.n12 B 0.6034f
C43 VP.n13 B 0.01045f
C44 VP.t2 B 1.59166f
C45 VP.n14 B 0.600418f
C46 VP.n15 B 0.035689f
C47 VTAIL.t6 B 0.322136f
C48 VTAIL.t11 B 0.322136f
C49 VTAIL.n0 B 2.85592f
C50 VTAIL.n1 B 0.329298f
C51 VTAIL.t4 B 3.64731f
C52 VTAIL.n2 B 0.463478f
C53 VTAIL.t2 B 0.322136f
C54 VTAIL.t3 B 0.322136f
C55 VTAIL.n3 B 2.85592f
C56 VTAIL.n4 B 1.89834f
C57 VTAIL.t10 B 0.322136f
C58 VTAIL.t9 B 0.322136f
C59 VTAIL.n5 B 2.85592f
C60 VTAIL.n6 B 1.89834f
C61 VTAIL.t7 B 3.64733f
C62 VTAIL.n7 B 0.463456f
C63 VTAIL.t1 B 0.322136f
C64 VTAIL.t5 B 0.322136f
C65 VTAIL.n8 B 2.85592f
C66 VTAIL.n9 B 0.376311f
C67 VTAIL.t0 B 3.64731f
C68 VTAIL.n10 B 1.91688f
C69 VTAIL.t8 B 3.64731f
C70 VTAIL.n11 B 1.89527f
C71 VDD2.t2 B 3.6828f
C72 VDD2.t0 B 0.316746f
C73 VDD2.t3 B 0.316746f
C74 VDD2.n0 B 2.88057f
C75 VDD2.n1 B 2.25342f
C76 VDD2.t1 B 3.67971f
C77 VDD2.n2 B 2.50634f
C78 VDD2.t4 B 0.316746f
C79 VDD2.t5 B 0.316746f
C80 VDD2.n3 B 2.88054f
C81 VN.n0 B 0.188686f
C82 VN.t5 B 1.58784f
C83 VN.n1 B 0.579333f
C84 VN.t0 B 1.5682f
C85 VN.n2 B 0.598321f
C86 VN.n3 B 0.010296f
C87 VN.t3 B 1.5682f
C88 VN.n4 B 0.59157f
C89 VN.n5 B 0.035163f
C90 VN.n6 B 0.188686f
C91 VN.t4 B 1.58784f
C92 VN.n7 B 0.579333f
C93 VN.t2 B 1.5682f
C94 VN.n8 B 0.598321f
C95 VN.n9 B 0.010296f
C96 VN.t1 B 1.5682f
C97 VN.n10 B 0.59157f
C98 VN.n11 B 2.1372f
.ends

