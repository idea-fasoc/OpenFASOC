* NGSPICE file created from diff_pair_sample_1283.ext - technology: sky130A

.subckt diff_pair_sample_1283 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=5.1675 pd=27.28 as=0 ps=0 w=13.25 l=1.1
X1 VTAIL.t14 VN.t0 VDD2.t5 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=2.18625 ps=13.58 w=13.25 l=1.1
X2 VDD1.t7 VP.t0 VTAIL.t6 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=5.1675 ps=27.28 w=13.25 l=1.1
X3 VTAIL.t4 VP.t1 VDD1.t6 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=5.1675 pd=27.28 as=2.18625 ps=13.58 w=13.25 l=1.1
X4 B.t8 B.t6 B.t7 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=5.1675 pd=27.28 as=0 ps=0 w=13.25 l=1.1
X5 B.t5 B.t3 B.t4 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=5.1675 pd=27.28 as=0 ps=0 w=13.25 l=1.1
X6 VDD1.t5 VP.t2 VTAIL.t15 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=5.1675 ps=27.28 w=13.25 l=1.1
X7 VDD2.t6 VN.t1 VTAIL.t13 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=2.18625 ps=13.58 w=13.25 l=1.1
X8 VDD2.t3 VN.t2 VTAIL.t12 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=5.1675 ps=27.28 w=13.25 l=1.1
X9 VTAIL.t11 VN.t3 VDD2.t4 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=5.1675 pd=27.28 as=2.18625 ps=13.58 w=13.25 l=1.1
X10 VTAIL.t5 VP.t3 VDD1.t4 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=2.18625 ps=13.58 w=13.25 l=1.1
X11 VTAIL.t10 VN.t4 VDD2.t2 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=2.18625 ps=13.58 w=13.25 l=1.1
X12 B.t2 B.t0 B.t1 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=5.1675 pd=27.28 as=0 ps=0 w=13.25 l=1.1
X13 VTAIL.t0 VP.t4 VDD1.t3 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=2.18625 ps=13.58 w=13.25 l=1.1
X14 VDD2.t1 VN.t5 VTAIL.t9 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=2.18625 ps=13.58 w=13.25 l=1.1
X15 VDD1.t2 VP.t5 VTAIL.t2 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=2.18625 ps=13.58 w=13.25 l=1.1
X16 VTAIL.t3 VP.t6 VDD1.t1 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=5.1675 pd=27.28 as=2.18625 ps=13.58 w=13.25 l=1.1
X17 VDD2.t0 VN.t6 VTAIL.t8 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=5.1675 ps=27.28 w=13.25 l=1.1
X18 VDD1.t0 VP.t7 VTAIL.t1 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=2.18625 pd=13.58 as=2.18625 ps=13.58 w=13.25 l=1.1
X19 VTAIL.t7 VN.t7 VDD2.t7 w_n2400_n3618# sky130_fd_pr__pfet_01v8 ad=5.1675 pd=27.28 as=2.18625 ps=13.58 w=13.25 l=1.1
R0 B.n452 B.n451 585
R1 B.n453 B.n70 585
R2 B.n455 B.n454 585
R3 B.n456 B.n69 585
R4 B.n458 B.n457 585
R5 B.n459 B.n68 585
R6 B.n461 B.n460 585
R7 B.n462 B.n67 585
R8 B.n464 B.n463 585
R9 B.n465 B.n66 585
R10 B.n467 B.n466 585
R11 B.n468 B.n65 585
R12 B.n470 B.n469 585
R13 B.n471 B.n64 585
R14 B.n473 B.n472 585
R15 B.n474 B.n63 585
R16 B.n476 B.n475 585
R17 B.n477 B.n62 585
R18 B.n479 B.n478 585
R19 B.n480 B.n61 585
R20 B.n482 B.n481 585
R21 B.n483 B.n60 585
R22 B.n485 B.n484 585
R23 B.n486 B.n59 585
R24 B.n488 B.n487 585
R25 B.n489 B.n58 585
R26 B.n491 B.n490 585
R27 B.n492 B.n57 585
R28 B.n494 B.n493 585
R29 B.n495 B.n56 585
R30 B.n497 B.n496 585
R31 B.n498 B.n55 585
R32 B.n500 B.n499 585
R33 B.n501 B.n54 585
R34 B.n503 B.n502 585
R35 B.n504 B.n53 585
R36 B.n506 B.n505 585
R37 B.n507 B.n52 585
R38 B.n509 B.n508 585
R39 B.n510 B.n51 585
R40 B.n512 B.n511 585
R41 B.n513 B.n50 585
R42 B.n515 B.n514 585
R43 B.n516 B.n49 585
R44 B.n518 B.n517 585
R45 B.n520 B.n519 585
R46 B.n521 B.n45 585
R47 B.n523 B.n522 585
R48 B.n524 B.n44 585
R49 B.n526 B.n525 585
R50 B.n527 B.n43 585
R51 B.n529 B.n528 585
R52 B.n530 B.n42 585
R53 B.n532 B.n531 585
R54 B.n533 B.n39 585
R55 B.n536 B.n535 585
R56 B.n537 B.n38 585
R57 B.n539 B.n538 585
R58 B.n540 B.n37 585
R59 B.n542 B.n541 585
R60 B.n543 B.n36 585
R61 B.n545 B.n544 585
R62 B.n546 B.n35 585
R63 B.n548 B.n547 585
R64 B.n549 B.n34 585
R65 B.n551 B.n550 585
R66 B.n552 B.n33 585
R67 B.n554 B.n553 585
R68 B.n555 B.n32 585
R69 B.n557 B.n556 585
R70 B.n558 B.n31 585
R71 B.n560 B.n559 585
R72 B.n561 B.n30 585
R73 B.n563 B.n562 585
R74 B.n564 B.n29 585
R75 B.n566 B.n565 585
R76 B.n567 B.n28 585
R77 B.n569 B.n568 585
R78 B.n570 B.n27 585
R79 B.n572 B.n571 585
R80 B.n573 B.n26 585
R81 B.n575 B.n574 585
R82 B.n576 B.n25 585
R83 B.n578 B.n577 585
R84 B.n579 B.n24 585
R85 B.n581 B.n580 585
R86 B.n582 B.n23 585
R87 B.n584 B.n583 585
R88 B.n585 B.n22 585
R89 B.n587 B.n586 585
R90 B.n588 B.n21 585
R91 B.n590 B.n589 585
R92 B.n591 B.n20 585
R93 B.n593 B.n592 585
R94 B.n594 B.n19 585
R95 B.n596 B.n595 585
R96 B.n597 B.n18 585
R97 B.n599 B.n598 585
R98 B.n600 B.n17 585
R99 B.n602 B.n601 585
R100 B.n450 B.n71 585
R101 B.n449 B.n448 585
R102 B.n447 B.n72 585
R103 B.n446 B.n445 585
R104 B.n444 B.n73 585
R105 B.n443 B.n442 585
R106 B.n441 B.n74 585
R107 B.n440 B.n439 585
R108 B.n438 B.n75 585
R109 B.n437 B.n436 585
R110 B.n435 B.n76 585
R111 B.n434 B.n433 585
R112 B.n432 B.n77 585
R113 B.n431 B.n430 585
R114 B.n429 B.n78 585
R115 B.n428 B.n427 585
R116 B.n426 B.n79 585
R117 B.n425 B.n424 585
R118 B.n423 B.n80 585
R119 B.n422 B.n421 585
R120 B.n420 B.n81 585
R121 B.n419 B.n418 585
R122 B.n417 B.n82 585
R123 B.n416 B.n415 585
R124 B.n414 B.n83 585
R125 B.n413 B.n412 585
R126 B.n411 B.n84 585
R127 B.n410 B.n409 585
R128 B.n408 B.n85 585
R129 B.n407 B.n406 585
R130 B.n405 B.n86 585
R131 B.n404 B.n403 585
R132 B.n402 B.n87 585
R133 B.n401 B.n400 585
R134 B.n399 B.n88 585
R135 B.n398 B.n397 585
R136 B.n396 B.n89 585
R137 B.n395 B.n394 585
R138 B.n393 B.n90 585
R139 B.n392 B.n391 585
R140 B.n390 B.n91 585
R141 B.n389 B.n388 585
R142 B.n387 B.n92 585
R143 B.n386 B.n385 585
R144 B.n384 B.n93 585
R145 B.n383 B.n382 585
R146 B.n381 B.n94 585
R147 B.n380 B.n379 585
R148 B.n378 B.n95 585
R149 B.n377 B.n376 585
R150 B.n375 B.n96 585
R151 B.n374 B.n373 585
R152 B.n372 B.n97 585
R153 B.n371 B.n370 585
R154 B.n369 B.n98 585
R155 B.n368 B.n367 585
R156 B.n366 B.n99 585
R157 B.n365 B.n364 585
R158 B.n363 B.n100 585
R159 B.n212 B.n211 585
R160 B.n213 B.n154 585
R161 B.n215 B.n214 585
R162 B.n216 B.n153 585
R163 B.n218 B.n217 585
R164 B.n219 B.n152 585
R165 B.n221 B.n220 585
R166 B.n222 B.n151 585
R167 B.n224 B.n223 585
R168 B.n225 B.n150 585
R169 B.n227 B.n226 585
R170 B.n228 B.n149 585
R171 B.n230 B.n229 585
R172 B.n231 B.n148 585
R173 B.n233 B.n232 585
R174 B.n234 B.n147 585
R175 B.n236 B.n235 585
R176 B.n237 B.n146 585
R177 B.n239 B.n238 585
R178 B.n240 B.n145 585
R179 B.n242 B.n241 585
R180 B.n243 B.n144 585
R181 B.n245 B.n244 585
R182 B.n246 B.n143 585
R183 B.n248 B.n247 585
R184 B.n249 B.n142 585
R185 B.n251 B.n250 585
R186 B.n252 B.n141 585
R187 B.n254 B.n253 585
R188 B.n255 B.n140 585
R189 B.n257 B.n256 585
R190 B.n258 B.n139 585
R191 B.n260 B.n259 585
R192 B.n261 B.n138 585
R193 B.n263 B.n262 585
R194 B.n264 B.n137 585
R195 B.n266 B.n265 585
R196 B.n267 B.n136 585
R197 B.n269 B.n268 585
R198 B.n270 B.n135 585
R199 B.n272 B.n271 585
R200 B.n273 B.n134 585
R201 B.n275 B.n274 585
R202 B.n276 B.n133 585
R203 B.n278 B.n277 585
R204 B.n280 B.n279 585
R205 B.n281 B.n129 585
R206 B.n283 B.n282 585
R207 B.n284 B.n128 585
R208 B.n286 B.n285 585
R209 B.n287 B.n127 585
R210 B.n289 B.n288 585
R211 B.n290 B.n126 585
R212 B.n292 B.n291 585
R213 B.n293 B.n123 585
R214 B.n296 B.n295 585
R215 B.n297 B.n122 585
R216 B.n299 B.n298 585
R217 B.n300 B.n121 585
R218 B.n302 B.n301 585
R219 B.n303 B.n120 585
R220 B.n305 B.n304 585
R221 B.n306 B.n119 585
R222 B.n308 B.n307 585
R223 B.n309 B.n118 585
R224 B.n311 B.n310 585
R225 B.n312 B.n117 585
R226 B.n314 B.n313 585
R227 B.n315 B.n116 585
R228 B.n317 B.n316 585
R229 B.n318 B.n115 585
R230 B.n320 B.n319 585
R231 B.n321 B.n114 585
R232 B.n323 B.n322 585
R233 B.n324 B.n113 585
R234 B.n326 B.n325 585
R235 B.n327 B.n112 585
R236 B.n329 B.n328 585
R237 B.n330 B.n111 585
R238 B.n332 B.n331 585
R239 B.n333 B.n110 585
R240 B.n335 B.n334 585
R241 B.n336 B.n109 585
R242 B.n338 B.n337 585
R243 B.n339 B.n108 585
R244 B.n341 B.n340 585
R245 B.n342 B.n107 585
R246 B.n344 B.n343 585
R247 B.n345 B.n106 585
R248 B.n347 B.n346 585
R249 B.n348 B.n105 585
R250 B.n350 B.n349 585
R251 B.n351 B.n104 585
R252 B.n353 B.n352 585
R253 B.n354 B.n103 585
R254 B.n356 B.n355 585
R255 B.n357 B.n102 585
R256 B.n359 B.n358 585
R257 B.n360 B.n101 585
R258 B.n362 B.n361 585
R259 B.n210 B.n155 585
R260 B.n209 B.n208 585
R261 B.n207 B.n156 585
R262 B.n206 B.n205 585
R263 B.n204 B.n157 585
R264 B.n203 B.n202 585
R265 B.n201 B.n158 585
R266 B.n200 B.n199 585
R267 B.n198 B.n159 585
R268 B.n197 B.n196 585
R269 B.n195 B.n160 585
R270 B.n194 B.n193 585
R271 B.n192 B.n161 585
R272 B.n191 B.n190 585
R273 B.n189 B.n162 585
R274 B.n188 B.n187 585
R275 B.n186 B.n163 585
R276 B.n185 B.n184 585
R277 B.n183 B.n164 585
R278 B.n182 B.n181 585
R279 B.n180 B.n165 585
R280 B.n179 B.n178 585
R281 B.n177 B.n166 585
R282 B.n176 B.n175 585
R283 B.n174 B.n167 585
R284 B.n173 B.n172 585
R285 B.n171 B.n168 585
R286 B.n170 B.n169 585
R287 B.n2 B.n0 585
R288 B.n645 B.n1 585
R289 B.n644 B.n643 585
R290 B.n642 B.n3 585
R291 B.n641 B.n640 585
R292 B.n639 B.n4 585
R293 B.n638 B.n637 585
R294 B.n636 B.n5 585
R295 B.n635 B.n634 585
R296 B.n633 B.n6 585
R297 B.n632 B.n631 585
R298 B.n630 B.n7 585
R299 B.n629 B.n628 585
R300 B.n627 B.n8 585
R301 B.n626 B.n625 585
R302 B.n624 B.n9 585
R303 B.n623 B.n622 585
R304 B.n621 B.n10 585
R305 B.n620 B.n619 585
R306 B.n618 B.n11 585
R307 B.n617 B.n616 585
R308 B.n615 B.n12 585
R309 B.n614 B.n613 585
R310 B.n612 B.n13 585
R311 B.n611 B.n610 585
R312 B.n609 B.n14 585
R313 B.n608 B.n607 585
R314 B.n606 B.n15 585
R315 B.n605 B.n604 585
R316 B.n603 B.n16 585
R317 B.n647 B.n646 585
R318 B.n212 B.n155 535.745
R319 B.n603 B.n602 535.745
R320 B.n363 B.n362 535.745
R321 B.n452 B.n71 535.745
R322 B.n124 B.t6 493.856
R323 B.n130 B.t0 493.856
R324 B.n40 B.t3 493.856
R325 B.n46 B.t9 493.856
R326 B.n208 B.n155 163.367
R327 B.n208 B.n207 163.367
R328 B.n207 B.n206 163.367
R329 B.n206 B.n157 163.367
R330 B.n202 B.n157 163.367
R331 B.n202 B.n201 163.367
R332 B.n201 B.n200 163.367
R333 B.n200 B.n159 163.367
R334 B.n196 B.n159 163.367
R335 B.n196 B.n195 163.367
R336 B.n195 B.n194 163.367
R337 B.n194 B.n161 163.367
R338 B.n190 B.n161 163.367
R339 B.n190 B.n189 163.367
R340 B.n189 B.n188 163.367
R341 B.n188 B.n163 163.367
R342 B.n184 B.n163 163.367
R343 B.n184 B.n183 163.367
R344 B.n183 B.n182 163.367
R345 B.n182 B.n165 163.367
R346 B.n178 B.n165 163.367
R347 B.n178 B.n177 163.367
R348 B.n177 B.n176 163.367
R349 B.n176 B.n167 163.367
R350 B.n172 B.n167 163.367
R351 B.n172 B.n171 163.367
R352 B.n171 B.n170 163.367
R353 B.n170 B.n2 163.367
R354 B.n646 B.n2 163.367
R355 B.n646 B.n645 163.367
R356 B.n645 B.n644 163.367
R357 B.n644 B.n3 163.367
R358 B.n640 B.n3 163.367
R359 B.n640 B.n639 163.367
R360 B.n639 B.n638 163.367
R361 B.n638 B.n5 163.367
R362 B.n634 B.n5 163.367
R363 B.n634 B.n633 163.367
R364 B.n633 B.n632 163.367
R365 B.n632 B.n7 163.367
R366 B.n628 B.n7 163.367
R367 B.n628 B.n627 163.367
R368 B.n627 B.n626 163.367
R369 B.n626 B.n9 163.367
R370 B.n622 B.n9 163.367
R371 B.n622 B.n621 163.367
R372 B.n621 B.n620 163.367
R373 B.n620 B.n11 163.367
R374 B.n616 B.n11 163.367
R375 B.n616 B.n615 163.367
R376 B.n615 B.n614 163.367
R377 B.n614 B.n13 163.367
R378 B.n610 B.n13 163.367
R379 B.n610 B.n609 163.367
R380 B.n609 B.n608 163.367
R381 B.n608 B.n15 163.367
R382 B.n604 B.n15 163.367
R383 B.n604 B.n603 163.367
R384 B.n213 B.n212 163.367
R385 B.n214 B.n213 163.367
R386 B.n214 B.n153 163.367
R387 B.n218 B.n153 163.367
R388 B.n219 B.n218 163.367
R389 B.n220 B.n219 163.367
R390 B.n220 B.n151 163.367
R391 B.n224 B.n151 163.367
R392 B.n225 B.n224 163.367
R393 B.n226 B.n225 163.367
R394 B.n226 B.n149 163.367
R395 B.n230 B.n149 163.367
R396 B.n231 B.n230 163.367
R397 B.n232 B.n231 163.367
R398 B.n232 B.n147 163.367
R399 B.n236 B.n147 163.367
R400 B.n237 B.n236 163.367
R401 B.n238 B.n237 163.367
R402 B.n238 B.n145 163.367
R403 B.n242 B.n145 163.367
R404 B.n243 B.n242 163.367
R405 B.n244 B.n243 163.367
R406 B.n244 B.n143 163.367
R407 B.n248 B.n143 163.367
R408 B.n249 B.n248 163.367
R409 B.n250 B.n249 163.367
R410 B.n250 B.n141 163.367
R411 B.n254 B.n141 163.367
R412 B.n255 B.n254 163.367
R413 B.n256 B.n255 163.367
R414 B.n256 B.n139 163.367
R415 B.n260 B.n139 163.367
R416 B.n261 B.n260 163.367
R417 B.n262 B.n261 163.367
R418 B.n262 B.n137 163.367
R419 B.n266 B.n137 163.367
R420 B.n267 B.n266 163.367
R421 B.n268 B.n267 163.367
R422 B.n268 B.n135 163.367
R423 B.n272 B.n135 163.367
R424 B.n273 B.n272 163.367
R425 B.n274 B.n273 163.367
R426 B.n274 B.n133 163.367
R427 B.n278 B.n133 163.367
R428 B.n279 B.n278 163.367
R429 B.n279 B.n129 163.367
R430 B.n283 B.n129 163.367
R431 B.n284 B.n283 163.367
R432 B.n285 B.n284 163.367
R433 B.n285 B.n127 163.367
R434 B.n289 B.n127 163.367
R435 B.n290 B.n289 163.367
R436 B.n291 B.n290 163.367
R437 B.n291 B.n123 163.367
R438 B.n296 B.n123 163.367
R439 B.n297 B.n296 163.367
R440 B.n298 B.n297 163.367
R441 B.n298 B.n121 163.367
R442 B.n302 B.n121 163.367
R443 B.n303 B.n302 163.367
R444 B.n304 B.n303 163.367
R445 B.n304 B.n119 163.367
R446 B.n308 B.n119 163.367
R447 B.n309 B.n308 163.367
R448 B.n310 B.n309 163.367
R449 B.n310 B.n117 163.367
R450 B.n314 B.n117 163.367
R451 B.n315 B.n314 163.367
R452 B.n316 B.n315 163.367
R453 B.n316 B.n115 163.367
R454 B.n320 B.n115 163.367
R455 B.n321 B.n320 163.367
R456 B.n322 B.n321 163.367
R457 B.n322 B.n113 163.367
R458 B.n326 B.n113 163.367
R459 B.n327 B.n326 163.367
R460 B.n328 B.n327 163.367
R461 B.n328 B.n111 163.367
R462 B.n332 B.n111 163.367
R463 B.n333 B.n332 163.367
R464 B.n334 B.n333 163.367
R465 B.n334 B.n109 163.367
R466 B.n338 B.n109 163.367
R467 B.n339 B.n338 163.367
R468 B.n340 B.n339 163.367
R469 B.n340 B.n107 163.367
R470 B.n344 B.n107 163.367
R471 B.n345 B.n344 163.367
R472 B.n346 B.n345 163.367
R473 B.n346 B.n105 163.367
R474 B.n350 B.n105 163.367
R475 B.n351 B.n350 163.367
R476 B.n352 B.n351 163.367
R477 B.n352 B.n103 163.367
R478 B.n356 B.n103 163.367
R479 B.n357 B.n356 163.367
R480 B.n358 B.n357 163.367
R481 B.n358 B.n101 163.367
R482 B.n362 B.n101 163.367
R483 B.n364 B.n363 163.367
R484 B.n364 B.n99 163.367
R485 B.n368 B.n99 163.367
R486 B.n369 B.n368 163.367
R487 B.n370 B.n369 163.367
R488 B.n370 B.n97 163.367
R489 B.n374 B.n97 163.367
R490 B.n375 B.n374 163.367
R491 B.n376 B.n375 163.367
R492 B.n376 B.n95 163.367
R493 B.n380 B.n95 163.367
R494 B.n381 B.n380 163.367
R495 B.n382 B.n381 163.367
R496 B.n382 B.n93 163.367
R497 B.n386 B.n93 163.367
R498 B.n387 B.n386 163.367
R499 B.n388 B.n387 163.367
R500 B.n388 B.n91 163.367
R501 B.n392 B.n91 163.367
R502 B.n393 B.n392 163.367
R503 B.n394 B.n393 163.367
R504 B.n394 B.n89 163.367
R505 B.n398 B.n89 163.367
R506 B.n399 B.n398 163.367
R507 B.n400 B.n399 163.367
R508 B.n400 B.n87 163.367
R509 B.n404 B.n87 163.367
R510 B.n405 B.n404 163.367
R511 B.n406 B.n405 163.367
R512 B.n406 B.n85 163.367
R513 B.n410 B.n85 163.367
R514 B.n411 B.n410 163.367
R515 B.n412 B.n411 163.367
R516 B.n412 B.n83 163.367
R517 B.n416 B.n83 163.367
R518 B.n417 B.n416 163.367
R519 B.n418 B.n417 163.367
R520 B.n418 B.n81 163.367
R521 B.n422 B.n81 163.367
R522 B.n423 B.n422 163.367
R523 B.n424 B.n423 163.367
R524 B.n424 B.n79 163.367
R525 B.n428 B.n79 163.367
R526 B.n429 B.n428 163.367
R527 B.n430 B.n429 163.367
R528 B.n430 B.n77 163.367
R529 B.n434 B.n77 163.367
R530 B.n435 B.n434 163.367
R531 B.n436 B.n435 163.367
R532 B.n436 B.n75 163.367
R533 B.n440 B.n75 163.367
R534 B.n441 B.n440 163.367
R535 B.n442 B.n441 163.367
R536 B.n442 B.n73 163.367
R537 B.n446 B.n73 163.367
R538 B.n447 B.n446 163.367
R539 B.n448 B.n447 163.367
R540 B.n448 B.n71 163.367
R541 B.n602 B.n17 163.367
R542 B.n598 B.n17 163.367
R543 B.n598 B.n597 163.367
R544 B.n597 B.n596 163.367
R545 B.n596 B.n19 163.367
R546 B.n592 B.n19 163.367
R547 B.n592 B.n591 163.367
R548 B.n591 B.n590 163.367
R549 B.n590 B.n21 163.367
R550 B.n586 B.n21 163.367
R551 B.n586 B.n585 163.367
R552 B.n585 B.n584 163.367
R553 B.n584 B.n23 163.367
R554 B.n580 B.n23 163.367
R555 B.n580 B.n579 163.367
R556 B.n579 B.n578 163.367
R557 B.n578 B.n25 163.367
R558 B.n574 B.n25 163.367
R559 B.n574 B.n573 163.367
R560 B.n573 B.n572 163.367
R561 B.n572 B.n27 163.367
R562 B.n568 B.n27 163.367
R563 B.n568 B.n567 163.367
R564 B.n567 B.n566 163.367
R565 B.n566 B.n29 163.367
R566 B.n562 B.n29 163.367
R567 B.n562 B.n561 163.367
R568 B.n561 B.n560 163.367
R569 B.n560 B.n31 163.367
R570 B.n556 B.n31 163.367
R571 B.n556 B.n555 163.367
R572 B.n555 B.n554 163.367
R573 B.n554 B.n33 163.367
R574 B.n550 B.n33 163.367
R575 B.n550 B.n549 163.367
R576 B.n549 B.n548 163.367
R577 B.n548 B.n35 163.367
R578 B.n544 B.n35 163.367
R579 B.n544 B.n543 163.367
R580 B.n543 B.n542 163.367
R581 B.n542 B.n37 163.367
R582 B.n538 B.n37 163.367
R583 B.n538 B.n537 163.367
R584 B.n537 B.n536 163.367
R585 B.n536 B.n39 163.367
R586 B.n531 B.n39 163.367
R587 B.n531 B.n530 163.367
R588 B.n530 B.n529 163.367
R589 B.n529 B.n43 163.367
R590 B.n525 B.n43 163.367
R591 B.n525 B.n524 163.367
R592 B.n524 B.n523 163.367
R593 B.n523 B.n45 163.367
R594 B.n519 B.n45 163.367
R595 B.n519 B.n518 163.367
R596 B.n518 B.n49 163.367
R597 B.n514 B.n49 163.367
R598 B.n514 B.n513 163.367
R599 B.n513 B.n512 163.367
R600 B.n512 B.n51 163.367
R601 B.n508 B.n51 163.367
R602 B.n508 B.n507 163.367
R603 B.n507 B.n506 163.367
R604 B.n506 B.n53 163.367
R605 B.n502 B.n53 163.367
R606 B.n502 B.n501 163.367
R607 B.n501 B.n500 163.367
R608 B.n500 B.n55 163.367
R609 B.n496 B.n55 163.367
R610 B.n496 B.n495 163.367
R611 B.n495 B.n494 163.367
R612 B.n494 B.n57 163.367
R613 B.n490 B.n57 163.367
R614 B.n490 B.n489 163.367
R615 B.n489 B.n488 163.367
R616 B.n488 B.n59 163.367
R617 B.n484 B.n59 163.367
R618 B.n484 B.n483 163.367
R619 B.n483 B.n482 163.367
R620 B.n482 B.n61 163.367
R621 B.n478 B.n61 163.367
R622 B.n478 B.n477 163.367
R623 B.n477 B.n476 163.367
R624 B.n476 B.n63 163.367
R625 B.n472 B.n63 163.367
R626 B.n472 B.n471 163.367
R627 B.n471 B.n470 163.367
R628 B.n470 B.n65 163.367
R629 B.n466 B.n65 163.367
R630 B.n466 B.n465 163.367
R631 B.n465 B.n464 163.367
R632 B.n464 B.n67 163.367
R633 B.n460 B.n67 163.367
R634 B.n460 B.n459 163.367
R635 B.n459 B.n458 163.367
R636 B.n458 B.n69 163.367
R637 B.n454 B.n69 163.367
R638 B.n454 B.n453 163.367
R639 B.n453 B.n452 163.367
R640 B.n124 B.t8 140.981
R641 B.n46 B.t10 140.981
R642 B.n130 B.t2 140.964
R643 B.n40 B.t4 140.964
R644 B.n125 B.t7 113.246
R645 B.n47 B.t11 113.246
R646 B.n131 B.t1 113.231
R647 B.n41 B.t5 113.231
R648 B.n294 B.n125 59.5399
R649 B.n132 B.n131 59.5399
R650 B.n534 B.n41 59.5399
R651 B.n48 B.n47 59.5399
R652 B.n601 B.n16 34.8103
R653 B.n451 B.n450 34.8103
R654 B.n361 B.n100 34.8103
R655 B.n211 B.n210 34.8103
R656 B.n125 B.n124 27.7338
R657 B.n131 B.n130 27.7338
R658 B.n41 B.n40 27.7338
R659 B.n47 B.n46 27.7338
R660 B B.n647 18.0485
R661 B.n601 B.n600 10.6151
R662 B.n600 B.n599 10.6151
R663 B.n599 B.n18 10.6151
R664 B.n595 B.n18 10.6151
R665 B.n595 B.n594 10.6151
R666 B.n594 B.n593 10.6151
R667 B.n593 B.n20 10.6151
R668 B.n589 B.n20 10.6151
R669 B.n589 B.n588 10.6151
R670 B.n588 B.n587 10.6151
R671 B.n587 B.n22 10.6151
R672 B.n583 B.n22 10.6151
R673 B.n583 B.n582 10.6151
R674 B.n582 B.n581 10.6151
R675 B.n581 B.n24 10.6151
R676 B.n577 B.n24 10.6151
R677 B.n577 B.n576 10.6151
R678 B.n576 B.n575 10.6151
R679 B.n575 B.n26 10.6151
R680 B.n571 B.n26 10.6151
R681 B.n571 B.n570 10.6151
R682 B.n570 B.n569 10.6151
R683 B.n569 B.n28 10.6151
R684 B.n565 B.n28 10.6151
R685 B.n565 B.n564 10.6151
R686 B.n564 B.n563 10.6151
R687 B.n563 B.n30 10.6151
R688 B.n559 B.n30 10.6151
R689 B.n559 B.n558 10.6151
R690 B.n558 B.n557 10.6151
R691 B.n557 B.n32 10.6151
R692 B.n553 B.n32 10.6151
R693 B.n553 B.n552 10.6151
R694 B.n552 B.n551 10.6151
R695 B.n551 B.n34 10.6151
R696 B.n547 B.n34 10.6151
R697 B.n547 B.n546 10.6151
R698 B.n546 B.n545 10.6151
R699 B.n545 B.n36 10.6151
R700 B.n541 B.n36 10.6151
R701 B.n541 B.n540 10.6151
R702 B.n540 B.n539 10.6151
R703 B.n539 B.n38 10.6151
R704 B.n535 B.n38 10.6151
R705 B.n533 B.n532 10.6151
R706 B.n532 B.n42 10.6151
R707 B.n528 B.n42 10.6151
R708 B.n528 B.n527 10.6151
R709 B.n527 B.n526 10.6151
R710 B.n526 B.n44 10.6151
R711 B.n522 B.n44 10.6151
R712 B.n522 B.n521 10.6151
R713 B.n521 B.n520 10.6151
R714 B.n517 B.n516 10.6151
R715 B.n516 B.n515 10.6151
R716 B.n515 B.n50 10.6151
R717 B.n511 B.n50 10.6151
R718 B.n511 B.n510 10.6151
R719 B.n510 B.n509 10.6151
R720 B.n509 B.n52 10.6151
R721 B.n505 B.n52 10.6151
R722 B.n505 B.n504 10.6151
R723 B.n504 B.n503 10.6151
R724 B.n503 B.n54 10.6151
R725 B.n499 B.n54 10.6151
R726 B.n499 B.n498 10.6151
R727 B.n498 B.n497 10.6151
R728 B.n497 B.n56 10.6151
R729 B.n493 B.n56 10.6151
R730 B.n493 B.n492 10.6151
R731 B.n492 B.n491 10.6151
R732 B.n491 B.n58 10.6151
R733 B.n487 B.n58 10.6151
R734 B.n487 B.n486 10.6151
R735 B.n486 B.n485 10.6151
R736 B.n485 B.n60 10.6151
R737 B.n481 B.n60 10.6151
R738 B.n481 B.n480 10.6151
R739 B.n480 B.n479 10.6151
R740 B.n479 B.n62 10.6151
R741 B.n475 B.n62 10.6151
R742 B.n475 B.n474 10.6151
R743 B.n474 B.n473 10.6151
R744 B.n473 B.n64 10.6151
R745 B.n469 B.n64 10.6151
R746 B.n469 B.n468 10.6151
R747 B.n468 B.n467 10.6151
R748 B.n467 B.n66 10.6151
R749 B.n463 B.n66 10.6151
R750 B.n463 B.n462 10.6151
R751 B.n462 B.n461 10.6151
R752 B.n461 B.n68 10.6151
R753 B.n457 B.n68 10.6151
R754 B.n457 B.n456 10.6151
R755 B.n456 B.n455 10.6151
R756 B.n455 B.n70 10.6151
R757 B.n451 B.n70 10.6151
R758 B.n365 B.n100 10.6151
R759 B.n366 B.n365 10.6151
R760 B.n367 B.n366 10.6151
R761 B.n367 B.n98 10.6151
R762 B.n371 B.n98 10.6151
R763 B.n372 B.n371 10.6151
R764 B.n373 B.n372 10.6151
R765 B.n373 B.n96 10.6151
R766 B.n377 B.n96 10.6151
R767 B.n378 B.n377 10.6151
R768 B.n379 B.n378 10.6151
R769 B.n379 B.n94 10.6151
R770 B.n383 B.n94 10.6151
R771 B.n384 B.n383 10.6151
R772 B.n385 B.n384 10.6151
R773 B.n385 B.n92 10.6151
R774 B.n389 B.n92 10.6151
R775 B.n390 B.n389 10.6151
R776 B.n391 B.n390 10.6151
R777 B.n391 B.n90 10.6151
R778 B.n395 B.n90 10.6151
R779 B.n396 B.n395 10.6151
R780 B.n397 B.n396 10.6151
R781 B.n397 B.n88 10.6151
R782 B.n401 B.n88 10.6151
R783 B.n402 B.n401 10.6151
R784 B.n403 B.n402 10.6151
R785 B.n403 B.n86 10.6151
R786 B.n407 B.n86 10.6151
R787 B.n408 B.n407 10.6151
R788 B.n409 B.n408 10.6151
R789 B.n409 B.n84 10.6151
R790 B.n413 B.n84 10.6151
R791 B.n414 B.n413 10.6151
R792 B.n415 B.n414 10.6151
R793 B.n415 B.n82 10.6151
R794 B.n419 B.n82 10.6151
R795 B.n420 B.n419 10.6151
R796 B.n421 B.n420 10.6151
R797 B.n421 B.n80 10.6151
R798 B.n425 B.n80 10.6151
R799 B.n426 B.n425 10.6151
R800 B.n427 B.n426 10.6151
R801 B.n427 B.n78 10.6151
R802 B.n431 B.n78 10.6151
R803 B.n432 B.n431 10.6151
R804 B.n433 B.n432 10.6151
R805 B.n433 B.n76 10.6151
R806 B.n437 B.n76 10.6151
R807 B.n438 B.n437 10.6151
R808 B.n439 B.n438 10.6151
R809 B.n439 B.n74 10.6151
R810 B.n443 B.n74 10.6151
R811 B.n444 B.n443 10.6151
R812 B.n445 B.n444 10.6151
R813 B.n445 B.n72 10.6151
R814 B.n449 B.n72 10.6151
R815 B.n450 B.n449 10.6151
R816 B.n211 B.n154 10.6151
R817 B.n215 B.n154 10.6151
R818 B.n216 B.n215 10.6151
R819 B.n217 B.n216 10.6151
R820 B.n217 B.n152 10.6151
R821 B.n221 B.n152 10.6151
R822 B.n222 B.n221 10.6151
R823 B.n223 B.n222 10.6151
R824 B.n223 B.n150 10.6151
R825 B.n227 B.n150 10.6151
R826 B.n228 B.n227 10.6151
R827 B.n229 B.n228 10.6151
R828 B.n229 B.n148 10.6151
R829 B.n233 B.n148 10.6151
R830 B.n234 B.n233 10.6151
R831 B.n235 B.n234 10.6151
R832 B.n235 B.n146 10.6151
R833 B.n239 B.n146 10.6151
R834 B.n240 B.n239 10.6151
R835 B.n241 B.n240 10.6151
R836 B.n241 B.n144 10.6151
R837 B.n245 B.n144 10.6151
R838 B.n246 B.n245 10.6151
R839 B.n247 B.n246 10.6151
R840 B.n247 B.n142 10.6151
R841 B.n251 B.n142 10.6151
R842 B.n252 B.n251 10.6151
R843 B.n253 B.n252 10.6151
R844 B.n253 B.n140 10.6151
R845 B.n257 B.n140 10.6151
R846 B.n258 B.n257 10.6151
R847 B.n259 B.n258 10.6151
R848 B.n259 B.n138 10.6151
R849 B.n263 B.n138 10.6151
R850 B.n264 B.n263 10.6151
R851 B.n265 B.n264 10.6151
R852 B.n265 B.n136 10.6151
R853 B.n269 B.n136 10.6151
R854 B.n270 B.n269 10.6151
R855 B.n271 B.n270 10.6151
R856 B.n271 B.n134 10.6151
R857 B.n275 B.n134 10.6151
R858 B.n276 B.n275 10.6151
R859 B.n277 B.n276 10.6151
R860 B.n281 B.n280 10.6151
R861 B.n282 B.n281 10.6151
R862 B.n282 B.n128 10.6151
R863 B.n286 B.n128 10.6151
R864 B.n287 B.n286 10.6151
R865 B.n288 B.n287 10.6151
R866 B.n288 B.n126 10.6151
R867 B.n292 B.n126 10.6151
R868 B.n293 B.n292 10.6151
R869 B.n295 B.n122 10.6151
R870 B.n299 B.n122 10.6151
R871 B.n300 B.n299 10.6151
R872 B.n301 B.n300 10.6151
R873 B.n301 B.n120 10.6151
R874 B.n305 B.n120 10.6151
R875 B.n306 B.n305 10.6151
R876 B.n307 B.n306 10.6151
R877 B.n307 B.n118 10.6151
R878 B.n311 B.n118 10.6151
R879 B.n312 B.n311 10.6151
R880 B.n313 B.n312 10.6151
R881 B.n313 B.n116 10.6151
R882 B.n317 B.n116 10.6151
R883 B.n318 B.n317 10.6151
R884 B.n319 B.n318 10.6151
R885 B.n319 B.n114 10.6151
R886 B.n323 B.n114 10.6151
R887 B.n324 B.n323 10.6151
R888 B.n325 B.n324 10.6151
R889 B.n325 B.n112 10.6151
R890 B.n329 B.n112 10.6151
R891 B.n330 B.n329 10.6151
R892 B.n331 B.n330 10.6151
R893 B.n331 B.n110 10.6151
R894 B.n335 B.n110 10.6151
R895 B.n336 B.n335 10.6151
R896 B.n337 B.n336 10.6151
R897 B.n337 B.n108 10.6151
R898 B.n341 B.n108 10.6151
R899 B.n342 B.n341 10.6151
R900 B.n343 B.n342 10.6151
R901 B.n343 B.n106 10.6151
R902 B.n347 B.n106 10.6151
R903 B.n348 B.n347 10.6151
R904 B.n349 B.n348 10.6151
R905 B.n349 B.n104 10.6151
R906 B.n353 B.n104 10.6151
R907 B.n354 B.n353 10.6151
R908 B.n355 B.n354 10.6151
R909 B.n355 B.n102 10.6151
R910 B.n359 B.n102 10.6151
R911 B.n360 B.n359 10.6151
R912 B.n361 B.n360 10.6151
R913 B.n210 B.n209 10.6151
R914 B.n209 B.n156 10.6151
R915 B.n205 B.n156 10.6151
R916 B.n205 B.n204 10.6151
R917 B.n204 B.n203 10.6151
R918 B.n203 B.n158 10.6151
R919 B.n199 B.n158 10.6151
R920 B.n199 B.n198 10.6151
R921 B.n198 B.n197 10.6151
R922 B.n197 B.n160 10.6151
R923 B.n193 B.n160 10.6151
R924 B.n193 B.n192 10.6151
R925 B.n192 B.n191 10.6151
R926 B.n191 B.n162 10.6151
R927 B.n187 B.n162 10.6151
R928 B.n187 B.n186 10.6151
R929 B.n186 B.n185 10.6151
R930 B.n185 B.n164 10.6151
R931 B.n181 B.n164 10.6151
R932 B.n181 B.n180 10.6151
R933 B.n180 B.n179 10.6151
R934 B.n179 B.n166 10.6151
R935 B.n175 B.n166 10.6151
R936 B.n175 B.n174 10.6151
R937 B.n174 B.n173 10.6151
R938 B.n173 B.n168 10.6151
R939 B.n169 B.n168 10.6151
R940 B.n169 B.n0 10.6151
R941 B.n643 B.n1 10.6151
R942 B.n643 B.n642 10.6151
R943 B.n642 B.n641 10.6151
R944 B.n641 B.n4 10.6151
R945 B.n637 B.n4 10.6151
R946 B.n637 B.n636 10.6151
R947 B.n636 B.n635 10.6151
R948 B.n635 B.n6 10.6151
R949 B.n631 B.n6 10.6151
R950 B.n631 B.n630 10.6151
R951 B.n630 B.n629 10.6151
R952 B.n629 B.n8 10.6151
R953 B.n625 B.n8 10.6151
R954 B.n625 B.n624 10.6151
R955 B.n624 B.n623 10.6151
R956 B.n623 B.n10 10.6151
R957 B.n619 B.n10 10.6151
R958 B.n619 B.n618 10.6151
R959 B.n618 B.n617 10.6151
R960 B.n617 B.n12 10.6151
R961 B.n613 B.n12 10.6151
R962 B.n613 B.n612 10.6151
R963 B.n612 B.n611 10.6151
R964 B.n611 B.n14 10.6151
R965 B.n607 B.n14 10.6151
R966 B.n607 B.n606 10.6151
R967 B.n606 B.n605 10.6151
R968 B.n605 B.n16 10.6151
R969 B.n535 B.n534 9.36635
R970 B.n517 B.n48 9.36635
R971 B.n277 B.n132 9.36635
R972 B.n295 B.n294 9.36635
R973 B.n647 B.n0 2.81026
R974 B.n647 B.n1 2.81026
R975 B.n534 B.n533 1.24928
R976 B.n520 B.n48 1.24928
R977 B.n280 B.n132 1.24928
R978 B.n294 B.n293 1.24928
R979 VN.n3 VN.t7 348.825
R980 VN.n16 VN.t2 348.825
R981 VN.n11 VN.t6 326.226
R982 VN.n24 VN.t3 326.226
R983 VN.n4 VN.t1 290.296
R984 VN.n1 VN.t4 290.296
R985 VN.n17 VN.t0 290.296
R986 VN.n14 VN.t5 290.296
R987 VN.n23 VN.n13 161.3
R988 VN.n22 VN.n21 161.3
R989 VN.n20 VN.n19 161.3
R990 VN.n18 VN.n15 161.3
R991 VN.n10 VN.n0 161.3
R992 VN.n9 VN.n8 161.3
R993 VN.n7 VN.n6 161.3
R994 VN.n5 VN.n2 161.3
R995 VN.n25 VN.n24 80.6037
R996 VN.n12 VN.n11 80.6037
R997 VN.n6 VN.n5 56.5193
R998 VN.n19 VN.n18 56.5193
R999 VN.n11 VN.n10 48.9345
R1000 VN.n24 VN.n23 48.9345
R1001 VN VN.n25 45.2718
R1002 VN.n4 VN.n3 33.9754
R1003 VN.n17 VN.n16 33.9754
R1004 VN.n16 VN.n15 28.3407
R1005 VN.n3 VN.n2 28.3407
R1006 VN.n10 VN.n9 24.4675
R1007 VN.n23 VN.n22 24.4675
R1008 VN.n5 VN.n4 22.7548
R1009 VN.n6 VN.n1 22.7548
R1010 VN.n18 VN.n17 22.7548
R1011 VN.n19 VN.n14 22.7548
R1012 VN.n9 VN.n1 1.71319
R1013 VN.n22 VN.n14 1.71319
R1014 VN.n25 VN.n13 0.285035
R1015 VN.n12 VN.n0 0.285035
R1016 VN.n21 VN.n13 0.189894
R1017 VN.n21 VN.n20 0.189894
R1018 VN.n20 VN.n15 0.189894
R1019 VN.n7 VN.n2 0.189894
R1020 VN.n8 VN.n7 0.189894
R1021 VN.n8 VN.n0 0.189894
R1022 VN VN.n12 0.146778
R1023 VDD2.n2 VDD2.n1 74.1654
R1024 VDD2.n2 VDD2.n0 74.1654
R1025 VDD2 VDD2.n5 74.1624
R1026 VDD2.n4 VDD2.n3 73.6044
R1027 VDD2.n4 VDD2.n2 40.6851
R1028 VDD2.n5 VDD2.t5 2.45371
R1029 VDD2.n5 VDD2.t3 2.45371
R1030 VDD2.n3 VDD2.t4 2.45371
R1031 VDD2.n3 VDD2.t1 2.45371
R1032 VDD2.n1 VDD2.t2 2.45371
R1033 VDD2.n1 VDD2.t0 2.45371
R1034 VDD2.n0 VDD2.t7 2.45371
R1035 VDD2.n0 VDD2.t6 2.45371
R1036 VDD2 VDD2.n4 0.675069
R1037 VTAIL.n11 VTAIL.t4 59.3788
R1038 VTAIL.n10 VTAIL.t12 59.3788
R1039 VTAIL.n7 VTAIL.t11 59.3788
R1040 VTAIL.n15 VTAIL.t8 59.3786
R1041 VTAIL.n2 VTAIL.t7 59.3786
R1042 VTAIL.n3 VTAIL.t15 59.3786
R1043 VTAIL.n6 VTAIL.t3 59.3786
R1044 VTAIL.n14 VTAIL.t6 59.3786
R1045 VTAIL.n13 VTAIL.n12 56.9256
R1046 VTAIL.n9 VTAIL.n8 56.9256
R1047 VTAIL.n1 VTAIL.n0 56.9255
R1048 VTAIL.n5 VTAIL.n4 56.9255
R1049 VTAIL.n15 VTAIL.n14 25.0221
R1050 VTAIL.n7 VTAIL.n6 25.0221
R1051 VTAIL.n0 VTAIL.t13 2.45371
R1052 VTAIL.n0 VTAIL.t10 2.45371
R1053 VTAIL.n4 VTAIL.t1 2.45371
R1054 VTAIL.n4 VTAIL.t0 2.45371
R1055 VTAIL.n12 VTAIL.t2 2.45371
R1056 VTAIL.n12 VTAIL.t5 2.45371
R1057 VTAIL.n8 VTAIL.t9 2.45371
R1058 VTAIL.n8 VTAIL.t14 2.45371
R1059 VTAIL.n9 VTAIL.n7 1.23326
R1060 VTAIL.n10 VTAIL.n9 1.23326
R1061 VTAIL.n13 VTAIL.n11 1.23326
R1062 VTAIL.n14 VTAIL.n13 1.23326
R1063 VTAIL.n6 VTAIL.n5 1.23326
R1064 VTAIL.n5 VTAIL.n3 1.23326
R1065 VTAIL.n2 VTAIL.n1 1.23326
R1066 VTAIL VTAIL.n15 1.17507
R1067 VTAIL.n11 VTAIL.n10 0.470328
R1068 VTAIL.n3 VTAIL.n2 0.470328
R1069 VTAIL VTAIL.n1 0.0586897
R1070 VP.n7 VP.t1 348.825
R1071 VP.n17 VP.t6 326.226
R1072 VP.n29 VP.t2 326.226
R1073 VP.n15 VP.t0 326.226
R1074 VP.n22 VP.t7 290.296
R1075 VP.n1 VP.t4 290.296
R1076 VP.n5 VP.t3 290.296
R1077 VP.n8 VP.t5 290.296
R1078 VP.n9 VP.n6 161.3
R1079 VP.n11 VP.n10 161.3
R1080 VP.n13 VP.n12 161.3
R1081 VP.n14 VP.n4 161.3
R1082 VP.n28 VP.n0 161.3
R1083 VP.n27 VP.n26 161.3
R1084 VP.n25 VP.n24 161.3
R1085 VP.n23 VP.n2 161.3
R1086 VP.n21 VP.n20 161.3
R1087 VP.n19 VP.n3 161.3
R1088 VP.n16 VP.n15 80.6037
R1089 VP.n30 VP.n29 80.6037
R1090 VP.n18 VP.n17 80.6037
R1091 VP.n24 VP.n23 56.5193
R1092 VP.n10 VP.n9 56.5193
R1093 VP.n17 VP.n3 48.9345
R1094 VP.n29 VP.n28 48.9345
R1095 VP.n15 VP.n14 48.9345
R1096 VP.n18 VP.n16 44.9862
R1097 VP.n8 VP.n7 33.9754
R1098 VP.n7 VP.n6 28.3407
R1099 VP.n21 VP.n3 24.4675
R1100 VP.n28 VP.n27 24.4675
R1101 VP.n14 VP.n13 24.4675
R1102 VP.n23 VP.n22 22.7548
R1103 VP.n24 VP.n1 22.7548
R1104 VP.n10 VP.n5 22.7548
R1105 VP.n9 VP.n8 22.7548
R1106 VP.n22 VP.n21 1.71319
R1107 VP.n27 VP.n1 1.71319
R1108 VP.n13 VP.n5 1.71319
R1109 VP.n16 VP.n4 0.285035
R1110 VP.n19 VP.n18 0.285035
R1111 VP.n30 VP.n0 0.285035
R1112 VP.n11 VP.n6 0.189894
R1113 VP.n12 VP.n11 0.189894
R1114 VP.n12 VP.n4 0.189894
R1115 VP.n20 VP.n19 0.189894
R1116 VP.n20 VP.n2 0.189894
R1117 VP.n25 VP.n2 0.189894
R1118 VP.n26 VP.n25 0.189894
R1119 VP.n26 VP.n0 0.189894
R1120 VP VP.n30 0.146778
R1121 VDD1 VDD1.n0 74.279
R1122 VDD1.n3 VDD1.n2 74.1654
R1123 VDD1.n3 VDD1.n1 74.1654
R1124 VDD1.n5 VDD1.n4 73.6042
R1125 VDD1.n5 VDD1.n3 41.2681
R1126 VDD1.n4 VDD1.t4 2.45371
R1127 VDD1.n4 VDD1.t7 2.45371
R1128 VDD1.n0 VDD1.t6 2.45371
R1129 VDD1.n0 VDD1.t2 2.45371
R1130 VDD1.n2 VDD1.t3 2.45371
R1131 VDD1.n2 VDD1.t5 2.45371
R1132 VDD1.n1 VDD1.t1 2.45371
R1133 VDD1.n1 VDD1.t0 2.45371
R1134 VDD1 VDD1.n5 0.55869
C0 VDD1 w_n2400_n3618# 1.48529f
C1 VDD2 VDD1 1.02651f
C2 VTAIL VP 7.31028f
C3 B w_n2400_n3618# 8.16989f
C4 VN VDD1 0.149072f
C5 B VDD2 1.27498f
C6 VN B 0.890067f
C7 VDD2 w_n2400_n3618# 1.53688f
C8 VDD1 VP 7.642291f
C9 VTAIL VDD1 9.95439f
C10 VN w_n2400_n3618# 4.48416f
C11 B VP 1.39696f
C12 VN VDD2 7.43189f
C13 B VTAIL 4.499701f
C14 VP w_n2400_n3618# 4.79131f
C15 VTAIL w_n2400_n3618# 4.46331f
C16 VDD2 VP 0.360111f
C17 VDD2 VTAIL 9.99875f
C18 VN VP 6.05934f
C19 B VDD1 1.22593f
C20 VN VTAIL 7.29617f
C21 VDD2 VSUBS 1.437061f
C22 VDD1 VSUBS 1.816301f
C23 VTAIL VSUBS 1.092595f
C24 VN VSUBS 5.0948f
C25 VP VSUBS 2.117257f
C26 B VSUBS 3.436909f
C27 w_n2400_n3618# VSUBS 0.106704p
C28 VDD1.t6 VSUBS 0.270129f
C29 VDD1.t2 VSUBS 0.270129f
C30 VDD1.n0 VSUBS 2.15158f
C31 VDD1.t1 VSUBS 0.270129f
C32 VDD1.t0 VSUBS 0.270129f
C33 VDD1.n1 VSUBS 2.15052f
C34 VDD1.t3 VSUBS 0.270129f
C35 VDD1.t5 VSUBS 0.270129f
C36 VDD1.n2 VSUBS 2.15052f
C37 VDD1.n3 VSUBS 3.16961f
C38 VDD1.t4 VSUBS 0.270129f
C39 VDD1.t7 VSUBS 0.270129f
C40 VDD1.n4 VSUBS 2.14559f
C41 VDD1.n5 VSUBS 2.91533f
C42 VP.n0 VSUBS 0.060002f
C43 VP.t4 VSUBS 1.79049f
C44 VP.n1 VSUBS 0.653605f
C45 VP.n2 VSUBS 0.044967f
C46 VP.t7 VSUBS 1.79049f
C47 VP.n3 VSUBS 0.053902f
C48 VP.n4 VSUBS 0.060002f
C49 VP.t0 VSUBS 1.86627f
C50 VP.t3 VSUBS 1.79049f
C51 VP.n5 VSUBS 0.653605f
C52 VP.n6 VSUBS 0.233463f
C53 VP.t5 VSUBS 1.79049f
C54 VP.t1 VSUBS 1.91426f
C55 VP.n7 VSUBS 0.713401f
C56 VP.n8 VSUBS 0.72355f
C57 VP.n9 VSUBS 0.062745f
C58 VP.n10 VSUBS 0.062745f
C59 VP.n11 VSUBS 0.044967f
C60 VP.n12 VSUBS 0.044967f
C61 VP.n13 VSUBS 0.045325f
C62 VP.n14 VSUBS 0.053902f
C63 VP.n15 VSUBS 0.729922f
C64 VP.n16 VSUBS 2.09192f
C65 VP.t6 VSUBS 1.86627f
C66 VP.n17 VSUBS 0.729922f
C67 VP.n18 VSUBS 2.12785f
C68 VP.n19 VSUBS 0.060002f
C69 VP.n20 VSUBS 0.044967f
C70 VP.n21 VSUBS 0.045325f
C71 VP.n22 VSUBS 0.653605f
C72 VP.n23 VSUBS 0.062745f
C73 VP.n24 VSUBS 0.062745f
C74 VP.n25 VSUBS 0.044967f
C75 VP.n26 VSUBS 0.044967f
C76 VP.n27 VSUBS 0.045325f
C77 VP.n28 VSUBS 0.053902f
C78 VP.t2 VSUBS 1.86627f
C79 VP.n29 VSUBS 0.729922f
C80 VP.n30 VSUBS 0.042113f
C81 VTAIL.t13 VSUBS 0.252352f
C82 VTAIL.t10 VSUBS 0.252352f
C83 VTAIL.n0 VSUBS 1.87152f
C84 VTAIL.n1 VSUBS 0.658478f
C85 VTAIL.t7 VSUBS 2.46442f
C86 VTAIL.n2 VSUBS 0.78578f
C87 VTAIL.t15 VSUBS 2.46442f
C88 VTAIL.n3 VSUBS 0.78578f
C89 VTAIL.t1 VSUBS 0.252352f
C90 VTAIL.t0 VSUBS 0.252352f
C91 VTAIL.n4 VSUBS 1.87152f
C92 VTAIL.n5 VSUBS 0.749695f
C93 VTAIL.t3 VSUBS 2.46442f
C94 VTAIL.n6 VSUBS 2.05947f
C95 VTAIL.t11 VSUBS 2.46442f
C96 VTAIL.n7 VSUBS 2.05946f
C97 VTAIL.t9 VSUBS 0.252352f
C98 VTAIL.t14 VSUBS 0.252352f
C99 VTAIL.n8 VSUBS 1.87152f
C100 VTAIL.n9 VSUBS 0.749691f
C101 VTAIL.t12 VSUBS 2.46442f
C102 VTAIL.n10 VSUBS 0.785772f
C103 VTAIL.t4 VSUBS 2.46442f
C104 VTAIL.n11 VSUBS 0.785772f
C105 VTAIL.t2 VSUBS 0.252352f
C106 VTAIL.t5 VSUBS 0.252352f
C107 VTAIL.n12 VSUBS 1.87152f
C108 VTAIL.n13 VSUBS 0.749691f
C109 VTAIL.t6 VSUBS 2.46442f
C110 VTAIL.n14 VSUBS 2.05947f
C111 VTAIL.t8 VSUBS 2.46442f
C112 VTAIL.n15 VSUBS 2.05495f
C113 VDD2.t7 VSUBS 0.268514f
C114 VDD2.t6 VSUBS 0.268514f
C115 VDD2.n0 VSUBS 2.13765f
C116 VDD2.t2 VSUBS 0.268514f
C117 VDD2.t0 VSUBS 0.268514f
C118 VDD2.n1 VSUBS 2.13765f
C119 VDD2.n2 VSUBS 3.09631f
C120 VDD2.t4 VSUBS 0.268514f
C121 VDD2.t1 VSUBS 0.268514f
C122 VDD2.n3 VSUBS 2.13276f
C123 VDD2.n4 VSUBS 2.86712f
C124 VDD2.t5 VSUBS 0.268514f
C125 VDD2.t3 VSUBS 0.268514f
C126 VDD2.n5 VSUBS 2.13761f
C127 VN.n0 VSUBS 0.058695f
C128 VN.t4 VSUBS 1.7515f
C129 VN.n1 VSUBS 0.639372f
C130 VN.n2 VSUBS 0.228379f
C131 VN.t1 VSUBS 1.7515f
C132 VN.t7 VSUBS 1.87257f
C133 VN.n3 VSUBS 0.697866f
C134 VN.n4 VSUBS 0.707794f
C135 VN.n5 VSUBS 0.061378f
C136 VN.n6 VSUBS 0.061378f
C137 VN.n7 VSUBS 0.043987f
C138 VN.n8 VSUBS 0.043987f
C139 VN.n9 VSUBS 0.044338f
C140 VN.n10 VSUBS 0.052728f
C141 VN.t6 VSUBS 1.82563f
C142 VN.n11 VSUBS 0.714027f
C143 VN.n12 VSUBS 0.041196f
C144 VN.n13 VSUBS 0.058695f
C145 VN.t5 VSUBS 1.7515f
C146 VN.n14 VSUBS 0.639372f
C147 VN.n15 VSUBS 0.228379f
C148 VN.t0 VSUBS 1.7515f
C149 VN.t2 VSUBS 1.87257f
C150 VN.n16 VSUBS 0.697866f
C151 VN.n17 VSUBS 0.707794f
C152 VN.n18 VSUBS 0.061378f
C153 VN.n19 VSUBS 0.061378f
C154 VN.n20 VSUBS 0.043987f
C155 VN.n21 VSUBS 0.043987f
C156 VN.n22 VSUBS 0.044338f
C157 VN.n23 VSUBS 0.052728f
C158 VN.t3 VSUBS 1.82563f
C159 VN.n24 VSUBS 0.714027f
C160 VN.n25 VSUBS 2.07076f
C161 B.n0 VSUBS 0.004826f
C162 B.n1 VSUBS 0.004826f
C163 B.n2 VSUBS 0.007632f
C164 B.n3 VSUBS 0.007632f
C165 B.n4 VSUBS 0.007632f
C166 B.n5 VSUBS 0.007632f
C167 B.n6 VSUBS 0.007632f
C168 B.n7 VSUBS 0.007632f
C169 B.n8 VSUBS 0.007632f
C170 B.n9 VSUBS 0.007632f
C171 B.n10 VSUBS 0.007632f
C172 B.n11 VSUBS 0.007632f
C173 B.n12 VSUBS 0.007632f
C174 B.n13 VSUBS 0.007632f
C175 B.n14 VSUBS 0.007632f
C176 B.n15 VSUBS 0.007632f
C177 B.n16 VSUBS 0.018187f
C178 B.n17 VSUBS 0.007632f
C179 B.n18 VSUBS 0.007632f
C180 B.n19 VSUBS 0.007632f
C181 B.n20 VSUBS 0.007632f
C182 B.n21 VSUBS 0.007632f
C183 B.n22 VSUBS 0.007632f
C184 B.n23 VSUBS 0.007632f
C185 B.n24 VSUBS 0.007632f
C186 B.n25 VSUBS 0.007632f
C187 B.n26 VSUBS 0.007632f
C188 B.n27 VSUBS 0.007632f
C189 B.n28 VSUBS 0.007632f
C190 B.n29 VSUBS 0.007632f
C191 B.n30 VSUBS 0.007632f
C192 B.n31 VSUBS 0.007632f
C193 B.n32 VSUBS 0.007632f
C194 B.n33 VSUBS 0.007632f
C195 B.n34 VSUBS 0.007632f
C196 B.n35 VSUBS 0.007632f
C197 B.n36 VSUBS 0.007632f
C198 B.n37 VSUBS 0.007632f
C199 B.n38 VSUBS 0.007632f
C200 B.n39 VSUBS 0.007632f
C201 B.t5 VSUBS 0.475556f
C202 B.t4 VSUBS 0.487499f
C203 B.t3 VSUBS 0.6736f
C204 B.n40 VSUBS 0.191998f
C205 B.n41 VSUBS 0.071586f
C206 B.n42 VSUBS 0.007632f
C207 B.n43 VSUBS 0.007632f
C208 B.n44 VSUBS 0.007632f
C209 B.n45 VSUBS 0.007632f
C210 B.t11 VSUBS 0.475546f
C211 B.t10 VSUBS 0.487489f
C212 B.t9 VSUBS 0.6736f
C213 B.n46 VSUBS 0.192008f
C214 B.n47 VSUBS 0.071597f
C215 B.n48 VSUBS 0.017682f
C216 B.n49 VSUBS 0.007632f
C217 B.n50 VSUBS 0.007632f
C218 B.n51 VSUBS 0.007632f
C219 B.n52 VSUBS 0.007632f
C220 B.n53 VSUBS 0.007632f
C221 B.n54 VSUBS 0.007632f
C222 B.n55 VSUBS 0.007632f
C223 B.n56 VSUBS 0.007632f
C224 B.n57 VSUBS 0.007632f
C225 B.n58 VSUBS 0.007632f
C226 B.n59 VSUBS 0.007632f
C227 B.n60 VSUBS 0.007632f
C228 B.n61 VSUBS 0.007632f
C229 B.n62 VSUBS 0.007632f
C230 B.n63 VSUBS 0.007632f
C231 B.n64 VSUBS 0.007632f
C232 B.n65 VSUBS 0.007632f
C233 B.n66 VSUBS 0.007632f
C234 B.n67 VSUBS 0.007632f
C235 B.n68 VSUBS 0.007632f
C236 B.n69 VSUBS 0.007632f
C237 B.n70 VSUBS 0.007632f
C238 B.n71 VSUBS 0.018187f
C239 B.n72 VSUBS 0.007632f
C240 B.n73 VSUBS 0.007632f
C241 B.n74 VSUBS 0.007632f
C242 B.n75 VSUBS 0.007632f
C243 B.n76 VSUBS 0.007632f
C244 B.n77 VSUBS 0.007632f
C245 B.n78 VSUBS 0.007632f
C246 B.n79 VSUBS 0.007632f
C247 B.n80 VSUBS 0.007632f
C248 B.n81 VSUBS 0.007632f
C249 B.n82 VSUBS 0.007632f
C250 B.n83 VSUBS 0.007632f
C251 B.n84 VSUBS 0.007632f
C252 B.n85 VSUBS 0.007632f
C253 B.n86 VSUBS 0.007632f
C254 B.n87 VSUBS 0.007632f
C255 B.n88 VSUBS 0.007632f
C256 B.n89 VSUBS 0.007632f
C257 B.n90 VSUBS 0.007632f
C258 B.n91 VSUBS 0.007632f
C259 B.n92 VSUBS 0.007632f
C260 B.n93 VSUBS 0.007632f
C261 B.n94 VSUBS 0.007632f
C262 B.n95 VSUBS 0.007632f
C263 B.n96 VSUBS 0.007632f
C264 B.n97 VSUBS 0.007632f
C265 B.n98 VSUBS 0.007632f
C266 B.n99 VSUBS 0.007632f
C267 B.n100 VSUBS 0.018187f
C268 B.n101 VSUBS 0.007632f
C269 B.n102 VSUBS 0.007632f
C270 B.n103 VSUBS 0.007632f
C271 B.n104 VSUBS 0.007632f
C272 B.n105 VSUBS 0.007632f
C273 B.n106 VSUBS 0.007632f
C274 B.n107 VSUBS 0.007632f
C275 B.n108 VSUBS 0.007632f
C276 B.n109 VSUBS 0.007632f
C277 B.n110 VSUBS 0.007632f
C278 B.n111 VSUBS 0.007632f
C279 B.n112 VSUBS 0.007632f
C280 B.n113 VSUBS 0.007632f
C281 B.n114 VSUBS 0.007632f
C282 B.n115 VSUBS 0.007632f
C283 B.n116 VSUBS 0.007632f
C284 B.n117 VSUBS 0.007632f
C285 B.n118 VSUBS 0.007632f
C286 B.n119 VSUBS 0.007632f
C287 B.n120 VSUBS 0.007632f
C288 B.n121 VSUBS 0.007632f
C289 B.n122 VSUBS 0.007632f
C290 B.n123 VSUBS 0.007632f
C291 B.t7 VSUBS 0.475546f
C292 B.t8 VSUBS 0.487489f
C293 B.t6 VSUBS 0.6736f
C294 B.n124 VSUBS 0.192008f
C295 B.n125 VSUBS 0.071597f
C296 B.n126 VSUBS 0.007632f
C297 B.n127 VSUBS 0.007632f
C298 B.n128 VSUBS 0.007632f
C299 B.n129 VSUBS 0.007632f
C300 B.t1 VSUBS 0.475556f
C301 B.t2 VSUBS 0.487499f
C302 B.t0 VSUBS 0.6736f
C303 B.n130 VSUBS 0.191998f
C304 B.n131 VSUBS 0.071586f
C305 B.n132 VSUBS 0.017682f
C306 B.n133 VSUBS 0.007632f
C307 B.n134 VSUBS 0.007632f
C308 B.n135 VSUBS 0.007632f
C309 B.n136 VSUBS 0.007632f
C310 B.n137 VSUBS 0.007632f
C311 B.n138 VSUBS 0.007632f
C312 B.n139 VSUBS 0.007632f
C313 B.n140 VSUBS 0.007632f
C314 B.n141 VSUBS 0.007632f
C315 B.n142 VSUBS 0.007632f
C316 B.n143 VSUBS 0.007632f
C317 B.n144 VSUBS 0.007632f
C318 B.n145 VSUBS 0.007632f
C319 B.n146 VSUBS 0.007632f
C320 B.n147 VSUBS 0.007632f
C321 B.n148 VSUBS 0.007632f
C322 B.n149 VSUBS 0.007632f
C323 B.n150 VSUBS 0.007632f
C324 B.n151 VSUBS 0.007632f
C325 B.n152 VSUBS 0.007632f
C326 B.n153 VSUBS 0.007632f
C327 B.n154 VSUBS 0.007632f
C328 B.n155 VSUBS 0.018187f
C329 B.n156 VSUBS 0.007632f
C330 B.n157 VSUBS 0.007632f
C331 B.n158 VSUBS 0.007632f
C332 B.n159 VSUBS 0.007632f
C333 B.n160 VSUBS 0.007632f
C334 B.n161 VSUBS 0.007632f
C335 B.n162 VSUBS 0.007632f
C336 B.n163 VSUBS 0.007632f
C337 B.n164 VSUBS 0.007632f
C338 B.n165 VSUBS 0.007632f
C339 B.n166 VSUBS 0.007632f
C340 B.n167 VSUBS 0.007632f
C341 B.n168 VSUBS 0.007632f
C342 B.n169 VSUBS 0.007632f
C343 B.n170 VSUBS 0.007632f
C344 B.n171 VSUBS 0.007632f
C345 B.n172 VSUBS 0.007632f
C346 B.n173 VSUBS 0.007632f
C347 B.n174 VSUBS 0.007632f
C348 B.n175 VSUBS 0.007632f
C349 B.n176 VSUBS 0.007632f
C350 B.n177 VSUBS 0.007632f
C351 B.n178 VSUBS 0.007632f
C352 B.n179 VSUBS 0.007632f
C353 B.n180 VSUBS 0.007632f
C354 B.n181 VSUBS 0.007632f
C355 B.n182 VSUBS 0.007632f
C356 B.n183 VSUBS 0.007632f
C357 B.n184 VSUBS 0.007632f
C358 B.n185 VSUBS 0.007632f
C359 B.n186 VSUBS 0.007632f
C360 B.n187 VSUBS 0.007632f
C361 B.n188 VSUBS 0.007632f
C362 B.n189 VSUBS 0.007632f
C363 B.n190 VSUBS 0.007632f
C364 B.n191 VSUBS 0.007632f
C365 B.n192 VSUBS 0.007632f
C366 B.n193 VSUBS 0.007632f
C367 B.n194 VSUBS 0.007632f
C368 B.n195 VSUBS 0.007632f
C369 B.n196 VSUBS 0.007632f
C370 B.n197 VSUBS 0.007632f
C371 B.n198 VSUBS 0.007632f
C372 B.n199 VSUBS 0.007632f
C373 B.n200 VSUBS 0.007632f
C374 B.n201 VSUBS 0.007632f
C375 B.n202 VSUBS 0.007632f
C376 B.n203 VSUBS 0.007632f
C377 B.n204 VSUBS 0.007632f
C378 B.n205 VSUBS 0.007632f
C379 B.n206 VSUBS 0.007632f
C380 B.n207 VSUBS 0.007632f
C381 B.n208 VSUBS 0.007632f
C382 B.n209 VSUBS 0.007632f
C383 B.n210 VSUBS 0.018187f
C384 B.n211 VSUBS 0.019075f
C385 B.n212 VSUBS 0.019075f
C386 B.n213 VSUBS 0.007632f
C387 B.n214 VSUBS 0.007632f
C388 B.n215 VSUBS 0.007632f
C389 B.n216 VSUBS 0.007632f
C390 B.n217 VSUBS 0.007632f
C391 B.n218 VSUBS 0.007632f
C392 B.n219 VSUBS 0.007632f
C393 B.n220 VSUBS 0.007632f
C394 B.n221 VSUBS 0.007632f
C395 B.n222 VSUBS 0.007632f
C396 B.n223 VSUBS 0.007632f
C397 B.n224 VSUBS 0.007632f
C398 B.n225 VSUBS 0.007632f
C399 B.n226 VSUBS 0.007632f
C400 B.n227 VSUBS 0.007632f
C401 B.n228 VSUBS 0.007632f
C402 B.n229 VSUBS 0.007632f
C403 B.n230 VSUBS 0.007632f
C404 B.n231 VSUBS 0.007632f
C405 B.n232 VSUBS 0.007632f
C406 B.n233 VSUBS 0.007632f
C407 B.n234 VSUBS 0.007632f
C408 B.n235 VSUBS 0.007632f
C409 B.n236 VSUBS 0.007632f
C410 B.n237 VSUBS 0.007632f
C411 B.n238 VSUBS 0.007632f
C412 B.n239 VSUBS 0.007632f
C413 B.n240 VSUBS 0.007632f
C414 B.n241 VSUBS 0.007632f
C415 B.n242 VSUBS 0.007632f
C416 B.n243 VSUBS 0.007632f
C417 B.n244 VSUBS 0.007632f
C418 B.n245 VSUBS 0.007632f
C419 B.n246 VSUBS 0.007632f
C420 B.n247 VSUBS 0.007632f
C421 B.n248 VSUBS 0.007632f
C422 B.n249 VSUBS 0.007632f
C423 B.n250 VSUBS 0.007632f
C424 B.n251 VSUBS 0.007632f
C425 B.n252 VSUBS 0.007632f
C426 B.n253 VSUBS 0.007632f
C427 B.n254 VSUBS 0.007632f
C428 B.n255 VSUBS 0.007632f
C429 B.n256 VSUBS 0.007632f
C430 B.n257 VSUBS 0.007632f
C431 B.n258 VSUBS 0.007632f
C432 B.n259 VSUBS 0.007632f
C433 B.n260 VSUBS 0.007632f
C434 B.n261 VSUBS 0.007632f
C435 B.n262 VSUBS 0.007632f
C436 B.n263 VSUBS 0.007632f
C437 B.n264 VSUBS 0.007632f
C438 B.n265 VSUBS 0.007632f
C439 B.n266 VSUBS 0.007632f
C440 B.n267 VSUBS 0.007632f
C441 B.n268 VSUBS 0.007632f
C442 B.n269 VSUBS 0.007632f
C443 B.n270 VSUBS 0.007632f
C444 B.n271 VSUBS 0.007632f
C445 B.n272 VSUBS 0.007632f
C446 B.n273 VSUBS 0.007632f
C447 B.n274 VSUBS 0.007632f
C448 B.n275 VSUBS 0.007632f
C449 B.n276 VSUBS 0.007632f
C450 B.n277 VSUBS 0.007183f
C451 B.n278 VSUBS 0.007632f
C452 B.n279 VSUBS 0.007632f
C453 B.n280 VSUBS 0.004265f
C454 B.n281 VSUBS 0.007632f
C455 B.n282 VSUBS 0.007632f
C456 B.n283 VSUBS 0.007632f
C457 B.n284 VSUBS 0.007632f
C458 B.n285 VSUBS 0.007632f
C459 B.n286 VSUBS 0.007632f
C460 B.n287 VSUBS 0.007632f
C461 B.n288 VSUBS 0.007632f
C462 B.n289 VSUBS 0.007632f
C463 B.n290 VSUBS 0.007632f
C464 B.n291 VSUBS 0.007632f
C465 B.n292 VSUBS 0.007632f
C466 B.n293 VSUBS 0.004265f
C467 B.n294 VSUBS 0.017682f
C468 B.n295 VSUBS 0.007183f
C469 B.n296 VSUBS 0.007632f
C470 B.n297 VSUBS 0.007632f
C471 B.n298 VSUBS 0.007632f
C472 B.n299 VSUBS 0.007632f
C473 B.n300 VSUBS 0.007632f
C474 B.n301 VSUBS 0.007632f
C475 B.n302 VSUBS 0.007632f
C476 B.n303 VSUBS 0.007632f
C477 B.n304 VSUBS 0.007632f
C478 B.n305 VSUBS 0.007632f
C479 B.n306 VSUBS 0.007632f
C480 B.n307 VSUBS 0.007632f
C481 B.n308 VSUBS 0.007632f
C482 B.n309 VSUBS 0.007632f
C483 B.n310 VSUBS 0.007632f
C484 B.n311 VSUBS 0.007632f
C485 B.n312 VSUBS 0.007632f
C486 B.n313 VSUBS 0.007632f
C487 B.n314 VSUBS 0.007632f
C488 B.n315 VSUBS 0.007632f
C489 B.n316 VSUBS 0.007632f
C490 B.n317 VSUBS 0.007632f
C491 B.n318 VSUBS 0.007632f
C492 B.n319 VSUBS 0.007632f
C493 B.n320 VSUBS 0.007632f
C494 B.n321 VSUBS 0.007632f
C495 B.n322 VSUBS 0.007632f
C496 B.n323 VSUBS 0.007632f
C497 B.n324 VSUBS 0.007632f
C498 B.n325 VSUBS 0.007632f
C499 B.n326 VSUBS 0.007632f
C500 B.n327 VSUBS 0.007632f
C501 B.n328 VSUBS 0.007632f
C502 B.n329 VSUBS 0.007632f
C503 B.n330 VSUBS 0.007632f
C504 B.n331 VSUBS 0.007632f
C505 B.n332 VSUBS 0.007632f
C506 B.n333 VSUBS 0.007632f
C507 B.n334 VSUBS 0.007632f
C508 B.n335 VSUBS 0.007632f
C509 B.n336 VSUBS 0.007632f
C510 B.n337 VSUBS 0.007632f
C511 B.n338 VSUBS 0.007632f
C512 B.n339 VSUBS 0.007632f
C513 B.n340 VSUBS 0.007632f
C514 B.n341 VSUBS 0.007632f
C515 B.n342 VSUBS 0.007632f
C516 B.n343 VSUBS 0.007632f
C517 B.n344 VSUBS 0.007632f
C518 B.n345 VSUBS 0.007632f
C519 B.n346 VSUBS 0.007632f
C520 B.n347 VSUBS 0.007632f
C521 B.n348 VSUBS 0.007632f
C522 B.n349 VSUBS 0.007632f
C523 B.n350 VSUBS 0.007632f
C524 B.n351 VSUBS 0.007632f
C525 B.n352 VSUBS 0.007632f
C526 B.n353 VSUBS 0.007632f
C527 B.n354 VSUBS 0.007632f
C528 B.n355 VSUBS 0.007632f
C529 B.n356 VSUBS 0.007632f
C530 B.n357 VSUBS 0.007632f
C531 B.n358 VSUBS 0.007632f
C532 B.n359 VSUBS 0.007632f
C533 B.n360 VSUBS 0.007632f
C534 B.n361 VSUBS 0.019075f
C535 B.n362 VSUBS 0.019075f
C536 B.n363 VSUBS 0.018187f
C537 B.n364 VSUBS 0.007632f
C538 B.n365 VSUBS 0.007632f
C539 B.n366 VSUBS 0.007632f
C540 B.n367 VSUBS 0.007632f
C541 B.n368 VSUBS 0.007632f
C542 B.n369 VSUBS 0.007632f
C543 B.n370 VSUBS 0.007632f
C544 B.n371 VSUBS 0.007632f
C545 B.n372 VSUBS 0.007632f
C546 B.n373 VSUBS 0.007632f
C547 B.n374 VSUBS 0.007632f
C548 B.n375 VSUBS 0.007632f
C549 B.n376 VSUBS 0.007632f
C550 B.n377 VSUBS 0.007632f
C551 B.n378 VSUBS 0.007632f
C552 B.n379 VSUBS 0.007632f
C553 B.n380 VSUBS 0.007632f
C554 B.n381 VSUBS 0.007632f
C555 B.n382 VSUBS 0.007632f
C556 B.n383 VSUBS 0.007632f
C557 B.n384 VSUBS 0.007632f
C558 B.n385 VSUBS 0.007632f
C559 B.n386 VSUBS 0.007632f
C560 B.n387 VSUBS 0.007632f
C561 B.n388 VSUBS 0.007632f
C562 B.n389 VSUBS 0.007632f
C563 B.n390 VSUBS 0.007632f
C564 B.n391 VSUBS 0.007632f
C565 B.n392 VSUBS 0.007632f
C566 B.n393 VSUBS 0.007632f
C567 B.n394 VSUBS 0.007632f
C568 B.n395 VSUBS 0.007632f
C569 B.n396 VSUBS 0.007632f
C570 B.n397 VSUBS 0.007632f
C571 B.n398 VSUBS 0.007632f
C572 B.n399 VSUBS 0.007632f
C573 B.n400 VSUBS 0.007632f
C574 B.n401 VSUBS 0.007632f
C575 B.n402 VSUBS 0.007632f
C576 B.n403 VSUBS 0.007632f
C577 B.n404 VSUBS 0.007632f
C578 B.n405 VSUBS 0.007632f
C579 B.n406 VSUBS 0.007632f
C580 B.n407 VSUBS 0.007632f
C581 B.n408 VSUBS 0.007632f
C582 B.n409 VSUBS 0.007632f
C583 B.n410 VSUBS 0.007632f
C584 B.n411 VSUBS 0.007632f
C585 B.n412 VSUBS 0.007632f
C586 B.n413 VSUBS 0.007632f
C587 B.n414 VSUBS 0.007632f
C588 B.n415 VSUBS 0.007632f
C589 B.n416 VSUBS 0.007632f
C590 B.n417 VSUBS 0.007632f
C591 B.n418 VSUBS 0.007632f
C592 B.n419 VSUBS 0.007632f
C593 B.n420 VSUBS 0.007632f
C594 B.n421 VSUBS 0.007632f
C595 B.n422 VSUBS 0.007632f
C596 B.n423 VSUBS 0.007632f
C597 B.n424 VSUBS 0.007632f
C598 B.n425 VSUBS 0.007632f
C599 B.n426 VSUBS 0.007632f
C600 B.n427 VSUBS 0.007632f
C601 B.n428 VSUBS 0.007632f
C602 B.n429 VSUBS 0.007632f
C603 B.n430 VSUBS 0.007632f
C604 B.n431 VSUBS 0.007632f
C605 B.n432 VSUBS 0.007632f
C606 B.n433 VSUBS 0.007632f
C607 B.n434 VSUBS 0.007632f
C608 B.n435 VSUBS 0.007632f
C609 B.n436 VSUBS 0.007632f
C610 B.n437 VSUBS 0.007632f
C611 B.n438 VSUBS 0.007632f
C612 B.n439 VSUBS 0.007632f
C613 B.n440 VSUBS 0.007632f
C614 B.n441 VSUBS 0.007632f
C615 B.n442 VSUBS 0.007632f
C616 B.n443 VSUBS 0.007632f
C617 B.n444 VSUBS 0.007632f
C618 B.n445 VSUBS 0.007632f
C619 B.n446 VSUBS 0.007632f
C620 B.n447 VSUBS 0.007632f
C621 B.n448 VSUBS 0.007632f
C622 B.n449 VSUBS 0.007632f
C623 B.n450 VSUBS 0.019033f
C624 B.n451 VSUBS 0.018228f
C625 B.n452 VSUBS 0.019075f
C626 B.n453 VSUBS 0.007632f
C627 B.n454 VSUBS 0.007632f
C628 B.n455 VSUBS 0.007632f
C629 B.n456 VSUBS 0.007632f
C630 B.n457 VSUBS 0.007632f
C631 B.n458 VSUBS 0.007632f
C632 B.n459 VSUBS 0.007632f
C633 B.n460 VSUBS 0.007632f
C634 B.n461 VSUBS 0.007632f
C635 B.n462 VSUBS 0.007632f
C636 B.n463 VSUBS 0.007632f
C637 B.n464 VSUBS 0.007632f
C638 B.n465 VSUBS 0.007632f
C639 B.n466 VSUBS 0.007632f
C640 B.n467 VSUBS 0.007632f
C641 B.n468 VSUBS 0.007632f
C642 B.n469 VSUBS 0.007632f
C643 B.n470 VSUBS 0.007632f
C644 B.n471 VSUBS 0.007632f
C645 B.n472 VSUBS 0.007632f
C646 B.n473 VSUBS 0.007632f
C647 B.n474 VSUBS 0.007632f
C648 B.n475 VSUBS 0.007632f
C649 B.n476 VSUBS 0.007632f
C650 B.n477 VSUBS 0.007632f
C651 B.n478 VSUBS 0.007632f
C652 B.n479 VSUBS 0.007632f
C653 B.n480 VSUBS 0.007632f
C654 B.n481 VSUBS 0.007632f
C655 B.n482 VSUBS 0.007632f
C656 B.n483 VSUBS 0.007632f
C657 B.n484 VSUBS 0.007632f
C658 B.n485 VSUBS 0.007632f
C659 B.n486 VSUBS 0.007632f
C660 B.n487 VSUBS 0.007632f
C661 B.n488 VSUBS 0.007632f
C662 B.n489 VSUBS 0.007632f
C663 B.n490 VSUBS 0.007632f
C664 B.n491 VSUBS 0.007632f
C665 B.n492 VSUBS 0.007632f
C666 B.n493 VSUBS 0.007632f
C667 B.n494 VSUBS 0.007632f
C668 B.n495 VSUBS 0.007632f
C669 B.n496 VSUBS 0.007632f
C670 B.n497 VSUBS 0.007632f
C671 B.n498 VSUBS 0.007632f
C672 B.n499 VSUBS 0.007632f
C673 B.n500 VSUBS 0.007632f
C674 B.n501 VSUBS 0.007632f
C675 B.n502 VSUBS 0.007632f
C676 B.n503 VSUBS 0.007632f
C677 B.n504 VSUBS 0.007632f
C678 B.n505 VSUBS 0.007632f
C679 B.n506 VSUBS 0.007632f
C680 B.n507 VSUBS 0.007632f
C681 B.n508 VSUBS 0.007632f
C682 B.n509 VSUBS 0.007632f
C683 B.n510 VSUBS 0.007632f
C684 B.n511 VSUBS 0.007632f
C685 B.n512 VSUBS 0.007632f
C686 B.n513 VSUBS 0.007632f
C687 B.n514 VSUBS 0.007632f
C688 B.n515 VSUBS 0.007632f
C689 B.n516 VSUBS 0.007632f
C690 B.n517 VSUBS 0.007183f
C691 B.n518 VSUBS 0.007632f
C692 B.n519 VSUBS 0.007632f
C693 B.n520 VSUBS 0.004265f
C694 B.n521 VSUBS 0.007632f
C695 B.n522 VSUBS 0.007632f
C696 B.n523 VSUBS 0.007632f
C697 B.n524 VSUBS 0.007632f
C698 B.n525 VSUBS 0.007632f
C699 B.n526 VSUBS 0.007632f
C700 B.n527 VSUBS 0.007632f
C701 B.n528 VSUBS 0.007632f
C702 B.n529 VSUBS 0.007632f
C703 B.n530 VSUBS 0.007632f
C704 B.n531 VSUBS 0.007632f
C705 B.n532 VSUBS 0.007632f
C706 B.n533 VSUBS 0.004265f
C707 B.n534 VSUBS 0.017682f
C708 B.n535 VSUBS 0.007183f
C709 B.n536 VSUBS 0.007632f
C710 B.n537 VSUBS 0.007632f
C711 B.n538 VSUBS 0.007632f
C712 B.n539 VSUBS 0.007632f
C713 B.n540 VSUBS 0.007632f
C714 B.n541 VSUBS 0.007632f
C715 B.n542 VSUBS 0.007632f
C716 B.n543 VSUBS 0.007632f
C717 B.n544 VSUBS 0.007632f
C718 B.n545 VSUBS 0.007632f
C719 B.n546 VSUBS 0.007632f
C720 B.n547 VSUBS 0.007632f
C721 B.n548 VSUBS 0.007632f
C722 B.n549 VSUBS 0.007632f
C723 B.n550 VSUBS 0.007632f
C724 B.n551 VSUBS 0.007632f
C725 B.n552 VSUBS 0.007632f
C726 B.n553 VSUBS 0.007632f
C727 B.n554 VSUBS 0.007632f
C728 B.n555 VSUBS 0.007632f
C729 B.n556 VSUBS 0.007632f
C730 B.n557 VSUBS 0.007632f
C731 B.n558 VSUBS 0.007632f
C732 B.n559 VSUBS 0.007632f
C733 B.n560 VSUBS 0.007632f
C734 B.n561 VSUBS 0.007632f
C735 B.n562 VSUBS 0.007632f
C736 B.n563 VSUBS 0.007632f
C737 B.n564 VSUBS 0.007632f
C738 B.n565 VSUBS 0.007632f
C739 B.n566 VSUBS 0.007632f
C740 B.n567 VSUBS 0.007632f
C741 B.n568 VSUBS 0.007632f
C742 B.n569 VSUBS 0.007632f
C743 B.n570 VSUBS 0.007632f
C744 B.n571 VSUBS 0.007632f
C745 B.n572 VSUBS 0.007632f
C746 B.n573 VSUBS 0.007632f
C747 B.n574 VSUBS 0.007632f
C748 B.n575 VSUBS 0.007632f
C749 B.n576 VSUBS 0.007632f
C750 B.n577 VSUBS 0.007632f
C751 B.n578 VSUBS 0.007632f
C752 B.n579 VSUBS 0.007632f
C753 B.n580 VSUBS 0.007632f
C754 B.n581 VSUBS 0.007632f
C755 B.n582 VSUBS 0.007632f
C756 B.n583 VSUBS 0.007632f
C757 B.n584 VSUBS 0.007632f
C758 B.n585 VSUBS 0.007632f
C759 B.n586 VSUBS 0.007632f
C760 B.n587 VSUBS 0.007632f
C761 B.n588 VSUBS 0.007632f
C762 B.n589 VSUBS 0.007632f
C763 B.n590 VSUBS 0.007632f
C764 B.n591 VSUBS 0.007632f
C765 B.n592 VSUBS 0.007632f
C766 B.n593 VSUBS 0.007632f
C767 B.n594 VSUBS 0.007632f
C768 B.n595 VSUBS 0.007632f
C769 B.n596 VSUBS 0.007632f
C770 B.n597 VSUBS 0.007632f
C771 B.n598 VSUBS 0.007632f
C772 B.n599 VSUBS 0.007632f
C773 B.n600 VSUBS 0.007632f
C774 B.n601 VSUBS 0.019075f
C775 B.n602 VSUBS 0.019075f
C776 B.n603 VSUBS 0.018187f
C777 B.n604 VSUBS 0.007632f
C778 B.n605 VSUBS 0.007632f
C779 B.n606 VSUBS 0.007632f
C780 B.n607 VSUBS 0.007632f
C781 B.n608 VSUBS 0.007632f
C782 B.n609 VSUBS 0.007632f
C783 B.n610 VSUBS 0.007632f
C784 B.n611 VSUBS 0.007632f
C785 B.n612 VSUBS 0.007632f
C786 B.n613 VSUBS 0.007632f
C787 B.n614 VSUBS 0.007632f
C788 B.n615 VSUBS 0.007632f
C789 B.n616 VSUBS 0.007632f
C790 B.n617 VSUBS 0.007632f
C791 B.n618 VSUBS 0.007632f
C792 B.n619 VSUBS 0.007632f
C793 B.n620 VSUBS 0.007632f
C794 B.n621 VSUBS 0.007632f
C795 B.n622 VSUBS 0.007632f
C796 B.n623 VSUBS 0.007632f
C797 B.n624 VSUBS 0.007632f
C798 B.n625 VSUBS 0.007632f
C799 B.n626 VSUBS 0.007632f
C800 B.n627 VSUBS 0.007632f
C801 B.n628 VSUBS 0.007632f
C802 B.n629 VSUBS 0.007632f
C803 B.n630 VSUBS 0.007632f
C804 B.n631 VSUBS 0.007632f
C805 B.n632 VSUBS 0.007632f
C806 B.n633 VSUBS 0.007632f
C807 B.n634 VSUBS 0.007632f
C808 B.n635 VSUBS 0.007632f
C809 B.n636 VSUBS 0.007632f
C810 B.n637 VSUBS 0.007632f
C811 B.n638 VSUBS 0.007632f
C812 B.n639 VSUBS 0.007632f
C813 B.n640 VSUBS 0.007632f
C814 B.n641 VSUBS 0.007632f
C815 B.n642 VSUBS 0.007632f
C816 B.n643 VSUBS 0.007632f
C817 B.n644 VSUBS 0.007632f
C818 B.n645 VSUBS 0.007632f
C819 B.n646 VSUBS 0.007632f
C820 B.n647 VSUBS 0.017281f
.ends

