* NGSPICE file created from diff_pair_sample_1134.ext - technology: sky130A

.subckt diff_pair_sample_1134 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3595 pd=14.63 as=5.577 ps=29.38 w=14.3 l=0.34
X1 VTAIL.t4 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=5.577 pd=29.38 as=2.3595 ps=14.63 w=14.3 l=0.34
X2 VTAIL.t1 VP.t0 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.577 pd=29.38 as=2.3595 ps=14.63 w=14.3 l=0.34
X3 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=5.577 pd=29.38 as=0 ps=0 w=14.3 l=0.34
X4 VTAIL.t2 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.577 pd=29.38 as=2.3595 ps=14.63 w=14.3 l=0.34
X5 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3595 pd=14.63 as=5.577 ps=29.38 w=14.3 l=0.34
X6 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=5.577 pd=29.38 as=0 ps=0 w=14.3 l=0.34
X7 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=5.577 pd=29.38 as=0 ps=0 w=14.3 l=0.34
X8 VDD1.t0 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3595 pd=14.63 as=5.577 ps=29.38 w=14.3 l=0.34
X9 VTAIL.t5 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.577 pd=29.38 as=2.3595 ps=14.63 w=14.3 l=0.34
X10 VDD2.t0 VN.t3 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3595 pd=14.63 as=5.577 ps=29.38 w=14.3 l=0.34
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.577 pd=29.38 as=0 ps=0 w=14.3 l=0.34
R0 VN.n0 VN.t3 1154.67
R1 VN.n0 VN.t1 1154.67
R2 VN.n1 VN.t0 1154.67
R3 VN.n1 VN.t2 1154.67
R4 VN VN.n1 202.863
R5 VN VN.n0 161.351
R6 VTAIL.n5 VTAIL.t1 46.0595
R7 VTAIL.n4 VTAIL.t6 46.0595
R8 VTAIL.n3 VTAIL.t5 46.0595
R9 VTAIL.n7 VTAIL.t7 46.0594
R10 VTAIL.n0 VTAIL.t4 46.0594
R11 VTAIL.n1 VTAIL.t3 46.0594
R12 VTAIL.n2 VTAIL.t2 46.0594
R13 VTAIL.n6 VTAIL.t0 46.0594
R14 VTAIL.n7 VTAIL.n6 25.2893
R15 VTAIL.n3 VTAIL.n2 25.2893
R16 VTAIL.n4 VTAIL.n3 0.578086
R17 VTAIL.n6 VTAIL.n5 0.578086
R18 VTAIL.n2 VTAIL.n1 0.578086
R19 VTAIL.n5 VTAIL.n4 0.470328
R20 VTAIL.n1 VTAIL.n0 0.470328
R21 VTAIL VTAIL.n0 0.347483
R22 VTAIL VTAIL.n7 0.231103
R23 VDD2.n2 VDD2.n0 99.1459
R24 VDD2.n2 VDD2.n1 61.3536
R25 VDD2.n1 VDD2.t1 1.38512
R26 VDD2.n1 VDD2.t3 1.38512
R27 VDD2.n0 VDD2.t2 1.38512
R28 VDD2.n0 VDD2.t0 1.38512
R29 VDD2 VDD2.n2 0.0586897
R30 B.n147 B.t11 1225.7
R31 B.n139 B.t15 1225.7
R32 B.n55 B.t4 1225.7
R33 B.n61 B.t8 1225.7
R34 B.n445 B.n444 585
R35 B.n447 B.n87 585
R36 B.n450 B.n449 585
R37 B.n451 B.n86 585
R38 B.n453 B.n452 585
R39 B.n455 B.n85 585
R40 B.n458 B.n457 585
R41 B.n459 B.n84 585
R42 B.n461 B.n460 585
R43 B.n463 B.n83 585
R44 B.n466 B.n465 585
R45 B.n467 B.n82 585
R46 B.n469 B.n468 585
R47 B.n471 B.n81 585
R48 B.n474 B.n473 585
R49 B.n475 B.n80 585
R50 B.n477 B.n476 585
R51 B.n479 B.n79 585
R52 B.n482 B.n481 585
R53 B.n483 B.n78 585
R54 B.n485 B.n484 585
R55 B.n487 B.n77 585
R56 B.n490 B.n489 585
R57 B.n491 B.n76 585
R58 B.n493 B.n492 585
R59 B.n495 B.n75 585
R60 B.n498 B.n497 585
R61 B.n499 B.n74 585
R62 B.n501 B.n500 585
R63 B.n503 B.n73 585
R64 B.n506 B.n505 585
R65 B.n507 B.n72 585
R66 B.n509 B.n508 585
R67 B.n511 B.n71 585
R68 B.n514 B.n513 585
R69 B.n515 B.n70 585
R70 B.n517 B.n516 585
R71 B.n519 B.n69 585
R72 B.n522 B.n521 585
R73 B.n523 B.n68 585
R74 B.n525 B.n524 585
R75 B.n527 B.n67 585
R76 B.n530 B.n529 585
R77 B.n531 B.n66 585
R78 B.n533 B.n532 585
R79 B.n535 B.n65 585
R80 B.n537 B.n536 585
R81 B.n539 B.n538 585
R82 B.n542 B.n541 585
R83 B.n543 B.n60 585
R84 B.n545 B.n544 585
R85 B.n547 B.n59 585
R86 B.n550 B.n549 585
R87 B.n551 B.n58 585
R88 B.n553 B.n552 585
R89 B.n555 B.n57 585
R90 B.n558 B.n557 585
R91 B.n559 B.n54 585
R92 B.n562 B.n561 585
R93 B.n564 B.n53 585
R94 B.n567 B.n566 585
R95 B.n568 B.n52 585
R96 B.n570 B.n569 585
R97 B.n572 B.n51 585
R98 B.n575 B.n574 585
R99 B.n576 B.n50 585
R100 B.n578 B.n577 585
R101 B.n580 B.n49 585
R102 B.n583 B.n582 585
R103 B.n584 B.n48 585
R104 B.n586 B.n585 585
R105 B.n588 B.n47 585
R106 B.n591 B.n590 585
R107 B.n592 B.n46 585
R108 B.n594 B.n593 585
R109 B.n596 B.n45 585
R110 B.n599 B.n598 585
R111 B.n600 B.n44 585
R112 B.n602 B.n601 585
R113 B.n604 B.n43 585
R114 B.n607 B.n606 585
R115 B.n608 B.n42 585
R116 B.n610 B.n609 585
R117 B.n612 B.n41 585
R118 B.n615 B.n614 585
R119 B.n616 B.n40 585
R120 B.n618 B.n617 585
R121 B.n620 B.n39 585
R122 B.n623 B.n622 585
R123 B.n624 B.n38 585
R124 B.n626 B.n625 585
R125 B.n628 B.n37 585
R126 B.n631 B.n630 585
R127 B.n632 B.n36 585
R128 B.n634 B.n633 585
R129 B.n636 B.n35 585
R130 B.n639 B.n638 585
R131 B.n640 B.n34 585
R132 B.n642 B.n641 585
R133 B.n644 B.n33 585
R134 B.n647 B.n646 585
R135 B.n648 B.n32 585
R136 B.n650 B.n649 585
R137 B.n652 B.n31 585
R138 B.n655 B.n654 585
R139 B.n656 B.n30 585
R140 B.n443 B.n28 585
R141 B.n659 B.n28 585
R142 B.n442 B.n27 585
R143 B.n660 B.n27 585
R144 B.n441 B.n26 585
R145 B.n661 B.n26 585
R146 B.n440 B.n439 585
R147 B.n439 B.n22 585
R148 B.n438 B.n21 585
R149 B.n667 B.n21 585
R150 B.n437 B.n20 585
R151 B.n668 B.n20 585
R152 B.n436 B.n19 585
R153 B.n669 B.n19 585
R154 B.n435 B.n434 585
R155 B.n434 B.n15 585
R156 B.n433 B.n14 585
R157 B.n675 B.n14 585
R158 B.n432 B.n13 585
R159 B.n676 B.n13 585
R160 B.n431 B.n12 585
R161 B.n677 B.n12 585
R162 B.n430 B.n429 585
R163 B.n429 B.n11 585
R164 B.n428 B.n7 585
R165 B.n683 B.n7 585
R166 B.n427 B.n6 585
R167 B.n684 B.n6 585
R168 B.n426 B.n5 585
R169 B.n685 B.n5 585
R170 B.n425 B.n424 585
R171 B.n424 B.n4 585
R172 B.n423 B.n88 585
R173 B.n423 B.n422 585
R174 B.n412 B.n89 585
R175 B.n415 B.n89 585
R176 B.n414 B.n413 585
R177 B.n416 B.n414 585
R178 B.n411 B.n93 585
R179 B.n97 B.n93 585
R180 B.n410 B.n409 585
R181 B.n409 B.n408 585
R182 B.n95 B.n94 585
R183 B.n96 B.n95 585
R184 B.n401 B.n400 585
R185 B.n402 B.n401 585
R186 B.n399 B.n102 585
R187 B.n102 B.n101 585
R188 B.n398 B.n397 585
R189 B.n397 B.n396 585
R190 B.n104 B.n103 585
R191 B.n105 B.n104 585
R192 B.n389 B.n388 585
R193 B.n390 B.n389 585
R194 B.n387 B.n110 585
R195 B.n110 B.n109 585
R196 B.n386 B.n385 585
R197 B.n385 B.n384 585
R198 B.n381 B.n114 585
R199 B.n380 B.n379 585
R200 B.n377 B.n115 585
R201 B.n377 B.n113 585
R202 B.n376 B.n375 585
R203 B.n374 B.n373 585
R204 B.n372 B.n117 585
R205 B.n370 B.n369 585
R206 B.n368 B.n118 585
R207 B.n367 B.n366 585
R208 B.n364 B.n119 585
R209 B.n362 B.n361 585
R210 B.n360 B.n120 585
R211 B.n359 B.n358 585
R212 B.n356 B.n121 585
R213 B.n354 B.n353 585
R214 B.n352 B.n122 585
R215 B.n351 B.n350 585
R216 B.n348 B.n123 585
R217 B.n346 B.n345 585
R218 B.n344 B.n124 585
R219 B.n343 B.n342 585
R220 B.n340 B.n125 585
R221 B.n338 B.n337 585
R222 B.n336 B.n126 585
R223 B.n335 B.n334 585
R224 B.n332 B.n127 585
R225 B.n330 B.n329 585
R226 B.n328 B.n128 585
R227 B.n327 B.n326 585
R228 B.n324 B.n129 585
R229 B.n322 B.n321 585
R230 B.n320 B.n130 585
R231 B.n319 B.n318 585
R232 B.n316 B.n131 585
R233 B.n314 B.n313 585
R234 B.n312 B.n132 585
R235 B.n311 B.n310 585
R236 B.n308 B.n133 585
R237 B.n306 B.n305 585
R238 B.n304 B.n134 585
R239 B.n303 B.n302 585
R240 B.n300 B.n135 585
R241 B.n298 B.n297 585
R242 B.n296 B.n136 585
R243 B.n295 B.n294 585
R244 B.n292 B.n137 585
R245 B.n290 B.n289 585
R246 B.n288 B.n138 585
R247 B.n286 B.n285 585
R248 B.n283 B.n141 585
R249 B.n281 B.n280 585
R250 B.n279 B.n142 585
R251 B.n278 B.n277 585
R252 B.n275 B.n143 585
R253 B.n273 B.n272 585
R254 B.n271 B.n144 585
R255 B.n270 B.n269 585
R256 B.n267 B.n145 585
R257 B.n265 B.n264 585
R258 B.n263 B.n146 585
R259 B.n262 B.n261 585
R260 B.n259 B.n150 585
R261 B.n257 B.n256 585
R262 B.n255 B.n151 585
R263 B.n254 B.n253 585
R264 B.n251 B.n152 585
R265 B.n249 B.n248 585
R266 B.n247 B.n153 585
R267 B.n246 B.n245 585
R268 B.n243 B.n154 585
R269 B.n241 B.n240 585
R270 B.n239 B.n155 585
R271 B.n238 B.n237 585
R272 B.n235 B.n156 585
R273 B.n233 B.n232 585
R274 B.n231 B.n157 585
R275 B.n230 B.n229 585
R276 B.n227 B.n158 585
R277 B.n225 B.n224 585
R278 B.n223 B.n159 585
R279 B.n222 B.n221 585
R280 B.n219 B.n160 585
R281 B.n217 B.n216 585
R282 B.n215 B.n161 585
R283 B.n214 B.n213 585
R284 B.n211 B.n162 585
R285 B.n209 B.n208 585
R286 B.n207 B.n163 585
R287 B.n206 B.n205 585
R288 B.n203 B.n164 585
R289 B.n201 B.n200 585
R290 B.n199 B.n165 585
R291 B.n198 B.n197 585
R292 B.n195 B.n166 585
R293 B.n193 B.n192 585
R294 B.n191 B.n167 585
R295 B.n190 B.n189 585
R296 B.n187 B.n168 585
R297 B.n185 B.n184 585
R298 B.n183 B.n169 585
R299 B.n182 B.n181 585
R300 B.n179 B.n170 585
R301 B.n177 B.n176 585
R302 B.n175 B.n171 585
R303 B.n174 B.n173 585
R304 B.n112 B.n111 585
R305 B.n113 B.n112 585
R306 B.n383 B.n382 585
R307 B.n384 B.n383 585
R308 B.n108 B.n107 585
R309 B.n109 B.n108 585
R310 B.n392 B.n391 585
R311 B.n391 B.n390 585
R312 B.n393 B.n106 585
R313 B.n106 B.n105 585
R314 B.n395 B.n394 585
R315 B.n396 B.n395 585
R316 B.n100 B.n99 585
R317 B.n101 B.n100 585
R318 B.n404 B.n403 585
R319 B.n403 B.n402 585
R320 B.n405 B.n98 585
R321 B.n98 B.n96 585
R322 B.n407 B.n406 585
R323 B.n408 B.n407 585
R324 B.n92 B.n91 585
R325 B.n97 B.n92 585
R326 B.n418 B.n417 585
R327 B.n417 B.n416 585
R328 B.n419 B.n90 585
R329 B.n415 B.n90 585
R330 B.n421 B.n420 585
R331 B.n422 B.n421 585
R332 B.n2 B.n0 585
R333 B.n4 B.n2 585
R334 B.n3 B.n1 585
R335 B.n684 B.n3 585
R336 B.n682 B.n681 585
R337 B.n683 B.n682 585
R338 B.n680 B.n8 585
R339 B.n11 B.n8 585
R340 B.n679 B.n678 585
R341 B.n678 B.n677 585
R342 B.n10 B.n9 585
R343 B.n676 B.n10 585
R344 B.n674 B.n673 585
R345 B.n675 B.n674 585
R346 B.n672 B.n16 585
R347 B.n16 B.n15 585
R348 B.n671 B.n670 585
R349 B.n670 B.n669 585
R350 B.n18 B.n17 585
R351 B.n668 B.n18 585
R352 B.n666 B.n665 585
R353 B.n667 B.n666 585
R354 B.n664 B.n23 585
R355 B.n23 B.n22 585
R356 B.n663 B.n662 585
R357 B.n662 B.n661 585
R358 B.n25 B.n24 585
R359 B.n660 B.n25 585
R360 B.n658 B.n657 585
R361 B.n659 B.n658 585
R362 B.n687 B.n686 585
R363 B.n686 B.n685 585
R364 B.n383 B.n114 540.549
R365 B.n658 B.n30 540.549
R366 B.n385 B.n112 540.549
R367 B.n445 B.n28 540.549
R368 B.n446 B.n29 256.663
R369 B.n448 B.n29 256.663
R370 B.n454 B.n29 256.663
R371 B.n456 B.n29 256.663
R372 B.n462 B.n29 256.663
R373 B.n464 B.n29 256.663
R374 B.n470 B.n29 256.663
R375 B.n472 B.n29 256.663
R376 B.n478 B.n29 256.663
R377 B.n480 B.n29 256.663
R378 B.n486 B.n29 256.663
R379 B.n488 B.n29 256.663
R380 B.n494 B.n29 256.663
R381 B.n496 B.n29 256.663
R382 B.n502 B.n29 256.663
R383 B.n504 B.n29 256.663
R384 B.n510 B.n29 256.663
R385 B.n512 B.n29 256.663
R386 B.n518 B.n29 256.663
R387 B.n520 B.n29 256.663
R388 B.n526 B.n29 256.663
R389 B.n528 B.n29 256.663
R390 B.n534 B.n29 256.663
R391 B.n64 B.n29 256.663
R392 B.n540 B.n29 256.663
R393 B.n546 B.n29 256.663
R394 B.n548 B.n29 256.663
R395 B.n554 B.n29 256.663
R396 B.n556 B.n29 256.663
R397 B.n563 B.n29 256.663
R398 B.n565 B.n29 256.663
R399 B.n571 B.n29 256.663
R400 B.n573 B.n29 256.663
R401 B.n579 B.n29 256.663
R402 B.n581 B.n29 256.663
R403 B.n587 B.n29 256.663
R404 B.n589 B.n29 256.663
R405 B.n595 B.n29 256.663
R406 B.n597 B.n29 256.663
R407 B.n603 B.n29 256.663
R408 B.n605 B.n29 256.663
R409 B.n611 B.n29 256.663
R410 B.n613 B.n29 256.663
R411 B.n619 B.n29 256.663
R412 B.n621 B.n29 256.663
R413 B.n627 B.n29 256.663
R414 B.n629 B.n29 256.663
R415 B.n635 B.n29 256.663
R416 B.n637 B.n29 256.663
R417 B.n643 B.n29 256.663
R418 B.n645 B.n29 256.663
R419 B.n651 B.n29 256.663
R420 B.n653 B.n29 256.663
R421 B.n378 B.n113 256.663
R422 B.n116 B.n113 256.663
R423 B.n371 B.n113 256.663
R424 B.n365 B.n113 256.663
R425 B.n363 B.n113 256.663
R426 B.n357 B.n113 256.663
R427 B.n355 B.n113 256.663
R428 B.n349 B.n113 256.663
R429 B.n347 B.n113 256.663
R430 B.n341 B.n113 256.663
R431 B.n339 B.n113 256.663
R432 B.n333 B.n113 256.663
R433 B.n331 B.n113 256.663
R434 B.n325 B.n113 256.663
R435 B.n323 B.n113 256.663
R436 B.n317 B.n113 256.663
R437 B.n315 B.n113 256.663
R438 B.n309 B.n113 256.663
R439 B.n307 B.n113 256.663
R440 B.n301 B.n113 256.663
R441 B.n299 B.n113 256.663
R442 B.n293 B.n113 256.663
R443 B.n291 B.n113 256.663
R444 B.n284 B.n113 256.663
R445 B.n282 B.n113 256.663
R446 B.n276 B.n113 256.663
R447 B.n274 B.n113 256.663
R448 B.n268 B.n113 256.663
R449 B.n266 B.n113 256.663
R450 B.n260 B.n113 256.663
R451 B.n258 B.n113 256.663
R452 B.n252 B.n113 256.663
R453 B.n250 B.n113 256.663
R454 B.n244 B.n113 256.663
R455 B.n242 B.n113 256.663
R456 B.n236 B.n113 256.663
R457 B.n234 B.n113 256.663
R458 B.n228 B.n113 256.663
R459 B.n226 B.n113 256.663
R460 B.n220 B.n113 256.663
R461 B.n218 B.n113 256.663
R462 B.n212 B.n113 256.663
R463 B.n210 B.n113 256.663
R464 B.n204 B.n113 256.663
R465 B.n202 B.n113 256.663
R466 B.n196 B.n113 256.663
R467 B.n194 B.n113 256.663
R468 B.n188 B.n113 256.663
R469 B.n186 B.n113 256.663
R470 B.n180 B.n113 256.663
R471 B.n178 B.n113 256.663
R472 B.n172 B.n113 256.663
R473 B.n383 B.n108 163.367
R474 B.n391 B.n108 163.367
R475 B.n391 B.n106 163.367
R476 B.n395 B.n106 163.367
R477 B.n395 B.n100 163.367
R478 B.n403 B.n100 163.367
R479 B.n403 B.n98 163.367
R480 B.n407 B.n98 163.367
R481 B.n407 B.n92 163.367
R482 B.n417 B.n92 163.367
R483 B.n417 B.n90 163.367
R484 B.n421 B.n90 163.367
R485 B.n421 B.n2 163.367
R486 B.n686 B.n2 163.367
R487 B.n686 B.n3 163.367
R488 B.n682 B.n3 163.367
R489 B.n682 B.n8 163.367
R490 B.n678 B.n8 163.367
R491 B.n678 B.n10 163.367
R492 B.n674 B.n10 163.367
R493 B.n674 B.n16 163.367
R494 B.n670 B.n16 163.367
R495 B.n670 B.n18 163.367
R496 B.n666 B.n18 163.367
R497 B.n666 B.n23 163.367
R498 B.n662 B.n23 163.367
R499 B.n662 B.n25 163.367
R500 B.n658 B.n25 163.367
R501 B.n379 B.n377 163.367
R502 B.n377 B.n376 163.367
R503 B.n373 B.n372 163.367
R504 B.n370 B.n118 163.367
R505 B.n366 B.n364 163.367
R506 B.n362 B.n120 163.367
R507 B.n358 B.n356 163.367
R508 B.n354 B.n122 163.367
R509 B.n350 B.n348 163.367
R510 B.n346 B.n124 163.367
R511 B.n342 B.n340 163.367
R512 B.n338 B.n126 163.367
R513 B.n334 B.n332 163.367
R514 B.n330 B.n128 163.367
R515 B.n326 B.n324 163.367
R516 B.n322 B.n130 163.367
R517 B.n318 B.n316 163.367
R518 B.n314 B.n132 163.367
R519 B.n310 B.n308 163.367
R520 B.n306 B.n134 163.367
R521 B.n302 B.n300 163.367
R522 B.n298 B.n136 163.367
R523 B.n294 B.n292 163.367
R524 B.n290 B.n138 163.367
R525 B.n285 B.n283 163.367
R526 B.n281 B.n142 163.367
R527 B.n277 B.n275 163.367
R528 B.n273 B.n144 163.367
R529 B.n269 B.n267 163.367
R530 B.n265 B.n146 163.367
R531 B.n261 B.n259 163.367
R532 B.n257 B.n151 163.367
R533 B.n253 B.n251 163.367
R534 B.n249 B.n153 163.367
R535 B.n245 B.n243 163.367
R536 B.n241 B.n155 163.367
R537 B.n237 B.n235 163.367
R538 B.n233 B.n157 163.367
R539 B.n229 B.n227 163.367
R540 B.n225 B.n159 163.367
R541 B.n221 B.n219 163.367
R542 B.n217 B.n161 163.367
R543 B.n213 B.n211 163.367
R544 B.n209 B.n163 163.367
R545 B.n205 B.n203 163.367
R546 B.n201 B.n165 163.367
R547 B.n197 B.n195 163.367
R548 B.n193 B.n167 163.367
R549 B.n189 B.n187 163.367
R550 B.n185 B.n169 163.367
R551 B.n181 B.n179 163.367
R552 B.n177 B.n171 163.367
R553 B.n173 B.n112 163.367
R554 B.n385 B.n110 163.367
R555 B.n389 B.n110 163.367
R556 B.n389 B.n104 163.367
R557 B.n397 B.n104 163.367
R558 B.n397 B.n102 163.367
R559 B.n401 B.n102 163.367
R560 B.n401 B.n95 163.367
R561 B.n409 B.n95 163.367
R562 B.n409 B.n93 163.367
R563 B.n414 B.n93 163.367
R564 B.n414 B.n89 163.367
R565 B.n423 B.n89 163.367
R566 B.n424 B.n423 163.367
R567 B.n424 B.n5 163.367
R568 B.n6 B.n5 163.367
R569 B.n7 B.n6 163.367
R570 B.n429 B.n7 163.367
R571 B.n429 B.n12 163.367
R572 B.n13 B.n12 163.367
R573 B.n14 B.n13 163.367
R574 B.n434 B.n14 163.367
R575 B.n434 B.n19 163.367
R576 B.n20 B.n19 163.367
R577 B.n21 B.n20 163.367
R578 B.n439 B.n21 163.367
R579 B.n439 B.n26 163.367
R580 B.n27 B.n26 163.367
R581 B.n28 B.n27 163.367
R582 B.n654 B.n652 163.367
R583 B.n650 B.n32 163.367
R584 B.n646 B.n644 163.367
R585 B.n642 B.n34 163.367
R586 B.n638 B.n636 163.367
R587 B.n634 B.n36 163.367
R588 B.n630 B.n628 163.367
R589 B.n626 B.n38 163.367
R590 B.n622 B.n620 163.367
R591 B.n618 B.n40 163.367
R592 B.n614 B.n612 163.367
R593 B.n610 B.n42 163.367
R594 B.n606 B.n604 163.367
R595 B.n602 B.n44 163.367
R596 B.n598 B.n596 163.367
R597 B.n594 B.n46 163.367
R598 B.n590 B.n588 163.367
R599 B.n586 B.n48 163.367
R600 B.n582 B.n580 163.367
R601 B.n578 B.n50 163.367
R602 B.n574 B.n572 163.367
R603 B.n570 B.n52 163.367
R604 B.n566 B.n564 163.367
R605 B.n562 B.n54 163.367
R606 B.n557 B.n555 163.367
R607 B.n553 B.n58 163.367
R608 B.n549 B.n547 163.367
R609 B.n545 B.n60 163.367
R610 B.n541 B.n539 163.367
R611 B.n536 B.n535 163.367
R612 B.n533 B.n66 163.367
R613 B.n529 B.n527 163.367
R614 B.n525 B.n68 163.367
R615 B.n521 B.n519 163.367
R616 B.n517 B.n70 163.367
R617 B.n513 B.n511 163.367
R618 B.n509 B.n72 163.367
R619 B.n505 B.n503 163.367
R620 B.n501 B.n74 163.367
R621 B.n497 B.n495 163.367
R622 B.n493 B.n76 163.367
R623 B.n489 B.n487 163.367
R624 B.n485 B.n78 163.367
R625 B.n481 B.n479 163.367
R626 B.n477 B.n80 163.367
R627 B.n473 B.n471 163.367
R628 B.n469 B.n82 163.367
R629 B.n465 B.n463 163.367
R630 B.n461 B.n84 163.367
R631 B.n457 B.n455 163.367
R632 B.n453 B.n86 163.367
R633 B.n449 B.n447 163.367
R634 B.n147 B.t14 80.9098
R635 B.n61 B.t9 80.9098
R636 B.n139 B.t17 80.8911
R637 B.n55 B.t6 80.8911
R638 B.n378 B.n114 71.676
R639 B.n376 B.n116 71.676
R640 B.n372 B.n371 71.676
R641 B.n365 B.n118 71.676
R642 B.n364 B.n363 71.676
R643 B.n357 B.n120 71.676
R644 B.n356 B.n355 71.676
R645 B.n349 B.n122 71.676
R646 B.n348 B.n347 71.676
R647 B.n341 B.n124 71.676
R648 B.n340 B.n339 71.676
R649 B.n333 B.n126 71.676
R650 B.n332 B.n331 71.676
R651 B.n325 B.n128 71.676
R652 B.n324 B.n323 71.676
R653 B.n317 B.n130 71.676
R654 B.n316 B.n315 71.676
R655 B.n309 B.n132 71.676
R656 B.n308 B.n307 71.676
R657 B.n301 B.n134 71.676
R658 B.n300 B.n299 71.676
R659 B.n293 B.n136 71.676
R660 B.n292 B.n291 71.676
R661 B.n284 B.n138 71.676
R662 B.n283 B.n282 71.676
R663 B.n276 B.n142 71.676
R664 B.n275 B.n274 71.676
R665 B.n268 B.n144 71.676
R666 B.n267 B.n266 71.676
R667 B.n260 B.n146 71.676
R668 B.n259 B.n258 71.676
R669 B.n252 B.n151 71.676
R670 B.n251 B.n250 71.676
R671 B.n244 B.n153 71.676
R672 B.n243 B.n242 71.676
R673 B.n236 B.n155 71.676
R674 B.n235 B.n234 71.676
R675 B.n228 B.n157 71.676
R676 B.n227 B.n226 71.676
R677 B.n220 B.n159 71.676
R678 B.n219 B.n218 71.676
R679 B.n212 B.n161 71.676
R680 B.n211 B.n210 71.676
R681 B.n204 B.n163 71.676
R682 B.n203 B.n202 71.676
R683 B.n196 B.n165 71.676
R684 B.n195 B.n194 71.676
R685 B.n188 B.n167 71.676
R686 B.n187 B.n186 71.676
R687 B.n180 B.n169 71.676
R688 B.n179 B.n178 71.676
R689 B.n172 B.n171 71.676
R690 B.n653 B.n30 71.676
R691 B.n652 B.n651 71.676
R692 B.n645 B.n32 71.676
R693 B.n644 B.n643 71.676
R694 B.n637 B.n34 71.676
R695 B.n636 B.n635 71.676
R696 B.n629 B.n36 71.676
R697 B.n628 B.n627 71.676
R698 B.n621 B.n38 71.676
R699 B.n620 B.n619 71.676
R700 B.n613 B.n40 71.676
R701 B.n612 B.n611 71.676
R702 B.n605 B.n42 71.676
R703 B.n604 B.n603 71.676
R704 B.n597 B.n44 71.676
R705 B.n596 B.n595 71.676
R706 B.n589 B.n46 71.676
R707 B.n588 B.n587 71.676
R708 B.n581 B.n48 71.676
R709 B.n580 B.n579 71.676
R710 B.n573 B.n50 71.676
R711 B.n572 B.n571 71.676
R712 B.n565 B.n52 71.676
R713 B.n564 B.n563 71.676
R714 B.n556 B.n54 71.676
R715 B.n555 B.n554 71.676
R716 B.n548 B.n58 71.676
R717 B.n547 B.n546 71.676
R718 B.n540 B.n60 71.676
R719 B.n539 B.n64 71.676
R720 B.n535 B.n534 71.676
R721 B.n528 B.n66 71.676
R722 B.n527 B.n526 71.676
R723 B.n520 B.n68 71.676
R724 B.n519 B.n518 71.676
R725 B.n512 B.n70 71.676
R726 B.n511 B.n510 71.676
R727 B.n504 B.n72 71.676
R728 B.n503 B.n502 71.676
R729 B.n496 B.n74 71.676
R730 B.n495 B.n494 71.676
R731 B.n488 B.n76 71.676
R732 B.n487 B.n486 71.676
R733 B.n480 B.n78 71.676
R734 B.n479 B.n478 71.676
R735 B.n472 B.n80 71.676
R736 B.n471 B.n470 71.676
R737 B.n464 B.n82 71.676
R738 B.n463 B.n462 71.676
R739 B.n456 B.n84 71.676
R740 B.n455 B.n454 71.676
R741 B.n448 B.n86 71.676
R742 B.n447 B.n446 71.676
R743 B.n446 B.n445 71.676
R744 B.n449 B.n448 71.676
R745 B.n454 B.n453 71.676
R746 B.n457 B.n456 71.676
R747 B.n462 B.n461 71.676
R748 B.n465 B.n464 71.676
R749 B.n470 B.n469 71.676
R750 B.n473 B.n472 71.676
R751 B.n478 B.n477 71.676
R752 B.n481 B.n480 71.676
R753 B.n486 B.n485 71.676
R754 B.n489 B.n488 71.676
R755 B.n494 B.n493 71.676
R756 B.n497 B.n496 71.676
R757 B.n502 B.n501 71.676
R758 B.n505 B.n504 71.676
R759 B.n510 B.n509 71.676
R760 B.n513 B.n512 71.676
R761 B.n518 B.n517 71.676
R762 B.n521 B.n520 71.676
R763 B.n526 B.n525 71.676
R764 B.n529 B.n528 71.676
R765 B.n534 B.n533 71.676
R766 B.n536 B.n64 71.676
R767 B.n541 B.n540 71.676
R768 B.n546 B.n545 71.676
R769 B.n549 B.n548 71.676
R770 B.n554 B.n553 71.676
R771 B.n557 B.n556 71.676
R772 B.n563 B.n562 71.676
R773 B.n566 B.n565 71.676
R774 B.n571 B.n570 71.676
R775 B.n574 B.n573 71.676
R776 B.n579 B.n578 71.676
R777 B.n582 B.n581 71.676
R778 B.n587 B.n586 71.676
R779 B.n590 B.n589 71.676
R780 B.n595 B.n594 71.676
R781 B.n598 B.n597 71.676
R782 B.n603 B.n602 71.676
R783 B.n606 B.n605 71.676
R784 B.n611 B.n610 71.676
R785 B.n614 B.n613 71.676
R786 B.n619 B.n618 71.676
R787 B.n622 B.n621 71.676
R788 B.n627 B.n626 71.676
R789 B.n630 B.n629 71.676
R790 B.n635 B.n634 71.676
R791 B.n638 B.n637 71.676
R792 B.n643 B.n642 71.676
R793 B.n646 B.n645 71.676
R794 B.n651 B.n650 71.676
R795 B.n654 B.n653 71.676
R796 B.n379 B.n378 71.676
R797 B.n373 B.n116 71.676
R798 B.n371 B.n370 71.676
R799 B.n366 B.n365 71.676
R800 B.n363 B.n362 71.676
R801 B.n358 B.n357 71.676
R802 B.n355 B.n354 71.676
R803 B.n350 B.n349 71.676
R804 B.n347 B.n346 71.676
R805 B.n342 B.n341 71.676
R806 B.n339 B.n338 71.676
R807 B.n334 B.n333 71.676
R808 B.n331 B.n330 71.676
R809 B.n326 B.n325 71.676
R810 B.n323 B.n322 71.676
R811 B.n318 B.n317 71.676
R812 B.n315 B.n314 71.676
R813 B.n310 B.n309 71.676
R814 B.n307 B.n306 71.676
R815 B.n302 B.n301 71.676
R816 B.n299 B.n298 71.676
R817 B.n294 B.n293 71.676
R818 B.n291 B.n290 71.676
R819 B.n285 B.n284 71.676
R820 B.n282 B.n281 71.676
R821 B.n277 B.n276 71.676
R822 B.n274 B.n273 71.676
R823 B.n269 B.n268 71.676
R824 B.n266 B.n265 71.676
R825 B.n261 B.n260 71.676
R826 B.n258 B.n257 71.676
R827 B.n253 B.n252 71.676
R828 B.n250 B.n249 71.676
R829 B.n245 B.n244 71.676
R830 B.n242 B.n241 71.676
R831 B.n237 B.n236 71.676
R832 B.n234 B.n233 71.676
R833 B.n229 B.n228 71.676
R834 B.n226 B.n225 71.676
R835 B.n221 B.n220 71.676
R836 B.n218 B.n217 71.676
R837 B.n213 B.n212 71.676
R838 B.n210 B.n209 71.676
R839 B.n205 B.n204 71.676
R840 B.n202 B.n201 71.676
R841 B.n197 B.n196 71.676
R842 B.n194 B.n193 71.676
R843 B.n189 B.n188 71.676
R844 B.n186 B.n185 71.676
R845 B.n181 B.n180 71.676
R846 B.n178 B.n177 71.676
R847 B.n173 B.n172 71.676
R848 B.n384 B.n113 70.1715
R849 B.n659 B.n29 70.1715
R850 B.n148 B.t13 67.9159
R851 B.n62 B.t10 67.9159
R852 B.n140 B.t16 67.8972
R853 B.n56 B.t7 67.8972
R854 B.n149 B.n148 59.5399
R855 B.n287 B.n140 59.5399
R856 B.n560 B.n56 59.5399
R857 B.n63 B.n62 59.5399
R858 B.n384 B.n109 38.1735
R859 B.n390 B.n109 38.1735
R860 B.n390 B.n105 38.1735
R861 B.n396 B.n105 38.1735
R862 B.n402 B.n101 38.1735
R863 B.n402 B.n96 38.1735
R864 B.n408 B.n96 38.1735
R865 B.n408 B.n97 38.1735
R866 B.n416 B.n415 38.1735
R867 B.n422 B.n4 38.1735
R868 B.n685 B.n4 38.1735
R869 B.n685 B.n684 38.1735
R870 B.n684 B.n683 38.1735
R871 B.n677 B.n11 38.1735
R872 B.n676 B.n675 38.1735
R873 B.n675 B.n15 38.1735
R874 B.n669 B.n15 38.1735
R875 B.n669 B.n668 38.1735
R876 B.n667 B.n22 38.1735
R877 B.n661 B.n22 38.1735
R878 B.n661 B.n660 38.1735
R879 B.n660 B.n659 38.1735
R880 B.n657 B.n656 35.1225
R881 B.n444 B.n443 35.1225
R882 B.n386 B.n111 35.1225
R883 B.n382 B.n381 35.1225
R884 B.t12 B.n101 28.0689
R885 B.n668 B.t5 28.0689
R886 B.n422 B.t3 22.4552
R887 B.n683 B.t1 22.4552
R888 B.n416 B.t2 21.3325
R889 B.n677 B.t0 21.3325
R890 B B.n687 18.0485
R891 B.n97 B.t2 16.8415
R892 B.t0 B.n676 16.8415
R893 B.n415 B.t3 15.7188
R894 B.n11 B.t1 15.7188
R895 B.n148 B.n147 12.9944
R896 B.n140 B.n139 12.9944
R897 B.n56 B.n55 12.9944
R898 B.n62 B.n61 12.9944
R899 B.n656 B.n655 10.6151
R900 B.n655 B.n31 10.6151
R901 B.n649 B.n31 10.6151
R902 B.n649 B.n648 10.6151
R903 B.n648 B.n647 10.6151
R904 B.n647 B.n33 10.6151
R905 B.n641 B.n33 10.6151
R906 B.n641 B.n640 10.6151
R907 B.n640 B.n639 10.6151
R908 B.n639 B.n35 10.6151
R909 B.n633 B.n35 10.6151
R910 B.n633 B.n632 10.6151
R911 B.n632 B.n631 10.6151
R912 B.n631 B.n37 10.6151
R913 B.n625 B.n37 10.6151
R914 B.n625 B.n624 10.6151
R915 B.n624 B.n623 10.6151
R916 B.n623 B.n39 10.6151
R917 B.n617 B.n39 10.6151
R918 B.n617 B.n616 10.6151
R919 B.n616 B.n615 10.6151
R920 B.n615 B.n41 10.6151
R921 B.n609 B.n41 10.6151
R922 B.n609 B.n608 10.6151
R923 B.n608 B.n607 10.6151
R924 B.n607 B.n43 10.6151
R925 B.n601 B.n43 10.6151
R926 B.n601 B.n600 10.6151
R927 B.n600 B.n599 10.6151
R928 B.n599 B.n45 10.6151
R929 B.n593 B.n45 10.6151
R930 B.n593 B.n592 10.6151
R931 B.n592 B.n591 10.6151
R932 B.n591 B.n47 10.6151
R933 B.n585 B.n47 10.6151
R934 B.n585 B.n584 10.6151
R935 B.n584 B.n583 10.6151
R936 B.n583 B.n49 10.6151
R937 B.n577 B.n49 10.6151
R938 B.n577 B.n576 10.6151
R939 B.n576 B.n575 10.6151
R940 B.n575 B.n51 10.6151
R941 B.n569 B.n51 10.6151
R942 B.n569 B.n568 10.6151
R943 B.n568 B.n567 10.6151
R944 B.n567 B.n53 10.6151
R945 B.n561 B.n53 10.6151
R946 B.n559 B.n558 10.6151
R947 B.n558 B.n57 10.6151
R948 B.n552 B.n57 10.6151
R949 B.n552 B.n551 10.6151
R950 B.n551 B.n550 10.6151
R951 B.n550 B.n59 10.6151
R952 B.n544 B.n59 10.6151
R953 B.n544 B.n543 10.6151
R954 B.n543 B.n542 10.6151
R955 B.n538 B.n537 10.6151
R956 B.n537 B.n65 10.6151
R957 B.n532 B.n65 10.6151
R958 B.n532 B.n531 10.6151
R959 B.n531 B.n530 10.6151
R960 B.n530 B.n67 10.6151
R961 B.n524 B.n67 10.6151
R962 B.n524 B.n523 10.6151
R963 B.n523 B.n522 10.6151
R964 B.n522 B.n69 10.6151
R965 B.n516 B.n69 10.6151
R966 B.n516 B.n515 10.6151
R967 B.n515 B.n514 10.6151
R968 B.n514 B.n71 10.6151
R969 B.n508 B.n71 10.6151
R970 B.n508 B.n507 10.6151
R971 B.n507 B.n506 10.6151
R972 B.n506 B.n73 10.6151
R973 B.n500 B.n73 10.6151
R974 B.n500 B.n499 10.6151
R975 B.n499 B.n498 10.6151
R976 B.n498 B.n75 10.6151
R977 B.n492 B.n75 10.6151
R978 B.n492 B.n491 10.6151
R979 B.n491 B.n490 10.6151
R980 B.n490 B.n77 10.6151
R981 B.n484 B.n77 10.6151
R982 B.n484 B.n483 10.6151
R983 B.n483 B.n482 10.6151
R984 B.n482 B.n79 10.6151
R985 B.n476 B.n79 10.6151
R986 B.n476 B.n475 10.6151
R987 B.n475 B.n474 10.6151
R988 B.n474 B.n81 10.6151
R989 B.n468 B.n81 10.6151
R990 B.n468 B.n467 10.6151
R991 B.n467 B.n466 10.6151
R992 B.n466 B.n83 10.6151
R993 B.n460 B.n83 10.6151
R994 B.n460 B.n459 10.6151
R995 B.n459 B.n458 10.6151
R996 B.n458 B.n85 10.6151
R997 B.n452 B.n85 10.6151
R998 B.n452 B.n451 10.6151
R999 B.n451 B.n450 10.6151
R1000 B.n450 B.n87 10.6151
R1001 B.n444 B.n87 10.6151
R1002 B.n387 B.n386 10.6151
R1003 B.n388 B.n387 10.6151
R1004 B.n388 B.n103 10.6151
R1005 B.n398 B.n103 10.6151
R1006 B.n399 B.n398 10.6151
R1007 B.n400 B.n399 10.6151
R1008 B.n400 B.n94 10.6151
R1009 B.n410 B.n94 10.6151
R1010 B.n411 B.n410 10.6151
R1011 B.n413 B.n411 10.6151
R1012 B.n413 B.n412 10.6151
R1013 B.n412 B.n88 10.6151
R1014 B.n425 B.n88 10.6151
R1015 B.n426 B.n425 10.6151
R1016 B.n427 B.n426 10.6151
R1017 B.n428 B.n427 10.6151
R1018 B.n430 B.n428 10.6151
R1019 B.n431 B.n430 10.6151
R1020 B.n432 B.n431 10.6151
R1021 B.n433 B.n432 10.6151
R1022 B.n435 B.n433 10.6151
R1023 B.n436 B.n435 10.6151
R1024 B.n437 B.n436 10.6151
R1025 B.n438 B.n437 10.6151
R1026 B.n440 B.n438 10.6151
R1027 B.n441 B.n440 10.6151
R1028 B.n442 B.n441 10.6151
R1029 B.n443 B.n442 10.6151
R1030 B.n381 B.n380 10.6151
R1031 B.n380 B.n115 10.6151
R1032 B.n375 B.n115 10.6151
R1033 B.n375 B.n374 10.6151
R1034 B.n374 B.n117 10.6151
R1035 B.n369 B.n117 10.6151
R1036 B.n369 B.n368 10.6151
R1037 B.n368 B.n367 10.6151
R1038 B.n367 B.n119 10.6151
R1039 B.n361 B.n119 10.6151
R1040 B.n361 B.n360 10.6151
R1041 B.n360 B.n359 10.6151
R1042 B.n359 B.n121 10.6151
R1043 B.n353 B.n121 10.6151
R1044 B.n353 B.n352 10.6151
R1045 B.n352 B.n351 10.6151
R1046 B.n351 B.n123 10.6151
R1047 B.n345 B.n123 10.6151
R1048 B.n345 B.n344 10.6151
R1049 B.n344 B.n343 10.6151
R1050 B.n343 B.n125 10.6151
R1051 B.n337 B.n125 10.6151
R1052 B.n337 B.n336 10.6151
R1053 B.n336 B.n335 10.6151
R1054 B.n335 B.n127 10.6151
R1055 B.n329 B.n127 10.6151
R1056 B.n329 B.n328 10.6151
R1057 B.n328 B.n327 10.6151
R1058 B.n327 B.n129 10.6151
R1059 B.n321 B.n129 10.6151
R1060 B.n321 B.n320 10.6151
R1061 B.n320 B.n319 10.6151
R1062 B.n319 B.n131 10.6151
R1063 B.n313 B.n131 10.6151
R1064 B.n313 B.n312 10.6151
R1065 B.n312 B.n311 10.6151
R1066 B.n311 B.n133 10.6151
R1067 B.n305 B.n133 10.6151
R1068 B.n305 B.n304 10.6151
R1069 B.n304 B.n303 10.6151
R1070 B.n303 B.n135 10.6151
R1071 B.n297 B.n135 10.6151
R1072 B.n297 B.n296 10.6151
R1073 B.n296 B.n295 10.6151
R1074 B.n295 B.n137 10.6151
R1075 B.n289 B.n137 10.6151
R1076 B.n289 B.n288 10.6151
R1077 B.n286 B.n141 10.6151
R1078 B.n280 B.n141 10.6151
R1079 B.n280 B.n279 10.6151
R1080 B.n279 B.n278 10.6151
R1081 B.n278 B.n143 10.6151
R1082 B.n272 B.n143 10.6151
R1083 B.n272 B.n271 10.6151
R1084 B.n271 B.n270 10.6151
R1085 B.n270 B.n145 10.6151
R1086 B.n264 B.n263 10.6151
R1087 B.n263 B.n262 10.6151
R1088 B.n262 B.n150 10.6151
R1089 B.n256 B.n150 10.6151
R1090 B.n256 B.n255 10.6151
R1091 B.n255 B.n254 10.6151
R1092 B.n254 B.n152 10.6151
R1093 B.n248 B.n152 10.6151
R1094 B.n248 B.n247 10.6151
R1095 B.n247 B.n246 10.6151
R1096 B.n246 B.n154 10.6151
R1097 B.n240 B.n154 10.6151
R1098 B.n240 B.n239 10.6151
R1099 B.n239 B.n238 10.6151
R1100 B.n238 B.n156 10.6151
R1101 B.n232 B.n156 10.6151
R1102 B.n232 B.n231 10.6151
R1103 B.n231 B.n230 10.6151
R1104 B.n230 B.n158 10.6151
R1105 B.n224 B.n158 10.6151
R1106 B.n224 B.n223 10.6151
R1107 B.n223 B.n222 10.6151
R1108 B.n222 B.n160 10.6151
R1109 B.n216 B.n160 10.6151
R1110 B.n216 B.n215 10.6151
R1111 B.n215 B.n214 10.6151
R1112 B.n214 B.n162 10.6151
R1113 B.n208 B.n162 10.6151
R1114 B.n208 B.n207 10.6151
R1115 B.n207 B.n206 10.6151
R1116 B.n206 B.n164 10.6151
R1117 B.n200 B.n164 10.6151
R1118 B.n200 B.n199 10.6151
R1119 B.n199 B.n198 10.6151
R1120 B.n198 B.n166 10.6151
R1121 B.n192 B.n166 10.6151
R1122 B.n192 B.n191 10.6151
R1123 B.n191 B.n190 10.6151
R1124 B.n190 B.n168 10.6151
R1125 B.n184 B.n168 10.6151
R1126 B.n184 B.n183 10.6151
R1127 B.n183 B.n182 10.6151
R1128 B.n182 B.n170 10.6151
R1129 B.n176 B.n170 10.6151
R1130 B.n176 B.n175 10.6151
R1131 B.n175 B.n174 10.6151
R1132 B.n174 B.n111 10.6151
R1133 B.n382 B.n107 10.6151
R1134 B.n392 B.n107 10.6151
R1135 B.n393 B.n392 10.6151
R1136 B.n394 B.n393 10.6151
R1137 B.n394 B.n99 10.6151
R1138 B.n404 B.n99 10.6151
R1139 B.n405 B.n404 10.6151
R1140 B.n406 B.n405 10.6151
R1141 B.n406 B.n91 10.6151
R1142 B.n418 B.n91 10.6151
R1143 B.n419 B.n418 10.6151
R1144 B.n420 B.n419 10.6151
R1145 B.n420 B.n0 10.6151
R1146 B.n681 B.n1 10.6151
R1147 B.n681 B.n680 10.6151
R1148 B.n680 B.n679 10.6151
R1149 B.n679 B.n9 10.6151
R1150 B.n673 B.n9 10.6151
R1151 B.n673 B.n672 10.6151
R1152 B.n672 B.n671 10.6151
R1153 B.n671 B.n17 10.6151
R1154 B.n665 B.n17 10.6151
R1155 B.n665 B.n664 10.6151
R1156 B.n664 B.n663 10.6151
R1157 B.n663 B.n24 10.6151
R1158 B.n657 B.n24 10.6151
R1159 B.n396 B.t12 10.1051
R1160 B.t5 B.n667 10.1051
R1161 B.n561 B.n560 8.74196
R1162 B.n538 B.n63 8.74196
R1163 B.n288 B.n287 8.74196
R1164 B.n264 B.n149 8.74196
R1165 B.n687 B.n0 2.81026
R1166 B.n687 B.n1 2.81026
R1167 B.n560 B.n559 1.87367
R1168 B.n542 B.n63 1.87367
R1169 B.n287 B.n286 1.87367
R1170 B.n149 B.n145 1.87367
R1171 VP.n1 VP.t2 1154.67
R1172 VP.n1 VP.t1 1154.67
R1173 VP.n0 VP.t3 1154.67
R1174 VP.n0 VP.t0 1154.67
R1175 VP.n2 VP.n0 202.482
R1176 VP.n2 VP.n1 161.3
R1177 VP VP.n2 0.0516364
R1178 VDD1 VDD1.n1 99.6707
R1179 VDD1 VDD1.n0 61.4118
R1180 VDD1.n0 VDD1.t3 1.38512
R1181 VDD1.n0 VDD1.t0 1.38512
R1182 VDD1.n1 VDD1.t2 1.38512
R1183 VDD1.n1 VDD1.t1 1.38512
C0 VN VDD2 2.58944f
C1 VTAIL VDD1 10.456901f
C2 VDD2 VP 0.251304f
C3 VTAIL VN 1.97694f
C4 VTAIL VP 1.99105f
C5 VTAIL VDD2 10.496f
C6 VN VDD1 0.147764f
C7 VDD1 VP 2.69282f
C8 VDD1 VDD2 0.486883f
C9 VN VP 4.9835f
C10 VDD2 B 2.679163f
C11 VDD1 B 7.07894f
C12 VTAIL B 9.819319f
C13 VN B 7.89013f
C14 VP B 4.28721f
C15 VDD1.t3 B 0.366001f
C16 VDD1.t0 B 0.366001f
C17 VDD1.n0 B 3.30168f
C18 VDD1.t2 B 0.366001f
C19 VDD1.t1 B 0.366001f
C20 VDD1.n1 B 4.10404f
C21 VP.t0 B 0.676702f
C22 VP.t3 B 0.676702f
C23 VP.n0 B 0.919281f
C24 VP.t1 B 0.676702f
C25 VP.t2 B 0.676702f
C26 VP.n1 B 0.522028f
C27 VP.n2 B 3.5257f
C28 VDD2.t2 B 0.366551f
C29 VDD2.t0 B 0.366551f
C30 VDD2.n0 B 4.07834f
C31 VDD2.t1 B 0.366551f
C32 VDD2.t3 B 0.366551f
C33 VDD2.n1 B 3.30631f
C34 VDD2.n2 B 4.18179f
C35 VTAIL.t4 B 1.95175f
C36 VTAIL.n0 B 0.246503f
C37 VTAIL.t3 B 1.95175f
C38 VTAIL.n1 B 0.257993f
C39 VTAIL.t2 B 1.95175f
C40 VTAIL.n2 B 1.0885f
C41 VTAIL.t5 B 1.95176f
C42 VTAIL.n3 B 1.08849f
C43 VTAIL.t6 B 1.95176f
C44 VTAIL.n4 B 0.257979f
C45 VTAIL.t1 B 1.95176f
C46 VTAIL.n5 B 0.257979f
C47 VTAIL.t0 B 1.95175f
C48 VTAIL.n6 B 1.0885f
C49 VTAIL.t7 B 1.95175f
C50 VTAIL.n7 B 1.07122f
C51 VN.t1 B 0.662049f
C52 VN.t3 B 0.662049f
C53 VN.n0 B 0.51074f
C54 VN.t2 B 0.662049f
C55 VN.t0 B 0.662049f
C56 VN.n1 B 0.908624f
.ends

