* NGSPICE file created from diff_pair_sample_0652.ext - technology: sky130A

.subckt diff_pair_sample_0652 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7626 pd=35.46 as=0 ps=0 w=17.34 l=3.91
X1 VDD2.t5 VN.t0 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=6.7626 pd=35.46 as=2.8611 ps=17.67 w=17.34 l=3.91
X2 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=6.7626 pd=35.46 as=0 ps=0 w=17.34 l=3.91
X3 VTAIL.t5 VP.t0 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8611 pd=17.67 as=2.8611 ps=17.67 w=17.34 l=3.91
X4 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.7626 pd=35.46 as=0 ps=0 w=17.34 l=3.91
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7626 pd=35.46 as=0 ps=0 w=17.34 l=3.91
X6 VDD1.t4 VP.t1 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7626 pd=35.46 as=2.8611 ps=17.67 w=17.34 l=3.91
X7 VTAIL.t10 VN.t1 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8611 pd=17.67 as=2.8611 ps=17.67 w=17.34 l=3.91
X8 VDD2.t3 VN.t2 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8611 pd=17.67 as=6.7626 ps=35.46 w=17.34 l=3.91
X9 VDD1.t3 VP.t2 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8611 pd=17.67 as=6.7626 ps=35.46 w=17.34 l=3.91
X10 VTAIL.t9 VN.t3 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8611 pd=17.67 as=2.8611 ps=17.67 w=17.34 l=3.91
X11 VTAIL.t3 VP.t3 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8611 pd=17.67 as=2.8611 ps=17.67 w=17.34 l=3.91
X12 VDD1.t1 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8611 pd=17.67 as=6.7626 ps=35.46 w=17.34 l=3.91
X13 VDD2.t1 VN.t4 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=6.7626 pd=35.46 as=2.8611 ps=17.67 w=17.34 l=3.91
X14 VDD1.t0 VP.t5 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=6.7626 pd=35.46 as=2.8611 ps=17.67 w=17.34 l=3.91
X15 VDD2.t0 VN.t5 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.8611 pd=17.67 as=6.7626 ps=35.46 w=17.34 l=3.91
R0 B.n851 B.n850 585
R1 B.n853 B.n173 585
R2 B.n856 B.n855 585
R3 B.n857 B.n172 585
R4 B.n859 B.n858 585
R5 B.n861 B.n171 585
R6 B.n864 B.n863 585
R7 B.n865 B.n170 585
R8 B.n867 B.n866 585
R9 B.n869 B.n169 585
R10 B.n872 B.n871 585
R11 B.n873 B.n168 585
R12 B.n875 B.n874 585
R13 B.n877 B.n167 585
R14 B.n880 B.n879 585
R15 B.n881 B.n166 585
R16 B.n883 B.n882 585
R17 B.n885 B.n165 585
R18 B.n888 B.n887 585
R19 B.n889 B.n164 585
R20 B.n891 B.n890 585
R21 B.n893 B.n163 585
R22 B.n896 B.n895 585
R23 B.n897 B.n162 585
R24 B.n899 B.n898 585
R25 B.n901 B.n161 585
R26 B.n904 B.n903 585
R27 B.n905 B.n160 585
R28 B.n907 B.n906 585
R29 B.n909 B.n159 585
R30 B.n912 B.n911 585
R31 B.n913 B.n158 585
R32 B.n915 B.n914 585
R33 B.n917 B.n157 585
R34 B.n920 B.n919 585
R35 B.n921 B.n156 585
R36 B.n923 B.n922 585
R37 B.n925 B.n155 585
R38 B.n928 B.n927 585
R39 B.n929 B.n154 585
R40 B.n931 B.n930 585
R41 B.n933 B.n153 585
R42 B.n936 B.n935 585
R43 B.n937 B.n152 585
R44 B.n939 B.n938 585
R45 B.n941 B.n151 585
R46 B.n944 B.n943 585
R47 B.n945 B.n150 585
R48 B.n947 B.n946 585
R49 B.n949 B.n149 585
R50 B.n952 B.n951 585
R51 B.n953 B.n148 585
R52 B.n955 B.n954 585
R53 B.n957 B.n147 585
R54 B.n960 B.n959 585
R55 B.n961 B.n143 585
R56 B.n963 B.n962 585
R57 B.n965 B.n142 585
R58 B.n968 B.n967 585
R59 B.n969 B.n141 585
R60 B.n971 B.n970 585
R61 B.n973 B.n140 585
R62 B.n976 B.n975 585
R63 B.n977 B.n139 585
R64 B.n979 B.n978 585
R65 B.n981 B.n138 585
R66 B.n984 B.n983 585
R67 B.n986 B.n135 585
R68 B.n988 B.n987 585
R69 B.n990 B.n134 585
R70 B.n993 B.n992 585
R71 B.n994 B.n133 585
R72 B.n996 B.n995 585
R73 B.n998 B.n132 585
R74 B.n1001 B.n1000 585
R75 B.n1002 B.n131 585
R76 B.n1004 B.n1003 585
R77 B.n1006 B.n130 585
R78 B.n1009 B.n1008 585
R79 B.n1010 B.n129 585
R80 B.n1012 B.n1011 585
R81 B.n1014 B.n128 585
R82 B.n1017 B.n1016 585
R83 B.n1018 B.n127 585
R84 B.n1020 B.n1019 585
R85 B.n1022 B.n126 585
R86 B.n1025 B.n1024 585
R87 B.n1026 B.n125 585
R88 B.n1028 B.n1027 585
R89 B.n1030 B.n124 585
R90 B.n1033 B.n1032 585
R91 B.n1034 B.n123 585
R92 B.n1036 B.n1035 585
R93 B.n1038 B.n122 585
R94 B.n1041 B.n1040 585
R95 B.n1042 B.n121 585
R96 B.n1044 B.n1043 585
R97 B.n1046 B.n120 585
R98 B.n1049 B.n1048 585
R99 B.n1050 B.n119 585
R100 B.n1052 B.n1051 585
R101 B.n1054 B.n118 585
R102 B.n1057 B.n1056 585
R103 B.n1058 B.n117 585
R104 B.n1060 B.n1059 585
R105 B.n1062 B.n116 585
R106 B.n1065 B.n1064 585
R107 B.n1066 B.n115 585
R108 B.n1068 B.n1067 585
R109 B.n1070 B.n114 585
R110 B.n1073 B.n1072 585
R111 B.n1074 B.n113 585
R112 B.n1076 B.n1075 585
R113 B.n1078 B.n112 585
R114 B.n1081 B.n1080 585
R115 B.n1082 B.n111 585
R116 B.n1084 B.n1083 585
R117 B.n1086 B.n110 585
R118 B.n1089 B.n1088 585
R119 B.n1090 B.n109 585
R120 B.n1092 B.n1091 585
R121 B.n1094 B.n108 585
R122 B.n1097 B.n1096 585
R123 B.n1098 B.n107 585
R124 B.n849 B.n105 585
R125 B.n1101 B.n105 585
R126 B.n848 B.n104 585
R127 B.n1102 B.n104 585
R128 B.n847 B.n103 585
R129 B.n1103 B.n103 585
R130 B.n846 B.n845 585
R131 B.n845 B.n99 585
R132 B.n844 B.n98 585
R133 B.n1109 B.n98 585
R134 B.n843 B.n97 585
R135 B.n1110 B.n97 585
R136 B.n842 B.n96 585
R137 B.n1111 B.n96 585
R138 B.n841 B.n840 585
R139 B.n840 B.n92 585
R140 B.n839 B.n91 585
R141 B.n1117 B.n91 585
R142 B.n838 B.n90 585
R143 B.n1118 B.n90 585
R144 B.n837 B.n89 585
R145 B.n1119 B.n89 585
R146 B.n836 B.n835 585
R147 B.n835 B.n85 585
R148 B.n834 B.n84 585
R149 B.n1125 B.n84 585
R150 B.n833 B.n83 585
R151 B.n1126 B.n83 585
R152 B.n832 B.n82 585
R153 B.n1127 B.n82 585
R154 B.n831 B.n830 585
R155 B.n830 B.n78 585
R156 B.n829 B.n77 585
R157 B.n1133 B.n77 585
R158 B.n828 B.n76 585
R159 B.n1134 B.n76 585
R160 B.n827 B.n75 585
R161 B.n1135 B.n75 585
R162 B.n826 B.n825 585
R163 B.n825 B.n71 585
R164 B.n824 B.n70 585
R165 B.n1141 B.n70 585
R166 B.n823 B.n69 585
R167 B.n1142 B.n69 585
R168 B.n822 B.n68 585
R169 B.n1143 B.n68 585
R170 B.n821 B.n820 585
R171 B.n820 B.n64 585
R172 B.n819 B.n63 585
R173 B.n1149 B.n63 585
R174 B.n818 B.n62 585
R175 B.n1150 B.n62 585
R176 B.n817 B.n61 585
R177 B.n1151 B.n61 585
R178 B.n816 B.n815 585
R179 B.n815 B.n57 585
R180 B.n814 B.n56 585
R181 B.n1157 B.n56 585
R182 B.n813 B.n55 585
R183 B.n1158 B.n55 585
R184 B.n812 B.n54 585
R185 B.n1159 B.n54 585
R186 B.n811 B.n810 585
R187 B.n810 B.n50 585
R188 B.n809 B.n49 585
R189 B.n1165 B.n49 585
R190 B.n808 B.n48 585
R191 B.n1166 B.n48 585
R192 B.n807 B.n47 585
R193 B.n1167 B.n47 585
R194 B.n806 B.n805 585
R195 B.n805 B.n43 585
R196 B.n804 B.n42 585
R197 B.n1173 B.n42 585
R198 B.n803 B.n41 585
R199 B.n1174 B.n41 585
R200 B.n802 B.n40 585
R201 B.n1175 B.n40 585
R202 B.n801 B.n800 585
R203 B.n800 B.n36 585
R204 B.n799 B.n35 585
R205 B.n1181 B.n35 585
R206 B.n798 B.n34 585
R207 B.n1182 B.n34 585
R208 B.n797 B.n33 585
R209 B.n1183 B.n33 585
R210 B.n796 B.n795 585
R211 B.n795 B.n29 585
R212 B.n794 B.n28 585
R213 B.n1189 B.n28 585
R214 B.n793 B.n27 585
R215 B.n1190 B.n27 585
R216 B.n792 B.n26 585
R217 B.n1191 B.n26 585
R218 B.n791 B.n790 585
R219 B.n790 B.n22 585
R220 B.n789 B.n21 585
R221 B.n1197 B.n21 585
R222 B.n788 B.n20 585
R223 B.n1198 B.n20 585
R224 B.n787 B.n19 585
R225 B.n1199 B.n19 585
R226 B.n786 B.n785 585
R227 B.n785 B.n15 585
R228 B.n784 B.n14 585
R229 B.n1205 B.n14 585
R230 B.n783 B.n13 585
R231 B.n1206 B.n13 585
R232 B.n782 B.n12 585
R233 B.n1207 B.n12 585
R234 B.n781 B.n780 585
R235 B.n780 B.n8 585
R236 B.n779 B.n7 585
R237 B.n1213 B.n7 585
R238 B.n778 B.n6 585
R239 B.n1214 B.n6 585
R240 B.n777 B.n5 585
R241 B.n1215 B.n5 585
R242 B.n776 B.n775 585
R243 B.n775 B.n4 585
R244 B.n774 B.n174 585
R245 B.n774 B.n773 585
R246 B.n764 B.n175 585
R247 B.n176 B.n175 585
R248 B.n766 B.n765 585
R249 B.n767 B.n766 585
R250 B.n763 B.n181 585
R251 B.n181 B.n180 585
R252 B.n762 B.n761 585
R253 B.n761 B.n760 585
R254 B.n183 B.n182 585
R255 B.n184 B.n183 585
R256 B.n753 B.n752 585
R257 B.n754 B.n753 585
R258 B.n751 B.n189 585
R259 B.n189 B.n188 585
R260 B.n750 B.n749 585
R261 B.n749 B.n748 585
R262 B.n191 B.n190 585
R263 B.n192 B.n191 585
R264 B.n741 B.n740 585
R265 B.n742 B.n741 585
R266 B.n739 B.n197 585
R267 B.n197 B.n196 585
R268 B.n738 B.n737 585
R269 B.n737 B.n736 585
R270 B.n199 B.n198 585
R271 B.n200 B.n199 585
R272 B.n729 B.n728 585
R273 B.n730 B.n729 585
R274 B.n727 B.n205 585
R275 B.n205 B.n204 585
R276 B.n726 B.n725 585
R277 B.n725 B.n724 585
R278 B.n207 B.n206 585
R279 B.n208 B.n207 585
R280 B.n717 B.n716 585
R281 B.n718 B.n717 585
R282 B.n715 B.n212 585
R283 B.n216 B.n212 585
R284 B.n714 B.n713 585
R285 B.n713 B.n712 585
R286 B.n214 B.n213 585
R287 B.n215 B.n214 585
R288 B.n705 B.n704 585
R289 B.n706 B.n705 585
R290 B.n703 B.n221 585
R291 B.n221 B.n220 585
R292 B.n702 B.n701 585
R293 B.n701 B.n700 585
R294 B.n223 B.n222 585
R295 B.n224 B.n223 585
R296 B.n693 B.n692 585
R297 B.n694 B.n693 585
R298 B.n691 B.n229 585
R299 B.n229 B.n228 585
R300 B.n690 B.n689 585
R301 B.n689 B.n688 585
R302 B.n231 B.n230 585
R303 B.n232 B.n231 585
R304 B.n681 B.n680 585
R305 B.n682 B.n681 585
R306 B.n679 B.n236 585
R307 B.n240 B.n236 585
R308 B.n678 B.n677 585
R309 B.n677 B.n676 585
R310 B.n238 B.n237 585
R311 B.n239 B.n238 585
R312 B.n669 B.n668 585
R313 B.n670 B.n669 585
R314 B.n667 B.n245 585
R315 B.n245 B.n244 585
R316 B.n666 B.n665 585
R317 B.n665 B.n664 585
R318 B.n247 B.n246 585
R319 B.n248 B.n247 585
R320 B.n657 B.n656 585
R321 B.n658 B.n657 585
R322 B.n655 B.n253 585
R323 B.n253 B.n252 585
R324 B.n654 B.n653 585
R325 B.n653 B.n652 585
R326 B.n255 B.n254 585
R327 B.n256 B.n255 585
R328 B.n645 B.n644 585
R329 B.n646 B.n645 585
R330 B.n643 B.n261 585
R331 B.n261 B.n260 585
R332 B.n642 B.n641 585
R333 B.n641 B.n640 585
R334 B.n263 B.n262 585
R335 B.n264 B.n263 585
R336 B.n633 B.n632 585
R337 B.n634 B.n633 585
R338 B.n631 B.n268 585
R339 B.n272 B.n268 585
R340 B.n630 B.n629 585
R341 B.n629 B.n628 585
R342 B.n270 B.n269 585
R343 B.n271 B.n270 585
R344 B.n621 B.n620 585
R345 B.n622 B.n621 585
R346 B.n619 B.n277 585
R347 B.n277 B.n276 585
R348 B.n618 B.n617 585
R349 B.n617 B.n616 585
R350 B.n279 B.n278 585
R351 B.n280 B.n279 585
R352 B.n609 B.n608 585
R353 B.n610 B.n609 585
R354 B.n607 B.n285 585
R355 B.n285 B.n284 585
R356 B.n606 B.n605 585
R357 B.n605 B.n604 585
R358 B.n601 B.n289 585
R359 B.n600 B.n599 585
R360 B.n597 B.n290 585
R361 B.n597 B.n288 585
R362 B.n596 B.n595 585
R363 B.n594 B.n593 585
R364 B.n592 B.n292 585
R365 B.n590 B.n589 585
R366 B.n588 B.n293 585
R367 B.n587 B.n586 585
R368 B.n584 B.n294 585
R369 B.n582 B.n581 585
R370 B.n580 B.n295 585
R371 B.n579 B.n578 585
R372 B.n576 B.n296 585
R373 B.n574 B.n573 585
R374 B.n572 B.n297 585
R375 B.n571 B.n570 585
R376 B.n568 B.n298 585
R377 B.n566 B.n565 585
R378 B.n564 B.n299 585
R379 B.n563 B.n562 585
R380 B.n560 B.n300 585
R381 B.n558 B.n557 585
R382 B.n556 B.n301 585
R383 B.n555 B.n554 585
R384 B.n552 B.n302 585
R385 B.n550 B.n549 585
R386 B.n548 B.n303 585
R387 B.n547 B.n546 585
R388 B.n544 B.n304 585
R389 B.n542 B.n541 585
R390 B.n540 B.n305 585
R391 B.n539 B.n538 585
R392 B.n536 B.n306 585
R393 B.n534 B.n533 585
R394 B.n532 B.n307 585
R395 B.n531 B.n530 585
R396 B.n528 B.n308 585
R397 B.n526 B.n525 585
R398 B.n524 B.n309 585
R399 B.n523 B.n522 585
R400 B.n520 B.n310 585
R401 B.n518 B.n517 585
R402 B.n516 B.n311 585
R403 B.n515 B.n514 585
R404 B.n512 B.n312 585
R405 B.n510 B.n509 585
R406 B.n508 B.n313 585
R407 B.n507 B.n506 585
R408 B.n504 B.n314 585
R409 B.n502 B.n501 585
R410 B.n500 B.n315 585
R411 B.n499 B.n498 585
R412 B.n496 B.n316 585
R413 B.n494 B.n493 585
R414 B.n492 B.n317 585
R415 B.n491 B.n490 585
R416 B.n488 B.n487 585
R417 B.n486 B.n485 585
R418 B.n484 B.n322 585
R419 B.n482 B.n481 585
R420 B.n480 B.n323 585
R421 B.n479 B.n478 585
R422 B.n476 B.n324 585
R423 B.n474 B.n473 585
R424 B.n472 B.n325 585
R425 B.n471 B.n470 585
R426 B.n468 B.n467 585
R427 B.n466 B.n465 585
R428 B.n464 B.n330 585
R429 B.n462 B.n461 585
R430 B.n460 B.n331 585
R431 B.n459 B.n458 585
R432 B.n456 B.n332 585
R433 B.n454 B.n453 585
R434 B.n452 B.n333 585
R435 B.n451 B.n450 585
R436 B.n448 B.n334 585
R437 B.n446 B.n445 585
R438 B.n444 B.n335 585
R439 B.n443 B.n442 585
R440 B.n440 B.n336 585
R441 B.n438 B.n437 585
R442 B.n436 B.n337 585
R443 B.n435 B.n434 585
R444 B.n432 B.n338 585
R445 B.n430 B.n429 585
R446 B.n428 B.n339 585
R447 B.n427 B.n426 585
R448 B.n424 B.n340 585
R449 B.n422 B.n421 585
R450 B.n420 B.n341 585
R451 B.n419 B.n418 585
R452 B.n416 B.n342 585
R453 B.n414 B.n413 585
R454 B.n412 B.n343 585
R455 B.n411 B.n410 585
R456 B.n408 B.n344 585
R457 B.n406 B.n405 585
R458 B.n404 B.n345 585
R459 B.n403 B.n402 585
R460 B.n400 B.n346 585
R461 B.n398 B.n397 585
R462 B.n396 B.n347 585
R463 B.n395 B.n394 585
R464 B.n392 B.n348 585
R465 B.n390 B.n389 585
R466 B.n388 B.n349 585
R467 B.n387 B.n386 585
R468 B.n384 B.n350 585
R469 B.n382 B.n381 585
R470 B.n380 B.n351 585
R471 B.n379 B.n378 585
R472 B.n376 B.n352 585
R473 B.n374 B.n373 585
R474 B.n372 B.n353 585
R475 B.n371 B.n370 585
R476 B.n368 B.n354 585
R477 B.n366 B.n365 585
R478 B.n364 B.n355 585
R479 B.n363 B.n362 585
R480 B.n360 B.n356 585
R481 B.n358 B.n357 585
R482 B.n287 B.n286 585
R483 B.n288 B.n287 585
R484 B.n603 B.n602 585
R485 B.n604 B.n603 585
R486 B.n283 B.n282 585
R487 B.n284 B.n283 585
R488 B.n612 B.n611 585
R489 B.n611 B.n610 585
R490 B.n613 B.n281 585
R491 B.n281 B.n280 585
R492 B.n615 B.n614 585
R493 B.n616 B.n615 585
R494 B.n275 B.n274 585
R495 B.n276 B.n275 585
R496 B.n624 B.n623 585
R497 B.n623 B.n622 585
R498 B.n625 B.n273 585
R499 B.n273 B.n271 585
R500 B.n627 B.n626 585
R501 B.n628 B.n627 585
R502 B.n267 B.n266 585
R503 B.n272 B.n267 585
R504 B.n636 B.n635 585
R505 B.n635 B.n634 585
R506 B.n637 B.n265 585
R507 B.n265 B.n264 585
R508 B.n639 B.n638 585
R509 B.n640 B.n639 585
R510 B.n259 B.n258 585
R511 B.n260 B.n259 585
R512 B.n648 B.n647 585
R513 B.n647 B.n646 585
R514 B.n649 B.n257 585
R515 B.n257 B.n256 585
R516 B.n651 B.n650 585
R517 B.n652 B.n651 585
R518 B.n251 B.n250 585
R519 B.n252 B.n251 585
R520 B.n660 B.n659 585
R521 B.n659 B.n658 585
R522 B.n661 B.n249 585
R523 B.n249 B.n248 585
R524 B.n663 B.n662 585
R525 B.n664 B.n663 585
R526 B.n243 B.n242 585
R527 B.n244 B.n243 585
R528 B.n672 B.n671 585
R529 B.n671 B.n670 585
R530 B.n673 B.n241 585
R531 B.n241 B.n239 585
R532 B.n675 B.n674 585
R533 B.n676 B.n675 585
R534 B.n235 B.n234 585
R535 B.n240 B.n235 585
R536 B.n684 B.n683 585
R537 B.n683 B.n682 585
R538 B.n685 B.n233 585
R539 B.n233 B.n232 585
R540 B.n687 B.n686 585
R541 B.n688 B.n687 585
R542 B.n227 B.n226 585
R543 B.n228 B.n227 585
R544 B.n696 B.n695 585
R545 B.n695 B.n694 585
R546 B.n697 B.n225 585
R547 B.n225 B.n224 585
R548 B.n699 B.n698 585
R549 B.n700 B.n699 585
R550 B.n219 B.n218 585
R551 B.n220 B.n219 585
R552 B.n708 B.n707 585
R553 B.n707 B.n706 585
R554 B.n709 B.n217 585
R555 B.n217 B.n215 585
R556 B.n711 B.n710 585
R557 B.n712 B.n711 585
R558 B.n211 B.n210 585
R559 B.n216 B.n211 585
R560 B.n720 B.n719 585
R561 B.n719 B.n718 585
R562 B.n721 B.n209 585
R563 B.n209 B.n208 585
R564 B.n723 B.n722 585
R565 B.n724 B.n723 585
R566 B.n203 B.n202 585
R567 B.n204 B.n203 585
R568 B.n732 B.n731 585
R569 B.n731 B.n730 585
R570 B.n733 B.n201 585
R571 B.n201 B.n200 585
R572 B.n735 B.n734 585
R573 B.n736 B.n735 585
R574 B.n195 B.n194 585
R575 B.n196 B.n195 585
R576 B.n744 B.n743 585
R577 B.n743 B.n742 585
R578 B.n745 B.n193 585
R579 B.n193 B.n192 585
R580 B.n747 B.n746 585
R581 B.n748 B.n747 585
R582 B.n187 B.n186 585
R583 B.n188 B.n187 585
R584 B.n756 B.n755 585
R585 B.n755 B.n754 585
R586 B.n757 B.n185 585
R587 B.n185 B.n184 585
R588 B.n759 B.n758 585
R589 B.n760 B.n759 585
R590 B.n179 B.n178 585
R591 B.n180 B.n179 585
R592 B.n769 B.n768 585
R593 B.n768 B.n767 585
R594 B.n770 B.n177 585
R595 B.n177 B.n176 585
R596 B.n772 B.n771 585
R597 B.n773 B.n772 585
R598 B.n2 B.n0 585
R599 B.n4 B.n2 585
R600 B.n3 B.n1 585
R601 B.n1214 B.n3 585
R602 B.n1212 B.n1211 585
R603 B.n1213 B.n1212 585
R604 B.n1210 B.n9 585
R605 B.n9 B.n8 585
R606 B.n1209 B.n1208 585
R607 B.n1208 B.n1207 585
R608 B.n11 B.n10 585
R609 B.n1206 B.n11 585
R610 B.n1204 B.n1203 585
R611 B.n1205 B.n1204 585
R612 B.n1202 B.n16 585
R613 B.n16 B.n15 585
R614 B.n1201 B.n1200 585
R615 B.n1200 B.n1199 585
R616 B.n18 B.n17 585
R617 B.n1198 B.n18 585
R618 B.n1196 B.n1195 585
R619 B.n1197 B.n1196 585
R620 B.n1194 B.n23 585
R621 B.n23 B.n22 585
R622 B.n1193 B.n1192 585
R623 B.n1192 B.n1191 585
R624 B.n25 B.n24 585
R625 B.n1190 B.n25 585
R626 B.n1188 B.n1187 585
R627 B.n1189 B.n1188 585
R628 B.n1186 B.n30 585
R629 B.n30 B.n29 585
R630 B.n1185 B.n1184 585
R631 B.n1184 B.n1183 585
R632 B.n32 B.n31 585
R633 B.n1182 B.n32 585
R634 B.n1180 B.n1179 585
R635 B.n1181 B.n1180 585
R636 B.n1178 B.n37 585
R637 B.n37 B.n36 585
R638 B.n1177 B.n1176 585
R639 B.n1176 B.n1175 585
R640 B.n39 B.n38 585
R641 B.n1174 B.n39 585
R642 B.n1172 B.n1171 585
R643 B.n1173 B.n1172 585
R644 B.n1170 B.n44 585
R645 B.n44 B.n43 585
R646 B.n1169 B.n1168 585
R647 B.n1168 B.n1167 585
R648 B.n46 B.n45 585
R649 B.n1166 B.n46 585
R650 B.n1164 B.n1163 585
R651 B.n1165 B.n1164 585
R652 B.n1162 B.n51 585
R653 B.n51 B.n50 585
R654 B.n1161 B.n1160 585
R655 B.n1160 B.n1159 585
R656 B.n53 B.n52 585
R657 B.n1158 B.n53 585
R658 B.n1156 B.n1155 585
R659 B.n1157 B.n1156 585
R660 B.n1154 B.n58 585
R661 B.n58 B.n57 585
R662 B.n1153 B.n1152 585
R663 B.n1152 B.n1151 585
R664 B.n60 B.n59 585
R665 B.n1150 B.n60 585
R666 B.n1148 B.n1147 585
R667 B.n1149 B.n1148 585
R668 B.n1146 B.n65 585
R669 B.n65 B.n64 585
R670 B.n1145 B.n1144 585
R671 B.n1144 B.n1143 585
R672 B.n67 B.n66 585
R673 B.n1142 B.n67 585
R674 B.n1140 B.n1139 585
R675 B.n1141 B.n1140 585
R676 B.n1138 B.n72 585
R677 B.n72 B.n71 585
R678 B.n1137 B.n1136 585
R679 B.n1136 B.n1135 585
R680 B.n74 B.n73 585
R681 B.n1134 B.n74 585
R682 B.n1132 B.n1131 585
R683 B.n1133 B.n1132 585
R684 B.n1130 B.n79 585
R685 B.n79 B.n78 585
R686 B.n1129 B.n1128 585
R687 B.n1128 B.n1127 585
R688 B.n81 B.n80 585
R689 B.n1126 B.n81 585
R690 B.n1124 B.n1123 585
R691 B.n1125 B.n1124 585
R692 B.n1122 B.n86 585
R693 B.n86 B.n85 585
R694 B.n1121 B.n1120 585
R695 B.n1120 B.n1119 585
R696 B.n88 B.n87 585
R697 B.n1118 B.n88 585
R698 B.n1116 B.n1115 585
R699 B.n1117 B.n1116 585
R700 B.n1114 B.n93 585
R701 B.n93 B.n92 585
R702 B.n1113 B.n1112 585
R703 B.n1112 B.n1111 585
R704 B.n95 B.n94 585
R705 B.n1110 B.n95 585
R706 B.n1108 B.n1107 585
R707 B.n1109 B.n1108 585
R708 B.n1106 B.n100 585
R709 B.n100 B.n99 585
R710 B.n1105 B.n1104 585
R711 B.n1104 B.n1103 585
R712 B.n102 B.n101 585
R713 B.n1102 B.n102 585
R714 B.n1100 B.n1099 585
R715 B.n1101 B.n1100 585
R716 B.n1217 B.n1216 585
R717 B.n1216 B.n1215 585
R718 B.n603 B.n289 516.524
R719 B.n1100 B.n107 516.524
R720 B.n605 B.n287 516.524
R721 B.n851 B.n105 516.524
R722 B.n326 B.t14 316.305
R723 B.n318 B.t10 316.305
R724 B.n136 B.t17 316.305
R725 B.n144 B.t6 316.305
R726 B.n852 B.n106 256.663
R727 B.n854 B.n106 256.663
R728 B.n860 B.n106 256.663
R729 B.n862 B.n106 256.663
R730 B.n868 B.n106 256.663
R731 B.n870 B.n106 256.663
R732 B.n876 B.n106 256.663
R733 B.n878 B.n106 256.663
R734 B.n884 B.n106 256.663
R735 B.n886 B.n106 256.663
R736 B.n892 B.n106 256.663
R737 B.n894 B.n106 256.663
R738 B.n900 B.n106 256.663
R739 B.n902 B.n106 256.663
R740 B.n908 B.n106 256.663
R741 B.n910 B.n106 256.663
R742 B.n916 B.n106 256.663
R743 B.n918 B.n106 256.663
R744 B.n924 B.n106 256.663
R745 B.n926 B.n106 256.663
R746 B.n932 B.n106 256.663
R747 B.n934 B.n106 256.663
R748 B.n940 B.n106 256.663
R749 B.n942 B.n106 256.663
R750 B.n948 B.n106 256.663
R751 B.n950 B.n106 256.663
R752 B.n956 B.n106 256.663
R753 B.n958 B.n106 256.663
R754 B.n964 B.n106 256.663
R755 B.n966 B.n106 256.663
R756 B.n972 B.n106 256.663
R757 B.n974 B.n106 256.663
R758 B.n980 B.n106 256.663
R759 B.n982 B.n106 256.663
R760 B.n989 B.n106 256.663
R761 B.n991 B.n106 256.663
R762 B.n997 B.n106 256.663
R763 B.n999 B.n106 256.663
R764 B.n1005 B.n106 256.663
R765 B.n1007 B.n106 256.663
R766 B.n1013 B.n106 256.663
R767 B.n1015 B.n106 256.663
R768 B.n1021 B.n106 256.663
R769 B.n1023 B.n106 256.663
R770 B.n1029 B.n106 256.663
R771 B.n1031 B.n106 256.663
R772 B.n1037 B.n106 256.663
R773 B.n1039 B.n106 256.663
R774 B.n1045 B.n106 256.663
R775 B.n1047 B.n106 256.663
R776 B.n1053 B.n106 256.663
R777 B.n1055 B.n106 256.663
R778 B.n1061 B.n106 256.663
R779 B.n1063 B.n106 256.663
R780 B.n1069 B.n106 256.663
R781 B.n1071 B.n106 256.663
R782 B.n1077 B.n106 256.663
R783 B.n1079 B.n106 256.663
R784 B.n1085 B.n106 256.663
R785 B.n1087 B.n106 256.663
R786 B.n1093 B.n106 256.663
R787 B.n1095 B.n106 256.663
R788 B.n598 B.n288 256.663
R789 B.n291 B.n288 256.663
R790 B.n591 B.n288 256.663
R791 B.n585 B.n288 256.663
R792 B.n583 B.n288 256.663
R793 B.n577 B.n288 256.663
R794 B.n575 B.n288 256.663
R795 B.n569 B.n288 256.663
R796 B.n567 B.n288 256.663
R797 B.n561 B.n288 256.663
R798 B.n559 B.n288 256.663
R799 B.n553 B.n288 256.663
R800 B.n551 B.n288 256.663
R801 B.n545 B.n288 256.663
R802 B.n543 B.n288 256.663
R803 B.n537 B.n288 256.663
R804 B.n535 B.n288 256.663
R805 B.n529 B.n288 256.663
R806 B.n527 B.n288 256.663
R807 B.n521 B.n288 256.663
R808 B.n519 B.n288 256.663
R809 B.n513 B.n288 256.663
R810 B.n511 B.n288 256.663
R811 B.n505 B.n288 256.663
R812 B.n503 B.n288 256.663
R813 B.n497 B.n288 256.663
R814 B.n495 B.n288 256.663
R815 B.n489 B.n288 256.663
R816 B.n321 B.n288 256.663
R817 B.n483 B.n288 256.663
R818 B.n477 B.n288 256.663
R819 B.n475 B.n288 256.663
R820 B.n469 B.n288 256.663
R821 B.n329 B.n288 256.663
R822 B.n463 B.n288 256.663
R823 B.n457 B.n288 256.663
R824 B.n455 B.n288 256.663
R825 B.n449 B.n288 256.663
R826 B.n447 B.n288 256.663
R827 B.n441 B.n288 256.663
R828 B.n439 B.n288 256.663
R829 B.n433 B.n288 256.663
R830 B.n431 B.n288 256.663
R831 B.n425 B.n288 256.663
R832 B.n423 B.n288 256.663
R833 B.n417 B.n288 256.663
R834 B.n415 B.n288 256.663
R835 B.n409 B.n288 256.663
R836 B.n407 B.n288 256.663
R837 B.n401 B.n288 256.663
R838 B.n399 B.n288 256.663
R839 B.n393 B.n288 256.663
R840 B.n391 B.n288 256.663
R841 B.n385 B.n288 256.663
R842 B.n383 B.n288 256.663
R843 B.n377 B.n288 256.663
R844 B.n375 B.n288 256.663
R845 B.n369 B.n288 256.663
R846 B.n367 B.n288 256.663
R847 B.n361 B.n288 256.663
R848 B.n359 B.n288 256.663
R849 B.n603 B.n283 163.367
R850 B.n611 B.n283 163.367
R851 B.n611 B.n281 163.367
R852 B.n615 B.n281 163.367
R853 B.n615 B.n275 163.367
R854 B.n623 B.n275 163.367
R855 B.n623 B.n273 163.367
R856 B.n627 B.n273 163.367
R857 B.n627 B.n267 163.367
R858 B.n635 B.n267 163.367
R859 B.n635 B.n265 163.367
R860 B.n639 B.n265 163.367
R861 B.n639 B.n259 163.367
R862 B.n647 B.n259 163.367
R863 B.n647 B.n257 163.367
R864 B.n651 B.n257 163.367
R865 B.n651 B.n251 163.367
R866 B.n659 B.n251 163.367
R867 B.n659 B.n249 163.367
R868 B.n663 B.n249 163.367
R869 B.n663 B.n243 163.367
R870 B.n671 B.n243 163.367
R871 B.n671 B.n241 163.367
R872 B.n675 B.n241 163.367
R873 B.n675 B.n235 163.367
R874 B.n683 B.n235 163.367
R875 B.n683 B.n233 163.367
R876 B.n687 B.n233 163.367
R877 B.n687 B.n227 163.367
R878 B.n695 B.n227 163.367
R879 B.n695 B.n225 163.367
R880 B.n699 B.n225 163.367
R881 B.n699 B.n219 163.367
R882 B.n707 B.n219 163.367
R883 B.n707 B.n217 163.367
R884 B.n711 B.n217 163.367
R885 B.n711 B.n211 163.367
R886 B.n719 B.n211 163.367
R887 B.n719 B.n209 163.367
R888 B.n723 B.n209 163.367
R889 B.n723 B.n203 163.367
R890 B.n731 B.n203 163.367
R891 B.n731 B.n201 163.367
R892 B.n735 B.n201 163.367
R893 B.n735 B.n195 163.367
R894 B.n743 B.n195 163.367
R895 B.n743 B.n193 163.367
R896 B.n747 B.n193 163.367
R897 B.n747 B.n187 163.367
R898 B.n755 B.n187 163.367
R899 B.n755 B.n185 163.367
R900 B.n759 B.n185 163.367
R901 B.n759 B.n179 163.367
R902 B.n768 B.n179 163.367
R903 B.n768 B.n177 163.367
R904 B.n772 B.n177 163.367
R905 B.n772 B.n2 163.367
R906 B.n1216 B.n2 163.367
R907 B.n1216 B.n3 163.367
R908 B.n1212 B.n3 163.367
R909 B.n1212 B.n9 163.367
R910 B.n1208 B.n9 163.367
R911 B.n1208 B.n11 163.367
R912 B.n1204 B.n11 163.367
R913 B.n1204 B.n16 163.367
R914 B.n1200 B.n16 163.367
R915 B.n1200 B.n18 163.367
R916 B.n1196 B.n18 163.367
R917 B.n1196 B.n23 163.367
R918 B.n1192 B.n23 163.367
R919 B.n1192 B.n25 163.367
R920 B.n1188 B.n25 163.367
R921 B.n1188 B.n30 163.367
R922 B.n1184 B.n30 163.367
R923 B.n1184 B.n32 163.367
R924 B.n1180 B.n32 163.367
R925 B.n1180 B.n37 163.367
R926 B.n1176 B.n37 163.367
R927 B.n1176 B.n39 163.367
R928 B.n1172 B.n39 163.367
R929 B.n1172 B.n44 163.367
R930 B.n1168 B.n44 163.367
R931 B.n1168 B.n46 163.367
R932 B.n1164 B.n46 163.367
R933 B.n1164 B.n51 163.367
R934 B.n1160 B.n51 163.367
R935 B.n1160 B.n53 163.367
R936 B.n1156 B.n53 163.367
R937 B.n1156 B.n58 163.367
R938 B.n1152 B.n58 163.367
R939 B.n1152 B.n60 163.367
R940 B.n1148 B.n60 163.367
R941 B.n1148 B.n65 163.367
R942 B.n1144 B.n65 163.367
R943 B.n1144 B.n67 163.367
R944 B.n1140 B.n67 163.367
R945 B.n1140 B.n72 163.367
R946 B.n1136 B.n72 163.367
R947 B.n1136 B.n74 163.367
R948 B.n1132 B.n74 163.367
R949 B.n1132 B.n79 163.367
R950 B.n1128 B.n79 163.367
R951 B.n1128 B.n81 163.367
R952 B.n1124 B.n81 163.367
R953 B.n1124 B.n86 163.367
R954 B.n1120 B.n86 163.367
R955 B.n1120 B.n88 163.367
R956 B.n1116 B.n88 163.367
R957 B.n1116 B.n93 163.367
R958 B.n1112 B.n93 163.367
R959 B.n1112 B.n95 163.367
R960 B.n1108 B.n95 163.367
R961 B.n1108 B.n100 163.367
R962 B.n1104 B.n100 163.367
R963 B.n1104 B.n102 163.367
R964 B.n1100 B.n102 163.367
R965 B.n599 B.n597 163.367
R966 B.n597 B.n596 163.367
R967 B.n593 B.n592 163.367
R968 B.n590 B.n293 163.367
R969 B.n586 B.n584 163.367
R970 B.n582 B.n295 163.367
R971 B.n578 B.n576 163.367
R972 B.n574 B.n297 163.367
R973 B.n570 B.n568 163.367
R974 B.n566 B.n299 163.367
R975 B.n562 B.n560 163.367
R976 B.n558 B.n301 163.367
R977 B.n554 B.n552 163.367
R978 B.n550 B.n303 163.367
R979 B.n546 B.n544 163.367
R980 B.n542 B.n305 163.367
R981 B.n538 B.n536 163.367
R982 B.n534 B.n307 163.367
R983 B.n530 B.n528 163.367
R984 B.n526 B.n309 163.367
R985 B.n522 B.n520 163.367
R986 B.n518 B.n311 163.367
R987 B.n514 B.n512 163.367
R988 B.n510 B.n313 163.367
R989 B.n506 B.n504 163.367
R990 B.n502 B.n315 163.367
R991 B.n498 B.n496 163.367
R992 B.n494 B.n317 163.367
R993 B.n490 B.n488 163.367
R994 B.n485 B.n484 163.367
R995 B.n482 B.n323 163.367
R996 B.n478 B.n476 163.367
R997 B.n474 B.n325 163.367
R998 B.n470 B.n468 163.367
R999 B.n465 B.n464 163.367
R1000 B.n462 B.n331 163.367
R1001 B.n458 B.n456 163.367
R1002 B.n454 B.n333 163.367
R1003 B.n450 B.n448 163.367
R1004 B.n446 B.n335 163.367
R1005 B.n442 B.n440 163.367
R1006 B.n438 B.n337 163.367
R1007 B.n434 B.n432 163.367
R1008 B.n430 B.n339 163.367
R1009 B.n426 B.n424 163.367
R1010 B.n422 B.n341 163.367
R1011 B.n418 B.n416 163.367
R1012 B.n414 B.n343 163.367
R1013 B.n410 B.n408 163.367
R1014 B.n406 B.n345 163.367
R1015 B.n402 B.n400 163.367
R1016 B.n398 B.n347 163.367
R1017 B.n394 B.n392 163.367
R1018 B.n390 B.n349 163.367
R1019 B.n386 B.n384 163.367
R1020 B.n382 B.n351 163.367
R1021 B.n378 B.n376 163.367
R1022 B.n374 B.n353 163.367
R1023 B.n370 B.n368 163.367
R1024 B.n366 B.n355 163.367
R1025 B.n362 B.n360 163.367
R1026 B.n358 B.n287 163.367
R1027 B.n605 B.n285 163.367
R1028 B.n609 B.n285 163.367
R1029 B.n609 B.n279 163.367
R1030 B.n617 B.n279 163.367
R1031 B.n617 B.n277 163.367
R1032 B.n621 B.n277 163.367
R1033 B.n621 B.n270 163.367
R1034 B.n629 B.n270 163.367
R1035 B.n629 B.n268 163.367
R1036 B.n633 B.n268 163.367
R1037 B.n633 B.n263 163.367
R1038 B.n641 B.n263 163.367
R1039 B.n641 B.n261 163.367
R1040 B.n645 B.n261 163.367
R1041 B.n645 B.n255 163.367
R1042 B.n653 B.n255 163.367
R1043 B.n653 B.n253 163.367
R1044 B.n657 B.n253 163.367
R1045 B.n657 B.n247 163.367
R1046 B.n665 B.n247 163.367
R1047 B.n665 B.n245 163.367
R1048 B.n669 B.n245 163.367
R1049 B.n669 B.n238 163.367
R1050 B.n677 B.n238 163.367
R1051 B.n677 B.n236 163.367
R1052 B.n681 B.n236 163.367
R1053 B.n681 B.n231 163.367
R1054 B.n689 B.n231 163.367
R1055 B.n689 B.n229 163.367
R1056 B.n693 B.n229 163.367
R1057 B.n693 B.n223 163.367
R1058 B.n701 B.n223 163.367
R1059 B.n701 B.n221 163.367
R1060 B.n705 B.n221 163.367
R1061 B.n705 B.n214 163.367
R1062 B.n713 B.n214 163.367
R1063 B.n713 B.n212 163.367
R1064 B.n717 B.n212 163.367
R1065 B.n717 B.n207 163.367
R1066 B.n725 B.n207 163.367
R1067 B.n725 B.n205 163.367
R1068 B.n729 B.n205 163.367
R1069 B.n729 B.n199 163.367
R1070 B.n737 B.n199 163.367
R1071 B.n737 B.n197 163.367
R1072 B.n741 B.n197 163.367
R1073 B.n741 B.n191 163.367
R1074 B.n749 B.n191 163.367
R1075 B.n749 B.n189 163.367
R1076 B.n753 B.n189 163.367
R1077 B.n753 B.n183 163.367
R1078 B.n761 B.n183 163.367
R1079 B.n761 B.n181 163.367
R1080 B.n766 B.n181 163.367
R1081 B.n766 B.n175 163.367
R1082 B.n774 B.n175 163.367
R1083 B.n775 B.n774 163.367
R1084 B.n775 B.n5 163.367
R1085 B.n6 B.n5 163.367
R1086 B.n7 B.n6 163.367
R1087 B.n780 B.n7 163.367
R1088 B.n780 B.n12 163.367
R1089 B.n13 B.n12 163.367
R1090 B.n14 B.n13 163.367
R1091 B.n785 B.n14 163.367
R1092 B.n785 B.n19 163.367
R1093 B.n20 B.n19 163.367
R1094 B.n21 B.n20 163.367
R1095 B.n790 B.n21 163.367
R1096 B.n790 B.n26 163.367
R1097 B.n27 B.n26 163.367
R1098 B.n28 B.n27 163.367
R1099 B.n795 B.n28 163.367
R1100 B.n795 B.n33 163.367
R1101 B.n34 B.n33 163.367
R1102 B.n35 B.n34 163.367
R1103 B.n800 B.n35 163.367
R1104 B.n800 B.n40 163.367
R1105 B.n41 B.n40 163.367
R1106 B.n42 B.n41 163.367
R1107 B.n805 B.n42 163.367
R1108 B.n805 B.n47 163.367
R1109 B.n48 B.n47 163.367
R1110 B.n49 B.n48 163.367
R1111 B.n810 B.n49 163.367
R1112 B.n810 B.n54 163.367
R1113 B.n55 B.n54 163.367
R1114 B.n56 B.n55 163.367
R1115 B.n815 B.n56 163.367
R1116 B.n815 B.n61 163.367
R1117 B.n62 B.n61 163.367
R1118 B.n63 B.n62 163.367
R1119 B.n820 B.n63 163.367
R1120 B.n820 B.n68 163.367
R1121 B.n69 B.n68 163.367
R1122 B.n70 B.n69 163.367
R1123 B.n825 B.n70 163.367
R1124 B.n825 B.n75 163.367
R1125 B.n76 B.n75 163.367
R1126 B.n77 B.n76 163.367
R1127 B.n830 B.n77 163.367
R1128 B.n830 B.n82 163.367
R1129 B.n83 B.n82 163.367
R1130 B.n84 B.n83 163.367
R1131 B.n835 B.n84 163.367
R1132 B.n835 B.n89 163.367
R1133 B.n90 B.n89 163.367
R1134 B.n91 B.n90 163.367
R1135 B.n840 B.n91 163.367
R1136 B.n840 B.n96 163.367
R1137 B.n97 B.n96 163.367
R1138 B.n98 B.n97 163.367
R1139 B.n845 B.n98 163.367
R1140 B.n845 B.n103 163.367
R1141 B.n104 B.n103 163.367
R1142 B.n105 B.n104 163.367
R1143 B.n1096 B.n1094 163.367
R1144 B.n1092 B.n109 163.367
R1145 B.n1088 B.n1086 163.367
R1146 B.n1084 B.n111 163.367
R1147 B.n1080 B.n1078 163.367
R1148 B.n1076 B.n113 163.367
R1149 B.n1072 B.n1070 163.367
R1150 B.n1068 B.n115 163.367
R1151 B.n1064 B.n1062 163.367
R1152 B.n1060 B.n117 163.367
R1153 B.n1056 B.n1054 163.367
R1154 B.n1052 B.n119 163.367
R1155 B.n1048 B.n1046 163.367
R1156 B.n1044 B.n121 163.367
R1157 B.n1040 B.n1038 163.367
R1158 B.n1036 B.n123 163.367
R1159 B.n1032 B.n1030 163.367
R1160 B.n1028 B.n125 163.367
R1161 B.n1024 B.n1022 163.367
R1162 B.n1020 B.n127 163.367
R1163 B.n1016 B.n1014 163.367
R1164 B.n1012 B.n129 163.367
R1165 B.n1008 B.n1006 163.367
R1166 B.n1004 B.n131 163.367
R1167 B.n1000 B.n998 163.367
R1168 B.n996 B.n133 163.367
R1169 B.n992 B.n990 163.367
R1170 B.n988 B.n135 163.367
R1171 B.n983 B.n981 163.367
R1172 B.n979 B.n139 163.367
R1173 B.n975 B.n973 163.367
R1174 B.n971 B.n141 163.367
R1175 B.n967 B.n965 163.367
R1176 B.n963 B.n143 163.367
R1177 B.n959 B.n957 163.367
R1178 B.n955 B.n148 163.367
R1179 B.n951 B.n949 163.367
R1180 B.n947 B.n150 163.367
R1181 B.n943 B.n941 163.367
R1182 B.n939 B.n152 163.367
R1183 B.n935 B.n933 163.367
R1184 B.n931 B.n154 163.367
R1185 B.n927 B.n925 163.367
R1186 B.n923 B.n156 163.367
R1187 B.n919 B.n917 163.367
R1188 B.n915 B.n158 163.367
R1189 B.n911 B.n909 163.367
R1190 B.n907 B.n160 163.367
R1191 B.n903 B.n901 163.367
R1192 B.n899 B.n162 163.367
R1193 B.n895 B.n893 163.367
R1194 B.n891 B.n164 163.367
R1195 B.n887 B.n885 163.367
R1196 B.n883 B.n166 163.367
R1197 B.n879 B.n877 163.367
R1198 B.n875 B.n168 163.367
R1199 B.n871 B.n869 163.367
R1200 B.n867 B.n170 163.367
R1201 B.n863 B.n861 163.367
R1202 B.n859 B.n172 163.367
R1203 B.n855 B.n853 163.367
R1204 B.n326 B.t16 156.113
R1205 B.n144 B.t8 156.113
R1206 B.n318 B.t13 156.09
R1207 B.n136 B.t18 156.09
R1208 B.n327 B.n326 82.2308
R1209 B.n319 B.n318 82.2308
R1210 B.n137 B.n136 82.2308
R1211 B.n145 B.n144 82.2308
R1212 B.n327 B.t15 73.8832
R1213 B.n145 B.t9 73.8832
R1214 B.n319 B.t12 73.8605
R1215 B.n137 B.t19 73.8605
R1216 B.n598 B.n289 71.676
R1217 B.n596 B.n291 71.676
R1218 B.n592 B.n591 71.676
R1219 B.n585 B.n293 71.676
R1220 B.n584 B.n583 71.676
R1221 B.n577 B.n295 71.676
R1222 B.n576 B.n575 71.676
R1223 B.n569 B.n297 71.676
R1224 B.n568 B.n567 71.676
R1225 B.n561 B.n299 71.676
R1226 B.n560 B.n559 71.676
R1227 B.n553 B.n301 71.676
R1228 B.n552 B.n551 71.676
R1229 B.n545 B.n303 71.676
R1230 B.n544 B.n543 71.676
R1231 B.n537 B.n305 71.676
R1232 B.n536 B.n535 71.676
R1233 B.n529 B.n307 71.676
R1234 B.n528 B.n527 71.676
R1235 B.n521 B.n309 71.676
R1236 B.n520 B.n519 71.676
R1237 B.n513 B.n311 71.676
R1238 B.n512 B.n511 71.676
R1239 B.n505 B.n313 71.676
R1240 B.n504 B.n503 71.676
R1241 B.n497 B.n315 71.676
R1242 B.n496 B.n495 71.676
R1243 B.n489 B.n317 71.676
R1244 B.n488 B.n321 71.676
R1245 B.n484 B.n483 71.676
R1246 B.n477 B.n323 71.676
R1247 B.n476 B.n475 71.676
R1248 B.n469 B.n325 71.676
R1249 B.n468 B.n329 71.676
R1250 B.n464 B.n463 71.676
R1251 B.n457 B.n331 71.676
R1252 B.n456 B.n455 71.676
R1253 B.n449 B.n333 71.676
R1254 B.n448 B.n447 71.676
R1255 B.n441 B.n335 71.676
R1256 B.n440 B.n439 71.676
R1257 B.n433 B.n337 71.676
R1258 B.n432 B.n431 71.676
R1259 B.n425 B.n339 71.676
R1260 B.n424 B.n423 71.676
R1261 B.n417 B.n341 71.676
R1262 B.n416 B.n415 71.676
R1263 B.n409 B.n343 71.676
R1264 B.n408 B.n407 71.676
R1265 B.n401 B.n345 71.676
R1266 B.n400 B.n399 71.676
R1267 B.n393 B.n347 71.676
R1268 B.n392 B.n391 71.676
R1269 B.n385 B.n349 71.676
R1270 B.n384 B.n383 71.676
R1271 B.n377 B.n351 71.676
R1272 B.n376 B.n375 71.676
R1273 B.n369 B.n353 71.676
R1274 B.n368 B.n367 71.676
R1275 B.n361 B.n355 71.676
R1276 B.n360 B.n359 71.676
R1277 B.n1095 B.n107 71.676
R1278 B.n1094 B.n1093 71.676
R1279 B.n1087 B.n109 71.676
R1280 B.n1086 B.n1085 71.676
R1281 B.n1079 B.n111 71.676
R1282 B.n1078 B.n1077 71.676
R1283 B.n1071 B.n113 71.676
R1284 B.n1070 B.n1069 71.676
R1285 B.n1063 B.n115 71.676
R1286 B.n1062 B.n1061 71.676
R1287 B.n1055 B.n117 71.676
R1288 B.n1054 B.n1053 71.676
R1289 B.n1047 B.n119 71.676
R1290 B.n1046 B.n1045 71.676
R1291 B.n1039 B.n121 71.676
R1292 B.n1038 B.n1037 71.676
R1293 B.n1031 B.n123 71.676
R1294 B.n1030 B.n1029 71.676
R1295 B.n1023 B.n125 71.676
R1296 B.n1022 B.n1021 71.676
R1297 B.n1015 B.n127 71.676
R1298 B.n1014 B.n1013 71.676
R1299 B.n1007 B.n129 71.676
R1300 B.n1006 B.n1005 71.676
R1301 B.n999 B.n131 71.676
R1302 B.n998 B.n997 71.676
R1303 B.n991 B.n133 71.676
R1304 B.n990 B.n989 71.676
R1305 B.n982 B.n135 71.676
R1306 B.n981 B.n980 71.676
R1307 B.n974 B.n139 71.676
R1308 B.n973 B.n972 71.676
R1309 B.n966 B.n141 71.676
R1310 B.n965 B.n964 71.676
R1311 B.n958 B.n143 71.676
R1312 B.n957 B.n956 71.676
R1313 B.n950 B.n148 71.676
R1314 B.n949 B.n948 71.676
R1315 B.n942 B.n150 71.676
R1316 B.n941 B.n940 71.676
R1317 B.n934 B.n152 71.676
R1318 B.n933 B.n932 71.676
R1319 B.n926 B.n154 71.676
R1320 B.n925 B.n924 71.676
R1321 B.n918 B.n156 71.676
R1322 B.n917 B.n916 71.676
R1323 B.n910 B.n158 71.676
R1324 B.n909 B.n908 71.676
R1325 B.n902 B.n160 71.676
R1326 B.n901 B.n900 71.676
R1327 B.n894 B.n162 71.676
R1328 B.n893 B.n892 71.676
R1329 B.n886 B.n164 71.676
R1330 B.n885 B.n884 71.676
R1331 B.n878 B.n166 71.676
R1332 B.n877 B.n876 71.676
R1333 B.n870 B.n168 71.676
R1334 B.n869 B.n868 71.676
R1335 B.n862 B.n170 71.676
R1336 B.n861 B.n860 71.676
R1337 B.n854 B.n172 71.676
R1338 B.n853 B.n852 71.676
R1339 B.n852 B.n851 71.676
R1340 B.n855 B.n854 71.676
R1341 B.n860 B.n859 71.676
R1342 B.n863 B.n862 71.676
R1343 B.n868 B.n867 71.676
R1344 B.n871 B.n870 71.676
R1345 B.n876 B.n875 71.676
R1346 B.n879 B.n878 71.676
R1347 B.n884 B.n883 71.676
R1348 B.n887 B.n886 71.676
R1349 B.n892 B.n891 71.676
R1350 B.n895 B.n894 71.676
R1351 B.n900 B.n899 71.676
R1352 B.n903 B.n902 71.676
R1353 B.n908 B.n907 71.676
R1354 B.n911 B.n910 71.676
R1355 B.n916 B.n915 71.676
R1356 B.n919 B.n918 71.676
R1357 B.n924 B.n923 71.676
R1358 B.n927 B.n926 71.676
R1359 B.n932 B.n931 71.676
R1360 B.n935 B.n934 71.676
R1361 B.n940 B.n939 71.676
R1362 B.n943 B.n942 71.676
R1363 B.n948 B.n947 71.676
R1364 B.n951 B.n950 71.676
R1365 B.n956 B.n955 71.676
R1366 B.n959 B.n958 71.676
R1367 B.n964 B.n963 71.676
R1368 B.n967 B.n966 71.676
R1369 B.n972 B.n971 71.676
R1370 B.n975 B.n974 71.676
R1371 B.n980 B.n979 71.676
R1372 B.n983 B.n982 71.676
R1373 B.n989 B.n988 71.676
R1374 B.n992 B.n991 71.676
R1375 B.n997 B.n996 71.676
R1376 B.n1000 B.n999 71.676
R1377 B.n1005 B.n1004 71.676
R1378 B.n1008 B.n1007 71.676
R1379 B.n1013 B.n1012 71.676
R1380 B.n1016 B.n1015 71.676
R1381 B.n1021 B.n1020 71.676
R1382 B.n1024 B.n1023 71.676
R1383 B.n1029 B.n1028 71.676
R1384 B.n1032 B.n1031 71.676
R1385 B.n1037 B.n1036 71.676
R1386 B.n1040 B.n1039 71.676
R1387 B.n1045 B.n1044 71.676
R1388 B.n1048 B.n1047 71.676
R1389 B.n1053 B.n1052 71.676
R1390 B.n1056 B.n1055 71.676
R1391 B.n1061 B.n1060 71.676
R1392 B.n1064 B.n1063 71.676
R1393 B.n1069 B.n1068 71.676
R1394 B.n1072 B.n1071 71.676
R1395 B.n1077 B.n1076 71.676
R1396 B.n1080 B.n1079 71.676
R1397 B.n1085 B.n1084 71.676
R1398 B.n1088 B.n1087 71.676
R1399 B.n1093 B.n1092 71.676
R1400 B.n1096 B.n1095 71.676
R1401 B.n599 B.n598 71.676
R1402 B.n593 B.n291 71.676
R1403 B.n591 B.n590 71.676
R1404 B.n586 B.n585 71.676
R1405 B.n583 B.n582 71.676
R1406 B.n578 B.n577 71.676
R1407 B.n575 B.n574 71.676
R1408 B.n570 B.n569 71.676
R1409 B.n567 B.n566 71.676
R1410 B.n562 B.n561 71.676
R1411 B.n559 B.n558 71.676
R1412 B.n554 B.n553 71.676
R1413 B.n551 B.n550 71.676
R1414 B.n546 B.n545 71.676
R1415 B.n543 B.n542 71.676
R1416 B.n538 B.n537 71.676
R1417 B.n535 B.n534 71.676
R1418 B.n530 B.n529 71.676
R1419 B.n527 B.n526 71.676
R1420 B.n522 B.n521 71.676
R1421 B.n519 B.n518 71.676
R1422 B.n514 B.n513 71.676
R1423 B.n511 B.n510 71.676
R1424 B.n506 B.n505 71.676
R1425 B.n503 B.n502 71.676
R1426 B.n498 B.n497 71.676
R1427 B.n495 B.n494 71.676
R1428 B.n490 B.n489 71.676
R1429 B.n485 B.n321 71.676
R1430 B.n483 B.n482 71.676
R1431 B.n478 B.n477 71.676
R1432 B.n475 B.n474 71.676
R1433 B.n470 B.n469 71.676
R1434 B.n465 B.n329 71.676
R1435 B.n463 B.n462 71.676
R1436 B.n458 B.n457 71.676
R1437 B.n455 B.n454 71.676
R1438 B.n450 B.n449 71.676
R1439 B.n447 B.n446 71.676
R1440 B.n442 B.n441 71.676
R1441 B.n439 B.n438 71.676
R1442 B.n434 B.n433 71.676
R1443 B.n431 B.n430 71.676
R1444 B.n426 B.n425 71.676
R1445 B.n423 B.n422 71.676
R1446 B.n418 B.n417 71.676
R1447 B.n415 B.n414 71.676
R1448 B.n410 B.n409 71.676
R1449 B.n407 B.n406 71.676
R1450 B.n402 B.n401 71.676
R1451 B.n399 B.n398 71.676
R1452 B.n394 B.n393 71.676
R1453 B.n391 B.n390 71.676
R1454 B.n386 B.n385 71.676
R1455 B.n383 B.n382 71.676
R1456 B.n378 B.n377 71.676
R1457 B.n375 B.n374 71.676
R1458 B.n370 B.n369 71.676
R1459 B.n367 B.n366 71.676
R1460 B.n362 B.n361 71.676
R1461 B.n359 B.n358 71.676
R1462 B.n604 B.n288 59.828
R1463 B.n1101 B.n106 59.828
R1464 B.n328 B.n327 59.5399
R1465 B.n320 B.n319 59.5399
R1466 B.n985 B.n137 59.5399
R1467 B.n146 B.n145 59.5399
R1468 B.n1099 B.n1098 33.5615
R1469 B.n850 B.n849 33.5615
R1470 B.n606 B.n286 33.5615
R1471 B.n602 B.n601 33.5615
R1472 B.n604 B.n284 33.0759
R1473 B.n610 B.n284 33.0759
R1474 B.n610 B.n280 33.0759
R1475 B.n616 B.n280 33.0759
R1476 B.n616 B.n276 33.0759
R1477 B.n622 B.n276 33.0759
R1478 B.n622 B.n271 33.0759
R1479 B.n628 B.n271 33.0759
R1480 B.n628 B.n272 33.0759
R1481 B.n634 B.n264 33.0759
R1482 B.n640 B.n264 33.0759
R1483 B.n640 B.n260 33.0759
R1484 B.n646 B.n260 33.0759
R1485 B.n646 B.n256 33.0759
R1486 B.n652 B.n256 33.0759
R1487 B.n652 B.n252 33.0759
R1488 B.n658 B.n252 33.0759
R1489 B.n658 B.n248 33.0759
R1490 B.n664 B.n248 33.0759
R1491 B.n664 B.n244 33.0759
R1492 B.n670 B.n244 33.0759
R1493 B.n670 B.n239 33.0759
R1494 B.n676 B.n239 33.0759
R1495 B.n676 B.n240 33.0759
R1496 B.n682 B.n232 33.0759
R1497 B.n688 B.n232 33.0759
R1498 B.n688 B.n228 33.0759
R1499 B.n694 B.n228 33.0759
R1500 B.n694 B.n224 33.0759
R1501 B.n700 B.n224 33.0759
R1502 B.n700 B.n220 33.0759
R1503 B.n706 B.n220 33.0759
R1504 B.n706 B.n215 33.0759
R1505 B.n712 B.n215 33.0759
R1506 B.n712 B.n216 33.0759
R1507 B.n718 B.n208 33.0759
R1508 B.n724 B.n208 33.0759
R1509 B.n724 B.n204 33.0759
R1510 B.n730 B.n204 33.0759
R1511 B.n730 B.n200 33.0759
R1512 B.n736 B.n200 33.0759
R1513 B.n736 B.n196 33.0759
R1514 B.n742 B.n196 33.0759
R1515 B.n742 B.n192 33.0759
R1516 B.n748 B.n192 33.0759
R1517 B.n748 B.n188 33.0759
R1518 B.n754 B.n188 33.0759
R1519 B.n760 B.n184 33.0759
R1520 B.n760 B.n180 33.0759
R1521 B.n767 B.n180 33.0759
R1522 B.n767 B.n176 33.0759
R1523 B.n773 B.n176 33.0759
R1524 B.n773 B.n4 33.0759
R1525 B.n1215 B.n4 33.0759
R1526 B.n1215 B.n1214 33.0759
R1527 B.n1214 B.n1213 33.0759
R1528 B.n1213 B.n8 33.0759
R1529 B.n1207 B.n8 33.0759
R1530 B.n1207 B.n1206 33.0759
R1531 B.n1206 B.n1205 33.0759
R1532 B.n1205 B.n15 33.0759
R1533 B.n1199 B.n1198 33.0759
R1534 B.n1198 B.n1197 33.0759
R1535 B.n1197 B.n22 33.0759
R1536 B.n1191 B.n22 33.0759
R1537 B.n1191 B.n1190 33.0759
R1538 B.n1190 B.n1189 33.0759
R1539 B.n1189 B.n29 33.0759
R1540 B.n1183 B.n29 33.0759
R1541 B.n1183 B.n1182 33.0759
R1542 B.n1182 B.n1181 33.0759
R1543 B.n1181 B.n36 33.0759
R1544 B.n1175 B.n36 33.0759
R1545 B.n1174 B.n1173 33.0759
R1546 B.n1173 B.n43 33.0759
R1547 B.n1167 B.n43 33.0759
R1548 B.n1167 B.n1166 33.0759
R1549 B.n1166 B.n1165 33.0759
R1550 B.n1165 B.n50 33.0759
R1551 B.n1159 B.n50 33.0759
R1552 B.n1159 B.n1158 33.0759
R1553 B.n1158 B.n1157 33.0759
R1554 B.n1157 B.n57 33.0759
R1555 B.n1151 B.n57 33.0759
R1556 B.n1150 B.n1149 33.0759
R1557 B.n1149 B.n64 33.0759
R1558 B.n1143 B.n64 33.0759
R1559 B.n1143 B.n1142 33.0759
R1560 B.n1142 B.n1141 33.0759
R1561 B.n1141 B.n71 33.0759
R1562 B.n1135 B.n71 33.0759
R1563 B.n1135 B.n1134 33.0759
R1564 B.n1134 B.n1133 33.0759
R1565 B.n1133 B.n78 33.0759
R1566 B.n1127 B.n78 33.0759
R1567 B.n1127 B.n1126 33.0759
R1568 B.n1126 B.n1125 33.0759
R1569 B.n1125 B.n85 33.0759
R1570 B.n1119 B.n85 33.0759
R1571 B.n1118 B.n1117 33.0759
R1572 B.n1117 B.n92 33.0759
R1573 B.n1111 B.n92 33.0759
R1574 B.n1111 B.n1110 33.0759
R1575 B.n1110 B.n1109 33.0759
R1576 B.n1109 B.n99 33.0759
R1577 B.n1103 B.n99 33.0759
R1578 B.n1103 B.n1102 33.0759
R1579 B.n1102 B.n1101 33.0759
R1580 B.t2 B.n184 27.7255
R1581 B.t1 B.n15 27.7255
R1582 B.n682 B.t3 25.7799
R1583 B.n1151 B.t0 25.7799
R1584 B.n216 B.t5 22.8614
R1585 B.t4 B.n1174 22.8614
R1586 B B.n1217 18.0485
R1587 B.n272 B.t11 17.9974
R1588 B.t7 B.n1118 17.9974
R1589 B.n634 B.t11 15.079
R1590 B.n1119 B.t7 15.079
R1591 B.n1098 B.n1097 10.6151
R1592 B.n1097 B.n108 10.6151
R1593 B.n1091 B.n108 10.6151
R1594 B.n1091 B.n1090 10.6151
R1595 B.n1090 B.n1089 10.6151
R1596 B.n1089 B.n110 10.6151
R1597 B.n1083 B.n110 10.6151
R1598 B.n1083 B.n1082 10.6151
R1599 B.n1082 B.n1081 10.6151
R1600 B.n1081 B.n112 10.6151
R1601 B.n1075 B.n112 10.6151
R1602 B.n1075 B.n1074 10.6151
R1603 B.n1074 B.n1073 10.6151
R1604 B.n1073 B.n114 10.6151
R1605 B.n1067 B.n114 10.6151
R1606 B.n1067 B.n1066 10.6151
R1607 B.n1066 B.n1065 10.6151
R1608 B.n1065 B.n116 10.6151
R1609 B.n1059 B.n116 10.6151
R1610 B.n1059 B.n1058 10.6151
R1611 B.n1058 B.n1057 10.6151
R1612 B.n1057 B.n118 10.6151
R1613 B.n1051 B.n118 10.6151
R1614 B.n1051 B.n1050 10.6151
R1615 B.n1050 B.n1049 10.6151
R1616 B.n1049 B.n120 10.6151
R1617 B.n1043 B.n120 10.6151
R1618 B.n1043 B.n1042 10.6151
R1619 B.n1042 B.n1041 10.6151
R1620 B.n1041 B.n122 10.6151
R1621 B.n1035 B.n122 10.6151
R1622 B.n1035 B.n1034 10.6151
R1623 B.n1034 B.n1033 10.6151
R1624 B.n1033 B.n124 10.6151
R1625 B.n1027 B.n124 10.6151
R1626 B.n1027 B.n1026 10.6151
R1627 B.n1026 B.n1025 10.6151
R1628 B.n1025 B.n126 10.6151
R1629 B.n1019 B.n126 10.6151
R1630 B.n1019 B.n1018 10.6151
R1631 B.n1018 B.n1017 10.6151
R1632 B.n1017 B.n128 10.6151
R1633 B.n1011 B.n128 10.6151
R1634 B.n1011 B.n1010 10.6151
R1635 B.n1010 B.n1009 10.6151
R1636 B.n1009 B.n130 10.6151
R1637 B.n1003 B.n130 10.6151
R1638 B.n1003 B.n1002 10.6151
R1639 B.n1002 B.n1001 10.6151
R1640 B.n1001 B.n132 10.6151
R1641 B.n995 B.n132 10.6151
R1642 B.n995 B.n994 10.6151
R1643 B.n994 B.n993 10.6151
R1644 B.n993 B.n134 10.6151
R1645 B.n987 B.n134 10.6151
R1646 B.n987 B.n986 10.6151
R1647 B.n984 B.n138 10.6151
R1648 B.n978 B.n138 10.6151
R1649 B.n978 B.n977 10.6151
R1650 B.n977 B.n976 10.6151
R1651 B.n976 B.n140 10.6151
R1652 B.n970 B.n140 10.6151
R1653 B.n970 B.n969 10.6151
R1654 B.n969 B.n968 10.6151
R1655 B.n968 B.n142 10.6151
R1656 B.n962 B.n961 10.6151
R1657 B.n961 B.n960 10.6151
R1658 B.n960 B.n147 10.6151
R1659 B.n954 B.n147 10.6151
R1660 B.n954 B.n953 10.6151
R1661 B.n953 B.n952 10.6151
R1662 B.n952 B.n149 10.6151
R1663 B.n946 B.n149 10.6151
R1664 B.n946 B.n945 10.6151
R1665 B.n945 B.n944 10.6151
R1666 B.n944 B.n151 10.6151
R1667 B.n938 B.n151 10.6151
R1668 B.n938 B.n937 10.6151
R1669 B.n937 B.n936 10.6151
R1670 B.n936 B.n153 10.6151
R1671 B.n930 B.n153 10.6151
R1672 B.n930 B.n929 10.6151
R1673 B.n929 B.n928 10.6151
R1674 B.n928 B.n155 10.6151
R1675 B.n922 B.n155 10.6151
R1676 B.n922 B.n921 10.6151
R1677 B.n921 B.n920 10.6151
R1678 B.n920 B.n157 10.6151
R1679 B.n914 B.n157 10.6151
R1680 B.n914 B.n913 10.6151
R1681 B.n913 B.n912 10.6151
R1682 B.n912 B.n159 10.6151
R1683 B.n906 B.n159 10.6151
R1684 B.n906 B.n905 10.6151
R1685 B.n905 B.n904 10.6151
R1686 B.n904 B.n161 10.6151
R1687 B.n898 B.n161 10.6151
R1688 B.n898 B.n897 10.6151
R1689 B.n897 B.n896 10.6151
R1690 B.n896 B.n163 10.6151
R1691 B.n890 B.n163 10.6151
R1692 B.n890 B.n889 10.6151
R1693 B.n889 B.n888 10.6151
R1694 B.n888 B.n165 10.6151
R1695 B.n882 B.n165 10.6151
R1696 B.n882 B.n881 10.6151
R1697 B.n881 B.n880 10.6151
R1698 B.n880 B.n167 10.6151
R1699 B.n874 B.n167 10.6151
R1700 B.n874 B.n873 10.6151
R1701 B.n873 B.n872 10.6151
R1702 B.n872 B.n169 10.6151
R1703 B.n866 B.n169 10.6151
R1704 B.n866 B.n865 10.6151
R1705 B.n865 B.n864 10.6151
R1706 B.n864 B.n171 10.6151
R1707 B.n858 B.n171 10.6151
R1708 B.n858 B.n857 10.6151
R1709 B.n857 B.n856 10.6151
R1710 B.n856 B.n173 10.6151
R1711 B.n850 B.n173 10.6151
R1712 B.n607 B.n606 10.6151
R1713 B.n608 B.n607 10.6151
R1714 B.n608 B.n278 10.6151
R1715 B.n618 B.n278 10.6151
R1716 B.n619 B.n618 10.6151
R1717 B.n620 B.n619 10.6151
R1718 B.n620 B.n269 10.6151
R1719 B.n630 B.n269 10.6151
R1720 B.n631 B.n630 10.6151
R1721 B.n632 B.n631 10.6151
R1722 B.n632 B.n262 10.6151
R1723 B.n642 B.n262 10.6151
R1724 B.n643 B.n642 10.6151
R1725 B.n644 B.n643 10.6151
R1726 B.n644 B.n254 10.6151
R1727 B.n654 B.n254 10.6151
R1728 B.n655 B.n654 10.6151
R1729 B.n656 B.n655 10.6151
R1730 B.n656 B.n246 10.6151
R1731 B.n666 B.n246 10.6151
R1732 B.n667 B.n666 10.6151
R1733 B.n668 B.n667 10.6151
R1734 B.n668 B.n237 10.6151
R1735 B.n678 B.n237 10.6151
R1736 B.n679 B.n678 10.6151
R1737 B.n680 B.n679 10.6151
R1738 B.n680 B.n230 10.6151
R1739 B.n690 B.n230 10.6151
R1740 B.n691 B.n690 10.6151
R1741 B.n692 B.n691 10.6151
R1742 B.n692 B.n222 10.6151
R1743 B.n702 B.n222 10.6151
R1744 B.n703 B.n702 10.6151
R1745 B.n704 B.n703 10.6151
R1746 B.n704 B.n213 10.6151
R1747 B.n714 B.n213 10.6151
R1748 B.n715 B.n714 10.6151
R1749 B.n716 B.n715 10.6151
R1750 B.n716 B.n206 10.6151
R1751 B.n726 B.n206 10.6151
R1752 B.n727 B.n726 10.6151
R1753 B.n728 B.n727 10.6151
R1754 B.n728 B.n198 10.6151
R1755 B.n738 B.n198 10.6151
R1756 B.n739 B.n738 10.6151
R1757 B.n740 B.n739 10.6151
R1758 B.n740 B.n190 10.6151
R1759 B.n750 B.n190 10.6151
R1760 B.n751 B.n750 10.6151
R1761 B.n752 B.n751 10.6151
R1762 B.n752 B.n182 10.6151
R1763 B.n762 B.n182 10.6151
R1764 B.n763 B.n762 10.6151
R1765 B.n765 B.n763 10.6151
R1766 B.n765 B.n764 10.6151
R1767 B.n764 B.n174 10.6151
R1768 B.n776 B.n174 10.6151
R1769 B.n777 B.n776 10.6151
R1770 B.n778 B.n777 10.6151
R1771 B.n779 B.n778 10.6151
R1772 B.n781 B.n779 10.6151
R1773 B.n782 B.n781 10.6151
R1774 B.n783 B.n782 10.6151
R1775 B.n784 B.n783 10.6151
R1776 B.n786 B.n784 10.6151
R1777 B.n787 B.n786 10.6151
R1778 B.n788 B.n787 10.6151
R1779 B.n789 B.n788 10.6151
R1780 B.n791 B.n789 10.6151
R1781 B.n792 B.n791 10.6151
R1782 B.n793 B.n792 10.6151
R1783 B.n794 B.n793 10.6151
R1784 B.n796 B.n794 10.6151
R1785 B.n797 B.n796 10.6151
R1786 B.n798 B.n797 10.6151
R1787 B.n799 B.n798 10.6151
R1788 B.n801 B.n799 10.6151
R1789 B.n802 B.n801 10.6151
R1790 B.n803 B.n802 10.6151
R1791 B.n804 B.n803 10.6151
R1792 B.n806 B.n804 10.6151
R1793 B.n807 B.n806 10.6151
R1794 B.n808 B.n807 10.6151
R1795 B.n809 B.n808 10.6151
R1796 B.n811 B.n809 10.6151
R1797 B.n812 B.n811 10.6151
R1798 B.n813 B.n812 10.6151
R1799 B.n814 B.n813 10.6151
R1800 B.n816 B.n814 10.6151
R1801 B.n817 B.n816 10.6151
R1802 B.n818 B.n817 10.6151
R1803 B.n819 B.n818 10.6151
R1804 B.n821 B.n819 10.6151
R1805 B.n822 B.n821 10.6151
R1806 B.n823 B.n822 10.6151
R1807 B.n824 B.n823 10.6151
R1808 B.n826 B.n824 10.6151
R1809 B.n827 B.n826 10.6151
R1810 B.n828 B.n827 10.6151
R1811 B.n829 B.n828 10.6151
R1812 B.n831 B.n829 10.6151
R1813 B.n832 B.n831 10.6151
R1814 B.n833 B.n832 10.6151
R1815 B.n834 B.n833 10.6151
R1816 B.n836 B.n834 10.6151
R1817 B.n837 B.n836 10.6151
R1818 B.n838 B.n837 10.6151
R1819 B.n839 B.n838 10.6151
R1820 B.n841 B.n839 10.6151
R1821 B.n842 B.n841 10.6151
R1822 B.n843 B.n842 10.6151
R1823 B.n844 B.n843 10.6151
R1824 B.n846 B.n844 10.6151
R1825 B.n847 B.n846 10.6151
R1826 B.n848 B.n847 10.6151
R1827 B.n849 B.n848 10.6151
R1828 B.n601 B.n600 10.6151
R1829 B.n600 B.n290 10.6151
R1830 B.n595 B.n290 10.6151
R1831 B.n595 B.n594 10.6151
R1832 B.n594 B.n292 10.6151
R1833 B.n589 B.n292 10.6151
R1834 B.n589 B.n588 10.6151
R1835 B.n588 B.n587 10.6151
R1836 B.n587 B.n294 10.6151
R1837 B.n581 B.n294 10.6151
R1838 B.n581 B.n580 10.6151
R1839 B.n580 B.n579 10.6151
R1840 B.n579 B.n296 10.6151
R1841 B.n573 B.n296 10.6151
R1842 B.n573 B.n572 10.6151
R1843 B.n572 B.n571 10.6151
R1844 B.n571 B.n298 10.6151
R1845 B.n565 B.n298 10.6151
R1846 B.n565 B.n564 10.6151
R1847 B.n564 B.n563 10.6151
R1848 B.n563 B.n300 10.6151
R1849 B.n557 B.n300 10.6151
R1850 B.n557 B.n556 10.6151
R1851 B.n556 B.n555 10.6151
R1852 B.n555 B.n302 10.6151
R1853 B.n549 B.n302 10.6151
R1854 B.n549 B.n548 10.6151
R1855 B.n548 B.n547 10.6151
R1856 B.n547 B.n304 10.6151
R1857 B.n541 B.n304 10.6151
R1858 B.n541 B.n540 10.6151
R1859 B.n540 B.n539 10.6151
R1860 B.n539 B.n306 10.6151
R1861 B.n533 B.n306 10.6151
R1862 B.n533 B.n532 10.6151
R1863 B.n532 B.n531 10.6151
R1864 B.n531 B.n308 10.6151
R1865 B.n525 B.n308 10.6151
R1866 B.n525 B.n524 10.6151
R1867 B.n524 B.n523 10.6151
R1868 B.n523 B.n310 10.6151
R1869 B.n517 B.n310 10.6151
R1870 B.n517 B.n516 10.6151
R1871 B.n516 B.n515 10.6151
R1872 B.n515 B.n312 10.6151
R1873 B.n509 B.n312 10.6151
R1874 B.n509 B.n508 10.6151
R1875 B.n508 B.n507 10.6151
R1876 B.n507 B.n314 10.6151
R1877 B.n501 B.n314 10.6151
R1878 B.n501 B.n500 10.6151
R1879 B.n500 B.n499 10.6151
R1880 B.n499 B.n316 10.6151
R1881 B.n493 B.n316 10.6151
R1882 B.n493 B.n492 10.6151
R1883 B.n492 B.n491 10.6151
R1884 B.n487 B.n486 10.6151
R1885 B.n486 B.n322 10.6151
R1886 B.n481 B.n322 10.6151
R1887 B.n481 B.n480 10.6151
R1888 B.n480 B.n479 10.6151
R1889 B.n479 B.n324 10.6151
R1890 B.n473 B.n324 10.6151
R1891 B.n473 B.n472 10.6151
R1892 B.n472 B.n471 10.6151
R1893 B.n467 B.n466 10.6151
R1894 B.n466 B.n330 10.6151
R1895 B.n461 B.n330 10.6151
R1896 B.n461 B.n460 10.6151
R1897 B.n460 B.n459 10.6151
R1898 B.n459 B.n332 10.6151
R1899 B.n453 B.n332 10.6151
R1900 B.n453 B.n452 10.6151
R1901 B.n452 B.n451 10.6151
R1902 B.n451 B.n334 10.6151
R1903 B.n445 B.n334 10.6151
R1904 B.n445 B.n444 10.6151
R1905 B.n444 B.n443 10.6151
R1906 B.n443 B.n336 10.6151
R1907 B.n437 B.n336 10.6151
R1908 B.n437 B.n436 10.6151
R1909 B.n436 B.n435 10.6151
R1910 B.n435 B.n338 10.6151
R1911 B.n429 B.n338 10.6151
R1912 B.n429 B.n428 10.6151
R1913 B.n428 B.n427 10.6151
R1914 B.n427 B.n340 10.6151
R1915 B.n421 B.n340 10.6151
R1916 B.n421 B.n420 10.6151
R1917 B.n420 B.n419 10.6151
R1918 B.n419 B.n342 10.6151
R1919 B.n413 B.n342 10.6151
R1920 B.n413 B.n412 10.6151
R1921 B.n412 B.n411 10.6151
R1922 B.n411 B.n344 10.6151
R1923 B.n405 B.n344 10.6151
R1924 B.n405 B.n404 10.6151
R1925 B.n404 B.n403 10.6151
R1926 B.n403 B.n346 10.6151
R1927 B.n397 B.n346 10.6151
R1928 B.n397 B.n396 10.6151
R1929 B.n396 B.n395 10.6151
R1930 B.n395 B.n348 10.6151
R1931 B.n389 B.n348 10.6151
R1932 B.n389 B.n388 10.6151
R1933 B.n388 B.n387 10.6151
R1934 B.n387 B.n350 10.6151
R1935 B.n381 B.n350 10.6151
R1936 B.n381 B.n380 10.6151
R1937 B.n380 B.n379 10.6151
R1938 B.n379 B.n352 10.6151
R1939 B.n373 B.n352 10.6151
R1940 B.n373 B.n372 10.6151
R1941 B.n372 B.n371 10.6151
R1942 B.n371 B.n354 10.6151
R1943 B.n365 B.n354 10.6151
R1944 B.n365 B.n364 10.6151
R1945 B.n364 B.n363 10.6151
R1946 B.n363 B.n356 10.6151
R1947 B.n357 B.n356 10.6151
R1948 B.n357 B.n286 10.6151
R1949 B.n602 B.n282 10.6151
R1950 B.n612 B.n282 10.6151
R1951 B.n613 B.n612 10.6151
R1952 B.n614 B.n613 10.6151
R1953 B.n614 B.n274 10.6151
R1954 B.n624 B.n274 10.6151
R1955 B.n625 B.n624 10.6151
R1956 B.n626 B.n625 10.6151
R1957 B.n626 B.n266 10.6151
R1958 B.n636 B.n266 10.6151
R1959 B.n637 B.n636 10.6151
R1960 B.n638 B.n637 10.6151
R1961 B.n638 B.n258 10.6151
R1962 B.n648 B.n258 10.6151
R1963 B.n649 B.n648 10.6151
R1964 B.n650 B.n649 10.6151
R1965 B.n650 B.n250 10.6151
R1966 B.n660 B.n250 10.6151
R1967 B.n661 B.n660 10.6151
R1968 B.n662 B.n661 10.6151
R1969 B.n662 B.n242 10.6151
R1970 B.n672 B.n242 10.6151
R1971 B.n673 B.n672 10.6151
R1972 B.n674 B.n673 10.6151
R1973 B.n674 B.n234 10.6151
R1974 B.n684 B.n234 10.6151
R1975 B.n685 B.n684 10.6151
R1976 B.n686 B.n685 10.6151
R1977 B.n686 B.n226 10.6151
R1978 B.n696 B.n226 10.6151
R1979 B.n697 B.n696 10.6151
R1980 B.n698 B.n697 10.6151
R1981 B.n698 B.n218 10.6151
R1982 B.n708 B.n218 10.6151
R1983 B.n709 B.n708 10.6151
R1984 B.n710 B.n709 10.6151
R1985 B.n710 B.n210 10.6151
R1986 B.n720 B.n210 10.6151
R1987 B.n721 B.n720 10.6151
R1988 B.n722 B.n721 10.6151
R1989 B.n722 B.n202 10.6151
R1990 B.n732 B.n202 10.6151
R1991 B.n733 B.n732 10.6151
R1992 B.n734 B.n733 10.6151
R1993 B.n734 B.n194 10.6151
R1994 B.n744 B.n194 10.6151
R1995 B.n745 B.n744 10.6151
R1996 B.n746 B.n745 10.6151
R1997 B.n746 B.n186 10.6151
R1998 B.n756 B.n186 10.6151
R1999 B.n757 B.n756 10.6151
R2000 B.n758 B.n757 10.6151
R2001 B.n758 B.n178 10.6151
R2002 B.n769 B.n178 10.6151
R2003 B.n770 B.n769 10.6151
R2004 B.n771 B.n770 10.6151
R2005 B.n771 B.n0 10.6151
R2006 B.n1211 B.n1 10.6151
R2007 B.n1211 B.n1210 10.6151
R2008 B.n1210 B.n1209 10.6151
R2009 B.n1209 B.n10 10.6151
R2010 B.n1203 B.n10 10.6151
R2011 B.n1203 B.n1202 10.6151
R2012 B.n1202 B.n1201 10.6151
R2013 B.n1201 B.n17 10.6151
R2014 B.n1195 B.n17 10.6151
R2015 B.n1195 B.n1194 10.6151
R2016 B.n1194 B.n1193 10.6151
R2017 B.n1193 B.n24 10.6151
R2018 B.n1187 B.n24 10.6151
R2019 B.n1187 B.n1186 10.6151
R2020 B.n1186 B.n1185 10.6151
R2021 B.n1185 B.n31 10.6151
R2022 B.n1179 B.n31 10.6151
R2023 B.n1179 B.n1178 10.6151
R2024 B.n1178 B.n1177 10.6151
R2025 B.n1177 B.n38 10.6151
R2026 B.n1171 B.n38 10.6151
R2027 B.n1171 B.n1170 10.6151
R2028 B.n1170 B.n1169 10.6151
R2029 B.n1169 B.n45 10.6151
R2030 B.n1163 B.n45 10.6151
R2031 B.n1163 B.n1162 10.6151
R2032 B.n1162 B.n1161 10.6151
R2033 B.n1161 B.n52 10.6151
R2034 B.n1155 B.n52 10.6151
R2035 B.n1155 B.n1154 10.6151
R2036 B.n1154 B.n1153 10.6151
R2037 B.n1153 B.n59 10.6151
R2038 B.n1147 B.n59 10.6151
R2039 B.n1147 B.n1146 10.6151
R2040 B.n1146 B.n1145 10.6151
R2041 B.n1145 B.n66 10.6151
R2042 B.n1139 B.n66 10.6151
R2043 B.n1139 B.n1138 10.6151
R2044 B.n1138 B.n1137 10.6151
R2045 B.n1137 B.n73 10.6151
R2046 B.n1131 B.n73 10.6151
R2047 B.n1131 B.n1130 10.6151
R2048 B.n1130 B.n1129 10.6151
R2049 B.n1129 B.n80 10.6151
R2050 B.n1123 B.n80 10.6151
R2051 B.n1123 B.n1122 10.6151
R2052 B.n1122 B.n1121 10.6151
R2053 B.n1121 B.n87 10.6151
R2054 B.n1115 B.n87 10.6151
R2055 B.n1115 B.n1114 10.6151
R2056 B.n1114 B.n1113 10.6151
R2057 B.n1113 B.n94 10.6151
R2058 B.n1107 B.n94 10.6151
R2059 B.n1107 B.n1106 10.6151
R2060 B.n1106 B.n1105 10.6151
R2061 B.n1105 B.n101 10.6151
R2062 B.n1099 B.n101 10.6151
R2063 B.n718 B.t5 10.215
R2064 B.n1175 B.t4 10.215
R2065 B.n986 B.n985 9.36635
R2066 B.n962 B.n146 9.36635
R2067 B.n491 B.n320 9.36635
R2068 B.n467 B.n328 9.36635
R2069 B.n240 B.t3 7.29654
R2070 B.t0 B.n1150 7.29654
R2071 B.n754 B.t2 5.35093
R2072 B.n1199 B.t1 5.35093
R2073 B.n1217 B.n0 2.81026
R2074 B.n1217 B.n1 2.81026
R2075 B.n985 B.n984 1.24928
R2076 B.n146 B.n142 1.24928
R2077 B.n487 B.n320 1.24928
R2078 B.n471 B.n328 1.24928
R2079 VN.n37 VN.n20 161.3
R2080 VN.n36 VN.n35 161.3
R2081 VN.n34 VN.n21 161.3
R2082 VN.n33 VN.n32 161.3
R2083 VN.n31 VN.n22 161.3
R2084 VN.n30 VN.n29 161.3
R2085 VN.n28 VN.n23 161.3
R2086 VN.n27 VN.n26 161.3
R2087 VN.n17 VN.n0 161.3
R2088 VN.n16 VN.n15 161.3
R2089 VN.n14 VN.n1 161.3
R2090 VN.n13 VN.n12 161.3
R2091 VN.n11 VN.n2 161.3
R2092 VN.n10 VN.n9 161.3
R2093 VN.n8 VN.n3 161.3
R2094 VN.n7 VN.n6 161.3
R2095 VN.n4 VN.t0 138.994
R2096 VN.n24 VN.t2 138.994
R2097 VN.n5 VN.t3 106.879
R2098 VN.n18 VN.t5 106.879
R2099 VN.n25 VN.t1 106.879
R2100 VN.n38 VN.t4 106.879
R2101 VN.n5 VN.n4 63.0818
R2102 VN.n25 VN.n24 63.0818
R2103 VN.n19 VN.n18 58.2799
R2104 VN.n39 VN.n38 58.2799
R2105 VN VN.n39 58.1786
R2106 VN.n12 VN.n11 53.171
R2107 VN.n32 VN.n31 53.171
R2108 VN.n12 VN.n1 27.983
R2109 VN.n32 VN.n21 27.983
R2110 VN.n6 VN.n3 24.5923
R2111 VN.n10 VN.n3 24.5923
R2112 VN.n11 VN.n10 24.5923
R2113 VN.n16 VN.n1 24.5923
R2114 VN.n17 VN.n16 24.5923
R2115 VN.n31 VN.n30 24.5923
R2116 VN.n30 VN.n23 24.5923
R2117 VN.n26 VN.n23 24.5923
R2118 VN.n37 VN.n36 24.5923
R2119 VN.n36 VN.n21 24.5923
R2120 VN.n18 VN.n17 24.1005
R2121 VN.n38 VN.n37 24.1005
R2122 VN.n6 VN.n5 12.2964
R2123 VN.n26 VN.n25 12.2964
R2124 VN.n27 VN.n24 2.54055
R2125 VN.n7 VN.n4 2.54055
R2126 VN.n39 VN.n20 0.417304
R2127 VN.n19 VN.n0 0.417304
R2128 VN VN.n19 0.394524
R2129 VN.n35 VN.n20 0.189894
R2130 VN.n35 VN.n34 0.189894
R2131 VN.n34 VN.n33 0.189894
R2132 VN.n33 VN.n22 0.189894
R2133 VN.n29 VN.n22 0.189894
R2134 VN.n29 VN.n28 0.189894
R2135 VN.n28 VN.n27 0.189894
R2136 VN.n8 VN.n7 0.189894
R2137 VN.n9 VN.n8 0.189894
R2138 VN.n9 VN.n2 0.189894
R2139 VN.n13 VN.n2 0.189894
R2140 VN.n14 VN.n13 0.189894
R2141 VN.n15 VN.n14 0.189894
R2142 VN.n15 VN.n0 0.189894
R2143 VTAIL.n7 VTAIL.t7 48.656
R2144 VTAIL.n11 VTAIL.t8 48.6559
R2145 VTAIL.n2 VTAIL.t1 48.6559
R2146 VTAIL.n10 VTAIL.t0 48.6559
R2147 VTAIL.n9 VTAIL.n8 47.5142
R2148 VTAIL.n6 VTAIL.n5 47.5142
R2149 VTAIL.n1 VTAIL.n0 47.5139
R2150 VTAIL.n4 VTAIL.n3 47.5139
R2151 VTAIL.n6 VTAIL.n4 34.6255
R2152 VTAIL.n11 VTAIL.n10 30.9703
R2153 VTAIL.n7 VTAIL.n6 3.65567
R2154 VTAIL.n10 VTAIL.n9 3.65567
R2155 VTAIL.n4 VTAIL.n2 3.65567
R2156 VTAIL VTAIL.n11 2.68369
R2157 VTAIL.n9 VTAIL.n7 2.29791
R2158 VTAIL.n2 VTAIL.n1 2.29791
R2159 VTAIL.n0 VTAIL.t11 1.14237
R2160 VTAIL.n0 VTAIL.t9 1.14237
R2161 VTAIL.n3 VTAIL.t2 1.14237
R2162 VTAIL.n3 VTAIL.t5 1.14237
R2163 VTAIL.n8 VTAIL.t4 1.14237
R2164 VTAIL.n8 VTAIL.t3 1.14237
R2165 VTAIL.n5 VTAIL.t6 1.14237
R2166 VTAIL.n5 VTAIL.t10 1.14237
R2167 VTAIL VTAIL.n1 0.972483
R2168 VDD2.n1 VDD2.t5 68.0207
R2169 VDD2.n2 VDD2.t1 65.3348
R2170 VDD2.n1 VDD2.n0 65.0512
R2171 VDD2 VDD2.n3 65.0484
R2172 VDD2.n2 VDD2.n1 50.5429
R2173 VDD2 VDD2.n2 2.80007
R2174 VDD2.n3 VDD2.t4 1.14237
R2175 VDD2.n3 VDD2.t3 1.14237
R2176 VDD2.n0 VDD2.t2 1.14237
R2177 VDD2.n0 VDD2.t0 1.14237
R2178 VP.n15 VP.n14 161.3
R2179 VP.n16 VP.n11 161.3
R2180 VP.n18 VP.n17 161.3
R2181 VP.n19 VP.n10 161.3
R2182 VP.n21 VP.n20 161.3
R2183 VP.n22 VP.n9 161.3
R2184 VP.n24 VP.n23 161.3
R2185 VP.n25 VP.n8 161.3
R2186 VP.n54 VP.n0 161.3
R2187 VP.n53 VP.n52 161.3
R2188 VP.n51 VP.n1 161.3
R2189 VP.n50 VP.n49 161.3
R2190 VP.n48 VP.n2 161.3
R2191 VP.n47 VP.n46 161.3
R2192 VP.n45 VP.n3 161.3
R2193 VP.n44 VP.n43 161.3
R2194 VP.n41 VP.n4 161.3
R2195 VP.n40 VP.n39 161.3
R2196 VP.n38 VP.n5 161.3
R2197 VP.n37 VP.n36 161.3
R2198 VP.n35 VP.n6 161.3
R2199 VP.n34 VP.n33 161.3
R2200 VP.n32 VP.n7 161.3
R2201 VP.n31 VP.n30 161.3
R2202 VP.n12 VP.t5 138.994
R2203 VP.n29 VP.t1 106.879
R2204 VP.n42 VP.t0 106.879
R2205 VP.n55 VP.t2 106.879
R2206 VP.n26 VP.t4 106.879
R2207 VP.n13 VP.t3 106.879
R2208 VP.n13 VP.n12 63.0818
R2209 VP.n29 VP.n28 58.2799
R2210 VP.n56 VP.n55 58.2799
R2211 VP.n27 VP.n26 58.2799
R2212 VP.n28 VP.n27 58.1408
R2213 VP.n36 VP.n35 53.171
R2214 VP.n49 VP.n48 53.171
R2215 VP.n20 VP.n19 53.171
R2216 VP.n35 VP.n34 27.983
R2217 VP.n49 VP.n1 27.983
R2218 VP.n20 VP.n9 27.983
R2219 VP.n30 VP.n7 24.5923
R2220 VP.n34 VP.n7 24.5923
R2221 VP.n36 VP.n5 24.5923
R2222 VP.n40 VP.n5 24.5923
R2223 VP.n41 VP.n40 24.5923
R2224 VP.n43 VP.n3 24.5923
R2225 VP.n47 VP.n3 24.5923
R2226 VP.n48 VP.n47 24.5923
R2227 VP.n53 VP.n1 24.5923
R2228 VP.n54 VP.n53 24.5923
R2229 VP.n24 VP.n9 24.5923
R2230 VP.n25 VP.n24 24.5923
R2231 VP.n14 VP.n11 24.5923
R2232 VP.n18 VP.n11 24.5923
R2233 VP.n19 VP.n18 24.5923
R2234 VP.n30 VP.n29 24.1005
R2235 VP.n55 VP.n54 24.1005
R2236 VP.n26 VP.n25 24.1005
R2237 VP.n42 VP.n41 12.2964
R2238 VP.n43 VP.n42 12.2964
R2239 VP.n14 VP.n13 12.2964
R2240 VP.n15 VP.n12 2.54052
R2241 VP.n27 VP.n8 0.417304
R2242 VP.n31 VP.n28 0.417304
R2243 VP.n56 VP.n0 0.417304
R2244 VP VP.n56 0.394524
R2245 VP.n16 VP.n15 0.189894
R2246 VP.n17 VP.n16 0.189894
R2247 VP.n17 VP.n10 0.189894
R2248 VP.n21 VP.n10 0.189894
R2249 VP.n22 VP.n21 0.189894
R2250 VP.n23 VP.n22 0.189894
R2251 VP.n23 VP.n8 0.189894
R2252 VP.n32 VP.n31 0.189894
R2253 VP.n33 VP.n32 0.189894
R2254 VP.n33 VP.n6 0.189894
R2255 VP.n37 VP.n6 0.189894
R2256 VP.n38 VP.n37 0.189894
R2257 VP.n39 VP.n38 0.189894
R2258 VP.n39 VP.n4 0.189894
R2259 VP.n44 VP.n4 0.189894
R2260 VP.n45 VP.n44 0.189894
R2261 VP.n46 VP.n45 0.189894
R2262 VP.n46 VP.n2 0.189894
R2263 VP.n50 VP.n2 0.189894
R2264 VP.n51 VP.n50 0.189894
R2265 VP.n52 VP.n51 0.189894
R2266 VP.n52 VP.n0 0.189894
R2267 VDD1 VDD1.t0 68.1344
R2268 VDD1.n1 VDD1.t4 68.0207
R2269 VDD1.n1 VDD1.n0 65.0512
R2270 VDD1.n3 VDD1.n2 64.1928
R2271 VDD1.n3 VDD1.n1 52.9535
R2272 VDD1.n2 VDD1.t2 1.14237
R2273 VDD1.n2 VDD1.t1 1.14237
R2274 VDD1.n0 VDD1.t5 1.14237
R2275 VDD1.n0 VDD1.t3 1.14237
R2276 VDD1 VDD1.n3 0.856103
C0 VDD2 VN 10.1866f
C1 VDD1 VN 0.152893f
C2 VN VP 9.183741f
C3 VDD2 VTAIL 9.96174f
C4 VDD1 VTAIL 9.9019f
C5 VTAIL VP 10.4192f
C6 VTAIL VN 10.403901f
C7 VDD1 VDD2 1.91886f
C8 VDD2 VP 0.569119f
C9 VDD1 VP 10.6001f
C10 VDD2 B 7.932517f
C11 VDD1 B 8.317008f
C12 VTAIL B 10.828926f
C13 VN B 17.168642f
C14 VP B 15.847204f
C15 VDD1.t0 B 3.43453f
C16 VDD1.t4 B 3.43352f
C17 VDD1.t5 B 0.293406f
C18 VDD1.t3 B 0.293406f
C19 VDD1.n0 B 2.67868f
C20 VDD1.n1 B 3.39464f
C21 VDD1.t2 B 0.293406f
C22 VDD1.t1 B 0.293406f
C23 VDD1.n2 B 2.67215f
C24 VDD1.n3 B 3.04692f
C25 VP.n0 B 0.032139f
C26 VP.t2 B 3.18499f
C27 VP.n1 B 0.033324f
C28 VP.n2 B 0.017091f
C29 VP.n3 B 0.031694f
C30 VP.n4 B 0.017091f
C31 VP.t0 B 3.18499f
C32 VP.n5 B 0.031694f
C33 VP.n6 B 0.017091f
C34 VP.n7 B 0.031694f
C35 VP.n8 B 0.032139f
C36 VP.t4 B 3.18499f
C37 VP.n9 B 0.033324f
C38 VP.n10 B 0.017091f
C39 VP.n11 B 0.031694f
C40 VP.t5 B 3.47024f
C41 VP.n12 B 1.10955f
C42 VP.t3 B 3.18499f
C43 VP.n13 B 1.15974f
C44 VP.n14 B 0.023871f
C45 VP.n15 B 0.223372f
C46 VP.n16 B 0.017091f
C47 VP.n17 B 0.017091f
C48 VP.n18 B 0.031694f
C49 VP.n19 B 0.03018f
C50 VP.n20 B 0.017879f
C51 VP.n21 B 0.017091f
C52 VP.n22 B 0.017091f
C53 VP.n23 B 0.017091f
C54 VP.n24 B 0.031694f
C55 VP.n25 B 0.031381f
C56 VP.n26 B 1.17638f
C57 VP.n27 B 1.21904f
C58 VP.n28 B 1.22963f
C59 VP.t1 B 3.18499f
C60 VP.n29 B 1.17638f
C61 VP.n30 B 0.031381f
C62 VP.n31 B 0.032139f
C63 VP.n32 B 0.017091f
C64 VP.n33 B 0.017091f
C65 VP.n34 B 0.033324f
C66 VP.n35 B 0.017879f
C67 VP.n36 B 0.03018f
C68 VP.n37 B 0.017091f
C69 VP.n38 B 0.017091f
C70 VP.n39 B 0.017091f
C71 VP.n40 B 0.031694f
C72 VP.n41 B 0.023871f
C73 VP.n42 B 1.09812f
C74 VP.n43 B 0.023871f
C75 VP.n44 B 0.017091f
C76 VP.n45 B 0.017091f
C77 VP.n46 B 0.017091f
C78 VP.n47 B 0.031694f
C79 VP.n48 B 0.03018f
C80 VP.n49 B 0.017879f
C81 VP.n50 B 0.017091f
C82 VP.n51 B 0.017091f
C83 VP.n52 B 0.017091f
C84 VP.n53 B 0.031694f
C85 VP.n54 B 0.031381f
C86 VP.n55 B 1.17638f
C87 VP.n56 B 0.050205f
C88 VDD2.t5 B 3.39638f
C89 VDD2.t2 B 0.290232f
C90 VDD2.t0 B 0.290232f
C91 VDD2.n0 B 2.64971f
C92 VDD2.n1 B 3.21921f
C93 VDD2.t1 B 3.37984f
C94 VDD2.n2 B 3.01258f
C95 VDD2.t4 B 0.290232f
C96 VDD2.t3 B 0.290232f
C97 VDD2.n3 B 2.64967f
C98 VTAIL.t11 B 0.318111f
C99 VTAIL.t9 B 0.318111f
C100 VTAIL.n0 B 2.83243f
C101 VTAIL.n1 B 0.466528f
C102 VTAIL.t1 B 3.62063f
C103 VTAIL.n2 B 0.746621f
C104 VTAIL.t2 B 0.318111f
C105 VTAIL.t5 B 0.318111f
C106 VTAIL.n3 B 2.83243f
C107 VTAIL.n4 B 2.4758f
C108 VTAIL.t6 B 0.318111f
C109 VTAIL.t10 B 0.318111f
C110 VTAIL.n5 B 2.83244f
C111 VTAIL.n6 B 2.4758f
C112 VTAIL.t7 B 3.62066f
C113 VTAIL.n7 B 0.7466f
C114 VTAIL.t4 B 0.318111f
C115 VTAIL.t3 B 0.318111f
C116 VTAIL.n8 B 2.83244f
C117 VTAIL.n9 B 0.667241f
C118 VTAIL.t0 B 3.62063f
C119 VTAIL.n10 B 2.28175f
C120 VTAIL.t8 B 3.62063f
C121 VTAIL.n11 B 2.20904f
C122 VN.n0 B 0.031688f
C123 VN.t5 B 3.14031f
C124 VN.n1 B 0.032857f
C125 VN.n2 B 0.016851f
C126 VN.n3 B 0.031249f
C127 VN.t0 B 3.42155f
C128 VN.n4 B 1.09398f
C129 VN.t3 B 3.14031f
C130 VN.n5 B 1.14347f
C131 VN.n6 B 0.023536f
C132 VN.n7 B 0.220238f
C133 VN.n8 B 0.016851f
C134 VN.n9 B 0.016851f
C135 VN.n10 B 0.031249f
C136 VN.n11 B 0.029757f
C137 VN.n12 B 0.017628f
C138 VN.n13 B 0.016851f
C139 VN.n14 B 0.016851f
C140 VN.n15 B 0.016851f
C141 VN.n16 B 0.031249f
C142 VN.n17 B 0.030941f
C143 VN.n18 B 1.15988f
C144 VN.n19 B 0.049501f
C145 VN.n20 B 0.031688f
C146 VN.t4 B 3.14031f
C147 VN.n21 B 0.032857f
C148 VN.n22 B 0.016851f
C149 VN.n23 B 0.031249f
C150 VN.t2 B 3.42155f
C151 VN.n24 B 1.09398f
C152 VN.t1 B 3.14031f
C153 VN.n25 B 1.14347f
C154 VN.n26 B 0.023536f
C155 VN.n27 B 0.220238f
C156 VN.n28 B 0.016851f
C157 VN.n29 B 0.016851f
C158 VN.n30 B 0.031249f
C159 VN.n31 B 0.029757f
C160 VN.n32 B 0.017628f
C161 VN.n33 B 0.016851f
C162 VN.n34 B 0.016851f
C163 VN.n35 B 0.016851f
C164 VN.n36 B 0.031249f
C165 VN.n37 B 0.030941f
C166 VN.n38 B 1.15988f
C167 VN.n39 B 1.20586f
.ends

