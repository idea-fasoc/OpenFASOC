* NGSPICE file created from diff_pair_sample_1141.ext - technology: sky130A

.subckt diff_pair_sample_1141 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9932 pd=12.41 as=1.9932 ps=12.41 w=12.08 l=1.46
X1 VTAIL.t10 VN.t1 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9932 pd=12.41 as=1.9932 ps=12.41 w=12.08 l=1.46
X2 VDD1.t5 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7112 pd=24.94 as=1.9932 ps=12.41 w=12.08 l=1.46
X3 VDD2.t2 VN.t2 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7112 pd=24.94 as=1.9932 ps=12.41 w=12.08 l=1.46
X4 VDD2.t0 VN.t3 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=4.7112 pd=24.94 as=1.9932 ps=12.41 w=12.08 l=1.46
X5 VTAIL.t0 VP.t1 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.9932 pd=12.41 as=1.9932 ps=12.41 w=12.08 l=1.46
X6 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7112 pd=24.94 as=0 ps=0 w=12.08 l=1.46
X7 VDD2.t3 VN.t4 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9932 pd=12.41 as=4.7112 ps=24.94 w=12.08 l=1.46
X8 VDD2.t5 VN.t5 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9932 pd=12.41 as=4.7112 ps=24.94 w=12.08 l=1.46
X9 VDD1.t3 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.9932 pd=12.41 as=4.7112 ps=24.94 w=12.08 l=1.46
X10 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7112 pd=24.94 as=0 ps=0 w=12.08 l=1.46
X11 VTAIL.t2 VP.t3 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.9932 pd=12.41 as=1.9932 ps=12.41 w=12.08 l=1.46
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7112 pd=24.94 as=0 ps=0 w=12.08 l=1.46
X13 VDD1.t1 VP.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.9932 pd=12.41 as=4.7112 ps=24.94 w=12.08 l=1.46
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7112 pd=24.94 as=0 ps=0 w=12.08 l=1.46
X15 VDD1.t0 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.7112 pd=24.94 as=1.9932 ps=12.41 w=12.08 l=1.46
R0 VN.n3 VN.t2 236.121
R1 VN.n13 VN.t5 236.121
R2 VN.n2 VN.t1 199.404
R3 VN.n8 VN.t4 199.404
R4 VN.n12 VN.t0 199.404
R5 VN.n18 VN.t3 199.404
R6 VN.n9 VN.n8 171.63
R7 VN.n19 VN.n18 171.63
R8 VN.n17 VN.n10 161.3
R9 VN.n16 VN.n15 161.3
R10 VN.n14 VN.n11 161.3
R11 VN.n7 VN.n0 161.3
R12 VN.n6 VN.n5 161.3
R13 VN.n4 VN.n1 161.3
R14 VN.n6 VN.n1 50.7491
R15 VN.n16 VN.n11 50.7491
R16 VN VN.n19 44.6274
R17 VN.n3 VN.n2 41.9508
R18 VN.n13 VN.n12 41.9508
R19 VN.n7 VN.n6 30.405
R20 VN.n17 VN.n16 30.405
R21 VN.n2 VN.n1 24.5923
R22 VN.n12 VN.n11 24.5923
R23 VN.n14 VN.n13 17.3014
R24 VN.n4 VN.n3 17.3014
R25 VN.n8 VN.n7 14.2638
R26 VN.n18 VN.n17 14.2638
R27 VN.n19 VN.n10 0.189894
R28 VN.n15 VN.n10 0.189894
R29 VN.n15 VN.n14 0.189894
R30 VN.n5 VN.n4 0.189894
R31 VN.n5 VN.n0 0.189894
R32 VN.n9 VN.n0 0.189894
R33 VN VN.n9 0.0516364
R34 VDD2.n127 VDD2.n67 289.615
R35 VDD2.n60 VDD2.n0 289.615
R36 VDD2.n128 VDD2.n127 185
R37 VDD2.n126 VDD2.n125 185
R38 VDD2.n71 VDD2.n70 185
R39 VDD2.n120 VDD2.n119 185
R40 VDD2.n118 VDD2.n117 185
R41 VDD2.n75 VDD2.n74 185
R42 VDD2.n112 VDD2.n111 185
R43 VDD2.n110 VDD2.n77 185
R44 VDD2.n109 VDD2.n108 185
R45 VDD2.n80 VDD2.n78 185
R46 VDD2.n103 VDD2.n102 185
R47 VDD2.n101 VDD2.n100 185
R48 VDD2.n84 VDD2.n83 185
R49 VDD2.n95 VDD2.n94 185
R50 VDD2.n93 VDD2.n92 185
R51 VDD2.n88 VDD2.n87 185
R52 VDD2.n20 VDD2.n19 185
R53 VDD2.n25 VDD2.n24 185
R54 VDD2.n27 VDD2.n26 185
R55 VDD2.n16 VDD2.n15 185
R56 VDD2.n33 VDD2.n32 185
R57 VDD2.n35 VDD2.n34 185
R58 VDD2.n12 VDD2.n11 185
R59 VDD2.n42 VDD2.n41 185
R60 VDD2.n43 VDD2.n10 185
R61 VDD2.n45 VDD2.n44 185
R62 VDD2.n8 VDD2.n7 185
R63 VDD2.n51 VDD2.n50 185
R64 VDD2.n53 VDD2.n52 185
R65 VDD2.n4 VDD2.n3 185
R66 VDD2.n59 VDD2.n58 185
R67 VDD2.n61 VDD2.n60 185
R68 VDD2.n89 VDD2.t0 149.524
R69 VDD2.n21 VDD2.t2 149.524
R70 VDD2.n127 VDD2.n126 104.615
R71 VDD2.n126 VDD2.n70 104.615
R72 VDD2.n119 VDD2.n70 104.615
R73 VDD2.n119 VDD2.n118 104.615
R74 VDD2.n118 VDD2.n74 104.615
R75 VDD2.n111 VDD2.n74 104.615
R76 VDD2.n111 VDD2.n110 104.615
R77 VDD2.n110 VDD2.n109 104.615
R78 VDD2.n109 VDD2.n78 104.615
R79 VDD2.n102 VDD2.n78 104.615
R80 VDD2.n102 VDD2.n101 104.615
R81 VDD2.n101 VDD2.n83 104.615
R82 VDD2.n94 VDD2.n83 104.615
R83 VDD2.n94 VDD2.n93 104.615
R84 VDD2.n93 VDD2.n87 104.615
R85 VDD2.n25 VDD2.n19 104.615
R86 VDD2.n26 VDD2.n25 104.615
R87 VDD2.n26 VDD2.n15 104.615
R88 VDD2.n33 VDD2.n15 104.615
R89 VDD2.n34 VDD2.n33 104.615
R90 VDD2.n34 VDD2.n11 104.615
R91 VDD2.n42 VDD2.n11 104.615
R92 VDD2.n43 VDD2.n42 104.615
R93 VDD2.n44 VDD2.n43 104.615
R94 VDD2.n44 VDD2.n7 104.615
R95 VDD2.n51 VDD2.n7 104.615
R96 VDD2.n52 VDD2.n51 104.615
R97 VDD2.n52 VDD2.n3 104.615
R98 VDD2.n59 VDD2.n3 104.615
R99 VDD2.n60 VDD2.n59 104.615
R100 VDD2.n66 VDD2.n65 61.4344
R101 VDD2 VDD2.n133 61.4316
R102 VDD2.t0 VDD2.n87 52.3082
R103 VDD2.t2 VDD2.n19 52.3082
R104 VDD2.n66 VDD2.n64 49.1904
R105 VDD2.n132 VDD2.n131 48.0884
R106 VDD2.n132 VDD2.n66 39.1442
R107 VDD2.n112 VDD2.n77 13.1884
R108 VDD2.n45 VDD2.n10 13.1884
R109 VDD2.n113 VDD2.n75 12.8005
R110 VDD2.n108 VDD2.n79 12.8005
R111 VDD2.n41 VDD2.n40 12.8005
R112 VDD2.n46 VDD2.n8 12.8005
R113 VDD2.n117 VDD2.n116 12.0247
R114 VDD2.n107 VDD2.n80 12.0247
R115 VDD2.n39 VDD2.n12 12.0247
R116 VDD2.n50 VDD2.n49 12.0247
R117 VDD2.n120 VDD2.n73 11.249
R118 VDD2.n104 VDD2.n103 11.249
R119 VDD2.n36 VDD2.n35 11.249
R120 VDD2.n53 VDD2.n6 11.249
R121 VDD2.n121 VDD2.n71 10.4732
R122 VDD2.n100 VDD2.n82 10.4732
R123 VDD2.n32 VDD2.n14 10.4732
R124 VDD2.n54 VDD2.n4 10.4732
R125 VDD2.n89 VDD2.n88 10.2747
R126 VDD2.n21 VDD2.n20 10.2747
R127 VDD2.n125 VDD2.n124 9.69747
R128 VDD2.n99 VDD2.n84 9.69747
R129 VDD2.n31 VDD2.n16 9.69747
R130 VDD2.n58 VDD2.n57 9.69747
R131 VDD2.n131 VDD2.n130 9.45567
R132 VDD2.n64 VDD2.n63 9.45567
R133 VDD2.n91 VDD2.n90 9.3005
R134 VDD2.n86 VDD2.n85 9.3005
R135 VDD2.n97 VDD2.n96 9.3005
R136 VDD2.n99 VDD2.n98 9.3005
R137 VDD2.n82 VDD2.n81 9.3005
R138 VDD2.n105 VDD2.n104 9.3005
R139 VDD2.n107 VDD2.n106 9.3005
R140 VDD2.n79 VDD2.n76 9.3005
R141 VDD2.n130 VDD2.n129 9.3005
R142 VDD2.n69 VDD2.n68 9.3005
R143 VDD2.n124 VDD2.n123 9.3005
R144 VDD2.n122 VDD2.n121 9.3005
R145 VDD2.n73 VDD2.n72 9.3005
R146 VDD2.n116 VDD2.n115 9.3005
R147 VDD2.n114 VDD2.n113 9.3005
R148 VDD2.n63 VDD2.n62 9.3005
R149 VDD2.n2 VDD2.n1 9.3005
R150 VDD2.n57 VDD2.n56 9.3005
R151 VDD2.n55 VDD2.n54 9.3005
R152 VDD2.n6 VDD2.n5 9.3005
R153 VDD2.n49 VDD2.n48 9.3005
R154 VDD2.n47 VDD2.n46 9.3005
R155 VDD2.n23 VDD2.n22 9.3005
R156 VDD2.n18 VDD2.n17 9.3005
R157 VDD2.n29 VDD2.n28 9.3005
R158 VDD2.n31 VDD2.n30 9.3005
R159 VDD2.n14 VDD2.n13 9.3005
R160 VDD2.n37 VDD2.n36 9.3005
R161 VDD2.n39 VDD2.n38 9.3005
R162 VDD2.n40 VDD2.n9 9.3005
R163 VDD2.n128 VDD2.n69 8.92171
R164 VDD2.n96 VDD2.n95 8.92171
R165 VDD2.n28 VDD2.n27 8.92171
R166 VDD2.n61 VDD2.n2 8.92171
R167 VDD2.n129 VDD2.n67 8.14595
R168 VDD2.n92 VDD2.n86 8.14595
R169 VDD2.n24 VDD2.n18 8.14595
R170 VDD2.n62 VDD2.n0 8.14595
R171 VDD2.n91 VDD2.n88 7.3702
R172 VDD2.n23 VDD2.n20 7.3702
R173 VDD2.n131 VDD2.n67 5.81868
R174 VDD2.n92 VDD2.n91 5.81868
R175 VDD2.n24 VDD2.n23 5.81868
R176 VDD2.n64 VDD2.n0 5.81868
R177 VDD2.n129 VDD2.n128 5.04292
R178 VDD2.n95 VDD2.n86 5.04292
R179 VDD2.n27 VDD2.n18 5.04292
R180 VDD2.n62 VDD2.n61 5.04292
R181 VDD2.n125 VDD2.n69 4.26717
R182 VDD2.n96 VDD2.n84 4.26717
R183 VDD2.n28 VDD2.n16 4.26717
R184 VDD2.n58 VDD2.n2 4.26717
R185 VDD2.n124 VDD2.n71 3.49141
R186 VDD2.n100 VDD2.n99 3.49141
R187 VDD2.n32 VDD2.n31 3.49141
R188 VDD2.n57 VDD2.n4 3.49141
R189 VDD2.n90 VDD2.n89 2.84303
R190 VDD2.n22 VDD2.n21 2.84303
R191 VDD2.n121 VDD2.n120 2.71565
R192 VDD2.n103 VDD2.n82 2.71565
R193 VDD2.n35 VDD2.n14 2.71565
R194 VDD2.n54 VDD2.n53 2.71565
R195 VDD2.n117 VDD2.n73 1.93989
R196 VDD2.n104 VDD2.n80 1.93989
R197 VDD2.n36 VDD2.n12 1.93989
R198 VDD2.n50 VDD2.n6 1.93989
R199 VDD2.n133 VDD2.t4 1.63957
R200 VDD2.n133 VDD2.t5 1.63957
R201 VDD2.n65 VDD2.t1 1.63957
R202 VDD2.n65 VDD2.t3 1.63957
R203 VDD2 VDD2.n132 1.21602
R204 VDD2.n116 VDD2.n75 1.16414
R205 VDD2.n108 VDD2.n107 1.16414
R206 VDD2.n41 VDD2.n39 1.16414
R207 VDD2.n49 VDD2.n8 1.16414
R208 VDD2.n113 VDD2.n112 0.388379
R209 VDD2.n79 VDD2.n77 0.388379
R210 VDD2.n40 VDD2.n10 0.388379
R211 VDD2.n46 VDD2.n45 0.388379
R212 VDD2.n130 VDD2.n68 0.155672
R213 VDD2.n123 VDD2.n68 0.155672
R214 VDD2.n123 VDD2.n122 0.155672
R215 VDD2.n122 VDD2.n72 0.155672
R216 VDD2.n115 VDD2.n72 0.155672
R217 VDD2.n115 VDD2.n114 0.155672
R218 VDD2.n114 VDD2.n76 0.155672
R219 VDD2.n106 VDD2.n76 0.155672
R220 VDD2.n106 VDD2.n105 0.155672
R221 VDD2.n105 VDD2.n81 0.155672
R222 VDD2.n98 VDD2.n81 0.155672
R223 VDD2.n98 VDD2.n97 0.155672
R224 VDD2.n97 VDD2.n85 0.155672
R225 VDD2.n90 VDD2.n85 0.155672
R226 VDD2.n22 VDD2.n17 0.155672
R227 VDD2.n29 VDD2.n17 0.155672
R228 VDD2.n30 VDD2.n29 0.155672
R229 VDD2.n30 VDD2.n13 0.155672
R230 VDD2.n37 VDD2.n13 0.155672
R231 VDD2.n38 VDD2.n37 0.155672
R232 VDD2.n38 VDD2.n9 0.155672
R233 VDD2.n47 VDD2.n9 0.155672
R234 VDD2.n48 VDD2.n47 0.155672
R235 VDD2.n48 VDD2.n5 0.155672
R236 VDD2.n55 VDD2.n5 0.155672
R237 VDD2.n56 VDD2.n55 0.155672
R238 VDD2.n56 VDD2.n1 0.155672
R239 VDD2.n63 VDD2.n1 0.155672
R240 VTAIL.n266 VTAIL.n206 289.615
R241 VTAIL.n62 VTAIL.n2 289.615
R242 VTAIL.n200 VTAIL.n140 289.615
R243 VTAIL.n132 VTAIL.n72 289.615
R244 VTAIL.n226 VTAIL.n225 185
R245 VTAIL.n231 VTAIL.n230 185
R246 VTAIL.n233 VTAIL.n232 185
R247 VTAIL.n222 VTAIL.n221 185
R248 VTAIL.n239 VTAIL.n238 185
R249 VTAIL.n241 VTAIL.n240 185
R250 VTAIL.n218 VTAIL.n217 185
R251 VTAIL.n248 VTAIL.n247 185
R252 VTAIL.n249 VTAIL.n216 185
R253 VTAIL.n251 VTAIL.n250 185
R254 VTAIL.n214 VTAIL.n213 185
R255 VTAIL.n257 VTAIL.n256 185
R256 VTAIL.n259 VTAIL.n258 185
R257 VTAIL.n210 VTAIL.n209 185
R258 VTAIL.n265 VTAIL.n264 185
R259 VTAIL.n267 VTAIL.n266 185
R260 VTAIL.n22 VTAIL.n21 185
R261 VTAIL.n27 VTAIL.n26 185
R262 VTAIL.n29 VTAIL.n28 185
R263 VTAIL.n18 VTAIL.n17 185
R264 VTAIL.n35 VTAIL.n34 185
R265 VTAIL.n37 VTAIL.n36 185
R266 VTAIL.n14 VTAIL.n13 185
R267 VTAIL.n44 VTAIL.n43 185
R268 VTAIL.n45 VTAIL.n12 185
R269 VTAIL.n47 VTAIL.n46 185
R270 VTAIL.n10 VTAIL.n9 185
R271 VTAIL.n53 VTAIL.n52 185
R272 VTAIL.n55 VTAIL.n54 185
R273 VTAIL.n6 VTAIL.n5 185
R274 VTAIL.n61 VTAIL.n60 185
R275 VTAIL.n63 VTAIL.n62 185
R276 VTAIL.n201 VTAIL.n200 185
R277 VTAIL.n199 VTAIL.n198 185
R278 VTAIL.n144 VTAIL.n143 185
R279 VTAIL.n193 VTAIL.n192 185
R280 VTAIL.n191 VTAIL.n190 185
R281 VTAIL.n148 VTAIL.n147 185
R282 VTAIL.n185 VTAIL.n184 185
R283 VTAIL.n183 VTAIL.n150 185
R284 VTAIL.n182 VTAIL.n181 185
R285 VTAIL.n153 VTAIL.n151 185
R286 VTAIL.n176 VTAIL.n175 185
R287 VTAIL.n174 VTAIL.n173 185
R288 VTAIL.n157 VTAIL.n156 185
R289 VTAIL.n168 VTAIL.n167 185
R290 VTAIL.n166 VTAIL.n165 185
R291 VTAIL.n161 VTAIL.n160 185
R292 VTAIL.n133 VTAIL.n132 185
R293 VTAIL.n131 VTAIL.n130 185
R294 VTAIL.n76 VTAIL.n75 185
R295 VTAIL.n125 VTAIL.n124 185
R296 VTAIL.n123 VTAIL.n122 185
R297 VTAIL.n80 VTAIL.n79 185
R298 VTAIL.n117 VTAIL.n116 185
R299 VTAIL.n115 VTAIL.n82 185
R300 VTAIL.n114 VTAIL.n113 185
R301 VTAIL.n85 VTAIL.n83 185
R302 VTAIL.n108 VTAIL.n107 185
R303 VTAIL.n106 VTAIL.n105 185
R304 VTAIL.n89 VTAIL.n88 185
R305 VTAIL.n100 VTAIL.n99 185
R306 VTAIL.n98 VTAIL.n97 185
R307 VTAIL.n93 VTAIL.n92 185
R308 VTAIL.n227 VTAIL.t7 149.524
R309 VTAIL.n23 VTAIL.t3 149.524
R310 VTAIL.n162 VTAIL.t4 149.524
R311 VTAIL.n94 VTAIL.t6 149.524
R312 VTAIL.n231 VTAIL.n225 104.615
R313 VTAIL.n232 VTAIL.n231 104.615
R314 VTAIL.n232 VTAIL.n221 104.615
R315 VTAIL.n239 VTAIL.n221 104.615
R316 VTAIL.n240 VTAIL.n239 104.615
R317 VTAIL.n240 VTAIL.n217 104.615
R318 VTAIL.n248 VTAIL.n217 104.615
R319 VTAIL.n249 VTAIL.n248 104.615
R320 VTAIL.n250 VTAIL.n249 104.615
R321 VTAIL.n250 VTAIL.n213 104.615
R322 VTAIL.n257 VTAIL.n213 104.615
R323 VTAIL.n258 VTAIL.n257 104.615
R324 VTAIL.n258 VTAIL.n209 104.615
R325 VTAIL.n265 VTAIL.n209 104.615
R326 VTAIL.n266 VTAIL.n265 104.615
R327 VTAIL.n27 VTAIL.n21 104.615
R328 VTAIL.n28 VTAIL.n27 104.615
R329 VTAIL.n28 VTAIL.n17 104.615
R330 VTAIL.n35 VTAIL.n17 104.615
R331 VTAIL.n36 VTAIL.n35 104.615
R332 VTAIL.n36 VTAIL.n13 104.615
R333 VTAIL.n44 VTAIL.n13 104.615
R334 VTAIL.n45 VTAIL.n44 104.615
R335 VTAIL.n46 VTAIL.n45 104.615
R336 VTAIL.n46 VTAIL.n9 104.615
R337 VTAIL.n53 VTAIL.n9 104.615
R338 VTAIL.n54 VTAIL.n53 104.615
R339 VTAIL.n54 VTAIL.n5 104.615
R340 VTAIL.n61 VTAIL.n5 104.615
R341 VTAIL.n62 VTAIL.n61 104.615
R342 VTAIL.n200 VTAIL.n199 104.615
R343 VTAIL.n199 VTAIL.n143 104.615
R344 VTAIL.n192 VTAIL.n143 104.615
R345 VTAIL.n192 VTAIL.n191 104.615
R346 VTAIL.n191 VTAIL.n147 104.615
R347 VTAIL.n184 VTAIL.n147 104.615
R348 VTAIL.n184 VTAIL.n183 104.615
R349 VTAIL.n183 VTAIL.n182 104.615
R350 VTAIL.n182 VTAIL.n151 104.615
R351 VTAIL.n175 VTAIL.n151 104.615
R352 VTAIL.n175 VTAIL.n174 104.615
R353 VTAIL.n174 VTAIL.n156 104.615
R354 VTAIL.n167 VTAIL.n156 104.615
R355 VTAIL.n167 VTAIL.n166 104.615
R356 VTAIL.n166 VTAIL.n160 104.615
R357 VTAIL.n132 VTAIL.n131 104.615
R358 VTAIL.n131 VTAIL.n75 104.615
R359 VTAIL.n124 VTAIL.n75 104.615
R360 VTAIL.n124 VTAIL.n123 104.615
R361 VTAIL.n123 VTAIL.n79 104.615
R362 VTAIL.n116 VTAIL.n79 104.615
R363 VTAIL.n116 VTAIL.n115 104.615
R364 VTAIL.n115 VTAIL.n114 104.615
R365 VTAIL.n114 VTAIL.n83 104.615
R366 VTAIL.n107 VTAIL.n83 104.615
R367 VTAIL.n107 VTAIL.n106 104.615
R368 VTAIL.n106 VTAIL.n88 104.615
R369 VTAIL.n99 VTAIL.n88 104.615
R370 VTAIL.n99 VTAIL.n98 104.615
R371 VTAIL.n98 VTAIL.n92 104.615
R372 VTAIL.t7 VTAIL.n225 52.3082
R373 VTAIL.t3 VTAIL.n21 52.3082
R374 VTAIL.t4 VTAIL.n160 52.3082
R375 VTAIL.t6 VTAIL.n92 52.3082
R376 VTAIL.n139 VTAIL.n138 44.4254
R377 VTAIL.n71 VTAIL.n70 44.4254
R378 VTAIL.n1 VTAIL.n0 44.4252
R379 VTAIL.n69 VTAIL.n68 44.4252
R380 VTAIL.n271 VTAIL.n270 31.4096
R381 VTAIL.n67 VTAIL.n66 31.4096
R382 VTAIL.n205 VTAIL.n204 31.4096
R383 VTAIL.n137 VTAIL.n136 31.4096
R384 VTAIL.n71 VTAIL.n69 25.8669
R385 VTAIL.n271 VTAIL.n205 24.3238
R386 VTAIL.n251 VTAIL.n216 13.1884
R387 VTAIL.n47 VTAIL.n12 13.1884
R388 VTAIL.n185 VTAIL.n150 13.1884
R389 VTAIL.n117 VTAIL.n82 13.1884
R390 VTAIL.n247 VTAIL.n246 12.8005
R391 VTAIL.n252 VTAIL.n214 12.8005
R392 VTAIL.n43 VTAIL.n42 12.8005
R393 VTAIL.n48 VTAIL.n10 12.8005
R394 VTAIL.n186 VTAIL.n148 12.8005
R395 VTAIL.n181 VTAIL.n152 12.8005
R396 VTAIL.n118 VTAIL.n80 12.8005
R397 VTAIL.n113 VTAIL.n84 12.8005
R398 VTAIL.n245 VTAIL.n218 12.0247
R399 VTAIL.n256 VTAIL.n255 12.0247
R400 VTAIL.n41 VTAIL.n14 12.0247
R401 VTAIL.n52 VTAIL.n51 12.0247
R402 VTAIL.n190 VTAIL.n189 12.0247
R403 VTAIL.n180 VTAIL.n153 12.0247
R404 VTAIL.n122 VTAIL.n121 12.0247
R405 VTAIL.n112 VTAIL.n85 12.0247
R406 VTAIL.n242 VTAIL.n241 11.249
R407 VTAIL.n259 VTAIL.n212 11.249
R408 VTAIL.n38 VTAIL.n37 11.249
R409 VTAIL.n55 VTAIL.n8 11.249
R410 VTAIL.n193 VTAIL.n146 11.249
R411 VTAIL.n177 VTAIL.n176 11.249
R412 VTAIL.n125 VTAIL.n78 11.249
R413 VTAIL.n109 VTAIL.n108 11.249
R414 VTAIL.n238 VTAIL.n220 10.4732
R415 VTAIL.n260 VTAIL.n210 10.4732
R416 VTAIL.n34 VTAIL.n16 10.4732
R417 VTAIL.n56 VTAIL.n6 10.4732
R418 VTAIL.n194 VTAIL.n144 10.4732
R419 VTAIL.n173 VTAIL.n155 10.4732
R420 VTAIL.n126 VTAIL.n76 10.4732
R421 VTAIL.n105 VTAIL.n87 10.4732
R422 VTAIL.n227 VTAIL.n226 10.2747
R423 VTAIL.n23 VTAIL.n22 10.2747
R424 VTAIL.n162 VTAIL.n161 10.2747
R425 VTAIL.n94 VTAIL.n93 10.2747
R426 VTAIL.n237 VTAIL.n222 9.69747
R427 VTAIL.n264 VTAIL.n263 9.69747
R428 VTAIL.n33 VTAIL.n18 9.69747
R429 VTAIL.n60 VTAIL.n59 9.69747
R430 VTAIL.n198 VTAIL.n197 9.69747
R431 VTAIL.n172 VTAIL.n157 9.69747
R432 VTAIL.n130 VTAIL.n129 9.69747
R433 VTAIL.n104 VTAIL.n89 9.69747
R434 VTAIL.n270 VTAIL.n269 9.45567
R435 VTAIL.n66 VTAIL.n65 9.45567
R436 VTAIL.n204 VTAIL.n203 9.45567
R437 VTAIL.n136 VTAIL.n135 9.45567
R438 VTAIL.n269 VTAIL.n268 9.3005
R439 VTAIL.n208 VTAIL.n207 9.3005
R440 VTAIL.n263 VTAIL.n262 9.3005
R441 VTAIL.n261 VTAIL.n260 9.3005
R442 VTAIL.n212 VTAIL.n211 9.3005
R443 VTAIL.n255 VTAIL.n254 9.3005
R444 VTAIL.n253 VTAIL.n252 9.3005
R445 VTAIL.n229 VTAIL.n228 9.3005
R446 VTAIL.n224 VTAIL.n223 9.3005
R447 VTAIL.n235 VTAIL.n234 9.3005
R448 VTAIL.n237 VTAIL.n236 9.3005
R449 VTAIL.n220 VTAIL.n219 9.3005
R450 VTAIL.n243 VTAIL.n242 9.3005
R451 VTAIL.n245 VTAIL.n244 9.3005
R452 VTAIL.n246 VTAIL.n215 9.3005
R453 VTAIL.n65 VTAIL.n64 9.3005
R454 VTAIL.n4 VTAIL.n3 9.3005
R455 VTAIL.n59 VTAIL.n58 9.3005
R456 VTAIL.n57 VTAIL.n56 9.3005
R457 VTAIL.n8 VTAIL.n7 9.3005
R458 VTAIL.n51 VTAIL.n50 9.3005
R459 VTAIL.n49 VTAIL.n48 9.3005
R460 VTAIL.n25 VTAIL.n24 9.3005
R461 VTAIL.n20 VTAIL.n19 9.3005
R462 VTAIL.n31 VTAIL.n30 9.3005
R463 VTAIL.n33 VTAIL.n32 9.3005
R464 VTAIL.n16 VTAIL.n15 9.3005
R465 VTAIL.n39 VTAIL.n38 9.3005
R466 VTAIL.n41 VTAIL.n40 9.3005
R467 VTAIL.n42 VTAIL.n11 9.3005
R468 VTAIL.n164 VTAIL.n163 9.3005
R469 VTAIL.n159 VTAIL.n158 9.3005
R470 VTAIL.n170 VTAIL.n169 9.3005
R471 VTAIL.n172 VTAIL.n171 9.3005
R472 VTAIL.n155 VTAIL.n154 9.3005
R473 VTAIL.n178 VTAIL.n177 9.3005
R474 VTAIL.n180 VTAIL.n179 9.3005
R475 VTAIL.n152 VTAIL.n149 9.3005
R476 VTAIL.n203 VTAIL.n202 9.3005
R477 VTAIL.n142 VTAIL.n141 9.3005
R478 VTAIL.n197 VTAIL.n196 9.3005
R479 VTAIL.n195 VTAIL.n194 9.3005
R480 VTAIL.n146 VTAIL.n145 9.3005
R481 VTAIL.n189 VTAIL.n188 9.3005
R482 VTAIL.n187 VTAIL.n186 9.3005
R483 VTAIL.n96 VTAIL.n95 9.3005
R484 VTAIL.n91 VTAIL.n90 9.3005
R485 VTAIL.n102 VTAIL.n101 9.3005
R486 VTAIL.n104 VTAIL.n103 9.3005
R487 VTAIL.n87 VTAIL.n86 9.3005
R488 VTAIL.n110 VTAIL.n109 9.3005
R489 VTAIL.n112 VTAIL.n111 9.3005
R490 VTAIL.n84 VTAIL.n81 9.3005
R491 VTAIL.n135 VTAIL.n134 9.3005
R492 VTAIL.n74 VTAIL.n73 9.3005
R493 VTAIL.n129 VTAIL.n128 9.3005
R494 VTAIL.n127 VTAIL.n126 9.3005
R495 VTAIL.n78 VTAIL.n77 9.3005
R496 VTAIL.n121 VTAIL.n120 9.3005
R497 VTAIL.n119 VTAIL.n118 9.3005
R498 VTAIL.n234 VTAIL.n233 8.92171
R499 VTAIL.n267 VTAIL.n208 8.92171
R500 VTAIL.n30 VTAIL.n29 8.92171
R501 VTAIL.n63 VTAIL.n4 8.92171
R502 VTAIL.n201 VTAIL.n142 8.92171
R503 VTAIL.n169 VTAIL.n168 8.92171
R504 VTAIL.n133 VTAIL.n74 8.92171
R505 VTAIL.n101 VTAIL.n100 8.92171
R506 VTAIL.n230 VTAIL.n224 8.14595
R507 VTAIL.n268 VTAIL.n206 8.14595
R508 VTAIL.n26 VTAIL.n20 8.14595
R509 VTAIL.n64 VTAIL.n2 8.14595
R510 VTAIL.n202 VTAIL.n140 8.14595
R511 VTAIL.n165 VTAIL.n159 8.14595
R512 VTAIL.n134 VTAIL.n72 8.14595
R513 VTAIL.n97 VTAIL.n91 8.14595
R514 VTAIL.n229 VTAIL.n226 7.3702
R515 VTAIL.n25 VTAIL.n22 7.3702
R516 VTAIL.n164 VTAIL.n161 7.3702
R517 VTAIL.n96 VTAIL.n93 7.3702
R518 VTAIL.n230 VTAIL.n229 5.81868
R519 VTAIL.n270 VTAIL.n206 5.81868
R520 VTAIL.n26 VTAIL.n25 5.81868
R521 VTAIL.n66 VTAIL.n2 5.81868
R522 VTAIL.n204 VTAIL.n140 5.81868
R523 VTAIL.n165 VTAIL.n164 5.81868
R524 VTAIL.n136 VTAIL.n72 5.81868
R525 VTAIL.n97 VTAIL.n96 5.81868
R526 VTAIL.n233 VTAIL.n224 5.04292
R527 VTAIL.n268 VTAIL.n267 5.04292
R528 VTAIL.n29 VTAIL.n20 5.04292
R529 VTAIL.n64 VTAIL.n63 5.04292
R530 VTAIL.n202 VTAIL.n201 5.04292
R531 VTAIL.n168 VTAIL.n159 5.04292
R532 VTAIL.n134 VTAIL.n133 5.04292
R533 VTAIL.n100 VTAIL.n91 5.04292
R534 VTAIL.n234 VTAIL.n222 4.26717
R535 VTAIL.n264 VTAIL.n208 4.26717
R536 VTAIL.n30 VTAIL.n18 4.26717
R537 VTAIL.n60 VTAIL.n4 4.26717
R538 VTAIL.n198 VTAIL.n142 4.26717
R539 VTAIL.n169 VTAIL.n157 4.26717
R540 VTAIL.n130 VTAIL.n74 4.26717
R541 VTAIL.n101 VTAIL.n89 4.26717
R542 VTAIL.n238 VTAIL.n237 3.49141
R543 VTAIL.n263 VTAIL.n210 3.49141
R544 VTAIL.n34 VTAIL.n33 3.49141
R545 VTAIL.n59 VTAIL.n6 3.49141
R546 VTAIL.n197 VTAIL.n144 3.49141
R547 VTAIL.n173 VTAIL.n172 3.49141
R548 VTAIL.n129 VTAIL.n76 3.49141
R549 VTAIL.n105 VTAIL.n104 3.49141
R550 VTAIL.n228 VTAIL.n227 2.84303
R551 VTAIL.n24 VTAIL.n23 2.84303
R552 VTAIL.n163 VTAIL.n162 2.84303
R553 VTAIL.n95 VTAIL.n94 2.84303
R554 VTAIL.n241 VTAIL.n220 2.71565
R555 VTAIL.n260 VTAIL.n259 2.71565
R556 VTAIL.n37 VTAIL.n16 2.71565
R557 VTAIL.n56 VTAIL.n55 2.71565
R558 VTAIL.n194 VTAIL.n193 2.71565
R559 VTAIL.n176 VTAIL.n155 2.71565
R560 VTAIL.n126 VTAIL.n125 2.71565
R561 VTAIL.n108 VTAIL.n87 2.71565
R562 VTAIL.n242 VTAIL.n218 1.93989
R563 VTAIL.n256 VTAIL.n212 1.93989
R564 VTAIL.n38 VTAIL.n14 1.93989
R565 VTAIL.n52 VTAIL.n8 1.93989
R566 VTAIL.n190 VTAIL.n146 1.93989
R567 VTAIL.n177 VTAIL.n153 1.93989
R568 VTAIL.n122 VTAIL.n78 1.93989
R569 VTAIL.n109 VTAIL.n85 1.93989
R570 VTAIL.n0 VTAIL.t9 1.63957
R571 VTAIL.n0 VTAIL.t10 1.63957
R572 VTAIL.n68 VTAIL.t1 1.63957
R573 VTAIL.n68 VTAIL.t2 1.63957
R574 VTAIL.n138 VTAIL.t5 1.63957
R575 VTAIL.n138 VTAIL.t0 1.63957
R576 VTAIL.n70 VTAIL.t8 1.63957
R577 VTAIL.n70 VTAIL.t11 1.63957
R578 VTAIL.n137 VTAIL.n71 1.5436
R579 VTAIL.n205 VTAIL.n139 1.5436
R580 VTAIL.n69 VTAIL.n67 1.5436
R581 VTAIL.n139 VTAIL.n137 1.24188
R582 VTAIL.n67 VTAIL.n1 1.24188
R583 VTAIL.n247 VTAIL.n245 1.16414
R584 VTAIL.n255 VTAIL.n214 1.16414
R585 VTAIL.n43 VTAIL.n41 1.16414
R586 VTAIL.n51 VTAIL.n10 1.16414
R587 VTAIL.n189 VTAIL.n148 1.16414
R588 VTAIL.n181 VTAIL.n180 1.16414
R589 VTAIL.n121 VTAIL.n80 1.16414
R590 VTAIL.n113 VTAIL.n112 1.16414
R591 VTAIL VTAIL.n271 1.09964
R592 VTAIL VTAIL.n1 0.444466
R593 VTAIL.n246 VTAIL.n216 0.388379
R594 VTAIL.n252 VTAIL.n251 0.388379
R595 VTAIL.n42 VTAIL.n12 0.388379
R596 VTAIL.n48 VTAIL.n47 0.388379
R597 VTAIL.n186 VTAIL.n185 0.388379
R598 VTAIL.n152 VTAIL.n150 0.388379
R599 VTAIL.n118 VTAIL.n117 0.388379
R600 VTAIL.n84 VTAIL.n82 0.388379
R601 VTAIL.n228 VTAIL.n223 0.155672
R602 VTAIL.n235 VTAIL.n223 0.155672
R603 VTAIL.n236 VTAIL.n235 0.155672
R604 VTAIL.n236 VTAIL.n219 0.155672
R605 VTAIL.n243 VTAIL.n219 0.155672
R606 VTAIL.n244 VTAIL.n243 0.155672
R607 VTAIL.n244 VTAIL.n215 0.155672
R608 VTAIL.n253 VTAIL.n215 0.155672
R609 VTAIL.n254 VTAIL.n253 0.155672
R610 VTAIL.n254 VTAIL.n211 0.155672
R611 VTAIL.n261 VTAIL.n211 0.155672
R612 VTAIL.n262 VTAIL.n261 0.155672
R613 VTAIL.n262 VTAIL.n207 0.155672
R614 VTAIL.n269 VTAIL.n207 0.155672
R615 VTAIL.n24 VTAIL.n19 0.155672
R616 VTAIL.n31 VTAIL.n19 0.155672
R617 VTAIL.n32 VTAIL.n31 0.155672
R618 VTAIL.n32 VTAIL.n15 0.155672
R619 VTAIL.n39 VTAIL.n15 0.155672
R620 VTAIL.n40 VTAIL.n39 0.155672
R621 VTAIL.n40 VTAIL.n11 0.155672
R622 VTAIL.n49 VTAIL.n11 0.155672
R623 VTAIL.n50 VTAIL.n49 0.155672
R624 VTAIL.n50 VTAIL.n7 0.155672
R625 VTAIL.n57 VTAIL.n7 0.155672
R626 VTAIL.n58 VTAIL.n57 0.155672
R627 VTAIL.n58 VTAIL.n3 0.155672
R628 VTAIL.n65 VTAIL.n3 0.155672
R629 VTAIL.n203 VTAIL.n141 0.155672
R630 VTAIL.n196 VTAIL.n141 0.155672
R631 VTAIL.n196 VTAIL.n195 0.155672
R632 VTAIL.n195 VTAIL.n145 0.155672
R633 VTAIL.n188 VTAIL.n145 0.155672
R634 VTAIL.n188 VTAIL.n187 0.155672
R635 VTAIL.n187 VTAIL.n149 0.155672
R636 VTAIL.n179 VTAIL.n149 0.155672
R637 VTAIL.n179 VTAIL.n178 0.155672
R638 VTAIL.n178 VTAIL.n154 0.155672
R639 VTAIL.n171 VTAIL.n154 0.155672
R640 VTAIL.n171 VTAIL.n170 0.155672
R641 VTAIL.n170 VTAIL.n158 0.155672
R642 VTAIL.n163 VTAIL.n158 0.155672
R643 VTAIL.n135 VTAIL.n73 0.155672
R644 VTAIL.n128 VTAIL.n73 0.155672
R645 VTAIL.n128 VTAIL.n127 0.155672
R646 VTAIL.n127 VTAIL.n77 0.155672
R647 VTAIL.n120 VTAIL.n77 0.155672
R648 VTAIL.n120 VTAIL.n119 0.155672
R649 VTAIL.n119 VTAIL.n81 0.155672
R650 VTAIL.n111 VTAIL.n81 0.155672
R651 VTAIL.n111 VTAIL.n110 0.155672
R652 VTAIL.n110 VTAIL.n86 0.155672
R653 VTAIL.n103 VTAIL.n86 0.155672
R654 VTAIL.n103 VTAIL.n102 0.155672
R655 VTAIL.n102 VTAIL.n90 0.155672
R656 VTAIL.n95 VTAIL.n90 0.155672
R657 B.n711 B.n710 585
R658 B.n712 B.n711 585
R659 B.n291 B.n102 585
R660 B.n290 B.n289 585
R661 B.n288 B.n287 585
R662 B.n286 B.n285 585
R663 B.n284 B.n283 585
R664 B.n282 B.n281 585
R665 B.n280 B.n279 585
R666 B.n278 B.n277 585
R667 B.n276 B.n275 585
R668 B.n274 B.n273 585
R669 B.n272 B.n271 585
R670 B.n270 B.n269 585
R671 B.n268 B.n267 585
R672 B.n266 B.n265 585
R673 B.n264 B.n263 585
R674 B.n262 B.n261 585
R675 B.n260 B.n259 585
R676 B.n258 B.n257 585
R677 B.n256 B.n255 585
R678 B.n254 B.n253 585
R679 B.n252 B.n251 585
R680 B.n250 B.n249 585
R681 B.n248 B.n247 585
R682 B.n246 B.n245 585
R683 B.n244 B.n243 585
R684 B.n242 B.n241 585
R685 B.n240 B.n239 585
R686 B.n238 B.n237 585
R687 B.n236 B.n235 585
R688 B.n234 B.n233 585
R689 B.n232 B.n231 585
R690 B.n230 B.n229 585
R691 B.n228 B.n227 585
R692 B.n226 B.n225 585
R693 B.n224 B.n223 585
R694 B.n222 B.n221 585
R695 B.n220 B.n219 585
R696 B.n218 B.n217 585
R697 B.n216 B.n215 585
R698 B.n214 B.n213 585
R699 B.n212 B.n211 585
R700 B.n209 B.n208 585
R701 B.n207 B.n206 585
R702 B.n205 B.n204 585
R703 B.n203 B.n202 585
R704 B.n201 B.n200 585
R705 B.n199 B.n198 585
R706 B.n197 B.n196 585
R707 B.n195 B.n194 585
R708 B.n193 B.n192 585
R709 B.n191 B.n190 585
R710 B.n189 B.n188 585
R711 B.n187 B.n186 585
R712 B.n185 B.n184 585
R713 B.n183 B.n182 585
R714 B.n181 B.n180 585
R715 B.n179 B.n178 585
R716 B.n177 B.n176 585
R717 B.n175 B.n174 585
R718 B.n173 B.n172 585
R719 B.n171 B.n170 585
R720 B.n169 B.n168 585
R721 B.n167 B.n166 585
R722 B.n165 B.n164 585
R723 B.n163 B.n162 585
R724 B.n161 B.n160 585
R725 B.n159 B.n158 585
R726 B.n157 B.n156 585
R727 B.n155 B.n154 585
R728 B.n153 B.n152 585
R729 B.n151 B.n150 585
R730 B.n149 B.n148 585
R731 B.n147 B.n146 585
R732 B.n145 B.n144 585
R733 B.n143 B.n142 585
R734 B.n141 B.n140 585
R735 B.n139 B.n138 585
R736 B.n137 B.n136 585
R737 B.n135 B.n134 585
R738 B.n133 B.n132 585
R739 B.n131 B.n130 585
R740 B.n129 B.n128 585
R741 B.n127 B.n126 585
R742 B.n125 B.n124 585
R743 B.n123 B.n122 585
R744 B.n121 B.n120 585
R745 B.n119 B.n118 585
R746 B.n117 B.n116 585
R747 B.n115 B.n114 585
R748 B.n113 B.n112 585
R749 B.n111 B.n110 585
R750 B.n109 B.n108 585
R751 B.n709 B.n55 585
R752 B.n713 B.n55 585
R753 B.n708 B.n54 585
R754 B.n714 B.n54 585
R755 B.n707 B.n706 585
R756 B.n706 B.n50 585
R757 B.n705 B.n49 585
R758 B.n720 B.n49 585
R759 B.n704 B.n48 585
R760 B.n721 B.n48 585
R761 B.n703 B.n47 585
R762 B.n722 B.n47 585
R763 B.n702 B.n701 585
R764 B.n701 B.n43 585
R765 B.n700 B.n42 585
R766 B.n728 B.n42 585
R767 B.n699 B.n41 585
R768 B.n729 B.n41 585
R769 B.n698 B.n40 585
R770 B.n730 B.n40 585
R771 B.n697 B.n696 585
R772 B.n696 B.n36 585
R773 B.n695 B.n35 585
R774 B.n736 B.n35 585
R775 B.n694 B.n34 585
R776 B.n737 B.n34 585
R777 B.n693 B.n33 585
R778 B.n738 B.n33 585
R779 B.n692 B.n691 585
R780 B.n691 B.n32 585
R781 B.n690 B.n28 585
R782 B.n744 B.n28 585
R783 B.n689 B.n27 585
R784 B.n745 B.n27 585
R785 B.n688 B.n26 585
R786 B.n746 B.n26 585
R787 B.n687 B.n686 585
R788 B.n686 B.n22 585
R789 B.n685 B.n21 585
R790 B.n752 B.n21 585
R791 B.n684 B.n20 585
R792 B.n753 B.n20 585
R793 B.n683 B.n19 585
R794 B.n754 B.n19 585
R795 B.n682 B.n681 585
R796 B.n681 B.n15 585
R797 B.n680 B.n14 585
R798 B.n760 B.n14 585
R799 B.n679 B.n13 585
R800 B.n761 B.n13 585
R801 B.n678 B.n12 585
R802 B.n762 B.n12 585
R803 B.n677 B.n676 585
R804 B.n676 B.n8 585
R805 B.n675 B.n7 585
R806 B.n768 B.n7 585
R807 B.n674 B.n6 585
R808 B.n769 B.n6 585
R809 B.n673 B.n5 585
R810 B.n770 B.n5 585
R811 B.n672 B.n671 585
R812 B.n671 B.n4 585
R813 B.n670 B.n292 585
R814 B.n670 B.n669 585
R815 B.n660 B.n293 585
R816 B.n294 B.n293 585
R817 B.n662 B.n661 585
R818 B.n663 B.n662 585
R819 B.n659 B.n298 585
R820 B.n302 B.n298 585
R821 B.n658 B.n657 585
R822 B.n657 B.n656 585
R823 B.n300 B.n299 585
R824 B.n301 B.n300 585
R825 B.n649 B.n648 585
R826 B.n650 B.n649 585
R827 B.n647 B.n307 585
R828 B.n307 B.n306 585
R829 B.n646 B.n645 585
R830 B.n645 B.n644 585
R831 B.n309 B.n308 585
R832 B.n310 B.n309 585
R833 B.n637 B.n636 585
R834 B.n638 B.n637 585
R835 B.n635 B.n315 585
R836 B.n315 B.n314 585
R837 B.n634 B.n633 585
R838 B.n633 B.n632 585
R839 B.n317 B.n316 585
R840 B.n625 B.n317 585
R841 B.n624 B.n623 585
R842 B.n626 B.n624 585
R843 B.n622 B.n322 585
R844 B.n322 B.n321 585
R845 B.n621 B.n620 585
R846 B.n620 B.n619 585
R847 B.n324 B.n323 585
R848 B.n325 B.n324 585
R849 B.n612 B.n611 585
R850 B.n613 B.n612 585
R851 B.n610 B.n330 585
R852 B.n330 B.n329 585
R853 B.n609 B.n608 585
R854 B.n608 B.n607 585
R855 B.n332 B.n331 585
R856 B.n333 B.n332 585
R857 B.n600 B.n599 585
R858 B.n601 B.n600 585
R859 B.n598 B.n338 585
R860 B.n338 B.n337 585
R861 B.n597 B.n596 585
R862 B.n596 B.n595 585
R863 B.n340 B.n339 585
R864 B.n341 B.n340 585
R865 B.n588 B.n587 585
R866 B.n589 B.n588 585
R867 B.n586 B.n346 585
R868 B.n346 B.n345 585
R869 B.n580 B.n579 585
R870 B.n578 B.n394 585
R871 B.n577 B.n393 585
R872 B.n582 B.n393 585
R873 B.n576 B.n575 585
R874 B.n574 B.n573 585
R875 B.n572 B.n571 585
R876 B.n570 B.n569 585
R877 B.n568 B.n567 585
R878 B.n566 B.n565 585
R879 B.n564 B.n563 585
R880 B.n562 B.n561 585
R881 B.n560 B.n559 585
R882 B.n558 B.n557 585
R883 B.n556 B.n555 585
R884 B.n554 B.n553 585
R885 B.n552 B.n551 585
R886 B.n550 B.n549 585
R887 B.n548 B.n547 585
R888 B.n546 B.n545 585
R889 B.n544 B.n543 585
R890 B.n542 B.n541 585
R891 B.n540 B.n539 585
R892 B.n538 B.n537 585
R893 B.n536 B.n535 585
R894 B.n534 B.n533 585
R895 B.n532 B.n531 585
R896 B.n530 B.n529 585
R897 B.n528 B.n527 585
R898 B.n526 B.n525 585
R899 B.n524 B.n523 585
R900 B.n522 B.n521 585
R901 B.n520 B.n519 585
R902 B.n518 B.n517 585
R903 B.n516 B.n515 585
R904 B.n514 B.n513 585
R905 B.n512 B.n511 585
R906 B.n510 B.n509 585
R907 B.n508 B.n507 585
R908 B.n506 B.n505 585
R909 B.n504 B.n503 585
R910 B.n502 B.n501 585
R911 B.n500 B.n499 585
R912 B.n497 B.n496 585
R913 B.n495 B.n494 585
R914 B.n493 B.n492 585
R915 B.n491 B.n490 585
R916 B.n489 B.n488 585
R917 B.n487 B.n486 585
R918 B.n485 B.n484 585
R919 B.n483 B.n482 585
R920 B.n481 B.n480 585
R921 B.n479 B.n478 585
R922 B.n477 B.n476 585
R923 B.n475 B.n474 585
R924 B.n473 B.n472 585
R925 B.n471 B.n470 585
R926 B.n469 B.n468 585
R927 B.n467 B.n466 585
R928 B.n465 B.n464 585
R929 B.n463 B.n462 585
R930 B.n461 B.n460 585
R931 B.n459 B.n458 585
R932 B.n457 B.n456 585
R933 B.n455 B.n454 585
R934 B.n453 B.n452 585
R935 B.n451 B.n450 585
R936 B.n449 B.n448 585
R937 B.n447 B.n446 585
R938 B.n445 B.n444 585
R939 B.n443 B.n442 585
R940 B.n441 B.n440 585
R941 B.n439 B.n438 585
R942 B.n437 B.n436 585
R943 B.n435 B.n434 585
R944 B.n433 B.n432 585
R945 B.n431 B.n430 585
R946 B.n429 B.n428 585
R947 B.n427 B.n426 585
R948 B.n425 B.n424 585
R949 B.n423 B.n422 585
R950 B.n421 B.n420 585
R951 B.n419 B.n418 585
R952 B.n417 B.n416 585
R953 B.n415 B.n414 585
R954 B.n413 B.n412 585
R955 B.n411 B.n410 585
R956 B.n409 B.n408 585
R957 B.n407 B.n406 585
R958 B.n405 B.n404 585
R959 B.n403 B.n402 585
R960 B.n401 B.n400 585
R961 B.n348 B.n347 585
R962 B.n585 B.n584 585
R963 B.n344 B.n343 585
R964 B.n345 B.n344 585
R965 B.n591 B.n590 585
R966 B.n590 B.n589 585
R967 B.n592 B.n342 585
R968 B.n342 B.n341 585
R969 B.n594 B.n593 585
R970 B.n595 B.n594 585
R971 B.n336 B.n335 585
R972 B.n337 B.n336 585
R973 B.n603 B.n602 585
R974 B.n602 B.n601 585
R975 B.n604 B.n334 585
R976 B.n334 B.n333 585
R977 B.n606 B.n605 585
R978 B.n607 B.n606 585
R979 B.n328 B.n327 585
R980 B.n329 B.n328 585
R981 B.n615 B.n614 585
R982 B.n614 B.n613 585
R983 B.n616 B.n326 585
R984 B.n326 B.n325 585
R985 B.n618 B.n617 585
R986 B.n619 B.n618 585
R987 B.n320 B.n319 585
R988 B.n321 B.n320 585
R989 B.n628 B.n627 585
R990 B.n627 B.n626 585
R991 B.n629 B.n318 585
R992 B.n625 B.n318 585
R993 B.n631 B.n630 585
R994 B.n632 B.n631 585
R995 B.n313 B.n312 585
R996 B.n314 B.n313 585
R997 B.n640 B.n639 585
R998 B.n639 B.n638 585
R999 B.n641 B.n311 585
R1000 B.n311 B.n310 585
R1001 B.n643 B.n642 585
R1002 B.n644 B.n643 585
R1003 B.n305 B.n304 585
R1004 B.n306 B.n305 585
R1005 B.n652 B.n651 585
R1006 B.n651 B.n650 585
R1007 B.n653 B.n303 585
R1008 B.n303 B.n301 585
R1009 B.n655 B.n654 585
R1010 B.n656 B.n655 585
R1011 B.n297 B.n296 585
R1012 B.n302 B.n297 585
R1013 B.n665 B.n664 585
R1014 B.n664 B.n663 585
R1015 B.n666 B.n295 585
R1016 B.n295 B.n294 585
R1017 B.n668 B.n667 585
R1018 B.n669 B.n668 585
R1019 B.n2 B.n0 585
R1020 B.n4 B.n2 585
R1021 B.n3 B.n1 585
R1022 B.n769 B.n3 585
R1023 B.n767 B.n766 585
R1024 B.n768 B.n767 585
R1025 B.n765 B.n9 585
R1026 B.n9 B.n8 585
R1027 B.n764 B.n763 585
R1028 B.n763 B.n762 585
R1029 B.n11 B.n10 585
R1030 B.n761 B.n11 585
R1031 B.n759 B.n758 585
R1032 B.n760 B.n759 585
R1033 B.n757 B.n16 585
R1034 B.n16 B.n15 585
R1035 B.n756 B.n755 585
R1036 B.n755 B.n754 585
R1037 B.n18 B.n17 585
R1038 B.n753 B.n18 585
R1039 B.n751 B.n750 585
R1040 B.n752 B.n751 585
R1041 B.n749 B.n23 585
R1042 B.n23 B.n22 585
R1043 B.n748 B.n747 585
R1044 B.n747 B.n746 585
R1045 B.n25 B.n24 585
R1046 B.n745 B.n25 585
R1047 B.n743 B.n742 585
R1048 B.n744 B.n743 585
R1049 B.n741 B.n29 585
R1050 B.n32 B.n29 585
R1051 B.n740 B.n739 585
R1052 B.n739 B.n738 585
R1053 B.n31 B.n30 585
R1054 B.n737 B.n31 585
R1055 B.n735 B.n734 585
R1056 B.n736 B.n735 585
R1057 B.n733 B.n37 585
R1058 B.n37 B.n36 585
R1059 B.n732 B.n731 585
R1060 B.n731 B.n730 585
R1061 B.n39 B.n38 585
R1062 B.n729 B.n39 585
R1063 B.n727 B.n726 585
R1064 B.n728 B.n727 585
R1065 B.n725 B.n44 585
R1066 B.n44 B.n43 585
R1067 B.n724 B.n723 585
R1068 B.n723 B.n722 585
R1069 B.n46 B.n45 585
R1070 B.n721 B.n46 585
R1071 B.n719 B.n718 585
R1072 B.n720 B.n719 585
R1073 B.n717 B.n51 585
R1074 B.n51 B.n50 585
R1075 B.n716 B.n715 585
R1076 B.n715 B.n714 585
R1077 B.n53 B.n52 585
R1078 B.n713 B.n53 585
R1079 B.n772 B.n771 585
R1080 B.n771 B.n770 585
R1081 B.n580 B.n344 550.159
R1082 B.n108 B.n53 550.159
R1083 B.n584 B.n346 550.159
R1084 B.n711 B.n55 550.159
R1085 B.n397 B.t6 404.69
R1086 B.n395 B.t17 404.69
R1087 B.n105 B.t10 404.69
R1088 B.n103 B.t14 404.69
R1089 B.n397 B.t9 318.274
R1090 B.n103 B.t15 318.274
R1091 B.n395 B.t19 318.274
R1092 B.n105 B.t12 318.274
R1093 B.n398 B.t8 283.56
R1094 B.n104 B.t16 283.56
R1095 B.n396 B.t18 283.56
R1096 B.n106 B.t13 283.56
R1097 B.n712 B.n101 256.663
R1098 B.n712 B.n100 256.663
R1099 B.n712 B.n99 256.663
R1100 B.n712 B.n98 256.663
R1101 B.n712 B.n97 256.663
R1102 B.n712 B.n96 256.663
R1103 B.n712 B.n95 256.663
R1104 B.n712 B.n94 256.663
R1105 B.n712 B.n93 256.663
R1106 B.n712 B.n92 256.663
R1107 B.n712 B.n91 256.663
R1108 B.n712 B.n90 256.663
R1109 B.n712 B.n89 256.663
R1110 B.n712 B.n88 256.663
R1111 B.n712 B.n87 256.663
R1112 B.n712 B.n86 256.663
R1113 B.n712 B.n85 256.663
R1114 B.n712 B.n84 256.663
R1115 B.n712 B.n83 256.663
R1116 B.n712 B.n82 256.663
R1117 B.n712 B.n81 256.663
R1118 B.n712 B.n80 256.663
R1119 B.n712 B.n79 256.663
R1120 B.n712 B.n78 256.663
R1121 B.n712 B.n77 256.663
R1122 B.n712 B.n76 256.663
R1123 B.n712 B.n75 256.663
R1124 B.n712 B.n74 256.663
R1125 B.n712 B.n73 256.663
R1126 B.n712 B.n72 256.663
R1127 B.n712 B.n71 256.663
R1128 B.n712 B.n70 256.663
R1129 B.n712 B.n69 256.663
R1130 B.n712 B.n68 256.663
R1131 B.n712 B.n67 256.663
R1132 B.n712 B.n66 256.663
R1133 B.n712 B.n65 256.663
R1134 B.n712 B.n64 256.663
R1135 B.n712 B.n63 256.663
R1136 B.n712 B.n62 256.663
R1137 B.n712 B.n61 256.663
R1138 B.n712 B.n60 256.663
R1139 B.n712 B.n59 256.663
R1140 B.n712 B.n58 256.663
R1141 B.n712 B.n57 256.663
R1142 B.n712 B.n56 256.663
R1143 B.n582 B.n581 256.663
R1144 B.n582 B.n349 256.663
R1145 B.n582 B.n350 256.663
R1146 B.n582 B.n351 256.663
R1147 B.n582 B.n352 256.663
R1148 B.n582 B.n353 256.663
R1149 B.n582 B.n354 256.663
R1150 B.n582 B.n355 256.663
R1151 B.n582 B.n356 256.663
R1152 B.n582 B.n357 256.663
R1153 B.n582 B.n358 256.663
R1154 B.n582 B.n359 256.663
R1155 B.n582 B.n360 256.663
R1156 B.n582 B.n361 256.663
R1157 B.n582 B.n362 256.663
R1158 B.n582 B.n363 256.663
R1159 B.n582 B.n364 256.663
R1160 B.n582 B.n365 256.663
R1161 B.n582 B.n366 256.663
R1162 B.n582 B.n367 256.663
R1163 B.n582 B.n368 256.663
R1164 B.n582 B.n369 256.663
R1165 B.n582 B.n370 256.663
R1166 B.n582 B.n371 256.663
R1167 B.n582 B.n372 256.663
R1168 B.n582 B.n373 256.663
R1169 B.n582 B.n374 256.663
R1170 B.n582 B.n375 256.663
R1171 B.n582 B.n376 256.663
R1172 B.n582 B.n377 256.663
R1173 B.n582 B.n378 256.663
R1174 B.n582 B.n379 256.663
R1175 B.n582 B.n380 256.663
R1176 B.n582 B.n381 256.663
R1177 B.n582 B.n382 256.663
R1178 B.n582 B.n383 256.663
R1179 B.n582 B.n384 256.663
R1180 B.n582 B.n385 256.663
R1181 B.n582 B.n386 256.663
R1182 B.n582 B.n387 256.663
R1183 B.n582 B.n388 256.663
R1184 B.n582 B.n389 256.663
R1185 B.n582 B.n390 256.663
R1186 B.n582 B.n391 256.663
R1187 B.n582 B.n392 256.663
R1188 B.n583 B.n582 256.663
R1189 B.n590 B.n344 163.367
R1190 B.n590 B.n342 163.367
R1191 B.n594 B.n342 163.367
R1192 B.n594 B.n336 163.367
R1193 B.n602 B.n336 163.367
R1194 B.n602 B.n334 163.367
R1195 B.n606 B.n334 163.367
R1196 B.n606 B.n328 163.367
R1197 B.n614 B.n328 163.367
R1198 B.n614 B.n326 163.367
R1199 B.n618 B.n326 163.367
R1200 B.n618 B.n320 163.367
R1201 B.n627 B.n320 163.367
R1202 B.n627 B.n318 163.367
R1203 B.n631 B.n318 163.367
R1204 B.n631 B.n313 163.367
R1205 B.n639 B.n313 163.367
R1206 B.n639 B.n311 163.367
R1207 B.n643 B.n311 163.367
R1208 B.n643 B.n305 163.367
R1209 B.n651 B.n305 163.367
R1210 B.n651 B.n303 163.367
R1211 B.n655 B.n303 163.367
R1212 B.n655 B.n297 163.367
R1213 B.n664 B.n297 163.367
R1214 B.n664 B.n295 163.367
R1215 B.n668 B.n295 163.367
R1216 B.n668 B.n2 163.367
R1217 B.n771 B.n2 163.367
R1218 B.n771 B.n3 163.367
R1219 B.n767 B.n3 163.367
R1220 B.n767 B.n9 163.367
R1221 B.n763 B.n9 163.367
R1222 B.n763 B.n11 163.367
R1223 B.n759 B.n11 163.367
R1224 B.n759 B.n16 163.367
R1225 B.n755 B.n16 163.367
R1226 B.n755 B.n18 163.367
R1227 B.n751 B.n18 163.367
R1228 B.n751 B.n23 163.367
R1229 B.n747 B.n23 163.367
R1230 B.n747 B.n25 163.367
R1231 B.n743 B.n25 163.367
R1232 B.n743 B.n29 163.367
R1233 B.n739 B.n29 163.367
R1234 B.n739 B.n31 163.367
R1235 B.n735 B.n31 163.367
R1236 B.n735 B.n37 163.367
R1237 B.n731 B.n37 163.367
R1238 B.n731 B.n39 163.367
R1239 B.n727 B.n39 163.367
R1240 B.n727 B.n44 163.367
R1241 B.n723 B.n44 163.367
R1242 B.n723 B.n46 163.367
R1243 B.n719 B.n46 163.367
R1244 B.n719 B.n51 163.367
R1245 B.n715 B.n51 163.367
R1246 B.n715 B.n53 163.367
R1247 B.n394 B.n393 163.367
R1248 B.n575 B.n393 163.367
R1249 B.n573 B.n572 163.367
R1250 B.n569 B.n568 163.367
R1251 B.n565 B.n564 163.367
R1252 B.n561 B.n560 163.367
R1253 B.n557 B.n556 163.367
R1254 B.n553 B.n552 163.367
R1255 B.n549 B.n548 163.367
R1256 B.n545 B.n544 163.367
R1257 B.n541 B.n540 163.367
R1258 B.n537 B.n536 163.367
R1259 B.n533 B.n532 163.367
R1260 B.n529 B.n528 163.367
R1261 B.n525 B.n524 163.367
R1262 B.n521 B.n520 163.367
R1263 B.n517 B.n516 163.367
R1264 B.n513 B.n512 163.367
R1265 B.n509 B.n508 163.367
R1266 B.n505 B.n504 163.367
R1267 B.n501 B.n500 163.367
R1268 B.n496 B.n495 163.367
R1269 B.n492 B.n491 163.367
R1270 B.n488 B.n487 163.367
R1271 B.n484 B.n483 163.367
R1272 B.n480 B.n479 163.367
R1273 B.n476 B.n475 163.367
R1274 B.n472 B.n471 163.367
R1275 B.n468 B.n467 163.367
R1276 B.n464 B.n463 163.367
R1277 B.n460 B.n459 163.367
R1278 B.n456 B.n455 163.367
R1279 B.n452 B.n451 163.367
R1280 B.n448 B.n447 163.367
R1281 B.n444 B.n443 163.367
R1282 B.n440 B.n439 163.367
R1283 B.n436 B.n435 163.367
R1284 B.n432 B.n431 163.367
R1285 B.n428 B.n427 163.367
R1286 B.n424 B.n423 163.367
R1287 B.n420 B.n419 163.367
R1288 B.n416 B.n415 163.367
R1289 B.n412 B.n411 163.367
R1290 B.n408 B.n407 163.367
R1291 B.n404 B.n403 163.367
R1292 B.n400 B.n348 163.367
R1293 B.n588 B.n346 163.367
R1294 B.n588 B.n340 163.367
R1295 B.n596 B.n340 163.367
R1296 B.n596 B.n338 163.367
R1297 B.n600 B.n338 163.367
R1298 B.n600 B.n332 163.367
R1299 B.n608 B.n332 163.367
R1300 B.n608 B.n330 163.367
R1301 B.n612 B.n330 163.367
R1302 B.n612 B.n324 163.367
R1303 B.n620 B.n324 163.367
R1304 B.n620 B.n322 163.367
R1305 B.n624 B.n322 163.367
R1306 B.n624 B.n317 163.367
R1307 B.n633 B.n317 163.367
R1308 B.n633 B.n315 163.367
R1309 B.n637 B.n315 163.367
R1310 B.n637 B.n309 163.367
R1311 B.n645 B.n309 163.367
R1312 B.n645 B.n307 163.367
R1313 B.n649 B.n307 163.367
R1314 B.n649 B.n300 163.367
R1315 B.n657 B.n300 163.367
R1316 B.n657 B.n298 163.367
R1317 B.n662 B.n298 163.367
R1318 B.n662 B.n293 163.367
R1319 B.n670 B.n293 163.367
R1320 B.n671 B.n670 163.367
R1321 B.n671 B.n5 163.367
R1322 B.n6 B.n5 163.367
R1323 B.n7 B.n6 163.367
R1324 B.n676 B.n7 163.367
R1325 B.n676 B.n12 163.367
R1326 B.n13 B.n12 163.367
R1327 B.n14 B.n13 163.367
R1328 B.n681 B.n14 163.367
R1329 B.n681 B.n19 163.367
R1330 B.n20 B.n19 163.367
R1331 B.n21 B.n20 163.367
R1332 B.n686 B.n21 163.367
R1333 B.n686 B.n26 163.367
R1334 B.n27 B.n26 163.367
R1335 B.n28 B.n27 163.367
R1336 B.n691 B.n28 163.367
R1337 B.n691 B.n33 163.367
R1338 B.n34 B.n33 163.367
R1339 B.n35 B.n34 163.367
R1340 B.n696 B.n35 163.367
R1341 B.n696 B.n40 163.367
R1342 B.n41 B.n40 163.367
R1343 B.n42 B.n41 163.367
R1344 B.n701 B.n42 163.367
R1345 B.n701 B.n47 163.367
R1346 B.n48 B.n47 163.367
R1347 B.n49 B.n48 163.367
R1348 B.n706 B.n49 163.367
R1349 B.n706 B.n54 163.367
R1350 B.n55 B.n54 163.367
R1351 B.n112 B.n111 163.367
R1352 B.n116 B.n115 163.367
R1353 B.n120 B.n119 163.367
R1354 B.n124 B.n123 163.367
R1355 B.n128 B.n127 163.367
R1356 B.n132 B.n131 163.367
R1357 B.n136 B.n135 163.367
R1358 B.n140 B.n139 163.367
R1359 B.n144 B.n143 163.367
R1360 B.n148 B.n147 163.367
R1361 B.n152 B.n151 163.367
R1362 B.n156 B.n155 163.367
R1363 B.n160 B.n159 163.367
R1364 B.n164 B.n163 163.367
R1365 B.n168 B.n167 163.367
R1366 B.n172 B.n171 163.367
R1367 B.n176 B.n175 163.367
R1368 B.n180 B.n179 163.367
R1369 B.n184 B.n183 163.367
R1370 B.n188 B.n187 163.367
R1371 B.n192 B.n191 163.367
R1372 B.n196 B.n195 163.367
R1373 B.n200 B.n199 163.367
R1374 B.n204 B.n203 163.367
R1375 B.n208 B.n207 163.367
R1376 B.n213 B.n212 163.367
R1377 B.n217 B.n216 163.367
R1378 B.n221 B.n220 163.367
R1379 B.n225 B.n224 163.367
R1380 B.n229 B.n228 163.367
R1381 B.n233 B.n232 163.367
R1382 B.n237 B.n236 163.367
R1383 B.n241 B.n240 163.367
R1384 B.n245 B.n244 163.367
R1385 B.n249 B.n248 163.367
R1386 B.n253 B.n252 163.367
R1387 B.n257 B.n256 163.367
R1388 B.n261 B.n260 163.367
R1389 B.n265 B.n264 163.367
R1390 B.n269 B.n268 163.367
R1391 B.n273 B.n272 163.367
R1392 B.n277 B.n276 163.367
R1393 B.n281 B.n280 163.367
R1394 B.n285 B.n284 163.367
R1395 B.n289 B.n288 163.367
R1396 B.n711 B.n102 163.367
R1397 B.n582 B.n345 85.5666
R1398 B.n713 B.n712 85.5666
R1399 B.n581 B.n580 71.676
R1400 B.n575 B.n349 71.676
R1401 B.n572 B.n350 71.676
R1402 B.n568 B.n351 71.676
R1403 B.n564 B.n352 71.676
R1404 B.n560 B.n353 71.676
R1405 B.n556 B.n354 71.676
R1406 B.n552 B.n355 71.676
R1407 B.n548 B.n356 71.676
R1408 B.n544 B.n357 71.676
R1409 B.n540 B.n358 71.676
R1410 B.n536 B.n359 71.676
R1411 B.n532 B.n360 71.676
R1412 B.n528 B.n361 71.676
R1413 B.n524 B.n362 71.676
R1414 B.n520 B.n363 71.676
R1415 B.n516 B.n364 71.676
R1416 B.n512 B.n365 71.676
R1417 B.n508 B.n366 71.676
R1418 B.n504 B.n367 71.676
R1419 B.n500 B.n368 71.676
R1420 B.n495 B.n369 71.676
R1421 B.n491 B.n370 71.676
R1422 B.n487 B.n371 71.676
R1423 B.n483 B.n372 71.676
R1424 B.n479 B.n373 71.676
R1425 B.n475 B.n374 71.676
R1426 B.n471 B.n375 71.676
R1427 B.n467 B.n376 71.676
R1428 B.n463 B.n377 71.676
R1429 B.n459 B.n378 71.676
R1430 B.n455 B.n379 71.676
R1431 B.n451 B.n380 71.676
R1432 B.n447 B.n381 71.676
R1433 B.n443 B.n382 71.676
R1434 B.n439 B.n383 71.676
R1435 B.n435 B.n384 71.676
R1436 B.n431 B.n385 71.676
R1437 B.n427 B.n386 71.676
R1438 B.n423 B.n387 71.676
R1439 B.n419 B.n388 71.676
R1440 B.n415 B.n389 71.676
R1441 B.n411 B.n390 71.676
R1442 B.n407 B.n391 71.676
R1443 B.n403 B.n392 71.676
R1444 B.n583 B.n348 71.676
R1445 B.n108 B.n56 71.676
R1446 B.n112 B.n57 71.676
R1447 B.n116 B.n58 71.676
R1448 B.n120 B.n59 71.676
R1449 B.n124 B.n60 71.676
R1450 B.n128 B.n61 71.676
R1451 B.n132 B.n62 71.676
R1452 B.n136 B.n63 71.676
R1453 B.n140 B.n64 71.676
R1454 B.n144 B.n65 71.676
R1455 B.n148 B.n66 71.676
R1456 B.n152 B.n67 71.676
R1457 B.n156 B.n68 71.676
R1458 B.n160 B.n69 71.676
R1459 B.n164 B.n70 71.676
R1460 B.n168 B.n71 71.676
R1461 B.n172 B.n72 71.676
R1462 B.n176 B.n73 71.676
R1463 B.n180 B.n74 71.676
R1464 B.n184 B.n75 71.676
R1465 B.n188 B.n76 71.676
R1466 B.n192 B.n77 71.676
R1467 B.n196 B.n78 71.676
R1468 B.n200 B.n79 71.676
R1469 B.n204 B.n80 71.676
R1470 B.n208 B.n81 71.676
R1471 B.n213 B.n82 71.676
R1472 B.n217 B.n83 71.676
R1473 B.n221 B.n84 71.676
R1474 B.n225 B.n85 71.676
R1475 B.n229 B.n86 71.676
R1476 B.n233 B.n87 71.676
R1477 B.n237 B.n88 71.676
R1478 B.n241 B.n89 71.676
R1479 B.n245 B.n90 71.676
R1480 B.n249 B.n91 71.676
R1481 B.n253 B.n92 71.676
R1482 B.n257 B.n93 71.676
R1483 B.n261 B.n94 71.676
R1484 B.n265 B.n95 71.676
R1485 B.n269 B.n96 71.676
R1486 B.n273 B.n97 71.676
R1487 B.n277 B.n98 71.676
R1488 B.n281 B.n99 71.676
R1489 B.n285 B.n100 71.676
R1490 B.n289 B.n101 71.676
R1491 B.n102 B.n101 71.676
R1492 B.n288 B.n100 71.676
R1493 B.n284 B.n99 71.676
R1494 B.n280 B.n98 71.676
R1495 B.n276 B.n97 71.676
R1496 B.n272 B.n96 71.676
R1497 B.n268 B.n95 71.676
R1498 B.n264 B.n94 71.676
R1499 B.n260 B.n93 71.676
R1500 B.n256 B.n92 71.676
R1501 B.n252 B.n91 71.676
R1502 B.n248 B.n90 71.676
R1503 B.n244 B.n89 71.676
R1504 B.n240 B.n88 71.676
R1505 B.n236 B.n87 71.676
R1506 B.n232 B.n86 71.676
R1507 B.n228 B.n85 71.676
R1508 B.n224 B.n84 71.676
R1509 B.n220 B.n83 71.676
R1510 B.n216 B.n82 71.676
R1511 B.n212 B.n81 71.676
R1512 B.n207 B.n80 71.676
R1513 B.n203 B.n79 71.676
R1514 B.n199 B.n78 71.676
R1515 B.n195 B.n77 71.676
R1516 B.n191 B.n76 71.676
R1517 B.n187 B.n75 71.676
R1518 B.n183 B.n74 71.676
R1519 B.n179 B.n73 71.676
R1520 B.n175 B.n72 71.676
R1521 B.n171 B.n71 71.676
R1522 B.n167 B.n70 71.676
R1523 B.n163 B.n69 71.676
R1524 B.n159 B.n68 71.676
R1525 B.n155 B.n67 71.676
R1526 B.n151 B.n66 71.676
R1527 B.n147 B.n65 71.676
R1528 B.n143 B.n64 71.676
R1529 B.n139 B.n63 71.676
R1530 B.n135 B.n62 71.676
R1531 B.n131 B.n61 71.676
R1532 B.n127 B.n60 71.676
R1533 B.n123 B.n59 71.676
R1534 B.n119 B.n58 71.676
R1535 B.n115 B.n57 71.676
R1536 B.n111 B.n56 71.676
R1537 B.n581 B.n394 71.676
R1538 B.n573 B.n349 71.676
R1539 B.n569 B.n350 71.676
R1540 B.n565 B.n351 71.676
R1541 B.n561 B.n352 71.676
R1542 B.n557 B.n353 71.676
R1543 B.n553 B.n354 71.676
R1544 B.n549 B.n355 71.676
R1545 B.n545 B.n356 71.676
R1546 B.n541 B.n357 71.676
R1547 B.n537 B.n358 71.676
R1548 B.n533 B.n359 71.676
R1549 B.n529 B.n360 71.676
R1550 B.n525 B.n361 71.676
R1551 B.n521 B.n362 71.676
R1552 B.n517 B.n363 71.676
R1553 B.n513 B.n364 71.676
R1554 B.n509 B.n365 71.676
R1555 B.n505 B.n366 71.676
R1556 B.n501 B.n367 71.676
R1557 B.n496 B.n368 71.676
R1558 B.n492 B.n369 71.676
R1559 B.n488 B.n370 71.676
R1560 B.n484 B.n371 71.676
R1561 B.n480 B.n372 71.676
R1562 B.n476 B.n373 71.676
R1563 B.n472 B.n374 71.676
R1564 B.n468 B.n375 71.676
R1565 B.n464 B.n376 71.676
R1566 B.n460 B.n377 71.676
R1567 B.n456 B.n378 71.676
R1568 B.n452 B.n379 71.676
R1569 B.n448 B.n380 71.676
R1570 B.n444 B.n381 71.676
R1571 B.n440 B.n382 71.676
R1572 B.n436 B.n383 71.676
R1573 B.n432 B.n384 71.676
R1574 B.n428 B.n385 71.676
R1575 B.n424 B.n386 71.676
R1576 B.n420 B.n387 71.676
R1577 B.n416 B.n388 71.676
R1578 B.n412 B.n389 71.676
R1579 B.n408 B.n390 71.676
R1580 B.n404 B.n391 71.676
R1581 B.n400 B.n392 71.676
R1582 B.n584 B.n583 71.676
R1583 B.n399 B.n398 59.5399
R1584 B.n498 B.n396 59.5399
R1585 B.n107 B.n106 59.5399
R1586 B.n210 B.n104 59.5399
R1587 B.n589 B.n345 43.1005
R1588 B.n589 B.n341 43.1005
R1589 B.n595 B.n341 43.1005
R1590 B.n595 B.n337 43.1005
R1591 B.n601 B.n337 43.1005
R1592 B.n607 B.n333 43.1005
R1593 B.n607 B.n329 43.1005
R1594 B.n613 B.n329 43.1005
R1595 B.n613 B.n325 43.1005
R1596 B.n619 B.n325 43.1005
R1597 B.n619 B.n321 43.1005
R1598 B.n626 B.n321 43.1005
R1599 B.n626 B.n625 43.1005
R1600 B.n632 B.n314 43.1005
R1601 B.n638 B.n314 43.1005
R1602 B.n638 B.n310 43.1005
R1603 B.n644 B.n310 43.1005
R1604 B.n650 B.n306 43.1005
R1605 B.n650 B.n301 43.1005
R1606 B.n656 B.n301 43.1005
R1607 B.n656 B.n302 43.1005
R1608 B.n663 B.n294 43.1005
R1609 B.n669 B.n294 43.1005
R1610 B.n669 B.n4 43.1005
R1611 B.n770 B.n4 43.1005
R1612 B.n770 B.n769 43.1005
R1613 B.n769 B.n768 43.1005
R1614 B.n768 B.n8 43.1005
R1615 B.n762 B.n8 43.1005
R1616 B.n761 B.n760 43.1005
R1617 B.n760 B.n15 43.1005
R1618 B.n754 B.n15 43.1005
R1619 B.n754 B.n753 43.1005
R1620 B.n752 B.n22 43.1005
R1621 B.n746 B.n22 43.1005
R1622 B.n746 B.n745 43.1005
R1623 B.n745 B.n744 43.1005
R1624 B.n738 B.n32 43.1005
R1625 B.n738 B.n737 43.1005
R1626 B.n737 B.n736 43.1005
R1627 B.n736 B.n36 43.1005
R1628 B.n730 B.n36 43.1005
R1629 B.n730 B.n729 43.1005
R1630 B.n729 B.n728 43.1005
R1631 B.n728 B.n43 43.1005
R1632 B.n722 B.n721 43.1005
R1633 B.n721 B.n720 43.1005
R1634 B.n720 B.n50 43.1005
R1635 B.n714 B.n50 43.1005
R1636 B.n714 B.n713 43.1005
R1637 B.n109 B.n52 35.7468
R1638 B.n710 B.n709 35.7468
R1639 B.n586 B.n585 35.7468
R1640 B.n579 B.n343 35.7468
R1641 B.n398 B.n397 34.7157
R1642 B.n396 B.n395 34.7157
R1643 B.n106 B.n105 34.7157
R1644 B.n104 B.n103 34.7157
R1645 B.n601 B.t7 32.9593
R1646 B.n632 B.t1 32.9593
R1647 B.n302 B.t3 32.9593
R1648 B.t5 B.n761 32.9593
R1649 B.n744 B.t4 32.9593
R1650 B.n722 B.t11 32.9593
R1651 B.n644 B.t2 21.5505
R1652 B.t2 B.n306 21.5505
R1653 B.n753 B.t0 21.5505
R1654 B.t0 B.n752 21.5505
R1655 B B.n772 18.0485
R1656 B.n110 B.n109 10.6151
R1657 B.n113 B.n110 10.6151
R1658 B.n114 B.n113 10.6151
R1659 B.n117 B.n114 10.6151
R1660 B.n118 B.n117 10.6151
R1661 B.n121 B.n118 10.6151
R1662 B.n122 B.n121 10.6151
R1663 B.n125 B.n122 10.6151
R1664 B.n126 B.n125 10.6151
R1665 B.n129 B.n126 10.6151
R1666 B.n130 B.n129 10.6151
R1667 B.n133 B.n130 10.6151
R1668 B.n134 B.n133 10.6151
R1669 B.n137 B.n134 10.6151
R1670 B.n138 B.n137 10.6151
R1671 B.n141 B.n138 10.6151
R1672 B.n142 B.n141 10.6151
R1673 B.n145 B.n142 10.6151
R1674 B.n146 B.n145 10.6151
R1675 B.n149 B.n146 10.6151
R1676 B.n150 B.n149 10.6151
R1677 B.n153 B.n150 10.6151
R1678 B.n154 B.n153 10.6151
R1679 B.n157 B.n154 10.6151
R1680 B.n158 B.n157 10.6151
R1681 B.n161 B.n158 10.6151
R1682 B.n162 B.n161 10.6151
R1683 B.n165 B.n162 10.6151
R1684 B.n166 B.n165 10.6151
R1685 B.n169 B.n166 10.6151
R1686 B.n170 B.n169 10.6151
R1687 B.n173 B.n170 10.6151
R1688 B.n174 B.n173 10.6151
R1689 B.n177 B.n174 10.6151
R1690 B.n178 B.n177 10.6151
R1691 B.n181 B.n178 10.6151
R1692 B.n182 B.n181 10.6151
R1693 B.n185 B.n182 10.6151
R1694 B.n186 B.n185 10.6151
R1695 B.n189 B.n186 10.6151
R1696 B.n190 B.n189 10.6151
R1697 B.n194 B.n193 10.6151
R1698 B.n197 B.n194 10.6151
R1699 B.n198 B.n197 10.6151
R1700 B.n201 B.n198 10.6151
R1701 B.n202 B.n201 10.6151
R1702 B.n205 B.n202 10.6151
R1703 B.n206 B.n205 10.6151
R1704 B.n209 B.n206 10.6151
R1705 B.n214 B.n211 10.6151
R1706 B.n215 B.n214 10.6151
R1707 B.n218 B.n215 10.6151
R1708 B.n219 B.n218 10.6151
R1709 B.n222 B.n219 10.6151
R1710 B.n223 B.n222 10.6151
R1711 B.n226 B.n223 10.6151
R1712 B.n227 B.n226 10.6151
R1713 B.n230 B.n227 10.6151
R1714 B.n231 B.n230 10.6151
R1715 B.n234 B.n231 10.6151
R1716 B.n235 B.n234 10.6151
R1717 B.n238 B.n235 10.6151
R1718 B.n239 B.n238 10.6151
R1719 B.n242 B.n239 10.6151
R1720 B.n243 B.n242 10.6151
R1721 B.n246 B.n243 10.6151
R1722 B.n247 B.n246 10.6151
R1723 B.n250 B.n247 10.6151
R1724 B.n251 B.n250 10.6151
R1725 B.n254 B.n251 10.6151
R1726 B.n255 B.n254 10.6151
R1727 B.n258 B.n255 10.6151
R1728 B.n259 B.n258 10.6151
R1729 B.n262 B.n259 10.6151
R1730 B.n263 B.n262 10.6151
R1731 B.n266 B.n263 10.6151
R1732 B.n267 B.n266 10.6151
R1733 B.n270 B.n267 10.6151
R1734 B.n271 B.n270 10.6151
R1735 B.n274 B.n271 10.6151
R1736 B.n275 B.n274 10.6151
R1737 B.n278 B.n275 10.6151
R1738 B.n279 B.n278 10.6151
R1739 B.n282 B.n279 10.6151
R1740 B.n283 B.n282 10.6151
R1741 B.n286 B.n283 10.6151
R1742 B.n287 B.n286 10.6151
R1743 B.n290 B.n287 10.6151
R1744 B.n291 B.n290 10.6151
R1745 B.n710 B.n291 10.6151
R1746 B.n587 B.n586 10.6151
R1747 B.n587 B.n339 10.6151
R1748 B.n597 B.n339 10.6151
R1749 B.n598 B.n597 10.6151
R1750 B.n599 B.n598 10.6151
R1751 B.n599 B.n331 10.6151
R1752 B.n609 B.n331 10.6151
R1753 B.n610 B.n609 10.6151
R1754 B.n611 B.n610 10.6151
R1755 B.n611 B.n323 10.6151
R1756 B.n621 B.n323 10.6151
R1757 B.n622 B.n621 10.6151
R1758 B.n623 B.n622 10.6151
R1759 B.n623 B.n316 10.6151
R1760 B.n634 B.n316 10.6151
R1761 B.n635 B.n634 10.6151
R1762 B.n636 B.n635 10.6151
R1763 B.n636 B.n308 10.6151
R1764 B.n646 B.n308 10.6151
R1765 B.n647 B.n646 10.6151
R1766 B.n648 B.n647 10.6151
R1767 B.n648 B.n299 10.6151
R1768 B.n658 B.n299 10.6151
R1769 B.n659 B.n658 10.6151
R1770 B.n661 B.n659 10.6151
R1771 B.n661 B.n660 10.6151
R1772 B.n660 B.n292 10.6151
R1773 B.n672 B.n292 10.6151
R1774 B.n673 B.n672 10.6151
R1775 B.n674 B.n673 10.6151
R1776 B.n675 B.n674 10.6151
R1777 B.n677 B.n675 10.6151
R1778 B.n678 B.n677 10.6151
R1779 B.n679 B.n678 10.6151
R1780 B.n680 B.n679 10.6151
R1781 B.n682 B.n680 10.6151
R1782 B.n683 B.n682 10.6151
R1783 B.n684 B.n683 10.6151
R1784 B.n685 B.n684 10.6151
R1785 B.n687 B.n685 10.6151
R1786 B.n688 B.n687 10.6151
R1787 B.n689 B.n688 10.6151
R1788 B.n690 B.n689 10.6151
R1789 B.n692 B.n690 10.6151
R1790 B.n693 B.n692 10.6151
R1791 B.n694 B.n693 10.6151
R1792 B.n695 B.n694 10.6151
R1793 B.n697 B.n695 10.6151
R1794 B.n698 B.n697 10.6151
R1795 B.n699 B.n698 10.6151
R1796 B.n700 B.n699 10.6151
R1797 B.n702 B.n700 10.6151
R1798 B.n703 B.n702 10.6151
R1799 B.n704 B.n703 10.6151
R1800 B.n705 B.n704 10.6151
R1801 B.n707 B.n705 10.6151
R1802 B.n708 B.n707 10.6151
R1803 B.n709 B.n708 10.6151
R1804 B.n579 B.n578 10.6151
R1805 B.n578 B.n577 10.6151
R1806 B.n577 B.n576 10.6151
R1807 B.n576 B.n574 10.6151
R1808 B.n574 B.n571 10.6151
R1809 B.n571 B.n570 10.6151
R1810 B.n570 B.n567 10.6151
R1811 B.n567 B.n566 10.6151
R1812 B.n566 B.n563 10.6151
R1813 B.n563 B.n562 10.6151
R1814 B.n562 B.n559 10.6151
R1815 B.n559 B.n558 10.6151
R1816 B.n558 B.n555 10.6151
R1817 B.n555 B.n554 10.6151
R1818 B.n554 B.n551 10.6151
R1819 B.n551 B.n550 10.6151
R1820 B.n550 B.n547 10.6151
R1821 B.n547 B.n546 10.6151
R1822 B.n546 B.n543 10.6151
R1823 B.n543 B.n542 10.6151
R1824 B.n542 B.n539 10.6151
R1825 B.n539 B.n538 10.6151
R1826 B.n538 B.n535 10.6151
R1827 B.n535 B.n534 10.6151
R1828 B.n534 B.n531 10.6151
R1829 B.n531 B.n530 10.6151
R1830 B.n530 B.n527 10.6151
R1831 B.n527 B.n526 10.6151
R1832 B.n526 B.n523 10.6151
R1833 B.n523 B.n522 10.6151
R1834 B.n522 B.n519 10.6151
R1835 B.n519 B.n518 10.6151
R1836 B.n518 B.n515 10.6151
R1837 B.n515 B.n514 10.6151
R1838 B.n514 B.n511 10.6151
R1839 B.n511 B.n510 10.6151
R1840 B.n510 B.n507 10.6151
R1841 B.n507 B.n506 10.6151
R1842 B.n506 B.n503 10.6151
R1843 B.n503 B.n502 10.6151
R1844 B.n502 B.n499 10.6151
R1845 B.n497 B.n494 10.6151
R1846 B.n494 B.n493 10.6151
R1847 B.n493 B.n490 10.6151
R1848 B.n490 B.n489 10.6151
R1849 B.n489 B.n486 10.6151
R1850 B.n486 B.n485 10.6151
R1851 B.n485 B.n482 10.6151
R1852 B.n482 B.n481 10.6151
R1853 B.n478 B.n477 10.6151
R1854 B.n477 B.n474 10.6151
R1855 B.n474 B.n473 10.6151
R1856 B.n473 B.n470 10.6151
R1857 B.n470 B.n469 10.6151
R1858 B.n469 B.n466 10.6151
R1859 B.n466 B.n465 10.6151
R1860 B.n465 B.n462 10.6151
R1861 B.n462 B.n461 10.6151
R1862 B.n461 B.n458 10.6151
R1863 B.n458 B.n457 10.6151
R1864 B.n457 B.n454 10.6151
R1865 B.n454 B.n453 10.6151
R1866 B.n453 B.n450 10.6151
R1867 B.n450 B.n449 10.6151
R1868 B.n449 B.n446 10.6151
R1869 B.n446 B.n445 10.6151
R1870 B.n445 B.n442 10.6151
R1871 B.n442 B.n441 10.6151
R1872 B.n441 B.n438 10.6151
R1873 B.n438 B.n437 10.6151
R1874 B.n437 B.n434 10.6151
R1875 B.n434 B.n433 10.6151
R1876 B.n433 B.n430 10.6151
R1877 B.n430 B.n429 10.6151
R1878 B.n429 B.n426 10.6151
R1879 B.n426 B.n425 10.6151
R1880 B.n425 B.n422 10.6151
R1881 B.n422 B.n421 10.6151
R1882 B.n421 B.n418 10.6151
R1883 B.n418 B.n417 10.6151
R1884 B.n417 B.n414 10.6151
R1885 B.n414 B.n413 10.6151
R1886 B.n413 B.n410 10.6151
R1887 B.n410 B.n409 10.6151
R1888 B.n409 B.n406 10.6151
R1889 B.n406 B.n405 10.6151
R1890 B.n405 B.n402 10.6151
R1891 B.n402 B.n401 10.6151
R1892 B.n401 B.n347 10.6151
R1893 B.n585 B.n347 10.6151
R1894 B.n591 B.n343 10.6151
R1895 B.n592 B.n591 10.6151
R1896 B.n593 B.n592 10.6151
R1897 B.n593 B.n335 10.6151
R1898 B.n603 B.n335 10.6151
R1899 B.n604 B.n603 10.6151
R1900 B.n605 B.n604 10.6151
R1901 B.n605 B.n327 10.6151
R1902 B.n615 B.n327 10.6151
R1903 B.n616 B.n615 10.6151
R1904 B.n617 B.n616 10.6151
R1905 B.n617 B.n319 10.6151
R1906 B.n628 B.n319 10.6151
R1907 B.n629 B.n628 10.6151
R1908 B.n630 B.n629 10.6151
R1909 B.n630 B.n312 10.6151
R1910 B.n640 B.n312 10.6151
R1911 B.n641 B.n640 10.6151
R1912 B.n642 B.n641 10.6151
R1913 B.n642 B.n304 10.6151
R1914 B.n652 B.n304 10.6151
R1915 B.n653 B.n652 10.6151
R1916 B.n654 B.n653 10.6151
R1917 B.n654 B.n296 10.6151
R1918 B.n665 B.n296 10.6151
R1919 B.n666 B.n665 10.6151
R1920 B.n667 B.n666 10.6151
R1921 B.n667 B.n0 10.6151
R1922 B.n766 B.n1 10.6151
R1923 B.n766 B.n765 10.6151
R1924 B.n765 B.n764 10.6151
R1925 B.n764 B.n10 10.6151
R1926 B.n758 B.n10 10.6151
R1927 B.n758 B.n757 10.6151
R1928 B.n757 B.n756 10.6151
R1929 B.n756 B.n17 10.6151
R1930 B.n750 B.n17 10.6151
R1931 B.n750 B.n749 10.6151
R1932 B.n749 B.n748 10.6151
R1933 B.n748 B.n24 10.6151
R1934 B.n742 B.n24 10.6151
R1935 B.n742 B.n741 10.6151
R1936 B.n741 B.n740 10.6151
R1937 B.n740 B.n30 10.6151
R1938 B.n734 B.n30 10.6151
R1939 B.n734 B.n733 10.6151
R1940 B.n733 B.n732 10.6151
R1941 B.n732 B.n38 10.6151
R1942 B.n726 B.n38 10.6151
R1943 B.n726 B.n725 10.6151
R1944 B.n725 B.n724 10.6151
R1945 B.n724 B.n45 10.6151
R1946 B.n718 B.n45 10.6151
R1947 B.n718 B.n717 10.6151
R1948 B.n717 B.n716 10.6151
R1949 B.n716 B.n52 10.6151
R1950 B.t7 B.n333 10.1417
R1951 B.n625 B.t1 10.1417
R1952 B.n663 B.t3 10.1417
R1953 B.n762 B.t5 10.1417
R1954 B.n32 B.t4 10.1417
R1955 B.t11 B.n43 10.1417
R1956 B.n193 B.n107 6.5566
R1957 B.n210 B.n209 6.5566
R1958 B.n498 B.n497 6.5566
R1959 B.n481 B.n399 6.5566
R1960 B.n190 B.n107 4.05904
R1961 B.n211 B.n210 4.05904
R1962 B.n499 B.n498 4.05904
R1963 B.n478 B.n399 4.05904
R1964 B.n772 B.n0 2.81026
R1965 B.n772 B.n1 2.81026
R1966 VP.n7 VP.t0 236.121
R1967 VP.n20 VP.t3 199.404
R1968 VP.n14 VP.t5 199.404
R1969 VP.n26 VP.t2 199.404
R1970 VP.n6 VP.t1 199.404
R1971 VP.n12 VP.t4 199.404
R1972 VP.n15 VP.n14 171.63
R1973 VP.n27 VP.n26 171.63
R1974 VP.n13 VP.n12 171.63
R1975 VP.n8 VP.n5 161.3
R1976 VP.n10 VP.n9 161.3
R1977 VP.n11 VP.n4 161.3
R1978 VP.n25 VP.n0 161.3
R1979 VP.n24 VP.n23 161.3
R1980 VP.n22 VP.n1 161.3
R1981 VP.n21 VP.n20 161.3
R1982 VP.n19 VP.n2 161.3
R1983 VP.n18 VP.n17 161.3
R1984 VP.n16 VP.n3 161.3
R1985 VP.n19 VP.n18 50.7491
R1986 VP.n24 VP.n1 50.7491
R1987 VP.n10 VP.n5 50.7491
R1988 VP.n15 VP.n13 44.2467
R1989 VP.n7 VP.n6 41.9508
R1990 VP.n18 VP.n3 30.405
R1991 VP.n25 VP.n24 30.405
R1992 VP.n11 VP.n10 30.405
R1993 VP.n20 VP.n19 24.5923
R1994 VP.n20 VP.n1 24.5923
R1995 VP.n6 VP.n5 24.5923
R1996 VP.n8 VP.n7 17.3014
R1997 VP.n14 VP.n3 14.2638
R1998 VP.n26 VP.n25 14.2638
R1999 VP.n12 VP.n11 14.2638
R2000 VP.n9 VP.n8 0.189894
R2001 VP.n9 VP.n4 0.189894
R2002 VP.n13 VP.n4 0.189894
R2003 VP.n16 VP.n15 0.189894
R2004 VP.n17 VP.n16 0.189894
R2005 VP.n17 VP.n2 0.189894
R2006 VP.n21 VP.n2 0.189894
R2007 VP.n22 VP.n21 0.189894
R2008 VP.n23 VP.n22 0.189894
R2009 VP.n23 VP.n0 0.189894
R2010 VP.n27 VP.n0 0.189894
R2011 VP VP.n27 0.0516364
R2012 VDD1.n60 VDD1.n0 289.615
R2013 VDD1.n125 VDD1.n65 289.615
R2014 VDD1.n61 VDD1.n60 185
R2015 VDD1.n59 VDD1.n58 185
R2016 VDD1.n4 VDD1.n3 185
R2017 VDD1.n53 VDD1.n52 185
R2018 VDD1.n51 VDD1.n50 185
R2019 VDD1.n8 VDD1.n7 185
R2020 VDD1.n45 VDD1.n44 185
R2021 VDD1.n43 VDD1.n10 185
R2022 VDD1.n42 VDD1.n41 185
R2023 VDD1.n13 VDD1.n11 185
R2024 VDD1.n36 VDD1.n35 185
R2025 VDD1.n34 VDD1.n33 185
R2026 VDD1.n17 VDD1.n16 185
R2027 VDD1.n28 VDD1.n27 185
R2028 VDD1.n26 VDD1.n25 185
R2029 VDD1.n21 VDD1.n20 185
R2030 VDD1.n85 VDD1.n84 185
R2031 VDD1.n90 VDD1.n89 185
R2032 VDD1.n92 VDD1.n91 185
R2033 VDD1.n81 VDD1.n80 185
R2034 VDD1.n98 VDD1.n97 185
R2035 VDD1.n100 VDD1.n99 185
R2036 VDD1.n77 VDD1.n76 185
R2037 VDD1.n107 VDD1.n106 185
R2038 VDD1.n108 VDD1.n75 185
R2039 VDD1.n110 VDD1.n109 185
R2040 VDD1.n73 VDD1.n72 185
R2041 VDD1.n116 VDD1.n115 185
R2042 VDD1.n118 VDD1.n117 185
R2043 VDD1.n69 VDD1.n68 185
R2044 VDD1.n124 VDD1.n123 185
R2045 VDD1.n126 VDD1.n125 185
R2046 VDD1.n22 VDD1.t5 149.524
R2047 VDD1.n86 VDD1.t0 149.524
R2048 VDD1.n60 VDD1.n59 104.615
R2049 VDD1.n59 VDD1.n3 104.615
R2050 VDD1.n52 VDD1.n3 104.615
R2051 VDD1.n52 VDD1.n51 104.615
R2052 VDD1.n51 VDD1.n7 104.615
R2053 VDD1.n44 VDD1.n7 104.615
R2054 VDD1.n44 VDD1.n43 104.615
R2055 VDD1.n43 VDD1.n42 104.615
R2056 VDD1.n42 VDD1.n11 104.615
R2057 VDD1.n35 VDD1.n11 104.615
R2058 VDD1.n35 VDD1.n34 104.615
R2059 VDD1.n34 VDD1.n16 104.615
R2060 VDD1.n27 VDD1.n16 104.615
R2061 VDD1.n27 VDD1.n26 104.615
R2062 VDD1.n26 VDD1.n20 104.615
R2063 VDD1.n90 VDD1.n84 104.615
R2064 VDD1.n91 VDD1.n90 104.615
R2065 VDD1.n91 VDD1.n80 104.615
R2066 VDD1.n98 VDD1.n80 104.615
R2067 VDD1.n99 VDD1.n98 104.615
R2068 VDD1.n99 VDD1.n76 104.615
R2069 VDD1.n107 VDD1.n76 104.615
R2070 VDD1.n108 VDD1.n107 104.615
R2071 VDD1.n109 VDD1.n108 104.615
R2072 VDD1.n109 VDD1.n72 104.615
R2073 VDD1.n116 VDD1.n72 104.615
R2074 VDD1.n117 VDD1.n116 104.615
R2075 VDD1.n117 VDD1.n68 104.615
R2076 VDD1.n124 VDD1.n68 104.615
R2077 VDD1.n125 VDD1.n124 104.615
R2078 VDD1.n131 VDD1.n130 61.4344
R2079 VDD1.n133 VDD1.n132 61.104
R2080 VDD1.t5 VDD1.n20 52.3082
R2081 VDD1.t0 VDD1.n84 52.3082
R2082 VDD1 VDD1.n64 49.3039
R2083 VDD1.n131 VDD1.n129 49.1904
R2084 VDD1.n133 VDD1.n131 40.4987
R2085 VDD1.n45 VDD1.n10 13.1884
R2086 VDD1.n110 VDD1.n75 13.1884
R2087 VDD1.n46 VDD1.n8 12.8005
R2088 VDD1.n41 VDD1.n12 12.8005
R2089 VDD1.n106 VDD1.n105 12.8005
R2090 VDD1.n111 VDD1.n73 12.8005
R2091 VDD1.n50 VDD1.n49 12.0247
R2092 VDD1.n40 VDD1.n13 12.0247
R2093 VDD1.n104 VDD1.n77 12.0247
R2094 VDD1.n115 VDD1.n114 12.0247
R2095 VDD1.n53 VDD1.n6 11.249
R2096 VDD1.n37 VDD1.n36 11.249
R2097 VDD1.n101 VDD1.n100 11.249
R2098 VDD1.n118 VDD1.n71 11.249
R2099 VDD1.n54 VDD1.n4 10.4732
R2100 VDD1.n33 VDD1.n15 10.4732
R2101 VDD1.n97 VDD1.n79 10.4732
R2102 VDD1.n119 VDD1.n69 10.4732
R2103 VDD1.n22 VDD1.n21 10.2747
R2104 VDD1.n86 VDD1.n85 10.2747
R2105 VDD1.n58 VDD1.n57 9.69747
R2106 VDD1.n32 VDD1.n17 9.69747
R2107 VDD1.n96 VDD1.n81 9.69747
R2108 VDD1.n123 VDD1.n122 9.69747
R2109 VDD1.n64 VDD1.n63 9.45567
R2110 VDD1.n129 VDD1.n128 9.45567
R2111 VDD1.n24 VDD1.n23 9.3005
R2112 VDD1.n19 VDD1.n18 9.3005
R2113 VDD1.n30 VDD1.n29 9.3005
R2114 VDD1.n32 VDD1.n31 9.3005
R2115 VDD1.n15 VDD1.n14 9.3005
R2116 VDD1.n38 VDD1.n37 9.3005
R2117 VDD1.n40 VDD1.n39 9.3005
R2118 VDD1.n12 VDD1.n9 9.3005
R2119 VDD1.n63 VDD1.n62 9.3005
R2120 VDD1.n2 VDD1.n1 9.3005
R2121 VDD1.n57 VDD1.n56 9.3005
R2122 VDD1.n55 VDD1.n54 9.3005
R2123 VDD1.n6 VDD1.n5 9.3005
R2124 VDD1.n49 VDD1.n48 9.3005
R2125 VDD1.n47 VDD1.n46 9.3005
R2126 VDD1.n128 VDD1.n127 9.3005
R2127 VDD1.n67 VDD1.n66 9.3005
R2128 VDD1.n122 VDD1.n121 9.3005
R2129 VDD1.n120 VDD1.n119 9.3005
R2130 VDD1.n71 VDD1.n70 9.3005
R2131 VDD1.n114 VDD1.n113 9.3005
R2132 VDD1.n112 VDD1.n111 9.3005
R2133 VDD1.n88 VDD1.n87 9.3005
R2134 VDD1.n83 VDD1.n82 9.3005
R2135 VDD1.n94 VDD1.n93 9.3005
R2136 VDD1.n96 VDD1.n95 9.3005
R2137 VDD1.n79 VDD1.n78 9.3005
R2138 VDD1.n102 VDD1.n101 9.3005
R2139 VDD1.n104 VDD1.n103 9.3005
R2140 VDD1.n105 VDD1.n74 9.3005
R2141 VDD1.n61 VDD1.n2 8.92171
R2142 VDD1.n29 VDD1.n28 8.92171
R2143 VDD1.n93 VDD1.n92 8.92171
R2144 VDD1.n126 VDD1.n67 8.92171
R2145 VDD1.n62 VDD1.n0 8.14595
R2146 VDD1.n25 VDD1.n19 8.14595
R2147 VDD1.n89 VDD1.n83 8.14595
R2148 VDD1.n127 VDD1.n65 8.14595
R2149 VDD1.n24 VDD1.n21 7.3702
R2150 VDD1.n88 VDD1.n85 7.3702
R2151 VDD1.n64 VDD1.n0 5.81868
R2152 VDD1.n25 VDD1.n24 5.81868
R2153 VDD1.n89 VDD1.n88 5.81868
R2154 VDD1.n129 VDD1.n65 5.81868
R2155 VDD1.n62 VDD1.n61 5.04292
R2156 VDD1.n28 VDD1.n19 5.04292
R2157 VDD1.n92 VDD1.n83 5.04292
R2158 VDD1.n127 VDD1.n126 5.04292
R2159 VDD1.n58 VDD1.n2 4.26717
R2160 VDD1.n29 VDD1.n17 4.26717
R2161 VDD1.n93 VDD1.n81 4.26717
R2162 VDD1.n123 VDD1.n67 4.26717
R2163 VDD1.n57 VDD1.n4 3.49141
R2164 VDD1.n33 VDD1.n32 3.49141
R2165 VDD1.n97 VDD1.n96 3.49141
R2166 VDD1.n122 VDD1.n69 3.49141
R2167 VDD1.n23 VDD1.n22 2.84303
R2168 VDD1.n87 VDD1.n86 2.84303
R2169 VDD1.n54 VDD1.n53 2.71565
R2170 VDD1.n36 VDD1.n15 2.71565
R2171 VDD1.n100 VDD1.n79 2.71565
R2172 VDD1.n119 VDD1.n118 2.71565
R2173 VDD1.n50 VDD1.n6 1.93989
R2174 VDD1.n37 VDD1.n13 1.93989
R2175 VDD1.n101 VDD1.n77 1.93989
R2176 VDD1.n115 VDD1.n71 1.93989
R2177 VDD1.n132 VDD1.t4 1.63957
R2178 VDD1.n132 VDD1.t1 1.63957
R2179 VDD1.n130 VDD1.t2 1.63957
R2180 VDD1.n130 VDD1.t3 1.63957
R2181 VDD1.n49 VDD1.n8 1.16414
R2182 VDD1.n41 VDD1.n40 1.16414
R2183 VDD1.n106 VDD1.n104 1.16414
R2184 VDD1.n114 VDD1.n73 1.16414
R2185 VDD1.n46 VDD1.n45 0.388379
R2186 VDD1.n12 VDD1.n10 0.388379
R2187 VDD1.n105 VDD1.n75 0.388379
R2188 VDD1.n111 VDD1.n110 0.388379
R2189 VDD1 VDD1.n133 0.328086
R2190 VDD1.n63 VDD1.n1 0.155672
R2191 VDD1.n56 VDD1.n1 0.155672
R2192 VDD1.n56 VDD1.n55 0.155672
R2193 VDD1.n55 VDD1.n5 0.155672
R2194 VDD1.n48 VDD1.n5 0.155672
R2195 VDD1.n48 VDD1.n47 0.155672
R2196 VDD1.n47 VDD1.n9 0.155672
R2197 VDD1.n39 VDD1.n9 0.155672
R2198 VDD1.n39 VDD1.n38 0.155672
R2199 VDD1.n38 VDD1.n14 0.155672
R2200 VDD1.n31 VDD1.n14 0.155672
R2201 VDD1.n31 VDD1.n30 0.155672
R2202 VDD1.n30 VDD1.n18 0.155672
R2203 VDD1.n23 VDD1.n18 0.155672
R2204 VDD1.n87 VDD1.n82 0.155672
R2205 VDD1.n94 VDD1.n82 0.155672
R2206 VDD1.n95 VDD1.n94 0.155672
R2207 VDD1.n95 VDD1.n78 0.155672
R2208 VDD1.n102 VDD1.n78 0.155672
R2209 VDD1.n103 VDD1.n102 0.155672
R2210 VDD1.n103 VDD1.n74 0.155672
R2211 VDD1.n112 VDD1.n74 0.155672
R2212 VDD1.n113 VDD1.n112 0.155672
R2213 VDD1.n113 VDD1.n70 0.155672
R2214 VDD1.n120 VDD1.n70 0.155672
R2215 VDD1.n121 VDD1.n120 0.155672
R2216 VDD1.n121 VDD1.n66 0.155672
R2217 VDD1.n128 VDD1.n66 0.155672
C0 VDD2 VP 0.362095f
C1 VDD1 VTAIL 8.06873f
C2 VN VTAIL 5.75766f
C3 VN VDD1 0.149465f
C4 VDD2 VTAIL 8.110129f
C5 VDD2 VDD1 0.99175f
C6 VN VDD2 5.86579f
C7 VTAIL VP 5.77209f
C8 VDD1 VP 6.07467f
C9 VN VP 5.82758f
C10 VDD2 B 5.099365f
C11 VDD1 B 5.163798f
C12 VTAIL B 7.035699f
C13 VN B 9.67434f
C14 VP B 8.053638f
C15 VDD1.n0 B 0.030323f
C16 VDD1.n1 B 0.021995f
C17 VDD1.n2 B 0.011819f
C18 VDD1.n3 B 0.027936f
C19 VDD1.n4 B 0.012514f
C20 VDD1.n5 B 0.021995f
C21 VDD1.n6 B 0.011819f
C22 VDD1.n7 B 0.027936f
C23 VDD1.n8 B 0.012514f
C24 VDD1.n9 B 0.021995f
C25 VDD1.n10 B 0.012167f
C26 VDD1.n11 B 0.027936f
C27 VDD1.n12 B 0.011819f
C28 VDD1.n13 B 0.012514f
C29 VDD1.n14 B 0.021995f
C30 VDD1.n15 B 0.011819f
C31 VDD1.n16 B 0.027936f
C32 VDD1.n17 B 0.012514f
C33 VDD1.n18 B 0.021995f
C34 VDD1.n19 B 0.011819f
C35 VDD1.n20 B 0.020952f
C36 VDD1.n21 B 0.019749f
C37 VDD1.t5 B 0.047192f
C38 VDD1.n22 B 0.159259f
C39 VDD1.n23 B 1.11745f
C40 VDD1.n24 B 0.011819f
C41 VDD1.n25 B 0.012514f
C42 VDD1.n26 B 0.027936f
C43 VDD1.n27 B 0.027936f
C44 VDD1.n28 B 0.012514f
C45 VDD1.n29 B 0.011819f
C46 VDD1.n30 B 0.021995f
C47 VDD1.n31 B 0.021995f
C48 VDD1.n32 B 0.011819f
C49 VDD1.n33 B 0.012514f
C50 VDD1.n34 B 0.027936f
C51 VDD1.n35 B 0.027936f
C52 VDD1.n36 B 0.012514f
C53 VDD1.n37 B 0.011819f
C54 VDD1.n38 B 0.021995f
C55 VDD1.n39 B 0.021995f
C56 VDD1.n40 B 0.011819f
C57 VDD1.n41 B 0.012514f
C58 VDD1.n42 B 0.027936f
C59 VDD1.n43 B 0.027936f
C60 VDD1.n44 B 0.027936f
C61 VDD1.n45 B 0.012167f
C62 VDD1.n46 B 0.011819f
C63 VDD1.n47 B 0.021995f
C64 VDD1.n48 B 0.021995f
C65 VDD1.n49 B 0.011819f
C66 VDD1.n50 B 0.012514f
C67 VDD1.n51 B 0.027936f
C68 VDD1.n52 B 0.027936f
C69 VDD1.n53 B 0.012514f
C70 VDD1.n54 B 0.011819f
C71 VDD1.n55 B 0.021995f
C72 VDD1.n56 B 0.021995f
C73 VDD1.n57 B 0.011819f
C74 VDD1.n58 B 0.012514f
C75 VDD1.n59 B 0.027936f
C76 VDD1.n60 B 0.059428f
C77 VDD1.n61 B 0.012514f
C78 VDD1.n62 B 0.011819f
C79 VDD1.n63 B 0.049639f
C80 VDD1.n64 B 0.051455f
C81 VDD1.n65 B 0.030323f
C82 VDD1.n66 B 0.021995f
C83 VDD1.n67 B 0.011819f
C84 VDD1.n68 B 0.027936f
C85 VDD1.n69 B 0.012514f
C86 VDD1.n70 B 0.021995f
C87 VDD1.n71 B 0.011819f
C88 VDD1.n72 B 0.027936f
C89 VDD1.n73 B 0.012514f
C90 VDD1.n74 B 0.021995f
C91 VDD1.n75 B 0.012167f
C92 VDD1.n76 B 0.027936f
C93 VDD1.n77 B 0.012514f
C94 VDD1.n78 B 0.021995f
C95 VDD1.n79 B 0.011819f
C96 VDD1.n80 B 0.027936f
C97 VDD1.n81 B 0.012514f
C98 VDD1.n82 B 0.021995f
C99 VDD1.n83 B 0.011819f
C100 VDD1.n84 B 0.020952f
C101 VDD1.n85 B 0.019749f
C102 VDD1.t0 B 0.047192f
C103 VDD1.n86 B 0.159259f
C104 VDD1.n87 B 1.11745f
C105 VDD1.n88 B 0.011819f
C106 VDD1.n89 B 0.012514f
C107 VDD1.n90 B 0.027936f
C108 VDD1.n91 B 0.027936f
C109 VDD1.n92 B 0.012514f
C110 VDD1.n93 B 0.011819f
C111 VDD1.n94 B 0.021995f
C112 VDD1.n95 B 0.021995f
C113 VDD1.n96 B 0.011819f
C114 VDD1.n97 B 0.012514f
C115 VDD1.n98 B 0.027936f
C116 VDD1.n99 B 0.027936f
C117 VDD1.n100 B 0.012514f
C118 VDD1.n101 B 0.011819f
C119 VDD1.n102 B 0.021995f
C120 VDD1.n103 B 0.021995f
C121 VDD1.n104 B 0.011819f
C122 VDD1.n105 B 0.011819f
C123 VDD1.n106 B 0.012514f
C124 VDD1.n107 B 0.027936f
C125 VDD1.n108 B 0.027936f
C126 VDD1.n109 B 0.027936f
C127 VDD1.n110 B 0.012167f
C128 VDD1.n111 B 0.011819f
C129 VDD1.n112 B 0.021995f
C130 VDD1.n113 B 0.021995f
C131 VDD1.n114 B 0.011819f
C132 VDD1.n115 B 0.012514f
C133 VDD1.n116 B 0.027936f
C134 VDD1.n117 B 0.027936f
C135 VDD1.n118 B 0.012514f
C136 VDD1.n119 B 0.011819f
C137 VDD1.n120 B 0.021995f
C138 VDD1.n121 B 0.021995f
C139 VDD1.n122 B 0.011819f
C140 VDD1.n123 B 0.012514f
C141 VDD1.n124 B 0.027936f
C142 VDD1.n125 B 0.059428f
C143 VDD1.n126 B 0.012514f
C144 VDD1.n127 B 0.011819f
C145 VDD1.n128 B 0.049639f
C146 VDD1.n129 B 0.050998f
C147 VDD1.t2 B 0.209966f
C148 VDD1.t3 B 0.209966f
C149 VDD1.n130 B 1.87251f
C150 VDD1.n131 B 2.01068f
C151 VDD1.t4 B 0.209966f
C152 VDD1.t1 B 0.209966f
C153 VDD1.n132 B 1.87076f
C154 VDD1.n133 B 2.179f
C155 VP.n0 B 0.033475f
C156 VP.t2 B 1.60892f
C157 VP.n1 B 0.060813f
C158 VP.n2 B 0.033475f
C159 VP.t3 B 1.60892f
C160 VP.n3 B 0.053658f
C161 VP.n4 B 0.033475f
C162 VP.t4 B 1.60892f
C163 VP.n5 B 0.060813f
C164 VP.t0 B 1.71956f
C165 VP.t1 B 1.60892f
C166 VP.n6 B 0.659598f
C167 VP.n7 B 0.648551f
C168 VP.n8 B 0.212902f
C169 VP.n9 B 0.033475f
C170 VP.n10 B 0.032057f
C171 VP.n11 B 0.053658f
C172 VP.n12 B 0.654912f
C173 VP.n13 B 1.50952f
C174 VP.t5 B 1.60892f
C175 VP.n14 B 0.654912f
C176 VP.n15 B 1.5368f
C177 VP.n16 B 0.033475f
C178 VP.n17 B 0.033475f
C179 VP.n18 B 0.032057f
C180 VP.n19 B 0.060813f
C181 VP.n20 B 0.613601f
C182 VP.n21 B 0.033475f
C183 VP.n22 B 0.033475f
C184 VP.n23 B 0.033475f
C185 VP.n24 B 0.032057f
C186 VP.n25 B 0.053658f
C187 VP.n26 B 0.654912f
C188 VP.n27 B 0.0306f
C189 VTAIL.t9 B 0.222855f
C190 VTAIL.t10 B 0.222855f
C191 VTAIL.n0 B 1.91431f
C192 VTAIL.n1 B 0.360643f
C193 VTAIL.n2 B 0.032184f
C194 VTAIL.n3 B 0.023346f
C195 VTAIL.n4 B 0.012545f
C196 VTAIL.n5 B 0.029651f
C197 VTAIL.n6 B 0.013283f
C198 VTAIL.n7 B 0.023346f
C199 VTAIL.n8 B 0.012545f
C200 VTAIL.n9 B 0.029651f
C201 VTAIL.n10 B 0.013283f
C202 VTAIL.n11 B 0.023346f
C203 VTAIL.n12 B 0.012914f
C204 VTAIL.n13 B 0.029651f
C205 VTAIL.n14 B 0.013283f
C206 VTAIL.n15 B 0.023346f
C207 VTAIL.n16 B 0.012545f
C208 VTAIL.n17 B 0.029651f
C209 VTAIL.n18 B 0.013283f
C210 VTAIL.n19 B 0.023346f
C211 VTAIL.n20 B 0.012545f
C212 VTAIL.n21 B 0.022239f
C213 VTAIL.n22 B 0.020961f
C214 VTAIL.t3 B 0.050089f
C215 VTAIL.n23 B 0.169035f
C216 VTAIL.n24 B 1.18605f
C217 VTAIL.n25 B 0.012545f
C218 VTAIL.n26 B 0.013283f
C219 VTAIL.n27 B 0.029651f
C220 VTAIL.n28 B 0.029651f
C221 VTAIL.n29 B 0.013283f
C222 VTAIL.n30 B 0.012545f
C223 VTAIL.n31 B 0.023346f
C224 VTAIL.n32 B 0.023346f
C225 VTAIL.n33 B 0.012545f
C226 VTAIL.n34 B 0.013283f
C227 VTAIL.n35 B 0.029651f
C228 VTAIL.n36 B 0.029651f
C229 VTAIL.n37 B 0.013283f
C230 VTAIL.n38 B 0.012545f
C231 VTAIL.n39 B 0.023346f
C232 VTAIL.n40 B 0.023346f
C233 VTAIL.n41 B 0.012545f
C234 VTAIL.n42 B 0.012545f
C235 VTAIL.n43 B 0.013283f
C236 VTAIL.n44 B 0.029651f
C237 VTAIL.n45 B 0.029651f
C238 VTAIL.n46 B 0.029651f
C239 VTAIL.n47 B 0.012914f
C240 VTAIL.n48 B 0.012545f
C241 VTAIL.n49 B 0.023346f
C242 VTAIL.n50 B 0.023346f
C243 VTAIL.n51 B 0.012545f
C244 VTAIL.n52 B 0.013283f
C245 VTAIL.n53 B 0.029651f
C246 VTAIL.n54 B 0.029651f
C247 VTAIL.n55 B 0.013283f
C248 VTAIL.n56 B 0.012545f
C249 VTAIL.n57 B 0.023346f
C250 VTAIL.n58 B 0.023346f
C251 VTAIL.n59 B 0.012545f
C252 VTAIL.n60 B 0.013283f
C253 VTAIL.n61 B 0.029651f
C254 VTAIL.n62 B 0.063076f
C255 VTAIL.n63 B 0.013283f
C256 VTAIL.n64 B 0.012545f
C257 VTAIL.n65 B 0.052686f
C258 VTAIL.n66 B 0.03514f
C259 VTAIL.n67 B 0.22868f
C260 VTAIL.t1 B 0.222855f
C261 VTAIL.t2 B 0.222855f
C262 VTAIL.n68 B 1.91431f
C263 VTAIL.n69 B 1.68259f
C264 VTAIL.t8 B 0.222855f
C265 VTAIL.t11 B 0.222855f
C266 VTAIL.n70 B 1.91432f
C267 VTAIL.n71 B 1.68258f
C268 VTAIL.n72 B 0.032184f
C269 VTAIL.n73 B 0.023346f
C270 VTAIL.n74 B 0.012545f
C271 VTAIL.n75 B 0.029651f
C272 VTAIL.n76 B 0.013283f
C273 VTAIL.n77 B 0.023346f
C274 VTAIL.n78 B 0.012545f
C275 VTAIL.n79 B 0.029651f
C276 VTAIL.n80 B 0.013283f
C277 VTAIL.n81 B 0.023346f
C278 VTAIL.n82 B 0.012914f
C279 VTAIL.n83 B 0.029651f
C280 VTAIL.n84 B 0.012545f
C281 VTAIL.n85 B 0.013283f
C282 VTAIL.n86 B 0.023346f
C283 VTAIL.n87 B 0.012545f
C284 VTAIL.n88 B 0.029651f
C285 VTAIL.n89 B 0.013283f
C286 VTAIL.n90 B 0.023346f
C287 VTAIL.n91 B 0.012545f
C288 VTAIL.n92 B 0.022239f
C289 VTAIL.n93 B 0.020961f
C290 VTAIL.t6 B 0.050089f
C291 VTAIL.n94 B 0.169035f
C292 VTAIL.n95 B 1.18605f
C293 VTAIL.n96 B 0.012545f
C294 VTAIL.n97 B 0.013283f
C295 VTAIL.n98 B 0.029651f
C296 VTAIL.n99 B 0.029651f
C297 VTAIL.n100 B 0.013283f
C298 VTAIL.n101 B 0.012545f
C299 VTAIL.n102 B 0.023346f
C300 VTAIL.n103 B 0.023346f
C301 VTAIL.n104 B 0.012545f
C302 VTAIL.n105 B 0.013283f
C303 VTAIL.n106 B 0.029651f
C304 VTAIL.n107 B 0.029651f
C305 VTAIL.n108 B 0.013283f
C306 VTAIL.n109 B 0.012545f
C307 VTAIL.n110 B 0.023346f
C308 VTAIL.n111 B 0.023346f
C309 VTAIL.n112 B 0.012545f
C310 VTAIL.n113 B 0.013283f
C311 VTAIL.n114 B 0.029651f
C312 VTAIL.n115 B 0.029651f
C313 VTAIL.n116 B 0.029651f
C314 VTAIL.n117 B 0.012914f
C315 VTAIL.n118 B 0.012545f
C316 VTAIL.n119 B 0.023346f
C317 VTAIL.n120 B 0.023346f
C318 VTAIL.n121 B 0.012545f
C319 VTAIL.n122 B 0.013283f
C320 VTAIL.n123 B 0.029651f
C321 VTAIL.n124 B 0.029651f
C322 VTAIL.n125 B 0.013283f
C323 VTAIL.n126 B 0.012545f
C324 VTAIL.n127 B 0.023346f
C325 VTAIL.n128 B 0.023346f
C326 VTAIL.n129 B 0.012545f
C327 VTAIL.n130 B 0.013283f
C328 VTAIL.n131 B 0.029651f
C329 VTAIL.n132 B 0.063076f
C330 VTAIL.n133 B 0.013283f
C331 VTAIL.n134 B 0.012545f
C332 VTAIL.n135 B 0.052686f
C333 VTAIL.n136 B 0.03514f
C334 VTAIL.n137 B 0.22868f
C335 VTAIL.t5 B 0.222855f
C336 VTAIL.t0 B 0.222855f
C337 VTAIL.n138 B 1.91432f
C338 VTAIL.n139 B 0.443314f
C339 VTAIL.n140 B 0.032184f
C340 VTAIL.n141 B 0.023346f
C341 VTAIL.n142 B 0.012545f
C342 VTAIL.n143 B 0.029651f
C343 VTAIL.n144 B 0.013283f
C344 VTAIL.n145 B 0.023346f
C345 VTAIL.n146 B 0.012545f
C346 VTAIL.n147 B 0.029651f
C347 VTAIL.n148 B 0.013283f
C348 VTAIL.n149 B 0.023346f
C349 VTAIL.n150 B 0.012914f
C350 VTAIL.n151 B 0.029651f
C351 VTAIL.n152 B 0.012545f
C352 VTAIL.n153 B 0.013283f
C353 VTAIL.n154 B 0.023346f
C354 VTAIL.n155 B 0.012545f
C355 VTAIL.n156 B 0.029651f
C356 VTAIL.n157 B 0.013283f
C357 VTAIL.n158 B 0.023346f
C358 VTAIL.n159 B 0.012545f
C359 VTAIL.n160 B 0.022239f
C360 VTAIL.n161 B 0.020961f
C361 VTAIL.t4 B 0.050089f
C362 VTAIL.n162 B 0.169035f
C363 VTAIL.n163 B 1.18605f
C364 VTAIL.n164 B 0.012545f
C365 VTAIL.n165 B 0.013283f
C366 VTAIL.n166 B 0.029651f
C367 VTAIL.n167 B 0.029651f
C368 VTAIL.n168 B 0.013283f
C369 VTAIL.n169 B 0.012545f
C370 VTAIL.n170 B 0.023346f
C371 VTAIL.n171 B 0.023346f
C372 VTAIL.n172 B 0.012545f
C373 VTAIL.n173 B 0.013283f
C374 VTAIL.n174 B 0.029651f
C375 VTAIL.n175 B 0.029651f
C376 VTAIL.n176 B 0.013283f
C377 VTAIL.n177 B 0.012545f
C378 VTAIL.n178 B 0.023346f
C379 VTAIL.n179 B 0.023346f
C380 VTAIL.n180 B 0.012545f
C381 VTAIL.n181 B 0.013283f
C382 VTAIL.n182 B 0.029651f
C383 VTAIL.n183 B 0.029651f
C384 VTAIL.n184 B 0.029651f
C385 VTAIL.n185 B 0.012914f
C386 VTAIL.n186 B 0.012545f
C387 VTAIL.n187 B 0.023346f
C388 VTAIL.n188 B 0.023346f
C389 VTAIL.n189 B 0.012545f
C390 VTAIL.n190 B 0.013283f
C391 VTAIL.n191 B 0.029651f
C392 VTAIL.n192 B 0.029651f
C393 VTAIL.n193 B 0.013283f
C394 VTAIL.n194 B 0.012545f
C395 VTAIL.n195 B 0.023346f
C396 VTAIL.n196 B 0.023346f
C397 VTAIL.n197 B 0.012545f
C398 VTAIL.n198 B 0.013283f
C399 VTAIL.n199 B 0.029651f
C400 VTAIL.n200 B 0.063076f
C401 VTAIL.n201 B 0.013283f
C402 VTAIL.n202 B 0.012545f
C403 VTAIL.n203 B 0.052686f
C404 VTAIL.n204 B 0.03514f
C405 VTAIL.n205 B 1.35187f
C406 VTAIL.n206 B 0.032184f
C407 VTAIL.n207 B 0.023346f
C408 VTAIL.n208 B 0.012545f
C409 VTAIL.n209 B 0.029651f
C410 VTAIL.n210 B 0.013283f
C411 VTAIL.n211 B 0.023346f
C412 VTAIL.n212 B 0.012545f
C413 VTAIL.n213 B 0.029651f
C414 VTAIL.n214 B 0.013283f
C415 VTAIL.n215 B 0.023346f
C416 VTAIL.n216 B 0.012914f
C417 VTAIL.n217 B 0.029651f
C418 VTAIL.n218 B 0.013283f
C419 VTAIL.n219 B 0.023346f
C420 VTAIL.n220 B 0.012545f
C421 VTAIL.n221 B 0.029651f
C422 VTAIL.n222 B 0.013283f
C423 VTAIL.n223 B 0.023346f
C424 VTAIL.n224 B 0.012545f
C425 VTAIL.n225 B 0.022239f
C426 VTAIL.n226 B 0.020961f
C427 VTAIL.t7 B 0.050089f
C428 VTAIL.n227 B 0.169035f
C429 VTAIL.n228 B 1.18605f
C430 VTAIL.n229 B 0.012545f
C431 VTAIL.n230 B 0.013283f
C432 VTAIL.n231 B 0.029651f
C433 VTAIL.n232 B 0.029651f
C434 VTAIL.n233 B 0.013283f
C435 VTAIL.n234 B 0.012545f
C436 VTAIL.n235 B 0.023346f
C437 VTAIL.n236 B 0.023346f
C438 VTAIL.n237 B 0.012545f
C439 VTAIL.n238 B 0.013283f
C440 VTAIL.n239 B 0.029651f
C441 VTAIL.n240 B 0.029651f
C442 VTAIL.n241 B 0.013283f
C443 VTAIL.n242 B 0.012545f
C444 VTAIL.n243 B 0.023346f
C445 VTAIL.n244 B 0.023346f
C446 VTAIL.n245 B 0.012545f
C447 VTAIL.n246 B 0.012545f
C448 VTAIL.n247 B 0.013283f
C449 VTAIL.n248 B 0.029651f
C450 VTAIL.n249 B 0.029651f
C451 VTAIL.n250 B 0.029651f
C452 VTAIL.n251 B 0.012914f
C453 VTAIL.n252 B 0.012545f
C454 VTAIL.n253 B 0.023346f
C455 VTAIL.n254 B 0.023346f
C456 VTAIL.n255 B 0.012545f
C457 VTAIL.n256 B 0.013283f
C458 VTAIL.n257 B 0.029651f
C459 VTAIL.n258 B 0.029651f
C460 VTAIL.n259 B 0.013283f
C461 VTAIL.n260 B 0.012545f
C462 VTAIL.n261 B 0.023346f
C463 VTAIL.n262 B 0.023346f
C464 VTAIL.n263 B 0.012545f
C465 VTAIL.n264 B 0.013283f
C466 VTAIL.n265 B 0.029651f
C467 VTAIL.n266 B 0.063076f
C468 VTAIL.n267 B 0.013283f
C469 VTAIL.n268 B 0.012545f
C470 VTAIL.n269 B 0.052686f
C471 VTAIL.n270 B 0.03514f
C472 VTAIL.n271 B 1.31847f
C473 VDD2.n0 B 0.030068f
C474 VDD2.n1 B 0.02181f
C475 VDD2.n2 B 0.01172f
C476 VDD2.n3 B 0.027701f
C477 VDD2.n4 B 0.012409f
C478 VDD2.n5 B 0.02181f
C479 VDD2.n6 B 0.01172f
C480 VDD2.n7 B 0.027701f
C481 VDD2.n8 B 0.012409f
C482 VDD2.n9 B 0.02181f
C483 VDD2.n10 B 0.012065f
C484 VDD2.n11 B 0.027701f
C485 VDD2.n12 B 0.012409f
C486 VDD2.n13 B 0.02181f
C487 VDD2.n14 B 0.01172f
C488 VDD2.n15 B 0.027701f
C489 VDD2.n16 B 0.012409f
C490 VDD2.n17 B 0.02181f
C491 VDD2.n18 B 0.01172f
C492 VDD2.n19 B 0.020776f
C493 VDD2.n20 B 0.019583f
C494 VDD2.t2 B 0.046796f
C495 VDD2.n21 B 0.157919f
C496 VDD2.n22 B 1.10805f
C497 VDD2.n23 B 0.01172f
C498 VDD2.n24 B 0.012409f
C499 VDD2.n25 B 0.027701f
C500 VDD2.n26 B 0.027701f
C501 VDD2.n27 B 0.012409f
C502 VDD2.n28 B 0.01172f
C503 VDD2.n29 B 0.02181f
C504 VDD2.n30 B 0.02181f
C505 VDD2.n31 B 0.01172f
C506 VDD2.n32 B 0.012409f
C507 VDD2.n33 B 0.027701f
C508 VDD2.n34 B 0.027701f
C509 VDD2.n35 B 0.012409f
C510 VDD2.n36 B 0.01172f
C511 VDD2.n37 B 0.02181f
C512 VDD2.n38 B 0.02181f
C513 VDD2.n39 B 0.01172f
C514 VDD2.n40 B 0.01172f
C515 VDD2.n41 B 0.012409f
C516 VDD2.n42 B 0.027701f
C517 VDD2.n43 B 0.027701f
C518 VDD2.n44 B 0.027701f
C519 VDD2.n45 B 0.012065f
C520 VDD2.n46 B 0.01172f
C521 VDD2.n47 B 0.02181f
C522 VDD2.n48 B 0.02181f
C523 VDD2.n49 B 0.01172f
C524 VDD2.n50 B 0.012409f
C525 VDD2.n51 B 0.027701f
C526 VDD2.n52 B 0.027701f
C527 VDD2.n53 B 0.012409f
C528 VDD2.n54 B 0.01172f
C529 VDD2.n55 B 0.02181f
C530 VDD2.n56 B 0.02181f
C531 VDD2.n57 B 0.01172f
C532 VDD2.n58 B 0.012409f
C533 VDD2.n59 B 0.027701f
C534 VDD2.n60 B 0.058928f
C535 VDD2.n61 B 0.012409f
C536 VDD2.n62 B 0.01172f
C537 VDD2.n63 B 0.049222f
C538 VDD2.n64 B 0.050569f
C539 VDD2.t1 B 0.2082f
C540 VDD2.t3 B 0.2082f
C541 VDD2.n65 B 1.85676f
C542 VDD2.n66 B 1.91062f
C543 VDD2.n67 B 0.030068f
C544 VDD2.n68 B 0.02181f
C545 VDD2.n69 B 0.01172f
C546 VDD2.n70 B 0.027701f
C547 VDD2.n71 B 0.012409f
C548 VDD2.n72 B 0.02181f
C549 VDD2.n73 B 0.01172f
C550 VDD2.n74 B 0.027701f
C551 VDD2.n75 B 0.012409f
C552 VDD2.n76 B 0.02181f
C553 VDD2.n77 B 0.012065f
C554 VDD2.n78 B 0.027701f
C555 VDD2.n79 B 0.01172f
C556 VDD2.n80 B 0.012409f
C557 VDD2.n81 B 0.02181f
C558 VDD2.n82 B 0.01172f
C559 VDD2.n83 B 0.027701f
C560 VDD2.n84 B 0.012409f
C561 VDD2.n85 B 0.02181f
C562 VDD2.n86 B 0.01172f
C563 VDD2.n87 B 0.020776f
C564 VDD2.n88 B 0.019583f
C565 VDD2.t0 B 0.046796f
C566 VDD2.n89 B 0.157919f
C567 VDD2.n90 B 1.10805f
C568 VDD2.n91 B 0.01172f
C569 VDD2.n92 B 0.012409f
C570 VDD2.n93 B 0.027701f
C571 VDD2.n94 B 0.027701f
C572 VDD2.n95 B 0.012409f
C573 VDD2.n96 B 0.01172f
C574 VDD2.n97 B 0.02181f
C575 VDD2.n98 B 0.02181f
C576 VDD2.n99 B 0.01172f
C577 VDD2.n100 B 0.012409f
C578 VDD2.n101 B 0.027701f
C579 VDD2.n102 B 0.027701f
C580 VDD2.n103 B 0.012409f
C581 VDD2.n104 B 0.01172f
C582 VDD2.n105 B 0.02181f
C583 VDD2.n106 B 0.02181f
C584 VDD2.n107 B 0.01172f
C585 VDD2.n108 B 0.012409f
C586 VDD2.n109 B 0.027701f
C587 VDD2.n110 B 0.027701f
C588 VDD2.n111 B 0.027701f
C589 VDD2.n112 B 0.012065f
C590 VDD2.n113 B 0.01172f
C591 VDD2.n114 B 0.02181f
C592 VDD2.n115 B 0.02181f
C593 VDD2.n116 B 0.01172f
C594 VDD2.n117 B 0.012409f
C595 VDD2.n118 B 0.027701f
C596 VDD2.n119 B 0.027701f
C597 VDD2.n120 B 0.012409f
C598 VDD2.n121 B 0.01172f
C599 VDD2.n122 B 0.02181f
C600 VDD2.n123 B 0.02181f
C601 VDD2.n124 B 0.01172f
C602 VDD2.n125 B 0.012409f
C603 VDD2.n126 B 0.027701f
C604 VDD2.n127 B 0.058928f
C605 VDD2.n128 B 0.012409f
C606 VDD2.n129 B 0.01172f
C607 VDD2.n130 B 0.049222f
C608 VDD2.n131 B 0.047898f
C609 VDD2.n132 B 1.96822f
C610 VDD2.t4 B 0.2082f
C611 VDD2.t5 B 0.2082f
C612 VDD2.n133 B 1.85674f
C613 VN.n0 B 0.033009f
C614 VN.t4 B 1.58652f
C615 VN.n1 B 0.059967f
C616 VN.t2 B 1.69563f
C617 VN.t1 B 1.58652f
C618 VN.n2 B 0.650416f
C619 VN.n3 B 0.639522f
C620 VN.n4 B 0.209938f
C621 VN.n5 B 0.033009f
C622 VN.n6 B 0.031611f
C623 VN.n7 B 0.052911f
C624 VN.n8 B 0.645795f
C625 VN.n9 B 0.030174f
C626 VN.n10 B 0.033009f
C627 VN.t3 B 1.58652f
C628 VN.n11 B 0.059967f
C629 VN.t5 B 1.69563f
C630 VN.t0 B 1.58652f
C631 VN.n12 B 0.650416f
C632 VN.n13 B 0.639522f
C633 VN.n14 B 0.209938f
C634 VN.n15 B 0.033009f
C635 VN.n16 B 0.031611f
C636 VN.n17 B 0.052911f
C637 VN.n18 B 0.645795f
C638 VN.n19 B 1.51011f
.ends

