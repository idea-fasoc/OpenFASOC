* NGSPICE file created from diff_pair_sample_0698.ext - technology: sky130A

.subckt diff_pair_sample_0698 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=2.98
X1 VDD2.t7 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=2.98
X2 VDD1.t6 VP.t1 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=2.98
X3 VTAIL.t13 VP.t2 VDD1.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=1.8678 ps=11.65 w=11.32 l=2.98
X4 VTAIL.t2 VN.t1 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=1.8678 ps=11.65 w=11.32 l=2.98
X5 VDD1.t4 VP.t3 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=4.4148 ps=23.42 w=11.32 l=2.98
X6 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=0 ps=0 w=11.32 l=2.98
X7 VTAIL.t0 VN.t2 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=1.8678 ps=11.65 w=11.32 l=2.98
X8 VDD1.t3 VP.t4 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=4.4148 ps=23.42 w=11.32 l=2.98
X9 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=0 ps=0 w=11.32 l=2.98
X10 VDD2.t4 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=4.4148 ps=23.42 w=11.32 l=2.98
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=0 ps=0 w=11.32 l=2.98
X12 VDD2.t3 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=2.98
X13 VTAIL.t11 VP.t5 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=1.8678 ps=11.65 w=11.32 l=2.98
X14 VDD2.t2 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=4.4148 ps=23.42 w=11.32 l=2.98
X15 VTAIL.t9 VP.t6 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=2.98
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.4148 pd=23.42 as=0 ps=0 w=11.32 l=2.98
X17 VTAIL.t5 VN.t6 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=2.98
X18 VTAIL.t15 VP.t7 VDD1.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=2.98
X19 VTAIL.t7 VN.t7 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=1.8678 pd=11.65 as=1.8678 ps=11.65 w=11.32 l=2.98
R0 VP.n21 VP.n20 161.3
R1 VP.n22 VP.n17 161.3
R2 VP.n24 VP.n23 161.3
R3 VP.n25 VP.n16 161.3
R4 VP.n27 VP.n26 161.3
R5 VP.n28 VP.n15 161.3
R6 VP.n30 VP.n29 161.3
R7 VP.n32 VP.n14 161.3
R8 VP.n34 VP.n33 161.3
R9 VP.n35 VP.n13 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n38 VP.n12 161.3
R12 VP.n40 VP.n39 161.3
R13 VP.n73 VP.n72 161.3
R14 VP.n71 VP.n1 161.3
R15 VP.n70 VP.n69 161.3
R16 VP.n68 VP.n2 161.3
R17 VP.n67 VP.n66 161.3
R18 VP.n65 VP.n3 161.3
R19 VP.n63 VP.n62 161.3
R20 VP.n61 VP.n4 161.3
R21 VP.n60 VP.n59 161.3
R22 VP.n58 VP.n5 161.3
R23 VP.n57 VP.n56 161.3
R24 VP.n55 VP.n6 161.3
R25 VP.n54 VP.n53 161.3
R26 VP.n51 VP.n7 161.3
R27 VP.n50 VP.n49 161.3
R28 VP.n48 VP.n8 161.3
R29 VP.n47 VP.n46 161.3
R30 VP.n45 VP.n9 161.3
R31 VP.n44 VP.n43 161.3
R32 VP.n18 VP.t2 123.234
R33 VP.n10 VP.t5 91.5481
R34 VP.n52 VP.t1 91.5481
R35 VP.n64 VP.t6 91.5481
R36 VP.n0 VP.t3 91.5481
R37 VP.n11 VP.t4 91.5481
R38 VP.n31 VP.t7 91.5481
R39 VP.n19 VP.t0 91.5481
R40 VP.n42 VP.n10 67.2516
R41 VP.n74 VP.n0 67.2516
R42 VP.n41 VP.n11 67.2516
R43 VP.n19 VP.n18 66.0815
R44 VP.n46 VP.n8 56.4773
R45 VP.n70 VP.n2 56.4773
R46 VP.n37 VP.n13 56.4773
R47 VP.n42 VP.n41 52.3173
R48 VP.n58 VP.n57 40.4106
R49 VP.n59 VP.n58 40.4106
R50 VP.n26 VP.n25 40.4106
R51 VP.n25 VP.n24 40.4106
R52 VP.n45 VP.n44 24.3439
R53 VP.n46 VP.n45 24.3439
R54 VP.n50 VP.n8 24.3439
R55 VP.n51 VP.n50 24.3439
R56 VP.n53 VP.n6 24.3439
R57 VP.n57 VP.n6 24.3439
R58 VP.n59 VP.n4 24.3439
R59 VP.n63 VP.n4 24.3439
R60 VP.n66 VP.n65 24.3439
R61 VP.n66 VP.n2 24.3439
R62 VP.n71 VP.n70 24.3439
R63 VP.n72 VP.n71 24.3439
R64 VP.n38 VP.n37 24.3439
R65 VP.n39 VP.n38 24.3439
R66 VP.n26 VP.n15 24.3439
R67 VP.n30 VP.n15 24.3439
R68 VP.n33 VP.n32 24.3439
R69 VP.n33 VP.n13 24.3439
R70 VP.n20 VP.n17 24.3439
R71 VP.n24 VP.n17 24.3439
R72 VP.n44 VP.n10 22.6399
R73 VP.n72 VP.n0 22.6399
R74 VP.n39 VP.n11 22.6399
R75 VP.n52 VP.n51 16.7975
R76 VP.n65 VP.n64 16.7975
R77 VP.n32 VP.n31 16.7975
R78 VP.n53 VP.n52 7.54696
R79 VP.n64 VP.n63 7.54696
R80 VP.n31 VP.n30 7.54696
R81 VP.n20 VP.n19 7.54696
R82 VP.n21 VP.n18 5.3732
R83 VP.n41 VP.n40 0.355081
R84 VP.n43 VP.n42 0.355081
R85 VP.n74 VP.n73 0.355081
R86 VP VP.n74 0.26685
R87 VP.n22 VP.n21 0.189894
R88 VP.n23 VP.n22 0.189894
R89 VP.n23 VP.n16 0.189894
R90 VP.n27 VP.n16 0.189894
R91 VP.n28 VP.n27 0.189894
R92 VP.n29 VP.n28 0.189894
R93 VP.n29 VP.n14 0.189894
R94 VP.n34 VP.n14 0.189894
R95 VP.n35 VP.n34 0.189894
R96 VP.n36 VP.n35 0.189894
R97 VP.n36 VP.n12 0.189894
R98 VP.n40 VP.n12 0.189894
R99 VP.n43 VP.n9 0.189894
R100 VP.n47 VP.n9 0.189894
R101 VP.n48 VP.n47 0.189894
R102 VP.n49 VP.n48 0.189894
R103 VP.n49 VP.n7 0.189894
R104 VP.n54 VP.n7 0.189894
R105 VP.n55 VP.n54 0.189894
R106 VP.n56 VP.n55 0.189894
R107 VP.n56 VP.n5 0.189894
R108 VP.n60 VP.n5 0.189894
R109 VP.n61 VP.n60 0.189894
R110 VP.n62 VP.n61 0.189894
R111 VP.n62 VP.n3 0.189894
R112 VP.n67 VP.n3 0.189894
R113 VP.n68 VP.n67 0.189894
R114 VP.n69 VP.n68 0.189894
R115 VP.n69 VP.n1 0.189894
R116 VP.n73 VP.n1 0.189894
R117 VTAIL.n498 VTAIL.n442 289.615
R118 VTAIL.n58 VTAIL.n2 289.615
R119 VTAIL.n120 VTAIL.n64 289.615
R120 VTAIL.n184 VTAIL.n128 289.615
R121 VTAIL.n436 VTAIL.n380 289.615
R122 VTAIL.n372 VTAIL.n316 289.615
R123 VTAIL.n310 VTAIL.n254 289.615
R124 VTAIL.n246 VTAIL.n190 289.615
R125 VTAIL.n463 VTAIL.n462 185
R126 VTAIL.n465 VTAIL.n464 185
R127 VTAIL.n458 VTAIL.n457 185
R128 VTAIL.n471 VTAIL.n470 185
R129 VTAIL.n473 VTAIL.n472 185
R130 VTAIL.n454 VTAIL.n453 185
R131 VTAIL.n480 VTAIL.n479 185
R132 VTAIL.n481 VTAIL.n452 185
R133 VTAIL.n483 VTAIL.n482 185
R134 VTAIL.n450 VTAIL.n449 185
R135 VTAIL.n489 VTAIL.n488 185
R136 VTAIL.n491 VTAIL.n490 185
R137 VTAIL.n446 VTAIL.n445 185
R138 VTAIL.n497 VTAIL.n496 185
R139 VTAIL.n499 VTAIL.n498 185
R140 VTAIL.n23 VTAIL.n22 185
R141 VTAIL.n25 VTAIL.n24 185
R142 VTAIL.n18 VTAIL.n17 185
R143 VTAIL.n31 VTAIL.n30 185
R144 VTAIL.n33 VTAIL.n32 185
R145 VTAIL.n14 VTAIL.n13 185
R146 VTAIL.n40 VTAIL.n39 185
R147 VTAIL.n41 VTAIL.n12 185
R148 VTAIL.n43 VTAIL.n42 185
R149 VTAIL.n10 VTAIL.n9 185
R150 VTAIL.n49 VTAIL.n48 185
R151 VTAIL.n51 VTAIL.n50 185
R152 VTAIL.n6 VTAIL.n5 185
R153 VTAIL.n57 VTAIL.n56 185
R154 VTAIL.n59 VTAIL.n58 185
R155 VTAIL.n85 VTAIL.n84 185
R156 VTAIL.n87 VTAIL.n86 185
R157 VTAIL.n80 VTAIL.n79 185
R158 VTAIL.n93 VTAIL.n92 185
R159 VTAIL.n95 VTAIL.n94 185
R160 VTAIL.n76 VTAIL.n75 185
R161 VTAIL.n102 VTAIL.n101 185
R162 VTAIL.n103 VTAIL.n74 185
R163 VTAIL.n105 VTAIL.n104 185
R164 VTAIL.n72 VTAIL.n71 185
R165 VTAIL.n111 VTAIL.n110 185
R166 VTAIL.n113 VTAIL.n112 185
R167 VTAIL.n68 VTAIL.n67 185
R168 VTAIL.n119 VTAIL.n118 185
R169 VTAIL.n121 VTAIL.n120 185
R170 VTAIL.n149 VTAIL.n148 185
R171 VTAIL.n151 VTAIL.n150 185
R172 VTAIL.n144 VTAIL.n143 185
R173 VTAIL.n157 VTAIL.n156 185
R174 VTAIL.n159 VTAIL.n158 185
R175 VTAIL.n140 VTAIL.n139 185
R176 VTAIL.n166 VTAIL.n165 185
R177 VTAIL.n167 VTAIL.n138 185
R178 VTAIL.n169 VTAIL.n168 185
R179 VTAIL.n136 VTAIL.n135 185
R180 VTAIL.n175 VTAIL.n174 185
R181 VTAIL.n177 VTAIL.n176 185
R182 VTAIL.n132 VTAIL.n131 185
R183 VTAIL.n183 VTAIL.n182 185
R184 VTAIL.n185 VTAIL.n184 185
R185 VTAIL.n437 VTAIL.n436 185
R186 VTAIL.n435 VTAIL.n434 185
R187 VTAIL.n384 VTAIL.n383 185
R188 VTAIL.n429 VTAIL.n428 185
R189 VTAIL.n427 VTAIL.n426 185
R190 VTAIL.n388 VTAIL.n387 185
R191 VTAIL.n392 VTAIL.n390 185
R192 VTAIL.n421 VTAIL.n420 185
R193 VTAIL.n419 VTAIL.n418 185
R194 VTAIL.n394 VTAIL.n393 185
R195 VTAIL.n413 VTAIL.n412 185
R196 VTAIL.n411 VTAIL.n410 185
R197 VTAIL.n398 VTAIL.n397 185
R198 VTAIL.n405 VTAIL.n404 185
R199 VTAIL.n403 VTAIL.n402 185
R200 VTAIL.n373 VTAIL.n372 185
R201 VTAIL.n371 VTAIL.n370 185
R202 VTAIL.n320 VTAIL.n319 185
R203 VTAIL.n365 VTAIL.n364 185
R204 VTAIL.n363 VTAIL.n362 185
R205 VTAIL.n324 VTAIL.n323 185
R206 VTAIL.n328 VTAIL.n326 185
R207 VTAIL.n357 VTAIL.n356 185
R208 VTAIL.n355 VTAIL.n354 185
R209 VTAIL.n330 VTAIL.n329 185
R210 VTAIL.n349 VTAIL.n348 185
R211 VTAIL.n347 VTAIL.n346 185
R212 VTAIL.n334 VTAIL.n333 185
R213 VTAIL.n341 VTAIL.n340 185
R214 VTAIL.n339 VTAIL.n338 185
R215 VTAIL.n311 VTAIL.n310 185
R216 VTAIL.n309 VTAIL.n308 185
R217 VTAIL.n258 VTAIL.n257 185
R218 VTAIL.n303 VTAIL.n302 185
R219 VTAIL.n301 VTAIL.n300 185
R220 VTAIL.n262 VTAIL.n261 185
R221 VTAIL.n266 VTAIL.n264 185
R222 VTAIL.n295 VTAIL.n294 185
R223 VTAIL.n293 VTAIL.n292 185
R224 VTAIL.n268 VTAIL.n267 185
R225 VTAIL.n287 VTAIL.n286 185
R226 VTAIL.n285 VTAIL.n284 185
R227 VTAIL.n272 VTAIL.n271 185
R228 VTAIL.n279 VTAIL.n278 185
R229 VTAIL.n277 VTAIL.n276 185
R230 VTAIL.n247 VTAIL.n246 185
R231 VTAIL.n245 VTAIL.n244 185
R232 VTAIL.n194 VTAIL.n193 185
R233 VTAIL.n239 VTAIL.n238 185
R234 VTAIL.n237 VTAIL.n236 185
R235 VTAIL.n198 VTAIL.n197 185
R236 VTAIL.n202 VTAIL.n200 185
R237 VTAIL.n231 VTAIL.n230 185
R238 VTAIL.n229 VTAIL.n228 185
R239 VTAIL.n204 VTAIL.n203 185
R240 VTAIL.n223 VTAIL.n222 185
R241 VTAIL.n221 VTAIL.n220 185
R242 VTAIL.n208 VTAIL.n207 185
R243 VTAIL.n215 VTAIL.n214 185
R244 VTAIL.n213 VTAIL.n212 185
R245 VTAIL.n461 VTAIL.t6 149.524
R246 VTAIL.n21 VTAIL.t0 149.524
R247 VTAIL.n83 VTAIL.t10 149.524
R248 VTAIL.n147 VTAIL.t11 149.524
R249 VTAIL.n401 VTAIL.t14 149.524
R250 VTAIL.n337 VTAIL.t13 149.524
R251 VTAIL.n275 VTAIL.t1 149.524
R252 VTAIL.n211 VTAIL.t2 149.524
R253 VTAIL.n464 VTAIL.n463 104.615
R254 VTAIL.n464 VTAIL.n457 104.615
R255 VTAIL.n471 VTAIL.n457 104.615
R256 VTAIL.n472 VTAIL.n471 104.615
R257 VTAIL.n472 VTAIL.n453 104.615
R258 VTAIL.n480 VTAIL.n453 104.615
R259 VTAIL.n481 VTAIL.n480 104.615
R260 VTAIL.n482 VTAIL.n481 104.615
R261 VTAIL.n482 VTAIL.n449 104.615
R262 VTAIL.n489 VTAIL.n449 104.615
R263 VTAIL.n490 VTAIL.n489 104.615
R264 VTAIL.n490 VTAIL.n445 104.615
R265 VTAIL.n497 VTAIL.n445 104.615
R266 VTAIL.n498 VTAIL.n497 104.615
R267 VTAIL.n24 VTAIL.n23 104.615
R268 VTAIL.n24 VTAIL.n17 104.615
R269 VTAIL.n31 VTAIL.n17 104.615
R270 VTAIL.n32 VTAIL.n31 104.615
R271 VTAIL.n32 VTAIL.n13 104.615
R272 VTAIL.n40 VTAIL.n13 104.615
R273 VTAIL.n41 VTAIL.n40 104.615
R274 VTAIL.n42 VTAIL.n41 104.615
R275 VTAIL.n42 VTAIL.n9 104.615
R276 VTAIL.n49 VTAIL.n9 104.615
R277 VTAIL.n50 VTAIL.n49 104.615
R278 VTAIL.n50 VTAIL.n5 104.615
R279 VTAIL.n57 VTAIL.n5 104.615
R280 VTAIL.n58 VTAIL.n57 104.615
R281 VTAIL.n86 VTAIL.n85 104.615
R282 VTAIL.n86 VTAIL.n79 104.615
R283 VTAIL.n93 VTAIL.n79 104.615
R284 VTAIL.n94 VTAIL.n93 104.615
R285 VTAIL.n94 VTAIL.n75 104.615
R286 VTAIL.n102 VTAIL.n75 104.615
R287 VTAIL.n103 VTAIL.n102 104.615
R288 VTAIL.n104 VTAIL.n103 104.615
R289 VTAIL.n104 VTAIL.n71 104.615
R290 VTAIL.n111 VTAIL.n71 104.615
R291 VTAIL.n112 VTAIL.n111 104.615
R292 VTAIL.n112 VTAIL.n67 104.615
R293 VTAIL.n119 VTAIL.n67 104.615
R294 VTAIL.n120 VTAIL.n119 104.615
R295 VTAIL.n150 VTAIL.n149 104.615
R296 VTAIL.n150 VTAIL.n143 104.615
R297 VTAIL.n157 VTAIL.n143 104.615
R298 VTAIL.n158 VTAIL.n157 104.615
R299 VTAIL.n158 VTAIL.n139 104.615
R300 VTAIL.n166 VTAIL.n139 104.615
R301 VTAIL.n167 VTAIL.n166 104.615
R302 VTAIL.n168 VTAIL.n167 104.615
R303 VTAIL.n168 VTAIL.n135 104.615
R304 VTAIL.n175 VTAIL.n135 104.615
R305 VTAIL.n176 VTAIL.n175 104.615
R306 VTAIL.n176 VTAIL.n131 104.615
R307 VTAIL.n183 VTAIL.n131 104.615
R308 VTAIL.n184 VTAIL.n183 104.615
R309 VTAIL.n436 VTAIL.n435 104.615
R310 VTAIL.n435 VTAIL.n383 104.615
R311 VTAIL.n428 VTAIL.n383 104.615
R312 VTAIL.n428 VTAIL.n427 104.615
R313 VTAIL.n427 VTAIL.n387 104.615
R314 VTAIL.n392 VTAIL.n387 104.615
R315 VTAIL.n420 VTAIL.n392 104.615
R316 VTAIL.n420 VTAIL.n419 104.615
R317 VTAIL.n419 VTAIL.n393 104.615
R318 VTAIL.n412 VTAIL.n393 104.615
R319 VTAIL.n412 VTAIL.n411 104.615
R320 VTAIL.n411 VTAIL.n397 104.615
R321 VTAIL.n404 VTAIL.n397 104.615
R322 VTAIL.n404 VTAIL.n403 104.615
R323 VTAIL.n372 VTAIL.n371 104.615
R324 VTAIL.n371 VTAIL.n319 104.615
R325 VTAIL.n364 VTAIL.n319 104.615
R326 VTAIL.n364 VTAIL.n363 104.615
R327 VTAIL.n363 VTAIL.n323 104.615
R328 VTAIL.n328 VTAIL.n323 104.615
R329 VTAIL.n356 VTAIL.n328 104.615
R330 VTAIL.n356 VTAIL.n355 104.615
R331 VTAIL.n355 VTAIL.n329 104.615
R332 VTAIL.n348 VTAIL.n329 104.615
R333 VTAIL.n348 VTAIL.n347 104.615
R334 VTAIL.n347 VTAIL.n333 104.615
R335 VTAIL.n340 VTAIL.n333 104.615
R336 VTAIL.n340 VTAIL.n339 104.615
R337 VTAIL.n310 VTAIL.n309 104.615
R338 VTAIL.n309 VTAIL.n257 104.615
R339 VTAIL.n302 VTAIL.n257 104.615
R340 VTAIL.n302 VTAIL.n301 104.615
R341 VTAIL.n301 VTAIL.n261 104.615
R342 VTAIL.n266 VTAIL.n261 104.615
R343 VTAIL.n294 VTAIL.n266 104.615
R344 VTAIL.n294 VTAIL.n293 104.615
R345 VTAIL.n293 VTAIL.n267 104.615
R346 VTAIL.n286 VTAIL.n267 104.615
R347 VTAIL.n286 VTAIL.n285 104.615
R348 VTAIL.n285 VTAIL.n271 104.615
R349 VTAIL.n278 VTAIL.n271 104.615
R350 VTAIL.n278 VTAIL.n277 104.615
R351 VTAIL.n246 VTAIL.n245 104.615
R352 VTAIL.n245 VTAIL.n193 104.615
R353 VTAIL.n238 VTAIL.n193 104.615
R354 VTAIL.n238 VTAIL.n237 104.615
R355 VTAIL.n237 VTAIL.n197 104.615
R356 VTAIL.n202 VTAIL.n197 104.615
R357 VTAIL.n230 VTAIL.n202 104.615
R358 VTAIL.n230 VTAIL.n229 104.615
R359 VTAIL.n229 VTAIL.n203 104.615
R360 VTAIL.n222 VTAIL.n203 104.615
R361 VTAIL.n222 VTAIL.n221 104.615
R362 VTAIL.n221 VTAIL.n207 104.615
R363 VTAIL.n214 VTAIL.n207 104.615
R364 VTAIL.n214 VTAIL.n213 104.615
R365 VTAIL.n463 VTAIL.t6 52.3082
R366 VTAIL.n23 VTAIL.t0 52.3082
R367 VTAIL.n85 VTAIL.t10 52.3082
R368 VTAIL.n149 VTAIL.t11 52.3082
R369 VTAIL.n403 VTAIL.t14 52.3082
R370 VTAIL.n339 VTAIL.t13 52.3082
R371 VTAIL.n277 VTAIL.t1 52.3082
R372 VTAIL.n213 VTAIL.t2 52.3082
R373 VTAIL.n379 VTAIL.n378 43.8596
R374 VTAIL.n253 VTAIL.n252 43.8596
R375 VTAIL.n1 VTAIL.n0 43.8594
R376 VTAIL.n127 VTAIL.n126 43.8594
R377 VTAIL.n503 VTAIL.n502 30.6338
R378 VTAIL.n63 VTAIL.n62 30.6338
R379 VTAIL.n125 VTAIL.n124 30.6338
R380 VTAIL.n189 VTAIL.n188 30.6338
R381 VTAIL.n441 VTAIL.n440 30.6338
R382 VTAIL.n377 VTAIL.n376 30.6338
R383 VTAIL.n315 VTAIL.n314 30.6338
R384 VTAIL.n251 VTAIL.n250 30.6338
R385 VTAIL.n503 VTAIL.n441 24.9789
R386 VTAIL.n251 VTAIL.n189 24.9789
R387 VTAIL.n483 VTAIL.n450 13.1884
R388 VTAIL.n43 VTAIL.n10 13.1884
R389 VTAIL.n105 VTAIL.n72 13.1884
R390 VTAIL.n169 VTAIL.n136 13.1884
R391 VTAIL.n390 VTAIL.n388 13.1884
R392 VTAIL.n326 VTAIL.n324 13.1884
R393 VTAIL.n264 VTAIL.n262 13.1884
R394 VTAIL.n200 VTAIL.n198 13.1884
R395 VTAIL.n484 VTAIL.n452 12.8005
R396 VTAIL.n488 VTAIL.n487 12.8005
R397 VTAIL.n44 VTAIL.n12 12.8005
R398 VTAIL.n48 VTAIL.n47 12.8005
R399 VTAIL.n106 VTAIL.n74 12.8005
R400 VTAIL.n110 VTAIL.n109 12.8005
R401 VTAIL.n170 VTAIL.n138 12.8005
R402 VTAIL.n174 VTAIL.n173 12.8005
R403 VTAIL.n426 VTAIL.n425 12.8005
R404 VTAIL.n422 VTAIL.n421 12.8005
R405 VTAIL.n362 VTAIL.n361 12.8005
R406 VTAIL.n358 VTAIL.n357 12.8005
R407 VTAIL.n300 VTAIL.n299 12.8005
R408 VTAIL.n296 VTAIL.n295 12.8005
R409 VTAIL.n236 VTAIL.n235 12.8005
R410 VTAIL.n232 VTAIL.n231 12.8005
R411 VTAIL.n479 VTAIL.n478 12.0247
R412 VTAIL.n491 VTAIL.n448 12.0247
R413 VTAIL.n39 VTAIL.n38 12.0247
R414 VTAIL.n51 VTAIL.n8 12.0247
R415 VTAIL.n101 VTAIL.n100 12.0247
R416 VTAIL.n113 VTAIL.n70 12.0247
R417 VTAIL.n165 VTAIL.n164 12.0247
R418 VTAIL.n177 VTAIL.n134 12.0247
R419 VTAIL.n429 VTAIL.n386 12.0247
R420 VTAIL.n418 VTAIL.n391 12.0247
R421 VTAIL.n365 VTAIL.n322 12.0247
R422 VTAIL.n354 VTAIL.n327 12.0247
R423 VTAIL.n303 VTAIL.n260 12.0247
R424 VTAIL.n292 VTAIL.n265 12.0247
R425 VTAIL.n239 VTAIL.n196 12.0247
R426 VTAIL.n228 VTAIL.n201 12.0247
R427 VTAIL.n477 VTAIL.n454 11.249
R428 VTAIL.n492 VTAIL.n446 11.249
R429 VTAIL.n37 VTAIL.n14 11.249
R430 VTAIL.n52 VTAIL.n6 11.249
R431 VTAIL.n99 VTAIL.n76 11.249
R432 VTAIL.n114 VTAIL.n68 11.249
R433 VTAIL.n163 VTAIL.n140 11.249
R434 VTAIL.n178 VTAIL.n132 11.249
R435 VTAIL.n430 VTAIL.n384 11.249
R436 VTAIL.n417 VTAIL.n394 11.249
R437 VTAIL.n366 VTAIL.n320 11.249
R438 VTAIL.n353 VTAIL.n330 11.249
R439 VTAIL.n304 VTAIL.n258 11.249
R440 VTAIL.n291 VTAIL.n268 11.249
R441 VTAIL.n240 VTAIL.n194 11.249
R442 VTAIL.n227 VTAIL.n204 11.249
R443 VTAIL.n474 VTAIL.n473 10.4732
R444 VTAIL.n496 VTAIL.n495 10.4732
R445 VTAIL.n34 VTAIL.n33 10.4732
R446 VTAIL.n56 VTAIL.n55 10.4732
R447 VTAIL.n96 VTAIL.n95 10.4732
R448 VTAIL.n118 VTAIL.n117 10.4732
R449 VTAIL.n160 VTAIL.n159 10.4732
R450 VTAIL.n182 VTAIL.n181 10.4732
R451 VTAIL.n434 VTAIL.n433 10.4732
R452 VTAIL.n414 VTAIL.n413 10.4732
R453 VTAIL.n370 VTAIL.n369 10.4732
R454 VTAIL.n350 VTAIL.n349 10.4732
R455 VTAIL.n308 VTAIL.n307 10.4732
R456 VTAIL.n288 VTAIL.n287 10.4732
R457 VTAIL.n244 VTAIL.n243 10.4732
R458 VTAIL.n224 VTAIL.n223 10.4732
R459 VTAIL.n462 VTAIL.n461 10.2747
R460 VTAIL.n22 VTAIL.n21 10.2747
R461 VTAIL.n84 VTAIL.n83 10.2747
R462 VTAIL.n148 VTAIL.n147 10.2747
R463 VTAIL.n402 VTAIL.n401 10.2747
R464 VTAIL.n338 VTAIL.n337 10.2747
R465 VTAIL.n276 VTAIL.n275 10.2747
R466 VTAIL.n212 VTAIL.n211 10.2747
R467 VTAIL.n470 VTAIL.n456 9.69747
R468 VTAIL.n499 VTAIL.n444 9.69747
R469 VTAIL.n30 VTAIL.n16 9.69747
R470 VTAIL.n59 VTAIL.n4 9.69747
R471 VTAIL.n92 VTAIL.n78 9.69747
R472 VTAIL.n121 VTAIL.n66 9.69747
R473 VTAIL.n156 VTAIL.n142 9.69747
R474 VTAIL.n185 VTAIL.n130 9.69747
R475 VTAIL.n437 VTAIL.n382 9.69747
R476 VTAIL.n410 VTAIL.n396 9.69747
R477 VTAIL.n373 VTAIL.n318 9.69747
R478 VTAIL.n346 VTAIL.n332 9.69747
R479 VTAIL.n311 VTAIL.n256 9.69747
R480 VTAIL.n284 VTAIL.n270 9.69747
R481 VTAIL.n247 VTAIL.n192 9.69747
R482 VTAIL.n220 VTAIL.n206 9.69747
R483 VTAIL.n502 VTAIL.n501 9.45567
R484 VTAIL.n62 VTAIL.n61 9.45567
R485 VTAIL.n124 VTAIL.n123 9.45567
R486 VTAIL.n188 VTAIL.n187 9.45567
R487 VTAIL.n440 VTAIL.n439 9.45567
R488 VTAIL.n376 VTAIL.n375 9.45567
R489 VTAIL.n314 VTAIL.n313 9.45567
R490 VTAIL.n250 VTAIL.n249 9.45567
R491 VTAIL.n501 VTAIL.n500 9.3005
R492 VTAIL.n444 VTAIL.n443 9.3005
R493 VTAIL.n495 VTAIL.n494 9.3005
R494 VTAIL.n493 VTAIL.n492 9.3005
R495 VTAIL.n448 VTAIL.n447 9.3005
R496 VTAIL.n487 VTAIL.n486 9.3005
R497 VTAIL.n460 VTAIL.n459 9.3005
R498 VTAIL.n467 VTAIL.n466 9.3005
R499 VTAIL.n469 VTAIL.n468 9.3005
R500 VTAIL.n456 VTAIL.n455 9.3005
R501 VTAIL.n475 VTAIL.n474 9.3005
R502 VTAIL.n477 VTAIL.n476 9.3005
R503 VTAIL.n478 VTAIL.n451 9.3005
R504 VTAIL.n485 VTAIL.n484 9.3005
R505 VTAIL.n61 VTAIL.n60 9.3005
R506 VTAIL.n4 VTAIL.n3 9.3005
R507 VTAIL.n55 VTAIL.n54 9.3005
R508 VTAIL.n53 VTAIL.n52 9.3005
R509 VTAIL.n8 VTAIL.n7 9.3005
R510 VTAIL.n47 VTAIL.n46 9.3005
R511 VTAIL.n20 VTAIL.n19 9.3005
R512 VTAIL.n27 VTAIL.n26 9.3005
R513 VTAIL.n29 VTAIL.n28 9.3005
R514 VTAIL.n16 VTAIL.n15 9.3005
R515 VTAIL.n35 VTAIL.n34 9.3005
R516 VTAIL.n37 VTAIL.n36 9.3005
R517 VTAIL.n38 VTAIL.n11 9.3005
R518 VTAIL.n45 VTAIL.n44 9.3005
R519 VTAIL.n123 VTAIL.n122 9.3005
R520 VTAIL.n66 VTAIL.n65 9.3005
R521 VTAIL.n117 VTAIL.n116 9.3005
R522 VTAIL.n115 VTAIL.n114 9.3005
R523 VTAIL.n70 VTAIL.n69 9.3005
R524 VTAIL.n109 VTAIL.n108 9.3005
R525 VTAIL.n82 VTAIL.n81 9.3005
R526 VTAIL.n89 VTAIL.n88 9.3005
R527 VTAIL.n91 VTAIL.n90 9.3005
R528 VTAIL.n78 VTAIL.n77 9.3005
R529 VTAIL.n97 VTAIL.n96 9.3005
R530 VTAIL.n99 VTAIL.n98 9.3005
R531 VTAIL.n100 VTAIL.n73 9.3005
R532 VTAIL.n107 VTAIL.n106 9.3005
R533 VTAIL.n187 VTAIL.n186 9.3005
R534 VTAIL.n130 VTAIL.n129 9.3005
R535 VTAIL.n181 VTAIL.n180 9.3005
R536 VTAIL.n179 VTAIL.n178 9.3005
R537 VTAIL.n134 VTAIL.n133 9.3005
R538 VTAIL.n173 VTAIL.n172 9.3005
R539 VTAIL.n146 VTAIL.n145 9.3005
R540 VTAIL.n153 VTAIL.n152 9.3005
R541 VTAIL.n155 VTAIL.n154 9.3005
R542 VTAIL.n142 VTAIL.n141 9.3005
R543 VTAIL.n161 VTAIL.n160 9.3005
R544 VTAIL.n163 VTAIL.n162 9.3005
R545 VTAIL.n164 VTAIL.n137 9.3005
R546 VTAIL.n171 VTAIL.n170 9.3005
R547 VTAIL.n400 VTAIL.n399 9.3005
R548 VTAIL.n407 VTAIL.n406 9.3005
R549 VTAIL.n409 VTAIL.n408 9.3005
R550 VTAIL.n396 VTAIL.n395 9.3005
R551 VTAIL.n415 VTAIL.n414 9.3005
R552 VTAIL.n417 VTAIL.n416 9.3005
R553 VTAIL.n391 VTAIL.n389 9.3005
R554 VTAIL.n423 VTAIL.n422 9.3005
R555 VTAIL.n439 VTAIL.n438 9.3005
R556 VTAIL.n382 VTAIL.n381 9.3005
R557 VTAIL.n433 VTAIL.n432 9.3005
R558 VTAIL.n431 VTAIL.n430 9.3005
R559 VTAIL.n386 VTAIL.n385 9.3005
R560 VTAIL.n425 VTAIL.n424 9.3005
R561 VTAIL.n336 VTAIL.n335 9.3005
R562 VTAIL.n343 VTAIL.n342 9.3005
R563 VTAIL.n345 VTAIL.n344 9.3005
R564 VTAIL.n332 VTAIL.n331 9.3005
R565 VTAIL.n351 VTAIL.n350 9.3005
R566 VTAIL.n353 VTAIL.n352 9.3005
R567 VTAIL.n327 VTAIL.n325 9.3005
R568 VTAIL.n359 VTAIL.n358 9.3005
R569 VTAIL.n375 VTAIL.n374 9.3005
R570 VTAIL.n318 VTAIL.n317 9.3005
R571 VTAIL.n369 VTAIL.n368 9.3005
R572 VTAIL.n367 VTAIL.n366 9.3005
R573 VTAIL.n322 VTAIL.n321 9.3005
R574 VTAIL.n361 VTAIL.n360 9.3005
R575 VTAIL.n274 VTAIL.n273 9.3005
R576 VTAIL.n281 VTAIL.n280 9.3005
R577 VTAIL.n283 VTAIL.n282 9.3005
R578 VTAIL.n270 VTAIL.n269 9.3005
R579 VTAIL.n289 VTAIL.n288 9.3005
R580 VTAIL.n291 VTAIL.n290 9.3005
R581 VTAIL.n265 VTAIL.n263 9.3005
R582 VTAIL.n297 VTAIL.n296 9.3005
R583 VTAIL.n313 VTAIL.n312 9.3005
R584 VTAIL.n256 VTAIL.n255 9.3005
R585 VTAIL.n307 VTAIL.n306 9.3005
R586 VTAIL.n305 VTAIL.n304 9.3005
R587 VTAIL.n260 VTAIL.n259 9.3005
R588 VTAIL.n299 VTAIL.n298 9.3005
R589 VTAIL.n210 VTAIL.n209 9.3005
R590 VTAIL.n217 VTAIL.n216 9.3005
R591 VTAIL.n219 VTAIL.n218 9.3005
R592 VTAIL.n206 VTAIL.n205 9.3005
R593 VTAIL.n225 VTAIL.n224 9.3005
R594 VTAIL.n227 VTAIL.n226 9.3005
R595 VTAIL.n201 VTAIL.n199 9.3005
R596 VTAIL.n233 VTAIL.n232 9.3005
R597 VTAIL.n249 VTAIL.n248 9.3005
R598 VTAIL.n192 VTAIL.n191 9.3005
R599 VTAIL.n243 VTAIL.n242 9.3005
R600 VTAIL.n241 VTAIL.n240 9.3005
R601 VTAIL.n196 VTAIL.n195 9.3005
R602 VTAIL.n235 VTAIL.n234 9.3005
R603 VTAIL.n469 VTAIL.n458 8.92171
R604 VTAIL.n500 VTAIL.n442 8.92171
R605 VTAIL.n29 VTAIL.n18 8.92171
R606 VTAIL.n60 VTAIL.n2 8.92171
R607 VTAIL.n91 VTAIL.n80 8.92171
R608 VTAIL.n122 VTAIL.n64 8.92171
R609 VTAIL.n155 VTAIL.n144 8.92171
R610 VTAIL.n186 VTAIL.n128 8.92171
R611 VTAIL.n438 VTAIL.n380 8.92171
R612 VTAIL.n409 VTAIL.n398 8.92171
R613 VTAIL.n374 VTAIL.n316 8.92171
R614 VTAIL.n345 VTAIL.n334 8.92171
R615 VTAIL.n312 VTAIL.n254 8.92171
R616 VTAIL.n283 VTAIL.n272 8.92171
R617 VTAIL.n248 VTAIL.n190 8.92171
R618 VTAIL.n219 VTAIL.n208 8.92171
R619 VTAIL.n466 VTAIL.n465 8.14595
R620 VTAIL.n26 VTAIL.n25 8.14595
R621 VTAIL.n88 VTAIL.n87 8.14595
R622 VTAIL.n152 VTAIL.n151 8.14595
R623 VTAIL.n406 VTAIL.n405 8.14595
R624 VTAIL.n342 VTAIL.n341 8.14595
R625 VTAIL.n280 VTAIL.n279 8.14595
R626 VTAIL.n216 VTAIL.n215 8.14595
R627 VTAIL.n462 VTAIL.n460 7.3702
R628 VTAIL.n22 VTAIL.n20 7.3702
R629 VTAIL.n84 VTAIL.n82 7.3702
R630 VTAIL.n148 VTAIL.n146 7.3702
R631 VTAIL.n402 VTAIL.n400 7.3702
R632 VTAIL.n338 VTAIL.n336 7.3702
R633 VTAIL.n276 VTAIL.n274 7.3702
R634 VTAIL.n212 VTAIL.n210 7.3702
R635 VTAIL.n465 VTAIL.n460 5.81868
R636 VTAIL.n25 VTAIL.n20 5.81868
R637 VTAIL.n87 VTAIL.n82 5.81868
R638 VTAIL.n151 VTAIL.n146 5.81868
R639 VTAIL.n405 VTAIL.n400 5.81868
R640 VTAIL.n341 VTAIL.n336 5.81868
R641 VTAIL.n279 VTAIL.n274 5.81868
R642 VTAIL.n215 VTAIL.n210 5.81868
R643 VTAIL.n466 VTAIL.n458 5.04292
R644 VTAIL.n502 VTAIL.n442 5.04292
R645 VTAIL.n26 VTAIL.n18 5.04292
R646 VTAIL.n62 VTAIL.n2 5.04292
R647 VTAIL.n88 VTAIL.n80 5.04292
R648 VTAIL.n124 VTAIL.n64 5.04292
R649 VTAIL.n152 VTAIL.n144 5.04292
R650 VTAIL.n188 VTAIL.n128 5.04292
R651 VTAIL.n440 VTAIL.n380 5.04292
R652 VTAIL.n406 VTAIL.n398 5.04292
R653 VTAIL.n376 VTAIL.n316 5.04292
R654 VTAIL.n342 VTAIL.n334 5.04292
R655 VTAIL.n314 VTAIL.n254 5.04292
R656 VTAIL.n280 VTAIL.n272 5.04292
R657 VTAIL.n250 VTAIL.n190 5.04292
R658 VTAIL.n216 VTAIL.n208 5.04292
R659 VTAIL.n470 VTAIL.n469 4.26717
R660 VTAIL.n500 VTAIL.n499 4.26717
R661 VTAIL.n30 VTAIL.n29 4.26717
R662 VTAIL.n60 VTAIL.n59 4.26717
R663 VTAIL.n92 VTAIL.n91 4.26717
R664 VTAIL.n122 VTAIL.n121 4.26717
R665 VTAIL.n156 VTAIL.n155 4.26717
R666 VTAIL.n186 VTAIL.n185 4.26717
R667 VTAIL.n438 VTAIL.n437 4.26717
R668 VTAIL.n410 VTAIL.n409 4.26717
R669 VTAIL.n374 VTAIL.n373 4.26717
R670 VTAIL.n346 VTAIL.n345 4.26717
R671 VTAIL.n312 VTAIL.n311 4.26717
R672 VTAIL.n284 VTAIL.n283 4.26717
R673 VTAIL.n248 VTAIL.n247 4.26717
R674 VTAIL.n220 VTAIL.n219 4.26717
R675 VTAIL.n473 VTAIL.n456 3.49141
R676 VTAIL.n496 VTAIL.n444 3.49141
R677 VTAIL.n33 VTAIL.n16 3.49141
R678 VTAIL.n56 VTAIL.n4 3.49141
R679 VTAIL.n95 VTAIL.n78 3.49141
R680 VTAIL.n118 VTAIL.n66 3.49141
R681 VTAIL.n159 VTAIL.n142 3.49141
R682 VTAIL.n182 VTAIL.n130 3.49141
R683 VTAIL.n434 VTAIL.n382 3.49141
R684 VTAIL.n413 VTAIL.n396 3.49141
R685 VTAIL.n370 VTAIL.n318 3.49141
R686 VTAIL.n349 VTAIL.n332 3.49141
R687 VTAIL.n308 VTAIL.n256 3.49141
R688 VTAIL.n287 VTAIL.n270 3.49141
R689 VTAIL.n244 VTAIL.n192 3.49141
R690 VTAIL.n223 VTAIL.n206 3.49141
R691 VTAIL.n253 VTAIL.n251 2.85395
R692 VTAIL.n315 VTAIL.n253 2.85395
R693 VTAIL.n379 VTAIL.n377 2.85395
R694 VTAIL.n441 VTAIL.n379 2.85395
R695 VTAIL.n189 VTAIL.n127 2.85395
R696 VTAIL.n127 VTAIL.n125 2.85395
R697 VTAIL.n63 VTAIL.n1 2.85395
R698 VTAIL.n461 VTAIL.n459 2.84303
R699 VTAIL.n21 VTAIL.n19 2.84303
R700 VTAIL.n83 VTAIL.n81 2.84303
R701 VTAIL.n147 VTAIL.n145 2.84303
R702 VTAIL.n401 VTAIL.n399 2.84303
R703 VTAIL.n337 VTAIL.n335 2.84303
R704 VTAIL.n275 VTAIL.n273 2.84303
R705 VTAIL.n211 VTAIL.n209 2.84303
R706 VTAIL VTAIL.n503 2.79576
R707 VTAIL.n474 VTAIL.n454 2.71565
R708 VTAIL.n495 VTAIL.n446 2.71565
R709 VTAIL.n34 VTAIL.n14 2.71565
R710 VTAIL.n55 VTAIL.n6 2.71565
R711 VTAIL.n96 VTAIL.n76 2.71565
R712 VTAIL.n117 VTAIL.n68 2.71565
R713 VTAIL.n160 VTAIL.n140 2.71565
R714 VTAIL.n181 VTAIL.n132 2.71565
R715 VTAIL.n433 VTAIL.n384 2.71565
R716 VTAIL.n414 VTAIL.n394 2.71565
R717 VTAIL.n369 VTAIL.n320 2.71565
R718 VTAIL.n350 VTAIL.n330 2.71565
R719 VTAIL.n307 VTAIL.n258 2.71565
R720 VTAIL.n288 VTAIL.n268 2.71565
R721 VTAIL.n243 VTAIL.n194 2.71565
R722 VTAIL.n224 VTAIL.n204 2.71565
R723 VTAIL.n479 VTAIL.n477 1.93989
R724 VTAIL.n492 VTAIL.n491 1.93989
R725 VTAIL.n39 VTAIL.n37 1.93989
R726 VTAIL.n52 VTAIL.n51 1.93989
R727 VTAIL.n101 VTAIL.n99 1.93989
R728 VTAIL.n114 VTAIL.n113 1.93989
R729 VTAIL.n165 VTAIL.n163 1.93989
R730 VTAIL.n178 VTAIL.n177 1.93989
R731 VTAIL.n430 VTAIL.n429 1.93989
R732 VTAIL.n418 VTAIL.n417 1.93989
R733 VTAIL.n366 VTAIL.n365 1.93989
R734 VTAIL.n354 VTAIL.n353 1.93989
R735 VTAIL.n304 VTAIL.n303 1.93989
R736 VTAIL.n292 VTAIL.n291 1.93989
R737 VTAIL.n240 VTAIL.n239 1.93989
R738 VTAIL.n228 VTAIL.n227 1.93989
R739 VTAIL.n0 VTAIL.t4 1.74962
R740 VTAIL.n0 VTAIL.t7 1.74962
R741 VTAIL.n126 VTAIL.t12 1.74962
R742 VTAIL.n126 VTAIL.t9 1.74962
R743 VTAIL.n378 VTAIL.t8 1.74962
R744 VTAIL.n378 VTAIL.t15 1.74962
R745 VTAIL.n252 VTAIL.t3 1.74962
R746 VTAIL.n252 VTAIL.t5 1.74962
R747 VTAIL.n478 VTAIL.n452 1.16414
R748 VTAIL.n488 VTAIL.n448 1.16414
R749 VTAIL.n38 VTAIL.n12 1.16414
R750 VTAIL.n48 VTAIL.n8 1.16414
R751 VTAIL.n100 VTAIL.n74 1.16414
R752 VTAIL.n110 VTAIL.n70 1.16414
R753 VTAIL.n164 VTAIL.n138 1.16414
R754 VTAIL.n174 VTAIL.n134 1.16414
R755 VTAIL.n426 VTAIL.n386 1.16414
R756 VTAIL.n421 VTAIL.n391 1.16414
R757 VTAIL.n362 VTAIL.n322 1.16414
R758 VTAIL.n357 VTAIL.n327 1.16414
R759 VTAIL.n300 VTAIL.n260 1.16414
R760 VTAIL.n295 VTAIL.n265 1.16414
R761 VTAIL.n236 VTAIL.n196 1.16414
R762 VTAIL.n231 VTAIL.n201 1.16414
R763 VTAIL.n377 VTAIL.n315 0.470328
R764 VTAIL.n125 VTAIL.n63 0.470328
R765 VTAIL.n484 VTAIL.n483 0.388379
R766 VTAIL.n487 VTAIL.n450 0.388379
R767 VTAIL.n44 VTAIL.n43 0.388379
R768 VTAIL.n47 VTAIL.n10 0.388379
R769 VTAIL.n106 VTAIL.n105 0.388379
R770 VTAIL.n109 VTAIL.n72 0.388379
R771 VTAIL.n170 VTAIL.n169 0.388379
R772 VTAIL.n173 VTAIL.n136 0.388379
R773 VTAIL.n425 VTAIL.n388 0.388379
R774 VTAIL.n422 VTAIL.n390 0.388379
R775 VTAIL.n361 VTAIL.n324 0.388379
R776 VTAIL.n358 VTAIL.n326 0.388379
R777 VTAIL.n299 VTAIL.n262 0.388379
R778 VTAIL.n296 VTAIL.n264 0.388379
R779 VTAIL.n235 VTAIL.n198 0.388379
R780 VTAIL.n232 VTAIL.n200 0.388379
R781 VTAIL.n467 VTAIL.n459 0.155672
R782 VTAIL.n468 VTAIL.n467 0.155672
R783 VTAIL.n468 VTAIL.n455 0.155672
R784 VTAIL.n475 VTAIL.n455 0.155672
R785 VTAIL.n476 VTAIL.n475 0.155672
R786 VTAIL.n476 VTAIL.n451 0.155672
R787 VTAIL.n485 VTAIL.n451 0.155672
R788 VTAIL.n486 VTAIL.n485 0.155672
R789 VTAIL.n486 VTAIL.n447 0.155672
R790 VTAIL.n493 VTAIL.n447 0.155672
R791 VTAIL.n494 VTAIL.n493 0.155672
R792 VTAIL.n494 VTAIL.n443 0.155672
R793 VTAIL.n501 VTAIL.n443 0.155672
R794 VTAIL.n27 VTAIL.n19 0.155672
R795 VTAIL.n28 VTAIL.n27 0.155672
R796 VTAIL.n28 VTAIL.n15 0.155672
R797 VTAIL.n35 VTAIL.n15 0.155672
R798 VTAIL.n36 VTAIL.n35 0.155672
R799 VTAIL.n36 VTAIL.n11 0.155672
R800 VTAIL.n45 VTAIL.n11 0.155672
R801 VTAIL.n46 VTAIL.n45 0.155672
R802 VTAIL.n46 VTAIL.n7 0.155672
R803 VTAIL.n53 VTAIL.n7 0.155672
R804 VTAIL.n54 VTAIL.n53 0.155672
R805 VTAIL.n54 VTAIL.n3 0.155672
R806 VTAIL.n61 VTAIL.n3 0.155672
R807 VTAIL.n89 VTAIL.n81 0.155672
R808 VTAIL.n90 VTAIL.n89 0.155672
R809 VTAIL.n90 VTAIL.n77 0.155672
R810 VTAIL.n97 VTAIL.n77 0.155672
R811 VTAIL.n98 VTAIL.n97 0.155672
R812 VTAIL.n98 VTAIL.n73 0.155672
R813 VTAIL.n107 VTAIL.n73 0.155672
R814 VTAIL.n108 VTAIL.n107 0.155672
R815 VTAIL.n108 VTAIL.n69 0.155672
R816 VTAIL.n115 VTAIL.n69 0.155672
R817 VTAIL.n116 VTAIL.n115 0.155672
R818 VTAIL.n116 VTAIL.n65 0.155672
R819 VTAIL.n123 VTAIL.n65 0.155672
R820 VTAIL.n153 VTAIL.n145 0.155672
R821 VTAIL.n154 VTAIL.n153 0.155672
R822 VTAIL.n154 VTAIL.n141 0.155672
R823 VTAIL.n161 VTAIL.n141 0.155672
R824 VTAIL.n162 VTAIL.n161 0.155672
R825 VTAIL.n162 VTAIL.n137 0.155672
R826 VTAIL.n171 VTAIL.n137 0.155672
R827 VTAIL.n172 VTAIL.n171 0.155672
R828 VTAIL.n172 VTAIL.n133 0.155672
R829 VTAIL.n179 VTAIL.n133 0.155672
R830 VTAIL.n180 VTAIL.n179 0.155672
R831 VTAIL.n180 VTAIL.n129 0.155672
R832 VTAIL.n187 VTAIL.n129 0.155672
R833 VTAIL.n439 VTAIL.n381 0.155672
R834 VTAIL.n432 VTAIL.n381 0.155672
R835 VTAIL.n432 VTAIL.n431 0.155672
R836 VTAIL.n431 VTAIL.n385 0.155672
R837 VTAIL.n424 VTAIL.n385 0.155672
R838 VTAIL.n424 VTAIL.n423 0.155672
R839 VTAIL.n423 VTAIL.n389 0.155672
R840 VTAIL.n416 VTAIL.n389 0.155672
R841 VTAIL.n416 VTAIL.n415 0.155672
R842 VTAIL.n415 VTAIL.n395 0.155672
R843 VTAIL.n408 VTAIL.n395 0.155672
R844 VTAIL.n408 VTAIL.n407 0.155672
R845 VTAIL.n407 VTAIL.n399 0.155672
R846 VTAIL.n375 VTAIL.n317 0.155672
R847 VTAIL.n368 VTAIL.n317 0.155672
R848 VTAIL.n368 VTAIL.n367 0.155672
R849 VTAIL.n367 VTAIL.n321 0.155672
R850 VTAIL.n360 VTAIL.n321 0.155672
R851 VTAIL.n360 VTAIL.n359 0.155672
R852 VTAIL.n359 VTAIL.n325 0.155672
R853 VTAIL.n352 VTAIL.n325 0.155672
R854 VTAIL.n352 VTAIL.n351 0.155672
R855 VTAIL.n351 VTAIL.n331 0.155672
R856 VTAIL.n344 VTAIL.n331 0.155672
R857 VTAIL.n344 VTAIL.n343 0.155672
R858 VTAIL.n343 VTAIL.n335 0.155672
R859 VTAIL.n313 VTAIL.n255 0.155672
R860 VTAIL.n306 VTAIL.n255 0.155672
R861 VTAIL.n306 VTAIL.n305 0.155672
R862 VTAIL.n305 VTAIL.n259 0.155672
R863 VTAIL.n298 VTAIL.n259 0.155672
R864 VTAIL.n298 VTAIL.n297 0.155672
R865 VTAIL.n297 VTAIL.n263 0.155672
R866 VTAIL.n290 VTAIL.n263 0.155672
R867 VTAIL.n290 VTAIL.n289 0.155672
R868 VTAIL.n289 VTAIL.n269 0.155672
R869 VTAIL.n282 VTAIL.n269 0.155672
R870 VTAIL.n282 VTAIL.n281 0.155672
R871 VTAIL.n281 VTAIL.n273 0.155672
R872 VTAIL.n249 VTAIL.n191 0.155672
R873 VTAIL.n242 VTAIL.n191 0.155672
R874 VTAIL.n242 VTAIL.n241 0.155672
R875 VTAIL.n241 VTAIL.n195 0.155672
R876 VTAIL.n234 VTAIL.n195 0.155672
R877 VTAIL.n234 VTAIL.n233 0.155672
R878 VTAIL.n233 VTAIL.n199 0.155672
R879 VTAIL.n226 VTAIL.n199 0.155672
R880 VTAIL.n226 VTAIL.n225 0.155672
R881 VTAIL.n225 VTAIL.n205 0.155672
R882 VTAIL.n218 VTAIL.n205 0.155672
R883 VTAIL.n218 VTAIL.n217 0.155672
R884 VTAIL.n217 VTAIL.n209 0.155672
R885 VTAIL VTAIL.n1 0.0586897
R886 VDD1 VDD1.n0 62.0233
R887 VDD1.n3 VDD1.n2 61.9096
R888 VDD1.n3 VDD1.n1 61.9096
R889 VDD1.n5 VDD1.n4 60.5382
R890 VDD1.n5 VDD1.n3 46.8974
R891 VDD1.n4 VDD1.t0 1.74962
R892 VDD1.n4 VDD1.t3 1.74962
R893 VDD1.n0 VDD1.t5 1.74962
R894 VDD1.n0 VDD1.t7 1.74962
R895 VDD1.n2 VDD1.t1 1.74962
R896 VDD1.n2 VDD1.t4 1.74962
R897 VDD1.n1 VDD1.t2 1.74962
R898 VDD1.n1 VDD1.t6 1.74962
R899 VDD1 VDD1.n5 1.36903
R900 B.n909 B.n908 585
R901 B.n910 B.n909 585
R902 B.n328 B.n149 585
R903 B.n327 B.n326 585
R904 B.n325 B.n324 585
R905 B.n323 B.n322 585
R906 B.n321 B.n320 585
R907 B.n319 B.n318 585
R908 B.n317 B.n316 585
R909 B.n315 B.n314 585
R910 B.n313 B.n312 585
R911 B.n311 B.n310 585
R912 B.n309 B.n308 585
R913 B.n307 B.n306 585
R914 B.n305 B.n304 585
R915 B.n303 B.n302 585
R916 B.n301 B.n300 585
R917 B.n299 B.n298 585
R918 B.n297 B.n296 585
R919 B.n295 B.n294 585
R920 B.n293 B.n292 585
R921 B.n291 B.n290 585
R922 B.n289 B.n288 585
R923 B.n287 B.n286 585
R924 B.n285 B.n284 585
R925 B.n283 B.n282 585
R926 B.n281 B.n280 585
R927 B.n279 B.n278 585
R928 B.n277 B.n276 585
R929 B.n275 B.n274 585
R930 B.n273 B.n272 585
R931 B.n271 B.n270 585
R932 B.n269 B.n268 585
R933 B.n267 B.n266 585
R934 B.n265 B.n264 585
R935 B.n263 B.n262 585
R936 B.n261 B.n260 585
R937 B.n259 B.n258 585
R938 B.n257 B.n256 585
R939 B.n255 B.n254 585
R940 B.n253 B.n252 585
R941 B.n250 B.n249 585
R942 B.n248 B.n247 585
R943 B.n246 B.n245 585
R944 B.n244 B.n243 585
R945 B.n242 B.n241 585
R946 B.n240 B.n239 585
R947 B.n238 B.n237 585
R948 B.n236 B.n235 585
R949 B.n234 B.n233 585
R950 B.n232 B.n231 585
R951 B.n230 B.n229 585
R952 B.n228 B.n227 585
R953 B.n226 B.n225 585
R954 B.n224 B.n223 585
R955 B.n222 B.n221 585
R956 B.n220 B.n219 585
R957 B.n218 B.n217 585
R958 B.n216 B.n215 585
R959 B.n214 B.n213 585
R960 B.n212 B.n211 585
R961 B.n210 B.n209 585
R962 B.n208 B.n207 585
R963 B.n206 B.n205 585
R964 B.n204 B.n203 585
R965 B.n202 B.n201 585
R966 B.n200 B.n199 585
R967 B.n198 B.n197 585
R968 B.n196 B.n195 585
R969 B.n194 B.n193 585
R970 B.n192 B.n191 585
R971 B.n190 B.n189 585
R972 B.n188 B.n187 585
R973 B.n186 B.n185 585
R974 B.n184 B.n183 585
R975 B.n182 B.n181 585
R976 B.n180 B.n179 585
R977 B.n178 B.n177 585
R978 B.n176 B.n175 585
R979 B.n174 B.n173 585
R980 B.n172 B.n171 585
R981 B.n170 B.n169 585
R982 B.n168 B.n167 585
R983 B.n166 B.n165 585
R984 B.n164 B.n163 585
R985 B.n162 B.n161 585
R986 B.n160 B.n159 585
R987 B.n158 B.n157 585
R988 B.n156 B.n155 585
R989 B.n103 B.n102 585
R990 B.n907 B.n104 585
R991 B.n911 B.n104 585
R992 B.n906 B.n905 585
R993 B.n905 B.n100 585
R994 B.n904 B.n99 585
R995 B.n917 B.n99 585
R996 B.n903 B.n98 585
R997 B.n918 B.n98 585
R998 B.n902 B.n97 585
R999 B.n919 B.n97 585
R1000 B.n901 B.n900 585
R1001 B.n900 B.n93 585
R1002 B.n899 B.n92 585
R1003 B.n925 B.n92 585
R1004 B.n898 B.n91 585
R1005 B.n926 B.n91 585
R1006 B.n897 B.n90 585
R1007 B.n927 B.n90 585
R1008 B.n896 B.n895 585
R1009 B.n895 B.n86 585
R1010 B.n894 B.n85 585
R1011 B.n933 B.n85 585
R1012 B.n893 B.n84 585
R1013 B.n934 B.n84 585
R1014 B.n892 B.n83 585
R1015 B.n935 B.n83 585
R1016 B.n891 B.n890 585
R1017 B.n890 B.n79 585
R1018 B.n889 B.n78 585
R1019 B.n941 B.n78 585
R1020 B.n888 B.n77 585
R1021 B.n942 B.n77 585
R1022 B.n887 B.n76 585
R1023 B.n943 B.n76 585
R1024 B.n886 B.n885 585
R1025 B.n885 B.n72 585
R1026 B.n884 B.n71 585
R1027 B.n949 B.n71 585
R1028 B.n883 B.n70 585
R1029 B.n950 B.n70 585
R1030 B.n882 B.n69 585
R1031 B.n951 B.n69 585
R1032 B.n881 B.n880 585
R1033 B.n880 B.n65 585
R1034 B.n879 B.n64 585
R1035 B.n957 B.n64 585
R1036 B.n878 B.n63 585
R1037 B.n958 B.n63 585
R1038 B.n877 B.n62 585
R1039 B.n959 B.n62 585
R1040 B.n876 B.n875 585
R1041 B.n875 B.n58 585
R1042 B.n874 B.n57 585
R1043 B.n965 B.n57 585
R1044 B.n873 B.n56 585
R1045 B.n966 B.n56 585
R1046 B.n872 B.n55 585
R1047 B.n967 B.n55 585
R1048 B.n871 B.n870 585
R1049 B.n870 B.n51 585
R1050 B.n869 B.n50 585
R1051 B.n973 B.n50 585
R1052 B.n868 B.n49 585
R1053 B.n974 B.n49 585
R1054 B.n867 B.n48 585
R1055 B.n975 B.n48 585
R1056 B.n866 B.n865 585
R1057 B.n865 B.n44 585
R1058 B.n864 B.n43 585
R1059 B.n981 B.n43 585
R1060 B.n863 B.n42 585
R1061 B.n982 B.n42 585
R1062 B.n862 B.n41 585
R1063 B.n983 B.n41 585
R1064 B.n861 B.n860 585
R1065 B.n860 B.n37 585
R1066 B.n859 B.n36 585
R1067 B.n989 B.n36 585
R1068 B.n858 B.n35 585
R1069 B.n990 B.n35 585
R1070 B.n857 B.n34 585
R1071 B.n991 B.n34 585
R1072 B.n856 B.n855 585
R1073 B.n855 B.n30 585
R1074 B.n854 B.n29 585
R1075 B.n997 B.n29 585
R1076 B.n853 B.n28 585
R1077 B.n998 B.n28 585
R1078 B.n852 B.n27 585
R1079 B.n999 B.n27 585
R1080 B.n851 B.n850 585
R1081 B.n850 B.n23 585
R1082 B.n849 B.n22 585
R1083 B.n1005 B.n22 585
R1084 B.n848 B.n21 585
R1085 B.n1006 B.n21 585
R1086 B.n847 B.n20 585
R1087 B.n1007 B.n20 585
R1088 B.n846 B.n845 585
R1089 B.n845 B.n16 585
R1090 B.n844 B.n15 585
R1091 B.n1013 B.n15 585
R1092 B.n843 B.n14 585
R1093 B.n1014 B.n14 585
R1094 B.n842 B.n13 585
R1095 B.n1015 B.n13 585
R1096 B.n841 B.n840 585
R1097 B.n840 B.n12 585
R1098 B.n839 B.n838 585
R1099 B.n839 B.n8 585
R1100 B.n837 B.n7 585
R1101 B.n1022 B.n7 585
R1102 B.n836 B.n6 585
R1103 B.n1023 B.n6 585
R1104 B.n835 B.n5 585
R1105 B.n1024 B.n5 585
R1106 B.n834 B.n833 585
R1107 B.n833 B.n4 585
R1108 B.n832 B.n329 585
R1109 B.n832 B.n831 585
R1110 B.n822 B.n330 585
R1111 B.n331 B.n330 585
R1112 B.n824 B.n823 585
R1113 B.n825 B.n824 585
R1114 B.n821 B.n336 585
R1115 B.n336 B.n335 585
R1116 B.n820 B.n819 585
R1117 B.n819 B.n818 585
R1118 B.n338 B.n337 585
R1119 B.n339 B.n338 585
R1120 B.n811 B.n810 585
R1121 B.n812 B.n811 585
R1122 B.n809 B.n344 585
R1123 B.n344 B.n343 585
R1124 B.n808 B.n807 585
R1125 B.n807 B.n806 585
R1126 B.n346 B.n345 585
R1127 B.n347 B.n346 585
R1128 B.n799 B.n798 585
R1129 B.n800 B.n799 585
R1130 B.n797 B.n352 585
R1131 B.n352 B.n351 585
R1132 B.n796 B.n795 585
R1133 B.n795 B.n794 585
R1134 B.n354 B.n353 585
R1135 B.n355 B.n354 585
R1136 B.n787 B.n786 585
R1137 B.n788 B.n787 585
R1138 B.n785 B.n360 585
R1139 B.n360 B.n359 585
R1140 B.n784 B.n783 585
R1141 B.n783 B.n782 585
R1142 B.n362 B.n361 585
R1143 B.n363 B.n362 585
R1144 B.n775 B.n774 585
R1145 B.n776 B.n775 585
R1146 B.n773 B.n368 585
R1147 B.n368 B.n367 585
R1148 B.n772 B.n771 585
R1149 B.n771 B.n770 585
R1150 B.n370 B.n369 585
R1151 B.n371 B.n370 585
R1152 B.n763 B.n762 585
R1153 B.n764 B.n763 585
R1154 B.n761 B.n376 585
R1155 B.n376 B.n375 585
R1156 B.n760 B.n759 585
R1157 B.n759 B.n758 585
R1158 B.n378 B.n377 585
R1159 B.n379 B.n378 585
R1160 B.n751 B.n750 585
R1161 B.n752 B.n751 585
R1162 B.n749 B.n384 585
R1163 B.n384 B.n383 585
R1164 B.n748 B.n747 585
R1165 B.n747 B.n746 585
R1166 B.n386 B.n385 585
R1167 B.n387 B.n386 585
R1168 B.n739 B.n738 585
R1169 B.n740 B.n739 585
R1170 B.n737 B.n392 585
R1171 B.n392 B.n391 585
R1172 B.n736 B.n735 585
R1173 B.n735 B.n734 585
R1174 B.n394 B.n393 585
R1175 B.n395 B.n394 585
R1176 B.n727 B.n726 585
R1177 B.n728 B.n727 585
R1178 B.n725 B.n400 585
R1179 B.n400 B.n399 585
R1180 B.n724 B.n723 585
R1181 B.n723 B.n722 585
R1182 B.n402 B.n401 585
R1183 B.n403 B.n402 585
R1184 B.n715 B.n714 585
R1185 B.n716 B.n715 585
R1186 B.n713 B.n408 585
R1187 B.n408 B.n407 585
R1188 B.n712 B.n711 585
R1189 B.n711 B.n710 585
R1190 B.n410 B.n409 585
R1191 B.n411 B.n410 585
R1192 B.n703 B.n702 585
R1193 B.n704 B.n703 585
R1194 B.n701 B.n416 585
R1195 B.n416 B.n415 585
R1196 B.n700 B.n699 585
R1197 B.n699 B.n698 585
R1198 B.n418 B.n417 585
R1199 B.n419 B.n418 585
R1200 B.n691 B.n690 585
R1201 B.n692 B.n691 585
R1202 B.n689 B.n423 585
R1203 B.n427 B.n423 585
R1204 B.n688 B.n687 585
R1205 B.n687 B.n686 585
R1206 B.n425 B.n424 585
R1207 B.n426 B.n425 585
R1208 B.n679 B.n678 585
R1209 B.n680 B.n679 585
R1210 B.n677 B.n432 585
R1211 B.n432 B.n431 585
R1212 B.n676 B.n675 585
R1213 B.n675 B.n674 585
R1214 B.n434 B.n433 585
R1215 B.n435 B.n434 585
R1216 B.n667 B.n666 585
R1217 B.n668 B.n667 585
R1218 B.n438 B.n437 585
R1219 B.n490 B.n488 585
R1220 B.n491 B.n487 585
R1221 B.n491 B.n439 585
R1222 B.n494 B.n493 585
R1223 B.n495 B.n486 585
R1224 B.n497 B.n496 585
R1225 B.n499 B.n485 585
R1226 B.n502 B.n501 585
R1227 B.n503 B.n484 585
R1228 B.n505 B.n504 585
R1229 B.n507 B.n483 585
R1230 B.n510 B.n509 585
R1231 B.n511 B.n482 585
R1232 B.n513 B.n512 585
R1233 B.n515 B.n481 585
R1234 B.n518 B.n517 585
R1235 B.n519 B.n480 585
R1236 B.n521 B.n520 585
R1237 B.n523 B.n479 585
R1238 B.n526 B.n525 585
R1239 B.n527 B.n478 585
R1240 B.n529 B.n528 585
R1241 B.n531 B.n477 585
R1242 B.n534 B.n533 585
R1243 B.n535 B.n476 585
R1244 B.n537 B.n536 585
R1245 B.n539 B.n475 585
R1246 B.n542 B.n541 585
R1247 B.n543 B.n474 585
R1248 B.n545 B.n544 585
R1249 B.n547 B.n473 585
R1250 B.n550 B.n549 585
R1251 B.n551 B.n472 585
R1252 B.n553 B.n552 585
R1253 B.n555 B.n471 585
R1254 B.n558 B.n557 585
R1255 B.n559 B.n470 585
R1256 B.n561 B.n560 585
R1257 B.n563 B.n469 585
R1258 B.n566 B.n565 585
R1259 B.n568 B.n466 585
R1260 B.n570 B.n569 585
R1261 B.n572 B.n465 585
R1262 B.n575 B.n574 585
R1263 B.n576 B.n464 585
R1264 B.n578 B.n577 585
R1265 B.n580 B.n463 585
R1266 B.n583 B.n582 585
R1267 B.n584 B.n460 585
R1268 B.n587 B.n586 585
R1269 B.n589 B.n459 585
R1270 B.n592 B.n591 585
R1271 B.n593 B.n458 585
R1272 B.n595 B.n594 585
R1273 B.n597 B.n457 585
R1274 B.n600 B.n599 585
R1275 B.n601 B.n456 585
R1276 B.n603 B.n602 585
R1277 B.n605 B.n455 585
R1278 B.n608 B.n607 585
R1279 B.n609 B.n454 585
R1280 B.n611 B.n610 585
R1281 B.n613 B.n453 585
R1282 B.n616 B.n615 585
R1283 B.n617 B.n452 585
R1284 B.n619 B.n618 585
R1285 B.n621 B.n451 585
R1286 B.n624 B.n623 585
R1287 B.n625 B.n450 585
R1288 B.n627 B.n626 585
R1289 B.n629 B.n449 585
R1290 B.n632 B.n631 585
R1291 B.n633 B.n448 585
R1292 B.n635 B.n634 585
R1293 B.n637 B.n447 585
R1294 B.n640 B.n639 585
R1295 B.n641 B.n446 585
R1296 B.n643 B.n642 585
R1297 B.n645 B.n445 585
R1298 B.n648 B.n647 585
R1299 B.n649 B.n444 585
R1300 B.n651 B.n650 585
R1301 B.n653 B.n443 585
R1302 B.n656 B.n655 585
R1303 B.n657 B.n442 585
R1304 B.n659 B.n658 585
R1305 B.n661 B.n441 585
R1306 B.n664 B.n663 585
R1307 B.n665 B.n440 585
R1308 B.n670 B.n669 585
R1309 B.n669 B.n668 585
R1310 B.n671 B.n436 585
R1311 B.n436 B.n435 585
R1312 B.n673 B.n672 585
R1313 B.n674 B.n673 585
R1314 B.n430 B.n429 585
R1315 B.n431 B.n430 585
R1316 B.n682 B.n681 585
R1317 B.n681 B.n680 585
R1318 B.n683 B.n428 585
R1319 B.n428 B.n426 585
R1320 B.n685 B.n684 585
R1321 B.n686 B.n685 585
R1322 B.n422 B.n421 585
R1323 B.n427 B.n422 585
R1324 B.n694 B.n693 585
R1325 B.n693 B.n692 585
R1326 B.n695 B.n420 585
R1327 B.n420 B.n419 585
R1328 B.n697 B.n696 585
R1329 B.n698 B.n697 585
R1330 B.n414 B.n413 585
R1331 B.n415 B.n414 585
R1332 B.n706 B.n705 585
R1333 B.n705 B.n704 585
R1334 B.n707 B.n412 585
R1335 B.n412 B.n411 585
R1336 B.n709 B.n708 585
R1337 B.n710 B.n709 585
R1338 B.n406 B.n405 585
R1339 B.n407 B.n406 585
R1340 B.n718 B.n717 585
R1341 B.n717 B.n716 585
R1342 B.n719 B.n404 585
R1343 B.n404 B.n403 585
R1344 B.n721 B.n720 585
R1345 B.n722 B.n721 585
R1346 B.n398 B.n397 585
R1347 B.n399 B.n398 585
R1348 B.n730 B.n729 585
R1349 B.n729 B.n728 585
R1350 B.n731 B.n396 585
R1351 B.n396 B.n395 585
R1352 B.n733 B.n732 585
R1353 B.n734 B.n733 585
R1354 B.n390 B.n389 585
R1355 B.n391 B.n390 585
R1356 B.n742 B.n741 585
R1357 B.n741 B.n740 585
R1358 B.n743 B.n388 585
R1359 B.n388 B.n387 585
R1360 B.n745 B.n744 585
R1361 B.n746 B.n745 585
R1362 B.n382 B.n381 585
R1363 B.n383 B.n382 585
R1364 B.n754 B.n753 585
R1365 B.n753 B.n752 585
R1366 B.n755 B.n380 585
R1367 B.n380 B.n379 585
R1368 B.n757 B.n756 585
R1369 B.n758 B.n757 585
R1370 B.n374 B.n373 585
R1371 B.n375 B.n374 585
R1372 B.n766 B.n765 585
R1373 B.n765 B.n764 585
R1374 B.n767 B.n372 585
R1375 B.n372 B.n371 585
R1376 B.n769 B.n768 585
R1377 B.n770 B.n769 585
R1378 B.n366 B.n365 585
R1379 B.n367 B.n366 585
R1380 B.n778 B.n777 585
R1381 B.n777 B.n776 585
R1382 B.n779 B.n364 585
R1383 B.n364 B.n363 585
R1384 B.n781 B.n780 585
R1385 B.n782 B.n781 585
R1386 B.n358 B.n357 585
R1387 B.n359 B.n358 585
R1388 B.n790 B.n789 585
R1389 B.n789 B.n788 585
R1390 B.n791 B.n356 585
R1391 B.n356 B.n355 585
R1392 B.n793 B.n792 585
R1393 B.n794 B.n793 585
R1394 B.n350 B.n349 585
R1395 B.n351 B.n350 585
R1396 B.n802 B.n801 585
R1397 B.n801 B.n800 585
R1398 B.n803 B.n348 585
R1399 B.n348 B.n347 585
R1400 B.n805 B.n804 585
R1401 B.n806 B.n805 585
R1402 B.n342 B.n341 585
R1403 B.n343 B.n342 585
R1404 B.n814 B.n813 585
R1405 B.n813 B.n812 585
R1406 B.n815 B.n340 585
R1407 B.n340 B.n339 585
R1408 B.n817 B.n816 585
R1409 B.n818 B.n817 585
R1410 B.n334 B.n333 585
R1411 B.n335 B.n334 585
R1412 B.n827 B.n826 585
R1413 B.n826 B.n825 585
R1414 B.n828 B.n332 585
R1415 B.n332 B.n331 585
R1416 B.n830 B.n829 585
R1417 B.n831 B.n830 585
R1418 B.n3 B.n0 585
R1419 B.n4 B.n3 585
R1420 B.n1021 B.n1 585
R1421 B.n1022 B.n1021 585
R1422 B.n1020 B.n1019 585
R1423 B.n1020 B.n8 585
R1424 B.n1018 B.n9 585
R1425 B.n12 B.n9 585
R1426 B.n1017 B.n1016 585
R1427 B.n1016 B.n1015 585
R1428 B.n11 B.n10 585
R1429 B.n1014 B.n11 585
R1430 B.n1012 B.n1011 585
R1431 B.n1013 B.n1012 585
R1432 B.n1010 B.n17 585
R1433 B.n17 B.n16 585
R1434 B.n1009 B.n1008 585
R1435 B.n1008 B.n1007 585
R1436 B.n19 B.n18 585
R1437 B.n1006 B.n19 585
R1438 B.n1004 B.n1003 585
R1439 B.n1005 B.n1004 585
R1440 B.n1002 B.n24 585
R1441 B.n24 B.n23 585
R1442 B.n1001 B.n1000 585
R1443 B.n1000 B.n999 585
R1444 B.n26 B.n25 585
R1445 B.n998 B.n26 585
R1446 B.n996 B.n995 585
R1447 B.n997 B.n996 585
R1448 B.n994 B.n31 585
R1449 B.n31 B.n30 585
R1450 B.n993 B.n992 585
R1451 B.n992 B.n991 585
R1452 B.n33 B.n32 585
R1453 B.n990 B.n33 585
R1454 B.n988 B.n987 585
R1455 B.n989 B.n988 585
R1456 B.n986 B.n38 585
R1457 B.n38 B.n37 585
R1458 B.n985 B.n984 585
R1459 B.n984 B.n983 585
R1460 B.n40 B.n39 585
R1461 B.n982 B.n40 585
R1462 B.n980 B.n979 585
R1463 B.n981 B.n980 585
R1464 B.n978 B.n45 585
R1465 B.n45 B.n44 585
R1466 B.n977 B.n976 585
R1467 B.n976 B.n975 585
R1468 B.n47 B.n46 585
R1469 B.n974 B.n47 585
R1470 B.n972 B.n971 585
R1471 B.n973 B.n972 585
R1472 B.n970 B.n52 585
R1473 B.n52 B.n51 585
R1474 B.n969 B.n968 585
R1475 B.n968 B.n967 585
R1476 B.n54 B.n53 585
R1477 B.n966 B.n54 585
R1478 B.n964 B.n963 585
R1479 B.n965 B.n964 585
R1480 B.n962 B.n59 585
R1481 B.n59 B.n58 585
R1482 B.n961 B.n960 585
R1483 B.n960 B.n959 585
R1484 B.n61 B.n60 585
R1485 B.n958 B.n61 585
R1486 B.n956 B.n955 585
R1487 B.n957 B.n956 585
R1488 B.n954 B.n66 585
R1489 B.n66 B.n65 585
R1490 B.n953 B.n952 585
R1491 B.n952 B.n951 585
R1492 B.n68 B.n67 585
R1493 B.n950 B.n68 585
R1494 B.n948 B.n947 585
R1495 B.n949 B.n948 585
R1496 B.n946 B.n73 585
R1497 B.n73 B.n72 585
R1498 B.n945 B.n944 585
R1499 B.n944 B.n943 585
R1500 B.n75 B.n74 585
R1501 B.n942 B.n75 585
R1502 B.n940 B.n939 585
R1503 B.n941 B.n940 585
R1504 B.n938 B.n80 585
R1505 B.n80 B.n79 585
R1506 B.n937 B.n936 585
R1507 B.n936 B.n935 585
R1508 B.n82 B.n81 585
R1509 B.n934 B.n82 585
R1510 B.n932 B.n931 585
R1511 B.n933 B.n932 585
R1512 B.n930 B.n87 585
R1513 B.n87 B.n86 585
R1514 B.n929 B.n928 585
R1515 B.n928 B.n927 585
R1516 B.n89 B.n88 585
R1517 B.n926 B.n89 585
R1518 B.n924 B.n923 585
R1519 B.n925 B.n924 585
R1520 B.n922 B.n94 585
R1521 B.n94 B.n93 585
R1522 B.n921 B.n920 585
R1523 B.n920 B.n919 585
R1524 B.n96 B.n95 585
R1525 B.n918 B.n96 585
R1526 B.n916 B.n915 585
R1527 B.n917 B.n916 585
R1528 B.n914 B.n101 585
R1529 B.n101 B.n100 585
R1530 B.n913 B.n912 585
R1531 B.n912 B.n911 585
R1532 B.n1025 B.n1024 585
R1533 B.n1023 B.n2 585
R1534 B.n912 B.n103 530.939
R1535 B.n909 B.n104 530.939
R1536 B.n667 B.n440 530.939
R1537 B.n669 B.n438 530.939
R1538 B.n150 B.t17 334.49
R1539 B.n461 B.t21 334.49
R1540 B.n152 B.t10 334.49
R1541 B.n467 B.t15 334.49
R1542 B.n152 B.t8 300.104
R1543 B.n150 B.t16 300.104
R1544 B.n461 B.t19 300.104
R1545 B.n467 B.t12 300.104
R1546 B.n151 B.t18 270.296
R1547 B.n462 B.t20 270.296
R1548 B.n153 B.t11 270.296
R1549 B.n468 B.t14 270.296
R1550 B.n910 B.n148 256.663
R1551 B.n910 B.n147 256.663
R1552 B.n910 B.n146 256.663
R1553 B.n910 B.n145 256.663
R1554 B.n910 B.n144 256.663
R1555 B.n910 B.n143 256.663
R1556 B.n910 B.n142 256.663
R1557 B.n910 B.n141 256.663
R1558 B.n910 B.n140 256.663
R1559 B.n910 B.n139 256.663
R1560 B.n910 B.n138 256.663
R1561 B.n910 B.n137 256.663
R1562 B.n910 B.n136 256.663
R1563 B.n910 B.n135 256.663
R1564 B.n910 B.n134 256.663
R1565 B.n910 B.n133 256.663
R1566 B.n910 B.n132 256.663
R1567 B.n910 B.n131 256.663
R1568 B.n910 B.n130 256.663
R1569 B.n910 B.n129 256.663
R1570 B.n910 B.n128 256.663
R1571 B.n910 B.n127 256.663
R1572 B.n910 B.n126 256.663
R1573 B.n910 B.n125 256.663
R1574 B.n910 B.n124 256.663
R1575 B.n910 B.n123 256.663
R1576 B.n910 B.n122 256.663
R1577 B.n910 B.n121 256.663
R1578 B.n910 B.n120 256.663
R1579 B.n910 B.n119 256.663
R1580 B.n910 B.n118 256.663
R1581 B.n910 B.n117 256.663
R1582 B.n910 B.n116 256.663
R1583 B.n910 B.n115 256.663
R1584 B.n910 B.n114 256.663
R1585 B.n910 B.n113 256.663
R1586 B.n910 B.n112 256.663
R1587 B.n910 B.n111 256.663
R1588 B.n910 B.n110 256.663
R1589 B.n910 B.n109 256.663
R1590 B.n910 B.n108 256.663
R1591 B.n910 B.n107 256.663
R1592 B.n910 B.n106 256.663
R1593 B.n910 B.n105 256.663
R1594 B.n489 B.n439 256.663
R1595 B.n492 B.n439 256.663
R1596 B.n498 B.n439 256.663
R1597 B.n500 B.n439 256.663
R1598 B.n506 B.n439 256.663
R1599 B.n508 B.n439 256.663
R1600 B.n514 B.n439 256.663
R1601 B.n516 B.n439 256.663
R1602 B.n522 B.n439 256.663
R1603 B.n524 B.n439 256.663
R1604 B.n530 B.n439 256.663
R1605 B.n532 B.n439 256.663
R1606 B.n538 B.n439 256.663
R1607 B.n540 B.n439 256.663
R1608 B.n546 B.n439 256.663
R1609 B.n548 B.n439 256.663
R1610 B.n554 B.n439 256.663
R1611 B.n556 B.n439 256.663
R1612 B.n562 B.n439 256.663
R1613 B.n564 B.n439 256.663
R1614 B.n571 B.n439 256.663
R1615 B.n573 B.n439 256.663
R1616 B.n579 B.n439 256.663
R1617 B.n581 B.n439 256.663
R1618 B.n588 B.n439 256.663
R1619 B.n590 B.n439 256.663
R1620 B.n596 B.n439 256.663
R1621 B.n598 B.n439 256.663
R1622 B.n604 B.n439 256.663
R1623 B.n606 B.n439 256.663
R1624 B.n612 B.n439 256.663
R1625 B.n614 B.n439 256.663
R1626 B.n620 B.n439 256.663
R1627 B.n622 B.n439 256.663
R1628 B.n628 B.n439 256.663
R1629 B.n630 B.n439 256.663
R1630 B.n636 B.n439 256.663
R1631 B.n638 B.n439 256.663
R1632 B.n644 B.n439 256.663
R1633 B.n646 B.n439 256.663
R1634 B.n652 B.n439 256.663
R1635 B.n654 B.n439 256.663
R1636 B.n660 B.n439 256.663
R1637 B.n662 B.n439 256.663
R1638 B.n1027 B.n1026 256.663
R1639 B.n157 B.n156 163.367
R1640 B.n161 B.n160 163.367
R1641 B.n165 B.n164 163.367
R1642 B.n169 B.n168 163.367
R1643 B.n173 B.n172 163.367
R1644 B.n177 B.n176 163.367
R1645 B.n181 B.n180 163.367
R1646 B.n185 B.n184 163.367
R1647 B.n189 B.n188 163.367
R1648 B.n193 B.n192 163.367
R1649 B.n197 B.n196 163.367
R1650 B.n201 B.n200 163.367
R1651 B.n205 B.n204 163.367
R1652 B.n209 B.n208 163.367
R1653 B.n213 B.n212 163.367
R1654 B.n217 B.n216 163.367
R1655 B.n221 B.n220 163.367
R1656 B.n225 B.n224 163.367
R1657 B.n229 B.n228 163.367
R1658 B.n233 B.n232 163.367
R1659 B.n237 B.n236 163.367
R1660 B.n241 B.n240 163.367
R1661 B.n245 B.n244 163.367
R1662 B.n249 B.n248 163.367
R1663 B.n254 B.n253 163.367
R1664 B.n258 B.n257 163.367
R1665 B.n262 B.n261 163.367
R1666 B.n266 B.n265 163.367
R1667 B.n270 B.n269 163.367
R1668 B.n274 B.n273 163.367
R1669 B.n278 B.n277 163.367
R1670 B.n282 B.n281 163.367
R1671 B.n286 B.n285 163.367
R1672 B.n290 B.n289 163.367
R1673 B.n294 B.n293 163.367
R1674 B.n298 B.n297 163.367
R1675 B.n302 B.n301 163.367
R1676 B.n306 B.n305 163.367
R1677 B.n310 B.n309 163.367
R1678 B.n314 B.n313 163.367
R1679 B.n318 B.n317 163.367
R1680 B.n322 B.n321 163.367
R1681 B.n326 B.n325 163.367
R1682 B.n909 B.n149 163.367
R1683 B.n667 B.n434 163.367
R1684 B.n675 B.n434 163.367
R1685 B.n675 B.n432 163.367
R1686 B.n679 B.n432 163.367
R1687 B.n679 B.n425 163.367
R1688 B.n687 B.n425 163.367
R1689 B.n687 B.n423 163.367
R1690 B.n691 B.n423 163.367
R1691 B.n691 B.n418 163.367
R1692 B.n699 B.n418 163.367
R1693 B.n699 B.n416 163.367
R1694 B.n703 B.n416 163.367
R1695 B.n703 B.n410 163.367
R1696 B.n711 B.n410 163.367
R1697 B.n711 B.n408 163.367
R1698 B.n715 B.n408 163.367
R1699 B.n715 B.n402 163.367
R1700 B.n723 B.n402 163.367
R1701 B.n723 B.n400 163.367
R1702 B.n727 B.n400 163.367
R1703 B.n727 B.n394 163.367
R1704 B.n735 B.n394 163.367
R1705 B.n735 B.n392 163.367
R1706 B.n739 B.n392 163.367
R1707 B.n739 B.n386 163.367
R1708 B.n747 B.n386 163.367
R1709 B.n747 B.n384 163.367
R1710 B.n751 B.n384 163.367
R1711 B.n751 B.n378 163.367
R1712 B.n759 B.n378 163.367
R1713 B.n759 B.n376 163.367
R1714 B.n763 B.n376 163.367
R1715 B.n763 B.n370 163.367
R1716 B.n771 B.n370 163.367
R1717 B.n771 B.n368 163.367
R1718 B.n775 B.n368 163.367
R1719 B.n775 B.n362 163.367
R1720 B.n783 B.n362 163.367
R1721 B.n783 B.n360 163.367
R1722 B.n787 B.n360 163.367
R1723 B.n787 B.n354 163.367
R1724 B.n795 B.n354 163.367
R1725 B.n795 B.n352 163.367
R1726 B.n799 B.n352 163.367
R1727 B.n799 B.n346 163.367
R1728 B.n807 B.n346 163.367
R1729 B.n807 B.n344 163.367
R1730 B.n811 B.n344 163.367
R1731 B.n811 B.n338 163.367
R1732 B.n819 B.n338 163.367
R1733 B.n819 B.n336 163.367
R1734 B.n824 B.n336 163.367
R1735 B.n824 B.n330 163.367
R1736 B.n832 B.n330 163.367
R1737 B.n833 B.n832 163.367
R1738 B.n833 B.n5 163.367
R1739 B.n6 B.n5 163.367
R1740 B.n7 B.n6 163.367
R1741 B.n839 B.n7 163.367
R1742 B.n840 B.n839 163.367
R1743 B.n840 B.n13 163.367
R1744 B.n14 B.n13 163.367
R1745 B.n15 B.n14 163.367
R1746 B.n845 B.n15 163.367
R1747 B.n845 B.n20 163.367
R1748 B.n21 B.n20 163.367
R1749 B.n22 B.n21 163.367
R1750 B.n850 B.n22 163.367
R1751 B.n850 B.n27 163.367
R1752 B.n28 B.n27 163.367
R1753 B.n29 B.n28 163.367
R1754 B.n855 B.n29 163.367
R1755 B.n855 B.n34 163.367
R1756 B.n35 B.n34 163.367
R1757 B.n36 B.n35 163.367
R1758 B.n860 B.n36 163.367
R1759 B.n860 B.n41 163.367
R1760 B.n42 B.n41 163.367
R1761 B.n43 B.n42 163.367
R1762 B.n865 B.n43 163.367
R1763 B.n865 B.n48 163.367
R1764 B.n49 B.n48 163.367
R1765 B.n50 B.n49 163.367
R1766 B.n870 B.n50 163.367
R1767 B.n870 B.n55 163.367
R1768 B.n56 B.n55 163.367
R1769 B.n57 B.n56 163.367
R1770 B.n875 B.n57 163.367
R1771 B.n875 B.n62 163.367
R1772 B.n63 B.n62 163.367
R1773 B.n64 B.n63 163.367
R1774 B.n880 B.n64 163.367
R1775 B.n880 B.n69 163.367
R1776 B.n70 B.n69 163.367
R1777 B.n71 B.n70 163.367
R1778 B.n885 B.n71 163.367
R1779 B.n885 B.n76 163.367
R1780 B.n77 B.n76 163.367
R1781 B.n78 B.n77 163.367
R1782 B.n890 B.n78 163.367
R1783 B.n890 B.n83 163.367
R1784 B.n84 B.n83 163.367
R1785 B.n85 B.n84 163.367
R1786 B.n895 B.n85 163.367
R1787 B.n895 B.n90 163.367
R1788 B.n91 B.n90 163.367
R1789 B.n92 B.n91 163.367
R1790 B.n900 B.n92 163.367
R1791 B.n900 B.n97 163.367
R1792 B.n98 B.n97 163.367
R1793 B.n99 B.n98 163.367
R1794 B.n905 B.n99 163.367
R1795 B.n905 B.n104 163.367
R1796 B.n491 B.n490 163.367
R1797 B.n493 B.n491 163.367
R1798 B.n497 B.n486 163.367
R1799 B.n501 B.n499 163.367
R1800 B.n505 B.n484 163.367
R1801 B.n509 B.n507 163.367
R1802 B.n513 B.n482 163.367
R1803 B.n517 B.n515 163.367
R1804 B.n521 B.n480 163.367
R1805 B.n525 B.n523 163.367
R1806 B.n529 B.n478 163.367
R1807 B.n533 B.n531 163.367
R1808 B.n537 B.n476 163.367
R1809 B.n541 B.n539 163.367
R1810 B.n545 B.n474 163.367
R1811 B.n549 B.n547 163.367
R1812 B.n553 B.n472 163.367
R1813 B.n557 B.n555 163.367
R1814 B.n561 B.n470 163.367
R1815 B.n565 B.n563 163.367
R1816 B.n570 B.n466 163.367
R1817 B.n574 B.n572 163.367
R1818 B.n578 B.n464 163.367
R1819 B.n582 B.n580 163.367
R1820 B.n587 B.n460 163.367
R1821 B.n591 B.n589 163.367
R1822 B.n595 B.n458 163.367
R1823 B.n599 B.n597 163.367
R1824 B.n603 B.n456 163.367
R1825 B.n607 B.n605 163.367
R1826 B.n611 B.n454 163.367
R1827 B.n615 B.n613 163.367
R1828 B.n619 B.n452 163.367
R1829 B.n623 B.n621 163.367
R1830 B.n627 B.n450 163.367
R1831 B.n631 B.n629 163.367
R1832 B.n635 B.n448 163.367
R1833 B.n639 B.n637 163.367
R1834 B.n643 B.n446 163.367
R1835 B.n647 B.n645 163.367
R1836 B.n651 B.n444 163.367
R1837 B.n655 B.n653 163.367
R1838 B.n659 B.n442 163.367
R1839 B.n663 B.n661 163.367
R1840 B.n669 B.n436 163.367
R1841 B.n673 B.n436 163.367
R1842 B.n673 B.n430 163.367
R1843 B.n681 B.n430 163.367
R1844 B.n681 B.n428 163.367
R1845 B.n685 B.n428 163.367
R1846 B.n685 B.n422 163.367
R1847 B.n693 B.n422 163.367
R1848 B.n693 B.n420 163.367
R1849 B.n697 B.n420 163.367
R1850 B.n697 B.n414 163.367
R1851 B.n705 B.n414 163.367
R1852 B.n705 B.n412 163.367
R1853 B.n709 B.n412 163.367
R1854 B.n709 B.n406 163.367
R1855 B.n717 B.n406 163.367
R1856 B.n717 B.n404 163.367
R1857 B.n721 B.n404 163.367
R1858 B.n721 B.n398 163.367
R1859 B.n729 B.n398 163.367
R1860 B.n729 B.n396 163.367
R1861 B.n733 B.n396 163.367
R1862 B.n733 B.n390 163.367
R1863 B.n741 B.n390 163.367
R1864 B.n741 B.n388 163.367
R1865 B.n745 B.n388 163.367
R1866 B.n745 B.n382 163.367
R1867 B.n753 B.n382 163.367
R1868 B.n753 B.n380 163.367
R1869 B.n757 B.n380 163.367
R1870 B.n757 B.n374 163.367
R1871 B.n765 B.n374 163.367
R1872 B.n765 B.n372 163.367
R1873 B.n769 B.n372 163.367
R1874 B.n769 B.n366 163.367
R1875 B.n777 B.n366 163.367
R1876 B.n777 B.n364 163.367
R1877 B.n781 B.n364 163.367
R1878 B.n781 B.n358 163.367
R1879 B.n789 B.n358 163.367
R1880 B.n789 B.n356 163.367
R1881 B.n793 B.n356 163.367
R1882 B.n793 B.n350 163.367
R1883 B.n801 B.n350 163.367
R1884 B.n801 B.n348 163.367
R1885 B.n805 B.n348 163.367
R1886 B.n805 B.n342 163.367
R1887 B.n813 B.n342 163.367
R1888 B.n813 B.n340 163.367
R1889 B.n817 B.n340 163.367
R1890 B.n817 B.n334 163.367
R1891 B.n826 B.n334 163.367
R1892 B.n826 B.n332 163.367
R1893 B.n830 B.n332 163.367
R1894 B.n830 B.n3 163.367
R1895 B.n1025 B.n3 163.367
R1896 B.n1021 B.n2 163.367
R1897 B.n1021 B.n1020 163.367
R1898 B.n1020 B.n9 163.367
R1899 B.n1016 B.n9 163.367
R1900 B.n1016 B.n11 163.367
R1901 B.n1012 B.n11 163.367
R1902 B.n1012 B.n17 163.367
R1903 B.n1008 B.n17 163.367
R1904 B.n1008 B.n19 163.367
R1905 B.n1004 B.n19 163.367
R1906 B.n1004 B.n24 163.367
R1907 B.n1000 B.n24 163.367
R1908 B.n1000 B.n26 163.367
R1909 B.n996 B.n26 163.367
R1910 B.n996 B.n31 163.367
R1911 B.n992 B.n31 163.367
R1912 B.n992 B.n33 163.367
R1913 B.n988 B.n33 163.367
R1914 B.n988 B.n38 163.367
R1915 B.n984 B.n38 163.367
R1916 B.n984 B.n40 163.367
R1917 B.n980 B.n40 163.367
R1918 B.n980 B.n45 163.367
R1919 B.n976 B.n45 163.367
R1920 B.n976 B.n47 163.367
R1921 B.n972 B.n47 163.367
R1922 B.n972 B.n52 163.367
R1923 B.n968 B.n52 163.367
R1924 B.n968 B.n54 163.367
R1925 B.n964 B.n54 163.367
R1926 B.n964 B.n59 163.367
R1927 B.n960 B.n59 163.367
R1928 B.n960 B.n61 163.367
R1929 B.n956 B.n61 163.367
R1930 B.n956 B.n66 163.367
R1931 B.n952 B.n66 163.367
R1932 B.n952 B.n68 163.367
R1933 B.n948 B.n68 163.367
R1934 B.n948 B.n73 163.367
R1935 B.n944 B.n73 163.367
R1936 B.n944 B.n75 163.367
R1937 B.n940 B.n75 163.367
R1938 B.n940 B.n80 163.367
R1939 B.n936 B.n80 163.367
R1940 B.n936 B.n82 163.367
R1941 B.n932 B.n82 163.367
R1942 B.n932 B.n87 163.367
R1943 B.n928 B.n87 163.367
R1944 B.n928 B.n89 163.367
R1945 B.n924 B.n89 163.367
R1946 B.n924 B.n94 163.367
R1947 B.n920 B.n94 163.367
R1948 B.n920 B.n96 163.367
R1949 B.n916 B.n96 163.367
R1950 B.n916 B.n101 163.367
R1951 B.n912 B.n101 163.367
R1952 B.n668 B.n439 94.7881
R1953 B.n911 B.n910 94.7881
R1954 B.n105 B.n103 71.676
R1955 B.n157 B.n106 71.676
R1956 B.n161 B.n107 71.676
R1957 B.n165 B.n108 71.676
R1958 B.n169 B.n109 71.676
R1959 B.n173 B.n110 71.676
R1960 B.n177 B.n111 71.676
R1961 B.n181 B.n112 71.676
R1962 B.n185 B.n113 71.676
R1963 B.n189 B.n114 71.676
R1964 B.n193 B.n115 71.676
R1965 B.n197 B.n116 71.676
R1966 B.n201 B.n117 71.676
R1967 B.n205 B.n118 71.676
R1968 B.n209 B.n119 71.676
R1969 B.n213 B.n120 71.676
R1970 B.n217 B.n121 71.676
R1971 B.n221 B.n122 71.676
R1972 B.n225 B.n123 71.676
R1973 B.n229 B.n124 71.676
R1974 B.n233 B.n125 71.676
R1975 B.n237 B.n126 71.676
R1976 B.n241 B.n127 71.676
R1977 B.n245 B.n128 71.676
R1978 B.n249 B.n129 71.676
R1979 B.n254 B.n130 71.676
R1980 B.n258 B.n131 71.676
R1981 B.n262 B.n132 71.676
R1982 B.n266 B.n133 71.676
R1983 B.n270 B.n134 71.676
R1984 B.n274 B.n135 71.676
R1985 B.n278 B.n136 71.676
R1986 B.n282 B.n137 71.676
R1987 B.n286 B.n138 71.676
R1988 B.n290 B.n139 71.676
R1989 B.n294 B.n140 71.676
R1990 B.n298 B.n141 71.676
R1991 B.n302 B.n142 71.676
R1992 B.n306 B.n143 71.676
R1993 B.n310 B.n144 71.676
R1994 B.n314 B.n145 71.676
R1995 B.n318 B.n146 71.676
R1996 B.n322 B.n147 71.676
R1997 B.n326 B.n148 71.676
R1998 B.n149 B.n148 71.676
R1999 B.n325 B.n147 71.676
R2000 B.n321 B.n146 71.676
R2001 B.n317 B.n145 71.676
R2002 B.n313 B.n144 71.676
R2003 B.n309 B.n143 71.676
R2004 B.n305 B.n142 71.676
R2005 B.n301 B.n141 71.676
R2006 B.n297 B.n140 71.676
R2007 B.n293 B.n139 71.676
R2008 B.n289 B.n138 71.676
R2009 B.n285 B.n137 71.676
R2010 B.n281 B.n136 71.676
R2011 B.n277 B.n135 71.676
R2012 B.n273 B.n134 71.676
R2013 B.n269 B.n133 71.676
R2014 B.n265 B.n132 71.676
R2015 B.n261 B.n131 71.676
R2016 B.n257 B.n130 71.676
R2017 B.n253 B.n129 71.676
R2018 B.n248 B.n128 71.676
R2019 B.n244 B.n127 71.676
R2020 B.n240 B.n126 71.676
R2021 B.n236 B.n125 71.676
R2022 B.n232 B.n124 71.676
R2023 B.n228 B.n123 71.676
R2024 B.n224 B.n122 71.676
R2025 B.n220 B.n121 71.676
R2026 B.n216 B.n120 71.676
R2027 B.n212 B.n119 71.676
R2028 B.n208 B.n118 71.676
R2029 B.n204 B.n117 71.676
R2030 B.n200 B.n116 71.676
R2031 B.n196 B.n115 71.676
R2032 B.n192 B.n114 71.676
R2033 B.n188 B.n113 71.676
R2034 B.n184 B.n112 71.676
R2035 B.n180 B.n111 71.676
R2036 B.n176 B.n110 71.676
R2037 B.n172 B.n109 71.676
R2038 B.n168 B.n108 71.676
R2039 B.n164 B.n107 71.676
R2040 B.n160 B.n106 71.676
R2041 B.n156 B.n105 71.676
R2042 B.n489 B.n438 71.676
R2043 B.n493 B.n492 71.676
R2044 B.n498 B.n497 71.676
R2045 B.n501 B.n500 71.676
R2046 B.n506 B.n505 71.676
R2047 B.n509 B.n508 71.676
R2048 B.n514 B.n513 71.676
R2049 B.n517 B.n516 71.676
R2050 B.n522 B.n521 71.676
R2051 B.n525 B.n524 71.676
R2052 B.n530 B.n529 71.676
R2053 B.n533 B.n532 71.676
R2054 B.n538 B.n537 71.676
R2055 B.n541 B.n540 71.676
R2056 B.n546 B.n545 71.676
R2057 B.n549 B.n548 71.676
R2058 B.n554 B.n553 71.676
R2059 B.n557 B.n556 71.676
R2060 B.n562 B.n561 71.676
R2061 B.n565 B.n564 71.676
R2062 B.n571 B.n570 71.676
R2063 B.n574 B.n573 71.676
R2064 B.n579 B.n578 71.676
R2065 B.n582 B.n581 71.676
R2066 B.n588 B.n587 71.676
R2067 B.n591 B.n590 71.676
R2068 B.n596 B.n595 71.676
R2069 B.n599 B.n598 71.676
R2070 B.n604 B.n603 71.676
R2071 B.n607 B.n606 71.676
R2072 B.n612 B.n611 71.676
R2073 B.n615 B.n614 71.676
R2074 B.n620 B.n619 71.676
R2075 B.n623 B.n622 71.676
R2076 B.n628 B.n627 71.676
R2077 B.n631 B.n630 71.676
R2078 B.n636 B.n635 71.676
R2079 B.n639 B.n638 71.676
R2080 B.n644 B.n643 71.676
R2081 B.n647 B.n646 71.676
R2082 B.n652 B.n651 71.676
R2083 B.n655 B.n654 71.676
R2084 B.n660 B.n659 71.676
R2085 B.n663 B.n662 71.676
R2086 B.n490 B.n489 71.676
R2087 B.n492 B.n486 71.676
R2088 B.n499 B.n498 71.676
R2089 B.n500 B.n484 71.676
R2090 B.n507 B.n506 71.676
R2091 B.n508 B.n482 71.676
R2092 B.n515 B.n514 71.676
R2093 B.n516 B.n480 71.676
R2094 B.n523 B.n522 71.676
R2095 B.n524 B.n478 71.676
R2096 B.n531 B.n530 71.676
R2097 B.n532 B.n476 71.676
R2098 B.n539 B.n538 71.676
R2099 B.n540 B.n474 71.676
R2100 B.n547 B.n546 71.676
R2101 B.n548 B.n472 71.676
R2102 B.n555 B.n554 71.676
R2103 B.n556 B.n470 71.676
R2104 B.n563 B.n562 71.676
R2105 B.n564 B.n466 71.676
R2106 B.n572 B.n571 71.676
R2107 B.n573 B.n464 71.676
R2108 B.n580 B.n579 71.676
R2109 B.n581 B.n460 71.676
R2110 B.n589 B.n588 71.676
R2111 B.n590 B.n458 71.676
R2112 B.n597 B.n596 71.676
R2113 B.n598 B.n456 71.676
R2114 B.n605 B.n604 71.676
R2115 B.n606 B.n454 71.676
R2116 B.n613 B.n612 71.676
R2117 B.n614 B.n452 71.676
R2118 B.n621 B.n620 71.676
R2119 B.n622 B.n450 71.676
R2120 B.n629 B.n628 71.676
R2121 B.n630 B.n448 71.676
R2122 B.n637 B.n636 71.676
R2123 B.n638 B.n446 71.676
R2124 B.n645 B.n644 71.676
R2125 B.n646 B.n444 71.676
R2126 B.n653 B.n652 71.676
R2127 B.n654 B.n442 71.676
R2128 B.n661 B.n660 71.676
R2129 B.n662 B.n440 71.676
R2130 B.n1026 B.n1025 71.676
R2131 B.n1026 B.n2 71.676
R2132 B.n153 B.n152 64.1944
R2133 B.n151 B.n150 64.1944
R2134 B.n462 B.n461 64.1944
R2135 B.n468 B.n467 64.1944
R2136 B.n154 B.n153 59.5399
R2137 B.n251 B.n151 59.5399
R2138 B.n585 B.n462 59.5399
R2139 B.n567 B.n468 59.5399
R2140 B.n668 B.n435 45.0743
R2141 B.n674 B.n435 45.0743
R2142 B.n674 B.n431 45.0743
R2143 B.n680 B.n431 45.0743
R2144 B.n680 B.n426 45.0743
R2145 B.n686 B.n426 45.0743
R2146 B.n686 B.n427 45.0743
R2147 B.n692 B.n419 45.0743
R2148 B.n698 B.n419 45.0743
R2149 B.n698 B.n415 45.0743
R2150 B.n704 B.n415 45.0743
R2151 B.n704 B.n411 45.0743
R2152 B.n710 B.n411 45.0743
R2153 B.n710 B.n407 45.0743
R2154 B.n716 B.n407 45.0743
R2155 B.n716 B.n403 45.0743
R2156 B.n722 B.n403 45.0743
R2157 B.n722 B.n399 45.0743
R2158 B.n728 B.n399 45.0743
R2159 B.n734 B.n395 45.0743
R2160 B.n734 B.n391 45.0743
R2161 B.n740 B.n391 45.0743
R2162 B.n740 B.n387 45.0743
R2163 B.n746 B.n387 45.0743
R2164 B.n746 B.n383 45.0743
R2165 B.n752 B.n383 45.0743
R2166 B.n752 B.n379 45.0743
R2167 B.n758 B.n379 45.0743
R2168 B.n764 B.n375 45.0743
R2169 B.n764 B.n371 45.0743
R2170 B.n770 B.n371 45.0743
R2171 B.n770 B.n367 45.0743
R2172 B.n776 B.n367 45.0743
R2173 B.n776 B.n363 45.0743
R2174 B.n782 B.n363 45.0743
R2175 B.n782 B.n359 45.0743
R2176 B.n788 B.n359 45.0743
R2177 B.n794 B.n355 45.0743
R2178 B.n794 B.n351 45.0743
R2179 B.n800 B.n351 45.0743
R2180 B.n800 B.n347 45.0743
R2181 B.n806 B.n347 45.0743
R2182 B.n806 B.n343 45.0743
R2183 B.n812 B.n343 45.0743
R2184 B.n812 B.n339 45.0743
R2185 B.n818 B.n339 45.0743
R2186 B.n825 B.n335 45.0743
R2187 B.n825 B.n331 45.0743
R2188 B.n831 B.n331 45.0743
R2189 B.n831 B.n4 45.0743
R2190 B.n1024 B.n4 45.0743
R2191 B.n1024 B.n1023 45.0743
R2192 B.n1023 B.n1022 45.0743
R2193 B.n1022 B.n8 45.0743
R2194 B.n12 B.n8 45.0743
R2195 B.n1015 B.n12 45.0743
R2196 B.n1015 B.n1014 45.0743
R2197 B.n1013 B.n16 45.0743
R2198 B.n1007 B.n16 45.0743
R2199 B.n1007 B.n1006 45.0743
R2200 B.n1006 B.n1005 45.0743
R2201 B.n1005 B.n23 45.0743
R2202 B.n999 B.n23 45.0743
R2203 B.n999 B.n998 45.0743
R2204 B.n998 B.n997 45.0743
R2205 B.n997 B.n30 45.0743
R2206 B.n991 B.n990 45.0743
R2207 B.n990 B.n989 45.0743
R2208 B.n989 B.n37 45.0743
R2209 B.n983 B.n37 45.0743
R2210 B.n983 B.n982 45.0743
R2211 B.n982 B.n981 45.0743
R2212 B.n981 B.n44 45.0743
R2213 B.n975 B.n44 45.0743
R2214 B.n975 B.n974 45.0743
R2215 B.n973 B.n51 45.0743
R2216 B.n967 B.n51 45.0743
R2217 B.n967 B.n966 45.0743
R2218 B.n966 B.n965 45.0743
R2219 B.n965 B.n58 45.0743
R2220 B.n959 B.n58 45.0743
R2221 B.n959 B.n958 45.0743
R2222 B.n958 B.n957 45.0743
R2223 B.n957 B.n65 45.0743
R2224 B.n951 B.n950 45.0743
R2225 B.n950 B.n949 45.0743
R2226 B.n949 B.n72 45.0743
R2227 B.n943 B.n72 45.0743
R2228 B.n943 B.n942 45.0743
R2229 B.n942 B.n941 45.0743
R2230 B.n941 B.n79 45.0743
R2231 B.n935 B.n79 45.0743
R2232 B.n935 B.n934 45.0743
R2233 B.n934 B.n933 45.0743
R2234 B.n933 B.n86 45.0743
R2235 B.n927 B.n86 45.0743
R2236 B.n926 B.n925 45.0743
R2237 B.n925 B.n93 45.0743
R2238 B.n919 B.n93 45.0743
R2239 B.n919 B.n918 45.0743
R2240 B.n918 B.n917 45.0743
R2241 B.n917 B.n100 45.0743
R2242 B.n911 B.n100 45.0743
R2243 B.t1 B.n335 43.7486
R2244 B.n1014 B.t0 43.7486
R2245 B.n427 B.t13 39.7715
R2246 B.t9 B.n926 39.7715
R2247 B.n728 B.t2 37.1201
R2248 B.n951 B.t6 37.1201
R2249 B.n670 B.n437 34.4981
R2250 B.n666 B.n665 34.4981
R2251 B.n908 B.n907 34.4981
R2252 B.n913 B.n102 34.4981
R2253 B.t5 B.n355 31.8173
R2254 B.t4 B.n30 31.8173
R2255 B.n758 B.t3 25.1888
R2256 B.t7 B.n973 25.1888
R2257 B.t3 B.n375 19.886
R2258 B.n974 B.t7 19.886
R2259 B B.n1027 18.0485
R2260 B.n788 B.t5 13.2575
R2261 B.n991 B.t4 13.2575
R2262 B.n671 B.n670 10.6151
R2263 B.n672 B.n671 10.6151
R2264 B.n672 B.n429 10.6151
R2265 B.n682 B.n429 10.6151
R2266 B.n683 B.n682 10.6151
R2267 B.n684 B.n683 10.6151
R2268 B.n684 B.n421 10.6151
R2269 B.n694 B.n421 10.6151
R2270 B.n695 B.n694 10.6151
R2271 B.n696 B.n695 10.6151
R2272 B.n696 B.n413 10.6151
R2273 B.n706 B.n413 10.6151
R2274 B.n707 B.n706 10.6151
R2275 B.n708 B.n707 10.6151
R2276 B.n708 B.n405 10.6151
R2277 B.n718 B.n405 10.6151
R2278 B.n719 B.n718 10.6151
R2279 B.n720 B.n719 10.6151
R2280 B.n720 B.n397 10.6151
R2281 B.n730 B.n397 10.6151
R2282 B.n731 B.n730 10.6151
R2283 B.n732 B.n731 10.6151
R2284 B.n732 B.n389 10.6151
R2285 B.n742 B.n389 10.6151
R2286 B.n743 B.n742 10.6151
R2287 B.n744 B.n743 10.6151
R2288 B.n744 B.n381 10.6151
R2289 B.n754 B.n381 10.6151
R2290 B.n755 B.n754 10.6151
R2291 B.n756 B.n755 10.6151
R2292 B.n756 B.n373 10.6151
R2293 B.n766 B.n373 10.6151
R2294 B.n767 B.n766 10.6151
R2295 B.n768 B.n767 10.6151
R2296 B.n768 B.n365 10.6151
R2297 B.n778 B.n365 10.6151
R2298 B.n779 B.n778 10.6151
R2299 B.n780 B.n779 10.6151
R2300 B.n780 B.n357 10.6151
R2301 B.n790 B.n357 10.6151
R2302 B.n791 B.n790 10.6151
R2303 B.n792 B.n791 10.6151
R2304 B.n792 B.n349 10.6151
R2305 B.n802 B.n349 10.6151
R2306 B.n803 B.n802 10.6151
R2307 B.n804 B.n803 10.6151
R2308 B.n804 B.n341 10.6151
R2309 B.n814 B.n341 10.6151
R2310 B.n815 B.n814 10.6151
R2311 B.n816 B.n815 10.6151
R2312 B.n816 B.n333 10.6151
R2313 B.n827 B.n333 10.6151
R2314 B.n828 B.n827 10.6151
R2315 B.n829 B.n828 10.6151
R2316 B.n829 B.n0 10.6151
R2317 B.n488 B.n437 10.6151
R2318 B.n488 B.n487 10.6151
R2319 B.n494 B.n487 10.6151
R2320 B.n495 B.n494 10.6151
R2321 B.n496 B.n495 10.6151
R2322 B.n496 B.n485 10.6151
R2323 B.n502 B.n485 10.6151
R2324 B.n503 B.n502 10.6151
R2325 B.n504 B.n503 10.6151
R2326 B.n504 B.n483 10.6151
R2327 B.n510 B.n483 10.6151
R2328 B.n511 B.n510 10.6151
R2329 B.n512 B.n511 10.6151
R2330 B.n512 B.n481 10.6151
R2331 B.n518 B.n481 10.6151
R2332 B.n519 B.n518 10.6151
R2333 B.n520 B.n519 10.6151
R2334 B.n520 B.n479 10.6151
R2335 B.n526 B.n479 10.6151
R2336 B.n527 B.n526 10.6151
R2337 B.n528 B.n527 10.6151
R2338 B.n528 B.n477 10.6151
R2339 B.n534 B.n477 10.6151
R2340 B.n535 B.n534 10.6151
R2341 B.n536 B.n535 10.6151
R2342 B.n536 B.n475 10.6151
R2343 B.n542 B.n475 10.6151
R2344 B.n543 B.n542 10.6151
R2345 B.n544 B.n543 10.6151
R2346 B.n544 B.n473 10.6151
R2347 B.n550 B.n473 10.6151
R2348 B.n551 B.n550 10.6151
R2349 B.n552 B.n551 10.6151
R2350 B.n552 B.n471 10.6151
R2351 B.n558 B.n471 10.6151
R2352 B.n559 B.n558 10.6151
R2353 B.n560 B.n559 10.6151
R2354 B.n560 B.n469 10.6151
R2355 B.n566 B.n469 10.6151
R2356 B.n569 B.n568 10.6151
R2357 B.n569 B.n465 10.6151
R2358 B.n575 B.n465 10.6151
R2359 B.n576 B.n575 10.6151
R2360 B.n577 B.n576 10.6151
R2361 B.n577 B.n463 10.6151
R2362 B.n583 B.n463 10.6151
R2363 B.n584 B.n583 10.6151
R2364 B.n586 B.n459 10.6151
R2365 B.n592 B.n459 10.6151
R2366 B.n593 B.n592 10.6151
R2367 B.n594 B.n593 10.6151
R2368 B.n594 B.n457 10.6151
R2369 B.n600 B.n457 10.6151
R2370 B.n601 B.n600 10.6151
R2371 B.n602 B.n601 10.6151
R2372 B.n602 B.n455 10.6151
R2373 B.n608 B.n455 10.6151
R2374 B.n609 B.n608 10.6151
R2375 B.n610 B.n609 10.6151
R2376 B.n610 B.n453 10.6151
R2377 B.n616 B.n453 10.6151
R2378 B.n617 B.n616 10.6151
R2379 B.n618 B.n617 10.6151
R2380 B.n618 B.n451 10.6151
R2381 B.n624 B.n451 10.6151
R2382 B.n625 B.n624 10.6151
R2383 B.n626 B.n625 10.6151
R2384 B.n626 B.n449 10.6151
R2385 B.n632 B.n449 10.6151
R2386 B.n633 B.n632 10.6151
R2387 B.n634 B.n633 10.6151
R2388 B.n634 B.n447 10.6151
R2389 B.n640 B.n447 10.6151
R2390 B.n641 B.n640 10.6151
R2391 B.n642 B.n641 10.6151
R2392 B.n642 B.n445 10.6151
R2393 B.n648 B.n445 10.6151
R2394 B.n649 B.n648 10.6151
R2395 B.n650 B.n649 10.6151
R2396 B.n650 B.n443 10.6151
R2397 B.n656 B.n443 10.6151
R2398 B.n657 B.n656 10.6151
R2399 B.n658 B.n657 10.6151
R2400 B.n658 B.n441 10.6151
R2401 B.n664 B.n441 10.6151
R2402 B.n665 B.n664 10.6151
R2403 B.n666 B.n433 10.6151
R2404 B.n676 B.n433 10.6151
R2405 B.n677 B.n676 10.6151
R2406 B.n678 B.n677 10.6151
R2407 B.n678 B.n424 10.6151
R2408 B.n688 B.n424 10.6151
R2409 B.n689 B.n688 10.6151
R2410 B.n690 B.n689 10.6151
R2411 B.n690 B.n417 10.6151
R2412 B.n700 B.n417 10.6151
R2413 B.n701 B.n700 10.6151
R2414 B.n702 B.n701 10.6151
R2415 B.n702 B.n409 10.6151
R2416 B.n712 B.n409 10.6151
R2417 B.n713 B.n712 10.6151
R2418 B.n714 B.n713 10.6151
R2419 B.n714 B.n401 10.6151
R2420 B.n724 B.n401 10.6151
R2421 B.n725 B.n724 10.6151
R2422 B.n726 B.n725 10.6151
R2423 B.n726 B.n393 10.6151
R2424 B.n736 B.n393 10.6151
R2425 B.n737 B.n736 10.6151
R2426 B.n738 B.n737 10.6151
R2427 B.n738 B.n385 10.6151
R2428 B.n748 B.n385 10.6151
R2429 B.n749 B.n748 10.6151
R2430 B.n750 B.n749 10.6151
R2431 B.n750 B.n377 10.6151
R2432 B.n760 B.n377 10.6151
R2433 B.n761 B.n760 10.6151
R2434 B.n762 B.n761 10.6151
R2435 B.n762 B.n369 10.6151
R2436 B.n772 B.n369 10.6151
R2437 B.n773 B.n772 10.6151
R2438 B.n774 B.n773 10.6151
R2439 B.n774 B.n361 10.6151
R2440 B.n784 B.n361 10.6151
R2441 B.n785 B.n784 10.6151
R2442 B.n786 B.n785 10.6151
R2443 B.n786 B.n353 10.6151
R2444 B.n796 B.n353 10.6151
R2445 B.n797 B.n796 10.6151
R2446 B.n798 B.n797 10.6151
R2447 B.n798 B.n345 10.6151
R2448 B.n808 B.n345 10.6151
R2449 B.n809 B.n808 10.6151
R2450 B.n810 B.n809 10.6151
R2451 B.n810 B.n337 10.6151
R2452 B.n820 B.n337 10.6151
R2453 B.n821 B.n820 10.6151
R2454 B.n823 B.n821 10.6151
R2455 B.n823 B.n822 10.6151
R2456 B.n822 B.n329 10.6151
R2457 B.n834 B.n329 10.6151
R2458 B.n835 B.n834 10.6151
R2459 B.n836 B.n835 10.6151
R2460 B.n837 B.n836 10.6151
R2461 B.n838 B.n837 10.6151
R2462 B.n841 B.n838 10.6151
R2463 B.n842 B.n841 10.6151
R2464 B.n843 B.n842 10.6151
R2465 B.n844 B.n843 10.6151
R2466 B.n846 B.n844 10.6151
R2467 B.n847 B.n846 10.6151
R2468 B.n848 B.n847 10.6151
R2469 B.n849 B.n848 10.6151
R2470 B.n851 B.n849 10.6151
R2471 B.n852 B.n851 10.6151
R2472 B.n853 B.n852 10.6151
R2473 B.n854 B.n853 10.6151
R2474 B.n856 B.n854 10.6151
R2475 B.n857 B.n856 10.6151
R2476 B.n858 B.n857 10.6151
R2477 B.n859 B.n858 10.6151
R2478 B.n861 B.n859 10.6151
R2479 B.n862 B.n861 10.6151
R2480 B.n863 B.n862 10.6151
R2481 B.n864 B.n863 10.6151
R2482 B.n866 B.n864 10.6151
R2483 B.n867 B.n866 10.6151
R2484 B.n868 B.n867 10.6151
R2485 B.n869 B.n868 10.6151
R2486 B.n871 B.n869 10.6151
R2487 B.n872 B.n871 10.6151
R2488 B.n873 B.n872 10.6151
R2489 B.n874 B.n873 10.6151
R2490 B.n876 B.n874 10.6151
R2491 B.n877 B.n876 10.6151
R2492 B.n878 B.n877 10.6151
R2493 B.n879 B.n878 10.6151
R2494 B.n881 B.n879 10.6151
R2495 B.n882 B.n881 10.6151
R2496 B.n883 B.n882 10.6151
R2497 B.n884 B.n883 10.6151
R2498 B.n886 B.n884 10.6151
R2499 B.n887 B.n886 10.6151
R2500 B.n888 B.n887 10.6151
R2501 B.n889 B.n888 10.6151
R2502 B.n891 B.n889 10.6151
R2503 B.n892 B.n891 10.6151
R2504 B.n893 B.n892 10.6151
R2505 B.n894 B.n893 10.6151
R2506 B.n896 B.n894 10.6151
R2507 B.n897 B.n896 10.6151
R2508 B.n898 B.n897 10.6151
R2509 B.n899 B.n898 10.6151
R2510 B.n901 B.n899 10.6151
R2511 B.n902 B.n901 10.6151
R2512 B.n903 B.n902 10.6151
R2513 B.n904 B.n903 10.6151
R2514 B.n906 B.n904 10.6151
R2515 B.n907 B.n906 10.6151
R2516 B.n1019 B.n1 10.6151
R2517 B.n1019 B.n1018 10.6151
R2518 B.n1018 B.n1017 10.6151
R2519 B.n1017 B.n10 10.6151
R2520 B.n1011 B.n10 10.6151
R2521 B.n1011 B.n1010 10.6151
R2522 B.n1010 B.n1009 10.6151
R2523 B.n1009 B.n18 10.6151
R2524 B.n1003 B.n18 10.6151
R2525 B.n1003 B.n1002 10.6151
R2526 B.n1002 B.n1001 10.6151
R2527 B.n1001 B.n25 10.6151
R2528 B.n995 B.n25 10.6151
R2529 B.n995 B.n994 10.6151
R2530 B.n994 B.n993 10.6151
R2531 B.n993 B.n32 10.6151
R2532 B.n987 B.n32 10.6151
R2533 B.n987 B.n986 10.6151
R2534 B.n986 B.n985 10.6151
R2535 B.n985 B.n39 10.6151
R2536 B.n979 B.n39 10.6151
R2537 B.n979 B.n978 10.6151
R2538 B.n978 B.n977 10.6151
R2539 B.n977 B.n46 10.6151
R2540 B.n971 B.n46 10.6151
R2541 B.n971 B.n970 10.6151
R2542 B.n970 B.n969 10.6151
R2543 B.n969 B.n53 10.6151
R2544 B.n963 B.n53 10.6151
R2545 B.n963 B.n962 10.6151
R2546 B.n962 B.n961 10.6151
R2547 B.n961 B.n60 10.6151
R2548 B.n955 B.n60 10.6151
R2549 B.n955 B.n954 10.6151
R2550 B.n954 B.n953 10.6151
R2551 B.n953 B.n67 10.6151
R2552 B.n947 B.n67 10.6151
R2553 B.n947 B.n946 10.6151
R2554 B.n946 B.n945 10.6151
R2555 B.n945 B.n74 10.6151
R2556 B.n939 B.n74 10.6151
R2557 B.n939 B.n938 10.6151
R2558 B.n938 B.n937 10.6151
R2559 B.n937 B.n81 10.6151
R2560 B.n931 B.n81 10.6151
R2561 B.n931 B.n930 10.6151
R2562 B.n930 B.n929 10.6151
R2563 B.n929 B.n88 10.6151
R2564 B.n923 B.n88 10.6151
R2565 B.n923 B.n922 10.6151
R2566 B.n922 B.n921 10.6151
R2567 B.n921 B.n95 10.6151
R2568 B.n915 B.n95 10.6151
R2569 B.n915 B.n914 10.6151
R2570 B.n914 B.n913 10.6151
R2571 B.n155 B.n102 10.6151
R2572 B.n158 B.n155 10.6151
R2573 B.n159 B.n158 10.6151
R2574 B.n162 B.n159 10.6151
R2575 B.n163 B.n162 10.6151
R2576 B.n166 B.n163 10.6151
R2577 B.n167 B.n166 10.6151
R2578 B.n170 B.n167 10.6151
R2579 B.n171 B.n170 10.6151
R2580 B.n174 B.n171 10.6151
R2581 B.n175 B.n174 10.6151
R2582 B.n178 B.n175 10.6151
R2583 B.n179 B.n178 10.6151
R2584 B.n182 B.n179 10.6151
R2585 B.n183 B.n182 10.6151
R2586 B.n186 B.n183 10.6151
R2587 B.n187 B.n186 10.6151
R2588 B.n190 B.n187 10.6151
R2589 B.n191 B.n190 10.6151
R2590 B.n194 B.n191 10.6151
R2591 B.n195 B.n194 10.6151
R2592 B.n198 B.n195 10.6151
R2593 B.n199 B.n198 10.6151
R2594 B.n202 B.n199 10.6151
R2595 B.n203 B.n202 10.6151
R2596 B.n206 B.n203 10.6151
R2597 B.n207 B.n206 10.6151
R2598 B.n210 B.n207 10.6151
R2599 B.n211 B.n210 10.6151
R2600 B.n214 B.n211 10.6151
R2601 B.n215 B.n214 10.6151
R2602 B.n218 B.n215 10.6151
R2603 B.n219 B.n218 10.6151
R2604 B.n222 B.n219 10.6151
R2605 B.n223 B.n222 10.6151
R2606 B.n226 B.n223 10.6151
R2607 B.n227 B.n226 10.6151
R2608 B.n230 B.n227 10.6151
R2609 B.n231 B.n230 10.6151
R2610 B.n235 B.n234 10.6151
R2611 B.n238 B.n235 10.6151
R2612 B.n239 B.n238 10.6151
R2613 B.n242 B.n239 10.6151
R2614 B.n243 B.n242 10.6151
R2615 B.n246 B.n243 10.6151
R2616 B.n247 B.n246 10.6151
R2617 B.n250 B.n247 10.6151
R2618 B.n255 B.n252 10.6151
R2619 B.n256 B.n255 10.6151
R2620 B.n259 B.n256 10.6151
R2621 B.n260 B.n259 10.6151
R2622 B.n263 B.n260 10.6151
R2623 B.n264 B.n263 10.6151
R2624 B.n267 B.n264 10.6151
R2625 B.n268 B.n267 10.6151
R2626 B.n271 B.n268 10.6151
R2627 B.n272 B.n271 10.6151
R2628 B.n275 B.n272 10.6151
R2629 B.n276 B.n275 10.6151
R2630 B.n279 B.n276 10.6151
R2631 B.n280 B.n279 10.6151
R2632 B.n283 B.n280 10.6151
R2633 B.n284 B.n283 10.6151
R2634 B.n287 B.n284 10.6151
R2635 B.n288 B.n287 10.6151
R2636 B.n291 B.n288 10.6151
R2637 B.n292 B.n291 10.6151
R2638 B.n295 B.n292 10.6151
R2639 B.n296 B.n295 10.6151
R2640 B.n299 B.n296 10.6151
R2641 B.n300 B.n299 10.6151
R2642 B.n303 B.n300 10.6151
R2643 B.n304 B.n303 10.6151
R2644 B.n307 B.n304 10.6151
R2645 B.n308 B.n307 10.6151
R2646 B.n311 B.n308 10.6151
R2647 B.n312 B.n311 10.6151
R2648 B.n315 B.n312 10.6151
R2649 B.n316 B.n315 10.6151
R2650 B.n319 B.n316 10.6151
R2651 B.n320 B.n319 10.6151
R2652 B.n323 B.n320 10.6151
R2653 B.n324 B.n323 10.6151
R2654 B.n327 B.n324 10.6151
R2655 B.n328 B.n327 10.6151
R2656 B.n908 B.n328 10.6151
R2657 B.n1027 B.n0 8.11757
R2658 B.n1027 B.n1 8.11757
R2659 B.t2 B.n395 7.9547
R2660 B.t6 B.n65 7.9547
R2661 B.n568 B.n567 6.5566
R2662 B.n585 B.n584 6.5566
R2663 B.n234 B.n154 6.5566
R2664 B.n251 B.n250 6.5566
R2665 B.n692 B.t13 5.3033
R2666 B.n927 B.t9 5.3033
R2667 B.n567 B.n566 4.05904
R2668 B.n586 B.n585 4.05904
R2669 B.n231 B.n154 4.05904
R2670 B.n252 B.n251 4.05904
R2671 B.n818 B.t1 1.3262
R2672 B.t0 B.n1013 1.3262
R2673 VN.n60 VN.n59 161.3
R2674 VN.n58 VN.n32 161.3
R2675 VN.n57 VN.n56 161.3
R2676 VN.n55 VN.n33 161.3
R2677 VN.n54 VN.n53 161.3
R2678 VN.n52 VN.n34 161.3
R2679 VN.n50 VN.n49 161.3
R2680 VN.n48 VN.n35 161.3
R2681 VN.n47 VN.n46 161.3
R2682 VN.n45 VN.n36 161.3
R2683 VN.n44 VN.n43 161.3
R2684 VN.n42 VN.n37 161.3
R2685 VN.n41 VN.n40 161.3
R2686 VN.n29 VN.n28 161.3
R2687 VN.n27 VN.n1 161.3
R2688 VN.n26 VN.n25 161.3
R2689 VN.n24 VN.n2 161.3
R2690 VN.n23 VN.n22 161.3
R2691 VN.n21 VN.n3 161.3
R2692 VN.n19 VN.n18 161.3
R2693 VN.n17 VN.n4 161.3
R2694 VN.n16 VN.n15 161.3
R2695 VN.n14 VN.n5 161.3
R2696 VN.n13 VN.n12 161.3
R2697 VN.n11 VN.n6 161.3
R2698 VN.n10 VN.n9 161.3
R2699 VN.n38 VN.t3 123.234
R2700 VN.n7 VN.t2 123.234
R2701 VN.n8 VN.t4 91.5481
R2702 VN.n20 VN.t7 91.5481
R2703 VN.n0 VN.t5 91.5481
R2704 VN.n39 VN.t6 91.5481
R2705 VN.n51 VN.t0 91.5481
R2706 VN.n31 VN.t1 91.5481
R2707 VN.n30 VN.n0 67.2516
R2708 VN.n61 VN.n31 67.2516
R2709 VN.n8 VN.n7 66.0815
R2710 VN.n39 VN.n38 66.0814
R2711 VN.n26 VN.n2 56.4773
R2712 VN.n57 VN.n33 56.4773
R2713 VN VN.n61 52.4828
R2714 VN.n14 VN.n13 40.4106
R2715 VN.n15 VN.n14 40.4106
R2716 VN.n45 VN.n44 40.4106
R2717 VN.n46 VN.n45 40.4106
R2718 VN.n9 VN.n6 24.3439
R2719 VN.n13 VN.n6 24.3439
R2720 VN.n15 VN.n4 24.3439
R2721 VN.n19 VN.n4 24.3439
R2722 VN.n22 VN.n21 24.3439
R2723 VN.n22 VN.n2 24.3439
R2724 VN.n27 VN.n26 24.3439
R2725 VN.n28 VN.n27 24.3439
R2726 VN.n44 VN.n37 24.3439
R2727 VN.n40 VN.n37 24.3439
R2728 VN.n53 VN.n33 24.3439
R2729 VN.n53 VN.n52 24.3439
R2730 VN.n50 VN.n35 24.3439
R2731 VN.n46 VN.n35 24.3439
R2732 VN.n59 VN.n58 24.3439
R2733 VN.n58 VN.n57 24.3439
R2734 VN.n28 VN.n0 22.6399
R2735 VN.n59 VN.n31 22.6399
R2736 VN.n21 VN.n20 16.7975
R2737 VN.n52 VN.n51 16.7975
R2738 VN.n9 VN.n8 7.54696
R2739 VN.n20 VN.n19 7.54696
R2740 VN.n40 VN.n39 7.54696
R2741 VN.n51 VN.n50 7.54696
R2742 VN.n10 VN.n7 5.37324
R2743 VN.n41 VN.n38 5.37324
R2744 VN.n61 VN.n60 0.355081
R2745 VN.n30 VN.n29 0.355081
R2746 VN VN.n30 0.26685
R2747 VN.n60 VN.n32 0.189894
R2748 VN.n56 VN.n32 0.189894
R2749 VN.n56 VN.n55 0.189894
R2750 VN.n55 VN.n54 0.189894
R2751 VN.n54 VN.n34 0.189894
R2752 VN.n49 VN.n34 0.189894
R2753 VN.n49 VN.n48 0.189894
R2754 VN.n48 VN.n47 0.189894
R2755 VN.n47 VN.n36 0.189894
R2756 VN.n43 VN.n36 0.189894
R2757 VN.n43 VN.n42 0.189894
R2758 VN.n42 VN.n41 0.189894
R2759 VN.n11 VN.n10 0.189894
R2760 VN.n12 VN.n11 0.189894
R2761 VN.n12 VN.n5 0.189894
R2762 VN.n16 VN.n5 0.189894
R2763 VN.n17 VN.n16 0.189894
R2764 VN.n18 VN.n17 0.189894
R2765 VN.n18 VN.n3 0.189894
R2766 VN.n23 VN.n3 0.189894
R2767 VN.n24 VN.n23 0.189894
R2768 VN.n25 VN.n24 0.189894
R2769 VN.n25 VN.n1 0.189894
R2770 VN.n29 VN.n1 0.189894
R2771 VDD2.n2 VDD2.n1 61.9096
R2772 VDD2.n2 VDD2.n0 61.9096
R2773 VDD2 VDD2.n5 61.9067
R2774 VDD2.n4 VDD2.n3 60.5384
R2775 VDD2.n4 VDD2.n2 46.3144
R2776 VDD2.n5 VDD2.t1 1.74962
R2777 VDD2.n5 VDD2.t4 1.74962
R2778 VDD2.n3 VDD2.t6 1.74962
R2779 VDD2.n3 VDD2.t7 1.74962
R2780 VDD2.n1 VDD2.t0 1.74962
R2781 VDD2.n1 VDD2.t2 1.74962
R2782 VDD2.n0 VDD2.t5 1.74962
R2783 VDD2.n0 VDD2.t3 1.74962
R2784 VDD2 VDD2.n4 1.48541
C0 VN VDD1 0.152201f
C1 VN VTAIL 8.995461f
C2 VTAIL VDD1 7.97259f
C3 VP VDD2 0.559893f
C4 VN VP 8.008639f
C5 VP VDD1 8.836329f
C6 VTAIL VP 9.00957f
C7 VN VDD2 8.43023f
C8 VDD1 VDD2 1.97617f
C9 VTAIL VDD2 8.02955f
C10 VDD2 B 5.655513f
C11 VDD1 B 6.136851f
C12 VTAIL B 10.33222f
C13 VN B 16.92587f
C14 VP B 15.555052f
C15 VDD2.t5 B 0.215397f
C16 VDD2.t3 B 0.215397f
C17 VDD2.n0 B 1.92259f
C18 VDD2.t0 B 0.215397f
C19 VDD2.t2 B 0.215397f
C20 VDD2.n1 B 1.92259f
C21 VDD2.n2 B 3.33103f
C22 VDD2.t6 B 0.215397f
C23 VDD2.t7 B 0.215397f
C24 VDD2.n3 B 1.91068f
C25 VDD2.n4 B 2.92045f
C26 VDD2.t1 B 0.215397f
C27 VDD2.t4 B 0.215397f
C28 VDD2.n5 B 1.92255f
C29 VN.t5 B 1.87427f
C30 VN.n0 B 0.747359f
C31 VN.n1 B 0.020427f
C32 VN.n2 B 0.033389f
C33 VN.n3 B 0.020427f
C34 VN.t7 B 1.87427f
C35 VN.n4 B 0.038262f
C36 VN.n5 B 0.020427f
C37 VN.n6 B 0.038262f
C38 VN.t2 B 2.08051f
C39 VN.n7 B 0.703065f
C40 VN.t4 B 1.87427f
C41 VN.n8 B 0.72435f
C42 VN.n9 B 0.025227f
C43 VN.n10 B 0.219465f
C44 VN.n11 B 0.020427f
C45 VN.n12 B 0.020427f
C46 VN.n13 B 0.040816f
C47 VN.n14 B 0.01653f
C48 VN.n15 B 0.040816f
C49 VN.n16 B 0.020427f
C50 VN.n17 B 0.020427f
C51 VN.n18 B 0.020427f
C52 VN.n19 B 0.025227f
C53 VN.n20 B 0.662603f
C54 VN.n21 B 0.032406f
C55 VN.n22 B 0.038262f
C56 VN.n23 B 0.020427f
C57 VN.n24 B 0.020427f
C58 VN.n25 B 0.020427f
C59 VN.n26 B 0.02651f
C60 VN.n27 B 0.038262f
C61 VN.n28 B 0.03694f
C62 VN.n29 B 0.032974f
C63 VN.n30 B 0.039711f
C64 VN.t1 B 1.87427f
C65 VN.n31 B 0.747359f
C66 VN.n32 B 0.020427f
C67 VN.n33 B 0.033389f
C68 VN.n34 B 0.020427f
C69 VN.t0 B 1.87427f
C70 VN.n35 B 0.038262f
C71 VN.n36 B 0.020427f
C72 VN.n37 B 0.038262f
C73 VN.t3 B 2.08051f
C74 VN.n38 B 0.703065f
C75 VN.t6 B 1.87427f
C76 VN.n39 B 0.72435f
C77 VN.n40 B 0.025227f
C78 VN.n41 B 0.219465f
C79 VN.n42 B 0.020427f
C80 VN.n43 B 0.020427f
C81 VN.n44 B 0.040816f
C82 VN.n45 B 0.01653f
C83 VN.n46 B 0.040816f
C84 VN.n47 B 0.020427f
C85 VN.n48 B 0.020427f
C86 VN.n49 B 0.020427f
C87 VN.n50 B 0.025227f
C88 VN.n51 B 0.662603f
C89 VN.n52 B 0.032406f
C90 VN.n53 B 0.038262f
C91 VN.n54 B 0.020427f
C92 VN.n55 B 0.020427f
C93 VN.n56 B 0.020427f
C94 VN.n57 B 0.02651f
C95 VN.n58 B 0.038262f
C96 VN.n59 B 0.03694f
C97 VN.n60 B 0.032974f
C98 VN.n61 B 1.23813f
C99 VDD1.t5 B 0.219461f
C100 VDD1.t7 B 0.219461f
C101 VDD1.n0 B 1.96006f
C102 VDD1.t2 B 0.219461f
C103 VDD1.t6 B 0.219461f
C104 VDD1.n1 B 1.95886f
C105 VDD1.t1 B 0.219461f
C106 VDD1.t4 B 0.219461f
C107 VDD1.n2 B 1.95886f
C108 VDD1.n3 B 3.44479f
C109 VDD1.t0 B 0.219461f
C110 VDD1.t3 B 0.219461f
C111 VDD1.n4 B 1.94672f
C112 VDD1.n5 B 3.00604f
C113 VTAIL.t4 B 0.181858f
C114 VTAIL.t7 B 0.181858f
C115 VTAIL.n0 B 1.55038f
C116 VTAIL.n1 B 0.394859f
C117 VTAIL.n2 B 0.026929f
C118 VTAIL.n3 B 0.02033f
C119 VTAIL.n4 B 0.010924f
C120 VTAIL.n5 B 0.025821f
C121 VTAIL.n6 B 0.011567f
C122 VTAIL.n7 B 0.02033f
C123 VTAIL.n8 B 0.010924f
C124 VTAIL.n9 B 0.025821f
C125 VTAIL.n10 B 0.011246f
C126 VTAIL.n11 B 0.02033f
C127 VTAIL.n12 B 0.011567f
C128 VTAIL.n13 B 0.025821f
C129 VTAIL.n14 B 0.011567f
C130 VTAIL.n15 B 0.02033f
C131 VTAIL.n16 B 0.010924f
C132 VTAIL.n17 B 0.025821f
C133 VTAIL.n18 B 0.011567f
C134 VTAIL.n19 B 0.964115f
C135 VTAIL.n20 B 0.010924f
C136 VTAIL.t0 B 0.043536f
C137 VTAIL.n21 B 0.141269f
C138 VTAIL.n22 B 0.018254f
C139 VTAIL.n23 B 0.019366f
C140 VTAIL.n24 B 0.025821f
C141 VTAIL.n25 B 0.011567f
C142 VTAIL.n26 B 0.010924f
C143 VTAIL.n27 B 0.02033f
C144 VTAIL.n28 B 0.02033f
C145 VTAIL.n29 B 0.010924f
C146 VTAIL.n30 B 0.011567f
C147 VTAIL.n31 B 0.025821f
C148 VTAIL.n32 B 0.025821f
C149 VTAIL.n33 B 0.011567f
C150 VTAIL.n34 B 0.010924f
C151 VTAIL.n35 B 0.02033f
C152 VTAIL.n36 B 0.02033f
C153 VTAIL.n37 B 0.010924f
C154 VTAIL.n38 B 0.010924f
C155 VTAIL.n39 B 0.011567f
C156 VTAIL.n40 B 0.025821f
C157 VTAIL.n41 B 0.025821f
C158 VTAIL.n42 B 0.025821f
C159 VTAIL.n43 B 0.011246f
C160 VTAIL.n44 B 0.010924f
C161 VTAIL.n45 B 0.02033f
C162 VTAIL.n46 B 0.02033f
C163 VTAIL.n47 B 0.010924f
C164 VTAIL.n48 B 0.011567f
C165 VTAIL.n49 B 0.025821f
C166 VTAIL.n50 B 0.025821f
C167 VTAIL.n51 B 0.011567f
C168 VTAIL.n52 B 0.010924f
C169 VTAIL.n53 B 0.02033f
C170 VTAIL.n54 B 0.02033f
C171 VTAIL.n55 B 0.010924f
C172 VTAIL.n56 B 0.011567f
C173 VTAIL.n57 B 0.025821f
C174 VTAIL.n58 B 0.052988f
C175 VTAIL.n59 B 0.011567f
C176 VTAIL.n60 B 0.010924f
C177 VTAIL.n61 B 0.04477f
C178 VTAIL.n62 B 0.02928f
C179 VTAIL.n63 B 0.233809f
C180 VTAIL.n64 B 0.026929f
C181 VTAIL.n65 B 0.02033f
C182 VTAIL.n66 B 0.010924f
C183 VTAIL.n67 B 0.025821f
C184 VTAIL.n68 B 0.011567f
C185 VTAIL.n69 B 0.02033f
C186 VTAIL.n70 B 0.010924f
C187 VTAIL.n71 B 0.025821f
C188 VTAIL.n72 B 0.011246f
C189 VTAIL.n73 B 0.02033f
C190 VTAIL.n74 B 0.011567f
C191 VTAIL.n75 B 0.025821f
C192 VTAIL.n76 B 0.011567f
C193 VTAIL.n77 B 0.02033f
C194 VTAIL.n78 B 0.010924f
C195 VTAIL.n79 B 0.025821f
C196 VTAIL.n80 B 0.011567f
C197 VTAIL.n81 B 0.964115f
C198 VTAIL.n82 B 0.010924f
C199 VTAIL.t10 B 0.043536f
C200 VTAIL.n83 B 0.141269f
C201 VTAIL.n84 B 0.018254f
C202 VTAIL.n85 B 0.019366f
C203 VTAIL.n86 B 0.025821f
C204 VTAIL.n87 B 0.011567f
C205 VTAIL.n88 B 0.010924f
C206 VTAIL.n89 B 0.02033f
C207 VTAIL.n90 B 0.02033f
C208 VTAIL.n91 B 0.010924f
C209 VTAIL.n92 B 0.011567f
C210 VTAIL.n93 B 0.025821f
C211 VTAIL.n94 B 0.025821f
C212 VTAIL.n95 B 0.011567f
C213 VTAIL.n96 B 0.010924f
C214 VTAIL.n97 B 0.02033f
C215 VTAIL.n98 B 0.02033f
C216 VTAIL.n99 B 0.010924f
C217 VTAIL.n100 B 0.010924f
C218 VTAIL.n101 B 0.011567f
C219 VTAIL.n102 B 0.025821f
C220 VTAIL.n103 B 0.025821f
C221 VTAIL.n104 B 0.025821f
C222 VTAIL.n105 B 0.011246f
C223 VTAIL.n106 B 0.010924f
C224 VTAIL.n107 B 0.02033f
C225 VTAIL.n108 B 0.02033f
C226 VTAIL.n109 B 0.010924f
C227 VTAIL.n110 B 0.011567f
C228 VTAIL.n111 B 0.025821f
C229 VTAIL.n112 B 0.025821f
C230 VTAIL.n113 B 0.011567f
C231 VTAIL.n114 B 0.010924f
C232 VTAIL.n115 B 0.02033f
C233 VTAIL.n116 B 0.02033f
C234 VTAIL.n117 B 0.010924f
C235 VTAIL.n118 B 0.011567f
C236 VTAIL.n119 B 0.025821f
C237 VTAIL.n120 B 0.052988f
C238 VTAIL.n121 B 0.011567f
C239 VTAIL.n122 B 0.010924f
C240 VTAIL.n123 B 0.04477f
C241 VTAIL.n124 B 0.02928f
C242 VTAIL.n125 B 0.233809f
C243 VTAIL.t12 B 0.181858f
C244 VTAIL.t9 B 0.181858f
C245 VTAIL.n126 B 1.55038f
C246 VTAIL.n127 B 0.577968f
C247 VTAIL.n128 B 0.026929f
C248 VTAIL.n129 B 0.02033f
C249 VTAIL.n130 B 0.010924f
C250 VTAIL.n131 B 0.025821f
C251 VTAIL.n132 B 0.011567f
C252 VTAIL.n133 B 0.02033f
C253 VTAIL.n134 B 0.010924f
C254 VTAIL.n135 B 0.025821f
C255 VTAIL.n136 B 0.011246f
C256 VTAIL.n137 B 0.02033f
C257 VTAIL.n138 B 0.011567f
C258 VTAIL.n139 B 0.025821f
C259 VTAIL.n140 B 0.011567f
C260 VTAIL.n141 B 0.02033f
C261 VTAIL.n142 B 0.010924f
C262 VTAIL.n143 B 0.025821f
C263 VTAIL.n144 B 0.011567f
C264 VTAIL.n145 B 0.964115f
C265 VTAIL.n146 B 0.010924f
C266 VTAIL.t11 B 0.043536f
C267 VTAIL.n147 B 0.141269f
C268 VTAIL.n148 B 0.018254f
C269 VTAIL.n149 B 0.019366f
C270 VTAIL.n150 B 0.025821f
C271 VTAIL.n151 B 0.011567f
C272 VTAIL.n152 B 0.010924f
C273 VTAIL.n153 B 0.02033f
C274 VTAIL.n154 B 0.02033f
C275 VTAIL.n155 B 0.010924f
C276 VTAIL.n156 B 0.011567f
C277 VTAIL.n157 B 0.025821f
C278 VTAIL.n158 B 0.025821f
C279 VTAIL.n159 B 0.011567f
C280 VTAIL.n160 B 0.010924f
C281 VTAIL.n161 B 0.02033f
C282 VTAIL.n162 B 0.02033f
C283 VTAIL.n163 B 0.010924f
C284 VTAIL.n164 B 0.010924f
C285 VTAIL.n165 B 0.011567f
C286 VTAIL.n166 B 0.025821f
C287 VTAIL.n167 B 0.025821f
C288 VTAIL.n168 B 0.025821f
C289 VTAIL.n169 B 0.011246f
C290 VTAIL.n170 B 0.010924f
C291 VTAIL.n171 B 0.02033f
C292 VTAIL.n172 B 0.02033f
C293 VTAIL.n173 B 0.010924f
C294 VTAIL.n174 B 0.011567f
C295 VTAIL.n175 B 0.025821f
C296 VTAIL.n176 B 0.025821f
C297 VTAIL.n177 B 0.011567f
C298 VTAIL.n178 B 0.010924f
C299 VTAIL.n179 B 0.02033f
C300 VTAIL.n180 B 0.02033f
C301 VTAIL.n181 B 0.010924f
C302 VTAIL.n182 B 0.011567f
C303 VTAIL.n183 B 0.025821f
C304 VTAIL.n184 B 0.052988f
C305 VTAIL.n185 B 0.011567f
C306 VTAIL.n186 B 0.010924f
C307 VTAIL.n187 B 0.04477f
C308 VTAIL.n188 B 0.02928f
C309 VTAIL.n189 B 1.30537f
C310 VTAIL.n190 B 0.026929f
C311 VTAIL.n191 B 0.02033f
C312 VTAIL.n192 B 0.010924f
C313 VTAIL.n193 B 0.025821f
C314 VTAIL.n194 B 0.011567f
C315 VTAIL.n195 B 0.02033f
C316 VTAIL.n196 B 0.010924f
C317 VTAIL.n197 B 0.025821f
C318 VTAIL.n198 B 0.011246f
C319 VTAIL.n199 B 0.02033f
C320 VTAIL.n200 B 0.011246f
C321 VTAIL.n201 B 0.010924f
C322 VTAIL.n202 B 0.025821f
C323 VTAIL.n203 B 0.025821f
C324 VTAIL.n204 B 0.011567f
C325 VTAIL.n205 B 0.02033f
C326 VTAIL.n206 B 0.010924f
C327 VTAIL.n207 B 0.025821f
C328 VTAIL.n208 B 0.011567f
C329 VTAIL.n209 B 0.964115f
C330 VTAIL.n210 B 0.010924f
C331 VTAIL.t2 B 0.043536f
C332 VTAIL.n211 B 0.141269f
C333 VTAIL.n212 B 0.018254f
C334 VTAIL.n213 B 0.019366f
C335 VTAIL.n214 B 0.025821f
C336 VTAIL.n215 B 0.011567f
C337 VTAIL.n216 B 0.010924f
C338 VTAIL.n217 B 0.02033f
C339 VTAIL.n218 B 0.02033f
C340 VTAIL.n219 B 0.010924f
C341 VTAIL.n220 B 0.011567f
C342 VTAIL.n221 B 0.025821f
C343 VTAIL.n222 B 0.025821f
C344 VTAIL.n223 B 0.011567f
C345 VTAIL.n224 B 0.010924f
C346 VTAIL.n225 B 0.02033f
C347 VTAIL.n226 B 0.02033f
C348 VTAIL.n227 B 0.010924f
C349 VTAIL.n228 B 0.011567f
C350 VTAIL.n229 B 0.025821f
C351 VTAIL.n230 B 0.025821f
C352 VTAIL.n231 B 0.011567f
C353 VTAIL.n232 B 0.010924f
C354 VTAIL.n233 B 0.02033f
C355 VTAIL.n234 B 0.02033f
C356 VTAIL.n235 B 0.010924f
C357 VTAIL.n236 B 0.011567f
C358 VTAIL.n237 B 0.025821f
C359 VTAIL.n238 B 0.025821f
C360 VTAIL.n239 B 0.011567f
C361 VTAIL.n240 B 0.010924f
C362 VTAIL.n241 B 0.02033f
C363 VTAIL.n242 B 0.02033f
C364 VTAIL.n243 B 0.010924f
C365 VTAIL.n244 B 0.011567f
C366 VTAIL.n245 B 0.025821f
C367 VTAIL.n246 B 0.052988f
C368 VTAIL.n247 B 0.011567f
C369 VTAIL.n248 B 0.010924f
C370 VTAIL.n249 B 0.04477f
C371 VTAIL.n250 B 0.02928f
C372 VTAIL.n251 B 1.30537f
C373 VTAIL.t3 B 0.181858f
C374 VTAIL.t5 B 0.181858f
C375 VTAIL.n252 B 1.55039f
C376 VTAIL.n253 B 0.577959f
C377 VTAIL.n254 B 0.026929f
C378 VTAIL.n255 B 0.02033f
C379 VTAIL.n256 B 0.010924f
C380 VTAIL.n257 B 0.025821f
C381 VTAIL.n258 B 0.011567f
C382 VTAIL.n259 B 0.02033f
C383 VTAIL.n260 B 0.010924f
C384 VTAIL.n261 B 0.025821f
C385 VTAIL.n262 B 0.011246f
C386 VTAIL.n263 B 0.02033f
C387 VTAIL.n264 B 0.011246f
C388 VTAIL.n265 B 0.010924f
C389 VTAIL.n266 B 0.025821f
C390 VTAIL.n267 B 0.025821f
C391 VTAIL.n268 B 0.011567f
C392 VTAIL.n269 B 0.02033f
C393 VTAIL.n270 B 0.010924f
C394 VTAIL.n271 B 0.025821f
C395 VTAIL.n272 B 0.011567f
C396 VTAIL.n273 B 0.964115f
C397 VTAIL.n274 B 0.010924f
C398 VTAIL.t1 B 0.043536f
C399 VTAIL.n275 B 0.141269f
C400 VTAIL.n276 B 0.018254f
C401 VTAIL.n277 B 0.019366f
C402 VTAIL.n278 B 0.025821f
C403 VTAIL.n279 B 0.011567f
C404 VTAIL.n280 B 0.010924f
C405 VTAIL.n281 B 0.02033f
C406 VTAIL.n282 B 0.02033f
C407 VTAIL.n283 B 0.010924f
C408 VTAIL.n284 B 0.011567f
C409 VTAIL.n285 B 0.025821f
C410 VTAIL.n286 B 0.025821f
C411 VTAIL.n287 B 0.011567f
C412 VTAIL.n288 B 0.010924f
C413 VTAIL.n289 B 0.02033f
C414 VTAIL.n290 B 0.02033f
C415 VTAIL.n291 B 0.010924f
C416 VTAIL.n292 B 0.011567f
C417 VTAIL.n293 B 0.025821f
C418 VTAIL.n294 B 0.025821f
C419 VTAIL.n295 B 0.011567f
C420 VTAIL.n296 B 0.010924f
C421 VTAIL.n297 B 0.02033f
C422 VTAIL.n298 B 0.02033f
C423 VTAIL.n299 B 0.010924f
C424 VTAIL.n300 B 0.011567f
C425 VTAIL.n301 B 0.025821f
C426 VTAIL.n302 B 0.025821f
C427 VTAIL.n303 B 0.011567f
C428 VTAIL.n304 B 0.010924f
C429 VTAIL.n305 B 0.02033f
C430 VTAIL.n306 B 0.02033f
C431 VTAIL.n307 B 0.010924f
C432 VTAIL.n308 B 0.011567f
C433 VTAIL.n309 B 0.025821f
C434 VTAIL.n310 B 0.052988f
C435 VTAIL.n311 B 0.011567f
C436 VTAIL.n312 B 0.010924f
C437 VTAIL.n313 B 0.04477f
C438 VTAIL.n314 B 0.02928f
C439 VTAIL.n315 B 0.233809f
C440 VTAIL.n316 B 0.026929f
C441 VTAIL.n317 B 0.02033f
C442 VTAIL.n318 B 0.010924f
C443 VTAIL.n319 B 0.025821f
C444 VTAIL.n320 B 0.011567f
C445 VTAIL.n321 B 0.02033f
C446 VTAIL.n322 B 0.010924f
C447 VTAIL.n323 B 0.025821f
C448 VTAIL.n324 B 0.011246f
C449 VTAIL.n325 B 0.02033f
C450 VTAIL.n326 B 0.011246f
C451 VTAIL.n327 B 0.010924f
C452 VTAIL.n328 B 0.025821f
C453 VTAIL.n329 B 0.025821f
C454 VTAIL.n330 B 0.011567f
C455 VTAIL.n331 B 0.02033f
C456 VTAIL.n332 B 0.010924f
C457 VTAIL.n333 B 0.025821f
C458 VTAIL.n334 B 0.011567f
C459 VTAIL.n335 B 0.964115f
C460 VTAIL.n336 B 0.010924f
C461 VTAIL.t13 B 0.043536f
C462 VTAIL.n337 B 0.141269f
C463 VTAIL.n338 B 0.018254f
C464 VTAIL.n339 B 0.019366f
C465 VTAIL.n340 B 0.025821f
C466 VTAIL.n341 B 0.011567f
C467 VTAIL.n342 B 0.010924f
C468 VTAIL.n343 B 0.02033f
C469 VTAIL.n344 B 0.02033f
C470 VTAIL.n345 B 0.010924f
C471 VTAIL.n346 B 0.011567f
C472 VTAIL.n347 B 0.025821f
C473 VTAIL.n348 B 0.025821f
C474 VTAIL.n349 B 0.011567f
C475 VTAIL.n350 B 0.010924f
C476 VTAIL.n351 B 0.02033f
C477 VTAIL.n352 B 0.02033f
C478 VTAIL.n353 B 0.010924f
C479 VTAIL.n354 B 0.011567f
C480 VTAIL.n355 B 0.025821f
C481 VTAIL.n356 B 0.025821f
C482 VTAIL.n357 B 0.011567f
C483 VTAIL.n358 B 0.010924f
C484 VTAIL.n359 B 0.02033f
C485 VTAIL.n360 B 0.02033f
C486 VTAIL.n361 B 0.010924f
C487 VTAIL.n362 B 0.011567f
C488 VTAIL.n363 B 0.025821f
C489 VTAIL.n364 B 0.025821f
C490 VTAIL.n365 B 0.011567f
C491 VTAIL.n366 B 0.010924f
C492 VTAIL.n367 B 0.02033f
C493 VTAIL.n368 B 0.02033f
C494 VTAIL.n369 B 0.010924f
C495 VTAIL.n370 B 0.011567f
C496 VTAIL.n371 B 0.025821f
C497 VTAIL.n372 B 0.052988f
C498 VTAIL.n373 B 0.011567f
C499 VTAIL.n374 B 0.010924f
C500 VTAIL.n375 B 0.04477f
C501 VTAIL.n376 B 0.02928f
C502 VTAIL.n377 B 0.233809f
C503 VTAIL.t8 B 0.181858f
C504 VTAIL.t15 B 0.181858f
C505 VTAIL.n378 B 1.55039f
C506 VTAIL.n379 B 0.577959f
C507 VTAIL.n380 B 0.026929f
C508 VTAIL.n381 B 0.02033f
C509 VTAIL.n382 B 0.010924f
C510 VTAIL.n383 B 0.025821f
C511 VTAIL.n384 B 0.011567f
C512 VTAIL.n385 B 0.02033f
C513 VTAIL.n386 B 0.010924f
C514 VTAIL.n387 B 0.025821f
C515 VTAIL.n388 B 0.011246f
C516 VTAIL.n389 B 0.02033f
C517 VTAIL.n390 B 0.011246f
C518 VTAIL.n391 B 0.010924f
C519 VTAIL.n392 B 0.025821f
C520 VTAIL.n393 B 0.025821f
C521 VTAIL.n394 B 0.011567f
C522 VTAIL.n395 B 0.02033f
C523 VTAIL.n396 B 0.010924f
C524 VTAIL.n397 B 0.025821f
C525 VTAIL.n398 B 0.011567f
C526 VTAIL.n399 B 0.964115f
C527 VTAIL.n400 B 0.010924f
C528 VTAIL.t14 B 0.043536f
C529 VTAIL.n401 B 0.141269f
C530 VTAIL.n402 B 0.018254f
C531 VTAIL.n403 B 0.019366f
C532 VTAIL.n404 B 0.025821f
C533 VTAIL.n405 B 0.011567f
C534 VTAIL.n406 B 0.010924f
C535 VTAIL.n407 B 0.02033f
C536 VTAIL.n408 B 0.02033f
C537 VTAIL.n409 B 0.010924f
C538 VTAIL.n410 B 0.011567f
C539 VTAIL.n411 B 0.025821f
C540 VTAIL.n412 B 0.025821f
C541 VTAIL.n413 B 0.011567f
C542 VTAIL.n414 B 0.010924f
C543 VTAIL.n415 B 0.02033f
C544 VTAIL.n416 B 0.02033f
C545 VTAIL.n417 B 0.010924f
C546 VTAIL.n418 B 0.011567f
C547 VTAIL.n419 B 0.025821f
C548 VTAIL.n420 B 0.025821f
C549 VTAIL.n421 B 0.011567f
C550 VTAIL.n422 B 0.010924f
C551 VTAIL.n423 B 0.02033f
C552 VTAIL.n424 B 0.02033f
C553 VTAIL.n425 B 0.010924f
C554 VTAIL.n426 B 0.011567f
C555 VTAIL.n427 B 0.025821f
C556 VTAIL.n428 B 0.025821f
C557 VTAIL.n429 B 0.011567f
C558 VTAIL.n430 B 0.010924f
C559 VTAIL.n431 B 0.02033f
C560 VTAIL.n432 B 0.02033f
C561 VTAIL.n433 B 0.010924f
C562 VTAIL.n434 B 0.011567f
C563 VTAIL.n435 B 0.025821f
C564 VTAIL.n436 B 0.052988f
C565 VTAIL.n437 B 0.011567f
C566 VTAIL.n438 B 0.010924f
C567 VTAIL.n439 B 0.04477f
C568 VTAIL.n440 B 0.02928f
C569 VTAIL.n441 B 1.30537f
C570 VTAIL.n442 B 0.026929f
C571 VTAIL.n443 B 0.02033f
C572 VTAIL.n444 B 0.010924f
C573 VTAIL.n445 B 0.025821f
C574 VTAIL.n446 B 0.011567f
C575 VTAIL.n447 B 0.02033f
C576 VTAIL.n448 B 0.010924f
C577 VTAIL.n449 B 0.025821f
C578 VTAIL.n450 B 0.011246f
C579 VTAIL.n451 B 0.02033f
C580 VTAIL.n452 B 0.011567f
C581 VTAIL.n453 B 0.025821f
C582 VTAIL.n454 B 0.011567f
C583 VTAIL.n455 B 0.02033f
C584 VTAIL.n456 B 0.010924f
C585 VTAIL.n457 B 0.025821f
C586 VTAIL.n458 B 0.011567f
C587 VTAIL.n459 B 0.964115f
C588 VTAIL.n460 B 0.010924f
C589 VTAIL.t6 B 0.043536f
C590 VTAIL.n461 B 0.141269f
C591 VTAIL.n462 B 0.018254f
C592 VTAIL.n463 B 0.019366f
C593 VTAIL.n464 B 0.025821f
C594 VTAIL.n465 B 0.011567f
C595 VTAIL.n466 B 0.010924f
C596 VTAIL.n467 B 0.02033f
C597 VTAIL.n468 B 0.02033f
C598 VTAIL.n469 B 0.010924f
C599 VTAIL.n470 B 0.011567f
C600 VTAIL.n471 B 0.025821f
C601 VTAIL.n472 B 0.025821f
C602 VTAIL.n473 B 0.011567f
C603 VTAIL.n474 B 0.010924f
C604 VTAIL.n475 B 0.02033f
C605 VTAIL.n476 B 0.02033f
C606 VTAIL.n477 B 0.010924f
C607 VTAIL.n478 B 0.010924f
C608 VTAIL.n479 B 0.011567f
C609 VTAIL.n480 B 0.025821f
C610 VTAIL.n481 B 0.025821f
C611 VTAIL.n482 B 0.025821f
C612 VTAIL.n483 B 0.011246f
C613 VTAIL.n484 B 0.010924f
C614 VTAIL.n485 B 0.02033f
C615 VTAIL.n486 B 0.02033f
C616 VTAIL.n487 B 0.010924f
C617 VTAIL.n488 B 0.011567f
C618 VTAIL.n489 B 0.025821f
C619 VTAIL.n490 B 0.025821f
C620 VTAIL.n491 B 0.011567f
C621 VTAIL.n492 B 0.010924f
C622 VTAIL.n493 B 0.02033f
C623 VTAIL.n494 B 0.02033f
C624 VTAIL.n495 B 0.010924f
C625 VTAIL.n496 B 0.011567f
C626 VTAIL.n497 B 0.025821f
C627 VTAIL.n498 B 0.052988f
C628 VTAIL.n499 B 0.011567f
C629 VTAIL.n500 B 0.010924f
C630 VTAIL.n501 B 0.04477f
C631 VTAIL.n502 B 0.02928f
C632 VTAIL.n503 B 1.30156f
C633 VP.t3 B 1.90594f
C634 VP.n0 B 0.759987f
C635 VP.n1 B 0.020772f
C636 VP.n2 B 0.033954f
C637 VP.n3 B 0.020772f
C638 VP.t6 B 1.90594f
C639 VP.n4 B 0.038909f
C640 VP.n5 B 0.020772f
C641 VP.n6 B 0.038909f
C642 VP.n7 B 0.020772f
C643 VP.t1 B 1.90594f
C644 VP.n8 B 0.033954f
C645 VP.n9 B 0.020772f
C646 VP.t5 B 1.90594f
C647 VP.n10 B 0.759987f
C648 VP.t4 B 1.90594f
C649 VP.n11 B 0.759987f
C650 VP.n12 B 0.020772f
C651 VP.n13 B 0.033954f
C652 VP.n14 B 0.020772f
C653 VP.t7 B 1.90594f
C654 VP.n15 B 0.038909f
C655 VP.n16 B 0.020772f
C656 VP.n17 B 0.038909f
C657 VP.t2 B 2.11566f
C658 VP.n18 B 0.714946f
C659 VP.t0 B 1.90594f
C660 VP.n19 B 0.73659f
C661 VP.n20 B 0.025653f
C662 VP.n21 B 0.223174f
C663 VP.n22 B 0.020772f
C664 VP.n23 B 0.020772f
C665 VP.n24 B 0.041506f
C666 VP.n25 B 0.016809f
C667 VP.n26 B 0.041506f
C668 VP.n27 B 0.020772f
C669 VP.n28 B 0.020772f
C670 VP.n29 B 0.020772f
C671 VP.n30 B 0.025653f
C672 VP.n31 B 0.673799f
C673 VP.n32 B 0.032953f
C674 VP.n33 B 0.038909f
C675 VP.n34 B 0.020772f
C676 VP.n35 B 0.020772f
C677 VP.n36 B 0.020772f
C678 VP.n37 B 0.026958f
C679 VP.n38 B 0.038909f
C680 VP.n39 B 0.037564f
C681 VP.n40 B 0.033532f
C682 VP.n41 B 1.25069f
C683 VP.n42 B 1.26492f
C684 VP.n43 B 0.033532f
C685 VP.n44 B 0.037564f
C686 VP.n45 B 0.038909f
C687 VP.n46 B 0.026958f
C688 VP.n47 B 0.020772f
C689 VP.n48 B 0.020772f
C690 VP.n49 B 0.020772f
C691 VP.n50 B 0.038909f
C692 VP.n51 B 0.032953f
C693 VP.n52 B 0.673799f
C694 VP.n53 B 0.025653f
C695 VP.n54 B 0.020772f
C696 VP.n55 B 0.020772f
C697 VP.n56 B 0.020772f
C698 VP.n57 B 0.041506f
C699 VP.n58 B 0.016809f
C700 VP.n59 B 0.041506f
C701 VP.n60 B 0.020772f
C702 VP.n61 B 0.020772f
C703 VP.n62 B 0.020772f
C704 VP.n63 B 0.025653f
C705 VP.n64 B 0.673799f
C706 VP.n65 B 0.032953f
C707 VP.n66 B 0.038909f
C708 VP.n67 B 0.020772f
C709 VP.n68 B 0.020772f
C710 VP.n69 B 0.020772f
C711 VP.n70 B 0.026958f
C712 VP.n71 B 0.038909f
C713 VP.n72 B 0.037564f
C714 VP.n73 B 0.033532f
C715 VP.n74 B 0.040382f
.ends

