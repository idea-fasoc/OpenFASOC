* NGSPICE file created from diff_pair_sample_1112.ext - technology: sky130A

.subckt diff_pair_sample_1112 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1730_n3240# sky130_fd_pr__pfet_01v8 ad=4.4304 pd=23.5 as=4.4304 ps=23.5 w=11.36 l=1.57
X1 B.t11 B.t9 B.t10 w_n1730_n3240# sky130_fd_pr__pfet_01v8 ad=4.4304 pd=23.5 as=0 ps=0 w=11.36 l=1.57
X2 B.t8 B.t6 B.t7 w_n1730_n3240# sky130_fd_pr__pfet_01v8 ad=4.4304 pd=23.5 as=0 ps=0 w=11.36 l=1.57
X3 VDD2.t0 VN.t1 VTAIL.t3 w_n1730_n3240# sky130_fd_pr__pfet_01v8 ad=4.4304 pd=23.5 as=4.4304 ps=23.5 w=11.36 l=1.57
X4 VDD1.t1 VP.t0 VTAIL.t0 w_n1730_n3240# sky130_fd_pr__pfet_01v8 ad=4.4304 pd=23.5 as=4.4304 ps=23.5 w=11.36 l=1.57
X5 B.t5 B.t3 B.t4 w_n1730_n3240# sky130_fd_pr__pfet_01v8 ad=4.4304 pd=23.5 as=0 ps=0 w=11.36 l=1.57
X6 B.t2 B.t0 B.t1 w_n1730_n3240# sky130_fd_pr__pfet_01v8 ad=4.4304 pd=23.5 as=0 ps=0 w=11.36 l=1.57
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n1730_n3240# sky130_fd_pr__pfet_01v8 ad=4.4304 pd=23.5 as=4.4304 ps=23.5 w=11.36 l=1.57
R0 VN VN.t1 321.731
R1 VN VN.t0 280.151
R2 VTAIL.n242 VTAIL.n186 756.745
R3 VTAIL.n56 VTAIL.n0 756.745
R4 VTAIL.n180 VTAIL.n124 756.745
R5 VTAIL.n118 VTAIL.n62 756.745
R6 VTAIL.n207 VTAIL.n206 585
R7 VTAIL.n209 VTAIL.n208 585
R8 VTAIL.n202 VTAIL.n201 585
R9 VTAIL.n215 VTAIL.n214 585
R10 VTAIL.n217 VTAIL.n216 585
R11 VTAIL.n198 VTAIL.n197 585
R12 VTAIL.n224 VTAIL.n223 585
R13 VTAIL.n225 VTAIL.n196 585
R14 VTAIL.n227 VTAIL.n226 585
R15 VTAIL.n194 VTAIL.n193 585
R16 VTAIL.n233 VTAIL.n232 585
R17 VTAIL.n235 VTAIL.n234 585
R18 VTAIL.n190 VTAIL.n189 585
R19 VTAIL.n241 VTAIL.n240 585
R20 VTAIL.n243 VTAIL.n242 585
R21 VTAIL.n21 VTAIL.n20 585
R22 VTAIL.n23 VTAIL.n22 585
R23 VTAIL.n16 VTAIL.n15 585
R24 VTAIL.n29 VTAIL.n28 585
R25 VTAIL.n31 VTAIL.n30 585
R26 VTAIL.n12 VTAIL.n11 585
R27 VTAIL.n38 VTAIL.n37 585
R28 VTAIL.n39 VTAIL.n10 585
R29 VTAIL.n41 VTAIL.n40 585
R30 VTAIL.n8 VTAIL.n7 585
R31 VTAIL.n47 VTAIL.n46 585
R32 VTAIL.n49 VTAIL.n48 585
R33 VTAIL.n4 VTAIL.n3 585
R34 VTAIL.n55 VTAIL.n54 585
R35 VTAIL.n57 VTAIL.n56 585
R36 VTAIL.n181 VTAIL.n180 585
R37 VTAIL.n179 VTAIL.n178 585
R38 VTAIL.n128 VTAIL.n127 585
R39 VTAIL.n173 VTAIL.n172 585
R40 VTAIL.n171 VTAIL.n170 585
R41 VTAIL.n132 VTAIL.n131 585
R42 VTAIL.n136 VTAIL.n134 585
R43 VTAIL.n165 VTAIL.n164 585
R44 VTAIL.n163 VTAIL.n162 585
R45 VTAIL.n138 VTAIL.n137 585
R46 VTAIL.n157 VTAIL.n156 585
R47 VTAIL.n155 VTAIL.n154 585
R48 VTAIL.n142 VTAIL.n141 585
R49 VTAIL.n149 VTAIL.n148 585
R50 VTAIL.n147 VTAIL.n146 585
R51 VTAIL.n119 VTAIL.n118 585
R52 VTAIL.n117 VTAIL.n116 585
R53 VTAIL.n66 VTAIL.n65 585
R54 VTAIL.n111 VTAIL.n110 585
R55 VTAIL.n109 VTAIL.n108 585
R56 VTAIL.n70 VTAIL.n69 585
R57 VTAIL.n74 VTAIL.n72 585
R58 VTAIL.n103 VTAIL.n102 585
R59 VTAIL.n101 VTAIL.n100 585
R60 VTAIL.n76 VTAIL.n75 585
R61 VTAIL.n95 VTAIL.n94 585
R62 VTAIL.n93 VTAIL.n92 585
R63 VTAIL.n80 VTAIL.n79 585
R64 VTAIL.n87 VTAIL.n86 585
R65 VTAIL.n85 VTAIL.n84 585
R66 VTAIL.n205 VTAIL.t2 329.036
R67 VTAIL.n19 VTAIL.t0 329.036
R68 VTAIL.n145 VTAIL.t1 329.036
R69 VTAIL.n83 VTAIL.t3 329.036
R70 VTAIL.n208 VTAIL.n207 171.744
R71 VTAIL.n208 VTAIL.n201 171.744
R72 VTAIL.n215 VTAIL.n201 171.744
R73 VTAIL.n216 VTAIL.n215 171.744
R74 VTAIL.n216 VTAIL.n197 171.744
R75 VTAIL.n224 VTAIL.n197 171.744
R76 VTAIL.n225 VTAIL.n224 171.744
R77 VTAIL.n226 VTAIL.n225 171.744
R78 VTAIL.n226 VTAIL.n193 171.744
R79 VTAIL.n233 VTAIL.n193 171.744
R80 VTAIL.n234 VTAIL.n233 171.744
R81 VTAIL.n234 VTAIL.n189 171.744
R82 VTAIL.n241 VTAIL.n189 171.744
R83 VTAIL.n242 VTAIL.n241 171.744
R84 VTAIL.n22 VTAIL.n21 171.744
R85 VTAIL.n22 VTAIL.n15 171.744
R86 VTAIL.n29 VTAIL.n15 171.744
R87 VTAIL.n30 VTAIL.n29 171.744
R88 VTAIL.n30 VTAIL.n11 171.744
R89 VTAIL.n38 VTAIL.n11 171.744
R90 VTAIL.n39 VTAIL.n38 171.744
R91 VTAIL.n40 VTAIL.n39 171.744
R92 VTAIL.n40 VTAIL.n7 171.744
R93 VTAIL.n47 VTAIL.n7 171.744
R94 VTAIL.n48 VTAIL.n47 171.744
R95 VTAIL.n48 VTAIL.n3 171.744
R96 VTAIL.n55 VTAIL.n3 171.744
R97 VTAIL.n56 VTAIL.n55 171.744
R98 VTAIL.n180 VTAIL.n179 171.744
R99 VTAIL.n179 VTAIL.n127 171.744
R100 VTAIL.n172 VTAIL.n127 171.744
R101 VTAIL.n172 VTAIL.n171 171.744
R102 VTAIL.n171 VTAIL.n131 171.744
R103 VTAIL.n136 VTAIL.n131 171.744
R104 VTAIL.n164 VTAIL.n136 171.744
R105 VTAIL.n164 VTAIL.n163 171.744
R106 VTAIL.n163 VTAIL.n137 171.744
R107 VTAIL.n156 VTAIL.n137 171.744
R108 VTAIL.n156 VTAIL.n155 171.744
R109 VTAIL.n155 VTAIL.n141 171.744
R110 VTAIL.n148 VTAIL.n141 171.744
R111 VTAIL.n148 VTAIL.n147 171.744
R112 VTAIL.n118 VTAIL.n117 171.744
R113 VTAIL.n117 VTAIL.n65 171.744
R114 VTAIL.n110 VTAIL.n65 171.744
R115 VTAIL.n110 VTAIL.n109 171.744
R116 VTAIL.n109 VTAIL.n69 171.744
R117 VTAIL.n74 VTAIL.n69 171.744
R118 VTAIL.n102 VTAIL.n74 171.744
R119 VTAIL.n102 VTAIL.n101 171.744
R120 VTAIL.n101 VTAIL.n75 171.744
R121 VTAIL.n94 VTAIL.n75 171.744
R122 VTAIL.n94 VTAIL.n93 171.744
R123 VTAIL.n93 VTAIL.n79 171.744
R124 VTAIL.n86 VTAIL.n79 171.744
R125 VTAIL.n86 VTAIL.n85 171.744
R126 VTAIL.n207 VTAIL.t2 85.8723
R127 VTAIL.n21 VTAIL.t0 85.8723
R128 VTAIL.n147 VTAIL.t1 85.8723
R129 VTAIL.n85 VTAIL.t3 85.8723
R130 VTAIL.n247 VTAIL.n246 31.4096
R131 VTAIL.n61 VTAIL.n60 31.4096
R132 VTAIL.n185 VTAIL.n184 31.4096
R133 VTAIL.n123 VTAIL.n122 31.4096
R134 VTAIL.n123 VTAIL.n61 25.4358
R135 VTAIL.n247 VTAIL.n185 23.7979
R136 VTAIL.n227 VTAIL.n194 13.1884
R137 VTAIL.n41 VTAIL.n8 13.1884
R138 VTAIL.n134 VTAIL.n132 13.1884
R139 VTAIL.n72 VTAIL.n70 13.1884
R140 VTAIL.n228 VTAIL.n196 12.8005
R141 VTAIL.n232 VTAIL.n231 12.8005
R142 VTAIL.n42 VTAIL.n10 12.8005
R143 VTAIL.n46 VTAIL.n45 12.8005
R144 VTAIL.n170 VTAIL.n169 12.8005
R145 VTAIL.n166 VTAIL.n165 12.8005
R146 VTAIL.n108 VTAIL.n107 12.8005
R147 VTAIL.n104 VTAIL.n103 12.8005
R148 VTAIL.n223 VTAIL.n222 12.0247
R149 VTAIL.n235 VTAIL.n192 12.0247
R150 VTAIL.n37 VTAIL.n36 12.0247
R151 VTAIL.n49 VTAIL.n6 12.0247
R152 VTAIL.n173 VTAIL.n130 12.0247
R153 VTAIL.n162 VTAIL.n135 12.0247
R154 VTAIL.n111 VTAIL.n68 12.0247
R155 VTAIL.n100 VTAIL.n73 12.0247
R156 VTAIL.n221 VTAIL.n198 11.249
R157 VTAIL.n236 VTAIL.n190 11.249
R158 VTAIL.n35 VTAIL.n12 11.249
R159 VTAIL.n50 VTAIL.n4 11.249
R160 VTAIL.n174 VTAIL.n128 11.249
R161 VTAIL.n161 VTAIL.n138 11.249
R162 VTAIL.n112 VTAIL.n66 11.249
R163 VTAIL.n99 VTAIL.n76 11.249
R164 VTAIL.n206 VTAIL.n205 10.7239
R165 VTAIL.n20 VTAIL.n19 10.7239
R166 VTAIL.n146 VTAIL.n145 10.7239
R167 VTAIL.n84 VTAIL.n83 10.7239
R168 VTAIL.n218 VTAIL.n217 10.4732
R169 VTAIL.n240 VTAIL.n239 10.4732
R170 VTAIL.n32 VTAIL.n31 10.4732
R171 VTAIL.n54 VTAIL.n53 10.4732
R172 VTAIL.n178 VTAIL.n177 10.4732
R173 VTAIL.n158 VTAIL.n157 10.4732
R174 VTAIL.n116 VTAIL.n115 10.4732
R175 VTAIL.n96 VTAIL.n95 10.4732
R176 VTAIL.n214 VTAIL.n200 9.69747
R177 VTAIL.n243 VTAIL.n188 9.69747
R178 VTAIL.n28 VTAIL.n14 9.69747
R179 VTAIL.n57 VTAIL.n2 9.69747
R180 VTAIL.n181 VTAIL.n126 9.69747
R181 VTAIL.n154 VTAIL.n140 9.69747
R182 VTAIL.n119 VTAIL.n64 9.69747
R183 VTAIL.n92 VTAIL.n78 9.69747
R184 VTAIL.n246 VTAIL.n245 9.45567
R185 VTAIL.n60 VTAIL.n59 9.45567
R186 VTAIL.n184 VTAIL.n183 9.45567
R187 VTAIL.n122 VTAIL.n121 9.45567
R188 VTAIL.n245 VTAIL.n244 9.3005
R189 VTAIL.n188 VTAIL.n187 9.3005
R190 VTAIL.n239 VTAIL.n238 9.3005
R191 VTAIL.n237 VTAIL.n236 9.3005
R192 VTAIL.n192 VTAIL.n191 9.3005
R193 VTAIL.n231 VTAIL.n230 9.3005
R194 VTAIL.n204 VTAIL.n203 9.3005
R195 VTAIL.n211 VTAIL.n210 9.3005
R196 VTAIL.n213 VTAIL.n212 9.3005
R197 VTAIL.n200 VTAIL.n199 9.3005
R198 VTAIL.n219 VTAIL.n218 9.3005
R199 VTAIL.n221 VTAIL.n220 9.3005
R200 VTAIL.n222 VTAIL.n195 9.3005
R201 VTAIL.n229 VTAIL.n228 9.3005
R202 VTAIL.n59 VTAIL.n58 9.3005
R203 VTAIL.n2 VTAIL.n1 9.3005
R204 VTAIL.n53 VTAIL.n52 9.3005
R205 VTAIL.n51 VTAIL.n50 9.3005
R206 VTAIL.n6 VTAIL.n5 9.3005
R207 VTAIL.n45 VTAIL.n44 9.3005
R208 VTAIL.n18 VTAIL.n17 9.3005
R209 VTAIL.n25 VTAIL.n24 9.3005
R210 VTAIL.n27 VTAIL.n26 9.3005
R211 VTAIL.n14 VTAIL.n13 9.3005
R212 VTAIL.n33 VTAIL.n32 9.3005
R213 VTAIL.n35 VTAIL.n34 9.3005
R214 VTAIL.n36 VTAIL.n9 9.3005
R215 VTAIL.n43 VTAIL.n42 9.3005
R216 VTAIL.n144 VTAIL.n143 9.3005
R217 VTAIL.n151 VTAIL.n150 9.3005
R218 VTAIL.n153 VTAIL.n152 9.3005
R219 VTAIL.n140 VTAIL.n139 9.3005
R220 VTAIL.n159 VTAIL.n158 9.3005
R221 VTAIL.n161 VTAIL.n160 9.3005
R222 VTAIL.n135 VTAIL.n133 9.3005
R223 VTAIL.n167 VTAIL.n166 9.3005
R224 VTAIL.n183 VTAIL.n182 9.3005
R225 VTAIL.n126 VTAIL.n125 9.3005
R226 VTAIL.n177 VTAIL.n176 9.3005
R227 VTAIL.n175 VTAIL.n174 9.3005
R228 VTAIL.n130 VTAIL.n129 9.3005
R229 VTAIL.n169 VTAIL.n168 9.3005
R230 VTAIL.n82 VTAIL.n81 9.3005
R231 VTAIL.n89 VTAIL.n88 9.3005
R232 VTAIL.n91 VTAIL.n90 9.3005
R233 VTAIL.n78 VTAIL.n77 9.3005
R234 VTAIL.n97 VTAIL.n96 9.3005
R235 VTAIL.n99 VTAIL.n98 9.3005
R236 VTAIL.n73 VTAIL.n71 9.3005
R237 VTAIL.n105 VTAIL.n104 9.3005
R238 VTAIL.n121 VTAIL.n120 9.3005
R239 VTAIL.n64 VTAIL.n63 9.3005
R240 VTAIL.n115 VTAIL.n114 9.3005
R241 VTAIL.n113 VTAIL.n112 9.3005
R242 VTAIL.n68 VTAIL.n67 9.3005
R243 VTAIL.n107 VTAIL.n106 9.3005
R244 VTAIL.n213 VTAIL.n202 8.92171
R245 VTAIL.n244 VTAIL.n186 8.92171
R246 VTAIL.n27 VTAIL.n16 8.92171
R247 VTAIL.n58 VTAIL.n0 8.92171
R248 VTAIL.n182 VTAIL.n124 8.92171
R249 VTAIL.n153 VTAIL.n142 8.92171
R250 VTAIL.n120 VTAIL.n62 8.92171
R251 VTAIL.n91 VTAIL.n80 8.92171
R252 VTAIL.n210 VTAIL.n209 8.14595
R253 VTAIL.n24 VTAIL.n23 8.14595
R254 VTAIL.n150 VTAIL.n149 8.14595
R255 VTAIL.n88 VTAIL.n87 8.14595
R256 VTAIL.n206 VTAIL.n204 7.3702
R257 VTAIL.n20 VTAIL.n18 7.3702
R258 VTAIL.n146 VTAIL.n144 7.3702
R259 VTAIL.n84 VTAIL.n82 7.3702
R260 VTAIL.n209 VTAIL.n204 5.81868
R261 VTAIL.n23 VTAIL.n18 5.81868
R262 VTAIL.n149 VTAIL.n144 5.81868
R263 VTAIL.n87 VTAIL.n82 5.81868
R264 VTAIL.n210 VTAIL.n202 5.04292
R265 VTAIL.n246 VTAIL.n186 5.04292
R266 VTAIL.n24 VTAIL.n16 5.04292
R267 VTAIL.n60 VTAIL.n0 5.04292
R268 VTAIL.n184 VTAIL.n124 5.04292
R269 VTAIL.n150 VTAIL.n142 5.04292
R270 VTAIL.n122 VTAIL.n62 5.04292
R271 VTAIL.n88 VTAIL.n80 5.04292
R272 VTAIL.n214 VTAIL.n213 4.26717
R273 VTAIL.n244 VTAIL.n243 4.26717
R274 VTAIL.n28 VTAIL.n27 4.26717
R275 VTAIL.n58 VTAIL.n57 4.26717
R276 VTAIL.n182 VTAIL.n181 4.26717
R277 VTAIL.n154 VTAIL.n153 4.26717
R278 VTAIL.n120 VTAIL.n119 4.26717
R279 VTAIL.n92 VTAIL.n91 4.26717
R280 VTAIL.n217 VTAIL.n200 3.49141
R281 VTAIL.n240 VTAIL.n188 3.49141
R282 VTAIL.n31 VTAIL.n14 3.49141
R283 VTAIL.n54 VTAIL.n2 3.49141
R284 VTAIL.n178 VTAIL.n126 3.49141
R285 VTAIL.n157 VTAIL.n140 3.49141
R286 VTAIL.n116 VTAIL.n64 3.49141
R287 VTAIL.n95 VTAIL.n78 3.49141
R288 VTAIL.n218 VTAIL.n198 2.71565
R289 VTAIL.n239 VTAIL.n190 2.71565
R290 VTAIL.n32 VTAIL.n12 2.71565
R291 VTAIL.n53 VTAIL.n4 2.71565
R292 VTAIL.n177 VTAIL.n128 2.71565
R293 VTAIL.n158 VTAIL.n138 2.71565
R294 VTAIL.n115 VTAIL.n66 2.71565
R295 VTAIL.n96 VTAIL.n76 2.71565
R296 VTAIL.n205 VTAIL.n203 2.41282
R297 VTAIL.n19 VTAIL.n17 2.41282
R298 VTAIL.n145 VTAIL.n143 2.41282
R299 VTAIL.n83 VTAIL.n81 2.41282
R300 VTAIL.n223 VTAIL.n221 1.93989
R301 VTAIL.n236 VTAIL.n235 1.93989
R302 VTAIL.n37 VTAIL.n35 1.93989
R303 VTAIL.n50 VTAIL.n49 1.93989
R304 VTAIL.n174 VTAIL.n173 1.93989
R305 VTAIL.n162 VTAIL.n161 1.93989
R306 VTAIL.n112 VTAIL.n111 1.93989
R307 VTAIL.n100 VTAIL.n99 1.93989
R308 VTAIL.n185 VTAIL.n123 1.28929
R309 VTAIL.n222 VTAIL.n196 1.16414
R310 VTAIL.n232 VTAIL.n192 1.16414
R311 VTAIL.n36 VTAIL.n10 1.16414
R312 VTAIL.n46 VTAIL.n6 1.16414
R313 VTAIL.n170 VTAIL.n130 1.16414
R314 VTAIL.n165 VTAIL.n135 1.16414
R315 VTAIL.n108 VTAIL.n68 1.16414
R316 VTAIL.n103 VTAIL.n73 1.16414
R317 VTAIL VTAIL.n61 0.938
R318 VTAIL.n228 VTAIL.n227 0.388379
R319 VTAIL.n231 VTAIL.n194 0.388379
R320 VTAIL.n42 VTAIL.n41 0.388379
R321 VTAIL.n45 VTAIL.n8 0.388379
R322 VTAIL.n169 VTAIL.n132 0.388379
R323 VTAIL.n166 VTAIL.n134 0.388379
R324 VTAIL.n107 VTAIL.n70 0.388379
R325 VTAIL.n104 VTAIL.n72 0.388379
R326 VTAIL VTAIL.n247 0.351793
R327 VTAIL.n211 VTAIL.n203 0.155672
R328 VTAIL.n212 VTAIL.n211 0.155672
R329 VTAIL.n212 VTAIL.n199 0.155672
R330 VTAIL.n219 VTAIL.n199 0.155672
R331 VTAIL.n220 VTAIL.n219 0.155672
R332 VTAIL.n220 VTAIL.n195 0.155672
R333 VTAIL.n229 VTAIL.n195 0.155672
R334 VTAIL.n230 VTAIL.n229 0.155672
R335 VTAIL.n230 VTAIL.n191 0.155672
R336 VTAIL.n237 VTAIL.n191 0.155672
R337 VTAIL.n238 VTAIL.n237 0.155672
R338 VTAIL.n238 VTAIL.n187 0.155672
R339 VTAIL.n245 VTAIL.n187 0.155672
R340 VTAIL.n25 VTAIL.n17 0.155672
R341 VTAIL.n26 VTAIL.n25 0.155672
R342 VTAIL.n26 VTAIL.n13 0.155672
R343 VTAIL.n33 VTAIL.n13 0.155672
R344 VTAIL.n34 VTAIL.n33 0.155672
R345 VTAIL.n34 VTAIL.n9 0.155672
R346 VTAIL.n43 VTAIL.n9 0.155672
R347 VTAIL.n44 VTAIL.n43 0.155672
R348 VTAIL.n44 VTAIL.n5 0.155672
R349 VTAIL.n51 VTAIL.n5 0.155672
R350 VTAIL.n52 VTAIL.n51 0.155672
R351 VTAIL.n52 VTAIL.n1 0.155672
R352 VTAIL.n59 VTAIL.n1 0.155672
R353 VTAIL.n183 VTAIL.n125 0.155672
R354 VTAIL.n176 VTAIL.n125 0.155672
R355 VTAIL.n176 VTAIL.n175 0.155672
R356 VTAIL.n175 VTAIL.n129 0.155672
R357 VTAIL.n168 VTAIL.n129 0.155672
R358 VTAIL.n168 VTAIL.n167 0.155672
R359 VTAIL.n167 VTAIL.n133 0.155672
R360 VTAIL.n160 VTAIL.n133 0.155672
R361 VTAIL.n160 VTAIL.n159 0.155672
R362 VTAIL.n159 VTAIL.n139 0.155672
R363 VTAIL.n152 VTAIL.n139 0.155672
R364 VTAIL.n152 VTAIL.n151 0.155672
R365 VTAIL.n151 VTAIL.n143 0.155672
R366 VTAIL.n121 VTAIL.n63 0.155672
R367 VTAIL.n114 VTAIL.n63 0.155672
R368 VTAIL.n114 VTAIL.n113 0.155672
R369 VTAIL.n113 VTAIL.n67 0.155672
R370 VTAIL.n106 VTAIL.n67 0.155672
R371 VTAIL.n106 VTAIL.n105 0.155672
R372 VTAIL.n105 VTAIL.n71 0.155672
R373 VTAIL.n98 VTAIL.n71 0.155672
R374 VTAIL.n98 VTAIL.n97 0.155672
R375 VTAIL.n97 VTAIL.n77 0.155672
R376 VTAIL.n90 VTAIL.n77 0.155672
R377 VTAIL.n90 VTAIL.n89 0.155672
R378 VTAIL.n89 VTAIL.n81 0.155672
R379 VDD2.n117 VDD2.n61 756.745
R380 VDD2.n56 VDD2.n0 756.745
R381 VDD2.n118 VDD2.n117 585
R382 VDD2.n116 VDD2.n115 585
R383 VDD2.n65 VDD2.n64 585
R384 VDD2.n110 VDD2.n109 585
R385 VDD2.n108 VDD2.n107 585
R386 VDD2.n69 VDD2.n68 585
R387 VDD2.n73 VDD2.n71 585
R388 VDD2.n102 VDD2.n101 585
R389 VDD2.n100 VDD2.n99 585
R390 VDD2.n75 VDD2.n74 585
R391 VDD2.n94 VDD2.n93 585
R392 VDD2.n92 VDD2.n91 585
R393 VDD2.n79 VDD2.n78 585
R394 VDD2.n86 VDD2.n85 585
R395 VDD2.n84 VDD2.n83 585
R396 VDD2.n21 VDD2.n20 585
R397 VDD2.n23 VDD2.n22 585
R398 VDD2.n16 VDD2.n15 585
R399 VDD2.n29 VDD2.n28 585
R400 VDD2.n31 VDD2.n30 585
R401 VDD2.n12 VDD2.n11 585
R402 VDD2.n38 VDD2.n37 585
R403 VDD2.n39 VDD2.n10 585
R404 VDD2.n41 VDD2.n40 585
R405 VDD2.n8 VDD2.n7 585
R406 VDD2.n47 VDD2.n46 585
R407 VDD2.n49 VDD2.n48 585
R408 VDD2.n4 VDD2.n3 585
R409 VDD2.n55 VDD2.n54 585
R410 VDD2.n57 VDD2.n56 585
R411 VDD2.n82 VDD2.t0 329.036
R412 VDD2.n19 VDD2.t1 329.036
R413 VDD2.n117 VDD2.n116 171.744
R414 VDD2.n116 VDD2.n64 171.744
R415 VDD2.n109 VDD2.n64 171.744
R416 VDD2.n109 VDD2.n108 171.744
R417 VDD2.n108 VDD2.n68 171.744
R418 VDD2.n73 VDD2.n68 171.744
R419 VDD2.n101 VDD2.n73 171.744
R420 VDD2.n101 VDD2.n100 171.744
R421 VDD2.n100 VDD2.n74 171.744
R422 VDD2.n93 VDD2.n74 171.744
R423 VDD2.n93 VDD2.n92 171.744
R424 VDD2.n92 VDD2.n78 171.744
R425 VDD2.n85 VDD2.n78 171.744
R426 VDD2.n85 VDD2.n84 171.744
R427 VDD2.n22 VDD2.n21 171.744
R428 VDD2.n22 VDD2.n15 171.744
R429 VDD2.n29 VDD2.n15 171.744
R430 VDD2.n30 VDD2.n29 171.744
R431 VDD2.n30 VDD2.n11 171.744
R432 VDD2.n38 VDD2.n11 171.744
R433 VDD2.n39 VDD2.n38 171.744
R434 VDD2.n40 VDD2.n39 171.744
R435 VDD2.n40 VDD2.n7 171.744
R436 VDD2.n47 VDD2.n7 171.744
R437 VDD2.n48 VDD2.n47 171.744
R438 VDD2.n48 VDD2.n3 171.744
R439 VDD2.n55 VDD2.n3 171.744
R440 VDD2.n56 VDD2.n55 171.744
R441 VDD2.n84 VDD2.t0 85.8723
R442 VDD2.n21 VDD2.t1 85.8723
R443 VDD2.n122 VDD2.n60 84.8168
R444 VDD2.n122 VDD2.n121 48.0884
R445 VDD2.n71 VDD2.n69 13.1884
R446 VDD2.n41 VDD2.n8 13.1884
R447 VDD2.n107 VDD2.n106 12.8005
R448 VDD2.n103 VDD2.n102 12.8005
R449 VDD2.n42 VDD2.n10 12.8005
R450 VDD2.n46 VDD2.n45 12.8005
R451 VDD2.n110 VDD2.n67 12.0247
R452 VDD2.n99 VDD2.n72 12.0247
R453 VDD2.n37 VDD2.n36 12.0247
R454 VDD2.n49 VDD2.n6 12.0247
R455 VDD2.n111 VDD2.n65 11.249
R456 VDD2.n98 VDD2.n75 11.249
R457 VDD2.n35 VDD2.n12 11.249
R458 VDD2.n50 VDD2.n4 11.249
R459 VDD2.n83 VDD2.n82 10.7239
R460 VDD2.n20 VDD2.n19 10.7239
R461 VDD2.n115 VDD2.n114 10.4732
R462 VDD2.n95 VDD2.n94 10.4732
R463 VDD2.n32 VDD2.n31 10.4732
R464 VDD2.n54 VDD2.n53 10.4732
R465 VDD2.n118 VDD2.n63 9.69747
R466 VDD2.n91 VDD2.n77 9.69747
R467 VDD2.n28 VDD2.n14 9.69747
R468 VDD2.n57 VDD2.n2 9.69747
R469 VDD2.n121 VDD2.n120 9.45567
R470 VDD2.n60 VDD2.n59 9.45567
R471 VDD2.n81 VDD2.n80 9.3005
R472 VDD2.n88 VDD2.n87 9.3005
R473 VDD2.n90 VDD2.n89 9.3005
R474 VDD2.n77 VDD2.n76 9.3005
R475 VDD2.n96 VDD2.n95 9.3005
R476 VDD2.n98 VDD2.n97 9.3005
R477 VDD2.n72 VDD2.n70 9.3005
R478 VDD2.n104 VDD2.n103 9.3005
R479 VDD2.n120 VDD2.n119 9.3005
R480 VDD2.n63 VDD2.n62 9.3005
R481 VDD2.n114 VDD2.n113 9.3005
R482 VDD2.n112 VDD2.n111 9.3005
R483 VDD2.n67 VDD2.n66 9.3005
R484 VDD2.n106 VDD2.n105 9.3005
R485 VDD2.n59 VDD2.n58 9.3005
R486 VDD2.n2 VDD2.n1 9.3005
R487 VDD2.n53 VDD2.n52 9.3005
R488 VDD2.n51 VDD2.n50 9.3005
R489 VDD2.n6 VDD2.n5 9.3005
R490 VDD2.n45 VDD2.n44 9.3005
R491 VDD2.n18 VDD2.n17 9.3005
R492 VDD2.n25 VDD2.n24 9.3005
R493 VDD2.n27 VDD2.n26 9.3005
R494 VDD2.n14 VDD2.n13 9.3005
R495 VDD2.n33 VDD2.n32 9.3005
R496 VDD2.n35 VDD2.n34 9.3005
R497 VDD2.n36 VDD2.n9 9.3005
R498 VDD2.n43 VDD2.n42 9.3005
R499 VDD2.n119 VDD2.n61 8.92171
R500 VDD2.n90 VDD2.n79 8.92171
R501 VDD2.n27 VDD2.n16 8.92171
R502 VDD2.n58 VDD2.n0 8.92171
R503 VDD2.n87 VDD2.n86 8.14595
R504 VDD2.n24 VDD2.n23 8.14595
R505 VDD2.n83 VDD2.n81 7.3702
R506 VDD2.n20 VDD2.n18 7.3702
R507 VDD2.n86 VDD2.n81 5.81868
R508 VDD2.n23 VDD2.n18 5.81868
R509 VDD2.n121 VDD2.n61 5.04292
R510 VDD2.n87 VDD2.n79 5.04292
R511 VDD2.n24 VDD2.n16 5.04292
R512 VDD2.n60 VDD2.n0 5.04292
R513 VDD2.n119 VDD2.n118 4.26717
R514 VDD2.n91 VDD2.n90 4.26717
R515 VDD2.n28 VDD2.n27 4.26717
R516 VDD2.n58 VDD2.n57 4.26717
R517 VDD2.n115 VDD2.n63 3.49141
R518 VDD2.n94 VDD2.n77 3.49141
R519 VDD2.n31 VDD2.n14 3.49141
R520 VDD2.n54 VDD2.n2 3.49141
R521 VDD2.n114 VDD2.n65 2.71565
R522 VDD2.n95 VDD2.n75 2.71565
R523 VDD2.n32 VDD2.n12 2.71565
R524 VDD2.n53 VDD2.n4 2.71565
R525 VDD2.n82 VDD2.n80 2.41282
R526 VDD2.n19 VDD2.n17 2.41282
R527 VDD2.n111 VDD2.n110 1.93989
R528 VDD2.n99 VDD2.n98 1.93989
R529 VDD2.n37 VDD2.n35 1.93989
R530 VDD2.n50 VDD2.n49 1.93989
R531 VDD2.n107 VDD2.n67 1.16414
R532 VDD2.n102 VDD2.n72 1.16414
R533 VDD2.n36 VDD2.n10 1.16414
R534 VDD2.n46 VDD2.n6 1.16414
R535 VDD2 VDD2.n122 0.468172
R536 VDD2.n106 VDD2.n69 0.388379
R537 VDD2.n103 VDD2.n71 0.388379
R538 VDD2.n42 VDD2.n41 0.388379
R539 VDD2.n45 VDD2.n8 0.388379
R540 VDD2.n120 VDD2.n62 0.155672
R541 VDD2.n113 VDD2.n62 0.155672
R542 VDD2.n113 VDD2.n112 0.155672
R543 VDD2.n112 VDD2.n66 0.155672
R544 VDD2.n105 VDD2.n66 0.155672
R545 VDD2.n105 VDD2.n104 0.155672
R546 VDD2.n104 VDD2.n70 0.155672
R547 VDD2.n97 VDD2.n70 0.155672
R548 VDD2.n97 VDD2.n96 0.155672
R549 VDD2.n96 VDD2.n76 0.155672
R550 VDD2.n89 VDD2.n76 0.155672
R551 VDD2.n89 VDD2.n88 0.155672
R552 VDD2.n88 VDD2.n80 0.155672
R553 VDD2.n25 VDD2.n17 0.155672
R554 VDD2.n26 VDD2.n25 0.155672
R555 VDD2.n26 VDD2.n13 0.155672
R556 VDD2.n33 VDD2.n13 0.155672
R557 VDD2.n34 VDD2.n33 0.155672
R558 VDD2.n34 VDD2.n9 0.155672
R559 VDD2.n43 VDD2.n9 0.155672
R560 VDD2.n44 VDD2.n43 0.155672
R561 VDD2.n44 VDD2.n5 0.155672
R562 VDD2.n51 VDD2.n5 0.155672
R563 VDD2.n52 VDD2.n51 0.155672
R564 VDD2.n52 VDD2.n1 0.155672
R565 VDD2.n59 VDD2.n1 0.155672
R566 B.n359 B.n60 585
R567 B.n361 B.n360 585
R568 B.n362 B.n59 585
R569 B.n364 B.n363 585
R570 B.n365 B.n58 585
R571 B.n367 B.n366 585
R572 B.n368 B.n57 585
R573 B.n370 B.n369 585
R574 B.n371 B.n56 585
R575 B.n373 B.n372 585
R576 B.n374 B.n55 585
R577 B.n376 B.n375 585
R578 B.n377 B.n54 585
R579 B.n379 B.n378 585
R580 B.n380 B.n53 585
R581 B.n382 B.n381 585
R582 B.n383 B.n52 585
R583 B.n385 B.n384 585
R584 B.n386 B.n51 585
R585 B.n388 B.n387 585
R586 B.n389 B.n50 585
R587 B.n391 B.n390 585
R588 B.n392 B.n49 585
R589 B.n394 B.n393 585
R590 B.n395 B.n48 585
R591 B.n397 B.n396 585
R592 B.n398 B.n47 585
R593 B.n400 B.n399 585
R594 B.n401 B.n46 585
R595 B.n403 B.n402 585
R596 B.n404 B.n45 585
R597 B.n406 B.n405 585
R598 B.n407 B.n44 585
R599 B.n409 B.n408 585
R600 B.n410 B.n43 585
R601 B.n412 B.n411 585
R602 B.n413 B.n42 585
R603 B.n415 B.n414 585
R604 B.n416 B.n41 585
R605 B.n418 B.n417 585
R606 B.n420 B.n419 585
R607 B.n421 B.n37 585
R608 B.n423 B.n422 585
R609 B.n424 B.n36 585
R610 B.n426 B.n425 585
R611 B.n427 B.n35 585
R612 B.n429 B.n428 585
R613 B.n430 B.n34 585
R614 B.n432 B.n431 585
R615 B.n434 B.n31 585
R616 B.n436 B.n435 585
R617 B.n437 B.n30 585
R618 B.n439 B.n438 585
R619 B.n440 B.n29 585
R620 B.n442 B.n441 585
R621 B.n443 B.n28 585
R622 B.n445 B.n444 585
R623 B.n446 B.n27 585
R624 B.n448 B.n447 585
R625 B.n449 B.n26 585
R626 B.n451 B.n450 585
R627 B.n452 B.n25 585
R628 B.n454 B.n453 585
R629 B.n455 B.n24 585
R630 B.n457 B.n456 585
R631 B.n458 B.n23 585
R632 B.n460 B.n459 585
R633 B.n461 B.n22 585
R634 B.n463 B.n462 585
R635 B.n464 B.n21 585
R636 B.n466 B.n465 585
R637 B.n467 B.n20 585
R638 B.n469 B.n468 585
R639 B.n470 B.n19 585
R640 B.n472 B.n471 585
R641 B.n473 B.n18 585
R642 B.n475 B.n474 585
R643 B.n476 B.n17 585
R644 B.n478 B.n477 585
R645 B.n479 B.n16 585
R646 B.n481 B.n480 585
R647 B.n482 B.n15 585
R648 B.n484 B.n483 585
R649 B.n485 B.n14 585
R650 B.n487 B.n486 585
R651 B.n488 B.n13 585
R652 B.n490 B.n489 585
R653 B.n491 B.n12 585
R654 B.n493 B.n492 585
R655 B.n358 B.n357 585
R656 B.n356 B.n61 585
R657 B.n355 B.n354 585
R658 B.n353 B.n62 585
R659 B.n352 B.n351 585
R660 B.n350 B.n63 585
R661 B.n349 B.n348 585
R662 B.n347 B.n64 585
R663 B.n346 B.n345 585
R664 B.n344 B.n65 585
R665 B.n343 B.n342 585
R666 B.n341 B.n66 585
R667 B.n340 B.n339 585
R668 B.n338 B.n67 585
R669 B.n337 B.n336 585
R670 B.n335 B.n68 585
R671 B.n334 B.n333 585
R672 B.n332 B.n69 585
R673 B.n331 B.n330 585
R674 B.n329 B.n70 585
R675 B.n328 B.n327 585
R676 B.n326 B.n71 585
R677 B.n325 B.n324 585
R678 B.n323 B.n72 585
R679 B.n322 B.n321 585
R680 B.n320 B.n73 585
R681 B.n319 B.n318 585
R682 B.n317 B.n74 585
R683 B.n316 B.n315 585
R684 B.n314 B.n75 585
R685 B.n313 B.n312 585
R686 B.n311 B.n76 585
R687 B.n310 B.n309 585
R688 B.n308 B.n77 585
R689 B.n307 B.n306 585
R690 B.n305 B.n78 585
R691 B.n304 B.n303 585
R692 B.n302 B.n79 585
R693 B.n301 B.n300 585
R694 B.n166 B.n165 585
R695 B.n167 B.n128 585
R696 B.n169 B.n168 585
R697 B.n170 B.n127 585
R698 B.n172 B.n171 585
R699 B.n173 B.n126 585
R700 B.n175 B.n174 585
R701 B.n176 B.n125 585
R702 B.n178 B.n177 585
R703 B.n179 B.n124 585
R704 B.n181 B.n180 585
R705 B.n182 B.n123 585
R706 B.n184 B.n183 585
R707 B.n185 B.n122 585
R708 B.n187 B.n186 585
R709 B.n188 B.n121 585
R710 B.n190 B.n189 585
R711 B.n191 B.n120 585
R712 B.n193 B.n192 585
R713 B.n194 B.n119 585
R714 B.n196 B.n195 585
R715 B.n197 B.n118 585
R716 B.n199 B.n198 585
R717 B.n200 B.n117 585
R718 B.n202 B.n201 585
R719 B.n203 B.n116 585
R720 B.n205 B.n204 585
R721 B.n206 B.n115 585
R722 B.n208 B.n207 585
R723 B.n209 B.n114 585
R724 B.n211 B.n210 585
R725 B.n212 B.n113 585
R726 B.n214 B.n213 585
R727 B.n215 B.n112 585
R728 B.n217 B.n216 585
R729 B.n218 B.n111 585
R730 B.n220 B.n219 585
R731 B.n221 B.n110 585
R732 B.n223 B.n222 585
R733 B.n224 B.n107 585
R734 B.n227 B.n226 585
R735 B.n228 B.n106 585
R736 B.n230 B.n229 585
R737 B.n231 B.n105 585
R738 B.n233 B.n232 585
R739 B.n234 B.n104 585
R740 B.n236 B.n235 585
R741 B.n237 B.n103 585
R742 B.n239 B.n238 585
R743 B.n241 B.n240 585
R744 B.n242 B.n99 585
R745 B.n244 B.n243 585
R746 B.n245 B.n98 585
R747 B.n247 B.n246 585
R748 B.n248 B.n97 585
R749 B.n250 B.n249 585
R750 B.n251 B.n96 585
R751 B.n253 B.n252 585
R752 B.n254 B.n95 585
R753 B.n256 B.n255 585
R754 B.n257 B.n94 585
R755 B.n259 B.n258 585
R756 B.n260 B.n93 585
R757 B.n262 B.n261 585
R758 B.n263 B.n92 585
R759 B.n265 B.n264 585
R760 B.n266 B.n91 585
R761 B.n268 B.n267 585
R762 B.n269 B.n90 585
R763 B.n271 B.n270 585
R764 B.n272 B.n89 585
R765 B.n274 B.n273 585
R766 B.n275 B.n88 585
R767 B.n277 B.n276 585
R768 B.n278 B.n87 585
R769 B.n280 B.n279 585
R770 B.n281 B.n86 585
R771 B.n283 B.n282 585
R772 B.n284 B.n85 585
R773 B.n286 B.n285 585
R774 B.n287 B.n84 585
R775 B.n289 B.n288 585
R776 B.n290 B.n83 585
R777 B.n292 B.n291 585
R778 B.n293 B.n82 585
R779 B.n295 B.n294 585
R780 B.n296 B.n81 585
R781 B.n298 B.n297 585
R782 B.n299 B.n80 585
R783 B.n164 B.n129 585
R784 B.n163 B.n162 585
R785 B.n161 B.n130 585
R786 B.n160 B.n159 585
R787 B.n158 B.n131 585
R788 B.n157 B.n156 585
R789 B.n155 B.n132 585
R790 B.n154 B.n153 585
R791 B.n152 B.n133 585
R792 B.n151 B.n150 585
R793 B.n149 B.n134 585
R794 B.n148 B.n147 585
R795 B.n146 B.n135 585
R796 B.n145 B.n144 585
R797 B.n143 B.n136 585
R798 B.n142 B.n141 585
R799 B.n140 B.n137 585
R800 B.n139 B.n138 585
R801 B.n2 B.n0 585
R802 B.n521 B.n1 585
R803 B.n520 B.n519 585
R804 B.n518 B.n3 585
R805 B.n517 B.n516 585
R806 B.n515 B.n4 585
R807 B.n514 B.n513 585
R808 B.n512 B.n5 585
R809 B.n511 B.n510 585
R810 B.n509 B.n6 585
R811 B.n508 B.n507 585
R812 B.n506 B.n7 585
R813 B.n505 B.n504 585
R814 B.n503 B.n8 585
R815 B.n502 B.n501 585
R816 B.n500 B.n9 585
R817 B.n499 B.n498 585
R818 B.n497 B.n10 585
R819 B.n496 B.n495 585
R820 B.n494 B.n11 585
R821 B.n523 B.n522 585
R822 B.n166 B.n129 550.159
R823 B.n492 B.n11 550.159
R824 B.n300 B.n299 550.159
R825 B.n359 B.n358 550.159
R826 B.n100 B.t5 400.909
R827 B.n38 B.t10 400.909
R828 B.n108 B.t8 400.909
R829 B.n32 B.t1 400.909
R830 B.n100 B.t3 380.072
R831 B.n108 B.t6 380.072
R832 B.n32 B.t0 380.072
R833 B.n38 B.t9 380.072
R834 B.n101 B.t4 364.06
R835 B.n39 B.t11 364.06
R836 B.n109 B.t7 364.06
R837 B.n33 B.t2 364.06
R838 B.n162 B.n129 163.367
R839 B.n162 B.n161 163.367
R840 B.n161 B.n160 163.367
R841 B.n160 B.n131 163.367
R842 B.n156 B.n131 163.367
R843 B.n156 B.n155 163.367
R844 B.n155 B.n154 163.367
R845 B.n154 B.n133 163.367
R846 B.n150 B.n133 163.367
R847 B.n150 B.n149 163.367
R848 B.n149 B.n148 163.367
R849 B.n148 B.n135 163.367
R850 B.n144 B.n135 163.367
R851 B.n144 B.n143 163.367
R852 B.n143 B.n142 163.367
R853 B.n142 B.n137 163.367
R854 B.n138 B.n137 163.367
R855 B.n138 B.n2 163.367
R856 B.n522 B.n2 163.367
R857 B.n522 B.n521 163.367
R858 B.n521 B.n520 163.367
R859 B.n520 B.n3 163.367
R860 B.n516 B.n3 163.367
R861 B.n516 B.n515 163.367
R862 B.n515 B.n514 163.367
R863 B.n514 B.n5 163.367
R864 B.n510 B.n5 163.367
R865 B.n510 B.n509 163.367
R866 B.n509 B.n508 163.367
R867 B.n508 B.n7 163.367
R868 B.n504 B.n7 163.367
R869 B.n504 B.n503 163.367
R870 B.n503 B.n502 163.367
R871 B.n502 B.n9 163.367
R872 B.n498 B.n9 163.367
R873 B.n498 B.n497 163.367
R874 B.n497 B.n496 163.367
R875 B.n496 B.n11 163.367
R876 B.n167 B.n166 163.367
R877 B.n168 B.n167 163.367
R878 B.n168 B.n127 163.367
R879 B.n172 B.n127 163.367
R880 B.n173 B.n172 163.367
R881 B.n174 B.n173 163.367
R882 B.n174 B.n125 163.367
R883 B.n178 B.n125 163.367
R884 B.n179 B.n178 163.367
R885 B.n180 B.n179 163.367
R886 B.n180 B.n123 163.367
R887 B.n184 B.n123 163.367
R888 B.n185 B.n184 163.367
R889 B.n186 B.n185 163.367
R890 B.n186 B.n121 163.367
R891 B.n190 B.n121 163.367
R892 B.n191 B.n190 163.367
R893 B.n192 B.n191 163.367
R894 B.n192 B.n119 163.367
R895 B.n196 B.n119 163.367
R896 B.n197 B.n196 163.367
R897 B.n198 B.n197 163.367
R898 B.n198 B.n117 163.367
R899 B.n202 B.n117 163.367
R900 B.n203 B.n202 163.367
R901 B.n204 B.n203 163.367
R902 B.n204 B.n115 163.367
R903 B.n208 B.n115 163.367
R904 B.n209 B.n208 163.367
R905 B.n210 B.n209 163.367
R906 B.n210 B.n113 163.367
R907 B.n214 B.n113 163.367
R908 B.n215 B.n214 163.367
R909 B.n216 B.n215 163.367
R910 B.n216 B.n111 163.367
R911 B.n220 B.n111 163.367
R912 B.n221 B.n220 163.367
R913 B.n222 B.n221 163.367
R914 B.n222 B.n107 163.367
R915 B.n227 B.n107 163.367
R916 B.n228 B.n227 163.367
R917 B.n229 B.n228 163.367
R918 B.n229 B.n105 163.367
R919 B.n233 B.n105 163.367
R920 B.n234 B.n233 163.367
R921 B.n235 B.n234 163.367
R922 B.n235 B.n103 163.367
R923 B.n239 B.n103 163.367
R924 B.n240 B.n239 163.367
R925 B.n240 B.n99 163.367
R926 B.n244 B.n99 163.367
R927 B.n245 B.n244 163.367
R928 B.n246 B.n245 163.367
R929 B.n246 B.n97 163.367
R930 B.n250 B.n97 163.367
R931 B.n251 B.n250 163.367
R932 B.n252 B.n251 163.367
R933 B.n252 B.n95 163.367
R934 B.n256 B.n95 163.367
R935 B.n257 B.n256 163.367
R936 B.n258 B.n257 163.367
R937 B.n258 B.n93 163.367
R938 B.n262 B.n93 163.367
R939 B.n263 B.n262 163.367
R940 B.n264 B.n263 163.367
R941 B.n264 B.n91 163.367
R942 B.n268 B.n91 163.367
R943 B.n269 B.n268 163.367
R944 B.n270 B.n269 163.367
R945 B.n270 B.n89 163.367
R946 B.n274 B.n89 163.367
R947 B.n275 B.n274 163.367
R948 B.n276 B.n275 163.367
R949 B.n276 B.n87 163.367
R950 B.n280 B.n87 163.367
R951 B.n281 B.n280 163.367
R952 B.n282 B.n281 163.367
R953 B.n282 B.n85 163.367
R954 B.n286 B.n85 163.367
R955 B.n287 B.n286 163.367
R956 B.n288 B.n287 163.367
R957 B.n288 B.n83 163.367
R958 B.n292 B.n83 163.367
R959 B.n293 B.n292 163.367
R960 B.n294 B.n293 163.367
R961 B.n294 B.n81 163.367
R962 B.n298 B.n81 163.367
R963 B.n299 B.n298 163.367
R964 B.n300 B.n79 163.367
R965 B.n304 B.n79 163.367
R966 B.n305 B.n304 163.367
R967 B.n306 B.n305 163.367
R968 B.n306 B.n77 163.367
R969 B.n310 B.n77 163.367
R970 B.n311 B.n310 163.367
R971 B.n312 B.n311 163.367
R972 B.n312 B.n75 163.367
R973 B.n316 B.n75 163.367
R974 B.n317 B.n316 163.367
R975 B.n318 B.n317 163.367
R976 B.n318 B.n73 163.367
R977 B.n322 B.n73 163.367
R978 B.n323 B.n322 163.367
R979 B.n324 B.n323 163.367
R980 B.n324 B.n71 163.367
R981 B.n328 B.n71 163.367
R982 B.n329 B.n328 163.367
R983 B.n330 B.n329 163.367
R984 B.n330 B.n69 163.367
R985 B.n334 B.n69 163.367
R986 B.n335 B.n334 163.367
R987 B.n336 B.n335 163.367
R988 B.n336 B.n67 163.367
R989 B.n340 B.n67 163.367
R990 B.n341 B.n340 163.367
R991 B.n342 B.n341 163.367
R992 B.n342 B.n65 163.367
R993 B.n346 B.n65 163.367
R994 B.n347 B.n346 163.367
R995 B.n348 B.n347 163.367
R996 B.n348 B.n63 163.367
R997 B.n352 B.n63 163.367
R998 B.n353 B.n352 163.367
R999 B.n354 B.n353 163.367
R1000 B.n354 B.n61 163.367
R1001 B.n358 B.n61 163.367
R1002 B.n492 B.n491 163.367
R1003 B.n491 B.n490 163.367
R1004 B.n490 B.n13 163.367
R1005 B.n486 B.n13 163.367
R1006 B.n486 B.n485 163.367
R1007 B.n485 B.n484 163.367
R1008 B.n484 B.n15 163.367
R1009 B.n480 B.n15 163.367
R1010 B.n480 B.n479 163.367
R1011 B.n479 B.n478 163.367
R1012 B.n478 B.n17 163.367
R1013 B.n474 B.n17 163.367
R1014 B.n474 B.n473 163.367
R1015 B.n473 B.n472 163.367
R1016 B.n472 B.n19 163.367
R1017 B.n468 B.n19 163.367
R1018 B.n468 B.n467 163.367
R1019 B.n467 B.n466 163.367
R1020 B.n466 B.n21 163.367
R1021 B.n462 B.n21 163.367
R1022 B.n462 B.n461 163.367
R1023 B.n461 B.n460 163.367
R1024 B.n460 B.n23 163.367
R1025 B.n456 B.n23 163.367
R1026 B.n456 B.n455 163.367
R1027 B.n455 B.n454 163.367
R1028 B.n454 B.n25 163.367
R1029 B.n450 B.n25 163.367
R1030 B.n450 B.n449 163.367
R1031 B.n449 B.n448 163.367
R1032 B.n448 B.n27 163.367
R1033 B.n444 B.n27 163.367
R1034 B.n444 B.n443 163.367
R1035 B.n443 B.n442 163.367
R1036 B.n442 B.n29 163.367
R1037 B.n438 B.n29 163.367
R1038 B.n438 B.n437 163.367
R1039 B.n437 B.n436 163.367
R1040 B.n436 B.n31 163.367
R1041 B.n431 B.n31 163.367
R1042 B.n431 B.n430 163.367
R1043 B.n430 B.n429 163.367
R1044 B.n429 B.n35 163.367
R1045 B.n425 B.n35 163.367
R1046 B.n425 B.n424 163.367
R1047 B.n424 B.n423 163.367
R1048 B.n423 B.n37 163.367
R1049 B.n419 B.n37 163.367
R1050 B.n419 B.n418 163.367
R1051 B.n418 B.n41 163.367
R1052 B.n414 B.n41 163.367
R1053 B.n414 B.n413 163.367
R1054 B.n413 B.n412 163.367
R1055 B.n412 B.n43 163.367
R1056 B.n408 B.n43 163.367
R1057 B.n408 B.n407 163.367
R1058 B.n407 B.n406 163.367
R1059 B.n406 B.n45 163.367
R1060 B.n402 B.n45 163.367
R1061 B.n402 B.n401 163.367
R1062 B.n401 B.n400 163.367
R1063 B.n400 B.n47 163.367
R1064 B.n396 B.n47 163.367
R1065 B.n396 B.n395 163.367
R1066 B.n395 B.n394 163.367
R1067 B.n394 B.n49 163.367
R1068 B.n390 B.n49 163.367
R1069 B.n390 B.n389 163.367
R1070 B.n389 B.n388 163.367
R1071 B.n388 B.n51 163.367
R1072 B.n384 B.n51 163.367
R1073 B.n384 B.n383 163.367
R1074 B.n383 B.n382 163.367
R1075 B.n382 B.n53 163.367
R1076 B.n378 B.n53 163.367
R1077 B.n378 B.n377 163.367
R1078 B.n377 B.n376 163.367
R1079 B.n376 B.n55 163.367
R1080 B.n372 B.n55 163.367
R1081 B.n372 B.n371 163.367
R1082 B.n371 B.n370 163.367
R1083 B.n370 B.n57 163.367
R1084 B.n366 B.n57 163.367
R1085 B.n366 B.n365 163.367
R1086 B.n365 B.n364 163.367
R1087 B.n364 B.n59 163.367
R1088 B.n360 B.n59 163.367
R1089 B.n360 B.n359 163.367
R1090 B.n102 B.n101 59.5399
R1091 B.n225 B.n109 59.5399
R1092 B.n433 B.n33 59.5399
R1093 B.n40 B.n39 59.5399
R1094 B.n101 B.n100 36.849
R1095 B.n109 B.n108 36.849
R1096 B.n33 B.n32 36.849
R1097 B.n39 B.n38 36.849
R1098 B.n494 B.n493 35.7468
R1099 B.n357 B.n60 35.7468
R1100 B.n301 B.n80 35.7468
R1101 B.n165 B.n164 35.7468
R1102 B B.n523 18.0485
R1103 B.n493 B.n12 10.6151
R1104 B.n489 B.n12 10.6151
R1105 B.n489 B.n488 10.6151
R1106 B.n488 B.n487 10.6151
R1107 B.n487 B.n14 10.6151
R1108 B.n483 B.n14 10.6151
R1109 B.n483 B.n482 10.6151
R1110 B.n482 B.n481 10.6151
R1111 B.n481 B.n16 10.6151
R1112 B.n477 B.n16 10.6151
R1113 B.n477 B.n476 10.6151
R1114 B.n476 B.n475 10.6151
R1115 B.n475 B.n18 10.6151
R1116 B.n471 B.n18 10.6151
R1117 B.n471 B.n470 10.6151
R1118 B.n470 B.n469 10.6151
R1119 B.n469 B.n20 10.6151
R1120 B.n465 B.n20 10.6151
R1121 B.n465 B.n464 10.6151
R1122 B.n464 B.n463 10.6151
R1123 B.n463 B.n22 10.6151
R1124 B.n459 B.n22 10.6151
R1125 B.n459 B.n458 10.6151
R1126 B.n458 B.n457 10.6151
R1127 B.n457 B.n24 10.6151
R1128 B.n453 B.n24 10.6151
R1129 B.n453 B.n452 10.6151
R1130 B.n452 B.n451 10.6151
R1131 B.n451 B.n26 10.6151
R1132 B.n447 B.n26 10.6151
R1133 B.n447 B.n446 10.6151
R1134 B.n446 B.n445 10.6151
R1135 B.n445 B.n28 10.6151
R1136 B.n441 B.n28 10.6151
R1137 B.n441 B.n440 10.6151
R1138 B.n440 B.n439 10.6151
R1139 B.n439 B.n30 10.6151
R1140 B.n435 B.n30 10.6151
R1141 B.n435 B.n434 10.6151
R1142 B.n432 B.n34 10.6151
R1143 B.n428 B.n34 10.6151
R1144 B.n428 B.n427 10.6151
R1145 B.n427 B.n426 10.6151
R1146 B.n426 B.n36 10.6151
R1147 B.n422 B.n36 10.6151
R1148 B.n422 B.n421 10.6151
R1149 B.n421 B.n420 10.6151
R1150 B.n417 B.n416 10.6151
R1151 B.n416 B.n415 10.6151
R1152 B.n415 B.n42 10.6151
R1153 B.n411 B.n42 10.6151
R1154 B.n411 B.n410 10.6151
R1155 B.n410 B.n409 10.6151
R1156 B.n409 B.n44 10.6151
R1157 B.n405 B.n44 10.6151
R1158 B.n405 B.n404 10.6151
R1159 B.n404 B.n403 10.6151
R1160 B.n403 B.n46 10.6151
R1161 B.n399 B.n46 10.6151
R1162 B.n399 B.n398 10.6151
R1163 B.n398 B.n397 10.6151
R1164 B.n397 B.n48 10.6151
R1165 B.n393 B.n48 10.6151
R1166 B.n393 B.n392 10.6151
R1167 B.n392 B.n391 10.6151
R1168 B.n391 B.n50 10.6151
R1169 B.n387 B.n50 10.6151
R1170 B.n387 B.n386 10.6151
R1171 B.n386 B.n385 10.6151
R1172 B.n385 B.n52 10.6151
R1173 B.n381 B.n52 10.6151
R1174 B.n381 B.n380 10.6151
R1175 B.n380 B.n379 10.6151
R1176 B.n379 B.n54 10.6151
R1177 B.n375 B.n54 10.6151
R1178 B.n375 B.n374 10.6151
R1179 B.n374 B.n373 10.6151
R1180 B.n373 B.n56 10.6151
R1181 B.n369 B.n56 10.6151
R1182 B.n369 B.n368 10.6151
R1183 B.n368 B.n367 10.6151
R1184 B.n367 B.n58 10.6151
R1185 B.n363 B.n58 10.6151
R1186 B.n363 B.n362 10.6151
R1187 B.n362 B.n361 10.6151
R1188 B.n361 B.n60 10.6151
R1189 B.n302 B.n301 10.6151
R1190 B.n303 B.n302 10.6151
R1191 B.n303 B.n78 10.6151
R1192 B.n307 B.n78 10.6151
R1193 B.n308 B.n307 10.6151
R1194 B.n309 B.n308 10.6151
R1195 B.n309 B.n76 10.6151
R1196 B.n313 B.n76 10.6151
R1197 B.n314 B.n313 10.6151
R1198 B.n315 B.n314 10.6151
R1199 B.n315 B.n74 10.6151
R1200 B.n319 B.n74 10.6151
R1201 B.n320 B.n319 10.6151
R1202 B.n321 B.n320 10.6151
R1203 B.n321 B.n72 10.6151
R1204 B.n325 B.n72 10.6151
R1205 B.n326 B.n325 10.6151
R1206 B.n327 B.n326 10.6151
R1207 B.n327 B.n70 10.6151
R1208 B.n331 B.n70 10.6151
R1209 B.n332 B.n331 10.6151
R1210 B.n333 B.n332 10.6151
R1211 B.n333 B.n68 10.6151
R1212 B.n337 B.n68 10.6151
R1213 B.n338 B.n337 10.6151
R1214 B.n339 B.n338 10.6151
R1215 B.n339 B.n66 10.6151
R1216 B.n343 B.n66 10.6151
R1217 B.n344 B.n343 10.6151
R1218 B.n345 B.n344 10.6151
R1219 B.n345 B.n64 10.6151
R1220 B.n349 B.n64 10.6151
R1221 B.n350 B.n349 10.6151
R1222 B.n351 B.n350 10.6151
R1223 B.n351 B.n62 10.6151
R1224 B.n355 B.n62 10.6151
R1225 B.n356 B.n355 10.6151
R1226 B.n357 B.n356 10.6151
R1227 B.n165 B.n128 10.6151
R1228 B.n169 B.n128 10.6151
R1229 B.n170 B.n169 10.6151
R1230 B.n171 B.n170 10.6151
R1231 B.n171 B.n126 10.6151
R1232 B.n175 B.n126 10.6151
R1233 B.n176 B.n175 10.6151
R1234 B.n177 B.n176 10.6151
R1235 B.n177 B.n124 10.6151
R1236 B.n181 B.n124 10.6151
R1237 B.n182 B.n181 10.6151
R1238 B.n183 B.n182 10.6151
R1239 B.n183 B.n122 10.6151
R1240 B.n187 B.n122 10.6151
R1241 B.n188 B.n187 10.6151
R1242 B.n189 B.n188 10.6151
R1243 B.n189 B.n120 10.6151
R1244 B.n193 B.n120 10.6151
R1245 B.n194 B.n193 10.6151
R1246 B.n195 B.n194 10.6151
R1247 B.n195 B.n118 10.6151
R1248 B.n199 B.n118 10.6151
R1249 B.n200 B.n199 10.6151
R1250 B.n201 B.n200 10.6151
R1251 B.n201 B.n116 10.6151
R1252 B.n205 B.n116 10.6151
R1253 B.n206 B.n205 10.6151
R1254 B.n207 B.n206 10.6151
R1255 B.n207 B.n114 10.6151
R1256 B.n211 B.n114 10.6151
R1257 B.n212 B.n211 10.6151
R1258 B.n213 B.n212 10.6151
R1259 B.n213 B.n112 10.6151
R1260 B.n217 B.n112 10.6151
R1261 B.n218 B.n217 10.6151
R1262 B.n219 B.n218 10.6151
R1263 B.n219 B.n110 10.6151
R1264 B.n223 B.n110 10.6151
R1265 B.n224 B.n223 10.6151
R1266 B.n226 B.n106 10.6151
R1267 B.n230 B.n106 10.6151
R1268 B.n231 B.n230 10.6151
R1269 B.n232 B.n231 10.6151
R1270 B.n232 B.n104 10.6151
R1271 B.n236 B.n104 10.6151
R1272 B.n237 B.n236 10.6151
R1273 B.n238 B.n237 10.6151
R1274 B.n242 B.n241 10.6151
R1275 B.n243 B.n242 10.6151
R1276 B.n243 B.n98 10.6151
R1277 B.n247 B.n98 10.6151
R1278 B.n248 B.n247 10.6151
R1279 B.n249 B.n248 10.6151
R1280 B.n249 B.n96 10.6151
R1281 B.n253 B.n96 10.6151
R1282 B.n254 B.n253 10.6151
R1283 B.n255 B.n254 10.6151
R1284 B.n255 B.n94 10.6151
R1285 B.n259 B.n94 10.6151
R1286 B.n260 B.n259 10.6151
R1287 B.n261 B.n260 10.6151
R1288 B.n261 B.n92 10.6151
R1289 B.n265 B.n92 10.6151
R1290 B.n266 B.n265 10.6151
R1291 B.n267 B.n266 10.6151
R1292 B.n267 B.n90 10.6151
R1293 B.n271 B.n90 10.6151
R1294 B.n272 B.n271 10.6151
R1295 B.n273 B.n272 10.6151
R1296 B.n273 B.n88 10.6151
R1297 B.n277 B.n88 10.6151
R1298 B.n278 B.n277 10.6151
R1299 B.n279 B.n278 10.6151
R1300 B.n279 B.n86 10.6151
R1301 B.n283 B.n86 10.6151
R1302 B.n284 B.n283 10.6151
R1303 B.n285 B.n284 10.6151
R1304 B.n285 B.n84 10.6151
R1305 B.n289 B.n84 10.6151
R1306 B.n290 B.n289 10.6151
R1307 B.n291 B.n290 10.6151
R1308 B.n291 B.n82 10.6151
R1309 B.n295 B.n82 10.6151
R1310 B.n296 B.n295 10.6151
R1311 B.n297 B.n296 10.6151
R1312 B.n297 B.n80 10.6151
R1313 B.n164 B.n163 10.6151
R1314 B.n163 B.n130 10.6151
R1315 B.n159 B.n130 10.6151
R1316 B.n159 B.n158 10.6151
R1317 B.n158 B.n157 10.6151
R1318 B.n157 B.n132 10.6151
R1319 B.n153 B.n132 10.6151
R1320 B.n153 B.n152 10.6151
R1321 B.n152 B.n151 10.6151
R1322 B.n151 B.n134 10.6151
R1323 B.n147 B.n134 10.6151
R1324 B.n147 B.n146 10.6151
R1325 B.n146 B.n145 10.6151
R1326 B.n145 B.n136 10.6151
R1327 B.n141 B.n136 10.6151
R1328 B.n141 B.n140 10.6151
R1329 B.n140 B.n139 10.6151
R1330 B.n139 B.n0 10.6151
R1331 B.n519 B.n1 10.6151
R1332 B.n519 B.n518 10.6151
R1333 B.n518 B.n517 10.6151
R1334 B.n517 B.n4 10.6151
R1335 B.n513 B.n4 10.6151
R1336 B.n513 B.n512 10.6151
R1337 B.n512 B.n511 10.6151
R1338 B.n511 B.n6 10.6151
R1339 B.n507 B.n6 10.6151
R1340 B.n507 B.n506 10.6151
R1341 B.n506 B.n505 10.6151
R1342 B.n505 B.n8 10.6151
R1343 B.n501 B.n8 10.6151
R1344 B.n501 B.n500 10.6151
R1345 B.n500 B.n499 10.6151
R1346 B.n499 B.n10 10.6151
R1347 B.n495 B.n10 10.6151
R1348 B.n495 B.n494 10.6151
R1349 B.n433 B.n432 6.5566
R1350 B.n420 B.n40 6.5566
R1351 B.n226 B.n225 6.5566
R1352 B.n238 B.n102 6.5566
R1353 B.n434 B.n433 4.05904
R1354 B.n417 B.n40 4.05904
R1355 B.n225 B.n224 4.05904
R1356 B.n241 B.n102 4.05904
R1357 B.n523 B.n0 2.81026
R1358 B.n523 B.n1 2.81026
R1359 VP.n0 VP.t1 321.445
R1360 VP.n0 VP.t0 280.005
R1361 VP VP.n0 0.146778
R1362 VDD1.n56 VDD1.n0 756.745
R1363 VDD1.n117 VDD1.n61 756.745
R1364 VDD1.n57 VDD1.n56 585
R1365 VDD1.n55 VDD1.n54 585
R1366 VDD1.n4 VDD1.n3 585
R1367 VDD1.n49 VDD1.n48 585
R1368 VDD1.n47 VDD1.n46 585
R1369 VDD1.n8 VDD1.n7 585
R1370 VDD1.n12 VDD1.n10 585
R1371 VDD1.n41 VDD1.n40 585
R1372 VDD1.n39 VDD1.n38 585
R1373 VDD1.n14 VDD1.n13 585
R1374 VDD1.n33 VDD1.n32 585
R1375 VDD1.n31 VDD1.n30 585
R1376 VDD1.n18 VDD1.n17 585
R1377 VDD1.n25 VDD1.n24 585
R1378 VDD1.n23 VDD1.n22 585
R1379 VDD1.n82 VDD1.n81 585
R1380 VDD1.n84 VDD1.n83 585
R1381 VDD1.n77 VDD1.n76 585
R1382 VDD1.n90 VDD1.n89 585
R1383 VDD1.n92 VDD1.n91 585
R1384 VDD1.n73 VDD1.n72 585
R1385 VDD1.n99 VDD1.n98 585
R1386 VDD1.n100 VDD1.n71 585
R1387 VDD1.n102 VDD1.n101 585
R1388 VDD1.n69 VDD1.n68 585
R1389 VDD1.n108 VDD1.n107 585
R1390 VDD1.n110 VDD1.n109 585
R1391 VDD1.n65 VDD1.n64 585
R1392 VDD1.n116 VDD1.n115 585
R1393 VDD1.n118 VDD1.n117 585
R1394 VDD1.n21 VDD1.t0 329.036
R1395 VDD1.n80 VDD1.t1 329.036
R1396 VDD1.n56 VDD1.n55 171.744
R1397 VDD1.n55 VDD1.n3 171.744
R1398 VDD1.n48 VDD1.n3 171.744
R1399 VDD1.n48 VDD1.n47 171.744
R1400 VDD1.n47 VDD1.n7 171.744
R1401 VDD1.n12 VDD1.n7 171.744
R1402 VDD1.n40 VDD1.n12 171.744
R1403 VDD1.n40 VDD1.n39 171.744
R1404 VDD1.n39 VDD1.n13 171.744
R1405 VDD1.n32 VDD1.n13 171.744
R1406 VDD1.n32 VDD1.n31 171.744
R1407 VDD1.n31 VDD1.n17 171.744
R1408 VDD1.n24 VDD1.n17 171.744
R1409 VDD1.n24 VDD1.n23 171.744
R1410 VDD1.n83 VDD1.n82 171.744
R1411 VDD1.n83 VDD1.n76 171.744
R1412 VDD1.n90 VDD1.n76 171.744
R1413 VDD1.n91 VDD1.n90 171.744
R1414 VDD1.n91 VDD1.n72 171.744
R1415 VDD1.n99 VDD1.n72 171.744
R1416 VDD1.n100 VDD1.n99 171.744
R1417 VDD1.n101 VDD1.n100 171.744
R1418 VDD1.n101 VDD1.n68 171.744
R1419 VDD1.n108 VDD1.n68 171.744
R1420 VDD1.n109 VDD1.n108 171.744
R1421 VDD1.n109 VDD1.n64 171.744
R1422 VDD1.n116 VDD1.n64 171.744
R1423 VDD1.n117 VDD1.n116 171.744
R1424 VDD1.n23 VDD1.t0 85.8723
R1425 VDD1.n82 VDD1.t1 85.8723
R1426 VDD1 VDD1.n121 85.7511
R1427 VDD1 VDD1.n60 48.556
R1428 VDD1.n10 VDD1.n8 13.1884
R1429 VDD1.n102 VDD1.n69 13.1884
R1430 VDD1.n46 VDD1.n45 12.8005
R1431 VDD1.n42 VDD1.n41 12.8005
R1432 VDD1.n103 VDD1.n71 12.8005
R1433 VDD1.n107 VDD1.n106 12.8005
R1434 VDD1.n49 VDD1.n6 12.0247
R1435 VDD1.n38 VDD1.n11 12.0247
R1436 VDD1.n98 VDD1.n97 12.0247
R1437 VDD1.n110 VDD1.n67 12.0247
R1438 VDD1.n50 VDD1.n4 11.249
R1439 VDD1.n37 VDD1.n14 11.249
R1440 VDD1.n96 VDD1.n73 11.249
R1441 VDD1.n111 VDD1.n65 11.249
R1442 VDD1.n22 VDD1.n21 10.7239
R1443 VDD1.n81 VDD1.n80 10.7239
R1444 VDD1.n54 VDD1.n53 10.4732
R1445 VDD1.n34 VDD1.n33 10.4732
R1446 VDD1.n93 VDD1.n92 10.4732
R1447 VDD1.n115 VDD1.n114 10.4732
R1448 VDD1.n57 VDD1.n2 9.69747
R1449 VDD1.n30 VDD1.n16 9.69747
R1450 VDD1.n89 VDD1.n75 9.69747
R1451 VDD1.n118 VDD1.n63 9.69747
R1452 VDD1.n60 VDD1.n59 9.45567
R1453 VDD1.n121 VDD1.n120 9.45567
R1454 VDD1.n20 VDD1.n19 9.3005
R1455 VDD1.n27 VDD1.n26 9.3005
R1456 VDD1.n29 VDD1.n28 9.3005
R1457 VDD1.n16 VDD1.n15 9.3005
R1458 VDD1.n35 VDD1.n34 9.3005
R1459 VDD1.n37 VDD1.n36 9.3005
R1460 VDD1.n11 VDD1.n9 9.3005
R1461 VDD1.n43 VDD1.n42 9.3005
R1462 VDD1.n59 VDD1.n58 9.3005
R1463 VDD1.n2 VDD1.n1 9.3005
R1464 VDD1.n53 VDD1.n52 9.3005
R1465 VDD1.n51 VDD1.n50 9.3005
R1466 VDD1.n6 VDD1.n5 9.3005
R1467 VDD1.n45 VDD1.n44 9.3005
R1468 VDD1.n120 VDD1.n119 9.3005
R1469 VDD1.n63 VDD1.n62 9.3005
R1470 VDD1.n114 VDD1.n113 9.3005
R1471 VDD1.n112 VDD1.n111 9.3005
R1472 VDD1.n67 VDD1.n66 9.3005
R1473 VDD1.n106 VDD1.n105 9.3005
R1474 VDD1.n79 VDD1.n78 9.3005
R1475 VDD1.n86 VDD1.n85 9.3005
R1476 VDD1.n88 VDD1.n87 9.3005
R1477 VDD1.n75 VDD1.n74 9.3005
R1478 VDD1.n94 VDD1.n93 9.3005
R1479 VDD1.n96 VDD1.n95 9.3005
R1480 VDD1.n97 VDD1.n70 9.3005
R1481 VDD1.n104 VDD1.n103 9.3005
R1482 VDD1.n58 VDD1.n0 8.92171
R1483 VDD1.n29 VDD1.n18 8.92171
R1484 VDD1.n88 VDD1.n77 8.92171
R1485 VDD1.n119 VDD1.n61 8.92171
R1486 VDD1.n26 VDD1.n25 8.14595
R1487 VDD1.n85 VDD1.n84 8.14595
R1488 VDD1.n22 VDD1.n20 7.3702
R1489 VDD1.n81 VDD1.n79 7.3702
R1490 VDD1.n25 VDD1.n20 5.81868
R1491 VDD1.n84 VDD1.n79 5.81868
R1492 VDD1.n60 VDD1.n0 5.04292
R1493 VDD1.n26 VDD1.n18 5.04292
R1494 VDD1.n85 VDD1.n77 5.04292
R1495 VDD1.n121 VDD1.n61 5.04292
R1496 VDD1.n58 VDD1.n57 4.26717
R1497 VDD1.n30 VDD1.n29 4.26717
R1498 VDD1.n89 VDD1.n88 4.26717
R1499 VDD1.n119 VDD1.n118 4.26717
R1500 VDD1.n54 VDD1.n2 3.49141
R1501 VDD1.n33 VDD1.n16 3.49141
R1502 VDD1.n92 VDD1.n75 3.49141
R1503 VDD1.n115 VDD1.n63 3.49141
R1504 VDD1.n53 VDD1.n4 2.71565
R1505 VDD1.n34 VDD1.n14 2.71565
R1506 VDD1.n93 VDD1.n73 2.71565
R1507 VDD1.n114 VDD1.n65 2.71565
R1508 VDD1.n21 VDD1.n19 2.41282
R1509 VDD1.n80 VDD1.n78 2.41282
R1510 VDD1.n50 VDD1.n49 1.93989
R1511 VDD1.n38 VDD1.n37 1.93989
R1512 VDD1.n98 VDD1.n96 1.93989
R1513 VDD1.n111 VDD1.n110 1.93989
R1514 VDD1.n46 VDD1.n6 1.16414
R1515 VDD1.n41 VDD1.n11 1.16414
R1516 VDD1.n97 VDD1.n71 1.16414
R1517 VDD1.n107 VDD1.n67 1.16414
R1518 VDD1.n45 VDD1.n8 0.388379
R1519 VDD1.n42 VDD1.n10 0.388379
R1520 VDD1.n103 VDD1.n102 0.388379
R1521 VDD1.n106 VDD1.n69 0.388379
R1522 VDD1.n59 VDD1.n1 0.155672
R1523 VDD1.n52 VDD1.n1 0.155672
R1524 VDD1.n52 VDD1.n51 0.155672
R1525 VDD1.n51 VDD1.n5 0.155672
R1526 VDD1.n44 VDD1.n5 0.155672
R1527 VDD1.n44 VDD1.n43 0.155672
R1528 VDD1.n43 VDD1.n9 0.155672
R1529 VDD1.n36 VDD1.n9 0.155672
R1530 VDD1.n36 VDD1.n35 0.155672
R1531 VDD1.n35 VDD1.n15 0.155672
R1532 VDD1.n28 VDD1.n15 0.155672
R1533 VDD1.n28 VDD1.n27 0.155672
R1534 VDD1.n27 VDD1.n19 0.155672
R1535 VDD1.n86 VDD1.n78 0.155672
R1536 VDD1.n87 VDD1.n86 0.155672
R1537 VDD1.n87 VDD1.n74 0.155672
R1538 VDD1.n94 VDD1.n74 0.155672
R1539 VDD1.n95 VDD1.n94 0.155672
R1540 VDD1.n95 VDD1.n70 0.155672
R1541 VDD1.n104 VDD1.n70 0.155672
R1542 VDD1.n105 VDD1.n104 0.155672
R1543 VDD1.n105 VDD1.n66 0.155672
R1544 VDD1.n112 VDD1.n66 0.155672
R1545 VDD1.n113 VDD1.n112 0.155672
R1546 VDD1.n113 VDD1.n62 0.155672
R1547 VDD1.n120 VDD1.n62 0.155672
C0 VDD1 VP 2.54219f
C1 VN w_n1730_n3240# 2.27637f
C2 VN B 0.87122f
C3 w_n1730_n3240# B 7.51614f
C4 VTAIL VP 2.04315f
C5 VDD2 VDD1 0.553925f
C6 VN VP 4.84762f
C7 w_n1730_n3240# VP 2.49452f
C8 VDD2 VTAIL 4.90609f
C9 B VP 1.22573f
C10 VN VDD2 2.40309f
C11 VDD2 w_n1730_n3240# 1.63428f
C12 VTAIL VDD1 4.86369f
C13 VDD2 B 1.53122f
C14 VN VDD1 0.147984f
C15 w_n1730_n3240# VDD1 1.62072f
C16 VDD2 VP 0.290179f
C17 VDD1 B 1.51024f
C18 VN VTAIL 2.02876f
C19 w_n1730_n3240# VTAIL 2.69322f
C20 VTAIL B 3.06148f
C21 VDD2 VSUBS 0.787717f
C22 VDD1 VSUBS 3.290816f
C23 VTAIL VSUBS 0.864945f
C24 VN VSUBS 7.36076f
C25 VP VSUBS 1.349382f
C26 B VSUBS 3.077708f
C27 w_n1730_n3240# VSUBS 69.068504f
C28 VDD1.n0 VSUBS 0.021521f
C29 VDD1.n1 VSUBS 0.02029f
C30 VDD1.n2 VSUBS 0.010903f
C31 VDD1.n3 VSUBS 0.025771f
C32 VDD1.n4 VSUBS 0.011544f
C33 VDD1.n5 VSUBS 0.02029f
C34 VDD1.n6 VSUBS 0.010903f
C35 VDD1.n7 VSUBS 0.025771f
C36 VDD1.n8 VSUBS 0.011224f
C37 VDD1.n9 VSUBS 0.02029f
C38 VDD1.n10 VSUBS 0.011224f
C39 VDD1.n11 VSUBS 0.010903f
C40 VDD1.n12 VSUBS 0.025771f
C41 VDD1.n13 VSUBS 0.025771f
C42 VDD1.n14 VSUBS 0.011544f
C43 VDD1.n15 VSUBS 0.02029f
C44 VDD1.n16 VSUBS 0.010903f
C45 VDD1.n17 VSUBS 0.025771f
C46 VDD1.n18 VSUBS 0.011544f
C47 VDD1.n19 VSUBS 0.940008f
C48 VDD1.n20 VSUBS 0.010903f
C49 VDD1.t0 VSUBS 0.055491f
C50 VDD1.n21 VSUBS 0.153925f
C51 VDD1.n22 VSUBS 0.019386f
C52 VDD1.n23 VSUBS 0.019328f
C53 VDD1.n24 VSUBS 0.025771f
C54 VDD1.n25 VSUBS 0.011544f
C55 VDD1.n26 VSUBS 0.010903f
C56 VDD1.n27 VSUBS 0.02029f
C57 VDD1.n28 VSUBS 0.02029f
C58 VDD1.n29 VSUBS 0.010903f
C59 VDD1.n30 VSUBS 0.011544f
C60 VDD1.n31 VSUBS 0.025771f
C61 VDD1.n32 VSUBS 0.025771f
C62 VDD1.n33 VSUBS 0.011544f
C63 VDD1.n34 VSUBS 0.010903f
C64 VDD1.n35 VSUBS 0.02029f
C65 VDD1.n36 VSUBS 0.02029f
C66 VDD1.n37 VSUBS 0.010903f
C67 VDD1.n38 VSUBS 0.011544f
C68 VDD1.n39 VSUBS 0.025771f
C69 VDD1.n40 VSUBS 0.025771f
C70 VDD1.n41 VSUBS 0.011544f
C71 VDD1.n42 VSUBS 0.010903f
C72 VDD1.n43 VSUBS 0.02029f
C73 VDD1.n44 VSUBS 0.02029f
C74 VDD1.n45 VSUBS 0.010903f
C75 VDD1.n46 VSUBS 0.011544f
C76 VDD1.n47 VSUBS 0.025771f
C77 VDD1.n48 VSUBS 0.025771f
C78 VDD1.n49 VSUBS 0.011544f
C79 VDD1.n50 VSUBS 0.010903f
C80 VDD1.n51 VSUBS 0.02029f
C81 VDD1.n52 VSUBS 0.02029f
C82 VDD1.n53 VSUBS 0.010903f
C83 VDD1.n54 VSUBS 0.011544f
C84 VDD1.n55 VSUBS 0.025771f
C85 VDD1.n56 VSUBS 0.059755f
C86 VDD1.n57 VSUBS 0.011544f
C87 VDD1.n58 VSUBS 0.010903f
C88 VDD1.n59 VSUBS 0.045791f
C89 VDD1.n60 VSUBS 0.044582f
C90 VDD1.n61 VSUBS 0.021521f
C91 VDD1.n62 VSUBS 0.02029f
C92 VDD1.n63 VSUBS 0.010903f
C93 VDD1.n64 VSUBS 0.025771f
C94 VDD1.n65 VSUBS 0.011544f
C95 VDD1.n66 VSUBS 0.02029f
C96 VDD1.n67 VSUBS 0.010903f
C97 VDD1.n68 VSUBS 0.025771f
C98 VDD1.n69 VSUBS 0.011224f
C99 VDD1.n70 VSUBS 0.02029f
C100 VDD1.n71 VSUBS 0.011544f
C101 VDD1.n72 VSUBS 0.025771f
C102 VDD1.n73 VSUBS 0.011544f
C103 VDD1.n74 VSUBS 0.02029f
C104 VDD1.n75 VSUBS 0.010903f
C105 VDD1.n76 VSUBS 0.025771f
C106 VDD1.n77 VSUBS 0.011544f
C107 VDD1.n78 VSUBS 0.940008f
C108 VDD1.n79 VSUBS 0.010903f
C109 VDD1.t1 VSUBS 0.055491f
C110 VDD1.n80 VSUBS 0.153925f
C111 VDD1.n81 VSUBS 0.019386f
C112 VDD1.n82 VSUBS 0.019328f
C113 VDD1.n83 VSUBS 0.025771f
C114 VDD1.n84 VSUBS 0.011544f
C115 VDD1.n85 VSUBS 0.010903f
C116 VDD1.n86 VSUBS 0.02029f
C117 VDD1.n87 VSUBS 0.02029f
C118 VDD1.n88 VSUBS 0.010903f
C119 VDD1.n89 VSUBS 0.011544f
C120 VDD1.n90 VSUBS 0.025771f
C121 VDD1.n91 VSUBS 0.025771f
C122 VDD1.n92 VSUBS 0.011544f
C123 VDD1.n93 VSUBS 0.010903f
C124 VDD1.n94 VSUBS 0.02029f
C125 VDD1.n95 VSUBS 0.02029f
C126 VDD1.n96 VSUBS 0.010903f
C127 VDD1.n97 VSUBS 0.010903f
C128 VDD1.n98 VSUBS 0.011544f
C129 VDD1.n99 VSUBS 0.025771f
C130 VDD1.n100 VSUBS 0.025771f
C131 VDD1.n101 VSUBS 0.025771f
C132 VDD1.n102 VSUBS 0.011224f
C133 VDD1.n103 VSUBS 0.010903f
C134 VDD1.n104 VSUBS 0.02029f
C135 VDD1.n105 VSUBS 0.02029f
C136 VDD1.n106 VSUBS 0.010903f
C137 VDD1.n107 VSUBS 0.011544f
C138 VDD1.n108 VSUBS 0.025771f
C139 VDD1.n109 VSUBS 0.025771f
C140 VDD1.n110 VSUBS 0.011544f
C141 VDD1.n111 VSUBS 0.010903f
C142 VDD1.n112 VSUBS 0.02029f
C143 VDD1.n113 VSUBS 0.02029f
C144 VDD1.n114 VSUBS 0.010903f
C145 VDD1.n115 VSUBS 0.011544f
C146 VDD1.n116 VSUBS 0.025771f
C147 VDD1.n117 VSUBS 0.059755f
C148 VDD1.n118 VSUBS 0.011544f
C149 VDD1.n119 VSUBS 0.010903f
C150 VDD1.n120 VSUBS 0.045791f
C151 VDD1.n121 VSUBS 0.56014f
C152 VP.t1 VSUBS 3.34006f
C153 VP.t0 VSUBS 2.96456f
C154 VP.n0 VSUBS 5.43887f
C155 B.n0 VSUBS 0.004295f
C156 B.n1 VSUBS 0.004295f
C157 B.n2 VSUBS 0.006792f
C158 B.n3 VSUBS 0.006792f
C159 B.n4 VSUBS 0.006792f
C160 B.n5 VSUBS 0.006792f
C161 B.n6 VSUBS 0.006792f
C162 B.n7 VSUBS 0.006792f
C163 B.n8 VSUBS 0.006792f
C164 B.n9 VSUBS 0.006792f
C165 B.n10 VSUBS 0.006792f
C166 B.n11 VSUBS 0.01637f
C167 B.n12 VSUBS 0.006792f
C168 B.n13 VSUBS 0.006792f
C169 B.n14 VSUBS 0.006792f
C170 B.n15 VSUBS 0.006792f
C171 B.n16 VSUBS 0.006792f
C172 B.n17 VSUBS 0.006792f
C173 B.n18 VSUBS 0.006792f
C174 B.n19 VSUBS 0.006792f
C175 B.n20 VSUBS 0.006792f
C176 B.n21 VSUBS 0.006792f
C177 B.n22 VSUBS 0.006792f
C178 B.n23 VSUBS 0.006792f
C179 B.n24 VSUBS 0.006792f
C180 B.n25 VSUBS 0.006792f
C181 B.n26 VSUBS 0.006792f
C182 B.n27 VSUBS 0.006792f
C183 B.n28 VSUBS 0.006792f
C184 B.n29 VSUBS 0.006792f
C185 B.n30 VSUBS 0.006792f
C186 B.n31 VSUBS 0.006792f
C187 B.t2 VSUBS 0.190972f
C188 B.t1 VSUBS 0.211363f
C189 B.t0 VSUBS 0.762487f
C190 B.n32 VSUBS 0.328533f
C191 B.n33 VSUBS 0.231538f
C192 B.n34 VSUBS 0.006792f
C193 B.n35 VSUBS 0.006792f
C194 B.n36 VSUBS 0.006792f
C195 B.n37 VSUBS 0.006792f
C196 B.t11 VSUBS 0.190975f
C197 B.t10 VSUBS 0.211366f
C198 B.t9 VSUBS 0.762487f
C199 B.n38 VSUBS 0.32853f
C200 B.n39 VSUBS 0.231535f
C201 B.n40 VSUBS 0.015736f
C202 B.n41 VSUBS 0.006792f
C203 B.n42 VSUBS 0.006792f
C204 B.n43 VSUBS 0.006792f
C205 B.n44 VSUBS 0.006792f
C206 B.n45 VSUBS 0.006792f
C207 B.n46 VSUBS 0.006792f
C208 B.n47 VSUBS 0.006792f
C209 B.n48 VSUBS 0.006792f
C210 B.n49 VSUBS 0.006792f
C211 B.n50 VSUBS 0.006792f
C212 B.n51 VSUBS 0.006792f
C213 B.n52 VSUBS 0.006792f
C214 B.n53 VSUBS 0.006792f
C215 B.n54 VSUBS 0.006792f
C216 B.n55 VSUBS 0.006792f
C217 B.n56 VSUBS 0.006792f
C218 B.n57 VSUBS 0.006792f
C219 B.n58 VSUBS 0.006792f
C220 B.n59 VSUBS 0.006792f
C221 B.n60 VSUBS 0.016656f
C222 B.n61 VSUBS 0.006792f
C223 B.n62 VSUBS 0.006792f
C224 B.n63 VSUBS 0.006792f
C225 B.n64 VSUBS 0.006792f
C226 B.n65 VSUBS 0.006792f
C227 B.n66 VSUBS 0.006792f
C228 B.n67 VSUBS 0.006792f
C229 B.n68 VSUBS 0.006792f
C230 B.n69 VSUBS 0.006792f
C231 B.n70 VSUBS 0.006792f
C232 B.n71 VSUBS 0.006792f
C233 B.n72 VSUBS 0.006792f
C234 B.n73 VSUBS 0.006792f
C235 B.n74 VSUBS 0.006792f
C236 B.n75 VSUBS 0.006792f
C237 B.n76 VSUBS 0.006792f
C238 B.n77 VSUBS 0.006792f
C239 B.n78 VSUBS 0.006792f
C240 B.n79 VSUBS 0.006792f
C241 B.n80 VSUBS 0.01739f
C242 B.n81 VSUBS 0.006792f
C243 B.n82 VSUBS 0.006792f
C244 B.n83 VSUBS 0.006792f
C245 B.n84 VSUBS 0.006792f
C246 B.n85 VSUBS 0.006792f
C247 B.n86 VSUBS 0.006792f
C248 B.n87 VSUBS 0.006792f
C249 B.n88 VSUBS 0.006792f
C250 B.n89 VSUBS 0.006792f
C251 B.n90 VSUBS 0.006792f
C252 B.n91 VSUBS 0.006792f
C253 B.n92 VSUBS 0.006792f
C254 B.n93 VSUBS 0.006792f
C255 B.n94 VSUBS 0.006792f
C256 B.n95 VSUBS 0.006792f
C257 B.n96 VSUBS 0.006792f
C258 B.n97 VSUBS 0.006792f
C259 B.n98 VSUBS 0.006792f
C260 B.n99 VSUBS 0.006792f
C261 B.t4 VSUBS 0.190975f
C262 B.t5 VSUBS 0.211366f
C263 B.t3 VSUBS 0.762487f
C264 B.n100 VSUBS 0.32853f
C265 B.n101 VSUBS 0.231535f
C266 B.n102 VSUBS 0.015736f
C267 B.n103 VSUBS 0.006792f
C268 B.n104 VSUBS 0.006792f
C269 B.n105 VSUBS 0.006792f
C270 B.n106 VSUBS 0.006792f
C271 B.n107 VSUBS 0.006792f
C272 B.t7 VSUBS 0.190972f
C273 B.t8 VSUBS 0.211363f
C274 B.t6 VSUBS 0.762487f
C275 B.n108 VSUBS 0.328533f
C276 B.n109 VSUBS 0.231538f
C277 B.n110 VSUBS 0.006792f
C278 B.n111 VSUBS 0.006792f
C279 B.n112 VSUBS 0.006792f
C280 B.n113 VSUBS 0.006792f
C281 B.n114 VSUBS 0.006792f
C282 B.n115 VSUBS 0.006792f
C283 B.n116 VSUBS 0.006792f
C284 B.n117 VSUBS 0.006792f
C285 B.n118 VSUBS 0.006792f
C286 B.n119 VSUBS 0.006792f
C287 B.n120 VSUBS 0.006792f
C288 B.n121 VSUBS 0.006792f
C289 B.n122 VSUBS 0.006792f
C290 B.n123 VSUBS 0.006792f
C291 B.n124 VSUBS 0.006792f
C292 B.n125 VSUBS 0.006792f
C293 B.n126 VSUBS 0.006792f
C294 B.n127 VSUBS 0.006792f
C295 B.n128 VSUBS 0.006792f
C296 B.n129 VSUBS 0.01637f
C297 B.n130 VSUBS 0.006792f
C298 B.n131 VSUBS 0.006792f
C299 B.n132 VSUBS 0.006792f
C300 B.n133 VSUBS 0.006792f
C301 B.n134 VSUBS 0.006792f
C302 B.n135 VSUBS 0.006792f
C303 B.n136 VSUBS 0.006792f
C304 B.n137 VSUBS 0.006792f
C305 B.n138 VSUBS 0.006792f
C306 B.n139 VSUBS 0.006792f
C307 B.n140 VSUBS 0.006792f
C308 B.n141 VSUBS 0.006792f
C309 B.n142 VSUBS 0.006792f
C310 B.n143 VSUBS 0.006792f
C311 B.n144 VSUBS 0.006792f
C312 B.n145 VSUBS 0.006792f
C313 B.n146 VSUBS 0.006792f
C314 B.n147 VSUBS 0.006792f
C315 B.n148 VSUBS 0.006792f
C316 B.n149 VSUBS 0.006792f
C317 B.n150 VSUBS 0.006792f
C318 B.n151 VSUBS 0.006792f
C319 B.n152 VSUBS 0.006792f
C320 B.n153 VSUBS 0.006792f
C321 B.n154 VSUBS 0.006792f
C322 B.n155 VSUBS 0.006792f
C323 B.n156 VSUBS 0.006792f
C324 B.n157 VSUBS 0.006792f
C325 B.n158 VSUBS 0.006792f
C326 B.n159 VSUBS 0.006792f
C327 B.n160 VSUBS 0.006792f
C328 B.n161 VSUBS 0.006792f
C329 B.n162 VSUBS 0.006792f
C330 B.n163 VSUBS 0.006792f
C331 B.n164 VSUBS 0.01637f
C332 B.n165 VSUBS 0.01739f
C333 B.n166 VSUBS 0.01739f
C334 B.n167 VSUBS 0.006792f
C335 B.n168 VSUBS 0.006792f
C336 B.n169 VSUBS 0.006792f
C337 B.n170 VSUBS 0.006792f
C338 B.n171 VSUBS 0.006792f
C339 B.n172 VSUBS 0.006792f
C340 B.n173 VSUBS 0.006792f
C341 B.n174 VSUBS 0.006792f
C342 B.n175 VSUBS 0.006792f
C343 B.n176 VSUBS 0.006792f
C344 B.n177 VSUBS 0.006792f
C345 B.n178 VSUBS 0.006792f
C346 B.n179 VSUBS 0.006792f
C347 B.n180 VSUBS 0.006792f
C348 B.n181 VSUBS 0.006792f
C349 B.n182 VSUBS 0.006792f
C350 B.n183 VSUBS 0.006792f
C351 B.n184 VSUBS 0.006792f
C352 B.n185 VSUBS 0.006792f
C353 B.n186 VSUBS 0.006792f
C354 B.n187 VSUBS 0.006792f
C355 B.n188 VSUBS 0.006792f
C356 B.n189 VSUBS 0.006792f
C357 B.n190 VSUBS 0.006792f
C358 B.n191 VSUBS 0.006792f
C359 B.n192 VSUBS 0.006792f
C360 B.n193 VSUBS 0.006792f
C361 B.n194 VSUBS 0.006792f
C362 B.n195 VSUBS 0.006792f
C363 B.n196 VSUBS 0.006792f
C364 B.n197 VSUBS 0.006792f
C365 B.n198 VSUBS 0.006792f
C366 B.n199 VSUBS 0.006792f
C367 B.n200 VSUBS 0.006792f
C368 B.n201 VSUBS 0.006792f
C369 B.n202 VSUBS 0.006792f
C370 B.n203 VSUBS 0.006792f
C371 B.n204 VSUBS 0.006792f
C372 B.n205 VSUBS 0.006792f
C373 B.n206 VSUBS 0.006792f
C374 B.n207 VSUBS 0.006792f
C375 B.n208 VSUBS 0.006792f
C376 B.n209 VSUBS 0.006792f
C377 B.n210 VSUBS 0.006792f
C378 B.n211 VSUBS 0.006792f
C379 B.n212 VSUBS 0.006792f
C380 B.n213 VSUBS 0.006792f
C381 B.n214 VSUBS 0.006792f
C382 B.n215 VSUBS 0.006792f
C383 B.n216 VSUBS 0.006792f
C384 B.n217 VSUBS 0.006792f
C385 B.n218 VSUBS 0.006792f
C386 B.n219 VSUBS 0.006792f
C387 B.n220 VSUBS 0.006792f
C388 B.n221 VSUBS 0.006792f
C389 B.n222 VSUBS 0.006792f
C390 B.n223 VSUBS 0.006792f
C391 B.n224 VSUBS 0.004694f
C392 B.n225 VSUBS 0.015736f
C393 B.n226 VSUBS 0.005493f
C394 B.n227 VSUBS 0.006792f
C395 B.n228 VSUBS 0.006792f
C396 B.n229 VSUBS 0.006792f
C397 B.n230 VSUBS 0.006792f
C398 B.n231 VSUBS 0.006792f
C399 B.n232 VSUBS 0.006792f
C400 B.n233 VSUBS 0.006792f
C401 B.n234 VSUBS 0.006792f
C402 B.n235 VSUBS 0.006792f
C403 B.n236 VSUBS 0.006792f
C404 B.n237 VSUBS 0.006792f
C405 B.n238 VSUBS 0.005493f
C406 B.n239 VSUBS 0.006792f
C407 B.n240 VSUBS 0.006792f
C408 B.n241 VSUBS 0.004694f
C409 B.n242 VSUBS 0.006792f
C410 B.n243 VSUBS 0.006792f
C411 B.n244 VSUBS 0.006792f
C412 B.n245 VSUBS 0.006792f
C413 B.n246 VSUBS 0.006792f
C414 B.n247 VSUBS 0.006792f
C415 B.n248 VSUBS 0.006792f
C416 B.n249 VSUBS 0.006792f
C417 B.n250 VSUBS 0.006792f
C418 B.n251 VSUBS 0.006792f
C419 B.n252 VSUBS 0.006792f
C420 B.n253 VSUBS 0.006792f
C421 B.n254 VSUBS 0.006792f
C422 B.n255 VSUBS 0.006792f
C423 B.n256 VSUBS 0.006792f
C424 B.n257 VSUBS 0.006792f
C425 B.n258 VSUBS 0.006792f
C426 B.n259 VSUBS 0.006792f
C427 B.n260 VSUBS 0.006792f
C428 B.n261 VSUBS 0.006792f
C429 B.n262 VSUBS 0.006792f
C430 B.n263 VSUBS 0.006792f
C431 B.n264 VSUBS 0.006792f
C432 B.n265 VSUBS 0.006792f
C433 B.n266 VSUBS 0.006792f
C434 B.n267 VSUBS 0.006792f
C435 B.n268 VSUBS 0.006792f
C436 B.n269 VSUBS 0.006792f
C437 B.n270 VSUBS 0.006792f
C438 B.n271 VSUBS 0.006792f
C439 B.n272 VSUBS 0.006792f
C440 B.n273 VSUBS 0.006792f
C441 B.n274 VSUBS 0.006792f
C442 B.n275 VSUBS 0.006792f
C443 B.n276 VSUBS 0.006792f
C444 B.n277 VSUBS 0.006792f
C445 B.n278 VSUBS 0.006792f
C446 B.n279 VSUBS 0.006792f
C447 B.n280 VSUBS 0.006792f
C448 B.n281 VSUBS 0.006792f
C449 B.n282 VSUBS 0.006792f
C450 B.n283 VSUBS 0.006792f
C451 B.n284 VSUBS 0.006792f
C452 B.n285 VSUBS 0.006792f
C453 B.n286 VSUBS 0.006792f
C454 B.n287 VSUBS 0.006792f
C455 B.n288 VSUBS 0.006792f
C456 B.n289 VSUBS 0.006792f
C457 B.n290 VSUBS 0.006792f
C458 B.n291 VSUBS 0.006792f
C459 B.n292 VSUBS 0.006792f
C460 B.n293 VSUBS 0.006792f
C461 B.n294 VSUBS 0.006792f
C462 B.n295 VSUBS 0.006792f
C463 B.n296 VSUBS 0.006792f
C464 B.n297 VSUBS 0.006792f
C465 B.n298 VSUBS 0.006792f
C466 B.n299 VSUBS 0.01739f
C467 B.n300 VSUBS 0.01637f
C468 B.n301 VSUBS 0.01637f
C469 B.n302 VSUBS 0.006792f
C470 B.n303 VSUBS 0.006792f
C471 B.n304 VSUBS 0.006792f
C472 B.n305 VSUBS 0.006792f
C473 B.n306 VSUBS 0.006792f
C474 B.n307 VSUBS 0.006792f
C475 B.n308 VSUBS 0.006792f
C476 B.n309 VSUBS 0.006792f
C477 B.n310 VSUBS 0.006792f
C478 B.n311 VSUBS 0.006792f
C479 B.n312 VSUBS 0.006792f
C480 B.n313 VSUBS 0.006792f
C481 B.n314 VSUBS 0.006792f
C482 B.n315 VSUBS 0.006792f
C483 B.n316 VSUBS 0.006792f
C484 B.n317 VSUBS 0.006792f
C485 B.n318 VSUBS 0.006792f
C486 B.n319 VSUBS 0.006792f
C487 B.n320 VSUBS 0.006792f
C488 B.n321 VSUBS 0.006792f
C489 B.n322 VSUBS 0.006792f
C490 B.n323 VSUBS 0.006792f
C491 B.n324 VSUBS 0.006792f
C492 B.n325 VSUBS 0.006792f
C493 B.n326 VSUBS 0.006792f
C494 B.n327 VSUBS 0.006792f
C495 B.n328 VSUBS 0.006792f
C496 B.n329 VSUBS 0.006792f
C497 B.n330 VSUBS 0.006792f
C498 B.n331 VSUBS 0.006792f
C499 B.n332 VSUBS 0.006792f
C500 B.n333 VSUBS 0.006792f
C501 B.n334 VSUBS 0.006792f
C502 B.n335 VSUBS 0.006792f
C503 B.n336 VSUBS 0.006792f
C504 B.n337 VSUBS 0.006792f
C505 B.n338 VSUBS 0.006792f
C506 B.n339 VSUBS 0.006792f
C507 B.n340 VSUBS 0.006792f
C508 B.n341 VSUBS 0.006792f
C509 B.n342 VSUBS 0.006792f
C510 B.n343 VSUBS 0.006792f
C511 B.n344 VSUBS 0.006792f
C512 B.n345 VSUBS 0.006792f
C513 B.n346 VSUBS 0.006792f
C514 B.n347 VSUBS 0.006792f
C515 B.n348 VSUBS 0.006792f
C516 B.n349 VSUBS 0.006792f
C517 B.n350 VSUBS 0.006792f
C518 B.n351 VSUBS 0.006792f
C519 B.n352 VSUBS 0.006792f
C520 B.n353 VSUBS 0.006792f
C521 B.n354 VSUBS 0.006792f
C522 B.n355 VSUBS 0.006792f
C523 B.n356 VSUBS 0.006792f
C524 B.n357 VSUBS 0.017104f
C525 B.n358 VSUBS 0.01637f
C526 B.n359 VSUBS 0.01739f
C527 B.n360 VSUBS 0.006792f
C528 B.n361 VSUBS 0.006792f
C529 B.n362 VSUBS 0.006792f
C530 B.n363 VSUBS 0.006792f
C531 B.n364 VSUBS 0.006792f
C532 B.n365 VSUBS 0.006792f
C533 B.n366 VSUBS 0.006792f
C534 B.n367 VSUBS 0.006792f
C535 B.n368 VSUBS 0.006792f
C536 B.n369 VSUBS 0.006792f
C537 B.n370 VSUBS 0.006792f
C538 B.n371 VSUBS 0.006792f
C539 B.n372 VSUBS 0.006792f
C540 B.n373 VSUBS 0.006792f
C541 B.n374 VSUBS 0.006792f
C542 B.n375 VSUBS 0.006792f
C543 B.n376 VSUBS 0.006792f
C544 B.n377 VSUBS 0.006792f
C545 B.n378 VSUBS 0.006792f
C546 B.n379 VSUBS 0.006792f
C547 B.n380 VSUBS 0.006792f
C548 B.n381 VSUBS 0.006792f
C549 B.n382 VSUBS 0.006792f
C550 B.n383 VSUBS 0.006792f
C551 B.n384 VSUBS 0.006792f
C552 B.n385 VSUBS 0.006792f
C553 B.n386 VSUBS 0.006792f
C554 B.n387 VSUBS 0.006792f
C555 B.n388 VSUBS 0.006792f
C556 B.n389 VSUBS 0.006792f
C557 B.n390 VSUBS 0.006792f
C558 B.n391 VSUBS 0.006792f
C559 B.n392 VSUBS 0.006792f
C560 B.n393 VSUBS 0.006792f
C561 B.n394 VSUBS 0.006792f
C562 B.n395 VSUBS 0.006792f
C563 B.n396 VSUBS 0.006792f
C564 B.n397 VSUBS 0.006792f
C565 B.n398 VSUBS 0.006792f
C566 B.n399 VSUBS 0.006792f
C567 B.n400 VSUBS 0.006792f
C568 B.n401 VSUBS 0.006792f
C569 B.n402 VSUBS 0.006792f
C570 B.n403 VSUBS 0.006792f
C571 B.n404 VSUBS 0.006792f
C572 B.n405 VSUBS 0.006792f
C573 B.n406 VSUBS 0.006792f
C574 B.n407 VSUBS 0.006792f
C575 B.n408 VSUBS 0.006792f
C576 B.n409 VSUBS 0.006792f
C577 B.n410 VSUBS 0.006792f
C578 B.n411 VSUBS 0.006792f
C579 B.n412 VSUBS 0.006792f
C580 B.n413 VSUBS 0.006792f
C581 B.n414 VSUBS 0.006792f
C582 B.n415 VSUBS 0.006792f
C583 B.n416 VSUBS 0.006792f
C584 B.n417 VSUBS 0.004694f
C585 B.n418 VSUBS 0.006792f
C586 B.n419 VSUBS 0.006792f
C587 B.n420 VSUBS 0.005493f
C588 B.n421 VSUBS 0.006792f
C589 B.n422 VSUBS 0.006792f
C590 B.n423 VSUBS 0.006792f
C591 B.n424 VSUBS 0.006792f
C592 B.n425 VSUBS 0.006792f
C593 B.n426 VSUBS 0.006792f
C594 B.n427 VSUBS 0.006792f
C595 B.n428 VSUBS 0.006792f
C596 B.n429 VSUBS 0.006792f
C597 B.n430 VSUBS 0.006792f
C598 B.n431 VSUBS 0.006792f
C599 B.n432 VSUBS 0.005493f
C600 B.n433 VSUBS 0.015736f
C601 B.n434 VSUBS 0.004694f
C602 B.n435 VSUBS 0.006792f
C603 B.n436 VSUBS 0.006792f
C604 B.n437 VSUBS 0.006792f
C605 B.n438 VSUBS 0.006792f
C606 B.n439 VSUBS 0.006792f
C607 B.n440 VSUBS 0.006792f
C608 B.n441 VSUBS 0.006792f
C609 B.n442 VSUBS 0.006792f
C610 B.n443 VSUBS 0.006792f
C611 B.n444 VSUBS 0.006792f
C612 B.n445 VSUBS 0.006792f
C613 B.n446 VSUBS 0.006792f
C614 B.n447 VSUBS 0.006792f
C615 B.n448 VSUBS 0.006792f
C616 B.n449 VSUBS 0.006792f
C617 B.n450 VSUBS 0.006792f
C618 B.n451 VSUBS 0.006792f
C619 B.n452 VSUBS 0.006792f
C620 B.n453 VSUBS 0.006792f
C621 B.n454 VSUBS 0.006792f
C622 B.n455 VSUBS 0.006792f
C623 B.n456 VSUBS 0.006792f
C624 B.n457 VSUBS 0.006792f
C625 B.n458 VSUBS 0.006792f
C626 B.n459 VSUBS 0.006792f
C627 B.n460 VSUBS 0.006792f
C628 B.n461 VSUBS 0.006792f
C629 B.n462 VSUBS 0.006792f
C630 B.n463 VSUBS 0.006792f
C631 B.n464 VSUBS 0.006792f
C632 B.n465 VSUBS 0.006792f
C633 B.n466 VSUBS 0.006792f
C634 B.n467 VSUBS 0.006792f
C635 B.n468 VSUBS 0.006792f
C636 B.n469 VSUBS 0.006792f
C637 B.n470 VSUBS 0.006792f
C638 B.n471 VSUBS 0.006792f
C639 B.n472 VSUBS 0.006792f
C640 B.n473 VSUBS 0.006792f
C641 B.n474 VSUBS 0.006792f
C642 B.n475 VSUBS 0.006792f
C643 B.n476 VSUBS 0.006792f
C644 B.n477 VSUBS 0.006792f
C645 B.n478 VSUBS 0.006792f
C646 B.n479 VSUBS 0.006792f
C647 B.n480 VSUBS 0.006792f
C648 B.n481 VSUBS 0.006792f
C649 B.n482 VSUBS 0.006792f
C650 B.n483 VSUBS 0.006792f
C651 B.n484 VSUBS 0.006792f
C652 B.n485 VSUBS 0.006792f
C653 B.n486 VSUBS 0.006792f
C654 B.n487 VSUBS 0.006792f
C655 B.n488 VSUBS 0.006792f
C656 B.n489 VSUBS 0.006792f
C657 B.n490 VSUBS 0.006792f
C658 B.n491 VSUBS 0.006792f
C659 B.n492 VSUBS 0.01739f
C660 B.n493 VSUBS 0.01739f
C661 B.n494 VSUBS 0.01637f
C662 B.n495 VSUBS 0.006792f
C663 B.n496 VSUBS 0.006792f
C664 B.n497 VSUBS 0.006792f
C665 B.n498 VSUBS 0.006792f
C666 B.n499 VSUBS 0.006792f
C667 B.n500 VSUBS 0.006792f
C668 B.n501 VSUBS 0.006792f
C669 B.n502 VSUBS 0.006792f
C670 B.n503 VSUBS 0.006792f
C671 B.n504 VSUBS 0.006792f
C672 B.n505 VSUBS 0.006792f
C673 B.n506 VSUBS 0.006792f
C674 B.n507 VSUBS 0.006792f
C675 B.n508 VSUBS 0.006792f
C676 B.n509 VSUBS 0.006792f
C677 B.n510 VSUBS 0.006792f
C678 B.n511 VSUBS 0.006792f
C679 B.n512 VSUBS 0.006792f
C680 B.n513 VSUBS 0.006792f
C681 B.n514 VSUBS 0.006792f
C682 B.n515 VSUBS 0.006792f
C683 B.n516 VSUBS 0.006792f
C684 B.n517 VSUBS 0.006792f
C685 B.n518 VSUBS 0.006792f
C686 B.n519 VSUBS 0.006792f
C687 B.n520 VSUBS 0.006792f
C688 B.n521 VSUBS 0.006792f
C689 B.n522 VSUBS 0.006792f
C690 B.n523 VSUBS 0.015379f
C691 VDD2.n0 VSUBS 0.021448f
C692 VDD2.n1 VSUBS 0.020221f
C693 VDD2.n2 VSUBS 0.010866f
C694 VDD2.n3 VSUBS 0.025682f
C695 VDD2.n4 VSUBS 0.011505f
C696 VDD2.n5 VSUBS 0.020221f
C697 VDD2.n6 VSUBS 0.010866f
C698 VDD2.n7 VSUBS 0.025682f
C699 VDD2.n8 VSUBS 0.011185f
C700 VDD2.n9 VSUBS 0.020221f
C701 VDD2.n10 VSUBS 0.011505f
C702 VDD2.n11 VSUBS 0.025682f
C703 VDD2.n12 VSUBS 0.011505f
C704 VDD2.n13 VSUBS 0.020221f
C705 VDD2.n14 VSUBS 0.010866f
C706 VDD2.n15 VSUBS 0.025682f
C707 VDD2.n16 VSUBS 0.011505f
C708 VDD2.n17 VSUBS 0.936792f
C709 VDD2.n18 VSUBS 0.010866f
C710 VDD2.t1 VSUBS 0.055301f
C711 VDD2.n19 VSUBS 0.153399f
C712 VDD2.n20 VSUBS 0.01932f
C713 VDD2.n21 VSUBS 0.019262f
C714 VDD2.n22 VSUBS 0.025682f
C715 VDD2.n23 VSUBS 0.011505f
C716 VDD2.n24 VSUBS 0.010866f
C717 VDD2.n25 VSUBS 0.020221f
C718 VDD2.n26 VSUBS 0.020221f
C719 VDD2.n27 VSUBS 0.010866f
C720 VDD2.n28 VSUBS 0.011505f
C721 VDD2.n29 VSUBS 0.025682f
C722 VDD2.n30 VSUBS 0.025682f
C723 VDD2.n31 VSUBS 0.011505f
C724 VDD2.n32 VSUBS 0.010866f
C725 VDD2.n33 VSUBS 0.020221f
C726 VDD2.n34 VSUBS 0.020221f
C727 VDD2.n35 VSUBS 0.010866f
C728 VDD2.n36 VSUBS 0.010866f
C729 VDD2.n37 VSUBS 0.011505f
C730 VDD2.n38 VSUBS 0.025682f
C731 VDD2.n39 VSUBS 0.025682f
C732 VDD2.n40 VSUBS 0.025682f
C733 VDD2.n41 VSUBS 0.011185f
C734 VDD2.n42 VSUBS 0.010866f
C735 VDD2.n43 VSUBS 0.020221f
C736 VDD2.n44 VSUBS 0.020221f
C737 VDD2.n45 VSUBS 0.010866f
C738 VDD2.n46 VSUBS 0.011505f
C739 VDD2.n47 VSUBS 0.025682f
C740 VDD2.n48 VSUBS 0.025682f
C741 VDD2.n49 VSUBS 0.011505f
C742 VDD2.n50 VSUBS 0.010866f
C743 VDD2.n51 VSUBS 0.020221f
C744 VDD2.n52 VSUBS 0.020221f
C745 VDD2.n53 VSUBS 0.010866f
C746 VDD2.n54 VSUBS 0.011505f
C747 VDD2.n55 VSUBS 0.025682f
C748 VDD2.n56 VSUBS 0.059551f
C749 VDD2.n57 VSUBS 0.011505f
C750 VDD2.n58 VSUBS 0.010866f
C751 VDD2.n59 VSUBS 0.045634f
C752 VDD2.n60 VSUBS 0.52578f
C753 VDD2.n61 VSUBS 0.021448f
C754 VDD2.n62 VSUBS 0.020221f
C755 VDD2.n63 VSUBS 0.010866f
C756 VDD2.n64 VSUBS 0.025682f
C757 VDD2.n65 VSUBS 0.011505f
C758 VDD2.n66 VSUBS 0.020221f
C759 VDD2.n67 VSUBS 0.010866f
C760 VDD2.n68 VSUBS 0.025682f
C761 VDD2.n69 VSUBS 0.011185f
C762 VDD2.n70 VSUBS 0.020221f
C763 VDD2.n71 VSUBS 0.011185f
C764 VDD2.n72 VSUBS 0.010866f
C765 VDD2.n73 VSUBS 0.025682f
C766 VDD2.n74 VSUBS 0.025682f
C767 VDD2.n75 VSUBS 0.011505f
C768 VDD2.n76 VSUBS 0.020221f
C769 VDD2.n77 VSUBS 0.010866f
C770 VDD2.n78 VSUBS 0.025682f
C771 VDD2.n79 VSUBS 0.011505f
C772 VDD2.n80 VSUBS 0.936792f
C773 VDD2.n81 VSUBS 0.010866f
C774 VDD2.t0 VSUBS 0.055301f
C775 VDD2.n82 VSUBS 0.153399f
C776 VDD2.n83 VSUBS 0.01932f
C777 VDD2.n84 VSUBS 0.019262f
C778 VDD2.n85 VSUBS 0.025682f
C779 VDD2.n86 VSUBS 0.011505f
C780 VDD2.n87 VSUBS 0.010866f
C781 VDD2.n88 VSUBS 0.020221f
C782 VDD2.n89 VSUBS 0.020221f
C783 VDD2.n90 VSUBS 0.010866f
C784 VDD2.n91 VSUBS 0.011505f
C785 VDD2.n92 VSUBS 0.025682f
C786 VDD2.n93 VSUBS 0.025682f
C787 VDD2.n94 VSUBS 0.011505f
C788 VDD2.n95 VSUBS 0.010866f
C789 VDD2.n96 VSUBS 0.020221f
C790 VDD2.n97 VSUBS 0.020221f
C791 VDD2.n98 VSUBS 0.010866f
C792 VDD2.n99 VSUBS 0.011505f
C793 VDD2.n100 VSUBS 0.025682f
C794 VDD2.n101 VSUBS 0.025682f
C795 VDD2.n102 VSUBS 0.011505f
C796 VDD2.n103 VSUBS 0.010866f
C797 VDD2.n104 VSUBS 0.020221f
C798 VDD2.n105 VSUBS 0.020221f
C799 VDD2.n106 VSUBS 0.010866f
C800 VDD2.n107 VSUBS 0.011505f
C801 VDD2.n108 VSUBS 0.025682f
C802 VDD2.n109 VSUBS 0.025682f
C803 VDD2.n110 VSUBS 0.011505f
C804 VDD2.n111 VSUBS 0.010866f
C805 VDD2.n112 VSUBS 0.020221f
C806 VDD2.n113 VSUBS 0.020221f
C807 VDD2.n114 VSUBS 0.010866f
C808 VDD2.n115 VSUBS 0.011505f
C809 VDD2.n116 VSUBS 0.025682f
C810 VDD2.n117 VSUBS 0.059551f
C811 VDD2.n118 VSUBS 0.011505f
C812 VDD2.n119 VSUBS 0.010866f
C813 VDD2.n120 VSUBS 0.045634f
C814 VDD2.n121 VSUBS 0.043768f
C815 VDD2.n122 VSUBS 2.24652f
C816 VTAIL.n0 VSUBS 0.030883f
C817 VTAIL.n1 VSUBS 0.029116f
C818 VTAIL.n2 VSUBS 0.015646f
C819 VTAIL.n3 VSUBS 0.03698f
C820 VTAIL.n4 VSUBS 0.016566f
C821 VTAIL.n5 VSUBS 0.029116f
C822 VTAIL.n6 VSUBS 0.015646f
C823 VTAIL.n7 VSUBS 0.03698f
C824 VTAIL.n8 VSUBS 0.016106f
C825 VTAIL.n9 VSUBS 0.029116f
C826 VTAIL.n10 VSUBS 0.016566f
C827 VTAIL.n11 VSUBS 0.03698f
C828 VTAIL.n12 VSUBS 0.016566f
C829 VTAIL.n13 VSUBS 0.029116f
C830 VTAIL.n14 VSUBS 0.015646f
C831 VTAIL.n15 VSUBS 0.03698f
C832 VTAIL.n16 VSUBS 0.016566f
C833 VTAIL.n17 VSUBS 1.34889f
C834 VTAIL.n18 VSUBS 0.015646f
C835 VTAIL.t0 VSUBS 0.079628f
C836 VTAIL.n19 VSUBS 0.220879f
C837 VTAIL.n20 VSUBS 0.027819f
C838 VTAIL.n21 VSUBS 0.027735f
C839 VTAIL.n22 VSUBS 0.03698f
C840 VTAIL.n23 VSUBS 0.016566f
C841 VTAIL.n24 VSUBS 0.015646f
C842 VTAIL.n25 VSUBS 0.029116f
C843 VTAIL.n26 VSUBS 0.029116f
C844 VTAIL.n27 VSUBS 0.015646f
C845 VTAIL.n28 VSUBS 0.016566f
C846 VTAIL.n29 VSUBS 0.03698f
C847 VTAIL.n30 VSUBS 0.03698f
C848 VTAIL.n31 VSUBS 0.016566f
C849 VTAIL.n32 VSUBS 0.015646f
C850 VTAIL.n33 VSUBS 0.029116f
C851 VTAIL.n34 VSUBS 0.029116f
C852 VTAIL.n35 VSUBS 0.015646f
C853 VTAIL.n36 VSUBS 0.015646f
C854 VTAIL.n37 VSUBS 0.016566f
C855 VTAIL.n38 VSUBS 0.03698f
C856 VTAIL.n39 VSUBS 0.03698f
C857 VTAIL.n40 VSUBS 0.03698f
C858 VTAIL.n41 VSUBS 0.016106f
C859 VTAIL.n42 VSUBS 0.015646f
C860 VTAIL.n43 VSUBS 0.029116f
C861 VTAIL.n44 VSUBS 0.029116f
C862 VTAIL.n45 VSUBS 0.015646f
C863 VTAIL.n46 VSUBS 0.016566f
C864 VTAIL.n47 VSUBS 0.03698f
C865 VTAIL.n48 VSUBS 0.03698f
C866 VTAIL.n49 VSUBS 0.016566f
C867 VTAIL.n50 VSUBS 0.015646f
C868 VTAIL.n51 VSUBS 0.029116f
C869 VTAIL.n52 VSUBS 0.029116f
C870 VTAIL.n53 VSUBS 0.015646f
C871 VTAIL.n54 VSUBS 0.016566f
C872 VTAIL.n55 VSUBS 0.03698f
C873 VTAIL.n56 VSUBS 0.085747f
C874 VTAIL.n57 VSUBS 0.016566f
C875 VTAIL.n58 VSUBS 0.015646f
C876 VTAIL.n59 VSUBS 0.065708f
C877 VTAIL.n60 VSUBS 0.042904f
C878 VTAIL.n61 VSUBS 1.73352f
C879 VTAIL.n62 VSUBS 0.030883f
C880 VTAIL.n63 VSUBS 0.029116f
C881 VTAIL.n64 VSUBS 0.015646f
C882 VTAIL.n65 VSUBS 0.03698f
C883 VTAIL.n66 VSUBS 0.016566f
C884 VTAIL.n67 VSUBS 0.029116f
C885 VTAIL.n68 VSUBS 0.015646f
C886 VTAIL.n69 VSUBS 0.03698f
C887 VTAIL.n70 VSUBS 0.016106f
C888 VTAIL.n71 VSUBS 0.029116f
C889 VTAIL.n72 VSUBS 0.016106f
C890 VTAIL.n73 VSUBS 0.015646f
C891 VTAIL.n74 VSUBS 0.03698f
C892 VTAIL.n75 VSUBS 0.03698f
C893 VTAIL.n76 VSUBS 0.016566f
C894 VTAIL.n77 VSUBS 0.029116f
C895 VTAIL.n78 VSUBS 0.015646f
C896 VTAIL.n79 VSUBS 0.03698f
C897 VTAIL.n80 VSUBS 0.016566f
C898 VTAIL.n81 VSUBS 1.34889f
C899 VTAIL.n82 VSUBS 0.015646f
C900 VTAIL.t3 VSUBS 0.079628f
C901 VTAIL.n83 VSUBS 0.220879f
C902 VTAIL.n84 VSUBS 0.027819f
C903 VTAIL.n85 VSUBS 0.027735f
C904 VTAIL.n86 VSUBS 0.03698f
C905 VTAIL.n87 VSUBS 0.016566f
C906 VTAIL.n88 VSUBS 0.015646f
C907 VTAIL.n89 VSUBS 0.029116f
C908 VTAIL.n90 VSUBS 0.029116f
C909 VTAIL.n91 VSUBS 0.015646f
C910 VTAIL.n92 VSUBS 0.016566f
C911 VTAIL.n93 VSUBS 0.03698f
C912 VTAIL.n94 VSUBS 0.03698f
C913 VTAIL.n95 VSUBS 0.016566f
C914 VTAIL.n96 VSUBS 0.015646f
C915 VTAIL.n97 VSUBS 0.029116f
C916 VTAIL.n98 VSUBS 0.029116f
C917 VTAIL.n99 VSUBS 0.015646f
C918 VTAIL.n100 VSUBS 0.016566f
C919 VTAIL.n101 VSUBS 0.03698f
C920 VTAIL.n102 VSUBS 0.03698f
C921 VTAIL.n103 VSUBS 0.016566f
C922 VTAIL.n104 VSUBS 0.015646f
C923 VTAIL.n105 VSUBS 0.029116f
C924 VTAIL.n106 VSUBS 0.029116f
C925 VTAIL.n107 VSUBS 0.015646f
C926 VTAIL.n108 VSUBS 0.016566f
C927 VTAIL.n109 VSUBS 0.03698f
C928 VTAIL.n110 VSUBS 0.03698f
C929 VTAIL.n111 VSUBS 0.016566f
C930 VTAIL.n112 VSUBS 0.015646f
C931 VTAIL.n113 VSUBS 0.029116f
C932 VTAIL.n114 VSUBS 0.029116f
C933 VTAIL.n115 VSUBS 0.015646f
C934 VTAIL.n116 VSUBS 0.016566f
C935 VTAIL.n117 VSUBS 0.03698f
C936 VTAIL.n118 VSUBS 0.085747f
C937 VTAIL.n119 VSUBS 0.016566f
C938 VTAIL.n120 VSUBS 0.015646f
C939 VTAIL.n121 VSUBS 0.065708f
C940 VTAIL.n122 VSUBS 0.042904f
C941 VTAIL.n123 VSUBS 1.76647f
C942 VTAIL.n124 VSUBS 0.030883f
C943 VTAIL.n125 VSUBS 0.029116f
C944 VTAIL.n126 VSUBS 0.015646f
C945 VTAIL.n127 VSUBS 0.03698f
C946 VTAIL.n128 VSUBS 0.016566f
C947 VTAIL.n129 VSUBS 0.029116f
C948 VTAIL.n130 VSUBS 0.015646f
C949 VTAIL.n131 VSUBS 0.03698f
C950 VTAIL.n132 VSUBS 0.016106f
C951 VTAIL.n133 VSUBS 0.029116f
C952 VTAIL.n134 VSUBS 0.016106f
C953 VTAIL.n135 VSUBS 0.015646f
C954 VTAIL.n136 VSUBS 0.03698f
C955 VTAIL.n137 VSUBS 0.03698f
C956 VTAIL.n138 VSUBS 0.016566f
C957 VTAIL.n139 VSUBS 0.029116f
C958 VTAIL.n140 VSUBS 0.015646f
C959 VTAIL.n141 VSUBS 0.03698f
C960 VTAIL.n142 VSUBS 0.016566f
C961 VTAIL.n143 VSUBS 1.34889f
C962 VTAIL.n144 VSUBS 0.015646f
C963 VTAIL.t1 VSUBS 0.079628f
C964 VTAIL.n145 VSUBS 0.220879f
C965 VTAIL.n146 VSUBS 0.027819f
C966 VTAIL.n147 VSUBS 0.027735f
C967 VTAIL.n148 VSUBS 0.03698f
C968 VTAIL.n149 VSUBS 0.016566f
C969 VTAIL.n150 VSUBS 0.015646f
C970 VTAIL.n151 VSUBS 0.029116f
C971 VTAIL.n152 VSUBS 0.029116f
C972 VTAIL.n153 VSUBS 0.015646f
C973 VTAIL.n154 VSUBS 0.016566f
C974 VTAIL.n155 VSUBS 0.03698f
C975 VTAIL.n156 VSUBS 0.03698f
C976 VTAIL.n157 VSUBS 0.016566f
C977 VTAIL.n158 VSUBS 0.015646f
C978 VTAIL.n159 VSUBS 0.029116f
C979 VTAIL.n160 VSUBS 0.029116f
C980 VTAIL.n161 VSUBS 0.015646f
C981 VTAIL.n162 VSUBS 0.016566f
C982 VTAIL.n163 VSUBS 0.03698f
C983 VTAIL.n164 VSUBS 0.03698f
C984 VTAIL.n165 VSUBS 0.016566f
C985 VTAIL.n166 VSUBS 0.015646f
C986 VTAIL.n167 VSUBS 0.029116f
C987 VTAIL.n168 VSUBS 0.029116f
C988 VTAIL.n169 VSUBS 0.015646f
C989 VTAIL.n170 VSUBS 0.016566f
C990 VTAIL.n171 VSUBS 0.03698f
C991 VTAIL.n172 VSUBS 0.03698f
C992 VTAIL.n173 VSUBS 0.016566f
C993 VTAIL.n174 VSUBS 0.015646f
C994 VTAIL.n175 VSUBS 0.029116f
C995 VTAIL.n176 VSUBS 0.029116f
C996 VTAIL.n177 VSUBS 0.015646f
C997 VTAIL.n178 VSUBS 0.016566f
C998 VTAIL.n179 VSUBS 0.03698f
C999 VTAIL.n180 VSUBS 0.085747f
C1000 VTAIL.n181 VSUBS 0.016566f
C1001 VTAIL.n182 VSUBS 0.015646f
C1002 VTAIL.n183 VSUBS 0.065708f
C1003 VTAIL.n184 VSUBS 0.042904f
C1004 VTAIL.n185 VSUBS 1.61281f
C1005 VTAIL.n186 VSUBS 0.030883f
C1006 VTAIL.n187 VSUBS 0.029116f
C1007 VTAIL.n188 VSUBS 0.015646f
C1008 VTAIL.n189 VSUBS 0.03698f
C1009 VTAIL.n190 VSUBS 0.016566f
C1010 VTAIL.n191 VSUBS 0.029116f
C1011 VTAIL.n192 VSUBS 0.015646f
C1012 VTAIL.n193 VSUBS 0.03698f
C1013 VTAIL.n194 VSUBS 0.016106f
C1014 VTAIL.n195 VSUBS 0.029116f
C1015 VTAIL.n196 VSUBS 0.016566f
C1016 VTAIL.n197 VSUBS 0.03698f
C1017 VTAIL.n198 VSUBS 0.016566f
C1018 VTAIL.n199 VSUBS 0.029116f
C1019 VTAIL.n200 VSUBS 0.015646f
C1020 VTAIL.n201 VSUBS 0.03698f
C1021 VTAIL.n202 VSUBS 0.016566f
C1022 VTAIL.n203 VSUBS 1.34889f
C1023 VTAIL.n204 VSUBS 0.015646f
C1024 VTAIL.t2 VSUBS 0.079628f
C1025 VTAIL.n205 VSUBS 0.220879f
C1026 VTAIL.n206 VSUBS 0.027819f
C1027 VTAIL.n207 VSUBS 0.027735f
C1028 VTAIL.n208 VSUBS 0.03698f
C1029 VTAIL.n209 VSUBS 0.016566f
C1030 VTAIL.n210 VSUBS 0.015646f
C1031 VTAIL.n211 VSUBS 0.029116f
C1032 VTAIL.n212 VSUBS 0.029116f
C1033 VTAIL.n213 VSUBS 0.015646f
C1034 VTAIL.n214 VSUBS 0.016566f
C1035 VTAIL.n215 VSUBS 0.03698f
C1036 VTAIL.n216 VSUBS 0.03698f
C1037 VTAIL.n217 VSUBS 0.016566f
C1038 VTAIL.n218 VSUBS 0.015646f
C1039 VTAIL.n219 VSUBS 0.029116f
C1040 VTAIL.n220 VSUBS 0.029116f
C1041 VTAIL.n221 VSUBS 0.015646f
C1042 VTAIL.n222 VSUBS 0.015646f
C1043 VTAIL.n223 VSUBS 0.016566f
C1044 VTAIL.n224 VSUBS 0.03698f
C1045 VTAIL.n225 VSUBS 0.03698f
C1046 VTAIL.n226 VSUBS 0.03698f
C1047 VTAIL.n227 VSUBS 0.016106f
C1048 VTAIL.n228 VSUBS 0.015646f
C1049 VTAIL.n229 VSUBS 0.029116f
C1050 VTAIL.n230 VSUBS 0.029116f
C1051 VTAIL.n231 VSUBS 0.015646f
C1052 VTAIL.n232 VSUBS 0.016566f
C1053 VTAIL.n233 VSUBS 0.03698f
C1054 VTAIL.n234 VSUBS 0.03698f
C1055 VTAIL.n235 VSUBS 0.016566f
C1056 VTAIL.n236 VSUBS 0.015646f
C1057 VTAIL.n237 VSUBS 0.029116f
C1058 VTAIL.n238 VSUBS 0.029116f
C1059 VTAIL.n239 VSUBS 0.015646f
C1060 VTAIL.n240 VSUBS 0.016566f
C1061 VTAIL.n241 VSUBS 0.03698f
C1062 VTAIL.n242 VSUBS 0.085747f
C1063 VTAIL.n243 VSUBS 0.016566f
C1064 VTAIL.n244 VSUBS 0.015646f
C1065 VTAIL.n245 VSUBS 0.065708f
C1066 VTAIL.n246 VSUBS 0.042904f
C1067 VTAIL.n247 VSUBS 1.52485f
C1068 VN.t0 VSUBS 2.87172f
C1069 VN.t1 VSUBS 3.24086f
.ends

