* NGSPICE file created from diff_pair_sample_0265.ext - technology: sky130A

.subckt diff_pair_sample_0265 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t17 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.8424 ps=5.1 w=2.16 l=2.89
X1 VTAIL.t14 VN.t1 VDD2.t8 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X2 VDD1.t9 VP.t0 VTAIL.t19 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.8424 ps=5.1 w=2.16 l=2.89
X3 VTAIL.t0 VP.t1 VDD1.t8 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X4 B.t11 B.t9 B.t10 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.8424 pd=5.1 as=0 ps=0 w=2.16 l=2.89
X5 VTAIL.t10 VN.t2 VDD2.t7 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X6 VDD2.t6 VN.t3 VTAIL.t11 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.8424 pd=5.1 as=0.3564 ps=2.49 w=2.16 l=2.89
X7 VDD1.t7 VP.t2 VTAIL.t1 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X8 VDD2.t5 VN.t4 VTAIL.t18 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.8424 ps=5.1 w=2.16 l=2.89
X9 VTAIL.t9 VN.t5 VDD2.t4 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X10 B.t8 B.t6 B.t7 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.8424 pd=5.1 as=0 ps=0 w=2.16 l=2.89
X11 VTAIL.t16 VN.t6 VDD2.t3 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X12 VTAIL.t3 VP.t3 VDD1.t6 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X13 VDD2.t2 VN.t7 VTAIL.t15 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X14 VTAIL.t5 VP.t4 VDD1.t5 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X15 VTAIL.t4 VP.t5 VDD1.t4 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X16 VDD1.t3 VP.t6 VTAIL.t8 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.8424 pd=5.1 as=0.3564 ps=2.49 w=2.16 l=2.89
X17 VDD1.t2 VP.t7 VTAIL.t6 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.8424 pd=5.1 as=0.3564 ps=2.49 w=2.16 l=2.89
X18 VDD2.t1 VN.t8 VTAIL.t13 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.8424 pd=5.1 as=0.3564 ps=2.49 w=2.16 l=2.89
X19 VDD2.t0 VN.t9 VTAIL.t12 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X20 VDD1.t1 VP.t8 VTAIL.t7 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.3564 ps=2.49 w=2.16 l=2.89
X21 VDD1.t0 VP.t9 VTAIL.t2 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.3564 pd=2.49 as=0.8424 ps=5.1 w=2.16 l=2.89
X22 B.t5 B.t3 B.t4 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.8424 pd=5.1 as=0 ps=0 w=2.16 l=2.89
X23 B.t2 B.t0 B.t1 w_n4834_n1400# sky130_fd_pr__pfet_01v8 ad=0.8424 pd=5.1 as=0 ps=0 w=2.16 l=2.89
R0 VN.n84 VN.n83 161.3
R1 VN.n82 VN.n44 161.3
R2 VN.n81 VN.n80 161.3
R3 VN.n79 VN.n45 161.3
R4 VN.n78 VN.n77 161.3
R5 VN.n76 VN.n46 161.3
R6 VN.n74 VN.n73 161.3
R7 VN.n72 VN.n47 161.3
R8 VN.n71 VN.n70 161.3
R9 VN.n69 VN.n48 161.3
R10 VN.n68 VN.n67 161.3
R11 VN.n66 VN.n49 161.3
R12 VN.n65 VN.n64 161.3
R13 VN.n63 VN.n50 161.3
R14 VN.n62 VN.n61 161.3
R15 VN.n60 VN.n51 161.3
R16 VN.n59 VN.n58 161.3
R17 VN.n57 VN.n52 161.3
R18 VN.n56 VN.n55 161.3
R19 VN.n41 VN.n40 161.3
R20 VN.n39 VN.n1 161.3
R21 VN.n38 VN.n37 161.3
R22 VN.n36 VN.n2 161.3
R23 VN.n35 VN.n34 161.3
R24 VN.n33 VN.n3 161.3
R25 VN.n31 VN.n30 161.3
R26 VN.n29 VN.n4 161.3
R27 VN.n28 VN.n27 161.3
R28 VN.n26 VN.n5 161.3
R29 VN.n25 VN.n24 161.3
R30 VN.n23 VN.n6 161.3
R31 VN.n22 VN.n21 161.3
R32 VN.n20 VN.n7 161.3
R33 VN.n19 VN.n18 161.3
R34 VN.n17 VN.n8 161.3
R35 VN.n16 VN.n15 161.3
R36 VN.n14 VN.n9 161.3
R37 VN.n13 VN.n12 161.3
R38 VN.n42 VN.n0 68.6047
R39 VN.n85 VN.n43 68.6047
R40 VN.n11 VN.n10 63.1738
R41 VN.n54 VN.n53 63.1738
R42 VN.n38 VN.n2 56.5617
R43 VN.n81 VN.n45 56.5617
R44 VN.n15 VN.n8 51.2335
R45 VN.n27 VN.n26 51.2335
R46 VN.n58 VN.n51 51.2335
R47 VN.n70 VN.n69 51.2335
R48 VN.n54 VN.t4 49.8399
R49 VN.n11 VN.t8 49.8399
R50 VN VN.n85 47.5209
R51 VN.n19 VN.n8 29.9206
R52 VN.n26 VN.n25 29.9206
R53 VN.n62 VN.n51 29.9206
R54 VN.n69 VN.n68 29.9206
R55 VN.n14 VN.n13 24.5923
R56 VN.n15 VN.n14 24.5923
R57 VN.n20 VN.n19 24.5923
R58 VN.n21 VN.n20 24.5923
R59 VN.n21 VN.n6 24.5923
R60 VN.n25 VN.n6 24.5923
R61 VN.n27 VN.n4 24.5923
R62 VN.n31 VN.n4 24.5923
R63 VN.n34 VN.n33 24.5923
R64 VN.n34 VN.n2 24.5923
R65 VN.n39 VN.n38 24.5923
R66 VN.n40 VN.n39 24.5923
R67 VN.n58 VN.n57 24.5923
R68 VN.n57 VN.n56 24.5923
R69 VN.n68 VN.n49 24.5923
R70 VN.n64 VN.n49 24.5923
R71 VN.n64 VN.n63 24.5923
R72 VN.n63 VN.n62 24.5923
R73 VN.n77 VN.n45 24.5923
R74 VN.n77 VN.n76 24.5923
R75 VN.n74 VN.n47 24.5923
R76 VN.n70 VN.n47 24.5923
R77 VN.n83 VN.n82 24.5923
R78 VN.n82 VN.n81 24.5923
R79 VN.n40 VN.n0 21.6413
R80 VN.n83 VN.n43 21.6413
R81 VN.n21 VN.t9 18.013
R82 VN.n10 VN.t6 18.013
R83 VN.n32 VN.t5 18.013
R84 VN.n0 VN.t0 18.013
R85 VN.n64 VN.t7 18.013
R86 VN.n53 VN.t2 18.013
R87 VN.n75 VN.t1 18.013
R88 VN.n43 VN.t3 18.013
R89 VN.n33 VN.n32 13.7719
R90 VN.n76 VN.n75 13.7719
R91 VN.n13 VN.n10 10.8209
R92 VN.n32 VN.n31 10.8209
R93 VN.n56 VN.n53 10.8209
R94 VN.n75 VN.n74 10.8209
R95 VN.n55 VN.n54 5.42647
R96 VN.n12 VN.n11 5.42647
R97 VN.n85 VN.n84 0.354861
R98 VN.n42 VN.n41 0.354861
R99 VN VN.n42 0.267071
R100 VN.n84 VN.n44 0.189894
R101 VN.n80 VN.n44 0.189894
R102 VN.n80 VN.n79 0.189894
R103 VN.n79 VN.n78 0.189894
R104 VN.n78 VN.n46 0.189894
R105 VN.n73 VN.n46 0.189894
R106 VN.n73 VN.n72 0.189894
R107 VN.n72 VN.n71 0.189894
R108 VN.n71 VN.n48 0.189894
R109 VN.n67 VN.n48 0.189894
R110 VN.n67 VN.n66 0.189894
R111 VN.n66 VN.n65 0.189894
R112 VN.n65 VN.n50 0.189894
R113 VN.n61 VN.n50 0.189894
R114 VN.n61 VN.n60 0.189894
R115 VN.n60 VN.n59 0.189894
R116 VN.n59 VN.n52 0.189894
R117 VN.n55 VN.n52 0.189894
R118 VN.n12 VN.n9 0.189894
R119 VN.n16 VN.n9 0.189894
R120 VN.n17 VN.n16 0.189894
R121 VN.n18 VN.n17 0.189894
R122 VN.n18 VN.n7 0.189894
R123 VN.n22 VN.n7 0.189894
R124 VN.n23 VN.n22 0.189894
R125 VN.n24 VN.n23 0.189894
R126 VN.n24 VN.n5 0.189894
R127 VN.n28 VN.n5 0.189894
R128 VN.n29 VN.n28 0.189894
R129 VN.n30 VN.n29 0.189894
R130 VN.n30 VN.n3 0.189894
R131 VN.n35 VN.n3 0.189894
R132 VN.n36 VN.n35 0.189894
R133 VN.n37 VN.n36 0.189894
R134 VN.n37 VN.n1 0.189894
R135 VN.n41 VN.n1 0.189894
R136 VTAIL.n17 VTAIL.t17 171.536
R137 VTAIL.n2 VTAIL.t19 171.536
R138 VTAIL.n16 VTAIL.t2 171.536
R139 VTAIL.n11 VTAIL.t18 171.536
R140 VTAIL.n15 VTAIL.n14 156.488
R141 VTAIL.n13 VTAIL.n12 156.488
R142 VTAIL.n10 VTAIL.n9 156.488
R143 VTAIL.n8 VTAIL.n7 156.488
R144 VTAIL.n19 VTAIL.n18 156.488
R145 VTAIL.n1 VTAIL.n0 156.488
R146 VTAIL.n4 VTAIL.n3 156.488
R147 VTAIL.n6 VTAIL.n5 156.488
R148 VTAIL.n8 VTAIL.n6 19.7807
R149 VTAIL.n17 VTAIL.n16 17.0048
R150 VTAIL.n18 VTAIL.t12 15.0491
R151 VTAIL.n18 VTAIL.t9 15.0491
R152 VTAIL.n0 VTAIL.t13 15.0491
R153 VTAIL.n0 VTAIL.t16 15.0491
R154 VTAIL.n3 VTAIL.t7 15.0491
R155 VTAIL.n3 VTAIL.t4 15.0491
R156 VTAIL.n5 VTAIL.t8 15.0491
R157 VTAIL.n5 VTAIL.t5 15.0491
R158 VTAIL.n14 VTAIL.t1 15.0491
R159 VTAIL.n14 VTAIL.t0 15.0491
R160 VTAIL.n12 VTAIL.t6 15.0491
R161 VTAIL.n12 VTAIL.t3 15.0491
R162 VTAIL.n9 VTAIL.t15 15.0491
R163 VTAIL.n9 VTAIL.t10 15.0491
R164 VTAIL.n7 VTAIL.t11 15.0491
R165 VTAIL.n7 VTAIL.t14 15.0491
R166 VTAIL.n10 VTAIL.n8 2.77636
R167 VTAIL.n11 VTAIL.n10 2.77636
R168 VTAIL.n15 VTAIL.n13 2.77636
R169 VTAIL.n16 VTAIL.n15 2.77636
R170 VTAIL.n6 VTAIL.n4 2.77636
R171 VTAIL.n4 VTAIL.n2 2.77636
R172 VTAIL.n19 VTAIL.n17 2.77636
R173 VTAIL VTAIL.n1 2.14059
R174 VTAIL.n13 VTAIL.n11 1.85826
R175 VTAIL.n2 VTAIL.n1 1.85826
R176 VTAIL VTAIL.n19 0.636276
R177 VDD2.n1 VDD2.t1 190.992
R178 VDD2.n4 VDD2.t6 188.215
R179 VDD2.n3 VDD2.n2 175.192
R180 VDD2 VDD2.n7 175.19
R181 VDD2.n6 VDD2.n5 173.167
R182 VDD2.n1 VDD2.n0 173.167
R183 VDD2.n4 VDD2.n3 38.7627
R184 VDD2.n7 VDD2.t7 15.0491
R185 VDD2.n7 VDD2.t5 15.0491
R186 VDD2.n5 VDD2.t8 15.0491
R187 VDD2.n5 VDD2.t2 15.0491
R188 VDD2.n2 VDD2.t4 15.0491
R189 VDD2.n2 VDD2.t9 15.0491
R190 VDD2.n0 VDD2.t3 15.0491
R191 VDD2.n0 VDD2.t0 15.0491
R192 VDD2.n6 VDD2.n4 2.77636
R193 VDD2 VDD2.n6 0.752655
R194 VDD2.n3 VDD2.n1 0.639119
R195 VP.n27 VP.n26 161.3
R196 VP.n28 VP.n23 161.3
R197 VP.n30 VP.n29 161.3
R198 VP.n31 VP.n22 161.3
R199 VP.n33 VP.n32 161.3
R200 VP.n34 VP.n21 161.3
R201 VP.n36 VP.n35 161.3
R202 VP.n37 VP.n20 161.3
R203 VP.n39 VP.n38 161.3
R204 VP.n40 VP.n19 161.3
R205 VP.n42 VP.n41 161.3
R206 VP.n43 VP.n18 161.3
R207 VP.n45 VP.n44 161.3
R208 VP.n47 VP.n17 161.3
R209 VP.n49 VP.n48 161.3
R210 VP.n50 VP.n16 161.3
R211 VP.n52 VP.n51 161.3
R212 VP.n53 VP.n15 161.3
R213 VP.n55 VP.n54 161.3
R214 VP.n97 VP.n96 161.3
R215 VP.n95 VP.n1 161.3
R216 VP.n94 VP.n93 161.3
R217 VP.n92 VP.n2 161.3
R218 VP.n91 VP.n90 161.3
R219 VP.n89 VP.n3 161.3
R220 VP.n87 VP.n86 161.3
R221 VP.n85 VP.n4 161.3
R222 VP.n84 VP.n83 161.3
R223 VP.n82 VP.n5 161.3
R224 VP.n81 VP.n80 161.3
R225 VP.n79 VP.n6 161.3
R226 VP.n78 VP.n77 161.3
R227 VP.n76 VP.n7 161.3
R228 VP.n75 VP.n74 161.3
R229 VP.n73 VP.n8 161.3
R230 VP.n72 VP.n71 161.3
R231 VP.n70 VP.n9 161.3
R232 VP.n69 VP.n68 161.3
R233 VP.n67 VP.n66 161.3
R234 VP.n65 VP.n11 161.3
R235 VP.n64 VP.n63 161.3
R236 VP.n62 VP.n12 161.3
R237 VP.n61 VP.n60 161.3
R238 VP.n59 VP.n13 161.3
R239 VP.n58 VP.n57 68.6047
R240 VP.n98 VP.n0 68.6047
R241 VP.n56 VP.n14 68.6047
R242 VP.n25 VP.n24 63.1738
R243 VP.n64 VP.n12 56.5617
R244 VP.n94 VP.n2 56.5617
R245 VP.n52 VP.n16 56.5617
R246 VP.n71 VP.n8 51.2335
R247 VP.n83 VP.n82 51.2335
R248 VP.n41 VP.n40 51.2335
R249 VP.n29 VP.n22 51.2335
R250 VP.n25 VP.t7 49.8397
R251 VP.n57 VP.n56 47.3556
R252 VP.n75 VP.n8 29.9206
R253 VP.n82 VP.n81 29.9206
R254 VP.n40 VP.n39 29.9206
R255 VP.n33 VP.n22 29.9206
R256 VP.n60 VP.n59 24.5923
R257 VP.n60 VP.n12 24.5923
R258 VP.n65 VP.n64 24.5923
R259 VP.n66 VP.n65 24.5923
R260 VP.n70 VP.n69 24.5923
R261 VP.n71 VP.n70 24.5923
R262 VP.n76 VP.n75 24.5923
R263 VP.n77 VP.n76 24.5923
R264 VP.n77 VP.n6 24.5923
R265 VP.n81 VP.n6 24.5923
R266 VP.n83 VP.n4 24.5923
R267 VP.n87 VP.n4 24.5923
R268 VP.n90 VP.n89 24.5923
R269 VP.n90 VP.n2 24.5923
R270 VP.n95 VP.n94 24.5923
R271 VP.n96 VP.n95 24.5923
R272 VP.n53 VP.n52 24.5923
R273 VP.n54 VP.n53 24.5923
R274 VP.n41 VP.n18 24.5923
R275 VP.n45 VP.n18 24.5923
R276 VP.n48 VP.n47 24.5923
R277 VP.n48 VP.n16 24.5923
R278 VP.n34 VP.n33 24.5923
R279 VP.n35 VP.n34 24.5923
R280 VP.n35 VP.n20 24.5923
R281 VP.n39 VP.n20 24.5923
R282 VP.n28 VP.n27 24.5923
R283 VP.n29 VP.n28 24.5923
R284 VP.n59 VP.n58 21.6413
R285 VP.n96 VP.n0 21.6413
R286 VP.n54 VP.n14 21.6413
R287 VP.n77 VP.t8 18.013
R288 VP.n58 VP.t6 18.013
R289 VP.n10 VP.t4 18.013
R290 VP.n88 VP.t5 18.013
R291 VP.n0 VP.t0 18.013
R292 VP.n35 VP.t2 18.013
R293 VP.n14 VP.t9 18.013
R294 VP.n46 VP.t1 18.013
R295 VP.n24 VP.t3 18.013
R296 VP.n66 VP.n10 13.7719
R297 VP.n89 VP.n88 13.7719
R298 VP.n47 VP.n46 13.7719
R299 VP.n69 VP.n10 10.8209
R300 VP.n88 VP.n87 10.8209
R301 VP.n46 VP.n45 10.8209
R302 VP.n27 VP.n24 10.8209
R303 VP.n26 VP.n25 5.42643
R304 VP.n56 VP.n55 0.354861
R305 VP.n57 VP.n13 0.354861
R306 VP.n98 VP.n97 0.354861
R307 VP VP.n98 0.267071
R308 VP.n26 VP.n23 0.189894
R309 VP.n30 VP.n23 0.189894
R310 VP.n31 VP.n30 0.189894
R311 VP.n32 VP.n31 0.189894
R312 VP.n32 VP.n21 0.189894
R313 VP.n36 VP.n21 0.189894
R314 VP.n37 VP.n36 0.189894
R315 VP.n38 VP.n37 0.189894
R316 VP.n38 VP.n19 0.189894
R317 VP.n42 VP.n19 0.189894
R318 VP.n43 VP.n42 0.189894
R319 VP.n44 VP.n43 0.189894
R320 VP.n44 VP.n17 0.189894
R321 VP.n49 VP.n17 0.189894
R322 VP.n50 VP.n49 0.189894
R323 VP.n51 VP.n50 0.189894
R324 VP.n51 VP.n15 0.189894
R325 VP.n55 VP.n15 0.189894
R326 VP.n61 VP.n13 0.189894
R327 VP.n62 VP.n61 0.189894
R328 VP.n63 VP.n62 0.189894
R329 VP.n63 VP.n11 0.189894
R330 VP.n67 VP.n11 0.189894
R331 VP.n68 VP.n67 0.189894
R332 VP.n68 VP.n9 0.189894
R333 VP.n72 VP.n9 0.189894
R334 VP.n73 VP.n72 0.189894
R335 VP.n74 VP.n73 0.189894
R336 VP.n74 VP.n7 0.189894
R337 VP.n78 VP.n7 0.189894
R338 VP.n79 VP.n78 0.189894
R339 VP.n80 VP.n79 0.189894
R340 VP.n80 VP.n5 0.189894
R341 VP.n84 VP.n5 0.189894
R342 VP.n85 VP.n84 0.189894
R343 VP.n86 VP.n85 0.189894
R344 VP.n86 VP.n3 0.189894
R345 VP.n91 VP.n3 0.189894
R346 VP.n92 VP.n91 0.189894
R347 VP.n93 VP.n92 0.189894
R348 VP.n93 VP.n1 0.189894
R349 VP.n97 VP.n1 0.189894
R350 VDD1.n3 VDD1.t3 190.992
R351 VDD1.n1 VDD1.t2 190.99
R352 VDD1.n5 VDD1.n4 175.192
R353 VDD1.n1 VDD1.n0 173.167
R354 VDD1.n7 VDD1.n6 173.167
R355 VDD1.n3 VDD1.n2 173.167
R356 VDD1.n7 VDD1.n5 40.7337
R357 VDD1.n6 VDD1.t8 15.0491
R358 VDD1.n6 VDD1.t0 15.0491
R359 VDD1.n0 VDD1.t6 15.0491
R360 VDD1.n0 VDD1.t7 15.0491
R361 VDD1.n4 VDD1.t4 15.0491
R362 VDD1.n4 VDD1.t9 15.0491
R363 VDD1.n2 VDD1.t5 15.0491
R364 VDD1.n2 VDD1.t1 15.0491
R365 VDD1 VDD1.n7 2.02421
R366 VDD1 VDD1.n1 0.752655
R367 VDD1.n5 VDD1.n3 0.639119
R368 B.n523 B.n522 585
R369 B.n524 B.n55 585
R370 B.n526 B.n525 585
R371 B.n527 B.n54 585
R372 B.n529 B.n528 585
R373 B.n530 B.n53 585
R374 B.n532 B.n531 585
R375 B.n533 B.n52 585
R376 B.n535 B.n534 585
R377 B.n536 B.n51 585
R378 B.n538 B.n537 585
R379 B.n539 B.n50 585
R380 B.n541 B.n540 585
R381 B.n543 B.n47 585
R382 B.n545 B.n544 585
R383 B.n546 B.n46 585
R384 B.n548 B.n547 585
R385 B.n549 B.n45 585
R386 B.n551 B.n550 585
R387 B.n552 B.n44 585
R388 B.n554 B.n553 585
R389 B.n555 B.n41 585
R390 B.n558 B.n557 585
R391 B.n559 B.n40 585
R392 B.n561 B.n560 585
R393 B.n562 B.n39 585
R394 B.n564 B.n563 585
R395 B.n565 B.n38 585
R396 B.n567 B.n566 585
R397 B.n568 B.n37 585
R398 B.n570 B.n569 585
R399 B.n571 B.n36 585
R400 B.n573 B.n572 585
R401 B.n574 B.n35 585
R402 B.n576 B.n575 585
R403 B.n521 B.n56 585
R404 B.n520 B.n519 585
R405 B.n518 B.n57 585
R406 B.n517 B.n516 585
R407 B.n515 B.n58 585
R408 B.n514 B.n513 585
R409 B.n512 B.n59 585
R410 B.n511 B.n510 585
R411 B.n509 B.n60 585
R412 B.n508 B.n507 585
R413 B.n506 B.n61 585
R414 B.n505 B.n504 585
R415 B.n503 B.n62 585
R416 B.n502 B.n501 585
R417 B.n500 B.n63 585
R418 B.n499 B.n498 585
R419 B.n497 B.n64 585
R420 B.n496 B.n495 585
R421 B.n494 B.n65 585
R422 B.n493 B.n492 585
R423 B.n491 B.n66 585
R424 B.n490 B.n489 585
R425 B.n488 B.n67 585
R426 B.n487 B.n486 585
R427 B.n485 B.n68 585
R428 B.n484 B.n483 585
R429 B.n482 B.n69 585
R430 B.n481 B.n480 585
R431 B.n479 B.n70 585
R432 B.n478 B.n477 585
R433 B.n476 B.n71 585
R434 B.n475 B.n474 585
R435 B.n473 B.n72 585
R436 B.n472 B.n471 585
R437 B.n470 B.n73 585
R438 B.n469 B.n468 585
R439 B.n467 B.n74 585
R440 B.n466 B.n465 585
R441 B.n464 B.n75 585
R442 B.n463 B.n462 585
R443 B.n461 B.n76 585
R444 B.n460 B.n459 585
R445 B.n458 B.n77 585
R446 B.n457 B.n456 585
R447 B.n455 B.n78 585
R448 B.n454 B.n453 585
R449 B.n452 B.n79 585
R450 B.n451 B.n450 585
R451 B.n449 B.n80 585
R452 B.n448 B.n447 585
R453 B.n446 B.n81 585
R454 B.n445 B.n444 585
R455 B.n443 B.n82 585
R456 B.n442 B.n441 585
R457 B.n440 B.n83 585
R458 B.n439 B.n438 585
R459 B.n437 B.n84 585
R460 B.n436 B.n435 585
R461 B.n434 B.n85 585
R462 B.n433 B.n432 585
R463 B.n431 B.n86 585
R464 B.n430 B.n429 585
R465 B.n428 B.n87 585
R466 B.n427 B.n426 585
R467 B.n425 B.n88 585
R468 B.n424 B.n423 585
R469 B.n422 B.n89 585
R470 B.n421 B.n420 585
R471 B.n419 B.n90 585
R472 B.n418 B.n417 585
R473 B.n416 B.n91 585
R474 B.n415 B.n414 585
R475 B.n413 B.n92 585
R476 B.n412 B.n411 585
R477 B.n410 B.n93 585
R478 B.n409 B.n408 585
R479 B.n407 B.n94 585
R480 B.n406 B.n405 585
R481 B.n404 B.n95 585
R482 B.n403 B.n402 585
R483 B.n401 B.n96 585
R484 B.n400 B.n399 585
R485 B.n398 B.n97 585
R486 B.n397 B.n396 585
R487 B.n395 B.n98 585
R488 B.n394 B.n393 585
R489 B.n392 B.n99 585
R490 B.n391 B.n390 585
R491 B.n389 B.n100 585
R492 B.n388 B.n387 585
R493 B.n386 B.n101 585
R494 B.n385 B.n384 585
R495 B.n383 B.n102 585
R496 B.n382 B.n381 585
R497 B.n380 B.n103 585
R498 B.n379 B.n378 585
R499 B.n377 B.n104 585
R500 B.n376 B.n375 585
R501 B.n374 B.n105 585
R502 B.n373 B.n372 585
R503 B.n371 B.n106 585
R504 B.n370 B.n369 585
R505 B.n368 B.n107 585
R506 B.n367 B.n366 585
R507 B.n365 B.n108 585
R508 B.n364 B.n363 585
R509 B.n362 B.n109 585
R510 B.n361 B.n360 585
R511 B.n359 B.n110 585
R512 B.n358 B.n357 585
R513 B.n356 B.n111 585
R514 B.n355 B.n354 585
R515 B.n353 B.n112 585
R516 B.n352 B.n351 585
R517 B.n350 B.n113 585
R518 B.n349 B.n348 585
R519 B.n347 B.n114 585
R520 B.n346 B.n345 585
R521 B.n344 B.n115 585
R522 B.n343 B.n342 585
R523 B.n341 B.n116 585
R524 B.n340 B.n339 585
R525 B.n338 B.n117 585
R526 B.n337 B.n336 585
R527 B.n335 B.n118 585
R528 B.n334 B.n333 585
R529 B.n332 B.n119 585
R530 B.n331 B.n330 585
R531 B.n329 B.n120 585
R532 B.n328 B.n327 585
R533 B.n326 B.n121 585
R534 B.n272 B.n143 585
R535 B.n274 B.n273 585
R536 B.n275 B.n142 585
R537 B.n277 B.n276 585
R538 B.n278 B.n141 585
R539 B.n280 B.n279 585
R540 B.n281 B.n140 585
R541 B.n283 B.n282 585
R542 B.n284 B.n139 585
R543 B.n286 B.n285 585
R544 B.n287 B.n138 585
R545 B.n289 B.n288 585
R546 B.n290 B.n135 585
R547 B.n293 B.n292 585
R548 B.n294 B.n134 585
R549 B.n296 B.n295 585
R550 B.n297 B.n133 585
R551 B.n299 B.n298 585
R552 B.n300 B.n132 585
R553 B.n302 B.n301 585
R554 B.n303 B.n131 585
R555 B.n305 B.n304 585
R556 B.n307 B.n306 585
R557 B.n308 B.n127 585
R558 B.n310 B.n309 585
R559 B.n311 B.n126 585
R560 B.n313 B.n312 585
R561 B.n314 B.n125 585
R562 B.n316 B.n315 585
R563 B.n317 B.n124 585
R564 B.n319 B.n318 585
R565 B.n320 B.n123 585
R566 B.n322 B.n321 585
R567 B.n323 B.n122 585
R568 B.n325 B.n324 585
R569 B.n271 B.n270 585
R570 B.n269 B.n144 585
R571 B.n268 B.n267 585
R572 B.n266 B.n145 585
R573 B.n265 B.n264 585
R574 B.n263 B.n146 585
R575 B.n262 B.n261 585
R576 B.n260 B.n147 585
R577 B.n259 B.n258 585
R578 B.n257 B.n148 585
R579 B.n256 B.n255 585
R580 B.n254 B.n149 585
R581 B.n253 B.n252 585
R582 B.n251 B.n150 585
R583 B.n250 B.n249 585
R584 B.n248 B.n151 585
R585 B.n247 B.n246 585
R586 B.n245 B.n152 585
R587 B.n244 B.n243 585
R588 B.n242 B.n153 585
R589 B.n241 B.n240 585
R590 B.n239 B.n154 585
R591 B.n238 B.n237 585
R592 B.n236 B.n155 585
R593 B.n235 B.n234 585
R594 B.n233 B.n156 585
R595 B.n232 B.n231 585
R596 B.n230 B.n157 585
R597 B.n229 B.n228 585
R598 B.n227 B.n158 585
R599 B.n226 B.n225 585
R600 B.n224 B.n159 585
R601 B.n223 B.n222 585
R602 B.n221 B.n160 585
R603 B.n220 B.n219 585
R604 B.n218 B.n161 585
R605 B.n217 B.n216 585
R606 B.n215 B.n162 585
R607 B.n214 B.n213 585
R608 B.n212 B.n163 585
R609 B.n211 B.n210 585
R610 B.n209 B.n164 585
R611 B.n208 B.n207 585
R612 B.n206 B.n165 585
R613 B.n205 B.n204 585
R614 B.n203 B.n166 585
R615 B.n202 B.n201 585
R616 B.n200 B.n167 585
R617 B.n199 B.n198 585
R618 B.n197 B.n168 585
R619 B.n196 B.n195 585
R620 B.n194 B.n169 585
R621 B.n193 B.n192 585
R622 B.n191 B.n170 585
R623 B.n190 B.n189 585
R624 B.n188 B.n171 585
R625 B.n187 B.n186 585
R626 B.n185 B.n172 585
R627 B.n184 B.n183 585
R628 B.n182 B.n173 585
R629 B.n181 B.n180 585
R630 B.n179 B.n174 585
R631 B.n178 B.n177 585
R632 B.n176 B.n175 585
R633 B.n2 B.n0 585
R634 B.n673 B.n1 585
R635 B.n672 B.n671 585
R636 B.n670 B.n3 585
R637 B.n669 B.n668 585
R638 B.n667 B.n4 585
R639 B.n666 B.n665 585
R640 B.n664 B.n5 585
R641 B.n663 B.n662 585
R642 B.n661 B.n6 585
R643 B.n660 B.n659 585
R644 B.n658 B.n7 585
R645 B.n657 B.n656 585
R646 B.n655 B.n8 585
R647 B.n654 B.n653 585
R648 B.n652 B.n9 585
R649 B.n651 B.n650 585
R650 B.n649 B.n10 585
R651 B.n648 B.n647 585
R652 B.n646 B.n11 585
R653 B.n645 B.n644 585
R654 B.n643 B.n12 585
R655 B.n642 B.n641 585
R656 B.n640 B.n13 585
R657 B.n639 B.n638 585
R658 B.n637 B.n14 585
R659 B.n636 B.n635 585
R660 B.n634 B.n15 585
R661 B.n633 B.n632 585
R662 B.n631 B.n16 585
R663 B.n630 B.n629 585
R664 B.n628 B.n17 585
R665 B.n627 B.n626 585
R666 B.n625 B.n18 585
R667 B.n624 B.n623 585
R668 B.n622 B.n19 585
R669 B.n621 B.n620 585
R670 B.n619 B.n20 585
R671 B.n618 B.n617 585
R672 B.n616 B.n21 585
R673 B.n615 B.n614 585
R674 B.n613 B.n22 585
R675 B.n612 B.n611 585
R676 B.n610 B.n23 585
R677 B.n609 B.n608 585
R678 B.n607 B.n24 585
R679 B.n606 B.n605 585
R680 B.n604 B.n25 585
R681 B.n603 B.n602 585
R682 B.n601 B.n26 585
R683 B.n600 B.n599 585
R684 B.n598 B.n27 585
R685 B.n597 B.n596 585
R686 B.n595 B.n28 585
R687 B.n594 B.n593 585
R688 B.n592 B.n29 585
R689 B.n591 B.n590 585
R690 B.n589 B.n30 585
R691 B.n588 B.n587 585
R692 B.n586 B.n31 585
R693 B.n585 B.n584 585
R694 B.n583 B.n32 585
R695 B.n582 B.n581 585
R696 B.n580 B.n33 585
R697 B.n579 B.n578 585
R698 B.n577 B.n34 585
R699 B.n675 B.n674 585
R700 B.n270 B.n143 482.89
R701 B.n577 B.n576 482.89
R702 B.n324 B.n121 482.89
R703 B.n522 B.n521 482.89
R704 B.n128 B.t2 234.794
R705 B.n48 B.t4 234.794
R706 B.n136 B.t8 234.794
R707 B.n42 B.t10 234.794
R708 B.n128 B.t0 226.458
R709 B.n136 B.t6 226.458
R710 B.n42 B.t9 226.458
R711 B.n48 B.t3 226.458
R712 B.n129 B.t1 172.345
R713 B.n49 B.t5 172.345
R714 B.n137 B.t7 172.345
R715 B.n43 B.t11 172.345
R716 B.n270 B.n269 163.367
R717 B.n269 B.n268 163.367
R718 B.n268 B.n145 163.367
R719 B.n264 B.n145 163.367
R720 B.n264 B.n263 163.367
R721 B.n263 B.n262 163.367
R722 B.n262 B.n147 163.367
R723 B.n258 B.n147 163.367
R724 B.n258 B.n257 163.367
R725 B.n257 B.n256 163.367
R726 B.n256 B.n149 163.367
R727 B.n252 B.n149 163.367
R728 B.n252 B.n251 163.367
R729 B.n251 B.n250 163.367
R730 B.n250 B.n151 163.367
R731 B.n246 B.n151 163.367
R732 B.n246 B.n245 163.367
R733 B.n245 B.n244 163.367
R734 B.n244 B.n153 163.367
R735 B.n240 B.n153 163.367
R736 B.n240 B.n239 163.367
R737 B.n239 B.n238 163.367
R738 B.n238 B.n155 163.367
R739 B.n234 B.n155 163.367
R740 B.n234 B.n233 163.367
R741 B.n233 B.n232 163.367
R742 B.n232 B.n157 163.367
R743 B.n228 B.n157 163.367
R744 B.n228 B.n227 163.367
R745 B.n227 B.n226 163.367
R746 B.n226 B.n159 163.367
R747 B.n222 B.n159 163.367
R748 B.n222 B.n221 163.367
R749 B.n221 B.n220 163.367
R750 B.n220 B.n161 163.367
R751 B.n216 B.n161 163.367
R752 B.n216 B.n215 163.367
R753 B.n215 B.n214 163.367
R754 B.n214 B.n163 163.367
R755 B.n210 B.n163 163.367
R756 B.n210 B.n209 163.367
R757 B.n209 B.n208 163.367
R758 B.n208 B.n165 163.367
R759 B.n204 B.n165 163.367
R760 B.n204 B.n203 163.367
R761 B.n203 B.n202 163.367
R762 B.n202 B.n167 163.367
R763 B.n198 B.n167 163.367
R764 B.n198 B.n197 163.367
R765 B.n197 B.n196 163.367
R766 B.n196 B.n169 163.367
R767 B.n192 B.n169 163.367
R768 B.n192 B.n191 163.367
R769 B.n191 B.n190 163.367
R770 B.n190 B.n171 163.367
R771 B.n186 B.n171 163.367
R772 B.n186 B.n185 163.367
R773 B.n185 B.n184 163.367
R774 B.n184 B.n173 163.367
R775 B.n180 B.n173 163.367
R776 B.n180 B.n179 163.367
R777 B.n179 B.n178 163.367
R778 B.n178 B.n175 163.367
R779 B.n175 B.n2 163.367
R780 B.n674 B.n2 163.367
R781 B.n674 B.n673 163.367
R782 B.n673 B.n672 163.367
R783 B.n672 B.n3 163.367
R784 B.n668 B.n3 163.367
R785 B.n668 B.n667 163.367
R786 B.n667 B.n666 163.367
R787 B.n666 B.n5 163.367
R788 B.n662 B.n5 163.367
R789 B.n662 B.n661 163.367
R790 B.n661 B.n660 163.367
R791 B.n660 B.n7 163.367
R792 B.n656 B.n7 163.367
R793 B.n656 B.n655 163.367
R794 B.n655 B.n654 163.367
R795 B.n654 B.n9 163.367
R796 B.n650 B.n9 163.367
R797 B.n650 B.n649 163.367
R798 B.n649 B.n648 163.367
R799 B.n648 B.n11 163.367
R800 B.n644 B.n11 163.367
R801 B.n644 B.n643 163.367
R802 B.n643 B.n642 163.367
R803 B.n642 B.n13 163.367
R804 B.n638 B.n13 163.367
R805 B.n638 B.n637 163.367
R806 B.n637 B.n636 163.367
R807 B.n636 B.n15 163.367
R808 B.n632 B.n15 163.367
R809 B.n632 B.n631 163.367
R810 B.n631 B.n630 163.367
R811 B.n630 B.n17 163.367
R812 B.n626 B.n17 163.367
R813 B.n626 B.n625 163.367
R814 B.n625 B.n624 163.367
R815 B.n624 B.n19 163.367
R816 B.n620 B.n19 163.367
R817 B.n620 B.n619 163.367
R818 B.n619 B.n618 163.367
R819 B.n618 B.n21 163.367
R820 B.n614 B.n21 163.367
R821 B.n614 B.n613 163.367
R822 B.n613 B.n612 163.367
R823 B.n612 B.n23 163.367
R824 B.n608 B.n23 163.367
R825 B.n608 B.n607 163.367
R826 B.n607 B.n606 163.367
R827 B.n606 B.n25 163.367
R828 B.n602 B.n25 163.367
R829 B.n602 B.n601 163.367
R830 B.n601 B.n600 163.367
R831 B.n600 B.n27 163.367
R832 B.n596 B.n27 163.367
R833 B.n596 B.n595 163.367
R834 B.n595 B.n594 163.367
R835 B.n594 B.n29 163.367
R836 B.n590 B.n29 163.367
R837 B.n590 B.n589 163.367
R838 B.n589 B.n588 163.367
R839 B.n588 B.n31 163.367
R840 B.n584 B.n31 163.367
R841 B.n584 B.n583 163.367
R842 B.n583 B.n582 163.367
R843 B.n582 B.n33 163.367
R844 B.n578 B.n33 163.367
R845 B.n578 B.n577 163.367
R846 B.n274 B.n143 163.367
R847 B.n275 B.n274 163.367
R848 B.n276 B.n275 163.367
R849 B.n276 B.n141 163.367
R850 B.n280 B.n141 163.367
R851 B.n281 B.n280 163.367
R852 B.n282 B.n281 163.367
R853 B.n282 B.n139 163.367
R854 B.n286 B.n139 163.367
R855 B.n287 B.n286 163.367
R856 B.n288 B.n287 163.367
R857 B.n288 B.n135 163.367
R858 B.n293 B.n135 163.367
R859 B.n294 B.n293 163.367
R860 B.n295 B.n294 163.367
R861 B.n295 B.n133 163.367
R862 B.n299 B.n133 163.367
R863 B.n300 B.n299 163.367
R864 B.n301 B.n300 163.367
R865 B.n301 B.n131 163.367
R866 B.n305 B.n131 163.367
R867 B.n306 B.n305 163.367
R868 B.n306 B.n127 163.367
R869 B.n310 B.n127 163.367
R870 B.n311 B.n310 163.367
R871 B.n312 B.n311 163.367
R872 B.n312 B.n125 163.367
R873 B.n316 B.n125 163.367
R874 B.n317 B.n316 163.367
R875 B.n318 B.n317 163.367
R876 B.n318 B.n123 163.367
R877 B.n322 B.n123 163.367
R878 B.n323 B.n322 163.367
R879 B.n324 B.n323 163.367
R880 B.n328 B.n121 163.367
R881 B.n329 B.n328 163.367
R882 B.n330 B.n329 163.367
R883 B.n330 B.n119 163.367
R884 B.n334 B.n119 163.367
R885 B.n335 B.n334 163.367
R886 B.n336 B.n335 163.367
R887 B.n336 B.n117 163.367
R888 B.n340 B.n117 163.367
R889 B.n341 B.n340 163.367
R890 B.n342 B.n341 163.367
R891 B.n342 B.n115 163.367
R892 B.n346 B.n115 163.367
R893 B.n347 B.n346 163.367
R894 B.n348 B.n347 163.367
R895 B.n348 B.n113 163.367
R896 B.n352 B.n113 163.367
R897 B.n353 B.n352 163.367
R898 B.n354 B.n353 163.367
R899 B.n354 B.n111 163.367
R900 B.n358 B.n111 163.367
R901 B.n359 B.n358 163.367
R902 B.n360 B.n359 163.367
R903 B.n360 B.n109 163.367
R904 B.n364 B.n109 163.367
R905 B.n365 B.n364 163.367
R906 B.n366 B.n365 163.367
R907 B.n366 B.n107 163.367
R908 B.n370 B.n107 163.367
R909 B.n371 B.n370 163.367
R910 B.n372 B.n371 163.367
R911 B.n372 B.n105 163.367
R912 B.n376 B.n105 163.367
R913 B.n377 B.n376 163.367
R914 B.n378 B.n377 163.367
R915 B.n378 B.n103 163.367
R916 B.n382 B.n103 163.367
R917 B.n383 B.n382 163.367
R918 B.n384 B.n383 163.367
R919 B.n384 B.n101 163.367
R920 B.n388 B.n101 163.367
R921 B.n389 B.n388 163.367
R922 B.n390 B.n389 163.367
R923 B.n390 B.n99 163.367
R924 B.n394 B.n99 163.367
R925 B.n395 B.n394 163.367
R926 B.n396 B.n395 163.367
R927 B.n396 B.n97 163.367
R928 B.n400 B.n97 163.367
R929 B.n401 B.n400 163.367
R930 B.n402 B.n401 163.367
R931 B.n402 B.n95 163.367
R932 B.n406 B.n95 163.367
R933 B.n407 B.n406 163.367
R934 B.n408 B.n407 163.367
R935 B.n408 B.n93 163.367
R936 B.n412 B.n93 163.367
R937 B.n413 B.n412 163.367
R938 B.n414 B.n413 163.367
R939 B.n414 B.n91 163.367
R940 B.n418 B.n91 163.367
R941 B.n419 B.n418 163.367
R942 B.n420 B.n419 163.367
R943 B.n420 B.n89 163.367
R944 B.n424 B.n89 163.367
R945 B.n425 B.n424 163.367
R946 B.n426 B.n425 163.367
R947 B.n426 B.n87 163.367
R948 B.n430 B.n87 163.367
R949 B.n431 B.n430 163.367
R950 B.n432 B.n431 163.367
R951 B.n432 B.n85 163.367
R952 B.n436 B.n85 163.367
R953 B.n437 B.n436 163.367
R954 B.n438 B.n437 163.367
R955 B.n438 B.n83 163.367
R956 B.n442 B.n83 163.367
R957 B.n443 B.n442 163.367
R958 B.n444 B.n443 163.367
R959 B.n444 B.n81 163.367
R960 B.n448 B.n81 163.367
R961 B.n449 B.n448 163.367
R962 B.n450 B.n449 163.367
R963 B.n450 B.n79 163.367
R964 B.n454 B.n79 163.367
R965 B.n455 B.n454 163.367
R966 B.n456 B.n455 163.367
R967 B.n456 B.n77 163.367
R968 B.n460 B.n77 163.367
R969 B.n461 B.n460 163.367
R970 B.n462 B.n461 163.367
R971 B.n462 B.n75 163.367
R972 B.n466 B.n75 163.367
R973 B.n467 B.n466 163.367
R974 B.n468 B.n467 163.367
R975 B.n468 B.n73 163.367
R976 B.n472 B.n73 163.367
R977 B.n473 B.n472 163.367
R978 B.n474 B.n473 163.367
R979 B.n474 B.n71 163.367
R980 B.n478 B.n71 163.367
R981 B.n479 B.n478 163.367
R982 B.n480 B.n479 163.367
R983 B.n480 B.n69 163.367
R984 B.n484 B.n69 163.367
R985 B.n485 B.n484 163.367
R986 B.n486 B.n485 163.367
R987 B.n486 B.n67 163.367
R988 B.n490 B.n67 163.367
R989 B.n491 B.n490 163.367
R990 B.n492 B.n491 163.367
R991 B.n492 B.n65 163.367
R992 B.n496 B.n65 163.367
R993 B.n497 B.n496 163.367
R994 B.n498 B.n497 163.367
R995 B.n498 B.n63 163.367
R996 B.n502 B.n63 163.367
R997 B.n503 B.n502 163.367
R998 B.n504 B.n503 163.367
R999 B.n504 B.n61 163.367
R1000 B.n508 B.n61 163.367
R1001 B.n509 B.n508 163.367
R1002 B.n510 B.n509 163.367
R1003 B.n510 B.n59 163.367
R1004 B.n514 B.n59 163.367
R1005 B.n515 B.n514 163.367
R1006 B.n516 B.n515 163.367
R1007 B.n516 B.n57 163.367
R1008 B.n520 B.n57 163.367
R1009 B.n521 B.n520 163.367
R1010 B.n576 B.n35 163.367
R1011 B.n572 B.n35 163.367
R1012 B.n572 B.n571 163.367
R1013 B.n571 B.n570 163.367
R1014 B.n570 B.n37 163.367
R1015 B.n566 B.n37 163.367
R1016 B.n566 B.n565 163.367
R1017 B.n565 B.n564 163.367
R1018 B.n564 B.n39 163.367
R1019 B.n560 B.n39 163.367
R1020 B.n560 B.n559 163.367
R1021 B.n559 B.n558 163.367
R1022 B.n558 B.n41 163.367
R1023 B.n553 B.n41 163.367
R1024 B.n553 B.n552 163.367
R1025 B.n552 B.n551 163.367
R1026 B.n551 B.n45 163.367
R1027 B.n547 B.n45 163.367
R1028 B.n547 B.n546 163.367
R1029 B.n546 B.n545 163.367
R1030 B.n545 B.n47 163.367
R1031 B.n540 B.n47 163.367
R1032 B.n540 B.n539 163.367
R1033 B.n539 B.n538 163.367
R1034 B.n538 B.n51 163.367
R1035 B.n534 B.n51 163.367
R1036 B.n534 B.n533 163.367
R1037 B.n533 B.n532 163.367
R1038 B.n532 B.n53 163.367
R1039 B.n528 B.n53 163.367
R1040 B.n528 B.n527 163.367
R1041 B.n527 B.n526 163.367
R1042 B.n526 B.n55 163.367
R1043 B.n522 B.n55 163.367
R1044 B.n129 B.n128 62.449
R1045 B.n137 B.n136 62.449
R1046 B.n43 B.n42 62.449
R1047 B.n49 B.n48 62.449
R1048 B.n130 B.n129 59.5399
R1049 B.n291 B.n137 59.5399
R1050 B.n556 B.n43 59.5399
R1051 B.n542 B.n49 59.5399
R1052 B.n575 B.n34 31.3761
R1053 B.n523 B.n56 31.3761
R1054 B.n326 B.n325 31.3761
R1055 B.n272 B.n271 31.3761
R1056 B B.n675 18.0485
R1057 B.n575 B.n574 10.6151
R1058 B.n574 B.n573 10.6151
R1059 B.n573 B.n36 10.6151
R1060 B.n569 B.n36 10.6151
R1061 B.n569 B.n568 10.6151
R1062 B.n568 B.n567 10.6151
R1063 B.n567 B.n38 10.6151
R1064 B.n563 B.n38 10.6151
R1065 B.n563 B.n562 10.6151
R1066 B.n562 B.n561 10.6151
R1067 B.n561 B.n40 10.6151
R1068 B.n557 B.n40 10.6151
R1069 B.n555 B.n554 10.6151
R1070 B.n554 B.n44 10.6151
R1071 B.n550 B.n44 10.6151
R1072 B.n550 B.n549 10.6151
R1073 B.n549 B.n548 10.6151
R1074 B.n548 B.n46 10.6151
R1075 B.n544 B.n46 10.6151
R1076 B.n544 B.n543 10.6151
R1077 B.n541 B.n50 10.6151
R1078 B.n537 B.n50 10.6151
R1079 B.n537 B.n536 10.6151
R1080 B.n536 B.n535 10.6151
R1081 B.n535 B.n52 10.6151
R1082 B.n531 B.n52 10.6151
R1083 B.n531 B.n530 10.6151
R1084 B.n530 B.n529 10.6151
R1085 B.n529 B.n54 10.6151
R1086 B.n525 B.n54 10.6151
R1087 B.n525 B.n524 10.6151
R1088 B.n524 B.n523 10.6151
R1089 B.n327 B.n326 10.6151
R1090 B.n327 B.n120 10.6151
R1091 B.n331 B.n120 10.6151
R1092 B.n332 B.n331 10.6151
R1093 B.n333 B.n332 10.6151
R1094 B.n333 B.n118 10.6151
R1095 B.n337 B.n118 10.6151
R1096 B.n338 B.n337 10.6151
R1097 B.n339 B.n338 10.6151
R1098 B.n339 B.n116 10.6151
R1099 B.n343 B.n116 10.6151
R1100 B.n344 B.n343 10.6151
R1101 B.n345 B.n344 10.6151
R1102 B.n345 B.n114 10.6151
R1103 B.n349 B.n114 10.6151
R1104 B.n350 B.n349 10.6151
R1105 B.n351 B.n350 10.6151
R1106 B.n351 B.n112 10.6151
R1107 B.n355 B.n112 10.6151
R1108 B.n356 B.n355 10.6151
R1109 B.n357 B.n356 10.6151
R1110 B.n357 B.n110 10.6151
R1111 B.n361 B.n110 10.6151
R1112 B.n362 B.n361 10.6151
R1113 B.n363 B.n362 10.6151
R1114 B.n363 B.n108 10.6151
R1115 B.n367 B.n108 10.6151
R1116 B.n368 B.n367 10.6151
R1117 B.n369 B.n368 10.6151
R1118 B.n369 B.n106 10.6151
R1119 B.n373 B.n106 10.6151
R1120 B.n374 B.n373 10.6151
R1121 B.n375 B.n374 10.6151
R1122 B.n375 B.n104 10.6151
R1123 B.n379 B.n104 10.6151
R1124 B.n380 B.n379 10.6151
R1125 B.n381 B.n380 10.6151
R1126 B.n381 B.n102 10.6151
R1127 B.n385 B.n102 10.6151
R1128 B.n386 B.n385 10.6151
R1129 B.n387 B.n386 10.6151
R1130 B.n387 B.n100 10.6151
R1131 B.n391 B.n100 10.6151
R1132 B.n392 B.n391 10.6151
R1133 B.n393 B.n392 10.6151
R1134 B.n393 B.n98 10.6151
R1135 B.n397 B.n98 10.6151
R1136 B.n398 B.n397 10.6151
R1137 B.n399 B.n398 10.6151
R1138 B.n399 B.n96 10.6151
R1139 B.n403 B.n96 10.6151
R1140 B.n404 B.n403 10.6151
R1141 B.n405 B.n404 10.6151
R1142 B.n405 B.n94 10.6151
R1143 B.n409 B.n94 10.6151
R1144 B.n410 B.n409 10.6151
R1145 B.n411 B.n410 10.6151
R1146 B.n411 B.n92 10.6151
R1147 B.n415 B.n92 10.6151
R1148 B.n416 B.n415 10.6151
R1149 B.n417 B.n416 10.6151
R1150 B.n417 B.n90 10.6151
R1151 B.n421 B.n90 10.6151
R1152 B.n422 B.n421 10.6151
R1153 B.n423 B.n422 10.6151
R1154 B.n423 B.n88 10.6151
R1155 B.n427 B.n88 10.6151
R1156 B.n428 B.n427 10.6151
R1157 B.n429 B.n428 10.6151
R1158 B.n429 B.n86 10.6151
R1159 B.n433 B.n86 10.6151
R1160 B.n434 B.n433 10.6151
R1161 B.n435 B.n434 10.6151
R1162 B.n435 B.n84 10.6151
R1163 B.n439 B.n84 10.6151
R1164 B.n440 B.n439 10.6151
R1165 B.n441 B.n440 10.6151
R1166 B.n441 B.n82 10.6151
R1167 B.n445 B.n82 10.6151
R1168 B.n446 B.n445 10.6151
R1169 B.n447 B.n446 10.6151
R1170 B.n447 B.n80 10.6151
R1171 B.n451 B.n80 10.6151
R1172 B.n452 B.n451 10.6151
R1173 B.n453 B.n452 10.6151
R1174 B.n453 B.n78 10.6151
R1175 B.n457 B.n78 10.6151
R1176 B.n458 B.n457 10.6151
R1177 B.n459 B.n458 10.6151
R1178 B.n459 B.n76 10.6151
R1179 B.n463 B.n76 10.6151
R1180 B.n464 B.n463 10.6151
R1181 B.n465 B.n464 10.6151
R1182 B.n465 B.n74 10.6151
R1183 B.n469 B.n74 10.6151
R1184 B.n470 B.n469 10.6151
R1185 B.n471 B.n470 10.6151
R1186 B.n471 B.n72 10.6151
R1187 B.n475 B.n72 10.6151
R1188 B.n476 B.n475 10.6151
R1189 B.n477 B.n476 10.6151
R1190 B.n477 B.n70 10.6151
R1191 B.n481 B.n70 10.6151
R1192 B.n482 B.n481 10.6151
R1193 B.n483 B.n482 10.6151
R1194 B.n483 B.n68 10.6151
R1195 B.n487 B.n68 10.6151
R1196 B.n488 B.n487 10.6151
R1197 B.n489 B.n488 10.6151
R1198 B.n489 B.n66 10.6151
R1199 B.n493 B.n66 10.6151
R1200 B.n494 B.n493 10.6151
R1201 B.n495 B.n494 10.6151
R1202 B.n495 B.n64 10.6151
R1203 B.n499 B.n64 10.6151
R1204 B.n500 B.n499 10.6151
R1205 B.n501 B.n500 10.6151
R1206 B.n501 B.n62 10.6151
R1207 B.n505 B.n62 10.6151
R1208 B.n506 B.n505 10.6151
R1209 B.n507 B.n506 10.6151
R1210 B.n507 B.n60 10.6151
R1211 B.n511 B.n60 10.6151
R1212 B.n512 B.n511 10.6151
R1213 B.n513 B.n512 10.6151
R1214 B.n513 B.n58 10.6151
R1215 B.n517 B.n58 10.6151
R1216 B.n518 B.n517 10.6151
R1217 B.n519 B.n518 10.6151
R1218 B.n519 B.n56 10.6151
R1219 B.n273 B.n272 10.6151
R1220 B.n273 B.n142 10.6151
R1221 B.n277 B.n142 10.6151
R1222 B.n278 B.n277 10.6151
R1223 B.n279 B.n278 10.6151
R1224 B.n279 B.n140 10.6151
R1225 B.n283 B.n140 10.6151
R1226 B.n284 B.n283 10.6151
R1227 B.n285 B.n284 10.6151
R1228 B.n285 B.n138 10.6151
R1229 B.n289 B.n138 10.6151
R1230 B.n290 B.n289 10.6151
R1231 B.n292 B.n134 10.6151
R1232 B.n296 B.n134 10.6151
R1233 B.n297 B.n296 10.6151
R1234 B.n298 B.n297 10.6151
R1235 B.n298 B.n132 10.6151
R1236 B.n302 B.n132 10.6151
R1237 B.n303 B.n302 10.6151
R1238 B.n304 B.n303 10.6151
R1239 B.n308 B.n307 10.6151
R1240 B.n309 B.n308 10.6151
R1241 B.n309 B.n126 10.6151
R1242 B.n313 B.n126 10.6151
R1243 B.n314 B.n313 10.6151
R1244 B.n315 B.n314 10.6151
R1245 B.n315 B.n124 10.6151
R1246 B.n319 B.n124 10.6151
R1247 B.n320 B.n319 10.6151
R1248 B.n321 B.n320 10.6151
R1249 B.n321 B.n122 10.6151
R1250 B.n325 B.n122 10.6151
R1251 B.n271 B.n144 10.6151
R1252 B.n267 B.n144 10.6151
R1253 B.n267 B.n266 10.6151
R1254 B.n266 B.n265 10.6151
R1255 B.n265 B.n146 10.6151
R1256 B.n261 B.n146 10.6151
R1257 B.n261 B.n260 10.6151
R1258 B.n260 B.n259 10.6151
R1259 B.n259 B.n148 10.6151
R1260 B.n255 B.n148 10.6151
R1261 B.n255 B.n254 10.6151
R1262 B.n254 B.n253 10.6151
R1263 B.n253 B.n150 10.6151
R1264 B.n249 B.n150 10.6151
R1265 B.n249 B.n248 10.6151
R1266 B.n248 B.n247 10.6151
R1267 B.n247 B.n152 10.6151
R1268 B.n243 B.n152 10.6151
R1269 B.n243 B.n242 10.6151
R1270 B.n242 B.n241 10.6151
R1271 B.n241 B.n154 10.6151
R1272 B.n237 B.n154 10.6151
R1273 B.n237 B.n236 10.6151
R1274 B.n236 B.n235 10.6151
R1275 B.n235 B.n156 10.6151
R1276 B.n231 B.n156 10.6151
R1277 B.n231 B.n230 10.6151
R1278 B.n230 B.n229 10.6151
R1279 B.n229 B.n158 10.6151
R1280 B.n225 B.n158 10.6151
R1281 B.n225 B.n224 10.6151
R1282 B.n224 B.n223 10.6151
R1283 B.n223 B.n160 10.6151
R1284 B.n219 B.n160 10.6151
R1285 B.n219 B.n218 10.6151
R1286 B.n218 B.n217 10.6151
R1287 B.n217 B.n162 10.6151
R1288 B.n213 B.n162 10.6151
R1289 B.n213 B.n212 10.6151
R1290 B.n212 B.n211 10.6151
R1291 B.n211 B.n164 10.6151
R1292 B.n207 B.n164 10.6151
R1293 B.n207 B.n206 10.6151
R1294 B.n206 B.n205 10.6151
R1295 B.n205 B.n166 10.6151
R1296 B.n201 B.n166 10.6151
R1297 B.n201 B.n200 10.6151
R1298 B.n200 B.n199 10.6151
R1299 B.n199 B.n168 10.6151
R1300 B.n195 B.n168 10.6151
R1301 B.n195 B.n194 10.6151
R1302 B.n194 B.n193 10.6151
R1303 B.n193 B.n170 10.6151
R1304 B.n189 B.n170 10.6151
R1305 B.n189 B.n188 10.6151
R1306 B.n188 B.n187 10.6151
R1307 B.n187 B.n172 10.6151
R1308 B.n183 B.n172 10.6151
R1309 B.n183 B.n182 10.6151
R1310 B.n182 B.n181 10.6151
R1311 B.n181 B.n174 10.6151
R1312 B.n177 B.n174 10.6151
R1313 B.n177 B.n176 10.6151
R1314 B.n176 B.n0 10.6151
R1315 B.n671 B.n1 10.6151
R1316 B.n671 B.n670 10.6151
R1317 B.n670 B.n669 10.6151
R1318 B.n669 B.n4 10.6151
R1319 B.n665 B.n4 10.6151
R1320 B.n665 B.n664 10.6151
R1321 B.n664 B.n663 10.6151
R1322 B.n663 B.n6 10.6151
R1323 B.n659 B.n6 10.6151
R1324 B.n659 B.n658 10.6151
R1325 B.n658 B.n657 10.6151
R1326 B.n657 B.n8 10.6151
R1327 B.n653 B.n8 10.6151
R1328 B.n653 B.n652 10.6151
R1329 B.n652 B.n651 10.6151
R1330 B.n651 B.n10 10.6151
R1331 B.n647 B.n10 10.6151
R1332 B.n647 B.n646 10.6151
R1333 B.n646 B.n645 10.6151
R1334 B.n645 B.n12 10.6151
R1335 B.n641 B.n12 10.6151
R1336 B.n641 B.n640 10.6151
R1337 B.n640 B.n639 10.6151
R1338 B.n639 B.n14 10.6151
R1339 B.n635 B.n14 10.6151
R1340 B.n635 B.n634 10.6151
R1341 B.n634 B.n633 10.6151
R1342 B.n633 B.n16 10.6151
R1343 B.n629 B.n16 10.6151
R1344 B.n629 B.n628 10.6151
R1345 B.n628 B.n627 10.6151
R1346 B.n627 B.n18 10.6151
R1347 B.n623 B.n18 10.6151
R1348 B.n623 B.n622 10.6151
R1349 B.n622 B.n621 10.6151
R1350 B.n621 B.n20 10.6151
R1351 B.n617 B.n20 10.6151
R1352 B.n617 B.n616 10.6151
R1353 B.n616 B.n615 10.6151
R1354 B.n615 B.n22 10.6151
R1355 B.n611 B.n22 10.6151
R1356 B.n611 B.n610 10.6151
R1357 B.n610 B.n609 10.6151
R1358 B.n609 B.n24 10.6151
R1359 B.n605 B.n24 10.6151
R1360 B.n605 B.n604 10.6151
R1361 B.n604 B.n603 10.6151
R1362 B.n603 B.n26 10.6151
R1363 B.n599 B.n26 10.6151
R1364 B.n599 B.n598 10.6151
R1365 B.n598 B.n597 10.6151
R1366 B.n597 B.n28 10.6151
R1367 B.n593 B.n28 10.6151
R1368 B.n593 B.n592 10.6151
R1369 B.n592 B.n591 10.6151
R1370 B.n591 B.n30 10.6151
R1371 B.n587 B.n30 10.6151
R1372 B.n587 B.n586 10.6151
R1373 B.n586 B.n585 10.6151
R1374 B.n585 B.n32 10.6151
R1375 B.n581 B.n32 10.6151
R1376 B.n581 B.n580 10.6151
R1377 B.n580 B.n579 10.6151
R1378 B.n579 B.n34 10.6151
R1379 B.n556 B.n555 6.5566
R1380 B.n543 B.n542 6.5566
R1381 B.n292 B.n291 6.5566
R1382 B.n304 B.n130 6.5566
R1383 B.n557 B.n556 4.05904
R1384 B.n542 B.n541 4.05904
R1385 B.n291 B.n290 4.05904
R1386 B.n307 B.n130 4.05904
R1387 B.n675 B.n0 2.81026
R1388 B.n675 B.n1 2.81026
C0 VTAIL VDD1 6.16625f
C1 VP B 2.32323f
C2 B w_n4834_n1400# 8.33391f
C3 VN B 1.26251f
C4 VP w_n4834_n1400# 10.8931f
C5 VN VP 7.0068f
C6 B VDD2 1.93966f
C7 VP VDD2 0.627797f
C8 B VDD1 1.81008f
C9 VN w_n4834_n1400# 10.266901f
C10 VP VDD1 2.85659f
C11 w_n4834_n1400# VDD2 2.37241f
C12 VN VDD2 2.3934f
C13 VTAIL B 1.50294f
C14 w_n4834_n1400# VDD1 2.21448f
C15 VN VDD1 0.160628f
C16 VTAIL VP 3.96568f
C17 VDD1 VDD2 2.36262f
C18 VTAIL w_n4834_n1400# 1.85025f
C19 VTAIL VN 3.95155f
C20 VTAIL VDD2 6.22149f
C21 VDD2 VSUBS 1.977645f
C22 VDD1 VSUBS 1.841978f
C23 VTAIL VSUBS 0.599448f
C24 VN VSUBS 8.332041f
C25 VP VSUBS 3.951606f
C26 B VSUBS 4.584121f
C27 w_n4834_n1400# VSUBS 86.2579f
C28 B.n0 VSUBS 0.006643f
C29 B.n1 VSUBS 0.006643f
C30 B.n2 VSUBS 0.010505f
C31 B.n3 VSUBS 0.010505f
C32 B.n4 VSUBS 0.010505f
C33 B.n5 VSUBS 0.010505f
C34 B.n6 VSUBS 0.010505f
C35 B.n7 VSUBS 0.010505f
C36 B.n8 VSUBS 0.010505f
C37 B.n9 VSUBS 0.010505f
C38 B.n10 VSUBS 0.010505f
C39 B.n11 VSUBS 0.010505f
C40 B.n12 VSUBS 0.010505f
C41 B.n13 VSUBS 0.010505f
C42 B.n14 VSUBS 0.010505f
C43 B.n15 VSUBS 0.010505f
C44 B.n16 VSUBS 0.010505f
C45 B.n17 VSUBS 0.010505f
C46 B.n18 VSUBS 0.010505f
C47 B.n19 VSUBS 0.010505f
C48 B.n20 VSUBS 0.010505f
C49 B.n21 VSUBS 0.010505f
C50 B.n22 VSUBS 0.010505f
C51 B.n23 VSUBS 0.010505f
C52 B.n24 VSUBS 0.010505f
C53 B.n25 VSUBS 0.010505f
C54 B.n26 VSUBS 0.010505f
C55 B.n27 VSUBS 0.010505f
C56 B.n28 VSUBS 0.010505f
C57 B.n29 VSUBS 0.010505f
C58 B.n30 VSUBS 0.010505f
C59 B.n31 VSUBS 0.010505f
C60 B.n32 VSUBS 0.010505f
C61 B.n33 VSUBS 0.010505f
C62 B.n34 VSUBS 0.023361f
C63 B.n35 VSUBS 0.010505f
C64 B.n36 VSUBS 0.010505f
C65 B.n37 VSUBS 0.010505f
C66 B.n38 VSUBS 0.010505f
C67 B.n39 VSUBS 0.010505f
C68 B.n40 VSUBS 0.010505f
C69 B.n41 VSUBS 0.010505f
C70 B.t11 VSUBS 0.071223f
C71 B.t10 VSUBS 0.091519f
C72 B.t9 VSUBS 0.461276f
C73 B.n42 VSUBS 0.113379f
C74 B.n43 VSUBS 0.091291f
C75 B.n44 VSUBS 0.010505f
C76 B.n45 VSUBS 0.010505f
C77 B.n46 VSUBS 0.010505f
C78 B.n47 VSUBS 0.010505f
C79 B.t5 VSUBS 0.071223f
C80 B.t4 VSUBS 0.091518f
C81 B.t3 VSUBS 0.461276f
C82 B.n48 VSUBS 0.113379f
C83 B.n49 VSUBS 0.091291f
C84 B.n50 VSUBS 0.010505f
C85 B.n51 VSUBS 0.010505f
C86 B.n52 VSUBS 0.010505f
C87 B.n53 VSUBS 0.010505f
C88 B.n54 VSUBS 0.010505f
C89 B.n55 VSUBS 0.010505f
C90 B.n56 VSUBS 0.024653f
C91 B.n57 VSUBS 0.010505f
C92 B.n58 VSUBS 0.010505f
C93 B.n59 VSUBS 0.010505f
C94 B.n60 VSUBS 0.010505f
C95 B.n61 VSUBS 0.010505f
C96 B.n62 VSUBS 0.010505f
C97 B.n63 VSUBS 0.010505f
C98 B.n64 VSUBS 0.010505f
C99 B.n65 VSUBS 0.010505f
C100 B.n66 VSUBS 0.010505f
C101 B.n67 VSUBS 0.010505f
C102 B.n68 VSUBS 0.010505f
C103 B.n69 VSUBS 0.010505f
C104 B.n70 VSUBS 0.010505f
C105 B.n71 VSUBS 0.010505f
C106 B.n72 VSUBS 0.010505f
C107 B.n73 VSUBS 0.010505f
C108 B.n74 VSUBS 0.010505f
C109 B.n75 VSUBS 0.010505f
C110 B.n76 VSUBS 0.010505f
C111 B.n77 VSUBS 0.010505f
C112 B.n78 VSUBS 0.010505f
C113 B.n79 VSUBS 0.010505f
C114 B.n80 VSUBS 0.010505f
C115 B.n81 VSUBS 0.010505f
C116 B.n82 VSUBS 0.010505f
C117 B.n83 VSUBS 0.010505f
C118 B.n84 VSUBS 0.010505f
C119 B.n85 VSUBS 0.010505f
C120 B.n86 VSUBS 0.010505f
C121 B.n87 VSUBS 0.010505f
C122 B.n88 VSUBS 0.010505f
C123 B.n89 VSUBS 0.010505f
C124 B.n90 VSUBS 0.010505f
C125 B.n91 VSUBS 0.010505f
C126 B.n92 VSUBS 0.010505f
C127 B.n93 VSUBS 0.010505f
C128 B.n94 VSUBS 0.010505f
C129 B.n95 VSUBS 0.010505f
C130 B.n96 VSUBS 0.010505f
C131 B.n97 VSUBS 0.010505f
C132 B.n98 VSUBS 0.010505f
C133 B.n99 VSUBS 0.010505f
C134 B.n100 VSUBS 0.010505f
C135 B.n101 VSUBS 0.010505f
C136 B.n102 VSUBS 0.010505f
C137 B.n103 VSUBS 0.010505f
C138 B.n104 VSUBS 0.010505f
C139 B.n105 VSUBS 0.010505f
C140 B.n106 VSUBS 0.010505f
C141 B.n107 VSUBS 0.010505f
C142 B.n108 VSUBS 0.010505f
C143 B.n109 VSUBS 0.010505f
C144 B.n110 VSUBS 0.010505f
C145 B.n111 VSUBS 0.010505f
C146 B.n112 VSUBS 0.010505f
C147 B.n113 VSUBS 0.010505f
C148 B.n114 VSUBS 0.010505f
C149 B.n115 VSUBS 0.010505f
C150 B.n116 VSUBS 0.010505f
C151 B.n117 VSUBS 0.010505f
C152 B.n118 VSUBS 0.010505f
C153 B.n119 VSUBS 0.010505f
C154 B.n120 VSUBS 0.010505f
C155 B.n121 VSUBS 0.023361f
C156 B.n122 VSUBS 0.010505f
C157 B.n123 VSUBS 0.010505f
C158 B.n124 VSUBS 0.010505f
C159 B.n125 VSUBS 0.010505f
C160 B.n126 VSUBS 0.010505f
C161 B.n127 VSUBS 0.010505f
C162 B.t1 VSUBS 0.071223f
C163 B.t2 VSUBS 0.091518f
C164 B.t0 VSUBS 0.461276f
C165 B.n128 VSUBS 0.113379f
C166 B.n129 VSUBS 0.091291f
C167 B.n130 VSUBS 0.024338f
C168 B.n131 VSUBS 0.010505f
C169 B.n132 VSUBS 0.010505f
C170 B.n133 VSUBS 0.010505f
C171 B.n134 VSUBS 0.010505f
C172 B.n135 VSUBS 0.010505f
C173 B.t7 VSUBS 0.071223f
C174 B.t8 VSUBS 0.091519f
C175 B.t6 VSUBS 0.461276f
C176 B.n136 VSUBS 0.113379f
C177 B.n137 VSUBS 0.091291f
C178 B.n138 VSUBS 0.010505f
C179 B.n139 VSUBS 0.010505f
C180 B.n140 VSUBS 0.010505f
C181 B.n141 VSUBS 0.010505f
C182 B.n142 VSUBS 0.010505f
C183 B.n143 VSUBS 0.024527f
C184 B.n144 VSUBS 0.010505f
C185 B.n145 VSUBS 0.010505f
C186 B.n146 VSUBS 0.010505f
C187 B.n147 VSUBS 0.010505f
C188 B.n148 VSUBS 0.010505f
C189 B.n149 VSUBS 0.010505f
C190 B.n150 VSUBS 0.010505f
C191 B.n151 VSUBS 0.010505f
C192 B.n152 VSUBS 0.010505f
C193 B.n153 VSUBS 0.010505f
C194 B.n154 VSUBS 0.010505f
C195 B.n155 VSUBS 0.010505f
C196 B.n156 VSUBS 0.010505f
C197 B.n157 VSUBS 0.010505f
C198 B.n158 VSUBS 0.010505f
C199 B.n159 VSUBS 0.010505f
C200 B.n160 VSUBS 0.010505f
C201 B.n161 VSUBS 0.010505f
C202 B.n162 VSUBS 0.010505f
C203 B.n163 VSUBS 0.010505f
C204 B.n164 VSUBS 0.010505f
C205 B.n165 VSUBS 0.010505f
C206 B.n166 VSUBS 0.010505f
C207 B.n167 VSUBS 0.010505f
C208 B.n168 VSUBS 0.010505f
C209 B.n169 VSUBS 0.010505f
C210 B.n170 VSUBS 0.010505f
C211 B.n171 VSUBS 0.010505f
C212 B.n172 VSUBS 0.010505f
C213 B.n173 VSUBS 0.010505f
C214 B.n174 VSUBS 0.010505f
C215 B.n175 VSUBS 0.010505f
C216 B.n176 VSUBS 0.010505f
C217 B.n177 VSUBS 0.010505f
C218 B.n178 VSUBS 0.010505f
C219 B.n179 VSUBS 0.010505f
C220 B.n180 VSUBS 0.010505f
C221 B.n181 VSUBS 0.010505f
C222 B.n182 VSUBS 0.010505f
C223 B.n183 VSUBS 0.010505f
C224 B.n184 VSUBS 0.010505f
C225 B.n185 VSUBS 0.010505f
C226 B.n186 VSUBS 0.010505f
C227 B.n187 VSUBS 0.010505f
C228 B.n188 VSUBS 0.010505f
C229 B.n189 VSUBS 0.010505f
C230 B.n190 VSUBS 0.010505f
C231 B.n191 VSUBS 0.010505f
C232 B.n192 VSUBS 0.010505f
C233 B.n193 VSUBS 0.010505f
C234 B.n194 VSUBS 0.010505f
C235 B.n195 VSUBS 0.010505f
C236 B.n196 VSUBS 0.010505f
C237 B.n197 VSUBS 0.010505f
C238 B.n198 VSUBS 0.010505f
C239 B.n199 VSUBS 0.010505f
C240 B.n200 VSUBS 0.010505f
C241 B.n201 VSUBS 0.010505f
C242 B.n202 VSUBS 0.010505f
C243 B.n203 VSUBS 0.010505f
C244 B.n204 VSUBS 0.010505f
C245 B.n205 VSUBS 0.010505f
C246 B.n206 VSUBS 0.010505f
C247 B.n207 VSUBS 0.010505f
C248 B.n208 VSUBS 0.010505f
C249 B.n209 VSUBS 0.010505f
C250 B.n210 VSUBS 0.010505f
C251 B.n211 VSUBS 0.010505f
C252 B.n212 VSUBS 0.010505f
C253 B.n213 VSUBS 0.010505f
C254 B.n214 VSUBS 0.010505f
C255 B.n215 VSUBS 0.010505f
C256 B.n216 VSUBS 0.010505f
C257 B.n217 VSUBS 0.010505f
C258 B.n218 VSUBS 0.010505f
C259 B.n219 VSUBS 0.010505f
C260 B.n220 VSUBS 0.010505f
C261 B.n221 VSUBS 0.010505f
C262 B.n222 VSUBS 0.010505f
C263 B.n223 VSUBS 0.010505f
C264 B.n224 VSUBS 0.010505f
C265 B.n225 VSUBS 0.010505f
C266 B.n226 VSUBS 0.010505f
C267 B.n227 VSUBS 0.010505f
C268 B.n228 VSUBS 0.010505f
C269 B.n229 VSUBS 0.010505f
C270 B.n230 VSUBS 0.010505f
C271 B.n231 VSUBS 0.010505f
C272 B.n232 VSUBS 0.010505f
C273 B.n233 VSUBS 0.010505f
C274 B.n234 VSUBS 0.010505f
C275 B.n235 VSUBS 0.010505f
C276 B.n236 VSUBS 0.010505f
C277 B.n237 VSUBS 0.010505f
C278 B.n238 VSUBS 0.010505f
C279 B.n239 VSUBS 0.010505f
C280 B.n240 VSUBS 0.010505f
C281 B.n241 VSUBS 0.010505f
C282 B.n242 VSUBS 0.010505f
C283 B.n243 VSUBS 0.010505f
C284 B.n244 VSUBS 0.010505f
C285 B.n245 VSUBS 0.010505f
C286 B.n246 VSUBS 0.010505f
C287 B.n247 VSUBS 0.010505f
C288 B.n248 VSUBS 0.010505f
C289 B.n249 VSUBS 0.010505f
C290 B.n250 VSUBS 0.010505f
C291 B.n251 VSUBS 0.010505f
C292 B.n252 VSUBS 0.010505f
C293 B.n253 VSUBS 0.010505f
C294 B.n254 VSUBS 0.010505f
C295 B.n255 VSUBS 0.010505f
C296 B.n256 VSUBS 0.010505f
C297 B.n257 VSUBS 0.010505f
C298 B.n258 VSUBS 0.010505f
C299 B.n259 VSUBS 0.010505f
C300 B.n260 VSUBS 0.010505f
C301 B.n261 VSUBS 0.010505f
C302 B.n262 VSUBS 0.010505f
C303 B.n263 VSUBS 0.010505f
C304 B.n264 VSUBS 0.010505f
C305 B.n265 VSUBS 0.010505f
C306 B.n266 VSUBS 0.010505f
C307 B.n267 VSUBS 0.010505f
C308 B.n268 VSUBS 0.010505f
C309 B.n269 VSUBS 0.010505f
C310 B.n270 VSUBS 0.023361f
C311 B.n271 VSUBS 0.023361f
C312 B.n272 VSUBS 0.024527f
C313 B.n273 VSUBS 0.010505f
C314 B.n274 VSUBS 0.010505f
C315 B.n275 VSUBS 0.010505f
C316 B.n276 VSUBS 0.010505f
C317 B.n277 VSUBS 0.010505f
C318 B.n278 VSUBS 0.010505f
C319 B.n279 VSUBS 0.010505f
C320 B.n280 VSUBS 0.010505f
C321 B.n281 VSUBS 0.010505f
C322 B.n282 VSUBS 0.010505f
C323 B.n283 VSUBS 0.010505f
C324 B.n284 VSUBS 0.010505f
C325 B.n285 VSUBS 0.010505f
C326 B.n286 VSUBS 0.010505f
C327 B.n287 VSUBS 0.010505f
C328 B.n288 VSUBS 0.010505f
C329 B.n289 VSUBS 0.010505f
C330 B.n290 VSUBS 0.007261f
C331 B.n291 VSUBS 0.024338f
C332 B.n292 VSUBS 0.008496f
C333 B.n293 VSUBS 0.010505f
C334 B.n294 VSUBS 0.010505f
C335 B.n295 VSUBS 0.010505f
C336 B.n296 VSUBS 0.010505f
C337 B.n297 VSUBS 0.010505f
C338 B.n298 VSUBS 0.010505f
C339 B.n299 VSUBS 0.010505f
C340 B.n300 VSUBS 0.010505f
C341 B.n301 VSUBS 0.010505f
C342 B.n302 VSUBS 0.010505f
C343 B.n303 VSUBS 0.010505f
C344 B.n304 VSUBS 0.008496f
C345 B.n305 VSUBS 0.010505f
C346 B.n306 VSUBS 0.010505f
C347 B.n307 VSUBS 0.007261f
C348 B.n308 VSUBS 0.010505f
C349 B.n309 VSUBS 0.010505f
C350 B.n310 VSUBS 0.010505f
C351 B.n311 VSUBS 0.010505f
C352 B.n312 VSUBS 0.010505f
C353 B.n313 VSUBS 0.010505f
C354 B.n314 VSUBS 0.010505f
C355 B.n315 VSUBS 0.010505f
C356 B.n316 VSUBS 0.010505f
C357 B.n317 VSUBS 0.010505f
C358 B.n318 VSUBS 0.010505f
C359 B.n319 VSUBS 0.010505f
C360 B.n320 VSUBS 0.010505f
C361 B.n321 VSUBS 0.010505f
C362 B.n322 VSUBS 0.010505f
C363 B.n323 VSUBS 0.010505f
C364 B.n324 VSUBS 0.024527f
C365 B.n325 VSUBS 0.024527f
C366 B.n326 VSUBS 0.023361f
C367 B.n327 VSUBS 0.010505f
C368 B.n328 VSUBS 0.010505f
C369 B.n329 VSUBS 0.010505f
C370 B.n330 VSUBS 0.010505f
C371 B.n331 VSUBS 0.010505f
C372 B.n332 VSUBS 0.010505f
C373 B.n333 VSUBS 0.010505f
C374 B.n334 VSUBS 0.010505f
C375 B.n335 VSUBS 0.010505f
C376 B.n336 VSUBS 0.010505f
C377 B.n337 VSUBS 0.010505f
C378 B.n338 VSUBS 0.010505f
C379 B.n339 VSUBS 0.010505f
C380 B.n340 VSUBS 0.010505f
C381 B.n341 VSUBS 0.010505f
C382 B.n342 VSUBS 0.010505f
C383 B.n343 VSUBS 0.010505f
C384 B.n344 VSUBS 0.010505f
C385 B.n345 VSUBS 0.010505f
C386 B.n346 VSUBS 0.010505f
C387 B.n347 VSUBS 0.010505f
C388 B.n348 VSUBS 0.010505f
C389 B.n349 VSUBS 0.010505f
C390 B.n350 VSUBS 0.010505f
C391 B.n351 VSUBS 0.010505f
C392 B.n352 VSUBS 0.010505f
C393 B.n353 VSUBS 0.010505f
C394 B.n354 VSUBS 0.010505f
C395 B.n355 VSUBS 0.010505f
C396 B.n356 VSUBS 0.010505f
C397 B.n357 VSUBS 0.010505f
C398 B.n358 VSUBS 0.010505f
C399 B.n359 VSUBS 0.010505f
C400 B.n360 VSUBS 0.010505f
C401 B.n361 VSUBS 0.010505f
C402 B.n362 VSUBS 0.010505f
C403 B.n363 VSUBS 0.010505f
C404 B.n364 VSUBS 0.010505f
C405 B.n365 VSUBS 0.010505f
C406 B.n366 VSUBS 0.010505f
C407 B.n367 VSUBS 0.010505f
C408 B.n368 VSUBS 0.010505f
C409 B.n369 VSUBS 0.010505f
C410 B.n370 VSUBS 0.010505f
C411 B.n371 VSUBS 0.010505f
C412 B.n372 VSUBS 0.010505f
C413 B.n373 VSUBS 0.010505f
C414 B.n374 VSUBS 0.010505f
C415 B.n375 VSUBS 0.010505f
C416 B.n376 VSUBS 0.010505f
C417 B.n377 VSUBS 0.010505f
C418 B.n378 VSUBS 0.010505f
C419 B.n379 VSUBS 0.010505f
C420 B.n380 VSUBS 0.010505f
C421 B.n381 VSUBS 0.010505f
C422 B.n382 VSUBS 0.010505f
C423 B.n383 VSUBS 0.010505f
C424 B.n384 VSUBS 0.010505f
C425 B.n385 VSUBS 0.010505f
C426 B.n386 VSUBS 0.010505f
C427 B.n387 VSUBS 0.010505f
C428 B.n388 VSUBS 0.010505f
C429 B.n389 VSUBS 0.010505f
C430 B.n390 VSUBS 0.010505f
C431 B.n391 VSUBS 0.010505f
C432 B.n392 VSUBS 0.010505f
C433 B.n393 VSUBS 0.010505f
C434 B.n394 VSUBS 0.010505f
C435 B.n395 VSUBS 0.010505f
C436 B.n396 VSUBS 0.010505f
C437 B.n397 VSUBS 0.010505f
C438 B.n398 VSUBS 0.010505f
C439 B.n399 VSUBS 0.010505f
C440 B.n400 VSUBS 0.010505f
C441 B.n401 VSUBS 0.010505f
C442 B.n402 VSUBS 0.010505f
C443 B.n403 VSUBS 0.010505f
C444 B.n404 VSUBS 0.010505f
C445 B.n405 VSUBS 0.010505f
C446 B.n406 VSUBS 0.010505f
C447 B.n407 VSUBS 0.010505f
C448 B.n408 VSUBS 0.010505f
C449 B.n409 VSUBS 0.010505f
C450 B.n410 VSUBS 0.010505f
C451 B.n411 VSUBS 0.010505f
C452 B.n412 VSUBS 0.010505f
C453 B.n413 VSUBS 0.010505f
C454 B.n414 VSUBS 0.010505f
C455 B.n415 VSUBS 0.010505f
C456 B.n416 VSUBS 0.010505f
C457 B.n417 VSUBS 0.010505f
C458 B.n418 VSUBS 0.010505f
C459 B.n419 VSUBS 0.010505f
C460 B.n420 VSUBS 0.010505f
C461 B.n421 VSUBS 0.010505f
C462 B.n422 VSUBS 0.010505f
C463 B.n423 VSUBS 0.010505f
C464 B.n424 VSUBS 0.010505f
C465 B.n425 VSUBS 0.010505f
C466 B.n426 VSUBS 0.010505f
C467 B.n427 VSUBS 0.010505f
C468 B.n428 VSUBS 0.010505f
C469 B.n429 VSUBS 0.010505f
C470 B.n430 VSUBS 0.010505f
C471 B.n431 VSUBS 0.010505f
C472 B.n432 VSUBS 0.010505f
C473 B.n433 VSUBS 0.010505f
C474 B.n434 VSUBS 0.010505f
C475 B.n435 VSUBS 0.010505f
C476 B.n436 VSUBS 0.010505f
C477 B.n437 VSUBS 0.010505f
C478 B.n438 VSUBS 0.010505f
C479 B.n439 VSUBS 0.010505f
C480 B.n440 VSUBS 0.010505f
C481 B.n441 VSUBS 0.010505f
C482 B.n442 VSUBS 0.010505f
C483 B.n443 VSUBS 0.010505f
C484 B.n444 VSUBS 0.010505f
C485 B.n445 VSUBS 0.010505f
C486 B.n446 VSUBS 0.010505f
C487 B.n447 VSUBS 0.010505f
C488 B.n448 VSUBS 0.010505f
C489 B.n449 VSUBS 0.010505f
C490 B.n450 VSUBS 0.010505f
C491 B.n451 VSUBS 0.010505f
C492 B.n452 VSUBS 0.010505f
C493 B.n453 VSUBS 0.010505f
C494 B.n454 VSUBS 0.010505f
C495 B.n455 VSUBS 0.010505f
C496 B.n456 VSUBS 0.010505f
C497 B.n457 VSUBS 0.010505f
C498 B.n458 VSUBS 0.010505f
C499 B.n459 VSUBS 0.010505f
C500 B.n460 VSUBS 0.010505f
C501 B.n461 VSUBS 0.010505f
C502 B.n462 VSUBS 0.010505f
C503 B.n463 VSUBS 0.010505f
C504 B.n464 VSUBS 0.010505f
C505 B.n465 VSUBS 0.010505f
C506 B.n466 VSUBS 0.010505f
C507 B.n467 VSUBS 0.010505f
C508 B.n468 VSUBS 0.010505f
C509 B.n469 VSUBS 0.010505f
C510 B.n470 VSUBS 0.010505f
C511 B.n471 VSUBS 0.010505f
C512 B.n472 VSUBS 0.010505f
C513 B.n473 VSUBS 0.010505f
C514 B.n474 VSUBS 0.010505f
C515 B.n475 VSUBS 0.010505f
C516 B.n476 VSUBS 0.010505f
C517 B.n477 VSUBS 0.010505f
C518 B.n478 VSUBS 0.010505f
C519 B.n479 VSUBS 0.010505f
C520 B.n480 VSUBS 0.010505f
C521 B.n481 VSUBS 0.010505f
C522 B.n482 VSUBS 0.010505f
C523 B.n483 VSUBS 0.010505f
C524 B.n484 VSUBS 0.010505f
C525 B.n485 VSUBS 0.010505f
C526 B.n486 VSUBS 0.010505f
C527 B.n487 VSUBS 0.010505f
C528 B.n488 VSUBS 0.010505f
C529 B.n489 VSUBS 0.010505f
C530 B.n490 VSUBS 0.010505f
C531 B.n491 VSUBS 0.010505f
C532 B.n492 VSUBS 0.010505f
C533 B.n493 VSUBS 0.010505f
C534 B.n494 VSUBS 0.010505f
C535 B.n495 VSUBS 0.010505f
C536 B.n496 VSUBS 0.010505f
C537 B.n497 VSUBS 0.010505f
C538 B.n498 VSUBS 0.010505f
C539 B.n499 VSUBS 0.010505f
C540 B.n500 VSUBS 0.010505f
C541 B.n501 VSUBS 0.010505f
C542 B.n502 VSUBS 0.010505f
C543 B.n503 VSUBS 0.010505f
C544 B.n504 VSUBS 0.010505f
C545 B.n505 VSUBS 0.010505f
C546 B.n506 VSUBS 0.010505f
C547 B.n507 VSUBS 0.010505f
C548 B.n508 VSUBS 0.010505f
C549 B.n509 VSUBS 0.010505f
C550 B.n510 VSUBS 0.010505f
C551 B.n511 VSUBS 0.010505f
C552 B.n512 VSUBS 0.010505f
C553 B.n513 VSUBS 0.010505f
C554 B.n514 VSUBS 0.010505f
C555 B.n515 VSUBS 0.010505f
C556 B.n516 VSUBS 0.010505f
C557 B.n517 VSUBS 0.010505f
C558 B.n518 VSUBS 0.010505f
C559 B.n519 VSUBS 0.010505f
C560 B.n520 VSUBS 0.010505f
C561 B.n521 VSUBS 0.023361f
C562 B.n522 VSUBS 0.024527f
C563 B.n523 VSUBS 0.023235f
C564 B.n524 VSUBS 0.010505f
C565 B.n525 VSUBS 0.010505f
C566 B.n526 VSUBS 0.010505f
C567 B.n527 VSUBS 0.010505f
C568 B.n528 VSUBS 0.010505f
C569 B.n529 VSUBS 0.010505f
C570 B.n530 VSUBS 0.010505f
C571 B.n531 VSUBS 0.010505f
C572 B.n532 VSUBS 0.010505f
C573 B.n533 VSUBS 0.010505f
C574 B.n534 VSUBS 0.010505f
C575 B.n535 VSUBS 0.010505f
C576 B.n536 VSUBS 0.010505f
C577 B.n537 VSUBS 0.010505f
C578 B.n538 VSUBS 0.010505f
C579 B.n539 VSUBS 0.010505f
C580 B.n540 VSUBS 0.010505f
C581 B.n541 VSUBS 0.007261f
C582 B.n542 VSUBS 0.024338f
C583 B.n543 VSUBS 0.008496f
C584 B.n544 VSUBS 0.010505f
C585 B.n545 VSUBS 0.010505f
C586 B.n546 VSUBS 0.010505f
C587 B.n547 VSUBS 0.010505f
C588 B.n548 VSUBS 0.010505f
C589 B.n549 VSUBS 0.010505f
C590 B.n550 VSUBS 0.010505f
C591 B.n551 VSUBS 0.010505f
C592 B.n552 VSUBS 0.010505f
C593 B.n553 VSUBS 0.010505f
C594 B.n554 VSUBS 0.010505f
C595 B.n555 VSUBS 0.008496f
C596 B.n556 VSUBS 0.024338f
C597 B.n557 VSUBS 0.007261f
C598 B.n558 VSUBS 0.010505f
C599 B.n559 VSUBS 0.010505f
C600 B.n560 VSUBS 0.010505f
C601 B.n561 VSUBS 0.010505f
C602 B.n562 VSUBS 0.010505f
C603 B.n563 VSUBS 0.010505f
C604 B.n564 VSUBS 0.010505f
C605 B.n565 VSUBS 0.010505f
C606 B.n566 VSUBS 0.010505f
C607 B.n567 VSUBS 0.010505f
C608 B.n568 VSUBS 0.010505f
C609 B.n569 VSUBS 0.010505f
C610 B.n570 VSUBS 0.010505f
C611 B.n571 VSUBS 0.010505f
C612 B.n572 VSUBS 0.010505f
C613 B.n573 VSUBS 0.010505f
C614 B.n574 VSUBS 0.010505f
C615 B.n575 VSUBS 0.024527f
C616 B.n576 VSUBS 0.024527f
C617 B.n577 VSUBS 0.023361f
C618 B.n578 VSUBS 0.010505f
C619 B.n579 VSUBS 0.010505f
C620 B.n580 VSUBS 0.010505f
C621 B.n581 VSUBS 0.010505f
C622 B.n582 VSUBS 0.010505f
C623 B.n583 VSUBS 0.010505f
C624 B.n584 VSUBS 0.010505f
C625 B.n585 VSUBS 0.010505f
C626 B.n586 VSUBS 0.010505f
C627 B.n587 VSUBS 0.010505f
C628 B.n588 VSUBS 0.010505f
C629 B.n589 VSUBS 0.010505f
C630 B.n590 VSUBS 0.010505f
C631 B.n591 VSUBS 0.010505f
C632 B.n592 VSUBS 0.010505f
C633 B.n593 VSUBS 0.010505f
C634 B.n594 VSUBS 0.010505f
C635 B.n595 VSUBS 0.010505f
C636 B.n596 VSUBS 0.010505f
C637 B.n597 VSUBS 0.010505f
C638 B.n598 VSUBS 0.010505f
C639 B.n599 VSUBS 0.010505f
C640 B.n600 VSUBS 0.010505f
C641 B.n601 VSUBS 0.010505f
C642 B.n602 VSUBS 0.010505f
C643 B.n603 VSUBS 0.010505f
C644 B.n604 VSUBS 0.010505f
C645 B.n605 VSUBS 0.010505f
C646 B.n606 VSUBS 0.010505f
C647 B.n607 VSUBS 0.010505f
C648 B.n608 VSUBS 0.010505f
C649 B.n609 VSUBS 0.010505f
C650 B.n610 VSUBS 0.010505f
C651 B.n611 VSUBS 0.010505f
C652 B.n612 VSUBS 0.010505f
C653 B.n613 VSUBS 0.010505f
C654 B.n614 VSUBS 0.010505f
C655 B.n615 VSUBS 0.010505f
C656 B.n616 VSUBS 0.010505f
C657 B.n617 VSUBS 0.010505f
C658 B.n618 VSUBS 0.010505f
C659 B.n619 VSUBS 0.010505f
C660 B.n620 VSUBS 0.010505f
C661 B.n621 VSUBS 0.010505f
C662 B.n622 VSUBS 0.010505f
C663 B.n623 VSUBS 0.010505f
C664 B.n624 VSUBS 0.010505f
C665 B.n625 VSUBS 0.010505f
C666 B.n626 VSUBS 0.010505f
C667 B.n627 VSUBS 0.010505f
C668 B.n628 VSUBS 0.010505f
C669 B.n629 VSUBS 0.010505f
C670 B.n630 VSUBS 0.010505f
C671 B.n631 VSUBS 0.010505f
C672 B.n632 VSUBS 0.010505f
C673 B.n633 VSUBS 0.010505f
C674 B.n634 VSUBS 0.010505f
C675 B.n635 VSUBS 0.010505f
C676 B.n636 VSUBS 0.010505f
C677 B.n637 VSUBS 0.010505f
C678 B.n638 VSUBS 0.010505f
C679 B.n639 VSUBS 0.010505f
C680 B.n640 VSUBS 0.010505f
C681 B.n641 VSUBS 0.010505f
C682 B.n642 VSUBS 0.010505f
C683 B.n643 VSUBS 0.010505f
C684 B.n644 VSUBS 0.010505f
C685 B.n645 VSUBS 0.010505f
C686 B.n646 VSUBS 0.010505f
C687 B.n647 VSUBS 0.010505f
C688 B.n648 VSUBS 0.010505f
C689 B.n649 VSUBS 0.010505f
C690 B.n650 VSUBS 0.010505f
C691 B.n651 VSUBS 0.010505f
C692 B.n652 VSUBS 0.010505f
C693 B.n653 VSUBS 0.010505f
C694 B.n654 VSUBS 0.010505f
C695 B.n655 VSUBS 0.010505f
C696 B.n656 VSUBS 0.010505f
C697 B.n657 VSUBS 0.010505f
C698 B.n658 VSUBS 0.010505f
C699 B.n659 VSUBS 0.010505f
C700 B.n660 VSUBS 0.010505f
C701 B.n661 VSUBS 0.010505f
C702 B.n662 VSUBS 0.010505f
C703 B.n663 VSUBS 0.010505f
C704 B.n664 VSUBS 0.010505f
C705 B.n665 VSUBS 0.010505f
C706 B.n666 VSUBS 0.010505f
C707 B.n667 VSUBS 0.010505f
C708 B.n668 VSUBS 0.010505f
C709 B.n669 VSUBS 0.010505f
C710 B.n670 VSUBS 0.010505f
C711 B.n671 VSUBS 0.010505f
C712 B.n672 VSUBS 0.010505f
C713 B.n673 VSUBS 0.010505f
C714 B.n674 VSUBS 0.010505f
C715 B.n675 VSUBS 0.023786f
C716 VDD1.t2 VSUBS 0.435949f
C717 VDD1.t6 VSUBS 0.062414f
C718 VDD1.t7 VSUBS 0.062414f
C719 VDD1.n0 VSUBS 0.285961f
C720 VDD1.n1 VSUBS 1.5796f
C721 VDD1.t3 VSUBS 0.435948f
C722 VDD1.t5 VSUBS 0.062414f
C723 VDD1.t1 VSUBS 0.062414f
C724 VDD1.n2 VSUBS 0.28596f
C725 VDD1.n3 VSUBS 1.56756f
C726 VDD1.t4 VSUBS 0.062414f
C727 VDD1.t9 VSUBS 0.062414f
C728 VDD1.n4 VSUBS 0.297319f
C729 VDD1.n5 VSUBS 3.89879f
C730 VDD1.t8 VSUBS 0.062414f
C731 VDD1.t0 VSUBS 0.062414f
C732 VDD1.n6 VSUBS 0.28596f
C733 VDD1.n7 VSUBS 3.80059f
C734 VP.t0 VSUBS 0.841278f
C735 VP.n0 VSUBS 0.605584f
C736 VP.n1 VSUBS 0.056865f
C737 VP.n2 VSUBS 0.095248f
C738 VP.n3 VSUBS 0.056865f
C739 VP.t5 VSUBS 0.841278f
C740 VP.n4 VSUBS 0.10545f
C741 VP.n5 VSUBS 0.056865f
C742 VP.n6 VSUBS 0.10545f
C743 VP.n7 VSUBS 0.056865f
C744 VP.t8 VSUBS 0.841278f
C745 VP.n8 VSUBS 0.055349f
C746 VP.n9 VSUBS 0.056865f
C747 VP.t4 VSUBS 0.841278f
C748 VP.n10 VSUBS 0.383657f
C749 VP.n11 VSUBS 0.056865f
C750 VP.n12 VSUBS 0.070075f
C751 VP.n13 VSUBS 0.091764f
C752 VP.t6 VSUBS 0.841278f
C753 VP.t9 VSUBS 0.841278f
C754 VP.n14 VSUBS 0.605584f
C755 VP.n15 VSUBS 0.056865f
C756 VP.n16 VSUBS 0.095248f
C757 VP.n17 VSUBS 0.056865f
C758 VP.t1 VSUBS 0.841278f
C759 VP.n18 VSUBS 0.10545f
C760 VP.n19 VSUBS 0.056865f
C761 VP.n20 VSUBS 0.10545f
C762 VP.n21 VSUBS 0.056865f
C763 VP.t2 VSUBS 0.841278f
C764 VP.n22 VSUBS 0.055349f
C765 VP.n23 VSUBS 0.056865f
C766 VP.t3 VSUBS 0.841278f
C767 VP.n24 VSUBS 0.556727f
C768 VP.t7 VSUBS 1.32416f
C769 VP.n25 VSUBS 0.556343f
C770 VP.n26 VSUBS 0.606097f
C771 VP.n27 VSUBS 0.076298f
C772 VP.n28 VSUBS 0.10545f
C773 VP.n29 VSUBS 0.102743f
C774 VP.n30 VSUBS 0.056865f
C775 VP.n31 VSUBS 0.056865f
C776 VP.n32 VSUBS 0.056865f
C777 VP.n33 VSUBS 0.112681f
C778 VP.n34 VSUBS 0.10545f
C779 VP.n35 VSUBS 0.437049f
C780 VP.n36 VSUBS 0.056865f
C781 VP.n37 VSUBS 0.056865f
C782 VP.n38 VSUBS 0.056865f
C783 VP.n39 VSUBS 0.112681f
C784 VP.n40 VSUBS 0.055349f
C785 VP.n41 VSUBS 0.102743f
C786 VP.n42 VSUBS 0.056865f
C787 VP.n43 VSUBS 0.056865f
C788 VP.n44 VSUBS 0.056865f
C789 VP.n45 VSUBS 0.076298f
C790 VP.n46 VSUBS 0.383657f
C791 VP.n47 VSUBS 0.082545f
C792 VP.n48 VSUBS 0.10545f
C793 VP.n49 VSUBS 0.056865f
C794 VP.n50 VSUBS 0.056865f
C795 VP.n51 VSUBS 0.056865f
C796 VP.n52 VSUBS 0.070075f
C797 VP.n53 VSUBS 0.10545f
C798 VP.n54 VSUBS 0.099203f
C799 VP.n55 VSUBS 0.091764f
C800 VP.n56 VSUBS 2.96126f
C801 VP.n57 VSUBS 3.00454f
C802 VP.n58 VSUBS 0.605584f
C803 VP.n59 VSUBS 0.099203f
C804 VP.n60 VSUBS 0.10545f
C805 VP.n61 VSUBS 0.056865f
C806 VP.n62 VSUBS 0.056865f
C807 VP.n63 VSUBS 0.056865f
C808 VP.n64 VSUBS 0.095248f
C809 VP.n65 VSUBS 0.10545f
C810 VP.n66 VSUBS 0.082545f
C811 VP.n67 VSUBS 0.056865f
C812 VP.n68 VSUBS 0.056865f
C813 VP.n69 VSUBS 0.076298f
C814 VP.n70 VSUBS 0.10545f
C815 VP.n71 VSUBS 0.102743f
C816 VP.n72 VSUBS 0.056865f
C817 VP.n73 VSUBS 0.056865f
C818 VP.n74 VSUBS 0.056865f
C819 VP.n75 VSUBS 0.112681f
C820 VP.n76 VSUBS 0.10545f
C821 VP.n77 VSUBS 0.437049f
C822 VP.n78 VSUBS 0.056865f
C823 VP.n79 VSUBS 0.056865f
C824 VP.n80 VSUBS 0.056865f
C825 VP.n81 VSUBS 0.112681f
C826 VP.n82 VSUBS 0.055349f
C827 VP.n83 VSUBS 0.102743f
C828 VP.n84 VSUBS 0.056865f
C829 VP.n85 VSUBS 0.056865f
C830 VP.n86 VSUBS 0.056865f
C831 VP.n87 VSUBS 0.076298f
C832 VP.n88 VSUBS 0.383657f
C833 VP.n89 VSUBS 0.082545f
C834 VP.n90 VSUBS 0.10545f
C835 VP.n91 VSUBS 0.056865f
C836 VP.n92 VSUBS 0.056865f
C837 VP.n93 VSUBS 0.056865f
C838 VP.n94 VSUBS 0.070075f
C839 VP.n95 VSUBS 0.10545f
C840 VP.n96 VSUBS 0.099203f
C841 VP.n97 VSUBS 0.091764f
C842 VP.n98 VSUBS 0.112298f
C843 VDD2.t1 VSUBS 0.430647f
C844 VDD2.t3 VSUBS 0.061654f
C845 VDD2.t0 VSUBS 0.061654f
C846 VDD2.n0 VSUBS 0.282483f
C847 VDD2.n1 VSUBS 1.5485f
C848 VDD2.t4 VSUBS 0.061654f
C849 VDD2.t9 VSUBS 0.061654f
C850 VDD2.n2 VSUBS 0.293704f
C851 VDD2.n3 VSUBS 3.67288f
C852 VDD2.t6 VSUBS 0.419532f
C853 VDD2.n4 VSUBS 3.59503f
C854 VDD2.t8 VSUBS 0.061654f
C855 VDD2.t2 VSUBS 0.061654f
C856 VDD2.n5 VSUBS 0.282484f
C857 VDD2.n6 VSUBS 0.806703f
C858 VDD2.t7 VSUBS 0.061654f
C859 VDD2.t5 VSUBS 0.061654f
C860 VDD2.n7 VSUBS 0.293679f
C861 VTAIL.t13 VSUBS 0.062841f
C862 VTAIL.t16 VSUBS 0.062841f
C863 VTAIL.n0 VSUBS 0.245638f
C864 VTAIL.n1 VSUBS 0.870201f
C865 VTAIL.t19 VSUBS 0.38595f
C866 VTAIL.n2 VSUBS 0.976695f
C867 VTAIL.t7 VSUBS 0.062841f
C868 VTAIL.t4 VSUBS 0.062841f
C869 VTAIL.n3 VSUBS 0.245638f
C870 VTAIL.n4 VSUBS 1.05454f
C871 VTAIL.t8 VSUBS 0.062841f
C872 VTAIL.t5 VSUBS 0.062841f
C873 VTAIL.n5 VSUBS 0.245638f
C874 VTAIL.n6 VSUBS 2.10483f
C875 VTAIL.t11 VSUBS 0.062841f
C876 VTAIL.t14 VSUBS 0.062841f
C877 VTAIL.n7 VSUBS 0.245639f
C878 VTAIL.n8 VSUBS 2.10483f
C879 VTAIL.t15 VSUBS 0.062841f
C880 VTAIL.t10 VSUBS 0.062841f
C881 VTAIL.n9 VSUBS 0.245639f
C882 VTAIL.n10 VSUBS 1.05454f
C883 VTAIL.t18 VSUBS 0.385952f
C884 VTAIL.n11 VSUBS 0.976693f
C885 VTAIL.t6 VSUBS 0.062841f
C886 VTAIL.t3 VSUBS 0.062841f
C887 VTAIL.n12 VSUBS 0.245639f
C888 VTAIL.n13 VSUBS 0.945622f
C889 VTAIL.t1 VSUBS 0.062841f
C890 VTAIL.t0 VSUBS 0.062841f
C891 VTAIL.n14 VSUBS 0.245639f
C892 VTAIL.n15 VSUBS 1.05454f
C893 VTAIL.t2 VSUBS 0.38595f
C894 VTAIL.n16 VSUBS 1.8066f
C895 VTAIL.t17 VSUBS 0.38595f
C896 VTAIL.n17 VSUBS 1.8066f
C897 VTAIL.t12 VSUBS 0.062841f
C898 VTAIL.t9 VSUBS 0.062841f
C899 VTAIL.n18 VSUBS 0.245638f
C900 VTAIL.n19 VSUBS 0.80066f
C901 VN.t0 VSUBS 0.733567f
C902 VN.n0 VSUBS 0.528049f
C903 VN.n1 VSUBS 0.049584f
C904 VN.n2 VSUBS 0.083053f
C905 VN.n3 VSUBS 0.049584f
C906 VN.t5 VSUBS 0.733567f
C907 VN.n4 VSUBS 0.091949f
C908 VN.n5 VSUBS 0.049584f
C909 VN.n6 VSUBS 0.091949f
C910 VN.n7 VSUBS 0.049584f
C911 VN.t9 VSUBS 0.733567f
C912 VN.n8 VSUBS 0.048262f
C913 VN.n9 VSUBS 0.049584f
C914 VN.t6 VSUBS 0.733567f
C915 VN.n10 VSUBS 0.485447f
C916 VN.t8 VSUBS 1.15462f
C917 VN.n11 VSUBS 0.485112f
C918 VN.n12 VSUBS 0.528495f
C919 VN.n13 VSUBS 0.066529f
C920 VN.n14 VSUBS 0.091949f
C921 VN.n15 VSUBS 0.089589f
C922 VN.n16 VSUBS 0.049584f
C923 VN.n17 VSUBS 0.049584f
C924 VN.n18 VSUBS 0.049584f
C925 VN.n19 VSUBS 0.098254f
C926 VN.n20 VSUBS 0.091949f
C927 VN.n21 VSUBS 0.381092f
C928 VN.n22 VSUBS 0.049584f
C929 VN.n23 VSUBS 0.049584f
C930 VN.n24 VSUBS 0.049584f
C931 VN.n25 VSUBS 0.098254f
C932 VN.n26 VSUBS 0.048262f
C933 VN.n27 VSUBS 0.089589f
C934 VN.n28 VSUBS 0.049584f
C935 VN.n29 VSUBS 0.049584f
C936 VN.n30 VSUBS 0.049584f
C937 VN.n31 VSUBS 0.066529f
C938 VN.n32 VSUBS 0.334536f
C939 VN.n33 VSUBS 0.071976f
C940 VN.n34 VSUBS 0.091949f
C941 VN.n35 VSUBS 0.049584f
C942 VN.n36 VSUBS 0.049584f
C943 VN.n37 VSUBS 0.049584f
C944 VN.n38 VSUBS 0.061103f
C945 VN.n39 VSUBS 0.091949f
C946 VN.n40 VSUBS 0.086502f
C947 VN.n41 VSUBS 0.080015f
C948 VN.n42 VSUBS 0.09792f
C949 VN.t3 VSUBS 0.733567f
C950 VN.n43 VSUBS 0.528049f
C951 VN.n44 VSUBS 0.049584f
C952 VN.n45 VSUBS 0.083053f
C953 VN.n46 VSUBS 0.049584f
C954 VN.t1 VSUBS 0.733567f
C955 VN.n47 VSUBS 0.091949f
C956 VN.n48 VSUBS 0.049584f
C957 VN.n49 VSUBS 0.091949f
C958 VN.n50 VSUBS 0.049584f
C959 VN.t7 VSUBS 0.733567f
C960 VN.n51 VSUBS 0.048262f
C961 VN.n52 VSUBS 0.049584f
C962 VN.t2 VSUBS 0.733567f
C963 VN.n53 VSUBS 0.485447f
C964 VN.t4 VSUBS 1.15462f
C965 VN.n54 VSUBS 0.485112f
C966 VN.n55 VSUBS 0.528495f
C967 VN.n56 VSUBS 0.066529f
C968 VN.n57 VSUBS 0.091949f
C969 VN.n58 VSUBS 0.089589f
C970 VN.n59 VSUBS 0.049584f
C971 VN.n60 VSUBS 0.049584f
C972 VN.n61 VSUBS 0.049584f
C973 VN.n62 VSUBS 0.098254f
C974 VN.n63 VSUBS 0.091949f
C975 VN.n64 VSUBS 0.381092f
C976 VN.n65 VSUBS 0.049584f
C977 VN.n66 VSUBS 0.049584f
C978 VN.n67 VSUBS 0.049584f
C979 VN.n68 VSUBS 0.098254f
C980 VN.n69 VSUBS 0.048262f
C981 VN.n70 VSUBS 0.089589f
C982 VN.n71 VSUBS 0.049584f
C983 VN.n72 VSUBS 0.049584f
C984 VN.n73 VSUBS 0.049584f
C985 VN.n74 VSUBS 0.066529f
C986 VN.n75 VSUBS 0.334536f
C987 VN.n76 VSUBS 0.071976f
C988 VN.n77 VSUBS 0.091949f
C989 VN.n78 VSUBS 0.049584f
C990 VN.n79 VSUBS 0.049584f
C991 VN.n80 VSUBS 0.049584f
C992 VN.n81 VSUBS 0.061103f
C993 VN.n82 VSUBS 0.091949f
C994 VN.n83 VSUBS 0.086502f
C995 VN.n84 VSUBS 0.080015f
C996 VN.n85 VSUBS 2.6028f
.ends

