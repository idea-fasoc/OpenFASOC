* NGSPICE file created from diff_pair_sample_1787.ext - technology: sky130A

.subckt diff_pair_sample_1787 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1254_n2516# sky130_fd_pr__pfet_01v8 ad=3.0108 pd=16.22 as=3.0108 ps=16.22 w=7.72 l=0.38
X1 VDD1.t1 VP.t0 VTAIL.t1 w_n1254_n2516# sky130_fd_pr__pfet_01v8 ad=3.0108 pd=16.22 as=3.0108 ps=16.22 w=7.72 l=0.38
X2 B.t11 B.t9 B.t10 w_n1254_n2516# sky130_fd_pr__pfet_01v8 ad=3.0108 pd=16.22 as=0 ps=0 w=7.72 l=0.38
X3 B.t8 B.t6 B.t7 w_n1254_n2516# sky130_fd_pr__pfet_01v8 ad=3.0108 pd=16.22 as=0 ps=0 w=7.72 l=0.38
X4 B.t5 B.t3 B.t4 w_n1254_n2516# sky130_fd_pr__pfet_01v8 ad=3.0108 pd=16.22 as=0 ps=0 w=7.72 l=0.38
X5 B.t2 B.t0 B.t1 w_n1254_n2516# sky130_fd_pr__pfet_01v8 ad=3.0108 pd=16.22 as=0 ps=0 w=7.72 l=0.38
X6 VDD2.t0 VN.t1 VTAIL.t3 w_n1254_n2516# sky130_fd_pr__pfet_01v8 ad=3.0108 pd=16.22 as=3.0108 ps=16.22 w=7.72 l=0.38
X7 VDD1.t0 VP.t1 VTAIL.t0 w_n1254_n2516# sky130_fd_pr__pfet_01v8 ad=3.0108 pd=16.22 as=3.0108 ps=16.22 w=7.72 l=0.38
R0 VN VN.t1 791.479
R1 VN VN.t0 755.606
R2 VTAIL.n2 VTAIL.t1 69.9623
R3 VTAIL.n1 VTAIL.t3 69.9622
R4 VTAIL.n3 VTAIL.t2 69.9621
R5 VTAIL.n0 VTAIL.t0 69.9621
R6 VTAIL.n1 VTAIL.n0 20.2634
R7 VTAIL.n3 VTAIL.n2 19.6514
R8 VTAIL.n2 VTAIL.n1 0.776362
R9 VTAIL VTAIL.n0 0.681535
R10 VTAIL VTAIL.n3 0.0953276
R11 VDD2.n0 VDD2.t1 118.197
R12 VDD2.n0 VDD2.t0 86.6411
R13 VDD2 VDD2.n0 0.211707
R14 VP.n0 VP.t0 791.097
R15 VP.n0 VP.t1 755.556
R16 VP VP.n0 0.0516364
R17 VDD1 VDD1.t0 118.874
R18 VDD1 VDD1.t1 86.8523
R19 B.n75 B.t6 699.823
R20 B.n81 B.t3 699.823
R21 B.n24 B.t0 699.823
R22 B.n31 B.t9 699.823
R23 B.n262 B.n261 585
R24 B.n263 B.n46 585
R25 B.n265 B.n264 585
R26 B.n266 B.n45 585
R27 B.n268 B.n267 585
R28 B.n269 B.n44 585
R29 B.n271 B.n270 585
R30 B.n272 B.n43 585
R31 B.n274 B.n273 585
R32 B.n275 B.n42 585
R33 B.n277 B.n276 585
R34 B.n278 B.n41 585
R35 B.n280 B.n279 585
R36 B.n281 B.n40 585
R37 B.n283 B.n282 585
R38 B.n284 B.n39 585
R39 B.n286 B.n285 585
R40 B.n287 B.n38 585
R41 B.n289 B.n288 585
R42 B.n290 B.n37 585
R43 B.n292 B.n291 585
R44 B.n293 B.n36 585
R45 B.n295 B.n294 585
R46 B.n296 B.n35 585
R47 B.n298 B.n297 585
R48 B.n299 B.n34 585
R49 B.n301 B.n300 585
R50 B.n302 B.n33 585
R51 B.n304 B.n303 585
R52 B.n306 B.n30 585
R53 B.n308 B.n307 585
R54 B.n309 B.n29 585
R55 B.n311 B.n310 585
R56 B.n312 B.n28 585
R57 B.n314 B.n313 585
R58 B.n315 B.n27 585
R59 B.n317 B.n316 585
R60 B.n318 B.n23 585
R61 B.n320 B.n319 585
R62 B.n321 B.n22 585
R63 B.n323 B.n322 585
R64 B.n324 B.n21 585
R65 B.n326 B.n325 585
R66 B.n327 B.n20 585
R67 B.n329 B.n328 585
R68 B.n330 B.n19 585
R69 B.n332 B.n331 585
R70 B.n333 B.n18 585
R71 B.n335 B.n334 585
R72 B.n336 B.n17 585
R73 B.n338 B.n337 585
R74 B.n339 B.n16 585
R75 B.n341 B.n340 585
R76 B.n342 B.n15 585
R77 B.n344 B.n343 585
R78 B.n345 B.n14 585
R79 B.n347 B.n346 585
R80 B.n348 B.n13 585
R81 B.n350 B.n349 585
R82 B.n351 B.n12 585
R83 B.n353 B.n352 585
R84 B.n354 B.n11 585
R85 B.n356 B.n355 585
R86 B.n357 B.n10 585
R87 B.n359 B.n358 585
R88 B.n360 B.n9 585
R89 B.n362 B.n361 585
R90 B.n363 B.n8 585
R91 B.n260 B.n47 585
R92 B.n259 B.n258 585
R93 B.n257 B.n48 585
R94 B.n256 B.n255 585
R95 B.n254 B.n49 585
R96 B.n253 B.n252 585
R97 B.n251 B.n50 585
R98 B.n250 B.n249 585
R99 B.n248 B.n51 585
R100 B.n247 B.n246 585
R101 B.n245 B.n52 585
R102 B.n244 B.n243 585
R103 B.n242 B.n53 585
R104 B.n241 B.n240 585
R105 B.n239 B.n54 585
R106 B.n238 B.n237 585
R107 B.n236 B.n55 585
R108 B.n235 B.n234 585
R109 B.n233 B.n56 585
R110 B.n232 B.n231 585
R111 B.n230 B.n57 585
R112 B.n229 B.n228 585
R113 B.n227 B.n58 585
R114 B.n226 B.n225 585
R115 B.n224 B.n59 585
R116 B.n121 B.n120 585
R117 B.n122 B.n97 585
R118 B.n124 B.n123 585
R119 B.n125 B.n96 585
R120 B.n127 B.n126 585
R121 B.n128 B.n95 585
R122 B.n130 B.n129 585
R123 B.n131 B.n94 585
R124 B.n133 B.n132 585
R125 B.n134 B.n93 585
R126 B.n136 B.n135 585
R127 B.n137 B.n92 585
R128 B.n139 B.n138 585
R129 B.n140 B.n91 585
R130 B.n142 B.n141 585
R131 B.n143 B.n90 585
R132 B.n145 B.n144 585
R133 B.n146 B.n89 585
R134 B.n148 B.n147 585
R135 B.n149 B.n88 585
R136 B.n151 B.n150 585
R137 B.n152 B.n87 585
R138 B.n154 B.n153 585
R139 B.n155 B.n86 585
R140 B.n157 B.n156 585
R141 B.n158 B.n85 585
R142 B.n160 B.n159 585
R143 B.n161 B.n84 585
R144 B.n163 B.n162 585
R145 B.n165 B.n164 585
R146 B.n166 B.n80 585
R147 B.n168 B.n167 585
R148 B.n169 B.n79 585
R149 B.n171 B.n170 585
R150 B.n172 B.n78 585
R151 B.n174 B.n173 585
R152 B.n175 B.n77 585
R153 B.n177 B.n176 585
R154 B.n178 B.n74 585
R155 B.n181 B.n180 585
R156 B.n182 B.n73 585
R157 B.n184 B.n183 585
R158 B.n185 B.n72 585
R159 B.n187 B.n186 585
R160 B.n188 B.n71 585
R161 B.n190 B.n189 585
R162 B.n191 B.n70 585
R163 B.n193 B.n192 585
R164 B.n194 B.n69 585
R165 B.n196 B.n195 585
R166 B.n197 B.n68 585
R167 B.n199 B.n198 585
R168 B.n200 B.n67 585
R169 B.n202 B.n201 585
R170 B.n203 B.n66 585
R171 B.n205 B.n204 585
R172 B.n206 B.n65 585
R173 B.n208 B.n207 585
R174 B.n209 B.n64 585
R175 B.n211 B.n210 585
R176 B.n212 B.n63 585
R177 B.n214 B.n213 585
R178 B.n215 B.n62 585
R179 B.n217 B.n216 585
R180 B.n218 B.n61 585
R181 B.n220 B.n219 585
R182 B.n221 B.n60 585
R183 B.n223 B.n222 585
R184 B.n119 B.n98 585
R185 B.n118 B.n117 585
R186 B.n116 B.n99 585
R187 B.n115 B.n114 585
R188 B.n113 B.n100 585
R189 B.n112 B.n111 585
R190 B.n110 B.n101 585
R191 B.n109 B.n108 585
R192 B.n107 B.n102 585
R193 B.n106 B.n105 585
R194 B.n104 B.n103 585
R195 B.n2 B.n0 585
R196 B.n381 B.n1 585
R197 B.n380 B.n379 585
R198 B.n378 B.n3 585
R199 B.n377 B.n376 585
R200 B.n375 B.n4 585
R201 B.n374 B.n373 585
R202 B.n372 B.n5 585
R203 B.n371 B.n370 585
R204 B.n369 B.n6 585
R205 B.n368 B.n367 585
R206 B.n366 B.n7 585
R207 B.n365 B.n364 585
R208 B.n383 B.n382 585
R209 B.n121 B.n98 526.135
R210 B.n364 B.n363 526.135
R211 B.n224 B.n223 526.135
R212 B.n261 B.n260 526.135
R213 B.n117 B.n98 163.367
R214 B.n117 B.n116 163.367
R215 B.n116 B.n115 163.367
R216 B.n115 B.n100 163.367
R217 B.n111 B.n100 163.367
R218 B.n111 B.n110 163.367
R219 B.n110 B.n109 163.367
R220 B.n109 B.n102 163.367
R221 B.n105 B.n102 163.367
R222 B.n105 B.n104 163.367
R223 B.n104 B.n2 163.367
R224 B.n382 B.n2 163.367
R225 B.n382 B.n381 163.367
R226 B.n381 B.n380 163.367
R227 B.n380 B.n3 163.367
R228 B.n376 B.n3 163.367
R229 B.n376 B.n375 163.367
R230 B.n375 B.n374 163.367
R231 B.n374 B.n5 163.367
R232 B.n370 B.n5 163.367
R233 B.n370 B.n369 163.367
R234 B.n369 B.n368 163.367
R235 B.n368 B.n7 163.367
R236 B.n364 B.n7 163.367
R237 B.n122 B.n121 163.367
R238 B.n123 B.n122 163.367
R239 B.n123 B.n96 163.367
R240 B.n127 B.n96 163.367
R241 B.n128 B.n127 163.367
R242 B.n129 B.n128 163.367
R243 B.n129 B.n94 163.367
R244 B.n133 B.n94 163.367
R245 B.n134 B.n133 163.367
R246 B.n135 B.n134 163.367
R247 B.n135 B.n92 163.367
R248 B.n139 B.n92 163.367
R249 B.n140 B.n139 163.367
R250 B.n141 B.n140 163.367
R251 B.n141 B.n90 163.367
R252 B.n145 B.n90 163.367
R253 B.n146 B.n145 163.367
R254 B.n147 B.n146 163.367
R255 B.n147 B.n88 163.367
R256 B.n151 B.n88 163.367
R257 B.n152 B.n151 163.367
R258 B.n153 B.n152 163.367
R259 B.n153 B.n86 163.367
R260 B.n157 B.n86 163.367
R261 B.n158 B.n157 163.367
R262 B.n159 B.n158 163.367
R263 B.n159 B.n84 163.367
R264 B.n163 B.n84 163.367
R265 B.n164 B.n163 163.367
R266 B.n164 B.n80 163.367
R267 B.n168 B.n80 163.367
R268 B.n169 B.n168 163.367
R269 B.n170 B.n169 163.367
R270 B.n170 B.n78 163.367
R271 B.n174 B.n78 163.367
R272 B.n175 B.n174 163.367
R273 B.n176 B.n175 163.367
R274 B.n176 B.n74 163.367
R275 B.n181 B.n74 163.367
R276 B.n182 B.n181 163.367
R277 B.n183 B.n182 163.367
R278 B.n183 B.n72 163.367
R279 B.n187 B.n72 163.367
R280 B.n188 B.n187 163.367
R281 B.n189 B.n188 163.367
R282 B.n189 B.n70 163.367
R283 B.n193 B.n70 163.367
R284 B.n194 B.n193 163.367
R285 B.n195 B.n194 163.367
R286 B.n195 B.n68 163.367
R287 B.n199 B.n68 163.367
R288 B.n200 B.n199 163.367
R289 B.n201 B.n200 163.367
R290 B.n201 B.n66 163.367
R291 B.n205 B.n66 163.367
R292 B.n206 B.n205 163.367
R293 B.n207 B.n206 163.367
R294 B.n207 B.n64 163.367
R295 B.n211 B.n64 163.367
R296 B.n212 B.n211 163.367
R297 B.n213 B.n212 163.367
R298 B.n213 B.n62 163.367
R299 B.n217 B.n62 163.367
R300 B.n218 B.n217 163.367
R301 B.n219 B.n218 163.367
R302 B.n219 B.n60 163.367
R303 B.n223 B.n60 163.367
R304 B.n225 B.n224 163.367
R305 B.n225 B.n58 163.367
R306 B.n229 B.n58 163.367
R307 B.n230 B.n229 163.367
R308 B.n231 B.n230 163.367
R309 B.n231 B.n56 163.367
R310 B.n235 B.n56 163.367
R311 B.n236 B.n235 163.367
R312 B.n237 B.n236 163.367
R313 B.n237 B.n54 163.367
R314 B.n241 B.n54 163.367
R315 B.n242 B.n241 163.367
R316 B.n243 B.n242 163.367
R317 B.n243 B.n52 163.367
R318 B.n247 B.n52 163.367
R319 B.n248 B.n247 163.367
R320 B.n249 B.n248 163.367
R321 B.n249 B.n50 163.367
R322 B.n253 B.n50 163.367
R323 B.n254 B.n253 163.367
R324 B.n255 B.n254 163.367
R325 B.n255 B.n48 163.367
R326 B.n259 B.n48 163.367
R327 B.n260 B.n259 163.367
R328 B.n363 B.n362 163.367
R329 B.n362 B.n9 163.367
R330 B.n358 B.n9 163.367
R331 B.n358 B.n357 163.367
R332 B.n357 B.n356 163.367
R333 B.n356 B.n11 163.367
R334 B.n352 B.n11 163.367
R335 B.n352 B.n351 163.367
R336 B.n351 B.n350 163.367
R337 B.n350 B.n13 163.367
R338 B.n346 B.n13 163.367
R339 B.n346 B.n345 163.367
R340 B.n345 B.n344 163.367
R341 B.n344 B.n15 163.367
R342 B.n340 B.n15 163.367
R343 B.n340 B.n339 163.367
R344 B.n339 B.n338 163.367
R345 B.n338 B.n17 163.367
R346 B.n334 B.n17 163.367
R347 B.n334 B.n333 163.367
R348 B.n333 B.n332 163.367
R349 B.n332 B.n19 163.367
R350 B.n328 B.n19 163.367
R351 B.n328 B.n327 163.367
R352 B.n327 B.n326 163.367
R353 B.n326 B.n21 163.367
R354 B.n322 B.n21 163.367
R355 B.n322 B.n321 163.367
R356 B.n321 B.n320 163.367
R357 B.n320 B.n23 163.367
R358 B.n316 B.n23 163.367
R359 B.n316 B.n315 163.367
R360 B.n315 B.n314 163.367
R361 B.n314 B.n28 163.367
R362 B.n310 B.n28 163.367
R363 B.n310 B.n309 163.367
R364 B.n309 B.n308 163.367
R365 B.n308 B.n30 163.367
R366 B.n303 B.n30 163.367
R367 B.n303 B.n302 163.367
R368 B.n302 B.n301 163.367
R369 B.n301 B.n34 163.367
R370 B.n297 B.n34 163.367
R371 B.n297 B.n296 163.367
R372 B.n296 B.n295 163.367
R373 B.n295 B.n36 163.367
R374 B.n291 B.n36 163.367
R375 B.n291 B.n290 163.367
R376 B.n290 B.n289 163.367
R377 B.n289 B.n38 163.367
R378 B.n285 B.n38 163.367
R379 B.n285 B.n284 163.367
R380 B.n284 B.n283 163.367
R381 B.n283 B.n40 163.367
R382 B.n279 B.n40 163.367
R383 B.n279 B.n278 163.367
R384 B.n278 B.n277 163.367
R385 B.n277 B.n42 163.367
R386 B.n273 B.n42 163.367
R387 B.n273 B.n272 163.367
R388 B.n272 B.n271 163.367
R389 B.n271 B.n44 163.367
R390 B.n267 B.n44 163.367
R391 B.n267 B.n266 163.367
R392 B.n266 B.n265 163.367
R393 B.n265 B.n46 163.367
R394 B.n261 B.n46 163.367
R395 B.n75 B.t8 127.341
R396 B.n31 B.t10 127.341
R397 B.n81 B.t5 127.334
R398 B.n24 B.t1 127.334
R399 B.n76 B.t7 113.573
R400 B.n32 B.t11 113.573
R401 B.n82 B.t4 113.564
R402 B.n25 B.t2 113.564
R403 B.n179 B.n76 59.5399
R404 B.n83 B.n82 59.5399
R405 B.n26 B.n25 59.5399
R406 B.n305 B.n32 59.5399
R407 B.n365 B.n8 34.1859
R408 B.n262 B.n47 34.1859
R409 B.n222 B.n59 34.1859
R410 B.n120 B.n119 34.1859
R411 B B.n383 18.0485
R412 B.n76 B.n75 13.7702
R413 B.n82 B.n81 13.7702
R414 B.n25 B.n24 13.7702
R415 B.n32 B.n31 13.7702
R416 B.n361 B.n8 10.6151
R417 B.n361 B.n360 10.6151
R418 B.n360 B.n359 10.6151
R419 B.n359 B.n10 10.6151
R420 B.n355 B.n10 10.6151
R421 B.n355 B.n354 10.6151
R422 B.n354 B.n353 10.6151
R423 B.n353 B.n12 10.6151
R424 B.n349 B.n12 10.6151
R425 B.n349 B.n348 10.6151
R426 B.n348 B.n347 10.6151
R427 B.n347 B.n14 10.6151
R428 B.n343 B.n14 10.6151
R429 B.n343 B.n342 10.6151
R430 B.n342 B.n341 10.6151
R431 B.n341 B.n16 10.6151
R432 B.n337 B.n16 10.6151
R433 B.n337 B.n336 10.6151
R434 B.n336 B.n335 10.6151
R435 B.n335 B.n18 10.6151
R436 B.n331 B.n18 10.6151
R437 B.n331 B.n330 10.6151
R438 B.n330 B.n329 10.6151
R439 B.n329 B.n20 10.6151
R440 B.n325 B.n20 10.6151
R441 B.n325 B.n324 10.6151
R442 B.n324 B.n323 10.6151
R443 B.n323 B.n22 10.6151
R444 B.n319 B.n318 10.6151
R445 B.n318 B.n317 10.6151
R446 B.n317 B.n27 10.6151
R447 B.n313 B.n27 10.6151
R448 B.n313 B.n312 10.6151
R449 B.n312 B.n311 10.6151
R450 B.n311 B.n29 10.6151
R451 B.n307 B.n29 10.6151
R452 B.n307 B.n306 10.6151
R453 B.n304 B.n33 10.6151
R454 B.n300 B.n33 10.6151
R455 B.n300 B.n299 10.6151
R456 B.n299 B.n298 10.6151
R457 B.n298 B.n35 10.6151
R458 B.n294 B.n35 10.6151
R459 B.n294 B.n293 10.6151
R460 B.n293 B.n292 10.6151
R461 B.n292 B.n37 10.6151
R462 B.n288 B.n37 10.6151
R463 B.n288 B.n287 10.6151
R464 B.n287 B.n286 10.6151
R465 B.n286 B.n39 10.6151
R466 B.n282 B.n39 10.6151
R467 B.n282 B.n281 10.6151
R468 B.n281 B.n280 10.6151
R469 B.n280 B.n41 10.6151
R470 B.n276 B.n41 10.6151
R471 B.n276 B.n275 10.6151
R472 B.n275 B.n274 10.6151
R473 B.n274 B.n43 10.6151
R474 B.n270 B.n43 10.6151
R475 B.n270 B.n269 10.6151
R476 B.n269 B.n268 10.6151
R477 B.n268 B.n45 10.6151
R478 B.n264 B.n45 10.6151
R479 B.n264 B.n263 10.6151
R480 B.n263 B.n262 10.6151
R481 B.n226 B.n59 10.6151
R482 B.n227 B.n226 10.6151
R483 B.n228 B.n227 10.6151
R484 B.n228 B.n57 10.6151
R485 B.n232 B.n57 10.6151
R486 B.n233 B.n232 10.6151
R487 B.n234 B.n233 10.6151
R488 B.n234 B.n55 10.6151
R489 B.n238 B.n55 10.6151
R490 B.n239 B.n238 10.6151
R491 B.n240 B.n239 10.6151
R492 B.n240 B.n53 10.6151
R493 B.n244 B.n53 10.6151
R494 B.n245 B.n244 10.6151
R495 B.n246 B.n245 10.6151
R496 B.n246 B.n51 10.6151
R497 B.n250 B.n51 10.6151
R498 B.n251 B.n250 10.6151
R499 B.n252 B.n251 10.6151
R500 B.n252 B.n49 10.6151
R501 B.n256 B.n49 10.6151
R502 B.n257 B.n256 10.6151
R503 B.n258 B.n257 10.6151
R504 B.n258 B.n47 10.6151
R505 B.n120 B.n97 10.6151
R506 B.n124 B.n97 10.6151
R507 B.n125 B.n124 10.6151
R508 B.n126 B.n125 10.6151
R509 B.n126 B.n95 10.6151
R510 B.n130 B.n95 10.6151
R511 B.n131 B.n130 10.6151
R512 B.n132 B.n131 10.6151
R513 B.n132 B.n93 10.6151
R514 B.n136 B.n93 10.6151
R515 B.n137 B.n136 10.6151
R516 B.n138 B.n137 10.6151
R517 B.n138 B.n91 10.6151
R518 B.n142 B.n91 10.6151
R519 B.n143 B.n142 10.6151
R520 B.n144 B.n143 10.6151
R521 B.n144 B.n89 10.6151
R522 B.n148 B.n89 10.6151
R523 B.n149 B.n148 10.6151
R524 B.n150 B.n149 10.6151
R525 B.n150 B.n87 10.6151
R526 B.n154 B.n87 10.6151
R527 B.n155 B.n154 10.6151
R528 B.n156 B.n155 10.6151
R529 B.n156 B.n85 10.6151
R530 B.n160 B.n85 10.6151
R531 B.n161 B.n160 10.6151
R532 B.n162 B.n161 10.6151
R533 B.n166 B.n165 10.6151
R534 B.n167 B.n166 10.6151
R535 B.n167 B.n79 10.6151
R536 B.n171 B.n79 10.6151
R537 B.n172 B.n171 10.6151
R538 B.n173 B.n172 10.6151
R539 B.n173 B.n77 10.6151
R540 B.n177 B.n77 10.6151
R541 B.n178 B.n177 10.6151
R542 B.n180 B.n73 10.6151
R543 B.n184 B.n73 10.6151
R544 B.n185 B.n184 10.6151
R545 B.n186 B.n185 10.6151
R546 B.n186 B.n71 10.6151
R547 B.n190 B.n71 10.6151
R548 B.n191 B.n190 10.6151
R549 B.n192 B.n191 10.6151
R550 B.n192 B.n69 10.6151
R551 B.n196 B.n69 10.6151
R552 B.n197 B.n196 10.6151
R553 B.n198 B.n197 10.6151
R554 B.n198 B.n67 10.6151
R555 B.n202 B.n67 10.6151
R556 B.n203 B.n202 10.6151
R557 B.n204 B.n203 10.6151
R558 B.n204 B.n65 10.6151
R559 B.n208 B.n65 10.6151
R560 B.n209 B.n208 10.6151
R561 B.n210 B.n209 10.6151
R562 B.n210 B.n63 10.6151
R563 B.n214 B.n63 10.6151
R564 B.n215 B.n214 10.6151
R565 B.n216 B.n215 10.6151
R566 B.n216 B.n61 10.6151
R567 B.n220 B.n61 10.6151
R568 B.n221 B.n220 10.6151
R569 B.n222 B.n221 10.6151
R570 B.n119 B.n118 10.6151
R571 B.n118 B.n99 10.6151
R572 B.n114 B.n99 10.6151
R573 B.n114 B.n113 10.6151
R574 B.n113 B.n112 10.6151
R575 B.n112 B.n101 10.6151
R576 B.n108 B.n101 10.6151
R577 B.n108 B.n107 10.6151
R578 B.n107 B.n106 10.6151
R579 B.n106 B.n103 10.6151
R580 B.n103 B.n0 10.6151
R581 B.n379 B.n1 10.6151
R582 B.n379 B.n378 10.6151
R583 B.n378 B.n377 10.6151
R584 B.n377 B.n4 10.6151
R585 B.n373 B.n4 10.6151
R586 B.n373 B.n372 10.6151
R587 B.n372 B.n371 10.6151
R588 B.n371 B.n6 10.6151
R589 B.n367 B.n6 10.6151
R590 B.n367 B.n366 10.6151
R591 B.n366 B.n365 10.6151
R592 B.n26 B.n22 8.74196
R593 B.n305 B.n304 8.74196
R594 B.n162 B.n83 8.74196
R595 B.n180 B.n179 8.74196
R596 B.n383 B.n0 2.81026
R597 B.n383 B.n1 2.81026
R598 B.n319 B.n26 1.87367
R599 B.n306 B.n305 1.87367
R600 B.n165 B.n83 1.87367
R601 B.n179 B.n178 1.87367
C0 VN VDD2 1.09481f
C1 VP VDD1 1.18417f
C2 VN VTAIL 0.729093f
C3 VDD1 B 1.05202f
C4 VP VDD2 0.240662f
C5 w_n1254_n2516# VDD1 1.21734f
C6 VP VTAIL 0.743597f
C7 VDD2 B 1.06443f
C8 VTAIL B 1.79274f
C9 w_n1254_n2516# VDD2 1.2188f
C10 w_n1254_n2516# VTAIL 2.24983f
C11 VN VP 3.62629f
C12 VN B 0.619572f
C13 VN w_n1254_n2516# 1.47446f
C14 VDD1 VDD2 0.431939f
C15 VTAIL VDD1 4.61166f
C16 VP B 0.865409f
C17 w_n1254_n2516# VP 1.62941f
C18 VTAIL VDD2 4.64484f
C19 w_n1254_n2516# B 5.21358f
C20 VN VDD1 0.14811f
C21 VDD2 VSUBS 0.576698f
C22 VDD1 VSUBS 2.956753f
C23 VTAIL VSUBS 0.224907f
C24 VN VSUBS 4.1239f
C25 VP VSUBS 0.856577f
C26 B VSUBS 1.898609f
C27 w_n1254_n2516# VSUBS 39.169895f
C28 B.n0 VSUBS 0.003961f
C29 B.n1 VSUBS 0.003961f
C30 B.n2 VSUBS 0.006263f
C31 B.n3 VSUBS 0.006263f
C32 B.n4 VSUBS 0.006263f
C33 B.n5 VSUBS 0.006263f
C34 B.n6 VSUBS 0.006263f
C35 B.n7 VSUBS 0.006263f
C36 B.n8 VSUBS 0.015683f
C37 B.n9 VSUBS 0.006263f
C38 B.n10 VSUBS 0.006263f
C39 B.n11 VSUBS 0.006263f
C40 B.n12 VSUBS 0.006263f
C41 B.n13 VSUBS 0.006263f
C42 B.n14 VSUBS 0.006263f
C43 B.n15 VSUBS 0.006263f
C44 B.n16 VSUBS 0.006263f
C45 B.n17 VSUBS 0.006263f
C46 B.n18 VSUBS 0.006263f
C47 B.n19 VSUBS 0.006263f
C48 B.n20 VSUBS 0.006263f
C49 B.n21 VSUBS 0.006263f
C50 B.n22 VSUBS 0.005711f
C51 B.n23 VSUBS 0.006263f
C52 B.t2 VSUBS 0.211814f
C53 B.t1 VSUBS 0.216865f
C54 B.t0 VSUBS 0.106776f
C55 B.n24 VSUBS 0.07685f
C56 B.n25 VSUBS 0.055647f
C57 B.n26 VSUBS 0.014512f
C58 B.n27 VSUBS 0.006263f
C59 B.n28 VSUBS 0.006263f
C60 B.n29 VSUBS 0.006263f
C61 B.n30 VSUBS 0.006263f
C62 B.t11 VSUBS 0.211812f
C63 B.t10 VSUBS 0.216864f
C64 B.t9 VSUBS 0.106776f
C65 B.n31 VSUBS 0.076851f
C66 B.n32 VSUBS 0.055649f
C67 B.n33 VSUBS 0.006263f
C68 B.n34 VSUBS 0.006263f
C69 B.n35 VSUBS 0.006263f
C70 B.n36 VSUBS 0.006263f
C71 B.n37 VSUBS 0.006263f
C72 B.n38 VSUBS 0.006263f
C73 B.n39 VSUBS 0.006263f
C74 B.n40 VSUBS 0.006263f
C75 B.n41 VSUBS 0.006263f
C76 B.n42 VSUBS 0.006263f
C77 B.n43 VSUBS 0.006263f
C78 B.n44 VSUBS 0.006263f
C79 B.n45 VSUBS 0.006263f
C80 B.n46 VSUBS 0.006263f
C81 B.n47 VSUBS 0.015235f
C82 B.n48 VSUBS 0.006263f
C83 B.n49 VSUBS 0.006263f
C84 B.n50 VSUBS 0.006263f
C85 B.n51 VSUBS 0.006263f
C86 B.n52 VSUBS 0.006263f
C87 B.n53 VSUBS 0.006263f
C88 B.n54 VSUBS 0.006263f
C89 B.n55 VSUBS 0.006263f
C90 B.n56 VSUBS 0.006263f
C91 B.n57 VSUBS 0.006263f
C92 B.n58 VSUBS 0.006263f
C93 B.n59 VSUBS 0.014528f
C94 B.n60 VSUBS 0.006263f
C95 B.n61 VSUBS 0.006263f
C96 B.n62 VSUBS 0.006263f
C97 B.n63 VSUBS 0.006263f
C98 B.n64 VSUBS 0.006263f
C99 B.n65 VSUBS 0.006263f
C100 B.n66 VSUBS 0.006263f
C101 B.n67 VSUBS 0.006263f
C102 B.n68 VSUBS 0.006263f
C103 B.n69 VSUBS 0.006263f
C104 B.n70 VSUBS 0.006263f
C105 B.n71 VSUBS 0.006263f
C106 B.n72 VSUBS 0.006263f
C107 B.n73 VSUBS 0.006263f
C108 B.n74 VSUBS 0.006263f
C109 B.t7 VSUBS 0.211812f
C110 B.t8 VSUBS 0.216864f
C111 B.t6 VSUBS 0.106776f
C112 B.n75 VSUBS 0.076851f
C113 B.n76 VSUBS 0.055649f
C114 B.n77 VSUBS 0.006263f
C115 B.n78 VSUBS 0.006263f
C116 B.n79 VSUBS 0.006263f
C117 B.n80 VSUBS 0.006263f
C118 B.t4 VSUBS 0.211814f
C119 B.t5 VSUBS 0.216865f
C120 B.t3 VSUBS 0.106776f
C121 B.n81 VSUBS 0.07685f
C122 B.n82 VSUBS 0.055647f
C123 B.n83 VSUBS 0.014512f
C124 B.n84 VSUBS 0.006263f
C125 B.n85 VSUBS 0.006263f
C126 B.n86 VSUBS 0.006263f
C127 B.n87 VSUBS 0.006263f
C128 B.n88 VSUBS 0.006263f
C129 B.n89 VSUBS 0.006263f
C130 B.n90 VSUBS 0.006263f
C131 B.n91 VSUBS 0.006263f
C132 B.n92 VSUBS 0.006263f
C133 B.n93 VSUBS 0.006263f
C134 B.n94 VSUBS 0.006263f
C135 B.n95 VSUBS 0.006263f
C136 B.n96 VSUBS 0.006263f
C137 B.n97 VSUBS 0.006263f
C138 B.n98 VSUBS 0.014528f
C139 B.n99 VSUBS 0.006263f
C140 B.n100 VSUBS 0.006263f
C141 B.n101 VSUBS 0.006263f
C142 B.n102 VSUBS 0.006263f
C143 B.n103 VSUBS 0.006263f
C144 B.n104 VSUBS 0.006263f
C145 B.n105 VSUBS 0.006263f
C146 B.n106 VSUBS 0.006263f
C147 B.n107 VSUBS 0.006263f
C148 B.n108 VSUBS 0.006263f
C149 B.n109 VSUBS 0.006263f
C150 B.n110 VSUBS 0.006263f
C151 B.n111 VSUBS 0.006263f
C152 B.n112 VSUBS 0.006263f
C153 B.n113 VSUBS 0.006263f
C154 B.n114 VSUBS 0.006263f
C155 B.n115 VSUBS 0.006263f
C156 B.n116 VSUBS 0.006263f
C157 B.n117 VSUBS 0.006263f
C158 B.n118 VSUBS 0.006263f
C159 B.n119 VSUBS 0.014528f
C160 B.n120 VSUBS 0.015683f
C161 B.n121 VSUBS 0.015683f
C162 B.n122 VSUBS 0.006263f
C163 B.n123 VSUBS 0.006263f
C164 B.n124 VSUBS 0.006263f
C165 B.n125 VSUBS 0.006263f
C166 B.n126 VSUBS 0.006263f
C167 B.n127 VSUBS 0.006263f
C168 B.n128 VSUBS 0.006263f
C169 B.n129 VSUBS 0.006263f
C170 B.n130 VSUBS 0.006263f
C171 B.n131 VSUBS 0.006263f
C172 B.n132 VSUBS 0.006263f
C173 B.n133 VSUBS 0.006263f
C174 B.n134 VSUBS 0.006263f
C175 B.n135 VSUBS 0.006263f
C176 B.n136 VSUBS 0.006263f
C177 B.n137 VSUBS 0.006263f
C178 B.n138 VSUBS 0.006263f
C179 B.n139 VSUBS 0.006263f
C180 B.n140 VSUBS 0.006263f
C181 B.n141 VSUBS 0.006263f
C182 B.n142 VSUBS 0.006263f
C183 B.n143 VSUBS 0.006263f
C184 B.n144 VSUBS 0.006263f
C185 B.n145 VSUBS 0.006263f
C186 B.n146 VSUBS 0.006263f
C187 B.n147 VSUBS 0.006263f
C188 B.n148 VSUBS 0.006263f
C189 B.n149 VSUBS 0.006263f
C190 B.n150 VSUBS 0.006263f
C191 B.n151 VSUBS 0.006263f
C192 B.n152 VSUBS 0.006263f
C193 B.n153 VSUBS 0.006263f
C194 B.n154 VSUBS 0.006263f
C195 B.n155 VSUBS 0.006263f
C196 B.n156 VSUBS 0.006263f
C197 B.n157 VSUBS 0.006263f
C198 B.n158 VSUBS 0.006263f
C199 B.n159 VSUBS 0.006263f
C200 B.n160 VSUBS 0.006263f
C201 B.n161 VSUBS 0.006263f
C202 B.n162 VSUBS 0.005711f
C203 B.n163 VSUBS 0.006263f
C204 B.n164 VSUBS 0.006263f
C205 B.n165 VSUBS 0.003684f
C206 B.n166 VSUBS 0.006263f
C207 B.n167 VSUBS 0.006263f
C208 B.n168 VSUBS 0.006263f
C209 B.n169 VSUBS 0.006263f
C210 B.n170 VSUBS 0.006263f
C211 B.n171 VSUBS 0.006263f
C212 B.n172 VSUBS 0.006263f
C213 B.n173 VSUBS 0.006263f
C214 B.n174 VSUBS 0.006263f
C215 B.n175 VSUBS 0.006263f
C216 B.n176 VSUBS 0.006263f
C217 B.n177 VSUBS 0.006263f
C218 B.n178 VSUBS 0.003684f
C219 B.n179 VSUBS 0.014512f
C220 B.n180 VSUBS 0.005711f
C221 B.n181 VSUBS 0.006263f
C222 B.n182 VSUBS 0.006263f
C223 B.n183 VSUBS 0.006263f
C224 B.n184 VSUBS 0.006263f
C225 B.n185 VSUBS 0.006263f
C226 B.n186 VSUBS 0.006263f
C227 B.n187 VSUBS 0.006263f
C228 B.n188 VSUBS 0.006263f
C229 B.n189 VSUBS 0.006263f
C230 B.n190 VSUBS 0.006263f
C231 B.n191 VSUBS 0.006263f
C232 B.n192 VSUBS 0.006263f
C233 B.n193 VSUBS 0.006263f
C234 B.n194 VSUBS 0.006263f
C235 B.n195 VSUBS 0.006263f
C236 B.n196 VSUBS 0.006263f
C237 B.n197 VSUBS 0.006263f
C238 B.n198 VSUBS 0.006263f
C239 B.n199 VSUBS 0.006263f
C240 B.n200 VSUBS 0.006263f
C241 B.n201 VSUBS 0.006263f
C242 B.n202 VSUBS 0.006263f
C243 B.n203 VSUBS 0.006263f
C244 B.n204 VSUBS 0.006263f
C245 B.n205 VSUBS 0.006263f
C246 B.n206 VSUBS 0.006263f
C247 B.n207 VSUBS 0.006263f
C248 B.n208 VSUBS 0.006263f
C249 B.n209 VSUBS 0.006263f
C250 B.n210 VSUBS 0.006263f
C251 B.n211 VSUBS 0.006263f
C252 B.n212 VSUBS 0.006263f
C253 B.n213 VSUBS 0.006263f
C254 B.n214 VSUBS 0.006263f
C255 B.n215 VSUBS 0.006263f
C256 B.n216 VSUBS 0.006263f
C257 B.n217 VSUBS 0.006263f
C258 B.n218 VSUBS 0.006263f
C259 B.n219 VSUBS 0.006263f
C260 B.n220 VSUBS 0.006263f
C261 B.n221 VSUBS 0.006263f
C262 B.n222 VSUBS 0.015683f
C263 B.n223 VSUBS 0.015683f
C264 B.n224 VSUBS 0.014528f
C265 B.n225 VSUBS 0.006263f
C266 B.n226 VSUBS 0.006263f
C267 B.n227 VSUBS 0.006263f
C268 B.n228 VSUBS 0.006263f
C269 B.n229 VSUBS 0.006263f
C270 B.n230 VSUBS 0.006263f
C271 B.n231 VSUBS 0.006263f
C272 B.n232 VSUBS 0.006263f
C273 B.n233 VSUBS 0.006263f
C274 B.n234 VSUBS 0.006263f
C275 B.n235 VSUBS 0.006263f
C276 B.n236 VSUBS 0.006263f
C277 B.n237 VSUBS 0.006263f
C278 B.n238 VSUBS 0.006263f
C279 B.n239 VSUBS 0.006263f
C280 B.n240 VSUBS 0.006263f
C281 B.n241 VSUBS 0.006263f
C282 B.n242 VSUBS 0.006263f
C283 B.n243 VSUBS 0.006263f
C284 B.n244 VSUBS 0.006263f
C285 B.n245 VSUBS 0.006263f
C286 B.n246 VSUBS 0.006263f
C287 B.n247 VSUBS 0.006263f
C288 B.n248 VSUBS 0.006263f
C289 B.n249 VSUBS 0.006263f
C290 B.n250 VSUBS 0.006263f
C291 B.n251 VSUBS 0.006263f
C292 B.n252 VSUBS 0.006263f
C293 B.n253 VSUBS 0.006263f
C294 B.n254 VSUBS 0.006263f
C295 B.n255 VSUBS 0.006263f
C296 B.n256 VSUBS 0.006263f
C297 B.n257 VSUBS 0.006263f
C298 B.n258 VSUBS 0.006263f
C299 B.n259 VSUBS 0.006263f
C300 B.n260 VSUBS 0.014528f
C301 B.n261 VSUBS 0.015683f
C302 B.n262 VSUBS 0.014976f
C303 B.n263 VSUBS 0.006263f
C304 B.n264 VSUBS 0.006263f
C305 B.n265 VSUBS 0.006263f
C306 B.n266 VSUBS 0.006263f
C307 B.n267 VSUBS 0.006263f
C308 B.n268 VSUBS 0.006263f
C309 B.n269 VSUBS 0.006263f
C310 B.n270 VSUBS 0.006263f
C311 B.n271 VSUBS 0.006263f
C312 B.n272 VSUBS 0.006263f
C313 B.n273 VSUBS 0.006263f
C314 B.n274 VSUBS 0.006263f
C315 B.n275 VSUBS 0.006263f
C316 B.n276 VSUBS 0.006263f
C317 B.n277 VSUBS 0.006263f
C318 B.n278 VSUBS 0.006263f
C319 B.n279 VSUBS 0.006263f
C320 B.n280 VSUBS 0.006263f
C321 B.n281 VSUBS 0.006263f
C322 B.n282 VSUBS 0.006263f
C323 B.n283 VSUBS 0.006263f
C324 B.n284 VSUBS 0.006263f
C325 B.n285 VSUBS 0.006263f
C326 B.n286 VSUBS 0.006263f
C327 B.n287 VSUBS 0.006263f
C328 B.n288 VSUBS 0.006263f
C329 B.n289 VSUBS 0.006263f
C330 B.n290 VSUBS 0.006263f
C331 B.n291 VSUBS 0.006263f
C332 B.n292 VSUBS 0.006263f
C333 B.n293 VSUBS 0.006263f
C334 B.n294 VSUBS 0.006263f
C335 B.n295 VSUBS 0.006263f
C336 B.n296 VSUBS 0.006263f
C337 B.n297 VSUBS 0.006263f
C338 B.n298 VSUBS 0.006263f
C339 B.n299 VSUBS 0.006263f
C340 B.n300 VSUBS 0.006263f
C341 B.n301 VSUBS 0.006263f
C342 B.n302 VSUBS 0.006263f
C343 B.n303 VSUBS 0.006263f
C344 B.n304 VSUBS 0.005711f
C345 B.n305 VSUBS 0.014512f
C346 B.n306 VSUBS 0.003684f
C347 B.n307 VSUBS 0.006263f
C348 B.n308 VSUBS 0.006263f
C349 B.n309 VSUBS 0.006263f
C350 B.n310 VSUBS 0.006263f
C351 B.n311 VSUBS 0.006263f
C352 B.n312 VSUBS 0.006263f
C353 B.n313 VSUBS 0.006263f
C354 B.n314 VSUBS 0.006263f
C355 B.n315 VSUBS 0.006263f
C356 B.n316 VSUBS 0.006263f
C357 B.n317 VSUBS 0.006263f
C358 B.n318 VSUBS 0.006263f
C359 B.n319 VSUBS 0.003684f
C360 B.n320 VSUBS 0.006263f
C361 B.n321 VSUBS 0.006263f
C362 B.n322 VSUBS 0.006263f
C363 B.n323 VSUBS 0.006263f
C364 B.n324 VSUBS 0.006263f
C365 B.n325 VSUBS 0.006263f
C366 B.n326 VSUBS 0.006263f
C367 B.n327 VSUBS 0.006263f
C368 B.n328 VSUBS 0.006263f
C369 B.n329 VSUBS 0.006263f
C370 B.n330 VSUBS 0.006263f
C371 B.n331 VSUBS 0.006263f
C372 B.n332 VSUBS 0.006263f
C373 B.n333 VSUBS 0.006263f
C374 B.n334 VSUBS 0.006263f
C375 B.n335 VSUBS 0.006263f
C376 B.n336 VSUBS 0.006263f
C377 B.n337 VSUBS 0.006263f
C378 B.n338 VSUBS 0.006263f
C379 B.n339 VSUBS 0.006263f
C380 B.n340 VSUBS 0.006263f
C381 B.n341 VSUBS 0.006263f
C382 B.n342 VSUBS 0.006263f
C383 B.n343 VSUBS 0.006263f
C384 B.n344 VSUBS 0.006263f
C385 B.n345 VSUBS 0.006263f
C386 B.n346 VSUBS 0.006263f
C387 B.n347 VSUBS 0.006263f
C388 B.n348 VSUBS 0.006263f
C389 B.n349 VSUBS 0.006263f
C390 B.n350 VSUBS 0.006263f
C391 B.n351 VSUBS 0.006263f
C392 B.n352 VSUBS 0.006263f
C393 B.n353 VSUBS 0.006263f
C394 B.n354 VSUBS 0.006263f
C395 B.n355 VSUBS 0.006263f
C396 B.n356 VSUBS 0.006263f
C397 B.n357 VSUBS 0.006263f
C398 B.n358 VSUBS 0.006263f
C399 B.n359 VSUBS 0.006263f
C400 B.n360 VSUBS 0.006263f
C401 B.n361 VSUBS 0.006263f
C402 B.n362 VSUBS 0.006263f
C403 B.n363 VSUBS 0.015683f
C404 B.n364 VSUBS 0.014528f
C405 B.n365 VSUBS 0.014528f
C406 B.n366 VSUBS 0.006263f
C407 B.n367 VSUBS 0.006263f
C408 B.n368 VSUBS 0.006263f
C409 B.n369 VSUBS 0.006263f
C410 B.n370 VSUBS 0.006263f
C411 B.n371 VSUBS 0.006263f
C412 B.n372 VSUBS 0.006263f
C413 B.n373 VSUBS 0.006263f
C414 B.n374 VSUBS 0.006263f
C415 B.n375 VSUBS 0.006263f
C416 B.n376 VSUBS 0.006263f
C417 B.n377 VSUBS 0.006263f
C418 B.n378 VSUBS 0.006263f
C419 B.n379 VSUBS 0.006263f
C420 B.n380 VSUBS 0.006263f
C421 B.n381 VSUBS 0.006263f
C422 B.n382 VSUBS 0.006263f
C423 B.n383 VSUBS 0.014182f
C424 VDD1.t1 VSUBS 1.01276f
C425 VDD1.t0 VSUBS 1.3114f
C426 VP.t0 VSUBS 0.447085f
C427 VP.t1 VSUBS 0.384444f
C428 VP.n0 VSUBS 2.76217f
C429 VDD2.t1 VSUBS 1.3144f
C430 VDD2.t0 VSUBS 1.02647f
C431 VDD2.n0 VSUBS 2.22864f
C432 VTAIL.t0 VSUBS 1.2796f
C433 VTAIL.n0 VSUBS 1.58706f
C434 VTAIL.t3 VSUBS 1.27961f
C435 VTAIL.n1 VSUBS 1.59453f
C436 VTAIL.t1 VSUBS 1.27961f
C437 VTAIL.n2 VSUBS 1.54625f
C438 VTAIL.t2 VSUBS 1.2796f
C439 VTAIL.n3 VSUBS 1.49253f
C440 VN.t0 VSUBS 0.378293f
C441 VN.t1 VSUBS 0.441787f
.ends

