* NGSPICE file created from diff_pair_sample_0248.ext - technology: sky130A

.subckt diff_pair_sample_0248 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=1.9344 pd=10.7 as=0 ps=0 w=4.96 l=1.28
X1 VTAIL.t19 VN.t0 VDD2.t5 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X2 VTAIL.t18 VN.t1 VDD2.t1 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X3 VDD2.t2 VN.t2 VTAIL.t17 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=1.9344 pd=10.7 as=0.8184 ps=5.29 w=4.96 l=1.28
X4 VTAIL.t4 VP.t0 VDD1.t9 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X5 VDD1.t8 VP.t1 VTAIL.t7 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X6 VDD2.t0 VN.t3 VTAIL.t16 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X7 VTAIL.t15 VN.t4 VDD2.t3 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X8 VDD2.t6 VN.t5 VTAIL.t14 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X9 VDD1.t7 VP.t2 VTAIL.t9 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=1.9344 pd=10.7 as=0.8184 ps=5.29 w=4.96 l=1.28
X10 VDD2.t7 VN.t6 VTAIL.t13 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=1.9344 ps=10.7 w=4.96 l=1.28
X11 VDD1.t6 VP.t3 VTAIL.t2 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=1.9344 ps=10.7 w=4.96 l=1.28
X12 B.t8 B.t6 B.t7 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=1.9344 pd=10.7 as=0 ps=0 w=4.96 l=1.28
X13 VTAIL.t8 VP.t4 VDD1.t5 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X14 VDD1.t4 VP.t5 VTAIL.t3 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=1.9344 pd=10.7 as=0.8184 ps=5.29 w=4.96 l=1.28
X15 VDD2.t8 VN.t7 VTAIL.t12 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=1.9344 pd=10.7 as=0.8184 ps=5.29 w=4.96 l=1.28
X16 VDD1.t3 VP.t6 VTAIL.t5 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X17 VTAIL.t6 VP.t7 VDD1.t2 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X18 VTAIL.t11 VN.t8 VDD2.t9 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X19 VDD2.t4 VN.t9 VTAIL.t10 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=1.9344 ps=10.7 w=4.96 l=1.28
X20 VTAIL.t1 VP.t8 VDD1.t1 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=0.8184 ps=5.29 w=4.96 l=1.28
X21 VDD1.t0 VP.t9 VTAIL.t0 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=0.8184 pd=5.29 as=1.9344 ps=10.7 w=4.96 l=1.28
X22 B.t5 B.t3 B.t4 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=1.9344 pd=10.7 as=0 ps=0 w=4.96 l=1.28
X23 B.t2 B.t0 B.t1 w_n2902_n1960# sky130_fd_pr__pfet_01v8 ad=1.9344 pd=10.7 as=0 ps=0 w=4.96 l=1.28
R0 B.n265 B.n264 585
R1 B.n263 B.n88 585
R2 B.n262 B.n261 585
R3 B.n260 B.n89 585
R4 B.n259 B.n258 585
R5 B.n257 B.n90 585
R6 B.n256 B.n255 585
R7 B.n254 B.n91 585
R8 B.n253 B.n252 585
R9 B.n251 B.n92 585
R10 B.n250 B.n249 585
R11 B.n248 B.n93 585
R12 B.n247 B.n246 585
R13 B.n245 B.n94 585
R14 B.n244 B.n243 585
R15 B.n242 B.n95 585
R16 B.n241 B.n240 585
R17 B.n239 B.n96 585
R18 B.n238 B.n237 585
R19 B.n236 B.n97 585
R20 B.n235 B.n234 585
R21 B.n232 B.n98 585
R22 B.n231 B.n230 585
R23 B.n229 B.n101 585
R24 B.n228 B.n227 585
R25 B.n226 B.n102 585
R26 B.n225 B.n224 585
R27 B.n223 B.n103 585
R28 B.n222 B.n221 585
R29 B.n220 B.n104 585
R30 B.n218 B.n217 585
R31 B.n216 B.n107 585
R32 B.n215 B.n214 585
R33 B.n213 B.n108 585
R34 B.n212 B.n211 585
R35 B.n210 B.n109 585
R36 B.n209 B.n208 585
R37 B.n207 B.n110 585
R38 B.n206 B.n205 585
R39 B.n204 B.n111 585
R40 B.n203 B.n202 585
R41 B.n201 B.n112 585
R42 B.n200 B.n199 585
R43 B.n198 B.n113 585
R44 B.n197 B.n196 585
R45 B.n195 B.n114 585
R46 B.n194 B.n193 585
R47 B.n192 B.n115 585
R48 B.n191 B.n190 585
R49 B.n189 B.n116 585
R50 B.n188 B.n187 585
R51 B.n266 B.n87 585
R52 B.n268 B.n267 585
R53 B.n269 B.n86 585
R54 B.n271 B.n270 585
R55 B.n272 B.n85 585
R56 B.n274 B.n273 585
R57 B.n275 B.n84 585
R58 B.n277 B.n276 585
R59 B.n278 B.n83 585
R60 B.n280 B.n279 585
R61 B.n281 B.n82 585
R62 B.n283 B.n282 585
R63 B.n284 B.n81 585
R64 B.n286 B.n285 585
R65 B.n287 B.n80 585
R66 B.n289 B.n288 585
R67 B.n290 B.n79 585
R68 B.n292 B.n291 585
R69 B.n293 B.n78 585
R70 B.n295 B.n294 585
R71 B.n296 B.n77 585
R72 B.n298 B.n297 585
R73 B.n299 B.n76 585
R74 B.n301 B.n300 585
R75 B.n302 B.n75 585
R76 B.n304 B.n303 585
R77 B.n305 B.n74 585
R78 B.n307 B.n306 585
R79 B.n308 B.n73 585
R80 B.n310 B.n309 585
R81 B.n311 B.n72 585
R82 B.n313 B.n312 585
R83 B.n314 B.n71 585
R84 B.n316 B.n315 585
R85 B.n317 B.n70 585
R86 B.n319 B.n318 585
R87 B.n320 B.n69 585
R88 B.n322 B.n321 585
R89 B.n323 B.n68 585
R90 B.n325 B.n324 585
R91 B.n326 B.n67 585
R92 B.n328 B.n327 585
R93 B.n329 B.n66 585
R94 B.n331 B.n330 585
R95 B.n332 B.n65 585
R96 B.n334 B.n333 585
R97 B.n335 B.n64 585
R98 B.n337 B.n336 585
R99 B.n338 B.n63 585
R100 B.n340 B.n339 585
R101 B.n341 B.n62 585
R102 B.n343 B.n342 585
R103 B.n344 B.n61 585
R104 B.n346 B.n345 585
R105 B.n347 B.n60 585
R106 B.n349 B.n348 585
R107 B.n350 B.n59 585
R108 B.n352 B.n351 585
R109 B.n353 B.n58 585
R110 B.n355 B.n354 585
R111 B.n356 B.n57 585
R112 B.n358 B.n357 585
R113 B.n359 B.n56 585
R114 B.n361 B.n360 585
R115 B.n362 B.n55 585
R116 B.n364 B.n363 585
R117 B.n365 B.n54 585
R118 B.n367 B.n366 585
R119 B.n368 B.n53 585
R120 B.n370 B.n369 585
R121 B.n371 B.n52 585
R122 B.n373 B.n372 585
R123 B.n374 B.n51 585
R124 B.n376 B.n375 585
R125 B.n453 B.n20 585
R126 B.n452 B.n451 585
R127 B.n450 B.n21 585
R128 B.n449 B.n448 585
R129 B.n447 B.n22 585
R130 B.n446 B.n445 585
R131 B.n444 B.n23 585
R132 B.n443 B.n442 585
R133 B.n441 B.n24 585
R134 B.n440 B.n439 585
R135 B.n438 B.n25 585
R136 B.n437 B.n436 585
R137 B.n435 B.n26 585
R138 B.n434 B.n433 585
R139 B.n432 B.n27 585
R140 B.n431 B.n430 585
R141 B.n429 B.n28 585
R142 B.n428 B.n427 585
R143 B.n426 B.n29 585
R144 B.n425 B.n424 585
R145 B.n423 B.n30 585
R146 B.n422 B.n421 585
R147 B.n420 B.n31 585
R148 B.n419 B.n418 585
R149 B.n417 B.n35 585
R150 B.n416 B.n415 585
R151 B.n414 B.n36 585
R152 B.n413 B.n412 585
R153 B.n411 B.n37 585
R154 B.n410 B.n409 585
R155 B.n407 B.n38 585
R156 B.n406 B.n405 585
R157 B.n404 B.n41 585
R158 B.n403 B.n402 585
R159 B.n401 B.n42 585
R160 B.n400 B.n399 585
R161 B.n398 B.n43 585
R162 B.n397 B.n396 585
R163 B.n395 B.n44 585
R164 B.n394 B.n393 585
R165 B.n392 B.n45 585
R166 B.n391 B.n390 585
R167 B.n389 B.n46 585
R168 B.n388 B.n387 585
R169 B.n386 B.n47 585
R170 B.n385 B.n384 585
R171 B.n383 B.n48 585
R172 B.n382 B.n381 585
R173 B.n380 B.n49 585
R174 B.n379 B.n378 585
R175 B.n377 B.n50 585
R176 B.n455 B.n454 585
R177 B.n456 B.n19 585
R178 B.n458 B.n457 585
R179 B.n459 B.n18 585
R180 B.n461 B.n460 585
R181 B.n462 B.n17 585
R182 B.n464 B.n463 585
R183 B.n465 B.n16 585
R184 B.n467 B.n466 585
R185 B.n468 B.n15 585
R186 B.n470 B.n469 585
R187 B.n471 B.n14 585
R188 B.n473 B.n472 585
R189 B.n474 B.n13 585
R190 B.n476 B.n475 585
R191 B.n477 B.n12 585
R192 B.n479 B.n478 585
R193 B.n480 B.n11 585
R194 B.n482 B.n481 585
R195 B.n483 B.n10 585
R196 B.n485 B.n484 585
R197 B.n486 B.n9 585
R198 B.n488 B.n487 585
R199 B.n489 B.n8 585
R200 B.n491 B.n490 585
R201 B.n492 B.n7 585
R202 B.n494 B.n493 585
R203 B.n495 B.n6 585
R204 B.n497 B.n496 585
R205 B.n498 B.n5 585
R206 B.n500 B.n499 585
R207 B.n501 B.n4 585
R208 B.n503 B.n502 585
R209 B.n504 B.n3 585
R210 B.n506 B.n505 585
R211 B.n507 B.n0 585
R212 B.n2 B.n1 585
R213 B.n135 B.n134 585
R214 B.n137 B.n136 585
R215 B.n138 B.n133 585
R216 B.n140 B.n139 585
R217 B.n141 B.n132 585
R218 B.n143 B.n142 585
R219 B.n144 B.n131 585
R220 B.n146 B.n145 585
R221 B.n147 B.n130 585
R222 B.n149 B.n148 585
R223 B.n150 B.n129 585
R224 B.n152 B.n151 585
R225 B.n153 B.n128 585
R226 B.n155 B.n154 585
R227 B.n156 B.n127 585
R228 B.n158 B.n157 585
R229 B.n159 B.n126 585
R230 B.n161 B.n160 585
R231 B.n162 B.n125 585
R232 B.n164 B.n163 585
R233 B.n165 B.n124 585
R234 B.n167 B.n166 585
R235 B.n168 B.n123 585
R236 B.n170 B.n169 585
R237 B.n171 B.n122 585
R238 B.n173 B.n172 585
R239 B.n174 B.n121 585
R240 B.n176 B.n175 585
R241 B.n177 B.n120 585
R242 B.n179 B.n178 585
R243 B.n180 B.n119 585
R244 B.n182 B.n181 585
R245 B.n183 B.n118 585
R246 B.n185 B.n184 585
R247 B.n186 B.n117 585
R248 B.n187 B.n186 535.745
R249 B.n266 B.n265 535.745
R250 B.n375 B.n50 535.745
R251 B.n454 B.n453 535.745
R252 B.n105 B.t3 297.902
R253 B.n99 B.t6 297.902
R254 B.n39 B.t0 297.902
R255 B.n32 B.t9 297.902
R256 B.n509 B.n508 256.663
R257 B.n508 B.n507 235.042
R258 B.n508 B.n2 235.042
R259 B.n187 B.n116 163.367
R260 B.n191 B.n116 163.367
R261 B.n192 B.n191 163.367
R262 B.n193 B.n192 163.367
R263 B.n193 B.n114 163.367
R264 B.n197 B.n114 163.367
R265 B.n198 B.n197 163.367
R266 B.n199 B.n198 163.367
R267 B.n199 B.n112 163.367
R268 B.n203 B.n112 163.367
R269 B.n204 B.n203 163.367
R270 B.n205 B.n204 163.367
R271 B.n205 B.n110 163.367
R272 B.n209 B.n110 163.367
R273 B.n210 B.n209 163.367
R274 B.n211 B.n210 163.367
R275 B.n211 B.n108 163.367
R276 B.n215 B.n108 163.367
R277 B.n216 B.n215 163.367
R278 B.n217 B.n216 163.367
R279 B.n217 B.n104 163.367
R280 B.n222 B.n104 163.367
R281 B.n223 B.n222 163.367
R282 B.n224 B.n223 163.367
R283 B.n224 B.n102 163.367
R284 B.n228 B.n102 163.367
R285 B.n229 B.n228 163.367
R286 B.n230 B.n229 163.367
R287 B.n230 B.n98 163.367
R288 B.n235 B.n98 163.367
R289 B.n236 B.n235 163.367
R290 B.n237 B.n236 163.367
R291 B.n237 B.n96 163.367
R292 B.n241 B.n96 163.367
R293 B.n242 B.n241 163.367
R294 B.n243 B.n242 163.367
R295 B.n243 B.n94 163.367
R296 B.n247 B.n94 163.367
R297 B.n248 B.n247 163.367
R298 B.n249 B.n248 163.367
R299 B.n249 B.n92 163.367
R300 B.n253 B.n92 163.367
R301 B.n254 B.n253 163.367
R302 B.n255 B.n254 163.367
R303 B.n255 B.n90 163.367
R304 B.n259 B.n90 163.367
R305 B.n260 B.n259 163.367
R306 B.n261 B.n260 163.367
R307 B.n261 B.n88 163.367
R308 B.n265 B.n88 163.367
R309 B.n375 B.n374 163.367
R310 B.n374 B.n373 163.367
R311 B.n373 B.n52 163.367
R312 B.n369 B.n52 163.367
R313 B.n369 B.n368 163.367
R314 B.n368 B.n367 163.367
R315 B.n367 B.n54 163.367
R316 B.n363 B.n54 163.367
R317 B.n363 B.n362 163.367
R318 B.n362 B.n361 163.367
R319 B.n361 B.n56 163.367
R320 B.n357 B.n56 163.367
R321 B.n357 B.n356 163.367
R322 B.n356 B.n355 163.367
R323 B.n355 B.n58 163.367
R324 B.n351 B.n58 163.367
R325 B.n351 B.n350 163.367
R326 B.n350 B.n349 163.367
R327 B.n349 B.n60 163.367
R328 B.n345 B.n60 163.367
R329 B.n345 B.n344 163.367
R330 B.n344 B.n343 163.367
R331 B.n343 B.n62 163.367
R332 B.n339 B.n62 163.367
R333 B.n339 B.n338 163.367
R334 B.n338 B.n337 163.367
R335 B.n337 B.n64 163.367
R336 B.n333 B.n64 163.367
R337 B.n333 B.n332 163.367
R338 B.n332 B.n331 163.367
R339 B.n331 B.n66 163.367
R340 B.n327 B.n66 163.367
R341 B.n327 B.n326 163.367
R342 B.n326 B.n325 163.367
R343 B.n325 B.n68 163.367
R344 B.n321 B.n68 163.367
R345 B.n321 B.n320 163.367
R346 B.n320 B.n319 163.367
R347 B.n319 B.n70 163.367
R348 B.n315 B.n70 163.367
R349 B.n315 B.n314 163.367
R350 B.n314 B.n313 163.367
R351 B.n313 B.n72 163.367
R352 B.n309 B.n72 163.367
R353 B.n309 B.n308 163.367
R354 B.n308 B.n307 163.367
R355 B.n307 B.n74 163.367
R356 B.n303 B.n74 163.367
R357 B.n303 B.n302 163.367
R358 B.n302 B.n301 163.367
R359 B.n301 B.n76 163.367
R360 B.n297 B.n76 163.367
R361 B.n297 B.n296 163.367
R362 B.n296 B.n295 163.367
R363 B.n295 B.n78 163.367
R364 B.n291 B.n78 163.367
R365 B.n291 B.n290 163.367
R366 B.n290 B.n289 163.367
R367 B.n289 B.n80 163.367
R368 B.n285 B.n80 163.367
R369 B.n285 B.n284 163.367
R370 B.n284 B.n283 163.367
R371 B.n283 B.n82 163.367
R372 B.n279 B.n82 163.367
R373 B.n279 B.n278 163.367
R374 B.n278 B.n277 163.367
R375 B.n277 B.n84 163.367
R376 B.n273 B.n84 163.367
R377 B.n273 B.n272 163.367
R378 B.n272 B.n271 163.367
R379 B.n271 B.n86 163.367
R380 B.n267 B.n86 163.367
R381 B.n267 B.n266 163.367
R382 B.n453 B.n452 163.367
R383 B.n452 B.n21 163.367
R384 B.n448 B.n21 163.367
R385 B.n448 B.n447 163.367
R386 B.n447 B.n446 163.367
R387 B.n446 B.n23 163.367
R388 B.n442 B.n23 163.367
R389 B.n442 B.n441 163.367
R390 B.n441 B.n440 163.367
R391 B.n440 B.n25 163.367
R392 B.n436 B.n25 163.367
R393 B.n436 B.n435 163.367
R394 B.n435 B.n434 163.367
R395 B.n434 B.n27 163.367
R396 B.n430 B.n27 163.367
R397 B.n430 B.n429 163.367
R398 B.n429 B.n428 163.367
R399 B.n428 B.n29 163.367
R400 B.n424 B.n29 163.367
R401 B.n424 B.n423 163.367
R402 B.n423 B.n422 163.367
R403 B.n422 B.n31 163.367
R404 B.n418 B.n31 163.367
R405 B.n418 B.n417 163.367
R406 B.n417 B.n416 163.367
R407 B.n416 B.n36 163.367
R408 B.n412 B.n36 163.367
R409 B.n412 B.n411 163.367
R410 B.n411 B.n410 163.367
R411 B.n410 B.n38 163.367
R412 B.n405 B.n38 163.367
R413 B.n405 B.n404 163.367
R414 B.n404 B.n403 163.367
R415 B.n403 B.n42 163.367
R416 B.n399 B.n42 163.367
R417 B.n399 B.n398 163.367
R418 B.n398 B.n397 163.367
R419 B.n397 B.n44 163.367
R420 B.n393 B.n44 163.367
R421 B.n393 B.n392 163.367
R422 B.n392 B.n391 163.367
R423 B.n391 B.n46 163.367
R424 B.n387 B.n46 163.367
R425 B.n387 B.n386 163.367
R426 B.n386 B.n385 163.367
R427 B.n385 B.n48 163.367
R428 B.n381 B.n48 163.367
R429 B.n381 B.n380 163.367
R430 B.n380 B.n379 163.367
R431 B.n379 B.n50 163.367
R432 B.n454 B.n19 163.367
R433 B.n458 B.n19 163.367
R434 B.n459 B.n458 163.367
R435 B.n460 B.n459 163.367
R436 B.n460 B.n17 163.367
R437 B.n464 B.n17 163.367
R438 B.n465 B.n464 163.367
R439 B.n466 B.n465 163.367
R440 B.n466 B.n15 163.367
R441 B.n470 B.n15 163.367
R442 B.n471 B.n470 163.367
R443 B.n472 B.n471 163.367
R444 B.n472 B.n13 163.367
R445 B.n476 B.n13 163.367
R446 B.n477 B.n476 163.367
R447 B.n478 B.n477 163.367
R448 B.n478 B.n11 163.367
R449 B.n482 B.n11 163.367
R450 B.n483 B.n482 163.367
R451 B.n484 B.n483 163.367
R452 B.n484 B.n9 163.367
R453 B.n488 B.n9 163.367
R454 B.n489 B.n488 163.367
R455 B.n490 B.n489 163.367
R456 B.n490 B.n7 163.367
R457 B.n494 B.n7 163.367
R458 B.n495 B.n494 163.367
R459 B.n496 B.n495 163.367
R460 B.n496 B.n5 163.367
R461 B.n500 B.n5 163.367
R462 B.n501 B.n500 163.367
R463 B.n502 B.n501 163.367
R464 B.n502 B.n3 163.367
R465 B.n506 B.n3 163.367
R466 B.n507 B.n506 163.367
R467 B.n134 B.n2 163.367
R468 B.n137 B.n134 163.367
R469 B.n138 B.n137 163.367
R470 B.n139 B.n138 163.367
R471 B.n139 B.n132 163.367
R472 B.n143 B.n132 163.367
R473 B.n144 B.n143 163.367
R474 B.n145 B.n144 163.367
R475 B.n145 B.n130 163.367
R476 B.n149 B.n130 163.367
R477 B.n150 B.n149 163.367
R478 B.n151 B.n150 163.367
R479 B.n151 B.n128 163.367
R480 B.n155 B.n128 163.367
R481 B.n156 B.n155 163.367
R482 B.n157 B.n156 163.367
R483 B.n157 B.n126 163.367
R484 B.n161 B.n126 163.367
R485 B.n162 B.n161 163.367
R486 B.n163 B.n162 163.367
R487 B.n163 B.n124 163.367
R488 B.n167 B.n124 163.367
R489 B.n168 B.n167 163.367
R490 B.n169 B.n168 163.367
R491 B.n169 B.n122 163.367
R492 B.n173 B.n122 163.367
R493 B.n174 B.n173 163.367
R494 B.n175 B.n174 163.367
R495 B.n175 B.n120 163.367
R496 B.n179 B.n120 163.367
R497 B.n180 B.n179 163.367
R498 B.n181 B.n180 163.367
R499 B.n181 B.n118 163.367
R500 B.n185 B.n118 163.367
R501 B.n186 B.n185 163.367
R502 B.n99 B.t7 149.674
R503 B.n39 B.t2 149.674
R504 B.n105 B.t4 149.671
R505 B.n32 B.t11 149.671
R506 B.n100 B.t8 118.451
R507 B.n40 B.t1 118.451
R508 B.n106 B.t5 118.447
R509 B.n33 B.t10 118.447
R510 B.n219 B.n106 59.5399
R511 B.n233 B.n100 59.5399
R512 B.n408 B.n40 59.5399
R513 B.n34 B.n33 59.5399
R514 B.n455 B.n20 34.8103
R515 B.n377 B.n376 34.8103
R516 B.n264 B.n87 34.8103
R517 B.n188 B.n117 34.8103
R518 B.n106 B.n105 31.2247
R519 B.n100 B.n99 31.2247
R520 B.n40 B.n39 31.2247
R521 B.n33 B.n32 31.2247
R522 B B.n509 18.0485
R523 B.n456 B.n455 10.6151
R524 B.n457 B.n456 10.6151
R525 B.n457 B.n18 10.6151
R526 B.n461 B.n18 10.6151
R527 B.n462 B.n461 10.6151
R528 B.n463 B.n462 10.6151
R529 B.n463 B.n16 10.6151
R530 B.n467 B.n16 10.6151
R531 B.n468 B.n467 10.6151
R532 B.n469 B.n468 10.6151
R533 B.n469 B.n14 10.6151
R534 B.n473 B.n14 10.6151
R535 B.n474 B.n473 10.6151
R536 B.n475 B.n474 10.6151
R537 B.n475 B.n12 10.6151
R538 B.n479 B.n12 10.6151
R539 B.n480 B.n479 10.6151
R540 B.n481 B.n480 10.6151
R541 B.n481 B.n10 10.6151
R542 B.n485 B.n10 10.6151
R543 B.n486 B.n485 10.6151
R544 B.n487 B.n486 10.6151
R545 B.n487 B.n8 10.6151
R546 B.n491 B.n8 10.6151
R547 B.n492 B.n491 10.6151
R548 B.n493 B.n492 10.6151
R549 B.n493 B.n6 10.6151
R550 B.n497 B.n6 10.6151
R551 B.n498 B.n497 10.6151
R552 B.n499 B.n498 10.6151
R553 B.n499 B.n4 10.6151
R554 B.n503 B.n4 10.6151
R555 B.n504 B.n503 10.6151
R556 B.n505 B.n504 10.6151
R557 B.n505 B.n0 10.6151
R558 B.n451 B.n20 10.6151
R559 B.n451 B.n450 10.6151
R560 B.n450 B.n449 10.6151
R561 B.n449 B.n22 10.6151
R562 B.n445 B.n22 10.6151
R563 B.n445 B.n444 10.6151
R564 B.n444 B.n443 10.6151
R565 B.n443 B.n24 10.6151
R566 B.n439 B.n24 10.6151
R567 B.n439 B.n438 10.6151
R568 B.n438 B.n437 10.6151
R569 B.n437 B.n26 10.6151
R570 B.n433 B.n26 10.6151
R571 B.n433 B.n432 10.6151
R572 B.n432 B.n431 10.6151
R573 B.n431 B.n28 10.6151
R574 B.n427 B.n28 10.6151
R575 B.n427 B.n426 10.6151
R576 B.n426 B.n425 10.6151
R577 B.n425 B.n30 10.6151
R578 B.n421 B.n420 10.6151
R579 B.n420 B.n419 10.6151
R580 B.n419 B.n35 10.6151
R581 B.n415 B.n35 10.6151
R582 B.n415 B.n414 10.6151
R583 B.n414 B.n413 10.6151
R584 B.n413 B.n37 10.6151
R585 B.n409 B.n37 10.6151
R586 B.n407 B.n406 10.6151
R587 B.n406 B.n41 10.6151
R588 B.n402 B.n41 10.6151
R589 B.n402 B.n401 10.6151
R590 B.n401 B.n400 10.6151
R591 B.n400 B.n43 10.6151
R592 B.n396 B.n43 10.6151
R593 B.n396 B.n395 10.6151
R594 B.n395 B.n394 10.6151
R595 B.n394 B.n45 10.6151
R596 B.n390 B.n45 10.6151
R597 B.n390 B.n389 10.6151
R598 B.n389 B.n388 10.6151
R599 B.n388 B.n47 10.6151
R600 B.n384 B.n47 10.6151
R601 B.n384 B.n383 10.6151
R602 B.n383 B.n382 10.6151
R603 B.n382 B.n49 10.6151
R604 B.n378 B.n49 10.6151
R605 B.n378 B.n377 10.6151
R606 B.n376 B.n51 10.6151
R607 B.n372 B.n51 10.6151
R608 B.n372 B.n371 10.6151
R609 B.n371 B.n370 10.6151
R610 B.n370 B.n53 10.6151
R611 B.n366 B.n53 10.6151
R612 B.n366 B.n365 10.6151
R613 B.n365 B.n364 10.6151
R614 B.n364 B.n55 10.6151
R615 B.n360 B.n55 10.6151
R616 B.n360 B.n359 10.6151
R617 B.n359 B.n358 10.6151
R618 B.n358 B.n57 10.6151
R619 B.n354 B.n57 10.6151
R620 B.n354 B.n353 10.6151
R621 B.n353 B.n352 10.6151
R622 B.n352 B.n59 10.6151
R623 B.n348 B.n59 10.6151
R624 B.n348 B.n347 10.6151
R625 B.n347 B.n346 10.6151
R626 B.n346 B.n61 10.6151
R627 B.n342 B.n61 10.6151
R628 B.n342 B.n341 10.6151
R629 B.n341 B.n340 10.6151
R630 B.n340 B.n63 10.6151
R631 B.n336 B.n63 10.6151
R632 B.n336 B.n335 10.6151
R633 B.n335 B.n334 10.6151
R634 B.n334 B.n65 10.6151
R635 B.n330 B.n65 10.6151
R636 B.n330 B.n329 10.6151
R637 B.n329 B.n328 10.6151
R638 B.n328 B.n67 10.6151
R639 B.n324 B.n67 10.6151
R640 B.n324 B.n323 10.6151
R641 B.n323 B.n322 10.6151
R642 B.n322 B.n69 10.6151
R643 B.n318 B.n69 10.6151
R644 B.n318 B.n317 10.6151
R645 B.n317 B.n316 10.6151
R646 B.n316 B.n71 10.6151
R647 B.n312 B.n71 10.6151
R648 B.n312 B.n311 10.6151
R649 B.n311 B.n310 10.6151
R650 B.n310 B.n73 10.6151
R651 B.n306 B.n73 10.6151
R652 B.n306 B.n305 10.6151
R653 B.n305 B.n304 10.6151
R654 B.n304 B.n75 10.6151
R655 B.n300 B.n75 10.6151
R656 B.n300 B.n299 10.6151
R657 B.n299 B.n298 10.6151
R658 B.n298 B.n77 10.6151
R659 B.n294 B.n77 10.6151
R660 B.n294 B.n293 10.6151
R661 B.n293 B.n292 10.6151
R662 B.n292 B.n79 10.6151
R663 B.n288 B.n79 10.6151
R664 B.n288 B.n287 10.6151
R665 B.n287 B.n286 10.6151
R666 B.n286 B.n81 10.6151
R667 B.n282 B.n81 10.6151
R668 B.n282 B.n281 10.6151
R669 B.n281 B.n280 10.6151
R670 B.n280 B.n83 10.6151
R671 B.n276 B.n83 10.6151
R672 B.n276 B.n275 10.6151
R673 B.n275 B.n274 10.6151
R674 B.n274 B.n85 10.6151
R675 B.n270 B.n85 10.6151
R676 B.n270 B.n269 10.6151
R677 B.n269 B.n268 10.6151
R678 B.n268 B.n87 10.6151
R679 B.n135 B.n1 10.6151
R680 B.n136 B.n135 10.6151
R681 B.n136 B.n133 10.6151
R682 B.n140 B.n133 10.6151
R683 B.n141 B.n140 10.6151
R684 B.n142 B.n141 10.6151
R685 B.n142 B.n131 10.6151
R686 B.n146 B.n131 10.6151
R687 B.n147 B.n146 10.6151
R688 B.n148 B.n147 10.6151
R689 B.n148 B.n129 10.6151
R690 B.n152 B.n129 10.6151
R691 B.n153 B.n152 10.6151
R692 B.n154 B.n153 10.6151
R693 B.n154 B.n127 10.6151
R694 B.n158 B.n127 10.6151
R695 B.n159 B.n158 10.6151
R696 B.n160 B.n159 10.6151
R697 B.n160 B.n125 10.6151
R698 B.n164 B.n125 10.6151
R699 B.n165 B.n164 10.6151
R700 B.n166 B.n165 10.6151
R701 B.n166 B.n123 10.6151
R702 B.n170 B.n123 10.6151
R703 B.n171 B.n170 10.6151
R704 B.n172 B.n171 10.6151
R705 B.n172 B.n121 10.6151
R706 B.n176 B.n121 10.6151
R707 B.n177 B.n176 10.6151
R708 B.n178 B.n177 10.6151
R709 B.n178 B.n119 10.6151
R710 B.n182 B.n119 10.6151
R711 B.n183 B.n182 10.6151
R712 B.n184 B.n183 10.6151
R713 B.n184 B.n117 10.6151
R714 B.n189 B.n188 10.6151
R715 B.n190 B.n189 10.6151
R716 B.n190 B.n115 10.6151
R717 B.n194 B.n115 10.6151
R718 B.n195 B.n194 10.6151
R719 B.n196 B.n195 10.6151
R720 B.n196 B.n113 10.6151
R721 B.n200 B.n113 10.6151
R722 B.n201 B.n200 10.6151
R723 B.n202 B.n201 10.6151
R724 B.n202 B.n111 10.6151
R725 B.n206 B.n111 10.6151
R726 B.n207 B.n206 10.6151
R727 B.n208 B.n207 10.6151
R728 B.n208 B.n109 10.6151
R729 B.n212 B.n109 10.6151
R730 B.n213 B.n212 10.6151
R731 B.n214 B.n213 10.6151
R732 B.n214 B.n107 10.6151
R733 B.n218 B.n107 10.6151
R734 B.n221 B.n220 10.6151
R735 B.n221 B.n103 10.6151
R736 B.n225 B.n103 10.6151
R737 B.n226 B.n225 10.6151
R738 B.n227 B.n226 10.6151
R739 B.n227 B.n101 10.6151
R740 B.n231 B.n101 10.6151
R741 B.n232 B.n231 10.6151
R742 B.n234 B.n97 10.6151
R743 B.n238 B.n97 10.6151
R744 B.n239 B.n238 10.6151
R745 B.n240 B.n239 10.6151
R746 B.n240 B.n95 10.6151
R747 B.n244 B.n95 10.6151
R748 B.n245 B.n244 10.6151
R749 B.n246 B.n245 10.6151
R750 B.n246 B.n93 10.6151
R751 B.n250 B.n93 10.6151
R752 B.n251 B.n250 10.6151
R753 B.n252 B.n251 10.6151
R754 B.n252 B.n91 10.6151
R755 B.n256 B.n91 10.6151
R756 B.n257 B.n256 10.6151
R757 B.n258 B.n257 10.6151
R758 B.n258 B.n89 10.6151
R759 B.n262 B.n89 10.6151
R760 B.n263 B.n262 10.6151
R761 B.n264 B.n263 10.6151
R762 B.n509 B.n0 8.11757
R763 B.n509 B.n1 8.11757
R764 B.n421 B.n34 6.5566
R765 B.n409 B.n408 6.5566
R766 B.n220 B.n219 6.5566
R767 B.n233 B.n232 6.5566
R768 B.n34 B.n30 4.05904
R769 B.n408 B.n407 4.05904
R770 B.n219 B.n218 4.05904
R771 B.n234 B.n233 4.05904
R772 VN.n24 VN.n23 175.071
R773 VN.n49 VN.n48 175.071
R774 VN.n47 VN.n25 161.3
R775 VN.n46 VN.n45 161.3
R776 VN.n44 VN.n26 161.3
R777 VN.n43 VN.n42 161.3
R778 VN.n41 VN.n27 161.3
R779 VN.n40 VN.n39 161.3
R780 VN.n38 VN.n29 161.3
R781 VN.n37 VN.n36 161.3
R782 VN.n35 VN.n30 161.3
R783 VN.n34 VN.n33 161.3
R784 VN.n22 VN.n0 161.3
R785 VN.n21 VN.n20 161.3
R786 VN.n19 VN.n1 161.3
R787 VN.n18 VN.n17 161.3
R788 VN.n15 VN.n2 161.3
R789 VN.n14 VN.n13 161.3
R790 VN.n12 VN.n3 161.3
R791 VN.n11 VN.n10 161.3
R792 VN.n9 VN.n4 161.3
R793 VN.n8 VN.n7 161.3
R794 VN.n6 VN.t2 121.617
R795 VN.n32 VN.t6 121.617
R796 VN.n3 VN.t5 93.388
R797 VN.n5 VN.t1 93.388
R798 VN.n16 VN.t0 93.388
R799 VN.n23 VN.t9 93.388
R800 VN.n29 VN.t3 93.388
R801 VN.n31 VN.t4 93.388
R802 VN.n28 VN.t8 93.388
R803 VN.n48 VN.t7 93.388
R804 VN.n6 VN.n5 59.8719
R805 VN.n32 VN.n31 59.8719
R806 VN.n10 VN.n9 56.5617
R807 VN.n15 VN.n14 56.5617
R808 VN.n36 VN.n35 56.5617
R809 VN.n41 VN.n40 56.5617
R810 VN.n21 VN.n1 48.8116
R811 VN.n46 VN.n26 48.8116
R812 VN VN.n49 40.8698
R813 VN.n22 VN.n21 32.3425
R814 VN.n47 VN.n46 32.3425
R815 VN.n33 VN.n32 27.4672
R816 VN.n7 VN.n6 27.4672
R817 VN.n9 VN.n8 24.5923
R818 VN.n10 VN.n3 24.5923
R819 VN.n14 VN.n3 24.5923
R820 VN.n17 VN.n15 24.5923
R821 VN.n35 VN.n34 24.5923
R822 VN.n40 VN.n29 24.5923
R823 VN.n36 VN.n29 24.5923
R824 VN.n42 VN.n41 24.5923
R825 VN.n16 VN.n1 19.1821
R826 VN.n28 VN.n26 19.1821
R827 VN.n23 VN.n22 10.8209
R828 VN.n48 VN.n47 10.8209
R829 VN.n8 VN.n5 5.4107
R830 VN.n17 VN.n16 5.4107
R831 VN.n34 VN.n31 5.4107
R832 VN.n42 VN.n28 5.4107
R833 VN.n49 VN.n25 0.189894
R834 VN.n45 VN.n25 0.189894
R835 VN.n45 VN.n44 0.189894
R836 VN.n44 VN.n43 0.189894
R837 VN.n43 VN.n27 0.189894
R838 VN.n39 VN.n27 0.189894
R839 VN.n39 VN.n38 0.189894
R840 VN.n38 VN.n37 0.189894
R841 VN.n37 VN.n30 0.189894
R842 VN.n33 VN.n30 0.189894
R843 VN.n7 VN.n4 0.189894
R844 VN.n11 VN.n4 0.189894
R845 VN.n12 VN.n11 0.189894
R846 VN.n13 VN.n12 0.189894
R847 VN.n13 VN.n2 0.189894
R848 VN.n18 VN.n2 0.189894
R849 VN.n19 VN.n18 0.189894
R850 VN.n20 VN.n19 0.189894
R851 VN.n20 VN.n0 0.189894
R852 VN.n24 VN.n0 0.189894
R853 VN VN.n24 0.0516364
R854 VDD2.n1 VDD2.t2 109.157
R855 VDD2.n4 VDD2.t8 107.769
R856 VDD2.n3 VDD2.n2 102.201
R857 VDD2 VDD2.n7 102.2
R858 VDD2.n6 VDD2.n5 101.216
R859 VDD2.n1 VDD2.n0 101.216
R860 VDD2.n4 VDD2.n3 34.5838
R861 VDD2.n7 VDD2.t3 6.55393
R862 VDD2.n7 VDD2.t7 6.55393
R863 VDD2.n5 VDD2.t9 6.55393
R864 VDD2.n5 VDD2.t0 6.55393
R865 VDD2.n2 VDD2.t5 6.55393
R866 VDD2.n2 VDD2.t4 6.55393
R867 VDD2.n0 VDD2.t1 6.55393
R868 VDD2.n0 VDD2.t6 6.55393
R869 VDD2.n6 VDD2.n4 1.38843
R870 VDD2 VDD2.n6 0.405672
R871 VDD2.n3 VDD2.n1 0.292137
R872 VTAIL.n11 VTAIL.t13 91.0911
R873 VTAIL.n17 VTAIL.t10 91.091
R874 VTAIL.n2 VTAIL.t0 91.091
R875 VTAIL.n16 VTAIL.t2 91.091
R876 VTAIL.n15 VTAIL.n14 84.5378
R877 VTAIL.n13 VTAIL.n12 84.5378
R878 VTAIL.n10 VTAIL.n9 84.5378
R879 VTAIL.n8 VTAIL.n7 84.5378
R880 VTAIL.n19 VTAIL.n18 84.5375
R881 VTAIL.n1 VTAIL.n0 84.5375
R882 VTAIL.n4 VTAIL.n3 84.5375
R883 VTAIL.n6 VTAIL.n5 84.5375
R884 VTAIL.n8 VTAIL.n6 19.4186
R885 VTAIL.n17 VTAIL.n16 18.0307
R886 VTAIL.n18 VTAIL.t14 6.55393
R887 VTAIL.n18 VTAIL.t19 6.55393
R888 VTAIL.n0 VTAIL.t17 6.55393
R889 VTAIL.n0 VTAIL.t18 6.55393
R890 VTAIL.n3 VTAIL.t7 6.55393
R891 VTAIL.n3 VTAIL.t6 6.55393
R892 VTAIL.n5 VTAIL.t9 6.55393
R893 VTAIL.n5 VTAIL.t4 6.55393
R894 VTAIL.n14 VTAIL.t5 6.55393
R895 VTAIL.n14 VTAIL.t8 6.55393
R896 VTAIL.n12 VTAIL.t3 6.55393
R897 VTAIL.n12 VTAIL.t1 6.55393
R898 VTAIL.n9 VTAIL.t16 6.55393
R899 VTAIL.n9 VTAIL.t15 6.55393
R900 VTAIL.n7 VTAIL.t12 6.55393
R901 VTAIL.n7 VTAIL.t11 6.55393
R902 VTAIL.n10 VTAIL.n8 1.38843
R903 VTAIL.n11 VTAIL.n10 1.38843
R904 VTAIL.n15 VTAIL.n13 1.38843
R905 VTAIL.n16 VTAIL.n15 1.38843
R906 VTAIL.n6 VTAIL.n4 1.38843
R907 VTAIL.n4 VTAIL.n2 1.38843
R908 VTAIL.n19 VTAIL.n17 1.38843
R909 VTAIL.n13 VTAIL.n11 1.16429
R910 VTAIL.n2 VTAIL.n1 1.16429
R911 VTAIL VTAIL.n1 1.09964
R912 VTAIL VTAIL.n19 0.289293
R913 VP.n33 VP.n7 175.071
R914 VP.n56 VP.n55 175.071
R915 VP.n32 VP.n31 175.071
R916 VP.n16 VP.n15 161.3
R917 VP.n17 VP.n12 161.3
R918 VP.n19 VP.n18 161.3
R919 VP.n20 VP.n11 161.3
R920 VP.n22 VP.n21 161.3
R921 VP.n23 VP.n10 161.3
R922 VP.n26 VP.n25 161.3
R923 VP.n27 VP.n9 161.3
R924 VP.n29 VP.n28 161.3
R925 VP.n30 VP.n8 161.3
R926 VP.n54 VP.n0 161.3
R927 VP.n53 VP.n52 161.3
R928 VP.n51 VP.n1 161.3
R929 VP.n50 VP.n49 161.3
R930 VP.n47 VP.n2 161.3
R931 VP.n46 VP.n45 161.3
R932 VP.n44 VP.n3 161.3
R933 VP.n43 VP.n42 161.3
R934 VP.n41 VP.n4 161.3
R935 VP.n40 VP.n39 161.3
R936 VP.n38 VP.n37 161.3
R937 VP.n36 VP.n6 161.3
R938 VP.n35 VP.n34 161.3
R939 VP.n14 VP.t5 121.617
R940 VP.n3 VP.t1 93.388
R941 VP.n7 VP.t2 93.388
R942 VP.n5 VP.t0 93.388
R943 VP.n48 VP.t7 93.388
R944 VP.n55 VP.t9 93.388
R945 VP.n11 VP.t6 93.388
R946 VP.n31 VP.t3 93.388
R947 VP.n24 VP.t4 93.388
R948 VP.n13 VP.t8 93.388
R949 VP.n14 VP.n13 59.8719
R950 VP.n42 VP.n41 56.5617
R951 VP.n47 VP.n46 56.5617
R952 VP.n23 VP.n22 56.5617
R953 VP.n18 VP.n17 56.5617
R954 VP.n37 VP.n36 48.8116
R955 VP.n53 VP.n1 48.8116
R956 VP.n29 VP.n9 48.8116
R957 VP.n33 VP.n32 40.4891
R958 VP.n36 VP.n35 32.3425
R959 VP.n54 VP.n53 32.3425
R960 VP.n30 VP.n29 32.3425
R961 VP.n15 VP.n14 27.4672
R962 VP.n41 VP.n40 24.5923
R963 VP.n42 VP.n3 24.5923
R964 VP.n46 VP.n3 24.5923
R965 VP.n49 VP.n47 24.5923
R966 VP.n25 VP.n23 24.5923
R967 VP.n18 VP.n11 24.5923
R968 VP.n22 VP.n11 24.5923
R969 VP.n17 VP.n16 24.5923
R970 VP.n37 VP.n5 19.1821
R971 VP.n48 VP.n1 19.1821
R972 VP.n24 VP.n9 19.1821
R973 VP.n35 VP.n7 10.8209
R974 VP.n55 VP.n54 10.8209
R975 VP.n31 VP.n30 10.8209
R976 VP.n40 VP.n5 5.4107
R977 VP.n49 VP.n48 5.4107
R978 VP.n25 VP.n24 5.4107
R979 VP.n16 VP.n13 5.4107
R980 VP.n15 VP.n12 0.189894
R981 VP.n19 VP.n12 0.189894
R982 VP.n20 VP.n19 0.189894
R983 VP.n21 VP.n20 0.189894
R984 VP.n21 VP.n10 0.189894
R985 VP.n26 VP.n10 0.189894
R986 VP.n27 VP.n26 0.189894
R987 VP.n28 VP.n27 0.189894
R988 VP.n28 VP.n8 0.189894
R989 VP.n32 VP.n8 0.189894
R990 VP.n34 VP.n33 0.189894
R991 VP.n34 VP.n6 0.189894
R992 VP.n38 VP.n6 0.189894
R993 VP.n39 VP.n38 0.189894
R994 VP.n39 VP.n4 0.189894
R995 VP.n43 VP.n4 0.189894
R996 VP.n44 VP.n43 0.189894
R997 VP.n45 VP.n44 0.189894
R998 VP.n45 VP.n2 0.189894
R999 VP.n50 VP.n2 0.189894
R1000 VP.n51 VP.n50 0.189894
R1001 VP.n52 VP.n51 0.189894
R1002 VP.n52 VP.n0 0.189894
R1003 VP.n56 VP.n0 0.189894
R1004 VP VP.n56 0.0516364
R1005 VDD1.n1 VDD1.t4 109.157
R1006 VDD1.n3 VDD1.t7 109.157
R1007 VDD1.n5 VDD1.n4 102.201
R1008 VDD1.n1 VDD1.n0 101.216
R1009 VDD1.n7 VDD1.n6 101.216
R1010 VDD1.n3 VDD1.n2 101.216
R1011 VDD1.n7 VDD1.n5 35.8608
R1012 VDD1.n6 VDD1.t5 6.55393
R1013 VDD1.n6 VDD1.t6 6.55393
R1014 VDD1.n0 VDD1.t1 6.55393
R1015 VDD1.n0 VDD1.t3 6.55393
R1016 VDD1.n4 VDD1.t2 6.55393
R1017 VDD1.n4 VDD1.t0 6.55393
R1018 VDD1.n2 VDD1.t9 6.55393
R1019 VDD1.n2 VDD1.t8 6.55393
R1020 VDD1 VDD1.n7 0.983259
R1021 VDD1 VDD1.n1 0.405672
R1022 VDD1.n5 VDD1.n3 0.292137
C0 VN w_n2902_n1960# 5.6764f
C1 w_n2902_n1960# B 6.35733f
C2 VDD1 w_n2902_n1960# 1.7748f
C3 VP VTAIL 4.4082f
C4 VP VDD2 0.419032f
C5 w_n2902_n1960# VTAIL 1.9999f
C6 VN B 0.888265f
C7 w_n2902_n1960# VDD2 1.8495f
C8 VDD1 VN 0.150662f
C9 VDD1 B 1.41911f
C10 VN VTAIL 4.39395f
C11 B VTAIL 1.69628f
C12 VN VDD2 3.89927f
C13 VDD2 B 1.48569f
C14 VDD1 VTAIL 6.58675f
C15 VDD1 VDD2 1.32984f
C16 VP w_n2902_n1960# 6.05007f
C17 VDD2 VTAIL 6.62954f
C18 VP VN 5.14694f
C19 VP B 1.5094f
C20 VDD1 VP 4.16107f
C21 VDD2 VSUBS 1.222228f
C22 VDD1 VSUBS 1.162834f
C23 VTAIL VSUBS 0.480683f
C24 VN VSUBS 5.21597f
C25 VP VSUBS 2.118443f
C26 B VSUBS 2.967847f
C27 w_n2902_n1960# VSUBS 71.2847f
C28 VDD1.t4 VSUBS 0.791386f
C29 VDD1.t1 VSUBS 0.092202f
C30 VDD1.t3 VSUBS 0.092202f
C31 VDD1.n0 VSUBS 0.578175f
C32 VDD1.n1 VSUBS 1.00685f
C33 VDD1.t7 VSUBS 0.791383f
C34 VDD1.t9 VSUBS 0.092202f
C35 VDD1.t8 VSUBS 0.092202f
C36 VDD1.n2 VSUBS 0.578173f
C37 VDD1.n3 VSUBS 1.00012f
C38 VDD1.t2 VSUBS 0.092202f
C39 VDD1.t0 VSUBS 0.092202f
C40 VDD1.n4 VSUBS 0.583466f
C41 VDD1.n5 VSUBS 1.93314f
C42 VDD1.t5 VSUBS 0.092202f
C43 VDD1.t6 VSUBS 0.092202f
C44 VDD1.n6 VSUBS 0.578172f
C45 VDD1.n7 VSUBS 2.11631f
C46 VP.n0 VSUBS 0.051715f
C47 VP.t9 VSUBS 0.858293f
C48 VP.n1 VSUBS 0.085485f
C49 VP.n2 VSUBS 0.051715f
C50 VP.t1 VSUBS 0.858293f
C51 VP.n3 VSUBS 0.402611f
C52 VP.n4 VSUBS 0.051715f
C53 VP.t0 VSUBS 0.858293f
C54 VP.n5 VSUBS 0.354054f
C55 VP.n6 VSUBS 0.051715f
C56 VP.t2 VSUBS 0.858293f
C57 VP.n7 VSUBS 0.442411f
C58 VP.n8 VSUBS 0.051715f
C59 VP.t3 VSUBS 0.858293f
C60 VP.n9 VSUBS 0.085485f
C61 VP.n10 VSUBS 0.051715f
C62 VP.t6 VSUBS 0.858293f
C63 VP.n11 VSUBS 0.402611f
C64 VP.n12 VSUBS 0.051715f
C65 VP.t8 VSUBS 0.858293f
C66 VP.n13 VSUBS 0.424021f
C67 VP.t5 VSUBS 0.977486f
C68 VP.n14 VSUBS 0.465119f
C69 VP.n15 VSUBS 0.270588f
C70 VP.n16 VSUBS 0.058973f
C71 VP.n17 VSUBS 0.067306f
C72 VP.n18 VSUBS 0.083045f
C73 VP.n19 VSUBS 0.051715f
C74 VP.n20 VSUBS 0.051715f
C75 VP.n21 VSUBS 0.051715f
C76 VP.n22 VSUBS 0.083045f
C77 VP.n23 VSUBS 0.067306f
C78 VP.t4 VSUBS 0.858293f
C79 VP.n24 VSUBS 0.354054f
C80 VP.n25 VSUBS 0.058973f
C81 VP.n26 VSUBS 0.051715f
C82 VP.n27 VSUBS 0.051715f
C83 VP.n28 VSUBS 0.051715f
C84 VP.n29 VSUBS 0.046736f
C85 VP.n30 VSUBS 0.077103f
C86 VP.n31 VSUBS 0.442411f
C87 VP.n32 VSUBS 2.01411f
C88 VP.n33 VSUBS 2.06016f
C89 VP.n34 VSUBS 0.051715f
C90 VP.n35 VSUBS 0.077103f
C91 VP.n36 VSUBS 0.046736f
C92 VP.n37 VSUBS 0.085485f
C93 VP.n38 VSUBS 0.051715f
C94 VP.n39 VSUBS 0.051715f
C95 VP.n40 VSUBS 0.058973f
C96 VP.n41 VSUBS 0.067306f
C97 VP.n42 VSUBS 0.083045f
C98 VP.n43 VSUBS 0.051715f
C99 VP.n44 VSUBS 0.051715f
C100 VP.n45 VSUBS 0.051715f
C101 VP.n46 VSUBS 0.083045f
C102 VP.n47 VSUBS 0.067306f
C103 VP.t7 VSUBS 0.858293f
C104 VP.n48 VSUBS 0.354054f
C105 VP.n49 VSUBS 0.058973f
C106 VP.n50 VSUBS 0.051715f
C107 VP.n51 VSUBS 0.051715f
C108 VP.n52 VSUBS 0.051715f
C109 VP.n53 VSUBS 0.046736f
C110 VP.n54 VSUBS 0.077103f
C111 VP.n55 VSUBS 0.442411f
C112 VP.n56 VSUBS 0.047621f
C113 VTAIL.t17 VSUBS 0.109142f
C114 VTAIL.t18 VSUBS 0.109142f
C115 VTAIL.n0 VSUBS 0.601598f
C116 VTAIL.n1 VSUBS 0.672952f
C117 VTAIL.t0 VSUBS 0.842413f
C118 VTAIL.n2 VSUBS 0.755708f
C119 VTAIL.t7 VSUBS 0.109142f
C120 VTAIL.t6 VSUBS 0.109142f
C121 VTAIL.n3 VSUBS 0.601598f
C122 VTAIL.n4 VSUBS 0.718974f
C123 VTAIL.t9 VSUBS 0.109142f
C124 VTAIL.t4 VSUBS 0.109142f
C125 VTAIL.n5 VSUBS 0.601598f
C126 VTAIL.n6 VSUBS 1.60541f
C127 VTAIL.t12 VSUBS 0.109142f
C128 VTAIL.t11 VSUBS 0.109142f
C129 VTAIL.n7 VSUBS 0.601602f
C130 VTAIL.n8 VSUBS 1.6054f
C131 VTAIL.t16 VSUBS 0.109142f
C132 VTAIL.t15 VSUBS 0.109142f
C133 VTAIL.n9 VSUBS 0.601602f
C134 VTAIL.n10 VSUBS 0.718971f
C135 VTAIL.t13 VSUBS 0.842418f
C136 VTAIL.n11 VSUBS 0.755704f
C137 VTAIL.t3 VSUBS 0.109142f
C138 VTAIL.t1 VSUBS 0.109142f
C139 VTAIL.n12 VSUBS 0.601602f
C140 VTAIL.n13 VSUBS 0.69886f
C141 VTAIL.t5 VSUBS 0.109142f
C142 VTAIL.t8 VSUBS 0.109142f
C143 VTAIL.n14 VSUBS 0.601602f
C144 VTAIL.n15 VSUBS 0.718971f
C145 VTAIL.t2 VSUBS 0.842413f
C146 VTAIL.n16 VSUBS 1.53772f
C147 VTAIL.t10 VSUBS 0.842413f
C148 VTAIL.n17 VSUBS 1.53772f
C149 VTAIL.t14 VSUBS 0.109142f
C150 VTAIL.t19 VSUBS 0.109142f
C151 VTAIL.n18 VSUBS 0.601598f
C152 VTAIL.n19 VSUBS 0.620354f
C153 VDD2.t2 VSUBS 0.77564f
C154 VDD2.t1 VSUBS 0.090368f
C155 VDD2.t6 VSUBS 0.090368f
C156 VDD2.n0 VSUBS 0.566671f
C157 VDD2.n1 VSUBS 0.980223f
C158 VDD2.t5 VSUBS 0.090368f
C159 VDD2.t4 VSUBS 0.090368f
C160 VDD2.n2 VSUBS 0.57186f
C161 VDD2.n3 VSUBS 1.81466f
C162 VDD2.t8 VSUBS 0.769182f
C163 VDD2.n4 VSUBS 2.04002f
C164 VDD2.t9 VSUBS 0.090368f
C165 VDD2.t0 VSUBS 0.090368f
C166 VDD2.n5 VSUBS 0.566673f
C167 VDD2.n6 VSUBS 0.485072f
C168 VDD2.t3 VSUBS 0.090368f
C169 VDD2.t7 VSUBS 0.090368f
C170 VDD2.n7 VSUBS 0.571837f
C171 VN.n0 VSUBS 0.049704f
C172 VN.t9 VSUBS 0.82492f
C173 VN.n1 VSUBS 0.082161f
C174 VN.n2 VSUBS 0.049704f
C175 VN.t5 VSUBS 0.82492f
C176 VN.n3 VSUBS 0.386956f
C177 VN.n4 VSUBS 0.049704f
C178 VN.t1 VSUBS 0.82492f
C179 VN.n5 VSUBS 0.407534f
C180 VN.t2 VSUBS 0.939479f
C181 VN.n6 VSUBS 0.447034f
C182 VN.n7 VSUBS 0.260067f
C183 VN.n8 VSUBS 0.05668f
C184 VN.n9 VSUBS 0.064689f
C185 VN.n10 VSUBS 0.079816f
C186 VN.n11 VSUBS 0.049704f
C187 VN.n12 VSUBS 0.049704f
C188 VN.n13 VSUBS 0.049704f
C189 VN.n14 VSUBS 0.079816f
C190 VN.n15 VSUBS 0.064689f
C191 VN.t0 VSUBS 0.82492f
C192 VN.n16 VSUBS 0.340287f
C193 VN.n17 VSUBS 0.05668f
C194 VN.n18 VSUBS 0.049704f
C195 VN.n19 VSUBS 0.049704f
C196 VN.n20 VSUBS 0.049704f
C197 VN.n21 VSUBS 0.044919f
C198 VN.n22 VSUBS 0.074105f
C199 VN.n23 VSUBS 0.425209f
C200 VN.n24 VSUBS 0.045769f
C201 VN.n25 VSUBS 0.049704f
C202 VN.t7 VSUBS 0.82492f
C203 VN.n26 VSUBS 0.082161f
C204 VN.n27 VSUBS 0.049704f
C205 VN.t8 VSUBS 0.82492f
C206 VN.n28 VSUBS 0.340287f
C207 VN.t3 VSUBS 0.82492f
C208 VN.n29 VSUBS 0.386956f
C209 VN.n30 VSUBS 0.049704f
C210 VN.t4 VSUBS 0.82492f
C211 VN.n31 VSUBS 0.407534f
C212 VN.t6 VSUBS 0.939479f
C213 VN.n32 VSUBS 0.447034f
C214 VN.n33 VSUBS 0.260067f
C215 VN.n34 VSUBS 0.05668f
C216 VN.n35 VSUBS 0.064689f
C217 VN.n36 VSUBS 0.079816f
C218 VN.n37 VSUBS 0.049704f
C219 VN.n38 VSUBS 0.049704f
C220 VN.n39 VSUBS 0.049704f
C221 VN.n40 VSUBS 0.079816f
C222 VN.n41 VSUBS 0.064689f
C223 VN.n42 VSUBS 0.05668f
C224 VN.n43 VSUBS 0.049704f
C225 VN.n44 VSUBS 0.049704f
C226 VN.n45 VSUBS 0.049704f
C227 VN.n46 VSUBS 0.044919f
C228 VN.n47 VSUBS 0.074105f
C229 VN.n48 VSUBS 0.425209f
C230 VN.n49 VSUBS 1.9685f
C231 B.n0 VSUBS 0.005937f
C232 B.n1 VSUBS 0.005937f
C233 B.n2 VSUBS 0.00878f
C234 B.n3 VSUBS 0.006729f
C235 B.n4 VSUBS 0.006729f
C236 B.n5 VSUBS 0.006729f
C237 B.n6 VSUBS 0.006729f
C238 B.n7 VSUBS 0.006729f
C239 B.n8 VSUBS 0.006729f
C240 B.n9 VSUBS 0.006729f
C241 B.n10 VSUBS 0.006729f
C242 B.n11 VSUBS 0.006729f
C243 B.n12 VSUBS 0.006729f
C244 B.n13 VSUBS 0.006729f
C245 B.n14 VSUBS 0.006729f
C246 B.n15 VSUBS 0.006729f
C247 B.n16 VSUBS 0.006729f
C248 B.n17 VSUBS 0.006729f
C249 B.n18 VSUBS 0.006729f
C250 B.n19 VSUBS 0.006729f
C251 B.n20 VSUBS 0.016671f
C252 B.n21 VSUBS 0.006729f
C253 B.n22 VSUBS 0.006729f
C254 B.n23 VSUBS 0.006729f
C255 B.n24 VSUBS 0.006729f
C256 B.n25 VSUBS 0.006729f
C257 B.n26 VSUBS 0.006729f
C258 B.n27 VSUBS 0.006729f
C259 B.n28 VSUBS 0.006729f
C260 B.n29 VSUBS 0.006729f
C261 B.n30 VSUBS 0.004651f
C262 B.n31 VSUBS 0.006729f
C263 B.t10 VSUBS 0.13282f
C264 B.t11 VSUBS 0.143788f
C265 B.t9 VSUBS 0.280111f
C266 B.n32 VSUBS 0.086016f
C267 B.n33 VSUBS 0.062172f
C268 B.n34 VSUBS 0.015589f
C269 B.n35 VSUBS 0.006729f
C270 B.n36 VSUBS 0.006729f
C271 B.n37 VSUBS 0.006729f
C272 B.n38 VSUBS 0.006729f
C273 B.t1 VSUBS 0.13282f
C274 B.t2 VSUBS 0.143788f
C275 B.t0 VSUBS 0.280111f
C276 B.n39 VSUBS 0.086016f
C277 B.n40 VSUBS 0.062172f
C278 B.n41 VSUBS 0.006729f
C279 B.n42 VSUBS 0.006729f
C280 B.n43 VSUBS 0.006729f
C281 B.n44 VSUBS 0.006729f
C282 B.n45 VSUBS 0.006729f
C283 B.n46 VSUBS 0.006729f
C284 B.n47 VSUBS 0.006729f
C285 B.n48 VSUBS 0.006729f
C286 B.n49 VSUBS 0.006729f
C287 B.n50 VSUBS 0.016671f
C288 B.n51 VSUBS 0.006729f
C289 B.n52 VSUBS 0.006729f
C290 B.n53 VSUBS 0.006729f
C291 B.n54 VSUBS 0.006729f
C292 B.n55 VSUBS 0.006729f
C293 B.n56 VSUBS 0.006729f
C294 B.n57 VSUBS 0.006729f
C295 B.n58 VSUBS 0.006729f
C296 B.n59 VSUBS 0.006729f
C297 B.n60 VSUBS 0.006729f
C298 B.n61 VSUBS 0.006729f
C299 B.n62 VSUBS 0.006729f
C300 B.n63 VSUBS 0.006729f
C301 B.n64 VSUBS 0.006729f
C302 B.n65 VSUBS 0.006729f
C303 B.n66 VSUBS 0.006729f
C304 B.n67 VSUBS 0.006729f
C305 B.n68 VSUBS 0.006729f
C306 B.n69 VSUBS 0.006729f
C307 B.n70 VSUBS 0.006729f
C308 B.n71 VSUBS 0.006729f
C309 B.n72 VSUBS 0.006729f
C310 B.n73 VSUBS 0.006729f
C311 B.n74 VSUBS 0.006729f
C312 B.n75 VSUBS 0.006729f
C313 B.n76 VSUBS 0.006729f
C314 B.n77 VSUBS 0.006729f
C315 B.n78 VSUBS 0.006729f
C316 B.n79 VSUBS 0.006729f
C317 B.n80 VSUBS 0.006729f
C318 B.n81 VSUBS 0.006729f
C319 B.n82 VSUBS 0.006729f
C320 B.n83 VSUBS 0.006729f
C321 B.n84 VSUBS 0.006729f
C322 B.n85 VSUBS 0.006729f
C323 B.n86 VSUBS 0.006729f
C324 B.n87 VSUBS 0.016926f
C325 B.n88 VSUBS 0.006729f
C326 B.n89 VSUBS 0.006729f
C327 B.n90 VSUBS 0.006729f
C328 B.n91 VSUBS 0.006729f
C329 B.n92 VSUBS 0.006729f
C330 B.n93 VSUBS 0.006729f
C331 B.n94 VSUBS 0.006729f
C332 B.n95 VSUBS 0.006729f
C333 B.n96 VSUBS 0.006729f
C334 B.n97 VSUBS 0.006729f
C335 B.n98 VSUBS 0.006729f
C336 B.t8 VSUBS 0.13282f
C337 B.t7 VSUBS 0.143788f
C338 B.t6 VSUBS 0.280111f
C339 B.n99 VSUBS 0.086016f
C340 B.n100 VSUBS 0.062172f
C341 B.n101 VSUBS 0.006729f
C342 B.n102 VSUBS 0.006729f
C343 B.n103 VSUBS 0.006729f
C344 B.n104 VSUBS 0.006729f
C345 B.t5 VSUBS 0.13282f
C346 B.t4 VSUBS 0.143788f
C347 B.t3 VSUBS 0.280111f
C348 B.n105 VSUBS 0.086016f
C349 B.n106 VSUBS 0.062172f
C350 B.n107 VSUBS 0.006729f
C351 B.n108 VSUBS 0.006729f
C352 B.n109 VSUBS 0.006729f
C353 B.n110 VSUBS 0.006729f
C354 B.n111 VSUBS 0.006729f
C355 B.n112 VSUBS 0.006729f
C356 B.n113 VSUBS 0.006729f
C357 B.n114 VSUBS 0.006729f
C358 B.n115 VSUBS 0.006729f
C359 B.n116 VSUBS 0.006729f
C360 B.n117 VSUBS 0.01618f
C361 B.n118 VSUBS 0.006729f
C362 B.n119 VSUBS 0.006729f
C363 B.n120 VSUBS 0.006729f
C364 B.n121 VSUBS 0.006729f
C365 B.n122 VSUBS 0.006729f
C366 B.n123 VSUBS 0.006729f
C367 B.n124 VSUBS 0.006729f
C368 B.n125 VSUBS 0.006729f
C369 B.n126 VSUBS 0.006729f
C370 B.n127 VSUBS 0.006729f
C371 B.n128 VSUBS 0.006729f
C372 B.n129 VSUBS 0.006729f
C373 B.n130 VSUBS 0.006729f
C374 B.n131 VSUBS 0.006729f
C375 B.n132 VSUBS 0.006729f
C376 B.n133 VSUBS 0.006729f
C377 B.n134 VSUBS 0.006729f
C378 B.n135 VSUBS 0.006729f
C379 B.n136 VSUBS 0.006729f
C380 B.n137 VSUBS 0.006729f
C381 B.n138 VSUBS 0.006729f
C382 B.n139 VSUBS 0.006729f
C383 B.n140 VSUBS 0.006729f
C384 B.n141 VSUBS 0.006729f
C385 B.n142 VSUBS 0.006729f
C386 B.n143 VSUBS 0.006729f
C387 B.n144 VSUBS 0.006729f
C388 B.n145 VSUBS 0.006729f
C389 B.n146 VSUBS 0.006729f
C390 B.n147 VSUBS 0.006729f
C391 B.n148 VSUBS 0.006729f
C392 B.n149 VSUBS 0.006729f
C393 B.n150 VSUBS 0.006729f
C394 B.n151 VSUBS 0.006729f
C395 B.n152 VSUBS 0.006729f
C396 B.n153 VSUBS 0.006729f
C397 B.n154 VSUBS 0.006729f
C398 B.n155 VSUBS 0.006729f
C399 B.n156 VSUBS 0.006729f
C400 B.n157 VSUBS 0.006729f
C401 B.n158 VSUBS 0.006729f
C402 B.n159 VSUBS 0.006729f
C403 B.n160 VSUBS 0.006729f
C404 B.n161 VSUBS 0.006729f
C405 B.n162 VSUBS 0.006729f
C406 B.n163 VSUBS 0.006729f
C407 B.n164 VSUBS 0.006729f
C408 B.n165 VSUBS 0.006729f
C409 B.n166 VSUBS 0.006729f
C410 B.n167 VSUBS 0.006729f
C411 B.n168 VSUBS 0.006729f
C412 B.n169 VSUBS 0.006729f
C413 B.n170 VSUBS 0.006729f
C414 B.n171 VSUBS 0.006729f
C415 B.n172 VSUBS 0.006729f
C416 B.n173 VSUBS 0.006729f
C417 B.n174 VSUBS 0.006729f
C418 B.n175 VSUBS 0.006729f
C419 B.n176 VSUBS 0.006729f
C420 B.n177 VSUBS 0.006729f
C421 B.n178 VSUBS 0.006729f
C422 B.n179 VSUBS 0.006729f
C423 B.n180 VSUBS 0.006729f
C424 B.n181 VSUBS 0.006729f
C425 B.n182 VSUBS 0.006729f
C426 B.n183 VSUBS 0.006729f
C427 B.n184 VSUBS 0.006729f
C428 B.n185 VSUBS 0.006729f
C429 B.n186 VSUBS 0.01618f
C430 B.n187 VSUBS 0.016671f
C431 B.n188 VSUBS 0.016671f
C432 B.n189 VSUBS 0.006729f
C433 B.n190 VSUBS 0.006729f
C434 B.n191 VSUBS 0.006729f
C435 B.n192 VSUBS 0.006729f
C436 B.n193 VSUBS 0.006729f
C437 B.n194 VSUBS 0.006729f
C438 B.n195 VSUBS 0.006729f
C439 B.n196 VSUBS 0.006729f
C440 B.n197 VSUBS 0.006729f
C441 B.n198 VSUBS 0.006729f
C442 B.n199 VSUBS 0.006729f
C443 B.n200 VSUBS 0.006729f
C444 B.n201 VSUBS 0.006729f
C445 B.n202 VSUBS 0.006729f
C446 B.n203 VSUBS 0.006729f
C447 B.n204 VSUBS 0.006729f
C448 B.n205 VSUBS 0.006729f
C449 B.n206 VSUBS 0.006729f
C450 B.n207 VSUBS 0.006729f
C451 B.n208 VSUBS 0.006729f
C452 B.n209 VSUBS 0.006729f
C453 B.n210 VSUBS 0.006729f
C454 B.n211 VSUBS 0.006729f
C455 B.n212 VSUBS 0.006729f
C456 B.n213 VSUBS 0.006729f
C457 B.n214 VSUBS 0.006729f
C458 B.n215 VSUBS 0.006729f
C459 B.n216 VSUBS 0.006729f
C460 B.n217 VSUBS 0.006729f
C461 B.n218 VSUBS 0.004651f
C462 B.n219 VSUBS 0.015589f
C463 B.n220 VSUBS 0.005442f
C464 B.n221 VSUBS 0.006729f
C465 B.n222 VSUBS 0.006729f
C466 B.n223 VSUBS 0.006729f
C467 B.n224 VSUBS 0.006729f
C468 B.n225 VSUBS 0.006729f
C469 B.n226 VSUBS 0.006729f
C470 B.n227 VSUBS 0.006729f
C471 B.n228 VSUBS 0.006729f
C472 B.n229 VSUBS 0.006729f
C473 B.n230 VSUBS 0.006729f
C474 B.n231 VSUBS 0.006729f
C475 B.n232 VSUBS 0.005442f
C476 B.n233 VSUBS 0.015589f
C477 B.n234 VSUBS 0.004651f
C478 B.n235 VSUBS 0.006729f
C479 B.n236 VSUBS 0.006729f
C480 B.n237 VSUBS 0.006729f
C481 B.n238 VSUBS 0.006729f
C482 B.n239 VSUBS 0.006729f
C483 B.n240 VSUBS 0.006729f
C484 B.n241 VSUBS 0.006729f
C485 B.n242 VSUBS 0.006729f
C486 B.n243 VSUBS 0.006729f
C487 B.n244 VSUBS 0.006729f
C488 B.n245 VSUBS 0.006729f
C489 B.n246 VSUBS 0.006729f
C490 B.n247 VSUBS 0.006729f
C491 B.n248 VSUBS 0.006729f
C492 B.n249 VSUBS 0.006729f
C493 B.n250 VSUBS 0.006729f
C494 B.n251 VSUBS 0.006729f
C495 B.n252 VSUBS 0.006729f
C496 B.n253 VSUBS 0.006729f
C497 B.n254 VSUBS 0.006729f
C498 B.n255 VSUBS 0.006729f
C499 B.n256 VSUBS 0.006729f
C500 B.n257 VSUBS 0.006729f
C501 B.n258 VSUBS 0.006729f
C502 B.n259 VSUBS 0.006729f
C503 B.n260 VSUBS 0.006729f
C504 B.n261 VSUBS 0.006729f
C505 B.n262 VSUBS 0.006729f
C506 B.n263 VSUBS 0.006729f
C507 B.n264 VSUBS 0.015925f
C508 B.n265 VSUBS 0.016671f
C509 B.n266 VSUBS 0.01618f
C510 B.n267 VSUBS 0.006729f
C511 B.n268 VSUBS 0.006729f
C512 B.n269 VSUBS 0.006729f
C513 B.n270 VSUBS 0.006729f
C514 B.n271 VSUBS 0.006729f
C515 B.n272 VSUBS 0.006729f
C516 B.n273 VSUBS 0.006729f
C517 B.n274 VSUBS 0.006729f
C518 B.n275 VSUBS 0.006729f
C519 B.n276 VSUBS 0.006729f
C520 B.n277 VSUBS 0.006729f
C521 B.n278 VSUBS 0.006729f
C522 B.n279 VSUBS 0.006729f
C523 B.n280 VSUBS 0.006729f
C524 B.n281 VSUBS 0.006729f
C525 B.n282 VSUBS 0.006729f
C526 B.n283 VSUBS 0.006729f
C527 B.n284 VSUBS 0.006729f
C528 B.n285 VSUBS 0.006729f
C529 B.n286 VSUBS 0.006729f
C530 B.n287 VSUBS 0.006729f
C531 B.n288 VSUBS 0.006729f
C532 B.n289 VSUBS 0.006729f
C533 B.n290 VSUBS 0.006729f
C534 B.n291 VSUBS 0.006729f
C535 B.n292 VSUBS 0.006729f
C536 B.n293 VSUBS 0.006729f
C537 B.n294 VSUBS 0.006729f
C538 B.n295 VSUBS 0.006729f
C539 B.n296 VSUBS 0.006729f
C540 B.n297 VSUBS 0.006729f
C541 B.n298 VSUBS 0.006729f
C542 B.n299 VSUBS 0.006729f
C543 B.n300 VSUBS 0.006729f
C544 B.n301 VSUBS 0.006729f
C545 B.n302 VSUBS 0.006729f
C546 B.n303 VSUBS 0.006729f
C547 B.n304 VSUBS 0.006729f
C548 B.n305 VSUBS 0.006729f
C549 B.n306 VSUBS 0.006729f
C550 B.n307 VSUBS 0.006729f
C551 B.n308 VSUBS 0.006729f
C552 B.n309 VSUBS 0.006729f
C553 B.n310 VSUBS 0.006729f
C554 B.n311 VSUBS 0.006729f
C555 B.n312 VSUBS 0.006729f
C556 B.n313 VSUBS 0.006729f
C557 B.n314 VSUBS 0.006729f
C558 B.n315 VSUBS 0.006729f
C559 B.n316 VSUBS 0.006729f
C560 B.n317 VSUBS 0.006729f
C561 B.n318 VSUBS 0.006729f
C562 B.n319 VSUBS 0.006729f
C563 B.n320 VSUBS 0.006729f
C564 B.n321 VSUBS 0.006729f
C565 B.n322 VSUBS 0.006729f
C566 B.n323 VSUBS 0.006729f
C567 B.n324 VSUBS 0.006729f
C568 B.n325 VSUBS 0.006729f
C569 B.n326 VSUBS 0.006729f
C570 B.n327 VSUBS 0.006729f
C571 B.n328 VSUBS 0.006729f
C572 B.n329 VSUBS 0.006729f
C573 B.n330 VSUBS 0.006729f
C574 B.n331 VSUBS 0.006729f
C575 B.n332 VSUBS 0.006729f
C576 B.n333 VSUBS 0.006729f
C577 B.n334 VSUBS 0.006729f
C578 B.n335 VSUBS 0.006729f
C579 B.n336 VSUBS 0.006729f
C580 B.n337 VSUBS 0.006729f
C581 B.n338 VSUBS 0.006729f
C582 B.n339 VSUBS 0.006729f
C583 B.n340 VSUBS 0.006729f
C584 B.n341 VSUBS 0.006729f
C585 B.n342 VSUBS 0.006729f
C586 B.n343 VSUBS 0.006729f
C587 B.n344 VSUBS 0.006729f
C588 B.n345 VSUBS 0.006729f
C589 B.n346 VSUBS 0.006729f
C590 B.n347 VSUBS 0.006729f
C591 B.n348 VSUBS 0.006729f
C592 B.n349 VSUBS 0.006729f
C593 B.n350 VSUBS 0.006729f
C594 B.n351 VSUBS 0.006729f
C595 B.n352 VSUBS 0.006729f
C596 B.n353 VSUBS 0.006729f
C597 B.n354 VSUBS 0.006729f
C598 B.n355 VSUBS 0.006729f
C599 B.n356 VSUBS 0.006729f
C600 B.n357 VSUBS 0.006729f
C601 B.n358 VSUBS 0.006729f
C602 B.n359 VSUBS 0.006729f
C603 B.n360 VSUBS 0.006729f
C604 B.n361 VSUBS 0.006729f
C605 B.n362 VSUBS 0.006729f
C606 B.n363 VSUBS 0.006729f
C607 B.n364 VSUBS 0.006729f
C608 B.n365 VSUBS 0.006729f
C609 B.n366 VSUBS 0.006729f
C610 B.n367 VSUBS 0.006729f
C611 B.n368 VSUBS 0.006729f
C612 B.n369 VSUBS 0.006729f
C613 B.n370 VSUBS 0.006729f
C614 B.n371 VSUBS 0.006729f
C615 B.n372 VSUBS 0.006729f
C616 B.n373 VSUBS 0.006729f
C617 B.n374 VSUBS 0.006729f
C618 B.n375 VSUBS 0.01618f
C619 B.n376 VSUBS 0.01618f
C620 B.n377 VSUBS 0.016671f
C621 B.n378 VSUBS 0.006729f
C622 B.n379 VSUBS 0.006729f
C623 B.n380 VSUBS 0.006729f
C624 B.n381 VSUBS 0.006729f
C625 B.n382 VSUBS 0.006729f
C626 B.n383 VSUBS 0.006729f
C627 B.n384 VSUBS 0.006729f
C628 B.n385 VSUBS 0.006729f
C629 B.n386 VSUBS 0.006729f
C630 B.n387 VSUBS 0.006729f
C631 B.n388 VSUBS 0.006729f
C632 B.n389 VSUBS 0.006729f
C633 B.n390 VSUBS 0.006729f
C634 B.n391 VSUBS 0.006729f
C635 B.n392 VSUBS 0.006729f
C636 B.n393 VSUBS 0.006729f
C637 B.n394 VSUBS 0.006729f
C638 B.n395 VSUBS 0.006729f
C639 B.n396 VSUBS 0.006729f
C640 B.n397 VSUBS 0.006729f
C641 B.n398 VSUBS 0.006729f
C642 B.n399 VSUBS 0.006729f
C643 B.n400 VSUBS 0.006729f
C644 B.n401 VSUBS 0.006729f
C645 B.n402 VSUBS 0.006729f
C646 B.n403 VSUBS 0.006729f
C647 B.n404 VSUBS 0.006729f
C648 B.n405 VSUBS 0.006729f
C649 B.n406 VSUBS 0.006729f
C650 B.n407 VSUBS 0.004651f
C651 B.n408 VSUBS 0.015589f
C652 B.n409 VSUBS 0.005442f
C653 B.n410 VSUBS 0.006729f
C654 B.n411 VSUBS 0.006729f
C655 B.n412 VSUBS 0.006729f
C656 B.n413 VSUBS 0.006729f
C657 B.n414 VSUBS 0.006729f
C658 B.n415 VSUBS 0.006729f
C659 B.n416 VSUBS 0.006729f
C660 B.n417 VSUBS 0.006729f
C661 B.n418 VSUBS 0.006729f
C662 B.n419 VSUBS 0.006729f
C663 B.n420 VSUBS 0.006729f
C664 B.n421 VSUBS 0.005442f
C665 B.n422 VSUBS 0.006729f
C666 B.n423 VSUBS 0.006729f
C667 B.n424 VSUBS 0.006729f
C668 B.n425 VSUBS 0.006729f
C669 B.n426 VSUBS 0.006729f
C670 B.n427 VSUBS 0.006729f
C671 B.n428 VSUBS 0.006729f
C672 B.n429 VSUBS 0.006729f
C673 B.n430 VSUBS 0.006729f
C674 B.n431 VSUBS 0.006729f
C675 B.n432 VSUBS 0.006729f
C676 B.n433 VSUBS 0.006729f
C677 B.n434 VSUBS 0.006729f
C678 B.n435 VSUBS 0.006729f
C679 B.n436 VSUBS 0.006729f
C680 B.n437 VSUBS 0.006729f
C681 B.n438 VSUBS 0.006729f
C682 B.n439 VSUBS 0.006729f
C683 B.n440 VSUBS 0.006729f
C684 B.n441 VSUBS 0.006729f
C685 B.n442 VSUBS 0.006729f
C686 B.n443 VSUBS 0.006729f
C687 B.n444 VSUBS 0.006729f
C688 B.n445 VSUBS 0.006729f
C689 B.n446 VSUBS 0.006729f
C690 B.n447 VSUBS 0.006729f
C691 B.n448 VSUBS 0.006729f
C692 B.n449 VSUBS 0.006729f
C693 B.n450 VSUBS 0.006729f
C694 B.n451 VSUBS 0.006729f
C695 B.n452 VSUBS 0.006729f
C696 B.n453 VSUBS 0.016671f
C697 B.n454 VSUBS 0.01618f
C698 B.n455 VSUBS 0.01618f
C699 B.n456 VSUBS 0.006729f
C700 B.n457 VSUBS 0.006729f
C701 B.n458 VSUBS 0.006729f
C702 B.n459 VSUBS 0.006729f
C703 B.n460 VSUBS 0.006729f
C704 B.n461 VSUBS 0.006729f
C705 B.n462 VSUBS 0.006729f
C706 B.n463 VSUBS 0.006729f
C707 B.n464 VSUBS 0.006729f
C708 B.n465 VSUBS 0.006729f
C709 B.n466 VSUBS 0.006729f
C710 B.n467 VSUBS 0.006729f
C711 B.n468 VSUBS 0.006729f
C712 B.n469 VSUBS 0.006729f
C713 B.n470 VSUBS 0.006729f
C714 B.n471 VSUBS 0.006729f
C715 B.n472 VSUBS 0.006729f
C716 B.n473 VSUBS 0.006729f
C717 B.n474 VSUBS 0.006729f
C718 B.n475 VSUBS 0.006729f
C719 B.n476 VSUBS 0.006729f
C720 B.n477 VSUBS 0.006729f
C721 B.n478 VSUBS 0.006729f
C722 B.n479 VSUBS 0.006729f
C723 B.n480 VSUBS 0.006729f
C724 B.n481 VSUBS 0.006729f
C725 B.n482 VSUBS 0.006729f
C726 B.n483 VSUBS 0.006729f
C727 B.n484 VSUBS 0.006729f
C728 B.n485 VSUBS 0.006729f
C729 B.n486 VSUBS 0.006729f
C730 B.n487 VSUBS 0.006729f
C731 B.n488 VSUBS 0.006729f
C732 B.n489 VSUBS 0.006729f
C733 B.n490 VSUBS 0.006729f
C734 B.n491 VSUBS 0.006729f
C735 B.n492 VSUBS 0.006729f
C736 B.n493 VSUBS 0.006729f
C737 B.n494 VSUBS 0.006729f
C738 B.n495 VSUBS 0.006729f
C739 B.n496 VSUBS 0.006729f
C740 B.n497 VSUBS 0.006729f
C741 B.n498 VSUBS 0.006729f
C742 B.n499 VSUBS 0.006729f
C743 B.n500 VSUBS 0.006729f
C744 B.n501 VSUBS 0.006729f
C745 B.n502 VSUBS 0.006729f
C746 B.n503 VSUBS 0.006729f
C747 B.n504 VSUBS 0.006729f
C748 B.n505 VSUBS 0.006729f
C749 B.n506 VSUBS 0.006729f
C750 B.n507 VSUBS 0.00878f
C751 B.n508 VSUBS 0.009353f
C752 B.n509 VSUBS 0.0186f
.ends

