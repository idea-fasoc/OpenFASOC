* NGSPICE file created from diff_pair_sample_1251.ext - technology: sky130A

.subckt diff_pair_sample_1251 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=0 ps=0 w=14.6 l=3.85
X1 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=0 ps=0 w=14.6 l=3.85
X2 VDD1.t7 VP.t0 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=5.694 ps=29.98 w=14.6 l=3.85
X3 VTAIL.t9 VP.t1 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=3.85
X4 VTAIL.t10 VP.t2 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=2.409 ps=14.93 w=14.6 l=3.85
X5 VTAIL.t11 VP.t3 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=3.85
X6 VTAIL.t3 VN.t0 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=2.409 ps=14.93 w=14.6 l=3.85
X7 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=0 ps=0 w=14.6 l=3.85
X8 VDD1.t3 VP.t4 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=5.694 ps=29.98 w=14.6 l=3.85
X9 VTAIL.t2 VN.t1 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=3.85
X10 VDD2.t5 VN.t2 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=3.85
X11 VDD2.t4 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=5.694 ps=29.98 w=14.6 l=3.85
X12 VDD1.t2 VP.t5 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=3.85
X13 VDD2.t3 VN.t4 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=3.85
X14 VTAIL.t0 VN.t5 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=2.409 ps=14.93 w=14.6 l=3.85
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=0 ps=0 w=14.6 l=3.85
X16 VTAIL.t14 VP.t6 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.694 pd=29.98 as=2.409 ps=14.93 w=14.6 l=3.85
X17 VDD2.t1 VN.t6 VTAIL.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=5.694 ps=29.98 w=14.6 l=3.85
X18 VTAIL.t4 VN.t7 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=3.85
X19 VDD1.t0 VP.t7 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.409 pd=14.93 as=2.409 ps=14.93 w=14.6 l=3.85
R0 B.n1108 B.n1107 585
R1 B.n399 B.n180 585
R2 B.n398 B.n397 585
R3 B.n396 B.n395 585
R4 B.n394 B.n393 585
R5 B.n392 B.n391 585
R6 B.n390 B.n389 585
R7 B.n388 B.n387 585
R8 B.n386 B.n385 585
R9 B.n384 B.n383 585
R10 B.n382 B.n381 585
R11 B.n380 B.n379 585
R12 B.n378 B.n377 585
R13 B.n376 B.n375 585
R14 B.n374 B.n373 585
R15 B.n372 B.n371 585
R16 B.n370 B.n369 585
R17 B.n368 B.n367 585
R18 B.n366 B.n365 585
R19 B.n364 B.n363 585
R20 B.n362 B.n361 585
R21 B.n360 B.n359 585
R22 B.n358 B.n357 585
R23 B.n356 B.n355 585
R24 B.n354 B.n353 585
R25 B.n352 B.n351 585
R26 B.n350 B.n349 585
R27 B.n348 B.n347 585
R28 B.n346 B.n345 585
R29 B.n344 B.n343 585
R30 B.n342 B.n341 585
R31 B.n340 B.n339 585
R32 B.n338 B.n337 585
R33 B.n336 B.n335 585
R34 B.n334 B.n333 585
R35 B.n332 B.n331 585
R36 B.n330 B.n329 585
R37 B.n328 B.n327 585
R38 B.n326 B.n325 585
R39 B.n324 B.n323 585
R40 B.n322 B.n321 585
R41 B.n320 B.n319 585
R42 B.n318 B.n317 585
R43 B.n316 B.n315 585
R44 B.n314 B.n313 585
R45 B.n312 B.n311 585
R46 B.n310 B.n309 585
R47 B.n308 B.n307 585
R48 B.n306 B.n305 585
R49 B.n303 B.n302 585
R50 B.n301 B.n300 585
R51 B.n299 B.n298 585
R52 B.n297 B.n296 585
R53 B.n295 B.n294 585
R54 B.n293 B.n292 585
R55 B.n291 B.n290 585
R56 B.n289 B.n288 585
R57 B.n287 B.n286 585
R58 B.n285 B.n284 585
R59 B.n282 B.n281 585
R60 B.n280 B.n279 585
R61 B.n278 B.n277 585
R62 B.n276 B.n275 585
R63 B.n274 B.n273 585
R64 B.n272 B.n271 585
R65 B.n270 B.n269 585
R66 B.n268 B.n267 585
R67 B.n266 B.n265 585
R68 B.n264 B.n263 585
R69 B.n262 B.n261 585
R70 B.n260 B.n259 585
R71 B.n258 B.n257 585
R72 B.n256 B.n255 585
R73 B.n254 B.n253 585
R74 B.n252 B.n251 585
R75 B.n250 B.n249 585
R76 B.n248 B.n247 585
R77 B.n246 B.n245 585
R78 B.n244 B.n243 585
R79 B.n242 B.n241 585
R80 B.n240 B.n239 585
R81 B.n238 B.n237 585
R82 B.n236 B.n235 585
R83 B.n234 B.n233 585
R84 B.n232 B.n231 585
R85 B.n230 B.n229 585
R86 B.n228 B.n227 585
R87 B.n226 B.n225 585
R88 B.n224 B.n223 585
R89 B.n222 B.n221 585
R90 B.n220 B.n219 585
R91 B.n218 B.n217 585
R92 B.n216 B.n215 585
R93 B.n214 B.n213 585
R94 B.n212 B.n211 585
R95 B.n210 B.n209 585
R96 B.n208 B.n207 585
R97 B.n206 B.n205 585
R98 B.n204 B.n203 585
R99 B.n202 B.n201 585
R100 B.n200 B.n199 585
R101 B.n198 B.n197 585
R102 B.n196 B.n195 585
R103 B.n194 B.n193 585
R104 B.n192 B.n191 585
R105 B.n190 B.n189 585
R106 B.n188 B.n187 585
R107 B.n186 B.n185 585
R108 B.n1106 B.n126 585
R109 B.n1111 B.n126 585
R110 B.n1105 B.n125 585
R111 B.n1112 B.n125 585
R112 B.n1104 B.n1103 585
R113 B.n1103 B.n121 585
R114 B.n1102 B.n120 585
R115 B.n1118 B.n120 585
R116 B.n1101 B.n119 585
R117 B.n1119 B.n119 585
R118 B.n1100 B.n118 585
R119 B.n1120 B.n118 585
R120 B.n1099 B.n1098 585
R121 B.n1098 B.n114 585
R122 B.n1097 B.n113 585
R123 B.n1126 B.n113 585
R124 B.n1096 B.n112 585
R125 B.n1127 B.n112 585
R126 B.n1095 B.n111 585
R127 B.n1128 B.n111 585
R128 B.n1094 B.n1093 585
R129 B.n1093 B.n107 585
R130 B.n1092 B.n106 585
R131 B.n1134 B.n106 585
R132 B.n1091 B.n105 585
R133 B.n1135 B.n105 585
R134 B.n1090 B.n104 585
R135 B.n1136 B.n104 585
R136 B.n1089 B.n1088 585
R137 B.n1088 B.n100 585
R138 B.n1087 B.n99 585
R139 B.n1142 B.n99 585
R140 B.n1086 B.n98 585
R141 B.n1143 B.n98 585
R142 B.n1085 B.n97 585
R143 B.n1144 B.n97 585
R144 B.n1084 B.n1083 585
R145 B.n1083 B.n93 585
R146 B.n1082 B.n92 585
R147 B.n1150 B.n92 585
R148 B.n1081 B.n91 585
R149 B.n1151 B.n91 585
R150 B.n1080 B.n90 585
R151 B.n1152 B.n90 585
R152 B.n1079 B.n1078 585
R153 B.n1078 B.n86 585
R154 B.n1077 B.n85 585
R155 B.n1158 B.n85 585
R156 B.n1076 B.n84 585
R157 B.n1159 B.n84 585
R158 B.n1075 B.n83 585
R159 B.n1160 B.n83 585
R160 B.n1074 B.n1073 585
R161 B.n1073 B.n79 585
R162 B.n1072 B.n78 585
R163 B.n1166 B.n78 585
R164 B.n1071 B.n77 585
R165 B.n1167 B.n77 585
R166 B.n1070 B.n76 585
R167 B.n1168 B.n76 585
R168 B.n1069 B.n1068 585
R169 B.n1068 B.n72 585
R170 B.n1067 B.n71 585
R171 B.n1174 B.n71 585
R172 B.n1066 B.n70 585
R173 B.n1175 B.n70 585
R174 B.n1065 B.n69 585
R175 B.n1176 B.n69 585
R176 B.n1064 B.n1063 585
R177 B.n1063 B.n65 585
R178 B.n1062 B.n64 585
R179 B.n1182 B.n64 585
R180 B.n1061 B.n63 585
R181 B.n1183 B.n63 585
R182 B.n1060 B.n62 585
R183 B.n1184 B.n62 585
R184 B.n1059 B.n1058 585
R185 B.n1058 B.n58 585
R186 B.n1057 B.n57 585
R187 B.n1190 B.n57 585
R188 B.n1056 B.n56 585
R189 B.n1191 B.n56 585
R190 B.n1055 B.n55 585
R191 B.n1192 B.n55 585
R192 B.n1054 B.n1053 585
R193 B.n1053 B.n51 585
R194 B.n1052 B.n50 585
R195 B.n1198 B.n50 585
R196 B.n1051 B.n49 585
R197 B.n1199 B.n49 585
R198 B.n1050 B.n48 585
R199 B.n1200 B.n48 585
R200 B.n1049 B.n1048 585
R201 B.n1048 B.n44 585
R202 B.n1047 B.n43 585
R203 B.n1206 B.n43 585
R204 B.n1046 B.n42 585
R205 B.n1207 B.n42 585
R206 B.n1045 B.n41 585
R207 B.n1208 B.n41 585
R208 B.n1044 B.n1043 585
R209 B.n1043 B.n37 585
R210 B.n1042 B.n36 585
R211 B.n1214 B.n36 585
R212 B.n1041 B.n35 585
R213 B.n1215 B.n35 585
R214 B.n1040 B.n34 585
R215 B.n1216 B.n34 585
R216 B.n1039 B.n1038 585
R217 B.n1038 B.n30 585
R218 B.n1037 B.n29 585
R219 B.n1222 B.n29 585
R220 B.n1036 B.n28 585
R221 B.n1223 B.n28 585
R222 B.n1035 B.n27 585
R223 B.n1224 B.n27 585
R224 B.n1034 B.n1033 585
R225 B.n1033 B.n23 585
R226 B.n1032 B.n22 585
R227 B.n1230 B.n22 585
R228 B.n1031 B.n21 585
R229 B.n1231 B.n21 585
R230 B.n1030 B.n20 585
R231 B.n1232 B.n20 585
R232 B.n1029 B.n1028 585
R233 B.n1028 B.n16 585
R234 B.n1027 B.n15 585
R235 B.n1238 B.n15 585
R236 B.n1026 B.n14 585
R237 B.n1239 B.n14 585
R238 B.n1025 B.n13 585
R239 B.n1240 B.n13 585
R240 B.n1024 B.n1023 585
R241 B.n1023 B.n12 585
R242 B.n1022 B.n1021 585
R243 B.n1022 B.n8 585
R244 B.n1020 B.n7 585
R245 B.n1247 B.n7 585
R246 B.n1019 B.n6 585
R247 B.n1248 B.n6 585
R248 B.n1018 B.n5 585
R249 B.n1249 B.n5 585
R250 B.n1017 B.n1016 585
R251 B.n1016 B.n4 585
R252 B.n1015 B.n400 585
R253 B.n1015 B.n1014 585
R254 B.n1005 B.n401 585
R255 B.n402 B.n401 585
R256 B.n1007 B.n1006 585
R257 B.n1008 B.n1007 585
R258 B.n1004 B.n407 585
R259 B.n407 B.n406 585
R260 B.n1003 B.n1002 585
R261 B.n1002 B.n1001 585
R262 B.n409 B.n408 585
R263 B.n410 B.n409 585
R264 B.n994 B.n993 585
R265 B.n995 B.n994 585
R266 B.n992 B.n415 585
R267 B.n415 B.n414 585
R268 B.n991 B.n990 585
R269 B.n990 B.n989 585
R270 B.n417 B.n416 585
R271 B.n418 B.n417 585
R272 B.n982 B.n981 585
R273 B.n983 B.n982 585
R274 B.n980 B.n423 585
R275 B.n423 B.n422 585
R276 B.n979 B.n978 585
R277 B.n978 B.n977 585
R278 B.n425 B.n424 585
R279 B.n426 B.n425 585
R280 B.n970 B.n969 585
R281 B.n971 B.n970 585
R282 B.n968 B.n431 585
R283 B.n431 B.n430 585
R284 B.n967 B.n966 585
R285 B.n966 B.n965 585
R286 B.n433 B.n432 585
R287 B.n434 B.n433 585
R288 B.n958 B.n957 585
R289 B.n959 B.n958 585
R290 B.n956 B.n439 585
R291 B.n439 B.n438 585
R292 B.n955 B.n954 585
R293 B.n954 B.n953 585
R294 B.n441 B.n440 585
R295 B.n442 B.n441 585
R296 B.n946 B.n945 585
R297 B.n947 B.n946 585
R298 B.n944 B.n447 585
R299 B.n447 B.n446 585
R300 B.n943 B.n942 585
R301 B.n942 B.n941 585
R302 B.n449 B.n448 585
R303 B.n450 B.n449 585
R304 B.n934 B.n933 585
R305 B.n935 B.n934 585
R306 B.n932 B.n455 585
R307 B.n455 B.n454 585
R308 B.n931 B.n930 585
R309 B.n930 B.n929 585
R310 B.n457 B.n456 585
R311 B.n458 B.n457 585
R312 B.n922 B.n921 585
R313 B.n923 B.n922 585
R314 B.n920 B.n463 585
R315 B.n463 B.n462 585
R316 B.n919 B.n918 585
R317 B.n918 B.n917 585
R318 B.n465 B.n464 585
R319 B.n466 B.n465 585
R320 B.n910 B.n909 585
R321 B.n911 B.n910 585
R322 B.n908 B.n471 585
R323 B.n471 B.n470 585
R324 B.n907 B.n906 585
R325 B.n906 B.n905 585
R326 B.n473 B.n472 585
R327 B.n474 B.n473 585
R328 B.n898 B.n897 585
R329 B.n899 B.n898 585
R330 B.n896 B.n479 585
R331 B.n479 B.n478 585
R332 B.n895 B.n894 585
R333 B.n894 B.n893 585
R334 B.n481 B.n480 585
R335 B.n482 B.n481 585
R336 B.n886 B.n885 585
R337 B.n887 B.n886 585
R338 B.n884 B.n486 585
R339 B.n490 B.n486 585
R340 B.n883 B.n882 585
R341 B.n882 B.n881 585
R342 B.n488 B.n487 585
R343 B.n489 B.n488 585
R344 B.n874 B.n873 585
R345 B.n875 B.n874 585
R346 B.n872 B.n495 585
R347 B.n495 B.n494 585
R348 B.n871 B.n870 585
R349 B.n870 B.n869 585
R350 B.n497 B.n496 585
R351 B.n498 B.n497 585
R352 B.n862 B.n861 585
R353 B.n863 B.n862 585
R354 B.n860 B.n503 585
R355 B.n503 B.n502 585
R356 B.n859 B.n858 585
R357 B.n858 B.n857 585
R358 B.n505 B.n504 585
R359 B.n506 B.n505 585
R360 B.n850 B.n849 585
R361 B.n851 B.n850 585
R362 B.n848 B.n511 585
R363 B.n511 B.n510 585
R364 B.n847 B.n846 585
R365 B.n846 B.n845 585
R366 B.n513 B.n512 585
R367 B.n514 B.n513 585
R368 B.n838 B.n837 585
R369 B.n839 B.n838 585
R370 B.n836 B.n519 585
R371 B.n519 B.n518 585
R372 B.n835 B.n834 585
R373 B.n834 B.n833 585
R374 B.n521 B.n520 585
R375 B.n522 B.n521 585
R376 B.n826 B.n825 585
R377 B.n827 B.n826 585
R378 B.n824 B.n527 585
R379 B.n527 B.n526 585
R380 B.n823 B.n822 585
R381 B.n822 B.n821 585
R382 B.n529 B.n528 585
R383 B.n530 B.n529 585
R384 B.n814 B.n813 585
R385 B.n815 B.n814 585
R386 B.n812 B.n535 585
R387 B.n535 B.n534 585
R388 B.n807 B.n806 585
R389 B.n805 B.n591 585
R390 B.n804 B.n590 585
R391 B.n809 B.n590 585
R392 B.n803 B.n802 585
R393 B.n801 B.n800 585
R394 B.n799 B.n798 585
R395 B.n797 B.n796 585
R396 B.n795 B.n794 585
R397 B.n793 B.n792 585
R398 B.n791 B.n790 585
R399 B.n789 B.n788 585
R400 B.n787 B.n786 585
R401 B.n785 B.n784 585
R402 B.n783 B.n782 585
R403 B.n781 B.n780 585
R404 B.n779 B.n778 585
R405 B.n777 B.n776 585
R406 B.n775 B.n774 585
R407 B.n773 B.n772 585
R408 B.n771 B.n770 585
R409 B.n769 B.n768 585
R410 B.n767 B.n766 585
R411 B.n765 B.n764 585
R412 B.n763 B.n762 585
R413 B.n761 B.n760 585
R414 B.n759 B.n758 585
R415 B.n757 B.n756 585
R416 B.n755 B.n754 585
R417 B.n753 B.n752 585
R418 B.n751 B.n750 585
R419 B.n749 B.n748 585
R420 B.n747 B.n746 585
R421 B.n745 B.n744 585
R422 B.n743 B.n742 585
R423 B.n741 B.n740 585
R424 B.n739 B.n738 585
R425 B.n737 B.n736 585
R426 B.n735 B.n734 585
R427 B.n733 B.n732 585
R428 B.n731 B.n730 585
R429 B.n729 B.n728 585
R430 B.n727 B.n726 585
R431 B.n725 B.n724 585
R432 B.n723 B.n722 585
R433 B.n721 B.n720 585
R434 B.n719 B.n718 585
R435 B.n717 B.n716 585
R436 B.n715 B.n714 585
R437 B.n713 B.n712 585
R438 B.n711 B.n710 585
R439 B.n709 B.n708 585
R440 B.n707 B.n706 585
R441 B.n705 B.n704 585
R442 B.n703 B.n702 585
R443 B.n701 B.n700 585
R444 B.n699 B.n698 585
R445 B.n697 B.n696 585
R446 B.n695 B.n694 585
R447 B.n693 B.n692 585
R448 B.n691 B.n690 585
R449 B.n689 B.n688 585
R450 B.n687 B.n686 585
R451 B.n685 B.n684 585
R452 B.n683 B.n682 585
R453 B.n681 B.n680 585
R454 B.n679 B.n678 585
R455 B.n677 B.n676 585
R456 B.n675 B.n674 585
R457 B.n673 B.n672 585
R458 B.n671 B.n670 585
R459 B.n669 B.n668 585
R460 B.n667 B.n666 585
R461 B.n665 B.n664 585
R462 B.n663 B.n662 585
R463 B.n661 B.n660 585
R464 B.n659 B.n658 585
R465 B.n657 B.n656 585
R466 B.n655 B.n654 585
R467 B.n653 B.n652 585
R468 B.n651 B.n650 585
R469 B.n649 B.n648 585
R470 B.n647 B.n646 585
R471 B.n645 B.n644 585
R472 B.n643 B.n642 585
R473 B.n641 B.n640 585
R474 B.n639 B.n638 585
R475 B.n637 B.n636 585
R476 B.n635 B.n634 585
R477 B.n633 B.n632 585
R478 B.n631 B.n630 585
R479 B.n629 B.n628 585
R480 B.n627 B.n626 585
R481 B.n625 B.n624 585
R482 B.n623 B.n622 585
R483 B.n621 B.n620 585
R484 B.n619 B.n618 585
R485 B.n617 B.n616 585
R486 B.n615 B.n614 585
R487 B.n613 B.n612 585
R488 B.n611 B.n610 585
R489 B.n609 B.n608 585
R490 B.n607 B.n606 585
R491 B.n605 B.n604 585
R492 B.n603 B.n602 585
R493 B.n601 B.n600 585
R494 B.n599 B.n598 585
R495 B.n537 B.n536 585
R496 B.n811 B.n810 585
R497 B.n810 B.n809 585
R498 B.n533 B.n532 585
R499 B.n534 B.n533 585
R500 B.n817 B.n816 585
R501 B.n816 B.n815 585
R502 B.n818 B.n531 585
R503 B.n531 B.n530 585
R504 B.n820 B.n819 585
R505 B.n821 B.n820 585
R506 B.n525 B.n524 585
R507 B.n526 B.n525 585
R508 B.n829 B.n828 585
R509 B.n828 B.n827 585
R510 B.n830 B.n523 585
R511 B.n523 B.n522 585
R512 B.n832 B.n831 585
R513 B.n833 B.n832 585
R514 B.n517 B.n516 585
R515 B.n518 B.n517 585
R516 B.n841 B.n840 585
R517 B.n840 B.n839 585
R518 B.n842 B.n515 585
R519 B.n515 B.n514 585
R520 B.n844 B.n843 585
R521 B.n845 B.n844 585
R522 B.n509 B.n508 585
R523 B.n510 B.n509 585
R524 B.n853 B.n852 585
R525 B.n852 B.n851 585
R526 B.n854 B.n507 585
R527 B.n507 B.n506 585
R528 B.n856 B.n855 585
R529 B.n857 B.n856 585
R530 B.n501 B.n500 585
R531 B.n502 B.n501 585
R532 B.n865 B.n864 585
R533 B.n864 B.n863 585
R534 B.n866 B.n499 585
R535 B.n499 B.n498 585
R536 B.n868 B.n867 585
R537 B.n869 B.n868 585
R538 B.n493 B.n492 585
R539 B.n494 B.n493 585
R540 B.n877 B.n876 585
R541 B.n876 B.n875 585
R542 B.n878 B.n491 585
R543 B.n491 B.n489 585
R544 B.n880 B.n879 585
R545 B.n881 B.n880 585
R546 B.n485 B.n484 585
R547 B.n490 B.n485 585
R548 B.n889 B.n888 585
R549 B.n888 B.n887 585
R550 B.n890 B.n483 585
R551 B.n483 B.n482 585
R552 B.n892 B.n891 585
R553 B.n893 B.n892 585
R554 B.n477 B.n476 585
R555 B.n478 B.n477 585
R556 B.n901 B.n900 585
R557 B.n900 B.n899 585
R558 B.n902 B.n475 585
R559 B.n475 B.n474 585
R560 B.n904 B.n903 585
R561 B.n905 B.n904 585
R562 B.n469 B.n468 585
R563 B.n470 B.n469 585
R564 B.n913 B.n912 585
R565 B.n912 B.n911 585
R566 B.n914 B.n467 585
R567 B.n467 B.n466 585
R568 B.n916 B.n915 585
R569 B.n917 B.n916 585
R570 B.n461 B.n460 585
R571 B.n462 B.n461 585
R572 B.n925 B.n924 585
R573 B.n924 B.n923 585
R574 B.n926 B.n459 585
R575 B.n459 B.n458 585
R576 B.n928 B.n927 585
R577 B.n929 B.n928 585
R578 B.n453 B.n452 585
R579 B.n454 B.n453 585
R580 B.n937 B.n936 585
R581 B.n936 B.n935 585
R582 B.n938 B.n451 585
R583 B.n451 B.n450 585
R584 B.n940 B.n939 585
R585 B.n941 B.n940 585
R586 B.n445 B.n444 585
R587 B.n446 B.n445 585
R588 B.n949 B.n948 585
R589 B.n948 B.n947 585
R590 B.n950 B.n443 585
R591 B.n443 B.n442 585
R592 B.n952 B.n951 585
R593 B.n953 B.n952 585
R594 B.n437 B.n436 585
R595 B.n438 B.n437 585
R596 B.n961 B.n960 585
R597 B.n960 B.n959 585
R598 B.n962 B.n435 585
R599 B.n435 B.n434 585
R600 B.n964 B.n963 585
R601 B.n965 B.n964 585
R602 B.n429 B.n428 585
R603 B.n430 B.n429 585
R604 B.n973 B.n972 585
R605 B.n972 B.n971 585
R606 B.n974 B.n427 585
R607 B.n427 B.n426 585
R608 B.n976 B.n975 585
R609 B.n977 B.n976 585
R610 B.n421 B.n420 585
R611 B.n422 B.n421 585
R612 B.n985 B.n984 585
R613 B.n984 B.n983 585
R614 B.n986 B.n419 585
R615 B.n419 B.n418 585
R616 B.n988 B.n987 585
R617 B.n989 B.n988 585
R618 B.n413 B.n412 585
R619 B.n414 B.n413 585
R620 B.n997 B.n996 585
R621 B.n996 B.n995 585
R622 B.n998 B.n411 585
R623 B.n411 B.n410 585
R624 B.n1000 B.n999 585
R625 B.n1001 B.n1000 585
R626 B.n405 B.n404 585
R627 B.n406 B.n405 585
R628 B.n1010 B.n1009 585
R629 B.n1009 B.n1008 585
R630 B.n1011 B.n403 585
R631 B.n403 B.n402 585
R632 B.n1013 B.n1012 585
R633 B.n1014 B.n1013 585
R634 B.n3 B.n0 585
R635 B.n4 B.n3 585
R636 B.n1246 B.n1 585
R637 B.n1247 B.n1246 585
R638 B.n1245 B.n1244 585
R639 B.n1245 B.n8 585
R640 B.n1243 B.n9 585
R641 B.n12 B.n9 585
R642 B.n1242 B.n1241 585
R643 B.n1241 B.n1240 585
R644 B.n11 B.n10 585
R645 B.n1239 B.n11 585
R646 B.n1237 B.n1236 585
R647 B.n1238 B.n1237 585
R648 B.n1235 B.n17 585
R649 B.n17 B.n16 585
R650 B.n1234 B.n1233 585
R651 B.n1233 B.n1232 585
R652 B.n19 B.n18 585
R653 B.n1231 B.n19 585
R654 B.n1229 B.n1228 585
R655 B.n1230 B.n1229 585
R656 B.n1227 B.n24 585
R657 B.n24 B.n23 585
R658 B.n1226 B.n1225 585
R659 B.n1225 B.n1224 585
R660 B.n26 B.n25 585
R661 B.n1223 B.n26 585
R662 B.n1221 B.n1220 585
R663 B.n1222 B.n1221 585
R664 B.n1219 B.n31 585
R665 B.n31 B.n30 585
R666 B.n1218 B.n1217 585
R667 B.n1217 B.n1216 585
R668 B.n33 B.n32 585
R669 B.n1215 B.n33 585
R670 B.n1213 B.n1212 585
R671 B.n1214 B.n1213 585
R672 B.n1211 B.n38 585
R673 B.n38 B.n37 585
R674 B.n1210 B.n1209 585
R675 B.n1209 B.n1208 585
R676 B.n40 B.n39 585
R677 B.n1207 B.n40 585
R678 B.n1205 B.n1204 585
R679 B.n1206 B.n1205 585
R680 B.n1203 B.n45 585
R681 B.n45 B.n44 585
R682 B.n1202 B.n1201 585
R683 B.n1201 B.n1200 585
R684 B.n47 B.n46 585
R685 B.n1199 B.n47 585
R686 B.n1197 B.n1196 585
R687 B.n1198 B.n1197 585
R688 B.n1195 B.n52 585
R689 B.n52 B.n51 585
R690 B.n1194 B.n1193 585
R691 B.n1193 B.n1192 585
R692 B.n54 B.n53 585
R693 B.n1191 B.n54 585
R694 B.n1189 B.n1188 585
R695 B.n1190 B.n1189 585
R696 B.n1187 B.n59 585
R697 B.n59 B.n58 585
R698 B.n1186 B.n1185 585
R699 B.n1185 B.n1184 585
R700 B.n61 B.n60 585
R701 B.n1183 B.n61 585
R702 B.n1181 B.n1180 585
R703 B.n1182 B.n1181 585
R704 B.n1179 B.n66 585
R705 B.n66 B.n65 585
R706 B.n1178 B.n1177 585
R707 B.n1177 B.n1176 585
R708 B.n68 B.n67 585
R709 B.n1175 B.n68 585
R710 B.n1173 B.n1172 585
R711 B.n1174 B.n1173 585
R712 B.n1171 B.n73 585
R713 B.n73 B.n72 585
R714 B.n1170 B.n1169 585
R715 B.n1169 B.n1168 585
R716 B.n75 B.n74 585
R717 B.n1167 B.n75 585
R718 B.n1165 B.n1164 585
R719 B.n1166 B.n1165 585
R720 B.n1163 B.n80 585
R721 B.n80 B.n79 585
R722 B.n1162 B.n1161 585
R723 B.n1161 B.n1160 585
R724 B.n82 B.n81 585
R725 B.n1159 B.n82 585
R726 B.n1157 B.n1156 585
R727 B.n1158 B.n1157 585
R728 B.n1155 B.n87 585
R729 B.n87 B.n86 585
R730 B.n1154 B.n1153 585
R731 B.n1153 B.n1152 585
R732 B.n89 B.n88 585
R733 B.n1151 B.n89 585
R734 B.n1149 B.n1148 585
R735 B.n1150 B.n1149 585
R736 B.n1147 B.n94 585
R737 B.n94 B.n93 585
R738 B.n1146 B.n1145 585
R739 B.n1145 B.n1144 585
R740 B.n96 B.n95 585
R741 B.n1143 B.n96 585
R742 B.n1141 B.n1140 585
R743 B.n1142 B.n1141 585
R744 B.n1139 B.n101 585
R745 B.n101 B.n100 585
R746 B.n1138 B.n1137 585
R747 B.n1137 B.n1136 585
R748 B.n103 B.n102 585
R749 B.n1135 B.n103 585
R750 B.n1133 B.n1132 585
R751 B.n1134 B.n1133 585
R752 B.n1131 B.n108 585
R753 B.n108 B.n107 585
R754 B.n1130 B.n1129 585
R755 B.n1129 B.n1128 585
R756 B.n110 B.n109 585
R757 B.n1127 B.n110 585
R758 B.n1125 B.n1124 585
R759 B.n1126 B.n1125 585
R760 B.n1123 B.n115 585
R761 B.n115 B.n114 585
R762 B.n1122 B.n1121 585
R763 B.n1121 B.n1120 585
R764 B.n117 B.n116 585
R765 B.n1119 B.n117 585
R766 B.n1117 B.n1116 585
R767 B.n1118 B.n1117 585
R768 B.n1115 B.n122 585
R769 B.n122 B.n121 585
R770 B.n1114 B.n1113 585
R771 B.n1113 B.n1112 585
R772 B.n124 B.n123 585
R773 B.n1111 B.n124 585
R774 B.n1250 B.n1249 585
R775 B.n1248 B.n2 585
R776 B.n185 B.n124 521.33
R777 B.n1108 B.n126 521.33
R778 B.n810 B.n535 521.33
R779 B.n807 B.n533 521.33
R780 B.n183 B.t12 300.774
R781 B.n181 B.t19 300.774
R782 B.n595 B.t16 300.774
R783 B.n592 B.t8 300.774
R784 B.n1110 B.n1109 256.663
R785 B.n1110 B.n179 256.663
R786 B.n1110 B.n178 256.663
R787 B.n1110 B.n177 256.663
R788 B.n1110 B.n176 256.663
R789 B.n1110 B.n175 256.663
R790 B.n1110 B.n174 256.663
R791 B.n1110 B.n173 256.663
R792 B.n1110 B.n172 256.663
R793 B.n1110 B.n171 256.663
R794 B.n1110 B.n170 256.663
R795 B.n1110 B.n169 256.663
R796 B.n1110 B.n168 256.663
R797 B.n1110 B.n167 256.663
R798 B.n1110 B.n166 256.663
R799 B.n1110 B.n165 256.663
R800 B.n1110 B.n164 256.663
R801 B.n1110 B.n163 256.663
R802 B.n1110 B.n162 256.663
R803 B.n1110 B.n161 256.663
R804 B.n1110 B.n160 256.663
R805 B.n1110 B.n159 256.663
R806 B.n1110 B.n158 256.663
R807 B.n1110 B.n157 256.663
R808 B.n1110 B.n156 256.663
R809 B.n1110 B.n155 256.663
R810 B.n1110 B.n154 256.663
R811 B.n1110 B.n153 256.663
R812 B.n1110 B.n152 256.663
R813 B.n1110 B.n151 256.663
R814 B.n1110 B.n150 256.663
R815 B.n1110 B.n149 256.663
R816 B.n1110 B.n148 256.663
R817 B.n1110 B.n147 256.663
R818 B.n1110 B.n146 256.663
R819 B.n1110 B.n145 256.663
R820 B.n1110 B.n144 256.663
R821 B.n1110 B.n143 256.663
R822 B.n1110 B.n142 256.663
R823 B.n1110 B.n141 256.663
R824 B.n1110 B.n140 256.663
R825 B.n1110 B.n139 256.663
R826 B.n1110 B.n138 256.663
R827 B.n1110 B.n137 256.663
R828 B.n1110 B.n136 256.663
R829 B.n1110 B.n135 256.663
R830 B.n1110 B.n134 256.663
R831 B.n1110 B.n133 256.663
R832 B.n1110 B.n132 256.663
R833 B.n1110 B.n131 256.663
R834 B.n1110 B.n130 256.663
R835 B.n1110 B.n129 256.663
R836 B.n1110 B.n128 256.663
R837 B.n1110 B.n127 256.663
R838 B.n809 B.n808 256.663
R839 B.n809 B.n538 256.663
R840 B.n809 B.n539 256.663
R841 B.n809 B.n540 256.663
R842 B.n809 B.n541 256.663
R843 B.n809 B.n542 256.663
R844 B.n809 B.n543 256.663
R845 B.n809 B.n544 256.663
R846 B.n809 B.n545 256.663
R847 B.n809 B.n546 256.663
R848 B.n809 B.n547 256.663
R849 B.n809 B.n548 256.663
R850 B.n809 B.n549 256.663
R851 B.n809 B.n550 256.663
R852 B.n809 B.n551 256.663
R853 B.n809 B.n552 256.663
R854 B.n809 B.n553 256.663
R855 B.n809 B.n554 256.663
R856 B.n809 B.n555 256.663
R857 B.n809 B.n556 256.663
R858 B.n809 B.n557 256.663
R859 B.n809 B.n558 256.663
R860 B.n809 B.n559 256.663
R861 B.n809 B.n560 256.663
R862 B.n809 B.n561 256.663
R863 B.n809 B.n562 256.663
R864 B.n809 B.n563 256.663
R865 B.n809 B.n564 256.663
R866 B.n809 B.n565 256.663
R867 B.n809 B.n566 256.663
R868 B.n809 B.n567 256.663
R869 B.n809 B.n568 256.663
R870 B.n809 B.n569 256.663
R871 B.n809 B.n570 256.663
R872 B.n809 B.n571 256.663
R873 B.n809 B.n572 256.663
R874 B.n809 B.n573 256.663
R875 B.n809 B.n574 256.663
R876 B.n809 B.n575 256.663
R877 B.n809 B.n576 256.663
R878 B.n809 B.n577 256.663
R879 B.n809 B.n578 256.663
R880 B.n809 B.n579 256.663
R881 B.n809 B.n580 256.663
R882 B.n809 B.n581 256.663
R883 B.n809 B.n582 256.663
R884 B.n809 B.n583 256.663
R885 B.n809 B.n584 256.663
R886 B.n809 B.n585 256.663
R887 B.n809 B.n586 256.663
R888 B.n809 B.n587 256.663
R889 B.n809 B.n588 256.663
R890 B.n809 B.n589 256.663
R891 B.n1252 B.n1251 256.663
R892 B.n189 B.n188 163.367
R893 B.n193 B.n192 163.367
R894 B.n197 B.n196 163.367
R895 B.n201 B.n200 163.367
R896 B.n205 B.n204 163.367
R897 B.n209 B.n208 163.367
R898 B.n213 B.n212 163.367
R899 B.n217 B.n216 163.367
R900 B.n221 B.n220 163.367
R901 B.n225 B.n224 163.367
R902 B.n229 B.n228 163.367
R903 B.n233 B.n232 163.367
R904 B.n237 B.n236 163.367
R905 B.n241 B.n240 163.367
R906 B.n245 B.n244 163.367
R907 B.n249 B.n248 163.367
R908 B.n253 B.n252 163.367
R909 B.n257 B.n256 163.367
R910 B.n261 B.n260 163.367
R911 B.n265 B.n264 163.367
R912 B.n269 B.n268 163.367
R913 B.n273 B.n272 163.367
R914 B.n277 B.n276 163.367
R915 B.n281 B.n280 163.367
R916 B.n286 B.n285 163.367
R917 B.n290 B.n289 163.367
R918 B.n294 B.n293 163.367
R919 B.n298 B.n297 163.367
R920 B.n302 B.n301 163.367
R921 B.n307 B.n306 163.367
R922 B.n311 B.n310 163.367
R923 B.n315 B.n314 163.367
R924 B.n319 B.n318 163.367
R925 B.n323 B.n322 163.367
R926 B.n327 B.n326 163.367
R927 B.n331 B.n330 163.367
R928 B.n335 B.n334 163.367
R929 B.n339 B.n338 163.367
R930 B.n343 B.n342 163.367
R931 B.n347 B.n346 163.367
R932 B.n351 B.n350 163.367
R933 B.n355 B.n354 163.367
R934 B.n359 B.n358 163.367
R935 B.n363 B.n362 163.367
R936 B.n367 B.n366 163.367
R937 B.n371 B.n370 163.367
R938 B.n375 B.n374 163.367
R939 B.n379 B.n378 163.367
R940 B.n383 B.n382 163.367
R941 B.n387 B.n386 163.367
R942 B.n391 B.n390 163.367
R943 B.n395 B.n394 163.367
R944 B.n397 B.n180 163.367
R945 B.n814 B.n535 163.367
R946 B.n814 B.n529 163.367
R947 B.n822 B.n529 163.367
R948 B.n822 B.n527 163.367
R949 B.n826 B.n527 163.367
R950 B.n826 B.n521 163.367
R951 B.n834 B.n521 163.367
R952 B.n834 B.n519 163.367
R953 B.n838 B.n519 163.367
R954 B.n838 B.n513 163.367
R955 B.n846 B.n513 163.367
R956 B.n846 B.n511 163.367
R957 B.n850 B.n511 163.367
R958 B.n850 B.n505 163.367
R959 B.n858 B.n505 163.367
R960 B.n858 B.n503 163.367
R961 B.n862 B.n503 163.367
R962 B.n862 B.n497 163.367
R963 B.n870 B.n497 163.367
R964 B.n870 B.n495 163.367
R965 B.n874 B.n495 163.367
R966 B.n874 B.n488 163.367
R967 B.n882 B.n488 163.367
R968 B.n882 B.n486 163.367
R969 B.n886 B.n486 163.367
R970 B.n886 B.n481 163.367
R971 B.n894 B.n481 163.367
R972 B.n894 B.n479 163.367
R973 B.n898 B.n479 163.367
R974 B.n898 B.n473 163.367
R975 B.n906 B.n473 163.367
R976 B.n906 B.n471 163.367
R977 B.n910 B.n471 163.367
R978 B.n910 B.n465 163.367
R979 B.n918 B.n465 163.367
R980 B.n918 B.n463 163.367
R981 B.n922 B.n463 163.367
R982 B.n922 B.n457 163.367
R983 B.n930 B.n457 163.367
R984 B.n930 B.n455 163.367
R985 B.n934 B.n455 163.367
R986 B.n934 B.n449 163.367
R987 B.n942 B.n449 163.367
R988 B.n942 B.n447 163.367
R989 B.n946 B.n447 163.367
R990 B.n946 B.n441 163.367
R991 B.n954 B.n441 163.367
R992 B.n954 B.n439 163.367
R993 B.n958 B.n439 163.367
R994 B.n958 B.n433 163.367
R995 B.n966 B.n433 163.367
R996 B.n966 B.n431 163.367
R997 B.n970 B.n431 163.367
R998 B.n970 B.n425 163.367
R999 B.n978 B.n425 163.367
R1000 B.n978 B.n423 163.367
R1001 B.n982 B.n423 163.367
R1002 B.n982 B.n417 163.367
R1003 B.n990 B.n417 163.367
R1004 B.n990 B.n415 163.367
R1005 B.n994 B.n415 163.367
R1006 B.n994 B.n409 163.367
R1007 B.n1002 B.n409 163.367
R1008 B.n1002 B.n407 163.367
R1009 B.n1007 B.n407 163.367
R1010 B.n1007 B.n401 163.367
R1011 B.n1015 B.n401 163.367
R1012 B.n1016 B.n1015 163.367
R1013 B.n1016 B.n5 163.367
R1014 B.n6 B.n5 163.367
R1015 B.n7 B.n6 163.367
R1016 B.n1022 B.n7 163.367
R1017 B.n1023 B.n1022 163.367
R1018 B.n1023 B.n13 163.367
R1019 B.n14 B.n13 163.367
R1020 B.n15 B.n14 163.367
R1021 B.n1028 B.n15 163.367
R1022 B.n1028 B.n20 163.367
R1023 B.n21 B.n20 163.367
R1024 B.n22 B.n21 163.367
R1025 B.n1033 B.n22 163.367
R1026 B.n1033 B.n27 163.367
R1027 B.n28 B.n27 163.367
R1028 B.n29 B.n28 163.367
R1029 B.n1038 B.n29 163.367
R1030 B.n1038 B.n34 163.367
R1031 B.n35 B.n34 163.367
R1032 B.n36 B.n35 163.367
R1033 B.n1043 B.n36 163.367
R1034 B.n1043 B.n41 163.367
R1035 B.n42 B.n41 163.367
R1036 B.n43 B.n42 163.367
R1037 B.n1048 B.n43 163.367
R1038 B.n1048 B.n48 163.367
R1039 B.n49 B.n48 163.367
R1040 B.n50 B.n49 163.367
R1041 B.n1053 B.n50 163.367
R1042 B.n1053 B.n55 163.367
R1043 B.n56 B.n55 163.367
R1044 B.n57 B.n56 163.367
R1045 B.n1058 B.n57 163.367
R1046 B.n1058 B.n62 163.367
R1047 B.n63 B.n62 163.367
R1048 B.n64 B.n63 163.367
R1049 B.n1063 B.n64 163.367
R1050 B.n1063 B.n69 163.367
R1051 B.n70 B.n69 163.367
R1052 B.n71 B.n70 163.367
R1053 B.n1068 B.n71 163.367
R1054 B.n1068 B.n76 163.367
R1055 B.n77 B.n76 163.367
R1056 B.n78 B.n77 163.367
R1057 B.n1073 B.n78 163.367
R1058 B.n1073 B.n83 163.367
R1059 B.n84 B.n83 163.367
R1060 B.n85 B.n84 163.367
R1061 B.n1078 B.n85 163.367
R1062 B.n1078 B.n90 163.367
R1063 B.n91 B.n90 163.367
R1064 B.n92 B.n91 163.367
R1065 B.n1083 B.n92 163.367
R1066 B.n1083 B.n97 163.367
R1067 B.n98 B.n97 163.367
R1068 B.n99 B.n98 163.367
R1069 B.n1088 B.n99 163.367
R1070 B.n1088 B.n104 163.367
R1071 B.n105 B.n104 163.367
R1072 B.n106 B.n105 163.367
R1073 B.n1093 B.n106 163.367
R1074 B.n1093 B.n111 163.367
R1075 B.n112 B.n111 163.367
R1076 B.n113 B.n112 163.367
R1077 B.n1098 B.n113 163.367
R1078 B.n1098 B.n118 163.367
R1079 B.n119 B.n118 163.367
R1080 B.n120 B.n119 163.367
R1081 B.n1103 B.n120 163.367
R1082 B.n1103 B.n125 163.367
R1083 B.n126 B.n125 163.367
R1084 B.n591 B.n590 163.367
R1085 B.n802 B.n590 163.367
R1086 B.n800 B.n799 163.367
R1087 B.n796 B.n795 163.367
R1088 B.n792 B.n791 163.367
R1089 B.n788 B.n787 163.367
R1090 B.n784 B.n783 163.367
R1091 B.n780 B.n779 163.367
R1092 B.n776 B.n775 163.367
R1093 B.n772 B.n771 163.367
R1094 B.n768 B.n767 163.367
R1095 B.n764 B.n763 163.367
R1096 B.n760 B.n759 163.367
R1097 B.n756 B.n755 163.367
R1098 B.n752 B.n751 163.367
R1099 B.n748 B.n747 163.367
R1100 B.n744 B.n743 163.367
R1101 B.n740 B.n739 163.367
R1102 B.n736 B.n735 163.367
R1103 B.n732 B.n731 163.367
R1104 B.n728 B.n727 163.367
R1105 B.n724 B.n723 163.367
R1106 B.n720 B.n719 163.367
R1107 B.n716 B.n715 163.367
R1108 B.n712 B.n711 163.367
R1109 B.n708 B.n707 163.367
R1110 B.n704 B.n703 163.367
R1111 B.n700 B.n699 163.367
R1112 B.n696 B.n695 163.367
R1113 B.n692 B.n691 163.367
R1114 B.n688 B.n687 163.367
R1115 B.n684 B.n683 163.367
R1116 B.n680 B.n679 163.367
R1117 B.n676 B.n675 163.367
R1118 B.n672 B.n671 163.367
R1119 B.n668 B.n667 163.367
R1120 B.n664 B.n663 163.367
R1121 B.n660 B.n659 163.367
R1122 B.n656 B.n655 163.367
R1123 B.n652 B.n651 163.367
R1124 B.n648 B.n647 163.367
R1125 B.n644 B.n643 163.367
R1126 B.n640 B.n639 163.367
R1127 B.n636 B.n635 163.367
R1128 B.n632 B.n631 163.367
R1129 B.n628 B.n627 163.367
R1130 B.n624 B.n623 163.367
R1131 B.n620 B.n619 163.367
R1132 B.n616 B.n615 163.367
R1133 B.n612 B.n611 163.367
R1134 B.n608 B.n607 163.367
R1135 B.n604 B.n603 163.367
R1136 B.n600 B.n599 163.367
R1137 B.n810 B.n537 163.367
R1138 B.n816 B.n533 163.367
R1139 B.n816 B.n531 163.367
R1140 B.n820 B.n531 163.367
R1141 B.n820 B.n525 163.367
R1142 B.n828 B.n525 163.367
R1143 B.n828 B.n523 163.367
R1144 B.n832 B.n523 163.367
R1145 B.n832 B.n517 163.367
R1146 B.n840 B.n517 163.367
R1147 B.n840 B.n515 163.367
R1148 B.n844 B.n515 163.367
R1149 B.n844 B.n509 163.367
R1150 B.n852 B.n509 163.367
R1151 B.n852 B.n507 163.367
R1152 B.n856 B.n507 163.367
R1153 B.n856 B.n501 163.367
R1154 B.n864 B.n501 163.367
R1155 B.n864 B.n499 163.367
R1156 B.n868 B.n499 163.367
R1157 B.n868 B.n493 163.367
R1158 B.n876 B.n493 163.367
R1159 B.n876 B.n491 163.367
R1160 B.n880 B.n491 163.367
R1161 B.n880 B.n485 163.367
R1162 B.n888 B.n485 163.367
R1163 B.n888 B.n483 163.367
R1164 B.n892 B.n483 163.367
R1165 B.n892 B.n477 163.367
R1166 B.n900 B.n477 163.367
R1167 B.n900 B.n475 163.367
R1168 B.n904 B.n475 163.367
R1169 B.n904 B.n469 163.367
R1170 B.n912 B.n469 163.367
R1171 B.n912 B.n467 163.367
R1172 B.n916 B.n467 163.367
R1173 B.n916 B.n461 163.367
R1174 B.n924 B.n461 163.367
R1175 B.n924 B.n459 163.367
R1176 B.n928 B.n459 163.367
R1177 B.n928 B.n453 163.367
R1178 B.n936 B.n453 163.367
R1179 B.n936 B.n451 163.367
R1180 B.n940 B.n451 163.367
R1181 B.n940 B.n445 163.367
R1182 B.n948 B.n445 163.367
R1183 B.n948 B.n443 163.367
R1184 B.n952 B.n443 163.367
R1185 B.n952 B.n437 163.367
R1186 B.n960 B.n437 163.367
R1187 B.n960 B.n435 163.367
R1188 B.n964 B.n435 163.367
R1189 B.n964 B.n429 163.367
R1190 B.n972 B.n429 163.367
R1191 B.n972 B.n427 163.367
R1192 B.n976 B.n427 163.367
R1193 B.n976 B.n421 163.367
R1194 B.n984 B.n421 163.367
R1195 B.n984 B.n419 163.367
R1196 B.n988 B.n419 163.367
R1197 B.n988 B.n413 163.367
R1198 B.n996 B.n413 163.367
R1199 B.n996 B.n411 163.367
R1200 B.n1000 B.n411 163.367
R1201 B.n1000 B.n405 163.367
R1202 B.n1009 B.n405 163.367
R1203 B.n1009 B.n403 163.367
R1204 B.n1013 B.n403 163.367
R1205 B.n1013 B.n3 163.367
R1206 B.n1250 B.n3 163.367
R1207 B.n1246 B.n2 163.367
R1208 B.n1246 B.n1245 163.367
R1209 B.n1245 B.n9 163.367
R1210 B.n1241 B.n9 163.367
R1211 B.n1241 B.n11 163.367
R1212 B.n1237 B.n11 163.367
R1213 B.n1237 B.n17 163.367
R1214 B.n1233 B.n17 163.367
R1215 B.n1233 B.n19 163.367
R1216 B.n1229 B.n19 163.367
R1217 B.n1229 B.n24 163.367
R1218 B.n1225 B.n24 163.367
R1219 B.n1225 B.n26 163.367
R1220 B.n1221 B.n26 163.367
R1221 B.n1221 B.n31 163.367
R1222 B.n1217 B.n31 163.367
R1223 B.n1217 B.n33 163.367
R1224 B.n1213 B.n33 163.367
R1225 B.n1213 B.n38 163.367
R1226 B.n1209 B.n38 163.367
R1227 B.n1209 B.n40 163.367
R1228 B.n1205 B.n40 163.367
R1229 B.n1205 B.n45 163.367
R1230 B.n1201 B.n45 163.367
R1231 B.n1201 B.n47 163.367
R1232 B.n1197 B.n47 163.367
R1233 B.n1197 B.n52 163.367
R1234 B.n1193 B.n52 163.367
R1235 B.n1193 B.n54 163.367
R1236 B.n1189 B.n54 163.367
R1237 B.n1189 B.n59 163.367
R1238 B.n1185 B.n59 163.367
R1239 B.n1185 B.n61 163.367
R1240 B.n1181 B.n61 163.367
R1241 B.n1181 B.n66 163.367
R1242 B.n1177 B.n66 163.367
R1243 B.n1177 B.n68 163.367
R1244 B.n1173 B.n68 163.367
R1245 B.n1173 B.n73 163.367
R1246 B.n1169 B.n73 163.367
R1247 B.n1169 B.n75 163.367
R1248 B.n1165 B.n75 163.367
R1249 B.n1165 B.n80 163.367
R1250 B.n1161 B.n80 163.367
R1251 B.n1161 B.n82 163.367
R1252 B.n1157 B.n82 163.367
R1253 B.n1157 B.n87 163.367
R1254 B.n1153 B.n87 163.367
R1255 B.n1153 B.n89 163.367
R1256 B.n1149 B.n89 163.367
R1257 B.n1149 B.n94 163.367
R1258 B.n1145 B.n94 163.367
R1259 B.n1145 B.n96 163.367
R1260 B.n1141 B.n96 163.367
R1261 B.n1141 B.n101 163.367
R1262 B.n1137 B.n101 163.367
R1263 B.n1137 B.n103 163.367
R1264 B.n1133 B.n103 163.367
R1265 B.n1133 B.n108 163.367
R1266 B.n1129 B.n108 163.367
R1267 B.n1129 B.n110 163.367
R1268 B.n1125 B.n110 163.367
R1269 B.n1125 B.n115 163.367
R1270 B.n1121 B.n115 163.367
R1271 B.n1121 B.n117 163.367
R1272 B.n1117 B.n117 163.367
R1273 B.n1117 B.n122 163.367
R1274 B.n1113 B.n122 163.367
R1275 B.n1113 B.n124 163.367
R1276 B.n181 B.t20 154.773
R1277 B.n595 B.t18 154.773
R1278 B.n183 B.t14 154.754
R1279 B.n592 B.t11 154.754
R1280 B.n184 B.n183 81.0672
R1281 B.n182 B.n181 81.0672
R1282 B.n596 B.n595 81.0672
R1283 B.n593 B.n592 81.0672
R1284 B.n182 B.t21 73.7056
R1285 B.n596 B.t17 73.7056
R1286 B.n184 B.t15 73.6869
R1287 B.n593 B.t10 73.6869
R1288 B.n185 B.n127 71.676
R1289 B.n189 B.n128 71.676
R1290 B.n193 B.n129 71.676
R1291 B.n197 B.n130 71.676
R1292 B.n201 B.n131 71.676
R1293 B.n205 B.n132 71.676
R1294 B.n209 B.n133 71.676
R1295 B.n213 B.n134 71.676
R1296 B.n217 B.n135 71.676
R1297 B.n221 B.n136 71.676
R1298 B.n225 B.n137 71.676
R1299 B.n229 B.n138 71.676
R1300 B.n233 B.n139 71.676
R1301 B.n237 B.n140 71.676
R1302 B.n241 B.n141 71.676
R1303 B.n245 B.n142 71.676
R1304 B.n249 B.n143 71.676
R1305 B.n253 B.n144 71.676
R1306 B.n257 B.n145 71.676
R1307 B.n261 B.n146 71.676
R1308 B.n265 B.n147 71.676
R1309 B.n269 B.n148 71.676
R1310 B.n273 B.n149 71.676
R1311 B.n277 B.n150 71.676
R1312 B.n281 B.n151 71.676
R1313 B.n286 B.n152 71.676
R1314 B.n290 B.n153 71.676
R1315 B.n294 B.n154 71.676
R1316 B.n298 B.n155 71.676
R1317 B.n302 B.n156 71.676
R1318 B.n307 B.n157 71.676
R1319 B.n311 B.n158 71.676
R1320 B.n315 B.n159 71.676
R1321 B.n319 B.n160 71.676
R1322 B.n323 B.n161 71.676
R1323 B.n327 B.n162 71.676
R1324 B.n331 B.n163 71.676
R1325 B.n335 B.n164 71.676
R1326 B.n339 B.n165 71.676
R1327 B.n343 B.n166 71.676
R1328 B.n347 B.n167 71.676
R1329 B.n351 B.n168 71.676
R1330 B.n355 B.n169 71.676
R1331 B.n359 B.n170 71.676
R1332 B.n363 B.n171 71.676
R1333 B.n367 B.n172 71.676
R1334 B.n371 B.n173 71.676
R1335 B.n375 B.n174 71.676
R1336 B.n379 B.n175 71.676
R1337 B.n383 B.n176 71.676
R1338 B.n387 B.n177 71.676
R1339 B.n391 B.n178 71.676
R1340 B.n395 B.n179 71.676
R1341 B.n1109 B.n180 71.676
R1342 B.n1109 B.n1108 71.676
R1343 B.n397 B.n179 71.676
R1344 B.n394 B.n178 71.676
R1345 B.n390 B.n177 71.676
R1346 B.n386 B.n176 71.676
R1347 B.n382 B.n175 71.676
R1348 B.n378 B.n174 71.676
R1349 B.n374 B.n173 71.676
R1350 B.n370 B.n172 71.676
R1351 B.n366 B.n171 71.676
R1352 B.n362 B.n170 71.676
R1353 B.n358 B.n169 71.676
R1354 B.n354 B.n168 71.676
R1355 B.n350 B.n167 71.676
R1356 B.n346 B.n166 71.676
R1357 B.n342 B.n165 71.676
R1358 B.n338 B.n164 71.676
R1359 B.n334 B.n163 71.676
R1360 B.n330 B.n162 71.676
R1361 B.n326 B.n161 71.676
R1362 B.n322 B.n160 71.676
R1363 B.n318 B.n159 71.676
R1364 B.n314 B.n158 71.676
R1365 B.n310 B.n157 71.676
R1366 B.n306 B.n156 71.676
R1367 B.n301 B.n155 71.676
R1368 B.n297 B.n154 71.676
R1369 B.n293 B.n153 71.676
R1370 B.n289 B.n152 71.676
R1371 B.n285 B.n151 71.676
R1372 B.n280 B.n150 71.676
R1373 B.n276 B.n149 71.676
R1374 B.n272 B.n148 71.676
R1375 B.n268 B.n147 71.676
R1376 B.n264 B.n146 71.676
R1377 B.n260 B.n145 71.676
R1378 B.n256 B.n144 71.676
R1379 B.n252 B.n143 71.676
R1380 B.n248 B.n142 71.676
R1381 B.n244 B.n141 71.676
R1382 B.n240 B.n140 71.676
R1383 B.n236 B.n139 71.676
R1384 B.n232 B.n138 71.676
R1385 B.n228 B.n137 71.676
R1386 B.n224 B.n136 71.676
R1387 B.n220 B.n135 71.676
R1388 B.n216 B.n134 71.676
R1389 B.n212 B.n133 71.676
R1390 B.n208 B.n132 71.676
R1391 B.n204 B.n131 71.676
R1392 B.n200 B.n130 71.676
R1393 B.n196 B.n129 71.676
R1394 B.n192 B.n128 71.676
R1395 B.n188 B.n127 71.676
R1396 B.n808 B.n807 71.676
R1397 B.n802 B.n538 71.676
R1398 B.n799 B.n539 71.676
R1399 B.n795 B.n540 71.676
R1400 B.n791 B.n541 71.676
R1401 B.n787 B.n542 71.676
R1402 B.n783 B.n543 71.676
R1403 B.n779 B.n544 71.676
R1404 B.n775 B.n545 71.676
R1405 B.n771 B.n546 71.676
R1406 B.n767 B.n547 71.676
R1407 B.n763 B.n548 71.676
R1408 B.n759 B.n549 71.676
R1409 B.n755 B.n550 71.676
R1410 B.n751 B.n551 71.676
R1411 B.n747 B.n552 71.676
R1412 B.n743 B.n553 71.676
R1413 B.n739 B.n554 71.676
R1414 B.n735 B.n555 71.676
R1415 B.n731 B.n556 71.676
R1416 B.n727 B.n557 71.676
R1417 B.n723 B.n558 71.676
R1418 B.n719 B.n559 71.676
R1419 B.n715 B.n560 71.676
R1420 B.n711 B.n561 71.676
R1421 B.n707 B.n562 71.676
R1422 B.n703 B.n563 71.676
R1423 B.n699 B.n564 71.676
R1424 B.n695 B.n565 71.676
R1425 B.n691 B.n566 71.676
R1426 B.n687 B.n567 71.676
R1427 B.n683 B.n568 71.676
R1428 B.n679 B.n569 71.676
R1429 B.n675 B.n570 71.676
R1430 B.n671 B.n571 71.676
R1431 B.n667 B.n572 71.676
R1432 B.n663 B.n573 71.676
R1433 B.n659 B.n574 71.676
R1434 B.n655 B.n575 71.676
R1435 B.n651 B.n576 71.676
R1436 B.n647 B.n577 71.676
R1437 B.n643 B.n578 71.676
R1438 B.n639 B.n579 71.676
R1439 B.n635 B.n580 71.676
R1440 B.n631 B.n581 71.676
R1441 B.n627 B.n582 71.676
R1442 B.n623 B.n583 71.676
R1443 B.n619 B.n584 71.676
R1444 B.n615 B.n585 71.676
R1445 B.n611 B.n586 71.676
R1446 B.n607 B.n587 71.676
R1447 B.n603 B.n588 71.676
R1448 B.n599 B.n589 71.676
R1449 B.n808 B.n591 71.676
R1450 B.n800 B.n538 71.676
R1451 B.n796 B.n539 71.676
R1452 B.n792 B.n540 71.676
R1453 B.n788 B.n541 71.676
R1454 B.n784 B.n542 71.676
R1455 B.n780 B.n543 71.676
R1456 B.n776 B.n544 71.676
R1457 B.n772 B.n545 71.676
R1458 B.n768 B.n546 71.676
R1459 B.n764 B.n547 71.676
R1460 B.n760 B.n548 71.676
R1461 B.n756 B.n549 71.676
R1462 B.n752 B.n550 71.676
R1463 B.n748 B.n551 71.676
R1464 B.n744 B.n552 71.676
R1465 B.n740 B.n553 71.676
R1466 B.n736 B.n554 71.676
R1467 B.n732 B.n555 71.676
R1468 B.n728 B.n556 71.676
R1469 B.n724 B.n557 71.676
R1470 B.n720 B.n558 71.676
R1471 B.n716 B.n559 71.676
R1472 B.n712 B.n560 71.676
R1473 B.n708 B.n561 71.676
R1474 B.n704 B.n562 71.676
R1475 B.n700 B.n563 71.676
R1476 B.n696 B.n564 71.676
R1477 B.n692 B.n565 71.676
R1478 B.n688 B.n566 71.676
R1479 B.n684 B.n567 71.676
R1480 B.n680 B.n568 71.676
R1481 B.n676 B.n569 71.676
R1482 B.n672 B.n570 71.676
R1483 B.n668 B.n571 71.676
R1484 B.n664 B.n572 71.676
R1485 B.n660 B.n573 71.676
R1486 B.n656 B.n574 71.676
R1487 B.n652 B.n575 71.676
R1488 B.n648 B.n576 71.676
R1489 B.n644 B.n577 71.676
R1490 B.n640 B.n578 71.676
R1491 B.n636 B.n579 71.676
R1492 B.n632 B.n580 71.676
R1493 B.n628 B.n581 71.676
R1494 B.n624 B.n582 71.676
R1495 B.n620 B.n583 71.676
R1496 B.n616 B.n584 71.676
R1497 B.n612 B.n585 71.676
R1498 B.n608 B.n586 71.676
R1499 B.n604 B.n587 71.676
R1500 B.n600 B.n588 71.676
R1501 B.n589 B.n537 71.676
R1502 B.n1251 B.n1250 71.676
R1503 B.n1251 B.n2 71.676
R1504 B.n809 B.n534 71.3967
R1505 B.n1111 B.n1110 71.3967
R1506 B.n283 B.n184 59.5399
R1507 B.n304 B.n182 59.5399
R1508 B.n597 B.n596 59.5399
R1509 B.n594 B.n593 59.5399
R1510 B.n815 B.n534 37.6357
R1511 B.n815 B.n530 37.6357
R1512 B.n821 B.n530 37.6357
R1513 B.n821 B.n526 37.6357
R1514 B.n827 B.n526 37.6357
R1515 B.n827 B.n522 37.6357
R1516 B.n833 B.n522 37.6357
R1517 B.n833 B.n518 37.6357
R1518 B.n839 B.n518 37.6357
R1519 B.n845 B.n514 37.6357
R1520 B.n845 B.n510 37.6357
R1521 B.n851 B.n510 37.6357
R1522 B.n851 B.n506 37.6357
R1523 B.n857 B.n506 37.6357
R1524 B.n857 B.n502 37.6357
R1525 B.n863 B.n502 37.6357
R1526 B.n863 B.n498 37.6357
R1527 B.n869 B.n498 37.6357
R1528 B.n869 B.n494 37.6357
R1529 B.n875 B.n494 37.6357
R1530 B.n875 B.n489 37.6357
R1531 B.n881 B.n489 37.6357
R1532 B.n881 B.n490 37.6357
R1533 B.n887 B.n482 37.6357
R1534 B.n893 B.n482 37.6357
R1535 B.n893 B.n478 37.6357
R1536 B.n899 B.n478 37.6357
R1537 B.n899 B.n474 37.6357
R1538 B.n905 B.n474 37.6357
R1539 B.n905 B.n470 37.6357
R1540 B.n911 B.n470 37.6357
R1541 B.n911 B.n466 37.6357
R1542 B.n917 B.n466 37.6357
R1543 B.n917 B.n462 37.6357
R1544 B.n923 B.n462 37.6357
R1545 B.n929 B.n458 37.6357
R1546 B.n929 B.n454 37.6357
R1547 B.n935 B.n454 37.6357
R1548 B.n935 B.n450 37.6357
R1549 B.n941 B.n450 37.6357
R1550 B.n941 B.n446 37.6357
R1551 B.n947 B.n446 37.6357
R1552 B.n947 B.n442 37.6357
R1553 B.n953 B.n442 37.6357
R1554 B.n953 B.n438 37.6357
R1555 B.n959 B.n438 37.6357
R1556 B.n965 B.n434 37.6357
R1557 B.n965 B.n430 37.6357
R1558 B.n971 B.n430 37.6357
R1559 B.n971 B.n426 37.6357
R1560 B.n977 B.n426 37.6357
R1561 B.n977 B.n422 37.6357
R1562 B.n983 B.n422 37.6357
R1563 B.n983 B.n418 37.6357
R1564 B.n989 B.n418 37.6357
R1565 B.n989 B.n414 37.6357
R1566 B.n995 B.n414 37.6357
R1567 B.n1001 B.n410 37.6357
R1568 B.n1001 B.n406 37.6357
R1569 B.n1008 B.n406 37.6357
R1570 B.n1008 B.n402 37.6357
R1571 B.n1014 B.n402 37.6357
R1572 B.n1014 B.n4 37.6357
R1573 B.n1249 B.n4 37.6357
R1574 B.n1249 B.n1248 37.6357
R1575 B.n1248 B.n1247 37.6357
R1576 B.n1247 B.n8 37.6357
R1577 B.n12 B.n8 37.6357
R1578 B.n1240 B.n12 37.6357
R1579 B.n1240 B.n1239 37.6357
R1580 B.n1239 B.n1238 37.6357
R1581 B.n1238 B.n16 37.6357
R1582 B.n1232 B.n1231 37.6357
R1583 B.n1231 B.n1230 37.6357
R1584 B.n1230 B.n23 37.6357
R1585 B.n1224 B.n23 37.6357
R1586 B.n1224 B.n1223 37.6357
R1587 B.n1223 B.n1222 37.6357
R1588 B.n1222 B.n30 37.6357
R1589 B.n1216 B.n30 37.6357
R1590 B.n1216 B.n1215 37.6357
R1591 B.n1215 B.n1214 37.6357
R1592 B.n1214 B.n37 37.6357
R1593 B.n1208 B.n1207 37.6357
R1594 B.n1207 B.n1206 37.6357
R1595 B.n1206 B.n44 37.6357
R1596 B.n1200 B.n44 37.6357
R1597 B.n1200 B.n1199 37.6357
R1598 B.n1199 B.n1198 37.6357
R1599 B.n1198 B.n51 37.6357
R1600 B.n1192 B.n51 37.6357
R1601 B.n1192 B.n1191 37.6357
R1602 B.n1191 B.n1190 37.6357
R1603 B.n1190 B.n58 37.6357
R1604 B.n1184 B.n1183 37.6357
R1605 B.n1183 B.n1182 37.6357
R1606 B.n1182 B.n65 37.6357
R1607 B.n1176 B.n65 37.6357
R1608 B.n1176 B.n1175 37.6357
R1609 B.n1175 B.n1174 37.6357
R1610 B.n1174 B.n72 37.6357
R1611 B.n1168 B.n72 37.6357
R1612 B.n1168 B.n1167 37.6357
R1613 B.n1167 B.n1166 37.6357
R1614 B.n1166 B.n79 37.6357
R1615 B.n1160 B.n79 37.6357
R1616 B.n1159 B.n1158 37.6357
R1617 B.n1158 B.n86 37.6357
R1618 B.n1152 B.n86 37.6357
R1619 B.n1152 B.n1151 37.6357
R1620 B.n1151 B.n1150 37.6357
R1621 B.n1150 B.n93 37.6357
R1622 B.n1144 B.n93 37.6357
R1623 B.n1144 B.n1143 37.6357
R1624 B.n1143 B.n1142 37.6357
R1625 B.n1142 B.n100 37.6357
R1626 B.n1136 B.n100 37.6357
R1627 B.n1136 B.n1135 37.6357
R1628 B.n1135 B.n1134 37.6357
R1629 B.n1134 B.n107 37.6357
R1630 B.n1128 B.n1127 37.6357
R1631 B.n1127 B.n1126 37.6357
R1632 B.n1126 B.n114 37.6357
R1633 B.n1120 B.n114 37.6357
R1634 B.n1120 B.n1119 37.6357
R1635 B.n1119 B.n1118 37.6357
R1636 B.n1118 B.n121 37.6357
R1637 B.n1112 B.n121 37.6357
R1638 B.n1112 B.n1111 37.6357
R1639 B.n806 B.n532 33.8737
R1640 B.n812 B.n811 33.8737
R1641 B.n1107 B.n1106 33.8737
R1642 B.n186 B.n123 33.8737
R1643 B.n490 B.t4 32.6546
R1644 B.t6 B.n1159 32.6546
R1645 B.t7 B.n458 31.5477
R1646 B.t5 B.n58 31.5477
R1647 B.n995 B.t1 28.2269
R1648 B.n1232 B.t0 28.2269
R1649 B.t9 B.n514 23.7992
R1650 B.t13 B.n107 23.7992
R1651 B.t2 B.n434 20.4785
R1652 B.t3 B.n37 20.4785
R1653 B B.n1252 18.0485
R1654 B.n959 B.t2 17.1577
R1655 B.n1208 B.t3 17.1577
R1656 B.n839 B.t9 13.837
R1657 B.n1128 B.t13 13.837
R1658 B.n817 B.n532 10.6151
R1659 B.n818 B.n817 10.6151
R1660 B.n819 B.n818 10.6151
R1661 B.n819 B.n524 10.6151
R1662 B.n829 B.n524 10.6151
R1663 B.n830 B.n829 10.6151
R1664 B.n831 B.n830 10.6151
R1665 B.n831 B.n516 10.6151
R1666 B.n841 B.n516 10.6151
R1667 B.n842 B.n841 10.6151
R1668 B.n843 B.n842 10.6151
R1669 B.n843 B.n508 10.6151
R1670 B.n853 B.n508 10.6151
R1671 B.n854 B.n853 10.6151
R1672 B.n855 B.n854 10.6151
R1673 B.n855 B.n500 10.6151
R1674 B.n865 B.n500 10.6151
R1675 B.n866 B.n865 10.6151
R1676 B.n867 B.n866 10.6151
R1677 B.n867 B.n492 10.6151
R1678 B.n877 B.n492 10.6151
R1679 B.n878 B.n877 10.6151
R1680 B.n879 B.n878 10.6151
R1681 B.n879 B.n484 10.6151
R1682 B.n889 B.n484 10.6151
R1683 B.n890 B.n889 10.6151
R1684 B.n891 B.n890 10.6151
R1685 B.n891 B.n476 10.6151
R1686 B.n901 B.n476 10.6151
R1687 B.n902 B.n901 10.6151
R1688 B.n903 B.n902 10.6151
R1689 B.n903 B.n468 10.6151
R1690 B.n913 B.n468 10.6151
R1691 B.n914 B.n913 10.6151
R1692 B.n915 B.n914 10.6151
R1693 B.n915 B.n460 10.6151
R1694 B.n925 B.n460 10.6151
R1695 B.n926 B.n925 10.6151
R1696 B.n927 B.n926 10.6151
R1697 B.n927 B.n452 10.6151
R1698 B.n937 B.n452 10.6151
R1699 B.n938 B.n937 10.6151
R1700 B.n939 B.n938 10.6151
R1701 B.n939 B.n444 10.6151
R1702 B.n949 B.n444 10.6151
R1703 B.n950 B.n949 10.6151
R1704 B.n951 B.n950 10.6151
R1705 B.n951 B.n436 10.6151
R1706 B.n961 B.n436 10.6151
R1707 B.n962 B.n961 10.6151
R1708 B.n963 B.n962 10.6151
R1709 B.n963 B.n428 10.6151
R1710 B.n973 B.n428 10.6151
R1711 B.n974 B.n973 10.6151
R1712 B.n975 B.n974 10.6151
R1713 B.n975 B.n420 10.6151
R1714 B.n985 B.n420 10.6151
R1715 B.n986 B.n985 10.6151
R1716 B.n987 B.n986 10.6151
R1717 B.n987 B.n412 10.6151
R1718 B.n997 B.n412 10.6151
R1719 B.n998 B.n997 10.6151
R1720 B.n999 B.n998 10.6151
R1721 B.n999 B.n404 10.6151
R1722 B.n1010 B.n404 10.6151
R1723 B.n1011 B.n1010 10.6151
R1724 B.n1012 B.n1011 10.6151
R1725 B.n1012 B.n0 10.6151
R1726 B.n806 B.n805 10.6151
R1727 B.n805 B.n804 10.6151
R1728 B.n804 B.n803 10.6151
R1729 B.n803 B.n801 10.6151
R1730 B.n801 B.n798 10.6151
R1731 B.n798 B.n797 10.6151
R1732 B.n797 B.n794 10.6151
R1733 B.n794 B.n793 10.6151
R1734 B.n793 B.n790 10.6151
R1735 B.n790 B.n789 10.6151
R1736 B.n789 B.n786 10.6151
R1737 B.n786 B.n785 10.6151
R1738 B.n785 B.n782 10.6151
R1739 B.n782 B.n781 10.6151
R1740 B.n781 B.n778 10.6151
R1741 B.n778 B.n777 10.6151
R1742 B.n777 B.n774 10.6151
R1743 B.n774 B.n773 10.6151
R1744 B.n773 B.n770 10.6151
R1745 B.n770 B.n769 10.6151
R1746 B.n769 B.n766 10.6151
R1747 B.n766 B.n765 10.6151
R1748 B.n765 B.n762 10.6151
R1749 B.n762 B.n761 10.6151
R1750 B.n761 B.n758 10.6151
R1751 B.n758 B.n757 10.6151
R1752 B.n757 B.n754 10.6151
R1753 B.n754 B.n753 10.6151
R1754 B.n753 B.n750 10.6151
R1755 B.n750 B.n749 10.6151
R1756 B.n749 B.n746 10.6151
R1757 B.n746 B.n745 10.6151
R1758 B.n745 B.n742 10.6151
R1759 B.n742 B.n741 10.6151
R1760 B.n741 B.n738 10.6151
R1761 B.n738 B.n737 10.6151
R1762 B.n737 B.n734 10.6151
R1763 B.n734 B.n733 10.6151
R1764 B.n733 B.n730 10.6151
R1765 B.n730 B.n729 10.6151
R1766 B.n729 B.n726 10.6151
R1767 B.n726 B.n725 10.6151
R1768 B.n725 B.n722 10.6151
R1769 B.n722 B.n721 10.6151
R1770 B.n721 B.n718 10.6151
R1771 B.n718 B.n717 10.6151
R1772 B.n717 B.n714 10.6151
R1773 B.n714 B.n713 10.6151
R1774 B.n710 B.n709 10.6151
R1775 B.n709 B.n706 10.6151
R1776 B.n706 B.n705 10.6151
R1777 B.n705 B.n702 10.6151
R1778 B.n702 B.n701 10.6151
R1779 B.n701 B.n698 10.6151
R1780 B.n698 B.n697 10.6151
R1781 B.n697 B.n694 10.6151
R1782 B.n694 B.n693 10.6151
R1783 B.n690 B.n689 10.6151
R1784 B.n689 B.n686 10.6151
R1785 B.n686 B.n685 10.6151
R1786 B.n685 B.n682 10.6151
R1787 B.n682 B.n681 10.6151
R1788 B.n681 B.n678 10.6151
R1789 B.n678 B.n677 10.6151
R1790 B.n677 B.n674 10.6151
R1791 B.n674 B.n673 10.6151
R1792 B.n673 B.n670 10.6151
R1793 B.n670 B.n669 10.6151
R1794 B.n669 B.n666 10.6151
R1795 B.n666 B.n665 10.6151
R1796 B.n665 B.n662 10.6151
R1797 B.n662 B.n661 10.6151
R1798 B.n661 B.n658 10.6151
R1799 B.n658 B.n657 10.6151
R1800 B.n657 B.n654 10.6151
R1801 B.n654 B.n653 10.6151
R1802 B.n653 B.n650 10.6151
R1803 B.n650 B.n649 10.6151
R1804 B.n649 B.n646 10.6151
R1805 B.n646 B.n645 10.6151
R1806 B.n645 B.n642 10.6151
R1807 B.n642 B.n641 10.6151
R1808 B.n641 B.n638 10.6151
R1809 B.n638 B.n637 10.6151
R1810 B.n637 B.n634 10.6151
R1811 B.n634 B.n633 10.6151
R1812 B.n633 B.n630 10.6151
R1813 B.n630 B.n629 10.6151
R1814 B.n629 B.n626 10.6151
R1815 B.n626 B.n625 10.6151
R1816 B.n625 B.n622 10.6151
R1817 B.n622 B.n621 10.6151
R1818 B.n621 B.n618 10.6151
R1819 B.n618 B.n617 10.6151
R1820 B.n617 B.n614 10.6151
R1821 B.n614 B.n613 10.6151
R1822 B.n613 B.n610 10.6151
R1823 B.n610 B.n609 10.6151
R1824 B.n609 B.n606 10.6151
R1825 B.n606 B.n605 10.6151
R1826 B.n605 B.n602 10.6151
R1827 B.n602 B.n601 10.6151
R1828 B.n601 B.n598 10.6151
R1829 B.n598 B.n536 10.6151
R1830 B.n811 B.n536 10.6151
R1831 B.n813 B.n812 10.6151
R1832 B.n813 B.n528 10.6151
R1833 B.n823 B.n528 10.6151
R1834 B.n824 B.n823 10.6151
R1835 B.n825 B.n824 10.6151
R1836 B.n825 B.n520 10.6151
R1837 B.n835 B.n520 10.6151
R1838 B.n836 B.n835 10.6151
R1839 B.n837 B.n836 10.6151
R1840 B.n837 B.n512 10.6151
R1841 B.n847 B.n512 10.6151
R1842 B.n848 B.n847 10.6151
R1843 B.n849 B.n848 10.6151
R1844 B.n849 B.n504 10.6151
R1845 B.n859 B.n504 10.6151
R1846 B.n860 B.n859 10.6151
R1847 B.n861 B.n860 10.6151
R1848 B.n861 B.n496 10.6151
R1849 B.n871 B.n496 10.6151
R1850 B.n872 B.n871 10.6151
R1851 B.n873 B.n872 10.6151
R1852 B.n873 B.n487 10.6151
R1853 B.n883 B.n487 10.6151
R1854 B.n884 B.n883 10.6151
R1855 B.n885 B.n884 10.6151
R1856 B.n885 B.n480 10.6151
R1857 B.n895 B.n480 10.6151
R1858 B.n896 B.n895 10.6151
R1859 B.n897 B.n896 10.6151
R1860 B.n897 B.n472 10.6151
R1861 B.n907 B.n472 10.6151
R1862 B.n908 B.n907 10.6151
R1863 B.n909 B.n908 10.6151
R1864 B.n909 B.n464 10.6151
R1865 B.n919 B.n464 10.6151
R1866 B.n920 B.n919 10.6151
R1867 B.n921 B.n920 10.6151
R1868 B.n921 B.n456 10.6151
R1869 B.n931 B.n456 10.6151
R1870 B.n932 B.n931 10.6151
R1871 B.n933 B.n932 10.6151
R1872 B.n933 B.n448 10.6151
R1873 B.n943 B.n448 10.6151
R1874 B.n944 B.n943 10.6151
R1875 B.n945 B.n944 10.6151
R1876 B.n945 B.n440 10.6151
R1877 B.n955 B.n440 10.6151
R1878 B.n956 B.n955 10.6151
R1879 B.n957 B.n956 10.6151
R1880 B.n957 B.n432 10.6151
R1881 B.n967 B.n432 10.6151
R1882 B.n968 B.n967 10.6151
R1883 B.n969 B.n968 10.6151
R1884 B.n969 B.n424 10.6151
R1885 B.n979 B.n424 10.6151
R1886 B.n980 B.n979 10.6151
R1887 B.n981 B.n980 10.6151
R1888 B.n981 B.n416 10.6151
R1889 B.n991 B.n416 10.6151
R1890 B.n992 B.n991 10.6151
R1891 B.n993 B.n992 10.6151
R1892 B.n993 B.n408 10.6151
R1893 B.n1003 B.n408 10.6151
R1894 B.n1004 B.n1003 10.6151
R1895 B.n1006 B.n1004 10.6151
R1896 B.n1006 B.n1005 10.6151
R1897 B.n1005 B.n400 10.6151
R1898 B.n1017 B.n400 10.6151
R1899 B.n1018 B.n1017 10.6151
R1900 B.n1019 B.n1018 10.6151
R1901 B.n1020 B.n1019 10.6151
R1902 B.n1021 B.n1020 10.6151
R1903 B.n1024 B.n1021 10.6151
R1904 B.n1025 B.n1024 10.6151
R1905 B.n1026 B.n1025 10.6151
R1906 B.n1027 B.n1026 10.6151
R1907 B.n1029 B.n1027 10.6151
R1908 B.n1030 B.n1029 10.6151
R1909 B.n1031 B.n1030 10.6151
R1910 B.n1032 B.n1031 10.6151
R1911 B.n1034 B.n1032 10.6151
R1912 B.n1035 B.n1034 10.6151
R1913 B.n1036 B.n1035 10.6151
R1914 B.n1037 B.n1036 10.6151
R1915 B.n1039 B.n1037 10.6151
R1916 B.n1040 B.n1039 10.6151
R1917 B.n1041 B.n1040 10.6151
R1918 B.n1042 B.n1041 10.6151
R1919 B.n1044 B.n1042 10.6151
R1920 B.n1045 B.n1044 10.6151
R1921 B.n1046 B.n1045 10.6151
R1922 B.n1047 B.n1046 10.6151
R1923 B.n1049 B.n1047 10.6151
R1924 B.n1050 B.n1049 10.6151
R1925 B.n1051 B.n1050 10.6151
R1926 B.n1052 B.n1051 10.6151
R1927 B.n1054 B.n1052 10.6151
R1928 B.n1055 B.n1054 10.6151
R1929 B.n1056 B.n1055 10.6151
R1930 B.n1057 B.n1056 10.6151
R1931 B.n1059 B.n1057 10.6151
R1932 B.n1060 B.n1059 10.6151
R1933 B.n1061 B.n1060 10.6151
R1934 B.n1062 B.n1061 10.6151
R1935 B.n1064 B.n1062 10.6151
R1936 B.n1065 B.n1064 10.6151
R1937 B.n1066 B.n1065 10.6151
R1938 B.n1067 B.n1066 10.6151
R1939 B.n1069 B.n1067 10.6151
R1940 B.n1070 B.n1069 10.6151
R1941 B.n1071 B.n1070 10.6151
R1942 B.n1072 B.n1071 10.6151
R1943 B.n1074 B.n1072 10.6151
R1944 B.n1075 B.n1074 10.6151
R1945 B.n1076 B.n1075 10.6151
R1946 B.n1077 B.n1076 10.6151
R1947 B.n1079 B.n1077 10.6151
R1948 B.n1080 B.n1079 10.6151
R1949 B.n1081 B.n1080 10.6151
R1950 B.n1082 B.n1081 10.6151
R1951 B.n1084 B.n1082 10.6151
R1952 B.n1085 B.n1084 10.6151
R1953 B.n1086 B.n1085 10.6151
R1954 B.n1087 B.n1086 10.6151
R1955 B.n1089 B.n1087 10.6151
R1956 B.n1090 B.n1089 10.6151
R1957 B.n1091 B.n1090 10.6151
R1958 B.n1092 B.n1091 10.6151
R1959 B.n1094 B.n1092 10.6151
R1960 B.n1095 B.n1094 10.6151
R1961 B.n1096 B.n1095 10.6151
R1962 B.n1097 B.n1096 10.6151
R1963 B.n1099 B.n1097 10.6151
R1964 B.n1100 B.n1099 10.6151
R1965 B.n1101 B.n1100 10.6151
R1966 B.n1102 B.n1101 10.6151
R1967 B.n1104 B.n1102 10.6151
R1968 B.n1105 B.n1104 10.6151
R1969 B.n1106 B.n1105 10.6151
R1970 B.n1244 B.n1 10.6151
R1971 B.n1244 B.n1243 10.6151
R1972 B.n1243 B.n1242 10.6151
R1973 B.n1242 B.n10 10.6151
R1974 B.n1236 B.n10 10.6151
R1975 B.n1236 B.n1235 10.6151
R1976 B.n1235 B.n1234 10.6151
R1977 B.n1234 B.n18 10.6151
R1978 B.n1228 B.n18 10.6151
R1979 B.n1228 B.n1227 10.6151
R1980 B.n1227 B.n1226 10.6151
R1981 B.n1226 B.n25 10.6151
R1982 B.n1220 B.n25 10.6151
R1983 B.n1220 B.n1219 10.6151
R1984 B.n1219 B.n1218 10.6151
R1985 B.n1218 B.n32 10.6151
R1986 B.n1212 B.n32 10.6151
R1987 B.n1212 B.n1211 10.6151
R1988 B.n1211 B.n1210 10.6151
R1989 B.n1210 B.n39 10.6151
R1990 B.n1204 B.n39 10.6151
R1991 B.n1204 B.n1203 10.6151
R1992 B.n1203 B.n1202 10.6151
R1993 B.n1202 B.n46 10.6151
R1994 B.n1196 B.n46 10.6151
R1995 B.n1196 B.n1195 10.6151
R1996 B.n1195 B.n1194 10.6151
R1997 B.n1194 B.n53 10.6151
R1998 B.n1188 B.n53 10.6151
R1999 B.n1188 B.n1187 10.6151
R2000 B.n1187 B.n1186 10.6151
R2001 B.n1186 B.n60 10.6151
R2002 B.n1180 B.n60 10.6151
R2003 B.n1180 B.n1179 10.6151
R2004 B.n1179 B.n1178 10.6151
R2005 B.n1178 B.n67 10.6151
R2006 B.n1172 B.n67 10.6151
R2007 B.n1172 B.n1171 10.6151
R2008 B.n1171 B.n1170 10.6151
R2009 B.n1170 B.n74 10.6151
R2010 B.n1164 B.n74 10.6151
R2011 B.n1164 B.n1163 10.6151
R2012 B.n1163 B.n1162 10.6151
R2013 B.n1162 B.n81 10.6151
R2014 B.n1156 B.n81 10.6151
R2015 B.n1156 B.n1155 10.6151
R2016 B.n1155 B.n1154 10.6151
R2017 B.n1154 B.n88 10.6151
R2018 B.n1148 B.n88 10.6151
R2019 B.n1148 B.n1147 10.6151
R2020 B.n1147 B.n1146 10.6151
R2021 B.n1146 B.n95 10.6151
R2022 B.n1140 B.n95 10.6151
R2023 B.n1140 B.n1139 10.6151
R2024 B.n1139 B.n1138 10.6151
R2025 B.n1138 B.n102 10.6151
R2026 B.n1132 B.n102 10.6151
R2027 B.n1132 B.n1131 10.6151
R2028 B.n1131 B.n1130 10.6151
R2029 B.n1130 B.n109 10.6151
R2030 B.n1124 B.n109 10.6151
R2031 B.n1124 B.n1123 10.6151
R2032 B.n1123 B.n1122 10.6151
R2033 B.n1122 B.n116 10.6151
R2034 B.n1116 B.n116 10.6151
R2035 B.n1116 B.n1115 10.6151
R2036 B.n1115 B.n1114 10.6151
R2037 B.n1114 B.n123 10.6151
R2038 B.n187 B.n186 10.6151
R2039 B.n190 B.n187 10.6151
R2040 B.n191 B.n190 10.6151
R2041 B.n194 B.n191 10.6151
R2042 B.n195 B.n194 10.6151
R2043 B.n198 B.n195 10.6151
R2044 B.n199 B.n198 10.6151
R2045 B.n202 B.n199 10.6151
R2046 B.n203 B.n202 10.6151
R2047 B.n206 B.n203 10.6151
R2048 B.n207 B.n206 10.6151
R2049 B.n210 B.n207 10.6151
R2050 B.n211 B.n210 10.6151
R2051 B.n214 B.n211 10.6151
R2052 B.n215 B.n214 10.6151
R2053 B.n218 B.n215 10.6151
R2054 B.n219 B.n218 10.6151
R2055 B.n222 B.n219 10.6151
R2056 B.n223 B.n222 10.6151
R2057 B.n226 B.n223 10.6151
R2058 B.n227 B.n226 10.6151
R2059 B.n230 B.n227 10.6151
R2060 B.n231 B.n230 10.6151
R2061 B.n234 B.n231 10.6151
R2062 B.n235 B.n234 10.6151
R2063 B.n238 B.n235 10.6151
R2064 B.n239 B.n238 10.6151
R2065 B.n242 B.n239 10.6151
R2066 B.n243 B.n242 10.6151
R2067 B.n246 B.n243 10.6151
R2068 B.n247 B.n246 10.6151
R2069 B.n250 B.n247 10.6151
R2070 B.n251 B.n250 10.6151
R2071 B.n254 B.n251 10.6151
R2072 B.n255 B.n254 10.6151
R2073 B.n258 B.n255 10.6151
R2074 B.n259 B.n258 10.6151
R2075 B.n262 B.n259 10.6151
R2076 B.n263 B.n262 10.6151
R2077 B.n266 B.n263 10.6151
R2078 B.n267 B.n266 10.6151
R2079 B.n270 B.n267 10.6151
R2080 B.n271 B.n270 10.6151
R2081 B.n274 B.n271 10.6151
R2082 B.n275 B.n274 10.6151
R2083 B.n278 B.n275 10.6151
R2084 B.n279 B.n278 10.6151
R2085 B.n282 B.n279 10.6151
R2086 B.n287 B.n284 10.6151
R2087 B.n288 B.n287 10.6151
R2088 B.n291 B.n288 10.6151
R2089 B.n292 B.n291 10.6151
R2090 B.n295 B.n292 10.6151
R2091 B.n296 B.n295 10.6151
R2092 B.n299 B.n296 10.6151
R2093 B.n300 B.n299 10.6151
R2094 B.n303 B.n300 10.6151
R2095 B.n308 B.n305 10.6151
R2096 B.n309 B.n308 10.6151
R2097 B.n312 B.n309 10.6151
R2098 B.n313 B.n312 10.6151
R2099 B.n316 B.n313 10.6151
R2100 B.n317 B.n316 10.6151
R2101 B.n320 B.n317 10.6151
R2102 B.n321 B.n320 10.6151
R2103 B.n324 B.n321 10.6151
R2104 B.n325 B.n324 10.6151
R2105 B.n328 B.n325 10.6151
R2106 B.n329 B.n328 10.6151
R2107 B.n332 B.n329 10.6151
R2108 B.n333 B.n332 10.6151
R2109 B.n336 B.n333 10.6151
R2110 B.n337 B.n336 10.6151
R2111 B.n340 B.n337 10.6151
R2112 B.n341 B.n340 10.6151
R2113 B.n344 B.n341 10.6151
R2114 B.n345 B.n344 10.6151
R2115 B.n348 B.n345 10.6151
R2116 B.n349 B.n348 10.6151
R2117 B.n352 B.n349 10.6151
R2118 B.n353 B.n352 10.6151
R2119 B.n356 B.n353 10.6151
R2120 B.n357 B.n356 10.6151
R2121 B.n360 B.n357 10.6151
R2122 B.n361 B.n360 10.6151
R2123 B.n364 B.n361 10.6151
R2124 B.n365 B.n364 10.6151
R2125 B.n368 B.n365 10.6151
R2126 B.n369 B.n368 10.6151
R2127 B.n372 B.n369 10.6151
R2128 B.n373 B.n372 10.6151
R2129 B.n376 B.n373 10.6151
R2130 B.n377 B.n376 10.6151
R2131 B.n380 B.n377 10.6151
R2132 B.n381 B.n380 10.6151
R2133 B.n384 B.n381 10.6151
R2134 B.n385 B.n384 10.6151
R2135 B.n388 B.n385 10.6151
R2136 B.n389 B.n388 10.6151
R2137 B.n392 B.n389 10.6151
R2138 B.n393 B.n392 10.6151
R2139 B.n396 B.n393 10.6151
R2140 B.n398 B.n396 10.6151
R2141 B.n399 B.n398 10.6151
R2142 B.n1107 B.n399 10.6151
R2143 B.t1 B.n410 9.4093
R2144 B.t0 B.n16 9.4093
R2145 B.n713 B.n594 9.36635
R2146 B.n690 B.n597 9.36635
R2147 B.n283 B.n282 9.36635
R2148 B.n305 B.n304 9.36635
R2149 B.n1252 B.n0 8.11757
R2150 B.n1252 B.n1 8.11757
R2151 B.n923 B.t7 6.08855
R2152 B.n1184 B.t5 6.08855
R2153 B.n887 B.t4 4.98163
R2154 B.n1160 B.t6 4.98163
R2155 B.n710 B.n594 1.24928
R2156 B.n693 B.n597 1.24928
R2157 B.n284 B.n283 1.24928
R2158 B.n304 B.n303 1.24928
R2159 VP.n26 VP.n25 161.3
R2160 VP.n27 VP.n22 161.3
R2161 VP.n29 VP.n28 161.3
R2162 VP.n30 VP.n21 161.3
R2163 VP.n32 VP.n31 161.3
R2164 VP.n33 VP.n20 161.3
R2165 VP.n35 VP.n34 161.3
R2166 VP.n36 VP.n19 161.3
R2167 VP.n39 VP.n38 161.3
R2168 VP.n40 VP.n18 161.3
R2169 VP.n42 VP.n41 161.3
R2170 VP.n43 VP.n17 161.3
R2171 VP.n45 VP.n44 161.3
R2172 VP.n46 VP.n16 161.3
R2173 VP.n48 VP.n47 161.3
R2174 VP.n49 VP.n15 161.3
R2175 VP.n51 VP.n50 161.3
R2176 VP.n95 VP.n94 161.3
R2177 VP.n93 VP.n1 161.3
R2178 VP.n92 VP.n91 161.3
R2179 VP.n90 VP.n2 161.3
R2180 VP.n89 VP.n88 161.3
R2181 VP.n87 VP.n3 161.3
R2182 VP.n86 VP.n85 161.3
R2183 VP.n84 VP.n4 161.3
R2184 VP.n83 VP.n82 161.3
R2185 VP.n80 VP.n5 161.3
R2186 VP.n79 VP.n78 161.3
R2187 VP.n77 VP.n6 161.3
R2188 VP.n76 VP.n75 161.3
R2189 VP.n74 VP.n7 161.3
R2190 VP.n73 VP.n72 161.3
R2191 VP.n71 VP.n8 161.3
R2192 VP.n70 VP.n69 161.3
R2193 VP.n67 VP.n9 161.3
R2194 VP.n66 VP.n65 161.3
R2195 VP.n64 VP.n10 161.3
R2196 VP.n63 VP.n62 161.3
R2197 VP.n61 VP.n11 161.3
R2198 VP.n60 VP.n59 161.3
R2199 VP.n58 VP.n12 161.3
R2200 VP.n57 VP.n56 161.3
R2201 VP.n55 VP.n13 161.3
R2202 VP.n23 VP.t6 123.796
R2203 VP.n54 VP.t2 91.3927
R2204 VP.n68 VP.t7 91.3927
R2205 VP.n81 VP.t1 91.3927
R2206 VP.n0 VP.t4 91.3927
R2207 VP.n14 VP.t0 91.3927
R2208 VP.n37 VP.t3 91.3927
R2209 VP.n24 VP.t5 91.3927
R2210 VP.n54 VP.n53 89.2619
R2211 VP.n96 VP.n0 89.2619
R2212 VP.n52 VP.n14 89.2619
R2213 VP.n53 VP.n52 58.7495
R2214 VP.n24 VP.n23 58.6002
R2215 VP.n75 VP.n74 56.5617
R2216 VP.n31 VP.n30 56.5617
R2217 VP.n62 VP.n61 47.3584
R2218 VP.n88 VP.n87 47.3584
R2219 VP.n44 VP.n43 47.3584
R2220 VP.n61 VP.n60 33.7956
R2221 VP.n88 VP.n2 33.7956
R2222 VP.n44 VP.n16 33.7956
R2223 VP.n56 VP.n55 24.5923
R2224 VP.n56 VP.n12 24.5923
R2225 VP.n60 VP.n12 24.5923
R2226 VP.n62 VP.n10 24.5923
R2227 VP.n66 VP.n10 24.5923
R2228 VP.n67 VP.n66 24.5923
R2229 VP.n69 VP.n8 24.5923
R2230 VP.n73 VP.n8 24.5923
R2231 VP.n74 VP.n73 24.5923
R2232 VP.n75 VP.n6 24.5923
R2233 VP.n79 VP.n6 24.5923
R2234 VP.n80 VP.n79 24.5923
R2235 VP.n82 VP.n4 24.5923
R2236 VP.n86 VP.n4 24.5923
R2237 VP.n87 VP.n86 24.5923
R2238 VP.n92 VP.n2 24.5923
R2239 VP.n93 VP.n92 24.5923
R2240 VP.n94 VP.n93 24.5923
R2241 VP.n48 VP.n16 24.5923
R2242 VP.n49 VP.n48 24.5923
R2243 VP.n50 VP.n49 24.5923
R2244 VP.n31 VP.n20 24.5923
R2245 VP.n35 VP.n20 24.5923
R2246 VP.n36 VP.n35 24.5923
R2247 VP.n38 VP.n18 24.5923
R2248 VP.n42 VP.n18 24.5923
R2249 VP.n43 VP.n42 24.5923
R2250 VP.n25 VP.n22 24.5923
R2251 VP.n29 VP.n22 24.5923
R2252 VP.n30 VP.n29 24.5923
R2253 VP.n69 VP.n68 16.7229
R2254 VP.n81 VP.n80 16.7229
R2255 VP.n37 VP.n36 16.7229
R2256 VP.n25 VP.n24 16.7229
R2257 VP.n68 VP.n67 7.86989
R2258 VP.n82 VP.n81 7.86989
R2259 VP.n38 VP.n37 7.86989
R2260 VP.n26 VP.n23 2.49643
R2261 VP.n55 VP.n54 0.984173
R2262 VP.n94 VP.n0 0.984173
R2263 VP.n50 VP.n14 0.984173
R2264 VP.n52 VP.n51 0.354861
R2265 VP.n53 VP.n13 0.354861
R2266 VP.n96 VP.n95 0.354861
R2267 VP VP.n96 0.267071
R2268 VP.n27 VP.n26 0.189894
R2269 VP.n28 VP.n27 0.189894
R2270 VP.n28 VP.n21 0.189894
R2271 VP.n32 VP.n21 0.189894
R2272 VP.n33 VP.n32 0.189894
R2273 VP.n34 VP.n33 0.189894
R2274 VP.n34 VP.n19 0.189894
R2275 VP.n39 VP.n19 0.189894
R2276 VP.n40 VP.n39 0.189894
R2277 VP.n41 VP.n40 0.189894
R2278 VP.n41 VP.n17 0.189894
R2279 VP.n45 VP.n17 0.189894
R2280 VP.n46 VP.n45 0.189894
R2281 VP.n47 VP.n46 0.189894
R2282 VP.n47 VP.n15 0.189894
R2283 VP.n51 VP.n15 0.189894
R2284 VP.n57 VP.n13 0.189894
R2285 VP.n58 VP.n57 0.189894
R2286 VP.n59 VP.n58 0.189894
R2287 VP.n59 VP.n11 0.189894
R2288 VP.n63 VP.n11 0.189894
R2289 VP.n64 VP.n63 0.189894
R2290 VP.n65 VP.n64 0.189894
R2291 VP.n65 VP.n9 0.189894
R2292 VP.n70 VP.n9 0.189894
R2293 VP.n71 VP.n70 0.189894
R2294 VP.n72 VP.n71 0.189894
R2295 VP.n72 VP.n7 0.189894
R2296 VP.n76 VP.n7 0.189894
R2297 VP.n77 VP.n76 0.189894
R2298 VP.n78 VP.n77 0.189894
R2299 VP.n78 VP.n5 0.189894
R2300 VP.n83 VP.n5 0.189894
R2301 VP.n84 VP.n83 0.189894
R2302 VP.n85 VP.n84 0.189894
R2303 VP.n85 VP.n3 0.189894
R2304 VP.n89 VP.n3 0.189894
R2305 VP.n90 VP.n89 0.189894
R2306 VP.n91 VP.n90 0.189894
R2307 VP.n91 VP.n1 0.189894
R2308 VP.n95 VP.n1 0.189894
R2309 VTAIL.n11 VTAIL.t14 45.2741
R2310 VTAIL.n10 VTAIL.t1 45.2741
R2311 VTAIL.n7 VTAIL.t3 45.2741
R2312 VTAIL.n14 VTAIL.t8 45.2741
R2313 VTAIL.n15 VTAIL.t5 45.2739
R2314 VTAIL.n2 VTAIL.t0 45.2739
R2315 VTAIL.n3 VTAIL.t12 45.2739
R2316 VTAIL.n6 VTAIL.t10 45.2739
R2317 VTAIL.n13 VTAIL.n12 43.9179
R2318 VTAIL.n9 VTAIL.n8 43.9179
R2319 VTAIL.n1 VTAIL.n0 43.9179
R2320 VTAIL.n5 VTAIL.n4 43.9179
R2321 VTAIL.n15 VTAIL.n14 28.5565
R2322 VTAIL.n7 VTAIL.n6 28.5565
R2323 VTAIL.n9 VTAIL.n7 3.60395
R2324 VTAIL.n10 VTAIL.n9 3.60395
R2325 VTAIL.n13 VTAIL.n11 3.60395
R2326 VTAIL.n14 VTAIL.n13 3.60395
R2327 VTAIL.n6 VTAIL.n5 3.60395
R2328 VTAIL.n5 VTAIL.n3 3.60395
R2329 VTAIL.n2 VTAIL.n1 3.60395
R2330 VTAIL VTAIL.n15 3.54576
R2331 VTAIL.n0 VTAIL.t6 1.35666
R2332 VTAIL.n0 VTAIL.t4 1.35666
R2333 VTAIL.n4 VTAIL.t15 1.35666
R2334 VTAIL.n4 VTAIL.t9 1.35666
R2335 VTAIL.n12 VTAIL.t13 1.35666
R2336 VTAIL.n12 VTAIL.t11 1.35666
R2337 VTAIL.n8 VTAIL.t7 1.35666
R2338 VTAIL.n8 VTAIL.t2 1.35666
R2339 VTAIL.n11 VTAIL.n10 0.470328
R2340 VTAIL.n3 VTAIL.n2 0.470328
R2341 VTAIL VTAIL.n1 0.0586897
R2342 VDD1 VDD1.n0 62.4566
R2343 VDD1.n3 VDD1.n2 62.3431
R2344 VDD1.n3 VDD1.n1 62.3431
R2345 VDD1.n5 VDD1.n4 60.5967
R2346 VDD1.n5 VDD1.n3 53.1
R2347 VDD1 VDD1.n5 1.74403
R2348 VDD1.n4 VDD1.t4 1.35666
R2349 VDD1.n4 VDD1.t7 1.35666
R2350 VDD1.n0 VDD1.t1 1.35666
R2351 VDD1.n0 VDD1.t2 1.35666
R2352 VDD1.n2 VDD1.t6 1.35666
R2353 VDD1.n2 VDD1.t3 1.35666
R2354 VDD1.n1 VDD1.t5 1.35666
R2355 VDD1.n1 VDD1.t0 1.35666
R2356 VN.n76 VN.n75 161.3
R2357 VN.n74 VN.n40 161.3
R2358 VN.n73 VN.n72 161.3
R2359 VN.n71 VN.n41 161.3
R2360 VN.n70 VN.n69 161.3
R2361 VN.n68 VN.n42 161.3
R2362 VN.n67 VN.n66 161.3
R2363 VN.n65 VN.n43 161.3
R2364 VN.n64 VN.n63 161.3
R2365 VN.n61 VN.n44 161.3
R2366 VN.n60 VN.n59 161.3
R2367 VN.n58 VN.n45 161.3
R2368 VN.n57 VN.n56 161.3
R2369 VN.n55 VN.n46 161.3
R2370 VN.n54 VN.n53 161.3
R2371 VN.n52 VN.n47 161.3
R2372 VN.n51 VN.n50 161.3
R2373 VN.n37 VN.n36 161.3
R2374 VN.n35 VN.n1 161.3
R2375 VN.n34 VN.n33 161.3
R2376 VN.n32 VN.n2 161.3
R2377 VN.n31 VN.n30 161.3
R2378 VN.n29 VN.n3 161.3
R2379 VN.n28 VN.n27 161.3
R2380 VN.n26 VN.n4 161.3
R2381 VN.n25 VN.n24 161.3
R2382 VN.n22 VN.n5 161.3
R2383 VN.n21 VN.n20 161.3
R2384 VN.n19 VN.n6 161.3
R2385 VN.n18 VN.n17 161.3
R2386 VN.n16 VN.n7 161.3
R2387 VN.n15 VN.n14 161.3
R2388 VN.n13 VN.n8 161.3
R2389 VN.n12 VN.n11 161.3
R2390 VN.n48 VN.t3 123.796
R2391 VN.n9 VN.t5 123.796
R2392 VN.n10 VN.t2 91.3927
R2393 VN.n23 VN.t7 91.3927
R2394 VN.n0 VN.t6 91.3927
R2395 VN.n49 VN.t1 91.3927
R2396 VN.n62 VN.t4 91.3927
R2397 VN.n39 VN.t0 91.3927
R2398 VN.n38 VN.n0 89.2619
R2399 VN.n77 VN.n39 89.2619
R2400 VN VN.n77 58.9148
R2401 VN.n10 VN.n9 58.6002
R2402 VN.n49 VN.n48 58.6002
R2403 VN.n17 VN.n16 56.5617
R2404 VN.n56 VN.n55 56.5617
R2405 VN.n30 VN.n29 47.3584
R2406 VN.n69 VN.n68 47.3584
R2407 VN.n30 VN.n2 33.7956
R2408 VN.n69 VN.n41 33.7956
R2409 VN.n11 VN.n8 24.5923
R2410 VN.n15 VN.n8 24.5923
R2411 VN.n16 VN.n15 24.5923
R2412 VN.n17 VN.n6 24.5923
R2413 VN.n21 VN.n6 24.5923
R2414 VN.n22 VN.n21 24.5923
R2415 VN.n24 VN.n4 24.5923
R2416 VN.n28 VN.n4 24.5923
R2417 VN.n29 VN.n28 24.5923
R2418 VN.n34 VN.n2 24.5923
R2419 VN.n35 VN.n34 24.5923
R2420 VN.n36 VN.n35 24.5923
R2421 VN.n55 VN.n54 24.5923
R2422 VN.n54 VN.n47 24.5923
R2423 VN.n50 VN.n47 24.5923
R2424 VN.n68 VN.n67 24.5923
R2425 VN.n67 VN.n43 24.5923
R2426 VN.n63 VN.n43 24.5923
R2427 VN.n61 VN.n60 24.5923
R2428 VN.n60 VN.n45 24.5923
R2429 VN.n56 VN.n45 24.5923
R2430 VN.n75 VN.n74 24.5923
R2431 VN.n74 VN.n73 24.5923
R2432 VN.n73 VN.n41 24.5923
R2433 VN.n11 VN.n10 16.7229
R2434 VN.n23 VN.n22 16.7229
R2435 VN.n50 VN.n49 16.7229
R2436 VN.n62 VN.n61 16.7229
R2437 VN.n24 VN.n23 7.86989
R2438 VN.n63 VN.n62 7.86989
R2439 VN.n12 VN.n9 2.49644
R2440 VN.n51 VN.n48 2.49644
R2441 VN.n36 VN.n0 0.984173
R2442 VN.n75 VN.n39 0.984173
R2443 VN.n77 VN.n76 0.354861
R2444 VN.n38 VN.n37 0.354861
R2445 VN VN.n38 0.267071
R2446 VN.n76 VN.n40 0.189894
R2447 VN.n72 VN.n40 0.189894
R2448 VN.n72 VN.n71 0.189894
R2449 VN.n71 VN.n70 0.189894
R2450 VN.n70 VN.n42 0.189894
R2451 VN.n66 VN.n42 0.189894
R2452 VN.n66 VN.n65 0.189894
R2453 VN.n65 VN.n64 0.189894
R2454 VN.n64 VN.n44 0.189894
R2455 VN.n59 VN.n44 0.189894
R2456 VN.n59 VN.n58 0.189894
R2457 VN.n58 VN.n57 0.189894
R2458 VN.n57 VN.n46 0.189894
R2459 VN.n53 VN.n46 0.189894
R2460 VN.n53 VN.n52 0.189894
R2461 VN.n52 VN.n51 0.189894
R2462 VN.n13 VN.n12 0.189894
R2463 VN.n14 VN.n13 0.189894
R2464 VN.n14 VN.n7 0.189894
R2465 VN.n18 VN.n7 0.189894
R2466 VN.n19 VN.n18 0.189894
R2467 VN.n20 VN.n19 0.189894
R2468 VN.n20 VN.n5 0.189894
R2469 VN.n25 VN.n5 0.189894
R2470 VN.n26 VN.n25 0.189894
R2471 VN.n27 VN.n26 0.189894
R2472 VN.n27 VN.n3 0.189894
R2473 VN.n31 VN.n3 0.189894
R2474 VN.n32 VN.n31 0.189894
R2475 VN.n33 VN.n32 0.189894
R2476 VN.n33 VN.n1 0.189894
R2477 VN.n37 VN.n1 0.189894
R2478 VDD2.n2 VDD2.n1 62.3431
R2479 VDD2.n2 VDD2.n0 62.3431
R2480 VDD2 VDD2.n5 62.3403
R2481 VDD2.n4 VDD2.n3 60.5967
R2482 VDD2.n4 VDD2.n2 52.517
R2483 VDD2 VDD2.n4 1.86041
R2484 VDD2.n5 VDD2.t6 1.35666
R2485 VDD2.n5 VDD2.t4 1.35666
R2486 VDD2.n3 VDD2.t7 1.35666
R2487 VDD2.n3 VDD2.t3 1.35666
R2488 VDD2.n1 VDD2.t0 1.35666
R2489 VDD2.n1 VDD2.t1 1.35666
R2490 VDD2.n0 VDD2.t2 1.35666
R2491 VDD2.n0 VDD2.t5 1.35666
C0 VP VN 9.66664f
C1 VP VDD1 11.6822f
C2 VP VDD2 0.652814f
C3 VN VDD1 0.154117f
C4 VP VTAIL 11.8826f
C5 VN VDD2 11.1855f
C6 VDD1 VDD2 2.42493f
C7 VN VTAIL 11.868501f
C8 VTAIL VDD1 9.352309f
C9 VTAIL VDD2 9.41511f
C10 VDD2 B 6.84858f
C11 VDD1 B 7.423349f
C12 VTAIL B 12.901874f
C13 VN B 20.52042f
C14 VP B 19.165575f
C15 VDD2.t2 B 0.309506f
C16 VDD2.t5 B 0.309506f
C17 VDD2.n0 B 2.80613f
C18 VDD2.t0 B 0.309506f
C19 VDD2.t1 B 0.309506f
C20 VDD2.n1 B 2.80613f
C21 VDD2.n2 B 4.47975f
C22 VDD2.t7 B 0.309506f
C23 VDD2.t3 B 0.309506f
C24 VDD2.n3 B 2.78651f
C25 VDD2.n4 B 3.84768f
C26 VDD2.t6 B 0.309506f
C27 VDD2.t4 B 0.309506f
C28 VDD2.n5 B 2.80608f
C29 VN.t6 B 2.56464f
C30 VN.n0 B 0.951325f
C31 VN.n1 B 0.016661f
C32 VN.n2 B 0.033472f
C33 VN.n3 B 0.016661f
C34 VN.n4 B 0.030896f
C35 VN.n5 B 0.016661f
C36 VN.t7 B 2.56464f
C37 VN.n6 B 0.030896f
C38 VN.n7 B 0.016661f
C39 VN.n8 B 0.030896f
C40 VN.t5 B 2.83233f
C41 VN.n9 B 0.908471f
C42 VN.t2 B 2.56464f
C43 VN.n10 B 0.952665f
C44 VN.n11 B 0.026015f
C45 VN.n12 B 0.21566f
C46 VN.n13 B 0.016661f
C47 VN.n14 B 0.016661f
C48 VN.n15 B 0.030896f
C49 VN.n16 B 0.024219f
C50 VN.n17 B 0.024219f
C51 VN.n18 B 0.016661f
C52 VN.n19 B 0.016661f
C53 VN.n20 B 0.016661f
C54 VN.n21 B 0.030896f
C55 VN.n22 B 0.026015f
C56 VN.n23 B 0.890107f
C57 VN.n24 B 0.020524f
C58 VN.n25 B 0.016661f
C59 VN.n26 B 0.016661f
C60 VN.n27 B 0.016661f
C61 VN.n28 B 0.030896f
C62 VN.n29 B 0.031336f
C63 VN.n30 B 0.014527f
C64 VN.n31 B 0.016661f
C65 VN.n32 B 0.016661f
C66 VN.n33 B 0.016661f
C67 VN.n34 B 0.030896f
C68 VN.n35 B 0.030896f
C69 VN.n36 B 0.016254f
C70 VN.n37 B 0.026886f
C71 VN.n38 B 0.05249f
C72 VN.t0 B 2.56464f
C73 VN.n39 B 0.951325f
C74 VN.n40 B 0.016661f
C75 VN.n41 B 0.033472f
C76 VN.n42 B 0.016661f
C77 VN.n43 B 0.030896f
C78 VN.n44 B 0.016661f
C79 VN.t4 B 2.56464f
C80 VN.n45 B 0.030896f
C81 VN.n46 B 0.016661f
C82 VN.n47 B 0.030896f
C83 VN.t3 B 2.83233f
C84 VN.n48 B 0.908471f
C85 VN.t1 B 2.56464f
C86 VN.n49 B 0.952665f
C87 VN.n50 B 0.026015f
C88 VN.n51 B 0.21566f
C89 VN.n52 B 0.016661f
C90 VN.n53 B 0.016661f
C91 VN.n54 B 0.030896f
C92 VN.n55 B 0.024219f
C93 VN.n56 B 0.024219f
C94 VN.n57 B 0.016661f
C95 VN.n58 B 0.016661f
C96 VN.n59 B 0.016661f
C97 VN.n60 B 0.030896f
C98 VN.n61 B 0.026015f
C99 VN.n62 B 0.890107f
C100 VN.n63 B 0.020524f
C101 VN.n64 B 0.016661f
C102 VN.n65 B 0.016661f
C103 VN.n66 B 0.016661f
C104 VN.n67 B 0.030896f
C105 VN.n68 B 0.031336f
C106 VN.n69 B 0.014527f
C107 VN.n70 B 0.016661f
C108 VN.n71 B 0.016661f
C109 VN.n72 B 0.016661f
C110 VN.n73 B 0.030896f
C111 VN.n74 B 0.030896f
C112 VN.n75 B 0.016254f
C113 VN.n76 B 0.026886f
C114 VN.n77 B 1.2046f
C115 VDD1.t1 B 0.314878f
C116 VDD1.t2 B 0.314878f
C117 VDD1.n0 B 2.85638f
C118 VDD1.t5 B 0.314878f
C119 VDD1.t0 B 0.314878f
C120 VDD1.n1 B 2.85484f
C121 VDD1.t6 B 0.314878f
C122 VDD1.t3 B 0.314878f
C123 VDD1.n2 B 2.85484f
C124 VDD1.n3 B 4.61356f
C125 VDD1.t4 B 0.314878f
C126 VDD1.t7 B 0.314878f
C127 VDD1.n4 B 2.83487f
C128 VDD1.n5 B 3.94898f
C129 VTAIL.t6 B 0.2307f
C130 VTAIL.t4 B 0.2307f
C131 VTAIL.n0 B 2.01427f
C132 VTAIL.n1 B 0.440496f
C133 VTAIL.t0 B 2.57117f
C134 VTAIL.n2 B 0.539299f
C135 VTAIL.t12 B 2.57117f
C136 VTAIL.n3 B 0.539299f
C137 VTAIL.t15 B 0.2307f
C138 VTAIL.t9 B 0.2307f
C139 VTAIL.n4 B 2.01427f
C140 VTAIL.n5 B 0.668921f
C141 VTAIL.t10 B 2.57117f
C142 VTAIL.n6 B 1.82377f
C143 VTAIL.t3 B 2.57118f
C144 VTAIL.n7 B 1.82376f
C145 VTAIL.t7 B 0.2307f
C146 VTAIL.t2 B 0.2307f
C147 VTAIL.n8 B 2.01427f
C148 VTAIL.n9 B 0.668922f
C149 VTAIL.t1 B 2.57118f
C150 VTAIL.n10 B 0.539293f
C151 VTAIL.t14 B 2.57118f
C152 VTAIL.n11 B 0.539293f
C153 VTAIL.t13 B 0.2307f
C154 VTAIL.t11 B 0.2307f
C155 VTAIL.n12 B 2.01427f
C156 VTAIL.n13 B 0.668922f
C157 VTAIL.t8 B 2.57118f
C158 VTAIL.n14 B 1.82376f
C159 VTAIL.t5 B 2.57117f
C160 VTAIL.n15 B 1.82002f
C161 VP.t4 B 2.6056f
C162 VP.n0 B 0.966517f
C163 VP.n1 B 0.016927f
C164 VP.n2 B 0.034006f
C165 VP.n3 B 0.016927f
C166 VP.n4 B 0.03139f
C167 VP.n5 B 0.016927f
C168 VP.t1 B 2.6056f
C169 VP.n6 B 0.03139f
C170 VP.n7 B 0.016927f
C171 VP.n8 B 0.03139f
C172 VP.n9 B 0.016927f
C173 VP.t7 B 2.6056f
C174 VP.n10 B 0.03139f
C175 VP.n11 B 0.016927f
C176 VP.n12 B 0.03139f
C177 VP.n13 B 0.027316f
C178 VP.t2 B 2.6056f
C179 VP.t0 B 2.6056f
C180 VP.n14 B 0.966517f
C181 VP.n15 B 0.016927f
C182 VP.n16 B 0.034006f
C183 VP.n17 B 0.016927f
C184 VP.n18 B 0.03139f
C185 VP.n19 B 0.016927f
C186 VP.t3 B 2.6056f
C187 VP.n20 B 0.03139f
C188 VP.n21 B 0.016927f
C189 VP.n22 B 0.03139f
C190 VP.t6 B 2.87756f
C191 VP.n23 B 0.922979f
C192 VP.t5 B 2.6056f
C193 VP.n24 B 0.967878f
C194 VP.n25 B 0.026431f
C195 VP.n26 B 0.219104f
C196 VP.n27 B 0.016927f
C197 VP.n28 B 0.016927f
C198 VP.n29 B 0.03139f
C199 VP.n30 B 0.024606f
C200 VP.n31 B 0.024606f
C201 VP.n32 B 0.016927f
C202 VP.n33 B 0.016927f
C203 VP.n34 B 0.016927f
C204 VP.n35 B 0.03139f
C205 VP.n36 B 0.026431f
C206 VP.n37 B 0.904322f
C207 VP.n38 B 0.020852f
C208 VP.n39 B 0.016927f
C209 VP.n40 B 0.016927f
C210 VP.n41 B 0.016927f
C211 VP.n42 B 0.03139f
C212 VP.n43 B 0.031837f
C213 VP.n44 B 0.014759f
C214 VP.n45 B 0.016927f
C215 VP.n46 B 0.016927f
C216 VP.n47 B 0.016927f
C217 VP.n48 B 0.03139f
C218 VP.n49 B 0.03139f
C219 VP.n50 B 0.016513f
C220 VP.n51 B 0.027316f
C221 VP.n52 B 1.21727f
C222 VP.n53 B 1.22765f
C223 VP.n54 B 0.966517f
C224 VP.n55 B 0.016513f
C225 VP.n56 B 0.03139f
C226 VP.n57 B 0.016927f
C227 VP.n58 B 0.016927f
C228 VP.n59 B 0.016927f
C229 VP.n60 B 0.034006f
C230 VP.n61 B 0.014759f
C231 VP.n62 B 0.031837f
C232 VP.n63 B 0.016927f
C233 VP.n64 B 0.016927f
C234 VP.n65 B 0.016927f
C235 VP.n66 B 0.03139f
C236 VP.n67 B 0.020852f
C237 VP.n68 B 0.904322f
C238 VP.n69 B 0.026431f
C239 VP.n70 B 0.016927f
C240 VP.n71 B 0.016927f
C241 VP.n72 B 0.016927f
C242 VP.n73 B 0.03139f
C243 VP.n74 B 0.024606f
C244 VP.n75 B 0.024606f
C245 VP.n76 B 0.016927f
C246 VP.n77 B 0.016927f
C247 VP.n78 B 0.016927f
C248 VP.n79 B 0.03139f
C249 VP.n80 B 0.026431f
C250 VP.n81 B 0.904322f
C251 VP.n82 B 0.020852f
C252 VP.n83 B 0.016927f
C253 VP.n84 B 0.016927f
C254 VP.n85 B 0.016927f
C255 VP.n86 B 0.03139f
C256 VP.n87 B 0.031837f
C257 VP.n88 B 0.014759f
C258 VP.n89 B 0.016927f
C259 VP.n90 B 0.016927f
C260 VP.n91 B 0.016927f
C261 VP.n92 B 0.03139f
C262 VP.n93 B 0.03139f
C263 VP.n94 B 0.016513f
C264 VP.n95 B 0.027316f
C265 VP.n96 B 0.053328f
.ends

