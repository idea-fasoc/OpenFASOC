* NGSPICE file created from diff_pair_sample_0720.ext - technology: sky130A

.subckt diff_pair_sample_0720 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.72745 pd=16.86 as=2.72745 ps=16.86 w=16.53 l=3.73
X1 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=6.4467 pd=33.84 as=0 ps=0 w=16.53 l=3.73
X2 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4467 pd=33.84 as=2.72745 ps=16.86 w=16.53 l=3.73
X3 VDD2.t4 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.4467 pd=33.84 as=2.72745 ps=16.86 w=16.53 l=3.73
X4 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=6.4467 pd=33.84 as=0 ps=0 w=16.53 l=3.73
X5 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=6.4467 pd=33.84 as=0 ps=0 w=16.53 l=3.73
X6 VDD1.t4 VP.t1 VTAIL.t10 B.t0 sky130_fd_pr__nfet_01v8 ad=2.72745 pd=16.86 as=6.4467 ps=33.84 w=16.53 l=3.73
X7 VTAIL.t1 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.72745 pd=16.86 as=2.72745 ps=16.86 w=16.53 l=3.73
X8 VDD1.t3 VP.t2 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=6.4467 pd=33.84 as=2.72745 ps=16.86 w=16.53 l=3.73
X9 VTAIL.t4 VN.t3 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.72745 pd=16.86 as=2.72745 ps=16.86 w=16.53 l=3.73
X10 VDD2.t1 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.72745 pd=16.86 as=6.4467 ps=33.84 w=16.53 l=3.73
X11 VTAIL.t8 VP.t3 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.72745 pd=16.86 as=2.72745 ps=16.86 w=16.53 l=3.73
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.4467 pd=33.84 as=0 ps=0 w=16.53 l=3.73
X13 VDD1.t0 VP.t4 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.72745 pd=16.86 as=6.4467 ps=33.84 w=16.53 l=3.73
X14 VDD2.t0 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.72745 pd=16.86 as=6.4467 ps=33.84 w=16.53 l=3.73
X15 VDD1.t1 VP.t5 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=6.4467 pd=33.84 as=2.72745 ps=16.86 w=16.53 l=3.73
R0 VP.n16 VP.n13 161.3
R1 VP.n18 VP.n17 161.3
R2 VP.n19 VP.n12 161.3
R3 VP.n21 VP.n20 161.3
R4 VP.n22 VP.n11 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n10 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n56 VP.n55 161.3
R9 VP.n54 VP.n1 161.3
R10 VP.n53 VP.n52 161.3
R11 VP.n51 VP.n2 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n48 VP.n3 161.3
R14 VP.n47 VP.n46 161.3
R15 VP.n45 VP.n4 161.3
R16 VP.n44 VP.n43 161.3
R17 VP.n42 VP.n5 161.3
R18 VP.n41 VP.n40 161.3
R19 VP.n39 VP.n6 161.3
R20 VP.n38 VP.n37 161.3
R21 VP.n36 VP.n7 161.3
R22 VP.n35 VP.n34 161.3
R23 VP.n33 VP.n8 161.3
R24 VP.n32 VP.n31 161.3
R25 VP.n15 VP.t2 139.721
R26 VP.n43 VP.t3 106.802
R27 VP.n30 VP.t5 106.802
R28 VP.n0 VP.t1 106.802
R29 VP.n14 VP.t0 106.802
R30 VP.n9 VP.t4 106.802
R31 VP.n30 VP.n29 87.1314
R32 VP.n57 VP.n0 87.1314
R33 VP.n28 VP.n9 87.1314
R34 VP.n29 VP.n28 56.5751
R35 VP.n15 VP.n14 50.484
R36 VP.n37 VP.n36 43.4072
R37 VP.n49 VP.n2 43.4072
R38 VP.n20 VP.n11 43.4072
R39 VP.n37 VP.n6 37.5796
R40 VP.n49 VP.n48 37.5796
R41 VP.n20 VP.n19 37.5796
R42 VP.n31 VP.n8 24.4675
R43 VP.n35 VP.n8 24.4675
R44 VP.n36 VP.n35 24.4675
R45 VP.n41 VP.n6 24.4675
R46 VP.n42 VP.n41 24.4675
R47 VP.n43 VP.n42 24.4675
R48 VP.n43 VP.n4 24.4675
R49 VP.n47 VP.n4 24.4675
R50 VP.n48 VP.n47 24.4675
R51 VP.n53 VP.n2 24.4675
R52 VP.n54 VP.n53 24.4675
R53 VP.n55 VP.n54 24.4675
R54 VP.n24 VP.n11 24.4675
R55 VP.n25 VP.n24 24.4675
R56 VP.n26 VP.n25 24.4675
R57 VP.n14 VP.n13 24.4675
R58 VP.n18 VP.n13 24.4675
R59 VP.n19 VP.n18 24.4675
R60 VP.n31 VP.n30 2.93654
R61 VP.n55 VP.n0 2.93654
R62 VP.n26 VP.n9 2.93654
R63 VP.n16 VP.n15 2.46264
R64 VP.n28 VP.n27 0.354971
R65 VP.n32 VP.n29 0.354971
R66 VP.n57 VP.n56 0.354971
R67 VP VP.n57 0.26696
R68 VP.n17 VP.n16 0.189894
R69 VP.n17 VP.n12 0.189894
R70 VP.n21 VP.n12 0.189894
R71 VP.n22 VP.n21 0.189894
R72 VP.n23 VP.n22 0.189894
R73 VP.n23 VP.n10 0.189894
R74 VP.n27 VP.n10 0.189894
R75 VP.n33 VP.n32 0.189894
R76 VP.n34 VP.n33 0.189894
R77 VP.n34 VP.n7 0.189894
R78 VP.n38 VP.n7 0.189894
R79 VP.n39 VP.n38 0.189894
R80 VP.n40 VP.n39 0.189894
R81 VP.n40 VP.n5 0.189894
R82 VP.n44 VP.n5 0.189894
R83 VP.n45 VP.n44 0.189894
R84 VP.n46 VP.n45 0.189894
R85 VP.n46 VP.n3 0.189894
R86 VP.n50 VP.n3 0.189894
R87 VP.n51 VP.n50 0.189894
R88 VP.n52 VP.n51 0.189894
R89 VP.n52 VP.n1 0.189894
R90 VP.n56 VP.n1 0.189894
R91 VDD1 VDD1.t3 66.3761
R92 VDD1.n1 VDD1.t1 66.2623
R93 VDD1.n1 VDD1.n0 63.3145
R94 VDD1.n3 VDD1.n2 62.4949
R95 VDD1.n3 VDD1.n1 51.6733
R96 VDD1.n2 VDD1.t2 1.19832
R97 VDD1.n2 VDD1.t0 1.19832
R98 VDD1.n0 VDD1.t5 1.19832
R99 VDD1.n0 VDD1.t4 1.19832
R100 VDD1 VDD1.n3 0.81731
R101 VTAIL.n7 VTAIL.t0 47.0141
R102 VTAIL.n11 VTAIL.t5 47.0139
R103 VTAIL.n2 VTAIL.t10 47.0139
R104 VTAIL.n10 VTAIL.t7 47.0139
R105 VTAIL.n9 VTAIL.n8 45.8163
R106 VTAIL.n6 VTAIL.n5 45.8163
R107 VTAIL.n1 VTAIL.n0 45.8161
R108 VTAIL.n4 VTAIL.n3 45.8161
R109 VTAIL.n6 VTAIL.n4 33.6169
R110 VTAIL.n11 VTAIL.n10 30.1169
R111 VTAIL.n7 VTAIL.n6 3.5005
R112 VTAIL.n10 VTAIL.n9 3.5005
R113 VTAIL.n4 VTAIL.n2 3.5005
R114 VTAIL VTAIL.n11 2.56731
R115 VTAIL.n9 VTAIL.n7 2.22033
R116 VTAIL.n2 VTAIL.n1 2.22033
R117 VTAIL.n0 VTAIL.t3 1.19832
R118 VTAIL.n0 VTAIL.t4 1.19832
R119 VTAIL.n3 VTAIL.t6 1.19832
R120 VTAIL.n3 VTAIL.t8 1.19832
R121 VTAIL.n8 VTAIL.t9 1.19832
R122 VTAIL.n8 VTAIL.t11 1.19832
R123 VTAIL.n5 VTAIL.t2 1.19832
R124 VTAIL.n5 VTAIL.t1 1.19832
R125 VTAIL VTAIL.n1 0.93369
R126 B.n1056 B.n1055 585
R127 B.n1057 B.n1056 585
R128 B.n402 B.n163 585
R129 B.n401 B.n400 585
R130 B.n399 B.n398 585
R131 B.n397 B.n396 585
R132 B.n395 B.n394 585
R133 B.n393 B.n392 585
R134 B.n391 B.n390 585
R135 B.n389 B.n388 585
R136 B.n387 B.n386 585
R137 B.n385 B.n384 585
R138 B.n383 B.n382 585
R139 B.n381 B.n380 585
R140 B.n379 B.n378 585
R141 B.n377 B.n376 585
R142 B.n375 B.n374 585
R143 B.n373 B.n372 585
R144 B.n371 B.n370 585
R145 B.n369 B.n368 585
R146 B.n367 B.n366 585
R147 B.n365 B.n364 585
R148 B.n363 B.n362 585
R149 B.n361 B.n360 585
R150 B.n359 B.n358 585
R151 B.n357 B.n356 585
R152 B.n355 B.n354 585
R153 B.n353 B.n352 585
R154 B.n351 B.n350 585
R155 B.n349 B.n348 585
R156 B.n347 B.n346 585
R157 B.n345 B.n344 585
R158 B.n343 B.n342 585
R159 B.n341 B.n340 585
R160 B.n339 B.n338 585
R161 B.n337 B.n336 585
R162 B.n335 B.n334 585
R163 B.n333 B.n332 585
R164 B.n331 B.n330 585
R165 B.n329 B.n328 585
R166 B.n327 B.n326 585
R167 B.n325 B.n324 585
R168 B.n323 B.n322 585
R169 B.n321 B.n320 585
R170 B.n319 B.n318 585
R171 B.n317 B.n316 585
R172 B.n315 B.n314 585
R173 B.n313 B.n312 585
R174 B.n311 B.n310 585
R175 B.n309 B.n308 585
R176 B.n307 B.n306 585
R177 B.n305 B.n304 585
R178 B.n303 B.n302 585
R179 B.n301 B.n300 585
R180 B.n299 B.n298 585
R181 B.n297 B.n296 585
R182 B.n295 B.n294 585
R183 B.n293 B.n292 585
R184 B.n291 B.n290 585
R185 B.n289 B.n288 585
R186 B.n287 B.n286 585
R187 B.n285 B.n284 585
R188 B.n283 B.n282 585
R189 B.n281 B.n280 585
R190 B.n279 B.n278 585
R191 B.n276 B.n275 585
R192 B.n274 B.n273 585
R193 B.n272 B.n271 585
R194 B.n270 B.n269 585
R195 B.n268 B.n267 585
R196 B.n266 B.n265 585
R197 B.n264 B.n263 585
R198 B.n262 B.n261 585
R199 B.n260 B.n259 585
R200 B.n258 B.n257 585
R201 B.n256 B.n255 585
R202 B.n254 B.n253 585
R203 B.n252 B.n251 585
R204 B.n250 B.n249 585
R205 B.n248 B.n247 585
R206 B.n246 B.n245 585
R207 B.n244 B.n243 585
R208 B.n242 B.n241 585
R209 B.n240 B.n239 585
R210 B.n238 B.n237 585
R211 B.n236 B.n235 585
R212 B.n234 B.n233 585
R213 B.n232 B.n231 585
R214 B.n230 B.n229 585
R215 B.n228 B.n227 585
R216 B.n226 B.n225 585
R217 B.n224 B.n223 585
R218 B.n222 B.n221 585
R219 B.n220 B.n219 585
R220 B.n218 B.n217 585
R221 B.n216 B.n215 585
R222 B.n214 B.n213 585
R223 B.n212 B.n211 585
R224 B.n210 B.n209 585
R225 B.n208 B.n207 585
R226 B.n206 B.n205 585
R227 B.n204 B.n203 585
R228 B.n202 B.n201 585
R229 B.n200 B.n199 585
R230 B.n198 B.n197 585
R231 B.n196 B.n195 585
R232 B.n194 B.n193 585
R233 B.n192 B.n191 585
R234 B.n190 B.n189 585
R235 B.n188 B.n187 585
R236 B.n186 B.n185 585
R237 B.n184 B.n183 585
R238 B.n182 B.n181 585
R239 B.n180 B.n179 585
R240 B.n178 B.n177 585
R241 B.n176 B.n175 585
R242 B.n174 B.n173 585
R243 B.n172 B.n171 585
R244 B.n170 B.n169 585
R245 B.n102 B.n101 585
R246 B.n1054 B.n103 585
R247 B.n1058 B.n103 585
R248 B.n1053 B.n1052 585
R249 B.n1052 B.n99 585
R250 B.n1051 B.n98 585
R251 B.n1064 B.n98 585
R252 B.n1050 B.n97 585
R253 B.n1065 B.n97 585
R254 B.n1049 B.n96 585
R255 B.n1066 B.n96 585
R256 B.n1048 B.n1047 585
R257 B.n1047 B.n92 585
R258 B.n1046 B.n91 585
R259 B.n1072 B.n91 585
R260 B.n1045 B.n90 585
R261 B.n1073 B.n90 585
R262 B.n1044 B.n89 585
R263 B.n1074 B.n89 585
R264 B.n1043 B.n1042 585
R265 B.n1042 B.n88 585
R266 B.n1041 B.n84 585
R267 B.n1080 B.n84 585
R268 B.n1040 B.n83 585
R269 B.n1081 B.n83 585
R270 B.n1039 B.n82 585
R271 B.n1082 B.n82 585
R272 B.n1038 B.n1037 585
R273 B.n1037 B.n78 585
R274 B.n1036 B.n77 585
R275 B.n1088 B.n77 585
R276 B.n1035 B.n76 585
R277 B.n1089 B.n76 585
R278 B.n1034 B.n75 585
R279 B.n1090 B.n75 585
R280 B.n1033 B.n1032 585
R281 B.n1032 B.n71 585
R282 B.n1031 B.n70 585
R283 B.n1096 B.n70 585
R284 B.n1030 B.n69 585
R285 B.n1097 B.n69 585
R286 B.n1029 B.n68 585
R287 B.n1098 B.n68 585
R288 B.n1028 B.n1027 585
R289 B.n1027 B.n64 585
R290 B.n1026 B.n63 585
R291 B.n1104 B.n63 585
R292 B.n1025 B.n62 585
R293 B.n1105 B.n62 585
R294 B.n1024 B.n61 585
R295 B.n1106 B.n61 585
R296 B.n1023 B.n1022 585
R297 B.n1022 B.n57 585
R298 B.n1021 B.n56 585
R299 B.n1112 B.n56 585
R300 B.n1020 B.n55 585
R301 B.n1113 B.n55 585
R302 B.n1019 B.n54 585
R303 B.n1114 B.n54 585
R304 B.n1018 B.n1017 585
R305 B.n1017 B.n50 585
R306 B.n1016 B.n49 585
R307 B.n1120 B.n49 585
R308 B.n1015 B.n48 585
R309 B.n1121 B.n48 585
R310 B.n1014 B.n47 585
R311 B.n1122 B.n47 585
R312 B.n1013 B.n1012 585
R313 B.n1012 B.n43 585
R314 B.n1011 B.n42 585
R315 B.n1128 B.n42 585
R316 B.n1010 B.n41 585
R317 B.n1129 B.n41 585
R318 B.n1009 B.n40 585
R319 B.n1130 B.n40 585
R320 B.n1008 B.n1007 585
R321 B.n1007 B.n36 585
R322 B.n1006 B.n35 585
R323 B.n1136 B.n35 585
R324 B.n1005 B.n34 585
R325 B.n1137 B.n34 585
R326 B.n1004 B.n33 585
R327 B.n1138 B.n33 585
R328 B.n1003 B.n1002 585
R329 B.n1002 B.n29 585
R330 B.n1001 B.n28 585
R331 B.n1144 B.n28 585
R332 B.n1000 B.n27 585
R333 B.n1145 B.n27 585
R334 B.n999 B.n26 585
R335 B.n1146 B.n26 585
R336 B.n998 B.n997 585
R337 B.n997 B.n22 585
R338 B.n996 B.n21 585
R339 B.n1152 B.n21 585
R340 B.n995 B.n20 585
R341 B.n1153 B.n20 585
R342 B.n994 B.n19 585
R343 B.n1154 B.n19 585
R344 B.n993 B.n992 585
R345 B.n992 B.n15 585
R346 B.n991 B.n14 585
R347 B.n1160 B.n14 585
R348 B.n990 B.n13 585
R349 B.n1161 B.n13 585
R350 B.n989 B.n12 585
R351 B.n1162 B.n12 585
R352 B.n988 B.n987 585
R353 B.n987 B.n8 585
R354 B.n986 B.n7 585
R355 B.n1168 B.n7 585
R356 B.n985 B.n6 585
R357 B.n1169 B.n6 585
R358 B.n984 B.n5 585
R359 B.n1170 B.n5 585
R360 B.n983 B.n982 585
R361 B.n982 B.n4 585
R362 B.n981 B.n403 585
R363 B.n981 B.n980 585
R364 B.n971 B.n404 585
R365 B.n405 B.n404 585
R366 B.n973 B.n972 585
R367 B.n974 B.n973 585
R368 B.n970 B.n410 585
R369 B.n410 B.n409 585
R370 B.n969 B.n968 585
R371 B.n968 B.n967 585
R372 B.n412 B.n411 585
R373 B.n413 B.n412 585
R374 B.n960 B.n959 585
R375 B.n961 B.n960 585
R376 B.n958 B.n418 585
R377 B.n418 B.n417 585
R378 B.n957 B.n956 585
R379 B.n956 B.n955 585
R380 B.n420 B.n419 585
R381 B.n421 B.n420 585
R382 B.n948 B.n947 585
R383 B.n949 B.n948 585
R384 B.n946 B.n426 585
R385 B.n426 B.n425 585
R386 B.n945 B.n944 585
R387 B.n944 B.n943 585
R388 B.n428 B.n427 585
R389 B.n429 B.n428 585
R390 B.n936 B.n935 585
R391 B.n937 B.n936 585
R392 B.n934 B.n434 585
R393 B.n434 B.n433 585
R394 B.n933 B.n932 585
R395 B.n932 B.n931 585
R396 B.n436 B.n435 585
R397 B.n437 B.n436 585
R398 B.n924 B.n923 585
R399 B.n925 B.n924 585
R400 B.n922 B.n442 585
R401 B.n442 B.n441 585
R402 B.n921 B.n920 585
R403 B.n920 B.n919 585
R404 B.n444 B.n443 585
R405 B.n445 B.n444 585
R406 B.n912 B.n911 585
R407 B.n913 B.n912 585
R408 B.n910 B.n450 585
R409 B.n450 B.n449 585
R410 B.n909 B.n908 585
R411 B.n908 B.n907 585
R412 B.n452 B.n451 585
R413 B.n453 B.n452 585
R414 B.n900 B.n899 585
R415 B.n901 B.n900 585
R416 B.n898 B.n458 585
R417 B.n458 B.n457 585
R418 B.n897 B.n896 585
R419 B.n896 B.n895 585
R420 B.n460 B.n459 585
R421 B.n461 B.n460 585
R422 B.n888 B.n887 585
R423 B.n889 B.n888 585
R424 B.n886 B.n466 585
R425 B.n466 B.n465 585
R426 B.n885 B.n884 585
R427 B.n884 B.n883 585
R428 B.n468 B.n467 585
R429 B.n469 B.n468 585
R430 B.n876 B.n875 585
R431 B.n877 B.n876 585
R432 B.n874 B.n474 585
R433 B.n474 B.n473 585
R434 B.n873 B.n872 585
R435 B.n872 B.n871 585
R436 B.n476 B.n475 585
R437 B.n477 B.n476 585
R438 B.n864 B.n863 585
R439 B.n865 B.n864 585
R440 B.n862 B.n482 585
R441 B.n482 B.n481 585
R442 B.n861 B.n860 585
R443 B.n860 B.n859 585
R444 B.n484 B.n483 585
R445 B.n485 B.n484 585
R446 B.n852 B.n851 585
R447 B.n853 B.n852 585
R448 B.n850 B.n490 585
R449 B.n490 B.n489 585
R450 B.n849 B.n848 585
R451 B.n848 B.n847 585
R452 B.n492 B.n491 585
R453 B.n840 B.n492 585
R454 B.n839 B.n838 585
R455 B.n841 B.n839 585
R456 B.n837 B.n497 585
R457 B.n497 B.n496 585
R458 B.n836 B.n835 585
R459 B.n835 B.n834 585
R460 B.n499 B.n498 585
R461 B.n500 B.n499 585
R462 B.n827 B.n826 585
R463 B.n828 B.n827 585
R464 B.n825 B.n505 585
R465 B.n505 B.n504 585
R466 B.n824 B.n823 585
R467 B.n823 B.n822 585
R468 B.n507 B.n506 585
R469 B.n508 B.n507 585
R470 B.n815 B.n814 585
R471 B.n816 B.n815 585
R472 B.n511 B.n510 585
R473 B.n576 B.n575 585
R474 B.n577 B.n573 585
R475 B.n573 B.n512 585
R476 B.n579 B.n578 585
R477 B.n581 B.n572 585
R478 B.n584 B.n583 585
R479 B.n585 B.n571 585
R480 B.n587 B.n586 585
R481 B.n589 B.n570 585
R482 B.n592 B.n591 585
R483 B.n593 B.n569 585
R484 B.n595 B.n594 585
R485 B.n597 B.n568 585
R486 B.n600 B.n599 585
R487 B.n601 B.n567 585
R488 B.n603 B.n602 585
R489 B.n605 B.n566 585
R490 B.n608 B.n607 585
R491 B.n609 B.n565 585
R492 B.n611 B.n610 585
R493 B.n613 B.n564 585
R494 B.n616 B.n615 585
R495 B.n617 B.n563 585
R496 B.n619 B.n618 585
R497 B.n621 B.n562 585
R498 B.n624 B.n623 585
R499 B.n625 B.n561 585
R500 B.n627 B.n626 585
R501 B.n629 B.n560 585
R502 B.n632 B.n631 585
R503 B.n633 B.n559 585
R504 B.n635 B.n634 585
R505 B.n637 B.n558 585
R506 B.n640 B.n639 585
R507 B.n641 B.n557 585
R508 B.n643 B.n642 585
R509 B.n645 B.n556 585
R510 B.n648 B.n647 585
R511 B.n649 B.n555 585
R512 B.n651 B.n650 585
R513 B.n653 B.n554 585
R514 B.n656 B.n655 585
R515 B.n657 B.n553 585
R516 B.n659 B.n658 585
R517 B.n661 B.n552 585
R518 B.n664 B.n663 585
R519 B.n665 B.n551 585
R520 B.n667 B.n666 585
R521 B.n669 B.n550 585
R522 B.n672 B.n671 585
R523 B.n673 B.n549 585
R524 B.n675 B.n674 585
R525 B.n677 B.n548 585
R526 B.n680 B.n679 585
R527 B.n681 B.n545 585
R528 B.n684 B.n683 585
R529 B.n686 B.n544 585
R530 B.n689 B.n688 585
R531 B.n690 B.n543 585
R532 B.n692 B.n691 585
R533 B.n694 B.n542 585
R534 B.n697 B.n696 585
R535 B.n698 B.n541 585
R536 B.n703 B.n702 585
R537 B.n705 B.n540 585
R538 B.n708 B.n707 585
R539 B.n709 B.n539 585
R540 B.n711 B.n710 585
R541 B.n713 B.n538 585
R542 B.n716 B.n715 585
R543 B.n717 B.n537 585
R544 B.n719 B.n718 585
R545 B.n721 B.n536 585
R546 B.n724 B.n723 585
R547 B.n725 B.n535 585
R548 B.n727 B.n726 585
R549 B.n729 B.n534 585
R550 B.n732 B.n731 585
R551 B.n733 B.n533 585
R552 B.n735 B.n734 585
R553 B.n737 B.n532 585
R554 B.n740 B.n739 585
R555 B.n741 B.n531 585
R556 B.n743 B.n742 585
R557 B.n745 B.n530 585
R558 B.n748 B.n747 585
R559 B.n749 B.n529 585
R560 B.n751 B.n750 585
R561 B.n753 B.n528 585
R562 B.n756 B.n755 585
R563 B.n757 B.n527 585
R564 B.n759 B.n758 585
R565 B.n761 B.n526 585
R566 B.n764 B.n763 585
R567 B.n765 B.n525 585
R568 B.n767 B.n766 585
R569 B.n769 B.n524 585
R570 B.n772 B.n771 585
R571 B.n773 B.n523 585
R572 B.n775 B.n774 585
R573 B.n777 B.n522 585
R574 B.n780 B.n779 585
R575 B.n781 B.n521 585
R576 B.n783 B.n782 585
R577 B.n785 B.n520 585
R578 B.n788 B.n787 585
R579 B.n789 B.n519 585
R580 B.n791 B.n790 585
R581 B.n793 B.n518 585
R582 B.n796 B.n795 585
R583 B.n797 B.n517 585
R584 B.n799 B.n798 585
R585 B.n801 B.n516 585
R586 B.n804 B.n803 585
R587 B.n805 B.n515 585
R588 B.n807 B.n806 585
R589 B.n809 B.n514 585
R590 B.n812 B.n811 585
R591 B.n813 B.n513 585
R592 B.n818 B.n817 585
R593 B.n817 B.n816 585
R594 B.n819 B.n509 585
R595 B.n509 B.n508 585
R596 B.n821 B.n820 585
R597 B.n822 B.n821 585
R598 B.n503 B.n502 585
R599 B.n504 B.n503 585
R600 B.n830 B.n829 585
R601 B.n829 B.n828 585
R602 B.n831 B.n501 585
R603 B.n501 B.n500 585
R604 B.n833 B.n832 585
R605 B.n834 B.n833 585
R606 B.n495 B.n494 585
R607 B.n496 B.n495 585
R608 B.n843 B.n842 585
R609 B.n842 B.n841 585
R610 B.n844 B.n493 585
R611 B.n840 B.n493 585
R612 B.n846 B.n845 585
R613 B.n847 B.n846 585
R614 B.n488 B.n487 585
R615 B.n489 B.n488 585
R616 B.n855 B.n854 585
R617 B.n854 B.n853 585
R618 B.n856 B.n486 585
R619 B.n486 B.n485 585
R620 B.n858 B.n857 585
R621 B.n859 B.n858 585
R622 B.n480 B.n479 585
R623 B.n481 B.n480 585
R624 B.n867 B.n866 585
R625 B.n866 B.n865 585
R626 B.n868 B.n478 585
R627 B.n478 B.n477 585
R628 B.n870 B.n869 585
R629 B.n871 B.n870 585
R630 B.n472 B.n471 585
R631 B.n473 B.n472 585
R632 B.n879 B.n878 585
R633 B.n878 B.n877 585
R634 B.n880 B.n470 585
R635 B.n470 B.n469 585
R636 B.n882 B.n881 585
R637 B.n883 B.n882 585
R638 B.n464 B.n463 585
R639 B.n465 B.n464 585
R640 B.n891 B.n890 585
R641 B.n890 B.n889 585
R642 B.n892 B.n462 585
R643 B.n462 B.n461 585
R644 B.n894 B.n893 585
R645 B.n895 B.n894 585
R646 B.n456 B.n455 585
R647 B.n457 B.n456 585
R648 B.n903 B.n902 585
R649 B.n902 B.n901 585
R650 B.n904 B.n454 585
R651 B.n454 B.n453 585
R652 B.n906 B.n905 585
R653 B.n907 B.n906 585
R654 B.n448 B.n447 585
R655 B.n449 B.n448 585
R656 B.n915 B.n914 585
R657 B.n914 B.n913 585
R658 B.n916 B.n446 585
R659 B.n446 B.n445 585
R660 B.n918 B.n917 585
R661 B.n919 B.n918 585
R662 B.n440 B.n439 585
R663 B.n441 B.n440 585
R664 B.n927 B.n926 585
R665 B.n926 B.n925 585
R666 B.n928 B.n438 585
R667 B.n438 B.n437 585
R668 B.n930 B.n929 585
R669 B.n931 B.n930 585
R670 B.n432 B.n431 585
R671 B.n433 B.n432 585
R672 B.n939 B.n938 585
R673 B.n938 B.n937 585
R674 B.n940 B.n430 585
R675 B.n430 B.n429 585
R676 B.n942 B.n941 585
R677 B.n943 B.n942 585
R678 B.n424 B.n423 585
R679 B.n425 B.n424 585
R680 B.n951 B.n950 585
R681 B.n950 B.n949 585
R682 B.n952 B.n422 585
R683 B.n422 B.n421 585
R684 B.n954 B.n953 585
R685 B.n955 B.n954 585
R686 B.n416 B.n415 585
R687 B.n417 B.n416 585
R688 B.n963 B.n962 585
R689 B.n962 B.n961 585
R690 B.n964 B.n414 585
R691 B.n414 B.n413 585
R692 B.n966 B.n965 585
R693 B.n967 B.n966 585
R694 B.n408 B.n407 585
R695 B.n409 B.n408 585
R696 B.n976 B.n975 585
R697 B.n975 B.n974 585
R698 B.n977 B.n406 585
R699 B.n406 B.n405 585
R700 B.n979 B.n978 585
R701 B.n980 B.n979 585
R702 B.n2 B.n0 585
R703 B.n4 B.n2 585
R704 B.n3 B.n1 585
R705 B.n1169 B.n3 585
R706 B.n1167 B.n1166 585
R707 B.n1168 B.n1167 585
R708 B.n1165 B.n9 585
R709 B.n9 B.n8 585
R710 B.n1164 B.n1163 585
R711 B.n1163 B.n1162 585
R712 B.n11 B.n10 585
R713 B.n1161 B.n11 585
R714 B.n1159 B.n1158 585
R715 B.n1160 B.n1159 585
R716 B.n1157 B.n16 585
R717 B.n16 B.n15 585
R718 B.n1156 B.n1155 585
R719 B.n1155 B.n1154 585
R720 B.n18 B.n17 585
R721 B.n1153 B.n18 585
R722 B.n1151 B.n1150 585
R723 B.n1152 B.n1151 585
R724 B.n1149 B.n23 585
R725 B.n23 B.n22 585
R726 B.n1148 B.n1147 585
R727 B.n1147 B.n1146 585
R728 B.n25 B.n24 585
R729 B.n1145 B.n25 585
R730 B.n1143 B.n1142 585
R731 B.n1144 B.n1143 585
R732 B.n1141 B.n30 585
R733 B.n30 B.n29 585
R734 B.n1140 B.n1139 585
R735 B.n1139 B.n1138 585
R736 B.n32 B.n31 585
R737 B.n1137 B.n32 585
R738 B.n1135 B.n1134 585
R739 B.n1136 B.n1135 585
R740 B.n1133 B.n37 585
R741 B.n37 B.n36 585
R742 B.n1132 B.n1131 585
R743 B.n1131 B.n1130 585
R744 B.n39 B.n38 585
R745 B.n1129 B.n39 585
R746 B.n1127 B.n1126 585
R747 B.n1128 B.n1127 585
R748 B.n1125 B.n44 585
R749 B.n44 B.n43 585
R750 B.n1124 B.n1123 585
R751 B.n1123 B.n1122 585
R752 B.n46 B.n45 585
R753 B.n1121 B.n46 585
R754 B.n1119 B.n1118 585
R755 B.n1120 B.n1119 585
R756 B.n1117 B.n51 585
R757 B.n51 B.n50 585
R758 B.n1116 B.n1115 585
R759 B.n1115 B.n1114 585
R760 B.n53 B.n52 585
R761 B.n1113 B.n53 585
R762 B.n1111 B.n1110 585
R763 B.n1112 B.n1111 585
R764 B.n1109 B.n58 585
R765 B.n58 B.n57 585
R766 B.n1108 B.n1107 585
R767 B.n1107 B.n1106 585
R768 B.n60 B.n59 585
R769 B.n1105 B.n60 585
R770 B.n1103 B.n1102 585
R771 B.n1104 B.n1103 585
R772 B.n1101 B.n65 585
R773 B.n65 B.n64 585
R774 B.n1100 B.n1099 585
R775 B.n1099 B.n1098 585
R776 B.n67 B.n66 585
R777 B.n1097 B.n67 585
R778 B.n1095 B.n1094 585
R779 B.n1096 B.n1095 585
R780 B.n1093 B.n72 585
R781 B.n72 B.n71 585
R782 B.n1092 B.n1091 585
R783 B.n1091 B.n1090 585
R784 B.n74 B.n73 585
R785 B.n1089 B.n74 585
R786 B.n1087 B.n1086 585
R787 B.n1088 B.n1087 585
R788 B.n1085 B.n79 585
R789 B.n79 B.n78 585
R790 B.n1084 B.n1083 585
R791 B.n1083 B.n1082 585
R792 B.n81 B.n80 585
R793 B.n1081 B.n81 585
R794 B.n1079 B.n1078 585
R795 B.n1080 B.n1079 585
R796 B.n1077 B.n85 585
R797 B.n88 B.n85 585
R798 B.n1076 B.n1075 585
R799 B.n1075 B.n1074 585
R800 B.n87 B.n86 585
R801 B.n1073 B.n87 585
R802 B.n1071 B.n1070 585
R803 B.n1072 B.n1071 585
R804 B.n1069 B.n93 585
R805 B.n93 B.n92 585
R806 B.n1068 B.n1067 585
R807 B.n1067 B.n1066 585
R808 B.n95 B.n94 585
R809 B.n1065 B.n95 585
R810 B.n1063 B.n1062 585
R811 B.n1064 B.n1063 585
R812 B.n1061 B.n100 585
R813 B.n100 B.n99 585
R814 B.n1060 B.n1059 585
R815 B.n1059 B.n1058 585
R816 B.n1172 B.n1171 585
R817 B.n1171 B.n1170 585
R818 B.n817 B.n511 516.524
R819 B.n1059 B.n102 516.524
R820 B.n815 B.n513 516.524
R821 B.n1056 B.n103 516.524
R822 B.n699 B.t13 316.091
R823 B.n546 B.t17 316.091
R824 B.n167 B.t6 316.091
R825 B.n164 B.t10 316.091
R826 B.n1057 B.n162 256.663
R827 B.n1057 B.n161 256.663
R828 B.n1057 B.n160 256.663
R829 B.n1057 B.n159 256.663
R830 B.n1057 B.n158 256.663
R831 B.n1057 B.n157 256.663
R832 B.n1057 B.n156 256.663
R833 B.n1057 B.n155 256.663
R834 B.n1057 B.n154 256.663
R835 B.n1057 B.n153 256.663
R836 B.n1057 B.n152 256.663
R837 B.n1057 B.n151 256.663
R838 B.n1057 B.n150 256.663
R839 B.n1057 B.n149 256.663
R840 B.n1057 B.n148 256.663
R841 B.n1057 B.n147 256.663
R842 B.n1057 B.n146 256.663
R843 B.n1057 B.n145 256.663
R844 B.n1057 B.n144 256.663
R845 B.n1057 B.n143 256.663
R846 B.n1057 B.n142 256.663
R847 B.n1057 B.n141 256.663
R848 B.n1057 B.n140 256.663
R849 B.n1057 B.n139 256.663
R850 B.n1057 B.n138 256.663
R851 B.n1057 B.n137 256.663
R852 B.n1057 B.n136 256.663
R853 B.n1057 B.n135 256.663
R854 B.n1057 B.n134 256.663
R855 B.n1057 B.n133 256.663
R856 B.n1057 B.n132 256.663
R857 B.n1057 B.n131 256.663
R858 B.n1057 B.n130 256.663
R859 B.n1057 B.n129 256.663
R860 B.n1057 B.n128 256.663
R861 B.n1057 B.n127 256.663
R862 B.n1057 B.n126 256.663
R863 B.n1057 B.n125 256.663
R864 B.n1057 B.n124 256.663
R865 B.n1057 B.n123 256.663
R866 B.n1057 B.n122 256.663
R867 B.n1057 B.n121 256.663
R868 B.n1057 B.n120 256.663
R869 B.n1057 B.n119 256.663
R870 B.n1057 B.n118 256.663
R871 B.n1057 B.n117 256.663
R872 B.n1057 B.n116 256.663
R873 B.n1057 B.n115 256.663
R874 B.n1057 B.n114 256.663
R875 B.n1057 B.n113 256.663
R876 B.n1057 B.n112 256.663
R877 B.n1057 B.n111 256.663
R878 B.n1057 B.n110 256.663
R879 B.n1057 B.n109 256.663
R880 B.n1057 B.n108 256.663
R881 B.n1057 B.n107 256.663
R882 B.n1057 B.n106 256.663
R883 B.n1057 B.n105 256.663
R884 B.n1057 B.n104 256.663
R885 B.n574 B.n512 256.663
R886 B.n580 B.n512 256.663
R887 B.n582 B.n512 256.663
R888 B.n588 B.n512 256.663
R889 B.n590 B.n512 256.663
R890 B.n596 B.n512 256.663
R891 B.n598 B.n512 256.663
R892 B.n604 B.n512 256.663
R893 B.n606 B.n512 256.663
R894 B.n612 B.n512 256.663
R895 B.n614 B.n512 256.663
R896 B.n620 B.n512 256.663
R897 B.n622 B.n512 256.663
R898 B.n628 B.n512 256.663
R899 B.n630 B.n512 256.663
R900 B.n636 B.n512 256.663
R901 B.n638 B.n512 256.663
R902 B.n644 B.n512 256.663
R903 B.n646 B.n512 256.663
R904 B.n652 B.n512 256.663
R905 B.n654 B.n512 256.663
R906 B.n660 B.n512 256.663
R907 B.n662 B.n512 256.663
R908 B.n668 B.n512 256.663
R909 B.n670 B.n512 256.663
R910 B.n676 B.n512 256.663
R911 B.n678 B.n512 256.663
R912 B.n685 B.n512 256.663
R913 B.n687 B.n512 256.663
R914 B.n693 B.n512 256.663
R915 B.n695 B.n512 256.663
R916 B.n704 B.n512 256.663
R917 B.n706 B.n512 256.663
R918 B.n712 B.n512 256.663
R919 B.n714 B.n512 256.663
R920 B.n720 B.n512 256.663
R921 B.n722 B.n512 256.663
R922 B.n728 B.n512 256.663
R923 B.n730 B.n512 256.663
R924 B.n736 B.n512 256.663
R925 B.n738 B.n512 256.663
R926 B.n744 B.n512 256.663
R927 B.n746 B.n512 256.663
R928 B.n752 B.n512 256.663
R929 B.n754 B.n512 256.663
R930 B.n760 B.n512 256.663
R931 B.n762 B.n512 256.663
R932 B.n768 B.n512 256.663
R933 B.n770 B.n512 256.663
R934 B.n776 B.n512 256.663
R935 B.n778 B.n512 256.663
R936 B.n784 B.n512 256.663
R937 B.n786 B.n512 256.663
R938 B.n792 B.n512 256.663
R939 B.n794 B.n512 256.663
R940 B.n800 B.n512 256.663
R941 B.n802 B.n512 256.663
R942 B.n808 B.n512 256.663
R943 B.n810 B.n512 256.663
R944 B.n817 B.n509 163.367
R945 B.n821 B.n509 163.367
R946 B.n821 B.n503 163.367
R947 B.n829 B.n503 163.367
R948 B.n829 B.n501 163.367
R949 B.n833 B.n501 163.367
R950 B.n833 B.n495 163.367
R951 B.n842 B.n495 163.367
R952 B.n842 B.n493 163.367
R953 B.n846 B.n493 163.367
R954 B.n846 B.n488 163.367
R955 B.n854 B.n488 163.367
R956 B.n854 B.n486 163.367
R957 B.n858 B.n486 163.367
R958 B.n858 B.n480 163.367
R959 B.n866 B.n480 163.367
R960 B.n866 B.n478 163.367
R961 B.n870 B.n478 163.367
R962 B.n870 B.n472 163.367
R963 B.n878 B.n472 163.367
R964 B.n878 B.n470 163.367
R965 B.n882 B.n470 163.367
R966 B.n882 B.n464 163.367
R967 B.n890 B.n464 163.367
R968 B.n890 B.n462 163.367
R969 B.n894 B.n462 163.367
R970 B.n894 B.n456 163.367
R971 B.n902 B.n456 163.367
R972 B.n902 B.n454 163.367
R973 B.n906 B.n454 163.367
R974 B.n906 B.n448 163.367
R975 B.n914 B.n448 163.367
R976 B.n914 B.n446 163.367
R977 B.n918 B.n446 163.367
R978 B.n918 B.n440 163.367
R979 B.n926 B.n440 163.367
R980 B.n926 B.n438 163.367
R981 B.n930 B.n438 163.367
R982 B.n930 B.n432 163.367
R983 B.n938 B.n432 163.367
R984 B.n938 B.n430 163.367
R985 B.n942 B.n430 163.367
R986 B.n942 B.n424 163.367
R987 B.n950 B.n424 163.367
R988 B.n950 B.n422 163.367
R989 B.n954 B.n422 163.367
R990 B.n954 B.n416 163.367
R991 B.n962 B.n416 163.367
R992 B.n962 B.n414 163.367
R993 B.n966 B.n414 163.367
R994 B.n966 B.n408 163.367
R995 B.n975 B.n408 163.367
R996 B.n975 B.n406 163.367
R997 B.n979 B.n406 163.367
R998 B.n979 B.n2 163.367
R999 B.n1171 B.n2 163.367
R1000 B.n1171 B.n3 163.367
R1001 B.n1167 B.n3 163.367
R1002 B.n1167 B.n9 163.367
R1003 B.n1163 B.n9 163.367
R1004 B.n1163 B.n11 163.367
R1005 B.n1159 B.n11 163.367
R1006 B.n1159 B.n16 163.367
R1007 B.n1155 B.n16 163.367
R1008 B.n1155 B.n18 163.367
R1009 B.n1151 B.n18 163.367
R1010 B.n1151 B.n23 163.367
R1011 B.n1147 B.n23 163.367
R1012 B.n1147 B.n25 163.367
R1013 B.n1143 B.n25 163.367
R1014 B.n1143 B.n30 163.367
R1015 B.n1139 B.n30 163.367
R1016 B.n1139 B.n32 163.367
R1017 B.n1135 B.n32 163.367
R1018 B.n1135 B.n37 163.367
R1019 B.n1131 B.n37 163.367
R1020 B.n1131 B.n39 163.367
R1021 B.n1127 B.n39 163.367
R1022 B.n1127 B.n44 163.367
R1023 B.n1123 B.n44 163.367
R1024 B.n1123 B.n46 163.367
R1025 B.n1119 B.n46 163.367
R1026 B.n1119 B.n51 163.367
R1027 B.n1115 B.n51 163.367
R1028 B.n1115 B.n53 163.367
R1029 B.n1111 B.n53 163.367
R1030 B.n1111 B.n58 163.367
R1031 B.n1107 B.n58 163.367
R1032 B.n1107 B.n60 163.367
R1033 B.n1103 B.n60 163.367
R1034 B.n1103 B.n65 163.367
R1035 B.n1099 B.n65 163.367
R1036 B.n1099 B.n67 163.367
R1037 B.n1095 B.n67 163.367
R1038 B.n1095 B.n72 163.367
R1039 B.n1091 B.n72 163.367
R1040 B.n1091 B.n74 163.367
R1041 B.n1087 B.n74 163.367
R1042 B.n1087 B.n79 163.367
R1043 B.n1083 B.n79 163.367
R1044 B.n1083 B.n81 163.367
R1045 B.n1079 B.n81 163.367
R1046 B.n1079 B.n85 163.367
R1047 B.n1075 B.n85 163.367
R1048 B.n1075 B.n87 163.367
R1049 B.n1071 B.n87 163.367
R1050 B.n1071 B.n93 163.367
R1051 B.n1067 B.n93 163.367
R1052 B.n1067 B.n95 163.367
R1053 B.n1063 B.n95 163.367
R1054 B.n1063 B.n100 163.367
R1055 B.n1059 B.n100 163.367
R1056 B.n575 B.n573 163.367
R1057 B.n579 B.n573 163.367
R1058 B.n583 B.n581 163.367
R1059 B.n587 B.n571 163.367
R1060 B.n591 B.n589 163.367
R1061 B.n595 B.n569 163.367
R1062 B.n599 B.n597 163.367
R1063 B.n603 B.n567 163.367
R1064 B.n607 B.n605 163.367
R1065 B.n611 B.n565 163.367
R1066 B.n615 B.n613 163.367
R1067 B.n619 B.n563 163.367
R1068 B.n623 B.n621 163.367
R1069 B.n627 B.n561 163.367
R1070 B.n631 B.n629 163.367
R1071 B.n635 B.n559 163.367
R1072 B.n639 B.n637 163.367
R1073 B.n643 B.n557 163.367
R1074 B.n647 B.n645 163.367
R1075 B.n651 B.n555 163.367
R1076 B.n655 B.n653 163.367
R1077 B.n659 B.n553 163.367
R1078 B.n663 B.n661 163.367
R1079 B.n667 B.n551 163.367
R1080 B.n671 B.n669 163.367
R1081 B.n675 B.n549 163.367
R1082 B.n679 B.n677 163.367
R1083 B.n684 B.n545 163.367
R1084 B.n688 B.n686 163.367
R1085 B.n692 B.n543 163.367
R1086 B.n696 B.n694 163.367
R1087 B.n703 B.n541 163.367
R1088 B.n707 B.n705 163.367
R1089 B.n711 B.n539 163.367
R1090 B.n715 B.n713 163.367
R1091 B.n719 B.n537 163.367
R1092 B.n723 B.n721 163.367
R1093 B.n727 B.n535 163.367
R1094 B.n731 B.n729 163.367
R1095 B.n735 B.n533 163.367
R1096 B.n739 B.n737 163.367
R1097 B.n743 B.n531 163.367
R1098 B.n747 B.n745 163.367
R1099 B.n751 B.n529 163.367
R1100 B.n755 B.n753 163.367
R1101 B.n759 B.n527 163.367
R1102 B.n763 B.n761 163.367
R1103 B.n767 B.n525 163.367
R1104 B.n771 B.n769 163.367
R1105 B.n775 B.n523 163.367
R1106 B.n779 B.n777 163.367
R1107 B.n783 B.n521 163.367
R1108 B.n787 B.n785 163.367
R1109 B.n791 B.n519 163.367
R1110 B.n795 B.n793 163.367
R1111 B.n799 B.n517 163.367
R1112 B.n803 B.n801 163.367
R1113 B.n807 B.n515 163.367
R1114 B.n811 B.n809 163.367
R1115 B.n815 B.n507 163.367
R1116 B.n823 B.n507 163.367
R1117 B.n823 B.n505 163.367
R1118 B.n827 B.n505 163.367
R1119 B.n827 B.n499 163.367
R1120 B.n835 B.n499 163.367
R1121 B.n835 B.n497 163.367
R1122 B.n839 B.n497 163.367
R1123 B.n839 B.n492 163.367
R1124 B.n848 B.n492 163.367
R1125 B.n848 B.n490 163.367
R1126 B.n852 B.n490 163.367
R1127 B.n852 B.n484 163.367
R1128 B.n860 B.n484 163.367
R1129 B.n860 B.n482 163.367
R1130 B.n864 B.n482 163.367
R1131 B.n864 B.n476 163.367
R1132 B.n872 B.n476 163.367
R1133 B.n872 B.n474 163.367
R1134 B.n876 B.n474 163.367
R1135 B.n876 B.n468 163.367
R1136 B.n884 B.n468 163.367
R1137 B.n884 B.n466 163.367
R1138 B.n888 B.n466 163.367
R1139 B.n888 B.n460 163.367
R1140 B.n896 B.n460 163.367
R1141 B.n896 B.n458 163.367
R1142 B.n900 B.n458 163.367
R1143 B.n900 B.n452 163.367
R1144 B.n908 B.n452 163.367
R1145 B.n908 B.n450 163.367
R1146 B.n912 B.n450 163.367
R1147 B.n912 B.n444 163.367
R1148 B.n920 B.n444 163.367
R1149 B.n920 B.n442 163.367
R1150 B.n924 B.n442 163.367
R1151 B.n924 B.n436 163.367
R1152 B.n932 B.n436 163.367
R1153 B.n932 B.n434 163.367
R1154 B.n936 B.n434 163.367
R1155 B.n936 B.n428 163.367
R1156 B.n944 B.n428 163.367
R1157 B.n944 B.n426 163.367
R1158 B.n948 B.n426 163.367
R1159 B.n948 B.n420 163.367
R1160 B.n956 B.n420 163.367
R1161 B.n956 B.n418 163.367
R1162 B.n960 B.n418 163.367
R1163 B.n960 B.n412 163.367
R1164 B.n968 B.n412 163.367
R1165 B.n968 B.n410 163.367
R1166 B.n973 B.n410 163.367
R1167 B.n973 B.n404 163.367
R1168 B.n981 B.n404 163.367
R1169 B.n982 B.n981 163.367
R1170 B.n982 B.n5 163.367
R1171 B.n6 B.n5 163.367
R1172 B.n7 B.n6 163.367
R1173 B.n987 B.n7 163.367
R1174 B.n987 B.n12 163.367
R1175 B.n13 B.n12 163.367
R1176 B.n14 B.n13 163.367
R1177 B.n992 B.n14 163.367
R1178 B.n992 B.n19 163.367
R1179 B.n20 B.n19 163.367
R1180 B.n21 B.n20 163.367
R1181 B.n997 B.n21 163.367
R1182 B.n997 B.n26 163.367
R1183 B.n27 B.n26 163.367
R1184 B.n28 B.n27 163.367
R1185 B.n1002 B.n28 163.367
R1186 B.n1002 B.n33 163.367
R1187 B.n34 B.n33 163.367
R1188 B.n35 B.n34 163.367
R1189 B.n1007 B.n35 163.367
R1190 B.n1007 B.n40 163.367
R1191 B.n41 B.n40 163.367
R1192 B.n42 B.n41 163.367
R1193 B.n1012 B.n42 163.367
R1194 B.n1012 B.n47 163.367
R1195 B.n48 B.n47 163.367
R1196 B.n49 B.n48 163.367
R1197 B.n1017 B.n49 163.367
R1198 B.n1017 B.n54 163.367
R1199 B.n55 B.n54 163.367
R1200 B.n56 B.n55 163.367
R1201 B.n1022 B.n56 163.367
R1202 B.n1022 B.n61 163.367
R1203 B.n62 B.n61 163.367
R1204 B.n63 B.n62 163.367
R1205 B.n1027 B.n63 163.367
R1206 B.n1027 B.n68 163.367
R1207 B.n69 B.n68 163.367
R1208 B.n70 B.n69 163.367
R1209 B.n1032 B.n70 163.367
R1210 B.n1032 B.n75 163.367
R1211 B.n76 B.n75 163.367
R1212 B.n77 B.n76 163.367
R1213 B.n1037 B.n77 163.367
R1214 B.n1037 B.n82 163.367
R1215 B.n83 B.n82 163.367
R1216 B.n84 B.n83 163.367
R1217 B.n1042 B.n84 163.367
R1218 B.n1042 B.n89 163.367
R1219 B.n90 B.n89 163.367
R1220 B.n91 B.n90 163.367
R1221 B.n1047 B.n91 163.367
R1222 B.n1047 B.n96 163.367
R1223 B.n97 B.n96 163.367
R1224 B.n98 B.n97 163.367
R1225 B.n1052 B.n98 163.367
R1226 B.n1052 B.n103 163.367
R1227 B.n171 B.n170 163.367
R1228 B.n175 B.n174 163.367
R1229 B.n179 B.n178 163.367
R1230 B.n183 B.n182 163.367
R1231 B.n187 B.n186 163.367
R1232 B.n191 B.n190 163.367
R1233 B.n195 B.n194 163.367
R1234 B.n199 B.n198 163.367
R1235 B.n203 B.n202 163.367
R1236 B.n207 B.n206 163.367
R1237 B.n211 B.n210 163.367
R1238 B.n215 B.n214 163.367
R1239 B.n219 B.n218 163.367
R1240 B.n223 B.n222 163.367
R1241 B.n227 B.n226 163.367
R1242 B.n231 B.n230 163.367
R1243 B.n235 B.n234 163.367
R1244 B.n239 B.n238 163.367
R1245 B.n243 B.n242 163.367
R1246 B.n247 B.n246 163.367
R1247 B.n251 B.n250 163.367
R1248 B.n255 B.n254 163.367
R1249 B.n259 B.n258 163.367
R1250 B.n263 B.n262 163.367
R1251 B.n267 B.n266 163.367
R1252 B.n271 B.n270 163.367
R1253 B.n275 B.n274 163.367
R1254 B.n280 B.n279 163.367
R1255 B.n284 B.n283 163.367
R1256 B.n288 B.n287 163.367
R1257 B.n292 B.n291 163.367
R1258 B.n296 B.n295 163.367
R1259 B.n300 B.n299 163.367
R1260 B.n304 B.n303 163.367
R1261 B.n308 B.n307 163.367
R1262 B.n312 B.n311 163.367
R1263 B.n316 B.n315 163.367
R1264 B.n320 B.n319 163.367
R1265 B.n324 B.n323 163.367
R1266 B.n328 B.n327 163.367
R1267 B.n332 B.n331 163.367
R1268 B.n336 B.n335 163.367
R1269 B.n340 B.n339 163.367
R1270 B.n344 B.n343 163.367
R1271 B.n348 B.n347 163.367
R1272 B.n352 B.n351 163.367
R1273 B.n356 B.n355 163.367
R1274 B.n360 B.n359 163.367
R1275 B.n364 B.n363 163.367
R1276 B.n368 B.n367 163.367
R1277 B.n372 B.n371 163.367
R1278 B.n376 B.n375 163.367
R1279 B.n380 B.n379 163.367
R1280 B.n384 B.n383 163.367
R1281 B.n388 B.n387 163.367
R1282 B.n392 B.n391 163.367
R1283 B.n396 B.n395 163.367
R1284 B.n400 B.n399 163.367
R1285 B.n1056 B.n163 163.367
R1286 B.n699 B.t16 150.156
R1287 B.n164 B.t11 150.156
R1288 B.n546 B.t19 150.135
R1289 B.n167 B.t8 150.135
R1290 B.n700 B.n699 78.7399
R1291 B.n547 B.n546 78.7399
R1292 B.n168 B.n167 78.7399
R1293 B.n165 B.n164 78.7399
R1294 B.n574 B.n511 71.676
R1295 B.n580 B.n579 71.676
R1296 B.n583 B.n582 71.676
R1297 B.n588 B.n587 71.676
R1298 B.n591 B.n590 71.676
R1299 B.n596 B.n595 71.676
R1300 B.n599 B.n598 71.676
R1301 B.n604 B.n603 71.676
R1302 B.n607 B.n606 71.676
R1303 B.n612 B.n611 71.676
R1304 B.n615 B.n614 71.676
R1305 B.n620 B.n619 71.676
R1306 B.n623 B.n622 71.676
R1307 B.n628 B.n627 71.676
R1308 B.n631 B.n630 71.676
R1309 B.n636 B.n635 71.676
R1310 B.n639 B.n638 71.676
R1311 B.n644 B.n643 71.676
R1312 B.n647 B.n646 71.676
R1313 B.n652 B.n651 71.676
R1314 B.n655 B.n654 71.676
R1315 B.n660 B.n659 71.676
R1316 B.n663 B.n662 71.676
R1317 B.n668 B.n667 71.676
R1318 B.n671 B.n670 71.676
R1319 B.n676 B.n675 71.676
R1320 B.n679 B.n678 71.676
R1321 B.n685 B.n684 71.676
R1322 B.n688 B.n687 71.676
R1323 B.n693 B.n692 71.676
R1324 B.n696 B.n695 71.676
R1325 B.n704 B.n703 71.676
R1326 B.n707 B.n706 71.676
R1327 B.n712 B.n711 71.676
R1328 B.n715 B.n714 71.676
R1329 B.n720 B.n719 71.676
R1330 B.n723 B.n722 71.676
R1331 B.n728 B.n727 71.676
R1332 B.n731 B.n730 71.676
R1333 B.n736 B.n735 71.676
R1334 B.n739 B.n738 71.676
R1335 B.n744 B.n743 71.676
R1336 B.n747 B.n746 71.676
R1337 B.n752 B.n751 71.676
R1338 B.n755 B.n754 71.676
R1339 B.n760 B.n759 71.676
R1340 B.n763 B.n762 71.676
R1341 B.n768 B.n767 71.676
R1342 B.n771 B.n770 71.676
R1343 B.n776 B.n775 71.676
R1344 B.n779 B.n778 71.676
R1345 B.n784 B.n783 71.676
R1346 B.n787 B.n786 71.676
R1347 B.n792 B.n791 71.676
R1348 B.n795 B.n794 71.676
R1349 B.n800 B.n799 71.676
R1350 B.n803 B.n802 71.676
R1351 B.n808 B.n807 71.676
R1352 B.n811 B.n810 71.676
R1353 B.n104 B.n102 71.676
R1354 B.n171 B.n105 71.676
R1355 B.n175 B.n106 71.676
R1356 B.n179 B.n107 71.676
R1357 B.n183 B.n108 71.676
R1358 B.n187 B.n109 71.676
R1359 B.n191 B.n110 71.676
R1360 B.n195 B.n111 71.676
R1361 B.n199 B.n112 71.676
R1362 B.n203 B.n113 71.676
R1363 B.n207 B.n114 71.676
R1364 B.n211 B.n115 71.676
R1365 B.n215 B.n116 71.676
R1366 B.n219 B.n117 71.676
R1367 B.n223 B.n118 71.676
R1368 B.n227 B.n119 71.676
R1369 B.n231 B.n120 71.676
R1370 B.n235 B.n121 71.676
R1371 B.n239 B.n122 71.676
R1372 B.n243 B.n123 71.676
R1373 B.n247 B.n124 71.676
R1374 B.n251 B.n125 71.676
R1375 B.n255 B.n126 71.676
R1376 B.n259 B.n127 71.676
R1377 B.n263 B.n128 71.676
R1378 B.n267 B.n129 71.676
R1379 B.n271 B.n130 71.676
R1380 B.n275 B.n131 71.676
R1381 B.n280 B.n132 71.676
R1382 B.n284 B.n133 71.676
R1383 B.n288 B.n134 71.676
R1384 B.n292 B.n135 71.676
R1385 B.n296 B.n136 71.676
R1386 B.n300 B.n137 71.676
R1387 B.n304 B.n138 71.676
R1388 B.n308 B.n139 71.676
R1389 B.n312 B.n140 71.676
R1390 B.n316 B.n141 71.676
R1391 B.n320 B.n142 71.676
R1392 B.n324 B.n143 71.676
R1393 B.n328 B.n144 71.676
R1394 B.n332 B.n145 71.676
R1395 B.n336 B.n146 71.676
R1396 B.n340 B.n147 71.676
R1397 B.n344 B.n148 71.676
R1398 B.n348 B.n149 71.676
R1399 B.n352 B.n150 71.676
R1400 B.n356 B.n151 71.676
R1401 B.n360 B.n152 71.676
R1402 B.n364 B.n153 71.676
R1403 B.n368 B.n154 71.676
R1404 B.n372 B.n155 71.676
R1405 B.n376 B.n156 71.676
R1406 B.n380 B.n157 71.676
R1407 B.n384 B.n158 71.676
R1408 B.n388 B.n159 71.676
R1409 B.n392 B.n160 71.676
R1410 B.n396 B.n161 71.676
R1411 B.n400 B.n162 71.676
R1412 B.n163 B.n162 71.676
R1413 B.n399 B.n161 71.676
R1414 B.n395 B.n160 71.676
R1415 B.n391 B.n159 71.676
R1416 B.n387 B.n158 71.676
R1417 B.n383 B.n157 71.676
R1418 B.n379 B.n156 71.676
R1419 B.n375 B.n155 71.676
R1420 B.n371 B.n154 71.676
R1421 B.n367 B.n153 71.676
R1422 B.n363 B.n152 71.676
R1423 B.n359 B.n151 71.676
R1424 B.n355 B.n150 71.676
R1425 B.n351 B.n149 71.676
R1426 B.n347 B.n148 71.676
R1427 B.n343 B.n147 71.676
R1428 B.n339 B.n146 71.676
R1429 B.n335 B.n145 71.676
R1430 B.n331 B.n144 71.676
R1431 B.n327 B.n143 71.676
R1432 B.n323 B.n142 71.676
R1433 B.n319 B.n141 71.676
R1434 B.n315 B.n140 71.676
R1435 B.n311 B.n139 71.676
R1436 B.n307 B.n138 71.676
R1437 B.n303 B.n137 71.676
R1438 B.n299 B.n136 71.676
R1439 B.n295 B.n135 71.676
R1440 B.n291 B.n134 71.676
R1441 B.n287 B.n133 71.676
R1442 B.n283 B.n132 71.676
R1443 B.n279 B.n131 71.676
R1444 B.n274 B.n130 71.676
R1445 B.n270 B.n129 71.676
R1446 B.n266 B.n128 71.676
R1447 B.n262 B.n127 71.676
R1448 B.n258 B.n126 71.676
R1449 B.n254 B.n125 71.676
R1450 B.n250 B.n124 71.676
R1451 B.n246 B.n123 71.676
R1452 B.n242 B.n122 71.676
R1453 B.n238 B.n121 71.676
R1454 B.n234 B.n120 71.676
R1455 B.n230 B.n119 71.676
R1456 B.n226 B.n118 71.676
R1457 B.n222 B.n117 71.676
R1458 B.n218 B.n116 71.676
R1459 B.n214 B.n115 71.676
R1460 B.n210 B.n114 71.676
R1461 B.n206 B.n113 71.676
R1462 B.n202 B.n112 71.676
R1463 B.n198 B.n111 71.676
R1464 B.n194 B.n110 71.676
R1465 B.n190 B.n109 71.676
R1466 B.n186 B.n108 71.676
R1467 B.n182 B.n107 71.676
R1468 B.n178 B.n106 71.676
R1469 B.n174 B.n105 71.676
R1470 B.n170 B.n104 71.676
R1471 B.n575 B.n574 71.676
R1472 B.n581 B.n580 71.676
R1473 B.n582 B.n571 71.676
R1474 B.n589 B.n588 71.676
R1475 B.n590 B.n569 71.676
R1476 B.n597 B.n596 71.676
R1477 B.n598 B.n567 71.676
R1478 B.n605 B.n604 71.676
R1479 B.n606 B.n565 71.676
R1480 B.n613 B.n612 71.676
R1481 B.n614 B.n563 71.676
R1482 B.n621 B.n620 71.676
R1483 B.n622 B.n561 71.676
R1484 B.n629 B.n628 71.676
R1485 B.n630 B.n559 71.676
R1486 B.n637 B.n636 71.676
R1487 B.n638 B.n557 71.676
R1488 B.n645 B.n644 71.676
R1489 B.n646 B.n555 71.676
R1490 B.n653 B.n652 71.676
R1491 B.n654 B.n553 71.676
R1492 B.n661 B.n660 71.676
R1493 B.n662 B.n551 71.676
R1494 B.n669 B.n668 71.676
R1495 B.n670 B.n549 71.676
R1496 B.n677 B.n676 71.676
R1497 B.n678 B.n545 71.676
R1498 B.n686 B.n685 71.676
R1499 B.n687 B.n543 71.676
R1500 B.n694 B.n693 71.676
R1501 B.n695 B.n541 71.676
R1502 B.n705 B.n704 71.676
R1503 B.n706 B.n539 71.676
R1504 B.n713 B.n712 71.676
R1505 B.n714 B.n537 71.676
R1506 B.n721 B.n720 71.676
R1507 B.n722 B.n535 71.676
R1508 B.n729 B.n728 71.676
R1509 B.n730 B.n533 71.676
R1510 B.n737 B.n736 71.676
R1511 B.n738 B.n531 71.676
R1512 B.n745 B.n744 71.676
R1513 B.n746 B.n529 71.676
R1514 B.n753 B.n752 71.676
R1515 B.n754 B.n527 71.676
R1516 B.n761 B.n760 71.676
R1517 B.n762 B.n525 71.676
R1518 B.n769 B.n768 71.676
R1519 B.n770 B.n523 71.676
R1520 B.n777 B.n776 71.676
R1521 B.n778 B.n521 71.676
R1522 B.n785 B.n784 71.676
R1523 B.n786 B.n519 71.676
R1524 B.n793 B.n792 71.676
R1525 B.n794 B.n517 71.676
R1526 B.n801 B.n800 71.676
R1527 B.n802 B.n515 71.676
R1528 B.n809 B.n808 71.676
R1529 B.n810 B.n513 71.676
R1530 B.n700 B.t15 71.4169
R1531 B.n165 B.t12 71.4169
R1532 B.n547 B.t18 71.3952
R1533 B.n168 B.t9 71.3952
R1534 B.n701 B.n700 59.5399
R1535 B.n682 B.n547 59.5399
R1536 B.n277 B.n168 59.5399
R1537 B.n166 B.n165 59.5399
R1538 B.n816 B.n512 58.0147
R1539 B.n1058 B.n1057 58.0147
R1540 B.n816 B.n508 34.3046
R1541 B.n822 B.n508 34.3046
R1542 B.n822 B.n504 34.3046
R1543 B.n828 B.n504 34.3046
R1544 B.n828 B.n500 34.3046
R1545 B.n834 B.n500 34.3046
R1546 B.n834 B.n496 34.3046
R1547 B.n841 B.n496 34.3046
R1548 B.n841 B.n840 34.3046
R1549 B.n847 B.n489 34.3046
R1550 B.n853 B.n489 34.3046
R1551 B.n853 B.n485 34.3046
R1552 B.n859 B.n485 34.3046
R1553 B.n859 B.n481 34.3046
R1554 B.n865 B.n481 34.3046
R1555 B.n865 B.n477 34.3046
R1556 B.n871 B.n477 34.3046
R1557 B.n871 B.n473 34.3046
R1558 B.n877 B.n473 34.3046
R1559 B.n877 B.n469 34.3046
R1560 B.n883 B.n469 34.3046
R1561 B.n883 B.n465 34.3046
R1562 B.n889 B.n465 34.3046
R1563 B.n895 B.n461 34.3046
R1564 B.n895 B.n457 34.3046
R1565 B.n901 B.n457 34.3046
R1566 B.n901 B.n453 34.3046
R1567 B.n907 B.n453 34.3046
R1568 B.n907 B.n449 34.3046
R1569 B.n913 B.n449 34.3046
R1570 B.n913 B.n445 34.3046
R1571 B.n919 B.n445 34.3046
R1572 B.n919 B.n441 34.3046
R1573 B.n925 B.n441 34.3046
R1574 B.n931 B.n437 34.3046
R1575 B.n931 B.n433 34.3046
R1576 B.n937 B.n433 34.3046
R1577 B.n937 B.n429 34.3046
R1578 B.n943 B.n429 34.3046
R1579 B.n943 B.n425 34.3046
R1580 B.n949 B.n425 34.3046
R1581 B.n949 B.n421 34.3046
R1582 B.n955 B.n421 34.3046
R1583 B.n955 B.n417 34.3046
R1584 B.n961 B.n417 34.3046
R1585 B.n967 B.n413 34.3046
R1586 B.n967 B.n409 34.3046
R1587 B.n974 B.n409 34.3046
R1588 B.n974 B.n405 34.3046
R1589 B.n980 B.n405 34.3046
R1590 B.n980 B.n4 34.3046
R1591 B.n1170 B.n4 34.3046
R1592 B.n1170 B.n1169 34.3046
R1593 B.n1169 B.n1168 34.3046
R1594 B.n1168 B.n8 34.3046
R1595 B.n1162 B.n8 34.3046
R1596 B.n1162 B.n1161 34.3046
R1597 B.n1161 B.n1160 34.3046
R1598 B.n1160 B.n15 34.3046
R1599 B.n1154 B.n1153 34.3046
R1600 B.n1153 B.n1152 34.3046
R1601 B.n1152 B.n22 34.3046
R1602 B.n1146 B.n22 34.3046
R1603 B.n1146 B.n1145 34.3046
R1604 B.n1145 B.n1144 34.3046
R1605 B.n1144 B.n29 34.3046
R1606 B.n1138 B.n29 34.3046
R1607 B.n1138 B.n1137 34.3046
R1608 B.n1137 B.n1136 34.3046
R1609 B.n1136 B.n36 34.3046
R1610 B.n1130 B.n1129 34.3046
R1611 B.n1129 B.n1128 34.3046
R1612 B.n1128 B.n43 34.3046
R1613 B.n1122 B.n43 34.3046
R1614 B.n1122 B.n1121 34.3046
R1615 B.n1121 B.n1120 34.3046
R1616 B.n1120 B.n50 34.3046
R1617 B.n1114 B.n50 34.3046
R1618 B.n1114 B.n1113 34.3046
R1619 B.n1113 B.n1112 34.3046
R1620 B.n1112 B.n57 34.3046
R1621 B.n1106 B.n1105 34.3046
R1622 B.n1105 B.n1104 34.3046
R1623 B.n1104 B.n64 34.3046
R1624 B.n1098 B.n64 34.3046
R1625 B.n1098 B.n1097 34.3046
R1626 B.n1097 B.n1096 34.3046
R1627 B.n1096 B.n71 34.3046
R1628 B.n1090 B.n71 34.3046
R1629 B.n1090 B.n1089 34.3046
R1630 B.n1089 B.n1088 34.3046
R1631 B.n1088 B.n78 34.3046
R1632 B.n1082 B.n78 34.3046
R1633 B.n1082 B.n1081 34.3046
R1634 B.n1081 B.n1080 34.3046
R1635 B.n1074 B.n88 34.3046
R1636 B.n1074 B.n1073 34.3046
R1637 B.n1073 B.n1072 34.3046
R1638 B.n1072 B.n92 34.3046
R1639 B.n1066 B.n92 34.3046
R1640 B.n1066 B.n1065 34.3046
R1641 B.n1065 B.n1064 34.3046
R1642 B.n1064 B.n99 34.3046
R1643 B.n1058 B.n99 34.3046
R1644 B.n1060 B.n101 33.5615
R1645 B.n1055 B.n1054 33.5615
R1646 B.n814 B.n813 33.5615
R1647 B.n818 B.n510 33.5615
R1648 B.n847 B.t14 20.6838
R1649 B.n1080 B.t7 20.6838
R1650 B.t0 B.n413 19.6749
R1651 B.t3 B.n15 19.6749
R1652 B.n889 B.t2 18.6659
R1653 B.n1106 B.t5 18.6659
R1654 B B.n1172 18.0485
R1655 B.t1 B.n437 17.657
R1656 B.t4 B.n36 17.657
R1657 B.n925 B.t1 16.6481
R1658 B.n1130 B.t4 16.6481
R1659 B.t2 B.n461 15.6391
R1660 B.t5 B.n57 15.6391
R1661 B.n961 B.t0 14.6302
R1662 B.n1154 B.t3 14.6302
R1663 B.n840 B.t14 13.6212
R1664 B.n88 B.t7 13.6212
R1665 B.n169 B.n101 10.6151
R1666 B.n172 B.n169 10.6151
R1667 B.n173 B.n172 10.6151
R1668 B.n176 B.n173 10.6151
R1669 B.n177 B.n176 10.6151
R1670 B.n180 B.n177 10.6151
R1671 B.n181 B.n180 10.6151
R1672 B.n184 B.n181 10.6151
R1673 B.n185 B.n184 10.6151
R1674 B.n188 B.n185 10.6151
R1675 B.n189 B.n188 10.6151
R1676 B.n192 B.n189 10.6151
R1677 B.n193 B.n192 10.6151
R1678 B.n196 B.n193 10.6151
R1679 B.n197 B.n196 10.6151
R1680 B.n200 B.n197 10.6151
R1681 B.n201 B.n200 10.6151
R1682 B.n204 B.n201 10.6151
R1683 B.n205 B.n204 10.6151
R1684 B.n208 B.n205 10.6151
R1685 B.n209 B.n208 10.6151
R1686 B.n212 B.n209 10.6151
R1687 B.n213 B.n212 10.6151
R1688 B.n216 B.n213 10.6151
R1689 B.n217 B.n216 10.6151
R1690 B.n220 B.n217 10.6151
R1691 B.n221 B.n220 10.6151
R1692 B.n224 B.n221 10.6151
R1693 B.n225 B.n224 10.6151
R1694 B.n228 B.n225 10.6151
R1695 B.n229 B.n228 10.6151
R1696 B.n232 B.n229 10.6151
R1697 B.n233 B.n232 10.6151
R1698 B.n236 B.n233 10.6151
R1699 B.n237 B.n236 10.6151
R1700 B.n240 B.n237 10.6151
R1701 B.n241 B.n240 10.6151
R1702 B.n244 B.n241 10.6151
R1703 B.n245 B.n244 10.6151
R1704 B.n248 B.n245 10.6151
R1705 B.n249 B.n248 10.6151
R1706 B.n252 B.n249 10.6151
R1707 B.n253 B.n252 10.6151
R1708 B.n256 B.n253 10.6151
R1709 B.n257 B.n256 10.6151
R1710 B.n260 B.n257 10.6151
R1711 B.n261 B.n260 10.6151
R1712 B.n264 B.n261 10.6151
R1713 B.n265 B.n264 10.6151
R1714 B.n268 B.n265 10.6151
R1715 B.n269 B.n268 10.6151
R1716 B.n272 B.n269 10.6151
R1717 B.n273 B.n272 10.6151
R1718 B.n276 B.n273 10.6151
R1719 B.n281 B.n278 10.6151
R1720 B.n282 B.n281 10.6151
R1721 B.n285 B.n282 10.6151
R1722 B.n286 B.n285 10.6151
R1723 B.n289 B.n286 10.6151
R1724 B.n290 B.n289 10.6151
R1725 B.n293 B.n290 10.6151
R1726 B.n294 B.n293 10.6151
R1727 B.n298 B.n297 10.6151
R1728 B.n301 B.n298 10.6151
R1729 B.n302 B.n301 10.6151
R1730 B.n305 B.n302 10.6151
R1731 B.n306 B.n305 10.6151
R1732 B.n309 B.n306 10.6151
R1733 B.n310 B.n309 10.6151
R1734 B.n313 B.n310 10.6151
R1735 B.n314 B.n313 10.6151
R1736 B.n317 B.n314 10.6151
R1737 B.n318 B.n317 10.6151
R1738 B.n321 B.n318 10.6151
R1739 B.n322 B.n321 10.6151
R1740 B.n325 B.n322 10.6151
R1741 B.n326 B.n325 10.6151
R1742 B.n329 B.n326 10.6151
R1743 B.n330 B.n329 10.6151
R1744 B.n333 B.n330 10.6151
R1745 B.n334 B.n333 10.6151
R1746 B.n337 B.n334 10.6151
R1747 B.n338 B.n337 10.6151
R1748 B.n341 B.n338 10.6151
R1749 B.n342 B.n341 10.6151
R1750 B.n345 B.n342 10.6151
R1751 B.n346 B.n345 10.6151
R1752 B.n349 B.n346 10.6151
R1753 B.n350 B.n349 10.6151
R1754 B.n353 B.n350 10.6151
R1755 B.n354 B.n353 10.6151
R1756 B.n357 B.n354 10.6151
R1757 B.n358 B.n357 10.6151
R1758 B.n361 B.n358 10.6151
R1759 B.n362 B.n361 10.6151
R1760 B.n365 B.n362 10.6151
R1761 B.n366 B.n365 10.6151
R1762 B.n369 B.n366 10.6151
R1763 B.n370 B.n369 10.6151
R1764 B.n373 B.n370 10.6151
R1765 B.n374 B.n373 10.6151
R1766 B.n377 B.n374 10.6151
R1767 B.n378 B.n377 10.6151
R1768 B.n381 B.n378 10.6151
R1769 B.n382 B.n381 10.6151
R1770 B.n385 B.n382 10.6151
R1771 B.n386 B.n385 10.6151
R1772 B.n389 B.n386 10.6151
R1773 B.n390 B.n389 10.6151
R1774 B.n393 B.n390 10.6151
R1775 B.n394 B.n393 10.6151
R1776 B.n397 B.n394 10.6151
R1777 B.n398 B.n397 10.6151
R1778 B.n401 B.n398 10.6151
R1779 B.n402 B.n401 10.6151
R1780 B.n1055 B.n402 10.6151
R1781 B.n814 B.n506 10.6151
R1782 B.n824 B.n506 10.6151
R1783 B.n825 B.n824 10.6151
R1784 B.n826 B.n825 10.6151
R1785 B.n826 B.n498 10.6151
R1786 B.n836 B.n498 10.6151
R1787 B.n837 B.n836 10.6151
R1788 B.n838 B.n837 10.6151
R1789 B.n838 B.n491 10.6151
R1790 B.n849 B.n491 10.6151
R1791 B.n850 B.n849 10.6151
R1792 B.n851 B.n850 10.6151
R1793 B.n851 B.n483 10.6151
R1794 B.n861 B.n483 10.6151
R1795 B.n862 B.n861 10.6151
R1796 B.n863 B.n862 10.6151
R1797 B.n863 B.n475 10.6151
R1798 B.n873 B.n475 10.6151
R1799 B.n874 B.n873 10.6151
R1800 B.n875 B.n874 10.6151
R1801 B.n875 B.n467 10.6151
R1802 B.n885 B.n467 10.6151
R1803 B.n886 B.n885 10.6151
R1804 B.n887 B.n886 10.6151
R1805 B.n887 B.n459 10.6151
R1806 B.n897 B.n459 10.6151
R1807 B.n898 B.n897 10.6151
R1808 B.n899 B.n898 10.6151
R1809 B.n899 B.n451 10.6151
R1810 B.n909 B.n451 10.6151
R1811 B.n910 B.n909 10.6151
R1812 B.n911 B.n910 10.6151
R1813 B.n911 B.n443 10.6151
R1814 B.n921 B.n443 10.6151
R1815 B.n922 B.n921 10.6151
R1816 B.n923 B.n922 10.6151
R1817 B.n923 B.n435 10.6151
R1818 B.n933 B.n435 10.6151
R1819 B.n934 B.n933 10.6151
R1820 B.n935 B.n934 10.6151
R1821 B.n935 B.n427 10.6151
R1822 B.n945 B.n427 10.6151
R1823 B.n946 B.n945 10.6151
R1824 B.n947 B.n946 10.6151
R1825 B.n947 B.n419 10.6151
R1826 B.n957 B.n419 10.6151
R1827 B.n958 B.n957 10.6151
R1828 B.n959 B.n958 10.6151
R1829 B.n959 B.n411 10.6151
R1830 B.n969 B.n411 10.6151
R1831 B.n970 B.n969 10.6151
R1832 B.n972 B.n970 10.6151
R1833 B.n972 B.n971 10.6151
R1834 B.n971 B.n403 10.6151
R1835 B.n983 B.n403 10.6151
R1836 B.n984 B.n983 10.6151
R1837 B.n985 B.n984 10.6151
R1838 B.n986 B.n985 10.6151
R1839 B.n988 B.n986 10.6151
R1840 B.n989 B.n988 10.6151
R1841 B.n990 B.n989 10.6151
R1842 B.n991 B.n990 10.6151
R1843 B.n993 B.n991 10.6151
R1844 B.n994 B.n993 10.6151
R1845 B.n995 B.n994 10.6151
R1846 B.n996 B.n995 10.6151
R1847 B.n998 B.n996 10.6151
R1848 B.n999 B.n998 10.6151
R1849 B.n1000 B.n999 10.6151
R1850 B.n1001 B.n1000 10.6151
R1851 B.n1003 B.n1001 10.6151
R1852 B.n1004 B.n1003 10.6151
R1853 B.n1005 B.n1004 10.6151
R1854 B.n1006 B.n1005 10.6151
R1855 B.n1008 B.n1006 10.6151
R1856 B.n1009 B.n1008 10.6151
R1857 B.n1010 B.n1009 10.6151
R1858 B.n1011 B.n1010 10.6151
R1859 B.n1013 B.n1011 10.6151
R1860 B.n1014 B.n1013 10.6151
R1861 B.n1015 B.n1014 10.6151
R1862 B.n1016 B.n1015 10.6151
R1863 B.n1018 B.n1016 10.6151
R1864 B.n1019 B.n1018 10.6151
R1865 B.n1020 B.n1019 10.6151
R1866 B.n1021 B.n1020 10.6151
R1867 B.n1023 B.n1021 10.6151
R1868 B.n1024 B.n1023 10.6151
R1869 B.n1025 B.n1024 10.6151
R1870 B.n1026 B.n1025 10.6151
R1871 B.n1028 B.n1026 10.6151
R1872 B.n1029 B.n1028 10.6151
R1873 B.n1030 B.n1029 10.6151
R1874 B.n1031 B.n1030 10.6151
R1875 B.n1033 B.n1031 10.6151
R1876 B.n1034 B.n1033 10.6151
R1877 B.n1035 B.n1034 10.6151
R1878 B.n1036 B.n1035 10.6151
R1879 B.n1038 B.n1036 10.6151
R1880 B.n1039 B.n1038 10.6151
R1881 B.n1040 B.n1039 10.6151
R1882 B.n1041 B.n1040 10.6151
R1883 B.n1043 B.n1041 10.6151
R1884 B.n1044 B.n1043 10.6151
R1885 B.n1045 B.n1044 10.6151
R1886 B.n1046 B.n1045 10.6151
R1887 B.n1048 B.n1046 10.6151
R1888 B.n1049 B.n1048 10.6151
R1889 B.n1050 B.n1049 10.6151
R1890 B.n1051 B.n1050 10.6151
R1891 B.n1053 B.n1051 10.6151
R1892 B.n1054 B.n1053 10.6151
R1893 B.n576 B.n510 10.6151
R1894 B.n577 B.n576 10.6151
R1895 B.n578 B.n577 10.6151
R1896 B.n578 B.n572 10.6151
R1897 B.n584 B.n572 10.6151
R1898 B.n585 B.n584 10.6151
R1899 B.n586 B.n585 10.6151
R1900 B.n586 B.n570 10.6151
R1901 B.n592 B.n570 10.6151
R1902 B.n593 B.n592 10.6151
R1903 B.n594 B.n593 10.6151
R1904 B.n594 B.n568 10.6151
R1905 B.n600 B.n568 10.6151
R1906 B.n601 B.n600 10.6151
R1907 B.n602 B.n601 10.6151
R1908 B.n602 B.n566 10.6151
R1909 B.n608 B.n566 10.6151
R1910 B.n609 B.n608 10.6151
R1911 B.n610 B.n609 10.6151
R1912 B.n610 B.n564 10.6151
R1913 B.n616 B.n564 10.6151
R1914 B.n617 B.n616 10.6151
R1915 B.n618 B.n617 10.6151
R1916 B.n618 B.n562 10.6151
R1917 B.n624 B.n562 10.6151
R1918 B.n625 B.n624 10.6151
R1919 B.n626 B.n625 10.6151
R1920 B.n626 B.n560 10.6151
R1921 B.n632 B.n560 10.6151
R1922 B.n633 B.n632 10.6151
R1923 B.n634 B.n633 10.6151
R1924 B.n634 B.n558 10.6151
R1925 B.n640 B.n558 10.6151
R1926 B.n641 B.n640 10.6151
R1927 B.n642 B.n641 10.6151
R1928 B.n642 B.n556 10.6151
R1929 B.n648 B.n556 10.6151
R1930 B.n649 B.n648 10.6151
R1931 B.n650 B.n649 10.6151
R1932 B.n650 B.n554 10.6151
R1933 B.n656 B.n554 10.6151
R1934 B.n657 B.n656 10.6151
R1935 B.n658 B.n657 10.6151
R1936 B.n658 B.n552 10.6151
R1937 B.n664 B.n552 10.6151
R1938 B.n665 B.n664 10.6151
R1939 B.n666 B.n665 10.6151
R1940 B.n666 B.n550 10.6151
R1941 B.n672 B.n550 10.6151
R1942 B.n673 B.n672 10.6151
R1943 B.n674 B.n673 10.6151
R1944 B.n674 B.n548 10.6151
R1945 B.n680 B.n548 10.6151
R1946 B.n681 B.n680 10.6151
R1947 B.n683 B.n544 10.6151
R1948 B.n689 B.n544 10.6151
R1949 B.n690 B.n689 10.6151
R1950 B.n691 B.n690 10.6151
R1951 B.n691 B.n542 10.6151
R1952 B.n697 B.n542 10.6151
R1953 B.n698 B.n697 10.6151
R1954 B.n702 B.n698 10.6151
R1955 B.n708 B.n540 10.6151
R1956 B.n709 B.n708 10.6151
R1957 B.n710 B.n709 10.6151
R1958 B.n710 B.n538 10.6151
R1959 B.n716 B.n538 10.6151
R1960 B.n717 B.n716 10.6151
R1961 B.n718 B.n717 10.6151
R1962 B.n718 B.n536 10.6151
R1963 B.n724 B.n536 10.6151
R1964 B.n725 B.n724 10.6151
R1965 B.n726 B.n725 10.6151
R1966 B.n726 B.n534 10.6151
R1967 B.n732 B.n534 10.6151
R1968 B.n733 B.n732 10.6151
R1969 B.n734 B.n733 10.6151
R1970 B.n734 B.n532 10.6151
R1971 B.n740 B.n532 10.6151
R1972 B.n741 B.n740 10.6151
R1973 B.n742 B.n741 10.6151
R1974 B.n742 B.n530 10.6151
R1975 B.n748 B.n530 10.6151
R1976 B.n749 B.n748 10.6151
R1977 B.n750 B.n749 10.6151
R1978 B.n750 B.n528 10.6151
R1979 B.n756 B.n528 10.6151
R1980 B.n757 B.n756 10.6151
R1981 B.n758 B.n757 10.6151
R1982 B.n758 B.n526 10.6151
R1983 B.n764 B.n526 10.6151
R1984 B.n765 B.n764 10.6151
R1985 B.n766 B.n765 10.6151
R1986 B.n766 B.n524 10.6151
R1987 B.n772 B.n524 10.6151
R1988 B.n773 B.n772 10.6151
R1989 B.n774 B.n773 10.6151
R1990 B.n774 B.n522 10.6151
R1991 B.n780 B.n522 10.6151
R1992 B.n781 B.n780 10.6151
R1993 B.n782 B.n781 10.6151
R1994 B.n782 B.n520 10.6151
R1995 B.n788 B.n520 10.6151
R1996 B.n789 B.n788 10.6151
R1997 B.n790 B.n789 10.6151
R1998 B.n790 B.n518 10.6151
R1999 B.n796 B.n518 10.6151
R2000 B.n797 B.n796 10.6151
R2001 B.n798 B.n797 10.6151
R2002 B.n798 B.n516 10.6151
R2003 B.n804 B.n516 10.6151
R2004 B.n805 B.n804 10.6151
R2005 B.n806 B.n805 10.6151
R2006 B.n806 B.n514 10.6151
R2007 B.n812 B.n514 10.6151
R2008 B.n813 B.n812 10.6151
R2009 B.n819 B.n818 10.6151
R2010 B.n820 B.n819 10.6151
R2011 B.n820 B.n502 10.6151
R2012 B.n830 B.n502 10.6151
R2013 B.n831 B.n830 10.6151
R2014 B.n832 B.n831 10.6151
R2015 B.n832 B.n494 10.6151
R2016 B.n843 B.n494 10.6151
R2017 B.n844 B.n843 10.6151
R2018 B.n845 B.n844 10.6151
R2019 B.n845 B.n487 10.6151
R2020 B.n855 B.n487 10.6151
R2021 B.n856 B.n855 10.6151
R2022 B.n857 B.n856 10.6151
R2023 B.n857 B.n479 10.6151
R2024 B.n867 B.n479 10.6151
R2025 B.n868 B.n867 10.6151
R2026 B.n869 B.n868 10.6151
R2027 B.n869 B.n471 10.6151
R2028 B.n879 B.n471 10.6151
R2029 B.n880 B.n879 10.6151
R2030 B.n881 B.n880 10.6151
R2031 B.n881 B.n463 10.6151
R2032 B.n891 B.n463 10.6151
R2033 B.n892 B.n891 10.6151
R2034 B.n893 B.n892 10.6151
R2035 B.n893 B.n455 10.6151
R2036 B.n903 B.n455 10.6151
R2037 B.n904 B.n903 10.6151
R2038 B.n905 B.n904 10.6151
R2039 B.n905 B.n447 10.6151
R2040 B.n915 B.n447 10.6151
R2041 B.n916 B.n915 10.6151
R2042 B.n917 B.n916 10.6151
R2043 B.n917 B.n439 10.6151
R2044 B.n927 B.n439 10.6151
R2045 B.n928 B.n927 10.6151
R2046 B.n929 B.n928 10.6151
R2047 B.n929 B.n431 10.6151
R2048 B.n939 B.n431 10.6151
R2049 B.n940 B.n939 10.6151
R2050 B.n941 B.n940 10.6151
R2051 B.n941 B.n423 10.6151
R2052 B.n951 B.n423 10.6151
R2053 B.n952 B.n951 10.6151
R2054 B.n953 B.n952 10.6151
R2055 B.n953 B.n415 10.6151
R2056 B.n963 B.n415 10.6151
R2057 B.n964 B.n963 10.6151
R2058 B.n965 B.n964 10.6151
R2059 B.n965 B.n407 10.6151
R2060 B.n976 B.n407 10.6151
R2061 B.n977 B.n976 10.6151
R2062 B.n978 B.n977 10.6151
R2063 B.n978 B.n0 10.6151
R2064 B.n1166 B.n1 10.6151
R2065 B.n1166 B.n1165 10.6151
R2066 B.n1165 B.n1164 10.6151
R2067 B.n1164 B.n10 10.6151
R2068 B.n1158 B.n10 10.6151
R2069 B.n1158 B.n1157 10.6151
R2070 B.n1157 B.n1156 10.6151
R2071 B.n1156 B.n17 10.6151
R2072 B.n1150 B.n17 10.6151
R2073 B.n1150 B.n1149 10.6151
R2074 B.n1149 B.n1148 10.6151
R2075 B.n1148 B.n24 10.6151
R2076 B.n1142 B.n24 10.6151
R2077 B.n1142 B.n1141 10.6151
R2078 B.n1141 B.n1140 10.6151
R2079 B.n1140 B.n31 10.6151
R2080 B.n1134 B.n31 10.6151
R2081 B.n1134 B.n1133 10.6151
R2082 B.n1133 B.n1132 10.6151
R2083 B.n1132 B.n38 10.6151
R2084 B.n1126 B.n38 10.6151
R2085 B.n1126 B.n1125 10.6151
R2086 B.n1125 B.n1124 10.6151
R2087 B.n1124 B.n45 10.6151
R2088 B.n1118 B.n45 10.6151
R2089 B.n1118 B.n1117 10.6151
R2090 B.n1117 B.n1116 10.6151
R2091 B.n1116 B.n52 10.6151
R2092 B.n1110 B.n52 10.6151
R2093 B.n1110 B.n1109 10.6151
R2094 B.n1109 B.n1108 10.6151
R2095 B.n1108 B.n59 10.6151
R2096 B.n1102 B.n59 10.6151
R2097 B.n1102 B.n1101 10.6151
R2098 B.n1101 B.n1100 10.6151
R2099 B.n1100 B.n66 10.6151
R2100 B.n1094 B.n66 10.6151
R2101 B.n1094 B.n1093 10.6151
R2102 B.n1093 B.n1092 10.6151
R2103 B.n1092 B.n73 10.6151
R2104 B.n1086 B.n73 10.6151
R2105 B.n1086 B.n1085 10.6151
R2106 B.n1085 B.n1084 10.6151
R2107 B.n1084 B.n80 10.6151
R2108 B.n1078 B.n80 10.6151
R2109 B.n1078 B.n1077 10.6151
R2110 B.n1077 B.n1076 10.6151
R2111 B.n1076 B.n86 10.6151
R2112 B.n1070 B.n86 10.6151
R2113 B.n1070 B.n1069 10.6151
R2114 B.n1069 B.n1068 10.6151
R2115 B.n1068 B.n94 10.6151
R2116 B.n1062 B.n94 10.6151
R2117 B.n1062 B.n1061 10.6151
R2118 B.n1061 B.n1060 10.6151
R2119 B.n278 B.n277 6.5566
R2120 B.n294 B.n166 6.5566
R2121 B.n683 B.n682 6.5566
R2122 B.n702 B.n701 6.5566
R2123 B.n277 B.n276 4.05904
R2124 B.n297 B.n166 4.05904
R2125 B.n682 B.n681 4.05904
R2126 B.n701 B.n540 4.05904
R2127 B.n1172 B.n0 2.81026
R2128 B.n1172 B.n1 2.81026
R2129 VN.n38 VN.n37 161.3
R2130 VN.n36 VN.n21 161.3
R2131 VN.n35 VN.n34 161.3
R2132 VN.n33 VN.n22 161.3
R2133 VN.n32 VN.n31 161.3
R2134 VN.n30 VN.n23 161.3
R2135 VN.n29 VN.n28 161.3
R2136 VN.n27 VN.n24 161.3
R2137 VN.n18 VN.n17 161.3
R2138 VN.n16 VN.n1 161.3
R2139 VN.n15 VN.n14 161.3
R2140 VN.n13 VN.n2 161.3
R2141 VN.n12 VN.n11 161.3
R2142 VN.n10 VN.n3 161.3
R2143 VN.n9 VN.n8 161.3
R2144 VN.n7 VN.n4 161.3
R2145 VN.n26 VN.t4 139.722
R2146 VN.n6 VN.t0 139.722
R2147 VN.n5 VN.t3 106.802
R2148 VN.n0 VN.t5 106.802
R2149 VN.n25 VN.t2 106.802
R2150 VN.n20 VN.t1 106.802
R2151 VN.n19 VN.n0 87.1314
R2152 VN.n39 VN.n20 87.1314
R2153 VN VN.n39 56.7404
R2154 VN.n6 VN.n5 50.484
R2155 VN.n26 VN.n25 50.484
R2156 VN.n11 VN.n2 43.4072
R2157 VN.n31 VN.n22 43.4072
R2158 VN.n11 VN.n10 37.5796
R2159 VN.n31 VN.n30 37.5796
R2160 VN.n5 VN.n4 24.4675
R2161 VN.n9 VN.n4 24.4675
R2162 VN.n10 VN.n9 24.4675
R2163 VN.n15 VN.n2 24.4675
R2164 VN.n16 VN.n15 24.4675
R2165 VN.n17 VN.n16 24.4675
R2166 VN.n30 VN.n29 24.4675
R2167 VN.n29 VN.n24 24.4675
R2168 VN.n25 VN.n24 24.4675
R2169 VN.n37 VN.n36 24.4675
R2170 VN.n36 VN.n35 24.4675
R2171 VN.n35 VN.n22 24.4675
R2172 VN.n17 VN.n0 2.93654
R2173 VN.n37 VN.n20 2.93654
R2174 VN.n27 VN.n26 2.46264
R2175 VN.n7 VN.n6 2.46264
R2176 VN.n39 VN.n38 0.354971
R2177 VN.n19 VN.n18 0.354971
R2178 VN VN.n19 0.26696
R2179 VN.n38 VN.n21 0.189894
R2180 VN.n34 VN.n21 0.189894
R2181 VN.n34 VN.n33 0.189894
R2182 VN.n33 VN.n32 0.189894
R2183 VN.n32 VN.n23 0.189894
R2184 VN.n28 VN.n23 0.189894
R2185 VN.n28 VN.n27 0.189894
R2186 VN.n8 VN.n7 0.189894
R2187 VN.n8 VN.n3 0.189894
R2188 VN.n12 VN.n3 0.189894
R2189 VN.n13 VN.n12 0.189894
R2190 VN.n14 VN.n13 0.189894
R2191 VN.n14 VN.n1 0.189894
R2192 VN.n18 VN.n1 0.189894
R2193 VDD2.n1 VDD2.t5 66.2623
R2194 VDD2.n2 VDD2.t4 63.6929
R2195 VDD2.n1 VDD2.n0 63.3145
R2196 VDD2 VDD2.n3 63.3117
R2197 VDD2.n2 VDD2.n1 49.3403
R2198 VDD2 VDD2.n2 2.68369
R2199 VDD2.n3 VDD2.t3 1.19832
R2200 VDD2.n3 VDD2.t1 1.19832
R2201 VDD2.n0 VDD2.t2 1.19832
R2202 VDD2.n0 VDD2.t0 1.19832
C0 VDD2 VDD1 1.84724f
C1 VTAIL VN 9.88729f
C2 VP VN 8.86583f
C3 VDD1 VTAIL 9.57772f
C4 VDD2 VTAIL 9.636331f
C5 VP VDD1 10.0713f
C6 VDD1 VN 0.152134f
C7 VP VDD2 0.553782f
C8 VDD2 VN 9.67275f
C9 VP VTAIL 9.90205f
C10 VDD2 B 7.641905f
C11 VDD1 B 8.02273f
C12 VTAIL B 10.378037f
C13 VN B 16.56811f
C14 VP B 15.242352f
C15 VDD2.t5 B 3.22296f
C16 VDD2.t2 B 0.276272f
C17 VDD2.t0 B 0.276272f
C18 VDD2.n0 B 2.51582f
C19 VDD2.n1 B 3.10815f
C20 VDD2.t4 B 3.20695f
C21 VDD2.n2 B 2.9172f
C22 VDD2.t3 B 0.276272f
C23 VDD2.t1 B 0.276272f
C24 VDD2.n3 B 2.51579f
C25 VN.t5 B 2.97525f
C26 VN.n0 B 1.09319f
C27 VN.n1 B 0.017573f
C28 VN.n2 B 0.034303f
C29 VN.n3 B 0.017573f
C30 VN.n4 B 0.032752f
C31 VN.t3 B 2.97525f
C32 VN.n5 B 1.10038f
C33 VN.t0 B 3.25025f
C34 VN.n6 B 1.04698f
C35 VN.n7 B 0.224361f
C36 VN.n8 B 0.017573f
C37 VN.n9 B 0.032752f
C38 VN.n10 B 0.035346f
C39 VN.n11 B 0.01441f
C40 VN.n12 B 0.017573f
C41 VN.n13 B 0.017573f
C42 VN.n14 B 0.017573f
C43 VN.n15 B 0.032752f
C44 VN.n16 B 0.032752f
C45 VN.n17 B 0.018522f
C46 VN.n18 B 0.028363f
C47 VN.n19 B 0.053274f
C48 VN.t1 B 2.97525f
C49 VN.n20 B 1.09319f
C50 VN.n21 B 0.017573f
C51 VN.n22 B 0.034303f
C52 VN.n23 B 0.017573f
C53 VN.n24 B 0.032752f
C54 VN.t4 B 3.25025f
C55 VN.t2 B 2.97525f
C56 VN.n25 B 1.10038f
C57 VN.n26 B 1.04698f
C58 VN.n27 B 0.224361f
C59 VN.n28 B 0.017573f
C60 VN.n29 B 0.032752f
C61 VN.n30 B 0.035346f
C62 VN.n31 B 0.01441f
C63 VN.n32 B 0.017573f
C64 VN.n33 B 0.017573f
C65 VN.n34 B 0.017573f
C66 VN.n35 B 0.032752f
C67 VN.n36 B 0.032752f
C68 VN.n37 B 0.018522f
C69 VN.n38 B 0.028363f
C70 VN.n39 B 1.20592f
C71 VTAIL.t3 B 0.304084f
C72 VTAIL.t4 B 0.304084f
C73 VTAIL.n0 B 2.69462f
C74 VTAIL.n1 B 0.462887f
C75 VTAIL.t10 B 3.44191f
C76 VTAIL.n2 B 0.737461f
C77 VTAIL.t6 B 0.304084f
C78 VTAIL.t8 B 0.304084f
C79 VTAIL.n3 B 2.69462f
C80 VTAIL.n4 B 2.39911f
C81 VTAIL.t2 B 0.304084f
C82 VTAIL.t1 B 0.304084f
C83 VTAIL.n5 B 2.69463f
C84 VTAIL.n6 B 2.39911f
C85 VTAIL.t0 B 3.44191f
C86 VTAIL.n7 B 0.737458f
C87 VTAIL.t9 B 0.304084f
C88 VTAIL.t11 B 0.304084f
C89 VTAIL.n8 B 2.69463f
C90 VTAIL.n9 B 0.655421f
C91 VTAIL.t7 B 3.44191f
C92 VTAIL.n10 B 2.21861f
C93 VTAIL.t5 B 3.44191f
C94 VTAIL.n11 B 2.14861f
C95 VDD1.t3 B 3.2775f
C96 VDD1.t1 B 3.2765f
C97 VDD1.t5 B 0.280861f
C98 VDD1.t4 B 0.280861f
C99 VDD1.n0 B 2.55761f
C100 VDD1.n1 B 3.29574f
C101 VDD1.t2 B 0.280861f
C102 VDD1.t0 B 0.280861f
C103 VDD1.n2 B 2.55134f
C104 VDD1.n3 B 2.9652f
C105 VP.t1 B 3.01963f
C106 VP.n0 B 1.10949f
C107 VP.n1 B 0.017835f
C108 VP.n2 B 0.034814f
C109 VP.n3 B 0.017835f
C110 VP.n4 B 0.03324f
C111 VP.n5 B 0.017835f
C112 VP.t3 B 3.01963f
C113 VP.n6 B 0.035873f
C114 VP.n7 B 0.017835f
C115 VP.n8 B 0.03324f
C116 VP.t4 B 3.01963f
C117 VP.n9 B 1.10949f
C118 VP.n10 B 0.017835f
C119 VP.n11 B 0.034814f
C120 VP.n12 B 0.017835f
C121 VP.n13 B 0.03324f
C122 VP.t2 B 3.29873f
C123 VP.t0 B 3.01963f
C124 VP.n14 B 1.11679f
C125 VP.n15 B 1.06259f
C126 VP.n16 B 0.227708f
C127 VP.n17 B 0.017835f
C128 VP.n18 B 0.03324f
C129 VP.n19 B 0.035873f
C130 VP.n20 B 0.014625f
C131 VP.n21 B 0.017835f
C132 VP.n22 B 0.017835f
C133 VP.n23 B 0.017835f
C134 VP.n24 B 0.03324f
C135 VP.n25 B 0.03324f
C136 VP.n26 B 0.018799f
C137 VP.n27 B 0.028786f
C138 VP.n28 B 1.2169f
C139 VP.n29 B 1.22823f
C140 VP.t5 B 3.01963f
C141 VP.n30 B 1.10949f
C142 VP.n31 B 0.018799f
C143 VP.n32 B 0.028786f
C144 VP.n33 B 0.017835f
C145 VP.n34 B 0.017835f
C146 VP.n35 B 0.03324f
C147 VP.n36 B 0.034814f
C148 VP.n37 B 0.014625f
C149 VP.n38 B 0.017835f
C150 VP.n39 B 0.017835f
C151 VP.n40 B 0.017835f
C152 VP.n41 B 0.03324f
C153 VP.n42 B 0.03324f
C154 VP.n43 B 1.0605f
C155 VP.n44 B 0.017835f
C156 VP.n45 B 0.017835f
C157 VP.n46 B 0.017835f
C158 VP.n47 B 0.03324f
C159 VP.n48 B 0.035873f
C160 VP.n49 B 0.014625f
C161 VP.n50 B 0.017835f
C162 VP.n51 B 0.017835f
C163 VP.n52 B 0.017835f
C164 VP.n53 B 0.03324f
C165 VP.n54 B 0.03324f
C166 VP.n55 B 0.018799f
C167 VP.n56 B 0.028786f
C168 VP.n57 B 0.054068f
.ends

