* NGSPICE file created from diff_pair_sample_1479.ext - technology: sky130A

.subckt diff_pair_sample_1479 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.4 as=0 ps=0 w=2.31 l=3.96
X1 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.4 as=0 ps=0 w=2.31 l=3.96
X2 VDD2.t1 VN.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.4 as=0.9009 ps=5.4 w=2.31 l=3.96
X3 VDD1.t1 VP.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.4 as=0.9009 ps=5.4 w=2.31 l=3.96
X4 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.4 as=0 ps=0 w=2.31 l=3.96
X5 VDD2.t0 VN.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.4 as=0.9009 ps=5.4 w=2.31 l=3.96
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.4 as=0.9009 ps=5.4 w=2.31 l=3.96
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9009 pd=5.4 as=0 ps=0 w=2.31 l=3.96
R0 B.n460 B.n459 585
R1 B.n156 B.n81 585
R2 B.n155 B.n154 585
R3 B.n153 B.n152 585
R4 B.n151 B.n150 585
R5 B.n149 B.n148 585
R6 B.n147 B.n146 585
R7 B.n145 B.n144 585
R8 B.n143 B.n142 585
R9 B.n141 B.n140 585
R10 B.n139 B.n138 585
R11 B.n137 B.n136 585
R12 B.n135 B.n134 585
R13 B.n132 B.n131 585
R14 B.n130 B.n129 585
R15 B.n128 B.n127 585
R16 B.n126 B.n125 585
R17 B.n124 B.n123 585
R18 B.n122 B.n121 585
R19 B.n120 B.n119 585
R20 B.n118 B.n117 585
R21 B.n116 B.n115 585
R22 B.n114 B.n113 585
R23 B.n111 B.n110 585
R24 B.n109 B.n108 585
R25 B.n107 B.n106 585
R26 B.n105 B.n104 585
R27 B.n103 B.n102 585
R28 B.n101 B.n100 585
R29 B.n99 B.n98 585
R30 B.n97 B.n96 585
R31 B.n95 B.n94 585
R32 B.n93 B.n92 585
R33 B.n91 B.n90 585
R34 B.n89 B.n88 585
R35 B.n87 B.n86 585
R36 B.n458 B.n63 585
R37 B.n463 B.n63 585
R38 B.n457 B.n62 585
R39 B.n464 B.n62 585
R40 B.n456 B.n455 585
R41 B.n455 B.n58 585
R42 B.n454 B.n57 585
R43 B.n470 B.n57 585
R44 B.n453 B.n56 585
R45 B.n471 B.n56 585
R46 B.n452 B.n55 585
R47 B.n472 B.n55 585
R48 B.n451 B.n450 585
R49 B.n450 B.n51 585
R50 B.n449 B.n50 585
R51 B.n478 B.n50 585
R52 B.n448 B.n49 585
R53 B.n479 B.n49 585
R54 B.n447 B.n48 585
R55 B.n480 B.n48 585
R56 B.n446 B.n445 585
R57 B.n445 B.n44 585
R58 B.n444 B.n43 585
R59 B.n486 B.n43 585
R60 B.n443 B.n42 585
R61 B.n487 B.n42 585
R62 B.n442 B.n41 585
R63 B.n488 B.n41 585
R64 B.n441 B.n440 585
R65 B.n440 B.n37 585
R66 B.n439 B.n36 585
R67 B.n494 B.n36 585
R68 B.n438 B.n35 585
R69 B.n495 B.n35 585
R70 B.n437 B.n34 585
R71 B.n496 B.n34 585
R72 B.n436 B.n435 585
R73 B.n435 B.n30 585
R74 B.n434 B.n29 585
R75 B.n502 B.n29 585
R76 B.n433 B.n28 585
R77 B.n503 B.n28 585
R78 B.n432 B.n27 585
R79 B.n504 B.n27 585
R80 B.n431 B.n430 585
R81 B.n430 B.n23 585
R82 B.n429 B.n22 585
R83 B.n510 B.n22 585
R84 B.n428 B.n21 585
R85 B.n511 B.n21 585
R86 B.n427 B.n20 585
R87 B.n512 B.n20 585
R88 B.n426 B.n425 585
R89 B.n425 B.n16 585
R90 B.n424 B.n15 585
R91 B.n518 B.n15 585
R92 B.n423 B.n14 585
R93 B.n519 B.n14 585
R94 B.n422 B.n13 585
R95 B.n520 B.n13 585
R96 B.n421 B.n420 585
R97 B.n420 B.n12 585
R98 B.n419 B.n418 585
R99 B.n419 B.n8 585
R100 B.n417 B.n7 585
R101 B.n527 B.n7 585
R102 B.n416 B.n6 585
R103 B.n528 B.n6 585
R104 B.n415 B.n5 585
R105 B.n529 B.n5 585
R106 B.n414 B.n413 585
R107 B.n413 B.n4 585
R108 B.n412 B.n157 585
R109 B.n412 B.n411 585
R110 B.n402 B.n158 585
R111 B.n159 B.n158 585
R112 B.n404 B.n403 585
R113 B.n405 B.n404 585
R114 B.n401 B.n164 585
R115 B.n164 B.n163 585
R116 B.n400 B.n399 585
R117 B.n399 B.n398 585
R118 B.n166 B.n165 585
R119 B.n167 B.n166 585
R120 B.n391 B.n390 585
R121 B.n392 B.n391 585
R122 B.n389 B.n172 585
R123 B.n172 B.n171 585
R124 B.n388 B.n387 585
R125 B.n387 B.n386 585
R126 B.n174 B.n173 585
R127 B.n175 B.n174 585
R128 B.n379 B.n378 585
R129 B.n380 B.n379 585
R130 B.n377 B.n180 585
R131 B.n180 B.n179 585
R132 B.n376 B.n375 585
R133 B.n375 B.n374 585
R134 B.n182 B.n181 585
R135 B.n183 B.n182 585
R136 B.n367 B.n366 585
R137 B.n368 B.n367 585
R138 B.n365 B.n188 585
R139 B.n188 B.n187 585
R140 B.n364 B.n363 585
R141 B.n363 B.n362 585
R142 B.n190 B.n189 585
R143 B.n191 B.n190 585
R144 B.n355 B.n354 585
R145 B.n356 B.n355 585
R146 B.n353 B.n196 585
R147 B.n196 B.n195 585
R148 B.n352 B.n351 585
R149 B.n351 B.n350 585
R150 B.n198 B.n197 585
R151 B.n199 B.n198 585
R152 B.n343 B.n342 585
R153 B.n344 B.n343 585
R154 B.n341 B.n204 585
R155 B.n204 B.n203 585
R156 B.n340 B.n339 585
R157 B.n339 B.n338 585
R158 B.n206 B.n205 585
R159 B.n207 B.n206 585
R160 B.n331 B.n330 585
R161 B.n332 B.n331 585
R162 B.n329 B.n212 585
R163 B.n212 B.n211 585
R164 B.n328 B.n327 585
R165 B.n327 B.n326 585
R166 B.n214 B.n213 585
R167 B.n215 B.n214 585
R168 B.n319 B.n318 585
R169 B.n320 B.n319 585
R170 B.n317 B.n220 585
R171 B.n220 B.n219 585
R172 B.n312 B.n311 585
R173 B.n310 B.n240 585
R174 B.n309 B.n239 585
R175 B.n314 B.n239 585
R176 B.n308 B.n307 585
R177 B.n306 B.n305 585
R178 B.n304 B.n303 585
R179 B.n302 B.n301 585
R180 B.n300 B.n299 585
R181 B.n298 B.n297 585
R182 B.n296 B.n295 585
R183 B.n294 B.n293 585
R184 B.n292 B.n291 585
R185 B.n290 B.n289 585
R186 B.n288 B.n287 585
R187 B.n286 B.n285 585
R188 B.n284 B.n283 585
R189 B.n282 B.n281 585
R190 B.n280 B.n279 585
R191 B.n278 B.n277 585
R192 B.n276 B.n275 585
R193 B.n274 B.n273 585
R194 B.n272 B.n271 585
R195 B.n270 B.n269 585
R196 B.n268 B.n267 585
R197 B.n266 B.n265 585
R198 B.n264 B.n263 585
R199 B.n262 B.n261 585
R200 B.n260 B.n259 585
R201 B.n258 B.n257 585
R202 B.n256 B.n255 585
R203 B.n254 B.n253 585
R204 B.n252 B.n251 585
R205 B.n250 B.n249 585
R206 B.n248 B.n247 585
R207 B.n222 B.n221 585
R208 B.n316 B.n315 585
R209 B.n315 B.n314 585
R210 B.n218 B.n217 585
R211 B.n219 B.n218 585
R212 B.n322 B.n321 585
R213 B.n321 B.n320 585
R214 B.n323 B.n216 585
R215 B.n216 B.n215 585
R216 B.n325 B.n324 585
R217 B.n326 B.n325 585
R218 B.n210 B.n209 585
R219 B.n211 B.n210 585
R220 B.n334 B.n333 585
R221 B.n333 B.n332 585
R222 B.n335 B.n208 585
R223 B.n208 B.n207 585
R224 B.n337 B.n336 585
R225 B.n338 B.n337 585
R226 B.n202 B.n201 585
R227 B.n203 B.n202 585
R228 B.n346 B.n345 585
R229 B.n345 B.n344 585
R230 B.n347 B.n200 585
R231 B.n200 B.n199 585
R232 B.n349 B.n348 585
R233 B.n350 B.n349 585
R234 B.n194 B.n193 585
R235 B.n195 B.n194 585
R236 B.n358 B.n357 585
R237 B.n357 B.n356 585
R238 B.n359 B.n192 585
R239 B.n192 B.n191 585
R240 B.n361 B.n360 585
R241 B.n362 B.n361 585
R242 B.n186 B.n185 585
R243 B.n187 B.n186 585
R244 B.n370 B.n369 585
R245 B.n369 B.n368 585
R246 B.n371 B.n184 585
R247 B.n184 B.n183 585
R248 B.n373 B.n372 585
R249 B.n374 B.n373 585
R250 B.n178 B.n177 585
R251 B.n179 B.n178 585
R252 B.n382 B.n381 585
R253 B.n381 B.n380 585
R254 B.n383 B.n176 585
R255 B.n176 B.n175 585
R256 B.n385 B.n384 585
R257 B.n386 B.n385 585
R258 B.n170 B.n169 585
R259 B.n171 B.n170 585
R260 B.n394 B.n393 585
R261 B.n393 B.n392 585
R262 B.n395 B.n168 585
R263 B.n168 B.n167 585
R264 B.n397 B.n396 585
R265 B.n398 B.n397 585
R266 B.n162 B.n161 585
R267 B.n163 B.n162 585
R268 B.n407 B.n406 585
R269 B.n406 B.n405 585
R270 B.n408 B.n160 585
R271 B.n160 B.n159 585
R272 B.n410 B.n409 585
R273 B.n411 B.n410 585
R274 B.n3 B.n0 585
R275 B.n4 B.n3 585
R276 B.n526 B.n1 585
R277 B.n527 B.n526 585
R278 B.n525 B.n524 585
R279 B.n525 B.n8 585
R280 B.n523 B.n9 585
R281 B.n12 B.n9 585
R282 B.n522 B.n521 585
R283 B.n521 B.n520 585
R284 B.n11 B.n10 585
R285 B.n519 B.n11 585
R286 B.n517 B.n516 585
R287 B.n518 B.n517 585
R288 B.n515 B.n17 585
R289 B.n17 B.n16 585
R290 B.n514 B.n513 585
R291 B.n513 B.n512 585
R292 B.n19 B.n18 585
R293 B.n511 B.n19 585
R294 B.n509 B.n508 585
R295 B.n510 B.n509 585
R296 B.n507 B.n24 585
R297 B.n24 B.n23 585
R298 B.n506 B.n505 585
R299 B.n505 B.n504 585
R300 B.n26 B.n25 585
R301 B.n503 B.n26 585
R302 B.n501 B.n500 585
R303 B.n502 B.n501 585
R304 B.n499 B.n31 585
R305 B.n31 B.n30 585
R306 B.n498 B.n497 585
R307 B.n497 B.n496 585
R308 B.n33 B.n32 585
R309 B.n495 B.n33 585
R310 B.n493 B.n492 585
R311 B.n494 B.n493 585
R312 B.n491 B.n38 585
R313 B.n38 B.n37 585
R314 B.n490 B.n489 585
R315 B.n489 B.n488 585
R316 B.n40 B.n39 585
R317 B.n487 B.n40 585
R318 B.n485 B.n484 585
R319 B.n486 B.n485 585
R320 B.n483 B.n45 585
R321 B.n45 B.n44 585
R322 B.n482 B.n481 585
R323 B.n481 B.n480 585
R324 B.n47 B.n46 585
R325 B.n479 B.n47 585
R326 B.n477 B.n476 585
R327 B.n478 B.n477 585
R328 B.n475 B.n52 585
R329 B.n52 B.n51 585
R330 B.n474 B.n473 585
R331 B.n473 B.n472 585
R332 B.n54 B.n53 585
R333 B.n471 B.n54 585
R334 B.n469 B.n468 585
R335 B.n470 B.n469 585
R336 B.n467 B.n59 585
R337 B.n59 B.n58 585
R338 B.n466 B.n465 585
R339 B.n465 B.n464 585
R340 B.n61 B.n60 585
R341 B.n463 B.n61 585
R342 B.n530 B.n529 585
R343 B.n528 B.n2 585
R344 B.n86 B.n61 458.866
R345 B.n460 B.n63 458.866
R346 B.n315 B.n220 458.866
R347 B.n312 B.n218 458.866
R348 B.n462 B.n461 256.663
R349 B.n462 B.n80 256.663
R350 B.n462 B.n79 256.663
R351 B.n462 B.n78 256.663
R352 B.n462 B.n77 256.663
R353 B.n462 B.n76 256.663
R354 B.n462 B.n75 256.663
R355 B.n462 B.n74 256.663
R356 B.n462 B.n73 256.663
R357 B.n462 B.n72 256.663
R358 B.n462 B.n71 256.663
R359 B.n462 B.n70 256.663
R360 B.n462 B.n69 256.663
R361 B.n462 B.n68 256.663
R362 B.n462 B.n67 256.663
R363 B.n462 B.n66 256.663
R364 B.n462 B.n65 256.663
R365 B.n462 B.n64 256.663
R366 B.n314 B.n313 256.663
R367 B.n314 B.n223 256.663
R368 B.n314 B.n224 256.663
R369 B.n314 B.n225 256.663
R370 B.n314 B.n226 256.663
R371 B.n314 B.n227 256.663
R372 B.n314 B.n228 256.663
R373 B.n314 B.n229 256.663
R374 B.n314 B.n230 256.663
R375 B.n314 B.n231 256.663
R376 B.n314 B.n232 256.663
R377 B.n314 B.n233 256.663
R378 B.n314 B.n234 256.663
R379 B.n314 B.n235 256.663
R380 B.n314 B.n236 256.663
R381 B.n314 B.n237 256.663
R382 B.n314 B.n238 256.663
R383 B.n532 B.n531 256.663
R384 B.n84 B.t2 223.522
R385 B.n82 B.t6 223.522
R386 B.n244 B.t13 223.522
R387 B.n241 B.t9 223.522
R388 B.n82 B.t7 170.613
R389 B.n244 B.t15 170.613
R390 B.n84 B.t4 170.613
R391 B.n241 B.t12 170.613
R392 B.n314 B.n219 163.876
R393 B.n463 B.n462 163.876
R394 B.n90 B.n89 163.367
R395 B.n94 B.n93 163.367
R396 B.n98 B.n97 163.367
R397 B.n102 B.n101 163.367
R398 B.n106 B.n105 163.367
R399 B.n110 B.n109 163.367
R400 B.n115 B.n114 163.367
R401 B.n119 B.n118 163.367
R402 B.n123 B.n122 163.367
R403 B.n127 B.n126 163.367
R404 B.n131 B.n130 163.367
R405 B.n136 B.n135 163.367
R406 B.n140 B.n139 163.367
R407 B.n144 B.n143 163.367
R408 B.n148 B.n147 163.367
R409 B.n152 B.n151 163.367
R410 B.n154 B.n81 163.367
R411 B.n319 B.n220 163.367
R412 B.n319 B.n214 163.367
R413 B.n327 B.n214 163.367
R414 B.n327 B.n212 163.367
R415 B.n331 B.n212 163.367
R416 B.n331 B.n206 163.367
R417 B.n339 B.n206 163.367
R418 B.n339 B.n204 163.367
R419 B.n343 B.n204 163.367
R420 B.n343 B.n198 163.367
R421 B.n351 B.n198 163.367
R422 B.n351 B.n196 163.367
R423 B.n355 B.n196 163.367
R424 B.n355 B.n190 163.367
R425 B.n363 B.n190 163.367
R426 B.n363 B.n188 163.367
R427 B.n367 B.n188 163.367
R428 B.n367 B.n182 163.367
R429 B.n375 B.n182 163.367
R430 B.n375 B.n180 163.367
R431 B.n379 B.n180 163.367
R432 B.n379 B.n174 163.367
R433 B.n387 B.n174 163.367
R434 B.n387 B.n172 163.367
R435 B.n391 B.n172 163.367
R436 B.n391 B.n166 163.367
R437 B.n399 B.n166 163.367
R438 B.n399 B.n164 163.367
R439 B.n404 B.n164 163.367
R440 B.n404 B.n158 163.367
R441 B.n412 B.n158 163.367
R442 B.n413 B.n412 163.367
R443 B.n413 B.n5 163.367
R444 B.n6 B.n5 163.367
R445 B.n7 B.n6 163.367
R446 B.n419 B.n7 163.367
R447 B.n420 B.n419 163.367
R448 B.n420 B.n13 163.367
R449 B.n14 B.n13 163.367
R450 B.n15 B.n14 163.367
R451 B.n425 B.n15 163.367
R452 B.n425 B.n20 163.367
R453 B.n21 B.n20 163.367
R454 B.n22 B.n21 163.367
R455 B.n430 B.n22 163.367
R456 B.n430 B.n27 163.367
R457 B.n28 B.n27 163.367
R458 B.n29 B.n28 163.367
R459 B.n435 B.n29 163.367
R460 B.n435 B.n34 163.367
R461 B.n35 B.n34 163.367
R462 B.n36 B.n35 163.367
R463 B.n440 B.n36 163.367
R464 B.n440 B.n41 163.367
R465 B.n42 B.n41 163.367
R466 B.n43 B.n42 163.367
R467 B.n445 B.n43 163.367
R468 B.n445 B.n48 163.367
R469 B.n49 B.n48 163.367
R470 B.n50 B.n49 163.367
R471 B.n450 B.n50 163.367
R472 B.n450 B.n55 163.367
R473 B.n56 B.n55 163.367
R474 B.n57 B.n56 163.367
R475 B.n455 B.n57 163.367
R476 B.n455 B.n62 163.367
R477 B.n63 B.n62 163.367
R478 B.n240 B.n239 163.367
R479 B.n307 B.n239 163.367
R480 B.n305 B.n304 163.367
R481 B.n301 B.n300 163.367
R482 B.n297 B.n296 163.367
R483 B.n293 B.n292 163.367
R484 B.n289 B.n288 163.367
R485 B.n285 B.n284 163.367
R486 B.n281 B.n280 163.367
R487 B.n277 B.n276 163.367
R488 B.n273 B.n272 163.367
R489 B.n269 B.n268 163.367
R490 B.n265 B.n264 163.367
R491 B.n261 B.n260 163.367
R492 B.n257 B.n256 163.367
R493 B.n253 B.n252 163.367
R494 B.n249 B.n248 163.367
R495 B.n315 B.n222 163.367
R496 B.n321 B.n218 163.367
R497 B.n321 B.n216 163.367
R498 B.n325 B.n216 163.367
R499 B.n325 B.n210 163.367
R500 B.n333 B.n210 163.367
R501 B.n333 B.n208 163.367
R502 B.n337 B.n208 163.367
R503 B.n337 B.n202 163.367
R504 B.n345 B.n202 163.367
R505 B.n345 B.n200 163.367
R506 B.n349 B.n200 163.367
R507 B.n349 B.n194 163.367
R508 B.n357 B.n194 163.367
R509 B.n357 B.n192 163.367
R510 B.n361 B.n192 163.367
R511 B.n361 B.n186 163.367
R512 B.n369 B.n186 163.367
R513 B.n369 B.n184 163.367
R514 B.n373 B.n184 163.367
R515 B.n373 B.n178 163.367
R516 B.n381 B.n178 163.367
R517 B.n381 B.n176 163.367
R518 B.n385 B.n176 163.367
R519 B.n385 B.n170 163.367
R520 B.n393 B.n170 163.367
R521 B.n393 B.n168 163.367
R522 B.n397 B.n168 163.367
R523 B.n397 B.n162 163.367
R524 B.n406 B.n162 163.367
R525 B.n406 B.n160 163.367
R526 B.n410 B.n160 163.367
R527 B.n410 B.n3 163.367
R528 B.n530 B.n3 163.367
R529 B.n526 B.n2 163.367
R530 B.n526 B.n525 163.367
R531 B.n525 B.n9 163.367
R532 B.n521 B.n9 163.367
R533 B.n521 B.n11 163.367
R534 B.n517 B.n11 163.367
R535 B.n517 B.n17 163.367
R536 B.n513 B.n17 163.367
R537 B.n513 B.n19 163.367
R538 B.n509 B.n19 163.367
R539 B.n509 B.n24 163.367
R540 B.n505 B.n24 163.367
R541 B.n505 B.n26 163.367
R542 B.n501 B.n26 163.367
R543 B.n501 B.n31 163.367
R544 B.n497 B.n31 163.367
R545 B.n497 B.n33 163.367
R546 B.n493 B.n33 163.367
R547 B.n493 B.n38 163.367
R548 B.n489 B.n38 163.367
R549 B.n489 B.n40 163.367
R550 B.n485 B.n40 163.367
R551 B.n485 B.n45 163.367
R552 B.n481 B.n45 163.367
R553 B.n481 B.n47 163.367
R554 B.n477 B.n47 163.367
R555 B.n477 B.n52 163.367
R556 B.n473 B.n52 163.367
R557 B.n473 B.n54 163.367
R558 B.n469 B.n54 163.367
R559 B.n469 B.n59 163.367
R560 B.n465 B.n59 163.367
R561 B.n465 B.n61 163.367
R562 B.n320 B.n219 98.6162
R563 B.n320 B.n215 98.6162
R564 B.n326 B.n215 98.6162
R565 B.n326 B.n211 98.6162
R566 B.n332 B.n211 98.6162
R567 B.n332 B.n207 98.6162
R568 B.n338 B.n207 98.6162
R569 B.n338 B.n203 98.6162
R570 B.n344 B.n203 98.6162
R571 B.n350 B.n199 98.6162
R572 B.n350 B.n195 98.6162
R573 B.n356 B.n195 98.6162
R574 B.n356 B.n191 98.6162
R575 B.n362 B.n191 98.6162
R576 B.n362 B.n187 98.6162
R577 B.n368 B.n187 98.6162
R578 B.n368 B.n183 98.6162
R579 B.n374 B.n183 98.6162
R580 B.n374 B.n179 98.6162
R581 B.n380 B.n179 98.6162
R582 B.n380 B.n175 98.6162
R583 B.n386 B.n175 98.6162
R584 B.n386 B.n171 98.6162
R585 B.n392 B.n171 98.6162
R586 B.n398 B.n167 98.6162
R587 B.n398 B.n163 98.6162
R588 B.n405 B.n163 98.6162
R589 B.n405 B.n159 98.6162
R590 B.n411 B.n159 98.6162
R591 B.n411 B.n4 98.6162
R592 B.n529 B.n4 98.6162
R593 B.n529 B.n528 98.6162
R594 B.n528 B.n527 98.6162
R595 B.n527 B.n8 98.6162
R596 B.n12 B.n8 98.6162
R597 B.n520 B.n12 98.6162
R598 B.n520 B.n519 98.6162
R599 B.n519 B.n518 98.6162
R600 B.n518 B.n16 98.6162
R601 B.n512 B.n511 98.6162
R602 B.n511 B.n510 98.6162
R603 B.n510 B.n23 98.6162
R604 B.n504 B.n23 98.6162
R605 B.n504 B.n503 98.6162
R606 B.n503 B.n502 98.6162
R607 B.n502 B.n30 98.6162
R608 B.n496 B.n30 98.6162
R609 B.n496 B.n495 98.6162
R610 B.n495 B.n494 98.6162
R611 B.n494 B.n37 98.6162
R612 B.n488 B.n37 98.6162
R613 B.n488 B.n487 98.6162
R614 B.n487 B.n486 98.6162
R615 B.n486 B.n44 98.6162
R616 B.n480 B.n479 98.6162
R617 B.n479 B.n478 98.6162
R618 B.n478 B.n51 98.6162
R619 B.n472 B.n51 98.6162
R620 B.n472 B.n471 98.6162
R621 B.n471 B.n470 98.6162
R622 B.n470 B.n58 98.6162
R623 B.n464 B.n58 98.6162
R624 B.n464 B.n463 98.6162
R625 B.n83 B.t8 87.4125
R626 B.n245 B.t14 87.4125
R627 B.n85 B.t5 87.4123
R628 B.n242 B.t11 87.4123
R629 B.n85 B.n84 83.2005
R630 B.n83 B.n82 83.2005
R631 B.n245 B.n244 83.2005
R632 B.n242 B.n241 83.2005
R633 B.n344 B.t10 75.4125
R634 B.n480 B.t3 75.4125
R635 B.n86 B.n64 71.676
R636 B.n90 B.n65 71.676
R637 B.n94 B.n66 71.676
R638 B.n98 B.n67 71.676
R639 B.n102 B.n68 71.676
R640 B.n106 B.n69 71.676
R641 B.n110 B.n70 71.676
R642 B.n115 B.n71 71.676
R643 B.n119 B.n72 71.676
R644 B.n123 B.n73 71.676
R645 B.n127 B.n74 71.676
R646 B.n131 B.n75 71.676
R647 B.n136 B.n76 71.676
R648 B.n140 B.n77 71.676
R649 B.n144 B.n78 71.676
R650 B.n148 B.n79 71.676
R651 B.n152 B.n80 71.676
R652 B.n461 B.n81 71.676
R653 B.n461 B.n460 71.676
R654 B.n154 B.n80 71.676
R655 B.n151 B.n79 71.676
R656 B.n147 B.n78 71.676
R657 B.n143 B.n77 71.676
R658 B.n139 B.n76 71.676
R659 B.n135 B.n75 71.676
R660 B.n130 B.n74 71.676
R661 B.n126 B.n73 71.676
R662 B.n122 B.n72 71.676
R663 B.n118 B.n71 71.676
R664 B.n114 B.n70 71.676
R665 B.n109 B.n69 71.676
R666 B.n105 B.n68 71.676
R667 B.n101 B.n67 71.676
R668 B.n97 B.n66 71.676
R669 B.n93 B.n65 71.676
R670 B.n89 B.n64 71.676
R671 B.n313 B.n312 71.676
R672 B.n307 B.n223 71.676
R673 B.n304 B.n224 71.676
R674 B.n300 B.n225 71.676
R675 B.n296 B.n226 71.676
R676 B.n292 B.n227 71.676
R677 B.n288 B.n228 71.676
R678 B.n284 B.n229 71.676
R679 B.n280 B.n230 71.676
R680 B.n276 B.n231 71.676
R681 B.n272 B.n232 71.676
R682 B.n268 B.n233 71.676
R683 B.n264 B.n234 71.676
R684 B.n260 B.n235 71.676
R685 B.n256 B.n236 71.676
R686 B.n252 B.n237 71.676
R687 B.n248 B.n238 71.676
R688 B.n313 B.n240 71.676
R689 B.n305 B.n223 71.676
R690 B.n301 B.n224 71.676
R691 B.n297 B.n225 71.676
R692 B.n293 B.n226 71.676
R693 B.n289 B.n227 71.676
R694 B.n285 B.n228 71.676
R695 B.n281 B.n229 71.676
R696 B.n277 B.n230 71.676
R697 B.n273 B.n231 71.676
R698 B.n269 B.n232 71.676
R699 B.n265 B.n233 71.676
R700 B.n261 B.n234 71.676
R701 B.n257 B.n235 71.676
R702 B.n253 B.n236 71.676
R703 B.n249 B.n237 71.676
R704 B.n238 B.n222 71.676
R705 B.n531 B.n530 71.676
R706 B.n531 B.n2 71.676
R707 B.n112 B.n85 59.5399
R708 B.n133 B.n83 59.5399
R709 B.n246 B.n245 59.5399
R710 B.n243 B.n242 59.5399
R711 B.n392 B.t0 58.0097
R712 B.n512 B.t1 58.0097
R713 B.t0 B.n167 40.607
R714 B.t1 B.n16 40.607
R715 B.n311 B.n217 29.8151
R716 B.n317 B.n316 29.8151
R717 B.n459 B.n458 29.8151
R718 B.n87 B.n60 29.8151
R719 B.t10 B.n199 23.2042
R720 B.t3 B.n44 23.2042
R721 B B.n532 18.0485
R722 B.n322 B.n217 10.6151
R723 B.n323 B.n322 10.6151
R724 B.n324 B.n323 10.6151
R725 B.n324 B.n209 10.6151
R726 B.n334 B.n209 10.6151
R727 B.n335 B.n334 10.6151
R728 B.n336 B.n335 10.6151
R729 B.n336 B.n201 10.6151
R730 B.n346 B.n201 10.6151
R731 B.n347 B.n346 10.6151
R732 B.n348 B.n347 10.6151
R733 B.n348 B.n193 10.6151
R734 B.n358 B.n193 10.6151
R735 B.n359 B.n358 10.6151
R736 B.n360 B.n359 10.6151
R737 B.n360 B.n185 10.6151
R738 B.n370 B.n185 10.6151
R739 B.n371 B.n370 10.6151
R740 B.n372 B.n371 10.6151
R741 B.n372 B.n177 10.6151
R742 B.n382 B.n177 10.6151
R743 B.n383 B.n382 10.6151
R744 B.n384 B.n383 10.6151
R745 B.n384 B.n169 10.6151
R746 B.n394 B.n169 10.6151
R747 B.n395 B.n394 10.6151
R748 B.n396 B.n395 10.6151
R749 B.n396 B.n161 10.6151
R750 B.n407 B.n161 10.6151
R751 B.n408 B.n407 10.6151
R752 B.n409 B.n408 10.6151
R753 B.n409 B.n0 10.6151
R754 B.n311 B.n310 10.6151
R755 B.n310 B.n309 10.6151
R756 B.n309 B.n308 10.6151
R757 B.n308 B.n306 10.6151
R758 B.n306 B.n303 10.6151
R759 B.n303 B.n302 10.6151
R760 B.n302 B.n299 10.6151
R761 B.n299 B.n298 10.6151
R762 B.n298 B.n295 10.6151
R763 B.n295 B.n294 10.6151
R764 B.n294 B.n291 10.6151
R765 B.n291 B.n290 10.6151
R766 B.n287 B.n286 10.6151
R767 B.n286 B.n283 10.6151
R768 B.n283 B.n282 10.6151
R769 B.n282 B.n279 10.6151
R770 B.n279 B.n278 10.6151
R771 B.n278 B.n275 10.6151
R772 B.n275 B.n274 10.6151
R773 B.n274 B.n271 10.6151
R774 B.n271 B.n270 10.6151
R775 B.n267 B.n266 10.6151
R776 B.n266 B.n263 10.6151
R777 B.n263 B.n262 10.6151
R778 B.n262 B.n259 10.6151
R779 B.n259 B.n258 10.6151
R780 B.n258 B.n255 10.6151
R781 B.n255 B.n254 10.6151
R782 B.n254 B.n251 10.6151
R783 B.n251 B.n250 10.6151
R784 B.n250 B.n247 10.6151
R785 B.n247 B.n221 10.6151
R786 B.n316 B.n221 10.6151
R787 B.n318 B.n317 10.6151
R788 B.n318 B.n213 10.6151
R789 B.n328 B.n213 10.6151
R790 B.n329 B.n328 10.6151
R791 B.n330 B.n329 10.6151
R792 B.n330 B.n205 10.6151
R793 B.n340 B.n205 10.6151
R794 B.n341 B.n340 10.6151
R795 B.n342 B.n341 10.6151
R796 B.n342 B.n197 10.6151
R797 B.n352 B.n197 10.6151
R798 B.n353 B.n352 10.6151
R799 B.n354 B.n353 10.6151
R800 B.n354 B.n189 10.6151
R801 B.n364 B.n189 10.6151
R802 B.n365 B.n364 10.6151
R803 B.n366 B.n365 10.6151
R804 B.n366 B.n181 10.6151
R805 B.n376 B.n181 10.6151
R806 B.n377 B.n376 10.6151
R807 B.n378 B.n377 10.6151
R808 B.n378 B.n173 10.6151
R809 B.n388 B.n173 10.6151
R810 B.n389 B.n388 10.6151
R811 B.n390 B.n389 10.6151
R812 B.n390 B.n165 10.6151
R813 B.n400 B.n165 10.6151
R814 B.n401 B.n400 10.6151
R815 B.n403 B.n401 10.6151
R816 B.n403 B.n402 10.6151
R817 B.n402 B.n157 10.6151
R818 B.n414 B.n157 10.6151
R819 B.n415 B.n414 10.6151
R820 B.n416 B.n415 10.6151
R821 B.n417 B.n416 10.6151
R822 B.n418 B.n417 10.6151
R823 B.n421 B.n418 10.6151
R824 B.n422 B.n421 10.6151
R825 B.n423 B.n422 10.6151
R826 B.n424 B.n423 10.6151
R827 B.n426 B.n424 10.6151
R828 B.n427 B.n426 10.6151
R829 B.n428 B.n427 10.6151
R830 B.n429 B.n428 10.6151
R831 B.n431 B.n429 10.6151
R832 B.n432 B.n431 10.6151
R833 B.n433 B.n432 10.6151
R834 B.n434 B.n433 10.6151
R835 B.n436 B.n434 10.6151
R836 B.n437 B.n436 10.6151
R837 B.n438 B.n437 10.6151
R838 B.n439 B.n438 10.6151
R839 B.n441 B.n439 10.6151
R840 B.n442 B.n441 10.6151
R841 B.n443 B.n442 10.6151
R842 B.n444 B.n443 10.6151
R843 B.n446 B.n444 10.6151
R844 B.n447 B.n446 10.6151
R845 B.n448 B.n447 10.6151
R846 B.n449 B.n448 10.6151
R847 B.n451 B.n449 10.6151
R848 B.n452 B.n451 10.6151
R849 B.n453 B.n452 10.6151
R850 B.n454 B.n453 10.6151
R851 B.n456 B.n454 10.6151
R852 B.n457 B.n456 10.6151
R853 B.n458 B.n457 10.6151
R854 B.n524 B.n1 10.6151
R855 B.n524 B.n523 10.6151
R856 B.n523 B.n522 10.6151
R857 B.n522 B.n10 10.6151
R858 B.n516 B.n10 10.6151
R859 B.n516 B.n515 10.6151
R860 B.n515 B.n514 10.6151
R861 B.n514 B.n18 10.6151
R862 B.n508 B.n18 10.6151
R863 B.n508 B.n507 10.6151
R864 B.n507 B.n506 10.6151
R865 B.n506 B.n25 10.6151
R866 B.n500 B.n25 10.6151
R867 B.n500 B.n499 10.6151
R868 B.n499 B.n498 10.6151
R869 B.n498 B.n32 10.6151
R870 B.n492 B.n32 10.6151
R871 B.n492 B.n491 10.6151
R872 B.n491 B.n490 10.6151
R873 B.n490 B.n39 10.6151
R874 B.n484 B.n39 10.6151
R875 B.n484 B.n483 10.6151
R876 B.n483 B.n482 10.6151
R877 B.n482 B.n46 10.6151
R878 B.n476 B.n46 10.6151
R879 B.n476 B.n475 10.6151
R880 B.n475 B.n474 10.6151
R881 B.n474 B.n53 10.6151
R882 B.n468 B.n53 10.6151
R883 B.n468 B.n467 10.6151
R884 B.n467 B.n466 10.6151
R885 B.n466 B.n60 10.6151
R886 B.n88 B.n87 10.6151
R887 B.n91 B.n88 10.6151
R888 B.n92 B.n91 10.6151
R889 B.n95 B.n92 10.6151
R890 B.n96 B.n95 10.6151
R891 B.n99 B.n96 10.6151
R892 B.n100 B.n99 10.6151
R893 B.n103 B.n100 10.6151
R894 B.n104 B.n103 10.6151
R895 B.n107 B.n104 10.6151
R896 B.n108 B.n107 10.6151
R897 B.n111 B.n108 10.6151
R898 B.n116 B.n113 10.6151
R899 B.n117 B.n116 10.6151
R900 B.n120 B.n117 10.6151
R901 B.n121 B.n120 10.6151
R902 B.n124 B.n121 10.6151
R903 B.n125 B.n124 10.6151
R904 B.n128 B.n125 10.6151
R905 B.n129 B.n128 10.6151
R906 B.n132 B.n129 10.6151
R907 B.n137 B.n134 10.6151
R908 B.n138 B.n137 10.6151
R909 B.n141 B.n138 10.6151
R910 B.n142 B.n141 10.6151
R911 B.n145 B.n142 10.6151
R912 B.n146 B.n145 10.6151
R913 B.n149 B.n146 10.6151
R914 B.n150 B.n149 10.6151
R915 B.n153 B.n150 10.6151
R916 B.n155 B.n153 10.6151
R917 B.n156 B.n155 10.6151
R918 B.n459 B.n156 10.6151
R919 B.n290 B.n243 9.36635
R920 B.n267 B.n246 9.36635
R921 B.n112 B.n111 9.36635
R922 B.n134 B.n133 9.36635
R923 B.n532 B.n0 8.11757
R924 B.n532 B.n1 8.11757
R925 B.n287 B.n243 1.24928
R926 B.n270 B.n246 1.24928
R927 B.n113 B.n112 1.24928
R928 B.n133 B.n132 1.24928
R929 VN VN.t1 89.8303
R930 VN VN.t0 49.7167
R931 VTAIL.n2 VTAIL.t3 82.6219
R932 VTAIL.n1 VTAIL.t1 82.6219
R933 VTAIL.n3 VTAIL.t0 82.6218
R934 VTAIL.n0 VTAIL.t2 82.6218
R935 VTAIL.n1 VTAIL.n0 21.7548
R936 VTAIL.n3 VTAIL.n2 18.0565
R937 VTAIL.n2 VTAIL.n1 2.31947
R938 VTAIL VTAIL.n0 1.45309
R939 VTAIL VTAIL.n3 0.866879
R940 VDD2.n0 VDD2.t1 132.347
R941 VDD2.n0 VDD2.t0 99.3007
R942 VDD2 VDD2.n0 0.983259
R943 VP.n0 VP.t1 90.018
R944 VP.n0 VP.t0 49.0959
R945 VP VP.n0 0.621237
R946 VDD1 VDD1.t1 133.798
R947 VDD1 VDD1.t0 100.284
C0 VN VTAIL 1.20824f
C1 VP VDD2 0.39618f
C2 VP VDD1 1.01781f
C3 VDD2 VDD1 0.827567f
C4 VP VTAIL 1.2225f
C5 VP VN 4.30617f
C6 VDD2 VTAIL 3.0149f
C7 VDD2 VN 0.777822f
C8 VDD1 VTAIL 2.95268f
C9 VDD1 VN 0.154628f
C10 VDD2 B 3.14801f
C11 VDD1 B 5.40717f
C12 VTAIL B 3.567771f
C13 VN B 9.29599f
C14 VP B 7.194712f
C15 VDD1.t0 B 0.282694f
C16 VDD1.t1 B 0.533948f
C17 VP.t1 B 1.42695f
C18 VP.t0 B 0.833044f
C19 VP.n0 B 1.93301f
C20 VDD2.t1 B 0.520789f
C21 VDD2.t0 B 0.286757f
C22 VDD2.n0 B 2.02655f
C23 VTAIL.t2 B 0.305475f
C24 VTAIL.n0 B 1.26349f
C25 VTAIL.t1 B 0.305476f
C26 VTAIL.n1 B 1.32428f
C27 VTAIL.t3 B 0.305476f
C28 VTAIL.n2 B 1.06477f
C29 VTAIL.t0 B 0.305475f
C30 VTAIL.n3 B 0.962845f
C31 VN.t0 B 0.830606f
C32 VN.t1 B 1.41502f
.ends

