* NGSPICE file created from diff_pair_sample_0899.ext - technology: sky130A

.subckt diff_pair_sample_0899 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t0 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.9087 pd=5.44 as=0.38445 ps=2.66 w=2.33 l=3.12
X1 VTAIL.t0 VP.t0 VDD1.t7 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.9087 pd=5.44 as=0.38445 ps=2.66 w=2.33 l=3.12
X2 VDD1.t6 VP.t1 VTAIL.t4 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.38445 ps=2.66 w=2.33 l=3.12
X3 B.t11 B.t9 B.t10 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.9087 pd=5.44 as=0 ps=0 w=2.33 l=3.12
X4 VDD2.t3 VN.t1 VTAIL.t14 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.9087 ps=5.44 w=2.33 l=3.12
X5 B.t8 B.t6 B.t7 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.9087 pd=5.44 as=0 ps=0 w=2.33 l=3.12
X6 VDD2.t7 VN.t2 VTAIL.t13 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.9087 ps=5.44 w=2.33 l=3.12
X7 B.t5 B.t3 B.t4 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.9087 pd=5.44 as=0 ps=0 w=2.33 l=3.12
X8 VTAIL.t2 VP.t2 VDD1.t5 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.38445 ps=2.66 w=2.33 l=3.12
X9 VTAIL.t12 VN.t3 VDD2.t6 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.38445 ps=2.66 w=2.33 l=3.12
X10 B.t2 B.t0 B.t1 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.9087 pd=5.44 as=0 ps=0 w=2.33 l=3.12
X11 VTAIL.t11 VN.t4 VDD2.t5 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.38445 ps=2.66 w=2.33 l=3.12
X12 VTAIL.t7 VP.t3 VDD1.t4 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.38445 ps=2.66 w=2.33 l=3.12
X13 VTAIL.t1 VP.t4 VDD1.t3 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.9087 pd=5.44 as=0.38445 ps=2.66 w=2.33 l=3.12
X14 VDD2.t1 VN.t5 VTAIL.t10 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.38445 ps=2.66 w=2.33 l=3.12
X15 VTAIL.t9 VN.t6 VDD2.t4 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.9087 pd=5.44 as=0.38445 ps=2.66 w=2.33 l=3.12
X16 VDD1.t2 VP.t5 VTAIL.t3 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.38445 ps=2.66 w=2.33 l=3.12
X17 VDD2.t2 VN.t7 VTAIL.t8 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.38445 ps=2.66 w=2.33 l=3.12
X18 VDD1.t1 VP.t6 VTAIL.t6 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.9087 ps=5.44 w=2.33 l=3.12
X19 VDD1.t0 VP.t7 VTAIL.t5 w_n4420_n1434# sky130_fd_pr__pfet_01v8 ad=0.38445 pd=2.66 as=0.9087 ps=5.44 w=2.33 l=3.12
R0 VN.n60 VN.n59 161.3
R1 VN.n58 VN.n32 161.3
R2 VN.n57 VN.n56 161.3
R3 VN.n55 VN.n33 161.3
R4 VN.n54 VN.n53 161.3
R5 VN.n52 VN.n34 161.3
R6 VN.n51 VN.n50 161.3
R7 VN.n49 VN.n48 161.3
R8 VN.n47 VN.n36 161.3
R9 VN.n46 VN.n45 161.3
R10 VN.n44 VN.n37 161.3
R11 VN.n43 VN.n42 161.3
R12 VN.n41 VN.n38 161.3
R13 VN.n29 VN.n28 161.3
R14 VN.n27 VN.n1 161.3
R15 VN.n26 VN.n25 161.3
R16 VN.n24 VN.n2 161.3
R17 VN.n23 VN.n22 161.3
R18 VN.n21 VN.n3 161.3
R19 VN.n20 VN.n19 161.3
R20 VN.n18 VN.n17 161.3
R21 VN.n16 VN.n5 161.3
R22 VN.n15 VN.n14 161.3
R23 VN.n13 VN.n6 161.3
R24 VN.n12 VN.n11 161.3
R25 VN.n10 VN.n7 161.3
R26 VN.n30 VN.n0 69.2705
R27 VN.n61 VN.n31 69.2705
R28 VN.n15 VN.n6 56.5193
R29 VN.n26 VN.n2 56.5193
R30 VN.n46 VN.n37 56.5193
R31 VN.n57 VN.n33 56.5193
R32 VN.n39 VN.t2 51.4115
R33 VN.n8 VN.t0 51.4115
R34 VN.n9 VN.n8 50.6608
R35 VN.n40 VN.n39 50.6608
R36 VN VN.n61 46.3314
R37 VN.n11 VN.n10 24.4675
R38 VN.n11 VN.n6 24.4675
R39 VN.n16 VN.n15 24.4675
R40 VN.n17 VN.n16 24.4675
R41 VN.n21 VN.n20 24.4675
R42 VN.n22 VN.n21 24.4675
R43 VN.n22 VN.n2 24.4675
R44 VN.n27 VN.n26 24.4675
R45 VN.n28 VN.n27 24.4675
R46 VN.n42 VN.n37 24.4675
R47 VN.n42 VN.n41 24.4675
R48 VN.n53 VN.n33 24.4675
R49 VN.n53 VN.n52 24.4675
R50 VN.n52 VN.n51 24.4675
R51 VN.n48 VN.n47 24.4675
R52 VN.n47 VN.n46 24.4675
R53 VN.n59 VN.n58 24.4675
R54 VN.n58 VN.n57 24.4675
R55 VN.n10 VN.n9 23.2442
R56 VN.n17 VN.n4 23.2442
R57 VN.n41 VN.n40 23.2442
R58 VN.n48 VN.n35 23.2442
R59 VN.n28 VN.n0 20.7975
R60 VN.n59 VN.n31 20.7975
R61 VN.n9 VN.t5 17.9983
R62 VN.n4 VN.t4 17.9983
R63 VN.n0 VN.t1 17.9983
R64 VN.n40 VN.t3 17.9983
R65 VN.n35 VN.t7 17.9983
R66 VN.n31 VN.t6 17.9983
R67 VN.n39 VN.n38 3.87633
R68 VN.n8 VN.n7 3.87633
R69 VN.n20 VN.n4 1.22385
R70 VN.n51 VN.n35 1.22385
R71 VN.n61 VN.n60 0.354971
R72 VN.n30 VN.n29 0.354971
R73 VN VN.n30 0.26696
R74 VN.n60 VN.n32 0.189894
R75 VN.n56 VN.n32 0.189894
R76 VN.n56 VN.n55 0.189894
R77 VN.n55 VN.n54 0.189894
R78 VN.n54 VN.n34 0.189894
R79 VN.n50 VN.n34 0.189894
R80 VN.n50 VN.n49 0.189894
R81 VN.n49 VN.n36 0.189894
R82 VN.n45 VN.n36 0.189894
R83 VN.n45 VN.n44 0.189894
R84 VN.n44 VN.n43 0.189894
R85 VN.n43 VN.n38 0.189894
R86 VN.n12 VN.n7 0.189894
R87 VN.n13 VN.n12 0.189894
R88 VN.n14 VN.n13 0.189894
R89 VN.n14 VN.n5 0.189894
R90 VN.n18 VN.n5 0.189894
R91 VN.n19 VN.n18 0.189894
R92 VN.n19 VN.n3 0.189894
R93 VN.n23 VN.n3 0.189894
R94 VN.n24 VN.n23 0.189894
R95 VN.n25 VN.n24 0.189894
R96 VN.n25 VN.n1 0.189894
R97 VN.n29 VN.n1 0.189894
R98 VDD2.n2 VDD2.n1 172.589
R99 VDD2.n2 VDD2.n0 172.589
R100 VDD2 VDD2.n5 172.587
R101 VDD2.n4 VDD2.n3 171.159
R102 VDD2.n4 VDD2.n2 39.1075
R103 VDD2.n5 VDD2.t6 13.9511
R104 VDD2.n5 VDD2.t7 13.9511
R105 VDD2.n3 VDD2.t4 13.9511
R106 VDD2.n3 VDD2.t2 13.9511
R107 VDD2.n1 VDD2.t5 13.9511
R108 VDD2.n1 VDD2.t3 13.9511
R109 VDD2.n0 VDD2.t0 13.9511
R110 VDD2.n0 VDD2.t1 13.9511
R111 VDD2 VDD2.n4 1.54576
R112 VTAIL.n14 VTAIL.t6 168.429
R113 VTAIL.n11 VTAIL.t1 168.429
R114 VTAIL.n10 VTAIL.t13 168.429
R115 VTAIL.n7 VTAIL.t9 168.429
R116 VTAIL.n15 VTAIL.t14 168.429
R117 VTAIL.n2 VTAIL.t15 168.429
R118 VTAIL.n3 VTAIL.t5 168.429
R119 VTAIL.n6 VTAIL.t0 168.429
R120 VTAIL.n13 VTAIL.n12 154.48
R121 VTAIL.n9 VTAIL.n8 154.48
R122 VTAIL.n1 VTAIL.n0 154.48
R123 VTAIL.n5 VTAIL.n4 154.48
R124 VTAIL.n15 VTAIL.n14 17.3496
R125 VTAIL.n7 VTAIL.n6 17.3496
R126 VTAIL.n0 VTAIL.t10 13.9511
R127 VTAIL.n0 VTAIL.t11 13.9511
R128 VTAIL.n4 VTAIL.t4 13.9511
R129 VTAIL.n4 VTAIL.t2 13.9511
R130 VTAIL.n12 VTAIL.t3 13.9511
R131 VTAIL.n12 VTAIL.t7 13.9511
R132 VTAIL.n8 VTAIL.t8 13.9511
R133 VTAIL.n8 VTAIL.t12 13.9511
R134 VTAIL.n9 VTAIL.n7 2.97464
R135 VTAIL.n10 VTAIL.n9 2.97464
R136 VTAIL.n13 VTAIL.n11 2.97464
R137 VTAIL.n14 VTAIL.n13 2.97464
R138 VTAIL.n6 VTAIL.n5 2.97464
R139 VTAIL.n5 VTAIL.n3 2.97464
R140 VTAIL.n2 VTAIL.n1 2.97464
R141 VTAIL VTAIL.n15 2.91645
R142 VTAIL.n11 VTAIL.n10 0.470328
R143 VTAIL.n3 VTAIL.n2 0.470328
R144 VTAIL VTAIL.n1 0.0586897
R145 VP.n21 VP.n18 161.3
R146 VP.n23 VP.n22 161.3
R147 VP.n24 VP.n17 161.3
R148 VP.n26 VP.n25 161.3
R149 VP.n27 VP.n16 161.3
R150 VP.n29 VP.n28 161.3
R151 VP.n31 VP.n30 161.3
R152 VP.n32 VP.n14 161.3
R153 VP.n34 VP.n33 161.3
R154 VP.n35 VP.n13 161.3
R155 VP.n37 VP.n36 161.3
R156 VP.n38 VP.n12 161.3
R157 VP.n40 VP.n39 161.3
R158 VP.n75 VP.n74 161.3
R159 VP.n73 VP.n1 161.3
R160 VP.n72 VP.n71 161.3
R161 VP.n70 VP.n2 161.3
R162 VP.n69 VP.n68 161.3
R163 VP.n67 VP.n3 161.3
R164 VP.n66 VP.n65 161.3
R165 VP.n64 VP.n63 161.3
R166 VP.n62 VP.n5 161.3
R167 VP.n61 VP.n60 161.3
R168 VP.n59 VP.n6 161.3
R169 VP.n58 VP.n57 161.3
R170 VP.n56 VP.n7 161.3
R171 VP.n54 VP.n53 161.3
R172 VP.n52 VP.n8 161.3
R173 VP.n51 VP.n50 161.3
R174 VP.n49 VP.n9 161.3
R175 VP.n48 VP.n47 161.3
R176 VP.n46 VP.n10 161.3
R177 VP.n45 VP.n44 161.3
R178 VP.n43 VP.n42 69.2705
R179 VP.n76 VP.n0 69.2705
R180 VP.n41 VP.n11 69.2705
R181 VP.n49 VP.n48 56.5193
R182 VP.n61 VP.n6 56.5193
R183 VP.n72 VP.n2 56.5193
R184 VP.n37 VP.n13 56.5193
R185 VP.n26 VP.n17 56.5193
R186 VP.n19 VP.t4 51.4112
R187 VP.n20 VP.n19 50.6608
R188 VP.n42 VP.n41 46.166
R189 VP.n44 VP.n10 24.4675
R190 VP.n48 VP.n10 24.4675
R191 VP.n50 VP.n49 24.4675
R192 VP.n50 VP.n8 24.4675
R193 VP.n54 VP.n8 24.4675
R194 VP.n57 VP.n56 24.4675
R195 VP.n57 VP.n6 24.4675
R196 VP.n62 VP.n61 24.4675
R197 VP.n63 VP.n62 24.4675
R198 VP.n67 VP.n66 24.4675
R199 VP.n68 VP.n67 24.4675
R200 VP.n68 VP.n2 24.4675
R201 VP.n73 VP.n72 24.4675
R202 VP.n74 VP.n73 24.4675
R203 VP.n38 VP.n37 24.4675
R204 VP.n39 VP.n38 24.4675
R205 VP.n27 VP.n26 24.4675
R206 VP.n28 VP.n27 24.4675
R207 VP.n32 VP.n31 24.4675
R208 VP.n33 VP.n32 24.4675
R209 VP.n33 VP.n13 24.4675
R210 VP.n22 VP.n21 24.4675
R211 VP.n22 VP.n17 24.4675
R212 VP.n56 VP.n55 23.2442
R213 VP.n63 VP.n4 23.2442
R214 VP.n28 VP.n15 23.2442
R215 VP.n21 VP.n20 23.2442
R216 VP.n44 VP.n43 20.7975
R217 VP.n74 VP.n0 20.7975
R218 VP.n39 VP.n11 20.7975
R219 VP.n43 VP.t0 17.9983
R220 VP.n55 VP.t1 17.9983
R221 VP.n4 VP.t2 17.9983
R222 VP.n0 VP.t7 17.9983
R223 VP.n11 VP.t6 17.9983
R224 VP.n15 VP.t3 17.9983
R225 VP.n20 VP.t5 17.9983
R226 VP.n19 VP.n18 3.87631
R227 VP.n55 VP.n54 1.22385
R228 VP.n66 VP.n4 1.22385
R229 VP.n31 VP.n15 1.22385
R230 VP.n41 VP.n40 0.354971
R231 VP.n45 VP.n42 0.354971
R232 VP.n76 VP.n75 0.354971
R233 VP VP.n76 0.26696
R234 VP.n23 VP.n18 0.189894
R235 VP.n24 VP.n23 0.189894
R236 VP.n25 VP.n24 0.189894
R237 VP.n25 VP.n16 0.189894
R238 VP.n29 VP.n16 0.189894
R239 VP.n30 VP.n29 0.189894
R240 VP.n30 VP.n14 0.189894
R241 VP.n34 VP.n14 0.189894
R242 VP.n35 VP.n34 0.189894
R243 VP.n36 VP.n35 0.189894
R244 VP.n36 VP.n12 0.189894
R245 VP.n40 VP.n12 0.189894
R246 VP.n46 VP.n45 0.189894
R247 VP.n47 VP.n46 0.189894
R248 VP.n47 VP.n9 0.189894
R249 VP.n51 VP.n9 0.189894
R250 VP.n52 VP.n51 0.189894
R251 VP.n53 VP.n52 0.189894
R252 VP.n53 VP.n7 0.189894
R253 VP.n58 VP.n7 0.189894
R254 VP.n59 VP.n58 0.189894
R255 VP.n60 VP.n59 0.189894
R256 VP.n60 VP.n5 0.189894
R257 VP.n64 VP.n5 0.189894
R258 VP.n65 VP.n64 0.189894
R259 VP.n65 VP.n3 0.189894
R260 VP.n69 VP.n3 0.189894
R261 VP.n70 VP.n69 0.189894
R262 VP.n71 VP.n70 0.189894
R263 VP.n71 VP.n1 0.189894
R264 VP.n75 VP.n1 0.189894
R265 VDD1 VDD1.n0 172.703
R266 VDD1.n3 VDD1.n2 172.589
R267 VDD1.n3 VDD1.n1 172.589
R268 VDD1.n5 VDD1.n4 171.159
R269 VDD1.n5 VDD1.n3 39.6905
R270 VDD1.n4 VDD1.t4 13.9511
R271 VDD1.n4 VDD1.t1 13.9511
R272 VDD1.n0 VDD1.t3 13.9511
R273 VDD1.n0 VDD1.t2 13.9511
R274 VDD1.n2 VDD1.t5 13.9511
R275 VDD1.n2 VDD1.t0 13.9511
R276 VDD1.n1 VDD1.t7 13.9511
R277 VDD1.n1 VDD1.t6 13.9511
R278 VDD1 VDD1.n5 1.42938
R279 B.n487 B.n486 585
R280 B.n488 B.n53 585
R281 B.n490 B.n489 585
R282 B.n491 B.n52 585
R283 B.n493 B.n492 585
R284 B.n494 B.n51 585
R285 B.n496 B.n495 585
R286 B.n497 B.n50 585
R287 B.n499 B.n498 585
R288 B.n500 B.n49 585
R289 B.n502 B.n501 585
R290 B.n503 B.n48 585
R291 B.n505 B.n504 585
R292 B.n507 B.n45 585
R293 B.n509 B.n508 585
R294 B.n510 B.n44 585
R295 B.n512 B.n511 585
R296 B.n513 B.n43 585
R297 B.n515 B.n514 585
R298 B.n516 B.n42 585
R299 B.n518 B.n517 585
R300 B.n519 B.n41 585
R301 B.n521 B.n520 585
R302 B.n523 B.n522 585
R303 B.n524 B.n37 585
R304 B.n526 B.n525 585
R305 B.n527 B.n36 585
R306 B.n529 B.n528 585
R307 B.n530 B.n35 585
R308 B.n532 B.n531 585
R309 B.n533 B.n34 585
R310 B.n535 B.n534 585
R311 B.n536 B.n33 585
R312 B.n538 B.n537 585
R313 B.n539 B.n32 585
R314 B.n541 B.n540 585
R315 B.n485 B.n54 585
R316 B.n484 B.n483 585
R317 B.n482 B.n55 585
R318 B.n481 B.n480 585
R319 B.n479 B.n56 585
R320 B.n478 B.n477 585
R321 B.n476 B.n57 585
R322 B.n475 B.n474 585
R323 B.n473 B.n58 585
R324 B.n472 B.n471 585
R325 B.n470 B.n59 585
R326 B.n469 B.n468 585
R327 B.n467 B.n60 585
R328 B.n466 B.n465 585
R329 B.n464 B.n61 585
R330 B.n463 B.n462 585
R331 B.n461 B.n62 585
R332 B.n460 B.n459 585
R333 B.n458 B.n63 585
R334 B.n457 B.n456 585
R335 B.n455 B.n64 585
R336 B.n454 B.n453 585
R337 B.n452 B.n65 585
R338 B.n451 B.n450 585
R339 B.n449 B.n66 585
R340 B.n448 B.n447 585
R341 B.n446 B.n67 585
R342 B.n445 B.n444 585
R343 B.n443 B.n68 585
R344 B.n442 B.n441 585
R345 B.n440 B.n69 585
R346 B.n439 B.n438 585
R347 B.n437 B.n70 585
R348 B.n436 B.n435 585
R349 B.n434 B.n71 585
R350 B.n433 B.n432 585
R351 B.n431 B.n72 585
R352 B.n430 B.n429 585
R353 B.n428 B.n73 585
R354 B.n427 B.n426 585
R355 B.n425 B.n74 585
R356 B.n424 B.n423 585
R357 B.n422 B.n75 585
R358 B.n421 B.n420 585
R359 B.n419 B.n76 585
R360 B.n418 B.n417 585
R361 B.n416 B.n77 585
R362 B.n415 B.n414 585
R363 B.n413 B.n78 585
R364 B.n412 B.n411 585
R365 B.n410 B.n79 585
R366 B.n409 B.n408 585
R367 B.n407 B.n80 585
R368 B.n406 B.n405 585
R369 B.n404 B.n81 585
R370 B.n403 B.n402 585
R371 B.n401 B.n82 585
R372 B.n400 B.n399 585
R373 B.n398 B.n83 585
R374 B.n397 B.n396 585
R375 B.n395 B.n84 585
R376 B.n394 B.n393 585
R377 B.n392 B.n85 585
R378 B.n391 B.n390 585
R379 B.n389 B.n86 585
R380 B.n388 B.n387 585
R381 B.n386 B.n87 585
R382 B.n385 B.n384 585
R383 B.n383 B.n88 585
R384 B.n382 B.n381 585
R385 B.n380 B.n89 585
R386 B.n379 B.n378 585
R387 B.n377 B.n90 585
R388 B.n376 B.n375 585
R389 B.n374 B.n91 585
R390 B.n373 B.n372 585
R391 B.n371 B.n92 585
R392 B.n370 B.n369 585
R393 B.n368 B.n93 585
R394 B.n367 B.n366 585
R395 B.n365 B.n94 585
R396 B.n364 B.n363 585
R397 B.n362 B.n95 585
R398 B.n361 B.n360 585
R399 B.n359 B.n96 585
R400 B.n358 B.n357 585
R401 B.n356 B.n97 585
R402 B.n355 B.n354 585
R403 B.n353 B.n98 585
R404 B.n352 B.n351 585
R405 B.n350 B.n99 585
R406 B.n349 B.n348 585
R407 B.n347 B.n100 585
R408 B.n346 B.n345 585
R409 B.n344 B.n101 585
R410 B.n343 B.n342 585
R411 B.n341 B.n102 585
R412 B.n340 B.n339 585
R413 B.n338 B.n103 585
R414 B.n337 B.n336 585
R415 B.n335 B.n104 585
R416 B.n334 B.n333 585
R417 B.n332 B.n105 585
R418 B.n331 B.n330 585
R419 B.n329 B.n106 585
R420 B.n328 B.n327 585
R421 B.n326 B.n107 585
R422 B.n325 B.n324 585
R423 B.n323 B.n108 585
R424 B.n322 B.n321 585
R425 B.n320 B.n109 585
R426 B.n319 B.n318 585
R427 B.n317 B.n110 585
R428 B.n316 B.n315 585
R429 B.n314 B.n111 585
R430 B.n313 B.n312 585
R431 B.n311 B.n112 585
R432 B.n310 B.n309 585
R433 B.n308 B.n113 585
R434 B.n253 B.n252 585
R435 B.n254 B.n135 585
R436 B.n256 B.n255 585
R437 B.n257 B.n134 585
R438 B.n259 B.n258 585
R439 B.n260 B.n133 585
R440 B.n262 B.n261 585
R441 B.n263 B.n132 585
R442 B.n265 B.n264 585
R443 B.n266 B.n131 585
R444 B.n268 B.n267 585
R445 B.n269 B.n130 585
R446 B.n271 B.n270 585
R447 B.n273 B.n127 585
R448 B.n275 B.n274 585
R449 B.n276 B.n126 585
R450 B.n278 B.n277 585
R451 B.n279 B.n125 585
R452 B.n281 B.n280 585
R453 B.n282 B.n124 585
R454 B.n284 B.n283 585
R455 B.n285 B.n123 585
R456 B.n287 B.n286 585
R457 B.n289 B.n288 585
R458 B.n290 B.n119 585
R459 B.n292 B.n291 585
R460 B.n293 B.n118 585
R461 B.n295 B.n294 585
R462 B.n296 B.n117 585
R463 B.n298 B.n297 585
R464 B.n299 B.n116 585
R465 B.n301 B.n300 585
R466 B.n302 B.n115 585
R467 B.n304 B.n303 585
R468 B.n305 B.n114 585
R469 B.n307 B.n306 585
R470 B.n251 B.n136 585
R471 B.n250 B.n249 585
R472 B.n248 B.n137 585
R473 B.n247 B.n246 585
R474 B.n245 B.n138 585
R475 B.n244 B.n243 585
R476 B.n242 B.n139 585
R477 B.n241 B.n240 585
R478 B.n239 B.n140 585
R479 B.n238 B.n237 585
R480 B.n236 B.n141 585
R481 B.n235 B.n234 585
R482 B.n233 B.n142 585
R483 B.n232 B.n231 585
R484 B.n230 B.n143 585
R485 B.n229 B.n228 585
R486 B.n227 B.n144 585
R487 B.n226 B.n225 585
R488 B.n224 B.n145 585
R489 B.n223 B.n222 585
R490 B.n221 B.n146 585
R491 B.n220 B.n219 585
R492 B.n218 B.n147 585
R493 B.n217 B.n216 585
R494 B.n215 B.n148 585
R495 B.n214 B.n213 585
R496 B.n212 B.n149 585
R497 B.n211 B.n210 585
R498 B.n209 B.n150 585
R499 B.n208 B.n207 585
R500 B.n206 B.n151 585
R501 B.n205 B.n204 585
R502 B.n203 B.n152 585
R503 B.n202 B.n201 585
R504 B.n200 B.n153 585
R505 B.n199 B.n198 585
R506 B.n197 B.n154 585
R507 B.n196 B.n195 585
R508 B.n194 B.n155 585
R509 B.n193 B.n192 585
R510 B.n191 B.n156 585
R511 B.n190 B.n189 585
R512 B.n188 B.n157 585
R513 B.n187 B.n186 585
R514 B.n185 B.n158 585
R515 B.n184 B.n183 585
R516 B.n182 B.n159 585
R517 B.n181 B.n180 585
R518 B.n179 B.n160 585
R519 B.n178 B.n177 585
R520 B.n176 B.n161 585
R521 B.n175 B.n174 585
R522 B.n173 B.n162 585
R523 B.n172 B.n171 585
R524 B.n170 B.n163 585
R525 B.n169 B.n168 585
R526 B.n167 B.n164 585
R527 B.n166 B.n165 585
R528 B.n2 B.n0 585
R529 B.n629 B.n1 585
R530 B.n628 B.n627 585
R531 B.n626 B.n3 585
R532 B.n625 B.n624 585
R533 B.n623 B.n4 585
R534 B.n622 B.n621 585
R535 B.n620 B.n5 585
R536 B.n619 B.n618 585
R537 B.n617 B.n6 585
R538 B.n616 B.n615 585
R539 B.n614 B.n7 585
R540 B.n613 B.n612 585
R541 B.n611 B.n8 585
R542 B.n610 B.n609 585
R543 B.n608 B.n9 585
R544 B.n607 B.n606 585
R545 B.n605 B.n10 585
R546 B.n604 B.n603 585
R547 B.n602 B.n11 585
R548 B.n601 B.n600 585
R549 B.n599 B.n12 585
R550 B.n598 B.n597 585
R551 B.n596 B.n13 585
R552 B.n595 B.n594 585
R553 B.n593 B.n14 585
R554 B.n592 B.n591 585
R555 B.n590 B.n15 585
R556 B.n589 B.n588 585
R557 B.n587 B.n16 585
R558 B.n586 B.n585 585
R559 B.n584 B.n17 585
R560 B.n583 B.n582 585
R561 B.n581 B.n18 585
R562 B.n580 B.n579 585
R563 B.n578 B.n19 585
R564 B.n577 B.n576 585
R565 B.n575 B.n20 585
R566 B.n574 B.n573 585
R567 B.n572 B.n21 585
R568 B.n571 B.n570 585
R569 B.n569 B.n22 585
R570 B.n568 B.n567 585
R571 B.n566 B.n23 585
R572 B.n565 B.n564 585
R573 B.n563 B.n24 585
R574 B.n562 B.n561 585
R575 B.n560 B.n25 585
R576 B.n559 B.n558 585
R577 B.n557 B.n26 585
R578 B.n556 B.n555 585
R579 B.n554 B.n27 585
R580 B.n553 B.n552 585
R581 B.n551 B.n28 585
R582 B.n550 B.n549 585
R583 B.n548 B.n29 585
R584 B.n547 B.n546 585
R585 B.n545 B.n30 585
R586 B.n544 B.n543 585
R587 B.n542 B.n31 585
R588 B.n631 B.n630 585
R589 B.n252 B.n251 468.476
R590 B.n540 B.n31 468.476
R591 B.n306 B.n113 468.476
R592 B.n486 B.n485 468.476
R593 B.n120 B.t5 241.454
R594 B.n46 B.t1 241.454
R595 B.n128 B.t11 241.453
R596 B.n38 B.t7 241.453
R597 B.n120 B.t3 226.714
R598 B.n128 B.t9 226.714
R599 B.n38 B.t6 226.714
R600 B.n46 B.t0 226.714
R601 B.n121 B.t4 174.544
R602 B.n47 B.t2 174.544
R603 B.n129 B.t10 174.544
R604 B.n39 B.t8 174.544
R605 B.n251 B.n250 163.367
R606 B.n250 B.n137 163.367
R607 B.n246 B.n137 163.367
R608 B.n246 B.n245 163.367
R609 B.n245 B.n244 163.367
R610 B.n244 B.n139 163.367
R611 B.n240 B.n139 163.367
R612 B.n240 B.n239 163.367
R613 B.n239 B.n238 163.367
R614 B.n238 B.n141 163.367
R615 B.n234 B.n141 163.367
R616 B.n234 B.n233 163.367
R617 B.n233 B.n232 163.367
R618 B.n232 B.n143 163.367
R619 B.n228 B.n143 163.367
R620 B.n228 B.n227 163.367
R621 B.n227 B.n226 163.367
R622 B.n226 B.n145 163.367
R623 B.n222 B.n145 163.367
R624 B.n222 B.n221 163.367
R625 B.n221 B.n220 163.367
R626 B.n220 B.n147 163.367
R627 B.n216 B.n147 163.367
R628 B.n216 B.n215 163.367
R629 B.n215 B.n214 163.367
R630 B.n214 B.n149 163.367
R631 B.n210 B.n149 163.367
R632 B.n210 B.n209 163.367
R633 B.n209 B.n208 163.367
R634 B.n208 B.n151 163.367
R635 B.n204 B.n151 163.367
R636 B.n204 B.n203 163.367
R637 B.n203 B.n202 163.367
R638 B.n202 B.n153 163.367
R639 B.n198 B.n153 163.367
R640 B.n198 B.n197 163.367
R641 B.n197 B.n196 163.367
R642 B.n196 B.n155 163.367
R643 B.n192 B.n155 163.367
R644 B.n192 B.n191 163.367
R645 B.n191 B.n190 163.367
R646 B.n190 B.n157 163.367
R647 B.n186 B.n157 163.367
R648 B.n186 B.n185 163.367
R649 B.n185 B.n184 163.367
R650 B.n184 B.n159 163.367
R651 B.n180 B.n159 163.367
R652 B.n180 B.n179 163.367
R653 B.n179 B.n178 163.367
R654 B.n178 B.n161 163.367
R655 B.n174 B.n161 163.367
R656 B.n174 B.n173 163.367
R657 B.n173 B.n172 163.367
R658 B.n172 B.n163 163.367
R659 B.n168 B.n163 163.367
R660 B.n168 B.n167 163.367
R661 B.n167 B.n166 163.367
R662 B.n166 B.n2 163.367
R663 B.n630 B.n2 163.367
R664 B.n630 B.n629 163.367
R665 B.n629 B.n628 163.367
R666 B.n628 B.n3 163.367
R667 B.n624 B.n3 163.367
R668 B.n624 B.n623 163.367
R669 B.n623 B.n622 163.367
R670 B.n622 B.n5 163.367
R671 B.n618 B.n5 163.367
R672 B.n618 B.n617 163.367
R673 B.n617 B.n616 163.367
R674 B.n616 B.n7 163.367
R675 B.n612 B.n7 163.367
R676 B.n612 B.n611 163.367
R677 B.n611 B.n610 163.367
R678 B.n610 B.n9 163.367
R679 B.n606 B.n9 163.367
R680 B.n606 B.n605 163.367
R681 B.n605 B.n604 163.367
R682 B.n604 B.n11 163.367
R683 B.n600 B.n11 163.367
R684 B.n600 B.n599 163.367
R685 B.n599 B.n598 163.367
R686 B.n598 B.n13 163.367
R687 B.n594 B.n13 163.367
R688 B.n594 B.n593 163.367
R689 B.n593 B.n592 163.367
R690 B.n592 B.n15 163.367
R691 B.n588 B.n15 163.367
R692 B.n588 B.n587 163.367
R693 B.n587 B.n586 163.367
R694 B.n586 B.n17 163.367
R695 B.n582 B.n17 163.367
R696 B.n582 B.n581 163.367
R697 B.n581 B.n580 163.367
R698 B.n580 B.n19 163.367
R699 B.n576 B.n19 163.367
R700 B.n576 B.n575 163.367
R701 B.n575 B.n574 163.367
R702 B.n574 B.n21 163.367
R703 B.n570 B.n21 163.367
R704 B.n570 B.n569 163.367
R705 B.n569 B.n568 163.367
R706 B.n568 B.n23 163.367
R707 B.n564 B.n23 163.367
R708 B.n564 B.n563 163.367
R709 B.n563 B.n562 163.367
R710 B.n562 B.n25 163.367
R711 B.n558 B.n25 163.367
R712 B.n558 B.n557 163.367
R713 B.n557 B.n556 163.367
R714 B.n556 B.n27 163.367
R715 B.n552 B.n27 163.367
R716 B.n552 B.n551 163.367
R717 B.n551 B.n550 163.367
R718 B.n550 B.n29 163.367
R719 B.n546 B.n29 163.367
R720 B.n546 B.n545 163.367
R721 B.n545 B.n544 163.367
R722 B.n544 B.n31 163.367
R723 B.n252 B.n135 163.367
R724 B.n256 B.n135 163.367
R725 B.n257 B.n256 163.367
R726 B.n258 B.n257 163.367
R727 B.n258 B.n133 163.367
R728 B.n262 B.n133 163.367
R729 B.n263 B.n262 163.367
R730 B.n264 B.n263 163.367
R731 B.n264 B.n131 163.367
R732 B.n268 B.n131 163.367
R733 B.n269 B.n268 163.367
R734 B.n270 B.n269 163.367
R735 B.n270 B.n127 163.367
R736 B.n275 B.n127 163.367
R737 B.n276 B.n275 163.367
R738 B.n277 B.n276 163.367
R739 B.n277 B.n125 163.367
R740 B.n281 B.n125 163.367
R741 B.n282 B.n281 163.367
R742 B.n283 B.n282 163.367
R743 B.n283 B.n123 163.367
R744 B.n287 B.n123 163.367
R745 B.n288 B.n287 163.367
R746 B.n288 B.n119 163.367
R747 B.n292 B.n119 163.367
R748 B.n293 B.n292 163.367
R749 B.n294 B.n293 163.367
R750 B.n294 B.n117 163.367
R751 B.n298 B.n117 163.367
R752 B.n299 B.n298 163.367
R753 B.n300 B.n299 163.367
R754 B.n300 B.n115 163.367
R755 B.n304 B.n115 163.367
R756 B.n305 B.n304 163.367
R757 B.n306 B.n305 163.367
R758 B.n310 B.n113 163.367
R759 B.n311 B.n310 163.367
R760 B.n312 B.n311 163.367
R761 B.n312 B.n111 163.367
R762 B.n316 B.n111 163.367
R763 B.n317 B.n316 163.367
R764 B.n318 B.n317 163.367
R765 B.n318 B.n109 163.367
R766 B.n322 B.n109 163.367
R767 B.n323 B.n322 163.367
R768 B.n324 B.n323 163.367
R769 B.n324 B.n107 163.367
R770 B.n328 B.n107 163.367
R771 B.n329 B.n328 163.367
R772 B.n330 B.n329 163.367
R773 B.n330 B.n105 163.367
R774 B.n334 B.n105 163.367
R775 B.n335 B.n334 163.367
R776 B.n336 B.n335 163.367
R777 B.n336 B.n103 163.367
R778 B.n340 B.n103 163.367
R779 B.n341 B.n340 163.367
R780 B.n342 B.n341 163.367
R781 B.n342 B.n101 163.367
R782 B.n346 B.n101 163.367
R783 B.n347 B.n346 163.367
R784 B.n348 B.n347 163.367
R785 B.n348 B.n99 163.367
R786 B.n352 B.n99 163.367
R787 B.n353 B.n352 163.367
R788 B.n354 B.n353 163.367
R789 B.n354 B.n97 163.367
R790 B.n358 B.n97 163.367
R791 B.n359 B.n358 163.367
R792 B.n360 B.n359 163.367
R793 B.n360 B.n95 163.367
R794 B.n364 B.n95 163.367
R795 B.n365 B.n364 163.367
R796 B.n366 B.n365 163.367
R797 B.n366 B.n93 163.367
R798 B.n370 B.n93 163.367
R799 B.n371 B.n370 163.367
R800 B.n372 B.n371 163.367
R801 B.n372 B.n91 163.367
R802 B.n376 B.n91 163.367
R803 B.n377 B.n376 163.367
R804 B.n378 B.n377 163.367
R805 B.n378 B.n89 163.367
R806 B.n382 B.n89 163.367
R807 B.n383 B.n382 163.367
R808 B.n384 B.n383 163.367
R809 B.n384 B.n87 163.367
R810 B.n388 B.n87 163.367
R811 B.n389 B.n388 163.367
R812 B.n390 B.n389 163.367
R813 B.n390 B.n85 163.367
R814 B.n394 B.n85 163.367
R815 B.n395 B.n394 163.367
R816 B.n396 B.n395 163.367
R817 B.n396 B.n83 163.367
R818 B.n400 B.n83 163.367
R819 B.n401 B.n400 163.367
R820 B.n402 B.n401 163.367
R821 B.n402 B.n81 163.367
R822 B.n406 B.n81 163.367
R823 B.n407 B.n406 163.367
R824 B.n408 B.n407 163.367
R825 B.n408 B.n79 163.367
R826 B.n412 B.n79 163.367
R827 B.n413 B.n412 163.367
R828 B.n414 B.n413 163.367
R829 B.n414 B.n77 163.367
R830 B.n418 B.n77 163.367
R831 B.n419 B.n418 163.367
R832 B.n420 B.n419 163.367
R833 B.n420 B.n75 163.367
R834 B.n424 B.n75 163.367
R835 B.n425 B.n424 163.367
R836 B.n426 B.n425 163.367
R837 B.n426 B.n73 163.367
R838 B.n430 B.n73 163.367
R839 B.n431 B.n430 163.367
R840 B.n432 B.n431 163.367
R841 B.n432 B.n71 163.367
R842 B.n436 B.n71 163.367
R843 B.n437 B.n436 163.367
R844 B.n438 B.n437 163.367
R845 B.n438 B.n69 163.367
R846 B.n442 B.n69 163.367
R847 B.n443 B.n442 163.367
R848 B.n444 B.n443 163.367
R849 B.n444 B.n67 163.367
R850 B.n448 B.n67 163.367
R851 B.n449 B.n448 163.367
R852 B.n450 B.n449 163.367
R853 B.n450 B.n65 163.367
R854 B.n454 B.n65 163.367
R855 B.n455 B.n454 163.367
R856 B.n456 B.n455 163.367
R857 B.n456 B.n63 163.367
R858 B.n460 B.n63 163.367
R859 B.n461 B.n460 163.367
R860 B.n462 B.n461 163.367
R861 B.n462 B.n61 163.367
R862 B.n466 B.n61 163.367
R863 B.n467 B.n466 163.367
R864 B.n468 B.n467 163.367
R865 B.n468 B.n59 163.367
R866 B.n472 B.n59 163.367
R867 B.n473 B.n472 163.367
R868 B.n474 B.n473 163.367
R869 B.n474 B.n57 163.367
R870 B.n478 B.n57 163.367
R871 B.n479 B.n478 163.367
R872 B.n480 B.n479 163.367
R873 B.n480 B.n55 163.367
R874 B.n484 B.n55 163.367
R875 B.n485 B.n484 163.367
R876 B.n540 B.n539 163.367
R877 B.n539 B.n538 163.367
R878 B.n538 B.n33 163.367
R879 B.n534 B.n33 163.367
R880 B.n534 B.n533 163.367
R881 B.n533 B.n532 163.367
R882 B.n532 B.n35 163.367
R883 B.n528 B.n35 163.367
R884 B.n528 B.n527 163.367
R885 B.n527 B.n526 163.367
R886 B.n526 B.n37 163.367
R887 B.n522 B.n37 163.367
R888 B.n522 B.n521 163.367
R889 B.n521 B.n41 163.367
R890 B.n517 B.n41 163.367
R891 B.n517 B.n516 163.367
R892 B.n516 B.n515 163.367
R893 B.n515 B.n43 163.367
R894 B.n511 B.n43 163.367
R895 B.n511 B.n510 163.367
R896 B.n510 B.n509 163.367
R897 B.n509 B.n45 163.367
R898 B.n504 B.n45 163.367
R899 B.n504 B.n503 163.367
R900 B.n503 B.n502 163.367
R901 B.n502 B.n49 163.367
R902 B.n498 B.n49 163.367
R903 B.n498 B.n497 163.367
R904 B.n497 B.n496 163.367
R905 B.n496 B.n51 163.367
R906 B.n492 B.n51 163.367
R907 B.n492 B.n491 163.367
R908 B.n491 B.n490 163.367
R909 B.n490 B.n53 163.367
R910 B.n486 B.n53 163.367
R911 B.n121 B.n120 66.9096
R912 B.n129 B.n128 66.9096
R913 B.n39 B.n38 66.9096
R914 B.n47 B.n46 66.9096
R915 B.n122 B.n121 59.5399
R916 B.n272 B.n129 59.5399
R917 B.n40 B.n39 59.5399
R918 B.n506 B.n47 59.5399
R919 B.n542 B.n541 30.4395
R920 B.n487 B.n54 30.4395
R921 B.n308 B.n307 30.4395
R922 B.n253 B.n136 30.4395
R923 B B.n631 18.0485
R924 B.n541 B.n32 10.6151
R925 B.n537 B.n32 10.6151
R926 B.n537 B.n536 10.6151
R927 B.n536 B.n535 10.6151
R928 B.n535 B.n34 10.6151
R929 B.n531 B.n34 10.6151
R930 B.n531 B.n530 10.6151
R931 B.n530 B.n529 10.6151
R932 B.n529 B.n36 10.6151
R933 B.n525 B.n36 10.6151
R934 B.n525 B.n524 10.6151
R935 B.n524 B.n523 10.6151
R936 B.n520 B.n519 10.6151
R937 B.n519 B.n518 10.6151
R938 B.n518 B.n42 10.6151
R939 B.n514 B.n42 10.6151
R940 B.n514 B.n513 10.6151
R941 B.n513 B.n512 10.6151
R942 B.n512 B.n44 10.6151
R943 B.n508 B.n44 10.6151
R944 B.n508 B.n507 10.6151
R945 B.n505 B.n48 10.6151
R946 B.n501 B.n48 10.6151
R947 B.n501 B.n500 10.6151
R948 B.n500 B.n499 10.6151
R949 B.n499 B.n50 10.6151
R950 B.n495 B.n50 10.6151
R951 B.n495 B.n494 10.6151
R952 B.n494 B.n493 10.6151
R953 B.n493 B.n52 10.6151
R954 B.n489 B.n52 10.6151
R955 B.n489 B.n488 10.6151
R956 B.n488 B.n487 10.6151
R957 B.n309 B.n308 10.6151
R958 B.n309 B.n112 10.6151
R959 B.n313 B.n112 10.6151
R960 B.n314 B.n313 10.6151
R961 B.n315 B.n314 10.6151
R962 B.n315 B.n110 10.6151
R963 B.n319 B.n110 10.6151
R964 B.n320 B.n319 10.6151
R965 B.n321 B.n320 10.6151
R966 B.n321 B.n108 10.6151
R967 B.n325 B.n108 10.6151
R968 B.n326 B.n325 10.6151
R969 B.n327 B.n326 10.6151
R970 B.n327 B.n106 10.6151
R971 B.n331 B.n106 10.6151
R972 B.n332 B.n331 10.6151
R973 B.n333 B.n332 10.6151
R974 B.n333 B.n104 10.6151
R975 B.n337 B.n104 10.6151
R976 B.n338 B.n337 10.6151
R977 B.n339 B.n338 10.6151
R978 B.n339 B.n102 10.6151
R979 B.n343 B.n102 10.6151
R980 B.n344 B.n343 10.6151
R981 B.n345 B.n344 10.6151
R982 B.n345 B.n100 10.6151
R983 B.n349 B.n100 10.6151
R984 B.n350 B.n349 10.6151
R985 B.n351 B.n350 10.6151
R986 B.n351 B.n98 10.6151
R987 B.n355 B.n98 10.6151
R988 B.n356 B.n355 10.6151
R989 B.n357 B.n356 10.6151
R990 B.n357 B.n96 10.6151
R991 B.n361 B.n96 10.6151
R992 B.n362 B.n361 10.6151
R993 B.n363 B.n362 10.6151
R994 B.n363 B.n94 10.6151
R995 B.n367 B.n94 10.6151
R996 B.n368 B.n367 10.6151
R997 B.n369 B.n368 10.6151
R998 B.n369 B.n92 10.6151
R999 B.n373 B.n92 10.6151
R1000 B.n374 B.n373 10.6151
R1001 B.n375 B.n374 10.6151
R1002 B.n375 B.n90 10.6151
R1003 B.n379 B.n90 10.6151
R1004 B.n380 B.n379 10.6151
R1005 B.n381 B.n380 10.6151
R1006 B.n381 B.n88 10.6151
R1007 B.n385 B.n88 10.6151
R1008 B.n386 B.n385 10.6151
R1009 B.n387 B.n386 10.6151
R1010 B.n387 B.n86 10.6151
R1011 B.n391 B.n86 10.6151
R1012 B.n392 B.n391 10.6151
R1013 B.n393 B.n392 10.6151
R1014 B.n393 B.n84 10.6151
R1015 B.n397 B.n84 10.6151
R1016 B.n398 B.n397 10.6151
R1017 B.n399 B.n398 10.6151
R1018 B.n399 B.n82 10.6151
R1019 B.n403 B.n82 10.6151
R1020 B.n404 B.n403 10.6151
R1021 B.n405 B.n404 10.6151
R1022 B.n405 B.n80 10.6151
R1023 B.n409 B.n80 10.6151
R1024 B.n410 B.n409 10.6151
R1025 B.n411 B.n410 10.6151
R1026 B.n411 B.n78 10.6151
R1027 B.n415 B.n78 10.6151
R1028 B.n416 B.n415 10.6151
R1029 B.n417 B.n416 10.6151
R1030 B.n417 B.n76 10.6151
R1031 B.n421 B.n76 10.6151
R1032 B.n422 B.n421 10.6151
R1033 B.n423 B.n422 10.6151
R1034 B.n423 B.n74 10.6151
R1035 B.n427 B.n74 10.6151
R1036 B.n428 B.n427 10.6151
R1037 B.n429 B.n428 10.6151
R1038 B.n429 B.n72 10.6151
R1039 B.n433 B.n72 10.6151
R1040 B.n434 B.n433 10.6151
R1041 B.n435 B.n434 10.6151
R1042 B.n435 B.n70 10.6151
R1043 B.n439 B.n70 10.6151
R1044 B.n440 B.n439 10.6151
R1045 B.n441 B.n440 10.6151
R1046 B.n441 B.n68 10.6151
R1047 B.n445 B.n68 10.6151
R1048 B.n446 B.n445 10.6151
R1049 B.n447 B.n446 10.6151
R1050 B.n447 B.n66 10.6151
R1051 B.n451 B.n66 10.6151
R1052 B.n452 B.n451 10.6151
R1053 B.n453 B.n452 10.6151
R1054 B.n453 B.n64 10.6151
R1055 B.n457 B.n64 10.6151
R1056 B.n458 B.n457 10.6151
R1057 B.n459 B.n458 10.6151
R1058 B.n459 B.n62 10.6151
R1059 B.n463 B.n62 10.6151
R1060 B.n464 B.n463 10.6151
R1061 B.n465 B.n464 10.6151
R1062 B.n465 B.n60 10.6151
R1063 B.n469 B.n60 10.6151
R1064 B.n470 B.n469 10.6151
R1065 B.n471 B.n470 10.6151
R1066 B.n471 B.n58 10.6151
R1067 B.n475 B.n58 10.6151
R1068 B.n476 B.n475 10.6151
R1069 B.n477 B.n476 10.6151
R1070 B.n477 B.n56 10.6151
R1071 B.n481 B.n56 10.6151
R1072 B.n482 B.n481 10.6151
R1073 B.n483 B.n482 10.6151
R1074 B.n483 B.n54 10.6151
R1075 B.n254 B.n253 10.6151
R1076 B.n255 B.n254 10.6151
R1077 B.n255 B.n134 10.6151
R1078 B.n259 B.n134 10.6151
R1079 B.n260 B.n259 10.6151
R1080 B.n261 B.n260 10.6151
R1081 B.n261 B.n132 10.6151
R1082 B.n265 B.n132 10.6151
R1083 B.n266 B.n265 10.6151
R1084 B.n267 B.n266 10.6151
R1085 B.n267 B.n130 10.6151
R1086 B.n271 B.n130 10.6151
R1087 B.n274 B.n273 10.6151
R1088 B.n274 B.n126 10.6151
R1089 B.n278 B.n126 10.6151
R1090 B.n279 B.n278 10.6151
R1091 B.n280 B.n279 10.6151
R1092 B.n280 B.n124 10.6151
R1093 B.n284 B.n124 10.6151
R1094 B.n285 B.n284 10.6151
R1095 B.n286 B.n285 10.6151
R1096 B.n290 B.n289 10.6151
R1097 B.n291 B.n290 10.6151
R1098 B.n291 B.n118 10.6151
R1099 B.n295 B.n118 10.6151
R1100 B.n296 B.n295 10.6151
R1101 B.n297 B.n296 10.6151
R1102 B.n297 B.n116 10.6151
R1103 B.n301 B.n116 10.6151
R1104 B.n302 B.n301 10.6151
R1105 B.n303 B.n302 10.6151
R1106 B.n303 B.n114 10.6151
R1107 B.n307 B.n114 10.6151
R1108 B.n249 B.n136 10.6151
R1109 B.n249 B.n248 10.6151
R1110 B.n248 B.n247 10.6151
R1111 B.n247 B.n138 10.6151
R1112 B.n243 B.n138 10.6151
R1113 B.n243 B.n242 10.6151
R1114 B.n242 B.n241 10.6151
R1115 B.n241 B.n140 10.6151
R1116 B.n237 B.n140 10.6151
R1117 B.n237 B.n236 10.6151
R1118 B.n236 B.n235 10.6151
R1119 B.n235 B.n142 10.6151
R1120 B.n231 B.n142 10.6151
R1121 B.n231 B.n230 10.6151
R1122 B.n230 B.n229 10.6151
R1123 B.n229 B.n144 10.6151
R1124 B.n225 B.n144 10.6151
R1125 B.n225 B.n224 10.6151
R1126 B.n224 B.n223 10.6151
R1127 B.n223 B.n146 10.6151
R1128 B.n219 B.n146 10.6151
R1129 B.n219 B.n218 10.6151
R1130 B.n218 B.n217 10.6151
R1131 B.n217 B.n148 10.6151
R1132 B.n213 B.n148 10.6151
R1133 B.n213 B.n212 10.6151
R1134 B.n212 B.n211 10.6151
R1135 B.n211 B.n150 10.6151
R1136 B.n207 B.n150 10.6151
R1137 B.n207 B.n206 10.6151
R1138 B.n206 B.n205 10.6151
R1139 B.n205 B.n152 10.6151
R1140 B.n201 B.n152 10.6151
R1141 B.n201 B.n200 10.6151
R1142 B.n200 B.n199 10.6151
R1143 B.n199 B.n154 10.6151
R1144 B.n195 B.n154 10.6151
R1145 B.n195 B.n194 10.6151
R1146 B.n194 B.n193 10.6151
R1147 B.n193 B.n156 10.6151
R1148 B.n189 B.n156 10.6151
R1149 B.n189 B.n188 10.6151
R1150 B.n188 B.n187 10.6151
R1151 B.n187 B.n158 10.6151
R1152 B.n183 B.n158 10.6151
R1153 B.n183 B.n182 10.6151
R1154 B.n182 B.n181 10.6151
R1155 B.n181 B.n160 10.6151
R1156 B.n177 B.n160 10.6151
R1157 B.n177 B.n176 10.6151
R1158 B.n176 B.n175 10.6151
R1159 B.n175 B.n162 10.6151
R1160 B.n171 B.n162 10.6151
R1161 B.n171 B.n170 10.6151
R1162 B.n170 B.n169 10.6151
R1163 B.n169 B.n164 10.6151
R1164 B.n165 B.n164 10.6151
R1165 B.n165 B.n0 10.6151
R1166 B.n627 B.n1 10.6151
R1167 B.n627 B.n626 10.6151
R1168 B.n626 B.n625 10.6151
R1169 B.n625 B.n4 10.6151
R1170 B.n621 B.n4 10.6151
R1171 B.n621 B.n620 10.6151
R1172 B.n620 B.n619 10.6151
R1173 B.n619 B.n6 10.6151
R1174 B.n615 B.n6 10.6151
R1175 B.n615 B.n614 10.6151
R1176 B.n614 B.n613 10.6151
R1177 B.n613 B.n8 10.6151
R1178 B.n609 B.n8 10.6151
R1179 B.n609 B.n608 10.6151
R1180 B.n608 B.n607 10.6151
R1181 B.n607 B.n10 10.6151
R1182 B.n603 B.n10 10.6151
R1183 B.n603 B.n602 10.6151
R1184 B.n602 B.n601 10.6151
R1185 B.n601 B.n12 10.6151
R1186 B.n597 B.n12 10.6151
R1187 B.n597 B.n596 10.6151
R1188 B.n596 B.n595 10.6151
R1189 B.n595 B.n14 10.6151
R1190 B.n591 B.n14 10.6151
R1191 B.n591 B.n590 10.6151
R1192 B.n590 B.n589 10.6151
R1193 B.n589 B.n16 10.6151
R1194 B.n585 B.n16 10.6151
R1195 B.n585 B.n584 10.6151
R1196 B.n584 B.n583 10.6151
R1197 B.n583 B.n18 10.6151
R1198 B.n579 B.n18 10.6151
R1199 B.n579 B.n578 10.6151
R1200 B.n578 B.n577 10.6151
R1201 B.n577 B.n20 10.6151
R1202 B.n573 B.n20 10.6151
R1203 B.n573 B.n572 10.6151
R1204 B.n572 B.n571 10.6151
R1205 B.n571 B.n22 10.6151
R1206 B.n567 B.n22 10.6151
R1207 B.n567 B.n566 10.6151
R1208 B.n566 B.n565 10.6151
R1209 B.n565 B.n24 10.6151
R1210 B.n561 B.n24 10.6151
R1211 B.n561 B.n560 10.6151
R1212 B.n560 B.n559 10.6151
R1213 B.n559 B.n26 10.6151
R1214 B.n555 B.n26 10.6151
R1215 B.n555 B.n554 10.6151
R1216 B.n554 B.n553 10.6151
R1217 B.n553 B.n28 10.6151
R1218 B.n549 B.n28 10.6151
R1219 B.n549 B.n548 10.6151
R1220 B.n548 B.n547 10.6151
R1221 B.n547 B.n30 10.6151
R1222 B.n543 B.n30 10.6151
R1223 B.n543 B.n542 10.6151
R1224 B.n523 B.n40 9.36635
R1225 B.n506 B.n505 9.36635
R1226 B.n272 B.n271 9.36635
R1227 B.n289 B.n122 9.36635
R1228 B.n631 B.n0 2.81026
R1229 B.n631 B.n1 2.81026
R1230 B.n520 B.n40 1.24928
R1231 B.n507 B.n506 1.24928
R1232 B.n273 B.n272 1.24928
R1233 B.n286 B.n122 1.24928
C0 VP w_n4420_n1434# 9.54649f
C1 VTAIL B 1.84989f
C2 VDD2 VN 2.11811f
C3 VDD1 VN 0.158294f
C4 VTAIL VP 3.45631f
C5 VDD2 w_n4420_n1434# 1.99735f
C6 VP B 2.20758f
C7 VDD1 w_n4420_n1434# 1.86149f
C8 VDD2 VTAIL 5.34477f
C9 VDD1 VTAIL 5.28686f
C10 VDD2 B 1.65912f
C11 VDD1 B 1.54637f
C12 VN w_n4420_n1434# 8.97471f
C13 VDD2 VP 0.581781f
C14 VDD1 VP 2.53849f
C15 VTAIL VN 3.44221f
C16 VN B 1.24096f
C17 VTAIL w_n4420_n1434# 2.07908f
C18 B w_n4420_n1434# 8.25456f
C19 VDD2 VDD1 2.04916f
C20 VP VN 6.5148f
C21 VDD2 VSUBS 1.740192f
C22 VDD1 VSUBS 2.50668f
C23 VTAIL VSUBS 0.634607f
C24 VN VSUBS 7.546821f
C25 VP VSUBS 3.514808f
C26 B VSUBS 4.473215f
C27 w_n4420_n1434# VSUBS 80.6738f
C28 B.n0 VSUBS 0.006619f
C29 B.n1 VSUBS 0.006619f
C30 B.n2 VSUBS 0.010468f
C31 B.n3 VSUBS 0.010468f
C32 B.n4 VSUBS 0.010468f
C33 B.n5 VSUBS 0.010468f
C34 B.n6 VSUBS 0.010468f
C35 B.n7 VSUBS 0.010468f
C36 B.n8 VSUBS 0.010468f
C37 B.n9 VSUBS 0.010468f
C38 B.n10 VSUBS 0.010468f
C39 B.n11 VSUBS 0.010468f
C40 B.n12 VSUBS 0.010468f
C41 B.n13 VSUBS 0.010468f
C42 B.n14 VSUBS 0.010468f
C43 B.n15 VSUBS 0.010468f
C44 B.n16 VSUBS 0.010468f
C45 B.n17 VSUBS 0.010468f
C46 B.n18 VSUBS 0.010468f
C47 B.n19 VSUBS 0.010468f
C48 B.n20 VSUBS 0.010468f
C49 B.n21 VSUBS 0.010468f
C50 B.n22 VSUBS 0.010468f
C51 B.n23 VSUBS 0.010468f
C52 B.n24 VSUBS 0.010468f
C53 B.n25 VSUBS 0.010468f
C54 B.n26 VSUBS 0.010468f
C55 B.n27 VSUBS 0.010468f
C56 B.n28 VSUBS 0.010468f
C57 B.n29 VSUBS 0.010468f
C58 B.n30 VSUBS 0.010468f
C59 B.n31 VSUBS 0.022897f
C60 B.n32 VSUBS 0.010468f
C61 B.n33 VSUBS 0.010468f
C62 B.n34 VSUBS 0.010468f
C63 B.n35 VSUBS 0.010468f
C64 B.n36 VSUBS 0.010468f
C65 B.n37 VSUBS 0.010468f
C66 B.t8 VSUBS 0.07765f
C67 B.t7 VSUBS 0.099814f
C68 B.t6 VSUBS 0.534866f
C69 B.n38 VSUBS 0.119777f
C70 B.n39 VSUBS 0.094915f
C71 B.n40 VSUBS 0.024253f
C72 B.n41 VSUBS 0.010468f
C73 B.n42 VSUBS 0.010468f
C74 B.n43 VSUBS 0.010468f
C75 B.n44 VSUBS 0.010468f
C76 B.n45 VSUBS 0.010468f
C77 B.t2 VSUBS 0.07765f
C78 B.t1 VSUBS 0.099814f
C79 B.t0 VSUBS 0.534866f
C80 B.n46 VSUBS 0.119777f
C81 B.n47 VSUBS 0.094915f
C82 B.n48 VSUBS 0.010468f
C83 B.n49 VSUBS 0.010468f
C84 B.n50 VSUBS 0.010468f
C85 B.n51 VSUBS 0.010468f
C86 B.n52 VSUBS 0.010468f
C87 B.n53 VSUBS 0.010468f
C88 B.n54 VSUBS 0.024224f
C89 B.n55 VSUBS 0.010468f
C90 B.n56 VSUBS 0.010468f
C91 B.n57 VSUBS 0.010468f
C92 B.n58 VSUBS 0.010468f
C93 B.n59 VSUBS 0.010468f
C94 B.n60 VSUBS 0.010468f
C95 B.n61 VSUBS 0.010468f
C96 B.n62 VSUBS 0.010468f
C97 B.n63 VSUBS 0.010468f
C98 B.n64 VSUBS 0.010468f
C99 B.n65 VSUBS 0.010468f
C100 B.n66 VSUBS 0.010468f
C101 B.n67 VSUBS 0.010468f
C102 B.n68 VSUBS 0.010468f
C103 B.n69 VSUBS 0.010468f
C104 B.n70 VSUBS 0.010468f
C105 B.n71 VSUBS 0.010468f
C106 B.n72 VSUBS 0.010468f
C107 B.n73 VSUBS 0.010468f
C108 B.n74 VSUBS 0.010468f
C109 B.n75 VSUBS 0.010468f
C110 B.n76 VSUBS 0.010468f
C111 B.n77 VSUBS 0.010468f
C112 B.n78 VSUBS 0.010468f
C113 B.n79 VSUBS 0.010468f
C114 B.n80 VSUBS 0.010468f
C115 B.n81 VSUBS 0.010468f
C116 B.n82 VSUBS 0.010468f
C117 B.n83 VSUBS 0.010468f
C118 B.n84 VSUBS 0.010468f
C119 B.n85 VSUBS 0.010468f
C120 B.n86 VSUBS 0.010468f
C121 B.n87 VSUBS 0.010468f
C122 B.n88 VSUBS 0.010468f
C123 B.n89 VSUBS 0.010468f
C124 B.n90 VSUBS 0.010468f
C125 B.n91 VSUBS 0.010468f
C126 B.n92 VSUBS 0.010468f
C127 B.n93 VSUBS 0.010468f
C128 B.n94 VSUBS 0.010468f
C129 B.n95 VSUBS 0.010468f
C130 B.n96 VSUBS 0.010468f
C131 B.n97 VSUBS 0.010468f
C132 B.n98 VSUBS 0.010468f
C133 B.n99 VSUBS 0.010468f
C134 B.n100 VSUBS 0.010468f
C135 B.n101 VSUBS 0.010468f
C136 B.n102 VSUBS 0.010468f
C137 B.n103 VSUBS 0.010468f
C138 B.n104 VSUBS 0.010468f
C139 B.n105 VSUBS 0.010468f
C140 B.n106 VSUBS 0.010468f
C141 B.n107 VSUBS 0.010468f
C142 B.n108 VSUBS 0.010468f
C143 B.n109 VSUBS 0.010468f
C144 B.n110 VSUBS 0.010468f
C145 B.n111 VSUBS 0.010468f
C146 B.n112 VSUBS 0.010468f
C147 B.n113 VSUBS 0.022897f
C148 B.n114 VSUBS 0.010468f
C149 B.n115 VSUBS 0.010468f
C150 B.n116 VSUBS 0.010468f
C151 B.n117 VSUBS 0.010468f
C152 B.n118 VSUBS 0.010468f
C153 B.n119 VSUBS 0.010468f
C154 B.t4 VSUBS 0.07765f
C155 B.t5 VSUBS 0.099814f
C156 B.t3 VSUBS 0.534866f
C157 B.n120 VSUBS 0.119777f
C158 B.n121 VSUBS 0.094915f
C159 B.n122 VSUBS 0.024253f
C160 B.n123 VSUBS 0.010468f
C161 B.n124 VSUBS 0.010468f
C162 B.n125 VSUBS 0.010468f
C163 B.n126 VSUBS 0.010468f
C164 B.n127 VSUBS 0.010468f
C165 B.t10 VSUBS 0.07765f
C166 B.t11 VSUBS 0.099814f
C167 B.t9 VSUBS 0.534866f
C168 B.n128 VSUBS 0.119777f
C169 B.n129 VSUBS 0.094915f
C170 B.n130 VSUBS 0.010468f
C171 B.n131 VSUBS 0.010468f
C172 B.n132 VSUBS 0.010468f
C173 B.n133 VSUBS 0.010468f
C174 B.n134 VSUBS 0.010468f
C175 B.n135 VSUBS 0.010468f
C176 B.n136 VSUBS 0.022897f
C177 B.n137 VSUBS 0.010468f
C178 B.n138 VSUBS 0.010468f
C179 B.n139 VSUBS 0.010468f
C180 B.n140 VSUBS 0.010468f
C181 B.n141 VSUBS 0.010468f
C182 B.n142 VSUBS 0.010468f
C183 B.n143 VSUBS 0.010468f
C184 B.n144 VSUBS 0.010468f
C185 B.n145 VSUBS 0.010468f
C186 B.n146 VSUBS 0.010468f
C187 B.n147 VSUBS 0.010468f
C188 B.n148 VSUBS 0.010468f
C189 B.n149 VSUBS 0.010468f
C190 B.n150 VSUBS 0.010468f
C191 B.n151 VSUBS 0.010468f
C192 B.n152 VSUBS 0.010468f
C193 B.n153 VSUBS 0.010468f
C194 B.n154 VSUBS 0.010468f
C195 B.n155 VSUBS 0.010468f
C196 B.n156 VSUBS 0.010468f
C197 B.n157 VSUBS 0.010468f
C198 B.n158 VSUBS 0.010468f
C199 B.n159 VSUBS 0.010468f
C200 B.n160 VSUBS 0.010468f
C201 B.n161 VSUBS 0.010468f
C202 B.n162 VSUBS 0.010468f
C203 B.n163 VSUBS 0.010468f
C204 B.n164 VSUBS 0.010468f
C205 B.n165 VSUBS 0.010468f
C206 B.n166 VSUBS 0.010468f
C207 B.n167 VSUBS 0.010468f
C208 B.n168 VSUBS 0.010468f
C209 B.n169 VSUBS 0.010468f
C210 B.n170 VSUBS 0.010468f
C211 B.n171 VSUBS 0.010468f
C212 B.n172 VSUBS 0.010468f
C213 B.n173 VSUBS 0.010468f
C214 B.n174 VSUBS 0.010468f
C215 B.n175 VSUBS 0.010468f
C216 B.n176 VSUBS 0.010468f
C217 B.n177 VSUBS 0.010468f
C218 B.n178 VSUBS 0.010468f
C219 B.n179 VSUBS 0.010468f
C220 B.n180 VSUBS 0.010468f
C221 B.n181 VSUBS 0.010468f
C222 B.n182 VSUBS 0.010468f
C223 B.n183 VSUBS 0.010468f
C224 B.n184 VSUBS 0.010468f
C225 B.n185 VSUBS 0.010468f
C226 B.n186 VSUBS 0.010468f
C227 B.n187 VSUBS 0.010468f
C228 B.n188 VSUBS 0.010468f
C229 B.n189 VSUBS 0.010468f
C230 B.n190 VSUBS 0.010468f
C231 B.n191 VSUBS 0.010468f
C232 B.n192 VSUBS 0.010468f
C233 B.n193 VSUBS 0.010468f
C234 B.n194 VSUBS 0.010468f
C235 B.n195 VSUBS 0.010468f
C236 B.n196 VSUBS 0.010468f
C237 B.n197 VSUBS 0.010468f
C238 B.n198 VSUBS 0.010468f
C239 B.n199 VSUBS 0.010468f
C240 B.n200 VSUBS 0.010468f
C241 B.n201 VSUBS 0.010468f
C242 B.n202 VSUBS 0.010468f
C243 B.n203 VSUBS 0.010468f
C244 B.n204 VSUBS 0.010468f
C245 B.n205 VSUBS 0.010468f
C246 B.n206 VSUBS 0.010468f
C247 B.n207 VSUBS 0.010468f
C248 B.n208 VSUBS 0.010468f
C249 B.n209 VSUBS 0.010468f
C250 B.n210 VSUBS 0.010468f
C251 B.n211 VSUBS 0.010468f
C252 B.n212 VSUBS 0.010468f
C253 B.n213 VSUBS 0.010468f
C254 B.n214 VSUBS 0.010468f
C255 B.n215 VSUBS 0.010468f
C256 B.n216 VSUBS 0.010468f
C257 B.n217 VSUBS 0.010468f
C258 B.n218 VSUBS 0.010468f
C259 B.n219 VSUBS 0.010468f
C260 B.n220 VSUBS 0.010468f
C261 B.n221 VSUBS 0.010468f
C262 B.n222 VSUBS 0.010468f
C263 B.n223 VSUBS 0.010468f
C264 B.n224 VSUBS 0.010468f
C265 B.n225 VSUBS 0.010468f
C266 B.n226 VSUBS 0.010468f
C267 B.n227 VSUBS 0.010468f
C268 B.n228 VSUBS 0.010468f
C269 B.n229 VSUBS 0.010468f
C270 B.n230 VSUBS 0.010468f
C271 B.n231 VSUBS 0.010468f
C272 B.n232 VSUBS 0.010468f
C273 B.n233 VSUBS 0.010468f
C274 B.n234 VSUBS 0.010468f
C275 B.n235 VSUBS 0.010468f
C276 B.n236 VSUBS 0.010468f
C277 B.n237 VSUBS 0.010468f
C278 B.n238 VSUBS 0.010468f
C279 B.n239 VSUBS 0.010468f
C280 B.n240 VSUBS 0.010468f
C281 B.n241 VSUBS 0.010468f
C282 B.n242 VSUBS 0.010468f
C283 B.n243 VSUBS 0.010468f
C284 B.n244 VSUBS 0.010468f
C285 B.n245 VSUBS 0.010468f
C286 B.n246 VSUBS 0.010468f
C287 B.n247 VSUBS 0.010468f
C288 B.n248 VSUBS 0.010468f
C289 B.n249 VSUBS 0.010468f
C290 B.n250 VSUBS 0.010468f
C291 B.n251 VSUBS 0.022897f
C292 B.n252 VSUBS 0.023901f
C293 B.n253 VSUBS 0.023901f
C294 B.n254 VSUBS 0.010468f
C295 B.n255 VSUBS 0.010468f
C296 B.n256 VSUBS 0.010468f
C297 B.n257 VSUBS 0.010468f
C298 B.n258 VSUBS 0.010468f
C299 B.n259 VSUBS 0.010468f
C300 B.n260 VSUBS 0.010468f
C301 B.n261 VSUBS 0.010468f
C302 B.n262 VSUBS 0.010468f
C303 B.n263 VSUBS 0.010468f
C304 B.n264 VSUBS 0.010468f
C305 B.n265 VSUBS 0.010468f
C306 B.n266 VSUBS 0.010468f
C307 B.n267 VSUBS 0.010468f
C308 B.n268 VSUBS 0.010468f
C309 B.n269 VSUBS 0.010468f
C310 B.n270 VSUBS 0.010468f
C311 B.n271 VSUBS 0.009852f
C312 B.n272 VSUBS 0.024253f
C313 B.n273 VSUBS 0.00585f
C314 B.n274 VSUBS 0.010468f
C315 B.n275 VSUBS 0.010468f
C316 B.n276 VSUBS 0.010468f
C317 B.n277 VSUBS 0.010468f
C318 B.n278 VSUBS 0.010468f
C319 B.n279 VSUBS 0.010468f
C320 B.n280 VSUBS 0.010468f
C321 B.n281 VSUBS 0.010468f
C322 B.n282 VSUBS 0.010468f
C323 B.n283 VSUBS 0.010468f
C324 B.n284 VSUBS 0.010468f
C325 B.n285 VSUBS 0.010468f
C326 B.n286 VSUBS 0.00585f
C327 B.n287 VSUBS 0.010468f
C328 B.n288 VSUBS 0.010468f
C329 B.n289 VSUBS 0.009852f
C330 B.n290 VSUBS 0.010468f
C331 B.n291 VSUBS 0.010468f
C332 B.n292 VSUBS 0.010468f
C333 B.n293 VSUBS 0.010468f
C334 B.n294 VSUBS 0.010468f
C335 B.n295 VSUBS 0.010468f
C336 B.n296 VSUBS 0.010468f
C337 B.n297 VSUBS 0.010468f
C338 B.n298 VSUBS 0.010468f
C339 B.n299 VSUBS 0.010468f
C340 B.n300 VSUBS 0.010468f
C341 B.n301 VSUBS 0.010468f
C342 B.n302 VSUBS 0.010468f
C343 B.n303 VSUBS 0.010468f
C344 B.n304 VSUBS 0.010468f
C345 B.n305 VSUBS 0.010468f
C346 B.n306 VSUBS 0.023901f
C347 B.n307 VSUBS 0.023901f
C348 B.n308 VSUBS 0.022897f
C349 B.n309 VSUBS 0.010468f
C350 B.n310 VSUBS 0.010468f
C351 B.n311 VSUBS 0.010468f
C352 B.n312 VSUBS 0.010468f
C353 B.n313 VSUBS 0.010468f
C354 B.n314 VSUBS 0.010468f
C355 B.n315 VSUBS 0.010468f
C356 B.n316 VSUBS 0.010468f
C357 B.n317 VSUBS 0.010468f
C358 B.n318 VSUBS 0.010468f
C359 B.n319 VSUBS 0.010468f
C360 B.n320 VSUBS 0.010468f
C361 B.n321 VSUBS 0.010468f
C362 B.n322 VSUBS 0.010468f
C363 B.n323 VSUBS 0.010468f
C364 B.n324 VSUBS 0.010468f
C365 B.n325 VSUBS 0.010468f
C366 B.n326 VSUBS 0.010468f
C367 B.n327 VSUBS 0.010468f
C368 B.n328 VSUBS 0.010468f
C369 B.n329 VSUBS 0.010468f
C370 B.n330 VSUBS 0.010468f
C371 B.n331 VSUBS 0.010468f
C372 B.n332 VSUBS 0.010468f
C373 B.n333 VSUBS 0.010468f
C374 B.n334 VSUBS 0.010468f
C375 B.n335 VSUBS 0.010468f
C376 B.n336 VSUBS 0.010468f
C377 B.n337 VSUBS 0.010468f
C378 B.n338 VSUBS 0.010468f
C379 B.n339 VSUBS 0.010468f
C380 B.n340 VSUBS 0.010468f
C381 B.n341 VSUBS 0.010468f
C382 B.n342 VSUBS 0.010468f
C383 B.n343 VSUBS 0.010468f
C384 B.n344 VSUBS 0.010468f
C385 B.n345 VSUBS 0.010468f
C386 B.n346 VSUBS 0.010468f
C387 B.n347 VSUBS 0.010468f
C388 B.n348 VSUBS 0.010468f
C389 B.n349 VSUBS 0.010468f
C390 B.n350 VSUBS 0.010468f
C391 B.n351 VSUBS 0.010468f
C392 B.n352 VSUBS 0.010468f
C393 B.n353 VSUBS 0.010468f
C394 B.n354 VSUBS 0.010468f
C395 B.n355 VSUBS 0.010468f
C396 B.n356 VSUBS 0.010468f
C397 B.n357 VSUBS 0.010468f
C398 B.n358 VSUBS 0.010468f
C399 B.n359 VSUBS 0.010468f
C400 B.n360 VSUBS 0.010468f
C401 B.n361 VSUBS 0.010468f
C402 B.n362 VSUBS 0.010468f
C403 B.n363 VSUBS 0.010468f
C404 B.n364 VSUBS 0.010468f
C405 B.n365 VSUBS 0.010468f
C406 B.n366 VSUBS 0.010468f
C407 B.n367 VSUBS 0.010468f
C408 B.n368 VSUBS 0.010468f
C409 B.n369 VSUBS 0.010468f
C410 B.n370 VSUBS 0.010468f
C411 B.n371 VSUBS 0.010468f
C412 B.n372 VSUBS 0.010468f
C413 B.n373 VSUBS 0.010468f
C414 B.n374 VSUBS 0.010468f
C415 B.n375 VSUBS 0.010468f
C416 B.n376 VSUBS 0.010468f
C417 B.n377 VSUBS 0.010468f
C418 B.n378 VSUBS 0.010468f
C419 B.n379 VSUBS 0.010468f
C420 B.n380 VSUBS 0.010468f
C421 B.n381 VSUBS 0.010468f
C422 B.n382 VSUBS 0.010468f
C423 B.n383 VSUBS 0.010468f
C424 B.n384 VSUBS 0.010468f
C425 B.n385 VSUBS 0.010468f
C426 B.n386 VSUBS 0.010468f
C427 B.n387 VSUBS 0.010468f
C428 B.n388 VSUBS 0.010468f
C429 B.n389 VSUBS 0.010468f
C430 B.n390 VSUBS 0.010468f
C431 B.n391 VSUBS 0.010468f
C432 B.n392 VSUBS 0.010468f
C433 B.n393 VSUBS 0.010468f
C434 B.n394 VSUBS 0.010468f
C435 B.n395 VSUBS 0.010468f
C436 B.n396 VSUBS 0.010468f
C437 B.n397 VSUBS 0.010468f
C438 B.n398 VSUBS 0.010468f
C439 B.n399 VSUBS 0.010468f
C440 B.n400 VSUBS 0.010468f
C441 B.n401 VSUBS 0.010468f
C442 B.n402 VSUBS 0.010468f
C443 B.n403 VSUBS 0.010468f
C444 B.n404 VSUBS 0.010468f
C445 B.n405 VSUBS 0.010468f
C446 B.n406 VSUBS 0.010468f
C447 B.n407 VSUBS 0.010468f
C448 B.n408 VSUBS 0.010468f
C449 B.n409 VSUBS 0.010468f
C450 B.n410 VSUBS 0.010468f
C451 B.n411 VSUBS 0.010468f
C452 B.n412 VSUBS 0.010468f
C453 B.n413 VSUBS 0.010468f
C454 B.n414 VSUBS 0.010468f
C455 B.n415 VSUBS 0.010468f
C456 B.n416 VSUBS 0.010468f
C457 B.n417 VSUBS 0.010468f
C458 B.n418 VSUBS 0.010468f
C459 B.n419 VSUBS 0.010468f
C460 B.n420 VSUBS 0.010468f
C461 B.n421 VSUBS 0.010468f
C462 B.n422 VSUBS 0.010468f
C463 B.n423 VSUBS 0.010468f
C464 B.n424 VSUBS 0.010468f
C465 B.n425 VSUBS 0.010468f
C466 B.n426 VSUBS 0.010468f
C467 B.n427 VSUBS 0.010468f
C468 B.n428 VSUBS 0.010468f
C469 B.n429 VSUBS 0.010468f
C470 B.n430 VSUBS 0.010468f
C471 B.n431 VSUBS 0.010468f
C472 B.n432 VSUBS 0.010468f
C473 B.n433 VSUBS 0.010468f
C474 B.n434 VSUBS 0.010468f
C475 B.n435 VSUBS 0.010468f
C476 B.n436 VSUBS 0.010468f
C477 B.n437 VSUBS 0.010468f
C478 B.n438 VSUBS 0.010468f
C479 B.n439 VSUBS 0.010468f
C480 B.n440 VSUBS 0.010468f
C481 B.n441 VSUBS 0.010468f
C482 B.n442 VSUBS 0.010468f
C483 B.n443 VSUBS 0.010468f
C484 B.n444 VSUBS 0.010468f
C485 B.n445 VSUBS 0.010468f
C486 B.n446 VSUBS 0.010468f
C487 B.n447 VSUBS 0.010468f
C488 B.n448 VSUBS 0.010468f
C489 B.n449 VSUBS 0.010468f
C490 B.n450 VSUBS 0.010468f
C491 B.n451 VSUBS 0.010468f
C492 B.n452 VSUBS 0.010468f
C493 B.n453 VSUBS 0.010468f
C494 B.n454 VSUBS 0.010468f
C495 B.n455 VSUBS 0.010468f
C496 B.n456 VSUBS 0.010468f
C497 B.n457 VSUBS 0.010468f
C498 B.n458 VSUBS 0.010468f
C499 B.n459 VSUBS 0.010468f
C500 B.n460 VSUBS 0.010468f
C501 B.n461 VSUBS 0.010468f
C502 B.n462 VSUBS 0.010468f
C503 B.n463 VSUBS 0.010468f
C504 B.n464 VSUBS 0.010468f
C505 B.n465 VSUBS 0.010468f
C506 B.n466 VSUBS 0.010468f
C507 B.n467 VSUBS 0.010468f
C508 B.n468 VSUBS 0.010468f
C509 B.n469 VSUBS 0.010468f
C510 B.n470 VSUBS 0.010468f
C511 B.n471 VSUBS 0.010468f
C512 B.n472 VSUBS 0.010468f
C513 B.n473 VSUBS 0.010468f
C514 B.n474 VSUBS 0.010468f
C515 B.n475 VSUBS 0.010468f
C516 B.n476 VSUBS 0.010468f
C517 B.n477 VSUBS 0.010468f
C518 B.n478 VSUBS 0.010468f
C519 B.n479 VSUBS 0.010468f
C520 B.n480 VSUBS 0.010468f
C521 B.n481 VSUBS 0.010468f
C522 B.n482 VSUBS 0.010468f
C523 B.n483 VSUBS 0.010468f
C524 B.n484 VSUBS 0.010468f
C525 B.n485 VSUBS 0.022897f
C526 B.n486 VSUBS 0.023901f
C527 B.n487 VSUBS 0.022574f
C528 B.n488 VSUBS 0.010468f
C529 B.n489 VSUBS 0.010468f
C530 B.n490 VSUBS 0.010468f
C531 B.n491 VSUBS 0.010468f
C532 B.n492 VSUBS 0.010468f
C533 B.n493 VSUBS 0.010468f
C534 B.n494 VSUBS 0.010468f
C535 B.n495 VSUBS 0.010468f
C536 B.n496 VSUBS 0.010468f
C537 B.n497 VSUBS 0.010468f
C538 B.n498 VSUBS 0.010468f
C539 B.n499 VSUBS 0.010468f
C540 B.n500 VSUBS 0.010468f
C541 B.n501 VSUBS 0.010468f
C542 B.n502 VSUBS 0.010468f
C543 B.n503 VSUBS 0.010468f
C544 B.n504 VSUBS 0.010468f
C545 B.n505 VSUBS 0.009852f
C546 B.n506 VSUBS 0.024253f
C547 B.n507 VSUBS 0.00585f
C548 B.n508 VSUBS 0.010468f
C549 B.n509 VSUBS 0.010468f
C550 B.n510 VSUBS 0.010468f
C551 B.n511 VSUBS 0.010468f
C552 B.n512 VSUBS 0.010468f
C553 B.n513 VSUBS 0.010468f
C554 B.n514 VSUBS 0.010468f
C555 B.n515 VSUBS 0.010468f
C556 B.n516 VSUBS 0.010468f
C557 B.n517 VSUBS 0.010468f
C558 B.n518 VSUBS 0.010468f
C559 B.n519 VSUBS 0.010468f
C560 B.n520 VSUBS 0.00585f
C561 B.n521 VSUBS 0.010468f
C562 B.n522 VSUBS 0.010468f
C563 B.n523 VSUBS 0.009852f
C564 B.n524 VSUBS 0.010468f
C565 B.n525 VSUBS 0.010468f
C566 B.n526 VSUBS 0.010468f
C567 B.n527 VSUBS 0.010468f
C568 B.n528 VSUBS 0.010468f
C569 B.n529 VSUBS 0.010468f
C570 B.n530 VSUBS 0.010468f
C571 B.n531 VSUBS 0.010468f
C572 B.n532 VSUBS 0.010468f
C573 B.n533 VSUBS 0.010468f
C574 B.n534 VSUBS 0.010468f
C575 B.n535 VSUBS 0.010468f
C576 B.n536 VSUBS 0.010468f
C577 B.n537 VSUBS 0.010468f
C578 B.n538 VSUBS 0.010468f
C579 B.n539 VSUBS 0.010468f
C580 B.n540 VSUBS 0.023901f
C581 B.n541 VSUBS 0.023901f
C582 B.n542 VSUBS 0.022897f
C583 B.n543 VSUBS 0.010468f
C584 B.n544 VSUBS 0.010468f
C585 B.n545 VSUBS 0.010468f
C586 B.n546 VSUBS 0.010468f
C587 B.n547 VSUBS 0.010468f
C588 B.n548 VSUBS 0.010468f
C589 B.n549 VSUBS 0.010468f
C590 B.n550 VSUBS 0.010468f
C591 B.n551 VSUBS 0.010468f
C592 B.n552 VSUBS 0.010468f
C593 B.n553 VSUBS 0.010468f
C594 B.n554 VSUBS 0.010468f
C595 B.n555 VSUBS 0.010468f
C596 B.n556 VSUBS 0.010468f
C597 B.n557 VSUBS 0.010468f
C598 B.n558 VSUBS 0.010468f
C599 B.n559 VSUBS 0.010468f
C600 B.n560 VSUBS 0.010468f
C601 B.n561 VSUBS 0.010468f
C602 B.n562 VSUBS 0.010468f
C603 B.n563 VSUBS 0.010468f
C604 B.n564 VSUBS 0.010468f
C605 B.n565 VSUBS 0.010468f
C606 B.n566 VSUBS 0.010468f
C607 B.n567 VSUBS 0.010468f
C608 B.n568 VSUBS 0.010468f
C609 B.n569 VSUBS 0.010468f
C610 B.n570 VSUBS 0.010468f
C611 B.n571 VSUBS 0.010468f
C612 B.n572 VSUBS 0.010468f
C613 B.n573 VSUBS 0.010468f
C614 B.n574 VSUBS 0.010468f
C615 B.n575 VSUBS 0.010468f
C616 B.n576 VSUBS 0.010468f
C617 B.n577 VSUBS 0.010468f
C618 B.n578 VSUBS 0.010468f
C619 B.n579 VSUBS 0.010468f
C620 B.n580 VSUBS 0.010468f
C621 B.n581 VSUBS 0.010468f
C622 B.n582 VSUBS 0.010468f
C623 B.n583 VSUBS 0.010468f
C624 B.n584 VSUBS 0.010468f
C625 B.n585 VSUBS 0.010468f
C626 B.n586 VSUBS 0.010468f
C627 B.n587 VSUBS 0.010468f
C628 B.n588 VSUBS 0.010468f
C629 B.n589 VSUBS 0.010468f
C630 B.n590 VSUBS 0.010468f
C631 B.n591 VSUBS 0.010468f
C632 B.n592 VSUBS 0.010468f
C633 B.n593 VSUBS 0.010468f
C634 B.n594 VSUBS 0.010468f
C635 B.n595 VSUBS 0.010468f
C636 B.n596 VSUBS 0.010468f
C637 B.n597 VSUBS 0.010468f
C638 B.n598 VSUBS 0.010468f
C639 B.n599 VSUBS 0.010468f
C640 B.n600 VSUBS 0.010468f
C641 B.n601 VSUBS 0.010468f
C642 B.n602 VSUBS 0.010468f
C643 B.n603 VSUBS 0.010468f
C644 B.n604 VSUBS 0.010468f
C645 B.n605 VSUBS 0.010468f
C646 B.n606 VSUBS 0.010468f
C647 B.n607 VSUBS 0.010468f
C648 B.n608 VSUBS 0.010468f
C649 B.n609 VSUBS 0.010468f
C650 B.n610 VSUBS 0.010468f
C651 B.n611 VSUBS 0.010468f
C652 B.n612 VSUBS 0.010468f
C653 B.n613 VSUBS 0.010468f
C654 B.n614 VSUBS 0.010468f
C655 B.n615 VSUBS 0.010468f
C656 B.n616 VSUBS 0.010468f
C657 B.n617 VSUBS 0.010468f
C658 B.n618 VSUBS 0.010468f
C659 B.n619 VSUBS 0.010468f
C660 B.n620 VSUBS 0.010468f
C661 B.n621 VSUBS 0.010468f
C662 B.n622 VSUBS 0.010468f
C663 B.n623 VSUBS 0.010468f
C664 B.n624 VSUBS 0.010468f
C665 B.n625 VSUBS 0.010468f
C666 B.n626 VSUBS 0.010468f
C667 B.n627 VSUBS 0.010468f
C668 B.n628 VSUBS 0.010468f
C669 B.n629 VSUBS 0.010468f
C670 B.n630 VSUBS 0.010468f
C671 B.n631 VSUBS 0.023703f
C672 VDD1.t3 VSUBS 0.057495f
C673 VDD1.t2 VSUBS 0.057495f
C674 VDD1.n0 VSUBS 0.265517f
C675 VDD1.t7 VSUBS 0.057495f
C676 VDD1.t6 VSUBS 0.057495f
C677 VDD1.n1 VSUBS 0.264881f
C678 VDD1.t5 VSUBS 0.057495f
C679 VDD1.t0 VSUBS 0.057495f
C680 VDD1.n2 VSUBS 0.264881f
C681 VDD1.n3 VSUBS 4.03466f
C682 VDD1.t4 VSUBS 0.057495f
C683 VDD1.t1 VSUBS 0.057495f
C684 VDD1.n4 VSUBS 0.258039f
C685 VDD1.n5 VSUBS 3.12449f
C686 VP.t7 VSUBS 0.96975f
C687 VP.n0 VSUBS 0.658699f
C688 VP.n1 VSUBS 0.055547f
C689 VP.n2 VSUBS 0.073349f
C690 VP.n3 VSUBS 0.055547f
C691 VP.t2 VSUBS 0.96975f
C692 VP.n4 VSUBS 0.428321f
C693 VP.n5 VSUBS 0.055547f
C694 VP.n6 VSUBS 0.081088f
C695 VP.n7 VSUBS 0.055547f
C696 VP.t1 VSUBS 0.96975f
C697 VP.n8 VSUBS 0.103525f
C698 VP.n9 VSUBS 0.055547f
C699 VP.n10 VSUBS 0.103525f
C700 VP.t6 VSUBS 0.96975f
C701 VP.n11 VSUBS 0.658699f
C702 VP.n12 VSUBS 0.055547f
C703 VP.n13 VSUBS 0.073349f
C704 VP.n14 VSUBS 0.055547f
C705 VP.t3 VSUBS 0.96975f
C706 VP.n15 VSUBS 0.428321f
C707 VP.n16 VSUBS 0.055547f
C708 VP.n17 VSUBS 0.081088f
C709 VP.n18 VSUBS 0.633578f
C710 VP.t5 VSUBS 0.96975f
C711 VP.t4 VSUBS 1.50736f
C712 VP.n19 VSUBS 0.617003f
C713 VP.n20 VSUBS 0.63431f
C714 VP.n21 VSUBS 0.100967f
C715 VP.n22 VSUBS 0.103525f
C716 VP.n23 VSUBS 0.055547f
C717 VP.n24 VSUBS 0.055547f
C718 VP.n25 VSUBS 0.055547f
C719 VP.n26 VSUBS 0.081088f
C720 VP.n27 VSUBS 0.103525f
C721 VP.n28 VSUBS 0.100967f
C722 VP.n29 VSUBS 0.055547f
C723 VP.n30 VSUBS 0.055547f
C724 VP.n31 VSUBS 0.054967f
C725 VP.n32 VSUBS 0.103525f
C726 VP.n33 VSUBS 0.103525f
C727 VP.n34 VSUBS 0.055547f
C728 VP.n35 VSUBS 0.055547f
C729 VP.n36 VSUBS 0.055547f
C730 VP.n37 VSUBS 0.088828f
C731 VP.n38 VSUBS 0.103525f
C732 VP.n39 VSUBS 0.095856f
C733 VP.n40 VSUBS 0.089651f
C734 VP.n41 VSUBS 2.79445f
C735 VP.n42 VSUBS 2.8377f
C736 VP.t0 VSUBS 0.96975f
C737 VP.n43 VSUBS 0.658699f
C738 VP.n44 VSUBS 0.095856f
C739 VP.n45 VSUBS 0.089651f
C740 VP.n46 VSUBS 0.055547f
C741 VP.n47 VSUBS 0.055547f
C742 VP.n48 VSUBS 0.088828f
C743 VP.n49 VSUBS 0.073349f
C744 VP.n50 VSUBS 0.103525f
C745 VP.n51 VSUBS 0.055547f
C746 VP.n52 VSUBS 0.055547f
C747 VP.n53 VSUBS 0.055547f
C748 VP.n54 VSUBS 0.054967f
C749 VP.n55 VSUBS 0.428321f
C750 VP.n56 VSUBS 0.100967f
C751 VP.n57 VSUBS 0.103525f
C752 VP.n58 VSUBS 0.055547f
C753 VP.n59 VSUBS 0.055547f
C754 VP.n60 VSUBS 0.055547f
C755 VP.n61 VSUBS 0.081088f
C756 VP.n62 VSUBS 0.103525f
C757 VP.n63 VSUBS 0.100967f
C758 VP.n64 VSUBS 0.055547f
C759 VP.n65 VSUBS 0.055547f
C760 VP.n66 VSUBS 0.054967f
C761 VP.n67 VSUBS 0.103525f
C762 VP.n68 VSUBS 0.103525f
C763 VP.n69 VSUBS 0.055547f
C764 VP.n70 VSUBS 0.055547f
C765 VP.n71 VSUBS 0.055547f
C766 VP.n72 VSUBS 0.088828f
C767 VP.n73 VSUBS 0.103525f
C768 VP.n74 VSUBS 0.095856f
C769 VP.n75 VSUBS 0.089651f
C770 VP.n76 VSUBS 0.115658f
C771 VTAIL.t10 VSUBS 0.064755f
C772 VTAIL.t11 VSUBS 0.064755f
C773 VTAIL.n0 VSUBS 0.246532f
C774 VTAIL.n1 VSUBS 0.754935f
C775 VTAIL.t15 VSUBS 0.393451f
C776 VTAIL.n2 VSUBS 0.831267f
C777 VTAIL.t5 VSUBS 0.393451f
C778 VTAIL.n3 VSUBS 0.831267f
C779 VTAIL.t4 VSUBS 0.064755f
C780 VTAIL.t2 VSUBS 0.064755f
C781 VTAIL.n4 VSUBS 0.246532f
C782 VTAIL.n5 VSUBS 1.08538f
C783 VTAIL.t0 VSUBS 0.393451f
C784 VTAIL.n6 VSUBS 1.82041f
C785 VTAIL.t9 VSUBS 0.393452f
C786 VTAIL.n7 VSUBS 1.82041f
C787 VTAIL.t8 VSUBS 0.064755f
C788 VTAIL.t12 VSUBS 0.064755f
C789 VTAIL.n8 VSUBS 0.246533f
C790 VTAIL.n9 VSUBS 1.08538f
C791 VTAIL.t13 VSUBS 0.393452f
C792 VTAIL.n10 VSUBS 0.831266f
C793 VTAIL.t1 VSUBS 0.393452f
C794 VTAIL.n11 VSUBS 0.831266f
C795 VTAIL.t3 VSUBS 0.064755f
C796 VTAIL.t7 VSUBS 0.064755f
C797 VTAIL.n12 VSUBS 0.246533f
C798 VTAIL.n13 VSUBS 1.08538f
C799 VTAIL.t6 VSUBS 0.393452f
C800 VTAIL.n14 VSUBS 1.82041f
C801 VTAIL.t14 VSUBS 0.393451f
C802 VTAIL.n15 VSUBS 1.81382f
C803 VDD2.t0 VSUBS 0.055805f
C804 VDD2.t1 VSUBS 0.055805f
C805 VDD2.n0 VSUBS 0.257095f
C806 VDD2.t5 VSUBS 0.055805f
C807 VDD2.t3 VSUBS 0.055805f
C808 VDD2.n1 VSUBS 0.257095f
C809 VDD2.n2 VSUBS 3.85303f
C810 VDD2.t4 VSUBS 0.055805f
C811 VDD2.t2 VSUBS 0.055805f
C812 VDD2.n3 VSUBS 0.250454f
C813 VDD2.n4 VSUBS 2.99511f
C814 VDD2.t6 VSUBS 0.055805f
C815 VDD2.t7 VSUBS 0.055805f
C816 VDD2.n5 VSUBS 0.257077f
C817 VN.t1 VSUBS 0.838812f
C818 VN.n0 VSUBS 0.56976f
C819 VN.n1 VSUBS 0.048047f
C820 VN.n2 VSUBS 0.063445f
C821 VN.n3 VSUBS 0.048047f
C822 VN.t4 VSUBS 0.838812f
C823 VN.n4 VSUBS 0.370488f
C824 VN.n5 VSUBS 0.048047f
C825 VN.n6 VSUBS 0.07014f
C826 VN.n7 VSUBS 0.54803f
C827 VN.t5 VSUBS 0.838812f
C828 VN.t0 VSUBS 1.30383f
C829 VN.n8 VSUBS 0.533693f
C830 VN.n9 VSUBS 0.548664f
C831 VN.n10 VSUBS 0.087334f
C832 VN.n11 VSUBS 0.089547f
C833 VN.n12 VSUBS 0.048047f
C834 VN.n13 VSUBS 0.048047f
C835 VN.n14 VSUBS 0.048047f
C836 VN.n15 VSUBS 0.07014f
C837 VN.n16 VSUBS 0.089547f
C838 VN.n17 VSUBS 0.087334f
C839 VN.n18 VSUBS 0.048047f
C840 VN.n19 VSUBS 0.048047f
C841 VN.n20 VSUBS 0.047545f
C842 VN.n21 VSUBS 0.089547f
C843 VN.n22 VSUBS 0.089547f
C844 VN.n23 VSUBS 0.048047f
C845 VN.n24 VSUBS 0.048047f
C846 VN.n25 VSUBS 0.048047f
C847 VN.n26 VSUBS 0.076834f
C848 VN.n27 VSUBS 0.089547f
C849 VN.n28 VSUBS 0.082913f
C850 VN.n29 VSUBS 0.077546f
C851 VN.n30 VSUBS 0.100042f
C852 VN.t6 VSUBS 0.838812f
C853 VN.n31 VSUBS 0.56976f
C854 VN.n32 VSUBS 0.048047f
C855 VN.n33 VSUBS 0.063445f
C856 VN.n34 VSUBS 0.048047f
C857 VN.t7 VSUBS 0.838812f
C858 VN.n35 VSUBS 0.370488f
C859 VN.n36 VSUBS 0.048047f
C860 VN.n37 VSUBS 0.07014f
C861 VN.n38 VSUBS 0.54803f
C862 VN.t3 VSUBS 0.838812f
C863 VN.t2 VSUBS 1.30383f
C864 VN.n39 VSUBS 0.533693f
C865 VN.n40 VSUBS 0.548664f
C866 VN.n41 VSUBS 0.087334f
C867 VN.n42 VSUBS 0.089547f
C868 VN.n43 VSUBS 0.048047f
C869 VN.n44 VSUBS 0.048047f
C870 VN.n45 VSUBS 0.048047f
C871 VN.n46 VSUBS 0.07014f
C872 VN.n47 VSUBS 0.089547f
C873 VN.n48 VSUBS 0.087334f
C874 VN.n49 VSUBS 0.048047f
C875 VN.n50 VSUBS 0.048047f
C876 VN.n51 VSUBS 0.047545f
C877 VN.n52 VSUBS 0.089547f
C878 VN.n53 VSUBS 0.089547f
C879 VN.n54 VSUBS 0.048047f
C880 VN.n55 VSUBS 0.048047f
C881 VN.n56 VSUBS 0.048047f
C882 VN.n57 VSUBS 0.076834f
C883 VN.n58 VSUBS 0.089547f
C884 VN.n59 VSUBS 0.082913f
C885 VN.n60 VSUBS 0.077546f
C886 VN.n61 VSUBS 2.43734f
.ends

