* NGSPICE file created from diff_pair_sample_0021.ext - technology: sky130A

.subckt diff_pair_sample_0021 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t7 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=2.2572 pd=14.01 as=5.3352 ps=28.14 w=13.68 l=0.75
X1 B.t11 B.t9 B.t10 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=5.3352 pd=28.14 as=0 ps=0 w=13.68 l=0.75
X2 VDD1.t3 VP.t0 VTAIL.t0 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=2.2572 pd=14.01 as=5.3352 ps=28.14 w=13.68 l=0.75
X3 B.t8 B.t6 B.t7 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=5.3352 pd=28.14 as=0 ps=0 w=13.68 l=0.75
X4 VDD2.t2 VN.t1 VTAIL.t5 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=2.2572 pd=14.01 as=5.3352 ps=28.14 w=13.68 l=0.75
X5 B.t5 B.t3 B.t4 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=5.3352 pd=28.14 as=0 ps=0 w=13.68 l=0.75
X6 VTAIL.t4 VN.t2 VDD2.t1 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=5.3352 pd=28.14 as=2.2572 ps=14.01 w=13.68 l=0.75
X7 VTAIL.t1 VP.t1 VDD1.t2 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=5.3352 pd=28.14 as=2.2572 ps=14.01 w=13.68 l=0.75
X8 VTAIL.t3 VP.t2 VDD1.t1 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=5.3352 pd=28.14 as=2.2572 ps=14.01 w=13.68 l=0.75
X9 B.t2 B.t0 B.t1 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=5.3352 pd=28.14 as=0 ps=0 w=13.68 l=0.75
X10 VTAIL.t6 VN.t3 VDD2.t0 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=5.3352 pd=28.14 as=2.2572 ps=14.01 w=13.68 l=0.75
X11 VDD1.t0 VP.t3 VTAIL.t2 w_n1618_n3704# sky130_fd_pr__pfet_01v8 ad=2.2572 pd=14.01 as=5.3352 ps=28.14 w=13.68 l=0.75
R0 VN.n0 VN.t3 512.958
R1 VN.n1 VN.t1 512.958
R2 VN.n0 VN.t0 512.909
R3 VN.n1 VN.t2 512.909
R4 VN VN.n1 86.914
R5 VN VN.n0 44.7132
R6 VTAIL.n5 VTAIL.t1 59.6676
R7 VTAIL.n4 VTAIL.t5 59.6676
R8 VTAIL.n3 VTAIL.t4 59.6676
R9 VTAIL.n7 VTAIL.t7 59.6674
R10 VTAIL.n0 VTAIL.t6 59.6674
R11 VTAIL.n1 VTAIL.t2 59.6674
R12 VTAIL.n2 VTAIL.t3 59.6674
R13 VTAIL.n6 VTAIL.t0 59.6674
R14 VTAIL.n7 VTAIL.n6 25.091
R15 VTAIL.n3 VTAIL.n2 25.091
R16 VTAIL.n4 VTAIL.n3 0.931535
R17 VTAIL.n6 VTAIL.n5 0.931535
R18 VTAIL.n2 VTAIL.n1 0.931535
R19 VTAIL VTAIL.n0 0.524207
R20 VTAIL.n5 VTAIL.n4 0.470328
R21 VTAIL.n1 VTAIL.n0 0.470328
R22 VTAIL VTAIL.n7 0.407828
R23 VDD2.n2 VDD2.n0 112.272
R24 VDD2.n2 VDD2.n1 73.9701
R25 VDD2.n1 VDD2.t1 2.3766
R26 VDD2.n1 VDD2.t2 2.3766
R27 VDD2.n0 VDD2.t0 2.3766
R28 VDD2.n0 VDD2.t3 2.3766
R29 VDD2 VDD2.n2 0.0586897
R30 B.n116 B.t0 641.976
R31 B.n108 B.t3 641.976
R32 B.n42 B.t9 641.976
R33 B.n34 B.t6 641.976
R34 B.n328 B.n327 585
R35 B.n326 B.n85 585
R36 B.n325 B.n324 585
R37 B.n323 B.n86 585
R38 B.n322 B.n321 585
R39 B.n320 B.n87 585
R40 B.n319 B.n318 585
R41 B.n317 B.n88 585
R42 B.n316 B.n315 585
R43 B.n314 B.n89 585
R44 B.n313 B.n312 585
R45 B.n311 B.n90 585
R46 B.n310 B.n309 585
R47 B.n308 B.n91 585
R48 B.n307 B.n306 585
R49 B.n305 B.n92 585
R50 B.n304 B.n303 585
R51 B.n302 B.n93 585
R52 B.n301 B.n300 585
R53 B.n299 B.n94 585
R54 B.n298 B.n297 585
R55 B.n296 B.n95 585
R56 B.n295 B.n294 585
R57 B.n293 B.n96 585
R58 B.n292 B.n291 585
R59 B.n290 B.n97 585
R60 B.n289 B.n288 585
R61 B.n287 B.n98 585
R62 B.n286 B.n285 585
R63 B.n284 B.n99 585
R64 B.n283 B.n282 585
R65 B.n281 B.n100 585
R66 B.n280 B.n279 585
R67 B.n278 B.n101 585
R68 B.n277 B.n276 585
R69 B.n275 B.n102 585
R70 B.n274 B.n273 585
R71 B.n272 B.n103 585
R72 B.n271 B.n270 585
R73 B.n269 B.n104 585
R74 B.n268 B.n267 585
R75 B.n266 B.n105 585
R76 B.n265 B.n264 585
R77 B.n263 B.n106 585
R78 B.n262 B.n261 585
R79 B.n260 B.n107 585
R80 B.n259 B.n258 585
R81 B.n257 B.n256 585
R82 B.n255 B.n111 585
R83 B.n254 B.n253 585
R84 B.n252 B.n112 585
R85 B.n251 B.n250 585
R86 B.n249 B.n113 585
R87 B.n248 B.n247 585
R88 B.n246 B.n114 585
R89 B.n245 B.n244 585
R90 B.n242 B.n115 585
R91 B.n241 B.n240 585
R92 B.n239 B.n118 585
R93 B.n238 B.n237 585
R94 B.n236 B.n119 585
R95 B.n235 B.n234 585
R96 B.n233 B.n120 585
R97 B.n232 B.n231 585
R98 B.n230 B.n121 585
R99 B.n229 B.n228 585
R100 B.n227 B.n122 585
R101 B.n226 B.n225 585
R102 B.n224 B.n123 585
R103 B.n223 B.n222 585
R104 B.n221 B.n124 585
R105 B.n220 B.n219 585
R106 B.n218 B.n125 585
R107 B.n217 B.n216 585
R108 B.n215 B.n126 585
R109 B.n214 B.n213 585
R110 B.n212 B.n127 585
R111 B.n211 B.n210 585
R112 B.n209 B.n128 585
R113 B.n208 B.n207 585
R114 B.n206 B.n129 585
R115 B.n205 B.n204 585
R116 B.n203 B.n130 585
R117 B.n202 B.n201 585
R118 B.n200 B.n131 585
R119 B.n199 B.n198 585
R120 B.n197 B.n132 585
R121 B.n196 B.n195 585
R122 B.n194 B.n133 585
R123 B.n193 B.n192 585
R124 B.n191 B.n134 585
R125 B.n190 B.n189 585
R126 B.n188 B.n135 585
R127 B.n187 B.n186 585
R128 B.n185 B.n136 585
R129 B.n184 B.n183 585
R130 B.n182 B.n137 585
R131 B.n181 B.n180 585
R132 B.n179 B.n138 585
R133 B.n178 B.n177 585
R134 B.n176 B.n139 585
R135 B.n175 B.n174 585
R136 B.n173 B.n140 585
R137 B.n329 B.n84 585
R138 B.n331 B.n330 585
R139 B.n332 B.n83 585
R140 B.n334 B.n333 585
R141 B.n335 B.n82 585
R142 B.n337 B.n336 585
R143 B.n338 B.n81 585
R144 B.n340 B.n339 585
R145 B.n341 B.n80 585
R146 B.n343 B.n342 585
R147 B.n344 B.n79 585
R148 B.n346 B.n345 585
R149 B.n347 B.n78 585
R150 B.n349 B.n348 585
R151 B.n350 B.n77 585
R152 B.n352 B.n351 585
R153 B.n353 B.n76 585
R154 B.n355 B.n354 585
R155 B.n356 B.n75 585
R156 B.n358 B.n357 585
R157 B.n359 B.n74 585
R158 B.n361 B.n360 585
R159 B.n362 B.n73 585
R160 B.n364 B.n363 585
R161 B.n365 B.n72 585
R162 B.n367 B.n366 585
R163 B.n368 B.n71 585
R164 B.n370 B.n369 585
R165 B.n371 B.n70 585
R166 B.n373 B.n372 585
R167 B.n374 B.n69 585
R168 B.n376 B.n375 585
R169 B.n377 B.n68 585
R170 B.n379 B.n378 585
R171 B.n380 B.n67 585
R172 B.n382 B.n381 585
R173 B.n538 B.n537 585
R174 B.n536 B.n11 585
R175 B.n535 B.n534 585
R176 B.n533 B.n12 585
R177 B.n532 B.n531 585
R178 B.n530 B.n13 585
R179 B.n529 B.n528 585
R180 B.n527 B.n14 585
R181 B.n526 B.n525 585
R182 B.n524 B.n15 585
R183 B.n523 B.n522 585
R184 B.n521 B.n16 585
R185 B.n520 B.n519 585
R186 B.n518 B.n17 585
R187 B.n517 B.n516 585
R188 B.n515 B.n18 585
R189 B.n514 B.n513 585
R190 B.n512 B.n19 585
R191 B.n511 B.n510 585
R192 B.n509 B.n20 585
R193 B.n508 B.n507 585
R194 B.n506 B.n21 585
R195 B.n505 B.n504 585
R196 B.n503 B.n22 585
R197 B.n502 B.n501 585
R198 B.n500 B.n23 585
R199 B.n499 B.n498 585
R200 B.n497 B.n24 585
R201 B.n496 B.n495 585
R202 B.n494 B.n25 585
R203 B.n493 B.n492 585
R204 B.n491 B.n26 585
R205 B.n490 B.n489 585
R206 B.n488 B.n27 585
R207 B.n487 B.n486 585
R208 B.n485 B.n28 585
R209 B.n484 B.n483 585
R210 B.n482 B.n29 585
R211 B.n481 B.n480 585
R212 B.n479 B.n30 585
R213 B.n478 B.n477 585
R214 B.n476 B.n31 585
R215 B.n475 B.n474 585
R216 B.n473 B.n32 585
R217 B.n472 B.n471 585
R218 B.n470 B.n33 585
R219 B.n469 B.n468 585
R220 B.n467 B.n466 585
R221 B.n465 B.n37 585
R222 B.n464 B.n463 585
R223 B.n462 B.n38 585
R224 B.n461 B.n460 585
R225 B.n459 B.n39 585
R226 B.n458 B.n457 585
R227 B.n456 B.n40 585
R228 B.n455 B.n454 585
R229 B.n452 B.n41 585
R230 B.n451 B.n450 585
R231 B.n449 B.n44 585
R232 B.n448 B.n447 585
R233 B.n446 B.n45 585
R234 B.n445 B.n444 585
R235 B.n443 B.n46 585
R236 B.n442 B.n441 585
R237 B.n440 B.n47 585
R238 B.n439 B.n438 585
R239 B.n437 B.n48 585
R240 B.n436 B.n435 585
R241 B.n434 B.n49 585
R242 B.n433 B.n432 585
R243 B.n431 B.n50 585
R244 B.n430 B.n429 585
R245 B.n428 B.n51 585
R246 B.n427 B.n426 585
R247 B.n425 B.n52 585
R248 B.n424 B.n423 585
R249 B.n422 B.n53 585
R250 B.n421 B.n420 585
R251 B.n419 B.n54 585
R252 B.n418 B.n417 585
R253 B.n416 B.n55 585
R254 B.n415 B.n414 585
R255 B.n413 B.n56 585
R256 B.n412 B.n411 585
R257 B.n410 B.n57 585
R258 B.n409 B.n408 585
R259 B.n407 B.n58 585
R260 B.n406 B.n405 585
R261 B.n404 B.n59 585
R262 B.n403 B.n402 585
R263 B.n401 B.n60 585
R264 B.n400 B.n399 585
R265 B.n398 B.n61 585
R266 B.n397 B.n396 585
R267 B.n395 B.n62 585
R268 B.n394 B.n393 585
R269 B.n392 B.n63 585
R270 B.n391 B.n390 585
R271 B.n389 B.n64 585
R272 B.n388 B.n387 585
R273 B.n386 B.n65 585
R274 B.n385 B.n384 585
R275 B.n383 B.n66 585
R276 B.n539 B.n10 585
R277 B.n541 B.n540 585
R278 B.n542 B.n9 585
R279 B.n544 B.n543 585
R280 B.n545 B.n8 585
R281 B.n547 B.n546 585
R282 B.n548 B.n7 585
R283 B.n550 B.n549 585
R284 B.n551 B.n6 585
R285 B.n553 B.n552 585
R286 B.n554 B.n5 585
R287 B.n556 B.n555 585
R288 B.n557 B.n4 585
R289 B.n559 B.n558 585
R290 B.n560 B.n3 585
R291 B.n562 B.n561 585
R292 B.n563 B.n0 585
R293 B.n2 B.n1 585
R294 B.n149 B.n148 585
R295 B.n151 B.n150 585
R296 B.n152 B.n147 585
R297 B.n154 B.n153 585
R298 B.n155 B.n146 585
R299 B.n157 B.n156 585
R300 B.n158 B.n145 585
R301 B.n160 B.n159 585
R302 B.n161 B.n144 585
R303 B.n163 B.n162 585
R304 B.n164 B.n143 585
R305 B.n166 B.n165 585
R306 B.n167 B.n142 585
R307 B.n169 B.n168 585
R308 B.n170 B.n141 585
R309 B.n172 B.n171 585
R310 B.n173 B.n172 497.305
R311 B.n329 B.n328 497.305
R312 B.n383 B.n382 497.305
R313 B.n539 B.n538 497.305
R314 B.n565 B.n564 256.663
R315 B.n564 B.n563 235.042
R316 B.n564 B.n2 235.042
R317 B.n174 B.n173 163.367
R318 B.n174 B.n139 163.367
R319 B.n178 B.n139 163.367
R320 B.n179 B.n178 163.367
R321 B.n180 B.n179 163.367
R322 B.n180 B.n137 163.367
R323 B.n184 B.n137 163.367
R324 B.n185 B.n184 163.367
R325 B.n186 B.n185 163.367
R326 B.n186 B.n135 163.367
R327 B.n190 B.n135 163.367
R328 B.n191 B.n190 163.367
R329 B.n192 B.n191 163.367
R330 B.n192 B.n133 163.367
R331 B.n196 B.n133 163.367
R332 B.n197 B.n196 163.367
R333 B.n198 B.n197 163.367
R334 B.n198 B.n131 163.367
R335 B.n202 B.n131 163.367
R336 B.n203 B.n202 163.367
R337 B.n204 B.n203 163.367
R338 B.n204 B.n129 163.367
R339 B.n208 B.n129 163.367
R340 B.n209 B.n208 163.367
R341 B.n210 B.n209 163.367
R342 B.n210 B.n127 163.367
R343 B.n214 B.n127 163.367
R344 B.n215 B.n214 163.367
R345 B.n216 B.n215 163.367
R346 B.n216 B.n125 163.367
R347 B.n220 B.n125 163.367
R348 B.n221 B.n220 163.367
R349 B.n222 B.n221 163.367
R350 B.n222 B.n123 163.367
R351 B.n226 B.n123 163.367
R352 B.n227 B.n226 163.367
R353 B.n228 B.n227 163.367
R354 B.n228 B.n121 163.367
R355 B.n232 B.n121 163.367
R356 B.n233 B.n232 163.367
R357 B.n234 B.n233 163.367
R358 B.n234 B.n119 163.367
R359 B.n238 B.n119 163.367
R360 B.n239 B.n238 163.367
R361 B.n240 B.n239 163.367
R362 B.n240 B.n115 163.367
R363 B.n245 B.n115 163.367
R364 B.n246 B.n245 163.367
R365 B.n247 B.n246 163.367
R366 B.n247 B.n113 163.367
R367 B.n251 B.n113 163.367
R368 B.n252 B.n251 163.367
R369 B.n253 B.n252 163.367
R370 B.n253 B.n111 163.367
R371 B.n257 B.n111 163.367
R372 B.n258 B.n257 163.367
R373 B.n258 B.n107 163.367
R374 B.n262 B.n107 163.367
R375 B.n263 B.n262 163.367
R376 B.n264 B.n263 163.367
R377 B.n264 B.n105 163.367
R378 B.n268 B.n105 163.367
R379 B.n269 B.n268 163.367
R380 B.n270 B.n269 163.367
R381 B.n270 B.n103 163.367
R382 B.n274 B.n103 163.367
R383 B.n275 B.n274 163.367
R384 B.n276 B.n275 163.367
R385 B.n276 B.n101 163.367
R386 B.n280 B.n101 163.367
R387 B.n281 B.n280 163.367
R388 B.n282 B.n281 163.367
R389 B.n282 B.n99 163.367
R390 B.n286 B.n99 163.367
R391 B.n287 B.n286 163.367
R392 B.n288 B.n287 163.367
R393 B.n288 B.n97 163.367
R394 B.n292 B.n97 163.367
R395 B.n293 B.n292 163.367
R396 B.n294 B.n293 163.367
R397 B.n294 B.n95 163.367
R398 B.n298 B.n95 163.367
R399 B.n299 B.n298 163.367
R400 B.n300 B.n299 163.367
R401 B.n300 B.n93 163.367
R402 B.n304 B.n93 163.367
R403 B.n305 B.n304 163.367
R404 B.n306 B.n305 163.367
R405 B.n306 B.n91 163.367
R406 B.n310 B.n91 163.367
R407 B.n311 B.n310 163.367
R408 B.n312 B.n311 163.367
R409 B.n312 B.n89 163.367
R410 B.n316 B.n89 163.367
R411 B.n317 B.n316 163.367
R412 B.n318 B.n317 163.367
R413 B.n318 B.n87 163.367
R414 B.n322 B.n87 163.367
R415 B.n323 B.n322 163.367
R416 B.n324 B.n323 163.367
R417 B.n324 B.n85 163.367
R418 B.n328 B.n85 163.367
R419 B.n382 B.n67 163.367
R420 B.n378 B.n67 163.367
R421 B.n378 B.n377 163.367
R422 B.n377 B.n376 163.367
R423 B.n376 B.n69 163.367
R424 B.n372 B.n69 163.367
R425 B.n372 B.n371 163.367
R426 B.n371 B.n370 163.367
R427 B.n370 B.n71 163.367
R428 B.n366 B.n71 163.367
R429 B.n366 B.n365 163.367
R430 B.n365 B.n364 163.367
R431 B.n364 B.n73 163.367
R432 B.n360 B.n73 163.367
R433 B.n360 B.n359 163.367
R434 B.n359 B.n358 163.367
R435 B.n358 B.n75 163.367
R436 B.n354 B.n75 163.367
R437 B.n354 B.n353 163.367
R438 B.n353 B.n352 163.367
R439 B.n352 B.n77 163.367
R440 B.n348 B.n77 163.367
R441 B.n348 B.n347 163.367
R442 B.n347 B.n346 163.367
R443 B.n346 B.n79 163.367
R444 B.n342 B.n79 163.367
R445 B.n342 B.n341 163.367
R446 B.n341 B.n340 163.367
R447 B.n340 B.n81 163.367
R448 B.n336 B.n81 163.367
R449 B.n336 B.n335 163.367
R450 B.n335 B.n334 163.367
R451 B.n334 B.n83 163.367
R452 B.n330 B.n83 163.367
R453 B.n330 B.n329 163.367
R454 B.n538 B.n11 163.367
R455 B.n534 B.n11 163.367
R456 B.n534 B.n533 163.367
R457 B.n533 B.n532 163.367
R458 B.n532 B.n13 163.367
R459 B.n528 B.n13 163.367
R460 B.n528 B.n527 163.367
R461 B.n527 B.n526 163.367
R462 B.n526 B.n15 163.367
R463 B.n522 B.n15 163.367
R464 B.n522 B.n521 163.367
R465 B.n521 B.n520 163.367
R466 B.n520 B.n17 163.367
R467 B.n516 B.n17 163.367
R468 B.n516 B.n515 163.367
R469 B.n515 B.n514 163.367
R470 B.n514 B.n19 163.367
R471 B.n510 B.n19 163.367
R472 B.n510 B.n509 163.367
R473 B.n509 B.n508 163.367
R474 B.n508 B.n21 163.367
R475 B.n504 B.n21 163.367
R476 B.n504 B.n503 163.367
R477 B.n503 B.n502 163.367
R478 B.n502 B.n23 163.367
R479 B.n498 B.n23 163.367
R480 B.n498 B.n497 163.367
R481 B.n497 B.n496 163.367
R482 B.n496 B.n25 163.367
R483 B.n492 B.n25 163.367
R484 B.n492 B.n491 163.367
R485 B.n491 B.n490 163.367
R486 B.n490 B.n27 163.367
R487 B.n486 B.n27 163.367
R488 B.n486 B.n485 163.367
R489 B.n485 B.n484 163.367
R490 B.n484 B.n29 163.367
R491 B.n480 B.n29 163.367
R492 B.n480 B.n479 163.367
R493 B.n479 B.n478 163.367
R494 B.n478 B.n31 163.367
R495 B.n474 B.n31 163.367
R496 B.n474 B.n473 163.367
R497 B.n473 B.n472 163.367
R498 B.n472 B.n33 163.367
R499 B.n468 B.n33 163.367
R500 B.n468 B.n467 163.367
R501 B.n467 B.n37 163.367
R502 B.n463 B.n37 163.367
R503 B.n463 B.n462 163.367
R504 B.n462 B.n461 163.367
R505 B.n461 B.n39 163.367
R506 B.n457 B.n39 163.367
R507 B.n457 B.n456 163.367
R508 B.n456 B.n455 163.367
R509 B.n455 B.n41 163.367
R510 B.n450 B.n41 163.367
R511 B.n450 B.n449 163.367
R512 B.n449 B.n448 163.367
R513 B.n448 B.n45 163.367
R514 B.n444 B.n45 163.367
R515 B.n444 B.n443 163.367
R516 B.n443 B.n442 163.367
R517 B.n442 B.n47 163.367
R518 B.n438 B.n47 163.367
R519 B.n438 B.n437 163.367
R520 B.n437 B.n436 163.367
R521 B.n436 B.n49 163.367
R522 B.n432 B.n49 163.367
R523 B.n432 B.n431 163.367
R524 B.n431 B.n430 163.367
R525 B.n430 B.n51 163.367
R526 B.n426 B.n51 163.367
R527 B.n426 B.n425 163.367
R528 B.n425 B.n424 163.367
R529 B.n424 B.n53 163.367
R530 B.n420 B.n53 163.367
R531 B.n420 B.n419 163.367
R532 B.n419 B.n418 163.367
R533 B.n418 B.n55 163.367
R534 B.n414 B.n55 163.367
R535 B.n414 B.n413 163.367
R536 B.n413 B.n412 163.367
R537 B.n412 B.n57 163.367
R538 B.n408 B.n57 163.367
R539 B.n408 B.n407 163.367
R540 B.n407 B.n406 163.367
R541 B.n406 B.n59 163.367
R542 B.n402 B.n59 163.367
R543 B.n402 B.n401 163.367
R544 B.n401 B.n400 163.367
R545 B.n400 B.n61 163.367
R546 B.n396 B.n61 163.367
R547 B.n396 B.n395 163.367
R548 B.n395 B.n394 163.367
R549 B.n394 B.n63 163.367
R550 B.n390 B.n63 163.367
R551 B.n390 B.n389 163.367
R552 B.n389 B.n388 163.367
R553 B.n388 B.n65 163.367
R554 B.n384 B.n65 163.367
R555 B.n384 B.n383 163.367
R556 B.n540 B.n539 163.367
R557 B.n540 B.n9 163.367
R558 B.n544 B.n9 163.367
R559 B.n545 B.n544 163.367
R560 B.n546 B.n545 163.367
R561 B.n546 B.n7 163.367
R562 B.n550 B.n7 163.367
R563 B.n551 B.n550 163.367
R564 B.n552 B.n551 163.367
R565 B.n552 B.n5 163.367
R566 B.n556 B.n5 163.367
R567 B.n557 B.n556 163.367
R568 B.n558 B.n557 163.367
R569 B.n558 B.n3 163.367
R570 B.n562 B.n3 163.367
R571 B.n563 B.n562 163.367
R572 B.n149 B.n2 163.367
R573 B.n150 B.n149 163.367
R574 B.n150 B.n147 163.367
R575 B.n154 B.n147 163.367
R576 B.n155 B.n154 163.367
R577 B.n156 B.n155 163.367
R578 B.n156 B.n145 163.367
R579 B.n160 B.n145 163.367
R580 B.n161 B.n160 163.367
R581 B.n162 B.n161 163.367
R582 B.n162 B.n143 163.367
R583 B.n166 B.n143 163.367
R584 B.n167 B.n166 163.367
R585 B.n168 B.n167 163.367
R586 B.n168 B.n141 163.367
R587 B.n172 B.n141 163.367
R588 B.n108 B.t4 129.267
R589 B.n42 B.t11 129.267
R590 B.n116 B.t1 129.25
R591 B.n34 B.t8 129.25
R592 B.n109 B.t5 108.32
R593 B.n43 B.t10 108.32
R594 B.n117 B.t2 108.303
R595 B.n35 B.t7 108.303
R596 B.n243 B.n117 59.5399
R597 B.n110 B.n109 59.5399
R598 B.n453 B.n43 59.5399
R599 B.n36 B.n35 59.5399
R600 B.n537 B.n10 32.3127
R601 B.n381 B.n66 32.3127
R602 B.n327 B.n84 32.3127
R603 B.n171 B.n140 32.3127
R604 B.n117 B.n116 20.946
R605 B.n109 B.n108 20.946
R606 B.n43 B.n42 20.946
R607 B.n35 B.n34 20.946
R608 B B.n565 18.0485
R609 B.n541 B.n10 10.6151
R610 B.n542 B.n541 10.6151
R611 B.n543 B.n542 10.6151
R612 B.n543 B.n8 10.6151
R613 B.n547 B.n8 10.6151
R614 B.n548 B.n547 10.6151
R615 B.n549 B.n548 10.6151
R616 B.n549 B.n6 10.6151
R617 B.n553 B.n6 10.6151
R618 B.n554 B.n553 10.6151
R619 B.n555 B.n554 10.6151
R620 B.n555 B.n4 10.6151
R621 B.n559 B.n4 10.6151
R622 B.n560 B.n559 10.6151
R623 B.n561 B.n560 10.6151
R624 B.n561 B.n0 10.6151
R625 B.n537 B.n536 10.6151
R626 B.n536 B.n535 10.6151
R627 B.n535 B.n12 10.6151
R628 B.n531 B.n12 10.6151
R629 B.n531 B.n530 10.6151
R630 B.n530 B.n529 10.6151
R631 B.n529 B.n14 10.6151
R632 B.n525 B.n14 10.6151
R633 B.n525 B.n524 10.6151
R634 B.n524 B.n523 10.6151
R635 B.n523 B.n16 10.6151
R636 B.n519 B.n16 10.6151
R637 B.n519 B.n518 10.6151
R638 B.n518 B.n517 10.6151
R639 B.n517 B.n18 10.6151
R640 B.n513 B.n18 10.6151
R641 B.n513 B.n512 10.6151
R642 B.n512 B.n511 10.6151
R643 B.n511 B.n20 10.6151
R644 B.n507 B.n20 10.6151
R645 B.n507 B.n506 10.6151
R646 B.n506 B.n505 10.6151
R647 B.n505 B.n22 10.6151
R648 B.n501 B.n22 10.6151
R649 B.n501 B.n500 10.6151
R650 B.n500 B.n499 10.6151
R651 B.n499 B.n24 10.6151
R652 B.n495 B.n24 10.6151
R653 B.n495 B.n494 10.6151
R654 B.n494 B.n493 10.6151
R655 B.n493 B.n26 10.6151
R656 B.n489 B.n26 10.6151
R657 B.n489 B.n488 10.6151
R658 B.n488 B.n487 10.6151
R659 B.n487 B.n28 10.6151
R660 B.n483 B.n28 10.6151
R661 B.n483 B.n482 10.6151
R662 B.n482 B.n481 10.6151
R663 B.n481 B.n30 10.6151
R664 B.n477 B.n30 10.6151
R665 B.n477 B.n476 10.6151
R666 B.n476 B.n475 10.6151
R667 B.n475 B.n32 10.6151
R668 B.n471 B.n32 10.6151
R669 B.n471 B.n470 10.6151
R670 B.n470 B.n469 10.6151
R671 B.n466 B.n465 10.6151
R672 B.n465 B.n464 10.6151
R673 B.n464 B.n38 10.6151
R674 B.n460 B.n38 10.6151
R675 B.n460 B.n459 10.6151
R676 B.n459 B.n458 10.6151
R677 B.n458 B.n40 10.6151
R678 B.n454 B.n40 10.6151
R679 B.n452 B.n451 10.6151
R680 B.n451 B.n44 10.6151
R681 B.n447 B.n44 10.6151
R682 B.n447 B.n446 10.6151
R683 B.n446 B.n445 10.6151
R684 B.n445 B.n46 10.6151
R685 B.n441 B.n46 10.6151
R686 B.n441 B.n440 10.6151
R687 B.n440 B.n439 10.6151
R688 B.n439 B.n48 10.6151
R689 B.n435 B.n48 10.6151
R690 B.n435 B.n434 10.6151
R691 B.n434 B.n433 10.6151
R692 B.n433 B.n50 10.6151
R693 B.n429 B.n50 10.6151
R694 B.n429 B.n428 10.6151
R695 B.n428 B.n427 10.6151
R696 B.n427 B.n52 10.6151
R697 B.n423 B.n52 10.6151
R698 B.n423 B.n422 10.6151
R699 B.n422 B.n421 10.6151
R700 B.n421 B.n54 10.6151
R701 B.n417 B.n54 10.6151
R702 B.n417 B.n416 10.6151
R703 B.n416 B.n415 10.6151
R704 B.n415 B.n56 10.6151
R705 B.n411 B.n56 10.6151
R706 B.n411 B.n410 10.6151
R707 B.n410 B.n409 10.6151
R708 B.n409 B.n58 10.6151
R709 B.n405 B.n58 10.6151
R710 B.n405 B.n404 10.6151
R711 B.n404 B.n403 10.6151
R712 B.n403 B.n60 10.6151
R713 B.n399 B.n60 10.6151
R714 B.n399 B.n398 10.6151
R715 B.n398 B.n397 10.6151
R716 B.n397 B.n62 10.6151
R717 B.n393 B.n62 10.6151
R718 B.n393 B.n392 10.6151
R719 B.n392 B.n391 10.6151
R720 B.n391 B.n64 10.6151
R721 B.n387 B.n64 10.6151
R722 B.n387 B.n386 10.6151
R723 B.n386 B.n385 10.6151
R724 B.n385 B.n66 10.6151
R725 B.n381 B.n380 10.6151
R726 B.n380 B.n379 10.6151
R727 B.n379 B.n68 10.6151
R728 B.n375 B.n68 10.6151
R729 B.n375 B.n374 10.6151
R730 B.n374 B.n373 10.6151
R731 B.n373 B.n70 10.6151
R732 B.n369 B.n70 10.6151
R733 B.n369 B.n368 10.6151
R734 B.n368 B.n367 10.6151
R735 B.n367 B.n72 10.6151
R736 B.n363 B.n72 10.6151
R737 B.n363 B.n362 10.6151
R738 B.n362 B.n361 10.6151
R739 B.n361 B.n74 10.6151
R740 B.n357 B.n74 10.6151
R741 B.n357 B.n356 10.6151
R742 B.n356 B.n355 10.6151
R743 B.n355 B.n76 10.6151
R744 B.n351 B.n76 10.6151
R745 B.n351 B.n350 10.6151
R746 B.n350 B.n349 10.6151
R747 B.n349 B.n78 10.6151
R748 B.n345 B.n78 10.6151
R749 B.n345 B.n344 10.6151
R750 B.n344 B.n343 10.6151
R751 B.n343 B.n80 10.6151
R752 B.n339 B.n80 10.6151
R753 B.n339 B.n338 10.6151
R754 B.n338 B.n337 10.6151
R755 B.n337 B.n82 10.6151
R756 B.n333 B.n82 10.6151
R757 B.n333 B.n332 10.6151
R758 B.n332 B.n331 10.6151
R759 B.n331 B.n84 10.6151
R760 B.n148 B.n1 10.6151
R761 B.n151 B.n148 10.6151
R762 B.n152 B.n151 10.6151
R763 B.n153 B.n152 10.6151
R764 B.n153 B.n146 10.6151
R765 B.n157 B.n146 10.6151
R766 B.n158 B.n157 10.6151
R767 B.n159 B.n158 10.6151
R768 B.n159 B.n144 10.6151
R769 B.n163 B.n144 10.6151
R770 B.n164 B.n163 10.6151
R771 B.n165 B.n164 10.6151
R772 B.n165 B.n142 10.6151
R773 B.n169 B.n142 10.6151
R774 B.n170 B.n169 10.6151
R775 B.n171 B.n170 10.6151
R776 B.n175 B.n140 10.6151
R777 B.n176 B.n175 10.6151
R778 B.n177 B.n176 10.6151
R779 B.n177 B.n138 10.6151
R780 B.n181 B.n138 10.6151
R781 B.n182 B.n181 10.6151
R782 B.n183 B.n182 10.6151
R783 B.n183 B.n136 10.6151
R784 B.n187 B.n136 10.6151
R785 B.n188 B.n187 10.6151
R786 B.n189 B.n188 10.6151
R787 B.n189 B.n134 10.6151
R788 B.n193 B.n134 10.6151
R789 B.n194 B.n193 10.6151
R790 B.n195 B.n194 10.6151
R791 B.n195 B.n132 10.6151
R792 B.n199 B.n132 10.6151
R793 B.n200 B.n199 10.6151
R794 B.n201 B.n200 10.6151
R795 B.n201 B.n130 10.6151
R796 B.n205 B.n130 10.6151
R797 B.n206 B.n205 10.6151
R798 B.n207 B.n206 10.6151
R799 B.n207 B.n128 10.6151
R800 B.n211 B.n128 10.6151
R801 B.n212 B.n211 10.6151
R802 B.n213 B.n212 10.6151
R803 B.n213 B.n126 10.6151
R804 B.n217 B.n126 10.6151
R805 B.n218 B.n217 10.6151
R806 B.n219 B.n218 10.6151
R807 B.n219 B.n124 10.6151
R808 B.n223 B.n124 10.6151
R809 B.n224 B.n223 10.6151
R810 B.n225 B.n224 10.6151
R811 B.n225 B.n122 10.6151
R812 B.n229 B.n122 10.6151
R813 B.n230 B.n229 10.6151
R814 B.n231 B.n230 10.6151
R815 B.n231 B.n120 10.6151
R816 B.n235 B.n120 10.6151
R817 B.n236 B.n235 10.6151
R818 B.n237 B.n236 10.6151
R819 B.n237 B.n118 10.6151
R820 B.n241 B.n118 10.6151
R821 B.n242 B.n241 10.6151
R822 B.n244 B.n114 10.6151
R823 B.n248 B.n114 10.6151
R824 B.n249 B.n248 10.6151
R825 B.n250 B.n249 10.6151
R826 B.n250 B.n112 10.6151
R827 B.n254 B.n112 10.6151
R828 B.n255 B.n254 10.6151
R829 B.n256 B.n255 10.6151
R830 B.n260 B.n259 10.6151
R831 B.n261 B.n260 10.6151
R832 B.n261 B.n106 10.6151
R833 B.n265 B.n106 10.6151
R834 B.n266 B.n265 10.6151
R835 B.n267 B.n266 10.6151
R836 B.n267 B.n104 10.6151
R837 B.n271 B.n104 10.6151
R838 B.n272 B.n271 10.6151
R839 B.n273 B.n272 10.6151
R840 B.n273 B.n102 10.6151
R841 B.n277 B.n102 10.6151
R842 B.n278 B.n277 10.6151
R843 B.n279 B.n278 10.6151
R844 B.n279 B.n100 10.6151
R845 B.n283 B.n100 10.6151
R846 B.n284 B.n283 10.6151
R847 B.n285 B.n284 10.6151
R848 B.n285 B.n98 10.6151
R849 B.n289 B.n98 10.6151
R850 B.n290 B.n289 10.6151
R851 B.n291 B.n290 10.6151
R852 B.n291 B.n96 10.6151
R853 B.n295 B.n96 10.6151
R854 B.n296 B.n295 10.6151
R855 B.n297 B.n296 10.6151
R856 B.n297 B.n94 10.6151
R857 B.n301 B.n94 10.6151
R858 B.n302 B.n301 10.6151
R859 B.n303 B.n302 10.6151
R860 B.n303 B.n92 10.6151
R861 B.n307 B.n92 10.6151
R862 B.n308 B.n307 10.6151
R863 B.n309 B.n308 10.6151
R864 B.n309 B.n90 10.6151
R865 B.n313 B.n90 10.6151
R866 B.n314 B.n313 10.6151
R867 B.n315 B.n314 10.6151
R868 B.n315 B.n88 10.6151
R869 B.n319 B.n88 10.6151
R870 B.n320 B.n319 10.6151
R871 B.n321 B.n320 10.6151
R872 B.n321 B.n86 10.6151
R873 B.n325 B.n86 10.6151
R874 B.n326 B.n325 10.6151
R875 B.n327 B.n326 10.6151
R876 B.n565 B.n0 8.11757
R877 B.n565 B.n1 8.11757
R878 B.n466 B.n36 6.5566
R879 B.n454 B.n453 6.5566
R880 B.n244 B.n243 6.5566
R881 B.n256 B.n110 6.5566
R882 B.n469 B.n36 4.05904
R883 B.n453 B.n452 4.05904
R884 B.n243 B.n242 4.05904
R885 B.n259 B.n110 4.05904
R886 VP.n1 VP.t1 512.958
R887 VP.n1 VP.t0 512.909
R888 VP.n3 VP.t2 491.962
R889 VP.n5 VP.t3 491.962
R890 VP.n6 VP.n5 161.3
R891 VP.n4 VP.n0 161.3
R892 VP.n3 VP.n2 161.3
R893 VP.n2 VP.n1 86.5333
R894 VP.n4 VP.n3 24.1005
R895 VP.n5 VP.n4 24.1005
R896 VP.n2 VP.n0 0.189894
R897 VP.n6 VP.n0 0.189894
R898 VP VP.n6 0.0516364
R899 VDD1 VDD1.n1 112.796
R900 VDD1 VDD1.n0 74.0283
R901 VDD1.n0 VDD1.t2 2.3766
R902 VDD1.n0 VDD1.t3 2.3766
R903 VDD1.n1 VDD1.t1 2.3766
R904 VDD1.n1 VDD1.t0 2.3766
C0 B w_n1618_n3704# 7.44017f
C1 B VDD2 1.00247f
C2 w_n1618_n3704# VN 2.43101f
C3 B VDD1 0.980232f
C4 VN VDD2 3.67661f
C5 B VTAIL 4.31326f
C6 VN VDD1 0.147469f
C7 VN VTAIL 3.22611f
C8 w_n1618_n3704# VP 2.63433f
C9 VP VDD2 0.276727f
C10 VP VDD1 3.8056f
C11 VTAIL VP 3.24022f
C12 B VN 0.778027f
C13 w_n1618_n3704# VDD2 1.13278f
C14 w_n1618_n3704# VDD1 1.11725f
C15 w_n1618_n3704# VTAIL 4.53509f
C16 VDD1 VDD2 0.577924f
C17 VTAIL VDD2 7.38701f
C18 B VP 1.10682f
C19 VTAIL VDD1 7.345201f
C20 VN VP 5.16703f
C21 VDD2 VSUBS 0.723633f
C22 VDD1 VSUBS 5.172149f
C23 VTAIL VSUBS 0.965182f
C24 VN VSUBS 5.88221f
C25 VP VSUBS 1.379848f
C26 B VSUBS 2.804844f
C27 w_n1618_n3704# VSUBS 73.6061f
C28 VDD1.t2 VSUBS 0.301188f
C29 VDD1.t3 VSUBS 0.301188f
C30 VDD1.n0 VSUBS 2.42139f
C31 VDD1.t1 VSUBS 0.301188f
C32 VDD1.t0 VSUBS 0.301188f
C33 VDD1.n1 VSUBS 3.13305f
C34 VP.n0 VSUBS 0.059227f
C35 VP.t0 VSUBS 1.75664f
C36 VP.t1 VSUBS 1.75672f
C37 VP.n1 VSUBS 2.5387f
C38 VP.n2 VSUBS 3.80561f
C39 VP.t2 VSUBS 1.7291f
C40 VP.n3 VSUBS 0.670092f
C41 VP.n4 VSUBS 0.01344f
C42 VP.t3 VSUBS 1.7291f
C43 VP.n5 VSUBS 0.670092f
C44 VP.n6 VSUBS 0.045898f
C45 B.n0 VSUBS 0.007009f
C46 B.n1 VSUBS 0.007009f
C47 B.n2 VSUBS 0.010366f
C48 B.n3 VSUBS 0.007944f
C49 B.n4 VSUBS 0.007944f
C50 B.n5 VSUBS 0.007944f
C51 B.n6 VSUBS 0.007944f
C52 B.n7 VSUBS 0.007944f
C53 B.n8 VSUBS 0.007944f
C54 B.n9 VSUBS 0.007944f
C55 B.n10 VSUBS 0.017775f
C56 B.n11 VSUBS 0.007944f
C57 B.n12 VSUBS 0.007944f
C58 B.n13 VSUBS 0.007944f
C59 B.n14 VSUBS 0.007944f
C60 B.n15 VSUBS 0.007944f
C61 B.n16 VSUBS 0.007944f
C62 B.n17 VSUBS 0.007944f
C63 B.n18 VSUBS 0.007944f
C64 B.n19 VSUBS 0.007944f
C65 B.n20 VSUBS 0.007944f
C66 B.n21 VSUBS 0.007944f
C67 B.n22 VSUBS 0.007944f
C68 B.n23 VSUBS 0.007944f
C69 B.n24 VSUBS 0.007944f
C70 B.n25 VSUBS 0.007944f
C71 B.n26 VSUBS 0.007944f
C72 B.n27 VSUBS 0.007944f
C73 B.n28 VSUBS 0.007944f
C74 B.n29 VSUBS 0.007944f
C75 B.n30 VSUBS 0.007944f
C76 B.n31 VSUBS 0.007944f
C77 B.n32 VSUBS 0.007944f
C78 B.n33 VSUBS 0.007944f
C79 B.t7 VSUBS 0.512592f
C80 B.t8 VSUBS 0.522573f
C81 B.t6 VSUBS 0.478674f
C82 B.n34 VSUBS 0.17398f
C83 B.n35 VSUBS 0.072918f
C84 B.n36 VSUBS 0.018405f
C85 B.n37 VSUBS 0.007944f
C86 B.n38 VSUBS 0.007944f
C87 B.n39 VSUBS 0.007944f
C88 B.n40 VSUBS 0.007944f
C89 B.n41 VSUBS 0.007944f
C90 B.t10 VSUBS 0.512579f
C91 B.t11 VSUBS 0.522561f
C92 B.t9 VSUBS 0.478674f
C93 B.n42 VSUBS 0.173992f
C94 B.n43 VSUBS 0.072931f
C95 B.n44 VSUBS 0.007944f
C96 B.n45 VSUBS 0.007944f
C97 B.n46 VSUBS 0.007944f
C98 B.n47 VSUBS 0.007944f
C99 B.n48 VSUBS 0.007944f
C100 B.n49 VSUBS 0.007944f
C101 B.n50 VSUBS 0.007944f
C102 B.n51 VSUBS 0.007944f
C103 B.n52 VSUBS 0.007944f
C104 B.n53 VSUBS 0.007944f
C105 B.n54 VSUBS 0.007944f
C106 B.n55 VSUBS 0.007944f
C107 B.n56 VSUBS 0.007944f
C108 B.n57 VSUBS 0.007944f
C109 B.n58 VSUBS 0.007944f
C110 B.n59 VSUBS 0.007944f
C111 B.n60 VSUBS 0.007944f
C112 B.n61 VSUBS 0.007944f
C113 B.n62 VSUBS 0.007944f
C114 B.n63 VSUBS 0.007944f
C115 B.n64 VSUBS 0.007944f
C116 B.n65 VSUBS 0.007944f
C117 B.n66 VSUBS 0.019141f
C118 B.n67 VSUBS 0.007944f
C119 B.n68 VSUBS 0.007944f
C120 B.n69 VSUBS 0.007944f
C121 B.n70 VSUBS 0.007944f
C122 B.n71 VSUBS 0.007944f
C123 B.n72 VSUBS 0.007944f
C124 B.n73 VSUBS 0.007944f
C125 B.n74 VSUBS 0.007944f
C126 B.n75 VSUBS 0.007944f
C127 B.n76 VSUBS 0.007944f
C128 B.n77 VSUBS 0.007944f
C129 B.n78 VSUBS 0.007944f
C130 B.n79 VSUBS 0.007944f
C131 B.n80 VSUBS 0.007944f
C132 B.n81 VSUBS 0.007944f
C133 B.n82 VSUBS 0.007944f
C134 B.n83 VSUBS 0.007944f
C135 B.n84 VSUBS 0.018724f
C136 B.n85 VSUBS 0.007944f
C137 B.n86 VSUBS 0.007944f
C138 B.n87 VSUBS 0.007944f
C139 B.n88 VSUBS 0.007944f
C140 B.n89 VSUBS 0.007944f
C141 B.n90 VSUBS 0.007944f
C142 B.n91 VSUBS 0.007944f
C143 B.n92 VSUBS 0.007944f
C144 B.n93 VSUBS 0.007944f
C145 B.n94 VSUBS 0.007944f
C146 B.n95 VSUBS 0.007944f
C147 B.n96 VSUBS 0.007944f
C148 B.n97 VSUBS 0.007944f
C149 B.n98 VSUBS 0.007944f
C150 B.n99 VSUBS 0.007944f
C151 B.n100 VSUBS 0.007944f
C152 B.n101 VSUBS 0.007944f
C153 B.n102 VSUBS 0.007944f
C154 B.n103 VSUBS 0.007944f
C155 B.n104 VSUBS 0.007944f
C156 B.n105 VSUBS 0.007944f
C157 B.n106 VSUBS 0.007944f
C158 B.n107 VSUBS 0.007944f
C159 B.t5 VSUBS 0.512579f
C160 B.t4 VSUBS 0.522561f
C161 B.t3 VSUBS 0.478674f
C162 B.n108 VSUBS 0.173992f
C163 B.n109 VSUBS 0.072931f
C164 B.n110 VSUBS 0.018405f
C165 B.n111 VSUBS 0.007944f
C166 B.n112 VSUBS 0.007944f
C167 B.n113 VSUBS 0.007944f
C168 B.n114 VSUBS 0.007944f
C169 B.n115 VSUBS 0.007944f
C170 B.t2 VSUBS 0.512592f
C171 B.t1 VSUBS 0.522573f
C172 B.t0 VSUBS 0.478674f
C173 B.n116 VSUBS 0.17398f
C174 B.n117 VSUBS 0.072918f
C175 B.n118 VSUBS 0.007944f
C176 B.n119 VSUBS 0.007944f
C177 B.n120 VSUBS 0.007944f
C178 B.n121 VSUBS 0.007944f
C179 B.n122 VSUBS 0.007944f
C180 B.n123 VSUBS 0.007944f
C181 B.n124 VSUBS 0.007944f
C182 B.n125 VSUBS 0.007944f
C183 B.n126 VSUBS 0.007944f
C184 B.n127 VSUBS 0.007944f
C185 B.n128 VSUBS 0.007944f
C186 B.n129 VSUBS 0.007944f
C187 B.n130 VSUBS 0.007944f
C188 B.n131 VSUBS 0.007944f
C189 B.n132 VSUBS 0.007944f
C190 B.n133 VSUBS 0.007944f
C191 B.n134 VSUBS 0.007944f
C192 B.n135 VSUBS 0.007944f
C193 B.n136 VSUBS 0.007944f
C194 B.n137 VSUBS 0.007944f
C195 B.n138 VSUBS 0.007944f
C196 B.n139 VSUBS 0.007944f
C197 B.n140 VSUBS 0.019141f
C198 B.n141 VSUBS 0.007944f
C199 B.n142 VSUBS 0.007944f
C200 B.n143 VSUBS 0.007944f
C201 B.n144 VSUBS 0.007944f
C202 B.n145 VSUBS 0.007944f
C203 B.n146 VSUBS 0.007944f
C204 B.n147 VSUBS 0.007944f
C205 B.n148 VSUBS 0.007944f
C206 B.n149 VSUBS 0.007944f
C207 B.n150 VSUBS 0.007944f
C208 B.n151 VSUBS 0.007944f
C209 B.n152 VSUBS 0.007944f
C210 B.n153 VSUBS 0.007944f
C211 B.n154 VSUBS 0.007944f
C212 B.n155 VSUBS 0.007944f
C213 B.n156 VSUBS 0.007944f
C214 B.n157 VSUBS 0.007944f
C215 B.n158 VSUBS 0.007944f
C216 B.n159 VSUBS 0.007944f
C217 B.n160 VSUBS 0.007944f
C218 B.n161 VSUBS 0.007944f
C219 B.n162 VSUBS 0.007944f
C220 B.n163 VSUBS 0.007944f
C221 B.n164 VSUBS 0.007944f
C222 B.n165 VSUBS 0.007944f
C223 B.n166 VSUBS 0.007944f
C224 B.n167 VSUBS 0.007944f
C225 B.n168 VSUBS 0.007944f
C226 B.n169 VSUBS 0.007944f
C227 B.n170 VSUBS 0.007944f
C228 B.n171 VSUBS 0.017775f
C229 B.n172 VSUBS 0.017775f
C230 B.n173 VSUBS 0.019141f
C231 B.n174 VSUBS 0.007944f
C232 B.n175 VSUBS 0.007944f
C233 B.n176 VSUBS 0.007944f
C234 B.n177 VSUBS 0.007944f
C235 B.n178 VSUBS 0.007944f
C236 B.n179 VSUBS 0.007944f
C237 B.n180 VSUBS 0.007944f
C238 B.n181 VSUBS 0.007944f
C239 B.n182 VSUBS 0.007944f
C240 B.n183 VSUBS 0.007944f
C241 B.n184 VSUBS 0.007944f
C242 B.n185 VSUBS 0.007944f
C243 B.n186 VSUBS 0.007944f
C244 B.n187 VSUBS 0.007944f
C245 B.n188 VSUBS 0.007944f
C246 B.n189 VSUBS 0.007944f
C247 B.n190 VSUBS 0.007944f
C248 B.n191 VSUBS 0.007944f
C249 B.n192 VSUBS 0.007944f
C250 B.n193 VSUBS 0.007944f
C251 B.n194 VSUBS 0.007944f
C252 B.n195 VSUBS 0.007944f
C253 B.n196 VSUBS 0.007944f
C254 B.n197 VSUBS 0.007944f
C255 B.n198 VSUBS 0.007944f
C256 B.n199 VSUBS 0.007944f
C257 B.n200 VSUBS 0.007944f
C258 B.n201 VSUBS 0.007944f
C259 B.n202 VSUBS 0.007944f
C260 B.n203 VSUBS 0.007944f
C261 B.n204 VSUBS 0.007944f
C262 B.n205 VSUBS 0.007944f
C263 B.n206 VSUBS 0.007944f
C264 B.n207 VSUBS 0.007944f
C265 B.n208 VSUBS 0.007944f
C266 B.n209 VSUBS 0.007944f
C267 B.n210 VSUBS 0.007944f
C268 B.n211 VSUBS 0.007944f
C269 B.n212 VSUBS 0.007944f
C270 B.n213 VSUBS 0.007944f
C271 B.n214 VSUBS 0.007944f
C272 B.n215 VSUBS 0.007944f
C273 B.n216 VSUBS 0.007944f
C274 B.n217 VSUBS 0.007944f
C275 B.n218 VSUBS 0.007944f
C276 B.n219 VSUBS 0.007944f
C277 B.n220 VSUBS 0.007944f
C278 B.n221 VSUBS 0.007944f
C279 B.n222 VSUBS 0.007944f
C280 B.n223 VSUBS 0.007944f
C281 B.n224 VSUBS 0.007944f
C282 B.n225 VSUBS 0.007944f
C283 B.n226 VSUBS 0.007944f
C284 B.n227 VSUBS 0.007944f
C285 B.n228 VSUBS 0.007944f
C286 B.n229 VSUBS 0.007944f
C287 B.n230 VSUBS 0.007944f
C288 B.n231 VSUBS 0.007944f
C289 B.n232 VSUBS 0.007944f
C290 B.n233 VSUBS 0.007944f
C291 B.n234 VSUBS 0.007944f
C292 B.n235 VSUBS 0.007944f
C293 B.n236 VSUBS 0.007944f
C294 B.n237 VSUBS 0.007944f
C295 B.n238 VSUBS 0.007944f
C296 B.n239 VSUBS 0.007944f
C297 B.n240 VSUBS 0.007944f
C298 B.n241 VSUBS 0.007944f
C299 B.n242 VSUBS 0.005491f
C300 B.n243 VSUBS 0.018405f
C301 B.n244 VSUBS 0.006425f
C302 B.n245 VSUBS 0.007944f
C303 B.n246 VSUBS 0.007944f
C304 B.n247 VSUBS 0.007944f
C305 B.n248 VSUBS 0.007944f
C306 B.n249 VSUBS 0.007944f
C307 B.n250 VSUBS 0.007944f
C308 B.n251 VSUBS 0.007944f
C309 B.n252 VSUBS 0.007944f
C310 B.n253 VSUBS 0.007944f
C311 B.n254 VSUBS 0.007944f
C312 B.n255 VSUBS 0.007944f
C313 B.n256 VSUBS 0.006425f
C314 B.n257 VSUBS 0.007944f
C315 B.n258 VSUBS 0.007944f
C316 B.n259 VSUBS 0.005491f
C317 B.n260 VSUBS 0.007944f
C318 B.n261 VSUBS 0.007944f
C319 B.n262 VSUBS 0.007944f
C320 B.n263 VSUBS 0.007944f
C321 B.n264 VSUBS 0.007944f
C322 B.n265 VSUBS 0.007944f
C323 B.n266 VSUBS 0.007944f
C324 B.n267 VSUBS 0.007944f
C325 B.n268 VSUBS 0.007944f
C326 B.n269 VSUBS 0.007944f
C327 B.n270 VSUBS 0.007944f
C328 B.n271 VSUBS 0.007944f
C329 B.n272 VSUBS 0.007944f
C330 B.n273 VSUBS 0.007944f
C331 B.n274 VSUBS 0.007944f
C332 B.n275 VSUBS 0.007944f
C333 B.n276 VSUBS 0.007944f
C334 B.n277 VSUBS 0.007944f
C335 B.n278 VSUBS 0.007944f
C336 B.n279 VSUBS 0.007944f
C337 B.n280 VSUBS 0.007944f
C338 B.n281 VSUBS 0.007944f
C339 B.n282 VSUBS 0.007944f
C340 B.n283 VSUBS 0.007944f
C341 B.n284 VSUBS 0.007944f
C342 B.n285 VSUBS 0.007944f
C343 B.n286 VSUBS 0.007944f
C344 B.n287 VSUBS 0.007944f
C345 B.n288 VSUBS 0.007944f
C346 B.n289 VSUBS 0.007944f
C347 B.n290 VSUBS 0.007944f
C348 B.n291 VSUBS 0.007944f
C349 B.n292 VSUBS 0.007944f
C350 B.n293 VSUBS 0.007944f
C351 B.n294 VSUBS 0.007944f
C352 B.n295 VSUBS 0.007944f
C353 B.n296 VSUBS 0.007944f
C354 B.n297 VSUBS 0.007944f
C355 B.n298 VSUBS 0.007944f
C356 B.n299 VSUBS 0.007944f
C357 B.n300 VSUBS 0.007944f
C358 B.n301 VSUBS 0.007944f
C359 B.n302 VSUBS 0.007944f
C360 B.n303 VSUBS 0.007944f
C361 B.n304 VSUBS 0.007944f
C362 B.n305 VSUBS 0.007944f
C363 B.n306 VSUBS 0.007944f
C364 B.n307 VSUBS 0.007944f
C365 B.n308 VSUBS 0.007944f
C366 B.n309 VSUBS 0.007944f
C367 B.n310 VSUBS 0.007944f
C368 B.n311 VSUBS 0.007944f
C369 B.n312 VSUBS 0.007944f
C370 B.n313 VSUBS 0.007944f
C371 B.n314 VSUBS 0.007944f
C372 B.n315 VSUBS 0.007944f
C373 B.n316 VSUBS 0.007944f
C374 B.n317 VSUBS 0.007944f
C375 B.n318 VSUBS 0.007944f
C376 B.n319 VSUBS 0.007944f
C377 B.n320 VSUBS 0.007944f
C378 B.n321 VSUBS 0.007944f
C379 B.n322 VSUBS 0.007944f
C380 B.n323 VSUBS 0.007944f
C381 B.n324 VSUBS 0.007944f
C382 B.n325 VSUBS 0.007944f
C383 B.n326 VSUBS 0.007944f
C384 B.n327 VSUBS 0.018192f
C385 B.n328 VSUBS 0.019141f
C386 B.n329 VSUBS 0.017775f
C387 B.n330 VSUBS 0.007944f
C388 B.n331 VSUBS 0.007944f
C389 B.n332 VSUBS 0.007944f
C390 B.n333 VSUBS 0.007944f
C391 B.n334 VSUBS 0.007944f
C392 B.n335 VSUBS 0.007944f
C393 B.n336 VSUBS 0.007944f
C394 B.n337 VSUBS 0.007944f
C395 B.n338 VSUBS 0.007944f
C396 B.n339 VSUBS 0.007944f
C397 B.n340 VSUBS 0.007944f
C398 B.n341 VSUBS 0.007944f
C399 B.n342 VSUBS 0.007944f
C400 B.n343 VSUBS 0.007944f
C401 B.n344 VSUBS 0.007944f
C402 B.n345 VSUBS 0.007944f
C403 B.n346 VSUBS 0.007944f
C404 B.n347 VSUBS 0.007944f
C405 B.n348 VSUBS 0.007944f
C406 B.n349 VSUBS 0.007944f
C407 B.n350 VSUBS 0.007944f
C408 B.n351 VSUBS 0.007944f
C409 B.n352 VSUBS 0.007944f
C410 B.n353 VSUBS 0.007944f
C411 B.n354 VSUBS 0.007944f
C412 B.n355 VSUBS 0.007944f
C413 B.n356 VSUBS 0.007944f
C414 B.n357 VSUBS 0.007944f
C415 B.n358 VSUBS 0.007944f
C416 B.n359 VSUBS 0.007944f
C417 B.n360 VSUBS 0.007944f
C418 B.n361 VSUBS 0.007944f
C419 B.n362 VSUBS 0.007944f
C420 B.n363 VSUBS 0.007944f
C421 B.n364 VSUBS 0.007944f
C422 B.n365 VSUBS 0.007944f
C423 B.n366 VSUBS 0.007944f
C424 B.n367 VSUBS 0.007944f
C425 B.n368 VSUBS 0.007944f
C426 B.n369 VSUBS 0.007944f
C427 B.n370 VSUBS 0.007944f
C428 B.n371 VSUBS 0.007944f
C429 B.n372 VSUBS 0.007944f
C430 B.n373 VSUBS 0.007944f
C431 B.n374 VSUBS 0.007944f
C432 B.n375 VSUBS 0.007944f
C433 B.n376 VSUBS 0.007944f
C434 B.n377 VSUBS 0.007944f
C435 B.n378 VSUBS 0.007944f
C436 B.n379 VSUBS 0.007944f
C437 B.n380 VSUBS 0.007944f
C438 B.n381 VSUBS 0.017775f
C439 B.n382 VSUBS 0.017775f
C440 B.n383 VSUBS 0.019141f
C441 B.n384 VSUBS 0.007944f
C442 B.n385 VSUBS 0.007944f
C443 B.n386 VSUBS 0.007944f
C444 B.n387 VSUBS 0.007944f
C445 B.n388 VSUBS 0.007944f
C446 B.n389 VSUBS 0.007944f
C447 B.n390 VSUBS 0.007944f
C448 B.n391 VSUBS 0.007944f
C449 B.n392 VSUBS 0.007944f
C450 B.n393 VSUBS 0.007944f
C451 B.n394 VSUBS 0.007944f
C452 B.n395 VSUBS 0.007944f
C453 B.n396 VSUBS 0.007944f
C454 B.n397 VSUBS 0.007944f
C455 B.n398 VSUBS 0.007944f
C456 B.n399 VSUBS 0.007944f
C457 B.n400 VSUBS 0.007944f
C458 B.n401 VSUBS 0.007944f
C459 B.n402 VSUBS 0.007944f
C460 B.n403 VSUBS 0.007944f
C461 B.n404 VSUBS 0.007944f
C462 B.n405 VSUBS 0.007944f
C463 B.n406 VSUBS 0.007944f
C464 B.n407 VSUBS 0.007944f
C465 B.n408 VSUBS 0.007944f
C466 B.n409 VSUBS 0.007944f
C467 B.n410 VSUBS 0.007944f
C468 B.n411 VSUBS 0.007944f
C469 B.n412 VSUBS 0.007944f
C470 B.n413 VSUBS 0.007944f
C471 B.n414 VSUBS 0.007944f
C472 B.n415 VSUBS 0.007944f
C473 B.n416 VSUBS 0.007944f
C474 B.n417 VSUBS 0.007944f
C475 B.n418 VSUBS 0.007944f
C476 B.n419 VSUBS 0.007944f
C477 B.n420 VSUBS 0.007944f
C478 B.n421 VSUBS 0.007944f
C479 B.n422 VSUBS 0.007944f
C480 B.n423 VSUBS 0.007944f
C481 B.n424 VSUBS 0.007944f
C482 B.n425 VSUBS 0.007944f
C483 B.n426 VSUBS 0.007944f
C484 B.n427 VSUBS 0.007944f
C485 B.n428 VSUBS 0.007944f
C486 B.n429 VSUBS 0.007944f
C487 B.n430 VSUBS 0.007944f
C488 B.n431 VSUBS 0.007944f
C489 B.n432 VSUBS 0.007944f
C490 B.n433 VSUBS 0.007944f
C491 B.n434 VSUBS 0.007944f
C492 B.n435 VSUBS 0.007944f
C493 B.n436 VSUBS 0.007944f
C494 B.n437 VSUBS 0.007944f
C495 B.n438 VSUBS 0.007944f
C496 B.n439 VSUBS 0.007944f
C497 B.n440 VSUBS 0.007944f
C498 B.n441 VSUBS 0.007944f
C499 B.n442 VSUBS 0.007944f
C500 B.n443 VSUBS 0.007944f
C501 B.n444 VSUBS 0.007944f
C502 B.n445 VSUBS 0.007944f
C503 B.n446 VSUBS 0.007944f
C504 B.n447 VSUBS 0.007944f
C505 B.n448 VSUBS 0.007944f
C506 B.n449 VSUBS 0.007944f
C507 B.n450 VSUBS 0.007944f
C508 B.n451 VSUBS 0.007944f
C509 B.n452 VSUBS 0.005491f
C510 B.n453 VSUBS 0.018405f
C511 B.n454 VSUBS 0.006425f
C512 B.n455 VSUBS 0.007944f
C513 B.n456 VSUBS 0.007944f
C514 B.n457 VSUBS 0.007944f
C515 B.n458 VSUBS 0.007944f
C516 B.n459 VSUBS 0.007944f
C517 B.n460 VSUBS 0.007944f
C518 B.n461 VSUBS 0.007944f
C519 B.n462 VSUBS 0.007944f
C520 B.n463 VSUBS 0.007944f
C521 B.n464 VSUBS 0.007944f
C522 B.n465 VSUBS 0.007944f
C523 B.n466 VSUBS 0.006425f
C524 B.n467 VSUBS 0.007944f
C525 B.n468 VSUBS 0.007944f
C526 B.n469 VSUBS 0.005491f
C527 B.n470 VSUBS 0.007944f
C528 B.n471 VSUBS 0.007944f
C529 B.n472 VSUBS 0.007944f
C530 B.n473 VSUBS 0.007944f
C531 B.n474 VSUBS 0.007944f
C532 B.n475 VSUBS 0.007944f
C533 B.n476 VSUBS 0.007944f
C534 B.n477 VSUBS 0.007944f
C535 B.n478 VSUBS 0.007944f
C536 B.n479 VSUBS 0.007944f
C537 B.n480 VSUBS 0.007944f
C538 B.n481 VSUBS 0.007944f
C539 B.n482 VSUBS 0.007944f
C540 B.n483 VSUBS 0.007944f
C541 B.n484 VSUBS 0.007944f
C542 B.n485 VSUBS 0.007944f
C543 B.n486 VSUBS 0.007944f
C544 B.n487 VSUBS 0.007944f
C545 B.n488 VSUBS 0.007944f
C546 B.n489 VSUBS 0.007944f
C547 B.n490 VSUBS 0.007944f
C548 B.n491 VSUBS 0.007944f
C549 B.n492 VSUBS 0.007944f
C550 B.n493 VSUBS 0.007944f
C551 B.n494 VSUBS 0.007944f
C552 B.n495 VSUBS 0.007944f
C553 B.n496 VSUBS 0.007944f
C554 B.n497 VSUBS 0.007944f
C555 B.n498 VSUBS 0.007944f
C556 B.n499 VSUBS 0.007944f
C557 B.n500 VSUBS 0.007944f
C558 B.n501 VSUBS 0.007944f
C559 B.n502 VSUBS 0.007944f
C560 B.n503 VSUBS 0.007944f
C561 B.n504 VSUBS 0.007944f
C562 B.n505 VSUBS 0.007944f
C563 B.n506 VSUBS 0.007944f
C564 B.n507 VSUBS 0.007944f
C565 B.n508 VSUBS 0.007944f
C566 B.n509 VSUBS 0.007944f
C567 B.n510 VSUBS 0.007944f
C568 B.n511 VSUBS 0.007944f
C569 B.n512 VSUBS 0.007944f
C570 B.n513 VSUBS 0.007944f
C571 B.n514 VSUBS 0.007944f
C572 B.n515 VSUBS 0.007944f
C573 B.n516 VSUBS 0.007944f
C574 B.n517 VSUBS 0.007944f
C575 B.n518 VSUBS 0.007944f
C576 B.n519 VSUBS 0.007944f
C577 B.n520 VSUBS 0.007944f
C578 B.n521 VSUBS 0.007944f
C579 B.n522 VSUBS 0.007944f
C580 B.n523 VSUBS 0.007944f
C581 B.n524 VSUBS 0.007944f
C582 B.n525 VSUBS 0.007944f
C583 B.n526 VSUBS 0.007944f
C584 B.n527 VSUBS 0.007944f
C585 B.n528 VSUBS 0.007944f
C586 B.n529 VSUBS 0.007944f
C587 B.n530 VSUBS 0.007944f
C588 B.n531 VSUBS 0.007944f
C589 B.n532 VSUBS 0.007944f
C590 B.n533 VSUBS 0.007944f
C591 B.n534 VSUBS 0.007944f
C592 B.n535 VSUBS 0.007944f
C593 B.n536 VSUBS 0.007944f
C594 B.n537 VSUBS 0.019141f
C595 B.n538 VSUBS 0.019141f
C596 B.n539 VSUBS 0.017775f
C597 B.n540 VSUBS 0.007944f
C598 B.n541 VSUBS 0.007944f
C599 B.n542 VSUBS 0.007944f
C600 B.n543 VSUBS 0.007944f
C601 B.n544 VSUBS 0.007944f
C602 B.n545 VSUBS 0.007944f
C603 B.n546 VSUBS 0.007944f
C604 B.n547 VSUBS 0.007944f
C605 B.n548 VSUBS 0.007944f
C606 B.n549 VSUBS 0.007944f
C607 B.n550 VSUBS 0.007944f
C608 B.n551 VSUBS 0.007944f
C609 B.n552 VSUBS 0.007944f
C610 B.n553 VSUBS 0.007944f
C611 B.n554 VSUBS 0.007944f
C612 B.n555 VSUBS 0.007944f
C613 B.n556 VSUBS 0.007944f
C614 B.n557 VSUBS 0.007944f
C615 B.n558 VSUBS 0.007944f
C616 B.n559 VSUBS 0.007944f
C617 B.n560 VSUBS 0.007944f
C618 B.n561 VSUBS 0.007944f
C619 B.n562 VSUBS 0.007944f
C620 B.n563 VSUBS 0.010366f
C621 B.n564 VSUBS 0.011043f
C622 B.n565 VSUBS 0.02196f
C623 VDD2.t0 VSUBS 0.304006f
C624 VDD2.t3 VSUBS 0.304006f
C625 VDD2.n0 VSUBS 3.13659f
C626 VDD2.t1 VSUBS 0.304006f
C627 VDD2.t2 VSUBS 0.304006f
C628 VDD2.n1 VSUBS 2.44356f
C629 VDD2.n2 VSUBS 4.21341f
C630 VTAIL.t6 VSUBS 2.43102f
C631 VTAIL.n0 VSUBS 0.674081f
C632 VTAIL.t2 VSUBS 2.43102f
C633 VTAIL.n1 VSUBS 0.703887f
C634 VTAIL.t3 VSUBS 2.43102f
C635 VTAIL.n2 VSUBS 1.90908f
C636 VTAIL.t4 VSUBS 2.43102f
C637 VTAIL.n3 VSUBS 1.90907f
C638 VTAIL.t5 VSUBS 2.43102f
C639 VTAIL.n4 VSUBS 0.703883f
C640 VTAIL.t1 VSUBS 2.43102f
C641 VTAIL.n5 VSUBS 0.703883f
C642 VTAIL.t0 VSUBS 2.43102f
C643 VTAIL.n6 VSUBS 1.90908f
C644 VTAIL.t7 VSUBS 2.43102f
C645 VTAIL.n7 VSUBS 1.87075f
C646 VN.t3 VSUBS 1.71148f
C647 VN.t0 VSUBS 1.71141f
C648 VN.n0 VSUBS 1.26563f
C649 VN.t1 VSUBS 1.71148f
C650 VN.t2 VSUBS 1.71141f
C651 VN.n1 VSUBS 2.49739f
.ends

