* NGSPICE file created from diff_pair_sample_1547.ext - technology: sky130A

.subckt diff_pair_sample_1547 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t4 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=1.353 pd=8.53 as=1.353 ps=8.53 w=8.2 l=2.7
X1 B.t11 B.t9 B.t10 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=3.198 pd=17.18 as=0 ps=0 w=8.2 l=2.7
X2 B.t8 B.t6 B.t7 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=3.198 pd=17.18 as=0 ps=0 w=8.2 l=2.7
X3 VDD2.t5 VN.t0 VTAIL.t4 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=3.198 pd=17.18 as=1.353 ps=8.53 w=8.2 l=2.7
X4 VTAIL.t5 VN.t1 VDD2.t4 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=1.353 pd=8.53 as=1.353 ps=8.53 w=8.2 l=2.7
X5 VDD1.t2 VP.t1 VTAIL.t10 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=1.353 pd=8.53 as=3.198 ps=17.18 w=8.2 l=2.7
X6 VTAIL.t9 VP.t2 VDD1.t1 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=1.353 pd=8.53 as=1.353 ps=8.53 w=8.2 l=2.7
X7 B.t5 B.t3 B.t4 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=3.198 pd=17.18 as=0 ps=0 w=8.2 l=2.7
X8 VDD2.t3 VN.t2 VTAIL.t2 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=1.353 pd=8.53 as=3.198 ps=17.18 w=8.2 l=2.7
X9 VDD2.t2 VN.t3 VTAIL.t0 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=3.198 pd=17.18 as=1.353 ps=8.53 w=8.2 l=2.7
X10 VDD1.t5 VP.t3 VTAIL.t8 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=3.198 pd=17.18 as=1.353 ps=8.53 w=8.2 l=2.7
X11 B.t2 B.t0 B.t1 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=3.198 pd=17.18 as=0 ps=0 w=8.2 l=2.7
X12 VDD2.t1 VN.t4 VTAIL.t1 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=1.353 pd=8.53 as=3.198 ps=17.18 w=8.2 l=2.7
X13 VDD1.t3 VP.t4 VTAIL.t7 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=1.353 pd=8.53 as=3.198 ps=17.18 w=8.2 l=2.7
X14 VTAIL.t3 VN.t5 VDD2.t0 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=1.353 pd=8.53 as=1.353 ps=8.53 w=8.2 l=2.7
X15 VDD1.t0 VP.t5 VTAIL.t6 w_n3394_n2608# sky130_fd_pr__pfet_01v8 ad=3.198 pd=17.18 as=1.353 ps=8.53 w=8.2 l=2.7
R0 VP.n13 VP.n12 161.3
R1 VP.n14 VP.n9 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n17 VP.n8 161.3
R4 VP.n19 VP.n18 161.3
R5 VP.n20 VP.n7 161.3
R6 VP.n43 VP.n0 161.3
R7 VP.n42 VP.n41 161.3
R8 VP.n40 VP.n1 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n37 VP.n2 161.3
R11 VP.n36 VP.n35 161.3
R12 VP.n34 VP.n3 161.3
R13 VP.n33 VP.n32 161.3
R14 VP.n31 VP.n4 161.3
R15 VP.n30 VP.n29 161.3
R16 VP.n28 VP.n5 161.3
R17 VP.n27 VP.n26 161.3
R18 VP.n25 VP.n6 161.3
R19 VP.n24 VP.n23 109.433
R20 VP.n45 VP.n44 109.433
R21 VP.n22 VP.n21 109.433
R22 VP.n11 VP.t5 106.007
R23 VP.n3 VP.t2 73.1931
R24 VP.n24 VP.t3 73.1931
R25 VP.n44 VP.t4 73.1931
R26 VP.n10 VP.t0 73.1931
R27 VP.n21 VP.t1 73.1931
R28 VP.n11 VP.n10 49.0351
R29 VP.n23 VP.n22 46.1019
R30 VP.n30 VP.n5 42.0302
R31 VP.n38 VP.n1 42.0302
R32 VP.n15 VP.n8 42.0302
R33 VP.n31 VP.n30 39.1239
R34 VP.n38 VP.n37 39.1239
R35 VP.n15 VP.n14 39.1239
R36 VP.n26 VP.n25 24.5923
R37 VP.n26 VP.n5 24.5923
R38 VP.n32 VP.n31 24.5923
R39 VP.n32 VP.n3 24.5923
R40 VP.n36 VP.n3 24.5923
R41 VP.n37 VP.n36 24.5923
R42 VP.n42 VP.n1 24.5923
R43 VP.n43 VP.n42 24.5923
R44 VP.n19 VP.n8 24.5923
R45 VP.n20 VP.n19 24.5923
R46 VP.n13 VP.n10 24.5923
R47 VP.n14 VP.n13 24.5923
R48 VP.n12 VP.n11 5.10935
R49 VP.n25 VP.n24 1.47601
R50 VP.n44 VP.n43 1.47601
R51 VP.n21 VP.n20 1.47601
R52 VP.n22 VP.n7 0.278335
R53 VP.n23 VP.n6 0.278335
R54 VP.n45 VP.n0 0.278335
R55 VP.n12 VP.n9 0.189894
R56 VP.n16 VP.n9 0.189894
R57 VP.n17 VP.n16 0.189894
R58 VP.n18 VP.n17 0.189894
R59 VP.n18 VP.n7 0.189894
R60 VP.n27 VP.n6 0.189894
R61 VP.n28 VP.n27 0.189894
R62 VP.n29 VP.n28 0.189894
R63 VP.n29 VP.n4 0.189894
R64 VP.n33 VP.n4 0.189894
R65 VP.n34 VP.n33 0.189894
R66 VP.n35 VP.n34 0.189894
R67 VP.n35 VP.n2 0.189894
R68 VP.n39 VP.n2 0.189894
R69 VP.n40 VP.n39 0.189894
R70 VP.n41 VP.n40 0.189894
R71 VP.n41 VP.n0 0.189894
R72 VP VP.n45 0.153485
R73 VDD1 VDD1.t0 88.0418
R74 VDD1.n1 VDD1.t5 87.9282
R75 VDD1.n1 VDD1.n0 82.658
R76 VDD1.n3 VDD1.n2 82.0604
R77 VDD1.n3 VDD1.n1 41.1625
R78 VDD1.n2 VDD1.t4 3.96452
R79 VDD1.n2 VDD1.t2 3.96452
R80 VDD1.n0 VDD1.t1 3.96452
R81 VDD1.n0 VDD1.t3 3.96452
R82 VDD1 VDD1.n3 0.595328
R83 VTAIL.n7 VTAIL.t2 69.3458
R84 VTAIL.n11 VTAIL.t1 69.3457
R85 VTAIL.n2 VTAIL.t7 69.3457
R86 VTAIL.n10 VTAIL.t10 69.3457
R87 VTAIL.n9 VTAIL.n8 65.3818
R88 VTAIL.n6 VTAIL.n5 65.3818
R89 VTAIL.n1 VTAIL.n0 65.3816
R90 VTAIL.n4 VTAIL.n3 65.3816
R91 VTAIL.n6 VTAIL.n4 24.66
R92 VTAIL.n11 VTAIL.n10 22.0479
R93 VTAIL.n0 VTAIL.t0 3.96452
R94 VTAIL.n0 VTAIL.t5 3.96452
R95 VTAIL.n3 VTAIL.t8 3.96452
R96 VTAIL.n3 VTAIL.t9 3.96452
R97 VTAIL.n8 VTAIL.t6 3.96452
R98 VTAIL.n8 VTAIL.t11 3.96452
R99 VTAIL.n5 VTAIL.t4 3.96452
R100 VTAIL.n5 VTAIL.t3 3.96452
R101 VTAIL.n7 VTAIL.n6 2.61257
R102 VTAIL.n10 VTAIL.n9 2.61257
R103 VTAIL.n4 VTAIL.n2 2.61257
R104 VTAIL VTAIL.n11 1.90136
R105 VTAIL.n9 VTAIL.n7 1.77636
R106 VTAIL.n2 VTAIL.n1 1.77636
R107 VTAIL VTAIL.n1 0.711707
R108 B.n337 B.n336 585
R109 B.n335 B.n108 585
R110 B.n334 B.n333 585
R111 B.n332 B.n109 585
R112 B.n331 B.n330 585
R113 B.n329 B.n110 585
R114 B.n328 B.n327 585
R115 B.n326 B.n111 585
R116 B.n325 B.n324 585
R117 B.n323 B.n112 585
R118 B.n322 B.n321 585
R119 B.n320 B.n113 585
R120 B.n319 B.n318 585
R121 B.n317 B.n114 585
R122 B.n316 B.n315 585
R123 B.n314 B.n115 585
R124 B.n313 B.n312 585
R125 B.n311 B.n116 585
R126 B.n310 B.n309 585
R127 B.n308 B.n117 585
R128 B.n307 B.n306 585
R129 B.n305 B.n118 585
R130 B.n304 B.n303 585
R131 B.n302 B.n119 585
R132 B.n301 B.n300 585
R133 B.n299 B.n120 585
R134 B.n298 B.n297 585
R135 B.n296 B.n121 585
R136 B.n295 B.n294 585
R137 B.n293 B.n122 585
R138 B.n291 B.n290 585
R139 B.n289 B.n125 585
R140 B.n288 B.n287 585
R141 B.n286 B.n126 585
R142 B.n285 B.n284 585
R143 B.n283 B.n127 585
R144 B.n282 B.n281 585
R145 B.n280 B.n128 585
R146 B.n279 B.n278 585
R147 B.n277 B.n129 585
R148 B.n276 B.n275 585
R149 B.n271 B.n130 585
R150 B.n270 B.n269 585
R151 B.n268 B.n131 585
R152 B.n267 B.n266 585
R153 B.n265 B.n132 585
R154 B.n264 B.n263 585
R155 B.n262 B.n133 585
R156 B.n261 B.n260 585
R157 B.n259 B.n134 585
R158 B.n258 B.n257 585
R159 B.n256 B.n135 585
R160 B.n255 B.n254 585
R161 B.n253 B.n136 585
R162 B.n252 B.n251 585
R163 B.n250 B.n137 585
R164 B.n249 B.n248 585
R165 B.n247 B.n138 585
R166 B.n246 B.n245 585
R167 B.n244 B.n139 585
R168 B.n243 B.n242 585
R169 B.n241 B.n140 585
R170 B.n240 B.n239 585
R171 B.n238 B.n141 585
R172 B.n237 B.n236 585
R173 B.n235 B.n142 585
R174 B.n234 B.n233 585
R175 B.n232 B.n143 585
R176 B.n231 B.n230 585
R177 B.n229 B.n144 585
R178 B.n338 B.n107 585
R179 B.n340 B.n339 585
R180 B.n341 B.n106 585
R181 B.n343 B.n342 585
R182 B.n344 B.n105 585
R183 B.n346 B.n345 585
R184 B.n347 B.n104 585
R185 B.n349 B.n348 585
R186 B.n350 B.n103 585
R187 B.n352 B.n351 585
R188 B.n353 B.n102 585
R189 B.n355 B.n354 585
R190 B.n356 B.n101 585
R191 B.n358 B.n357 585
R192 B.n359 B.n100 585
R193 B.n361 B.n360 585
R194 B.n362 B.n99 585
R195 B.n364 B.n363 585
R196 B.n365 B.n98 585
R197 B.n367 B.n366 585
R198 B.n368 B.n97 585
R199 B.n370 B.n369 585
R200 B.n371 B.n96 585
R201 B.n373 B.n372 585
R202 B.n374 B.n95 585
R203 B.n376 B.n375 585
R204 B.n377 B.n94 585
R205 B.n379 B.n378 585
R206 B.n380 B.n93 585
R207 B.n382 B.n381 585
R208 B.n383 B.n92 585
R209 B.n385 B.n384 585
R210 B.n386 B.n91 585
R211 B.n388 B.n387 585
R212 B.n389 B.n90 585
R213 B.n391 B.n390 585
R214 B.n392 B.n89 585
R215 B.n394 B.n393 585
R216 B.n395 B.n88 585
R217 B.n397 B.n396 585
R218 B.n398 B.n87 585
R219 B.n400 B.n399 585
R220 B.n401 B.n86 585
R221 B.n403 B.n402 585
R222 B.n404 B.n85 585
R223 B.n406 B.n405 585
R224 B.n407 B.n84 585
R225 B.n409 B.n408 585
R226 B.n410 B.n83 585
R227 B.n412 B.n411 585
R228 B.n413 B.n82 585
R229 B.n415 B.n414 585
R230 B.n416 B.n81 585
R231 B.n418 B.n417 585
R232 B.n419 B.n80 585
R233 B.n421 B.n420 585
R234 B.n422 B.n79 585
R235 B.n424 B.n423 585
R236 B.n425 B.n78 585
R237 B.n427 B.n426 585
R238 B.n428 B.n77 585
R239 B.n430 B.n429 585
R240 B.n431 B.n76 585
R241 B.n433 B.n432 585
R242 B.n434 B.n75 585
R243 B.n436 B.n435 585
R244 B.n437 B.n74 585
R245 B.n439 B.n438 585
R246 B.n440 B.n73 585
R247 B.n442 B.n441 585
R248 B.n443 B.n72 585
R249 B.n445 B.n444 585
R250 B.n446 B.n71 585
R251 B.n448 B.n447 585
R252 B.n449 B.n70 585
R253 B.n451 B.n450 585
R254 B.n452 B.n69 585
R255 B.n454 B.n453 585
R256 B.n455 B.n68 585
R257 B.n457 B.n456 585
R258 B.n458 B.n67 585
R259 B.n460 B.n459 585
R260 B.n461 B.n66 585
R261 B.n463 B.n462 585
R262 B.n464 B.n65 585
R263 B.n466 B.n465 585
R264 B.n467 B.n64 585
R265 B.n469 B.n468 585
R266 B.n575 B.n574 585
R267 B.n573 B.n24 585
R268 B.n572 B.n571 585
R269 B.n570 B.n25 585
R270 B.n569 B.n568 585
R271 B.n567 B.n26 585
R272 B.n566 B.n565 585
R273 B.n564 B.n27 585
R274 B.n563 B.n562 585
R275 B.n561 B.n28 585
R276 B.n560 B.n559 585
R277 B.n558 B.n29 585
R278 B.n557 B.n556 585
R279 B.n555 B.n30 585
R280 B.n554 B.n553 585
R281 B.n552 B.n31 585
R282 B.n551 B.n550 585
R283 B.n549 B.n32 585
R284 B.n548 B.n547 585
R285 B.n546 B.n33 585
R286 B.n545 B.n544 585
R287 B.n543 B.n34 585
R288 B.n542 B.n541 585
R289 B.n540 B.n35 585
R290 B.n539 B.n538 585
R291 B.n537 B.n36 585
R292 B.n536 B.n535 585
R293 B.n534 B.n37 585
R294 B.n533 B.n532 585
R295 B.n531 B.n38 585
R296 B.n530 B.n529 585
R297 B.n528 B.n39 585
R298 B.n527 B.n526 585
R299 B.n525 B.n43 585
R300 B.n524 B.n523 585
R301 B.n522 B.n44 585
R302 B.n521 B.n520 585
R303 B.n519 B.n45 585
R304 B.n518 B.n517 585
R305 B.n516 B.n46 585
R306 B.n514 B.n513 585
R307 B.n512 B.n49 585
R308 B.n511 B.n510 585
R309 B.n509 B.n50 585
R310 B.n508 B.n507 585
R311 B.n506 B.n51 585
R312 B.n505 B.n504 585
R313 B.n503 B.n52 585
R314 B.n502 B.n501 585
R315 B.n500 B.n53 585
R316 B.n499 B.n498 585
R317 B.n497 B.n54 585
R318 B.n496 B.n495 585
R319 B.n494 B.n55 585
R320 B.n493 B.n492 585
R321 B.n491 B.n56 585
R322 B.n490 B.n489 585
R323 B.n488 B.n57 585
R324 B.n487 B.n486 585
R325 B.n485 B.n58 585
R326 B.n484 B.n483 585
R327 B.n482 B.n59 585
R328 B.n481 B.n480 585
R329 B.n479 B.n60 585
R330 B.n478 B.n477 585
R331 B.n476 B.n61 585
R332 B.n475 B.n474 585
R333 B.n473 B.n62 585
R334 B.n472 B.n471 585
R335 B.n470 B.n63 585
R336 B.n576 B.n23 585
R337 B.n578 B.n577 585
R338 B.n579 B.n22 585
R339 B.n581 B.n580 585
R340 B.n582 B.n21 585
R341 B.n584 B.n583 585
R342 B.n585 B.n20 585
R343 B.n587 B.n586 585
R344 B.n588 B.n19 585
R345 B.n590 B.n589 585
R346 B.n591 B.n18 585
R347 B.n593 B.n592 585
R348 B.n594 B.n17 585
R349 B.n596 B.n595 585
R350 B.n597 B.n16 585
R351 B.n599 B.n598 585
R352 B.n600 B.n15 585
R353 B.n602 B.n601 585
R354 B.n603 B.n14 585
R355 B.n605 B.n604 585
R356 B.n606 B.n13 585
R357 B.n608 B.n607 585
R358 B.n609 B.n12 585
R359 B.n611 B.n610 585
R360 B.n612 B.n11 585
R361 B.n614 B.n613 585
R362 B.n615 B.n10 585
R363 B.n617 B.n616 585
R364 B.n618 B.n9 585
R365 B.n620 B.n619 585
R366 B.n621 B.n8 585
R367 B.n623 B.n622 585
R368 B.n624 B.n7 585
R369 B.n626 B.n625 585
R370 B.n627 B.n6 585
R371 B.n629 B.n628 585
R372 B.n630 B.n5 585
R373 B.n632 B.n631 585
R374 B.n633 B.n4 585
R375 B.n635 B.n634 585
R376 B.n636 B.n3 585
R377 B.n638 B.n637 585
R378 B.n639 B.n0 585
R379 B.n2 B.n1 585
R380 B.n166 B.n165 585
R381 B.n168 B.n167 585
R382 B.n169 B.n164 585
R383 B.n171 B.n170 585
R384 B.n172 B.n163 585
R385 B.n174 B.n173 585
R386 B.n175 B.n162 585
R387 B.n177 B.n176 585
R388 B.n178 B.n161 585
R389 B.n180 B.n179 585
R390 B.n181 B.n160 585
R391 B.n183 B.n182 585
R392 B.n184 B.n159 585
R393 B.n186 B.n185 585
R394 B.n187 B.n158 585
R395 B.n189 B.n188 585
R396 B.n190 B.n157 585
R397 B.n192 B.n191 585
R398 B.n193 B.n156 585
R399 B.n195 B.n194 585
R400 B.n196 B.n155 585
R401 B.n198 B.n197 585
R402 B.n199 B.n154 585
R403 B.n201 B.n200 585
R404 B.n202 B.n153 585
R405 B.n204 B.n203 585
R406 B.n205 B.n152 585
R407 B.n207 B.n206 585
R408 B.n208 B.n151 585
R409 B.n210 B.n209 585
R410 B.n211 B.n150 585
R411 B.n213 B.n212 585
R412 B.n214 B.n149 585
R413 B.n216 B.n215 585
R414 B.n217 B.n148 585
R415 B.n219 B.n218 585
R416 B.n220 B.n147 585
R417 B.n222 B.n221 585
R418 B.n223 B.n146 585
R419 B.n225 B.n224 585
R420 B.n226 B.n145 585
R421 B.n228 B.n227 585
R422 B.n227 B.n144 578.989
R423 B.n338 B.n337 578.989
R424 B.n470 B.n469 578.989
R425 B.n574 B.n23 578.989
R426 B.n272 B.t6 281.385
R427 B.n123 B.t3 281.385
R428 B.n47 B.t9 281.385
R429 B.n40 B.t0 281.385
R430 B.n641 B.n640 256.663
R431 B.n640 B.n639 235.042
R432 B.n640 B.n2 235.042
R433 B.n123 B.t4 168.065
R434 B.n47 B.t11 168.065
R435 B.n272 B.t7 168.056
R436 B.n40 B.t2 168.056
R437 B.n231 B.n144 163.367
R438 B.n232 B.n231 163.367
R439 B.n233 B.n232 163.367
R440 B.n233 B.n142 163.367
R441 B.n237 B.n142 163.367
R442 B.n238 B.n237 163.367
R443 B.n239 B.n238 163.367
R444 B.n239 B.n140 163.367
R445 B.n243 B.n140 163.367
R446 B.n244 B.n243 163.367
R447 B.n245 B.n244 163.367
R448 B.n245 B.n138 163.367
R449 B.n249 B.n138 163.367
R450 B.n250 B.n249 163.367
R451 B.n251 B.n250 163.367
R452 B.n251 B.n136 163.367
R453 B.n255 B.n136 163.367
R454 B.n256 B.n255 163.367
R455 B.n257 B.n256 163.367
R456 B.n257 B.n134 163.367
R457 B.n261 B.n134 163.367
R458 B.n262 B.n261 163.367
R459 B.n263 B.n262 163.367
R460 B.n263 B.n132 163.367
R461 B.n267 B.n132 163.367
R462 B.n268 B.n267 163.367
R463 B.n269 B.n268 163.367
R464 B.n269 B.n130 163.367
R465 B.n276 B.n130 163.367
R466 B.n277 B.n276 163.367
R467 B.n278 B.n277 163.367
R468 B.n278 B.n128 163.367
R469 B.n282 B.n128 163.367
R470 B.n283 B.n282 163.367
R471 B.n284 B.n283 163.367
R472 B.n284 B.n126 163.367
R473 B.n288 B.n126 163.367
R474 B.n289 B.n288 163.367
R475 B.n290 B.n289 163.367
R476 B.n290 B.n122 163.367
R477 B.n295 B.n122 163.367
R478 B.n296 B.n295 163.367
R479 B.n297 B.n296 163.367
R480 B.n297 B.n120 163.367
R481 B.n301 B.n120 163.367
R482 B.n302 B.n301 163.367
R483 B.n303 B.n302 163.367
R484 B.n303 B.n118 163.367
R485 B.n307 B.n118 163.367
R486 B.n308 B.n307 163.367
R487 B.n309 B.n308 163.367
R488 B.n309 B.n116 163.367
R489 B.n313 B.n116 163.367
R490 B.n314 B.n313 163.367
R491 B.n315 B.n314 163.367
R492 B.n315 B.n114 163.367
R493 B.n319 B.n114 163.367
R494 B.n320 B.n319 163.367
R495 B.n321 B.n320 163.367
R496 B.n321 B.n112 163.367
R497 B.n325 B.n112 163.367
R498 B.n326 B.n325 163.367
R499 B.n327 B.n326 163.367
R500 B.n327 B.n110 163.367
R501 B.n331 B.n110 163.367
R502 B.n332 B.n331 163.367
R503 B.n333 B.n332 163.367
R504 B.n333 B.n108 163.367
R505 B.n337 B.n108 163.367
R506 B.n469 B.n64 163.367
R507 B.n465 B.n64 163.367
R508 B.n465 B.n464 163.367
R509 B.n464 B.n463 163.367
R510 B.n463 B.n66 163.367
R511 B.n459 B.n66 163.367
R512 B.n459 B.n458 163.367
R513 B.n458 B.n457 163.367
R514 B.n457 B.n68 163.367
R515 B.n453 B.n68 163.367
R516 B.n453 B.n452 163.367
R517 B.n452 B.n451 163.367
R518 B.n451 B.n70 163.367
R519 B.n447 B.n70 163.367
R520 B.n447 B.n446 163.367
R521 B.n446 B.n445 163.367
R522 B.n445 B.n72 163.367
R523 B.n441 B.n72 163.367
R524 B.n441 B.n440 163.367
R525 B.n440 B.n439 163.367
R526 B.n439 B.n74 163.367
R527 B.n435 B.n74 163.367
R528 B.n435 B.n434 163.367
R529 B.n434 B.n433 163.367
R530 B.n433 B.n76 163.367
R531 B.n429 B.n76 163.367
R532 B.n429 B.n428 163.367
R533 B.n428 B.n427 163.367
R534 B.n427 B.n78 163.367
R535 B.n423 B.n78 163.367
R536 B.n423 B.n422 163.367
R537 B.n422 B.n421 163.367
R538 B.n421 B.n80 163.367
R539 B.n417 B.n80 163.367
R540 B.n417 B.n416 163.367
R541 B.n416 B.n415 163.367
R542 B.n415 B.n82 163.367
R543 B.n411 B.n82 163.367
R544 B.n411 B.n410 163.367
R545 B.n410 B.n409 163.367
R546 B.n409 B.n84 163.367
R547 B.n405 B.n84 163.367
R548 B.n405 B.n404 163.367
R549 B.n404 B.n403 163.367
R550 B.n403 B.n86 163.367
R551 B.n399 B.n86 163.367
R552 B.n399 B.n398 163.367
R553 B.n398 B.n397 163.367
R554 B.n397 B.n88 163.367
R555 B.n393 B.n88 163.367
R556 B.n393 B.n392 163.367
R557 B.n392 B.n391 163.367
R558 B.n391 B.n90 163.367
R559 B.n387 B.n90 163.367
R560 B.n387 B.n386 163.367
R561 B.n386 B.n385 163.367
R562 B.n385 B.n92 163.367
R563 B.n381 B.n92 163.367
R564 B.n381 B.n380 163.367
R565 B.n380 B.n379 163.367
R566 B.n379 B.n94 163.367
R567 B.n375 B.n94 163.367
R568 B.n375 B.n374 163.367
R569 B.n374 B.n373 163.367
R570 B.n373 B.n96 163.367
R571 B.n369 B.n96 163.367
R572 B.n369 B.n368 163.367
R573 B.n368 B.n367 163.367
R574 B.n367 B.n98 163.367
R575 B.n363 B.n98 163.367
R576 B.n363 B.n362 163.367
R577 B.n362 B.n361 163.367
R578 B.n361 B.n100 163.367
R579 B.n357 B.n100 163.367
R580 B.n357 B.n356 163.367
R581 B.n356 B.n355 163.367
R582 B.n355 B.n102 163.367
R583 B.n351 B.n102 163.367
R584 B.n351 B.n350 163.367
R585 B.n350 B.n349 163.367
R586 B.n349 B.n104 163.367
R587 B.n345 B.n104 163.367
R588 B.n345 B.n344 163.367
R589 B.n344 B.n343 163.367
R590 B.n343 B.n106 163.367
R591 B.n339 B.n106 163.367
R592 B.n339 B.n338 163.367
R593 B.n574 B.n573 163.367
R594 B.n573 B.n572 163.367
R595 B.n572 B.n25 163.367
R596 B.n568 B.n25 163.367
R597 B.n568 B.n567 163.367
R598 B.n567 B.n566 163.367
R599 B.n566 B.n27 163.367
R600 B.n562 B.n27 163.367
R601 B.n562 B.n561 163.367
R602 B.n561 B.n560 163.367
R603 B.n560 B.n29 163.367
R604 B.n556 B.n29 163.367
R605 B.n556 B.n555 163.367
R606 B.n555 B.n554 163.367
R607 B.n554 B.n31 163.367
R608 B.n550 B.n31 163.367
R609 B.n550 B.n549 163.367
R610 B.n549 B.n548 163.367
R611 B.n548 B.n33 163.367
R612 B.n544 B.n33 163.367
R613 B.n544 B.n543 163.367
R614 B.n543 B.n542 163.367
R615 B.n542 B.n35 163.367
R616 B.n538 B.n35 163.367
R617 B.n538 B.n537 163.367
R618 B.n537 B.n536 163.367
R619 B.n536 B.n37 163.367
R620 B.n532 B.n37 163.367
R621 B.n532 B.n531 163.367
R622 B.n531 B.n530 163.367
R623 B.n530 B.n39 163.367
R624 B.n526 B.n39 163.367
R625 B.n526 B.n525 163.367
R626 B.n525 B.n524 163.367
R627 B.n524 B.n44 163.367
R628 B.n520 B.n44 163.367
R629 B.n520 B.n519 163.367
R630 B.n519 B.n518 163.367
R631 B.n518 B.n46 163.367
R632 B.n513 B.n46 163.367
R633 B.n513 B.n512 163.367
R634 B.n512 B.n511 163.367
R635 B.n511 B.n50 163.367
R636 B.n507 B.n50 163.367
R637 B.n507 B.n506 163.367
R638 B.n506 B.n505 163.367
R639 B.n505 B.n52 163.367
R640 B.n501 B.n52 163.367
R641 B.n501 B.n500 163.367
R642 B.n500 B.n499 163.367
R643 B.n499 B.n54 163.367
R644 B.n495 B.n54 163.367
R645 B.n495 B.n494 163.367
R646 B.n494 B.n493 163.367
R647 B.n493 B.n56 163.367
R648 B.n489 B.n56 163.367
R649 B.n489 B.n488 163.367
R650 B.n488 B.n487 163.367
R651 B.n487 B.n58 163.367
R652 B.n483 B.n58 163.367
R653 B.n483 B.n482 163.367
R654 B.n482 B.n481 163.367
R655 B.n481 B.n60 163.367
R656 B.n477 B.n60 163.367
R657 B.n477 B.n476 163.367
R658 B.n476 B.n475 163.367
R659 B.n475 B.n62 163.367
R660 B.n471 B.n62 163.367
R661 B.n471 B.n470 163.367
R662 B.n578 B.n23 163.367
R663 B.n579 B.n578 163.367
R664 B.n580 B.n579 163.367
R665 B.n580 B.n21 163.367
R666 B.n584 B.n21 163.367
R667 B.n585 B.n584 163.367
R668 B.n586 B.n585 163.367
R669 B.n586 B.n19 163.367
R670 B.n590 B.n19 163.367
R671 B.n591 B.n590 163.367
R672 B.n592 B.n591 163.367
R673 B.n592 B.n17 163.367
R674 B.n596 B.n17 163.367
R675 B.n597 B.n596 163.367
R676 B.n598 B.n597 163.367
R677 B.n598 B.n15 163.367
R678 B.n602 B.n15 163.367
R679 B.n603 B.n602 163.367
R680 B.n604 B.n603 163.367
R681 B.n604 B.n13 163.367
R682 B.n608 B.n13 163.367
R683 B.n609 B.n608 163.367
R684 B.n610 B.n609 163.367
R685 B.n610 B.n11 163.367
R686 B.n614 B.n11 163.367
R687 B.n615 B.n614 163.367
R688 B.n616 B.n615 163.367
R689 B.n616 B.n9 163.367
R690 B.n620 B.n9 163.367
R691 B.n621 B.n620 163.367
R692 B.n622 B.n621 163.367
R693 B.n622 B.n7 163.367
R694 B.n626 B.n7 163.367
R695 B.n627 B.n626 163.367
R696 B.n628 B.n627 163.367
R697 B.n628 B.n5 163.367
R698 B.n632 B.n5 163.367
R699 B.n633 B.n632 163.367
R700 B.n634 B.n633 163.367
R701 B.n634 B.n3 163.367
R702 B.n638 B.n3 163.367
R703 B.n639 B.n638 163.367
R704 B.n166 B.n2 163.367
R705 B.n167 B.n166 163.367
R706 B.n167 B.n164 163.367
R707 B.n171 B.n164 163.367
R708 B.n172 B.n171 163.367
R709 B.n173 B.n172 163.367
R710 B.n173 B.n162 163.367
R711 B.n177 B.n162 163.367
R712 B.n178 B.n177 163.367
R713 B.n179 B.n178 163.367
R714 B.n179 B.n160 163.367
R715 B.n183 B.n160 163.367
R716 B.n184 B.n183 163.367
R717 B.n185 B.n184 163.367
R718 B.n185 B.n158 163.367
R719 B.n189 B.n158 163.367
R720 B.n190 B.n189 163.367
R721 B.n191 B.n190 163.367
R722 B.n191 B.n156 163.367
R723 B.n195 B.n156 163.367
R724 B.n196 B.n195 163.367
R725 B.n197 B.n196 163.367
R726 B.n197 B.n154 163.367
R727 B.n201 B.n154 163.367
R728 B.n202 B.n201 163.367
R729 B.n203 B.n202 163.367
R730 B.n203 B.n152 163.367
R731 B.n207 B.n152 163.367
R732 B.n208 B.n207 163.367
R733 B.n209 B.n208 163.367
R734 B.n209 B.n150 163.367
R735 B.n213 B.n150 163.367
R736 B.n214 B.n213 163.367
R737 B.n215 B.n214 163.367
R738 B.n215 B.n148 163.367
R739 B.n219 B.n148 163.367
R740 B.n220 B.n219 163.367
R741 B.n221 B.n220 163.367
R742 B.n221 B.n146 163.367
R743 B.n225 B.n146 163.367
R744 B.n226 B.n225 163.367
R745 B.n227 B.n226 163.367
R746 B.n124 B.t5 109.302
R747 B.n48 B.t10 109.302
R748 B.n273 B.t8 109.293
R749 B.n41 B.t1 109.293
R750 B.n274 B.n273 59.5399
R751 B.n292 B.n124 59.5399
R752 B.n515 B.n48 59.5399
R753 B.n42 B.n41 59.5399
R754 B.n273 B.n272 58.7641
R755 B.n124 B.n123 58.7641
R756 B.n48 B.n47 58.7641
R757 B.n41 B.n40 58.7641
R758 B.n576 B.n575 37.62
R759 B.n468 B.n63 37.62
R760 B.n336 B.n107 37.62
R761 B.n229 B.n228 37.62
R762 B B.n641 18.0485
R763 B.n577 B.n576 10.6151
R764 B.n577 B.n22 10.6151
R765 B.n581 B.n22 10.6151
R766 B.n582 B.n581 10.6151
R767 B.n583 B.n582 10.6151
R768 B.n583 B.n20 10.6151
R769 B.n587 B.n20 10.6151
R770 B.n588 B.n587 10.6151
R771 B.n589 B.n588 10.6151
R772 B.n589 B.n18 10.6151
R773 B.n593 B.n18 10.6151
R774 B.n594 B.n593 10.6151
R775 B.n595 B.n594 10.6151
R776 B.n595 B.n16 10.6151
R777 B.n599 B.n16 10.6151
R778 B.n600 B.n599 10.6151
R779 B.n601 B.n600 10.6151
R780 B.n601 B.n14 10.6151
R781 B.n605 B.n14 10.6151
R782 B.n606 B.n605 10.6151
R783 B.n607 B.n606 10.6151
R784 B.n607 B.n12 10.6151
R785 B.n611 B.n12 10.6151
R786 B.n612 B.n611 10.6151
R787 B.n613 B.n612 10.6151
R788 B.n613 B.n10 10.6151
R789 B.n617 B.n10 10.6151
R790 B.n618 B.n617 10.6151
R791 B.n619 B.n618 10.6151
R792 B.n619 B.n8 10.6151
R793 B.n623 B.n8 10.6151
R794 B.n624 B.n623 10.6151
R795 B.n625 B.n624 10.6151
R796 B.n625 B.n6 10.6151
R797 B.n629 B.n6 10.6151
R798 B.n630 B.n629 10.6151
R799 B.n631 B.n630 10.6151
R800 B.n631 B.n4 10.6151
R801 B.n635 B.n4 10.6151
R802 B.n636 B.n635 10.6151
R803 B.n637 B.n636 10.6151
R804 B.n637 B.n0 10.6151
R805 B.n575 B.n24 10.6151
R806 B.n571 B.n24 10.6151
R807 B.n571 B.n570 10.6151
R808 B.n570 B.n569 10.6151
R809 B.n569 B.n26 10.6151
R810 B.n565 B.n26 10.6151
R811 B.n565 B.n564 10.6151
R812 B.n564 B.n563 10.6151
R813 B.n563 B.n28 10.6151
R814 B.n559 B.n28 10.6151
R815 B.n559 B.n558 10.6151
R816 B.n558 B.n557 10.6151
R817 B.n557 B.n30 10.6151
R818 B.n553 B.n30 10.6151
R819 B.n553 B.n552 10.6151
R820 B.n552 B.n551 10.6151
R821 B.n551 B.n32 10.6151
R822 B.n547 B.n32 10.6151
R823 B.n547 B.n546 10.6151
R824 B.n546 B.n545 10.6151
R825 B.n545 B.n34 10.6151
R826 B.n541 B.n34 10.6151
R827 B.n541 B.n540 10.6151
R828 B.n540 B.n539 10.6151
R829 B.n539 B.n36 10.6151
R830 B.n535 B.n36 10.6151
R831 B.n535 B.n534 10.6151
R832 B.n534 B.n533 10.6151
R833 B.n533 B.n38 10.6151
R834 B.n529 B.n528 10.6151
R835 B.n528 B.n527 10.6151
R836 B.n527 B.n43 10.6151
R837 B.n523 B.n43 10.6151
R838 B.n523 B.n522 10.6151
R839 B.n522 B.n521 10.6151
R840 B.n521 B.n45 10.6151
R841 B.n517 B.n45 10.6151
R842 B.n517 B.n516 10.6151
R843 B.n514 B.n49 10.6151
R844 B.n510 B.n49 10.6151
R845 B.n510 B.n509 10.6151
R846 B.n509 B.n508 10.6151
R847 B.n508 B.n51 10.6151
R848 B.n504 B.n51 10.6151
R849 B.n504 B.n503 10.6151
R850 B.n503 B.n502 10.6151
R851 B.n502 B.n53 10.6151
R852 B.n498 B.n53 10.6151
R853 B.n498 B.n497 10.6151
R854 B.n497 B.n496 10.6151
R855 B.n496 B.n55 10.6151
R856 B.n492 B.n55 10.6151
R857 B.n492 B.n491 10.6151
R858 B.n491 B.n490 10.6151
R859 B.n490 B.n57 10.6151
R860 B.n486 B.n57 10.6151
R861 B.n486 B.n485 10.6151
R862 B.n485 B.n484 10.6151
R863 B.n484 B.n59 10.6151
R864 B.n480 B.n59 10.6151
R865 B.n480 B.n479 10.6151
R866 B.n479 B.n478 10.6151
R867 B.n478 B.n61 10.6151
R868 B.n474 B.n61 10.6151
R869 B.n474 B.n473 10.6151
R870 B.n473 B.n472 10.6151
R871 B.n472 B.n63 10.6151
R872 B.n468 B.n467 10.6151
R873 B.n467 B.n466 10.6151
R874 B.n466 B.n65 10.6151
R875 B.n462 B.n65 10.6151
R876 B.n462 B.n461 10.6151
R877 B.n461 B.n460 10.6151
R878 B.n460 B.n67 10.6151
R879 B.n456 B.n67 10.6151
R880 B.n456 B.n455 10.6151
R881 B.n455 B.n454 10.6151
R882 B.n454 B.n69 10.6151
R883 B.n450 B.n69 10.6151
R884 B.n450 B.n449 10.6151
R885 B.n449 B.n448 10.6151
R886 B.n448 B.n71 10.6151
R887 B.n444 B.n71 10.6151
R888 B.n444 B.n443 10.6151
R889 B.n443 B.n442 10.6151
R890 B.n442 B.n73 10.6151
R891 B.n438 B.n73 10.6151
R892 B.n438 B.n437 10.6151
R893 B.n437 B.n436 10.6151
R894 B.n436 B.n75 10.6151
R895 B.n432 B.n75 10.6151
R896 B.n432 B.n431 10.6151
R897 B.n431 B.n430 10.6151
R898 B.n430 B.n77 10.6151
R899 B.n426 B.n77 10.6151
R900 B.n426 B.n425 10.6151
R901 B.n425 B.n424 10.6151
R902 B.n424 B.n79 10.6151
R903 B.n420 B.n79 10.6151
R904 B.n420 B.n419 10.6151
R905 B.n419 B.n418 10.6151
R906 B.n418 B.n81 10.6151
R907 B.n414 B.n81 10.6151
R908 B.n414 B.n413 10.6151
R909 B.n413 B.n412 10.6151
R910 B.n412 B.n83 10.6151
R911 B.n408 B.n83 10.6151
R912 B.n408 B.n407 10.6151
R913 B.n407 B.n406 10.6151
R914 B.n406 B.n85 10.6151
R915 B.n402 B.n85 10.6151
R916 B.n402 B.n401 10.6151
R917 B.n401 B.n400 10.6151
R918 B.n400 B.n87 10.6151
R919 B.n396 B.n87 10.6151
R920 B.n396 B.n395 10.6151
R921 B.n395 B.n394 10.6151
R922 B.n394 B.n89 10.6151
R923 B.n390 B.n89 10.6151
R924 B.n390 B.n389 10.6151
R925 B.n389 B.n388 10.6151
R926 B.n388 B.n91 10.6151
R927 B.n384 B.n91 10.6151
R928 B.n384 B.n383 10.6151
R929 B.n383 B.n382 10.6151
R930 B.n382 B.n93 10.6151
R931 B.n378 B.n93 10.6151
R932 B.n378 B.n377 10.6151
R933 B.n377 B.n376 10.6151
R934 B.n376 B.n95 10.6151
R935 B.n372 B.n95 10.6151
R936 B.n372 B.n371 10.6151
R937 B.n371 B.n370 10.6151
R938 B.n370 B.n97 10.6151
R939 B.n366 B.n97 10.6151
R940 B.n366 B.n365 10.6151
R941 B.n365 B.n364 10.6151
R942 B.n364 B.n99 10.6151
R943 B.n360 B.n99 10.6151
R944 B.n360 B.n359 10.6151
R945 B.n359 B.n358 10.6151
R946 B.n358 B.n101 10.6151
R947 B.n354 B.n101 10.6151
R948 B.n354 B.n353 10.6151
R949 B.n353 B.n352 10.6151
R950 B.n352 B.n103 10.6151
R951 B.n348 B.n103 10.6151
R952 B.n348 B.n347 10.6151
R953 B.n347 B.n346 10.6151
R954 B.n346 B.n105 10.6151
R955 B.n342 B.n105 10.6151
R956 B.n342 B.n341 10.6151
R957 B.n341 B.n340 10.6151
R958 B.n340 B.n107 10.6151
R959 B.n165 B.n1 10.6151
R960 B.n168 B.n165 10.6151
R961 B.n169 B.n168 10.6151
R962 B.n170 B.n169 10.6151
R963 B.n170 B.n163 10.6151
R964 B.n174 B.n163 10.6151
R965 B.n175 B.n174 10.6151
R966 B.n176 B.n175 10.6151
R967 B.n176 B.n161 10.6151
R968 B.n180 B.n161 10.6151
R969 B.n181 B.n180 10.6151
R970 B.n182 B.n181 10.6151
R971 B.n182 B.n159 10.6151
R972 B.n186 B.n159 10.6151
R973 B.n187 B.n186 10.6151
R974 B.n188 B.n187 10.6151
R975 B.n188 B.n157 10.6151
R976 B.n192 B.n157 10.6151
R977 B.n193 B.n192 10.6151
R978 B.n194 B.n193 10.6151
R979 B.n194 B.n155 10.6151
R980 B.n198 B.n155 10.6151
R981 B.n199 B.n198 10.6151
R982 B.n200 B.n199 10.6151
R983 B.n200 B.n153 10.6151
R984 B.n204 B.n153 10.6151
R985 B.n205 B.n204 10.6151
R986 B.n206 B.n205 10.6151
R987 B.n206 B.n151 10.6151
R988 B.n210 B.n151 10.6151
R989 B.n211 B.n210 10.6151
R990 B.n212 B.n211 10.6151
R991 B.n212 B.n149 10.6151
R992 B.n216 B.n149 10.6151
R993 B.n217 B.n216 10.6151
R994 B.n218 B.n217 10.6151
R995 B.n218 B.n147 10.6151
R996 B.n222 B.n147 10.6151
R997 B.n223 B.n222 10.6151
R998 B.n224 B.n223 10.6151
R999 B.n224 B.n145 10.6151
R1000 B.n228 B.n145 10.6151
R1001 B.n230 B.n229 10.6151
R1002 B.n230 B.n143 10.6151
R1003 B.n234 B.n143 10.6151
R1004 B.n235 B.n234 10.6151
R1005 B.n236 B.n235 10.6151
R1006 B.n236 B.n141 10.6151
R1007 B.n240 B.n141 10.6151
R1008 B.n241 B.n240 10.6151
R1009 B.n242 B.n241 10.6151
R1010 B.n242 B.n139 10.6151
R1011 B.n246 B.n139 10.6151
R1012 B.n247 B.n246 10.6151
R1013 B.n248 B.n247 10.6151
R1014 B.n248 B.n137 10.6151
R1015 B.n252 B.n137 10.6151
R1016 B.n253 B.n252 10.6151
R1017 B.n254 B.n253 10.6151
R1018 B.n254 B.n135 10.6151
R1019 B.n258 B.n135 10.6151
R1020 B.n259 B.n258 10.6151
R1021 B.n260 B.n259 10.6151
R1022 B.n260 B.n133 10.6151
R1023 B.n264 B.n133 10.6151
R1024 B.n265 B.n264 10.6151
R1025 B.n266 B.n265 10.6151
R1026 B.n266 B.n131 10.6151
R1027 B.n270 B.n131 10.6151
R1028 B.n271 B.n270 10.6151
R1029 B.n275 B.n271 10.6151
R1030 B.n279 B.n129 10.6151
R1031 B.n280 B.n279 10.6151
R1032 B.n281 B.n280 10.6151
R1033 B.n281 B.n127 10.6151
R1034 B.n285 B.n127 10.6151
R1035 B.n286 B.n285 10.6151
R1036 B.n287 B.n286 10.6151
R1037 B.n287 B.n125 10.6151
R1038 B.n291 B.n125 10.6151
R1039 B.n294 B.n293 10.6151
R1040 B.n294 B.n121 10.6151
R1041 B.n298 B.n121 10.6151
R1042 B.n299 B.n298 10.6151
R1043 B.n300 B.n299 10.6151
R1044 B.n300 B.n119 10.6151
R1045 B.n304 B.n119 10.6151
R1046 B.n305 B.n304 10.6151
R1047 B.n306 B.n305 10.6151
R1048 B.n306 B.n117 10.6151
R1049 B.n310 B.n117 10.6151
R1050 B.n311 B.n310 10.6151
R1051 B.n312 B.n311 10.6151
R1052 B.n312 B.n115 10.6151
R1053 B.n316 B.n115 10.6151
R1054 B.n317 B.n316 10.6151
R1055 B.n318 B.n317 10.6151
R1056 B.n318 B.n113 10.6151
R1057 B.n322 B.n113 10.6151
R1058 B.n323 B.n322 10.6151
R1059 B.n324 B.n323 10.6151
R1060 B.n324 B.n111 10.6151
R1061 B.n328 B.n111 10.6151
R1062 B.n329 B.n328 10.6151
R1063 B.n330 B.n329 10.6151
R1064 B.n330 B.n109 10.6151
R1065 B.n334 B.n109 10.6151
R1066 B.n335 B.n334 10.6151
R1067 B.n336 B.n335 10.6151
R1068 B.n42 B.n38 9.36635
R1069 B.n515 B.n514 9.36635
R1070 B.n275 B.n274 9.36635
R1071 B.n293 B.n292 9.36635
R1072 B.n641 B.n0 8.11757
R1073 B.n641 B.n1 8.11757
R1074 B.n529 B.n42 1.24928
R1075 B.n516 B.n515 1.24928
R1076 B.n274 B.n129 1.24928
R1077 B.n292 B.n291 1.24928
R1078 VN.n29 VN.n16 161.3
R1079 VN.n28 VN.n27 161.3
R1080 VN.n26 VN.n17 161.3
R1081 VN.n25 VN.n24 161.3
R1082 VN.n23 VN.n18 161.3
R1083 VN.n22 VN.n21 161.3
R1084 VN.n13 VN.n0 161.3
R1085 VN.n12 VN.n11 161.3
R1086 VN.n10 VN.n1 161.3
R1087 VN.n9 VN.n8 161.3
R1088 VN.n7 VN.n2 161.3
R1089 VN.n6 VN.n5 161.3
R1090 VN.n15 VN.n14 109.433
R1091 VN.n31 VN.n30 109.433
R1092 VN.n4 VN.t3 106.007
R1093 VN.n20 VN.t2 106.007
R1094 VN.n3 VN.t1 73.1931
R1095 VN.n14 VN.t4 73.1931
R1096 VN.n19 VN.t5 73.1931
R1097 VN.n30 VN.t0 73.1931
R1098 VN.n20 VN.n19 49.0351
R1099 VN.n4 VN.n3 49.0351
R1100 VN VN.n31 46.3808
R1101 VN.n8 VN.n1 42.0302
R1102 VN.n24 VN.n17 42.0302
R1103 VN.n8 VN.n7 39.1239
R1104 VN.n24 VN.n23 39.1239
R1105 VN.n6 VN.n3 24.5923
R1106 VN.n7 VN.n6 24.5923
R1107 VN.n12 VN.n1 24.5923
R1108 VN.n13 VN.n12 24.5923
R1109 VN.n23 VN.n22 24.5923
R1110 VN.n22 VN.n19 24.5923
R1111 VN.n29 VN.n28 24.5923
R1112 VN.n28 VN.n17 24.5923
R1113 VN.n21 VN.n20 5.10935
R1114 VN.n5 VN.n4 5.10935
R1115 VN.n14 VN.n13 1.47601
R1116 VN.n30 VN.n29 1.47601
R1117 VN.n31 VN.n16 0.278335
R1118 VN.n15 VN.n0 0.278335
R1119 VN.n27 VN.n16 0.189894
R1120 VN.n27 VN.n26 0.189894
R1121 VN.n26 VN.n25 0.189894
R1122 VN.n25 VN.n18 0.189894
R1123 VN.n21 VN.n18 0.189894
R1124 VN.n5 VN.n2 0.189894
R1125 VN.n9 VN.n2 0.189894
R1126 VN.n10 VN.n9 0.189894
R1127 VN.n11 VN.n10 0.189894
R1128 VN.n11 VN.n0 0.189894
R1129 VN VN.n15 0.153485
R1130 VDD2.n1 VDD2.t2 87.9282
R1131 VDD2.n2 VDD2.t5 86.0246
R1132 VDD2.n1 VDD2.n0 82.658
R1133 VDD2 VDD2.n3 82.6553
R1134 VDD2.n2 VDD2.n1 39.2735
R1135 VDD2.n3 VDD2.t0 3.96452
R1136 VDD2.n3 VDD2.t3 3.96452
R1137 VDD2.n0 VDD2.t4 3.96452
R1138 VDD2.n0 VDD2.t1 3.96452
R1139 VDD2 VDD2.n2 2.01774
C0 VTAIL w_n3394_n2608# 2.44867f
C1 VN w_n3394_n2608# 6.38671f
C2 VDD1 w_n3394_n2608# 2.04903f
C3 VP VTAIL 5.11765f
C4 VDD2 w_n3394_n2608# 2.13727f
C5 VP VN 6.31807f
C6 VP VDD1 5.06585f
C7 B w_n3394_n2608# 8.748981f
C8 VN VTAIL 5.10343f
C9 VDD2 VP 0.466645f
C10 VDD1 VTAIL 6.39025f
C11 VDD2 VTAIL 6.44271f
C12 VDD1 VN 0.151018f
C13 VP B 1.88105f
C14 VDD2 VN 4.75275f
C15 VTAIL B 2.87759f
C16 VDD2 VDD1 1.4442f
C17 VN B 1.14747f
C18 VDD1 B 1.81818f
C19 VDD2 B 1.89467f
C20 VP w_n3394_n2608# 6.82578f
C21 VDD2 VSUBS 1.695576f
C22 VDD1 VSUBS 2.182886f
C23 VTAIL VSUBS 1.075086f
C24 VN VSUBS 5.81331f
C25 VP VSUBS 2.864029f
C26 B VSUBS 4.41458f
C27 w_n3394_n2608# VSUBS 0.109762p
C28 VDD2.t2 VSUBS 1.60864f
C29 VDD2.t4 VSUBS 0.166467f
C30 VDD2.t1 VSUBS 0.166467f
C31 VDD2.n0 VSUBS 1.21412f
C32 VDD2.n1 VSUBS 3.24965f
C33 VDD2.t5 VSUBS 1.59398f
C34 VDD2.n2 VSUBS 2.82638f
C35 VDD2.t0 VSUBS 0.166467f
C36 VDD2.t3 VSUBS 0.166467f
C37 VDD2.n3 VSUBS 1.21408f
C38 VN.n0 VSUBS 0.044283f
C39 VN.t4 VSUBS 1.99944f
C40 VN.n1 VSUBS 0.065862f
C41 VN.n2 VSUBS 0.03359f
C42 VN.t1 VSUBS 1.99944f
C43 VN.n3 VSUBS 0.843334f
C44 VN.t3 VSUBS 2.29124f
C45 VN.n4 VSUBS 0.796528f
C46 VN.n5 VSUBS 0.348749f
C47 VN.n6 VSUBS 0.06229f
C48 VN.n7 VSUBS 0.066859f
C49 VN.n8 VSUBS 0.027226f
C50 VN.n9 VSUBS 0.03359f
C51 VN.n10 VSUBS 0.03359f
C52 VN.n11 VSUBS 0.03359f
C53 VN.n12 VSUBS 0.06229f
C54 VN.n13 VSUBS 0.033384f
C55 VN.n14 VSUBS 0.826725f
C56 VN.n15 VSUBS 0.062177f
C57 VN.n16 VSUBS 0.044283f
C58 VN.t0 VSUBS 1.99944f
C59 VN.n17 VSUBS 0.065862f
C60 VN.n18 VSUBS 0.03359f
C61 VN.t5 VSUBS 1.99944f
C62 VN.n19 VSUBS 0.843334f
C63 VN.t2 VSUBS 2.29124f
C64 VN.n20 VSUBS 0.796528f
C65 VN.n21 VSUBS 0.348749f
C66 VN.n22 VSUBS 0.06229f
C67 VN.n23 VSUBS 0.066859f
C68 VN.n24 VSUBS 0.027226f
C69 VN.n25 VSUBS 0.03359f
C70 VN.n26 VSUBS 0.03359f
C71 VN.n27 VSUBS 0.03359f
C72 VN.n28 VSUBS 0.06229f
C73 VN.n29 VSUBS 0.033384f
C74 VN.n30 VSUBS 0.826725f
C75 VN.n31 VSUBS 1.67954f
C76 B.n0 VSUBS 0.006072f
C77 B.n1 VSUBS 0.006072f
C78 B.n2 VSUBS 0.00898f
C79 B.n3 VSUBS 0.006881f
C80 B.n4 VSUBS 0.006881f
C81 B.n5 VSUBS 0.006881f
C82 B.n6 VSUBS 0.006881f
C83 B.n7 VSUBS 0.006881f
C84 B.n8 VSUBS 0.006881f
C85 B.n9 VSUBS 0.006881f
C86 B.n10 VSUBS 0.006881f
C87 B.n11 VSUBS 0.006881f
C88 B.n12 VSUBS 0.006881f
C89 B.n13 VSUBS 0.006881f
C90 B.n14 VSUBS 0.006881f
C91 B.n15 VSUBS 0.006881f
C92 B.n16 VSUBS 0.006881f
C93 B.n17 VSUBS 0.006881f
C94 B.n18 VSUBS 0.006881f
C95 B.n19 VSUBS 0.006881f
C96 B.n20 VSUBS 0.006881f
C97 B.n21 VSUBS 0.006881f
C98 B.n22 VSUBS 0.006881f
C99 B.n23 VSUBS 0.017356f
C100 B.n24 VSUBS 0.006881f
C101 B.n25 VSUBS 0.006881f
C102 B.n26 VSUBS 0.006881f
C103 B.n27 VSUBS 0.006881f
C104 B.n28 VSUBS 0.006881f
C105 B.n29 VSUBS 0.006881f
C106 B.n30 VSUBS 0.006881f
C107 B.n31 VSUBS 0.006881f
C108 B.n32 VSUBS 0.006881f
C109 B.n33 VSUBS 0.006881f
C110 B.n34 VSUBS 0.006881f
C111 B.n35 VSUBS 0.006881f
C112 B.n36 VSUBS 0.006881f
C113 B.n37 VSUBS 0.006881f
C114 B.n38 VSUBS 0.006476f
C115 B.n39 VSUBS 0.006881f
C116 B.t1 VSUBS 0.249771f
C117 B.t2 VSUBS 0.271021f
C118 B.t0 VSUBS 1.01561f
C119 B.n40 VSUBS 0.14687f
C120 B.n41 VSUBS 0.070585f
C121 B.n42 VSUBS 0.015943f
C122 B.n43 VSUBS 0.006881f
C123 B.n44 VSUBS 0.006881f
C124 B.n45 VSUBS 0.006881f
C125 B.n46 VSUBS 0.006881f
C126 B.t10 VSUBS 0.249769f
C127 B.t11 VSUBS 0.271018f
C128 B.t9 VSUBS 1.01561f
C129 B.n47 VSUBS 0.146873f
C130 B.n48 VSUBS 0.070588f
C131 B.n49 VSUBS 0.006881f
C132 B.n50 VSUBS 0.006881f
C133 B.n51 VSUBS 0.006881f
C134 B.n52 VSUBS 0.006881f
C135 B.n53 VSUBS 0.006881f
C136 B.n54 VSUBS 0.006881f
C137 B.n55 VSUBS 0.006881f
C138 B.n56 VSUBS 0.006881f
C139 B.n57 VSUBS 0.006881f
C140 B.n58 VSUBS 0.006881f
C141 B.n59 VSUBS 0.006881f
C142 B.n60 VSUBS 0.006881f
C143 B.n61 VSUBS 0.006881f
C144 B.n62 VSUBS 0.006881f
C145 B.n63 VSUBS 0.018062f
C146 B.n64 VSUBS 0.006881f
C147 B.n65 VSUBS 0.006881f
C148 B.n66 VSUBS 0.006881f
C149 B.n67 VSUBS 0.006881f
C150 B.n68 VSUBS 0.006881f
C151 B.n69 VSUBS 0.006881f
C152 B.n70 VSUBS 0.006881f
C153 B.n71 VSUBS 0.006881f
C154 B.n72 VSUBS 0.006881f
C155 B.n73 VSUBS 0.006881f
C156 B.n74 VSUBS 0.006881f
C157 B.n75 VSUBS 0.006881f
C158 B.n76 VSUBS 0.006881f
C159 B.n77 VSUBS 0.006881f
C160 B.n78 VSUBS 0.006881f
C161 B.n79 VSUBS 0.006881f
C162 B.n80 VSUBS 0.006881f
C163 B.n81 VSUBS 0.006881f
C164 B.n82 VSUBS 0.006881f
C165 B.n83 VSUBS 0.006881f
C166 B.n84 VSUBS 0.006881f
C167 B.n85 VSUBS 0.006881f
C168 B.n86 VSUBS 0.006881f
C169 B.n87 VSUBS 0.006881f
C170 B.n88 VSUBS 0.006881f
C171 B.n89 VSUBS 0.006881f
C172 B.n90 VSUBS 0.006881f
C173 B.n91 VSUBS 0.006881f
C174 B.n92 VSUBS 0.006881f
C175 B.n93 VSUBS 0.006881f
C176 B.n94 VSUBS 0.006881f
C177 B.n95 VSUBS 0.006881f
C178 B.n96 VSUBS 0.006881f
C179 B.n97 VSUBS 0.006881f
C180 B.n98 VSUBS 0.006881f
C181 B.n99 VSUBS 0.006881f
C182 B.n100 VSUBS 0.006881f
C183 B.n101 VSUBS 0.006881f
C184 B.n102 VSUBS 0.006881f
C185 B.n103 VSUBS 0.006881f
C186 B.n104 VSUBS 0.006881f
C187 B.n105 VSUBS 0.006881f
C188 B.n106 VSUBS 0.006881f
C189 B.n107 VSUBS 0.018062f
C190 B.n108 VSUBS 0.006881f
C191 B.n109 VSUBS 0.006881f
C192 B.n110 VSUBS 0.006881f
C193 B.n111 VSUBS 0.006881f
C194 B.n112 VSUBS 0.006881f
C195 B.n113 VSUBS 0.006881f
C196 B.n114 VSUBS 0.006881f
C197 B.n115 VSUBS 0.006881f
C198 B.n116 VSUBS 0.006881f
C199 B.n117 VSUBS 0.006881f
C200 B.n118 VSUBS 0.006881f
C201 B.n119 VSUBS 0.006881f
C202 B.n120 VSUBS 0.006881f
C203 B.n121 VSUBS 0.006881f
C204 B.n122 VSUBS 0.006881f
C205 B.t5 VSUBS 0.249769f
C206 B.t4 VSUBS 0.271018f
C207 B.t3 VSUBS 1.01561f
C208 B.n123 VSUBS 0.146873f
C209 B.n124 VSUBS 0.070588f
C210 B.n125 VSUBS 0.006881f
C211 B.n126 VSUBS 0.006881f
C212 B.n127 VSUBS 0.006881f
C213 B.n128 VSUBS 0.006881f
C214 B.n129 VSUBS 0.003845f
C215 B.n130 VSUBS 0.006881f
C216 B.n131 VSUBS 0.006881f
C217 B.n132 VSUBS 0.006881f
C218 B.n133 VSUBS 0.006881f
C219 B.n134 VSUBS 0.006881f
C220 B.n135 VSUBS 0.006881f
C221 B.n136 VSUBS 0.006881f
C222 B.n137 VSUBS 0.006881f
C223 B.n138 VSUBS 0.006881f
C224 B.n139 VSUBS 0.006881f
C225 B.n140 VSUBS 0.006881f
C226 B.n141 VSUBS 0.006881f
C227 B.n142 VSUBS 0.006881f
C228 B.n143 VSUBS 0.006881f
C229 B.n144 VSUBS 0.018062f
C230 B.n145 VSUBS 0.006881f
C231 B.n146 VSUBS 0.006881f
C232 B.n147 VSUBS 0.006881f
C233 B.n148 VSUBS 0.006881f
C234 B.n149 VSUBS 0.006881f
C235 B.n150 VSUBS 0.006881f
C236 B.n151 VSUBS 0.006881f
C237 B.n152 VSUBS 0.006881f
C238 B.n153 VSUBS 0.006881f
C239 B.n154 VSUBS 0.006881f
C240 B.n155 VSUBS 0.006881f
C241 B.n156 VSUBS 0.006881f
C242 B.n157 VSUBS 0.006881f
C243 B.n158 VSUBS 0.006881f
C244 B.n159 VSUBS 0.006881f
C245 B.n160 VSUBS 0.006881f
C246 B.n161 VSUBS 0.006881f
C247 B.n162 VSUBS 0.006881f
C248 B.n163 VSUBS 0.006881f
C249 B.n164 VSUBS 0.006881f
C250 B.n165 VSUBS 0.006881f
C251 B.n166 VSUBS 0.006881f
C252 B.n167 VSUBS 0.006881f
C253 B.n168 VSUBS 0.006881f
C254 B.n169 VSUBS 0.006881f
C255 B.n170 VSUBS 0.006881f
C256 B.n171 VSUBS 0.006881f
C257 B.n172 VSUBS 0.006881f
C258 B.n173 VSUBS 0.006881f
C259 B.n174 VSUBS 0.006881f
C260 B.n175 VSUBS 0.006881f
C261 B.n176 VSUBS 0.006881f
C262 B.n177 VSUBS 0.006881f
C263 B.n178 VSUBS 0.006881f
C264 B.n179 VSUBS 0.006881f
C265 B.n180 VSUBS 0.006881f
C266 B.n181 VSUBS 0.006881f
C267 B.n182 VSUBS 0.006881f
C268 B.n183 VSUBS 0.006881f
C269 B.n184 VSUBS 0.006881f
C270 B.n185 VSUBS 0.006881f
C271 B.n186 VSUBS 0.006881f
C272 B.n187 VSUBS 0.006881f
C273 B.n188 VSUBS 0.006881f
C274 B.n189 VSUBS 0.006881f
C275 B.n190 VSUBS 0.006881f
C276 B.n191 VSUBS 0.006881f
C277 B.n192 VSUBS 0.006881f
C278 B.n193 VSUBS 0.006881f
C279 B.n194 VSUBS 0.006881f
C280 B.n195 VSUBS 0.006881f
C281 B.n196 VSUBS 0.006881f
C282 B.n197 VSUBS 0.006881f
C283 B.n198 VSUBS 0.006881f
C284 B.n199 VSUBS 0.006881f
C285 B.n200 VSUBS 0.006881f
C286 B.n201 VSUBS 0.006881f
C287 B.n202 VSUBS 0.006881f
C288 B.n203 VSUBS 0.006881f
C289 B.n204 VSUBS 0.006881f
C290 B.n205 VSUBS 0.006881f
C291 B.n206 VSUBS 0.006881f
C292 B.n207 VSUBS 0.006881f
C293 B.n208 VSUBS 0.006881f
C294 B.n209 VSUBS 0.006881f
C295 B.n210 VSUBS 0.006881f
C296 B.n211 VSUBS 0.006881f
C297 B.n212 VSUBS 0.006881f
C298 B.n213 VSUBS 0.006881f
C299 B.n214 VSUBS 0.006881f
C300 B.n215 VSUBS 0.006881f
C301 B.n216 VSUBS 0.006881f
C302 B.n217 VSUBS 0.006881f
C303 B.n218 VSUBS 0.006881f
C304 B.n219 VSUBS 0.006881f
C305 B.n220 VSUBS 0.006881f
C306 B.n221 VSUBS 0.006881f
C307 B.n222 VSUBS 0.006881f
C308 B.n223 VSUBS 0.006881f
C309 B.n224 VSUBS 0.006881f
C310 B.n225 VSUBS 0.006881f
C311 B.n226 VSUBS 0.006881f
C312 B.n227 VSUBS 0.017356f
C313 B.n228 VSUBS 0.017356f
C314 B.n229 VSUBS 0.018062f
C315 B.n230 VSUBS 0.006881f
C316 B.n231 VSUBS 0.006881f
C317 B.n232 VSUBS 0.006881f
C318 B.n233 VSUBS 0.006881f
C319 B.n234 VSUBS 0.006881f
C320 B.n235 VSUBS 0.006881f
C321 B.n236 VSUBS 0.006881f
C322 B.n237 VSUBS 0.006881f
C323 B.n238 VSUBS 0.006881f
C324 B.n239 VSUBS 0.006881f
C325 B.n240 VSUBS 0.006881f
C326 B.n241 VSUBS 0.006881f
C327 B.n242 VSUBS 0.006881f
C328 B.n243 VSUBS 0.006881f
C329 B.n244 VSUBS 0.006881f
C330 B.n245 VSUBS 0.006881f
C331 B.n246 VSUBS 0.006881f
C332 B.n247 VSUBS 0.006881f
C333 B.n248 VSUBS 0.006881f
C334 B.n249 VSUBS 0.006881f
C335 B.n250 VSUBS 0.006881f
C336 B.n251 VSUBS 0.006881f
C337 B.n252 VSUBS 0.006881f
C338 B.n253 VSUBS 0.006881f
C339 B.n254 VSUBS 0.006881f
C340 B.n255 VSUBS 0.006881f
C341 B.n256 VSUBS 0.006881f
C342 B.n257 VSUBS 0.006881f
C343 B.n258 VSUBS 0.006881f
C344 B.n259 VSUBS 0.006881f
C345 B.n260 VSUBS 0.006881f
C346 B.n261 VSUBS 0.006881f
C347 B.n262 VSUBS 0.006881f
C348 B.n263 VSUBS 0.006881f
C349 B.n264 VSUBS 0.006881f
C350 B.n265 VSUBS 0.006881f
C351 B.n266 VSUBS 0.006881f
C352 B.n267 VSUBS 0.006881f
C353 B.n268 VSUBS 0.006881f
C354 B.n269 VSUBS 0.006881f
C355 B.n270 VSUBS 0.006881f
C356 B.n271 VSUBS 0.006881f
C357 B.t8 VSUBS 0.249771f
C358 B.t7 VSUBS 0.271021f
C359 B.t6 VSUBS 1.01561f
C360 B.n272 VSUBS 0.14687f
C361 B.n273 VSUBS 0.070585f
C362 B.n274 VSUBS 0.015943f
C363 B.n275 VSUBS 0.006476f
C364 B.n276 VSUBS 0.006881f
C365 B.n277 VSUBS 0.006881f
C366 B.n278 VSUBS 0.006881f
C367 B.n279 VSUBS 0.006881f
C368 B.n280 VSUBS 0.006881f
C369 B.n281 VSUBS 0.006881f
C370 B.n282 VSUBS 0.006881f
C371 B.n283 VSUBS 0.006881f
C372 B.n284 VSUBS 0.006881f
C373 B.n285 VSUBS 0.006881f
C374 B.n286 VSUBS 0.006881f
C375 B.n287 VSUBS 0.006881f
C376 B.n288 VSUBS 0.006881f
C377 B.n289 VSUBS 0.006881f
C378 B.n290 VSUBS 0.006881f
C379 B.n291 VSUBS 0.003845f
C380 B.n292 VSUBS 0.015943f
C381 B.n293 VSUBS 0.006476f
C382 B.n294 VSUBS 0.006881f
C383 B.n295 VSUBS 0.006881f
C384 B.n296 VSUBS 0.006881f
C385 B.n297 VSUBS 0.006881f
C386 B.n298 VSUBS 0.006881f
C387 B.n299 VSUBS 0.006881f
C388 B.n300 VSUBS 0.006881f
C389 B.n301 VSUBS 0.006881f
C390 B.n302 VSUBS 0.006881f
C391 B.n303 VSUBS 0.006881f
C392 B.n304 VSUBS 0.006881f
C393 B.n305 VSUBS 0.006881f
C394 B.n306 VSUBS 0.006881f
C395 B.n307 VSUBS 0.006881f
C396 B.n308 VSUBS 0.006881f
C397 B.n309 VSUBS 0.006881f
C398 B.n310 VSUBS 0.006881f
C399 B.n311 VSUBS 0.006881f
C400 B.n312 VSUBS 0.006881f
C401 B.n313 VSUBS 0.006881f
C402 B.n314 VSUBS 0.006881f
C403 B.n315 VSUBS 0.006881f
C404 B.n316 VSUBS 0.006881f
C405 B.n317 VSUBS 0.006881f
C406 B.n318 VSUBS 0.006881f
C407 B.n319 VSUBS 0.006881f
C408 B.n320 VSUBS 0.006881f
C409 B.n321 VSUBS 0.006881f
C410 B.n322 VSUBS 0.006881f
C411 B.n323 VSUBS 0.006881f
C412 B.n324 VSUBS 0.006881f
C413 B.n325 VSUBS 0.006881f
C414 B.n326 VSUBS 0.006881f
C415 B.n327 VSUBS 0.006881f
C416 B.n328 VSUBS 0.006881f
C417 B.n329 VSUBS 0.006881f
C418 B.n330 VSUBS 0.006881f
C419 B.n331 VSUBS 0.006881f
C420 B.n332 VSUBS 0.006881f
C421 B.n333 VSUBS 0.006881f
C422 B.n334 VSUBS 0.006881f
C423 B.n335 VSUBS 0.006881f
C424 B.n336 VSUBS 0.017356f
C425 B.n337 VSUBS 0.018062f
C426 B.n338 VSUBS 0.017356f
C427 B.n339 VSUBS 0.006881f
C428 B.n340 VSUBS 0.006881f
C429 B.n341 VSUBS 0.006881f
C430 B.n342 VSUBS 0.006881f
C431 B.n343 VSUBS 0.006881f
C432 B.n344 VSUBS 0.006881f
C433 B.n345 VSUBS 0.006881f
C434 B.n346 VSUBS 0.006881f
C435 B.n347 VSUBS 0.006881f
C436 B.n348 VSUBS 0.006881f
C437 B.n349 VSUBS 0.006881f
C438 B.n350 VSUBS 0.006881f
C439 B.n351 VSUBS 0.006881f
C440 B.n352 VSUBS 0.006881f
C441 B.n353 VSUBS 0.006881f
C442 B.n354 VSUBS 0.006881f
C443 B.n355 VSUBS 0.006881f
C444 B.n356 VSUBS 0.006881f
C445 B.n357 VSUBS 0.006881f
C446 B.n358 VSUBS 0.006881f
C447 B.n359 VSUBS 0.006881f
C448 B.n360 VSUBS 0.006881f
C449 B.n361 VSUBS 0.006881f
C450 B.n362 VSUBS 0.006881f
C451 B.n363 VSUBS 0.006881f
C452 B.n364 VSUBS 0.006881f
C453 B.n365 VSUBS 0.006881f
C454 B.n366 VSUBS 0.006881f
C455 B.n367 VSUBS 0.006881f
C456 B.n368 VSUBS 0.006881f
C457 B.n369 VSUBS 0.006881f
C458 B.n370 VSUBS 0.006881f
C459 B.n371 VSUBS 0.006881f
C460 B.n372 VSUBS 0.006881f
C461 B.n373 VSUBS 0.006881f
C462 B.n374 VSUBS 0.006881f
C463 B.n375 VSUBS 0.006881f
C464 B.n376 VSUBS 0.006881f
C465 B.n377 VSUBS 0.006881f
C466 B.n378 VSUBS 0.006881f
C467 B.n379 VSUBS 0.006881f
C468 B.n380 VSUBS 0.006881f
C469 B.n381 VSUBS 0.006881f
C470 B.n382 VSUBS 0.006881f
C471 B.n383 VSUBS 0.006881f
C472 B.n384 VSUBS 0.006881f
C473 B.n385 VSUBS 0.006881f
C474 B.n386 VSUBS 0.006881f
C475 B.n387 VSUBS 0.006881f
C476 B.n388 VSUBS 0.006881f
C477 B.n389 VSUBS 0.006881f
C478 B.n390 VSUBS 0.006881f
C479 B.n391 VSUBS 0.006881f
C480 B.n392 VSUBS 0.006881f
C481 B.n393 VSUBS 0.006881f
C482 B.n394 VSUBS 0.006881f
C483 B.n395 VSUBS 0.006881f
C484 B.n396 VSUBS 0.006881f
C485 B.n397 VSUBS 0.006881f
C486 B.n398 VSUBS 0.006881f
C487 B.n399 VSUBS 0.006881f
C488 B.n400 VSUBS 0.006881f
C489 B.n401 VSUBS 0.006881f
C490 B.n402 VSUBS 0.006881f
C491 B.n403 VSUBS 0.006881f
C492 B.n404 VSUBS 0.006881f
C493 B.n405 VSUBS 0.006881f
C494 B.n406 VSUBS 0.006881f
C495 B.n407 VSUBS 0.006881f
C496 B.n408 VSUBS 0.006881f
C497 B.n409 VSUBS 0.006881f
C498 B.n410 VSUBS 0.006881f
C499 B.n411 VSUBS 0.006881f
C500 B.n412 VSUBS 0.006881f
C501 B.n413 VSUBS 0.006881f
C502 B.n414 VSUBS 0.006881f
C503 B.n415 VSUBS 0.006881f
C504 B.n416 VSUBS 0.006881f
C505 B.n417 VSUBS 0.006881f
C506 B.n418 VSUBS 0.006881f
C507 B.n419 VSUBS 0.006881f
C508 B.n420 VSUBS 0.006881f
C509 B.n421 VSUBS 0.006881f
C510 B.n422 VSUBS 0.006881f
C511 B.n423 VSUBS 0.006881f
C512 B.n424 VSUBS 0.006881f
C513 B.n425 VSUBS 0.006881f
C514 B.n426 VSUBS 0.006881f
C515 B.n427 VSUBS 0.006881f
C516 B.n428 VSUBS 0.006881f
C517 B.n429 VSUBS 0.006881f
C518 B.n430 VSUBS 0.006881f
C519 B.n431 VSUBS 0.006881f
C520 B.n432 VSUBS 0.006881f
C521 B.n433 VSUBS 0.006881f
C522 B.n434 VSUBS 0.006881f
C523 B.n435 VSUBS 0.006881f
C524 B.n436 VSUBS 0.006881f
C525 B.n437 VSUBS 0.006881f
C526 B.n438 VSUBS 0.006881f
C527 B.n439 VSUBS 0.006881f
C528 B.n440 VSUBS 0.006881f
C529 B.n441 VSUBS 0.006881f
C530 B.n442 VSUBS 0.006881f
C531 B.n443 VSUBS 0.006881f
C532 B.n444 VSUBS 0.006881f
C533 B.n445 VSUBS 0.006881f
C534 B.n446 VSUBS 0.006881f
C535 B.n447 VSUBS 0.006881f
C536 B.n448 VSUBS 0.006881f
C537 B.n449 VSUBS 0.006881f
C538 B.n450 VSUBS 0.006881f
C539 B.n451 VSUBS 0.006881f
C540 B.n452 VSUBS 0.006881f
C541 B.n453 VSUBS 0.006881f
C542 B.n454 VSUBS 0.006881f
C543 B.n455 VSUBS 0.006881f
C544 B.n456 VSUBS 0.006881f
C545 B.n457 VSUBS 0.006881f
C546 B.n458 VSUBS 0.006881f
C547 B.n459 VSUBS 0.006881f
C548 B.n460 VSUBS 0.006881f
C549 B.n461 VSUBS 0.006881f
C550 B.n462 VSUBS 0.006881f
C551 B.n463 VSUBS 0.006881f
C552 B.n464 VSUBS 0.006881f
C553 B.n465 VSUBS 0.006881f
C554 B.n466 VSUBS 0.006881f
C555 B.n467 VSUBS 0.006881f
C556 B.n468 VSUBS 0.017356f
C557 B.n469 VSUBS 0.017356f
C558 B.n470 VSUBS 0.018062f
C559 B.n471 VSUBS 0.006881f
C560 B.n472 VSUBS 0.006881f
C561 B.n473 VSUBS 0.006881f
C562 B.n474 VSUBS 0.006881f
C563 B.n475 VSUBS 0.006881f
C564 B.n476 VSUBS 0.006881f
C565 B.n477 VSUBS 0.006881f
C566 B.n478 VSUBS 0.006881f
C567 B.n479 VSUBS 0.006881f
C568 B.n480 VSUBS 0.006881f
C569 B.n481 VSUBS 0.006881f
C570 B.n482 VSUBS 0.006881f
C571 B.n483 VSUBS 0.006881f
C572 B.n484 VSUBS 0.006881f
C573 B.n485 VSUBS 0.006881f
C574 B.n486 VSUBS 0.006881f
C575 B.n487 VSUBS 0.006881f
C576 B.n488 VSUBS 0.006881f
C577 B.n489 VSUBS 0.006881f
C578 B.n490 VSUBS 0.006881f
C579 B.n491 VSUBS 0.006881f
C580 B.n492 VSUBS 0.006881f
C581 B.n493 VSUBS 0.006881f
C582 B.n494 VSUBS 0.006881f
C583 B.n495 VSUBS 0.006881f
C584 B.n496 VSUBS 0.006881f
C585 B.n497 VSUBS 0.006881f
C586 B.n498 VSUBS 0.006881f
C587 B.n499 VSUBS 0.006881f
C588 B.n500 VSUBS 0.006881f
C589 B.n501 VSUBS 0.006881f
C590 B.n502 VSUBS 0.006881f
C591 B.n503 VSUBS 0.006881f
C592 B.n504 VSUBS 0.006881f
C593 B.n505 VSUBS 0.006881f
C594 B.n506 VSUBS 0.006881f
C595 B.n507 VSUBS 0.006881f
C596 B.n508 VSUBS 0.006881f
C597 B.n509 VSUBS 0.006881f
C598 B.n510 VSUBS 0.006881f
C599 B.n511 VSUBS 0.006881f
C600 B.n512 VSUBS 0.006881f
C601 B.n513 VSUBS 0.006881f
C602 B.n514 VSUBS 0.006476f
C603 B.n515 VSUBS 0.015943f
C604 B.n516 VSUBS 0.003845f
C605 B.n517 VSUBS 0.006881f
C606 B.n518 VSUBS 0.006881f
C607 B.n519 VSUBS 0.006881f
C608 B.n520 VSUBS 0.006881f
C609 B.n521 VSUBS 0.006881f
C610 B.n522 VSUBS 0.006881f
C611 B.n523 VSUBS 0.006881f
C612 B.n524 VSUBS 0.006881f
C613 B.n525 VSUBS 0.006881f
C614 B.n526 VSUBS 0.006881f
C615 B.n527 VSUBS 0.006881f
C616 B.n528 VSUBS 0.006881f
C617 B.n529 VSUBS 0.003845f
C618 B.n530 VSUBS 0.006881f
C619 B.n531 VSUBS 0.006881f
C620 B.n532 VSUBS 0.006881f
C621 B.n533 VSUBS 0.006881f
C622 B.n534 VSUBS 0.006881f
C623 B.n535 VSUBS 0.006881f
C624 B.n536 VSUBS 0.006881f
C625 B.n537 VSUBS 0.006881f
C626 B.n538 VSUBS 0.006881f
C627 B.n539 VSUBS 0.006881f
C628 B.n540 VSUBS 0.006881f
C629 B.n541 VSUBS 0.006881f
C630 B.n542 VSUBS 0.006881f
C631 B.n543 VSUBS 0.006881f
C632 B.n544 VSUBS 0.006881f
C633 B.n545 VSUBS 0.006881f
C634 B.n546 VSUBS 0.006881f
C635 B.n547 VSUBS 0.006881f
C636 B.n548 VSUBS 0.006881f
C637 B.n549 VSUBS 0.006881f
C638 B.n550 VSUBS 0.006881f
C639 B.n551 VSUBS 0.006881f
C640 B.n552 VSUBS 0.006881f
C641 B.n553 VSUBS 0.006881f
C642 B.n554 VSUBS 0.006881f
C643 B.n555 VSUBS 0.006881f
C644 B.n556 VSUBS 0.006881f
C645 B.n557 VSUBS 0.006881f
C646 B.n558 VSUBS 0.006881f
C647 B.n559 VSUBS 0.006881f
C648 B.n560 VSUBS 0.006881f
C649 B.n561 VSUBS 0.006881f
C650 B.n562 VSUBS 0.006881f
C651 B.n563 VSUBS 0.006881f
C652 B.n564 VSUBS 0.006881f
C653 B.n565 VSUBS 0.006881f
C654 B.n566 VSUBS 0.006881f
C655 B.n567 VSUBS 0.006881f
C656 B.n568 VSUBS 0.006881f
C657 B.n569 VSUBS 0.006881f
C658 B.n570 VSUBS 0.006881f
C659 B.n571 VSUBS 0.006881f
C660 B.n572 VSUBS 0.006881f
C661 B.n573 VSUBS 0.006881f
C662 B.n574 VSUBS 0.018062f
C663 B.n575 VSUBS 0.018062f
C664 B.n576 VSUBS 0.017356f
C665 B.n577 VSUBS 0.006881f
C666 B.n578 VSUBS 0.006881f
C667 B.n579 VSUBS 0.006881f
C668 B.n580 VSUBS 0.006881f
C669 B.n581 VSUBS 0.006881f
C670 B.n582 VSUBS 0.006881f
C671 B.n583 VSUBS 0.006881f
C672 B.n584 VSUBS 0.006881f
C673 B.n585 VSUBS 0.006881f
C674 B.n586 VSUBS 0.006881f
C675 B.n587 VSUBS 0.006881f
C676 B.n588 VSUBS 0.006881f
C677 B.n589 VSUBS 0.006881f
C678 B.n590 VSUBS 0.006881f
C679 B.n591 VSUBS 0.006881f
C680 B.n592 VSUBS 0.006881f
C681 B.n593 VSUBS 0.006881f
C682 B.n594 VSUBS 0.006881f
C683 B.n595 VSUBS 0.006881f
C684 B.n596 VSUBS 0.006881f
C685 B.n597 VSUBS 0.006881f
C686 B.n598 VSUBS 0.006881f
C687 B.n599 VSUBS 0.006881f
C688 B.n600 VSUBS 0.006881f
C689 B.n601 VSUBS 0.006881f
C690 B.n602 VSUBS 0.006881f
C691 B.n603 VSUBS 0.006881f
C692 B.n604 VSUBS 0.006881f
C693 B.n605 VSUBS 0.006881f
C694 B.n606 VSUBS 0.006881f
C695 B.n607 VSUBS 0.006881f
C696 B.n608 VSUBS 0.006881f
C697 B.n609 VSUBS 0.006881f
C698 B.n610 VSUBS 0.006881f
C699 B.n611 VSUBS 0.006881f
C700 B.n612 VSUBS 0.006881f
C701 B.n613 VSUBS 0.006881f
C702 B.n614 VSUBS 0.006881f
C703 B.n615 VSUBS 0.006881f
C704 B.n616 VSUBS 0.006881f
C705 B.n617 VSUBS 0.006881f
C706 B.n618 VSUBS 0.006881f
C707 B.n619 VSUBS 0.006881f
C708 B.n620 VSUBS 0.006881f
C709 B.n621 VSUBS 0.006881f
C710 B.n622 VSUBS 0.006881f
C711 B.n623 VSUBS 0.006881f
C712 B.n624 VSUBS 0.006881f
C713 B.n625 VSUBS 0.006881f
C714 B.n626 VSUBS 0.006881f
C715 B.n627 VSUBS 0.006881f
C716 B.n628 VSUBS 0.006881f
C717 B.n629 VSUBS 0.006881f
C718 B.n630 VSUBS 0.006881f
C719 B.n631 VSUBS 0.006881f
C720 B.n632 VSUBS 0.006881f
C721 B.n633 VSUBS 0.006881f
C722 B.n634 VSUBS 0.006881f
C723 B.n635 VSUBS 0.006881f
C724 B.n636 VSUBS 0.006881f
C725 B.n637 VSUBS 0.006881f
C726 B.n638 VSUBS 0.006881f
C727 B.n639 VSUBS 0.00898f
C728 B.n640 VSUBS 0.009566f
C729 B.n641 VSUBS 0.019022f
C730 VTAIL.t0 VSUBS 0.2012f
C731 VTAIL.t5 VSUBS 0.2012f
C732 VTAIL.n0 VSUBS 1.32688f
C733 VTAIL.n1 VSUBS 0.873195f
C734 VTAIL.t7 VSUBS 1.77989f
C735 VTAIL.n2 VSUBS 1.15909f
C736 VTAIL.t8 VSUBS 0.2012f
C737 VTAIL.t9 VSUBS 0.2012f
C738 VTAIL.n3 VSUBS 1.32688f
C739 VTAIL.n4 VSUBS 2.5374f
C740 VTAIL.t4 VSUBS 0.2012f
C741 VTAIL.t3 VSUBS 0.2012f
C742 VTAIL.n5 VSUBS 1.32689f
C743 VTAIL.n6 VSUBS 2.53739f
C744 VTAIL.t2 VSUBS 1.7799f
C745 VTAIL.n7 VSUBS 1.15908f
C746 VTAIL.t6 VSUBS 0.2012f
C747 VTAIL.t11 VSUBS 0.2012f
C748 VTAIL.n8 VSUBS 1.32689f
C749 VTAIL.n9 VSUBS 1.06337f
C750 VTAIL.t10 VSUBS 1.77989f
C751 VTAIL.n10 VSUBS 2.37178f
C752 VTAIL.t1 VSUBS 1.77989f
C753 VTAIL.n11 VSUBS 2.30062f
C754 VDD1.t0 VSUBS 1.62234f
C755 VDD1.t5 VSUBS 1.62126f
C756 VDD1.t1 VSUBS 0.167774f
C757 VDD1.t3 VSUBS 0.167774f
C758 VDD1.n0 VSUBS 1.22364f
C759 VDD1.n1 VSUBS 3.40292f
C760 VDD1.t4 VSUBS 0.167774f
C761 VDD1.t2 VSUBS 0.167774f
C762 VDD1.n2 VSUBS 1.21841f
C763 VDD1.n3 VSUBS 2.84618f
C764 VP.n0 VSUBS 0.04575f
C765 VP.t4 VSUBS 2.06569f
C766 VP.n1 VSUBS 0.068044f
C767 VP.n2 VSUBS 0.034703f
C768 VP.t2 VSUBS 2.06569f
C769 VP.n3 VSUBS 0.782092f
C770 VP.n4 VSUBS 0.034703f
C771 VP.n5 VSUBS 0.068044f
C772 VP.n6 VSUBS 0.04575f
C773 VP.t3 VSUBS 2.06569f
C774 VP.n7 VSUBS 0.04575f
C775 VP.t1 VSUBS 2.06569f
C776 VP.n8 VSUBS 0.068044f
C777 VP.n9 VSUBS 0.034703f
C778 VP.t0 VSUBS 2.06569f
C779 VP.n10 VSUBS 0.871275f
C780 VP.t5 VSUBS 2.36715f
C781 VP.n11 VSUBS 0.822919f
C782 VP.n12 VSUBS 0.360304f
C783 VP.n13 VSUBS 0.064354f
C784 VP.n14 VSUBS 0.069074f
C785 VP.n15 VSUBS 0.028128f
C786 VP.n16 VSUBS 0.034703f
C787 VP.n17 VSUBS 0.034703f
C788 VP.n18 VSUBS 0.034703f
C789 VP.n19 VSUBS 0.064354f
C790 VP.n20 VSUBS 0.03449f
C791 VP.n21 VSUBS 0.854116f
C792 VP.n22 VSUBS 1.71629f
C793 VP.n23 VSUBS 1.74342f
C794 VP.n24 VSUBS 0.854116f
C795 VP.n25 VSUBS 0.03449f
C796 VP.n26 VSUBS 0.064354f
C797 VP.n27 VSUBS 0.034703f
C798 VP.n28 VSUBS 0.034703f
C799 VP.n29 VSUBS 0.034703f
C800 VP.n30 VSUBS 0.028128f
C801 VP.n31 VSUBS 0.069074f
C802 VP.n32 VSUBS 0.064354f
C803 VP.n33 VSUBS 0.034703f
C804 VP.n34 VSUBS 0.034703f
C805 VP.n35 VSUBS 0.034703f
C806 VP.n36 VSUBS 0.064354f
C807 VP.n37 VSUBS 0.069074f
C808 VP.n38 VSUBS 0.028128f
C809 VP.n39 VSUBS 0.034703f
C810 VP.n40 VSUBS 0.034703f
C811 VP.n41 VSUBS 0.034703f
C812 VP.n42 VSUBS 0.064354f
C813 VP.n43 VSUBS 0.03449f
C814 VP.n44 VSUBS 0.854116f
C815 VP.n45 VSUBS 0.064237f
.ends

