* NGSPICE file created from diff_pair_sample_1715.ext - technology: sky130A

.subckt diff_pair_sample_1715 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=1.1253 ps=7.15 w=6.82 l=3.86
X1 VTAIL.t5 VN.t0 VDD2.t5 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=1.1253 pd=7.15 as=1.1253 ps=7.15 w=6.82 l=3.86
X2 VTAIL.t8 VP.t1 VDD1.t4 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=1.1253 pd=7.15 as=1.1253 ps=7.15 w=6.82 l=3.86
X3 VDD2.t4 VN.t1 VTAIL.t0 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=1.1253 pd=7.15 as=2.6598 ps=14.42 w=6.82 l=3.86
X4 VDD1.t3 VP.t2 VTAIL.t7 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=1.1253 pd=7.15 as=2.6598 ps=14.42 w=6.82 l=3.86
X5 VDD2.t3 VN.t2 VTAIL.t1 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=1.1253 ps=7.15 w=6.82 l=3.86
X6 B.t11 B.t9 B.t10 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=0 ps=0 w=6.82 l=3.86
X7 VDD2.t2 VN.t3 VTAIL.t4 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=1.1253 ps=7.15 w=6.82 l=3.86
X8 VDD2.t1 VN.t4 VTAIL.t3 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=1.1253 pd=7.15 as=2.6598 ps=14.42 w=6.82 l=3.86
X9 VTAIL.t10 VP.t3 VDD1.t2 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=1.1253 pd=7.15 as=1.1253 ps=7.15 w=6.82 l=3.86
X10 B.t8 B.t6 B.t7 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=0 ps=0 w=6.82 l=3.86
X11 VDD1.t1 VP.t4 VTAIL.t6 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=1.1253 pd=7.15 as=2.6598 ps=14.42 w=6.82 l=3.86
X12 VTAIL.t2 VN.t5 VDD2.t0 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=1.1253 pd=7.15 as=1.1253 ps=7.15 w=6.82 l=3.86
X13 B.t5 B.t3 B.t4 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=0 ps=0 w=6.82 l=3.86
X14 VDD1.t0 VP.t5 VTAIL.t11 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=1.1253 ps=7.15 w=6.82 l=3.86
X15 B.t2 B.t0 B.t1 w_n4322_n2332# sky130_fd_pr__pfet_01v8 ad=2.6598 pd=14.42 as=0 ps=0 w=6.82 l=3.86
R0 VP.n15 VP.n14 161.3
R1 VP.n16 VP.n11 161.3
R2 VP.n18 VP.n17 161.3
R3 VP.n19 VP.n10 161.3
R4 VP.n21 VP.n20 161.3
R5 VP.n22 VP.n9 161.3
R6 VP.n24 VP.n23 161.3
R7 VP.n25 VP.n8 161.3
R8 VP.n54 VP.n0 161.3
R9 VP.n53 VP.n52 161.3
R10 VP.n51 VP.n1 161.3
R11 VP.n50 VP.n49 161.3
R12 VP.n48 VP.n2 161.3
R13 VP.n47 VP.n46 161.3
R14 VP.n45 VP.n3 161.3
R15 VP.n44 VP.n43 161.3
R16 VP.n41 VP.n4 161.3
R17 VP.n40 VP.n39 161.3
R18 VP.n38 VP.n5 161.3
R19 VP.n37 VP.n36 161.3
R20 VP.n35 VP.n6 161.3
R21 VP.n34 VP.n33 161.3
R22 VP.n32 VP.n7 161.3
R23 VP.n31 VP.n30 161.3
R24 VP.n12 VP.t0 74.7092
R25 VP.n13 VP.n12 62.6969
R26 VP.n29 VP.n28 60.5633
R27 VP.n56 VP.n55 60.5633
R28 VP.n27 VP.n26 60.5633
R29 VP.n36 VP.n35 55.5035
R30 VP.n49 VP.n48 55.5035
R31 VP.n20 VP.n19 55.5035
R32 VP.n28 VP.n27 49.924
R33 VP.n29 VP.t5 42.5813
R34 VP.n42 VP.t3 42.5813
R35 VP.n55 VP.t4 42.5813
R36 VP.n26 VP.t2 42.5813
R37 VP.n13 VP.t1 42.5813
R38 VP.n35 VP.n34 25.3177
R39 VP.n49 VP.n1 25.3177
R40 VP.n20 VP.n9 25.3177
R41 VP.n30 VP.n7 24.3439
R42 VP.n34 VP.n7 24.3439
R43 VP.n36 VP.n5 24.3439
R44 VP.n40 VP.n5 24.3439
R45 VP.n41 VP.n40 24.3439
R46 VP.n43 VP.n3 24.3439
R47 VP.n47 VP.n3 24.3439
R48 VP.n48 VP.n47 24.3439
R49 VP.n53 VP.n1 24.3439
R50 VP.n54 VP.n53 24.3439
R51 VP.n24 VP.n9 24.3439
R52 VP.n25 VP.n24 24.3439
R53 VP.n14 VP.n11 24.3439
R54 VP.n18 VP.n11 24.3439
R55 VP.n19 VP.n18 24.3439
R56 VP.n30 VP.n29 21.4227
R57 VP.n55 VP.n54 21.4227
R58 VP.n26 VP.n25 21.4227
R59 VP.n42 VP.n41 12.1722
R60 VP.n43 VP.n42 12.1722
R61 VP.n14 VP.n13 12.1722
R62 VP.n15 VP.n12 2.65071
R63 VP.n27 VP.n8 0.417764
R64 VP.n31 VP.n28 0.417764
R65 VP.n56 VP.n0 0.417764
R66 VP VP.n56 0.394061
R67 VP.n16 VP.n15 0.189894
R68 VP.n17 VP.n16 0.189894
R69 VP.n17 VP.n10 0.189894
R70 VP.n21 VP.n10 0.189894
R71 VP.n22 VP.n21 0.189894
R72 VP.n23 VP.n22 0.189894
R73 VP.n23 VP.n8 0.189894
R74 VP.n32 VP.n31 0.189894
R75 VP.n33 VP.n32 0.189894
R76 VP.n33 VP.n6 0.189894
R77 VP.n37 VP.n6 0.189894
R78 VP.n38 VP.n37 0.189894
R79 VP.n39 VP.n38 0.189894
R80 VP.n39 VP.n4 0.189894
R81 VP.n44 VP.n4 0.189894
R82 VP.n45 VP.n44 0.189894
R83 VP.n46 VP.n45 0.189894
R84 VP.n46 VP.n2 0.189894
R85 VP.n50 VP.n2 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n52 VP.n51 0.189894
R88 VP.n52 VP.n0 0.189894
R89 VTAIL.n7 VTAIL.t3 76.306
R90 VTAIL.n11 VTAIL.t0 76.3059
R91 VTAIL.n2 VTAIL.t6 76.3059
R92 VTAIL.n10 VTAIL.t7 76.3059
R93 VTAIL.n9 VTAIL.n8 71.5399
R94 VTAIL.n6 VTAIL.n5 71.5399
R95 VTAIL.n1 VTAIL.n0 71.5388
R96 VTAIL.n4 VTAIL.n3 71.5388
R97 VTAIL.n6 VTAIL.n4 25.4703
R98 VTAIL.n11 VTAIL.n10 21.8583
R99 VTAIL.n0 VTAIL.t4 4.76663
R100 VTAIL.n0 VTAIL.t5 4.76663
R101 VTAIL.n3 VTAIL.t11 4.76663
R102 VTAIL.n3 VTAIL.t10 4.76663
R103 VTAIL.n8 VTAIL.t9 4.76663
R104 VTAIL.n8 VTAIL.t8 4.76663
R105 VTAIL.n5 VTAIL.t1 4.76663
R106 VTAIL.n5 VTAIL.t2 4.76663
R107 VTAIL.n7 VTAIL.n6 3.61257
R108 VTAIL.n10 VTAIL.n9 3.61257
R109 VTAIL.n4 VTAIL.n2 3.61257
R110 VTAIL VTAIL.n11 2.65136
R111 VTAIL.n9 VTAIL.n7 2.27636
R112 VTAIL.n2 VTAIL.n1 2.27636
R113 VTAIL VTAIL.n1 0.961707
R114 VDD1 VDD1.t5 95.752
R115 VDD1.n1 VDD1.t0 95.6384
R116 VDD1.n1 VDD1.n0 89.0652
R117 VDD1.n3 VDD1.n2 88.2185
R118 VDD1.n3 VDD1.n1 43.7229
R119 VDD1.n2 VDD1.t4 4.76663
R120 VDD1.n2 VDD1.t3 4.76663
R121 VDD1.n0 VDD1.t2 4.76663
R122 VDD1.n0 VDD1.t1 4.76663
R123 VDD1 VDD1.n3 0.845328
R124 VN.n37 VN.n20 161.3
R125 VN.n36 VN.n35 161.3
R126 VN.n34 VN.n21 161.3
R127 VN.n33 VN.n32 161.3
R128 VN.n31 VN.n22 161.3
R129 VN.n30 VN.n29 161.3
R130 VN.n28 VN.n23 161.3
R131 VN.n27 VN.n26 161.3
R132 VN.n17 VN.n0 161.3
R133 VN.n16 VN.n15 161.3
R134 VN.n14 VN.n1 161.3
R135 VN.n13 VN.n12 161.3
R136 VN.n11 VN.n2 161.3
R137 VN.n10 VN.n9 161.3
R138 VN.n8 VN.n3 161.3
R139 VN.n7 VN.n6 161.3
R140 VN.n4 VN.t3 74.7096
R141 VN.n24 VN.t4 74.7096
R142 VN.n5 VN.n4 62.6969
R143 VN.n25 VN.n24 62.6969
R144 VN.n19 VN.n18 60.5633
R145 VN.n39 VN.n38 60.5633
R146 VN.n12 VN.n11 55.5035
R147 VN.n32 VN.n31 55.5035
R148 VN VN.n39 49.9622
R149 VN.n5 VN.t0 42.5813
R150 VN.n18 VN.t1 42.5813
R151 VN.n25 VN.t5 42.5813
R152 VN.n38 VN.t2 42.5813
R153 VN.n12 VN.n1 25.3177
R154 VN.n32 VN.n21 25.3177
R155 VN.n6 VN.n3 24.3439
R156 VN.n10 VN.n3 24.3439
R157 VN.n11 VN.n10 24.3439
R158 VN.n16 VN.n1 24.3439
R159 VN.n17 VN.n16 24.3439
R160 VN.n31 VN.n30 24.3439
R161 VN.n30 VN.n23 24.3439
R162 VN.n26 VN.n23 24.3439
R163 VN.n37 VN.n36 24.3439
R164 VN.n36 VN.n21 24.3439
R165 VN.n18 VN.n17 21.4227
R166 VN.n38 VN.n37 21.4227
R167 VN.n6 VN.n5 12.1722
R168 VN.n26 VN.n25 12.1722
R169 VN.n27 VN.n24 2.65074
R170 VN.n7 VN.n4 2.65074
R171 VN.n39 VN.n20 0.417764
R172 VN.n19 VN.n0 0.417764
R173 VN VN.n19 0.394061
R174 VN.n35 VN.n20 0.189894
R175 VN.n35 VN.n34 0.189894
R176 VN.n34 VN.n33 0.189894
R177 VN.n33 VN.n22 0.189894
R178 VN.n29 VN.n22 0.189894
R179 VN.n29 VN.n28 0.189894
R180 VN.n28 VN.n27 0.189894
R181 VN.n8 VN.n7 0.189894
R182 VN.n9 VN.n8 0.189894
R183 VN.n9 VN.n2 0.189894
R184 VN.n13 VN.n2 0.189894
R185 VN.n14 VN.n13 0.189894
R186 VN.n15 VN.n14 0.189894
R187 VN.n15 VN.n0 0.189894
R188 VDD2.n1 VDD2.t2 95.6384
R189 VDD2.n2 VDD2.t3 92.9848
R190 VDD2.n1 VDD2.n0 89.0652
R191 VDD2 VDD2.n3 89.0634
R192 VDD2.n2 VDD2.n1 41.3338
R193 VDD2.n3 VDD2.t0 4.76663
R194 VDD2.n3 VDD2.t1 4.76663
R195 VDD2.n0 VDD2.t5 4.76663
R196 VDD2.n0 VDD2.t4 4.76663
R197 VDD2 VDD2.n2 2.76774
R198 B.n366 B.n365 585
R199 B.n364 B.n125 585
R200 B.n363 B.n362 585
R201 B.n361 B.n126 585
R202 B.n360 B.n359 585
R203 B.n358 B.n127 585
R204 B.n357 B.n356 585
R205 B.n355 B.n128 585
R206 B.n354 B.n353 585
R207 B.n352 B.n129 585
R208 B.n351 B.n350 585
R209 B.n349 B.n130 585
R210 B.n348 B.n347 585
R211 B.n346 B.n131 585
R212 B.n345 B.n344 585
R213 B.n343 B.n132 585
R214 B.n342 B.n341 585
R215 B.n340 B.n133 585
R216 B.n339 B.n338 585
R217 B.n337 B.n134 585
R218 B.n336 B.n335 585
R219 B.n334 B.n135 585
R220 B.n333 B.n332 585
R221 B.n331 B.n136 585
R222 B.n330 B.n329 585
R223 B.n328 B.n137 585
R224 B.n327 B.n326 585
R225 B.n322 B.n138 585
R226 B.n321 B.n320 585
R227 B.n319 B.n139 585
R228 B.n318 B.n317 585
R229 B.n316 B.n140 585
R230 B.n315 B.n314 585
R231 B.n313 B.n141 585
R232 B.n312 B.n311 585
R233 B.n310 B.n142 585
R234 B.n308 B.n307 585
R235 B.n306 B.n145 585
R236 B.n305 B.n304 585
R237 B.n303 B.n146 585
R238 B.n302 B.n301 585
R239 B.n300 B.n147 585
R240 B.n299 B.n298 585
R241 B.n297 B.n148 585
R242 B.n296 B.n295 585
R243 B.n294 B.n149 585
R244 B.n293 B.n292 585
R245 B.n291 B.n150 585
R246 B.n290 B.n289 585
R247 B.n288 B.n151 585
R248 B.n287 B.n286 585
R249 B.n285 B.n152 585
R250 B.n284 B.n283 585
R251 B.n282 B.n153 585
R252 B.n281 B.n280 585
R253 B.n279 B.n154 585
R254 B.n278 B.n277 585
R255 B.n276 B.n155 585
R256 B.n275 B.n274 585
R257 B.n273 B.n156 585
R258 B.n272 B.n271 585
R259 B.n270 B.n157 585
R260 B.n367 B.n124 585
R261 B.n369 B.n368 585
R262 B.n370 B.n123 585
R263 B.n372 B.n371 585
R264 B.n373 B.n122 585
R265 B.n375 B.n374 585
R266 B.n376 B.n121 585
R267 B.n378 B.n377 585
R268 B.n379 B.n120 585
R269 B.n381 B.n380 585
R270 B.n382 B.n119 585
R271 B.n384 B.n383 585
R272 B.n385 B.n118 585
R273 B.n387 B.n386 585
R274 B.n388 B.n117 585
R275 B.n390 B.n389 585
R276 B.n391 B.n116 585
R277 B.n393 B.n392 585
R278 B.n394 B.n115 585
R279 B.n396 B.n395 585
R280 B.n397 B.n114 585
R281 B.n399 B.n398 585
R282 B.n400 B.n113 585
R283 B.n402 B.n401 585
R284 B.n403 B.n112 585
R285 B.n405 B.n404 585
R286 B.n406 B.n111 585
R287 B.n408 B.n407 585
R288 B.n409 B.n110 585
R289 B.n411 B.n410 585
R290 B.n412 B.n109 585
R291 B.n414 B.n413 585
R292 B.n415 B.n108 585
R293 B.n417 B.n416 585
R294 B.n418 B.n107 585
R295 B.n420 B.n419 585
R296 B.n421 B.n106 585
R297 B.n423 B.n422 585
R298 B.n424 B.n105 585
R299 B.n426 B.n425 585
R300 B.n427 B.n104 585
R301 B.n429 B.n428 585
R302 B.n430 B.n103 585
R303 B.n432 B.n431 585
R304 B.n433 B.n102 585
R305 B.n435 B.n434 585
R306 B.n436 B.n101 585
R307 B.n438 B.n437 585
R308 B.n439 B.n100 585
R309 B.n441 B.n440 585
R310 B.n442 B.n99 585
R311 B.n444 B.n443 585
R312 B.n445 B.n98 585
R313 B.n447 B.n446 585
R314 B.n448 B.n97 585
R315 B.n450 B.n449 585
R316 B.n451 B.n96 585
R317 B.n453 B.n452 585
R318 B.n454 B.n95 585
R319 B.n456 B.n455 585
R320 B.n457 B.n94 585
R321 B.n459 B.n458 585
R322 B.n460 B.n93 585
R323 B.n462 B.n461 585
R324 B.n463 B.n92 585
R325 B.n465 B.n464 585
R326 B.n466 B.n91 585
R327 B.n468 B.n467 585
R328 B.n469 B.n90 585
R329 B.n471 B.n470 585
R330 B.n472 B.n89 585
R331 B.n474 B.n473 585
R332 B.n475 B.n88 585
R333 B.n477 B.n476 585
R334 B.n478 B.n87 585
R335 B.n480 B.n479 585
R336 B.n481 B.n86 585
R337 B.n483 B.n482 585
R338 B.n484 B.n85 585
R339 B.n486 B.n485 585
R340 B.n487 B.n84 585
R341 B.n489 B.n488 585
R342 B.n490 B.n83 585
R343 B.n492 B.n491 585
R344 B.n493 B.n82 585
R345 B.n495 B.n494 585
R346 B.n496 B.n81 585
R347 B.n498 B.n497 585
R348 B.n499 B.n80 585
R349 B.n501 B.n500 585
R350 B.n502 B.n79 585
R351 B.n504 B.n503 585
R352 B.n505 B.n78 585
R353 B.n507 B.n506 585
R354 B.n508 B.n77 585
R355 B.n510 B.n509 585
R356 B.n511 B.n76 585
R357 B.n513 B.n512 585
R358 B.n514 B.n75 585
R359 B.n516 B.n515 585
R360 B.n517 B.n74 585
R361 B.n519 B.n518 585
R362 B.n520 B.n73 585
R363 B.n522 B.n521 585
R364 B.n523 B.n72 585
R365 B.n525 B.n524 585
R366 B.n526 B.n71 585
R367 B.n528 B.n527 585
R368 B.n529 B.n70 585
R369 B.n531 B.n530 585
R370 B.n532 B.n69 585
R371 B.n534 B.n533 585
R372 B.n535 B.n68 585
R373 B.n537 B.n536 585
R374 B.n538 B.n67 585
R375 B.n540 B.n539 585
R376 B.n634 B.n633 585
R377 B.n632 B.n31 585
R378 B.n631 B.n630 585
R379 B.n629 B.n32 585
R380 B.n628 B.n627 585
R381 B.n626 B.n33 585
R382 B.n625 B.n624 585
R383 B.n623 B.n34 585
R384 B.n622 B.n621 585
R385 B.n620 B.n35 585
R386 B.n619 B.n618 585
R387 B.n617 B.n36 585
R388 B.n616 B.n615 585
R389 B.n614 B.n37 585
R390 B.n613 B.n612 585
R391 B.n611 B.n38 585
R392 B.n610 B.n609 585
R393 B.n608 B.n39 585
R394 B.n607 B.n606 585
R395 B.n605 B.n40 585
R396 B.n604 B.n603 585
R397 B.n602 B.n41 585
R398 B.n601 B.n600 585
R399 B.n599 B.n42 585
R400 B.n598 B.n597 585
R401 B.n596 B.n43 585
R402 B.n594 B.n593 585
R403 B.n592 B.n46 585
R404 B.n591 B.n590 585
R405 B.n589 B.n47 585
R406 B.n588 B.n587 585
R407 B.n586 B.n48 585
R408 B.n585 B.n584 585
R409 B.n583 B.n49 585
R410 B.n582 B.n581 585
R411 B.n580 B.n50 585
R412 B.n579 B.n578 585
R413 B.n577 B.n51 585
R414 B.n576 B.n575 585
R415 B.n574 B.n55 585
R416 B.n573 B.n572 585
R417 B.n571 B.n56 585
R418 B.n570 B.n569 585
R419 B.n568 B.n57 585
R420 B.n567 B.n566 585
R421 B.n565 B.n58 585
R422 B.n564 B.n563 585
R423 B.n562 B.n59 585
R424 B.n561 B.n560 585
R425 B.n559 B.n60 585
R426 B.n558 B.n557 585
R427 B.n556 B.n61 585
R428 B.n555 B.n554 585
R429 B.n553 B.n62 585
R430 B.n552 B.n551 585
R431 B.n550 B.n63 585
R432 B.n549 B.n548 585
R433 B.n547 B.n64 585
R434 B.n546 B.n545 585
R435 B.n544 B.n65 585
R436 B.n543 B.n542 585
R437 B.n541 B.n66 585
R438 B.n635 B.n30 585
R439 B.n637 B.n636 585
R440 B.n638 B.n29 585
R441 B.n640 B.n639 585
R442 B.n641 B.n28 585
R443 B.n643 B.n642 585
R444 B.n644 B.n27 585
R445 B.n646 B.n645 585
R446 B.n647 B.n26 585
R447 B.n649 B.n648 585
R448 B.n650 B.n25 585
R449 B.n652 B.n651 585
R450 B.n653 B.n24 585
R451 B.n655 B.n654 585
R452 B.n656 B.n23 585
R453 B.n658 B.n657 585
R454 B.n659 B.n22 585
R455 B.n661 B.n660 585
R456 B.n662 B.n21 585
R457 B.n664 B.n663 585
R458 B.n665 B.n20 585
R459 B.n667 B.n666 585
R460 B.n668 B.n19 585
R461 B.n670 B.n669 585
R462 B.n671 B.n18 585
R463 B.n673 B.n672 585
R464 B.n674 B.n17 585
R465 B.n676 B.n675 585
R466 B.n677 B.n16 585
R467 B.n679 B.n678 585
R468 B.n680 B.n15 585
R469 B.n682 B.n681 585
R470 B.n683 B.n14 585
R471 B.n685 B.n684 585
R472 B.n686 B.n13 585
R473 B.n688 B.n687 585
R474 B.n689 B.n12 585
R475 B.n691 B.n690 585
R476 B.n692 B.n11 585
R477 B.n694 B.n693 585
R478 B.n695 B.n10 585
R479 B.n697 B.n696 585
R480 B.n698 B.n9 585
R481 B.n700 B.n699 585
R482 B.n701 B.n8 585
R483 B.n703 B.n702 585
R484 B.n704 B.n7 585
R485 B.n706 B.n705 585
R486 B.n707 B.n6 585
R487 B.n709 B.n708 585
R488 B.n710 B.n5 585
R489 B.n712 B.n711 585
R490 B.n713 B.n4 585
R491 B.n715 B.n714 585
R492 B.n716 B.n3 585
R493 B.n718 B.n717 585
R494 B.n719 B.n0 585
R495 B.n2 B.n1 585
R496 B.n186 B.n185 585
R497 B.n188 B.n187 585
R498 B.n189 B.n184 585
R499 B.n191 B.n190 585
R500 B.n192 B.n183 585
R501 B.n194 B.n193 585
R502 B.n195 B.n182 585
R503 B.n197 B.n196 585
R504 B.n198 B.n181 585
R505 B.n200 B.n199 585
R506 B.n201 B.n180 585
R507 B.n203 B.n202 585
R508 B.n204 B.n179 585
R509 B.n206 B.n205 585
R510 B.n207 B.n178 585
R511 B.n209 B.n208 585
R512 B.n210 B.n177 585
R513 B.n212 B.n211 585
R514 B.n213 B.n176 585
R515 B.n215 B.n214 585
R516 B.n216 B.n175 585
R517 B.n218 B.n217 585
R518 B.n219 B.n174 585
R519 B.n221 B.n220 585
R520 B.n222 B.n173 585
R521 B.n224 B.n223 585
R522 B.n225 B.n172 585
R523 B.n227 B.n226 585
R524 B.n228 B.n171 585
R525 B.n230 B.n229 585
R526 B.n231 B.n170 585
R527 B.n233 B.n232 585
R528 B.n234 B.n169 585
R529 B.n236 B.n235 585
R530 B.n237 B.n168 585
R531 B.n239 B.n238 585
R532 B.n240 B.n167 585
R533 B.n242 B.n241 585
R534 B.n243 B.n166 585
R535 B.n245 B.n244 585
R536 B.n246 B.n165 585
R537 B.n248 B.n247 585
R538 B.n249 B.n164 585
R539 B.n251 B.n250 585
R540 B.n252 B.n163 585
R541 B.n254 B.n253 585
R542 B.n255 B.n162 585
R543 B.n257 B.n256 585
R544 B.n258 B.n161 585
R545 B.n260 B.n259 585
R546 B.n261 B.n160 585
R547 B.n263 B.n262 585
R548 B.n264 B.n159 585
R549 B.n266 B.n265 585
R550 B.n267 B.n158 585
R551 B.n269 B.n268 585
R552 B.n270 B.n269 511.721
R553 B.n365 B.n124 511.721
R554 B.n539 B.n66 511.721
R555 B.n635 B.n634 511.721
R556 B.n721 B.n720 256.663
R557 B.n143 B.t0 251.97
R558 B.n323 B.t9 251.97
R559 B.n52 B.t6 251.97
R560 B.n44 B.t3 251.97
R561 B.n720 B.n719 235.042
R562 B.n720 B.n2 235.042
R563 B.n323 B.t10 191.388
R564 B.n52 B.t8 191.388
R565 B.n143 B.t1 191.381
R566 B.n44 B.t5 191.381
R567 B.n271 B.n270 163.367
R568 B.n271 B.n156 163.367
R569 B.n275 B.n156 163.367
R570 B.n276 B.n275 163.367
R571 B.n277 B.n276 163.367
R572 B.n277 B.n154 163.367
R573 B.n281 B.n154 163.367
R574 B.n282 B.n281 163.367
R575 B.n283 B.n282 163.367
R576 B.n283 B.n152 163.367
R577 B.n287 B.n152 163.367
R578 B.n288 B.n287 163.367
R579 B.n289 B.n288 163.367
R580 B.n289 B.n150 163.367
R581 B.n293 B.n150 163.367
R582 B.n294 B.n293 163.367
R583 B.n295 B.n294 163.367
R584 B.n295 B.n148 163.367
R585 B.n299 B.n148 163.367
R586 B.n300 B.n299 163.367
R587 B.n301 B.n300 163.367
R588 B.n301 B.n146 163.367
R589 B.n305 B.n146 163.367
R590 B.n306 B.n305 163.367
R591 B.n307 B.n306 163.367
R592 B.n307 B.n142 163.367
R593 B.n312 B.n142 163.367
R594 B.n313 B.n312 163.367
R595 B.n314 B.n313 163.367
R596 B.n314 B.n140 163.367
R597 B.n318 B.n140 163.367
R598 B.n319 B.n318 163.367
R599 B.n320 B.n319 163.367
R600 B.n320 B.n138 163.367
R601 B.n327 B.n138 163.367
R602 B.n328 B.n327 163.367
R603 B.n329 B.n328 163.367
R604 B.n329 B.n136 163.367
R605 B.n333 B.n136 163.367
R606 B.n334 B.n333 163.367
R607 B.n335 B.n334 163.367
R608 B.n335 B.n134 163.367
R609 B.n339 B.n134 163.367
R610 B.n340 B.n339 163.367
R611 B.n341 B.n340 163.367
R612 B.n341 B.n132 163.367
R613 B.n345 B.n132 163.367
R614 B.n346 B.n345 163.367
R615 B.n347 B.n346 163.367
R616 B.n347 B.n130 163.367
R617 B.n351 B.n130 163.367
R618 B.n352 B.n351 163.367
R619 B.n353 B.n352 163.367
R620 B.n353 B.n128 163.367
R621 B.n357 B.n128 163.367
R622 B.n358 B.n357 163.367
R623 B.n359 B.n358 163.367
R624 B.n359 B.n126 163.367
R625 B.n363 B.n126 163.367
R626 B.n364 B.n363 163.367
R627 B.n365 B.n364 163.367
R628 B.n539 B.n538 163.367
R629 B.n538 B.n537 163.367
R630 B.n537 B.n68 163.367
R631 B.n533 B.n68 163.367
R632 B.n533 B.n532 163.367
R633 B.n532 B.n531 163.367
R634 B.n531 B.n70 163.367
R635 B.n527 B.n70 163.367
R636 B.n527 B.n526 163.367
R637 B.n526 B.n525 163.367
R638 B.n525 B.n72 163.367
R639 B.n521 B.n72 163.367
R640 B.n521 B.n520 163.367
R641 B.n520 B.n519 163.367
R642 B.n519 B.n74 163.367
R643 B.n515 B.n74 163.367
R644 B.n515 B.n514 163.367
R645 B.n514 B.n513 163.367
R646 B.n513 B.n76 163.367
R647 B.n509 B.n76 163.367
R648 B.n509 B.n508 163.367
R649 B.n508 B.n507 163.367
R650 B.n507 B.n78 163.367
R651 B.n503 B.n78 163.367
R652 B.n503 B.n502 163.367
R653 B.n502 B.n501 163.367
R654 B.n501 B.n80 163.367
R655 B.n497 B.n80 163.367
R656 B.n497 B.n496 163.367
R657 B.n496 B.n495 163.367
R658 B.n495 B.n82 163.367
R659 B.n491 B.n82 163.367
R660 B.n491 B.n490 163.367
R661 B.n490 B.n489 163.367
R662 B.n489 B.n84 163.367
R663 B.n485 B.n84 163.367
R664 B.n485 B.n484 163.367
R665 B.n484 B.n483 163.367
R666 B.n483 B.n86 163.367
R667 B.n479 B.n86 163.367
R668 B.n479 B.n478 163.367
R669 B.n478 B.n477 163.367
R670 B.n477 B.n88 163.367
R671 B.n473 B.n88 163.367
R672 B.n473 B.n472 163.367
R673 B.n472 B.n471 163.367
R674 B.n471 B.n90 163.367
R675 B.n467 B.n90 163.367
R676 B.n467 B.n466 163.367
R677 B.n466 B.n465 163.367
R678 B.n465 B.n92 163.367
R679 B.n461 B.n92 163.367
R680 B.n461 B.n460 163.367
R681 B.n460 B.n459 163.367
R682 B.n459 B.n94 163.367
R683 B.n455 B.n94 163.367
R684 B.n455 B.n454 163.367
R685 B.n454 B.n453 163.367
R686 B.n453 B.n96 163.367
R687 B.n449 B.n96 163.367
R688 B.n449 B.n448 163.367
R689 B.n448 B.n447 163.367
R690 B.n447 B.n98 163.367
R691 B.n443 B.n98 163.367
R692 B.n443 B.n442 163.367
R693 B.n442 B.n441 163.367
R694 B.n441 B.n100 163.367
R695 B.n437 B.n100 163.367
R696 B.n437 B.n436 163.367
R697 B.n436 B.n435 163.367
R698 B.n435 B.n102 163.367
R699 B.n431 B.n102 163.367
R700 B.n431 B.n430 163.367
R701 B.n430 B.n429 163.367
R702 B.n429 B.n104 163.367
R703 B.n425 B.n104 163.367
R704 B.n425 B.n424 163.367
R705 B.n424 B.n423 163.367
R706 B.n423 B.n106 163.367
R707 B.n419 B.n106 163.367
R708 B.n419 B.n418 163.367
R709 B.n418 B.n417 163.367
R710 B.n417 B.n108 163.367
R711 B.n413 B.n108 163.367
R712 B.n413 B.n412 163.367
R713 B.n412 B.n411 163.367
R714 B.n411 B.n110 163.367
R715 B.n407 B.n110 163.367
R716 B.n407 B.n406 163.367
R717 B.n406 B.n405 163.367
R718 B.n405 B.n112 163.367
R719 B.n401 B.n112 163.367
R720 B.n401 B.n400 163.367
R721 B.n400 B.n399 163.367
R722 B.n399 B.n114 163.367
R723 B.n395 B.n114 163.367
R724 B.n395 B.n394 163.367
R725 B.n394 B.n393 163.367
R726 B.n393 B.n116 163.367
R727 B.n389 B.n116 163.367
R728 B.n389 B.n388 163.367
R729 B.n388 B.n387 163.367
R730 B.n387 B.n118 163.367
R731 B.n383 B.n118 163.367
R732 B.n383 B.n382 163.367
R733 B.n382 B.n381 163.367
R734 B.n381 B.n120 163.367
R735 B.n377 B.n120 163.367
R736 B.n377 B.n376 163.367
R737 B.n376 B.n375 163.367
R738 B.n375 B.n122 163.367
R739 B.n371 B.n122 163.367
R740 B.n371 B.n370 163.367
R741 B.n370 B.n369 163.367
R742 B.n369 B.n124 163.367
R743 B.n634 B.n31 163.367
R744 B.n630 B.n31 163.367
R745 B.n630 B.n629 163.367
R746 B.n629 B.n628 163.367
R747 B.n628 B.n33 163.367
R748 B.n624 B.n33 163.367
R749 B.n624 B.n623 163.367
R750 B.n623 B.n622 163.367
R751 B.n622 B.n35 163.367
R752 B.n618 B.n35 163.367
R753 B.n618 B.n617 163.367
R754 B.n617 B.n616 163.367
R755 B.n616 B.n37 163.367
R756 B.n612 B.n37 163.367
R757 B.n612 B.n611 163.367
R758 B.n611 B.n610 163.367
R759 B.n610 B.n39 163.367
R760 B.n606 B.n39 163.367
R761 B.n606 B.n605 163.367
R762 B.n605 B.n604 163.367
R763 B.n604 B.n41 163.367
R764 B.n600 B.n41 163.367
R765 B.n600 B.n599 163.367
R766 B.n599 B.n598 163.367
R767 B.n598 B.n43 163.367
R768 B.n593 B.n43 163.367
R769 B.n593 B.n592 163.367
R770 B.n592 B.n591 163.367
R771 B.n591 B.n47 163.367
R772 B.n587 B.n47 163.367
R773 B.n587 B.n586 163.367
R774 B.n586 B.n585 163.367
R775 B.n585 B.n49 163.367
R776 B.n581 B.n49 163.367
R777 B.n581 B.n580 163.367
R778 B.n580 B.n579 163.367
R779 B.n579 B.n51 163.367
R780 B.n575 B.n51 163.367
R781 B.n575 B.n574 163.367
R782 B.n574 B.n573 163.367
R783 B.n573 B.n56 163.367
R784 B.n569 B.n56 163.367
R785 B.n569 B.n568 163.367
R786 B.n568 B.n567 163.367
R787 B.n567 B.n58 163.367
R788 B.n563 B.n58 163.367
R789 B.n563 B.n562 163.367
R790 B.n562 B.n561 163.367
R791 B.n561 B.n60 163.367
R792 B.n557 B.n60 163.367
R793 B.n557 B.n556 163.367
R794 B.n556 B.n555 163.367
R795 B.n555 B.n62 163.367
R796 B.n551 B.n62 163.367
R797 B.n551 B.n550 163.367
R798 B.n550 B.n549 163.367
R799 B.n549 B.n64 163.367
R800 B.n545 B.n64 163.367
R801 B.n545 B.n544 163.367
R802 B.n544 B.n543 163.367
R803 B.n543 B.n66 163.367
R804 B.n636 B.n635 163.367
R805 B.n636 B.n29 163.367
R806 B.n640 B.n29 163.367
R807 B.n641 B.n640 163.367
R808 B.n642 B.n641 163.367
R809 B.n642 B.n27 163.367
R810 B.n646 B.n27 163.367
R811 B.n647 B.n646 163.367
R812 B.n648 B.n647 163.367
R813 B.n648 B.n25 163.367
R814 B.n652 B.n25 163.367
R815 B.n653 B.n652 163.367
R816 B.n654 B.n653 163.367
R817 B.n654 B.n23 163.367
R818 B.n658 B.n23 163.367
R819 B.n659 B.n658 163.367
R820 B.n660 B.n659 163.367
R821 B.n660 B.n21 163.367
R822 B.n664 B.n21 163.367
R823 B.n665 B.n664 163.367
R824 B.n666 B.n665 163.367
R825 B.n666 B.n19 163.367
R826 B.n670 B.n19 163.367
R827 B.n671 B.n670 163.367
R828 B.n672 B.n671 163.367
R829 B.n672 B.n17 163.367
R830 B.n676 B.n17 163.367
R831 B.n677 B.n676 163.367
R832 B.n678 B.n677 163.367
R833 B.n678 B.n15 163.367
R834 B.n682 B.n15 163.367
R835 B.n683 B.n682 163.367
R836 B.n684 B.n683 163.367
R837 B.n684 B.n13 163.367
R838 B.n688 B.n13 163.367
R839 B.n689 B.n688 163.367
R840 B.n690 B.n689 163.367
R841 B.n690 B.n11 163.367
R842 B.n694 B.n11 163.367
R843 B.n695 B.n694 163.367
R844 B.n696 B.n695 163.367
R845 B.n696 B.n9 163.367
R846 B.n700 B.n9 163.367
R847 B.n701 B.n700 163.367
R848 B.n702 B.n701 163.367
R849 B.n702 B.n7 163.367
R850 B.n706 B.n7 163.367
R851 B.n707 B.n706 163.367
R852 B.n708 B.n707 163.367
R853 B.n708 B.n5 163.367
R854 B.n712 B.n5 163.367
R855 B.n713 B.n712 163.367
R856 B.n714 B.n713 163.367
R857 B.n714 B.n3 163.367
R858 B.n718 B.n3 163.367
R859 B.n719 B.n718 163.367
R860 B.n186 B.n2 163.367
R861 B.n187 B.n186 163.367
R862 B.n187 B.n184 163.367
R863 B.n191 B.n184 163.367
R864 B.n192 B.n191 163.367
R865 B.n193 B.n192 163.367
R866 B.n193 B.n182 163.367
R867 B.n197 B.n182 163.367
R868 B.n198 B.n197 163.367
R869 B.n199 B.n198 163.367
R870 B.n199 B.n180 163.367
R871 B.n203 B.n180 163.367
R872 B.n204 B.n203 163.367
R873 B.n205 B.n204 163.367
R874 B.n205 B.n178 163.367
R875 B.n209 B.n178 163.367
R876 B.n210 B.n209 163.367
R877 B.n211 B.n210 163.367
R878 B.n211 B.n176 163.367
R879 B.n215 B.n176 163.367
R880 B.n216 B.n215 163.367
R881 B.n217 B.n216 163.367
R882 B.n217 B.n174 163.367
R883 B.n221 B.n174 163.367
R884 B.n222 B.n221 163.367
R885 B.n223 B.n222 163.367
R886 B.n223 B.n172 163.367
R887 B.n227 B.n172 163.367
R888 B.n228 B.n227 163.367
R889 B.n229 B.n228 163.367
R890 B.n229 B.n170 163.367
R891 B.n233 B.n170 163.367
R892 B.n234 B.n233 163.367
R893 B.n235 B.n234 163.367
R894 B.n235 B.n168 163.367
R895 B.n239 B.n168 163.367
R896 B.n240 B.n239 163.367
R897 B.n241 B.n240 163.367
R898 B.n241 B.n166 163.367
R899 B.n245 B.n166 163.367
R900 B.n246 B.n245 163.367
R901 B.n247 B.n246 163.367
R902 B.n247 B.n164 163.367
R903 B.n251 B.n164 163.367
R904 B.n252 B.n251 163.367
R905 B.n253 B.n252 163.367
R906 B.n253 B.n162 163.367
R907 B.n257 B.n162 163.367
R908 B.n258 B.n257 163.367
R909 B.n259 B.n258 163.367
R910 B.n259 B.n160 163.367
R911 B.n263 B.n160 163.367
R912 B.n264 B.n263 163.367
R913 B.n265 B.n264 163.367
R914 B.n265 B.n158 163.367
R915 B.n269 B.n158 163.367
R916 B.n324 B.t11 110.127
R917 B.n53 B.t7 110.127
R918 B.n144 B.t2 110.121
R919 B.n45 B.t4 110.121
R920 B.n144 B.n143 81.2611
R921 B.n324 B.n323 81.2611
R922 B.n53 B.n52 81.2611
R923 B.n45 B.n44 81.2611
R924 B.n309 B.n144 59.5399
R925 B.n325 B.n324 59.5399
R926 B.n54 B.n53 59.5399
R927 B.n595 B.n45 59.5399
R928 B.n633 B.n30 33.2493
R929 B.n541 B.n540 33.2493
R930 B.n367 B.n366 33.2493
R931 B.n268 B.n157 33.2493
R932 B B.n721 18.0485
R933 B.n637 B.n30 10.6151
R934 B.n638 B.n637 10.6151
R935 B.n639 B.n638 10.6151
R936 B.n639 B.n28 10.6151
R937 B.n643 B.n28 10.6151
R938 B.n644 B.n643 10.6151
R939 B.n645 B.n644 10.6151
R940 B.n645 B.n26 10.6151
R941 B.n649 B.n26 10.6151
R942 B.n650 B.n649 10.6151
R943 B.n651 B.n650 10.6151
R944 B.n651 B.n24 10.6151
R945 B.n655 B.n24 10.6151
R946 B.n656 B.n655 10.6151
R947 B.n657 B.n656 10.6151
R948 B.n657 B.n22 10.6151
R949 B.n661 B.n22 10.6151
R950 B.n662 B.n661 10.6151
R951 B.n663 B.n662 10.6151
R952 B.n663 B.n20 10.6151
R953 B.n667 B.n20 10.6151
R954 B.n668 B.n667 10.6151
R955 B.n669 B.n668 10.6151
R956 B.n669 B.n18 10.6151
R957 B.n673 B.n18 10.6151
R958 B.n674 B.n673 10.6151
R959 B.n675 B.n674 10.6151
R960 B.n675 B.n16 10.6151
R961 B.n679 B.n16 10.6151
R962 B.n680 B.n679 10.6151
R963 B.n681 B.n680 10.6151
R964 B.n681 B.n14 10.6151
R965 B.n685 B.n14 10.6151
R966 B.n686 B.n685 10.6151
R967 B.n687 B.n686 10.6151
R968 B.n687 B.n12 10.6151
R969 B.n691 B.n12 10.6151
R970 B.n692 B.n691 10.6151
R971 B.n693 B.n692 10.6151
R972 B.n693 B.n10 10.6151
R973 B.n697 B.n10 10.6151
R974 B.n698 B.n697 10.6151
R975 B.n699 B.n698 10.6151
R976 B.n699 B.n8 10.6151
R977 B.n703 B.n8 10.6151
R978 B.n704 B.n703 10.6151
R979 B.n705 B.n704 10.6151
R980 B.n705 B.n6 10.6151
R981 B.n709 B.n6 10.6151
R982 B.n710 B.n709 10.6151
R983 B.n711 B.n710 10.6151
R984 B.n711 B.n4 10.6151
R985 B.n715 B.n4 10.6151
R986 B.n716 B.n715 10.6151
R987 B.n717 B.n716 10.6151
R988 B.n717 B.n0 10.6151
R989 B.n633 B.n632 10.6151
R990 B.n632 B.n631 10.6151
R991 B.n631 B.n32 10.6151
R992 B.n627 B.n32 10.6151
R993 B.n627 B.n626 10.6151
R994 B.n626 B.n625 10.6151
R995 B.n625 B.n34 10.6151
R996 B.n621 B.n34 10.6151
R997 B.n621 B.n620 10.6151
R998 B.n620 B.n619 10.6151
R999 B.n619 B.n36 10.6151
R1000 B.n615 B.n36 10.6151
R1001 B.n615 B.n614 10.6151
R1002 B.n614 B.n613 10.6151
R1003 B.n613 B.n38 10.6151
R1004 B.n609 B.n38 10.6151
R1005 B.n609 B.n608 10.6151
R1006 B.n608 B.n607 10.6151
R1007 B.n607 B.n40 10.6151
R1008 B.n603 B.n40 10.6151
R1009 B.n603 B.n602 10.6151
R1010 B.n602 B.n601 10.6151
R1011 B.n601 B.n42 10.6151
R1012 B.n597 B.n42 10.6151
R1013 B.n597 B.n596 10.6151
R1014 B.n594 B.n46 10.6151
R1015 B.n590 B.n46 10.6151
R1016 B.n590 B.n589 10.6151
R1017 B.n589 B.n588 10.6151
R1018 B.n588 B.n48 10.6151
R1019 B.n584 B.n48 10.6151
R1020 B.n584 B.n583 10.6151
R1021 B.n583 B.n582 10.6151
R1022 B.n582 B.n50 10.6151
R1023 B.n578 B.n577 10.6151
R1024 B.n577 B.n576 10.6151
R1025 B.n576 B.n55 10.6151
R1026 B.n572 B.n55 10.6151
R1027 B.n572 B.n571 10.6151
R1028 B.n571 B.n570 10.6151
R1029 B.n570 B.n57 10.6151
R1030 B.n566 B.n57 10.6151
R1031 B.n566 B.n565 10.6151
R1032 B.n565 B.n564 10.6151
R1033 B.n564 B.n59 10.6151
R1034 B.n560 B.n59 10.6151
R1035 B.n560 B.n559 10.6151
R1036 B.n559 B.n558 10.6151
R1037 B.n558 B.n61 10.6151
R1038 B.n554 B.n61 10.6151
R1039 B.n554 B.n553 10.6151
R1040 B.n553 B.n552 10.6151
R1041 B.n552 B.n63 10.6151
R1042 B.n548 B.n63 10.6151
R1043 B.n548 B.n547 10.6151
R1044 B.n547 B.n546 10.6151
R1045 B.n546 B.n65 10.6151
R1046 B.n542 B.n65 10.6151
R1047 B.n542 B.n541 10.6151
R1048 B.n540 B.n67 10.6151
R1049 B.n536 B.n67 10.6151
R1050 B.n536 B.n535 10.6151
R1051 B.n535 B.n534 10.6151
R1052 B.n534 B.n69 10.6151
R1053 B.n530 B.n69 10.6151
R1054 B.n530 B.n529 10.6151
R1055 B.n529 B.n528 10.6151
R1056 B.n528 B.n71 10.6151
R1057 B.n524 B.n71 10.6151
R1058 B.n524 B.n523 10.6151
R1059 B.n523 B.n522 10.6151
R1060 B.n522 B.n73 10.6151
R1061 B.n518 B.n73 10.6151
R1062 B.n518 B.n517 10.6151
R1063 B.n517 B.n516 10.6151
R1064 B.n516 B.n75 10.6151
R1065 B.n512 B.n75 10.6151
R1066 B.n512 B.n511 10.6151
R1067 B.n511 B.n510 10.6151
R1068 B.n510 B.n77 10.6151
R1069 B.n506 B.n77 10.6151
R1070 B.n506 B.n505 10.6151
R1071 B.n505 B.n504 10.6151
R1072 B.n504 B.n79 10.6151
R1073 B.n500 B.n79 10.6151
R1074 B.n500 B.n499 10.6151
R1075 B.n499 B.n498 10.6151
R1076 B.n498 B.n81 10.6151
R1077 B.n494 B.n81 10.6151
R1078 B.n494 B.n493 10.6151
R1079 B.n493 B.n492 10.6151
R1080 B.n492 B.n83 10.6151
R1081 B.n488 B.n83 10.6151
R1082 B.n488 B.n487 10.6151
R1083 B.n487 B.n486 10.6151
R1084 B.n486 B.n85 10.6151
R1085 B.n482 B.n85 10.6151
R1086 B.n482 B.n481 10.6151
R1087 B.n481 B.n480 10.6151
R1088 B.n480 B.n87 10.6151
R1089 B.n476 B.n87 10.6151
R1090 B.n476 B.n475 10.6151
R1091 B.n475 B.n474 10.6151
R1092 B.n474 B.n89 10.6151
R1093 B.n470 B.n89 10.6151
R1094 B.n470 B.n469 10.6151
R1095 B.n469 B.n468 10.6151
R1096 B.n468 B.n91 10.6151
R1097 B.n464 B.n91 10.6151
R1098 B.n464 B.n463 10.6151
R1099 B.n463 B.n462 10.6151
R1100 B.n462 B.n93 10.6151
R1101 B.n458 B.n93 10.6151
R1102 B.n458 B.n457 10.6151
R1103 B.n457 B.n456 10.6151
R1104 B.n456 B.n95 10.6151
R1105 B.n452 B.n95 10.6151
R1106 B.n452 B.n451 10.6151
R1107 B.n451 B.n450 10.6151
R1108 B.n450 B.n97 10.6151
R1109 B.n446 B.n97 10.6151
R1110 B.n446 B.n445 10.6151
R1111 B.n445 B.n444 10.6151
R1112 B.n444 B.n99 10.6151
R1113 B.n440 B.n99 10.6151
R1114 B.n440 B.n439 10.6151
R1115 B.n439 B.n438 10.6151
R1116 B.n438 B.n101 10.6151
R1117 B.n434 B.n101 10.6151
R1118 B.n434 B.n433 10.6151
R1119 B.n433 B.n432 10.6151
R1120 B.n432 B.n103 10.6151
R1121 B.n428 B.n103 10.6151
R1122 B.n428 B.n427 10.6151
R1123 B.n427 B.n426 10.6151
R1124 B.n426 B.n105 10.6151
R1125 B.n422 B.n105 10.6151
R1126 B.n422 B.n421 10.6151
R1127 B.n421 B.n420 10.6151
R1128 B.n420 B.n107 10.6151
R1129 B.n416 B.n107 10.6151
R1130 B.n416 B.n415 10.6151
R1131 B.n415 B.n414 10.6151
R1132 B.n414 B.n109 10.6151
R1133 B.n410 B.n109 10.6151
R1134 B.n410 B.n409 10.6151
R1135 B.n409 B.n408 10.6151
R1136 B.n408 B.n111 10.6151
R1137 B.n404 B.n111 10.6151
R1138 B.n404 B.n403 10.6151
R1139 B.n403 B.n402 10.6151
R1140 B.n402 B.n113 10.6151
R1141 B.n398 B.n113 10.6151
R1142 B.n398 B.n397 10.6151
R1143 B.n397 B.n396 10.6151
R1144 B.n396 B.n115 10.6151
R1145 B.n392 B.n115 10.6151
R1146 B.n392 B.n391 10.6151
R1147 B.n391 B.n390 10.6151
R1148 B.n390 B.n117 10.6151
R1149 B.n386 B.n117 10.6151
R1150 B.n386 B.n385 10.6151
R1151 B.n385 B.n384 10.6151
R1152 B.n384 B.n119 10.6151
R1153 B.n380 B.n119 10.6151
R1154 B.n380 B.n379 10.6151
R1155 B.n379 B.n378 10.6151
R1156 B.n378 B.n121 10.6151
R1157 B.n374 B.n121 10.6151
R1158 B.n374 B.n373 10.6151
R1159 B.n373 B.n372 10.6151
R1160 B.n372 B.n123 10.6151
R1161 B.n368 B.n123 10.6151
R1162 B.n368 B.n367 10.6151
R1163 B.n185 B.n1 10.6151
R1164 B.n188 B.n185 10.6151
R1165 B.n189 B.n188 10.6151
R1166 B.n190 B.n189 10.6151
R1167 B.n190 B.n183 10.6151
R1168 B.n194 B.n183 10.6151
R1169 B.n195 B.n194 10.6151
R1170 B.n196 B.n195 10.6151
R1171 B.n196 B.n181 10.6151
R1172 B.n200 B.n181 10.6151
R1173 B.n201 B.n200 10.6151
R1174 B.n202 B.n201 10.6151
R1175 B.n202 B.n179 10.6151
R1176 B.n206 B.n179 10.6151
R1177 B.n207 B.n206 10.6151
R1178 B.n208 B.n207 10.6151
R1179 B.n208 B.n177 10.6151
R1180 B.n212 B.n177 10.6151
R1181 B.n213 B.n212 10.6151
R1182 B.n214 B.n213 10.6151
R1183 B.n214 B.n175 10.6151
R1184 B.n218 B.n175 10.6151
R1185 B.n219 B.n218 10.6151
R1186 B.n220 B.n219 10.6151
R1187 B.n220 B.n173 10.6151
R1188 B.n224 B.n173 10.6151
R1189 B.n225 B.n224 10.6151
R1190 B.n226 B.n225 10.6151
R1191 B.n226 B.n171 10.6151
R1192 B.n230 B.n171 10.6151
R1193 B.n231 B.n230 10.6151
R1194 B.n232 B.n231 10.6151
R1195 B.n232 B.n169 10.6151
R1196 B.n236 B.n169 10.6151
R1197 B.n237 B.n236 10.6151
R1198 B.n238 B.n237 10.6151
R1199 B.n238 B.n167 10.6151
R1200 B.n242 B.n167 10.6151
R1201 B.n243 B.n242 10.6151
R1202 B.n244 B.n243 10.6151
R1203 B.n244 B.n165 10.6151
R1204 B.n248 B.n165 10.6151
R1205 B.n249 B.n248 10.6151
R1206 B.n250 B.n249 10.6151
R1207 B.n250 B.n163 10.6151
R1208 B.n254 B.n163 10.6151
R1209 B.n255 B.n254 10.6151
R1210 B.n256 B.n255 10.6151
R1211 B.n256 B.n161 10.6151
R1212 B.n260 B.n161 10.6151
R1213 B.n261 B.n260 10.6151
R1214 B.n262 B.n261 10.6151
R1215 B.n262 B.n159 10.6151
R1216 B.n266 B.n159 10.6151
R1217 B.n267 B.n266 10.6151
R1218 B.n268 B.n267 10.6151
R1219 B.n272 B.n157 10.6151
R1220 B.n273 B.n272 10.6151
R1221 B.n274 B.n273 10.6151
R1222 B.n274 B.n155 10.6151
R1223 B.n278 B.n155 10.6151
R1224 B.n279 B.n278 10.6151
R1225 B.n280 B.n279 10.6151
R1226 B.n280 B.n153 10.6151
R1227 B.n284 B.n153 10.6151
R1228 B.n285 B.n284 10.6151
R1229 B.n286 B.n285 10.6151
R1230 B.n286 B.n151 10.6151
R1231 B.n290 B.n151 10.6151
R1232 B.n291 B.n290 10.6151
R1233 B.n292 B.n291 10.6151
R1234 B.n292 B.n149 10.6151
R1235 B.n296 B.n149 10.6151
R1236 B.n297 B.n296 10.6151
R1237 B.n298 B.n297 10.6151
R1238 B.n298 B.n147 10.6151
R1239 B.n302 B.n147 10.6151
R1240 B.n303 B.n302 10.6151
R1241 B.n304 B.n303 10.6151
R1242 B.n304 B.n145 10.6151
R1243 B.n308 B.n145 10.6151
R1244 B.n311 B.n310 10.6151
R1245 B.n311 B.n141 10.6151
R1246 B.n315 B.n141 10.6151
R1247 B.n316 B.n315 10.6151
R1248 B.n317 B.n316 10.6151
R1249 B.n317 B.n139 10.6151
R1250 B.n321 B.n139 10.6151
R1251 B.n322 B.n321 10.6151
R1252 B.n326 B.n322 10.6151
R1253 B.n330 B.n137 10.6151
R1254 B.n331 B.n330 10.6151
R1255 B.n332 B.n331 10.6151
R1256 B.n332 B.n135 10.6151
R1257 B.n336 B.n135 10.6151
R1258 B.n337 B.n336 10.6151
R1259 B.n338 B.n337 10.6151
R1260 B.n338 B.n133 10.6151
R1261 B.n342 B.n133 10.6151
R1262 B.n343 B.n342 10.6151
R1263 B.n344 B.n343 10.6151
R1264 B.n344 B.n131 10.6151
R1265 B.n348 B.n131 10.6151
R1266 B.n349 B.n348 10.6151
R1267 B.n350 B.n349 10.6151
R1268 B.n350 B.n129 10.6151
R1269 B.n354 B.n129 10.6151
R1270 B.n355 B.n354 10.6151
R1271 B.n356 B.n355 10.6151
R1272 B.n356 B.n127 10.6151
R1273 B.n360 B.n127 10.6151
R1274 B.n361 B.n360 10.6151
R1275 B.n362 B.n361 10.6151
R1276 B.n362 B.n125 10.6151
R1277 B.n366 B.n125 10.6151
R1278 B.n596 B.n595 9.36635
R1279 B.n578 B.n54 9.36635
R1280 B.n309 B.n308 9.36635
R1281 B.n325 B.n137 9.36635
R1282 B.n721 B.n0 8.11757
R1283 B.n721 B.n1 8.11757
R1284 B.n595 B.n594 1.24928
R1285 B.n54 B.n50 1.24928
R1286 B.n310 B.n309 1.24928
R1287 B.n326 B.n325 1.24928
C0 w_n4322_n2332# VDD1 2.24386f
C1 w_n4322_n2332# VN 8.41411f
C2 VP B 2.31071f
C3 VTAIL VDD1 6.55223f
C4 VTAIL VN 5.14897f
C5 VP VDD2 0.564281f
C6 B VDD2 2.10557f
C7 w_n4322_n2332# VP 8.9764f
C8 w_n4322_n2332# B 9.97025f
C9 VTAIL VP 5.16349f
C10 VN VDD1 0.152202f
C11 w_n4322_n2332# VDD2 2.36922f
C12 VTAIL B 2.91131f
C13 VTAIL VDD2 6.6133f
C14 w_n4322_n2332# VTAIL 2.39156f
C15 VP VDD1 4.65195f
C16 VN VP 7.20238f
C17 VDD1 B 2.00126f
C18 VN B 1.36558f
C19 VDD1 VDD2 1.89884f
C20 VN VDD2 4.24194f
C21 VDD2 VSUBS 2.120163f
C22 VDD1 VSUBS 2.6938f
C23 VTAIL VSUBS 0.840605f
C24 VN VSUBS 6.88096f
C25 VP VSUBS 3.544374f
C26 B VSUBS 5.445867f
C27 w_n4322_n2332# VSUBS 0.125459p
C28 B.n0 VSUBS 0.009273f
C29 B.n1 VSUBS 0.009273f
C30 B.n2 VSUBS 0.013714f
C31 B.n3 VSUBS 0.010509f
C32 B.n4 VSUBS 0.010509f
C33 B.n5 VSUBS 0.010509f
C34 B.n6 VSUBS 0.010509f
C35 B.n7 VSUBS 0.010509f
C36 B.n8 VSUBS 0.010509f
C37 B.n9 VSUBS 0.010509f
C38 B.n10 VSUBS 0.010509f
C39 B.n11 VSUBS 0.010509f
C40 B.n12 VSUBS 0.010509f
C41 B.n13 VSUBS 0.010509f
C42 B.n14 VSUBS 0.010509f
C43 B.n15 VSUBS 0.010509f
C44 B.n16 VSUBS 0.010509f
C45 B.n17 VSUBS 0.010509f
C46 B.n18 VSUBS 0.010509f
C47 B.n19 VSUBS 0.010509f
C48 B.n20 VSUBS 0.010509f
C49 B.n21 VSUBS 0.010509f
C50 B.n22 VSUBS 0.010509f
C51 B.n23 VSUBS 0.010509f
C52 B.n24 VSUBS 0.010509f
C53 B.n25 VSUBS 0.010509f
C54 B.n26 VSUBS 0.010509f
C55 B.n27 VSUBS 0.010509f
C56 B.n28 VSUBS 0.010509f
C57 B.n29 VSUBS 0.010509f
C58 B.n30 VSUBS 0.02457f
C59 B.n31 VSUBS 0.010509f
C60 B.n32 VSUBS 0.010509f
C61 B.n33 VSUBS 0.010509f
C62 B.n34 VSUBS 0.010509f
C63 B.n35 VSUBS 0.010509f
C64 B.n36 VSUBS 0.010509f
C65 B.n37 VSUBS 0.010509f
C66 B.n38 VSUBS 0.010509f
C67 B.n39 VSUBS 0.010509f
C68 B.n40 VSUBS 0.010509f
C69 B.n41 VSUBS 0.010509f
C70 B.n42 VSUBS 0.010509f
C71 B.n43 VSUBS 0.010509f
C72 B.t4 VSUBS 0.307049f
C73 B.t5 VSUBS 0.349306f
C74 B.t3 VSUBS 1.89224f
C75 B.n44 VSUBS 0.209969f
C76 B.n45 VSUBS 0.114512f
C77 B.n46 VSUBS 0.010509f
C78 B.n47 VSUBS 0.010509f
C79 B.n48 VSUBS 0.010509f
C80 B.n49 VSUBS 0.010509f
C81 B.n50 VSUBS 0.005873f
C82 B.n51 VSUBS 0.010509f
C83 B.t7 VSUBS 0.307047f
C84 B.t8 VSUBS 0.349304f
C85 B.t6 VSUBS 1.89224f
C86 B.n52 VSUBS 0.209971f
C87 B.n53 VSUBS 0.114513f
C88 B.n54 VSUBS 0.024349f
C89 B.n55 VSUBS 0.010509f
C90 B.n56 VSUBS 0.010509f
C91 B.n57 VSUBS 0.010509f
C92 B.n58 VSUBS 0.010509f
C93 B.n59 VSUBS 0.010509f
C94 B.n60 VSUBS 0.010509f
C95 B.n61 VSUBS 0.010509f
C96 B.n62 VSUBS 0.010509f
C97 B.n63 VSUBS 0.010509f
C98 B.n64 VSUBS 0.010509f
C99 B.n65 VSUBS 0.010509f
C100 B.n66 VSUBS 0.025194f
C101 B.n67 VSUBS 0.010509f
C102 B.n68 VSUBS 0.010509f
C103 B.n69 VSUBS 0.010509f
C104 B.n70 VSUBS 0.010509f
C105 B.n71 VSUBS 0.010509f
C106 B.n72 VSUBS 0.010509f
C107 B.n73 VSUBS 0.010509f
C108 B.n74 VSUBS 0.010509f
C109 B.n75 VSUBS 0.010509f
C110 B.n76 VSUBS 0.010509f
C111 B.n77 VSUBS 0.010509f
C112 B.n78 VSUBS 0.010509f
C113 B.n79 VSUBS 0.010509f
C114 B.n80 VSUBS 0.010509f
C115 B.n81 VSUBS 0.010509f
C116 B.n82 VSUBS 0.010509f
C117 B.n83 VSUBS 0.010509f
C118 B.n84 VSUBS 0.010509f
C119 B.n85 VSUBS 0.010509f
C120 B.n86 VSUBS 0.010509f
C121 B.n87 VSUBS 0.010509f
C122 B.n88 VSUBS 0.010509f
C123 B.n89 VSUBS 0.010509f
C124 B.n90 VSUBS 0.010509f
C125 B.n91 VSUBS 0.010509f
C126 B.n92 VSUBS 0.010509f
C127 B.n93 VSUBS 0.010509f
C128 B.n94 VSUBS 0.010509f
C129 B.n95 VSUBS 0.010509f
C130 B.n96 VSUBS 0.010509f
C131 B.n97 VSUBS 0.010509f
C132 B.n98 VSUBS 0.010509f
C133 B.n99 VSUBS 0.010509f
C134 B.n100 VSUBS 0.010509f
C135 B.n101 VSUBS 0.010509f
C136 B.n102 VSUBS 0.010509f
C137 B.n103 VSUBS 0.010509f
C138 B.n104 VSUBS 0.010509f
C139 B.n105 VSUBS 0.010509f
C140 B.n106 VSUBS 0.010509f
C141 B.n107 VSUBS 0.010509f
C142 B.n108 VSUBS 0.010509f
C143 B.n109 VSUBS 0.010509f
C144 B.n110 VSUBS 0.010509f
C145 B.n111 VSUBS 0.010509f
C146 B.n112 VSUBS 0.010509f
C147 B.n113 VSUBS 0.010509f
C148 B.n114 VSUBS 0.010509f
C149 B.n115 VSUBS 0.010509f
C150 B.n116 VSUBS 0.010509f
C151 B.n117 VSUBS 0.010509f
C152 B.n118 VSUBS 0.010509f
C153 B.n119 VSUBS 0.010509f
C154 B.n120 VSUBS 0.010509f
C155 B.n121 VSUBS 0.010509f
C156 B.n122 VSUBS 0.010509f
C157 B.n123 VSUBS 0.010509f
C158 B.n124 VSUBS 0.02457f
C159 B.n125 VSUBS 0.010509f
C160 B.n126 VSUBS 0.010509f
C161 B.n127 VSUBS 0.010509f
C162 B.n128 VSUBS 0.010509f
C163 B.n129 VSUBS 0.010509f
C164 B.n130 VSUBS 0.010509f
C165 B.n131 VSUBS 0.010509f
C166 B.n132 VSUBS 0.010509f
C167 B.n133 VSUBS 0.010509f
C168 B.n134 VSUBS 0.010509f
C169 B.n135 VSUBS 0.010509f
C170 B.n136 VSUBS 0.010509f
C171 B.n137 VSUBS 0.009891f
C172 B.n138 VSUBS 0.010509f
C173 B.n139 VSUBS 0.010509f
C174 B.n140 VSUBS 0.010509f
C175 B.n141 VSUBS 0.010509f
C176 B.n142 VSUBS 0.010509f
C177 B.t2 VSUBS 0.307049f
C178 B.t1 VSUBS 0.349306f
C179 B.t0 VSUBS 1.89224f
C180 B.n143 VSUBS 0.209969f
C181 B.n144 VSUBS 0.114512f
C182 B.n145 VSUBS 0.010509f
C183 B.n146 VSUBS 0.010509f
C184 B.n147 VSUBS 0.010509f
C185 B.n148 VSUBS 0.010509f
C186 B.n149 VSUBS 0.010509f
C187 B.n150 VSUBS 0.010509f
C188 B.n151 VSUBS 0.010509f
C189 B.n152 VSUBS 0.010509f
C190 B.n153 VSUBS 0.010509f
C191 B.n154 VSUBS 0.010509f
C192 B.n155 VSUBS 0.010509f
C193 B.n156 VSUBS 0.010509f
C194 B.n157 VSUBS 0.025194f
C195 B.n158 VSUBS 0.010509f
C196 B.n159 VSUBS 0.010509f
C197 B.n160 VSUBS 0.010509f
C198 B.n161 VSUBS 0.010509f
C199 B.n162 VSUBS 0.010509f
C200 B.n163 VSUBS 0.010509f
C201 B.n164 VSUBS 0.010509f
C202 B.n165 VSUBS 0.010509f
C203 B.n166 VSUBS 0.010509f
C204 B.n167 VSUBS 0.010509f
C205 B.n168 VSUBS 0.010509f
C206 B.n169 VSUBS 0.010509f
C207 B.n170 VSUBS 0.010509f
C208 B.n171 VSUBS 0.010509f
C209 B.n172 VSUBS 0.010509f
C210 B.n173 VSUBS 0.010509f
C211 B.n174 VSUBS 0.010509f
C212 B.n175 VSUBS 0.010509f
C213 B.n176 VSUBS 0.010509f
C214 B.n177 VSUBS 0.010509f
C215 B.n178 VSUBS 0.010509f
C216 B.n179 VSUBS 0.010509f
C217 B.n180 VSUBS 0.010509f
C218 B.n181 VSUBS 0.010509f
C219 B.n182 VSUBS 0.010509f
C220 B.n183 VSUBS 0.010509f
C221 B.n184 VSUBS 0.010509f
C222 B.n185 VSUBS 0.010509f
C223 B.n186 VSUBS 0.010509f
C224 B.n187 VSUBS 0.010509f
C225 B.n188 VSUBS 0.010509f
C226 B.n189 VSUBS 0.010509f
C227 B.n190 VSUBS 0.010509f
C228 B.n191 VSUBS 0.010509f
C229 B.n192 VSUBS 0.010509f
C230 B.n193 VSUBS 0.010509f
C231 B.n194 VSUBS 0.010509f
C232 B.n195 VSUBS 0.010509f
C233 B.n196 VSUBS 0.010509f
C234 B.n197 VSUBS 0.010509f
C235 B.n198 VSUBS 0.010509f
C236 B.n199 VSUBS 0.010509f
C237 B.n200 VSUBS 0.010509f
C238 B.n201 VSUBS 0.010509f
C239 B.n202 VSUBS 0.010509f
C240 B.n203 VSUBS 0.010509f
C241 B.n204 VSUBS 0.010509f
C242 B.n205 VSUBS 0.010509f
C243 B.n206 VSUBS 0.010509f
C244 B.n207 VSUBS 0.010509f
C245 B.n208 VSUBS 0.010509f
C246 B.n209 VSUBS 0.010509f
C247 B.n210 VSUBS 0.010509f
C248 B.n211 VSUBS 0.010509f
C249 B.n212 VSUBS 0.010509f
C250 B.n213 VSUBS 0.010509f
C251 B.n214 VSUBS 0.010509f
C252 B.n215 VSUBS 0.010509f
C253 B.n216 VSUBS 0.010509f
C254 B.n217 VSUBS 0.010509f
C255 B.n218 VSUBS 0.010509f
C256 B.n219 VSUBS 0.010509f
C257 B.n220 VSUBS 0.010509f
C258 B.n221 VSUBS 0.010509f
C259 B.n222 VSUBS 0.010509f
C260 B.n223 VSUBS 0.010509f
C261 B.n224 VSUBS 0.010509f
C262 B.n225 VSUBS 0.010509f
C263 B.n226 VSUBS 0.010509f
C264 B.n227 VSUBS 0.010509f
C265 B.n228 VSUBS 0.010509f
C266 B.n229 VSUBS 0.010509f
C267 B.n230 VSUBS 0.010509f
C268 B.n231 VSUBS 0.010509f
C269 B.n232 VSUBS 0.010509f
C270 B.n233 VSUBS 0.010509f
C271 B.n234 VSUBS 0.010509f
C272 B.n235 VSUBS 0.010509f
C273 B.n236 VSUBS 0.010509f
C274 B.n237 VSUBS 0.010509f
C275 B.n238 VSUBS 0.010509f
C276 B.n239 VSUBS 0.010509f
C277 B.n240 VSUBS 0.010509f
C278 B.n241 VSUBS 0.010509f
C279 B.n242 VSUBS 0.010509f
C280 B.n243 VSUBS 0.010509f
C281 B.n244 VSUBS 0.010509f
C282 B.n245 VSUBS 0.010509f
C283 B.n246 VSUBS 0.010509f
C284 B.n247 VSUBS 0.010509f
C285 B.n248 VSUBS 0.010509f
C286 B.n249 VSUBS 0.010509f
C287 B.n250 VSUBS 0.010509f
C288 B.n251 VSUBS 0.010509f
C289 B.n252 VSUBS 0.010509f
C290 B.n253 VSUBS 0.010509f
C291 B.n254 VSUBS 0.010509f
C292 B.n255 VSUBS 0.010509f
C293 B.n256 VSUBS 0.010509f
C294 B.n257 VSUBS 0.010509f
C295 B.n258 VSUBS 0.010509f
C296 B.n259 VSUBS 0.010509f
C297 B.n260 VSUBS 0.010509f
C298 B.n261 VSUBS 0.010509f
C299 B.n262 VSUBS 0.010509f
C300 B.n263 VSUBS 0.010509f
C301 B.n264 VSUBS 0.010509f
C302 B.n265 VSUBS 0.010509f
C303 B.n266 VSUBS 0.010509f
C304 B.n267 VSUBS 0.010509f
C305 B.n268 VSUBS 0.02457f
C306 B.n269 VSUBS 0.02457f
C307 B.n270 VSUBS 0.025194f
C308 B.n271 VSUBS 0.010509f
C309 B.n272 VSUBS 0.010509f
C310 B.n273 VSUBS 0.010509f
C311 B.n274 VSUBS 0.010509f
C312 B.n275 VSUBS 0.010509f
C313 B.n276 VSUBS 0.010509f
C314 B.n277 VSUBS 0.010509f
C315 B.n278 VSUBS 0.010509f
C316 B.n279 VSUBS 0.010509f
C317 B.n280 VSUBS 0.010509f
C318 B.n281 VSUBS 0.010509f
C319 B.n282 VSUBS 0.010509f
C320 B.n283 VSUBS 0.010509f
C321 B.n284 VSUBS 0.010509f
C322 B.n285 VSUBS 0.010509f
C323 B.n286 VSUBS 0.010509f
C324 B.n287 VSUBS 0.010509f
C325 B.n288 VSUBS 0.010509f
C326 B.n289 VSUBS 0.010509f
C327 B.n290 VSUBS 0.010509f
C328 B.n291 VSUBS 0.010509f
C329 B.n292 VSUBS 0.010509f
C330 B.n293 VSUBS 0.010509f
C331 B.n294 VSUBS 0.010509f
C332 B.n295 VSUBS 0.010509f
C333 B.n296 VSUBS 0.010509f
C334 B.n297 VSUBS 0.010509f
C335 B.n298 VSUBS 0.010509f
C336 B.n299 VSUBS 0.010509f
C337 B.n300 VSUBS 0.010509f
C338 B.n301 VSUBS 0.010509f
C339 B.n302 VSUBS 0.010509f
C340 B.n303 VSUBS 0.010509f
C341 B.n304 VSUBS 0.010509f
C342 B.n305 VSUBS 0.010509f
C343 B.n306 VSUBS 0.010509f
C344 B.n307 VSUBS 0.010509f
C345 B.n308 VSUBS 0.009891f
C346 B.n309 VSUBS 0.024349f
C347 B.n310 VSUBS 0.005873f
C348 B.n311 VSUBS 0.010509f
C349 B.n312 VSUBS 0.010509f
C350 B.n313 VSUBS 0.010509f
C351 B.n314 VSUBS 0.010509f
C352 B.n315 VSUBS 0.010509f
C353 B.n316 VSUBS 0.010509f
C354 B.n317 VSUBS 0.010509f
C355 B.n318 VSUBS 0.010509f
C356 B.n319 VSUBS 0.010509f
C357 B.n320 VSUBS 0.010509f
C358 B.n321 VSUBS 0.010509f
C359 B.n322 VSUBS 0.010509f
C360 B.t11 VSUBS 0.307047f
C361 B.t10 VSUBS 0.349304f
C362 B.t9 VSUBS 1.89224f
C363 B.n323 VSUBS 0.209971f
C364 B.n324 VSUBS 0.114513f
C365 B.n325 VSUBS 0.024349f
C366 B.n326 VSUBS 0.005873f
C367 B.n327 VSUBS 0.010509f
C368 B.n328 VSUBS 0.010509f
C369 B.n329 VSUBS 0.010509f
C370 B.n330 VSUBS 0.010509f
C371 B.n331 VSUBS 0.010509f
C372 B.n332 VSUBS 0.010509f
C373 B.n333 VSUBS 0.010509f
C374 B.n334 VSUBS 0.010509f
C375 B.n335 VSUBS 0.010509f
C376 B.n336 VSUBS 0.010509f
C377 B.n337 VSUBS 0.010509f
C378 B.n338 VSUBS 0.010509f
C379 B.n339 VSUBS 0.010509f
C380 B.n340 VSUBS 0.010509f
C381 B.n341 VSUBS 0.010509f
C382 B.n342 VSUBS 0.010509f
C383 B.n343 VSUBS 0.010509f
C384 B.n344 VSUBS 0.010509f
C385 B.n345 VSUBS 0.010509f
C386 B.n346 VSUBS 0.010509f
C387 B.n347 VSUBS 0.010509f
C388 B.n348 VSUBS 0.010509f
C389 B.n349 VSUBS 0.010509f
C390 B.n350 VSUBS 0.010509f
C391 B.n351 VSUBS 0.010509f
C392 B.n352 VSUBS 0.010509f
C393 B.n353 VSUBS 0.010509f
C394 B.n354 VSUBS 0.010509f
C395 B.n355 VSUBS 0.010509f
C396 B.n356 VSUBS 0.010509f
C397 B.n357 VSUBS 0.010509f
C398 B.n358 VSUBS 0.010509f
C399 B.n359 VSUBS 0.010509f
C400 B.n360 VSUBS 0.010509f
C401 B.n361 VSUBS 0.010509f
C402 B.n362 VSUBS 0.010509f
C403 B.n363 VSUBS 0.010509f
C404 B.n364 VSUBS 0.010509f
C405 B.n365 VSUBS 0.025194f
C406 B.n366 VSUBS 0.023975f
C407 B.n367 VSUBS 0.025789f
C408 B.n368 VSUBS 0.010509f
C409 B.n369 VSUBS 0.010509f
C410 B.n370 VSUBS 0.010509f
C411 B.n371 VSUBS 0.010509f
C412 B.n372 VSUBS 0.010509f
C413 B.n373 VSUBS 0.010509f
C414 B.n374 VSUBS 0.010509f
C415 B.n375 VSUBS 0.010509f
C416 B.n376 VSUBS 0.010509f
C417 B.n377 VSUBS 0.010509f
C418 B.n378 VSUBS 0.010509f
C419 B.n379 VSUBS 0.010509f
C420 B.n380 VSUBS 0.010509f
C421 B.n381 VSUBS 0.010509f
C422 B.n382 VSUBS 0.010509f
C423 B.n383 VSUBS 0.010509f
C424 B.n384 VSUBS 0.010509f
C425 B.n385 VSUBS 0.010509f
C426 B.n386 VSUBS 0.010509f
C427 B.n387 VSUBS 0.010509f
C428 B.n388 VSUBS 0.010509f
C429 B.n389 VSUBS 0.010509f
C430 B.n390 VSUBS 0.010509f
C431 B.n391 VSUBS 0.010509f
C432 B.n392 VSUBS 0.010509f
C433 B.n393 VSUBS 0.010509f
C434 B.n394 VSUBS 0.010509f
C435 B.n395 VSUBS 0.010509f
C436 B.n396 VSUBS 0.010509f
C437 B.n397 VSUBS 0.010509f
C438 B.n398 VSUBS 0.010509f
C439 B.n399 VSUBS 0.010509f
C440 B.n400 VSUBS 0.010509f
C441 B.n401 VSUBS 0.010509f
C442 B.n402 VSUBS 0.010509f
C443 B.n403 VSUBS 0.010509f
C444 B.n404 VSUBS 0.010509f
C445 B.n405 VSUBS 0.010509f
C446 B.n406 VSUBS 0.010509f
C447 B.n407 VSUBS 0.010509f
C448 B.n408 VSUBS 0.010509f
C449 B.n409 VSUBS 0.010509f
C450 B.n410 VSUBS 0.010509f
C451 B.n411 VSUBS 0.010509f
C452 B.n412 VSUBS 0.010509f
C453 B.n413 VSUBS 0.010509f
C454 B.n414 VSUBS 0.010509f
C455 B.n415 VSUBS 0.010509f
C456 B.n416 VSUBS 0.010509f
C457 B.n417 VSUBS 0.010509f
C458 B.n418 VSUBS 0.010509f
C459 B.n419 VSUBS 0.010509f
C460 B.n420 VSUBS 0.010509f
C461 B.n421 VSUBS 0.010509f
C462 B.n422 VSUBS 0.010509f
C463 B.n423 VSUBS 0.010509f
C464 B.n424 VSUBS 0.010509f
C465 B.n425 VSUBS 0.010509f
C466 B.n426 VSUBS 0.010509f
C467 B.n427 VSUBS 0.010509f
C468 B.n428 VSUBS 0.010509f
C469 B.n429 VSUBS 0.010509f
C470 B.n430 VSUBS 0.010509f
C471 B.n431 VSUBS 0.010509f
C472 B.n432 VSUBS 0.010509f
C473 B.n433 VSUBS 0.010509f
C474 B.n434 VSUBS 0.010509f
C475 B.n435 VSUBS 0.010509f
C476 B.n436 VSUBS 0.010509f
C477 B.n437 VSUBS 0.010509f
C478 B.n438 VSUBS 0.010509f
C479 B.n439 VSUBS 0.010509f
C480 B.n440 VSUBS 0.010509f
C481 B.n441 VSUBS 0.010509f
C482 B.n442 VSUBS 0.010509f
C483 B.n443 VSUBS 0.010509f
C484 B.n444 VSUBS 0.010509f
C485 B.n445 VSUBS 0.010509f
C486 B.n446 VSUBS 0.010509f
C487 B.n447 VSUBS 0.010509f
C488 B.n448 VSUBS 0.010509f
C489 B.n449 VSUBS 0.010509f
C490 B.n450 VSUBS 0.010509f
C491 B.n451 VSUBS 0.010509f
C492 B.n452 VSUBS 0.010509f
C493 B.n453 VSUBS 0.010509f
C494 B.n454 VSUBS 0.010509f
C495 B.n455 VSUBS 0.010509f
C496 B.n456 VSUBS 0.010509f
C497 B.n457 VSUBS 0.010509f
C498 B.n458 VSUBS 0.010509f
C499 B.n459 VSUBS 0.010509f
C500 B.n460 VSUBS 0.010509f
C501 B.n461 VSUBS 0.010509f
C502 B.n462 VSUBS 0.010509f
C503 B.n463 VSUBS 0.010509f
C504 B.n464 VSUBS 0.010509f
C505 B.n465 VSUBS 0.010509f
C506 B.n466 VSUBS 0.010509f
C507 B.n467 VSUBS 0.010509f
C508 B.n468 VSUBS 0.010509f
C509 B.n469 VSUBS 0.010509f
C510 B.n470 VSUBS 0.010509f
C511 B.n471 VSUBS 0.010509f
C512 B.n472 VSUBS 0.010509f
C513 B.n473 VSUBS 0.010509f
C514 B.n474 VSUBS 0.010509f
C515 B.n475 VSUBS 0.010509f
C516 B.n476 VSUBS 0.010509f
C517 B.n477 VSUBS 0.010509f
C518 B.n478 VSUBS 0.010509f
C519 B.n479 VSUBS 0.010509f
C520 B.n480 VSUBS 0.010509f
C521 B.n481 VSUBS 0.010509f
C522 B.n482 VSUBS 0.010509f
C523 B.n483 VSUBS 0.010509f
C524 B.n484 VSUBS 0.010509f
C525 B.n485 VSUBS 0.010509f
C526 B.n486 VSUBS 0.010509f
C527 B.n487 VSUBS 0.010509f
C528 B.n488 VSUBS 0.010509f
C529 B.n489 VSUBS 0.010509f
C530 B.n490 VSUBS 0.010509f
C531 B.n491 VSUBS 0.010509f
C532 B.n492 VSUBS 0.010509f
C533 B.n493 VSUBS 0.010509f
C534 B.n494 VSUBS 0.010509f
C535 B.n495 VSUBS 0.010509f
C536 B.n496 VSUBS 0.010509f
C537 B.n497 VSUBS 0.010509f
C538 B.n498 VSUBS 0.010509f
C539 B.n499 VSUBS 0.010509f
C540 B.n500 VSUBS 0.010509f
C541 B.n501 VSUBS 0.010509f
C542 B.n502 VSUBS 0.010509f
C543 B.n503 VSUBS 0.010509f
C544 B.n504 VSUBS 0.010509f
C545 B.n505 VSUBS 0.010509f
C546 B.n506 VSUBS 0.010509f
C547 B.n507 VSUBS 0.010509f
C548 B.n508 VSUBS 0.010509f
C549 B.n509 VSUBS 0.010509f
C550 B.n510 VSUBS 0.010509f
C551 B.n511 VSUBS 0.010509f
C552 B.n512 VSUBS 0.010509f
C553 B.n513 VSUBS 0.010509f
C554 B.n514 VSUBS 0.010509f
C555 B.n515 VSUBS 0.010509f
C556 B.n516 VSUBS 0.010509f
C557 B.n517 VSUBS 0.010509f
C558 B.n518 VSUBS 0.010509f
C559 B.n519 VSUBS 0.010509f
C560 B.n520 VSUBS 0.010509f
C561 B.n521 VSUBS 0.010509f
C562 B.n522 VSUBS 0.010509f
C563 B.n523 VSUBS 0.010509f
C564 B.n524 VSUBS 0.010509f
C565 B.n525 VSUBS 0.010509f
C566 B.n526 VSUBS 0.010509f
C567 B.n527 VSUBS 0.010509f
C568 B.n528 VSUBS 0.010509f
C569 B.n529 VSUBS 0.010509f
C570 B.n530 VSUBS 0.010509f
C571 B.n531 VSUBS 0.010509f
C572 B.n532 VSUBS 0.010509f
C573 B.n533 VSUBS 0.010509f
C574 B.n534 VSUBS 0.010509f
C575 B.n535 VSUBS 0.010509f
C576 B.n536 VSUBS 0.010509f
C577 B.n537 VSUBS 0.010509f
C578 B.n538 VSUBS 0.010509f
C579 B.n539 VSUBS 0.02457f
C580 B.n540 VSUBS 0.02457f
C581 B.n541 VSUBS 0.025194f
C582 B.n542 VSUBS 0.010509f
C583 B.n543 VSUBS 0.010509f
C584 B.n544 VSUBS 0.010509f
C585 B.n545 VSUBS 0.010509f
C586 B.n546 VSUBS 0.010509f
C587 B.n547 VSUBS 0.010509f
C588 B.n548 VSUBS 0.010509f
C589 B.n549 VSUBS 0.010509f
C590 B.n550 VSUBS 0.010509f
C591 B.n551 VSUBS 0.010509f
C592 B.n552 VSUBS 0.010509f
C593 B.n553 VSUBS 0.010509f
C594 B.n554 VSUBS 0.010509f
C595 B.n555 VSUBS 0.010509f
C596 B.n556 VSUBS 0.010509f
C597 B.n557 VSUBS 0.010509f
C598 B.n558 VSUBS 0.010509f
C599 B.n559 VSUBS 0.010509f
C600 B.n560 VSUBS 0.010509f
C601 B.n561 VSUBS 0.010509f
C602 B.n562 VSUBS 0.010509f
C603 B.n563 VSUBS 0.010509f
C604 B.n564 VSUBS 0.010509f
C605 B.n565 VSUBS 0.010509f
C606 B.n566 VSUBS 0.010509f
C607 B.n567 VSUBS 0.010509f
C608 B.n568 VSUBS 0.010509f
C609 B.n569 VSUBS 0.010509f
C610 B.n570 VSUBS 0.010509f
C611 B.n571 VSUBS 0.010509f
C612 B.n572 VSUBS 0.010509f
C613 B.n573 VSUBS 0.010509f
C614 B.n574 VSUBS 0.010509f
C615 B.n575 VSUBS 0.010509f
C616 B.n576 VSUBS 0.010509f
C617 B.n577 VSUBS 0.010509f
C618 B.n578 VSUBS 0.009891f
C619 B.n579 VSUBS 0.010509f
C620 B.n580 VSUBS 0.010509f
C621 B.n581 VSUBS 0.010509f
C622 B.n582 VSUBS 0.010509f
C623 B.n583 VSUBS 0.010509f
C624 B.n584 VSUBS 0.010509f
C625 B.n585 VSUBS 0.010509f
C626 B.n586 VSUBS 0.010509f
C627 B.n587 VSUBS 0.010509f
C628 B.n588 VSUBS 0.010509f
C629 B.n589 VSUBS 0.010509f
C630 B.n590 VSUBS 0.010509f
C631 B.n591 VSUBS 0.010509f
C632 B.n592 VSUBS 0.010509f
C633 B.n593 VSUBS 0.010509f
C634 B.n594 VSUBS 0.005873f
C635 B.n595 VSUBS 0.024349f
C636 B.n596 VSUBS 0.009891f
C637 B.n597 VSUBS 0.010509f
C638 B.n598 VSUBS 0.010509f
C639 B.n599 VSUBS 0.010509f
C640 B.n600 VSUBS 0.010509f
C641 B.n601 VSUBS 0.010509f
C642 B.n602 VSUBS 0.010509f
C643 B.n603 VSUBS 0.010509f
C644 B.n604 VSUBS 0.010509f
C645 B.n605 VSUBS 0.010509f
C646 B.n606 VSUBS 0.010509f
C647 B.n607 VSUBS 0.010509f
C648 B.n608 VSUBS 0.010509f
C649 B.n609 VSUBS 0.010509f
C650 B.n610 VSUBS 0.010509f
C651 B.n611 VSUBS 0.010509f
C652 B.n612 VSUBS 0.010509f
C653 B.n613 VSUBS 0.010509f
C654 B.n614 VSUBS 0.010509f
C655 B.n615 VSUBS 0.010509f
C656 B.n616 VSUBS 0.010509f
C657 B.n617 VSUBS 0.010509f
C658 B.n618 VSUBS 0.010509f
C659 B.n619 VSUBS 0.010509f
C660 B.n620 VSUBS 0.010509f
C661 B.n621 VSUBS 0.010509f
C662 B.n622 VSUBS 0.010509f
C663 B.n623 VSUBS 0.010509f
C664 B.n624 VSUBS 0.010509f
C665 B.n625 VSUBS 0.010509f
C666 B.n626 VSUBS 0.010509f
C667 B.n627 VSUBS 0.010509f
C668 B.n628 VSUBS 0.010509f
C669 B.n629 VSUBS 0.010509f
C670 B.n630 VSUBS 0.010509f
C671 B.n631 VSUBS 0.010509f
C672 B.n632 VSUBS 0.010509f
C673 B.n633 VSUBS 0.025194f
C674 B.n634 VSUBS 0.025194f
C675 B.n635 VSUBS 0.02457f
C676 B.n636 VSUBS 0.010509f
C677 B.n637 VSUBS 0.010509f
C678 B.n638 VSUBS 0.010509f
C679 B.n639 VSUBS 0.010509f
C680 B.n640 VSUBS 0.010509f
C681 B.n641 VSUBS 0.010509f
C682 B.n642 VSUBS 0.010509f
C683 B.n643 VSUBS 0.010509f
C684 B.n644 VSUBS 0.010509f
C685 B.n645 VSUBS 0.010509f
C686 B.n646 VSUBS 0.010509f
C687 B.n647 VSUBS 0.010509f
C688 B.n648 VSUBS 0.010509f
C689 B.n649 VSUBS 0.010509f
C690 B.n650 VSUBS 0.010509f
C691 B.n651 VSUBS 0.010509f
C692 B.n652 VSUBS 0.010509f
C693 B.n653 VSUBS 0.010509f
C694 B.n654 VSUBS 0.010509f
C695 B.n655 VSUBS 0.010509f
C696 B.n656 VSUBS 0.010509f
C697 B.n657 VSUBS 0.010509f
C698 B.n658 VSUBS 0.010509f
C699 B.n659 VSUBS 0.010509f
C700 B.n660 VSUBS 0.010509f
C701 B.n661 VSUBS 0.010509f
C702 B.n662 VSUBS 0.010509f
C703 B.n663 VSUBS 0.010509f
C704 B.n664 VSUBS 0.010509f
C705 B.n665 VSUBS 0.010509f
C706 B.n666 VSUBS 0.010509f
C707 B.n667 VSUBS 0.010509f
C708 B.n668 VSUBS 0.010509f
C709 B.n669 VSUBS 0.010509f
C710 B.n670 VSUBS 0.010509f
C711 B.n671 VSUBS 0.010509f
C712 B.n672 VSUBS 0.010509f
C713 B.n673 VSUBS 0.010509f
C714 B.n674 VSUBS 0.010509f
C715 B.n675 VSUBS 0.010509f
C716 B.n676 VSUBS 0.010509f
C717 B.n677 VSUBS 0.010509f
C718 B.n678 VSUBS 0.010509f
C719 B.n679 VSUBS 0.010509f
C720 B.n680 VSUBS 0.010509f
C721 B.n681 VSUBS 0.010509f
C722 B.n682 VSUBS 0.010509f
C723 B.n683 VSUBS 0.010509f
C724 B.n684 VSUBS 0.010509f
C725 B.n685 VSUBS 0.010509f
C726 B.n686 VSUBS 0.010509f
C727 B.n687 VSUBS 0.010509f
C728 B.n688 VSUBS 0.010509f
C729 B.n689 VSUBS 0.010509f
C730 B.n690 VSUBS 0.010509f
C731 B.n691 VSUBS 0.010509f
C732 B.n692 VSUBS 0.010509f
C733 B.n693 VSUBS 0.010509f
C734 B.n694 VSUBS 0.010509f
C735 B.n695 VSUBS 0.010509f
C736 B.n696 VSUBS 0.010509f
C737 B.n697 VSUBS 0.010509f
C738 B.n698 VSUBS 0.010509f
C739 B.n699 VSUBS 0.010509f
C740 B.n700 VSUBS 0.010509f
C741 B.n701 VSUBS 0.010509f
C742 B.n702 VSUBS 0.010509f
C743 B.n703 VSUBS 0.010509f
C744 B.n704 VSUBS 0.010509f
C745 B.n705 VSUBS 0.010509f
C746 B.n706 VSUBS 0.010509f
C747 B.n707 VSUBS 0.010509f
C748 B.n708 VSUBS 0.010509f
C749 B.n709 VSUBS 0.010509f
C750 B.n710 VSUBS 0.010509f
C751 B.n711 VSUBS 0.010509f
C752 B.n712 VSUBS 0.010509f
C753 B.n713 VSUBS 0.010509f
C754 B.n714 VSUBS 0.010509f
C755 B.n715 VSUBS 0.010509f
C756 B.n716 VSUBS 0.010509f
C757 B.n717 VSUBS 0.010509f
C758 B.n718 VSUBS 0.010509f
C759 B.n719 VSUBS 0.013714f
C760 B.n720 VSUBS 0.014609f
C761 B.n721 VSUBS 0.029051f
C762 VDD2.t2 VSUBS 1.5551f
C763 VDD2.t5 VSUBS 0.165408f
C764 VDD2.t4 VSUBS 0.165408f
C765 VDD2.n0 VSUBS 1.16337f
C766 VDD2.n1 VSUBS 4.32693f
C767 VDD2.t3 VSUBS 1.53162f
C768 VDD2.n2 VSUBS 3.59904f
C769 VDD2.t0 VSUBS 0.165408f
C770 VDD2.t1 VSUBS 0.165408f
C771 VDD2.n3 VSUBS 1.16333f
C772 VN.n0 VSUBS 0.057721f
C773 VN.t1 VSUBS 2.15262f
C774 VN.n1 VSUBS 0.058509f
C775 VN.n2 VSUBS 0.030677f
C776 VN.n3 VSUBS 0.057461f
C777 VN.t3 VSUBS 2.59333f
C778 VN.n4 VSUBS 0.866039f
C779 VN.t0 VSUBS 2.15262f
C780 VN.n5 VSUBS 0.894275f
C781 VN.n6 VSUBS 0.043276f
C782 VN.n7 VSUBS 0.40351f
C783 VN.n8 VSUBS 0.030677f
C784 VN.n9 VSUBS 0.030677f
C785 VN.n10 VSUBS 0.057461f
C786 VN.n11 VSUBS 0.053002f
C787 VN.n12 VSUBS 0.035907f
C788 VN.n13 VSUBS 0.030677f
C789 VN.n14 VSUBS 0.030677f
C790 VN.n15 VSUBS 0.030677f
C791 VN.n16 VSUBS 0.057461f
C792 VN.n17 VSUBS 0.054057f
C793 VN.n18 VSUBS 0.918119f
C794 VN.n19 VSUBS 0.094149f
C795 VN.n20 VSUBS 0.057721f
C796 VN.t2 VSUBS 2.15262f
C797 VN.n21 VSUBS 0.058509f
C798 VN.n22 VSUBS 0.030677f
C799 VN.n23 VSUBS 0.057461f
C800 VN.t4 VSUBS 2.59333f
C801 VN.n24 VSUBS 0.866039f
C802 VN.t5 VSUBS 2.15262f
C803 VN.n25 VSUBS 0.894275f
C804 VN.n26 VSUBS 0.043276f
C805 VN.n27 VSUBS 0.40351f
C806 VN.n28 VSUBS 0.030677f
C807 VN.n29 VSUBS 0.030677f
C808 VN.n30 VSUBS 0.057461f
C809 VN.n31 VSUBS 0.053002f
C810 VN.n32 VSUBS 0.035907f
C811 VN.n33 VSUBS 0.030677f
C812 VN.n34 VSUBS 0.030677f
C813 VN.n35 VSUBS 0.030677f
C814 VN.n36 VSUBS 0.057461f
C815 VN.n37 VSUBS 0.054057f
C816 VN.n38 VSUBS 0.918119f
C817 VN.n39 VSUBS 1.78605f
C818 VDD1.t5 VSUBS 1.56515f
C819 VDD1.t0 VSUBS 1.56384f
C820 VDD1.t2 VSUBS 0.166338f
C821 VDD1.t1 VSUBS 0.166338f
C822 VDD1.n0 VSUBS 1.16991f
C823 VDD1.n1 VSUBS 4.53911f
C824 VDD1.t4 VSUBS 0.166338f
C825 VDD1.t3 VSUBS 0.166338f
C826 VDD1.n2 VSUBS 1.1608f
C827 VDD1.n3 VSUBS 3.63923f
C828 VTAIL.t4 VSUBS 0.183897f
C829 VTAIL.t5 VSUBS 0.183897f
C830 VTAIL.n0 VSUBS 1.15585f
C831 VTAIL.n1 VSUBS 0.990314f
C832 VTAIL.t6 VSUBS 1.56535f
C833 VTAIL.n2 VSUBS 1.37381f
C834 VTAIL.t11 VSUBS 0.183897f
C835 VTAIL.t10 VSUBS 0.183897f
C836 VTAIL.n3 VSUBS 1.15585f
C837 VTAIL.n4 VSUBS 2.93577f
C838 VTAIL.t1 VSUBS 0.183897f
C839 VTAIL.t2 VSUBS 0.183897f
C840 VTAIL.n5 VSUBS 1.15586f
C841 VTAIL.n6 VSUBS 2.93575f
C842 VTAIL.t3 VSUBS 1.56536f
C843 VTAIL.n7 VSUBS 1.3738f
C844 VTAIL.t9 VSUBS 0.183897f
C845 VTAIL.t8 VSUBS 0.183897f
C846 VTAIL.n8 VSUBS 1.15586f
C847 VTAIL.n9 VSUBS 1.28176f
C848 VTAIL.t7 VSUBS 1.56535f
C849 VTAIL.n10 VSUBS 2.63066f
C850 VTAIL.t0 VSUBS 1.56535f
C851 VTAIL.n11 VSUBS 2.52498f
C852 VP.n0 VSUBS 0.065948f
C853 VP.t4 VSUBS 2.45945f
C854 VP.n1 VSUBS 0.066849f
C855 VP.n2 VSUBS 0.03505f
C856 VP.n3 VSUBS 0.065652f
C857 VP.n4 VSUBS 0.03505f
C858 VP.t3 VSUBS 2.45945f
C859 VP.n5 VSUBS 0.065652f
C860 VP.n6 VSUBS 0.03505f
C861 VP.n7 VSUBS 0.065652f
C862 VP.n8 VSUBS 0.065948f
C863 VP.t2 VSUBS 2.45945f
C864 VP.n9 VSUBS 0.066849f
C865 VP.n10 VSUBS 0.03505f
C866 VP.n11 VSUBS 0.065652f
C867 VP.t0 VSUBS 2.96298f
C868 VP.n12 VSUBS 0.989488f
C869 VP.t1 VSUBS 2.45945f
C870 VP.n13 VSUBS 1.02175f
C871 VP.n14 VSUBS 0.049445f
C872 VP.n15 VSUBS 0.461028f
C873 VP.n16 VSUBS 0.03505f
C874 VP.n17 VSUBS 0.03505f
C875 VP.n18 VSUBS 0.065652f
C876 VP.n19 VSUBS 0.060557f
C877 VP.n20 VSUBS 0.041025f
C878 VP.n21 VSUBS 0.03505f
C879 VP.n22 VSUBS 0.03505f
C880 VP.n23 VSUBS 0.03505f
C881 VP.n24 VSUBS 0.065652f
C882 VP.n25 VSUBS 0.061762f
C883 VP.n26 VSUBS 1.04899f
C884 VP.n27 VSUBS 2.03144f
C885 VP.n28 VSUBS 2.0566f
C886 VP.t5 VSUBS 2.45945f
C887 VP.n29 VSUBS 1.04899f
C888 VP.n30 VSUBS 0.061762f
C889 VP.n31 VSUBS 0.065948f
C890 VP.n32 VSUBS 0.03505f
C891 VP.n33 VSUBS 0.03505f
C892 VP.n34 VSUBS 0.066849f
C893 VP.n35 VSUBS 0.041025f
C894 VP.n36 VSUBS 0.060557f
C895 VP.n37 VSUBS 0.03505f
C896 VP.n38 VSUBS 0.03505f
C897 VP.n39 VSUBS 0.03505f
C898 VP.n40 VSUBS 0.065652f
C899 VP.n41 VSUBS 0.049445f
C900 VP.n42 VSUBS 0.894361f
C901 VP.n43 VSUBS 0.049445f
C902 VP.n44 VSUBS 0.03505f
C903 VP.n45 VSUBS 0.03505f
C904 VP.n46 VSUBS 0.03505f
C905 VP.n47 VSUBS 0.065652f
C906 VP.n48 VSUBS 0.060557f
C907 VP.n49 VSUBS 0.041026f
C908 VP.n50 VSUBS 0.03505f
C909 VP.n51 VSUBS 0.03505f
C910 VP.n52 VSUBS 0.03505f
C911 VP.n53 VSUBS 0.065652f
C912 VP.n54 VSUBS 0.061762f
C913 VP.n55 VSUBS 1.04899f
C914 VP.n56 VSUBS 0.107569f
.ends

