* NGSPICE file created from diff_pair_sample_0364.ext - technology: sky130A

.subckt diff_pair_sample_0364 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t12 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=2.97165 ps=18.34 w=18.01 l=0.98
X1 VTAIL.t1 VP.t0 VDD1.t7 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=7.0239 pd=36.8 as=2.97165 ps=18.34 w=18.01 l=0.98
X2 B.t11 B.t9 B.t10 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=7.0239 pd=36.8 as=0 ps=0 w=18.01 l=0.98
X3 VDD1.t6 VP.t1 VTAIL.t7 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=7.0239 ps=36.8 w=18.01 l=0.98
X4 VDD2.t6 VN.t1 VTAIL.t13 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=2.97165 ps=18.34 w=18.01 l=0.98
X5 VDD1.t5 VP.t2 VTAIL.t2 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=2.97165 ps=18.34 w=18.01 l=0.98
X6 VTAIL.t15 VN.t2 VDD2.t5 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=7.0239 pd=36.8 as=2.97165 ps=18.34 w=18.01 l=0.98
X7 VDD2.t4 VN.t3 VTAIL.t8 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=7.0239 ps=36.8 w=18.01 l=0.98
X8 B.t8 B.t6 B.t7 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=7.0239 pd=36.8 as=0 ps=0 w=18.01 l=0.98
X9 VDD1.t4 VP.t3 VTAIL.t4 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=2.97165 ps=18.34 w=18.01 l=0.98
X10 VTAIL.t10 VN.t4 VDD2.t3 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=7.0239 pd=36.8 as=2.97165 ps=18.34 w=18.01 l=0.98
X11 VTAIL.t6 VP.t4 VDD1.t3 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=7.0239 pd=36.8 as=2.97165 ps=18.34 w=18.01 l=0.98
X12 VTAIL.t0 VP.t5 VDD1.t2 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=2.97165 ps=18.34 w=18.01 l=0.98
X13 VDD1.t1 VP.t6 VTAIL.t3 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=7.0239 ps=36.8 w=18.01 l=0.98
X14 B.t5 B.t3 B.t4 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=7.0239 pd=36.8 as=0 ps=0 w=18.01 l=0.98
X15 VTAIL.t5 VP.t7 VDD1.t0 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=2.97165 ps=18.34 w=18.01 l=0.98
X16 VTAIL.t11 VN.t5 VDD2.t2 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=2.97165 ps=18.34 w=18.01 l=0.98
X17 VTAIL.t14 VN.t6 VDD2.t1 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=2.97165 ps=18.34 w=18.01 l=0.98
X18 VDD2.t0 VN.t7 VTAIL.t9 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=2.97165 pd=18.34 as=7.0239 ps=36.8 w=18.01 l=0.98
X19 B.t2 B.t0 B.t1 w_n2280_n4570# sky130_fd_pr__pfet_01v8 ad=7.0239 pd=36.8 as=0 ps=0 w=18.01 l=0.98
R0 VN.n2 VN.t2 498.265
R1 VN.n15 VN.t3 498.265
R2 VN.n11 VN.t7 483.231
R3 VN.n24 VN.t4 483.231
R4 VN.n3 VN.t0 442.899
R5 VN.n9 VN.t5 442.899
R6 VN.n16 VN.t6 442.899
R7 VN.n22 VN.t1 442.899
R8 VN.n23 VN.n13 161.3
R9 VN.n21 VN.n20 161.3
R10 VN.n19 VN.n14 161.3
R11 VN.n18 VN.n17 161.3
R12 VN.n10 VN.n0 161.3
R13 VN.n8 VN.n7 161.3
R14 VN.n6 VN.n1 161.3
R15 VN.n5 VN.n4 161.3
R16 VN.n25 VN.n24 80.6037
R17 VN.n12 VN.n11 80.6037
R18 VN.n11 VN.n10 55.2959
R19 VN.n24 VN.n23 55.2959
R20 VN VN.n25 48.34
R21 VN.n3 VN.n2 46.8653
R22 VN.n16 VN.n15 46.8653
R23 VN.n18 VN.n15 44.049
R24 VN.n5 VN.n2 44.049
R25 VN.n4 VN.n1 40.4934
R26 VN.n8 VN.n1 40.4934
R27 VN.n17 VN.n14 40.4934
R28 VN.n21 VN.n14 40.4934
R29 VN.n10 VN.n9 16.8827
R30 VN.n23 VN.n22 16.8827
R31 VN.n4 VN.n3 7.58527
R32 VN.n9 VN.n8 7.58527
R33 VN.n17 VN.n16 7.58527
R34 VN.n22 VN.n21 7.58527
R35 VN.n25 VN.n13 0.285035
R36 VN.n12 VN.n0 0.285035
R37 VN.n20 VN.n13 0.189894
R38 VN.n20 VN.n19 0.189894
R39 VN.n19 VN.n18 0.189894
R40 VN.n6 VN.n5 0.189894
R41 VN.n7 VN.n6 0.189894
R42 VN.n7 VN.n0 0.189894
R43 VN VN.n12 0.146778
R44 VTAIL.n11 VTAIL.t1 56.498
R45 VTAIL.n10 VTAIL.t8 56.498
R46 VTAIL.n7 VTAIL.t10 56.498
R47 VTAIL.n15 VTAIL.t9 56.4977
R48 VTAIL.n2 VTAIL.t15 56.4977
R49 VTAIL.n3 VTAIL.t3 56.4977
R50 VTAIL.n6 VTAIL.t6 56.4977
R51 VTAIL.n14 VTAIL.t7 56.4977
R52 VTAIL.n13 VTAIL.n12 54.6931
R53 VTAIL.n9 VTAIL.n8 54.6931
R54 VTAIL.n1 VTAIL.n0 54.6929
R55 VTAIL.n5 VTAIL.n4 54.6929
R56 VTAIL.n15 VTAIL.n14 29.0221
R57 VTAIL.n7 VTAIL.n6 29.0221
R58 VTAIL.n0 VTAIL.t12 1.80533
R59 VTAIL.n0 VTAIL.t11 1.80533
R60 VTAIL.n4 VTAIL.t4 1.80533
R61 VTAIL.n4 VTAIL.t5 1.80533
R62 VTAIL.n12 VTAIL.t2 1.80533
R63 VTAIL.n12 VTAIL.t0 1.80533
R64 VTAIL.n8 VTAIL.t13 1.80533
R65 VTAIL.n8 VTAIL.t14 1.80533
R66 VTAIL.n9 VTAIL.n7 1.12981
R67 VTAIL.n10 VTAIL.n9 1.12981
R68 VTAIL.n13 VTAIL.n11 1.12981
R69 VTAIL.n14 VTAIL.n13 1.12981
R70 VTAIL.n6 VTAIL.n5 1.12981
R71 VTAIL.n5 VTAIL.n3 1.12981
R72 VTAIL.n2 VTAIL.n1 1.12981
R73 VTAIL VTAIL.n15 1.07162
R74 VTAIL.n11 VTAIL.n10 0.470328
R75 VTAIL.n3 VTAIL.n2 0.470328
R76 VTAIL VTAIL.n1 0.0586897
R77 VDD2.n2 VDD2.n1 71.881
R78 VDD2.n2 VDD2.n0 71.881
R79 VDD2 VDD2.n5 71.8782
R80 VDD2.n4 VDD2.n3 71.3719
R81 VDD2.n4 VDD2.n2 44.3231
R82 VDD2.n5 VDD2.t1 1.80533
R83 VDD2.n5 VDD2.t4 1.80533
R84 VDD2.n3 VDD2.t3 1.80533
R85 VDD2.n3 VDD2.t6 1.80533
R86 VDD2.n1 VDD2.t2 1.80533
R87 VDD2.n1 VDD2.t0 1.80533
R88 VDD2.n0 VDD2.t5 1.80533
R89 VDD2.n0 VDD2.t7 1.80533
R90 VDD2 VDD2.n4 0.623345
R91 VP.n5 VP.t0 498.265
R92 VP.n17 VP.t4 483.231
R93 VP.n27 VP.t6 483.231
R94 VP.n14 VP.t1 483.231
R95 VP.n19 VP.t3 442.899
R96 VP.n25 VP.t7 442.899
R97 VP.n12 VP.t5 442.899
R98 VP.n6 VP.t2 442.899
R99 VP.n8 VP.n7 161.3
R100 VP.n9 VP.n4 161.3
R101 VP.n11 VP.n10 161.3
R102 VP.n13 VP.n3 161.3
R103 VP.n26 VP.n0 161.3
R104 VP.n24 VP.n23 161.3
R105 VP.n22 VP.n1 161.3
R106 VP.n21 VP.n20 161.3
R107 VP.n18 VP.n2 161.3
R108 VP.n15 VP.n14 80.6037
R109 VP.n28 VP.n27 80.6037
R110 VP.n17 VP.n16 80.6037
R111 VP.n18 VP.n17 55.2959
R112 VP.n27 VP.n26 55.2959
R113 VP.n14 VP.n13 55.2959
R114 VP.n16 VP.n15 48.0544
R115 VP.n6 VP.n5 46.8653
R116 VP.n8 VP.n5 44.049
R117 VP.n20 VP.n1 40.4934
R118 VP.n24 VP.n1 40.4934
R119 VP.n11 VP.n4 40.4934
R120 VP.n7 VP.n4 40.4934
R121 VP.n19 VP.n18 16.8827
R122 VP.n26 VP.n25 16.8827
R123 VP.n13 VP.n12 16.8827
R124 VP.n20 VP.n19 7.58527
R125 VP.n25 VP.n24 7.58527
R126 VP.n12 VP.n11 7.58527
R127 VP.n7 VP.n6 7.58527
R128 VP.n15 VP.n3 0.285035
R129 VP.n16 VP.n2 0.285035
R130 VP.n28 VP.n0 0.285035
R131 VP.n9 VP.n8 0.189894
R132 VP.n10 VP.n9 0.189894
R133 VP.n10 VP.n3 0.189894
R134 VP.n21 VP.n2 0.189894
R135 VP.n22 VP.n21 0.189894
R136 VP.n23 VP.n22 0.189894
R137 VP.n23 VP.n0 0.189894
R138 VP VP.n28 0.146778
R139 VDD1 VDD1.n0 71.9947
R140 VDD1.n3 VDD1.n2 71.881
R141 VDD1.n3 VDD1.n1 71.881
R142 VDD1.n5 VDD1.n4 71.3717
R143 VDD1.n5 VDD1.n3 44.9061
R144 VDD1.n4 VDD1.t2 1.80533
R145 VDD1.n4 VDD1.t6 1.80533
R146 VDD1.n0 VDD1.t7 1.80533
R147 VDD1.n0 VDD1.t5 1.80533
R148 VDD1.n2 VDD1.t0 1.80533
R149 VDD1.n2 VDD1.t1 1.80533
R150 VDD1.n1 VDD1.t3 1.80533
R151 VDD1.n1 VDD1.t4 1.80533
R152 VDD1 VDD1.n5 0.506965
R153 B.n317 B.t9 645.688
R154 B.n142 B.t0 645.688
R155 B.n52 B.t6 645.688
R156 B.n46 B.t3 645.688
R157 B.n425 B.n112 585
R158 B.n424 B.n423 585
R159 B.n422 B.n113 585
R160 B.n421 B.n420 585
R161 B.n419 B.n114 585
R162 B.n418 B.n417 585
R163 B.n416 B.n115 585
R164 B.n415 B.n414 585
R165 B.n413 B.n116 585
R166 B.n412 B.n411 585
R167 B.n410 B.n117 585
R168 B.n409 B.n408 585
R169 B.n407 B.n118 585
R170 B.n406 B.n405 585
R171 B.n404 B.n119 585
R172 B.n403 B.n402 585
R173 B.n401 B.n120 585
R174 B.n400 B.n399 585
R175 B.n398 B.n121 585
R176 B.n397 B.n396 585
R177 B.n395 B.n122 585
R178 B.n394 B.n393 585
R179 B.n392 B.n123 585
R180 B.n391 B.n390 585
R181 B.n389 B.n124 585
R182 B.n388 B.n387 585
R183 B.n386 B.n125 585
R184 B.n385 B.n384 585
R185 B.n383 B.n126 585
R186 B.n382 B.n381 585
R187 B.n380 B.n127 585
R188 B.n379 B.n378 585
R189 B.n377 B.n128 585
R190 B.n376 B.n375 585
R191 B.n374 B.n129 585
R192 B.n373 B.n372 585
R193 B.n371 B.n130 585
R194 B.n370 B.n369 585
R195 B.n368 B.n131 585
R196 B.n367 B.n366 585
R197 B.n365 B.n132 585
R198 B.n364 B.n363 585
R199 B.n362 B.n133 585
R200 B.n361 B.n360 585
R201 B.n359 B.n134 585
R202 B.n358 B.n357 585
R203 B.n356 B.n135 585
R204 B.n355 B.n354 585
R205 B.n353 B.n136 585
R206 B.n352 B.n351 585
R207 B.n350 B.n137 585
R208 B.n349 B.n348 585
R209 B.n347 B.n138 585
R210 B.n346 B.n345 585
R211 B.n344 B.n139 585
R212 B.n343 B.n342 585
R213 B.n341 B.n140 585
R214 B.n340 B.n339 585
R215 B.n338 B.n141 585
R216 B.n336 B.n335 585
R217 B.n334 B.n144 585
R218 B.n333 B.n332 585
R219 B.n331 B.n145 585
R220 B.n330 B.n329 585
R221 B.n328 B.n146 585
R222 B.n327 B.n326 585
R223 B.n325 B.n147 585
R224 B.n324 B.n323 585
R225 B.n322 B.n148 585
R226 B.n321 B.n320 585
R227 B.n316 B.n149 585
R228 B.n315 B.n314 585
R229 B.n313 B.n150 585
R230 B.n312 B.n311 585
R231 B.n310 B.n151 585
R232 B.n309 B.n308 585
R233 B.n307 B.n152 585
R234 B.n306 B.n305 585
R235 B.n304 B.n153 585
R236 B.n303 B.n302 585
R237 B.n301 B.n154 585
R238 B.n300 B.n299 585
R239 B.n298 B.n155 585
R240 B.n297 B.n296 585
R241 B.n295 B.n156 585
R242 B.n294 B.n293 585
R243 B.n292 B.n157 585
R244 B.n291 B.n290 585
R245 B.n289 B.n158 585
R246 B.n288 B.n287 585
R247 B.n286 B.n159 585
R248 B.n285 B.n284 585
R249 B.n283 B.n160 585
R250 B.n282 B.n281 585
R251 B.n280 B.n161 585
R252 B.n279 B.n278 585
R253 B.n277 B.n162 585
R254 B.n276 B.n275 585
R255 B.n274 B.n163 585
R256 B.n273 B.n272 585
R257 B.n271 B.n164 585
R258 B.n270 B.n269 585
R259 B.n268 B.n165 585
R260 B.n267 B.n266 585
R261 B.n265 B.n166 585
R262 B.n264 B.n263 585
R263 B.n262 B.n167 585
R264 B.n261 B.n260 585
R265 B.n259 B.n168 585
R266 B.n258 B.n257 585
R267 B.n256 B.n169 585
R268 B.n255 B.n254 585
R269 B.n253 B.n170 585
R270 B.n252 B.n251 585
R271 B.n250 B.n171 585
R272 B.n249 B.n248 585
R273 B.n247 B.n172 585
R274 B.n246 B.n245 585
R275 B.n244 B.n173 585
R276 B.n243 B.n242 585
R277 B.n241 B.n174 585
R278 B.n240 B.n239 585
R279 B.n238 B.n175 585
R280 B.n237 B.n236 585
R281 B.n235 B.n176 585
R282 B.n234 B.n233 585
R283 B.n232 B.n177 585
R284 B.n231 B.n230 585
R285 B.n427 B.n426 585
R286 B.n428 B.n111 585
R287 B.n430 B.n429 585
R288 B.n431 B.n110 585
R289 B.n433 B.n432 585
R290 B.n434 B.n109 585
R291 B.n436 B.n435 585
R292 B.n437 B.n108 585
R293 B.n439 B.n438 585
R294 B.n440 B.n107 585
R295 B.n442 B.n441 585
R296 B.n443 B.n106 585
R297 B.n445 B.n444 585
R298 B.n446 B.n105 585
R299 B.n448 B.n447 585
R300 B.n449 B.n104 585
R301 B.n451 B.n450 585
R302 B.n452 B.n103 585
R303 B.n454 B.n453 585
R304 B.n455 B.n102 585
R305 B.n457 B.n456 585
R306 B.n458 B.n101 585
R307 B.n460 B.n459 585
R308 B.n461 B.n100 585
R309 B.n463 B.n462 585
R310 B.n464 B.n99 585
R311 B.n466 B.n465 585
R312 B.n467 B.n98 585
R313 B.n469 B.n468 585
R314 B.n470 B.n97 585
R315 B.n472 B.n471 585
R316 B.n473 B.n96 585
R317 B.n475 B.n474 585
R318 B.n476 B.n95 585
R319 B.n478 B.n477 585
R320 B.n479 B.n94 585
R321 B.n481 B.n480 585
R322 B.n482 B.n93 585
R323 B.n484 B.n483 585
R324 B.n485 B.n92 585
R325 B.n487 B.n486 585
R326 B.n488 B.n91 585
R327 B.n490 B.n489 585
R328 B.n491 B.n90 585
R329 B.n493 B.n492 585
R330 B.n494 B.n89 585
R331 B.n496 B.n495 585
R332 B.n497 B.n88 585
R333 B.n499 B.n498 585
R334 B.n500 B.n87 585
R335 B.n502 B.n501 585
R336 B.n503 B.n86 585
R337 B.n505 B.n504 585
R338 B.n506 B.n85 585
R339 B.n508 B.n507 585
R340 B.n509 B.n84 585
R341 B.n703 B.n702 585
R342 B.n701 B.n16 585
R343 B.n700 B.n699 585
R344 B.n698 B.n17 585
R345 B.n697 B.n696 585
R346 B.n695 B.n18 585
R347 B.n694 B.n693 585
R348 B.n692 B.n19 585
R349 B.n691 B.n690 585
R350 B.n689 B.n20 585
R351 B.n688 B.n687 585
R352 B.n686 B.n21 585
R353 B.n685 B.n684 585
R354 B.n683 B.n22 585
R355 B.n682 B.n681 585
R356 B.n680 B.n23 585
R357 B.n679 B.n678 585
R358 B.n677 B.n24 585
R359 B.n676 B.n675 585
R360 B.n674 B.n25 585
R361 B.n673 B.n672 585
R362 B.n671 B.n26 585
R363 B.n670 B.n669 585
R364 B.n668 B.n27 585
R365 B.n667 B.n666 585
R366 B.n665 B.n28 585
R367 B.n664 B.n663 585
R368 B.n662 B.n29 585
R369 B.n661 B.n660 585
R370 B.n659 B.n30 585
R371 B.n658 B.n657 585
R372 B.n656 B.n31 585
R373 B.n655 B.n654 585
R374 B.n653 B.n32 585
R375 B.n652 B.n651 585
R376 B.n650 B.n33 585
R377 B.n649 B.n648 585
R378 B.n647 B.n34 585
R379 B.n646 B.n645 585
R380 B.n644 B.n35 585
R381 B.n643 B.n642 585
R382 B.n641 B.n36 585
R383 B.n640 B.n639 585
R384 B.n638 B.n37 585
R385 B.n637 B.n636 585
R386 B.n635 B.n38 585
R387 B.n634 B.n633 585
R388 B.n632 B.n39 585
R389 B.n631 B.n630 585
R390 B.n629 B.n40 585
R391 B.n628 B.n627 585
R392 B.n626 B.n41 585
R393 B.n625 B.n624 585
R394 B.n623 B.n42 585
R395 B.n622 B.n621 585
R396 B.n620 B.n43 585
R397 B.n619 B.n618 585
R398 B.n617 B.n44 585
R399 B.n616 B.n615 585
R400 B.n613 B.n45 585
R401 B.n612 B.n611 585
R402 B.n610 B.n48 585
R403 B.n609 B.n608 585
R404 B.n607 B.n49 585
R405 B.n606 B.n605 585
R406 B.n604 B.n50 585
R407 B.n603 B.n602 585
R408 B.n601 B.n51 585
R409 B.n600 B.n599 585
R410 B.n598 B.n597 585
R411 B.n596 B.n55 585
R412 B.n595 B.n594 585
R413 B.n593 B.n56 585
R414 B.n592 B.n591 585
R415 B.n590 B.n57 585
R416 B.n589 B.n588 585
R417 B.n587 B.n58 585
R418 B.n586 B.n585 585
R419 B.n584 B.n59 585
R420 B.n583 B.n582 585
R421 B.n581 B.n60 585
R422 B.n580 B.n579 585
R423 B.n578 B.n61 585
R424 B.n577 B.n576 585
R425 B.n575 B.n62 585
R426 B.n574 B.n573 585
R427 B.n572 B.n63 585
R428 B.n571 B.n570 585
R429 B.n569 B.n64 585
R430 B.n568 B.n567 585
R431 B.n566 B.n65 585
R432 B.n565 B.n564 585
R433 B.n563 B.n66 585
R434 B.n562 B.n561 585
R435 B.n560 B.n67 585
R436 B.n559 B.n558 585
R437 B.n557 B.n68 585
R438 B.n556 B.n555 585
R439 B.n554 B.n69 585
R440 B.n553 B.n552 585
R441 B.n551 B.n70 585
R442 B.n550 B.n549 585
R443 B.n548 B.n71 585
R444 B.n547 B.n546 585
R445 B.n545 B.n72 585
R446 B.n544 B.n543 585
R447 B.n542 B.n73 585
R448 B.n541 B.n540 585
R449 B.n539 B.n74 585
R450 B.n538 B.n537 585
R451 B.n536 B.n75 585
R452 B.n535 B.n534 585
R453 B.n533 B.n76 585
R454 B.n532 B.n531 585
R455 B.n530 B.n77 585
R456 B.n529 B.n528 585
R457 B.n527 B.n78 585
R458 B.n526 B.n525 585
R459 B.n524 B.n79 585
R460 B.n523 B.n522 585
R461 B.n521 B.n80 585
R462 B.n520 B.n519 585
R463 B.n518 B.n81 585
R464 B.n517 B.n516 585
R465 B.n515 B.n82 585
R466 B.n514 B.n513 585
R467 B.n512 B.n83 585
R468 B.n511 B.n510 585
R469 B.n704 B.n15 585
R470 B.n706 B.n705 585
R471 B.n707 B.n14 585
R472 B.n709 B.n708 585
R473 B.n710 B.n13 585
R474 B.n712 B.n711 585
R475 B.n713 B.n12 585
R476 B.n715 B.n714 585
R477 B.n716 B.n11 585
R478 B.n718 B.n717 585
R479 B.n719 B.n10 585
R480 B.n721 B.n720 585
R481 B.n722 B.n9 585
R482 B.n724 B.n723 585
R483 B.n725 B.n8 585
R484 B.n727 B.n726 585
R485 B.n728 B.n7 585
R486 B.n730 B.n729 585
R487 B.n731 B.n6 585
R488 B.n733 B.n732 585
R489 B.n734 B.n5 585
R490 B.n736 B.n735 585
R491 B.n737 B.n4 585
R492 B.n739 B.n738 585
R493 B.n740 B.n3 585
R494 B.n742 B.n741 585
R495 B.n743 B.n0 585
R496 B.n2 B.n1 585
R497 B.n192 B.n191 585
R498 B.n193 B.n190 585
R499 B.n195 B.n194 585
R500 B.n196 B.n189 585
R501 B.n198 B.n197 585
R502 B.n199 B.n188 585
R503 B.n201 B.n200 585
R504 B.n202 B.n187 585
R505 B.n204 B.n203 585
R506 B.n205 B.n186 585
R507 B.n207 B.n206 585
R508 B.n208 B.n185 585
R509 B.n210 B.n209 585
R510 B.n211 B.n184 585
R511 B.n213 B.n212 585
R512 B.n214 B.n183 585
R513 B.n216 B.n215 585
R514 B.n217 B.n182 585
R515 B.n219 B.n218 585
R516 B.n220 B.n181 585
R517 B.n222 B.n221 585
R518 B.n223 B.n180 585
R519 B.n225 B.n224 585
R520 B.n226 B.n179 585
R521 B.n228 B.n227 585
R522 B.n229 B.n178 585
R523 B.n230 B.n229 492.5
R524 B.n426 B.n425 492.5
R525 B.n510 B.n509 492.5
R526 B.n702 B.n15 492.5
R527 B.n745 B.n744 256.663
R528 B.n744 B.n743 235.042
R529 B.n744 B.n2 235.042
R530 B.n230 B.n177 163.367
R531 B.n234 B.n177 163.367
R532 B.n235 B.n234 163.367
R533 B.n236 B.n235 163.367
R534 B.n236 B.n175 163.367
R535 B.n240 B.n175 163.367
R536 B.n241 B.n240 163.367
R537 B.n242 B.n241 163.367
R538 B.n242 B.n173 163.367
R539 B.n246 B.n173 163.367
R540 B.n247 B.n246 163.367
R541 B.n248 B.n247 163.367
R542 B.n248 B.n171 163.367
R543 B.n252 B.n171 163.367
R544 B.n253 B.n252 163.367
R545 B.n254 B.n253 163.367
R546 B.n254 B.n169 163.367
R547 B.n258 B.n169 163.367
R548 B.n259 B.n258 163.367
R549 B.n260 B.n259 163.367
R550 B.n260 B.n167 163.367
R551 B.n264 B.n167 163.367
R552 B.n265 B.n264 163.367
R553 B.n266 B.n265 163.367
R554 B.n266 B.n165 163.367
R555 B.n270 B.n165 163.367
R556 B.n271 B.n270 163.367
R557 B.n272 B.n271 163.367
R558 B.n272 B.n163 163.367
R559 B.n276 B.n163 163.367
R560 B.n277 B.n276 163.367
R561 B.n278 B.n277 163.367
R562 B.n278 B.n161 163.367
R563 B.n282 B.n161 163.367
R564 B.n283 B.n282 163.367
R565 B.n284 B.n283 163.367
R566 B.n284 B.n159 163.367
R567 B.n288 B.n159 163.367
R568 B.n289 B.n288 163.367
R569 B.n290 B.n289 163.367
R570 B.n290 B.n157 163.367
R571 B.n294 B.n157 163.367
R572 B.n295 B.n294 163.367
R573 B.n296 B.n295 163.367
R574 B.n296 B.n155 163.367
R575 B.n300 B.n155 163.367
R576 B.n301 B.n300 163.367
R577 B.n302 B.n301 163.367
R578 B.n302 B.n153 163.367
R579 B.n306 B.n153 163.367
R580 B.n307 B.n306 163.367
R581 B.n308 B.n307 163.367
R582 B.n308 B.n151 163.367
R583 B.n312 B.n151 163.367
R584 B.n313 B.n312 163.367
R585 B.n314 B.n313 163.367
R586 B.n314 B.n149 163.367
R587 B.n321 B.n149 163.367
R588 B.n322 B.n321 163.367
R589 B.n323 B.n322 163.367
R590 B.n323 B.n147 163.367
R591 B.n327 B.n147 163.367
R592 B.n328 B.n327 163.367
R593 B.n329 B.n328 163.367
R594 B.n329 B.n145 163.367
R595 B.n333 B.n145 163.367
R596 B.n334 B.n333 163.367
R597 B.n335 B.n334 163.367
R598 B.n335 B.n141 163.367
R599 B.n340 B.n141 163.367
R600 B.n341 B.n340 163.367
R601 B.n342 B.n341 163.367
R602 B.n342 B.n139 163.367
R603 B.n346 B.n139 163.367
R604 B.n347 B.n346 163.367
R605 B.n348 B.n347 163.367
R606 B.n348 B.n137 163.367
R607 B.n352 B.n137 163.367
R608 B.n353 B.n352 163.367
R609 B.n354 B.n353 163.367
R610 B.n354 B.n135 163.367
R611 B.n358 B.n135 163.367
R612 B.n359 B.n358 163.367
R613 B.n360 B.n359 163.367
R614 B.n360 B.n133 163.367
R615 B.n364 B.n133 163.367
R616 B.n365 B.n364 163.367
R617 B.n366 B.n365 163.367
R618 B.n366 B.n131 163.367
R619 B.n370 B.n131 163.367
R620 B.n371 B.n370 163.367
R621 B.n372 B.n371 163.367
R622 B.n372 B.n129 163.367
R623 B.n376 B.n129 163.367
R624 B.n377 B.n376 163.367
R625 B.n378 B.n377 163.367
R626 B.n378 B.n127 163.367
R627 B.n382 B.n127 163.367
R628 B.n383 B.n382 163.367
R629 B.n384 B.n383 163.367
R630 B.n384 B.n125 163.367
R631 B.n388 B.n125 163.367
R632 B.n389 B.n388 163.367
R633 B.n390 B.n389 163.367
R634 B.n390 B.n123 163.367
R635 B.n394 B.n123 163.367
R636 B.n395 B.n394 163.367
R637 B.n396 B.n395 163.367
R638 B.n396 B.n121 163.367
R639 B.n400 B.n121 163.367
R640 B.n401 B.n400 163.367
R641 B.n402 B.n401 163.367
R642 B.n402 B.n119 163.367
R643 B.n406 B.n119 163.367
R644 B.n407 B.n406 163.367
R645 B.n408 B.n407 163.367
R646 B.n408 B.n117 163.367
R647 B.n412 B.n117 163.367
R648 B.n413 B.n412 163.367
R649 B.n414 B.n413 163.367
R650 B.n414 B.n115 163.367
R651 B.n418 B.n115 163.367
R652 B.n419 B.n418 163.367
R653 B.n420 B.n419 163.367
R654 B.n420 B.n113 163.367
R655 B.n424 B.n113 163.367
R656 B.n425 B.n424 163.367
R657 B.n509 B.n508 163.367
R658 B.n508 B.n85 163.367
R659 B.n504 B.n85 163.367
R660 B.n504 B.n503 163.367
R661 B.n503 B.n502 163.367
R662 B.n502 B.n87 163.367
R663 B.n498 B.n87 163.367
R664 B.n498 B.n497 163.367
R665 B.n497 B.n496 163.367
R666 B.n496 B.n89 163.367
R667 B.n492 B.n89 163.367
R668 B.n492 B.n491 163.367
R669 B.n491 B.n490 163.367
R670 B.n490 B.n91 163.367
R671 B.n486 B.n91 163.367
R672 B.n486 B.n485 163.367
R673 B.n485 B.n484 163.367
R674 B.n484 B.n93 163.367
R675 B.n480 B.n93 163.367
R676 B.n480 B.n479 163.367
R677 B.n479 B.n478 163.367
R678 B.n478 B.n95 163.367
R679 B.n474 B.n95 163.367
R680 B.n474 B.n473 163.367
R681 B.n473 B.n472 163.367
R682 B.n472 B.n97 163.367
R683 B.n468 B.n97 163.367
R684 B.n468 B.n467 163.367
R685 B.n467 B.n466 163.367
R686 B.n466 B.n99 163.367
R687 B.n462 B.n99 163.367
R688 B.n462 B.n461 163.367
R689 B.n461 B.n460 163.367
R690 B.n460 B.n101 163.367
R691 B.n456 B.n101 163.367
R692 B.n456 B.n455 163.367
R693 B.n455 B.n454 163.367
R694 B.n454 B.n103 163.367
R695 B.n450 B.n103 163.367
R696 B.n450 B.n449 163.367
R697 B.n449 B.n448 163.367
R698 B.n448 B.n105 163.367
R699 B.n444 B.n105 163.367
R700 B.n444 B.n443 163.367
R701 B.n443 B.n442 163.367
R702 B.n442 B.n107 163.367
R703 B.n438 B.n107 163.367
R704 B.n438 B.n437 163.367
R705 B.n437 B.n436 163.367
R706 B.n436 B.n109 163.367
R707 B.n432 B.n109 163.367
R708 B.n432 B.n431 163.367
R709 B.n431 B.n430 163.367
R710 B.n430 B.n111 163.367
R711 B.n426 B.n111 163.367
R712 B.n702 B.n701 163.367
R713 B.n701 B.n700 163.367
R714 B.n700 B.n17 163.367
R715 B.n696 B.n17 163.367
R716 B.n696 B.n695 163.367
R717 B.n695 B.n694 163.367
R718 B.n694 B.n19 163.367
R719 B.n690 B.n19 163.367
R720 B.n690 B.n689 163.367
R721 B.n689 B.n688 163.367
R722 B.n688 B.n21 163.367
R723 B.n684 B.n21 163.367
R724 B.n684 B.n683 163.367
R725 B.n683 B.n682 163.367
R726 B.n682 B.n23 163.367
R727 B.n678 B.n23 163.367
R728 B.n678 B.n677 163.367
R729 B.n677 B.n676 163.367
R730 B.n676 B.n25 163.367
R731 B.n672 B.n25 163.367
R732 B.n672 B.n671 163.367
R733 B.n671 B.n670 163.367
R734 B.n670 B.n27 163.367
R735 B.n666 B.n27 163.367
R736 B.n666 B.n665 163.367
R737 B.n665 B.n664 163.367
R738 B.n664 B.n29 163.367
R739 B.n660 B.n29 163.367
R740 B.n660 B.n659 163.367
R741 B.n659 B.n658 163.367
R742 B.n658 B.n31 163.367
R743 B.n654 B.n31 163.367
R744 B.n654 B.n653 163.367
R745 B.n653 B.n652 163.367
R746 B.n652 B.n33 163.367
R747 B.n648 B.n33 163.367
R748 B.n648 B.n647 163.367
R749 B.n647 B.n646 163.367
R750 B.n646 B.n35 163.367
R751 B.n642 B.n35 163.367
R752 B.n642 B.n641 163.367
R753 B.n641 B.n640 163.367
R754 B.n640 B.n37 163.367
R755 B.n636 B.n37 163.367
R756 B.n636 B.n635 163.367
R757 B.n635 B.n634 163.367
R758 B.n634 B.n39 163.367
R759 B.n630 B.n39 163.367
R760 B.n630 B.n629 163.367
R761 B.n629 B.n628 163.367
R762 B.n628 B.n41 163.367
R763 B.n624 B.n41 163.367
R764 B.n624 B.n623 163.367
R765 B.n623 B.n622 163.367
R766 B.n622 B.n43 163.367
R767 B.n618 B.n43 163.367
R768 B.n618 B.n617 163.367
R769 B.n617 B.n616 163.367
R770 B.n616 B.n45 163.367
R771 B.n611 B.n45 163.367
R772 B.n611 B.n610 163.367
R773 B.n610 B.n609 163.367
R774 B.n609 B.n49 163.367
R775 B.n605 B.n49 163.367
R776 B.n605 B.n604 163.367
R777 B.n604 B.n603 163.367
R778 B.n603 B.n51 163.367
R779 B.n599 B.n51 163.367
R780 B.n599 B.n598 163.367
R781 B.n598 B.n55 163.367
R782 B.n594 B.n55 163.367
R783 B.n594 B.n593 163.367
R784 B.n593 B.n592 163.367
R785 B.n592 B.n57 163.367
R786 B.n588 B.n57 163.367
R787 B.n588 B.n587 163.367
R788 B.n587 B.n586 163.367
R789 B.n586 B.n59 163.367
R790 B.n582 B.n59 163.367
R791 B.n582 B.n581 163.367
R792 B.n581 B.n580 163.367
R793 B.n580 B.n61 163.367
R794 B.n576 B.n61 163.367
R795 B.n576 B.n575 163.367
R796 B.n575 B.n574 163.367
R797 B.n574 B.n63 163.367
R798 B.n570 B.n63 163.367
R799 B.n570 B.n569 163.367
R800 B.n569 B.n568 163.367
R801 B.n568 B.n65 163.367
R802 B.n564 B.n65 163.367
R803 B.n564 B.n563 163.367
R804 B.n563 B.n562 163.367
R805 B.n562 B.n67 163.367
R806 B.n558 B.n67 163.367
R807 B.n558 B.n557 163.367
R808 B.n557 B.n556 163.367
R809 B.n556 B.n69 163.367
R810 B.n552 B.n69 163.367
R811 B.n552 B.n551 163.367
R812 B.n551 B.n550 163.367
R813 B.n550 B.n71 163.367
R814 B.n546 B.n71 163.367
R815 B.n546 B.n545 163.367
R816 B.n545 B.n544 163.367
R817 B.n544 B.n73 163.367
R818 B.n540 B.n73 163.367
R819 B.n540 B.n539 163.367
R820 B.n539 B.n538 163.367
R821 B.n538 B.n75 163.367
R822 B.n534 B.n75 163.367
R823 B.n534 B.n533 163.367
R824 B.n533 B.n532 163.367
R825 B.n532 B.n77 163.367
R826 B.n528 B.n77 163.367
R827 B.n528 B.n527 163.367
R828 B.n527 B.n526 163.367
R829 B.n526 B.n79 163.367
R830 B.n522 B.n79 163.367
R831 B.n522 B.n521 163.367
R832 B.n521 B.n520 163.367
R833 B.n520 B.n81 163.367
R834 B.n516 B.n81 163.367
R835 B.n516 B.n515 163.367
R836 B.n515 B.n514 163.367
R837 B.n514 B.n83 163.367
R838 B.n510 B.n83 163.367
R839 B.n706 B.n15 163.367
R840 B.n707 B.n706 163.367
R841 B.n708 B.n707 163.367
R842 B.n708 B.n13 163.367
R843 B.n712 B.n13 163.367
R844 B.n713 B.n712 163.367
R845 B.n714 B.n713 163.367
R846 B.n714 B.n11 163.367
R847 B.n718 B.n11 163.367
R848 B.n719 B.n718 163.367
R849 B.n720 B.n719 163.367
R850 B.n720 B.n9 163.367
R851 B.n724 B.n9 163.367
R852 B.n725 B.n724 163.367
R853 B.n726 B.n725 163.367
R854 B.n726 B.n7 163.367
R855 B.n730 B.n7 163.367
R856 B.n731 B.n730 163.367
R857 B.n732 B.n731 163.367
R858 B.n732 B.n5 163.367
R859 B.n736 B.n5 163.367
R860 B.n737 B.n736 163.367
R861 B.n738 B.n737 163.367
R862 B.n738 B.n3 163.367
R863 B.n742 B.n3 163.367
R864 B.n743 B.n742 163.367
R865 B.n192 B.n2 163.367
R866 B.n193 B.n192 163.367
R867 B.n194 B.n193 163.367
R868 B.n194 B.n189 163.367
R869 B.n198 B.n189 163.367
R870 B.n199 B.n198 163.367
R871 B.n200 B.n199 163.367
R872 B.n200 B.n187 163.367
R873 B.n204 B.n187 163.367
R874 B.n205 B.n204 163.367
R875 B.n206 B.n205 163.367
R876 B.n206 B.n185 163.367
R877 B.n210 B.n185 163.367
R878 B.n211 B.n210 163.367
R879 B.n212 B.n211 163.367
R880 B.n212 B.n183 163.367
R881 B.n216 B.n183 163.367
R882 B.n217 B.n216 163.367
R883 B.n218 B.n217 163.367
R884 B.n218 B.n181 163.367
R885 B.n222 B.n181 163.367
R886 B.n223 B.n222 163.367
R887 B.n224 B.n223 163.367
R888 B.n224 B.n179 163.367
R889 B.n228 B.n179 163.367
R890 B.n229 B.n228 163.367
R891 B.n142 B.t1 138.008
R892 B.n52 B.t8 138.008
R893 B.n317 B.t10 137.986
R894 B.n46 B.t5 137.986
R895 B.n143 B.t2 112.603
R896 B.n53 B.t7 112.603
R897 B.n318 B.t11 112.579
R898 B.n47 B.t4 112.579
R899 B.n319 B.n318 59.5399
R900 B.n337 B.n143 59.5399
R901 B.n54 B.n53 59.5399
R902 B.n614 B.n47 59.5399
R903 B.n704 B.n703 32.0005
R904 B.n511 B.n84 32.0005
R905 B.n427 B.n112 32.0005
R906 B.n231 B.n178 32.0005
R907 B.n318 B.n317 25.4066
R908 B.n143 B.n142 25.4066
R909 B.n53 B.n52 25.4066
R910 B.n47 B.n46 25.4066
R911 B B.n745 18.0485
R912 B.n705 B.n704 10.6151
R913 B.n705 B.n14 10.6151
R914 B.n709 B.n14 10.6151
R915 B.n710 B.n709 10.6151
R916 B.n711 B.n710 10.6151
R917 B.n711 B.n12 10.6151
R918 B.n715 B.n12 10.6151
R919 B.n716 B.n715 10.6151
R920 B.n717 B.n716 10.6151
R921 B.n717 B.n10 10.6151
R922 B.n721 B.n10 10.6151
R923 B.n722 B.n721 10.6151
R924 B.n723 B.n722 10.6151
R925 B.n723 B.n8 10.6151
R926 B.n727 B.n8 10.6151
R927 B.n728 B.n727 10.6151
R928 B.n729 B.n728 10.6151
R929 B.n729 B.n6 10.6151
R930 B.n733 B.n6 10.6151
R931 B.n734 B.n733 10.6151
R932 B.n735 B.n734 10.6151
R933 B.n735 B.n4 10.6151
R934 B.n739 B.n4 10.6151
R935 B.n740 B.n739 10.6151
R936 B.n741 B.n740 10.6151
R937 B.n741 B.n0 10.6151
R938 B.n703 B.n16 10.6151
R939 B.n699 B.n16 10.6151
R940 B.n699 B.n698 10.6151
R941 B.n698 B.n697 10.6151
R942 B.n697 B.n18 10.6151
R943 B.n693 B.n18 10.6151
R944 B.n693 B.n692 10.6151
R945 B.n692 B.n691 10.6151
R946 B.n691 B.n20 10.6151
R947 B.n687 B.n20 10.6151
R948 B.n687 B.n686 10.6151
R949 B.n686 B.n685 10.6151
R950 B.n685 B.n22 10.6151
R951 B.n681 B.n22 10.6151
R952 B.n681 B.n680 10.6151
R953 B.n680 B.n679 10.6151
R954 B.n679 B.n24 10.6151
R955 B.n675 B.n24 10.6151
R956 B.n675 B.n674 10.6151
R957 B.n674 B.n673 10.6151
R958 B.n673 B.n26 10.6151
R959 B.n669 B.n26 10.6151
R960 B.n669 B.n668 10.6151
R961 B.n668 B.n667 10.6151
R962 B.n667 B.n28 10.6151
R963 B.n663 B.n28 10.6151
R964 B.n663 B.n662 10.6151
R965 B.n662 B.n661 10.6151
R966 B.n661 B.n30 10.6151
R967 B.n657 B.n30 10.6151
R968 B.n657 B.n656 10.6151
R969 B.n656 B.n655 10.6151
R970 B.n655 B.n32 10.6151
R971 B.n651 B.n32 10.6151
R972 B.n651 B.n650 10.6151
R973 B.n650 B.n649 10.6151
R974 B.n649 B.n34 10.6151
R975 B.n645 B.n34 10.6151
R976 B.n645 B.n644 10.6151
R977 B.n644 B.n643 10.6151
R978 B.n643 B.n36 10.6151
R979 B.n639 B.n36 10.6151
R980 B.n639 B.n638 10.6151
R981 B.n638 B.n637 10.6151
R982 B.n637 B.n38 10.6151
R983 B.n633 B.n38 10.6151
R984 B.n633 B.n632 10.6151
R985 B.n632 B.n631 10.6151
R986 B.n631 B.n40 10.6151
R987 B.n627 B.n40 10.6151
R988 B.n627 B.n626 10.6151
R989 B.n626 B.n625 10.6151
R990 B.n625 B.n42 10.6151
R991 B.n621 B.n42 10.6151
R992 B.n621 B.n620 10.6151
R993 B.n620 B.n619 10.6151
R994 B.n619 B.n44 10.6151
R995 B.n615 B.n44 10.6151
R996 B.n613 B.n612 10.6151
R997 B.n612 B.n48 10.6151
R998 B.n608 B.n48 10.6151
R999 B.n608 B.n607 10.6151
R1000 B.n607 B.n606 10.6151
R1001 B.n606 B.n50 10.6151
R1002 B.n602 B.n50 10.6151
R1003 B.n602 B.n601 10.6151
R1004 B.n601 B.n600 10.6151
R1005 B.n597 B.n596 10.6151
R1006 B.n596 B.n595 10.6151
R1007 B.n595 B.n56 10.6151
R1008 B.n591 B.n56 10.6151
R1009 B.n591 B.n590 10.6151
R1010 B.n590 B.n589 10.6151
R1011 B.n589 B.n58 10.6151
R1012 B.n585 B.n58 10.6151
R1013 B.n585 B.n584 10.6151
R1014 B.n584 B.n583 10.6151
R1015 B.n583 B.n60 10.6151
R1016 B.n579 B.n60 10.6151
R1017 B.n579 B.n578 10.6151
R1018 B.n578 B.n577 10.6151
R1019 B.n577 B.n62 10.6151
R1020 B.n573 B.n62 10.6151
R1021 B.n573 B.n572 10.6151
R1022 B.n572 B.n571 10.6151
R1023 B.n571 B.n64 10.6151
R1024 B.n567 B.n64 10.6151
R1025 B.n567 B.n566 10.6151
R1026 B.n566 B.n565 10.6151
R1027 B.n565 B.n66 10.6151
R1028 B.n561 B.n66 10.6151
R1029 B.n561 B.n560 10.6151
R1030 B.n560 B.n559 10.6151
R1031 B.n559 B.n68 10.6151
R1032 B.n555 B.n68 10.6151
R1033 B.n555 B.n554 10.6151
R1034 B.n554 B.n553 10.6151
R1035 B.n553 B.n70 10.6151
R1036 B.n549 B.n70 10.6151
R1037 B.n549 B.n548 10.6151
R1038 B.n548 B.n547 10.6151
R1039 B.n547 B.n72 10.6151
R1040 B.n543 B.n72 10.6151
R1041 B.n543 B.n542 10.6151
R1042 B.n542 B.n541 10.6151
R1043 B.n541 B.n74 10.6151
R1044 B.n537 B.n74 10.6151
R1045 B.n537 B.n536 10.6151
R1046 B.n536 B.n535 10.6151
R1047 B.n535 B.n76 10.6151
R1048 B.n531 B.n76 10.6151
R1049 B.n531 B.n530 10.6151
R1050 B.n530 B.n529 10.6151
R1051 B.n529 B.n78 10.6151
R1052 B.n525 B.n78 10.6151
R1053 B.n525 B.n524 10.6151
R1054 B.n524 B.n523 10.6151
R1055 B.n523 B.n80 10.6151
R1056 B.n519 B.n80 10.6151
R1057 B.n519 B.n518 10.6151
R1058 B.n518 B.n517 10.6151
R1059 B.n517 B.n82 10.6151
R1060 B.n513 B.n82 10.6151
R1061 B.n513 B.n512 10.6151
R1062 B.n512 B.n511 10.6151
R1063 B.n507 B.n84 10.6151
R1064 B.n507 B.n506 10.6151
R1065 B.n506 B.n505 10.6151
R1066 B.n505 B.n86 10.6151
R1067 B.n501 B.n86 10.6151
R1068 B.n501 B.n500 10.6151
R1069 B.n500 B.n499 10.6151
R1070 B.n499 B.n88 10.6151
R1071 B.n495 B.n88 10.6151
R1072 B.n495 B.n494 10.6151
R1073 B.n494 B.n493 10.6151
R1074 B.n493 B.n90 10.6151
R1075 B.n489 B.n90 10.6151
R1076 B.n489 B.n488 10.6151
R1077 B.n488 B.n487 10.6151
R1078 B.n487 B.n92 10.6151
R1079 B.n483 B.n92 10.6151
R1080 B.n483 B.n482 10.6151
R1081 B.n482 B.n481 10.6151
R1082 B.n481 B.n94 10.6151
R1083 B.n477 B.n94 10.6151
R1084 B.n477 B.n476 10.6151
R1085 B.n476 B.n475 10.6151
R1086 B.n475 B.n96 10.6151
R1087 B.n471 B.n96 10.6151
R1088 B.n471 B.n470 10.6151
R1089 B.n470 B.n469 10.6151
R1090 B.n469 B.n98 10.6151
R1091 B.n465 B.n98 10.6151
R1092 B.n465 B.n464 10.6151
R1093 B.n464 B.n463 10.6151
R1094 B.n463 B.n100 10.6151
R1095 B.n459 B.n100 10.6151
R1096 B.n459 B.n458 10.6151
R1097 B.n458 B.n457 10.6151
R1098 B.n457 B.n102 10.6151
R1099 B.n453 B.n102 10.6151
R1100 B.n453 B.n452 10.6151
R1101 B.n452 B.n451 10.6151
R1102 B.n451 B.n104 10.6151
R1103 B.n447 B.n104 10.6151
R1104 B.n447 B.n446 10.6151
R1105 B.n446 B.n445 10.6151
R1106 B.n445 B.n106 10.6151
R1107 B.n441 B.n106 10.6151
R1108 B.n441 B.n440 10.6151
R1109 B.n440 B.n439 10.6151
R1110 B.n439 B.n108 10.6151
R1111 B.n435 B.n108 10.6151
R1112 B.n435 B.n434 10.6151
R1113 B.n434 B.n433 10.6151
R1114 B.n433 B.n110 10.6151
R1115 B.n429 B.n110 10.6151
R1116 B.n429 B.n428 10.6151
R1117 B.n428 B.n427 10.6151
R1118 B.n191 B.n1 10.6151
R1119 B.n191 B.n190 10.6151
R1120 B.n195 B.n190 10.6151
R1121 B.n196 B.n195 10.6151
R1122 B.n197 B.n196 10.6151
R1123 B.n197 B.n188 10.6151
R1124 B.n201 B.n188 10.6151
R1125 B.n202 B.n201 10.6151
R1126 B.n203 B.n202 10.6151
R1127 B.n203 B.n186 10.6151
R1128 B.n207 B.n186 10.6151
R1129 B.n208 B.n207 10.6151
R1130 B.n209 B.n208 10.6151
R1131 B.n209 B.n184 10.6151
R1132 B.n213 B.n184 10.6151
R1133 B.n214 B.n213 10.6151
R1134 B.n215 B.n214 10.6151
R1135 B.n215 B.n182 10.6151
R1136 B.n219 B.n182 10.6151
R1137 B.n220 B.n219 10.6151
R1138 B.n221 B.n220 10.6151
R1139 B.n221 B.n180 10.6151
R1140 B.n225 B.n180 10.6151
R1141 B.n226 B.n225 10.6151
R1142 B.n227 B.n226 10.6151
R1143 B.n227 B.n178 10.6151
R1144 B.n232 B.n231 10.6151
R1145 B.n233 B.n232 10.6151
R1146 B.n233 B.n176 10.6151
R1147 B.n237 B.n176 10.6151
R1148 B.n238 B.n237 10.6151
R1149 B.n239 B.n238 10.6151
R1150 B.n239 B.n174 10.6151
R1151 B.n243 B.n174 10.6151
R1152 B.n244 B.n243 10.6151
R1153 B.n245 B.n244 10.6151
R1154 B.n245 B.n172 10.6151
R1155 B.n249 B.n172 10.6151
R1156 B.n250 B.n249 10.6151
R1157 B.n251 B.n250 10.6151
R1158 B.n251 B.n170 10.6151
R1159 B.n255 B.n170 10.6151
R1160 B.n256 B.n255 10.6151
R1161 B.n257 B.n256 10.6151
R1162 B.n257 B.n168 10.6151
R1163 B.n261 B.n168 10.6151
R1164 B.n262 B.n261 10.6151
R1165 B.n263 B.n262 10.6151
R1166 B.n263 B.n166 10.6151
R1167 B.n267 B.n166 10.6151
R1168 B.n268 B.n267 10.6151
R1169 B.n269 B.n268 10.6151
R1170 B.n269 B.n164 10.6151
R1171 B.n273 B.n164 10.6151
R1172 B.n274 B.n273 10.6151
R1173 B.n275 B.n274 10.6151
R1174 B.n275 B.n162 10.6151
R1175 B.n279 B.n162 10.6151
R1176 B.n280 B.n279 10.6151
R1177 B.n281 B.n280 10.6151
R1178 B.n281 B.n160 10.6151
R1179 B.n285 B.n160 10.6151
R1180 B.n286 B.n285 10.6151
R1181 B.n287 B.n286 10.6151
R1182 B.n287 B.n158 10.6151
R1183 B.n291 B.n158 10.6151
R1184 B.n292 B.n291 10.6151
R1185 B.n293 B.n292 10.6151
R1186 B.n293 B.n156 10.6151
R1187 B.n297 B.n156 10.6151
R1188 B.n298 B.n297 10.6151
R1189 B.n299 B.n298 10.6151
R1190 B.n299 B.n154 10.6151
R1191 B.n303 B.n154 10.6151
R1192 B.n304 B.n303 10.6151
R1193 B.n305 B.n304 10.6151
R1194 B.n305 B.n152 10.6151
R1195 B.n309 B.n152 10.6151
R1196 B.n310 B.n309 10.6151
R1197 B.n311 B.n310 10.6151
R1198 B.n311 B.n150 10.6151
R1199 B.n315 B.n150 10.6151
R1200 B.n316 B.n315 10.6151
R1201 B.n320 B.n316 10.6151
R1202 B.n324 B.n148 10.6151
R1203 B.n325 B.n324 10.6151
R1204 B.n326 B.n325 10.6151
R1205 B.n326 B.n146 10.6151
R1206 B.n330 B.n146 10.6151
R1207 B.n331 B.n330 10.6151
R1208 B.n332 B.n331 10.6151
R1209 B.n332 B.n144 10.6151
R1210 B.n336 B.n144 10.6151
R1211 B.n339 B.n338 10.6151
R1212 B.n339 B.n140 10.6151
R1213 B.n343 B.n140 10.6151
R1214 B.n344 B.n343 10.6151
R1215 B.n345 B.n344 10.6151
R1216 B.n345 B.n138 10.6151
R1217 B.n349 B.n138 10.6151
R1218 B.n350 B.n349 10.6151
R1219 B.n351 B.n350 10.6151
R1220 B.n351 B.n136 10.6151
R1221 B.n355 B.n136 10.6151
R1222 B.n356 B.n355 10.6151
R1223 B.n357 B.n356 10.6151
R1224 B.n357 B.n134 10.6151
R1225 B.n361 B.n134 10.6151
R1226 B.n362 B.n361 10.6151
R1227 B.n363 B.n362 10.6151
R1228 B.n363 B.n132 10.6151
R1229 B.n367 B.n132 10.6151
R1230 B.n368 B.n367 10.6151
R1231 B.n369 B.n368 10.6151
R1232 B.n369 B.n130 10.6151
R1233 B.n373 B.n130 10.6151
R1234 B.n374 B.n373 10.6151
R1235 B.n375 B.n374 10.6151
R1236 B.n375 B.n128 10.6151
R1237 B.n379 B.n128 10.6151
R1238 B.n380 B.n379 10.6151
R1239 B.n381 B.n380 10.6151
R1240 B.n381 B.n126 10.6151
R1241 B.n385 B.n126 10.6151
R1242 B.n386 B.n385 10.6151
R1243 B.n387 B.n386 10.6151
R1244 B.n387 B.n124 10.6151
R1245 B.n391 B.n124 10.6151
R1246 B.n392 B.n391 10.6151
R1247 B.n393 B.n392 10.6151
R1248 B.n393 B.n122 10.6151
R1249 B.n397 B.n122 10.6151
R1250 B.n398 B.n397 10.6151
R1251 B.n399 B.n398 10.6151
R1252 B.n399 B.n120 10.6151
R1253 B.n403 B.n120 10.6151
R1254 B.n404 B.n403 10.6151
R1255 B.n405 B.n404 10.6151
R1256 B.n405 B.n118 10.6151
R1257 B.n409 B.n118 10.6151
R1258 B.n410 B.n409 10.6151
R1259 B.n411 B.n410 10.6151
R1260 B.n411 B.n116 10.6151
R1261 B.n415 B.n116 10.6151
R1262 B.n416 B.n415 10.6151
R1263 B.n417 B.n416 10.6151
R1264 B.n417 B.n114 10.6151
R1265 B.n421 B.n114 10.6151
R1266 B.n422 B.n421 10.6151
R1267 B.n423 B.n422 10.6151
R1268 B.n423 B.n112 10.6151
R1269 B.n615 B.n614 9.36635
R1270 B.n597 B.n54 9.36635
R1271 B.n320 B.n319 9.36635
R1272 B.n338 B.n337 9.36635
R1273 B.n745 B.n0 8.11757
R1274 B.n745 B.n1 8.11757
R1275 B.n614 B.n613 1.24928
R1276 B.n600 B.n54 1.24928
R1277 B.n319 B.n148 1.24928
R1278 B.n337 B.n336 1.24928
C0 B VP 1.39741f
C1 VN VDD1 0.148851f
C2 VN VDD2 9.48975f
C3 w_n2280_n4570# VDD1 1.56901f
C4 VN VTAIL 9.14348f
C5 w_n2280_n4570# VDD2 1.61549f
C6 VN B 0.917864f
C7 w_n2280_n4570# VTAIL 5.6167f
C8 VDD1 VDD2 0.966157f
C9 VN VP 6.79365f
C10 VTAIL VDD1 13.2723f
C11 w_n2280_n4570# B 9.32079f
C12 w_n2280_n4570# VP 4.58949f
C13 VTAIL VDD2 13.3158f
C14 B VDD1 1.31749f
C15 VDD1 VP 9.68766f
C16 B VDD2 1.36281f
C17 VTAIL B 5.75072f
C18 VP VDD2 0.347337f
C19 VTAIL VP 9.15759f
C20 VN w_n2280_n4570# 4.29827f
C21 VDD2 VSUBS 1.536978f
C22 VDD1 VSUBS 1.894059f
C23 VTAIL VSUBS 1.288252f
C24 VN VSUBS 5.33069f
C25 VP VSUBS 2.172647f
C26 B VSUBS 3.706042f
C27 w_n2280_n4570# VSUBS 0.127416p
C28 B.n0 VSUBS 0.006513f
C29 B.n1 VSUBS 0.006513f
C30 B.n2 VSUBS 0.009632f
C31 B.n3 VSUBS 0.007381f
C32 B.n4 VSUBS 0.007381f
C33 B.n5 VSUBS 0.007381f
C34 B.n6 VSUBS 0.007381f
C35 B.n7 VSUBS 0.007381f
C36 B.n8 VSUBS 0.007381f
C37 B.n9 VSUBS 0.007381f
C38 B.n10 VSUBS 0.007381f
C39 B.n11 VSUBS 0.007381f
C40 B.n12 VSUBS 0.007381f
C41 B.n13 VSUBS 0.007381f
C42 B.n14 VSUBS 0.007381f
C43 B.n15 VSUBS 0.016771f
C44 B.n16 VSUBS 0.007381f
C45 B.n17 VSUBS 0.007381f
C46 B.n18 VSUBS 0.007381f
C47 B.n19 VSUBS 0.007381f
C48 B.n20 VSUBS 0.007381f
C49 B.n21 VSUBS 0.007381f
C50 B.n22 VSUBS 0.007381f
C51 B.n23 VSUBS 0.007381f
C52 B.n24 VSUBS 0.007381f
C53 B.n25 VSUBS 0.007381f
C54 B.n26 VSUBS 0.007381f
C55 B.n27 VSUBS 0.007381f
C56 B.n28 VSUBS 0.007381f
C57 B.n29 VSUBS 0.007381f
C58 B.n30 VSUBS 0.007381f
C59 B.n31 VSUBS 0.007381f
C60 B.n32 VSUBS 0.007381f
C61 B.n33 VSUBS 0.007381f
C62 B.n34 VSUBS 0.007381f
C63 B.n35 VSUBS 0.007381f
C64 B.n36 VSUBS 0.007381f
C65 B.n37 VSUBS 0.007381f
C66 B.n38 VSUBS 0.007381f
C67 B.n39 VSUBS 0.007381f
C68 B.n40 VSUBS 0.007381f
C69 B.n41 VSUBS 0.007381f
C70 B.n42 VSUBS 0.007381f
C71 B.n43 VSUBS 0.007381f
C72 B.n44 VSUBS 0.007381f
C73 B.n45 VSUBS 0.007381f
C74 B.t4 VSUBS 0.641178f
C75 B.t5 VSUBS 0.651933f
C76 B.t3 VSUBS 0.766711f
C77 B.n46 VSUBS 0.232721f
C78 B.n47 VSUBS 0.068941f
C79 B.n48 VSUBS 0.007381f
C80 B.n49 VSUBS 0.007381f
C81 B.n50 VSUBS 0.007381f
C82 B.n51 VSUBS 0.007381f
C83 B.t7 VSUBS 0.641155f
C84 B.t8 VSUBS 0.651912f
C85 B.t6 VSUBS 0.766711f
C86 B.n52 VSUBS 0.232741f
C87 B.n53 VSUBS 0.068964f
C88 B.n54 VSUBS 0.017102f
C89 B.n55 VSUBS 0.007381f
C90 B.n56 VSUBS 0.007381f
C91 B.n57 VSUBS 0.007381f
C92 B.n58 VSUBS 0.007381f
C93 B.n59 VSUBS 0.007381f
C94 B.n60 VSUBS 0.007381f
C95 B.n61 VSUBS 0.007381f
C96 B.n62 VSUBS 0.007381f
C97 B.n63 VSUBS 0.007381f
C98 B.n64 VSUBS 0.007381f
C99 B.n65 VSUBS 0.007381f
C100 B.n66 VSUBS 0.007381f
C101 B.n67 VSUBS 0.007381f
C102 B.n68 VSUBS 0.007381f
C103 B.n69 VSUBS 0.007381f
C104 B.n70 VSUBS 0.007381f
C105 B.n71 VSUBS 0.007381f
C106 B.n72 VSUBS 0.007381f
C107 B.n73 VSUBS 0.007381f
C108 B.n74 VSUBS 0.007381f
C109 B.n75 VSUBS 0.007381f
C110 B.n76 VSUBS 0.007381f
C111 B.n77 VSUBS 0.007381f
C112 B.n78 VSUBS 0.007381f
C113 B.n79 VSUBS 0.007381f
C114 B.n80 VSUBS 0.007381f
C115 B.n81 VSUBS 0.007381f
C116 B.n82 VSUBS 0.007381f
C117 B.n83 VSUBS 0.007381f
C118 B.n84 VSUBS 0.016771f
C119 B.n85 VSUBS 0.007381f
C120 B.n86 VSUBS 0.007381f
C121 B.n87 VSUBS 0.007381f
C122 B.n88 VSUBS 0.007381f
C123 B.n89 VSUBS 0.007381f
C124 B.n90 VSUBS 0.007381f
C125 B.n91 VSUBS 0.007381f
C126 B.n92 VSUBS 0.007381f
C127 B.n93 VSUBS 0.007381f
C128 B.n94 VSUBS 0.007381f
C129 B.n95 VSUBS 0.007381f
C130 B.n96 VSUBS 0.007381f
C131 B.n97 VSUBS 0.007381f
C132 B.n98 VSUBS 0.007381f
C133 B.n99 VSUBS 0.007381f
C134 B.n100 VSUBS 0.007381f
C135 B.n101 VSUBS 0.007381f
C136 B.n102 VSUBS 0.007381f
C137 B.n103 VSUBS 0.007381f
C138 B.n104 VSUBS 0.007381f
C139 B.n105 VSUBS 0.007381f
C140 B.n106 VSUBS 0.007381f
C141 B.n107 VSUBS 0.007381f
C142 B.n108 VSUBS 0.007381f
C143 B.n109 VSUBS 0.007381f
C144 B.n110 VSUBS 0.007381f
C145 B.n111 VSUBS 0.007381f
C146 B.n112 VSUBS 0.016423f
C147 B.n113 VSUBS 0.007381f
C148 B.n114 VSUBS 0.007381f
C149 B.n115 VSUBS 0.007381f
C150 B.n116 VSUBS 0.007381f
C151 B.n117 VSUBS 0.007381f
C152 B.n118 VSUBS 0.007381f
C153 B.n119 VSUBS 0.007381f
C154 B.n120 VSUBS 0.007381f
C155 B.n121 VSUBS 0.007381f
C156 B.n122 VSUBS 0.007381f
C157 B.n123 VSUBS 0.007381f
C158 B.n124 VSUBS 0.007381f
C159 B.n125 VSUBS 0.007381f
C160 B.n126 VSUBS 0.007381f
C161 B.n127 VSUBS 0.007381f
C162 B.n128 VSUBS 0.007381f
C163 B.n129 VSUBS 0.007381f
C164 B.n130 VSUBS 0.007381f
C165 B.n131 VSUBS 0.007381f
C166 B.n132 VSUBS 0.007381f
C167 B.n133 VSUBS 0.007381f
C168 B.n134 VSUBS 0.007381f
C169 B.n135 VSUBS 0.007381f
C170 B.n136 VSUBS 0.007381f
C171 B.n137 VSUBS 0.007381f
C172 B.n138 VSUBS 0.007381f
C173 B.n139 VSUBS 0.007381f
C174 B.n140 VSUBS 0.007381f
C175 B.n141 VSUBS 0.007381f
C176 B.t2 VSUBS 0.641155f
C177 B.t1 VSUBS 0.651912f
C178 B.t0 VSUBS 0.766711f
C179 B.n142 VSUBS 0.232741f
C180 B.n143 VSUBS 0.068964f
C181 B.n144 VSUBS 0.007381f
C182 B.n145 VSUBS 0.007381f
C183 B.n146 VSUBS 0.007381f
C184 B.n147 VSUBS 0.007381f
C185 B.n148 VSUBS 0.004125f
C186 B.n149 VSUBS 0.007381f
C187 B.n150 VSUBS 0.007381f
C188 B.n151 VSUBS 0.007381f
C189 B.n152 VSUBS 0.007381f
C190 B.n153 VSUBS 0.007381f
C191 B.n154 VSUBS 0.007381f
C192 B.n155 VSUBS 0.007381f
C193 B.n156 VSUBS 0.007381f
C194 B.n157 VSUBS 0.007381f
C195 B.n158 VSUBS 0.007381f
C196 B.n159 VSUBS 0.007381f
C197 B.n160 VSUBS 0.007381f
C198 B.n161 VSUBS 0.007381f
C199 B.n162 VSUBS 0.007381f
C200 B.n163 VSUBS 0.007381f
C201 B.n164 VSUBS 0.007381f
C202 B.n165 VSUBS 0.007381f
C203 B.n166 VSUBS 0.007381f
C204 B.n167 VSUBS 0.007381f
C205 B.n168 VSUBS 0.007381f
C206 B.n169 VSUBS 0.007381f
C207 B.n170 VSUBS 0.007381f
C208 B.n171 VSUBS 0.007381f
C209 B.n172 VSUBS 0.007381f
C210 B.n173 VSUBS 0.007381f
C211 B.n174 VSUBS 0.007381f
C212 B.n175 VSUBS 0.007381f
C213 B.n176 VSUBS 0.007381f
C214 B.n177 VSUBS 0.007381f
C215 B.n178 VSUBS 0.016771f
C216 B.n179 VSUBS 0.007381f
C217 B.n180 VSUBS 0.007381f
C218 B.n181 VSUBS 0.007381f
C219 B.n182 VSUBS 0.007381f
C220 B.n183 VSUBS 0.007381f
C221 B.n184 VSUBS 0.007381f
C222 B.n185 VSUBS 0.007381f
C223 B.n186 VSUBS 0.007381f
C224 B.n187 VSUBS 0.007381f
C225 B.n188 VSUBS 0.007381f
C226 B.n189 VSUBS 0.007381f
C227 B.n190 VSUBS 0.007381f
C228 B.n191 VSUBS 0.007381f
C229 B.n192 VSUBS 0.007381f
C230 B.n193 VSUBS 0.007381f
C231 B.n194 VSUBS 0.007381f
C232 B.n195 VSUBS 0.007381f
C233 B.n196 VSUBS 0.007381f
C234 B.n197 VSUBS 0.007381f
C235 B.n198 VSUBS 0.007381f
C236 B.n199 VSUBS 0.007381f
C237 B.n200 VSUBS 0.007381f
C238 B.n201 VSUBS 0.007381f
C239 B.n202 VSUBS 0.007381f
C240 B.n203 VSUBS 0.007381f
C241 B.n204 VSUBS 0.007381f
C242 B.n205 VSUBS 0.007381f
C243 B.n206 VSUBS 0.007381f
C244 B.n207 VSUBS 0.007381f
C245 B.n208 VSUBS 0.007381f
C246 B.n209 VSUBS 0.007381f
C247 B.n210 VSUBS 0.007381f
C248 B.n211 VSUBS 0.007381f
C249 B.n212 VSUBS 0.007381f
C250 B.n213 VSUBS 0.007381f
C251 B.n214 VSUBS 0.007381f
C252 B.n215 VSUBS 0.007381f
C253 B.n216 VSUBS 0.007381f
C254 B.n217 VSUBS 0.007381f
C255 B.n218 VSUBS 0.007381f
C256 B.n219 VSUBS 0.007381f
C257 B.n220 VSUBS 0.007381f
C258 B.n221 VSUBS 0.007381f
C259 B.n222 VSUBS 0.007381f
C260 B.n223 VSUBS 0.007381f
C261 B.n224 VSUBS 0.007381f
C262 B.n225 VSUBS 0.007381f
C263 B.n226 VSUBS 0.007381f
C264 B.n227 VSUBS 0.007381f
C265 B.n228 VSUBS 0.007381f
C266 B.n229 VSUBS 0.016771f
C267 B.n230 VSUBS 0.017313f
C268 B.n231 VSUBS 0.017313f
C269 B.n232 VSUBS 0.007381f
C270 B.n233 VSUBS 0.007381f
C271 B.n234 VSUBS 0.007381f
C272 B.n235 VSUBS 0.007381f
C273 B.n236 VSUBS 0.007381f
C274 B.n237 VSUBS 0.007381f
C275 B.n238 VSUBS 0.007381f
C276 B.n239 VSUBS 0.007381f
C277 B.n240 VSUBS 0.007381f
C278 B.n241 VSUBS 0.007381f
C279 B.n242 VSUBS 0.007381f
C280 B.n243 VSUBS 0.007381f
C281 B.n244 VSUBS 0.007381f
C282 B.n245 VSUBS 0.007381f
C283 B.n246 VSUBS 0.007381f
C284 B.n247 VSUBS 0.007381f
C285 B.n248 VSUBS 0.007381f
C286 B.n249 VSUBS 0.007381f
C287 B.n250 VSUBS 0.007381f
C288 B.n251 VSUBS 0.007381f
C289 B.n252 VSUBS 0.007381f
C290 B.n253 VSUBS 0.007381f
C291 B.n254 VSUBS 0.007381f
C292 B.n255 VSUBS 0.007381f
C293 B.n256 VSUBS 0.007381f
C294 B.n257 VSUBS 0.007381f
C295 B.n258 VSUBS 0.007381f
C296 B.n259 VSUBS 0.007381f
C297 B.n260 VSUBS 0.007381f
C298 B.n261 VSUBS 0.007381f
C299 B.n262 VSUBS 0.007381f
C300 B.n263 VSUBS 0.007381f
C301 B.n264 VSUBS 0.007381f
C302 B.n265 VSUBS 0.007381f
C303 B.n266 VSUBS 0.007381f
C304 B.n267 VSUBS 0.007381f
C305 B.n268 VSUBS 0.007381f
C306 B.n269 VSUBS 0.007381f
C307 B.n270 VSUBS 0.007381f
C308 B.n271 VSUBS 0.007381f
C309 B.n272 VSUBS 0.007381f
C310 B.n273 VSUBS 0.007381f
C311 B.n274 VSUBS 0.007381f
C312 B.n275 VSUBS 0.007381f
C313 B.n276 VSUBS 0.007381f
C314 B.n277 VSUBS 0.007381f
C315 B.n278 VSUBS 0.007381f
C316 B.n279 VSUBS 0.007381f
C317 B.n280 VSUBS 0.007381f
C318 B.n281 VSUBS 0.007381f
C319 B.n282 VSUBS 0.007381f
C320 B.n283 VSUBS 0.007381f
C321 B.n284 VSUBS 0.007381f
C322 B.n285 VSUBS 0.007381f
C323 B.n286 VSUBS 0.007381f
C324 B.n287 VSUBS 0.007381f
C325 B.n288 VSUBS 0.007381f
C326 B.n289 VSUBS 0.007381f
C327 B.n290 VSUBS 0.007381f
C328 B.n291 VSUBS 0.007381f
C329 B.n292 VSUBS 0.007381f
C330 B.n293 VSUBS 0.007381f
C331 B.n294 VSUBS 0.007381f
C332 B.n295 VSUBS 0.007381f
C333 B.n296 VSUBS 0.007381f
C334 B.n297 VSUBS 0.007381f
C335 B.n298 VSUBS 0.007381f
C336 B.n299 VSUBS 0.007381f
C337 B.n300 VSUBS 0.007381f
C338 B.n301 VSUBS 0.007381f
C339 B.n302 VSUBS 0.007381f
C340 B.n303 VSUBS 0.007381f
C341 B.n304 VSUBS 0.007381f
C342 B.n305 VSUBS 0.007381f
C343 B.n306 VSUBS 0.007381f
C344 B.n307 VSUBS 0.007381f
C345 B.n308 VSUBS 0.007381f
C346 B.n309 VSUBS 0.007381f
C347 B.n310 VSUBS 0.007381f
C348 B.n311 VSUBS 0.007381f
C349 B.n312 VSUBS 0.007381f
C350 B.n313 VSUBS 0.007381f
C351 B.n314 VSUBS 0.007381f
C352 B.n315 VSUBS 0.007381f
C353 B.n316 VSUBS 0.007381f
C354 B.t11 VSUBS 0.641178f
C355 B.t10 VSUBS 0.651933f
C356 B.t9 VSUBS 0.766711f
C357 B.n317 VSUBS 0.232721f
C358 B.n318 VSUBS 0.068941f
C359 B.n319 VSUBS 0.017102f
C360 B.n320 VSUBS 0.006947f
C361 B.n321 VSUBS 0.007381f
C362 B.n322 VSUBS 0.007381f
C363 B.n323 VSUBS 0.007381f
C364 B.n324 VSUBS 0.007381f
C365 B.n325 VSUBS 0.007381f
C366 B.n326 VSUBS 0.007381f
C367 B.n327 VSUBS 0.007381f
C368 B.n328 VSUBS 0.007381f
C369 B.n329 VSUBS 0.007381f
C370 B.n330 VSUBS 0.007381f
C371 B.n331 VSUBS 0.007381f
C372 B.n332 VSUBS 0.007381f
C373 B.n333 VSUBS 0.007381f
C374 B.n334 VSUBS 0.007381f
C375 B.n335 VSUBS 0.007381f
C376 B.n336 VSUBS 0.004125f
C377 B.n337 VSUBS 0.017102f
C378 B.n338 VSUBS 0.006947f
C379 B.n339 VSUBS 0.007381f
C380 B.n340 VSUBS 0.007381f
C381 B.n341 VSUBS 0.007381f
C382 B.n342 VSUBS 0.007381f
C383 B.n343 VSUBS 0.007381f
C384 B.n344 VSUBS 0.007381f
C385 B.n345 VSUBS 0.007381f
C386 B.n346 VSUBS 0.007381f
C387 B.n347 VSUBS 0.007381f
C388 B.n348 VSUBS 0.007381f
C389 B.n349 VSUBS 0.007381f
C390 B.n350 VSUBS 0.007381f
C391 B.n351 VSUBS 0.007381f
C392 B.n352 VSUBS 0.007381f
C393 B.n353 VSUBS 0.007381f
C394 B.n354 VSUBS 0.007381f
C395 B.n355 VSUBS 0.007381f
C396 B.n356 VSUBS 0.007381f
C397 B.n357 VSUBS 0.007381f
C398 B.n358 VSUBS 0.007381f
C399 B.n359 VSUBS 0.007381f
C400 B.n360 VSUBS 0.007381f
C401 B.n361 VSUBS 0.007381f
C402 B.n362 VSUBS 0.007381f
C403 B.n363 VSUBS 0.007381f
C404 B.n364 VSUBS 0.007381f
C405 B.n365 VSUBS 0.007381f
C406 B.n366 VSUBS 0.007381f
C407 B.n367 VSUBS 0.007381f
C408 B.n368 VSUBS 0.007381f
C409 B.n369 VSUBS 0.007381f
C410 B.n370 VSUBS 0.007381f
C411 B.n371 VSUBS 0.007381f
C412 B.n372 VSUBS 0.007381f
C413 B.n373 VSUBS 0.007381f
C414 B.n374 VSUBS 0.007381f
C415 B.n375 VSUBS 0.007381f
C416 B.n376 VSUBS 0.007381f
C417 B.n377 VSUBS 0.007381f
C418 B.n378 VSUBS 0.007381f
C419 B.n379 VSUBS 0.007381f
C420 B.n380 VSUBS 0.007381f
C421 B.n381 VSUBS 0.007381f
C422 B.n382 VSUBS 0.007381f
C423 B.n383 VSUBS 0.007381f
C424 B.n384 VSUBS 0.007381f
C425 B.n385 VSUBS 0.007381f
C426 B.n386 VSUBS 0.007381f
C427 B.n387 VSUBS 0.007381f
C428 B.n388 VSUBS 0.007381f
C429 B.n389 VSUBS 0.007381f
C430 B.n390 VSUBS 0.007381f
C431 B.n391 VSUBS 0.007381f
C432 B.n392 VSUBS 0.007381f
C433 B.n393 VSUBS 0.007381f
C434 B.n394 VSUBS 0.007381f
C435 B.n395 VSUBS 0.007381f
C436 B.n396 VSUBS 0.007381f
C437 B.n397 VSUBS 0.007381f
C438 B.n398 VSUBS 0.007381f
C439 B.n399 VSUBS 0.007381f
C440 B.n400 VSUBS 0.007381f
C441 B.n401 VSUBS 0.007381f
C442 B.n402 VSUBS 0.007381f
C443 B.n403 VSUBS 0.007381f
C444 B.n404 VSUBS 0.007381f
C445 B.n405 VSUBS 0.007381f
C446 B.n406 VSUBS 0.007381f
C447 B.n407 VSUBS 0.007381f
C448 B.n408 VSUBS 0.007381f
C449 B.n409 VSUBS 0.007381f
C450 B.n410 VSUBS 0.007381f
C451 B.n411 VSUBS 0.007381f
C452 B.n412 VSUBS 0.007381f
C453 B.n413 VSUBS 0.007381f
C454 B.n414 VSUBS 0.007381f
C455 B.n415 VSUBS 0.007381f
C456 B.n416 VSUBS 0.007381f
C457 B.n417 VSUBS 0.007381f
C458 B.n418 VSUBS 0.007381f
C459 B.n419 VSUBS 0.007381f
C460 B.n420 VSUBS 0.007381f
C461 B.n421 VSUBS 0.007381f
C462 B.n422 VSUBS 0.007381f
C463 B.n423 VSUBS 0.007381f
C464 B.n424 VSUBS 0.007381f
C465 B.n425 VSUBS 0.017313f
C466 B.n426 VSUBS 0.016771f
C467 B.n427 VSUBS 0.017661f
C468 B.n428 VSUBS 0.007381f
C469 B.n429 VSUBS 0.007381f
C470 B.n430 VSUBS 0.007381f
C471 B.n431 VSUBS 0.007381f
C472 B.n432 VSUBS 0.007381f
C473 B.n433 VSUBS 0.007381f
C474 B.n434 VSUBS 0.007381f
C475 B.n435 VSUBS 0.007381f
C476 B.n436 VSUBS 0.007381f
C477 B.n437 VSUBS 0.007381f
C478 B.n438 VSUBS 0.007381f
C479 B.n439 VSUBS 0.007381f
C480 B.n440 VSUBS 0.007381f
C481 B.n441 VSUBS 0.007381f
C482 B.n442 VSUBS 0.007381f
C483 B.n443 VSUBS 0.007381f
C484 B.n444 VSUBS 0.007381f
C485 B.n445 VSUBS 0.007381f
C486 B.n446 VSUBS 0.007381f
C487 B.n447 VSUBS 0.007381f
C488 B.n448 VSUBS 0.007381f
C489 B.n449 VSUBS 0.007381f
C490 B.n450 VSUBS 0.007381f
C491 B.n451 VSUBS 0.007381f
C492 B.n452 VSUBS 0.007381f
C493 B.n453 VSUBS 0.007381f
C494 B.n454 VSUBS 0.007381f
C495 B.n455 VSUBS 0.007381f
C496 B.n456 VSUBS 0.007381f
C497 B.n457 VSUBS 0.007381f
C498 B.n458 VSUBS 0.007381f
C499 B.n459 VSUBS 0.007381f
C500 B.n460 VSUBS 0.007381f
C501 B.n461 VSUBS 0.007381f
C502 B.n462 VSUBS 0.007381f
C503 B.n463 VSUBS 0.007381f
C504 B.n464 VSUBS 0.007381f
C505 B.n465 VSUBS 0.007381f
C506 B.n466 VSUBS 0.007381f
C507 B.n467 VSUBS 0.007381f
C508 B.n468 VSUBS 0.007381f
C509 B.n469 VSUBS 0.007381f
C510 B.n470 VSUBS 0.007381f
C511 B.n471 VSUBS 0.007381f
C512 B.n472 VSUBS 0.007381f
C513 B.n473 VSUBS 0.007381f
C514 B.n474 VSUBS 0.007381f
C515 B.n475 VSUBS 0.007381f
C516 B.n476 VSUBS 0.007381f
C517 B.n477 VSUBS 0.007381f
C518 B.n478 VSUBS 0.007381f
C519 B.n479 VSUBS 0.007381f
C520 B.n480 VSUBS 0.007381f
C521 B.n481 VSUBS 0.007381f
C522 B.n482 VSUBS 0.007381f
C523 B.n483 VSUBS 0.007381f
C524 B.n484 VSUBS 0.007381f
C525 B.n485 VSUBS 0.007381f
C526 B.n486 VSUBS 0.007381f
C527 B.n487 VSUBS 0.007381f
C528 B.n488 VSUBS 0.007381f
C529 B.n489 VSUBS 0.007381f
C530 B.n490 VSUBS 0.007381f
C531 B.n491 VSUBS 0.007381f
C532 B.n492 VSUBS 0.007381f
C533 B.n493 VSUBS 0.007381f
C534 B.n494 VSUBS 0.007381f
C535 B.n495 VSUBS 0.007381f
C536 B.n496 VSUBS 0.007381f
C537 B.n497 VSUBS 0.007381f
C538 B.n498 VSUBS 0.007381f
C539 B.n499 VSUBS 0.007381f
C540 B.n500 VSUBS 0.007381f
C541 B.n501 VSUBS 0.007381f
C542 B.n502 VSUBS 0.007381f
C543 B.n503 VSUBS 0.007381f
C544 B.n504 VSUBS 0.007381f
C545 B.n505 VSUBS 0.007381f
C546 B.n506 VSUBS 0.007381f
C547 B.n507 VSUBS 0.007381f
C548 B.n508 VSUBS 0.007381f
C549 B.n509 VSUBS 0.016771f
C550 B.n510 VSUBS 0.017313f
C551 B.n511 VSUBS 0.017313f
C552 B.n512 VSUBS 0.007381f
C553 B.n513 VSUBS 0.007381f
C554 B.n514 VSUBS 0.007381f
C555 B.n515 VSUBS 0.007381f
C556 B.n516 VSUBS 0.007381f
C557 B.n517 VSUBS 0.007381f
C558 B.n518 VSUBS 0.007381f
C559 B.n519 VSUBS 0.007381f
C560 B.n520 VSUBS 0.007381f
C561 B.n521 VSUBS 0.007381f
C562 B.n522 VSUBS 0.007381f
C563 B.n523 VSUBS 0.007381f
C564 B.n524 VSUBS 0.007381f
C565 B.n525 VSUBS 0.007381f
C566 B.n526 VSUBS 0.007381f
C567 B.n527 VSUBS 0.007381f
C568 B.n528 VSUBS 0.007381f
C569 B.n529 VSUBS 0.007381f
C570 B.n530 VSUBS 0.007381f
C571 B.n531 VSUBS 0.007381f
C572 B.n532 VSUBS 0.007381f
C573 B.n533 VSUBS 0.007381f
C574 B.n534 VSUBS 0.007381f
C575 B.n535 VSUBS 0.007381f
C576 B.n536 VSUBS 0.007381f
C577 B.n537 VSUBS 0.007381f
C578 B.n538 VSUBS 0.007381f
C579 B.n539 VSUBS 0.007381f
C580 B.n540 VSUBS 0.007381f
C581 B.n541 VSUBS 0.007381f
C582 B.n542 VSUBS 0.007381f
C583 B.n543 VSUBS 0.007381f
C584 B.n544 VSUBS 0.007381f
C585 B.n545 VSUBS 0.007381f
C586 B.n546 VSUBS 0.007381f
C587 B.n547 VSUBS 0.007381f
C588 B.n548 VSUBS 0.007381f
C589 B.n549 VSUBS 0.007381f
C590 B.n550 VSUBS 0.007381f
C591 B.n551 VSUBS 0.007381f
C592 B.n552 VSUBS 0.007381f
C593 B.n553 VSUBS 0.007381f
C594 B.n554 VSUBS 0.007381f
C595 B.n555 VSUBS 0.007381f
C596 B.n556 VSUBS 0.007381f
C597 B.n557 VSUBS 0.007381f
C598 B.n558 VSUBS 0.007381f
C599 B.n559 VSUBS 0.007381f
C600 B.n560 VSUBS 0.007381f
C601 B.n561 VSUBS 0.007381f
C602 B.n562 VSUBS 0.007381f
C603 B.n563 VSUBS 0.007381f
C604 B.n564 VSUBS 0.007381f
C605 B.n565 VSUBS 0.007381f
C606 B.n566 VSUBS 0.007381f
C607 B.n567 VSUBS 0.007381f
C608 B.n568 VSUBS 0.007381f
C609 B.n569 VSUBS 0.007381f
C610 B.n570 VSUBS 0.007381f
C611 B.n571 VSUBS 0.007381f
C612 B.n572 VSUBS 0.007381f
C613 B.n573 VSUBS 0.007381f
C614 B.n574 VSUBS 0.007381f
C615 B.n575 VSUBS 0.007381f
C616 B.n576 VSUBS 0.007381f
C617 B.n577 VSUBS 0.007381f
C618 B.n578 VSUBS 0.007381f
C619 B.n579 VSUBS 0.007381f
C620 B.n580 VSUBS 0.007381f
C621 B.n581 VSUBS 0.007381f
C622 B.n582 VSUBS 0.007381f
C623 B.n583 VSUBS 0.007381f
C624 B.n584 VSUBS 0.007381f
C625 B.n585 VSUBS 0.007381f
C626 B.n586 VSUBS 0.007381f
C627 B.n587 VSUBS 0.007381f
C628 B.n588 VSUBS 0.007381f
C629 B.n589 VSUBS 0.007381f
C630 B.n590 VSUBS 0.007381f
C631 B.n591 VSUBS 0.007381f
C632 B.n592 VSUBS 0.007381f
C633 B.n593 VSUBS 0.007381f
C634 B.n594 VSUBS 0.007381f
C635 B.n595 VSUBS 0.007381f
C636 B.n596 VSUBS 0.007381f
C637 B.n597 VSUBS 0.006947f
C638 B.n598 VSUBS 0.007381f
C639 B.n599 VSUBS 0.007381f
C640 B.n600 VSUBS 0.004125f
C641 B.n601 VSUBS 0.007381f
C642 B.n602 VSUBS 0.007381f
C643 B.n603 VSUBS 0.007381f
C644 B.n604 VSUBS 0.007381f
C645 B.n605 VSUBS 0.007381f
C646 B.n606 VSUBS 0.007381f
C647 B.n607 VSUBS 0.007381f
C648 B.n608 VSUBS 0.007381f
C649 B.n609 VSUBS 0.007381f
C650 B.n610 VSUBS 0.007381f
C651 B.n611 VSUBS 0.007381f
C652 B.n612 VSUBS 0.007381f
C653 B.n613 VSUBS 0.004125f
C654 B.n614 VSUBS 0.017102f
C655 B.n615 VSUBS 0.006947f
C656 B.n616 VSUBS 0.007381f
C657 B.n617 VSUBS 0.007381f
C658 B.n618 VSUBS 0.007381f
C659 B.n619 VSUBS 0.007381f
C660 B.n620 VSUBS 0.007381f
C661 B.n621 VSUBS 0.007381f
C662 B.n622 VSUBS 0.007381f
C663 B.n623 VSUBS 0.007381f
C664 B.n624 VSUBS 0.007381f
C665 B.n625 VSUBS 0.007381f
C666 B.n626 VSUBS 0.007381f
C667 B.n627 VSUBS 0.007381f
C668 B.n628 VSUBS 0.007381f
C669 B.n629 VSUBS 0.007381f
C670 B.n630 VSUBS 0.007381f
C671 B.n631 VSUBS 0.007381f
C672 B.n632 VSUBS 0.007381f
C673 B.n633 VSUBS 0.007381f
C674 B.n634 VSUBS 0.007381f
C675 B.n635 VSUBS 0.007381f
C676 B.n636 VSUBS 0.007381f
C677 B.n637 VSUBS 0.007381f
C678 B.n638 VSUBS 0.007381f
C679 B.n639 VSUBS 0.007381f
C680 B.n640 VSUBS 0.007381f
C681 B.n641 VSUBS 0.007381f
C682 B.n642 VSUBS 0.007381f
C683 B.n643 VSUBS 0.007381f
C684 B.n644 VSUBS 0.007381f
C685 B.n645 VSUBS 0.007381f
C686 B.n646 VSUBS 0.007381f
C687 B.n647 VSUBS 0.007381f
C688 B.n648 VSUBS 0.007381f
C689 B.n649 VSUBS 0.007381f
C690 B.n650 VSUBS 0.007381f
C691 B.n651 VSUBS 0.007381f
C692 B.n652 VSUBS 0.007381f
C693 B.n653 VSUBS 0.007381f
C694 B.n654 VSUBS 0.007381f
C695 B.n655 VSUBS 0.007381f
C696 B.n656 VSUBS 0.007381f
C697 B.n657 VSUBS 0.007381f
C698 B.n658 VSUBS 0.007381f
C699 B.n659 VSUBS 0.007381f
C700 B.n660 VSUBS 0.007381f
C701 B.n661 VSUBS 0.007381f
C702 B.n662 VSUBS 0.007381f
C703 B.n663 VSUBS 0.007381f
C704 B.n664 VSUBS 0.007381f
C705 B.n665 VSUBS 0.007381f
C706 B.n666 VSUBS 0.007381f
C707 B.n667 VSUBS 0.007381f
C708 B.n668 VSUBS 0.007381f
C709 B.n669 VSUBS 0.007381f
C710 B.n670 VSUBS 0.007381f
C711 B.n671 VSUBS 0.007381f
C712 B.n672 VSUBS 0.007381f
C713 B.n673 VSUBS 0.007381f
C714 B.n674 VSUBS 0.007381f
C715 B.n675 VSUBS 0.007381f
C716 B.n676 VSUBS 0.007381f
C717 B.n677 VSUBS 0.007381f
C718 B.n678 VSUBS 0.007381f
C719 B.n679 VSUBS 0.007381f
C720 B.n680 VSUBS 0.007381f
C721 B.n681 VSUBS 0.007381f
C722 B.n682 VSUBS 0.007381f
C723 B.n683 VSUBS 0.007381f
C724 B.n684 VSUBS 0.007381f
C725 B.n685 VSUBS 0.007381f
C726 B.n686 VSUBS 0.007381f
C727 B.n687 VSUBS 0.007381f
C728 B.n688 VSUBS 0.007381f
C729 B.n689 VSUBS 0.007381f
C730 B.n690 VSUBS 0.007381f
C731 B.n691 VSUBS 0.007381f
C732 B.n692 VSUBS 0.007381f
C733 B.n693 VSUBS 0.007381f
C734 B.n694 VSUBS 0.007381f
C735 B.n695 VSUBS 0.007381f
C736 B.n696 VSUBS 0.007381f
C737 B.n697 VSUBS 0.007381f
C738 B.n698 VSUBS 0.007381f
C739 B.n699 VSUBS 0.007381f
C740 B.n700 VSUBS 0.007381f
C741 B.n701 VSUBS 0.007381f
C742 B.n702 VSUBS 0.017313f
C743 B.n703 VSUBS 0.017313f
C744 B.n704 VSUBS 0.016771f
C745 B.n705 VSUBS 0.007381f
C746 B.n706 VSUBS 0.007381f
C747 B.n707 VSUBS 0.007381f
C748 B.n708 VSUBS 0.007381f
C749 B.n709 VSUBS 0.007381f
C750 B.n710 VSUBS 0.007381f
C751 B.n711 VSUBS 0.007381f
C752 B.n712 VSUBS 0.007381f
C753 B.n713 VSUBS 0.007381f
C754 B.n714 VSUBS 0.007381f
C755 B.n715 VSUBS 0.007381f
C756 B.n716 VSUBS 0.007381f
C757 B.n717 VSUBS 0.007381f
C758 B.n718 VSUBS 0.007381f
C759 B.n719 VSUBS 0.007381f
C760 B.n720 VSUBS 0.007381f
C761 B.n721 VSUBS 0.007381f
C762 B.n722 VSUBS 0.007381f
C763 B.n723 VSUBS 0.007381f
C764 B.n724 VSUBS 0.007381f
C765 B.n725 VSUBS 0.007381f
C766 B.n726 VSUBS 0.007381f
C767 B.n727 VSUBS 0.007381f
C768 B.n728 VSUBS 0.007381f
C769 B.n729 VSUBS 0.007381f
C770 B.n730 VSUBS 0.007381f
C771 B.n731 VSUBS 0.007381f
C772 B.n732 VSUBS 0.007381f
C773 B.n733 VSUBS 0.007381f
C774 B.n734 VSUBS 0.007381f
C775 B.n735 VSUBS 0.007381f
C776 B.n736 VSUBS 0.007381f
C777 B.n737 VSUBS 0.007381f
C778 B.n738 VSUBS 0.007381f
C779 B.n739 VSUBS 0.007381f
C780 B.n740 VSUBS 0.007381f
C781 B.n741 VSUBS 0.007381f
C782 B.n742 VSUBS 0.007381f
C783 B.n743 VSUBS 0.009632f
C784 B.n744 VSUBS 0.010261f
C785 B.n745 VSUBS 0.020404f
C786 VDD1.t7 VSUBS 0.373431f
C787 VDD1.t5 VSUBS 0.373431f
C788 VDD1.n0 VSUBS 3.11899f
C789 VDD1.t3 VSUBS 0.373431f
C790 VDD1.t4 VSUBS 0.373431f
C791 VDD1.n1 VSUBS 3.11789f
C792 VDD1.t0 VSUBS 0.373431f
C793 VDD1.t1 VSUBS 0.373431f
C794 VDD1.n2 VSUBS 3.11789f
C795 VDD1.n3 VSUBS 3.47823f
C796 VDD1.t2 VSUBS 0.373431f
C797 VDD1.t6 VSUBS 0.373431f
C798 VDD1.n4 VSUBS 3.11322f
C799 VDD1.n5 VSUBS 3.31111f
C800 VP.n0 VSUBS 0.060255f
C801 VP.t7 VSUBS 2.19222f
C802 VP.n1 VSUBS 0.036505f
C803 VP.n2 VSUBS 0.060255f
C804 VP.t3 VSUBS 2.19222f
C805 VP.n3 VSUBS 0.060255f
C806 VP.t1 VSUBS 2.26002f
C807 VP.t5 VSUBS 2.19222f
C808 VP.n4 VSUBS 0.036505f
C809 VP.t0 VSUBS 2.28579f
C810 VP.n5 VSUBS 0.850514f
C811 VP.t2 VSUBS 2.19222f
C812 VP.n6 VSUBS 0.824634f
C813 VP.n7 VSUBS 0.061076f
C814 VP.n8 VSUBS 0.191105f
C815 VP.n9 VSUBS 0.045156f
C816 VP.n10 VSUBS 0.045156f
C817 VP.n11 VSUBS 0.061076f
C818 VP.n12 VSUBS 0.786066f
C819 VP.n13 VSUBS 0.060284f
C820 VP.n14 VSUBS 0.853631f
C821 VP.n15 VSUBS 2.32741f
C822 VP.n16 VSUBS 2.36119f
C823 VP.t4 VSUBS 2.26002f
C824 VP.n17 VSUBS 0.853631f
C825 VP.n18 VSUBS 0.060284f
C826 VP.n19 VSUBS 0.786066f
C827 VP.n20 VSUBS 0.061076f
C828 VP.n21 VSUBS 0.045156f
C829 VP.n22 VSUBS 0.045156f
C830 VP.n23 VSUBS 0.045156f
C831 VP.n24 VSUBS 0.061076f
C832 VP.n25 VSUBS 0.786066f
C833 VP.n26 VSUBS 0.060284f
C834 VP.t6 VSUBS 2.26002f
C835 VP.n27 VSUBS 0.853631f
C836 VP.n28 VSUBS 0.042291f
C837 VDD2.t5 VSUBS 0.371751f
C838 VDD2.t7 VSUBS 0.371751f
C839 VDD2.n0 VSUBS 3.10385f
C840 VDD2.t2 VSUBS 0.371751f
C841 VDD2.t0 VSUBS 0.371751f
C842 VDD2.n1 VSUBS 3.10385f
C843 VDD2.n2 VSUBS 3.40742f
C844 VDD2.t3 VSUBS 0.371751f
C845 VDD2.t6 VSUBS 0.371751f
C846 VDD2.n3 VSUBS 3.09922f
C847 VDD2.n4 VSUBS 3.26467f
C848 VDD2.t1 VSUBS 0.371751f
C849 VDD2.t4 VSUBS 0.371751f
C850 VDD2.n5 VSUBS 3.10381f
C851 VTAIL.t12 VSUBS 0.334289f
C852 VTAIL.t11 VSUBS 0.334289f
C853 VTAIL.n0 VSUBS 2.64992f
C854 VTAIL.n1 VSUBS 0.648608f
C855 VTAIL.t15 VSUBS 3.45852f
C856 VTAIL.n2 VSUBS 0.782862f
C857 VTAIL.t3 VSUBS 3.45852f
C858 VTAIL.n3 VSUBS 0.782862f
C859 VTAIL.t4 VSUBS 0.334289f
C860 VTAIL.t5 VSUBS 0.334289f
C861 VTAIL.n4 VSUBS 2.64992f
C862 VTAIL.n5 VSUBS 0.729676f
C863 VTAIL.t6 VSUBS 3.45852f
C864 VTAIL.n6 VSUBS 2.32692f
C865 VTAIL.t10 VSUBS 3.45853f
C866 VTAIL.n7 VSUBS 2.32691f
C867 VTAIL.t13 VSUBS 0.334289f
C868 VTAIL.t14 VSUBS 0.334289f
C869 VTAIL.n8 VSUBS 2.64993f
C870 VTAIL.n9 VSUBS 0.729671f
C871 VTAIL.t8 VSUBS 3.45853f
C872 VTAIL.n10 VSUBS 0.782856f
C873 VTAIL.t1 VSUBS 3.45853f
C874 VTAIL.n11 VSUBS 0.782856f
C875 VTAIL.t2 VSUBS 0.334289f
C876 VTAIL.t0 VSUBS 0.334289f
C877 VTAIL.n12 VSUBS 2.64993f
C878 VTAIL.n13 VSUBS 0.729671f
C879 VTAIL.t7 VSUBS 3.45852f
C880 VTAIL.n14 VSUBS 2.32692f
C881 VTAIL.t9 VSUBS 3.45852f
C882 VTAIL.n15 VSUBS 2.32251f
C883 VN.n0 VSUBS 0.058939f
C884 VN.t5 VSUBS 2.14432f
C885 VN.n1 VSUBS 0.035707f
C886 VN.t2 VSUBS 2.23584f
C887 VN.n2 VSUBS 0.831929f
C888 VN.t0 VSUBS 2.14432f
C889 VN.n3 VSUBS 0.806615f
C890 VN.n4 VSUBS 0.059741f
C891 VN.n5 VSUBS 0.186929f
C892 VN.n6 VSUBS 0.044169f
C893 VN.n7 VSUBS 0.044169f
C894 VN.n8 VSUBS 0.059741f
C895 VN.n9 VSUBS 0.768889f
C896 VN.n10 VSUBS 0.058967f
C897 VN.t7 VSUBS 2.21063f
C898 VN.n11 VSUBS 0.834978f
C899 VN.n12 VSUBS 0.041366f
C900 VN.n13 VSUBS 0.058939f
C901 VN.t1 VSUBS 2.14432f
C902 VN.n14 VSUBS 0.035707f
C903 VN.t3 VSUBS 2.23584f
C904 VN.n15 VSUBS 0.831929f
C905 VN.t6 VSUBS 2.14432f
C906 VN.n16 VSUBS 0.806615f
C907 VN.n17 VSUBS 0.059741f
C908 VN.n18 VSUBS 0.186929f
C909 VN.n19 VSUBS 0.044169f
C910 VN.n20 VSUBS 0.044169f
C911 VN.n21 VSUBS 0.059741f
C912 VN.n22 VSUBS 0.768889f
C913 VN.n23 VSUBS 0.058967f
C914 VN.t4 VSUBS 2.21063f
C915 VN.n24 VSUBS 0.834978f
C916 VN.n25 VSUBS 2.30079f
.ends

