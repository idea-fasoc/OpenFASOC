* NGSPICE file created from diff_pair_sample_1119.ext - technology: sky130A

.subckt diff_pair_sample_1119 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=2.88585 ps=17.82 w=17.49 l=3.82
X1 VTAIL.t3 VN.t0 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=2.88585 ps=17.82 w=17.49 l=3.82
X2 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=0 ps=0 w=17.49 l=3.82
X3 VTAIL.t1 VN.t1 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=2.88585 ps=17.82 w=17.49 l=3.82
X4 VTAIL.t10 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=2.88585 ps=17.82 w=17.49 l=3.82
X5 VTAIL.t5 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=2.88585 ps=17.82 w=17.49 l=3.82
X6 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=0 ps=0 w=17.49 l=3.82
X7 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=0 ps=0 w=17.49 l=3.82
X8 VTAIL.t13 VP.t2 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=2.88585 ps=17.82 w=17.49 l=3.82
X9 VTAIL.t6 VN.t3 VDD2.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=2.88585 ps=17.82 w=17.49 l=3.82
X10 VTAIL.t11 VP.t3 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=2.88585 ps=17.82 w=17.49 l=3.82
X11 VDD2.t3 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=6.8211 ps=35.76 w=17.49 l=3.82
X12 VDD1.t3 VP.t4 VTAIL.t15 B.t0 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=2.88585 ps=17.82 w=17.49 l=3.82
X13 VDD2.t2 VN.t5 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=6.8211 ps=35.76 w=17.49 l=3.82
X14 VDD2.t1 VN.t6 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=2.88585 ps=17.82 w=17.49 l=3.82
X15 VDD2.t0 VN.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=2.88585 ps=17.82 w=17.49 l=3.82
X16 VDD1.t2 VP.t5 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=6.8211 ps=35.76 w=17.49 l=3.82
X17 VDD1.t1 VP.t6 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.88585 pd=17.82 as=6.8211 ps=35.76 w=17.49 l=3.82
X18 VTAIL.t8 VP.t7 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=2.88585 ps=17.82 w=17.49 l=3.82
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.8211 pd=35.76 as=0 ps=0 w=17.49 l=3.82
R0 VP.n23 VP.n22 161.3
R1 VP.n24 VP.n19 161.3
R2 VP.n26 VP.n25 161.3
R3 VP.n27 VP.n18 161.3
R4 VP.n29 VP.n28 161.3
R5 VP.n30 VP.n17 161.3
R6 VP.n32 VP.n31 161.3
R7 VP.n33 VP.n16 161.3
R8 VP.n36 VP.n35 161.3
R9 VP.n37 VP.n15 161.3
R10 VP.n39 VP.n38 161.3
R11 VP.n40 VP.n14 161.3
R12 VP.n42 VP.n41 161.3
R13 VP.n43 VP.n13 161.3
R14 VP.n45 VP.n44 161.3
R15 VP.n46 VP.n12 161.3
R16 VP.n88 VP.n0 161.3
R17 VP.n87 VP.n86 161.3
R18 VP.n85 VP.n1 161.3
R19 VP.n84 VP.n83 161.3
R20 VP.n82 VP.n2 161.3
R21 VP.n81 VP.n80 161.3
R22 VP.n79 VP.n3 161.3
R23 VP.n78 VP.n77 161.3
R24 VP.n75 VP.n4 161.3
R25 VP.n74 VP.n73 161.3
R26 VP.n72 VP.n5 161.3
R27 VP.n71 VP.n70 161.3
R28 VP.n69 VP.n6 161.3
R29 VP.n68 VP.n67 161.3
R30 VP.n66 VP.n7 161.3
R31 VP.n65 VP.n64 161.3
R32 VP.n62 VP.n8 161.3
R33 VP.n61 VP.n60 161.3
R34 VP.n59 VP.n9 161.3
R35 VP.n58 VP.n57 161.3
R36 VP.n56 VP.n10 161.3
R37 VP.n55 VP.n54 161.3
R38 VP.n53 VP.n11 161.3
R39 VP.n52 VP.n51 161.3
R40 VP.n20 VP.t7 142.482
R41 VP.n50 VP.t3 110.344
R42 VP.n63 VP.t0 110.344
R43 VP.n76 VP.t2 110.344
R44 VP.n89 VP.t6 110.344
R45 VP.n47 VP.t5 110.344
R46 VP.n34 VP.t1 110.344
R47 VP.n21 VP.t4 110.344
R48 VP.n49 VP.n48 61.0116
R49 VP.n21 VP.n20 59.1721
R50 VP.n50 VP.n49 58.9381
R51 VP.n90 VP.n89 58.9381
R52 VP.n48 VP.n47 58.9381
R53 VP.n70 VP.n69 56.5193
R54 VP.n28 VP.n27 56.5193
R55 VP.n57 VP.n56 50.2061
R56 VP.n83 VP.n82 50.2061
R57 VP.n41 VP.n40 50.2061
R58 VP.n56 VP.n55 30.7807
R59 VP.n83 VP.n1 30.7807
R60 VP.n41 VP.n13 30.7807
R61 VP.n51 VP.n11 24.4675
R62 VP.n55 VP.n11 24.4675
R63 VP.n57 VP.n9 24.4675
R64 VP.n61 VP.n9 24.4675
R65 VP.n62 VP.n61 24.4675
R66 VP.n64 VP.n7 24.4675
R67 VP.n68 VP.n7 24.4675
R68 VP.n69 VP.n68 24.4675
R69 VP.n70 VP.n5 24.4675
R70 VP.n74 VP.n5 24.4675
R71 VP.n75 VP.n74 24.4675
R72 VP.n77 VP.n3 24.4675
R73 VP.n81 VP.n3 24.4675
R74 VP.n82 VP.n81 24.4675
R75 VP.n87 VP.n1 24.4675
R76 VP.n88 VP.n87 24.4675
R77 VP.n45 VP.n13 24.4675
R78 VP.n46 VP.n45 24.4675
R79 VP.n28 VP.n17 24.4675
R80 VP.n32 VP.n17 24.4675
R81 VP.n33 VP.n32 24.4675
R82 VP.n35 VP.n15 24.4675
R83 VP.n39 VP.n15 24.4675
R84 VP.n40 VP.n39 24.4675
R85 VP.n22 VP.n19 24.4675
R86 VP.n26 VP.n19 24.4675
R87 VP.n27 VP.n26 24.4675
R88 VP.n51 VP.n50 23.2442
R89 VP.n89 VP.n88 23.2442
R90 VP.n47 VP.n46 23.2442
R91 VP.n64 VP.n63 15.9041
R92 VP.n76 VP.n75 15.9041
R93 VP.n34 VP.n33 15.9041
R94 VP.n22 VP.n21 15.9041
R95 VP.n63 VP.n62 8.56395
R96 VP.n77 VP.n76 8.56395
R97 VP.n35 VP.n34 8.56395
R98 VP.n23 VP.n20 2.57334
R99 VP.n48 VP.n12 0.417535
R100 VP.n52 VP.n49 0.417535
R101 VP.n90 VP.n0 0.417535
R102 VP VP.n90 0.394291
R103 VP.n24 VP.n23 0.189894
R104 VP.n25 VP.n24 0.189894
R105 VP.n25 VP.n18 0.189894
R106 VP.n29 VP.n18 0.189894
R107 VP.n30 VP.n29 0.189894
R108 VP.n31 VP.n30 0.189894
R109 VP.n31 VP.n16 0.189894
R110 VP.n36 VP.n16 0.189894
R111 VP.n37 VP.n36 0.189894
R112 VP.n38 VP.n37 0.189894
R113 VP.n38 VP.n14 0.189894
R114 VP.n42 VP.n14 0.189894
R115 VP.n43 VP.n42 0.189894
R116 VP.n44 VP.n43 0.189894
R117 VP.n44 VP.n12 0.189894
R118 VP.n53 VP.n52 0.189894
R119 VP.n54 VP.n53 0.189894
R120 VP.n54 VP.n10 0.189894
R121 VP.n58 VP.n10 0.189894
R122 VP.n59 VP.n58 0.189894
R123 VP.n60 VP.n59 0.189894
R124 VP.n60 VP.n8 0.189894
R125 VP.n65 VP.n8 0.189894
R126 VP.n66 VP.n65 0.189894
R127 VP.n67 VP.n66 0.189894
R128 VP.n67 VP.n6 0.189894
R129 VP.n71 VP.n6 0.189894
R130 VP.n72 VP.n71 0.189894
R131 VP.n73 VP.n72 0.189894
R132 VP.n73 VP.n4 0.189894
R133 VP.n78 VP.n4 0.189894
R134 VP.n79 VP.n78 0.189894
R135 VP.n80 VP.n79 0.189894
R136 VP.n80 VP.n2 0.189894
R137 VP.n84 VP.n2 0.189894
R138 VP.n85 VP.n84 0.189894
R139 VP.n86 VP.n85 0.189894
R140 VP.n86 VP.n0 0.189894
R141 VTAIL.n786 VTAIL.n694 289.615
R142 VTAIL.n94 VTAIL.n2 289.615
R143 VTAIL.n192 VTAIL.n100 289.615
R144 VTAIL.n292 VTAIL.n200 289.615
R145 VTAIL.n688 VTAIL.n596 289.615
R146 VTAIL.n588 VTAIL.n496 289.615
R147 VTAIL.n490 VTAIL.n398 289.615
R148 VTAIL.n390 VTAIL.n298 289.615
R149 VTAIL.n727 VTAIL.n726 185
R150 VTAIL.n729 VTAIL.n728 185
R151 VTAIL.n722 VTAIL.n721 185
R152 VTAIL.n735 VTAIL.n734 185
R153 VTAIL.n737 VTAIL.n736 185
R154 VTAIL.n718 VTAIL.n717 185
R155 VTAIL.n743 VTAIL.n742 185
R156 VTAIL.n745 VTAIL.n744 185
R157 VTAIL.n714 VTAIL.n713 185
R158 VTAIL.n751 VTAIL.n750 185
R159 VTAIL.n753 VTAIL.n752 185
R160 VTAIL.n710 VTAIL.n709 185
R161 VTAIL.n759 VTAIL.n758 185
R162 VTAIL.n761 VTAIL.n760 185
R163 VTAIL.n706 VTAIL.n705 185
R164 VTAIL.n768 VTAIL.n767 185
R165 VTAIL.n769 VTAIL.n704 185
R166 VTAIL.n771 VTAIL.n770 185
R167 VTAIL.n702 VTAIL.n701 185
R168 VTAIL.n777 VTAIL.n776 185
R169 VTAIL.n779 VTAIL.n778 185
R170 VTAIL.n698 VTAIL.n697 185
R171 VTAIL.n785 VTAIL.n784 185
R172 VTAIL.n787 VTAIL.n786 185
R173 VTAIL.n35 VTAIL.n34 185
R174 VTAIL.n37 VTAIL.n36 185
R175 VTAIL.n30 VTAIL.n29 185
R176 VTAIL.n43 VTAIL.n42 185
R177 VTAIL.n45 VTAIL.n44 185
R178 VTAIL.n26 VTAIL.n25 185
R179 VTAIL.n51 VTAIL.n50 185
R180 VTAIL.n53 VTAIL.n52 185
R181 VTAIL.n22 VTAIL.n21 185
R182 VTAIL.n59 VTAIL.n58 185
R183 VTAIL.n61 VTAIL.n60 185
R184 VTAIL.n18 VTAIL.n17 185
R185 VTAIL.n67 VTAIL.n66 185
R186 VTAIL.n69 VTAIL.n68 185
R187 VTAIL.n14 VTAIL.n13 185
R188 VTAIL.n76 VTAIL.n75 185
R189 VTAIL.n77 VTAIL.n12 185
R190 VTAIL.n79 VTAIL.n78 185
R191 VTAIL.n10 VTAIL.n9 185
R192 VTAIL.n85 VTAIL.n84 185
R193 VTAIL.n87 VTAIL.n86 185
R194 VTAIL.n6 VTAIL.n5 185
R195 VTAIL.n93 VTAIL.n92 185
R196 VTAIL.n95 VTAIL.n94 185
R197 VTAIL.n133 VTAIL.n132 185
R198 VTAIL.n135 VTAIL.n134 185
R199 VTAIL.n128 VTAIL.n127 185
R200 VTAIL.n141 VTAIL.n140 185
R201 VTAIL.n143 VTAIL.n142 185
R202 VTAIL.n124 VTAIL.n123 185
R203 VTAIL.n149 VTAIL.n148 185
R204 VTAIL.n151 VTAIL.n150 185
R205 VTAIL.n120 VTAIL.n119 185
R206 VTAIL.n157 VTAIL.n156 185
R207 VTAIL.n159 VTAIL.n158 185
R208 VTAIL.n116 VTAIL.n115 185
R209 VTAIL.n165 VTAIL.n164 185
R210 VTAIL.n167 VTAIL.n166 185
R211 VTAIL.n112 VTAIL.n111 185
R212 VTAIL.n174 VTAIL.n173 185
R213 VTAIL.n175 VTAIL.n110 185
R214 VTAIL.n177 VTAIL.n176 185
R215 VTAIL.n108 VTAIL.n107 185
R216 VTAIL.n183 VTAIL.n182 185
R217 VTAIL.n185 VTAIL.n184 185
R218 VTAIL.n104 VTAIL.n103 185
R219 VTAIL.n191 VTAIL.n190 185
R220 VTAIL.n193 VTAIL.n192 185
R221 VTAIL.n233 VTAIL.n232 185
R222 VTAIL.n235 VTAIL.n234 185
R223 VTAIL.n228 VTAIL.n227 185
R224 VTAIL.n241 VTAIL.n240 185
R225 VTAIL.n243 VTAIL.n242 185
R226 VTAIL.n224 VTAIL.n223 185
R227 VTAIL.n249 VTAIL.n248 185
R228 VTAIL.n251 VTAIL.n250 185
R229 VTAIL.n220 VTAIL.n219 185
R230 VTAIL.n257 VTAIL.n256 185
R231 VTAIL.n259 VTAIL.n258 185
R232 VTAIL.n216 VTAIL.n215 185
R233 VTAIL.n265 VTAIL.n264 185
R234 VTAIL.n267 VTAIL.n266 185
R235 VTAIL.n212 VTAIL.n211 185
R236 VTAIL.n274 VTAIL.n273 185
R237 VTAIL.n275 VTAIL.n210 185
R238 VTAIL.n277 VTAIL.n276 185
R239 VTAIL.n208 VTAIL.n207 185
R240 VTAIL.n283 VTAIL.n282 185
R241 VTAIL.n285 VTAIL.n284 185
R242 VTAIL.n204 VTAIL.n203 185
R243 VTAIL.n291 VTAIL.n290 185
R244 VTAIL.n293 VTAIL.n292 185
R245 VTAIL.n689 VTAIL.n688 185
R246 VTAIL.n687 VTAIL.n686 185
R247 VTAIL.n600 VTAIL.n599 185
R248 VTAIL.n681 VTAIL.n680 185
R249 VTAIL.n679 VTAIL.n678 185
R250 VTAIL.n604 VTAIL.n603 185
R251 VTAIL.n608 VTAIL.n606 185
R252 VTAIL.n673 VTAIL.n672 185
R253 VTAIL.n671 VTAIL.n670 185
R254 VTAIL.n610 VTAIL.n609 185
R255 VTAIL.n665 VTAIL.n664 185
R256 VTAIL.n663 VTAIL.n662 185
R257 VTAIL.n614 VTAIL.n613 185
R258 VTAIL.n657 VTAIL.n656 185
R259 VTAIL.n655 VTAIL.n654 185
R260 VTAIL.n618 VTAIL.n617 185
R261 VTAIL.n649 VTAIL.n648 185
R262 VTAIL.n647 VTAIL.n646 185
R263 VTAIL.n622 VTAIL.n621 185
R264 VTAIL.n641 VTAIL.n640 185
R265 VTAIL.n639 VTAIL.n638 185
R266 VTAIL.n626 VTAIL.n625 185
R267 VTAIL.n633 VTAIL.n632 185
R268 VTAIL.n631 VTAIL.n630 185
R269 VTAIL.n589 VTAIL.n588 185
R270 VTAIL.n587 VTAIL.n586 185
R271 VTAIL.n500 VTAIL.n499 185
R272 VTAIL.n581 VTAIL.n580 185
R273 VTAIL.n579 VTAIL.n578 185
R274 VTAIL.n504 VTAIL.n503 185
R275 VTAIL.n508 VTAIL.n506 185
R276 VTAIL.n573 VTAIL.n572 185
R277 VTAIL.n571 VTAIL.n570 185
R278 VTAIL.n510 VTAIL.n509 185
R279 VTAIL.n565 VTAIL.n564 185
R280 VTAIL.n563 VTAIL.n562 185
R281 VTAIL.n514 VTAIL.n513 185
R282 VTAIL.n557 VTAIL.n556 185
R283 VTAIL.n555 VTAIL.n554 185
R284 VTAIL.n518 VTAIL.n517 185
R285 VTAIL.n549 VTAIL.n548 185
R286 VTAIL.n547 VTAIL.n546 185
R287 VTAIL.n522 VTAIL.n521 185
R288 VTAIL.n541 VTAIL.n540 185
R289 VTAIL.n539 VTAIL.n538 185
R290 VTAIL.n526 VTAIL.n525 185
R291 VTAIL.n533 VTAIL.n532 185
R292 VTAIL.n531 VTAIL.n530 185
R293 VTAIL.n491 VTAIL.n490 185
R294 VTAIL.n489 VTAIL.n488 185
R295 VTAIL.n402 VTAIL.n401 185
R296 VTAIL.n483 VTAIL.n482 185
R297 VTAIL.n481 VTAIL.n480 185
R298 VTAIL.n406 VTAIL.n405 185
R299 VTAIL.n410 VTAIL.n408 185
R300 VTAIL.n475 VTAIL.n474 185
R301 VTAIL.n473 VTAIL.n472 185
R302 VTAIL.n412 VTAIL.n411 185
R303 VTAIL.n467 VTAIL.n466 185
R304 VTAIL.n465 VTAIL.n464 185
R305 VTAIL.n416 VTAIL.n415 185
R306 VTAIL.n459 VTAIL.n458 185
R307 VTAIL.n457 VTAIL.n456 185
R308 VTAIL.n420 VTAIL.n419 185
R309 VTAIL.n451 VTAIL.n450 185
R310 VTAIL.n449 VTAIL.n448 185
R311 VTAIL.n424 VTAIL.n423 185
R312 VTAIL.n443 VTAIL.n442 185
R313 VTAIL.n441 VTAIL.n440 185
R314 VTAIL.n428 VTAIL.n427 185
R315 VTAIL.n435 VTAIL.n434 185
R316 VTAIL.n433 VTAIL.n432 185
R317 VTAIL.n391 VTAIL.n390 185
R318 VTAIL.n389 VTAIL.n388 185
R319 VTAIL.n302 VTAIL.n301 185
R320 VTAIL.n383 VTAIL.n382 185
R321 VTAIL.n381 VTAIL.n380 185
R322 VTAIL.n306 VTAIL.n305 185
R323 VTAIL.n310 VTAIL.n308 185
R324 VTAIL.n375 VTAIL.n374 185
R325 VTAIL.n373 VTAIL.n372 185
R326 VTAIL.n312 VTAIL.n311 185
R327 VTAIL.n367 VTAIL.n366 185
R328 VTAIL.n365 VTAIL.n364 185
R329 VTAIL.n316 VTAIL.n315 185
R330 VTAIL.n359 VTAIL.n358 185
R331 VTAIL.n357 VTAIL.n356 185
R332 VTAIL.n320 VTAIL.n319 185
R333 VTAIL.n351 VTAIL.n350 185
R334 VTAIL.n349 VTAIL.n348 185
R335 VTAIL.n324 VTAIL.n323 185
R336 VTAIL.n343 VTAIL.n342 185
R337 VTAIL.n341 VTAIL.n340 185
R338 VTAIL.n328 VTAIL.n327 185
R339 VTAIL.n335 VTAIL.n334 185
R340 VTAIL.n333 VTAIL.n332 185
R341 VTAIL.n725 VTAIL.t4 147.659
R342 VTAIL.n33 VTAIL.t1 147.659
R343 VTAIL.n131 VTAIL.t14 147.659
R344 VTAIL.n231 VTAIL.t11 147.659
R345 VTAIL.n629 VTAIL.t9 147.659
R346 VTAIL.n529 VTAIL.t8 147.659
R347 VTAIL.n431 VTAIL.t7 147.659
R348 VTAIL.n331 VTAIL.t5 147.659
R349 VTAIL.n728 VTAIL.n727 104.615
R350 VTAIL.n728 VTAIL.n721 104.615
R351 VTAIL.n735 VTAIL.n721 104.615
R352 VTAIL.n736 VTAIL.n735 104.615
R353 VTAIL.n736 VTAIL.n717 104.615
R354 VTAIL.n743 VTAIL.n717 104.615
R355 VTAIL.n744 VTAIL.n743 104.615
R356 VTAIL.n744 VTAIL.n713 104.615
R357 VTAIL.n751 VTAIL.n713 104.615
R358 VTAIL.n752 VTAIL.n751 104.615
R359 VTAIL.n752 VTAIL.n709 104.615
R360 VTAIL.n759 VTAIL.n709 104.615
R361 VTAIL.n760 VTAIL.n759 104.615
R362 VTAIL.n760 VTAIL.n705 104.615
R363 VTAIL.n768 VTAIL.n705 104.615
R364 VTAIL.n769 VTAIL.n768 104.615
R365 VTAIL.n770 VTAIL.n769 104.615
R366 VTAIL.n770 VTAIL.n701 104.615
R367 VTAIL.n777 VTAIL.n701 104.615
R368 VTAIL.n778 VTAIL.n777 104.615
R369 VTAIL.n778 VTAIL.n697 104.615
R370 VTAIL.n785 VTAIL.n697 104.615
R371 VTAIL.n786 VTAIL.n785 104.615
R372 VTAIL.n36 VTAIL.n35 104.615
R373 VTAIL.n36 VTAIL.n29 104.615
R374 VTAIL.n43 VTAIL.n29 104.615
R375 VTAIL.n44 VTAIL.n43 104.615
R376 VTAIL.n44 VTAIL.n25 104.615
R377 VTAIL.n51 VTAIL.n25 104.615
R378 VTAIL.n52 VTAIL.n51 104.615
R379 VTAIL.n52 VTAIL.n21 104.615
R380 VTAIL.n59 VTAIL.n21 104.615
R381 VTAIL.n60 VTAIL.n59 104.615
R382 VTAIL.n60 VTAIL.n17 104.615
R383 VTAIL.n67 VTAIL.n17 104.615
R384 VTAIL.n68 VTAIL.n67 104.615
R385 VTAIL.n68 VTAIL.n13 104.615
R386 VTAIL.n76 VTAIL.n13 104.615
R387 VTAIL.n77 VTAIL.n76 104.615
R388 VTAIL.n78 VTAIL.n77 104.615
R389 VTAIL.n78 VTAIL.n9 104.615
R390 VTAIL.n85 VTAIL.n9 104.615
R391 VTAIL.n86 VTAIL.n85 104.615
R392 VTAIL.n86 VTAIL.n5 104.615
R393 VTAIL.n93 VTAIL.n5 104.615
R394 VTAIL.n94 VTAIL.n93 104.615
R395 VTAIL.n134 VTAIL.n133 104.615
R396 VTAIL.n134 VTAIL.n127 104.615
R397 VTAIL.n141 VTAIL.n127 104.615
R398 VTAIL.n142 VTAIL.n141 104.615
R399 VTAIL.n142 VTAIL.n123 104.615
R400 VTAIL.n149 VTAIL.n123 104.615
R401 VTAIL.n150 VTAIL.n149 104.615
R402 VTAIL.n150 VTAIL.n119 104.615
R403 VTAIL.n157 VTAIL.n119 104.615
R404 VTAIL.n158 VTAIL.n157 104.615
R405 VTAIL.n158 VTAIL.n115 104.615
R406 VTAIL.n165 VTAIL.n115 104.615
R407 VTAIL.n166 VTAIL.n165 104.615
R408 VTAIL.n166 VTAIL.n111 104.615
R409 VTAIL.n174 VTAIL.n111 104.615
R410 VTAIL.n175 VTAIL.n174 104.615
R411 VTAIL.n176 VTAIL.n175 104.615
R412 VTAIL.n176 VTAIL.n107 104.615
R413 VTAIL.n183 VTAIL.n107 104.615
R414 VTAIL.n184 VTAIL.n183 104.615
R415 VTAIL.n184 VTAIL.n103 104.615
R416 VTAIL.n191 VTAIL.n103 104.615
R417 VTAIL.n192 VTAIL.n191 104.615
R418 VTAIL.n234 VTAIL.n233 104.615
R419 VTAIL.n234 VTAIL.n227 104.615
R420 VTAIL.n241 VTAIL.n227 104.615
R421 VTAIL.n242 VTAIL.n241 104.615
R422 VTAIL.n242 VTAIL.n223 104.615
R423 VTAIL.n249 VTAIL.n223 104.615
R424 VTAIL.n250 VTAIL.n249 104.615
R425 VTAIL.n250 VTAIL.n219 104.615
R426 VTAIL.n257 VTAIL.n219 104.615
R427 VTAIL.n258 VTAIL.n257 104.615
R428 VTAIL.n258 VTAIL.n215 104.615
R429 VTAIL.n265 VTAIL.n215 104.615
R430 VTAIL.n266 VTAIL.n265 104.615
R431 VTAIL.n266 VTAIL.n211 104.615
R432 VTAIL.n274 VTAIL.n211 104.615
R433 VTAIL.n275 VTAIL.n274 104.615
R434 VTAIL.n276 VTAIL.n275 104.615
R435 VTAIL.n276 VTAIL.n207 104.615
R436 VTAIL.n283 VTAIL.n207 104.615
R437 VTAIL.n284 VTAIL.n283 104.615
R438 VTAIL.n284 VTAIL.n203 104.615
R439 VTAIL.n291 VTAIL.n203 104.615
R440 VTAIL.n292 VTAIL.n291 104.615
R441 VTAIL.n688 VTAIL.n687 104.615
R442 VTAIL.n687 VTAIL.n599 104.615
R443 VTAIL.n680 VTAIL.n599 104.615
R444 VTAIL.n680 VTAIL.n679 104.615
R445 VTAIL.n679 VTAIL.n603 104.615
R446 VTAIL.n608 VTAIL.n603 104.615
R447 VTAIL.n672 VTAIL.n608 104.615
R448 VTAIL.n672 VTAIL.n671 104.615
R449 VTAIL.n671 VTAIL.n609 104.615
R450 VTAIL.n664 VTAIL.n609 104.615
R451 VTAIL.n664 VTAIL.n663 104.615
R452 VTAIL.n663 VTAIL.n613 104.615
R453 VTAIL.n656 VTAIL.n613 104.615
R454 VTAIL.n656 VTAIL.n655 104.615
R455 VTAIL.n655 VTAIL.n617 104.615
R456 VTAIL.n648 VTAIL.n617 104.615
R457 VTAIL.n648 VTAIL.n647 104.615
R458 VTAIL.n647 VTAIL.n621 104.615
R459 VTAIL.n640 VTAIL.n621 104.615
R460 VTAIL.n640 VTAIL.n639 104.615
R461 VTAIL.n639 VTAIL.n625 104.615
R462 VTAIL.n632 VTAIL.n625 104.615
R463 VTAIL.n632 VTAIL.n631 104.615
R464 VTAIL.n588 VTAIL.n587 104.615
R465 VTAIL.n587 VTAIL.n499 104.615
R466 VTAIL.n580 VTAIL.n499 104.615
R467 VTAIL.n580 VTAIL.n579 104.615
R468 VTAIL.n579 VTAIL.n503 104.615
R469 VTAIL.n508 VTAIL.n503 104.615
R470 VTAIL.n572 VTAIL.n508 104.615
R471 VTAIL.n572 VTAIL.n571 104.615
R472 VTAIL.n571 VTAIL.n509 104.615
R473 VTAIL.n564 VTAIL.n509 104.615
R474 VTAIL.n564 VTAIL.n563 104.615
R475 VTAIL.n563 VTAIL.n513 104.615
R476 VTAIL.n556 VTAIL.n513 104.615
R477 VTAIL.n556 VTAIL.n555 104.615
R478 VTAIL.n555 VTAIL.n517 104.615
R479 VTAIL.n548 VTAIL.n517 104.615
R480 VTAIL.n548 VTAIL.n547 104.615
R481 VTAIL.n547 VTAIL.n521 104.615
R482 VTAIL.n540 VTAIL.n521 104.615
R483 VTAIL.n540 VTAIL.n539 104.615
R484 VTAIL.n539 VTAIL.n525 104.615
R485 VTAIL.n532 VTAIL.n525 104.615
R486 VTAIL.n532 VTAIL.n531 104.615
R487 VTAIL.n490 VTAIL.n489 104.615
R488 VTAIL.n489 VTAIL.n401 104.615
R489 VTAIL.n482 VTAIL.n401 104.615
R490 VTAIL.n482 VTAIL.n481 104.615
R491 VTAIL.n481 VTAIL.n405 104.615
R492 VTAIL.n410 VTAIL.n405 104.615
R493 VTAIL.n474 VTAIL.n410 104.615
R494 VTAIL.n474 VTAIL.n473 104.615
R495 VTAIL.n473 VTAIL.n411 104.615
R496 VTAIL.n466 VTAIL.n411 104.615
R497 VTAIL.n466 VTAIL.n465 104.615
R498 VTAIL.n465 VTAIL.n415 104.615
R499 VTAIL.n458 VTAIL.n415 104.615
R500 VTAIL.n458 VTAIL.n457 104.615
R501 VTAIL.n457 VTAIL.n419 104.615
R502 VTAIL.n450 VTAIL.n419 104.615
R503 VTAIL.n450 VTAIL.n449 104.615
R504 VTAIL.n449 VTAIL.n423 104.615
R505 VTAIL.n442 VTAIL.n423 104.615
R506 VTAIL.n442 VTAIL.n441 104.615
R507 VTAIL.n441 VTAIL.n427 104.615
R508 VTAIL.n434 VTAIL.n427 104.615
R509 VTAIL.n434 VTAIL.n433 104.615
R510 VTAIL.n390 VTAIL.n389 104.615
R511 VTAIL.n389 VTAIL.n301 104.615
R512 VTAIL.n382 VTAIL.n301 104.615
R513 VTAIL.n382 VTAIL.n381 104.615
R514 VTAIL.n381 VTAIL.n305 104.615
R515 VTAIL.n310 VTAIL.n305 104.615
R516 VTAIL.n374 VTAIL.n310 104.615
R517 VTAIL.n374 VTAIL.n373 104.615
R518 VTAIL.n373 VTAIL.n311 104.615
R519 VTAIL.n366 VTAIL.n311 104.615
R520 VTAIL.n366 VTAIL.n365 104.615
R521 VTAIL.n365 VTAIL.n315 104.615
R522 VTAIL.n358 VTAIL.n315 104.615
R523 VTAIL.n358 VTAIL.n357 104.615
R524 VTAIL.n357 VTAIL.n319 104.615
R525 VTAIL.n350 VTAIL.n319 104.615
R526 VTAIL.n350 VTAIL.n349 104.615
R527 VTAIL.n349 VTAIL.n323 104.615
R528 VTAIL.n342 VTAIL.n323 104.615
R529 VTAIL.n342 VTAIL.n341 104.615
R530 VTAIL.n341 VTAIL.n327 104.615
R531 VTAIL.n334 VTAIL.n327 104.615
R532 VTAIL.n334 VTAIL.n333 104.615
R533 VTAIL.n727 VTAIL.t4 52.3082
R534 VTAIL.n35 VTAIL.t1 52.3082
R535 VTAIL.n133 VTAIL.t14 52.3082
R536 VTAIL.n233 VTAIL.t11 52.3082
R537 VTAIL.n631 VTAIL.t9 52.3082
R538 VTAIL.n531 VTAIL.t8 52.3082
R539 VTAIL.n433 VTAIL.t7 52.3082
R540 VTAIL.n333 VTAIL.t5 52.3082
R541 VTAIL.n595 VTAIL.n594 43.4215
R542 VTAIL.n397 VTAIL.n396 43.4215
R543 VTAIL.n1 VTAIL.n0 43.4214
R544 VTAIL.n199 VTAIL.n198 43.4214
R545 VTAIL.n791 VTAIL.n790 31.6035
R546 VTAIL.n99 VTAIL.n98 31.6035
R547 VTAIL.n197 VTAIL.n196 31.6035
R548 VTAIL.n297 VTAIL.n296 31.6035
R549 VTAIL.n693 VTAIL.n692 31.6035
R550 VTAIL.n593 VTAIL.n592 31.6035
R551 VTAIL.n495 VTAIL.n494 31.6035
R552 VTAIL.n395 VTAIL.n394 31.6035
R553 VTAIL.n791 VTAIL.n693 31.0221
R554 VTAIL.n395 VTAIL.n297 31.0221
R555 VTAIL.n726 VTAIL.n725 15.6677
R556 VTAIL.n34 VTAIL.n33 15.6677
R557 VTAIL.n132 VTAIL.n131 15.6677
R558 VTAIL.n232 VTAIL.n231 15.6677
R559 VTAIL.n630 VTAIL.n629 15.6677
R560 VTAIL.n530 VTAIL.n529 15.6677
R561 VTAIL.n432 VTAIL.n431 15.6677
R562 VTAIL.n332 VTAIL.n331 15.6677
R563 VTAIL.n771 VTAIL.n702 13.1884
R564 VTAIL.n79 VTAIL.n10 13.1884
R565 VTAIL.n177 VTAIL.n108 13.1884
R566 VTAIL.n277 VTAIL.n208 13.1884
R567 VTAIL.n606 VTAIL.n604 13.1884
R568 VTAIL.n506 VTAIL.n504 13.1884
R569 VTAIL.n408 VTAIL.n406 13.1884
R570 VTAIL.n308 VTAIL.n306 13.1884
R571 VTAIL.n729 VTAIL.n724 12.8005
R572 VTAIL.n772 VTAIL.n704 12.8005
R573 VTAIL.n776 VTAIL.n775 12.8005
R574 VTAIL.n37 VTAIL.n32 12.8005
R575 VTAIL.n80 VTAIL.n12 12.8005
R576 VTAIL.n84 VTAIL.n83 12.8005
R577 VTAIL.n135 VTAIL.n130 12.8005
R578 VTAIL.n178 VTAIL.n110 12.8005
R579 VTAIL.n182 VTAIL.n181 12.8005
R580 VTAIL.n235 VTAIL.n230 12.8005
R581 VTAIL.n278 VTAIL.n210 12.8005
R582 VTAIL.n282 VTAIL.n281 12.8005
R583 VTAIL.n678 VTAIL.n677 12.8005
R584 VTAIL.n674 VTAIL.n673 12.8005
R585 VTAIL.n633 VTAIL.n628 12.8005
R586 VTAIL.n578 VTAIL.n577 12.8005
R587 VTAIL.n574 VTAIL.n573 12.8005
R588 VTAIL.n533 VTAIL.n528 12.8005
R589 VTAIL.n480 VTAIL.n479 12.8005
R590 VTAIL.n476 VTAIL.n475 12.8005
R591 VTAIL.n435 VTAIL.n430 12.8005
R592 VTAIL.n380 VTAIL.n379 12.8005
R593 VTAIL.n376 VTAIL.n375 12.8005
R594 VTAIL.n335 VTAIL.n330 12.8005
R595 VTAIL.n730 VTAIL.n722 12.0247
R596 VTAIL.n767 VTAIL.n766 12.0247
R597 VTAIL.n779 VTAIL.n700 12.0247
R598 VTAIL.n38 VTAIL.n30 12.0247
R599 VTAIL.n75 VTAIL.n74 12.0247
R600 VTAIL.n87 VTAIL.n8 12.0247
R601 VTAIL.n136 VTAIL.n128 12.0247
R602 VTAIL.n173 VTAIL.n172 12.0247
R603 VTAIL.n185 VTAIL.n106 12.0247
R604 VTAIL.n236 VTAIL.n228 12.0247
R605 VTAIL.n273 VTAIL.n272 12.0247
R606 VTAIL.n285 VTAIL.n206 12.0247
R607 VTAIL.n681 VTAIL.n602 12.0247
R608 VTAIL.n670 VTAIL.n607 12.0247
R609 VTAIL.n634 VTAIL.n626 12.0247
R610 VTAIL.n581 VTAIL.n502 12.0247
R611 VTAIL.n570 VTAIL.n507 12.0247
R612 VTAIL.n534 VTAIL.n526 12.0247
R613 VTAIL.n483 VTAIL.n404 12.0247
R614 VTAIL.n472 VTAIL.n409 12.0247
R615 VTAIL.n436 VTAIL.n428 12.0247
R616 VTAIL.n383 VTAIL.n304 12.0247
R617 VTAIL.n372 VTAIL.n309 12.0247
R618 VTAIL.n336 VTAIL.n328 12.0247
R619 VTAIL.n734 VTAIL.n733 11.249
R620 VTAIL.n765 VTAIL.n706 11.249
R621 VTAIL.n780 VTAIL.n698 11.249
R622 VTAIL.n42 VTAIL.n41 11.249
R623 VTAIL.n73 VTAIL.n14 11.249
R624 VTAIL.n88 VTAIL.n6 11.249
R625 VTAIL.n140 VTAIL.n139 11.249
R626 VTAIL.n171 VTAIL.n112 11.249
R627 VTAIL.n186 VTAIL.n104 11.249
R628 VTAIL.n240 VTAIL.n239 11.249
R629 VTAIL.n271 VTAIL.n212 11.249
R630 VTAIL.n286 VTAIL.n204 11.249
R631 VTAIL.n682 VTAIL.n600 11.249
R632 VTAIL.n669 VTAIL.n610 11.249
R633 VTAIL.n638 VTAIL.n637 11.249
R634 VTAIL.n582 VTAIL.n500 11.249
R635 VTAIL.n569 VTAIL.n510 11.249
R636 VTAIL.n538 VTAIL.n537 11.249
R637 VTAIL.n484 VTAIL.n402 11.249
R638 VTAIL.n471 VTAIL.n412 11.249
R639 VTAIL.n440 VTAIL.n439 11.249
R640 VTAIL.n384 VTAIL.n302 11.249
R641 VTAIL.n371 VTAIL.n312 11.249
R642 VTAIL.n340 VTAIL.n339 11.249
R643 VTAIL.n737 VTAIL.n720 10.4732
R644 VTAIL.n762 VTAIL.n761 10.4732
R645 VTAIL.n784 VTAIL.n783 10.4732
R646 VTAIL.n45 VTAIL.n28 10.4732
R647 VTAIL.n70 VTAIL.n69 10.4732
R648 VTAIL.n92 VTAIL.n91 10.4732
R649 VTAIL.n143 VTAIL.n126 10.4732
R650 VTAIL.n168 VTAIL.n167 10.4732
R651 VTAIL.n190 VTAIL.n189 10.4732
R652 VTAIL.n243 VTAIL.n226 10.4732
R653 VTAIL.n268 VTAIL.n267 10.4732
R654 VTAIL.n290 VTAIL.n289 10.4732
R655 VTAIL.n686 VTAIL.n685 10.4732
R656 VTAIL.n666 VTAIL.n665 10.4732
R657 VTAIL.n641 VTAIL.n624 10.4732
R658 VTAIL.n586 VTAIL.n585 10.4732
R659 VTAIL.n566 VTAIL.n565 10.4732
R660 VTAIL.n541 VTAIL.n524 10.4732
R661 VTAIL.n488 VTAIL.n487 10.4732
R662 VTAIL.n468 VTAIL.n467 10.4732
R663 VTAIL.n443 VTAIL.n426 10.4732
R664 VTAIL.n388 VTAIL.n387 10.4732
R665 VTAIL.n368 VTAIL.n367 10.4732
R666 VTAIL.n343 VTAIL.n326 10.4732
R667 VTAIL.n738 VTAIL.n718 9.69747
R668 VTAIL.n758 VTAIL.n708 9.69747
R669 VTAIL.n787 VTAIL.n696 9.69747
R670 VTAIL.n46 VTAIL.n26 9.69747
R671 VTAIL.n66 VTAIL.n16 9.69747
R672 VTAIL.n95 VTAIL.n4 9.69747
R673 VTAIL.n144 VTAIL.n124 9.69747
R674 VTAIL.n164 VTAIL.n114 9.69747
R675 VTAIL.n193 VTAIL.n102 9.69747
R676 VTAIL.n244 VTAIL.n224 9.69747
R677 VTAIL.n264 VTAIL.n214 9.69747
R678 VTAIL.n293 VTAIL.n202 9.69747
R679 VTAIL.n689 VTAIL.n598 9.69747
R680 VTAIL.n662 VTAIL.n612 9.69747
R681 VTAIL.n642 VTAIL.n622 9.69747
R682 VTAIL.n589 VTAIL.n498 9.69747
R683 VTAIL.n562 VTAIL.n512 9.69747
R684 VTAIL.n542 VTAIL.n522 9.69747
R685 VTAIL.n491 VTAIL.n400 9.69747
R686 VTAIL.n464 VTAIL.n414 9.69747
R687 VTAIL.n444 VTAIL.n424 9.69747
R688 VTAIL.n391 VTAIL.n300 9.69747
R689 VTAIL.n364 VTAIL.n314 9.69747
R690 VTAIL.n344 VTAIL.n324 9.69747
R691 VTAIL.n790 VTAIL.n789 9.45567
R692 VTAIL.n98 VTAIL.n97 9.45567
R693 VTAIL.n196 VTAIL.n195 9.45567
R694 VTAIL.n296 VTAIL.n295 9.45567
R695 VTAIL.n692 VTAIL.n691 9.45567
R696 VTAIL.n592 VTAIL.n591 9.45567
R697 VTAIL.n494 VTAIL.n493 9.45567
R698 VTAIL.n394 VTAIL.n393 9.45567
R699 VTAIL.n789 VTAIL.n788 9.3005
R700 VTAIL.n696 VTAIL.n695 9.3005
R701 VTAIL.n783 VTAIL.n782 9.3005
R702 VTAIL.n781 VTAIL.n780 9.3005
R703 VTAIL.n700 VTAIL.n699 9.3005
R704 VTAIL.n775 VTAIL.n774 9.3005
R705 VTAIL.n747 VTAIL.n746 9.3005
R706 VTAIL.n716 VTAIL.n715 9.3005
R707 VTAIL.n741 VTAIL.n740 9.3005
R708 VTAIL.n739 VTAIL.n738 9.3005
R709 VTAIL.n720 VTAIL.n719 9.3005
R710 VTAIL.n733 VTAIL.n732 9.3005
R711 VTAIL.n731 VTAIL.n730 9.3005
R712 VTAIL.n724 VTAIL.n723 9.3005
R713 VTAIL.n749 VTAIL.n748 9.3005
R714 VTAIL.n712 VTAIL.n711 9.3005
R715 VTAIL.n755 VTAIL.n754 9.3005
R716 VTAIL.n757 VTAIL.n756 9.3005
R717 VTAIL.n708 VTAIL.n707 9.3005
R718 VTAIL.n763 VTAIL.n762 9.3005
R719 VTAIL.n765 VTAIL.n764 9.3005
R720 VTAIL.n766 VTAIL.n703 9.3005
R721 VTAIL.n773 VTAIL.n772 9.3005
R722 VTAIL.n97 VTAIL.n96 9.3005
R723 VTAIL.n4 VTAIL.n3 9.3005
R724 VTAIL.n91 VTAIL.n90 9.3005
R725 VTAIL.n89 VTAIL.n88 9.3005
R726 VTAIL.n8 VTAIL.n7 9.3005
R727 VTAIL.n83 VTAIL.n82 9.3005
R728 VTAIL.n55 VTAIL.n54 9.3005
R729 VTAIL.n24 VTAIL.n23 9.3005
R730 VTAIL.n49 VTAIL.n48 9.3005
R731 VTAIL.n47 VTAIL.n46 9.3005
R732 VTAIL.n28 VTAIL.n27 9.3005
R733 VTAIL.n41 VTAIL.n40 9.3005
R734 VTAIL.n39 VTAIL.n38 9.3005
R735 VTAIL.n32 VTAIL.n31 9.3005
R736 VTAIL.n57 VTAIL.n56 9.3005
R737 VTAIL.n20 VTAIL.n19 9.3005
R738 VTAIL.n63 VTAIL.n62 9.3005
R739 VTAIL.n65 VTAIL.n64 9.3005
R740 VTAIL.n16 VTAIL.n15 9.3005
R741 VTAIL.n71 VTAIL.n70 9.3005
R742 VTAIL.n73 VTAIL.n72 9.3005
R743 VTAIL.n74 VTAIL.n11 9.3005
R744 VTAIL.n81 VTAIL.n80 9.3005
R745 VTAIL.n195 VTAIL.n194 9.3005
R746 VTAIL.n102 VTAIL.n101 9.3005
R747 VTAIL.n189 VTAIL.n188 9.3005
R748 VTAIL.n187 VTAIL.n186 9.3005
R749 VTAIL.n106 VTAIL.n105 9.3005
R750 VTAIL.n181 VTAIL.n180 9.3005
R751 VTAIL.n153 VTAIL.n152 9.3005
R752 VTAIL.n122 VTAIL.n121 9.3005
R753 VTAIL.n147 VTAIL.n146 9.3005
R754 VTAIL.n145 VTAIL.n144 9.3005
R755 VTAIL.n126 VTAIL.n125 9.3005
R756 VTAIL.n139 VTAIL.n138 9.3005
R757 VTAIL.n137 VTAIL.n136 9.3005
R758 VTAIL.n130 VTAIL.n129 9.3005
R759 VTAIL.n155 VTAIL.n154 9.3005
R760 VTAIL.n118 VTAIL.n117 9.3005
R761 VTAIL.n161 VTAIL.n160 9.3005
R762 VTAIL.n163 VTAIL.n162 9.3005
R763 VTAIL.n114 VTAIL.n113 9.3005
R764 VTAIL.n169 VTAIL.n168 9.3005
R765 VTAIL.n171 VTAIL.n170 9.3005
R766 VTAIL.n172 VTAIL.n109 9.3005
R767 VTAIL.n179 VTAIL.n178 9.3005
R768 VTAIL.n295 VTAIL.n294 9.3005
R769 VTAIL.n202 VTAIL.n201 9.3005
R770 VTAIL.n289 VTAIL.n288 9.3005
R771 VTAIL.n287 VTAIL.n286 9.3005
R772 VTAIL.n206 VTAIL.n205 9.3005
R773 VTAIL.n281 VTAIL.n280 9.3005
R774 VTAIL.n253 VTAIL.n252 9.3005
R775 VTAIL.n222 VTAIL.n221 9.3005
R776 VTAIL.n247 VTAIL.n246 9.3005
R777 VTAIL.n245 VTAIL.n244 9.3005
R778 VTAIL.n226 VTAIL.n225 9.3005
R779 VTAIL.n239 VTAIL.n238 9.3005
R780 VTAIL.n237 VTAIL.n236 9.3005
R781 VTAIL.n230 VTAIL.n229 9.3005
R782 VTAIL.n255 VTAIL.n254 9.3005
R783 VTAIL.n218 VTAIL.n217 9.3005
R784 VTAIL.n261 VTAIL.n260 9.3005
R785 VTAIL.n263 VTAIL.n262 9.3005
R786 VTAIL.n214 VTAIL.n213 9.3005
R787 VTAIL.n269 VTAIL.n268 9.3005
R788 VTAIL.n271 VTAIL.n270 9.3005
R789 VTAIL.n272 VTAIL.n209 9.3005
R790 VTAIL.n279 VTAIL.n278 9.3005
R791 VTAIL.n616 VTAIL.n615 9.3005
R792 VTAIL.n659 VTAIL.n658 9.3005
R793 VTAIL.n661 VTAIL.n660 9.3005
R794 VTAIL.n612 VTAIL.n611 9.3005
R795 VTAIL.n667 VTAIL.n666 9.3005
R796 VTAIL.n669 VTAIL.n668 9.3005
R797 VTAIL.n607 VTAIL.n605 9.3005
R798 VTAIL.n675 VTAIL.n674 9.3005
R799 VTAIL.n691 VTAIL.n690 9.3005
R800 VTAIL.n598 VTAIL.n597 9.3005
R801 VTAIL.n685 VTAIL.n684 9.3005
R802 VTAIL.n683 VTAIL.n682 9.3005
R803 VTAIL.n602 VTAIL.n601 9.3005
R804 VTAIL.n677 VTAIL.n676 9.3005
R805 VTAIL.n653 VTAIL.n652 9.3005
R806 VTAIL.n651 VTAIL.n650 9.3005
R807 VTAIL.n620 VTAIL.n619 9.3005
R808 VTAIL.n645 VTAIL.n644 9.3005
R809 VTAIL.n643 VTAIL.n642 9.3005
R810 VTAIL.n624 VTAIL.n623 9.3005
R811 VTAIL.n637 VTAIL.n636 9.3005
R812 VTAIL.n635 VTAIL.n634 9.3005
R813 VTAIL.n628 VTAIL.n627 9.3005
R814 VTAIL.n516 VTAIL.n515 9.3005
R815 VTAIL.n559 VTAIL.n558 9.3005
R816 VTAIL.n561 VTAIL.n560 9.3005
R817 VTAIL.n512 VTAIL.n511 9.3005
R818 VTAIL.n567 VTAIL.n566 9.3005
R819 VTAIL.n569 VTAIL.n568 9.3005
R820 VTAIL.n507 VTAIL.n505 9.3005
R821 VTAIL.n575 VTAIL.n574 9.3005
R822 VTAIL.n591 VTAIL.n590 9.3005
R823 VTAIL.n498 VTAIL.n497 9.3005
R824 VTAIL.n585 VTAIL.n584 9.3005
R825 VTAIL.n583 VTAIL.n582 9.3005
R826 VTAIL.n502 VTAIL.n501 9.3005
R827 VTAIL.n577 VTAIL.n576 9.3005
R828 VTAIL.n553 VTAIL.n552 9.3005
R829 VTAIL.n551 VTAIL.n550 9.3005
R830 VTAIL.n520 VTAIL.n519 9.3005
R831 VTAIL.n545 VTAIL.n544 9.3005
R832 VTAIL.n543 VTAIL.n542 9.3005
R833 VTAIL.n524 VTAIL.n523 9.3005
R834 VTAIL.n537 VTAIL.n536 9.3005
R835 VTAIL.n535 VTAIL.n534 9.3005
R836 VTAIL.n528 VTAIL.n527 9.3005
R837 VTAIL.n418 VTAIL.n417 9.3005
R838 VTAIL.n461 VTAIL.n460 9.3005
R839 VTAIL.n463 VTAIL.n462 9.3005
R840 VTAIL.n414 VTAIL.n413 9.3005
R841 VTAIL.n469 VTAIL.n468 9.3005
R842 VTAIL.n471 VTAIL.n470 9.3005
R843 VTAIL.n409 VTAIL.n407 9.3005
R844 VTAIL.n477 VTAIL.n476 9.3005
R845 VTAIL.n493 VTAIL.n492 9.3005
R846 VTAIL.n400 VTAIL.n399 9.3005
R847 VTAIL.n487 VTAIL.n486 9.3005
R848 VTAIL.n485 VTAIL.n484 9.3005
R849 VTAIL.n404 VTAIL.n403 9.3005
R850 VTAIL.n479 VTAIL.n478 9.3005
R851 VTAIL.n455 VTAIL.n454 9.3005
R852 VTAIL.n453 VTAIL.n452 9.3005
R853 VTAIL.n422 VTAIL.n421 9.3005
R854 VTAIL.n447 VTAIL.n446 9.3005
R855 VTAIL.n445 VTAIL.n444 9.3005
R856 VTAIL.n426 VTAIL.n425 9.3005
R857 VTAIL.n439 VTAIL.n438 9.3005
R858 VTAIL.n437 VTAIL.n436 9.3005
R859 VTAIL.n430 VTAIL.n429 9.3005
R860 VTAIL.n318 VTAIL.n317 9.3005
R861 VTAIL.n361 VTAIL.n360 9.3005
R862 VTAIL.n363 VTAIL.n362 9.3005
R863 VTAIL.n314 VTAIL.n313 9.3005
R864 VTAIL.n369 VTAIL.n368 9.3005
R865 VTAIL.n371 VTAIL.n370 9.3005
R866 VTAIL.n309 VTAIL.n307 9.3005
R867 VTAIL.n377 VTAIL.n376 9.3005
R868 VTAIL.n393 VTAIL.n392 9.3005
R869 VTAIL.n300 VTAIL.n299 9.3005
R870 VTAIL.n387 VTAIL.n386 9.3005
R871 VTAIL.n385 VTAIL.n384 9.3005
R872 VTAIL.n304 VTAIL.n303 9.3005
R873 VTAIL.n379 VTAIL.n378 9.3005
R874 VTAIL.n355 VTAIL.n354 9.3005
R875 VTAIL.n353 VTAIL.n352 9.3005
R876 VTAIL.n322 VTAIL.n321 9.3005
R877 VTAIL.n347 VTAIL.n346 9.3005
R878 VTAIL.n345 VTAIL.n344 9.3005
R879 VTAIL.n326 VTAIL.n325 9.3005
R880 VTAIL.n339 VTAIL.n338 9.3005
R881 VTAIL.n337 VTAIL.n336 9.3005
R882 VTAIL.n330 VTAIL.n329 9.3005
R883 VTAIL.n742 VTAIL.n741 8.92171
R884 VTAIL.n757 VTAIL.n710 8.92171
R885 VTAIL.n788 VTAIL.n694 8.92171
R886 VTAIL.n50 VTAIL.n49 8.92171
R887 VTAIL.n65 VTAIL.n18 8.92171
R888 VTAIL.n96 VTAIL.n2 8.92171
R889 VTAIL.n148 VTAIL.n147 8.92171
R890 VTAIL.n163 VTAIL.n116 8.92171
R891 VTAIL.n194 VTAIL.n100 8.92171
R892 VTAIL.n248 VTAIL.n247 8.92171
R893 VTAIL.n263 VTAIL.n216 8.92171
R894 VTAIL.n294 VTAIL.n200 8.92171
R895 VTAIL.n690 VTAIL.n596 8.92171
R896 VTAIL.n661 VTAIL.n614 8.92171
R897 VTAIL.n646 VTAIL.n645 8.92171
R898 VTAIL.n590 VTAIL.n496 8.92171
R899 VTAIL.n561 VTAIL.n514 8.92171
R900 VTAIL.n546 VTAIL.n545 8.92171
R901 VTAIL.n492 VTAIL.n398 8.92171
R902 VTAIL.n463 VTAIL.n416 8.92171
R903 VTAIL.n448 VTAIL.n447 8.92171
R904 VTAIL.n392 VTAIL.n298 8.92171
R905 VTAIL.n363 VTAIL.n316 8.92171
R906 VTAIL.n348 VTAIL.n347 8.92171
R907 VTAIL.n745 VTAIL.n716 8.14595
R908 VTAIL.n754 VTAIL.n753 8.14595
R909 VTAIL.n53 VTAIL.n24 8.14595
R910 VTAIL.n62 VTAIL.n61 8.14595
R911 VTAIL.n151 VTAIL.n122 8.14595
R912 VTAIL.n160 VTAIL.n159 8.14595
R913 VTAIL.n251 VTAIL.n222 8.14595
R914 VTAIL.n260 VTAIL.n259 8.14595
R915 VTAIL.n658 VTAIL.n657 8.14595
R916 VTAIL.n649 VTAIL.n620 8.14595
R917 VTAIL.n558 VTAIL.n557 8.14595
R918 VTAIL.n549 VTAIL.n520 8.14595
R919 VTAIL.n460 VTAIL.n459 8.14595
R920 VTAIL.n451 VTAIL.n422 8.14595
R921 VTAIL.n360 VTAIL.n359 8.14595
R922 VTAIL.n351 VTAIL.n322 8.14595
R923 VTAIL.n746 VTAIL.n714 7.3702
R924 VTAIL.n750 VTAIL.n712 7.3702
R925 VTAIL.n54 VTAIL.n22 7.3702
R926 VTAIL.n58 VTAIL.n20 7.3702
R927 VTAIL.n152 VTAIL.n120 7.3702
R928 VTAIL.n156 VTAIL.n118 7.3702
R929 VTAIL.n252 VTAIL.n220 7.3702
R930 VTAIL.n256 VTAIL.n218 7.3702
R931 VTAIL.n654 VTAIL.n616 7.3702
R932 VTAIL.n650 VTAIL.n618 7.3702
R933 VTAIL.n554 VTAIL.n516 7.3702
R934 VTAIL.n550 VTAIL.n518 7.3702
R935 VTAIL.n456 VTAIL.n418 7.3702
R936 VTAIL.n452 VTAIL.n420 7.3702
R937 VTAIL.n356 VTAIL.n318 7.3702
R938 VTAIL.n352 VTAIL.n320 7.3702
R939 VTAIL.n749 VTAIL.n714 6.59444
R940 VTAIL.n750 VTAIL.n749 6.59444
R941 VTAIL.n57 VTAIL.n22 6.59444
R942 VTAIL.n58 VTAIL.n57 6.59444
R943 VTAIL.n155 VTAIL.n120 6.59444
R944 VTAIL.n156 VTAIL.n155 6.59444
R945 VTAIL.n255 VTAIL.n220 6.59444
R946 VTAIL.n256 VTAIL.n255 6.59444
R947 VTAIL.n654 VTAIL.n653 6.59444
R948 VTAIL.n653 VTAIL.n618 6.59444
R949 VTAIL.n554 VTAIL.n553 6.59444
R950 VTAIL.n553 VTAIL.n518 6.59444
R951 VTAIL.n456 VTAIL.n455 6.59444
R952 VTAIL.n455 VTAIL.n420 6.59444
R953 VTAIL.n356 VTAIL.n355 6.59444
R954 VTAIL.n355 VTAIL.n320 6.59444
R955 VTAIL.n746 VTAIL.n745 5.81868
R956 VTAIL.n753 VTAIL.n712 5.81868
R957 VTAIL.n54 VTAIL.n53 5.81868
R958 VTAIL.n61 VTAIL.n20 5.81868
R959 VTAIL.n152 VTAIL.n151 5.81868
R960 VTAIL.n159 VTAIL.n118 5.81868
R961 VTAIL.n252 VTAIL.n251 5.81868
R962 VTAIL.n259 VTAIL.n218 5.81868
R963 VTAIL.n657 VTAIL.n616 5.81868
R964 VTAIL.n650 VTAIL.n649 5.81868
R965 VTAIL.n557 VTAIL.n516 5.81868
R966 VTAIL.n550 VTAIL.n549 5.81868
R967 VTAIL.n459 VTAIL.n418 5.81868
R968 VTAIL.n452 VTAIL.n451 5.81868
R969 VTAIL.n359 VTAIL.n318 5.81868
R970 VTAIL.n352 VTAIL.n351 5.81868
R971 VTAIL.n742 VTAIL.n716 5.04292
R972 VTAIL.n754 VTAIL.n710 5.04292
R973 VTAIL.n790 VTAIL.n694 5.04292
R974 VTAIL.n50 VTAIL.n24 5.04292
R975 VTAIL.n62 VTAIL.n18 5.04292
R976 VTAIL.n98 VTAIL.n2 5.04292
R977 VTAIL.n148 VTAIL.n122 5.04292
R978 VTAIL.n160 VTAIL.n116 5.04292
R979 VTAIL.n196 VTAIL.n100 5.04292
R980 VTAIL.n248 VTAIL.n222 5.04292
R981 VTAIL.n260 VTAIL.n216 5.04292
R982 VTAIL.n296 VTAIL.n200 5.04292
R983 VTAIL.n692 VTAIL.n596 5.04292
R984 VTAIL.n658 VTAIL.n614 5.04292
R985 VTAIL.n646 VTAIL.n620 5.04292
R986 VTAIL.n592 VTAIL.n496 5.04292
R987 VTAIL.n558 VTAIL.n514 5.04292
R988 VTAIL.n546 VTAIL.n520 5.04292
R989 VTAIL.n494 VTAIL.n398 5.04292
R990 VTAIL.n460 VTAIL.n416 5.04292
R991 VTAIL.n448 VTAIL.n422 5.04292
R992 VTAIL.n394 VTAIL.n298 5.04292
R993 VTAIL.n360 VTAIL.n316 5.04292
R994 VTAIL.n348 VTAIL.n322 5.04292
R995 VTAIL.n725 VTAIL.n723 4.38563
R996 VTAIL.n33 VTAIL.n31 4.38563
R997 VTAIL.n131 VTAIL.n129 4.38563
R998 VTAIL.n231 VTAIL.n229 4.38563
R999 VTAIL.n629 VTAIL.n627 4.38563
R1000 VTAIL.n529 VTAIL.n527 4.38563
R1001 VTAIL.n431 VTAIL.n429 4.38563
R1002 VTAIL.n331 VTAIL.n329 4.38563
R1003 VTAIL.n741 VTAIL.n718 4.26717
R1004 VTAIL.n758 VTAIL.n757 4.26717
R1005 VTAIL.n788 VTAIL.n787 4.26717
R1006 VTAIL.n49 VTAIL.n26 4.26717
R1007 VTAIL.n66 VTAIL.n65 4.26717
R1008 VTAIL.n96 VTAIL.n95 4.26717
R1009 VTAIL.n147 VTAIL.n124 4.26717
R1010 VTAIL.n164 VTAIL.n163 4.26717
R1011 VTAIL.n194 VTAIL.n193 4.26717
R1012 VTAIL.n247 VTAIL.n224 4.26717
R1013 VTAIL.n264 VTAIL.n263 4.26717
R1014 VTAIL.n294 VTAIL.n293 4.26717
R1015 VTAIL.n690 VTAIL.n689 4.26717
R1016 VTAIL.n662 VTAIL.n661 4.26717
R1017 VTAIL.n645 VTAIL.n622 4.26717
R1018 VTAIL.n590 VTAIL.n589 4.26717
R1019 VTAIL.n562 VTAIL.n561 4.26717
R1020 VTAIL.n545 VTAIL.n522 4.26717
R1021 VTAIL.n492 VTAIL.n491 4.26717
R1022 VTAIL.n464 VTAIL.n463 4.26717
R1023 VTAIL.n447 VTAIL.n424 4.26717
R1024 VTAIL.n392 VTAIL.n391 4.26717
R1025 VTAIL.n364 VTAIL.n363 4.26717
R1026 VTAIL.n347 VTAIL.n324 4.26717
R1027 VTAIL.n397 VTAIL.n395 3.57809
R1028 VTAIL.n495 VTAIL.n397 3.57809
R1029 VTAIL.n595 VTAIL.n593 3.57809
R1030 VTAIL.n693 VTAIL.n595 3.57809
R1031 VTAIL.n297 VTAIL.n199 3.57809
R1032 VTAIL.n199 VTAIL.n197 3.57809
R1033 VTAIL.n99 VTAIL.n1 3.57809
R1034 VTAIL VTAIL.n791 3.5199
R1035 VTAIL.n738 VTAIL.n737 3.49141
R1036 VTAIL.n761 VTAIL.n708 3.49141
R1037 VTAIL.n784 VTAIL.n696 3.49141
R1038 VTAIL.n46 VTAIL.n45 3.49141
R1039 VTAIL.n69 VTAIL.n16 3.49141
R1040 VTAIL.n92 VTAIL.n4 3.49141
R1041 VTAIL.n144 VTAIL.n143 3.49141
R1042 VTAIL.n167 VTAIL.n114 3.49141
R1043 VTAIL.n190 VTAIL.n102 3.49141
R1044 VTAIL.n244 VTAIL.n243 3.49141
R1045 VTAIL.n267 VTAIL.n214 3.49141
R1046 VTAIL.n290 VTAIL.n202 3.49141
R1047 VTAIL.n686 VTAIL.n598 3.49141
R1048 VTAIL.n665 VTAIL.n612 3.49141
R1049 VTAIL.n642 VTAIL.n641 3.49141
R1050 VTAIL.n586 VTAIL.n498 3.49141
R1051 VTAIL.n565 VTAIL.n512 3.49141
R1052 VTAIL.n542 VTAIL.n541 3.49141
R1053 VTAIL.n488 VTAIL.n400 3.49141
R1054 VTAIL.n467 VTAIL.n414 3.49141
R1055 VTAIL.n444 VTAIL.n443 3.49141
R1056 VTAIL.n388 VTAIL.n300 3.49141
R1057 VTAIL.n367 VTAIL.n314 3.49141
R1058 VTAIL.n344 VTAIL.n343 3.49141
R1059 VTAIL.n734 VTAIL.n720 2.71565
R1060 VTAIL.n762 VTAIL.n706 2.71565
R1061 VTAIL.n783 VTAIL.n698 2.71565
R1062 VTAIL.n42 VTAIL.n28 2.71565
R1063 VTAIL.n70 VTAIL.n14 2.71565
R1064 VTAIL.n91 VTAIL.n6 2.71565
R1065 VTAIL.n140 VTAIL.n126 2.71565
R1066 VTAIL.n168 VTAIL.n112 2.71565
R1067 VTAIL.n189 VTAIL.n104 2.71565
R1068 VTAIL.n240 VTAIL.n226 2.71565
R1069 VTAIL.n268 VTAIL.n212 2.71565
R1070 VTAIL.n289 VTAIL.n204 2.71565
R1071 VTAIL.n685 VTAIL.n600 2.71565
R1072 VTAIL.n666 VTAIL.n610 2.71565
R1073 VTAIL.n638 VTAIL.n624 2.71565
R1074 VTAIL.n585 VTAIL.n500 2.71565
R1075 VTAIL.n566 VTAIL.n510 2.71565
R1076 VTAIL.n538 VTAIL.n524 2.71565
R1077 VTAIL.n487 VTAIL.n402 2.71565
R1078 VTAIL.n468 VTAIL.n412 2.71565
R1079 VTAIL.n440 VTAIL.n426 2.71565
R1080 VTAIL.n387 VTAIL.n302 2.71565
R1081 VTAIL.n368 VTAIL.n312 2.71565
R1082 VTAIL.n340 VTAIL.n326 2.71565
R1083 VTAIL.n733 VTAIL.n722 1.93989
R1084 VTAIL.n767 VTAIL.n765 1.93989
R1085 VTAIL.n780 VTAIL.n779 1.93989
R1086 VTAIL.n41 VTAIL.n30 1.93989
R1087 VTAIL.n75 VTAIL.n73 1.93989
R1088 VTAIL.n88 VTAIL.n87 1.93989
R1089 VTAIL.n139 VTAIL.n128 1.93989
R1090 VTAIL.n173 VTAIL.n171 1.93989
R1091 VTAIL.n186 VTAIL.n185 1.93989
R1092 VTAIL.n239 VTAIL.n228 1.93989
R1093 VTAIL.n273 VTAIL.n271 1.93989
R1094 VTAIL.n286 VTAIL.n285 1.93989
R1095 VTAIL.n682 VTAIL.n681 1.93989
R1096 VTAIL.n670 VTAIL.n669 1.93989
R1097 VTAIL.n637 VTAIL.n626 1.93989
R1098 VTAIL.n582 VTAIL.n581 1.93989
R1099 VTAIL.n570 VTAIL.n569 1.93989
R1100 VTAIL.n537 VTAIL.n526 1.93989
R1101 VTAIL.n484 VTAIL.n483 1.93989
R1102 VTAIL.n472 VTAIL.n471 1.93989
R1103 VTAIL.n439 VTAIL.n428 1.93989
R1104 VTAIL.n384 VTAIL.n383 1.93989
R1105 VTAIL.n372 VTAIL.n371 1.93989
R1106 VTAIL.n339 VTAIL.n328 1.93989
R1107 VTAIL.n730 VTAIL.n729 1.16414
R1108 VTAIL.n766 VTAIL.n704 1.16414
R1109 VTAIL.n776 VTAIL.n700 1.16414
R1110 VTAIL.n38 VTAIL.n37 1.16414
R1111 VTAIL.n74 VTAIL.n12 1.16414
R1112 VTAIL.n84 VTAIL.n8 1.16414
R1113 VTAIL.n136 VTAIL.n135 1.16414
R1114 VTAIL.n172 VTAIL.n110 1.16414
R1115 VTAIL.n182 VTAIL.n106 1.16414
R1116 VTAIL.n236 VTAIL.n235 1.16414
R1117 VTAIL.n272 VTAIL.n210 1.16414
R1118 VTAIL.n282 VTAIL.n206 1.16414
R1119 VTAIL.n678 VTAIL.n602 1.16414
R1120 VTAIL.n673 VTAIL.n607 1.16414
R1121 VTAIL.n634 VTAIL.n633 1.16414
R1122 VTAIL.n578 VTAIL.n502 1.16414
R1123 VTAIL.n573 VTAIL.n507 1.16414
R1124 VTAIL.n534 VTAIL.n533 1.16414
R1125 VTAIL.n480 VTAIL.n404 1.16414
R1126 VTAIL.n475 VTAIL.n409 1.16414
R1127 VTAIL.n436 VTAIL.n435 1.16414
R1128 VTAIL.n380 VTAIL.n304 1.16414
R1129 VTAIL.n375 VTAIL.n309 1.16414
R1130 VTAIL.n336 VTAIL.n335 1.16414
R1131 VTAIL.n0 VTAIL.t0 1.13258
R1132 VTAIL.n0 VTAIL.t3 1.13258
R1133 VTAIL.n198 VTAIL.t12 1.13258
R1134 VTAIL.n198 VTAIL.t13 1.13258
R1135 VTAIL.n594 VTAIL.t15 1.13258
R1136 VTAIL.n594 VTAIL.t10 1.13258
R1137 VTAIL.n396 VTAIL.t2 1.13258
R1138 VTAIL.n396 VTAIL.t6 1.13258
R1139 VTAIL.n593 VTAIL.n495 0.470328
R1140 VTAIL.n197 VTAIL.n99 0.470328
R1141 VTAIL.n726 VTAIL.n724 0.388379
R1142 VTAIL.n772 VTAIL.n771 0.388379
R1143 VTAIL.n775 VTAIL.n702 0.388379
R1144 VTAIL.n34 VTAIL.n32 0.388379
R1145 VTAIL.n80 VTAIL.n79 0.388379
R1146 VTAIL.n83 VTAIL.n10 0.388379
R1147 VTAIL.n132 VTAIL.n130 0.388379
R1148 VTAIL.n178 VTAIL.n177 0.388379
R1149 VTAIL.n181 VTAIL.n108 0.388379
R1150 VTAIL.n232 VTAIL.n230 0.388379
R1151 VTAIL.n278 VTAIL.n277 0.388379
R1152 VTAIL.n281 VTAIL.n208 0.388379
R1153 VTAIL.n677 VTAIL.n604 0.388379
R1154 VTAIL.n674 VTAIL.n606 0.388379
R1155 VTAIL.n630 VTAIL.n628 0.388379
R1156 VTAIL.n577 VTAIL.n504 0.388379
R1157 VTAIL.n574 VTAIL.n506 0.388379
R1158 VTAIL.n530 VTAIL.n528 0.388379
R1159 VTAIL.n479 VTAIL.n406 0.388379
R1160 VTAIL.n476 VTAIL.n408 0.388379
R1161 VTAIL.n432 VTAIL.n430 0.388379
R1162 VTAIL.n379 VTAIL.n306 0.388379
R1163 VTAIL.n376 VTAIL.n308 0.388379
R1164 VTAIL.n332 VTAIL.n330 0.388379
R1165 VTAIL.n731 VTAIL.n723 0.155672
R1166 VTAIL.n732 VTAIL.n731 0.155672
R1167 VTAIL.n732 VTAIL.n719 0.155672
R1168 VTAIL.n739 VTAIL.n719 0.155672
R1169 VTAIL.n740 VTAIL.n739 0.155672
R1170 VTAIL.n740 VTAIL.n715 0.155672
R1171 VTAIL.n747 VTAIL.n715 0.155672
R1172 VTAIL.n748 VTAIL.n747 0.155672
R1173 VTAIL.n748 VTAIL.n711 0.155672
R1174 VTAIL.n755 VTAIL.n711 0.155672
R1175 VTAIL.n756 VTAIL.n755 0.155672
R1176 VTAIL.n756 VTAIL.n707 0.155672
R1177 VTAIL.n763 VTAIL.n707 0.155672
R1178 VTAIL.n764 VTAIL.n763 0.155672
R1179 VTAIL.n764 VTAIL.n703 0.155672
R1180 VTAIL.n773 VTAIL.n703 0.155672
R1181 VTAIL.n774 VTAIL.n773 0.155672
R1182 VTAIL.n774 VTAIL.n699 0.155672
R1183 VTAIL.n781 VTAIL.n699 0.155672
R1184 VTAIL.n782 VTAIL.n781 0.155672
R1185 VTAIL.n782 VTAIL.n695 0.155672
R1186 VTAIL.n789 VTAIL.n695 0.155672
R1187 VTAIL.n39 VTAIL.n31 0.155672
R1188 VTAIL.n40 VTAIL.n39 0.155672
R1189 VTAIL.n40 VTAIL.n27 0.155672
R1190 VTAIL.n47 VTAIL.n27 0.155672
R1191 VTAIL.n48 VTAIL.n47 0.155672
R1192 VTAIL.n48 VTAIL.n23 0.155672
R1193 VTAIL.n55 VTAIL.n23 0.155672
R1194 VTAIL.n56 VTAIL.n55 0.155672
R1195 VTAIL.n56 VTAIL.n19 0.155672
R1196 VTAIL.n63 VTAIL.n19 0.155672
R1197 VTAIL.n64 VTAIL.n63 0.155672
R1198 VTAIL.n64 VTAIL.n15 0.155672
R1199 VTAIL.n71 VTAIL.n15 0.155672
R1200 VTAIL.n72 VTAIL.n71 0.155672
R1201 VTAIL.n72 VTAIL.n11 0.155672
R1202 VTAIL.n81 VTAIL.n11 0.155672
R1203 VTAIL.n82 VTAIL.n81 0.155672
R1204 VTAIL.n82 VTAIL.n7 0.155672
R1205 VTAIL.n89 VTAIL.n7 0.155672
R1206 VTAIL.n90 VTAIL.n89 0.155672
R1207 VTAIL.n90 VTAIL.n3 0.155672
R1208 VTAIL.n97 VTAIL.n3 0.155672
R1209 VTAIL.n137 VTAIL.n129 0.155672
R1210 VTAIL.n138 VTAIL.n137 0.155672
R1211 VTAIL.n138 VTAIL.n125 0.155672
R1212 VTAIL.n145 VTAIL.n125 0.155672
R1213 VTAIL.n146 VTAIL.n145 0.155672
R1214 VTAIL.n146 VTAIL.n121 0.155672
R1215 VTAIL.n153 VTAIL.n121 0.155672
R1216 VTAIL.n154 VTAIL.n153 0.155672
R1217 VTAIL.n154 VTAIL.n117 0.155672
R1218 VTAIL.n161 VTAIL.n117 0.155672
R1219 VTAIL.n162 VTAIL.n161 0.155672
R1220 VTAIL.n162 VTAIL.n113 0.155672
R1221 VTAIL.n169 VTAIL.n113 0.155672
R1222 VTAIL.n170 VTAIL.n169 0.155672
R1223 VTAIL.n170 VTAIL.n109 0.155672
R1224 VTAIL.n179 VTAIL.n109 0.155672
R1225 VTAIL.n180 VTAIL.n179 0.155672
R1226 VTAIL.n180 VTAIL.n105 0.155672
R1227 VTAIL.n187 VTAIL.n105 0.155672
R1228 VTAIL.n188 VTAIL.n187 0.155672
R1229 VTAIL.n188 VTAIL.n101 0.155672
R1230 VTAIL.n195 VTAIL.n101 0.155672
R1231 VTAIL.n237 VTAIL.n229 0.155672
R1232 VTAIL.n238 VTAIL.n237 0.155672
R1233 VTAIL.n238 VTAIL.n225 0.155672
R1234 VTAIL.n245 VTAIL.n225 0.155672
R1235 VTAIL.n246 VTAIL.n245 0.155672
R1236 VTAIL.n246 VTAIL.n221 0.155672
R1237 VTAIL.n253 VTAIL.n221 0.155672
R1238 VTAIL.n254 VTAIL.n253 0.155672
R1239 VTAIL.n254 VTAIL.n217 0.155672
R1240 VTAIL.n261 VTAIL.n217 0.155672
R1241 VTAIL.n262 VTAIL.n261 0.155672
R1242 VTAIL.n262 VTAIL.n213 0.155672
R1243 VTAIL.n269 VTAIL.n213 0.155672
R1244 VTAIL.n270 VTAIL.n269 0.155672
R1245 VTAIL.n270 VTAIL.n209 0.155672
R1246 VTAIL.n279 VTAIL.n209 0.155672
R1247 VTAIL.n280 VTAIL.n279 0.155672
R1248 VTAIL.n280 VTAIL.n205 0.155672
R1249 VTAIL.n287 VTAIL.n205 0.155672
R1250 VTAIL.n288 VTAIL.n287 0.155672
R1251 VTAIL.n288 VTAIL.n201 0.155672
R1252 VTAIL.n295 VTAIL.n201 0.155672
R1253 VTAIL.n691 VTAIL.n597 0.155672
R1254 VTAIL.n684 VTAIL.n597 0.155672
R1255 VTAIL.n684 VTAIL.n683 0.155672
R1256 VTAIL.n683 VTAIL.n601 0.155672
R1257 VTAIL.n676 VTAIL.n601 0.155672
R1258 VTAIL.n676 VTAIL.n675 0.155672
R1259 VTAIL.n675 VTAIL.n605 0.155672
R1260 VTAIL.n668 VTAIL.n605 0.155672
R1261 VTAIL.n668 VTAIL.n667 0.155672
R1262 VTAIL.n667 VTAIL.n611 0.155672
R1263 VTAIL.n660 VTAIL.n611 0.155672
R1264 VTAIL.n660 VTAIL.n659 0.155672
R1265 VTAIL.n659 VTAIL.n615 0.155672
R1266 VTAIL.n652 VTAIL.n615 0.155672
R1267 VTAIL.n652 VTAIL.n651 0.155672
R1268 VTAIL.n651 VTAIL.n619 0.155672
R1269 VTAIL.n644 VTAIL.n619 0.155672
R1270 VTAIL.n644 VTAIL.n643 0.155672
R1271 VTAIL.n643 VTAIL.n623 0.155672
R1272 VTAIL.n636 VTAIL.n623 0.155672
R1273 VTAIL.n636 VTAIL.n635 0.155672
R1274 VTAIL.n635 VTAIL.n627 0.155672
R1275 VTAIL.n591 VTAIL.n497 0.155672
R1276 VTAIL.n584 VTAIL.n497 0.155672
R1277 VTAIL.n584 VTAIL.n583 0.155672
R1278 VTAIL.n583 VTAIL.n501 0.155672
R1279 VTAIL.n576 VTAIL.n501 0.155672
R1280 VTAIL.n576 VTAIL.n575 0.155672
R1281 VTAIL.n575 VTAIL.n505 0.155672
R1282 VTAIL.n568 VTAIL.n505 0.155672
R1283 VTAIL.n568 VTAIL.n567 0.155672
R1284 VTAIL.n567 VTAIL.n511 0.155672
R1285 VTAIL.n560 VTAIL.n511 0.155672
R1286 VTAIL.n560 VTAIL.n559 0.155672
R1287 VTAIL.n559 VTAIL.n515 0.155672
R1288 VTAIL.n552 VTAIL.n515 0.155672
R1289 VTAIL.n552 VTAIL.n551 0.155672
R1290 VTAIL.n551 VTAIL.n519 0.155672
R1291 VTAIL.n544 VTAIL.n519 0.155672
R1292 VTAIL.n544 VTAIL.n543 0.155672
R1293 VTAIL.n543 VTAIL.n523 0.155672
R1294 VTAIL.n536 VTAIL.n523 0.155672
R1295 VTAIL.n536 VTAIL.n535 0.155672
R1296 VTAIL.n535 VTAIL.n527 0.155672
R1297 VTAIL.n493 VTAIL.n399 0.155672
R1298 VTAIL.n486 VTAIL.n399 0.155672
R1299 VTAIL.n486 VTAIL.n485 0.155672
R1300 VTAIL.n485 VTAIL.n403 0.155672
R1301 VTAIL.n478 VTAIL.n403 0.155672
R1302 VTAIL.n478 VTAIL.n477 0.155672
R1303 VTAIL.n477 VTAIL.n407 0.155672
R1304 VTAIL.n470 VTAIL.n407 0.155672
R1305 VTAIL.n470 VTAIL.n469 0.155672
R1306 VTAIL.n469 VTAIL.n413 0.155672
R1307 VTAIL.n462 VTAIL.n413 0.155672
R1308 VTAIL.n462 VTAIL.n461 0.155672
R1309 VTAIL.n461 VTAIL.n417 0.155672
R1310 VTAIL.n454 VTAIL.n417 0.155672
R1311 VTAIL.n454 VTAIL.n453 0.155672
R1312 VTAIL.n453 VTAIL.n421 0.155672
R1313 VTAIL.n446 VTAIL.n421 0.155672
R1314 VTAIL.n446 VTAIL.n445 0.155672
R1315 VTAIL.n445 VTAIL.n425 0.155672
R1316 VTAIL.n438 VTAIL.n425 0.155672
R1317 VTAIL.n438 VTAIL.n437 0.155672
R1318 VTAIL.n437 VTAIL.n429 0.155672
R1319 VTAIL.n393 VTAIL.n299 0.155672
R1320 VTAIL.n386 VTAIL.n299 0.155672
R1321 VTAIL.n386 VTAIL.n385 0.155672
R1322 VTAIL.n385 VTAIL.n303 0.155672
R1323 VTAIL.n378 VTAIL.n303 0.155672
R1324 VTAIL.n378 VTAIL.n377 0.155672
R1325 VTAIL.n377 VTAIL.n307 0.155672
R1326 VTAIL.n370 VTAIL.n307 0.155672
R1327 VTAIL.n370 VTAIL.n369 0.155672
R1328 VTAIL.n369 VTAIL.n313 0.155672
R1329 VTAIL.n362 VTAIL.n313 0.155672
R1330 VTAIL.n362 VTAIL.n361 0.155672
R1331 VTAIL.n361 VTAIL.n317 0.155672
R1332 VTAIL.n354 VTAIL.n317 0.155672
R1333 VTAIL.n354 VTAIL.n353 0.155672
R1334 VTAIL.n353 VTAIL.n321 0.155672
R1335 VTAIL.n346 VTAIL.n321 0.155672
R1336 VTAIL.n346 VTAIL.n345 0.155672
R1337 VTAIL.n345 VTAIL.n325 0.155672
R1338 VTAIL.n338 VTAIL.n325 0.155672
R1339 VTAIL.n338 VTAIL.n337 0.155672
R1340 VTAIL.n337 VTAIL.n329 0.155672
R1341 VTAIL VTAIL.n1 0.0586897
R1342 VDD1 VDD1.n0 61.9473
R1343 VDD1.n3 VDD1.n2 61.8336
R1344 VDD1.n3 VDD1.n1 61.8336
R1345 VDD1.n5 VDD1.n4 60.1001
R1346 VDD1.n5 VDD1.n3 55.475
R1347 VDD1 VDD1.n5 1.7311
R1348 VDD1.n4 VDD1.t6 1.13258
R1349 VDD1.n4 VDD1.t2 1.13258
R1350 VDD1.n0 VDD1.t0 1.13258
R1351 VDD1.n0 VDD1.t3 1.13258
R1352 VDD1.n2 VDD1.t5 1.13258
R1353 VDD1.n2 VDD1.t1 1.13258
R1354 VDD1.n1 VDD1.t4 1.13258
R1355 VDD1.n1 VDD1.t7 1.13258
R1356 B.n1191 B.n1190 585
R1357 B.n1192 B.n1191 585
R1358 B.n441 B.n188 585
R1359 B.n440 B.n439 585
R1360 B.n438 B.n437 585
R1361 B.n436 B.n435 585
R1362 B.n434 B.n433 585
R1363 B.n432 B.n431 585
R1364 B.n430 B.n429 585
R1365 B.n428 B.n427 585
R1366 B.n426 B.n425 585
R1367 B.n424 B.n423 585
R1368 B.n422 B.n421 585
R1369 B.n420 B.n419 585
R1370 B.n418 B.n417 585
R1371 B.n416 B.n415 585
R1372 B.n414 B.n413 585
R1373 B.n412 B.n411 585
R1374 B.n410 B.n409 585
R1375 B.n408 B.n407 585
R1376 B.n406 B.n405 585
R1377 B.n404 B.n403 585
R1378 B.n402 B.n401 585
R1379 B.n400 B.n399 585
R1380 B.n398 B.n397 585
R1381 B.n396 B.n395 585
R1382 B.n394 B.n393 585
R1383 B.n392 B.n391 585
R1384 B.n390 B.n389 585
R1385 B.n388 B.n387 585
R1386 B.n386 B.n385 585
R1387 B.n384 B.n383 585
R1388 B.n382 B.n381 585
R1389 B.n380 B.n379 585
R1390 B.n378 B.n377 585
R1391 B.n376 B.n375 585
R1392 B.n374 B.n373 585
R1393 B.n372 B.n371 585
R1394 B.n370 B.n369 585
R1395 B.n368 B.n367 585
R1396 B.n366 B.n365 585
R1397 B.n364 B.n363 585
R1398 B.n362 B.n361 585
R1399 B.n360 B.n359 585
R1400 B.n358 B.n357 585
R1401 B.n356 B.n355 585
R1402 B.n354 B.n353 585
R1403 B.n352 B.n351 585
R1404 B.n350 B.n349 585
R1405 B.n348 B.n347 585
R1406 B.n346 B.n345 585
R1407 B.n344 B.n343 585
R1408 B.n342 B.n341 585
R1409 B.n340 B.n339 585
R1410 B.n338 B.n337 585
R1411 B.n336 B.n335 585
R1412 B.n334 B.n333 585
R1413 B.n332 B.n331 585
R1414 B.n330 B.n329 585
R1415 B.n327 B.n326 585
R1416 B.n325 B.n324 585
R1417 B.n323 B.n322 585
R1418 B.n321 B.n320 585
R1419 B.n319 B.n318 585
R1420 B.n317 B.n316 585
R1421 B.n315 B.n314 585
R1422 B.n313 B.n312 585
R1423 B.n311 B.n310 585
R1424 B.n309 B.n308 585
R1425 B.n307 B.n306 585
R1426 B.n305 B.n304 585
R1427 B.n303 B.n302 585
R1428 B.n301 B.n300 585
R1429 B.n299 B.n298 585
R1430 B.n297 B.n296 585
R1431 B.n295 B.n294 585
R1432 B.n293 B.n292 585
R1433 B.n291 B.n290 585
R1434 B.n289 B.n288 585
R1435 B.n287 B.n286 585
R1436 B.n285 B.n284 585
R1437 B.n283 B.n282 585
R1438 B.n281 B.n280 585
R1439 B.n279 B.n278 585
R1440 B.n277 B.n276 585
R1441 B.n275 B.n274 585
R1442 B.n273 B.n272 585
R1443 B.n271 B.n270 585
R1444 B.n269 B.n268 585
R1445 B.n267 B.n266 585
R1446 B.n265 B.n264 585
R1447 B.n263 B.n262 585
R1448 B.n261 B.n260 585
R1449 B.n259 B.n258 585
R1450 B.n257 B.n256 585
R1451 B.n255 B.n254 585
R1452 B.n253 B.n252 585
R1453 B.n251 B.n250 585
R1454 B.n249 B.n248 585
R1455 B.n247 B.n246 585
R1456 B.n245 B.n244 585
R1457 B.n243 B.n242 585
R1458 B.n241 B.n240 585
R1459 B.n239 B.n238 585
R1460 B.n237 B.n236 585
R1461 B.n235 B.n234 585
R1462 B.n233 B.n232 585
R1463 B.n231 B.n230 585
R1464 B.n229 B.n228 585
R1465 B.n227 B.n226 585
R1466 B.n225 B.n224 585
R1467 B.n223 B.n222 585
R1468 B.n221 B.n220 585
R1469 B.n219 B.n218 585
R1470 B.n217 B.n216 585
R1471 B.n215 B.n214 585
R1472 B.n213 B.n212 585
R1473 B.n211 B.n210 585
R1474 B.n209 B.n208 585
R1475 B.n207 B.n206 585
R1476 B.n205 B.n204 585
R1477 B.n203 B.n202 585
R1478 B.n201 B.n200 585
R1479 B.n199 B.n198 585
R1480 B.n197 B.n196 585
R1481 B.n195 B.n194 585
R1482 B.n1189 B.n125 585
R1483 B.n1193 B.n125 585
R1484 B.n1188 B.n124 585
R1485 B.n1194 B.n124 585
R1486 B.n1187 B.n1186 585
R1487 B.n1186 B.n120 585
R1488 B.n1185 B.n119 585
R1489 B.n1200 B.n119 585
R1490 B.n1184 B.n118 585
R1491 B.n1201 B.n118 585
R1492 B.n1183 B.n117 585
R1493 B.n1202 B.n117 585
R1494 B.n1182 B.n1181 585
R1495 B.n1181 B.n113 585
R1496 B.n1180 B.n112 585
R1497 B.n1208 B.n112 585
R1498 B.n1179 B.n111 585
R1499 B.n1209 B.n111 585
R1500 B.n1178 B.n110 585
R1501 B.n1210 B.n110 585
R1502 B.n1177 B.n1176 585
R1503 B.n1176 B.n106 585
R1504 B.n1175 B.n105 585
R1505 B.n1216 B.n105 585
R1506 B.n1174 B.n104 585
R1507 B.n1217 B.n104 585
R1508 B.n1173 B.n103 585
R1509 B.n1218 B.n103 585
R1510 B.n1172 B.n1171 585
R1511 B.n1171 B.n99 585
R1512 B.n1170 B.n98 585
R1513 B.n1224 B.n98 585
R1514 B.n1169 B.n97 585
R1515 B.n1225 B.n97 585
R1516 B.n1168 B.n96 585
R1517 B.n1226 B.n96 585
R1518 B.n1167 B.n1166 585
R1519 B.n1166 B.n92 585
R1520 B.n1165 B.n91 585
R1521 B.n1232 B.n91 585
R1522 B.n1164 B.n90 585
R1523 B.n1233 B.n90 585
R1524 B.n1163 B.n89 585
R1525 B.n1234 B.n89 585
R1526 B.n1162 B.n1161 585
R1527 B.n1161 B.n85 585
R1528 B.n1160 B.n84 585
R1529 B.n1240 B.n84 585
R1530 B.n1159 B.n83 585
R1531 B.n1241 B.n83 585
R1532 B.n1158 B.n82 585
R1533 B.n1242 B.n82 585
R1534 B.n1157 B.n1156 585
R1535 B.n1156 B.n78 585
R1536 B.n1155 B.n77 585
R1537 B.n1248 B.n77 585
R1538 B.n1154 B.n76 585
R1539 B.n1249 B.n76 585
R1540 B.n1153 B.n75 585
R1541 B.n1250 B.n75 585
R1542 B.n1152 B.n1151 585
R1543 B.n1151 B.n71 585
R1544 B.n1150 B.n70 585
R1545 B.n1256 B.n70 585
R1546 B.n1149 B.n69 585
R1547 B.n1257 B.n69 585
R1548 B.n1148 B.n68 585
R1549 B.n1258 B.n68 585
R1550 B.n1147 B.n1146 585
R1551 B.n1146 B.n64 585
R1552 B.n1145 B.n63 585
R1553 B.n1264 B.n63 585
R1554 B.n1144 B.n62 585
R1555 B.n1265 B.n62 585
R1556 B.n1143 B.n61 585
R1557 B.n1266 B.n61 585
R1558 B.n1142 B.n1141 585
R1559 B.n1141 B.n57 585
R1560 B.n1140 B.n56 585
R1561 B.n1272 B.n56 585
R1562 B.n1139 B.n55 585
R1563 B.n1273 B.n55 585
R1564 B.n1138 B.n54 585
R1565 B.n1274 B.n54 585
R1566 B.n1137 B.n1136 585
R1567 B.n1136 B.n50 585
R1568 B.n1135 B.n49 585
R1569 B.n1280 B.n49 585
R1570 B.n1134 B.n48 585
R1571 B.n1281 B.n48 585
R1572 B.n1133 B.n47 585
R1573 B.n1282 B.n47 585
R1574 B.n1132 B.n1131 585
R1575 B.n1131 B.n43 585
R1576 B.n1130 B.n42 585
R1577 B.n1288 B.n42 585
R1578 B.n1129 B.n41 585
R1579 B.n1289 B.n41 585
R1580 B.n1128 B.n40 585
R1581 B.n1290 B.n40 585
R1582 B.n1127 B.n1126 585
R1583 B.n1126 B.n36 585
R1584 B.n1125 B.n35 585
R1585 B.n1296 B.n35 585
R1586 B.n1124 B.n34 585
R1587 B.n1297 B.n34 585
R1588 B.n1123 B.n33 585
R1589 B.n1298 B.n33 585
R1590 B.n1122 B.n1121 585
R1591 B.n1121 B.n29 585
R1592 B.n1120 B.n28 585
R1593 B.n1304 B.n28 585
R1594 B.n1119 B.n27 585
R1595 B.n1305 B.n27 585
R1596 B.n1118 B.n26 585
R1597 B.n1306 B.n26 585
R1598 B.n1117 B.n1116 585
R1599 B.n1116 B.n22 585
R1600 B.n1115 B.n21 585
R1601 B.n1312 B.n21 585
R1602 B.n1114 B.n20 585
R1603 B.n1313 B.n20 585
R1604 B.n1113 B.n19 585
R1605 B.n1314 B.n19 585
R1606 B.n1112 B.n1111 585
R1607 B.n1111 B.n15 585
R1608 B.n1110 B.n14 585
R1609 B.n1320 B.n14 585
R1610 B.n1109 B.n13 585
R1611 B.n1321 B.n13 585
R1612 B.n1108 B.n12 585
R1613 B.n1322 B.n12 585
R1614 B.n1107 B.n1106 585
R1615 B.n1106 B.n8 585
R1616 B.n1105 B.n7 585
R1617 B.n1328 B.n7 585
R1618 B.n1104 B.n6 585
R1619 B.n1329 B.n6 585
R1620 B.n1103 B.n5 585
R1621 B.n1330 B.n5 585
R1622 B.n1102 B.n1101 585
R1623 B.n1101 B.n4 585
R1624 B.n1100 B.n442 585
R1625 B.n1100 B.n1099 585
R1626 B.n1090 B.n443 585
R1627 B.n444 B.n443 585
R1628 B.n1092 B.n1091 585
R1629 B.n1093 B.n1092 585
R1630 B.n1089 B.n449 585
R1631 B.n449 B.n448 585
R1632 B.n1088 B.n1087 585
R1633 B.n1087 B.n1086 585
R1634 B.n451 B.n450 585
R1635 B.n452 B.n451 585
R1636 B.n1079 B.n1078 585
R1637 B.n1080 B.n1079 585
R1638 B.n1077 B.n457 585
R1639 B.n457 B.n456 585
R1640 B.n1076 B.n1075 585
R1641 B.n1075 B.n1074 585
R1642 B.n459 B.n458 585
R1643 B.n460 B.n459 585
R1644 B.n1067 B.n1066 585
R1645 B.n1068 B.n1067 585
R1646 B.n1065 B.n465 585
R1647 B.n465 B.n464 585
R1648 B.n1064 B.n1063 585
R1649 B.n1063 B.n1062 585
R1650 B.n467 B.n466 585
R1651 B.n468 B.n467 585
R1652 B.n1055 B.n1054 585
R1653 B.n1056 B.n1055 585
R1654 B.n1053 B.n473 585
R1655 B.n473 B.n472 585
R1656 B.n1052 B.n1051 585
R1657 B.n1051 B.n1050 585
R1658 B.n475 B.n474 585
R1659 B.n476 B.n475 585
R1660 B.n1043 B.n1042 585
R1661 B.n1044 B.n1043 585
R1662 B.n1041 B.n481 585
R1663 B.n481 B.n480 585
R1664 B.n1040 B.n1039 585
R1665 B.n1039 B.n1038 585
R1666 B.n483 B.n482 585
R1667 B.n484 B.n483 585
R1668 B.n1031 B.n1030 585
R1669 B.n1032 B.n1031 585
R1670 B.n1029 B.n489 585
R1671 B.n489 B.n488 585
R1672 B.n1028 B.n1027 585
R1673 B.n1027 B.n1026 585
R1674 B.n491 B.n490 585
R1675 B.n492 B.n491 585
R1676 B.n1019 B.n1018 585
R1677 B.n1020 B.n1019 585
R1678 B.n1017 B.n497 585
R1679 B.n497 B.n496 585
R1680 B.n1016 B.n1015 585
R1681 B.n1015 B.n1014 585
R1682 B.n499 B.n498 585
R1683 B.n500 B.n499 585
R1684 B.n1007 B.n1006 585
R1685 B.n1008 B.n1007 585
R1686 B.n1005 B.n504 585
R1687 B.n508 B.n504 585
R1688 B.n1004 B.n1003 585
R1689 B.n1003 B.n1002 585
R1690 B.n506 B.n505 585
R1691 B.n507 B.n506 585
R1692 B.n995 B.n994 585
R1693 B.n996 B.n995 585
R1694 B.n993 B.n513 585
R1695 B.n513 B.n512 585
R1696 B.n992 B.n991 585
R1697 B.n991 B.n990 585
R1698 B.n515 B.n514 585
R1699 B.n516 B.n515 585
R1700 B.n983 B.n982 585
R1701 B.n984 B.n983 585
R1702 B.n981 B.n521 585
R1703 B.n521 B.n520 585
R1704 B.n980 B.n979 585
R1705 B.n979 B.n978 585
R1706 B.n523 B.n522 585
R1707 B.n524 B.n523 585
R1708 B.n971 B.n970 585
R1709 B.n972 B.n971 585
R1710 B.n969 B.n528 585
R1711 B.n532 B.n528 585
R1712 B.n968 B.n967 585
R1713 B.n967 B.n966 585
R1714 B.n530 B.n529 585
R1715 B.n531 B.n530 585
R1716 B.n959 B.n958 585
R1717 B.n960 B.n959 585
R1718 B.n957 B.n537 585
R1719 B.n537 B.n536 585
R1720 B.n956 B.n955 585
R1721 B.n955 B.n954 585
R1722 B.n539 B.n538 585
R1723 B.n540 B.n539 585
R1724 B.n947 B.n946 585
R1725 B.n948 B.n947 585
R1726 B.n945 B.n545 585
R1727 B.n545 B.n544 585
R1728 B.n944 B.n943 585
R1729 B.n943 B.n942 585
R1730 B.n547 B.n546 585
R1731 B.n548 B.n547 585
R1732 B.n935 B.n934 585
R1733 B.n936 B.n935 585
R1734 B.n933 B.n553 585
R1735 B.n553 B.n552 585
R1736 B.n932 B.n931 585
R1737 B.n931 B.n930 585
R1738 B.n555 B.n554 585
R1739 B.n556 B.n555 585
R1740 B.n923 B.n922 585
R1741 B.n924 B.n923 585
R1742 B.n921 B.n561 585
R1743 B.n561 B.n560 585
R1744 B.n920 B.n919 585
R1745 B.n919 B.n918 585
R1746 B.n563 B.n562 585
R1747 B.n564 B.n563 585
R1748 B.n911 B.n910 585
R1749 B.n912 B.n911 585
R1750 B.n909 B.n569 585
R1751 B.n569 B.n568 585
R1752 B.n908 B.n907 585
R1753 B.n907 B.n906 585
R1754 B.n571 B.n570 585
R1755 B.n572 B.n571 585
R1756 B.n899 B.n898 585
R1757 B.n900 B.n899 585
R1758 B.n897 B.n577 585
R1759 B.n577 B.n576 585
R1760 B.n891 B.n890 585
R1761 B.n889 B.n641 585
R1762 B.n888 B.n640 585
R1763 B.n893 B.n640 585
R1764 B.n887 B.n886 585
R1765 B.n885 B.n884 585
R1766 B.n883 B.n882 585
R1767 B.n881 B.n880 585
R1768 B.n879 B.n878 585
R1769 B.n877 B.n876 585
R1770 B.n875 B.n874 585
R1771 B.n873 B.n872 585
R1772 B.n871 B.n870 585
R1773 B.n869 B.n868 585
R1774 B.n867 B.n866 585
R1775 B.n865 B.n864 585
R1776 B.n863 B.n862 585
R1777 B.n861 B.n860 585
R1778 B.n859 B.n858 585
R1779 B.n857 B.n856 585
R1780 B.n855 B.n854 585
R1781 B.n853 B.n852 585
R1782 B.n851 B.n850 585
R1783 B.n849 B.n848 585
R1784 B.n847 B.n846 585
R1785 B.n845 B.n844 585
R1786 B.n843 B.n842 585
R1787 B.n841 B.n840 585
R1788 B.n839 B.n838 585
R1789 B.n837 B.n836 585
R1790 B.n835 B.n834 585
R1791 B.n833 B.n832 585
R1792 B.n831 B.n830 585
R1793 B.n829 B.n828 585
R1794 B.n827 B.n826 585
R1795 B.n825 B.n824 585
R1796 B.n823 B.n822 585
R1797 B.n821 B.n820 585
R1798 B.n819 B.n818 585
R1799 B.n817 B.n816 585
R1800 B.n815 B.n814 585
R1801 B.n813 B.n812 585
R1802 B.n811 B.n810 585
R1803 B.n809 B.n808 585
R1804 B.n807 B.n806 585
R1805 B.n805 B.n804 585
R1806 B.n803 B.n802 585
R1807 B.n801 B.n800 585
R1808 B.n799 B.n798 585
R1809 B.n797 B.n796 585
R1810 B.n795 B.n794 585
R1811 B.n793 B.n792 585
R1812 B.n791 B.n790 585
R1813 B.n789 B.n788 585
R1814 B.n787 B.n786 585
R1815 B.n785 B.n784 585
R1816 B.n783 B.n782 585
R1817 B.n781 B.n780 585
R1818 B.n779 B.n778 585
R1819 B.n776 B.n775 585
R1820 B.n774 B.n773 585
R1821 B.n772 B.n771 585
R1822 B.n770 B.n769 585
R1823 B.n768 B.n767 585
R1824 B.n766 B.n765 585
R1825 B.n764 B.n763 585
R1826 B.n762 B.n761 585
R1827 B.n760 B.n759 585
R1828 B.n758 B.n757 585
R1829 B.n756 B.n755 585
R1830 B.n754 B.n753 585
R1831 B.n752 B.n751 585
R1832 B.n750 B.n749 585
R1833 B.n748 B.n747 585
R1834 B.n746 B.n745 585
R1835 B.n744 B.n743 585
R1836 B.n742 B.n741 585
R1837 B.n740 B.n739 585
R1838 B.n738 B.n737 585
R1839 B.n736 B.n735 585
R1840 B.n734 B.n733 585
R1841 B.n732 B.n731 585
R1842 B.n730 B.n729 585
R1843 B.n728 B.n727 585
R1844 B.n726 B.n725 585
R1845 B.n724 B.n723 585
R1846 B.n722 B.n721 585
R1847 B.n720 B.n719 585
R1848 B.n718 B.n717 585
R1849 B.n716 B.n715 585
R1850 B.n714 B.n713 585
R1851 B.n712 B.n711 585
R1852 B.n710 B.n709 585
R1853 B.n708 B.n707 585
R1854 B.n706 B.n705 585
R1855 B.n704 B.n703 585
R1856 B.n702 B.n701 585
R1857 B.n700 B.n699 585
R1858 B.n698 B.n697 585
R1859 B.n696 B.n695 585
R1860 B.n694 B.n693 585
R1861 B.n692 B.n691 585
R1862 B.n690 B.n689 585
R1863 B.n688 B.n687 585
R1864 B.n686 B.n685 585
R1865 B.n684 B.n683 585
R1866 B.n682 B.n681 585
R1867 B.n680 B.n679 585
R1868 B.n678 B.n677 585
R1869 B.n676 B.n675 585
R1870 B.n674 B.n673 585
R1871 B.n672 B.n671 585
R1872 B.n670 B.n669 585
R1873 B.n668 B.n667 585
R1874 B.n666 B.n665 585
R1875 B.n664 B.n663 585
R1876 B.n662 B.n661 585
R1877 B.n660 B.n659 585
R1878 B.n658 B.n657 585
R1879 B.n656 B.n655 585
R1880 B.n654 B.n653 585
R1881 B.n652 B.n651 585
R1882 B.n650 B.n649 585
R1883 B.n648 B.n647 585
R1884 B.n579 B.n578 585
R1885 B.n896 B.n895 585
R1886 B.n575 B.n574 585
R1887 B.n576 B.n575 585
R1888 B.n902 B.n901 585
R1889 B.n901 B.n900 585
R1890 B.n903 B.n573 585
R1891 B.n573 B.n572 585
R1892 B.n905 B.n904 585
R1893 B.n906 B.n905 585
R1894 B.n567 B.n566 585
R1895 B.n568 B.n567 585
R1896 B.n914 B.n913 585
R1897 B.n913 B.n912 585
R1898 B.n915 B.n565 585
R1899 B.n565 B.n564 585
R1900 B.n917 B.n916 585
R1901 B.n918 B.n917 585
R1902 B.n559 B.n558 585
R1903 B.n560 B.n559 585
R1904 B.n926 B.n925 585
R1905 B.n925 B.n924 585
R1906 B.n927 B.n557 585
R1907 B.n557 B.n556 585
R1908 B.n929 B.n928 585
R1909 B.n930 B.n929 585
R1910 B.n551 B.n550 585
R1911 B.n552 B.n551 585
R1912 B.n938 B.n937 585
R1913 B.n937 B.n936 585
R1914 B.n939 B.n549 585
R1915 B.n549 B.n548 585
R1916 B.n941 B.n940 585
R1917 B.n942 B.n941 585
R1918 B.n543 B.n542 585
R1919 B.n544 B.n543 585
R1920 B.n950 B.n949 585
R1921 B.n949 B.n948 585
R1922 B.n951 B.n541 585
R1923 B.n541 B.n540 585
R1924 B.n953 B.n952 585
R1925 B.n954 B.n953 585
R1926 B.n535 B.n534 585
R1927 B.n536 B.n535 585
R1928 B.n962 B.n961 585
R1929 B.n961 B.n960 585
R1930 B.n963 B.n533 585
R1931 B.n533 B.n531 585
R1932 B.n965 B.n964 585
R1933 B.n966 B.n965 585
R1934 B.n527 B.n526 585
R1935 B.n532 B.n527 585
R1936 B.n974 B.n973 585
R1937 B.n973 B.n972 585
R1938 B.n975 B.n525 585
R1939 B.n525 B.n524 585
R1940 B.n977 B.n976 585
R1941 B.n978 B.n977 585
R1942 B.n519 B.n518 585
R1943 B.n520 B.n519 585
R1944 B.n986 B.n985 585
R1945 B.n985 B.n984 585
R1946 B.n987 B.n517 585
R1947 B.n517 B.n516 585
R1948 B.n989 B.n988 585
R1949 B.n990 B.n989 585
R1950 B.n511 B.n510 585
R1951 B.n512 B.n511 585
R1952 B.n998 B.n997 585
R1953 B.n997 B.n996 585
R1954 B.n999 B.n509 585
R1955 B.n509 B.n507 585
R1956 B.n1001 B.n1000 585
R1957 B.n1002 B.n1001 585
R1958 B.n503 B.n502 585
R1959 B.n508 B.n503 585
R1960 B.n1010 B.n1009 585
R1961 B.n1009 B.n1008 585
R1962 B.n1011 B.n501 585
R1963 B.n501 B.n500 585
R1964 B.n1013 B.n1012 585
R1965 B.n1014 B.n1013 585
R1966 B.n495 B.n494 585
R1967 B.n496 B.n495 585
R1968 B.n1022 B.n1021 585
R1969 B.n1021 B.n1020 585
R1970 B.n1023 B.n493 585
R1971 B.n493 B.n492 585
R1972 B.n1025 B.n1024 585
R1973 B.n1026 B.n1025 585
R1974 B.n487 B.n486 585
R1975 B.n488 B.n487 585
R1976 B.n1034 B.n1033 585
R1977 B.n1033 B.n1032 585
R1978 B.n1035 B.n485 585
R1979 B.n485 B.n484 585
R1980 B.n1037 B.n1036 585
R1981 B.n1038 B.n1037 585
R1982 B.n479 B.n478 585
R1983 B.n480 B.n479 585
R1984 B.n1046 B.n1045 585
R1985 B.n1045 B.n1044 585
R1986 B.n1047 B.n477 585
R1987 B.n477 B.n476 585
R1988 B.n1049 B.n1048 585
R1989 B.n1050 B.n1049 585
R1990 B.n471 B.n470 585
R1991 B.n472 B.n471 585
R1992 B.n1058 B.n1057 585
R1993 B.n1057 B.n1056 585
R1994 B.n1059 B.n469 585
R1995 B.n469 B.n468 585
R1996 B.n1061 B.n1060 585
R1997 B.n1062 B.n1061 585
R1998 B.n463 B.n462 585
R1999 B.n464 B.n463 585
R2000 B.n1070 B.n1069 585
R2001 B.n1069 B.n1068 585
R2002 B.n1071 B.n461 585
R2003 B.n461 B.n460 585
R2004 B.n1073 B.n1072 585
R2005 B.n1074 B.n1073 585
R2006 B.n455 B.n454 585
R2007 B.n456 B.n455 585
R2008 B.n1082 B.n1081 585
R2009 B.n1081 B.n1080 585
R2010 B.n1083 B.n453 585
R2011 B.n453 B.n452 585
R2012 B.n1085 B.n1084 585
R2013 B.n1086 B.n1085 585
R2014 B.n447 B.n446 585
R2015 B.n448 B.n447 585
R2016 B.n1095 B.n1094 585
R2017 B.n1094 B.n1093 585
R2018 B.n1096 B.n445 585
R2019 B.n445 B.n444 585
R2020 B.n1098 B.n1097 585
R2021 B.n1099 B.n1098 585
R2022 B.n2 B.n0 585
R2023 B.n4 B.n2 585
R2024 B.n3 B.n1 585
R2025 B.n1329 B.n3 585
R2026 B.n1327 B.n1326 585
R2027 B.n1328 B.n1327 585
R2028 B.n1325 B.n9 585
R2029 B.n9 B.n8 585
R2030 B.n1324 B.n1323 585
R2031 B.n1323 B.n1322 585
R2032 B.n11 B.n10 585
R2033 B.n1321 B.n11 585
R2034 B.n1319 B.n1318 585
R2035 B.n1320 B.n1319 585
R2036 B.n1317 B.n16 585
R2037 B.n16 B.n15 585
R2038 B.n1316 B.n1315 585
R2039 B.n1315 B.n1314 585
R2040 B.n18 B.n17 585
R2041 B.n1313 B.n18 585
R2042 B.n1311 B.n1310 585
R2043 B.n1312 B.n1311 585
R2044 B.n1309 B.n23 585
R2045 B.n23 B.n22 585
R2046 B.n1308 B.n1307 585
R2047 B.n1307 B.n1306 585
R2048 B.n25 B.n24 585
R2049 B.n1305 B.n25 585
R2050 B.n1303 B.n1302 585
R2051 B.n1304 B.n1303 585
R2052 B.n1301 B.n30 585
R2053 B.n30 B.n29 585
R2054 B.n1300 B.n1299 585
R2055 B.n1299 B.n1298 585
R2056 B.n32 B.n31 585
R2057 B.n1297 B.n32 585
R2058 B.n1295 B.n1294 585
R2059 B.n1296 B.n1295 585
R2060 B.n1293 B.n37 585
R2061 B.n37 B.n36 585
R2062 B.n1292 B.n1291 585
R2063 B.n1291 B.n1290 585
R2064 B.n39 B.n38 585
R2065 B.n1289 B.n39 585
R2066 B.n1287 B.n1286 585
R2067 B.n1288 B.n1287 585
R2068 B.n1285 B.n44 585
R2069 B.n44 B.n43 585
R2070 B.n1284 B.n1283 585
R2071 B.n1283 B.n1282 585
R2072 B.n46 B.n45 585
R2073 B.n1281 B.n46 585
R2074 B.n1279 B.n1278 585
R2075 B.n1280 B.n1279 585
R2076 B.n1277 B.n51 585
R2077 B.n51 B.n50 585
R2078 B.n1276 B.n1275 585
R2079 B.n1275 B.n1274 585
R2080 B.n53 B.n52 585
R2081 B.n1273 B.n53 585
R2082 B.n1271 B.n1270 585
R2083 B.n1272 B.n1271 585
R2084 B.n1269 B.n58 585
R2085 B.n58 B.n57 585
R2086 B.n1268 B.n1267 585
R2087 B.n1267 B.n1266 585
R2088 B.n60 B.n59 585
R2089 B.n1265 B.n60 585
R2090 B.n1263 B.n1262 585
R2091 B.n1264 B.n1263 585
R2092 B.n1261 B.n65 585
R2093 B.n65 B.n64 585
R2094 B.n1260 B.n1259 585
R2095 B.n1259 B.n1258 585
R2096 B.n67 B.n66 585
R2097 B.n1257 B.n67 585
R2098 B.n1255 B.n1254 585
R2099 B.n1256 B.n1255 585
R2100 B.n1253 B.n72 585
R2101 B.n72 B.n71 585
R2102 B.n1252 B.n1251 585
R2103 B.n1251 B.n1250 585
R2104 B.n74 B.n73 585
R2105 B.n1249 B.n74 585
R2106 B.n1247 B.n1246 585
R2107 B.n1248 B.n1247 585
R2108 B.n1245 B.n79 585
R2109 B.n79 B.n78 585
R2110 B.n1244 B.n1243 585
R2111 B.n1243 B.n1242 585
R2112 B.n81 B.n80 585
R2113 B.n1241 B.n81 585
R2114 B.n1239 B.n1238 585
R2115 B.n1240 B.n1239 585
R2116 B.n1237 B.n86 585
R2117 B.n86 B.n85 585
R2118 B.n1236 B.n1235 585
R2119 B.n1235 B.n1234 585
R2120 B.n88 B.n87 585
R2121 B.n1233 B.n88 585
R2122 B.n1231 B.n1230 585
R2123 B.n1232 B.n1231 585
R2124 B.n1229 B.n93 585
R2125 B.n93 B.n92 585
R2126 B.n1228 B.n1227 585
R2127 B.n1227 B.n1226 585
R2128 B.n95 B.n94 585
R2129 B.n1225 B.n95 585
R2130 B.n1223 B.n1222 585
R2131 B.n1224 B.n1223 585
R2132 B.n1221 B.n100 585
R2133 B.n100 B.n99 585
R2134 B.n1220 B.n1219 585
R2135 B.n1219 B.n1218 585
R2136 B.n102 B.n101 585
R2137 B.n1217 B.n102 585
R2138 B.n1215 B.n1214 585
R2139 B.n1216 B.n1215 585
R2140 B.n1213 B.n107 585
R2141 B.n107 B.n106 585
R2142 B.n1212 B.n1211 585
R2143 B.n1211 B.n1210 585
R2144 B.n109 B.n108 585
R2145 B.n1209 B.n109 585
R2146 B.n1207 B.n1206 585
R2147 B.n1208 B.n1207 585
R2148 B.n1205 B.n114 585
R2149 B.n114 B.n113 585
R2150 B.n1204 B.n1203 585
R2151 B.n1203 B.n1202 585
R2152 B.n116 B.n115 585
R2153 B.n1201 B.n116 585
R2154 B.n1199 B.n1198 585
R2155 B.n1200 B.n1199 585
R2156 B.n1197 B.n121 585
R2157 B.n121 B.n120 585
R2158 B.n1196 B.n1195 585
R2159 B.n1195 B.n1194 585
R2160 B.n123 B.n122 585
R2161 B.n1193 B.n123 585
R2162 B.n1332 B.n1331 585
R2163 B.n1331 B.n1330 585
R2164 B.n891 B.n575 530.939
R2165 B.n194 B.n123 530.939
R2166 B.n895 B.n577 530.939
R2167 B.n1191 B.n125 530.939
R2168 B.n644 B.t11 457.161
R2169 B.n642 B.t14 457.161
R2170 B.n191 B.t20 457.161
R2171 B.n189 B.t17 457.161
R2172 B.n645 B.t10 376.678
R2173 B.n190 B.t18 376.678
R2174 B.n643 B.t13 376.678
R2175 B.n192 B.t21 376.678
R2176 B.n644 B.t8 319.702
R2177 B.n642 B.t12 319.702
R2178 B.n191 B.t19 319.702
R2179 B.n189 B.t15 319.702
R2180 B.n1192 B.n187 256.663
R2181 B.n1192 B.n186 256.663
R2182 B.n1192 B.n185 256.663
R2183 B.n1192 B.n184 256.663
R2184 B.n1192 B.n183 256.663
R2185 B.n1192 B.n182 256.663
R2186 B.n1192 B.n181 256.663
R2187 B.n1192 B.n180 256.663
R2188 B.n1192 B.n179 256.663
R2189 B.n1192 B.n178 256.663
R2190 B.n1192 B.n177 256.663
R2191 B.n1192 B.n176 256.663
R2192 B.n1192 B.n175 256.663
R2193 B.n1192 B.n174 256.663
R2194 B.n1192 B.n173 256.663
R2195 B.n1192 B.n172 256.663
R2196 B.n1192 B.n171 256.663
R2197 B.n1192 B.n170 256.663
R2198 B.n1192 B.n169 256.663
R2199 B.n1192 B.n168 256.663
R2200 B.n1192 B.n167 256.663
R2201 B.n1192 B.n166 256.663
R2202 B.n1192 B.n165 256.663
R2203 B.n1192 B.n164 256.663
R2204 B.n1192 B.n163 256.663
R2205 B.n1192 B.n162 256.663
R2206 B.n1192 B.n161 256.663
R2207 B.n1192 B.n160 256.663
R2208 B.n1192 B.n159 256.663
R2209 B.n1192 B.n158 256.663
R2210 B.n1192 B.n157 256.663
R2211 B.n1192 B.n156 256.663
R2212 B.n1192 B.n155 256.663
R2213 B.n1192 B.n154 256.663
R2214 B.n1192 B.n153 256.663
R2215 B.n1192 B.n152 256.663
R2216 B.n1192 B.n151 256.663
R2217 B.n1192 B.n150 256.663
R2218 B.n1192 B.n149 256.663
R2219 B.n1192 B.n148 256.663
R2220 B.n1192 B.n147 256.663
R2221 B.n1192 B.n146 256.663
R2222 B.n1192 B.n145 256.663
R2223 B.n1192 B.n144 256.663
R2224 B.n1192 B.n143 256.663
R2225 B.n1192 B.n142 256.663
R2226 B.n1192 B.n141 256.663
R2227 B.n1192 B.n140 256.663
R2228 B.n1192 B.n139 256.663
R2229 B.n1192 B.n138 256.663
R2230 B.n1192 B.n137 256.663
R2231 B.n1192 B.n136 256.663
R2232 B.n1192 B.n135 256.663
R2233 B.n1192 B.n134 256.663
R2234 B.n1192 B.n133 256.663
R2235 B.n1192 B.n132 256.663
R2236 B.n1192 B.n131 256.663
R2237 B.n1192 B.n130 256.663
R2238 B.n1192 B.n129 256.663
R2239 B.n1192 B.n128 256.663
R2240 B.n1192 B.n127 256.663
R2241 B.n1192 B.n126 256.663
R2242 B.n893 B.n892 256.663
R2243 B.n893 B.n580 256.663
R2244 B.n893 B.n581 256.663
R2245 B.n893 B.n582 256.663
R2246 B.n893 B.n583 256.663
R2247 B.n893 B.n584 256.663
R2248 B.n893 B.n585 256.663
R2249 B.n893 B.n586 256.663
R2250 B.n893 B.n587 256.663
R2251 B.n893 B.n588 256.663
R2252 B.n893 B.n589 256.663
R2253 B.n893 B.n590 256.663
R2254 B.n893 B.n591 256.663
R2255 B.n893 B.n592 256.663
R2256 B.n893 B.n593 256.663
R2257 B.n893 B.n594 256.663
R2258 B.n893 B.n595 256.663
R2259 B.n893 B.n596 256.663
R2260 B.n893 B.n597 256.663
R2261 B.n893 B.n598 256.663
R2262 B.n893 B.n599 256.663
R2263 B.n893 B.n600 256.663
R2264 B.n893 B.n601 256.663
R2265 B.n893 B.n602 256.663
R2266 B.n893 B.n603 256.663
R2267 B.n893 B.n604 256.663
R2268 B.n893 B.n605 256.663
R2269 B.n893 B.n606 256.663
R2270 B.n893 B.n607 256.663
R2271 B.n893 B.n608 256.663
R2272 B.n893 B.n609 256.663
R2273 B.n893 B.n610 256.663
R2274 B.n893 B.n611 256.663
R2275 B.n893 B.n612 256.663
R2276 B.n893 B.n613 256.663
R2277 B.n893 B.n614 256.663
R2278 B.n893 B.n615 256.663
R2279 B.n893 B.n616 256.663
R2280 B.n893 B.n617 256.663
R2281 B.n893 B.n618 256.663
R2282 B.n893 B.n619 256.663
R2283 B.n893 B.n620 256.663
R2284 B.n893 B.n621 256.663
R2285 B.n893 B.n622 256.663
R2286 B.n893 B.n623 256.663
R2287 B.n893 B.n624 256.663
R2288 B.n893 B.n625 256.663
R2289 B.n893 B.n626 256.663
R2290 B.n893 B.n627 256.663
R2291 B.n893 B.n628 256.663
R2292 B.n893 B.n629 256.663
R2293 B.n893 B.n630 256.663
R2294 B.n893 B.n631 256.663
R2295 B.n893 B.n632 256.663
R2296 B.n893 B.n633 256.663
R2297 B.n893 B.n634 256.663
R2298 B.n893 B.n635 256.663
R2299 B.n893 B.n636 256.663
R2300 B.n893 B.n637 256.663
R2301 B.n893 B.n638 256.663
R2302 B.n893 B.n639 256.663
R2303 B.n894 B.n893 256.663
R2304 B.n901 B.n575 163.367
R2305 B.n901 B.n573 163.367
R2306 B.n905 B.n573 163.367
R2307 B.n905 B.n567 163.367
R2308 B.n913 B.n567 163.367
R2309 B.n913 B.n565 163.367
R2310 B.n917 B.n565 163.367
R2311 B.n917 B.n559 163.367
R2312 B.n925 B.n559 163.367
R2313 B.n925 B.n557 163.367
R2314 B.n929 B.n557 163.367
R2315 B.n929 B.n551 163.367
R2316 B.n937 B.n551 163.367
R2317 B.n937 B.n549 163.367
R2318 B.n941 B.n549 163.367
R2319 B.n941 B.n543 163.367
R2320 B.n949 B.n543 163.367
R2321 B.n949 B.n541 163.367
R2322 B.n953 B.n541 163.367
R2323 B.n953 B.n535 163.367
R2324 B.n961 B.n535 163.367
R2325 B.n961 B.n533 163.367
R2326 B.n965 B.n533 163.367
R2327 B.n965 B.n527 163.367
R2328 B.n973 B.n527 163.367
R2329 B.n973 B.n525 163.367
R2330 B.n977 B.n525 163.367
R2331 B.n977 B.n519 163.367
R2332 B.n985 B.n519 163.367
R2333 B.n985 B.n517 163.367
R2334 B.n989 B.n517 163.367
R2335 B.n989 B.n511 163.367
R2336 B.n997 B.n511 163.367
R2337 B.n997 B.n509 163.367
R2338 B.n1001 B.n509 163.367
R2339 B.n1001 B.n503 163.367
R2340 B.n1009 B.n503 163.367
R2341 B.n1009 B.n501 163.367
R2342 B.n1013 B.n501 163.367
R2343 B.n1013 B.n495 163.367
R2344 B.n1021 B.n495 163.367
R2345 B.n1021 B.n493 163.367
R2346 B.n1025 B.n493 163.367
R2347 B.n1025 B.n487 163.367
R2348 B.n1033 B.n487 163.367
R2349 B.n1033 B.n485 163.367
R2350 B.n1037 B.n485 163.367
R2351 B.n1037 B.n479 163.367
R2352 B.n1045 B.n479 163.367
R2353 B.n1045 B.n477 163.367
R2354 B.n1049 B.n477 163.367
R2355 B.n1049 B.n471 163.367
R2356 B.n1057 B.n471 163.367
R2357 B.n1057 B.n469 163.367
R2358 B.n1061 B.n469 163.367
R2359 B.n1061 B.n463 163.367
R2360 B.n1069 B.n463 163.367
R2361 B.n1069 B.n461 163.367
R2362 B.n1073 B.n461 163.367
R2363 B.n1073 B.n455 163.367
R2364 B.n1081 B.n455 163.367
R2365 B.n1081 B.n453 163.367
R2366 B.n1085 B.n453 163.367
R2367 B.n1085 B.n447 163.367
R2368 B.n1094 B.n447 163.367
R2369 B.n1094 B.n445 163.367
R2370 B.n1098 B.n445 163.367
R2371 B.n1098 B.n2 163.367
R2372 B.n1331 B.n2 163.367
R2373 B.n1331 B.n3 163.367
R2374 B.n1327 B.n3 163.367
R2375 B.n1327 B.n9 163.367
R2376 B.n1323 B.n9 163.367
R2377 B.n1323 B.n11 163.367
R2378 B.n1319 B.n11 163.367
R2379 B.n1319 B.n16 163.367
R2380 B.n1315 B.n16 163.367
R2381 B.n1315 B.n18 163.367
R2382 B.n1311 B.n18 163.367
R2383 B.n1311 B.n23 163.367
R2384 B.n1307 B.n23 163.367
R2385 B.n1307 B.n25 163.367
R2386 B.n1303 B.n25 163.367
R2387 B.n1303 B.n30 163.367
R2388 B.n1299 B.n30 163.367
R2389 B.n1299 B.n32 163.367
R2390 B.n1295 B.n32 163.367
R2391 B.n1295 B.n37 163.367
R2392 B.n1291 B.n37 163.367
R2393 B.n1291 B.n39 163.367
R2394 B.n1287 B.n39 163.367
R2395 B.n1287 B.n44 163.367
R2396 B.n1283 B.n44 163.367
R2397 B.n1283 B.n46 163.367
R2398 B.n1279 B.n46 163.367
R2399 B.n1279 B.n51 163.367
R2400 B.n1275 B.n51 163.367
R2401 B.n1275 B.n53 163.367
R2402 B.n1271 B.n53 163.367
R2403 B.n1271 B.n58 163.367
R2404 B.n1267 B.n58 163.367
R2405 B.n1267 B.n60 163.367
R2406 B.n1263 B.n60 163.367
R2407 B.n1263 B.n65 163.367
R2408 B.n1259 B.n65 163.367
R2409 B.n1259 B.n67 163.367
R2410 B.n1255 B.n67 163.367
R2411 B.n1255 B.n72 163.367
R2412 B.n1251 B.n72 163.367
R2413 B.n1251 B.n74 163.367
R2414 B.n1247 B.n74 163.367
R2415 B.n1247 B.n79 163.367
R2416 B.n1243 B.n79 163.367
R2417 B.n1243 B.n81 163.367
R2418 B.n1239 B.n81 163.367
R2419 B.n1239 B.n86 163.367
R2420 B.n1235 B.n86 163.367
R2421 B.n1235 B.n88 163.367
R2422 B.n1231 B.n88 163.367
R2423 B.n1231 B.n93 163.367
R2424 B.n1227 B.n93 163.367
R2425 B.n1227 B.n95 163.367
R2426 B.n1223 B.n95 163.367
R2427 B.n1223 B.n100 163.367
R2428 B.n1219 B.n100 163.367
R2429 B.n1219 B.n102 163.367
R2430 B.n1215 B.n102 163.367
R2431 B.n1215 B.n107 163.367
R2432 B.n1211 B.n107 163.367
R2433 B.n1211 B.n109 163.367
R2434 B.n1207 B.n109 163.367
R2435 B.n1207 B.n114 163.367
R2436 B.n1203 B.n114 163.367
R2437 B.n1203 B.n116 163.367
R2438 B.n1199 B.n116 163.367
R2439 B.n1199 B.n121 163.367
R2440 B.n1195 B.n121 163.367
R2441 B.n1195 B.n123 163.367
R2442 B.n641 B.n640 163.367
R2443 B.n886 B.n640 163.367
R2444 B.n884 B.n883 163.367
R2445 B.n880 B.n879 163.367
R2446 B.n876 B.n875 163.367
R2447 B.n872 B.n871 163.367
R2448 B.n868 B.n867 163.367
R2449 B.n864 B.n863 163.367
R2450 B.n860 B.n859 163.367
R2451 B.n856 B.n855 163.367
R2452 B.n852 B.n851 163.367
R2453 B.n848 B.n847 163.367
R2454 B.n844 B.n843 163.367
R2455 B.n840 B.n839 163.367
R2456 B.n836 B.n835 163.367
R2457 B.n832 B.n831 163.367
R2458 B.n828 B.n827 163.367
R2459 B.n824 B.n823 163.367
R2460 B.n820 B.n819 163.367
R2461 B.n816 B.n815 163.367
R2462 B.n812 B.n811 163.367
R2463 B.n808 B.n807 163.367
R2464 B.n804 B.n803 163.367
R2465 B.n800 B.n799 163.367
R2466 B.n796 B.n795 163.367
R2467 B.n792 B.n791 163.367
R2468 B.n788 B.n787 163.367
R2469 B.n784 B.n783 163.367
R2470 B.n780 B.n779 163.367
R2471 B.n775 B.n774 163.367
R2472 B.n771 B.n770 163.367
R2473 B.n767 B.n766 163.367
R2474 B.n763 B.n762 163.367
R2475 B.n759 B.n758 163.367
R2476 B.n755 B.n754 163.367
R2477 B.n751 B.n750 163.367
R2478 B.n747 B.n746 163.367
R2479 B.n743 B.n742 163.367
R2480 B.n739 B.n738 163.367
R2481 B.n735 B.n734 163.367
R2482 B.n731 B.n730 163.367
R2483 B.n727 B.n726 163.367
R2484 B.n723 B.n722 163.367
R2485 B.n719 B.n718 163.367
R2486 B.n715 B.n714 163.367
R2487 B.n711 B.n710 163.367
R2488 B.n707 B.n706 163.367
R2489 B.n703 B.n702 163.367
R2490 B.n699 B.n698 163.367
R2491 B.n695 B.n694 163.367
R2492 B.n691 B.n690 163.367
R2493 B.n687 B.n686 163.367
R2494 B.n683 B.n682 163.367
R2495 B.n679 B.n678 163.367
R2496 B.n675 B.n674 163.367
R2497 B.n671 B.n670 163.367
R2498 B.n667 B.n666 163.367
R2499 B.n663 B.n662 163.367
R2500 B.n659 B.n658 163.367
R2501 B.n655 B.n654 163.367
R2502 B.n651 B.n650 163.367
R2503 B.n647 B.n579 163.367
R2504 B.n899 B.n577 163.367
R2505 B.n899 B.n571 163.367
R2506 B.n907 B.n571 163.367
R2507 B.n907 B.n569 163.367
R2508 B.n911 B.n569 163.367
R2509 B.n911 B.n563 163.367
R2510 B.n919 B.n563 163.367
R2511 B.n919 B.n561 163.367
R2512 B.n923 B.n561 163.367
R2513 B.n923 B.n555 163.367
R2514 B.n931 B.n555 163.367
R2515 B.n931 B.n553 163.367
R2516 B.n935 B.n553 163.367
R2517 B.n935 B.n547 163.367
R2518 B.n943 B.n547 163.367
R2519 B.n943 B.n545 163.367
R2520 B.n947 B.n545 163.367
R2521 B.n947 B.n539 163.367
R2522 B.n955 B.n539 163.367
R2523 B.n955 B.n537 163.367
R2524 B.n959 B.n537 163.367
R2525 B.n959 B.n530 163.367
R2526 B.n967 B.n530 163.367
R2527 B.n967 B.n528 163.367
R2528 B.n971 B.n528 163.367
R2529 B.n971 B.n523 163.367
R2530 B.n979 B.n523 163.367
R2531 B.n979 B.n521 163.367
R2532 B.n983 B.n521 163.367
R2533 B.n983 B.n515 163.367
R2534 B.n991 B.n515 163.367
R2535 B.n991 B.n513 163.367
R2536 B.n995 B.n513 163.367
R2537 B.n995 B.n506 163.367
R2538 B.n1003 B.n506 163.367
R2539 B.n1003 B.n504 163.367
R2540 B.n1007 B.n504 163.367
R2541 B.n1007 B.n499 163.367
R2542 B.n1015 B.n499 163.367
R2543 B.n1015 B.n497 163.367
R2544 B.n1019 B.n497 163.367
R2545 B.n1019 B.n491 163.367
R2546 B.n1027 B.n491 163.367
R2547 B.n1027 B.n489 163.367
R2548 B.n1031 B.n489 163.367
R2549 B.n1031 B.n483 163.367
R2550 B.n1039 B.n483 163.367
R2551 B.n1039 B.n481 163.367
R2552 B.n1043 B.n481 163.367
R2553 B.n1043 B.n475 163.367
R2554 B.n1051 B.n475 163.367
R2555 B.n1051 B.n473 163.367
R2556 B.n1055 B.n473 163.367
R2557 B.n1055 B.n467 163.367
R2558 B.n1063 B.n467 163.367
R2559 B.n1063 B.n465 163.367
R2560 B.n1067 B.n465 163.367
R2561 B.n1067 B.n459 163.367
R2562 B.n1075 B.n459 163.367
R2563 B.n1075 B.n457 163.367
R2564 B.n1079 B.n457 163.367
R2565 B.n1079 B.n451 163.367
R2566 B.n1087 B.n451 163.367
R2567 B.n1087 B.n449 163.367
R2568 B.n1092 B.n449 163.367
R2569 B.n1092 B.n443 163.367
R2570 B.n1100 B.n443 163.367
R2571 B.n1101 B.n1100 163.367
R2572 B.n1101 B.n5 163.367
R2573 B.n6 B.n5 163.367
R2574 B.n7 B.n6 163.367
R2575 B.n1106 B.n7 163.367
R2576 B.n1106 B.n12 163.367
R2577 B.n13 B.n12 163.367
R2578 B.n14 B.n13 163.367
R2579 B.n1111 B.n14 163.367
R2580 B.n1111 B.n19 163.367
R2581 B.n20 B.n19 163.367
R2582 B.n21 B.n20 163.367
R2583 B.n1116 B.n21 163.367
R2584 B.n1116 B.n26 163.367
R2585 B.n27 B.n26 163.367
R2586 B.n28 B.n27 163.367
R2587 B.n1121 B.n28 163.367
R2588 B.n1121 B.n33 163.367
R2589 B.n34 B.n33 163.367
R2590 B.n35 B.n34 163.367
R2591 B.n1126 B.n35 163.367
R2592 B.n1126 B.n40 163.367
R2593 B.n41 B.n40 163.367
R2594 B.n42 B.n41 163.367
R2595 B.n1131 B.n42 163.367
R2596 B.n1131 B.n47 163.367
R2597 B.n48 B.n47 163.367
R2598 B.n49 B.n48 163.367
R2599 B.n1136 B.n49 163.367
R2600 B.n1136 B.n54 163.367
R2601 B.n55 B.n54 163.367
R2602 B.n56 B.n55 163.367
R2603 B.n1141 B.n56 163.367
R2604 B.n1141 B.n61 163.367
R2605 B.n62 B.n61 163.367
R2606 B.n63 B.n62 163.367
R2607 B.n1146 B.n63 163.367
R2608 B.n1146 B.n68 163.367
R2609 B.n69 B.n68 163.367
R2610 B.n70 B.n69 163.367
R2611 B.n1151 B.n70 163.367
R2612 B.n1151 B.n75 163.367
R2613 B.n76 B.n75 163.367
R2614 B.n77 B.n76 163.367
R2615 B.n1156 B.n77 163.367
R2616 B.n1156 B.n82 163.367
R2617 B.n83 B.n82 163.367
R2618 B.n84 B.n83 163.367
R2619 B.n1161 B.n84 163.367
R2620 B.n1161 B.n89 163.367
R2621 B.n90 B.n89 163.367
R2622 B.n91 B.n90 163.367
R2623 B.n1166 B.n91 163.367
R2624 B.n1166 B.n96 163.367
R2625 B.n97 B.n96 163.367
R2626 B.n98 B.n97 163.367
R2627 B.n1171 B.n98 163.367
R2628 B.n1171 B.n103 163.367
R2629 B.n104 B.n103 163.367
R2630 B.n105 B.n104 163.367
R2631 B.n1176 B.n105 163.367
R2632 B.n1176 B.n110 163.367
R2633 B.n111 B.n110 163.367
R2634 B.n112 B.n111 163.367
R2635 B.n1181 B.n112 163.367
R2636 B.n1181 B.n117 163.367
R2637 B.n118 B.n117 163.367
R2638 B.n119 B.n118 163.367
R2639 B.n1186 B.n119 163.367
R2640 B.n1186 B.n124 163.367
R2641 B.n125 B.n124 163.367
R2642 B.n198 B.n197 163.367
R2643 B.n202 B.n201 163.367
R2644 B.n206 B.n205 163.367
R2645 B.n210 B.n209 163.367
R2646 B.n214 B.n213 163.367
R2647 B.n218 B.n217 163.367
R2648 B.n222 B.n221 163.367
R2649 B.n226 B.n225 163.367
R2650 B.n230 B.n229 163.367
R2651 B.n234 B.n233 163.367
R2652 B.n238 B.n237 163.367
R2653 B.n242 B.n241 163.367
R2654 B.n246 B.n245 163.367
R2655 B.n250 B.n249 163.367
R2656 B.n254 B.n253 163.367
R2657 B.n258 B.n257 163.367
R2658 B.n262 B.n261 163.367
R2659 B.n266 B.n265 163.367
R2660 B.n270 B.n269 163.367
R2661 B.n274 B.n273 163.367
R2662 B.n278 B.n277 163.367
R2663 B.n282 B.n281 163.367
R2664 B.n286 B.n285 163.367
R2665 B.n290 B.n289 163.367
R2666 B.n294 B.n293 163.367
R2667 B.n298 B.n297 163.367
R2668 B.n302 B.n301 163.367
R2669 B.n306 B.n305 163.367
R2670 B.n310 B.n309 163.367
R2671 B.n314 B.n313 163.367
R2672 B.n318 B.n317 163.367
R2673 B.n322 B.n321 163.367
R2674 B.n326 B.n325 163.367
R2675 B.n331 B.n330 163.367
R2676 B.n335 B.n334 163.367
R2677 B.n339 B.n338 163.367
R2678 B.n343 B.n342 163.367
R2679 B.n347 B.n346 163.367
R2680 B.n351 B.n350 163.367
R2681 B.n355 B.n354 163.367
R2682 B.n359 B.n358 163.367
R2683 B.n363 B.n362 163.367
R2684 B.n367 B.n366 163.367
R2685 B.n371 B.n370 163.367
R2686 B.n375 B.n374 163.367
R2687 B.n379 B.n378 163.367
R2688 B.n383 B.n382 163.367
R2689 B.n387 B.n386 163.367
R2690 B.n391 B.n390 163.367
R2691 B.n395 B.n394 163.367
R2692 B.n399 B.n398 163.367
R2693 B.n403 B.n402 163.367
R2694 B.n407 B.n406 163.367
R2695 B.n411 B.n410 163.367
R2696 B.n415 B.n414 163.367
R2697 B.n419 B.n418 163.367
R2698 B.n423 B.n422 163.367
R2699 B.n427 B.n426 163.367
R2700 B.n431 B.n430 163.367
R2701 B.n435 B.n434 163.367
R2702 B.n439 B.n438 163.367
R2703 B.n1191 B.n188 163.367
R2704 B.n645 B.n644 80.4853
R2705 B.n643 B.n642 80.4853
R2706 B.n192 B.n191 80.4853
R2707 B.n190 B.n189 80.4853
R2708 B.n892 B.n891 71.676
R2709 B.n886 B.n580 71.676
R2710 B.n883 B.n581 71.676
R2711 B.n879 B.n582 71.676
R2712 B.n875 B.n583 71.676
R2713 B.n871 B.n584 71.676
R2714 B.n867 B.n585 71.676
R2715 B.n863 B.n586 71.676
R2716 B.n859 B.n587 71.676
R2717 B.n855 B.n588 71.676
R2718 B.n851 B.n589 71.676
R2719 B.n847 B.n590 71.676
R2720 B.n843 B.n591 71.676
R2721 B.n839 B.n592 71.676
R2722 B.n835 B.n593 71.676
R2723 B.n831 B.n594 71.676
R2724 B.n827 B.n595 71.676
R2725 B.n823 B.n596 71.676
R2726 B.n819 B.n597 71.676
R2727 B.n815 B.n598 71.676
R2728 B.n811 B.n599 71.676
R2729 B.n807 B.n600 71.676
R2730 B.n803 B.n601 71.676
R2731 B.n799 B.n602 71.676
R2732 B.n795 B.n603 71.676
R2733 B.n791 B.n604 71.676
R2734 B.n787 B.n605 71.676
R2735 B.n783 B.n606 71.676
R2736 B.n779 B.n607 71.676
R2737 B.n774 B.n608 71.676
R2738 B.n770 B.n609 71.676
R2739 B.n766 B.n610 71.676
R2740 B.n762 B.n611 71.676
R2741 B.n758 B.n612 71.676
R2742 B.n754 B.n613 71.676
R2743 B.n750 B.n614 71.676
R2744 B.n746 B.n615 71.676
R2745 B.n742 B.n616 71.676
R2746 B.n738 B.n617 71.676
R2747 B.n734 B.n618 71.676
R2748 B.n730 B.n619 71.676
R2749 B.n726 B.n620 71.676
R2750 B.n722 B.n621 71.676
R2751 B.n718 B.n622 71.676
R2752 B.n714 B.n623 71.676
R2753 B.n710 B.n624 71.676
R2754 B.n706 B.n625 71.676
R2755 B.n702 B.n626 71.676
R2756 B.n698 B.n627 71.676
R2757 B.n694 B.n628 71.676
R2758 B.n690 B.n629 71.676
R2759 B.n686 B.n630 71.676
R2760 B.n682 B.n631 71.676
R2761 B.n678 B.n632 71.676
R2762 B.n674 B.n633 71.676
R2763 B.n670 B.n634 71.676
R2764 B.n666 B.n635 71.676
R2765 B.n662 B.n636 71.676
R2766 B.n658 B.n637 71.676
R2767 B.n654 B.n638 71.676
R2768 B.n650 B.n639 71.676
R2769 B.n894 B.n579 71.676
R2770 B.n194 B.n126 71.676
R2771 B.n198 B.n127 71.676
R2772 B.n202 B.n128 71.676
R2773 B.n206 B.n129 71.676
R2774 B.n210 B.n130 71.676
R2775 B.n214 B.n131 71.676
R2776 B.n218 B.n132 71.676
R2777 B.n222 B.n133 71.676
R2778 B.n226 B.n134 71.676
R2779 B.n230 B.n135 71.676
R2780 B.n234 B.n136 71.676
R2781 B.n238 B.n137 71.676
R2782 B.n242 B.n138 71.676
R2783 B.n246 B.n139 71.676
R2784 B.n250 B.n140 71.676
R2785 B.n254 B.n141 71.676
R2786 B.n258 B.n142 71.676
R2787 B.n262 B.n143 71.676
R2788 B.n266 B.n144 71.676
R2789 B.n270 B.n145 71.676
R2790 B.n274 B.n146 71.676
R2791 B.n278 B.n147 71.676
R2792 B.n282 B.n148 71.676
R2793 B.n286 B.n149 71.676
R2794 B.n290 B.n150 71.676
R2795 B.n294 B.n151 71.676
R2796 B.n298 B.n152 71.676
R2797 B.n302 B.n153 71.676
R2798 B.n306 B.n154 71.676
R2799 B.n310 B.n155 71.676
R2800 B.n314 B.n156 71.676
R2801 B.n318 B.n157 71.676
R2802 B.n322 B.n158 71.676
R2803 B.n326 B.n159 71.676
R2804 B.n331 B.n160 71.676
R2805 B.n335 B.n161 71.676
R2806 B.n339 B.n162 71.676
R2807 B.n343 B.n163 71.676
R2808 B.n347 B.n164 71.676
R2809 B.n351 B.n165 71.676
R2810 B.n355 B.n166 71.676
R2811 B.n359 B.n167 71.676
R2812 B.n363 B.n168 71.676
R2813 B.n367 B.n169 71.676
R2814 B.n371 B.n170 71.676
R2815 B.n375 B.n171 71.676
R2816 B.n379 B.n172 71.676
R2817 B.n383 B.n173 71.676
R2818 B.n387 B.n174 71.676
R2819 B.n391 B.n175 71.676
R2820 B.n395 B.n176 71.676
R2821 B.n399 B.n177 71.676
R2822 B.n403 B.n178 71.676
R2823 B.n407 B.n179 71.676
R2824 B.n411 B.n180 71.676
R2825 B.n415 B.n181 71.676
R2826 B.n419 B.n182 71.676
R2827 B.n423 B.n183 71.676
R2828 B.n427 B.n184 71.676
R2829 B.n431 B.n185 71.676
R2830 B.n435 B.n186 71.676
R2831 B.n439 B.n187 71.676
R2832 B.n188 B.n187 71.676
R2833 B.n438 B.n186 71.676
R2834 B.n434 B.n185 71.676
R2835 B.n430 B.n184 71.676
R2836 B.n426 B.n183 71.676
R2837 B.n422 B.n182 71.676
R2838 B.n418 B.n181 71.676
R2839 B.n414 B.n180 71.676
R2840 B.n410 B.n179 71.676
R2841 B.n406 B.n178 71.676
R2842 B.n402 B.n177 71.676
R2843 B.n398 B.n176 71.676
R2844 B.n394 B.n175 71.676
R2845 B.n390 B.n174 71.676
R2846 B.n386 B.n173 71.676
R2847 B.n382 B.n172 71.676
R2848 B.n378 B.n171 71.676
R2849 B.n374 B.n170 71.676
R2850 B.n370 B.n169 71.676
R2851 B.n366 B.n168 71.676
R2852 B.n362 B.n167 71.676
R2853 B.n358 B.n166 71.676
R2854 B.n354 B.n165 71.676
R2855 B.n350 B.n164 71.676
R2856 B.n346 B.n163 71.676
R2857 B.n342 B.n162 71.676
R2858 B.n338 B.n161 71.676
R2859 B.n334 B.n160 71.676
R2860 B.n330 B.n159 71.676
R2861 B.n325 B.n158 71.676
R2862 B.n321 B.n157 71.676
R2863 B.n317 B.n156 71.676
R2864 B.n313 B.n155 71.676
R2865 B.n309 B.n154 71.676
R2866 B.n305 B.n153 71.676
R2867 B.n301 B.n152 71.676
R2868 B.n297 B.n151 71.676
R2869 B.n293 B.n150 71.676
R2870 B.n289 B.n149 71.676
R2871 B.n285 B.n148 71.676
R2872 B.n281 B.n147 71.676
R2873 B.n277 B.n146 71.676
R2874 B.n273 B.n145 71.676
R2875 B.n269 B.n144 71.676
R2876 B.n265 B.n143 71.676
R2877 B.n261 B.n142 71.676
R2878 B.n257 B.n141 71.676
R2879 B.n253 B.n140 71.676
R2880 B.n249 B.n139 71.676
R2881 B.n245 B.n138 71.676
R2882 B.n241 B.n137 71.676
R2883 B.n237 B.n136 71.676
R2884 B.n233 B.n135 71.676
R2885 B.n229 B.n134 71.676
R2886 B.n225 B.n133 71.676
R2887 B.n221 B.n132 71.676
R2888 B.n217 B.n131 71.676
R2889 B.n213 B.n130 71.676
R2890 B.n209 B.n129 71.676
R2891 B.n205 B.n128 71.676
R2892 B.n201 B.n127 71.676
R2893 B.n197 B.n126 71.676
R2894 B.n892 B.n641 71.676
R2895 B.n884 B.n580 71.676
R2896 B.n880 B.n581 71.676
R2897 B.n876 B.n582 71.676
R2898 B.n872 B.n583 71.676
R2899 B.n868 B.n584 71.676
R2900 B.n864 B.n585 71.676
R2901 B.n860 B.n586 71.676
R2902 B.n856 B.n587 71.676
R2903 B.n852 B.n588 71.676
R2904 B.n848 B.n589 71.676
R2905 B.n844 B.n590 71.676
R2906 B.n840 B.n591 71.676
R2907 B.n836 B.n592 71.676
R2908 B.n832 B.n593 71.676
R2909 B.n828 B.n594 71.676
R2910 B.n824 B.n595 71.676
R2911 B.n820 B.n596 71.676
R2912 B.n816 B.n597 71.676
R2913 B.n812 B.n598 71.676
R2914 B.n808 B.n599 71.676
R2915 B.n804 B.n600 71.676
R2916 B.n800 B.n601 71.676
R2917 B.n796 B.n602 71.676
R2918 B.n792 B.n603 71.676
R2919 B.n788 B.n604 71.676
R2920 B.n784 B.n605 71.676
R2921 B.n780 B.n606 71.676
R2922 B.n775 B.n607 71.676
R2923 B.n771 B.n608 71.676
R2924 B.n767 B.n609 71.676
R2925 B.n763 B.n610 71.676
R2926 B.n759 B.n611 71.676
R2927 B.n755 B.n612 71.676
R2928 B.n751 B.n613 71.676
R2929 B.n747 B.n614 71.676
R2930 B.n743 B.n615 71.676
R2931 B.n739 B.n616 71.676
R2932 B.n735 B.n617 71.676
R2933 B.n731 B.n618 71.676
R2934 B.n727 B.n619 71.676
R2935 B.n723 B.n620 71.676
R2936 B.n719 B.n621 71.676
R2937 B.n715 B.n622 71.676
R2938 B.n711 B.n623 71.676
R2939 B.n707 B.n624 71.676
R2940 B.n703 B.n625 71.676
R2941 B.n699 B.n626 71.676
R2942 B.n695 B.n627 71.676
R2943 B.n691 B.n628 71.676
R2944 B.n687 B.n629 71.676
R2945 B.n683 B.n630 71.676
R2946 B.n679 B.n631 71.676
R2947 B.n675 B.n632 71.676
R2948 B.n671 B.n633 71.676
R2949 B.n667 B.n634 71.676
R2950 B.n663 B.n635 71.676
R2951 B.n659 B.n636 71.676
R2952 B.n655 B.n637 71.676
R2953 B.n651 B.n638 71.676
R2954 B.n647 B.n639 71.676
R2955 B.n895 B.n894 71.676
R2956 B.n893 B.n576 64.2658
R2957 B.n1193 B.n1192 64.2658
R2958 B.n646 B.n645 59.5399
R2959 B.n777 B.n643 59.5399
R2960 B.n193 B.n192 59.5399
R2961 B.n328 B.n190 59.5399
R2962 B.n195 B.n122 34.4981
R2963 B.n1190 B.n1189 34.4981
R2964 B.n897 B.n896 34.4981
R2965 B.n890 B.n574 34.4981
R2966 B.n900 B.n576 32.858
R2967 B.n900 B.n572 32.858
R2968 B.n906 B.n572 32.858
R2969 B.n906 B.n568 32.858
R2970 B.n912 B.n568 32.858
R2971 B.n912 B.n564 32.858
R2972 B.n918 B.n564 32.858
R2973 B.n918 B.n560 32.858
R2974 B.n924 B.n560 32.858
R2975 B.n930 B.n556 32.858
R2976 B.n930 B.n552 32.858
R2977 B.n936 B.n552 32.858
R2978 B.n936 B.n548 32.858
R2979 B.n942 B.n548 32.858
R2980 B.n942 B.n544 32.858
R2981 B.n948 B.n544 32.858
R2982 B.n948 B.n540 32.858
R2983 B.n954 B.n540 32.858
R2984 B.n954 B.n536 32.858
R2985 B.n960 B.n536 32.858
R2986 B.n960 B.n531 32.858
R2987 B.n966 B.n531 32.858
R2988 B.n966 B.n532 32.858
R2989 B.n972 B.n524 32.858
R2990 B.n978 B.n524 32.858
R2991 B.n978 B.n520 32.858
R2992 B.n984 B.n520 32.858
R2993 B.n984 B.n516 32.858
R2994 B.n990 B.n516 32.858
R2995 B.n990 B.n512 32.858
R2996 B.n996 B.n512 32.858
R2997 B.n996 B.n507 32.858
R2998 B.n1002 B.n507 32.858
R2999 B.n1002 B.n508 32.858
R3000 B.n1008 B.n500 32.858
R3001 B.n1014 B.n500 32.858
R3002 B.n1014 B.n496 32.858
R3003 B.n1020 B.n496 32.858
R3004 B.n1020 B.n492 32.858
R3005 B.n1026 B.n492 32.858
R3006 B.n1026 B.n488 32.858
R3007 B.n1032 B.n488 32.858
R3008 B.n1032 B.n484 32.858
R3009 B.n1038 B.n484 32.858
R3010 B.n1038 B.n480 32.858
R3011 B.n1044 B.n480 32.858
R3012 B.n1050 B.n476 32.858
R3013 B.n1050 B.n472 32.858
R3014 B.n1056 B.n472 32.858
R3015 B.n1056 B.n468 32.858
R3016 B.n1062 B.n468 32.858
R3017 B.n1062 B.n464 32.858
R3018 B.n1068 B.n464 32.858
R3019 B.n1068 B.n460 32.858
R3020 B.n1074 B.n460 32.858
R3021 B.n1074 B.n456 32.858
R3022 B.n1080 B.n456 32.858
R3023 B.n1086 B.n452 32.858
R3024 B.n1086 B.n448 32.858
R3025 B.n1093 B.n448 32.858
R3026 B.n1093 B.n444 32.858
R3027 B.n1099 B.n444 32.858
R3028 B.n1099 B.n4 32.858
R3029 B.n1330 B.n4 32.858
R3030 B.n1330 B.n1329 32.858
R3031 B.n1329 B.n1328 32.858
R3032 B.n1328 B.n8 32.858
R3033 B.n1322 B.n8 32.858
R3034 B.n1322 B.n1321 32.858
R3035 B.n1321 B.n1320 32.858
R3036 B.n1320 B.n15 32.858
R3037 B.n1314 B.n1313 32.858
R3038 B.n1313 B.n1312 32.858
R3039 B.n1312 B.n22 32.858
R3040 B.n1306 B.n22 32.858
R3041 B.n1306 B.n1305 32.858
R3042 B.n1305 B.n1304 32.858
R3043 B.n1304 B.n29 32.858
R3044 B.n1298 B.n29 32.858
R3045 B.n1298 B.n1297 32.858
R3046 B.n1297 B.n1296 32.858
R3047 B.n1296 B.n36 32.858
R3048 B.n1290 B.n1289 32.858
R3049 B.n1289 B.n1288 32.858
R3050 B.n1288 B.n43 32.858
R3051 B.n1282 B.n43 32.858
R3052 B.n1282 B.n1281 32.858
R3053 B.n1281 B.n1280 32.858
R3054 B.n1280 B.n50 32.858
R3055 B.n1274 B.n50 32.858
R3056 B.n1274 B.n1273 32.858
R3057 B.n1273 B.n1272 32.858
R3058 B.n1272 B.n57 32.858
R3059 B.n1266 B.n57 32.858
R3060 B.n1265 B.n1264 32.858
R3061 B.n1264 B.n64 32.858
R3062 B.n1258 B.n64 32.858
R3063 B.n1258 B.n1257 32.858
R3064 B.n1257 B.n1256 32.858
R3065 B.n1256 B.n71 32.858
R3066 B.n1250 B.n71 32.858
R3067 B.n1250 B.n1249 32.858
R3068 B.n1249 B.n1248 32.858
R3069 B.n1248 B.n78 32.858
R3070 B.n1242 B.n78 32.858
R3071 B.n1241 B.n1240 32.858
R3072 B.n1240 B.n85 32.858
R3073 B.n1234 B.n85 32.858
R3074 B.n1234 B.n1233 32.858
R3075 B.n1233 B.n1232 32.858
R3076 B.n1232 B.n92 32.858
R3077 B.n1226 B.n92 32.858
R3078 B.n1226 B.n1225 32.858
R3079 B.n1225 B.n1224 32.858
R3080 B.n1224 B.n99 32.858
R3081 B.n1218 B.n99 32.858
R3082 B.n1218 B.n1217 32.858
R3083 B.n1217 B.n1216 32.858
R3084 B.n1216 B.n106 32.858
R3085 B.n1210 B.n1209 32.858
R3086 B.n1209 B.n1208 32.858
R3087 B.n1208 B.n113 32.858
R3088 B.n1202 B.n113 32.858
R3089 B.n1202 B.n1201 32.858
R3090 B.n1201 B.n1200 32.858
R3091 B.n1200 B.n120 32.858
R3092 B.n1194 B.n120 32.858
R3093 B.n1194 B.n1193 32.858
R3094 B.t6 B.n476 29.9588
R3095 B.t0 B.n36 29.9588
R3096 B.n508 B.t2 28.9924
R3097 B.t3 B.n1265 28.9924
R3098 B.t9 B.n556 24.1604
R3099 B.t16 B.n106 24.1604
R3100 B.t7 B.n452 23.194
R3101 B.t1 B.n15 23.194
R3102 B.n532 B.t5 22.2276
R3103 B.t4 B.n1241 22.2276
R3104 B B.n1332 18.0485
R3105 B.n972 B.t5 10.6309
R3106 B.n1242 B.t4 10.6309
R3107 B.n196 B.n195 10.6151
R3108 B.n199 B.n196 10.6151
R3109 B.n200 B.n199 10.6151
R3110 B.n203 B.n200 10.6151
R3111 B.n204 B.n203 10.6151
R3112 B.n207 B.n204 10.6151
R3113 B.n208 B.n207 10.6151
R3114 B.n211 B.n208 10.6151
R3115 B.n212 B.n211 10.6151
R3116 B.n215 B.n212 10.6151
R3117 B.n216 B.n215 10.6151
R3118 B.n219 B.n216 10.6151
R3119 B.n220 B.n219 10.6151
R3120 B.n223 B.n220 10.6151
R3121 B.n224 B.n223 10.6151
R3122 B.n227 B.n224 10.6151
R3123 B.n228 B.n227 10.6151
R3124 B.n231 B.n228 10.6151
R3125 B.n232 B.n231 10.6151
R3126 B.n235 B.n232 10.6151
R3127 B.n236 B.n235 10.6151
R3128 B.n239 B.n236 10.6151
R3129 B.n240 B.n239 10.6151
R3130 B.n243 B.n240 10.6151
R3131 B.n244 B.n243 10.6151
R3132 B.n247 B.n244 10.6151
R3133 B.n248 B.n247 10.6151
R3134 B.n251 B.n248 10.6151
R3135 B.n252 B.n251 10.6151
R3136 B.n255 B.n252 10.6151
R3137 B.n256 B.n255 10.6151
R3138 B.n259 B.n256 10.6151
R3139 B.n260 B.n259 10.6151
R3140 B.n263 B.n260 10.6151
R3141 B.n264 B.n263 10.6151
R3142 B.n267 B.n264 10.6151
R3143 B.n268 B.n267 10.6151
R3144 B.n271 B.n268 10.6151
R3145 B.n272 B.n271 10.6151
R3146 B.n275 B.n272 10.6151
R3147 B.n276 B.n275 10.6151
R3148 B.n279 B.n276 10.6151
R3149 B.n280 B.n279 10.6151
R3150 B.n283 B.n280 10.6151
R3151 B.n284 B.n283 10.6151
R3152 B.n287 B.n284 10.6151
R3153 B.n288 B.n287 10.6151
R3154 B.n291 B.n288 10.6151
R3155 B.n292 B.n291 10.6151
R3156 B.n295 B.n292 10.6151
R3157 B.n296 B.n295 10.6151
R3158 B.n299 B.n296 10.6151
R3159 B.n300 B.n299 10.6151
R3160 B.n303 B.n300 10.6151
R3161 B.n304 B.n303 10.6151
R3162 B.n307 B.n304 10.6151
R3163 B.n308 B.n307 10.6151
R3164 B.n312 B.n311 10.6151
R3165 B.n315 B.n312 10.6151
R3166 B.n316 B.n315 10.6151
R3167 B.n319 B.n316 10.6151
R3168 B.n320 B.n319 10.6151
R3169 B.n323 B.n320 10.6151
R3170 B.n324 B.n323 10.6151
R3171 B.n327 B.n324 10.6151
R3172 B.n332 B.n329 10.6151
R3173 B.n333 B.n332 10.6151
R3174 B.n336 B.n333 10.6151
R3175 B.n337 B.n336 10.6151
R3176 B.n340 B.n337 10.6151
R3177 B.n341 B.n340 10.6151
R3178 B.n344 B.n341 10.6151
R3179 B.n345 B.n344 10.6151
R3180 B.n348 B.n345 10.6151
R3181 B.n349 B.n348 10.6151
R3182 B.n352 B.n349 10.6151
R3183 B.n353 B.n352 10.6151
R3184 B.n356 B.n353 10.6151
R3185 B.n357 B.n356 10.6151
R3186 B.n360 B.n357 10.6151
R3187 B.n361 B.n360 10.6151
R3188 B.n364 B.n361 10.6151
R3189 B.n365 B.n364 10.6151
R3190 B.n368 B.n365 10.6151
R3191 B.n369 B.n368 10.6151
R3192 B.n372 B.n369 10.6151
R3193 B.n373 B.n372 10.6151
R3194 B.n376 B.n373 10.6151
R3195 B.n377 B.n376 10.6151
R3196 B.n380 B.n377 10.6151
R3197 B.n381 B.n380 10.6151
R3198 B.n384 B.n381 10.6151
R3199 B.n385 B.n384 10.6151
R3200 B.n388 B.n385 10.6151
R3201 B.n389 B.n388 10.6151
R3202 B.n392 B.n389 10.6151
R3203 B.n393 B.n392 10.6151
R3204 B.n396 B.n393 10.6151
R3205 B.n397 B.n396 10.6151
R3206 B.n400 B.n397 10.6151
R3207 B.n401 B.n400 10.6151
R3208 B.n404 B.n401 10.6151
R3209 B.n405 B.n404 10.6151
R3210 B.n408 B.n405 10.6151
R3211 B.n409 B.n408 10.6151
R3212 B.n412 B.n409 10.6151
R3213 B.n413 B.n412 10.6151
R3214 B.n416 B.n413 10.6151
R3215 B.n417 B.n416 10.6151
R3216 B.n420 B.n417 10.6151
R3217 B.n421 B.n420 10.6151
R3218 B.n424 B.n421 10.6151
R3219 B.n425 B.n424 10.6151
R3220 B.n428 B.n425 10.6151
R3221 B.n429 B.n428 10.6151
R3222 B.n432 B.n429 10.6151
R3223 B.n433 B.n432 10.6151
R3224 B.n436 B.n433 10.6151
R3225 B.n437 B.n436 10.6151
R3226 B.n440 B.n437 10.6151
R3227 B.n441 B.n440 10.6151
R3228 B.n1190 B.n441 10.6151
R3229 B.n898 B.n897 10.6151
R3230 B.n898 B.n570 10.6151
R3231 B.n908 B.n570 10.6151
R3232 B.n909 B.n908 10.6151
R3233 B.n910 B.n909 10.6151
R3234 B.n910 B.n562 10.6151
R3235 B.n920 B.n562 10.6151
R3236 B.n921 B.n920 10.6151
R3237 B.n922 B.n921 10.6151
R3238 B.n922 B.n554 10.6151
R3239 B.n932 B.n554 10.6151
R3240 B.n933 B.n932 10.6151
R3241 B.n934 B.n933 10.6151
R3242 B.n934 B.n546 10.6151
R3243 B.n944 B.n546 10.6151
R3244 B.n945 B.n944 10.6151
R3245 B.n946 B.n945 10.6151
R3246 B.n946 B.n538 10.6151
R3247 B.n956 B.n538 10.6151
R3248 B.n957 B.n956 10.6151
R3249 B.n958 B.n957 10.6151
R3250 B.n958 B.n529 10.6151
R3251 B.n968 B.n529 10.6151
R3252 B.n969 B.n968 10.6151
R3253 B.n970 B.n969 10.6151
R3254 B.n970 B.n522 10.6151
R3255 B.n980 B.n522 10.6151
R3256 B.n981 B.n980 10.6151
R3257 B.n982 B.n981 10.6151
R3258 B.n982 B.n514 10.6151
R3259 B.n992 B.n514 10.6151
R3260 B.n993 B.n992 10.6151
R3261 B.n994 B.n993 10.6151
R3262 B.n994 B.n505 10.6151
R3263 B.n1004 B.n505 10.6151
R3264 B.n1005 B.n1004 10.6151
R3265 B.n1006 B.n1005 10.6151
R3266 B.n1006 B.n498 10.6151
R3267 B.n1016 B.n498 10.6151
R3268 B.n1017 B.n1016 10.6151
R3269 B.n1018 B.n1017 10.6151
R3270 B.n1018 B.n490 10.6151
R3271 B.n1028 B.n490 10.6151
R3272 B.n1029 B.n1028 10.6151
R3273 B.n1030 B.n1029 10.6151
R3274 B.n1030 B.n482 10.6151
R3275 B.n1040 B.n482 10.6151
R3276 B.n1041 B.n1040 10.6151
R3277 B.n1042 B.n1041 10.6151
R3278 B.n1042 B.n474 10.6151
R3279 B.n1052 B.n474 10.6151
R3280 B.n1053 B.n1052 10.6151
R3281 B.n1054 B.n1053 10.6151
R3282 B.n1054 B.n466 10.6151
R3283 B.n1064 B.n466 10.6151
R3284 B.n1065 B.n1064 10.6151
R3285 B.n1066 B.n1065 10.6151
R3286 B.n1066 B.n458 10.6151
R3287 B.n1076 B.n458 10.6151
R3288 B.n1077 B.n1076 10.6151
R3289 B.n1078 B.n1077 10.6151
R3290 B.n1078 B.n450 10.6151
R3291 B.n1088 B.n450 10.6151
R3292 B.n1089 B.n1088 10.6151
R3293 B.n1091 B.n1089 10.6151
R3294 B.n1091 B.n1090 10.6151
R3295 B.n1090 B.n442 10.6151
R3296 B.n1102 B.n442 10.6151
R3297 B.n1103 B.n1102 10.6151
R3298 B.n1104 B.n1103 10.6151
R3299 B.n1105 B.n1104 10.6151
R3300 B.n1107 B.n1105 10.6151
R3301 B.n1108 B.n1107 10.6151
R3302 B.n1109 B.n1108 10.6151
R3303 B.n1110 B.n1109 10.6151
R3304 B.n1112 B.n1110 10.6151
R3305 B.n1113 B.n1112 10.6151
R3306 B.n1114 B.n1113 10.6151
R3307 B.n1115 B.n1114 10.6151
R3308 B.n1117 B.n1115 10.6151
R3309 B.n1118 B.n1117 10.6151
R3310 B.n1119 B.n1118 10.6151
R3311 B.n1120 B.n1119 10.6151
R3312 B.n1122 B.n1120 10.6151
R3313 B.n1123 B.n1122 10.6151
R3314 B.n1124 B.n1123 10.6151
R3315 B.n1125 B.n1124 10.6151
R3316 B.n1127 B.n1125 10.6151
R3317 B.n1128 B.n1127 10.6151
R3318 B.n1129 B.n1128 10.6151
R3319 B.n1130 B.n1129 10.6151
R3320 B.n1132 B.n1130 10.6151
R3321 B.n1133 B.n1132 10.6151
R3322 B.n1134 B.n1133 10.6151
R3323 B.n1135 B.n1134 10.6151
R3324 B.n1137 B.n1135 10.6151
R3325 B.n1138 B.n1137 10.6151
R3326 B.n1139 B.n1138 10.6151
R3327 B.n1140 B.n1139 10.6151
R3328 B.n1142 B.n1140 10.6151
R3329 B.n1143 B.n1142 10.6151
R3330 B.n1144 B.n1143 10.6151
R3331 B.n1145 B.n1144 10.6151
R3332 B.n1147 B.n1145 10.6151
R3333 B.n1148 B.n1147 10.6151
R3334 B.n1149 B.n1148 10.6151
R3335 B.n1150 B.n1149 10.6151
R3336 B.n1152 B.n1150 10.6151
R3337 B.n1153 B.n1152 10.6151
R3338 B.n1154 B.n1153 10.6151
R3339 B.n1155 B.n1154 10.6151
R3340 B.n1157 B.n1155 10.6151
R3341 B.n1158 B.n1157 10.6151
R3342 B.n1159 B.n1158 10.6151
R3343 B.n1160 B.n1159 10.6151
R3344 B.n1162 B.n1160 10.6151
R3345 B.n1163 B.n1162 10.6151
R3346 B.n1164 B.n1163 10.6151
R3347 B.n1165 B.n1164 10.6151
R3348 B.n1167 B.n1165 10.6151
R3349 B.n1168 B.n1167 10.6151
R3350 B.n1169 B.n1168 10.6151
R3351 B.n1170 B.n1169 10.6151
R3352 B.n1172 B.n1170 10.6151
R3353 B.n1173 B.n1172 10.6151
R3354 B.n1174 B.n1173 10.6151
R3355 B.n1175 B.n1174 10.6151
R3356 B.n1177 B.n1175 10.6151
R3357 B.n1178 B.n1177 10.6151
R3358 B.n1179 B.n1178 10.6151
R3359 B.n1180 B.n1179 10.6151
R3360 B.n1182 B.n1180 10.6151
R3361 B.n1183 B.n1182 10.6151
R3362 B.n1184 B.n1183 10.6151
R3363 B.n1185 B.n1184 10.6151
R3364 B.n1187 B.n1185 10.6151
R3365 B.n1188 B.n1187 10.6151
R3366 B.n1189 B.n1188 10.6151
R3367 B.n890 B.n889 10.6151
R3368 B.n889 B.n888 10.6151
R3369 B.n888 B.n887 10.6151
R3370 B.n887 B.n885 10.6151
R3371 B.n885 B.n882 10.6151
R3372 B.n882 B.n881 10.6151
R3373 B.n881 B.n878 10.6151
R3374 B.n878 B.n877 10.6151
R3375 B.n877 B.n874 10.6151
R3376 B.n874 B.n873 10.6151
R3377 B.n873 B.n870 10.6151
R3378 B.n870 B.n869 10.6151
R3379 B.n869 B.n866 10.6151
R3380 B.n866 B.n865 10.6151
R3381 B.n865 B.n862 10.6151
R3382 B.n862 B.n861 10.6151
R3383 B.n861 B.n858 10.6151
R3384 B.n858 B.n857 10.6151
R3385 B.n857 B.n854 10.6151
R3386 B.n854 B.n853 10.6151
R3387 B.n853 B.n850 10.6151
R3388 B.n850 B.n849 10.6151
R3389 B.n849 B.n846 10.6151
R3390 B.n846 B.n845 10.6151
R3391 B.n845 B.n842 10.6151
R3392 B.n842 B.n841 10.6151
R3393 B.n841 B.n838 10.6151
R3394 B.n838 B.n837 10.6151
R3395 B.n837 B.n834 10.6151
R3396 B.n834 B.n833 10.6151
R3397 B.n833 B.n830 10.6151
R3398 B.n830 B.n829 10.6151
R3399 B.n829 B.n826 10.6151
R3400 B.n826 B.n825 10.6151
R3401 B.n825 B.n822 10.6151
R3402 B.n822 B.n821 10.6151
R3403 B.n821 B.n818 10.6151
R3404 B.n818 B.n817 10.6151
R3405 B.n817 B.n814 10.6151
R3406 B.n814 B.n813 10.6151
R3407 B.n813 B.n810 10.6151
R3408 B.n810 B.n809 10.6151
R3409 B.n809 B.n806 10.6151
R3410 B.n806 B.n805 10.6151
R3411 B.n805 B.n802 10.6151
R3412 B.n802 B.n801 10.6151
R3413 B.n801 B.n798 10.6151
R3414 B.n798 B.n797 10.6151
R3415 B.n797 B.n794 10.6151
R3416 B.n794 B.n793 10.6151
R3417 B.n793 B.n790 10.6151
R3418 B.n790 B.n789 10.6151
R3419 B.n789 B.n786 10.6151
R3420 B.n786 B.n785 10.6151
R3421 B.n785 B.n782 10.6151
R3422 B.n782 B.n781 10.6151
R3423 B.n781 B.n778 10.6151
R3424 B.n776 B.n773 10.6151
R3425 B.n773 B.n772 10.6151
R3426 B.n772 B.n769 10.6151
R3427 B.n769 B.n768 10.6151
R3428 B.n768 B.n765 10.6151
R3429 B.n765 B.n764 10.6151
R3430 B.n764 B.n761 10.6151
R3431 B.n761 B.n760 10.6151
R3432 B.n757 B.n756 10.6151
R3433 B.n756 B.n753 10.6151
R3434 B.n753 B.n752 10.6151
R3435 B.n752 B.n749 10.6151
R3436 B.n749 B.n748 10.6151
R3437 B.n748 B.n745 10.6151
R3438 B.n745 B.n744 10.6151
R3439 B.n744 B.n741 10.6151
R3440 B.n741 B.n740 10.6151
R3441 B.n740 B.n737 10.6151
R3442 B.n737 B.n736 10.6151
R3443 B.n736 B.n733 10.6151
R3444 B.n733 B.n732 10.6151
R3445 B.n732 B.n729 10.6151
R3446 B.n729 B.n728 10.6151
R3447 B.n728 B.n725 10.6151
R3448 B.n725 B.n724 10.6151
R3449 B.n724 B.n721 10.6151
R3450 B.n721 B.n720 10.6151
R3451 B.n720 B.n717 10.6151
R3452 B.n717 B.n716 10.6151
R3453 B.n716 B.n713 10.6151
R3454 B.n713 B.n712 10.6151
R3455 B.n712 B.n709 10.6151
R3456 B.n709 B.n708 10.6151
R3457 B.n708 B.n705 10.6151
R3458 B.n705 B.n704 10.6151
R3459 B.n704 B.n701 10.6151
R3460 B.n701 B.n700 10.6151
R3461 B.n700 B.n697 10.6151
R3462 B.n697 B.n696 10.6151
R3463 B.n696 B.n693 10.6151
R3464 B.n693 B.n692 10.6151
R3465 B.n692 B.n689 10.6151
R3466 B.n689 B.n688 10.6151
R3467 B.n688 B.n685 10.6151
R3468 B.n685 B.n684 10.6151
R3469 B.n684 B.n681 10.6151
R3470 B.n681 B.n680 10.6151
R3471 B.n680 B.n677 10.6151
R3472 B.n677 B.n676 10.6151
R3473 B.n676 B.n673 10.6151
R3474 B.n673 B.n672 10.6151
R3475 B.n672 B.n669 10.6151
R3476 B.n669 B.n668 10.6151
R3477 B.n668 B.n665 10.6151
R3478 B.n665 B.n664 10.6151
R3479 B.n664 B.n661 10.6151
R3480 B.n661 B.n660 10.6151
R3481 B.n660 B.n657 10.6151
R3482 B.n657 B.n656 10.6151
R3483 B.n656 B.n653 10.6151
R3484 B.n653 B.n652 10.6151
R3485 B.n652 B.n649 10.6151
R3486 B.n649 B.n648 10.6151
R3487 B.n648 B.n578 10.6151
R3488 B.n896 B.n578 10.6151
R3489 B.n902 B.n574 10.6151
R3490 B.n903 B.n902 10.6151
R3491 B.n904 B.n903 10.6151
R3492 B.n904 B.n566 10.6151
R3493 B.n914 B.n566 10.6151
R3494 B.n915 B.n914 10.6151
R3495 B.n916 B.n915 10.6151
R3496 B.n916 B.n558 10.6151
R3497 B.n926 B.n558 10.6151
R3498 B.n927 B.n926 10.6151
R3499 B.n928 B.n927 10.6151
R3500 B.n928 B.n550 10.6151
R3501 B.n938 B.n550 10.6151
R3502 B.n939 B.n938 10.6151
R3503 B.n940 B.n939 10.6151
R3504 B.n940 B.n542 10.6151
R3505 B.n950 B.n542 10.6151
R3506 B.n951 B.n950 10.6151
R3507 B.n952 B.n951 10.6151
R3508 B.n952 B.n534 10.6151
R3509 B.n962 B.n534 10.6151
R3510 B.n963 B.n962 10.6151
R3511 B.n964 B.n963 10.6151
R3512 B.n964 B.n526 10.6151
R3513 B.n974 B.n526 10.6151
R3514 B.n975 B.n974 10.6151
R3515 B.n976 B.n975 10.6151
R3516 B.n976 B.n518 10.6151
R3517 B.n986 B.n518 10.6151
R3518 B.n987 B.n986 10.6151
R3519 B.n988 B.n987 10.6151
R3520 B.n988 B.n510 10.6151
R3521 B.n998 B.n510 10.6151
R3522 B.n999 B.n998 10.6151
R3523 B.n1000 B.n999 10.6151
R3524 B.n1000 B.n502 10.6151
R3525 B.n1010 B.n502 10.6151
R3526 B.n1011 B.n1010 10.6151
R3527 B.n1012 B.n1011 10.6151
R3528 B.n1012 B.n494 10.6151
R3529 B.n1022 B.n494 10.6151
R3530 B.n1023 B.n1022 10.6151
R3531 B.n1024 B.n1023 10.6151
R3532 B.n1024 B.n486 10.6151
R3533 B.n1034 B.n486 10.6151
R3534 B.n1035 B.n1034 10.6151
R3535 B.n1036 B.n1035 10.6151
R3536 B.n1036 B.n478 10.6151
R3537 B.n1046 B.n478 10.6151
R3538 B.n1047 B.n1046 10.6151
R3539 B.n1048 B.n1047 10.6151
R3540 B.n1048 B.n470 10.6151
R3541 B.n1058 B.n470 10.6151
R3542 B.n1059 B.n1058 10.6151
R3543 B.n1060 B.n1059 10.6151
R3544 B.n1060 B.n462 10.6151
R3545 B.n1070 B.n462 10.6151
R3546 B.n1071 B.n1070 10.6151
R3547 B.n1072 B.n1071 10.6151
R3548 B.n1072 B.n454 10.6151
R3549 B.n1082 B.n454 10.6151
R3550 B.n1083 B.n1082 10.6151
R3551 B.n1084 B.n1083 10.6151
R3552 B.n1084 B.n446 10.6151
R3553 B.n1095 B.n446 10.6151
R3554 B.n1096 B.n1095 10.6151
R3555 B.n1097 B.n1096 10.6151
R3556 B.n1097 B.n0 10.6151
R3557 B.n1326 B.n1 10.6151
R3558 B.n1326 B.n1325 10.6151
R3559 B.n1325 B.n1324 10.6151
R3560 B.n1324 B.n10 10.6151
R3561 B.n1318 B.n10 10.6151
R3562 B.n1318 B.n1317 10.6151
R3563 B.n1317 B.n1316 10.6151
R3564 B.n1316 B.n17 10.6151
R3565 B.n1310 B.n17 10.6151
R3566 B.n1310 B.n1309 10.6151
R3567 B.n1309 B.n1308 10.6151
R3568 B.n1308 B.n24 10.6151
R3569 B.n1302 B.n24 10.6151
R3570 B.n1302 B.n1301 10.6151
R3571 B.n1301 B.n1300 10.6151
R3572 B.n1300 B.n31 10.6151
R3573 B.n1294 B.n31 10.6151
R3574 B.n1294 B.n1293 10.6151
R3575 B.n1293 B.n1292 10.6151
R3576 B.n1292 B.n38 10.6151
R3577 B.n1286 B.n38 10.6151
R3578 B.n1286 B.n1285 10.6151
R3579 B.n1285 B.n1284 10.6151
R3580 B.n1284 B.n45 10.6151
R3581 B.n1278 B.n45 10.6151
R3582 B.n1278 B.n1277 10.6151
R3583 B.n1277 B.n1276 10.6151
R3584 B.n1276 B.n52 10.6151
R3585 B.n1270 B.n52 10.6151
R3586 B.n1270 B.n1269 10.6151
R3587 B.n1269 B.n1268 10.6151
R3588 B.n1268 B.n59 10.6151
R3589 B.n1262 B.n59 10.6151
R3590 B.n1262 B.n1261 10.6151
R3591 B.n1261 B.n1260 10.6151
R3592 B.n1260 B.n66 10.6151
R3593 B.n1254 B.n66 10.6151
R3594 B.n1254 B.n1253 10.6151
R3595 B.n1253 B.n1252 10.6151
R3596 B.n1252 B.n73 10.6151
R3597 B.n1246 B.n73 10.6151
R3598 B.n1246 B.n1245 10.6151
R3599 B.n1245 B.n1244 10.6151
R3600 B.n1244 B.n80 10.6151
R3601 B.n1238 B.n80 10.6151
R3602 B.n1238 B.n1237 10.6151
R3603 B.n1237 B.n1236 10.6151
R3604 B.n1236 B.n87 10.6151
R3605 B.n1230 B.n87 10.6151
R3606 B.n1230 B.n1229 10.6151
R3607 B.n1229 B.n1228 10.6151
R3608 B.n1228 B.n94 10.6151
R3609 B.n1222 B.n94 10.6151
R3610 B.n1222 B.n1221 10.6151
R3611 B.n1221 B.n1220 10.6151
R3612 B.n1220 B.n101 10.6151
R3613 B.n1214 B.n101 10.6151
R3614 B.n1214 B.n1213 10.6151
R3615 B.n1213 B.n1212 10.6151
R3616 B.n1212 B.n108 10.6151
R3617 B.n1206 B.n108 10.6151
R3618 B.n1206 B.n1205 10.6151
R3619 B.n1205 B.n1204 10.6151
R3620 B.n1204 B.n115 10.6151
R3621 B.n1198 B.n115 10.6151
R3622 B.n1198 B.n1197 10.6151
R3623 B.n1197 B.n1196 10.6151
R3624 B.n1196 B.n122 10.6151
R3625 B.n1080 B.t7 9.66446
R3626 B.n1314 B.t1 9.66446
R3627 B.n924 B.t9 8.69806
R3628 B.n1210 B.t16 8.69806
R3629 B.n311 B.n193 6.5566
R3630 B.n328 B.n327 6.5566
R3631 B.n777 B.n776 6.5566
R3632 B.n760 B.n646 6.5566
R3633 B.n308 B.n193 4.05904
R3634 B.n329 B.n328 4.05904
R3635 B.n778 B.n777 4.05904
R3636 B.n757 B.n646 4.05904
R3637 B.n1008 B.t2 3.86608
R3638 B.n1266 B.t3 3.86608
R3639 B.n1044 B.t6 2.89969
R3640 B.n1290 B.t0 2.89969
R3641 B.n1332 B.n0 2.81026
R3642 B.n1332 B.n1 2.81026
R3643 VN.n71 VN.n37 161.3
R3644 VN.n70 VN.n69 161.3
R3645 VN.n68 VN.n38 161.3
R3646 VN.n67 VN.n66 161.3
R3647 VN.n65 VN.n39 161.3
R3648 VN.n64 VN.n63 161.3
R3649 VN.n62 VN.n40 161.3
R3650 VN.n61 VN.n60 161.3
R3651 VN.n58 VN.n41 161.3
R3652 VN.n57 VN.n56 161.3
R3653 VN.n55 VN.n42 161.3
R3654 VN.n54 VN.n53 161.3
R3655 VN.n52 VN.n43 161.3
R3656 VN.n51 VN.n50 161.3
R3657 VN.n49 VN.n44 161.3
R3658 VN.n48 VN.n47 161.3
R3659 VN.n34 VN.n0 161.3
R3660 VN.n33 VN.n32 161.3
R3661 VN.n31 VN.n1 161.3
R3662 VN.n30 VN.n29 161.3
R3663 VN.n28 VN.n2 161.3
R3664 VN.n27 VN.n26 161.3
R3665 VN.n25 VN.n3 161.3
R3666 VN.n24 VN.n23 161.3
R3667 VN.n21 VN.n4 161.3
R3668 VN.n20 VN.n19 161.3
R3669 VN.n18 VN.n5 161.3
R3670 VN.n17 VN.n16 161.3
R3671 VN.n15 VN.n6 161.3
R3672 VN.n14 VN.n13 161.3
R3673 VN.n12 VN.n7 161.3
R3674 VN.n11 VN.n10 161.3
R3675 VN.n8 VN.t1 142.483
R3676 VN.n45 VN.t5 142.483
R3677 VN.n9 VN.t7 110.344
R3678 VN.n22 VN.t0 110.344
R3679 VN.n35 VN.t4 110.344
R3680 VN.n46 VN.t3 110.344
R3681 VN.n59 VN.t6 110.344
R3682 VN.n72 VN.t2 110.344
R3683 VN VN.n73 61.0496
R3684 VN.n9 VN.n8 59.1721
R3685 VN.n46 VN.n45 59.1721
R3686 VN.n36 VN.n35 58.9381
R3687 VN.n73 VN.n72 58.9381
R3688 VN.n16 VN.n15 56.5193
R3689 VN.n53 VN.n52 56.5193
R3690 VN.n29 VN.n28 50.2061
R3691 VN.n66 VN.n65 50.2061
R3692 VN.n29 VN.n1 30.7807
R3693 VN.n66 VN.n38 30.7807
R3694 VN.n10 VN.n7 24.4675
R3695 VN.n14 VN.n7 24.4675
R3696 VN.n15 VN.n14 24.4675
R3697 VN.n16 VN.n5 24.4675
R3698 VN.n20 VN.n5 24.4675
R3699 VN.n21 VN.n20 24.4675
R3700 VN.n23 VN.n3 24.4675
R3701 VN.n27 VN.n3 24.4675
R3702 VN.n28 VN.n27 24.4675
R3703 VN.n33 VN.n1 24.4675
R3704 VN.n34 VN.n33 24.4675
R3705 VN.n52 VN.n51 24.4675
R3706 VN.n51 VN.n44 24.4675
R3707 VN.n47 VN.n44 24.4675
R3708 VN.n65 VN.n64 24.4675
R3709 VN.n64 VN.n40 24.4675
R3710 VN.n60 VN.n40 24.4675
R3711 VN.n58 VN.n57 24.4675
R3712 VN.n57 VN.n42 24.4675
R3713 VN.n53 VN.n42 24.4675
R3714 VN.n71 VN.n70 24.4675
R3715 VN.n70 VN.n38 24.4675
R3716 VN.n35 VN.n34 23.2442
R3717 VN.n72 VN.n71 23.2442
R3718 VN.n10 VN.n9 15.9041
R3719 VN.n22 VN.n21 15.9041
R3720 VN.n47 VN.n46 15.9041
R3721 VN.n59 VN.n58 15.9041
R3722 VN.n23 VN.n22 8.56395
R3723 VN.n60 VN.n59 8.56395
R3724 VN.n48 VN.n45 2.57337
R3725 VN.n11 VN.n8 2.57337
R3726 VN.n73 VN.n37 0.417535
R3727 VN.n36 VN.n0 0.417535
R3728 VN VN.n36 0.394291
R3729 VN.n69 VN.n37 0.189894
R3730 VN.n69 VN.n68 0.189894
R3731 VN.n68 VN.n67 0.189894
R3732 VN.n67 VN.n39 0.189894
R3733 VN.n63 VN.n39 0.189894
R3734 VN.n63 VN.n62 0.189894
R3735 VN.n62 VN.n61 0.189894
R3736 VN.n61 VN.n41 0.189894
R3737 VN.n56 VN.n41 0.189894
R3738 VN.n56 VN.n55 0.189894
R3739 VN.n55 VN.n54 0.189894
R3740 VN.n54 VN.n43 0.189894
R3741 VN.n50 VN.n43 0.189894
R3742 VN.n50 VN.n49 0.189894
R3743 VN.n49 VN.n48 0.189894
R3744 VN.n12 VN.n11 0.189894
R3745 VN.n13 VN.n12 0.189894
R3746 VN.n13 VN.n6 0.189894
R3747 VN.n17 VN.n6 0.189894
R3748 VN.n18 VN.n17 0.189894
R3749 VN.n19 VN.n18 0.189894
R3750 VN.n19 VN.n4 0.189894
R3751 VN.n24 VN.n4 0.189894
R3752 VN.n25 VN.n24 0.189894
R3753 VN.n26 VN.n25 0.189894
R3754 VN.n26 VN.n2 0.189894
R3755 VN.n30 VN.n2 0.189894
R3756 VN.n31 VN.n30 0.189894
R3757 VN.n32 VN.n31 0.189894
R3758 VN.n32 VN.n0 0.189894
R3759 VDD2.n2 VDD2.n1 61.8336
R3760 VDD2.n2 VDD2.n0 61.8336
R3761 VDD2 VDD2.n5 61.8308
R3762 VDD2.n4 VDD2.n3 60.1003
R3763 VDD2.n4 VDD2.n2 54.892
R3764 VDD2 VDD2.n4 1.84748
R3765 VDD2.n5 VDD2.t4 1.13258
R3766 VDD2.n5 VDD2.t2 1.13258
R3767 VDD2.n3 VDD2.t5 1.13258
R3768 VDD2.n3 VDD2.t1 1.13258
R3769 VDD2.n1 VDD2.t7 1.13258
R3770 VDD2.n1 VDD2.t3 1.13258
R3771 VDD2.n0 VDD2.t6 1.13258
R3772 VDD2.n0 VDD2.t0 1.13258
C0 VN VP 10.1749f
C1 VDD1 VN 0.153834f
C2 VTAIL VP 13.839f
C3 VDD1 VTAIL 10.135401f
C4 VDD2 VN 13.287701f
C5 VDD2 VTAIL 10.198f
C6 VDD1 VP 13.7813f
C7 VDD2 VP 0.649393f
C8 VDD1 VDD2 2.41002f
C9 VN VTAIL 13.8248f
C10 VDD2 B 7.021531f
C11 VDD1 B 7.587125f
C12 VTAIL B 14.635782f
C13 VN B 20.65579f
C14 VP B 19.271639f
C15 VDD2.t6 B 0.36629f
C16 VDD2.t0 B 0.36629f
C17 VDD2.n0 B 3.35118f
C18 VDD2.t7 B 0.36629f
C19 VDD2.t3 B 0.36629f
C20 VDD2.n1 B 3.35118f
C21 VDD2.n2 B 4.59663f
C22 VDD2.t5 B 0.36629f
C23 VDD2.t1 B 0.36629f
C24 VDD2.n3 B 3.33198f
C25 VDD2.n4 B 4.01649f
C26 VDD2.t4 B 0.36629f
C27 VDD2.t2 B 0.36629f
C28 VDD2.n5 B 3.35113f
C29 VN.n0 B 0.030613f
C30 VN.t4 B 2.98919f
C31 VN.n1 B 0.032604f
C32 VN.n2 B 0.016275f
C33 VN.n3 B 0.030332f
C34 VN.n4 B 0.016275f
C35 VN.t0 B 2.98919f
C36 VN.n5 B 0.030332f
C37 VN.n6 B 0.016275f
C38 VN.n7 B 0.030332f
C39 VN.t1 B 3.25069f
C40 VN.n8 B 1.04528f
C41 VN.t7 B 2.98919f
C42 VN.n9 B 1.09158f
C43 VN.n10 B 0.02509f
C44 VN.n11 B 0.211594f
C45 VN.n12 B 0.016275f
C46 VN.n13 B 0.016275f
C47 VN.n14 B 0.030332f
C48 VN.n15 B 0.023758f
C49 VN.n16 B 0.023758f
C50 VN.n17 B 0.016275f
C51 VN.n18 B 0.016275f
C52 VN.n19 B 0.016275f
C53 VN.n20 B 0.030332f
C54 VN.n21 B 0.02509f
C55 VN.n22 B 1.03073f
C56 VN.n23 B 0.020598f
C57 VN.n24 B 0.016275f
C58 VN.n25 B 0.016275f
C59 VN.n26 B 0.016275f
C60 VN.n27 B 0.030332f
C61 VN.n28 B 0.02987f
C62 VN.n29 B 0.015375f
C63 VN.n30 B 0.016275f
C64 VN.n31 B 0.016275f
C65 VN.n32 B 0.016275f
C66 VN.n33 B 0.030332f
C67 VN.n34 B 0.029583f
C68 VN.n35 B 1.10352f
C69 VN.n36 B 0.047995f
C70 VN.n37 B 0.030613f
C71 VN.t2 B 2.98919f
C72 VN.n38 B 0.032604f
C73 VN.n39 B 0.016275f
C74 VN.n40 B 0.030332f
C75 VN.n41 B 0.016275f
C76 VN.t6 B 2.98919f
C77 VN.n42 B 0.030332f
C78 VN.n43 B 0.016275f
C79 VN.n44 B 0.030332f
C80 VN.t5 B 3.25069f
C81 VN.n45 B 1.04528f
C82 VN.t3 B 2.98919f
C83 VN.n46 B 1.09158f
C84 VN.n47 B 0.02509f
C85 VN.n48 B 0.211594f
C86 VN.n49 B 0.016275f
C87 VN.n50 B 0.016275f
C88 VN.n51 B 0.030332f
C89 VN.n52 B 0.023758f
C90 VN.n53 B 0.023758f
C91 VN.n54 B 0.016275f
C92 VN.n55 B 0.016275f
C93 VN.n56 B 0.016275f
C94 VN.n57 B 0.030332f
C95 VN.n58 B 0.02509f
C96 VN.n59 B 1.03073f
C97 VN.n60 B 0.020598f
C98 VN.n61 B 0.016275f
C99 VN.n62 B 0.016275f
C100 VN.n63 B 0.016275f
C101 VN.n64 B 0.030332f
C102 VN.n65 B 0.02987f
C103 VN.n66 B 0.015375f
C104 VN.n67 B 0.016275f
C105 VN.n68 B 0.016275f
C106 VN.n69 B 0.016275f
C107 VN.n70 B 0.030332f
C108 VN.n71 B 0.029583f
C109 VN.n72 B 1.10352f
C110 VN.n73 B 1.23996f
C111 VDD1.t0 B 0.370547f
C112 VDD1.t3 B 0.370547f
C113 VDD1.n0 B 3.39165f
C114 VDD1.t4 B 0.370547f
C115 VDD1.t7 B 0.370547f
C116 VDD1.n1 B 3.39012f
C117 VDD1.t5 B 0.370547f
C118 VDD1.t1 B 0.370547f
C119 VDD1.n2 B 3.39012f
C120 VDD1.n3 B 4.705009f
C121 VDD1.t6 B 0.370547f
C122 VDD1.t2 B 0.370547f
C123 VDD1.n4 B 3.37069f
C124 VDD1.n5 B 4.09718f
C125 VTAIL.t0 B 0.265903f
C126 VTAIL.t3 B 0.265903f
C127 VTAIL.n0 B 2.35864f
C128 VTAIL.n1 B 0.419662f
C129 VTAIL.n2 B 0.026133f
C130 VTAIL.n3 B 0.019239f
C131 VTAIL.n4 B 0.010338f
C132 VTAIL.n5 B 0.024436f
C133 VTAIL.n6 B 0.010946f
C134 VTAIL.n7 B 0.019239f
C135 VTAIL.n8 B 0.010338f
C136 VTAIL.n9 B 0.024436f
C137 VTAIL.n10 B 0.010642f
C138 VTAIL.n11 B 0.019239f
C139 VTAIL.n12 B 0.010946f
C140 VTAIL.n13 B 0.024436f
C141 VTAIL.n14 B 0.010946f
C142 VTAIL.n15 B 0.019239f
C143 VTAIL.n16 B 0.010338f
C144 VTAIL.n17 B 0.024436f
C145 VTAIL.n18 B 0.010946f
C146 VTAIL.n19 B 0.019239f
C147 VTAIL.n20 B 0.010338f
C148 VTAIL.n21 B 0.024436f
C149 VTAIL.n22 B 0.010946f
C150 VTAIL.n23 B 0.019239f
C151 VTAIL.n24 B 0.010338f
C152 VTAIL.n25 B 0.024436f
C153 VTAIL.n26 B 0.010946f
C154 VTAIL.n27 B 0.019239f
C155 VTAIL.n28 B 0.010338f
C156 VTAIL.n29 B 0.024436f
C157 VTAIL.n30 B 0.010946f
C158 VTAIL.n31 B 1.47126f
C159 VTAIL.n32 B 0.010338f
C160 VTAIL.t1 B 0.040456f
C161 VTAIL.n33 B 0.137491f
C162 VTAIL.n34 B 0.014435f
C163 VTAIL.n35 B 0.018327f
C164 VTAIL.n36 B 0.024436f
C165 VTAIL.n37 B 0.010946f
C166 VTAIL.n38 B 0.010338f
C167 VTAIL.n39 B 0.019239f
C168 VTAIL.n40 B 0.019239f
C169 VTAIL.n41 B 0.010338f
C170 VTAIL.n42 B 0.010946f
C171 VTAIL.n43 B 0.024436f
C172 VTAIL.n44 B 0.024436f
C173 VTAIL.n45 B 0.010946f
C174 VTAIL.n46 B 0.010338f
C175 VTAIL.n47 B 0.019239f
C176 VTAIL.n48 B 0.019239f
C177 VTAIL.n49 B 0.010338f
C178 VTAIL.n50 B 0.010946f
C179 VTAIL.n51 B 0.024436f
C180 VTAIL.n52 B 0.024436f
C181 VTAIL.n53 B 0.010946f
C182 VTAIL.n54 B 0.010338f
C183 VTAIL.n55 B 0.019239f
C184 VTAIL.n56 B 0.019239f
C185 VTAIL.n57 B 0.010338f
C186 VTAIL.n58 B 0.010946f
C187 VTAIL.n59 B 0.024436f
C188 VTAIL.n60 B 0.024436f
C189 VTAIL.n61 B 0.010946f
C190 VTAIL.n62 B 0.010338f
C191 VTAIL.n63 B 0.019239f
C192 VTAIL.n64 B 0.019239f
C193 VTAIL.n65 B 0.010338f
C194 VTAIL.n66 B 0.010946f
C195 VTAIL.n67 B 0.024436f
C196 VTAIL.n68 B 0.024436f
C197 VTAIL.n69 B 0.010946f
C198 VTAIL.n70 B 0.010338f
C199 VTAIL.n71 B 0.019239f
C200 VTAIL.n72 B 0.019239f
C201 VTAIL.n73 B 0.010338f
C202 VTAIL.n74 B 0.010338f
C203 VTAIL.n75 B 0.010946f
C204 VTAIL.n76 B 0.024436f
C205 VTAIL.n77 B 0.024436f
C206 VTAIL.n78 B 0.024436f
C207 VTAIL.n79 B 0.010642f
C208 VTAIL.n80 B 0.010338f
C209 VTAIL.n81 B 0.019239f
C210 VTAIL.n82 B 0.019239f
C211 VTAIL.n83 B 0.010338f
C212 VTAIL.n84 B 0.010946f
C213 VTAIL.n85 B 0.024436f
C214 VTAIL.n86 B 0.024436f
C215 VTAIL.n87 B 0.010946f
C216 VTAIL.n88 B 0.010338f
C217 VTAIL.n89 B 0.019239f
C218 VTAIL.n90 B 0.019239f
C219 VTAIL.n91 B 0.010338f
C220 VTAIL.n92 B 0.010946f
C221 VTAIL.n93 B 0.024436f
C222 VTAIL.n94 B 0.051292f
C223 VTAIL.n95 B 0.010946f
C224 VTAIL.n96 B 0.010338f
C225 VTAIL.n97 B 0.043681f
C226 VTAIL.n98 B 0.02851f
C227 VTAIL.n99 B 0.266894f
C228 VTAIL.n100 B 0.026133f
C229 VTAIL.n101 B 0.019239f
C230 VTAIL.n102 B 0.010338f
C231 VTAIL.n103 B 0.024436f
C232 VTAIL.n104 B 0.010946f
C233 VTAIL.n105 B 0.019239f
C234 VTAIL.n106 B 0.010338f
C235 VTAIL.n107 B 0.024436f
C236 VTAIL.n108 B 0.010642f
C237 VTAIL.n109 B 0.019239f
C238 VTAIL.n110 B 0.010946f
C239 VTAIL.n111 B 0.024436f
C240 VTAIL.n112 B 0.010946f
C241 VTAIL.n113 B 0.019239f
C242 VTAIL.n114 B 0.010338f
C243 VTAIL.n115 B 0.024436f
C244 VTAIL.n116 B 0.010946f
C245 VTAIL.n117 B 0.019239f
C246 VTAIL.n118 B 0.010338f
C247 VTAIL.n119 B 0.024436f
C248 VTAIL.n120 B 0.010946f
C249 VTAIL.n121 B 0.019239f
C250 VTAIL.n122 B 0.010338f
C251 VTAIL.n123 B 0.024436f
C252 VTAIL.n124 B 0.010946f
C253 VTAIL.n125 B 0.019239f
C254 VTAIL.n126 B 0.010338f
C255 VTAIL.n127 B 0.024436f
C256 VTAIL.n128 B 0.010946f
C257 VTAIL.n129 B 1.47126f
C258 VTAIL.n130 B 0.010338f
C259 VTAIL.t14 B 0.040456f
C260 VTAIL.n131 B 0.137491f
C261 VTAIL.n132 B 0.014435f
C262 VTAIL.n133 B 0.018327f
C263 VTAIL.n134 B 0.024436f
C264 VTAIL.n135 B 0.010946f
C265 VTAIL.n136 B 0.010338f
C266 VTAIL.n137 B 0.019239f
C267 VTAIL.n138 B 0.019239f
C268 VTAIL.n139 B 0.010338f
C269 VTAIL.n140 B 0.010946f
C270 VTAIL.n141 B 0.024436f
C271 VTAIL.n142 B 0.024436f
C272 VTAIL.n143 B 0.010946f
C273 VTAIL.n144 B 0.010338f
C274 VTAIL.n145 B 0.019239f
C275 VTAIL.n146 B 0.019239f
C276 VTAIL.n147 B 0.010338f
C277 VTAIL.n148 B 0.010946f
C278 VTAIL.n149 B 0.024436f
C279 VTAIL.n150 B 0.024436f
C280 VTAIL.n151 B 0.010946f
C281 VTAIL.n152 B 0.010338f
C282 VTAIL.n153 B 0.019239f
C283 VTAIL.n154 B 0.019239f
C284 VTAIL.n155 B 0.010338f
C285 VTAIL.n156 B 0.010946f
C286 VTAIL.n157 B 0.024436f
C287 VTAIL.n158 B 0.024436f
C288 VTAIL.n159 B 0.010946f
C289 VTAIL.n160 B 0.010338f
C290 VTAIL.n161 B 0.019239f
C291 VTAIL.n162 B 0.019239f
C292 VTAIL.n163 B 0.010338f
C293 VTAIL.n164 B 0.010946f
C294 VTAIL.n165 B 0.024436f
C295 VTAIL.n166 B 0.024436f
C296 VTAIL.n167 B 0.010946f
C297 VTAIL.n168 B 0.010338f
C298 VTAIL.n169 B 0.019239f
C299 VTAIL.n170 B 0.019239f
C300 VTAIL.n171 B 0.010338f
C301 VTAIL.n172 B 0.010338f
C302 VTAIL.n173 B 0.010946f
C303 VTAIL.n174 B 0.024436f
C304 VTAIL.n175 B 0.024436f
C305 VTAIL.n176 B 0.024436f
C306 VTAIL.n177 B 0.010642f
C307 VTAIL.n178 B 0.010338f
C308 VTAIL.n179 B 0.019239f
C309 VTAIL.n180 B 0.019239f
C310 VTAIL.n181 B 0.010338f
C311 VTAIL.n182 B 0.010946f
C312 VTAIL.n183 B 0.024436f
C313 VTAIL.n184 B 0.024436f
C314 VTAIL.n185 B 0.010946f
C315 VTAIL.n186 B 0.010338f
C316 VTAIL.n187 B 0.019239f
C317 VTAIL.n188 B 0.019239f
C318 VTAIL.n189 B 0.010338f
C319 VTAIL.n190 B 0.010946f
C320 VTAIL.n191 B 0.024436f
C321 VTAIL.n192 B 0.051292f
C322 VTAIL.n193 B 0.010946f
C323 VTAIL.n194 B 0.010338f
C324 VTAIL.n195 B 0.043681f
C325 VTAIL.n196 B 0.02851f
C326 VTAIL.n197 B 0.266894f
C327 VTAIL.t12 B 0.265903f
C328 VTAIL.t13 B 0.265903f
C329 VTAIL.n198 B 2.35864f
C330 VTAIL.n199 B 0.637837f
C331 VTAIL.n200 B 0.026133f
C332 VTAIL.n201 B 0.019239f
C333 VTAIL.n202 B 0.010338f
C334 VTAIL.n203 B 0.024436f
C335 VTAIL.n204 B 0.010946f
C336 VTAIL.n205 B 0.019239f
C337 VTAIL.n206 B 0.010338f
C338 VTAIL.n207 B 0.024436f
C339 VTAIL.n208 B 0.010642f
C340 VTAIL.n209 B 0.019239f
C341 VTAIL.n210 B 0.010946f
C342 VTAIL.n211 B 0.024436f
C343 VTAIL.n212 B 0.010946f
C344 VTAIL.n213 B 0.019239f
C345 VTAIL.n214 B 0.010338f
C346 VTAIL.n215 B 0.024436f
C347 VTAIL.n216 B 0.010946f
C348 VTAIL.n217 B 0.019239f
C349 VTAIL.n218 B 0.010338f
C350 VTAIL.n219 B 0.024436f
C351 VTAIL.n220 B 0.010946f
C352 VTAIL.n221 B 0.019239f
C353 VTAIL.n222 B 0.010338f
C354 VTAIL.n223 B 0.024436f
C355 VTAIL.n224 B 0.010946f
C356 VTAIL.n225 B 0.019239f
C357 VTAIL.n226 B 0.010338f
C358 VTAIL.n227 B 0.024436f
C359 VTAIL.n228 B 0.010946f
C360 VTAIL.n229 B 1.47126f
C361 VTAIL.n230 B 0.010338f
C362 VTAIL.t11 B 0.040456f
C363 VTAIL.n231 B 0.137491f
C364 VTAIL.n232 B 0.014435f
C365 VTAIL.n233 B 0.018327f
C366 VTAIL.n234 B 0.024436f
C367 VTAIL.n235 B 0.010946f
C368 VTAIL.n236 B 0.010338f
C369 VTAIL.n237 B 0.019239f
C370 VTAIL.n238 B 0.019239f
C371 VTAIL.n239 B 0.010338f
C372 VTAIL.n240 B 0.010946f
C373 VTAIL.n241 B 0.024436f
C374 VTAIL.n242 B 0.024436f
C375 VTAIL.n243 B 0.010946f
C376 VTAIL.n244 B 0.010338f
C377 VTAIL.n245 B 0.019239f
C378 VTAIL.n246 B 0.019239f
C379 VTAIL.n247 B 0.010338f
C380 VTAIL.n248 B 0.010946f
C381 VTAIL.n249 B 0.024436f
C382 VTAIL.n250 B 0.024436f
C383 VTAIL.n251 B 0.010946f
C384 VTAIL.n252 B 0.010338f
C385 VTAIL.n253 B 0.019239f
C386 VTAIL.n254 B 0.019239f
C387 VTAIL.n255 B 0.010338f
C388 VTAIL.n256 B 0.010946f
C389 VTAIL.n257 B 0.024436f
C390 VTAIL.n258 B 0.024436f
C391 VTAIL.n259 B 0.010946f
C392 VTAIL.n260 B 0.010338f
C393 VTAIL.n261 B 0.019239f
C394 VTAIL.n262 B 0.019239f
C395 VTAIL.n263 B 0.010338f
C396 VTAIL.n264 B 0.010946f
C397 VTAIL.n265 B 0.024436f
C398 VTAIL.n266 B 0.024436f
C399 VTAIL.n267 B 0.010946f
C400 VTAIL.n268 B 0.010338f
C401 VTAIL.n269 B 0.019239f
C402 VTAIL.n270 B 0.019239f
C403 VTAIL.n271 B 0.010338f
C404 VTAIL.n272 B 0.010338f
C405 VTAIL.n273 B 0.010946f
C406 VTAIL.n274 B 0.024436f
C407 VTAIL.n275 B 0.024436f
C408 VTAIL.n276 B 0.024436f
C409 VTAIL.n277 B 0.010642f
C410 VTAIL.n278 B 0.010338f
C411 VTAIL.n279 B 0.019239f
C412 VTAIL.n280 B 0.019239f
C413 VTAIL.n281 B 0.010338f
C414 VTAIL.n282 B 0.010946f
C415 VTAIL.n283 B 0.024436f
C416 VTAIL.n284 B 0.024436f
C417 VTAIL.n285 B 0.010946f
C418 VTAIL.n286 B 0.010338f
C419 VTAIL.n287 B 0.019239f
C420 VTAIL.n288 B 0.019239f
C421 VTAIL.n289 B 0.010338f
C422 VTAIL.n290 B 0.010946f
C423 VTAIL.n291 B 0.024436f
C424 VTAIL.n292 B 0.051292f
C425 VTAIL.n293 B 0.010946f
C426 VTAIL.n294 B 0.010338f
C427 VTAIL.n295 B 0.043681f
C428 VTAIL.n296 B 0.02851f
C429 VTAIL.n297 B 1.65558f
C430 VTAIL.n298 B 0.026133f
C431 VTAIL.n299 B 0.019239f
C432 VTAIL.n300 B 0.010338f
C433 VTAIL.n301 B 0.024436f
C434 VTAIL.n302 B 0.010946f
C435 VTAIL.n303 B 0.019239f
C436 VTAIL.n304 B 0.010338f
C437 VTAIL.n305 B 0.024436f
C438 VTAIL.n306 B 0.010642f
C439 VTAIL.n307 B 0.019239f
C440 VTAIL.n308 B 0.010642f
C441 VTAIL.n309 B 0.010338f
C442 VTAIL.n310 B 0.024436f
C443 VTAIL.n311 B 0.024436f
C444 VTAIL.n312 B 0.010946f
C445 VTAIL.n313 B 0.019239f
C446 VTAIL.n314 B 0.010338f
C447 VTAIL.n315 B 0.024436f
C448 VTAIL.n316 B 0.010946f
C449 VTAIL.n317 B 0.019239f
C450 VTAIL.n318 B 0.010338f
C451 VTAIL.n319 B 0.024436f
C452 VTAIL.n320 B 0.010946f
C453 VTAIL.n321 B 0.019239f
C454 VTAIL.n322 B 0.010338f
C455 VTAIL.n323 B 0.024436f
C456 VTAIL.n324 B 0.010946f
C457 VTAIL.n325 B 0.019239f
C458 VTAIL.n326 B 0.010338f
C459 VTAIL.n327 B 0.024436f
C460 VTAIL.n328 B 0.010946f
C461 VTAIL.n329 B 1.47126f
C462 VTAIL.n330 B 0.010338f
C463 VTAIL.t5 B 0.040456f
C464 VTAIL.n331 B 0.137491f
C465 VTAIL.n332 B 0.014435f
C466 VTAIL.n333 B 0.018327f
C467 VTAIL.n334 B 0.024436f
C468 VTAIL.n335 B 0.010946f
C469 VTAIL.n336 B 0.010338f
C470 VTAIL.n337 B 0.019239f
C471 VTAIL.n338 B 0.019239f
C472 VTAIL.n339 B 0.010338f
C473 VTAIL.n340 B 0.010946f
C474 VTAIL.n341 B 0.024436f
C475 VTAIL.n342 B 0.024436f
C476 VTAIL.n343 B 0.010946f
C477 VTAIL.n344 B 0.010338f
C478 VTAIL.n345 B 0.019239f
C479 VTAIL.n346 B 0.019239f
C480 VTAIL.n347 B 0.010338f
C481 VTAIL.n348 B 0.010946f
C482 VTAIL.n349 B 0.024436f
C483 VTAIL.n350 B 0.024436f
C484 VTAIL.n351 B 0.010946f
C485 VTAIL.n352 B 0.010338f
C486 VTAIL.n353 B 0.019239f
C487 VTAIL.n354 B 0.019239f
C488 VTAIL.n355 B 0.010338f
C489 VTAIL.n356 B 0.010946f
C490 VTAIL.n357 B 0.024436f
C491 VTAIL.n358 B 0.024436f
C492 VTAIL.n359 B 0.010946f
C493 VTAIL.n360 B 0.010338f
C494 VTAIL.n361 B 0.019239f
C495 VTAIL.n362 B 0.019239f
C496 VTAIL.n363 B 0.010338f
C497 VTAIL.n364 B 0.010946f
C498 VTAIL.n365 B 0.024436f
C499 VTAIL.n366 B 0.024436f
C500 VTAIL.n367 B 0.010946f
C501 VTAIL.n368 B 0.010338f
C502 VTAIL.n369 B 0.019239f
C503 VTAIL.n370 B 0.019239f
C504 VTAIL.n371 B 0.010338f
C505 VTAIL.n372 B 0.010946f
C506 VTAIL.n373 B 0.024436f
C507 VTAIL.n374 B 0.024436f
C508 VTAIL.n375 B 0.010946f
C509 VTAIL.n376 B 0.010338f
C510 VTAIL.n377 B 0.019239f
C511 VTAIL.n378 B 0.019239f
C512 VTAIL.n379 B 0.010338f
C513 VTAIL.n380 B 0.010946f
C514 VTAIL.n381 B 0.024436f
C515 VTAIL.n382 B 0.024436f
C516 VTAIL.n383 B 0.010946f
C517 VTAIL.n384 B 0.010338f
C518 VTAIL.n385 B 0.019239f
C519 VTAIL.n386 B 0.019239f
C520 VTAIL.n387 B 0.010338f
C521 VTAIL.n388 B 0.010946f
C522 VTAIL.n389 B 0.024436f
C523 VTAIL.n390 B 0.051292f
C524 VTAIL.n391 B 0.010946f
C525 VTAIL.n392 B 0.010338f
C526 VTAIL.n393 B 0.043681f
C527 VTAIL.n394 B 0.02851f
C528 VTAIL.n395 B 1.65558f
C529 VTAIL.t2 B 0.265903f
C530 VTAIL.t6 B 0.265903f
C531 VTAIL.n396 B 2.35865f
C532 VTAIL.n397 B 0.637826f
C533 VTAIL.n398 B 0.026133f
C534 VTAIL.n399 B 0.019239f
C535 VTAIL.n400 B 0.010338f
C536 VTAIL.n401 B 0.024436f
C537 VTAIL.n402 B 0.010946f
C538 VTAIL.n403 B 0.019239f
C539 VTAIL.n404 B 0.010338f
C540 VTAIL.n405 B 0.024436f
C541 VTAIL.n406 B 0.010642f
C542 VTAIL.n407 B 0.019239f
C543 VTAIL.n408 B 0.010642f
C544 VTAIL.n409 B 0.010338f
C545 VTAIL.n410 B 0.024436f
C546 VTAIL.n411 B 0.024436f
C547 VTAIL.n412 B 0.010946f
C548 VTAIL.n413 B 0.019239f
C549 VTAIL.n414 B 0.010338f
C550 VTAIL.n415 B 0.024436f
C551 VTAIL.n416 B 0.010946f
C552 VTAIL.n417 B 0.019239f
C553 VTAIL.n418 B 0.010338f
C554 VTAIL.n419 B 0.024436f
C555 VTAIL.n420 B 0.010946f
C556 VTAIL.n421 B 0.019239f
C557 VTAIL.n422 B 0.010338f
C558 VTAIL.n423 B 0.024436f
C559 VTAIL.n424 B 0.010946f
C560 VTAIL.n425 B 0.019239f
C561 VTAIL.n426 B 0.010338f
C562 VTAIL.n427 B 0.024436f
C563 VTAIL.n428 B 0.010946f
C564 VTAIL.n429 B 1.47126f
C565 VTAIL.n430 B 0.010338f
C566 VTAIL.t7 B 0.040456f
C567 VTAIL.n431 B 0.137491f
C568 VTAIL.n432 B 0.014435f
C569 VTAIL.n433 B 0.018327f
C570 VTAIL.n434 B 0.024436f
C571 VTAIL.n435 B 0.010946f
C572 VTAIL.n436 B 0.010338f
C573 VTAIL.n437 B 0.019239f
C574 VTAIL.n438 B 0.019239f
C575 VTAIL.n439 B 0.010338f
C576 VTAIL.n440 B 0.010946f
C577 VTAIL.n441 B 0.024436f
C578 VTAIL.n442 B 0.024436f
C579 VTAIL.n443 B 0.010946f
C580 VTAIL.n444 B 0.010338f
C581 VTAIL.n445 B 0.019239f
C582 VTAIL.n446 B 0.019239f
C583 VTAIL.n447 B 0.010338f
C584 VTAIL.n448 B 0.010946f
C585 VTAIL.n449 B 0.024436f
C586 VTAIL.n450 B 0.024436f
C587 VTAIL.n451 B 0.010946f
C588 VTAIL.n452 B 0.010338f
C589 VTAIL.n453 B 0.019239f
C590 VTAIL.n454 B 0.019239f
C591 VTAIL.n455 B 0.010338f
C592 VTAIL.n456 B 0.010946f
C593 VTAIL.n457 B 0.024436f
C594 VTAIL.n458 B 0.024436f
C595 VTAIL.n459 B 0.010946f
C596 VTAIL.n460 B 0.010338f
C597 VTAIL.n461 B 0.019239f
C598 VTAIL.n462 B 0.019239f
C599 VTAIL.n463 B 0.010338f
C600 VTAIL.n464 B 0.010946f
C601 VTAIL.n465 B 0.024436f
C602 VTAIL.n466 B 0.024436f
C603 VTAIL.n467 B 0.010946f
C604 VTAIL.n468 B 0.010338f
C605 VTAIL.n469 B 0.019239f
C606 VTAIL.n470 B 0.019239f
C607 VTAIL.n471 B 0.010338f
C608 VTAIL.n472 B 0.010946f
C609 VTAIL.n473 B 0.024436f
C610 VTAIL.n474 B 0.024436f
C611 VTAIL.n475 B 0.010946f
C612 VTAIL.n476 B 0.010338f
C613 VTAIL.n477 B 0.019239f
C614 VTAIL.n478 B 0.019239f
C615 VTAIL.n479 B 0.010338f
C616 VTAIL.n480 B 0.010946f
C617 VTAIL.n481 B 0.024436f
C618 VTAIL.n482 B 0.024436f
C619 VTAIL.n483 B 0.010946f
C620 VTAIL.n484 B 0.010338f
C621 VTAIL.n485 B 0.019239f
C622 VTAIL.n486 B 0.019239f
C623 VTAIL.n487 B 0.010338f
C624 VTAIL.n488 B 0.010946f
C625 VTAIL.n489 B 0.024436f
C626 VTAIL.n490 B 0.051292f
C627 VTAIL.n491 B 0.010946f
C628 VTAIL.n492 B 0.010338f
C629 VTAIL.n493 B 0.043681f
C630 VTAIL.n494 B 0.02851f
C631 VTAIL.n495 B 0.266894f
C632 VTAIL.n496 B 0.026133f
C633 VTAIL.n497 B 0.019239f
C634 VTAIL.n498 B 0.010338f
C635 VTAIL.n499 B 0.024436f
C636 VTAIL.n500 B 0.010946f
C637 VTAIL.n501 B 0.019239f
C638 VTAIL.n502 B 0.010338f
C639 VTAIL.n503 B 0.024436f
C640 VTAIL.n504 B 0.010642f
C641 VTAIL.n505 B 0.019239f
C642 VTAIL.n506 B 0.010642f
C643 VTAIL.n507 B 0.010338f
C644 VTAIL.n508 B 0.024436f
C645 VTAIL.n509 B 0.024436f
C646 VTAIL.n510 B 0.010946f
C647 VTAIL.n511 B 0.019239f
C648 VTAIL.n512 B 0.010338f
C649 VTAIL.n513 B 0.024436f
C650 VTAIL.n514 B 0.010946f
C651 VTAIL.n515 B 0.019239f
C652 VTAIL.n516 B 0.010338f
C653 VTAIL.n517 B 0.024436f
C654 VTAIL.n518 B 0.010946f
C655 VTAIL.n519 B 0.019239f
C656 VTAIL.n520 B 0.010338f
C657 VTAIL.n521 B 0.024436f
C658 VTAIL.n522 B 0.010946f
C659 VTAIL.n523 B 0.019239f
C660 VTAIL.n524 B 0.010338f
C661 VTAIL.n525 B 0.024436f
C662 VTAIL.n526 B 0.010946f
C663 VTAIL.n527 B 1.47126f
C664 VTAIL.n528 B 0.010338f
C665 VTAIL.t8 B 0.040456f
C666 VTAIL.n529 B 0.137491f
C667 VTAIL.n530 B 0.014435f
C668 VTAIL.n531 B 0.018327f
C669 VTAIL.n532 B 0.024436f
C670 VTAIL.n533 B 0.010946f
C671 VTAIL.n534 B 0.010338f
C672 VTAIL.n535 B 0.019239f
C673 VTAIL.n536 B 0.019239f
C674 VTAIL.n537 B 0.010338f
C675 VTAIL.n538 B 0.010946f
C676 VTAIL.n539 B 0.024436f
C677 VTAIL.n540 B 0.024436f
C678 VTAIL.n541 B 0.010946f
C679 VTAIL.n542 B 0.010338f
C680 VTAIL.n543 B 0.019239f
C681 VTAIL.n544 B 0.019239f
C682 VTAIL.n545 B 0.010338f
C683 VTAIL.n546 B 0.010946f
C684 VTAIL.n547 B 0.024436f
C685 VTAIL.n548 B 0.024436f
C686 VTAIL.n549 B 0.010946f
C687 VTAIL.n550 B 0.010338f
C688 VTAIL.n551 B 0.019239f
C689 VTAIL.n552 B 0.019239f
C690 VTAIL.n553 B 0.010338f
C691 VTAIL.n554 B 0.010946f
C692 VTAIL.n555 B 0.024436f
C693 VTAIL.n556 B 0.024436f
C694 VTAIL.n557 B 0.010946f
C695 VTAIL.n558 B 0.010338f
C696 VTAIL.n559 B 0.019239f
C697 VTAIL.n560 B 0.019239f
C698 VTAIL.n561 B 0.010338f
C699 VTAIL.n562 B 0.010946f
C700 VTAIL.n563 B 0.024436f
C701 VTAIL.n564 B 0.024436f
C702 VTAIL.n565 B 0.010946f
C703 VTAIL.n566 B 0.010338f
C704 VTAIL.n567 B 0.019239f
C705 VTAIL.n568 B 0.019239f
C706 VTAIL.n569 B 0.010338f
C707 VTAIL.n570 B 0.010946f
C708 VTAIL.n571 B 0.024436f
C709 VTAIL.n572 B 0.024436f
C710 VTAIL.n573 B 0.010946f
C711 VTAIL.n574 B 0.010338f
C712 VTAIL.n575 B 0.019239f
C713 VTAIL.n576 B 0.019239f
C714 VTAIL.n577 B 0.010338f
C715 VTAIL.n578 B 0.010946f
C716 VTAIL.n579 B 0.024436f
C717 VTAIL.n580 B 0.024436f
C718 VTAIL.n581 B 0.010946f
C719 VTAIL.n582 B 0.010338f
C720 VTAIL.n583 B 0.019239f
C721 VTAIL.n584 B 0.019239f
C722 VTAIL.n585 B 0.010338f
C723 VTAIL.n586 B 0.010946f
C724 VTAIL.n587 B 0.024436f
C725 VTAIL.n588 B 0.051292f
C726 VTAIL.n589 B 0.010946f
C727 VTAIL.n590 B 0.010338f
C728 VTAIL.n591 B 0.043681f
C729 VTAIL.n592 B 0.02851f
C730 VTAIL.n593 B 0.266894f
C731 VTAIL.t15 B 0.265903f
C732 VTAIL.t10 B 0.265903f
C733 VTAIL.n594 B 2.35865f
C734 VTAIL.n595 B 0.637826f
C735 VTAIL.n596 B 0.026133f
C736 VTAIL.n597 B 0.019239f
C737 VTAIL.n598 B 0.010338f
C738 VTAIL.n599 B 0.024436f
C739 VTAIL.n600 B 0.010946f
C740 VTAIL.n601 B 0.019239f
C741 VTAIL.n602 B 0.010338f
C742 VTAIL.n603 B 0.024436f
C743 VTAIL.n604 B 0.010642f
C744 VTAIL.n605 B 0.019239f
C745 VTAIL.n606 B 0.010642f
C746 VTAIL.n607 B 0.010338f
C747 VTAIL.n608 B 0.024436f
C748 VTAIL.n609 B 0.024436f
C749 VTAIL.n610 B 0.010946f
C750 VTAIL.n611 B 0.019239f
C751 VTAIL.n612 B 0.010338f
C752 VTAIL.n613 B 0.024436f
C753 VTAIL.n614 B 0.010946f
C754 VTAIL.n615 B 0.019239f
C755 VTAIL.n616 B 0.010338f
C756 VTAIL.n617 B 0.024436f
C757 VTAIL.n618 B 0.010946f
C758 VTAIL.n619 B 0.019239f
C759 VTAIL.n620 B 0.010338f
C760 VTAIL.n621 B 0.024436f
C761 VTAIL.n622 B 0.010946f
C762 VTAIL.n623 B 0.019239f
C763 VTAIL.n624 B 0.010338f
C764 VTAIL.n625 B 0.024436f
C765 VTAIL.n626 B 0.010946f
C766 VTAIL.n627 B 1.47126f
C767 VTAIL.n628 B 0.010338f
C768 VTAIL.t9 B 0.040456f
C769 VTAIL.n629 B 0.137491f
C770 VTAIL.n630 B 0.014435f
C771 VTAIL.n631 B 0.018327f
C772 VTAIL.n632 B 0.024436f
C773 VTAIL.n633 B 0.010946f
C774 VTAIL.n634 B 0.010338f
C775 VTAIL.n635 B 0.019239f
C776 VTAIL.n636 B 0.019239f
C777 VTAIL.n637 B 0.010338f
C778 VTAIL.n638 B 0.010946f
C779 VTAIL.n639 B 0.024436f
C780 VTAIL.n640 B 0.024436f
C781 VTAIL.n641 B 0.010946f
C782 VTAIL.n642 B 0.010338f
C783 VTAIL.n643 B 0.019239f
C784 VTAIL.n644 B 0.019239f
C785 VTAIL.n645 B 0.010338f
C786 VTAIL.n646 B 0.010946f
C787 VTAIL.n647 B 0.024436f
C788 VTAIL.n648 B 0.024436f
C789 VTAIL.n649 B 0.010946f
C790 VTAIL.n650 B 0.010338f
C791 VTAIL.n651 B 0.019239f
C792 VTAIL.n652 B 0.019239f
C793 VTAIL.n653 B 0.010338f
C794 VTAIL.n654 B 0.010946f
C795 VTAIL.n655 B 0.024436f
C796 VTAIL.n656 B 0.024436f
C797 VTAIL.n657 B 0.010946f
C798 VTAIL.n658 B 0.010338f
C799 VTAIL.n659 B 0.019239f
C800 VTAIL.n660 B 0.019239f
C801 VTAIL.n661 B 0.010338f
C802 VTAIL.n662 B 0.010946f
C803 VTAIL.n663 B 0.024436f
C804 VTAIL.n664 B 0.024436f
C805 VTAIL.n665 B 0.010946f
C806 VTAIL.n666 B 0.010338f
C807 VTAIL.n667 B 0.019239f
C808 VTAIL.n668 B 0.019239f
C809 VTAIL.n669 B 0.010338f
C810 VTAIL.n670 B 0.010946f
C811 VTAIL.n671 B 0.024436f
C812 VTAIL.n672 B 0.024436f
C813 VTAIL.n673 B 0.010946f
C814 VTAIL.n674 B 0.010338f
C815 VTAIL.n675 B 0.019239f
C816 VTAIL.n676 B 0.019239f
C817 VTAIL.n677 B 0.010338f
C818 VTAIL.n678 B 0.010946f
C819 VTAIL.n679 B 0.024436f
C820 VTAIL.n680 B 0.024436f
C821 VTAIL.n681 B 0.010946f
C822 VTAIL.n682 B 0.010338f
C823 VTAIL.n683 B 0.019239f
C824 VTAIL.n684 B 0.019239f
C825 VTAIL.n685 B 0.010338f
C826 VTAIL.n686 B 0.010946f
C827 VTAIL.n687 B 0.024436f
C828 VTAIL.n688 B 0.051292f
C829 VTAIL.n689 B 0.010946f
C830 VTAIL.n690 B 0.010338f
C831 VTAIL.n691 B 0.043681f
C832 VTAIL.n692 B 0.02851f
C833 VTAIL.n693 B 1.65558f
C834 VTAIL.n694 B 0.026133f
C835 VTAIL.n695 B 0.019239f
C836 VTAIL.n696 B 0.010338f
C837 VTAIL.n697 B 0.024436f
C838 VTAIL.n698 B 0.010946f
C839 VTAIL.n699 B 0.019239f
C840 VTAIL.n700 B 0.010338f
C841 VTAIL.n701 B 0.024436f
C842 VTAIL.n702 B 0.010642f
C843 VTAIL.n703 B 0.019239f
C844 VTAIL.n704 B 0.010946f
C845 VTAIL.n705 B 0.024436f
C846 VTAIL.n706 B 0.010946f
C847 VTAIL.n707 B 0.019239f
C848 VTAIL.n708 B 0.010338f
C849 VTAIL.n709 B 0.024436f
C850 VTAIL.n710 B 0.010946f
C851 VTAIL.n711 B 0.019239f
C852 VTAIL.n712 B 0.010338f
C853 VTAIL.n713 B 0.024436f
C854 VTAIL.n714 B 0.010946f
C855 VTAIL.n715 B 0.019239f
C856 VTAIL.n716 B 0.010338f
C857 VTAIL.n717 B 0.024436f
C858 VTAIL.n718 B 0.010946f
C859 VTAIL.n719 B 0.019239f
C860 VTAIL.n720 B 0.010338f
C861 VTAIL.n721 B 0.024436f
C862 VTAIL.n722 B 0.010946f
C863 VTAIL.n723 B 1.47126f
C864 VTAIL.n724 B 0.010338f
C865 VTAIL.t4 B 0.040456f
C866 VTAIL.n725 B 0.137491f
C867 VTAIL.n726 B 0.014435f
C868 VTAIL.n727 B 0.018327f
C869 VTAIL.n728 B 0.024436f
C870 VTAIL.n729 B 0.010946f
C871 VTAIL.n730 B 0.010338f
C872 VTAIL.n731 B 0.019239f
C873 VTAIL.n732 B 0.019239f
C874 VTAIL.n733 B 0.010338f
C875 VTAIL.n734 B 0.010946f
C876 VTAIL.n735 B 0.024436f
C877 VTAIL.n736 B 0.024436f
C878 VTAIL.n737 B 0.010946f
C879 VTAIL.n738 B 0.010338f
C880 VTAIL.n739 B 0.019239f
C881 VTAIL.n740 B 0.019239f
C882 VTAIL.n741 B 0.010338f
C883 VTAIL.n742 B 0.010946f
C884 VTAIL.n743 B 0.024436f
C885 VTAIL.n744 B 0.024436f
C886 VTAIL.n745 B 0.010946f
C887 VTAIL.n746 B 0.010338f
C888 VTAIL.n747 B 0.019239f
C889 VTAIL.n748 B 0.019239f
C890 VTAIL.n749 B 0.010338f
C891 VTAIL.n750 B 0.010946f
C892 VTAIL.n751 B 0.024436f
C893 VTAIL.n752 B 0.024436f
C894 VTAIL.n753 B 0.010946f
C895 VTAIL.n754 B 0.010338f
C896 VTAIL.n755 B 0.019239f
C897 VTAIL.n756 B 0.019239f
C898 VTAIL.n757 B 0.010338f
C899 VTAIL.n758 B 0.010946f
C900 VTAIL.n759 B 0.024436f
C901 VTAIL.n760 B 0.024436f
C902 VTAIL.n761 B 0.010946f
C903 VTAIL.n762 B 0.010338f
C904 VTAIL.n763 B 0.019239f
C905 VTAIL.n764 B 0.019239f
C906 VTAIL.n765 B 0.010338f
C907 VTAIL.n766 B 0.010338f
C908 VTAIL.n767 B 0.010946f
C909 VTAIL.n768 B 0.024436f
C910 VTAIL.n769 B 0.024436f
C911 VTAIL.n770 B 0.024436f
C912 VTAIL.n771 B 0.010642f
C913 VTAIL.n772 B 0.010338f
C914 VTAIL.n773 B 0.019239f
C915 VTAIL.n774 B 0.019239f
C916 VTAIL.n775 B 0.010338f
C917 VTAIL.n776 B 0.010946f
C918 VTAIL.n777 B 0.024436f
C919 VTAIL.n778 B 0.024436f
C920 VTAIL.n779 B 0.010946f
C921 VTAIL.n780 B 0.010338f
C922 VTAIL.n781 B 0.019239f
C923 VTAIL.n782 B 0.019239f
C924 VTAIL.n783 B 0.010338f
C925 VTAIL.n784 B 0.010946f
C926 VTAIL.n785 B 0.024436f
C927 VTAIL.n786 B 0.051292f
C928 VTAIL.n787 B 0.010946f
C929 VTAIL.n788 B 0.010338f
C930 VTAIL.n789 B 0.043681f
C931 VTAIL.n790 B 0.02851f
C932 VTAIL.n791 B 1.65197f
C933 VP.n0 B 0.031042f
C934 VP.t6 B 3.03112f
C935 VP.n1 B 0.033062f
C936 VP.n2 B 0.016503f
C937 VP.n3 B 0.030758f
C938 VP.n4 B 0.016503f
C939 VP.t2 B 3.03112f
C940 VP.n5 B 0.030758f
C941 VP.n6 B 0.016503f
C942 VP.n7 B 0.030758f
C943 VP.n8 B 0.016503f
C944 VP.t0 B 3.03112f
C945 VP.n9 B 0.030758f
C946 VP.n10 B 0.016503f
C947 VP.n11 B 0.030758f
C948 VP.n12 B 0.031042f
C949 VP.t5 B 3.03112f
C950 VP.n13 B 0.033062f
C951 VP.n14 B 0.016503f
C952 VP.n15 B 0.030758f
C953 VP.n16 B 0.016503f
C954 VP.t1 B 3.03112f
C955 VP.n17 B 0.030758f
C956 VP.n18 B 0.016503f
C957 VP.n19 B 0.030758f
C958 VP.t7 B 3.29629f
C959 VP.n20 B 1.05994f
C960 VP.t4 B 3.03112f
C961 VP.n21 B 1.10689f
C962 VP.n22 B 0.025442f
C963 VP.n23 B 0.214563f
C964 VP.n24 B 0.016503f
C965 VP.n25 B 0.016503f
C966 VP.n26 B 0.030758f
C967 VP.n27 B 0.024092f
C968 VP.n28 B 0.024092f
C969 VP.n29 B 0.016503f
C970 VP.n30 B 0.016503f
C971 VP.n31 B 0.016503f
C972 VP.n32 B 0.030758f
C973 VP.n33 B 0.025442f
C974 VP.n34 B 1.04519f
C975 VP.n35 B 0.020886f
C976 VP.n36 B 0.016503f
C977 VP.n37 B 0.016503f
C978 VP.n38 B 0.016503f
C979 VP.n39 B 0.030758f
C980 VP.n40 B 0.030289f
C981 VP.n41 B 0.01559f
C982 VP.n42 B 0.016503f
C983 VP.n43 B 0.016503f
C984 VP.n44 B 0.016503f
C985 VP.n45 B 0.030758f
C986 VP.n46 B 0.029998f
C987 VP.n47 B 1.119f
C988 VP.n48 B 1.25363f
C989 VP.n49 B 1.26335f
C990 VP.t3 B 3.03112f
C991 VP.n50 B 1.119f
C992 VP.n51 B 0.029998f
C993 VP.n52 B 0.031042f
C994 VP.n53 B 0.016503f
C995 VP.n54 B 0.016503f
C996 VP.n55 B 0.033062f
C997 VP.n56 B 0.01559f
C998 VP.n57 B 0.030289f
C999 VP.n58 B 0.016503f
C1000 VP.n59 B 0.016503f
C1001 VP.n60 B 0.016503f
C1002 VP.n61 B 0.030758f
C1003 VP.n62 B 0.020886f
C1004 VP.n63 B 1.04519f
C1005 VP.n64 B 0.025442f
C1006 VP.n65 B 0.016503f
C1007 VP.n66 B 0.016503f
C1008 VP.n67 B 0.016503f
C1009 VP.n68 B 0.030758f
C1010 VP.n69 B 0.024092f
C1011 VP.n70 B 0.024092f
C1012 VP.n71 B 0.016503f
C1013 VP.n72 B 0.016503f
C1014 VP.n73 B 0.016503f
C1015 VP.n74 B 0.030758f
C1016 VP.n75 B 0.025442f
C1017 VP.n76 B 1.04519f
C1018 VP.n77 B 0.020886f
C1019 VP.n78 B 0.016503f
C1020 VP.n79 B 0.016503f
C1021 VP.n80 B 0.016503f
C1022 VP.n81 B 0.030758f
C1023 VP.n82 B 0.030289f
C1024 VP.n83 B 0.01559f
C1025 VP.n84 B 0.016503f
C1026 VP.n85 B 0.016503f
C1027 VP.n86 B 0.016503f
C1028 VP.n87 B 0.030758f
C1029 VP.n88 B 0.029998f
C1030 VP.n89 B 1.119f
C1031 VP.n90 B 0.048668f
.ends

