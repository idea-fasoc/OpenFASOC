* NGSPICE file created from diff_pair_sample_0574.ext - technology: sky130A

.subckt diff_pair_sample_0574 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VN.t0 VDD2.t2 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=3.0723 pd=18.95 as=3.0723 ps=18.95 w=18.62 l=0.77
X1 VDD2.t4 VN.t1 VTAIL.t9 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=7.2618 pd=38.02 as=3.0723 ps=18.95 w=18.62 l=0.77
X2 VDD1.t5 VP.t0 VTAIL.t3 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=7.2618 pd=38.02 as=3.0723 ps=18.95 w=18.62 l=0.77
X3 VTAIL.t8 VN.t2 VDD2.t1 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=3.0723 pd=18.95 as=3.0723 ps=18.95 w=18.62 l=0.77
X4 VDD2.t3 VN.t3 VTAIL.t7 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=3.0723 pd=18.95 as=7.2618 ps=38.02 w=18.62 l=0.77
X5 VDD2.t5 VN.t4 VTAIL.t6 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=7.2618 pd=38.02 as=3.0723 ps=18.95 w=18.62 l=0.77
X6 VDD2.t0 VN.t5 VTAIL.t5 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=3.0723 pd=18.95 as=7.2618 ps=38.02 w=18.62 l=0.77
X7 VDD1.t4 VP.t1 VTAIL.t0 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=7.2618 pd=38.02 as=3.0723 ps=18.95 w=18.62 l=0.77
X8 VDD1.t3 VP.t2 VTAIL.t11 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=3.0723 pd=18.95 as=7.2618 ps=38.02 w=18.62 l=0.77
X9 B.t11 B.t9 B.t10 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=7.2618 pd=38.02 as=0 ps=0 w=18.62 l=0.77
X10 VDD1.t2 VP.t3 VTAIL.t2 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=3.0723 pd=18.95 as=7.2618 ps=38.02 w=18.62 l=0.77
X11 VTAIL.t1 VP.t4 VDD1.t1 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=3.0723 pd=18.95 as=3.0723 ps=18.95 w=18.62 l=0.77
X12 B.t8 B.t6 B.t7 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=7.2618 pd=38.02 as=0 ps=0 w=18.62 l=0.77
X13 B.t5 B.t3 B.t4 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=7.2618 pd=38.02 as=0 ps=0 w=18.62 l=0.77
X14 VTAIL.t4 VP.t5 VDD1.t0 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=3.0723 pd=18.95 as=3.0723 ps=18.95 w=18.62 l=0.77
X15 B.t2 B.t0 B.t1 w_n1850_n4692# sky130_fd_pr__pfet_01v8 ad=7.2618 pd=38.02 as=0 ps=0 w=18.62 l=0.77
R0 VN.n1 VN.t4 656.734
R1 VN.n7 VN.t5 656.734
R2 VN.n2 VN.t0 633.799
R3 VN.n4 VN.t3 633.799
R4 VN.n8 VN.t2 633.799
R5 VN.n10 VN.t1 633.799
R6 VN.n5 VN.n4 161.3
R7 VN.n11 VN.n10 161.3
R8 VN.n9 VN.n6 161.3
R9 VN.n3 VN.n0 161.3
R10 VN VN.n11 46.9418
R11 VN.n7 VN.n6 44.8791
R12 VN.n1 VN.n0 44.8791
R13 VN.n4 VN.n3 31.4035
R14 VN.n10 VN.n9 31.4035
R15 VN.n2 VN.n1 18.8496
R16 VN.n8 VN.n7 18.8496
R17 VN.n3 VN.n2 16.7975
R18 VN.n9 VN.n8 16.7975
R19 VN.n11 VN.n6 0.189894
R20 VN.n5 VN.n0 0.189894
R21 VN VN.n5 0.0516364
R22 VDD2.n1 VDD2.t5 71.3218
R23 VDD2.n2 VDD2.t4 70.6661
R24 VDD2.n1 VDD2.n0 69.1019
R25 VDD2 VDD2.n3 69.0991
R26 VDD2.n2 VDD2.n1 42.8489
R27 VDD2.n3 VDD2.t1 1.7462
R28 VDD2.n3 VDD2.t0 1.7462
R29 VDD2.n0 VDD2.t2 1.7462
R30 VDD2.n0 VDD2.t3 1.7462
R31 VDD2 VDD2.n2 0.769897
R32 VTAIL.n7 VTAIL.t5 53.9873
R33 VTAIL.n10 VTAIL.t11 53.9871
R34 VTAIL.n11 VTAIL.t7 53.9871
R35 VTAIL.n2 VTAIL.t2 53.9871
R36 VTAIL.n9 VTAIL.n8 52.2416
R37 VTAIL.n6 VTAIL.n5 52.2416
R38 VTAIL.n1 VTAIL.n0 52.2414
R39 VTAIL.n4 VTAIL.n3 52.2414
R40 VTAIL.n6 VTAIL.n4 30.3152
R41 VTAIL.n11 VTAIL.n10 29.3669
R42 VTAIL.n0 VTAIL.t6 1.7462
R43 VTAIL.n0 VTAIL.t10 1.7462
R44 VTAIL.n3 VTAIL.t3 1.7462
R45 VTAIL.n3 VTAIL.t4 1.7462
R46 VTAIL.n8 VTAIL.t0 1.7462
R47 VTAIL.n8 VTAIL.t1 1.7462
R48 VTAIL.n5 VTAIL.t9 1.7462
R49 VTAIL.n5 VTAIL.t8 1.7462
R50 VTAIL.n7 VTAIL.n6 0.948776
R51 VTAIL.n10 VTAIL.n9 0.948776
R52 VTAIL.n4 VTAIL.n2 0.948776
R53 VTAIL.n9 VTAIL.n7 0.944465
R54 VTAIL.n2 VTAIL.n1 0.944465
R55 VTAIL VTAIL.n11 0.653517
R56 VTAIL VTAIL.n1 0.295759
R57 VP.n3 VP.t1 656.734
R58 VP.n8 VP.t0 633.799
R59 VP.n12 VP.t5 633.799
R60 VP.n14 VP.t3 633.799
R61 VP.n6 VP.t2 633.799
R62 VP.n4 VP.t4 633.799
R63 VP.n15 VP.n14 161.3
R64 VP.n5 VP.n2 161.3
R65 VP.n7 VP.n6 161.3
R66 VP.n13 VP.n0 161.3
R67 VP.n12 VP.n11 161.3
R68 VP.n10 VP.n1 161.3
R69 VP.n9 VP.n8 161.3
R70 VP.n9 VP.n7 46.5611
R71 VP.n3 VP.n2 44.8791
R72 VP.n8 VP.n1 31.4035
R73 VP.n14 VP.n13 31.4035
R74 VP.n6 VP.n5 31.4035
R75 VP.n4 VP.n3 18.8496
R76 VP.n12 VP.n1 16.7975
R77 VP.n13 VP.n12 16.7975
R78 VP.n5 VP.n4 16.7975
R79 VP.n7 VP.n2 0.189894
R80 VP.n10 VP.n9 0.189894
R81 VP.n11 VP.n10 0.189894
R82 VP.n11 VP.n0 0.189894
R83 VP.n15 VP.n0 0.189894
R84 VP VP.n15 0.0516364
R85 VDD1 VDD1.t4 71.4355
R86 VDD1.n1 VDD1.t5 71.3218
R87 VDD1.n1 VDD1.n0 69.1019
R88 VDD1.n3 VDD1.n2 68.9202
R89 VDD1.n3 VDD1.n1 43.9061
R90 VDD1.n2 VDD1.t1 1.7462
R91 VDD1.n2 VDD1.t3 1.7462
R92 VDD1.n0 VDD1.t0 1.7462
R93 VDD1.n0 VDD1.t2 1.7462
R94 VDD1 VDD1.n3 0.179379
R95 B.n136 B.t6 784.965
R96 B.n142 B.t0 784.965
R97 B.n44 B.t3 784.965
R98 B.n50 B.t9 784.965
R99 B.n480 B.n479 585
R100 B.n481 B.n82 585
R101 B.n483 B.n482 585
R102 B.n484 B.n81 585
R103 B.n486 B.n485 585
R104 B.n487 B.n80 585
R105 B.n489 B.n488 585
R106 B.n490 B.n79 585
R107 B.n492 B.n491 585
R108 B.n493 B.n78 585
R109 B.n495 B.n494 585
R110 B.n496 B.n77 585
R111 B.n498 B.n497 585
R112 B.n499 B.n76 585
R113 B.n501 B.n500 585
R114 B.n502 B.n75 585
R115 B.n504 B.n503 585
R116 B.n505 B.n74 585
R117 B.n507 B.n506 585
R118 B.n508 B.n73 585
R119 B.n510 B.n509 585
R120 B.n511 B.n72 585
R121 B.n513 B.n512 585
R122 B.n514 B.n71 585
R123 B.n516 B.n515 585
R124 B.n517 B.n70 585
R125 B.n519 B.n518 585
R126 B.n520 B.n69 585
R127 B.n522 B.n521 585
R128 B.n523 B.n68 585
R129 B.n525 B.n524 585
R130 B.n526 B.n67 585
R131 B.n528 B.n527 585
R132 B.n529 B.n66 585
R133 B.n531 B.n530 585
R134 B.n532 B.n65 585
R135 B.n534 B.n533 585
R136 B.n535 B.n64 585
R137 B.n537 B.n536 585
R138 B.n538 B.n63 585
R139 B.n540 B.n539 585
R140 B.n541 B.n62 585
R141 B.n543 B.n542 585
R142 B.n544 B.n61 585
R143 B.n546 B.n545 585
R144 B.n547 B.n60 585
R145 B.n549 B.n548 585
R146 B.n550 B.n59 585
R147 B.n552 B.n551 585
R148 B.n553 B.n58 585
R149 B.n555 B.n554 585
R150 B.n556 B.n57 585
R151 B.n558 B.n557 585
R152 B.n559 B.n56 585
R153 B.n561 B.n560 585
R154 B.n562 B.n55 585
R155 B.n564 B.n563 585
R156 B.n565 B.n54 585
R157 B.n567 B.n566 585
R158 B.n568 B.n53 585
R159 B.n570 B.n569 585
R160 B.n572 B.n571 585
R161 B.n573 B.n49 585
R162 B.n575 B.n574 585
R163 B.n576 B.n48 585
R164 B.n578 B.n577 585
R165 B.n579 B.n47 585
R166 B.n581 B.n580 585
R167 B.n582 B.n46 585
R168 B.n584 B.n583 585
R169 B.n585 B.n43 585
R170 B.n588 B.n587 585
R171 B.n589 B.n42 585
R172 B.n591 B.n590 585
R173 B.n592 B.n41 585
R174 B.n594 B.n593 585
R175 B.n595 B.n40 585
R176 B.n597 B.n596 585
R177 B.n598 B.n39 585
R178 B.n600 B.n599 585
R179 B.n601 B.n38 585
R180 B.n603 B.n602 585
R181 B.n604 B.n37 585
R182 B.n606 B.n605 585
R183 B.n607 B.n36 585
R184 B.n609 B.n608 585
R185 B.n610 B.n35 585
R186 B.n612 B.n611 585
R187 B.n613 B.n34 585
R188 B.n615 B.n614 585
R189 B.n616 B.n33 585
R190 B.n618 B.n617 585
R191 B.n619 B.n32 585
R192 B.n621 B.n620 585
R193 B.n622 B.n31 585
R194 B.n624 B.n623 585
R195 B.n625 B.n30 585
R196 B.n627 B.n626 585
R197 B.n628 B.n29 585
R198 B.n630 B.n629 585
R199 B.n631 B.n28 585
R200 B.n633 B.n632 585
R201 B.n634 B.n27 585
R202 B.n636 B.n635 585
R203 B.n637 B.n26 585
R204 B.n639 B.n638 585
R205 B.n640 B.n25 585
R206 B.n642 B.n641 585
R207 B.n643 B.n24 585
R208 B.n645 B.n644 585
R209 B.n646 B.n23 585
R210 B.n648 B.n647 585
R211 B.n649 B.n22 585
R212 B.n651 B.n650 585
R213 B.n652 B.n21 585
R214 B.n654 B.n653 585
R215 B.n655 B.n20 585
R216 B.n657 B.n656 585
R217 B.n658 B.n19 585
R218 B.n660 B.n659 585
R219 B.n661 B.n18 585
R220 B.n663 B.n662 585
R221 B.n664 B.n17 585
R222 B.n666 B.n665 585
R223 B.n667 B.n16 585
R224 B.n669 B.n668 585
R225 B.n670 B.n15 585
R226 B.n672 B.n671 585
R227 B.n673 B.n14 585
R228 B.n675 B.n674 585
R229 B.n676 B.n13 585
R230 B.n678 B.n677 585
R231 B.n478 B.n83 585
R232 B.n477 B.n476 585
R233 B.n475 B.n84 585
R234 B.n474 B.n473 585
R235 B.n472 B.n85 585
R236 B.n471 B.n470 585
R237 B.n469 B.n86 585
R238 B.n468 B.n467 585
R239 B.n466 B.n87 585
R240 B.n465 B.n464 585
R241 B.n463 B.n88 585
R242 B.n462 B.n461 585
R243 B.n460 B.n89 585
R244 B.n459 B.n458 585
R245 B.n457 B.n90 585
R246 B.n456 B.n455 585
R247 B.n454 B.n91 585
R248 B.n453 B.n452 585
R249 B.n451 B.n92 585
R250 B.n450 B.n449 585
R251 B.n448 B.n93 585
R252 B.n447 B.n446 585
R253 B.n445 B.n94 585
R254 B.n444 B.n443 585
R255 B.n442 B.n95 585
R256 B.n441 B.n440 585
R257 B.n439 B.n96 585
R258 B.n438 B.n437 585
R259 B.n436 B.n97 585
R260 B.n435 B.n434 585
R261 B.n433 B.n98 585
R262 B.n432 B.n431 585
R263 B.n430 B.n99 585
R264 B.n429 B.n428 585
R265 B.n427 B.n100 585
R266 B.n426 B.n425 585
R267 B.n424 B.n101 585
R268 B.n423 B.n422 585
R269 B.n421 B.n102 585
R270 B.n420 B.n419 585
R271 B.n418 B.n103 585
R272 B.n417 B.n416 585
R273 B.n415 B.n104 585
R274 B.n216 B.n215 585
R275 B.n217 B.n174 585
R276 B.n219 B.n218 585
R277 B.n220 B.n173 585
R278 B.n222 B.n221 585
R279 B.n223 B.n172 585
R280 B.n225 B.n224 585
R281 B.n226 B.n171 585
R282 B.n228 B.n227 585
R283 B.n229 B.n170 585
R284 B.n231 B.n230 585
R285 B.n232 B.n169 585
R286 B.n234 B.n233 585
R287 B.n235 B.n168 585
R288 B.n237 B.n236 585
R289 B.n238 B.n167 585
R290 B.n240 B.n239 585
R291 B.n241 B.n166 585
R292 B.n243 B.n242 585
R293 B.n244 B.n165 585
R294 B.n246 B.n245 585
R295 B.n247 B.n164 585
R296 B.n249 B.n248 585
R297 B.n250 B.n163 585
R298 B.n252 B.n251 585
R299 B.n253 B.n162 585
R300 B.n255 B.n254 585
R301 B.n256 B.n161 585
R302 B.n258 B.n257 585
R303 B.n259 B.n160 585
R304 B.n261 B.n260 585
R305 B.n262 B.n159 585
R306 B.n264 B.n263 585
R307 B.n265 B.n158 585
R308 B.n267 B.n266 585
R309 B.n268 B.n157 585
R310 B.n270 B.n269 585
R311 B.n271 B.n156 585
R312 B.n273 B.n272 585
R313 B.n274 B.n155 585
R314 B.n276 B.n275 585
R315 B.n277 B.n154 585
R316 B.n279 B.n278 585
R317 B.n280 B.n153 585
R318 B.n282 B.n281 585
R319 B.n283 B.n152 585
R320 B.n285 B.n284 585
R321 B.n286 B.n151 585
R322 B.n288 B.n287 585
R323 B.n289 B.n150 585
R324 B.n291 B.n290 585
R325 B.n292 B.n149 585
R326 B.n294 B.n293 585
R327 B.n295 B.n148 585
R328 B.n297 B.n296 585
R329 B.n298 B.n147 585
R330 B.n300 B.n299 585
R331 B.n301 B.n146 585
R332 B.n303 B.n302 585
R333 B.n304 B.n145 585
R334 B.n306 B.n305 585
R335 B.n308 B.n307 585
R336 B.n309 B.n141 585
R337 B.n311 B.n310 585
R338 B.n312 B.n140 585
R339 B.n314 B.n313 585
R340 B.n315 B.n139 585
R341 B.n317 B.n316 585
R342 B.n318 B.n138 585
R343 B.n320 B.n319 585
R344 B.n321 B.n135 585
R345 B.n324 B.n323 585
R346 B.n325 B.n134 585
R347 B.n327 B.n326 585
R348 B.n328 B.n133 585
R349 B.n330 B.n329 585
R350 B.n331 B.n132 585
R351 B.n333 B.n332 585
R352 B.n334 B.n131 585
R353 B.n336 B.n335 585
R354 B.n337 B.n130 585
R355 B.n339 B.n338 585
R356 B.n340 B.n129 585
R357 B.n342 B.n341 585
R358 B.n343 B.n128 585
R359 B.n345 B.n344 585
R360 B.n346 B.n127 585
R361 B.n348 B.n347 585
R362 B.n349 B.n126 585
R363 B.n351 B.n350 585
R364 B.n352 B.n125 585
R365 B.n354 B.n353 585
R366 B.n355 B.n124 585
R367 B.n357 B.n356 585
R368 B.n358 B.n123 585
R369 B.n360 B.n359 585
R370 B.n361 B.n122 585
R371 B.n363 B.n362 585
R372 B.n364 B.n121 585
R373 B.n366 B.n365 585
R374 B.n367 B.n120 585
R375 B.n369 B.n368 585
R376 B.n370 B.n119 585
R377 B.n372 B.n371 585
R378 B.n373 B.n118 585
R379 B.n375 B.n374 585
R380 B.n376 B.n117 585
R381 B.n378 B.n377 585
R382 B.n379 B.n116 585
R383 B.n381 B.n380 585
R384 B.n382 B.n115 585
R385 B.n384 B.n383 585
R386 B.n385 B.n114 585
R387 B.n387 B.n386 585
R388 B.n388 B.n113 585
R389 B.n390 B.n389 585
R390 B.n391 B.n112 585
R391 B.n393 B.n392 585
R392 B.n394 B.n111 585
R393 B.n396 B.n395 585
R394 B.n397 B.n110 585
R395 B.n399 B.n398 585
R396 B.n400 B.n109 585
R397 B.n402 B.n401 585
R398 B.n403 B.n108 585
R399 B.n405 B.n404 585
R400 B.n406 B.n107 585
R401 B.n408 B.n407 585
R402 B.n409 B.n106 585
R403 B.n411 B.n410 585
R404 B.n412 B.n105 585
R405 B.n414 B.n413 585
R406 B.n214 B.n175 585
R407 B.n213 B.n212 585
R408 B.n211 B.n176 585
R409 B.n210 B.n209 585
R410 B.n208 B.n177 585
R411 B.n207 B.n206 585
R412 B.n205 B.n178 585
R413 B.n204 B.n203 585
R414 B.n202 B.n179 585
R415 B.n201 B.n200 585
R416 B.n199 B.n180 585
R417 B.n198 B.n197 585
R418 B.n196 B.n181 585
R419 B.n195 B.n194 585
R420 B.n193 B.n182 585
R421 B.n192 B.n191 585
R422 B.n190 B.n183 585
R423 B.n189 B.n188 585
R424 B.n187 B.n184 585
R425 B.n186 B.n185 585
R426 B.n2 B.n0 585
R427 B.n709 B.n1 585
R428 B.n708 B.n707 585
R429 B.n706 B.n3 585
R430 B.n705 B.n704 585
R431 B.n703 B.n4 585
R432 B.n702 B.n701 585
R433 B.n700 B.n5 585
R434 B.n699 B.n698 585
R435 B.n697 B.n6 585
R436 B.n696 B.n695 585
R437 B.n694 B.n7 585
R438 B.n693 B.n692 585
R439 B.n691 B.n8 585
R440 B.n690 B.n689 585
R441 B.n688 B.n9 585
R442 B.n687 B.n686 585
R443 B.n685 B.n10 585
R444 B.n684 B.n683 585
R445 B.n682 B.n11 585
R446 B.n681 B.n680 585
R447 B.n679 B.n12 585
R448 B.n711 B.n710 585
R449 B.n216 B.n175 487.695
R450 B.n679 B.n678 487.695
R451 B.n415 B.n414 487.695
R452 B.n480 B.n83 487.695
R453 B.n212 B.n175 163.367
R454 B.n212 B.n211 163.367
R455 B.n211 B.n210 163.367
R456 B.n210 B.n177 163.367
R457 B.n206 B.n177 163.367
R458 B.n206 B.n205 163.367
R459 B.n205 B.n204 163.367
R460 B.n204 B.n179 163.367
R461 B.n200 B.n179 163.367
R462 B.n200 B.n199 163.367
R463 B.n199 B.n198 163.367
R464 B.n198 B.n181 163.367
R465 B.n194 B.n181 163.367
R466 B.n194 B.n193 163.367
R467 B.n193 B.n192 163.367
R468 B.n192 B.n183 163.367
R469 B.n188 B.n183 163.367
R470 B.n188 B.n187 163.367
R471 B.n187 B.n186 163.367
R472 B.n186 B.n2 163.367
R473 B.n710 B.n2 163.367
R474 B.n710 B.n709 163.367
R475 B.n709 B.n708 163.367
R476 B.n708 B.n3 163.367
R477 B.n704 B.n3 163.367
R478 B.n704 B.n703 163.367
R479 B.n703 B.n702 163.367
R480 B.n702 B.n5 163.367
R481 B.n698 B.n5 163.367
R482 B.n698 B.n697 163.367
R483 B.n697 B.n696 163.367
R484 B.n696 B.n7 163.367
R485 B.n692 B.n7 163.367
R486 B.n692 B.n691 163.367
R487 B.n691 B.n690 163.367
R488 B.n690 B.n9 163.367
R489 B.n686 B.n9 163.367
R490 B.n686 B.n685 163.367
R491 B.n685 B.n684 163.367
R492 B.n684 B.n11 163.367
R493 B.n680 B.n11 163.367
R494 B.n680 B.n679 163.367
R495 B.n217 B.n216 163.367
R496 B.n218 B.n217 163.367
R497 B.n218 B.n173 163.367
R498 B.n222 B.n173 163.367
R499 B.n223 B.n222 163.367
R500 B.n224 B.n223 163.367
R501 B.n224 B.n171 163.367
R502 B.n228 B.n171 163.367
R503 B.n229 B.n228 163.367
R504 B.n230 B.n229 163.367
R505 B.n230 B.n169 163.367
R506 B.n234 B.n169 163.367
R507 B.n235 B.n234 163.367
R508 B.n236 B.n235 163.367
R509 B.n236 B.n167 163.367
R510 B.n240 B.n167 163.367
R511 B.n241 B.n240 163.367
R512 B.n242 B.n241 163.367
R513 B.n242 B.n165 163.367
R514 B.n246 B.n165 163.367
R515 B.n247 B.n246 163.367
R516 B.n248 B.n247 163.367
R517 B.n248 B.n163 163.367
R518 B.n252 B.n163 163.367
R519 B.n253 B.n252 163.367
R520 B.n254 B.n253 163.367
R521 B.n254 B.n161 163.367
R522 B.n258 B.n161 163.367
R523 B.n259 B.n258 163.367
R524 B.n260 B.n259 163.367
R525 B.n260 B.n159 163.367
R526 B.n264 B.n159 163.367
R527 B.n265 B.n264 163.367
R528 B.n266 B.n265 163.367
R529 B.n266 B.n157 163.367
R530 B.n270 B.n157 163.367
R531 B.n271 B.n270 163.367
R532 B.n272 B.n271 163.367
R533 B.n272 B.n155 163.367
R534 B.n276 B.n155 163.367
R535 B.n277 B.n276 163.367
R536 B.n278 B.n277 163.367
R537 B.n278 B.n153 163.367
R538 B.n282 B.n153 163.367
R539 B.n283 B.n282 163.367
R540 B.n284 B.n283 163.367
R541 B.n284 B.n151 163.367
R542 B.n288 B.n151 163.367
R543 B.n289 B.n288 163.367
R544 B.n290 B.n289 163.367
R545 B.n290 B.n149 163.367
R546 B.n294 B.n149 163.367
R547 B.n295 B.n294 163.367
R548 B.n296 B.n295 163.367
R549 B.n296 B.n147 163.367
R550 B.n300 B.n147 163.367
R551 B.n301 B.n300 163.367
R552 B.n302 B.n301 163.367
R553 B.n302 B.n145 163.367
R554 B.n306 B.n145 163.367
R555 B.n307 B.n306 163.367
R556 B.n307 B.n141 163.367
R557 B.n311 B.n141 163.367
R558 B.n312 B.n311 163.367
R559 B.n313 B.n312 163.367
R560 B.n313 B.n139 163.367
R561 B.n317 B.n139 163.367
R562 B.n318 B.n317 163.367
R563 B.n319 B.n318 163.367
R564 B.n319 B.n135 163.367
R565 B.n324 B.n135 163.367
R566 B.n325 B.n324 163.367
R567 B.n326 B.n325 163.367
R568 B.n326 B.n133 163.367
R569 B.n330 B.n133 163.367
R570 B.n331 B.n330 163.367
R571 B.n332 B.n331 163.367
R572 B.n332 B.n131 163.367
R573 B.n336 B.n131 163.367
R574 B.n337 B.n336 163.367
R575 B.n338 B.n337 163.367
R576 B.n338 B.n129 163.367
R577 B.n342 B.n129 163.367
R578 B.n343 B.n342 163.367
R579 B.n344 B.n343 163.367
R580 B.n344 B.n127 163.367
R581 B.n348 B.n127 163.367
R582 B.n349 B.n348 163.367
R583 B.n350 B.n349 163.367
R584 B.n350 B.n125 163.367
R585 B.n354 B.n125 163.367
R586 B.n355 B.n354 163.367
R587 B.n356 B.n355 163.367
R588 B.n356 B.n123 163.367
R589 B.n360 B.n123 163.367
R590 B.n361 B.n360 163.367
R591 B.n362 B.n361 163.367
R592 B.n362 B.n121 163.367
R593 B.n366 B.n121 163.367
R594 B.n367 B.n366 163.367
R595 B.n368 B.n367 163.367
R596 B.n368 B.n119 163.367
R597 B.n372 B.n119 163.367
R598 B.n373 B.n372 163.367
R599 B.n374 B.n373 163.367
R600 B.n374 B.n117 163.367
R601 B.n378 B.n117 163.367
R602 B.n379 B.n378 163.367
R603 B.n380 B.n379 163.367
R604 B.n380 B.n115 163.367
R605 B.n384 B.n115 163.367
R606 B.n385 B.n384 163.367
R607 B.n386 B.n385 163.367
R608 B.n386 B.n113 163.367
R609 B.n390 B.n113 163.367
R610 B.n391 B.n390 163.367
R611 B.n392 B.n391 163.367
R612 B.n392 B.n111 163.367
R613 B.n396 B.n111 163.367
R614 B.n397 B.n396 163.367
R615 B.n398 B.n397 163.367
R616 B.n398 B.n109 163.367
R617 B.n402 B.n109 163.367
R618 B.n403 B.n402 163.367
R619 B.n404 B.n403 163.367
R620 B.n404 B.n107 163.367
R621 B.n408 B.n107 163.367
R622 B.n409 B.n408 163.367
R623 B.n410 B.n409 163.367
R624 B.n410 B.n105 163.367
R625 B.n414 B.n105 163.367
R626 B.n416 B.n415 163.367
R627 B.n416 B.n103 163.367
R628 B.n420 B.n103 163.367
R629 B.n421 B.n420 163.367
R630 B.n422 B.n421 163.367
R631 B.n422 B.n101 163.367
R632 B.n426 B.n101 163.367
R633 B.n427 B.n426 163.367
R634 B.n428 B.n427 163.367
R635 B.n428 B.n99 163.367
R636 B.n432 B.n99 163.367
R637 B.n433 B.n432 163.367
R638 B.n434 B.n433 163.367
R639 B.n434 B.n97 163.367
R640 B.n438 B.n97 163.367
R641 B.n439 B.n438 163.367
R642 B.n440 B.n439 163.367
R643 B.n440 B.n95 163.367
R644 B.n444 B.n95 163.367
R645 B.n445 B.n444 163.367
R646 B.n446 B.n445 163.367
R647 B.n446 B.n93 163.367
R648 B.n450 B.n93 163.367
R649 B.n451 B.n450 163.367
R650 B.n452 B.n451 163.367
R651 B.n452 B.n91 163.367
R652 B.n456 B.n91 163.367
R653 B.n457 B.n456 163.367
R654 B.n458 B.n457 163.367
R655 B.n458 B.n89 163.367
R656 B.n462 B.n89 163.367
R657 B.n463 B.n462 163.367
R658 B.n464 B.n463 163.367
R659 B.n464 B.n87 163.367
R660 B.n468 B.n87 163.367
R661 B.n469 B.n468 163.367
R662 B.n470 B.n469 163.367
R663 B.n470 B.n85 163.367
R664 B.n474 B.n85 163.367
R665 B.n475 B.n474 163.367
R666 B.n476 B.n475 163.367
R667 B.n476 B.n83 163.367
R668 B.n678 B.n13 163.367
R669 B.n674 B.n13 163.367
R670 B.n674 B.n673 163.367
R671 B.n673 B.n672 163.367
R672 B.n672 B.n15 163.367
R673 B.n668 B.n15 163.367
R674 B.n668 B.n667 163.367
R675 B.n667 B.n666 163.367
R676 B.n666 B.n17 163.367
R677 B.n662 B.n17 163.367
R678 B.n662 B.n661 163.367
R679 B.n661 B.n660 163.367
R680 B.n660 B.n19 163.367
R681 B.n656 B.n19 163.367
R682 B.n656 B.n655 163.367
R683 B.n655 B.n654 163.367
R684 B.n654 B.n21 163.367
R685 B.n650 B.n21 163.367
R686 B.n650 B.n649 163.367
R687 B.n649 B.n648 163.367
R688 B.n648 B.n23 163.367
R689 B.n644 B.n23 163.367
R690 B.n644 B.n643 163.367
R691 B.n643 B.n642 163.367
R692 B.n642 B.n25 163.367
R693 B.n638 B.n25 163.367
R694 B.n638 B.n637 163.367
R695 B.n637 B.n636 163.367
R696 B.n636 B.n27 163.367
R697 B.n632 B.n27 163.367
R698 B.n632 B.n631 163.367
R699 B.n631 B.n630 163.367
R700 B.n630 B.n29 163.367
R701 B.n626 B.n29 163.367
R702 B.n626 B.n625 163.367
R703 B.n625 B.n624 163.367
R704 B.n624 B.n31 163.367
R705 B.n620 B.n31 163.367
R706 B.n620 B.n619 163.367
R707 B.n619 B.n618 163.367
R708 B.n618 B.n33 163.367
R709 B.n614 B.n33 163.367
R710 B.n614 B.n613 163.367
R711 B.n613 B.n612 163.367
R712 B.n612 B.n35 163.367
R713 B.n608 B.n35 163.367
R714 B.n608 B.n607 163.367
R715 B.n607 B.n606 163.367
R716 B.n606 B.n37 163.367
R717 B.n602 B.n37 163.367
R718 B.n602 B.n601 163.367
R719 B.n601 B.n600 163.367
R720 B.n600 B.n39 163.367
R721 B.n596 B.n39 163.367
R722 B.n596 B.n595 163.367
R723 B.n595 B.n594 163.367
R724 B.n594 B.n41 163.367
R725 B.n590 B.n41 163.367
R726 B.n590 B.n589 163.367
R727 B.n589 B.n588 163.367
R728 B.n588 B.n43 163.367
R729 B.n583 B.n43 163.367
R730 B.n583 B.n582 163.367
R731 B.n582 B.n581 163.367
R732 B.n581 B.n47 163.367
R733 B.n577 B.n47 163.367
R734 B.n577 B.n576 163.367
R735 B.n576 B.n575 163.367
R736 B.n575 B.n49 163.367
R737 B.n571 B.n49 163.367
R738 B.n571 B.n570 163.367
R739 B.n570 B.n53 163.367
R740 B.n566 B.n53 163.367
R741 B.n566 B.n565 163.367
R742 B.n565 B.n564 163.367
R743 B.n564 B.n55 163.367
R744 B.n560 B.n55 163.367
R745 B.n560 B.n559 163.367
R746 B.n559 B.n558 163.367
R747 B.n558 B.n57 163.367
R748 B.n554 B.n57 163.367
R749 B.n554 B.n553 163.367
R750 B.n553 B.n552 163.367
R751 B.n552 B.n59 163.367
R752 B.n548 B.n59 163.367
R753 B.n548 B.n547 163.367
R754 B.n547 B.n546 163.367
R755 B.n546 B.n61 163.367
R756 B.n542 B.n61 163.367
R757 B.n542 B.n541 163.367
R758 B.n541 B.n540 163.367
R759 B.n540 B.n63 163.367
R760 B.n536 B.n63 163.367
R761 B.n536 B.n535 163.367
R762 B.n535 B.n534 163.367
R763 B.n534 B.n65 163.367
R764 B.n530 B.n65 163.367
R765 B.n530 B.n529 163.367
R766 B.n529 B.n528 163.367
R767 B.n528 B.n67 163.367
R768 B.n524 B.n67 163.367
R769 B.n524 B.n523 163.367
R770 B.n523 B.n522 163.367
R771 B.n522 B.n69 163.367
R772 B.n518 B.n69 163.367
R773 B.n518 B.n517 163.367
R774 B.n517 B.n516 163.367
R775 B.n516 B.n71 163.367
R776 B.n512 B.n71 163.367
R777 B.n512 B.n511 163.367
R778 B.n511 B.n510 163.367
R779 B.n510 B.n73 163.367
R780 B.n506 B.n73 163.367
R781 B.n506 B.n505 163.367
R782 B.n505 B.n504 163.367
R783 B.n504 B.n75 163.367
R784 B.n500 B.n75 163.367
R785 B.n500 B.n499 163.367
R786 B.n499 B.n498 163.367
R787 B.n498 B.n77 163.367
R788 B.n494 B.n77 163.367
R789 B.n494 B.n493 163.367
R790 B.n493 B.n492 163.367
R791 B.n492 B.n79 163.367
R792 B.n488 B.n79 163.367
R793 B.n488 B.n487 163.367
R794 B.n487 B.n486 163.367
R795 B.n486 B.n81 163.367
R796 B.n482 B.n81 163.367
R797 B.n482 B.n481 163.367
R798 B.n481 B.n480 163.367
R799 B.n136 B.t8 132.52
R800 B.n50 B.t10 132.52
R801 B.n142 B.t2 132.496
R802 B.n44 B.t4 132.496
R803 B.n137 B.t7 111.188
R804 B.n51 B.t11 111.188
R805 B.n143 B.t1 111.163
R806 B.n45 B.t5 111.163
R807 B.n322 B.n137 59.5399
R808 B.n144 B.n143 59.5399
R809 B.n586 B.n45 59.5399
R810 B.n52 B.n51 59.5399
R811 B.n677 B.n12 31.6883
R812 B.n479 B.n478 31.6883
R813 B.n413 B.n104 31.6883
R814 B.n215 B.n214 31.6883
R815 B.n137 B.n136 21.3338
R816 B.n143 B.n142 21.3338
R817 B.n45 B.n44 21.3338
R818 B.n51 B.n50 21.3338
R819 B B.n711 18.0485
R820 B.n677 B.n676 10.6151
R821 B.n676 B.n675 10.6151
R822 B.n675 B.n14 10.6151
R823 B.n671 B.n14 10.6151
R824 B.n671 B.n670 10.6151
R825 B.n670 B.n669 10.6151
R826 B.n669 B.n16 10.6151
R827 B.n665 B.n16 10.6151
R828 B.n665 B.n664 10.6151
R829 B.n664 B.n663 10.6151
R830 B.n663 B.n18 10.6151
R831 B.n659 B.n18 10.6151
R832 B.n659 B.n658 10.6151
R833 B.n658 B.n657 10.6151
R834 B.n657 B.n20 10.6151
R835 B.n653 B.n20 10.6151
R836 B.n653 B.n652 10.6151
R837 B.n652 B.n651 10.6151
R838 B.n651 B.n22 10.6151
R839 B.n647 B.n22 10.6151
R840 B.n647 B.n646 10.6151
R841 B.n646 B.n645 10.6151
R842 B.n645 B.n24 10.6151
R843 B.n641 B.n24 10.6151
R844 B.n641 B.n640 10.6151
R845 B.n640 B.n639 10.6151
R846 B.n639 B.n26 10.6151
R847 B.n635 B.n26 10.6151
R848 B.n635 B.n634 10.6151
R849 B.n634 B.n633 10.6151
R850 B.n633 B.n28 10.6151
R851 B.n629 B.n28 10.6151
R852 B.n629 B.n628 10.6151
R853 B.n628 B.n627 10.6151
R854 B.n627 B.n30 10.6151
R855 B.n623 B.n30 10.6151
R856 B.n623 B.n622 10.6151
R857 B.n622 B.n621 10.6151
R858 B.n621 B.n32 10.6151
R859 B.n617 B.n32 10.6151
R860 B.n617 B.n616 10.6151
R861 B.n616 B.n615 10.6151
R862 B.n615 B.n34 10.6151
R863 B.n611 B.n34 10.6151
R864 B.n611 B.n610 10.6151
R865 B.n610 B.n609 10.6151
R866 B.n609 B.n36 10.6151
R867 B.n605 B.n36 10.6151
R868 B.n605 B.n604 10.6151
R869 B.n604 B.n603 10.6151
R870 B.n603 B.n38 10.6151
R871 B.n599 B.n38 10.6151
R872 B.n599 B.n598 10.6151
R873 B.n598 B.n597 10.6151
R874 B.n597 B.n40 10.6151
R875 B.n593 B.n40 10.6151
R876 B.n593 B.n592 10.6151
R877 B.n592 B.n591 10.6151
R878 B.n591 B.n42 10.6151
R879 B.n587 B.n42 10.6151
R880 B.n585 B.n584 10.6151
R881 B.n584 B.n46 10.6151
R882 B.n580 B.n46 10.6151
R883 B.n580 B.n579 10.6151
R884 B.n579 B.n578 10.6151
R885 B.n578 B.n48 10.6151
R886 B.n574 B.n48 10.6151
R887 B.n574 B.n573 10.6151
R888 B.n573 B.n572 10.6151
R889 B.n569 B.n568 10.6151
R890 B.n568 B.n567 10.6151
R891 B.n567 B.n54 10.6151
R892 B.n563 B.n54 10.6151
R893 B.n563 B.n562 10.6151
R894 B.n562 B.n561 10.6151
R895 B.n561 B.n56 10.6151
R896 B.n557 B.n56 10.6151
R897 B.n557 B.n556 10.6151
R898 B.n556 B.n555 10.6151
R899 B.n555 B.n58 10.6151
R900 B.n551 B.n58 10.6151
R901 B.n551 B.n550 10.6151
R902 B.n550 B.n549 10.6151
R903 B.n549 B.n60 10.6151
R904 B.n545 B.n60 10.6151
R905 B.n545 B.n544 10.6151
R906 B.n544 B.n543 10.6151
R907 B.n543 B.n62 10.6151
R908 B.n539 B.n62 10.6151
R909 B.n539 B.n538 10.6151
R910 B.n538 B.n537 10.6151
R911 B.n537 B.n64 10.6151
R912 B.n533 B.n64 10.6151
R913 B.n533 B.n532 10.6151
R914 B.n532 B.n531 10.6151
R915 B.n531 B.n66 10.6151
R916 B.n527 B.n66 10.6151
R917 B.n527 B.n526 10.6151
R918 B.n526 B.n525 10.6151
R919 B.n525 B.n68 10.6151
R920 B.n521 B.n68 10.6151
R921 B.n521 B.n520 10.6151
R922 B.n520 B.n519 10.6151
R923 B.n519 B.n70 10.6151
R924 B.n515 B.n70 10.6151
R925 B.n515 B.n514 10.6151
R926 B.n514 B.n513 10.6151
R927 B.n513 B.n72 10.6151
R928 B.n509 B.n72 10.6151
R929 B.n509 B.n508 10.6151
R930 B.n508 B.n507 10.6151
R931 B.n507 B.n74 10.6151
R932 B.n503 B.n74 10.6151
R933 B.n503 B.n502 10.6151
R934 B.n502 B.n501 10.6151
R935 B.n501 B.n76 10.6151
R936 B.n497 B.n76 10.6151
R937 B.n497 B.n496 10.6151
R938 B.n496 B.n495 10.6151
R939 B.n495 B.n78 10.6151
R940 B.n491 B.n78 10.6151
R941 B.n491 B.n490 10.6151
R942 B.n490 B.n489 10.6151
R943 B.n489 B.n80 10.6151
R944 B.n485 B.n80 10.6151
R945 B.n485 B.n484 10.6151
R946 B.n484 B.n483 10.6151
R947 B.n483 B.n82 10.6151
R948 B.n479 B.n82 10.6151
R949 B.n417 B.n104 10.6151
R950 B.n418 B.n417 10.6151
R951 B.n419 B.n418 10.6151
R952 B.n419 B.n102 10.6151
R953 B.n423 B.n102 10.6151
R954 B.n424 B.n423 10.6151
R955 B.n425 B.n424 10.6151
R956 B.n425 B.n100 10.6151
R957 B.n429 B.n100 10.6151
R958 B.n430 B.n429 10.6151
R959 B.n431 B.n430 10.6151
R960 B.n431 B.n98 10.6151
R961 B.n435 B.n98 10.6151
R962 B.n436 B.n435 10.6151
R963 B.n437 B.n436 10.6151
R964 B.n437 B.n96 10.6151
R965 B.n441 B.n96 10.6151
R966 B.n442 B.n441 10.6151
R967 B.n443 B.n442 10.6151
R968 B.n443 B.n94 10.6151
R969 B.n447 B.n94 10.6151
R970 B.n448 B.n447 10.6151
R971 B.n449 B.n448 10.6151
R972 B.n449 B.n92 10.6151
R973 B.n453 B.n92 10.6151
R974 B.n454 B.n453 10.6151
R975 B.n455 B.n454 10.6151
R976 B.n455 B.n90 10.6151
R977 B.n459 B.n90 10.6151
R978 B.n460 B.n459 10.6151
R979 B.n461 B.n460 10.6151
R980 B.n461 B.n88 10.6151
R981 B.n465 B.n88 10.6151
R982 B.n466 B.n465 10.6151
R983 B.n467 B.n466 10.6151
R984 B.n467 B.n86 10.6151
R985 B.n471 B.n86 10.6151
R986 B.n472 B.n471 10.6151
R987 B.n473 B.n472 10.6151
R988 B.n473 B.n84 10.6151
R989 B.n477 B.n84 10.6151
R990 B.n478 B.n477 10.6151
R991 B.n215 B.n174 10.6151
R992 B.n219 B.n174 10.6151
R993 B.n220 B.n219 10.6151
R994 B.n221 B.n220 10.6151
R995 B.n221 B.n172 10.6151
R996 B.n225 B.n172 10.6151
R997 B.n226 B.n225 10.6151
R998 B.n227 B.n226 10.6151
R999 B.n227 B.n170 10.6151
R1000 B.n231 B.n170 10.6151
R1001 B.n232 B.n231 10.6151
R1002 B.n233 B.n232 10.6151
R1003 B.n233 B.n168 10.6151
R1004 B.n237 B.n168 10.6151
R1005 B.n238 B.n237 10.6151
R1006 B.n239 B.n238 10.6151
R1007 B.n239 B.n166 10.6151
R1008 B.n243 B.n166 10.6151
R1009 B.n244 B.n243 10.6151
R1010 B.n245 B.n244 10.6151
R1011 B.n245 B.n164 10.6151
R1012 B.n249 B.n164 10.6151
R1013 B.n250 B.n249 10.6151
R1014 B.n251 B.n250 10.6151
R1015 B.n251 B.n162 10.6151
R1016 B.n255 B.n162 10.6151
R1017 B.n256 B.n255 10.6151
R1018 B.n257 B.n256 10.6151
R1019 B.n257 B.n160 10.6151
R1020 B.n261 B.n160 10.6151
R1021 B.n262 B.n261 10.6151
R1022 B.n263 B.n262 10.6151
R1023 B.n263 B.n158 10.6151
R1024 B.n267 B.n158 10.6151
R1025 B.n268 B.n267 10.6151
R1026 B.n269 B.n268 10.6151
R1027 B.n269 B.n156 10.6151
R1028 B.n273 B.n156 10.6151
R1029 B.n274 B.n273 10.6151
R1030 B.n275 B.n274 10.6151
R1031 B.n275 B.n154 10.6151
R1032 B.n279 B.n154 10.6151
R1033 B.n280 B.n279 10.6151
R1034 B.n281 B.n280 10.6151
R1035 B.n281 B.n152 10.6151
R1036 B.n285 B.n152 10.6151
R1037 B.n286 B.n285 10.6151
R1038 B.n287 B.n286 10.6151
R1039 B.n287 B.n150 10.6151
R1040 B.n291 B.n150 10.6151
R1041 B.n292 B.n291 10.6151
R1042 B.n293 B.n292 10.6151
R1043 B.n293 B.n148 10.6151
R1044 B.n297 B.n148 10.6151
R1045 B.n298 B.n297 10.6151
R1046 B.n299 B.n298 10.6151
R1047 B.n299 B.n146 10.6151
R1048 B.n303 B.n146 10.6151
R1049 B.n304 B.n303 10.6151
R1050 B.n305 B.n304 10.6151
R1051 B.n309 B.n308 10.6151
R1052 B.n310 B.n309 10.6151
R1053 B.n310 B.n140 10.6151
R1054 B.n314 B.n140 10.6151
R1055 B.n315 B.n314 10.6151
R1056 B.n316 B.n315 10.6151
R1057 B.n316 B.n138 10.6151
R1058 B.n320 B.n138 10.6151
R1059 B.n321 B.n320 10.6151
R1060 B.n323 B.n134 10.6151
R1061 B.n327 B.n134 10.6151
R1062 B.n328 B.n327 10.6151
R1063 B.n329 B.n328 10.6151
R1064 B.n329 B.n132 10.6151
R1065 B.n333 B.n132 10.6151
R1066 B.n334 B.n333 10.6151
R1067 B.n335 B.n334 10.6151
R1068 B.n335 B.n130 10.6151
R1069 B.n339 B.n130 10.6151
R1070 B.n340 B.n339 10.6151
R1071 B.n341 B.n340 10.6151
R1072 B.n341 B.n128 10.6151
R1073 B.n345 B.n128 10.6151
R1074 B.n346 B.n345 10.6151
R1075 B.n347 B.n346 10.6151
R1076 B.n347 B.n126 10.6151
R1077 B.n351 B.n126 10.6151
R1078 B.n352 B.n351 10.6151
R1079 B.n353 B.n352 10.6151
R1080 B.n353 B.n124 10.6151
R1081 B.n357 B.n124 10.6151
R1082 B.n358 B.n357 10.6151
R1083 B.n359 B.n358 10.6151
R1084 B.n359 B.n122 10.6151
R1085 B.n363 B.n122 10.6151
R1086 B.n364 B.n363 10.6151
R1087 B.n365 B.n364 10.6151
R1088 B.n365 B.n120 10.6151
R1089 B.n369 B.n120 10.6151
R1090 B.n370 B.n369 10.6151
R1091 B.n371 B.n370 10.6151
R1092 B.n371 B.n118 10.6151
R1093 B.n375 B.n118 10.6151
R1094 B.n376 B.n375 10.6151
R1095 B.n377 B.n376 10.6151
R1096 B.n377 B.n116 10.6151
R1097 B.n381 B.n116 10.6151
R1098 B.n382 B.n381 10.6151
R1099 B.n383 B.n382 10.6151
R1100 B.n383 B.n114 10.6151
R1101 B.n387 B.n114 10.6151
R1102 B.n388 B.n387 10.6151
R1103 B.n389 B.n388 10.6151
R1104 B.n389 B.n112 10.6151
R1105 B.n393 B.n112 10.6151
R1106 B.n394 B.n393 10.6151
R1107 B.n395 B.n394 10.6151
R1108 B.n395 B.n110 10.6151
R1109 B.n399 B.n110 10.6151
R1110 B.n400 B.n399 10.6151
R1111 B.n401 B.n400 10.6151
R1112 B.n401 B.n108 10.6151
R1113 B.n405 B.n108 10.6151
R1114 B.n406 B.n405 10.6151
R1115 B.n407 B.n406 10.6151
R1116 B.n407 B.n106 10.6151
R1117 B.n411 B.n106 10.6151
R1118 B.n412 B.n411 10.6151
R1119 B.n413 B.n412 10.6151
R1120 B.n214 B.n213 10.6151
R1121 B.n213 B.n176 10.6151
R1122 B.n209 B.n176 10.6151
R1123 B.n209 B.n208 10.6151
R1124 B.n208 B.n207 10.6151
R1125 B.n207 B.n178 10.6151
R1126 B.n203 B.n178 10.6151
R1127 B.n203 B.n202 10.6151
R1128 B.n202 B.n201 10.6151
R1129 B.n201 B.n180 10.6151
R1130 B.n197 B.n180 10.6151
R1131 B.n197 B.n196 10.6151
R1132 B.n196 B.n195 10.6151
R1133 B.n195 B.n182 10.6151
R1134 B.n191 B.n182 10.6151
R1135 B.n191 B.n190 10.6151
R1136 B.n190 B.n189 10.6151
R1137 B.n189 B.n184 10.6151
R1138 B.n185 B.n184 10.6151
R1139 B.n185 B.n0 10.6151
R1140 B.n707 B.n1 10.6151
R1141 B.n707 B.n706 10.6151
R1142 B.n706 B.n705 10.6151
R1143 B.n705 B.n4 10.6151
R1144 B.n701 B.n4 10.6151
R1145 B.n701 B.n700 10.6151
R1146 B.n700 B.n699 10.6151
R1147 B.n699 B.n6 10.6151
R1148 B.n695 B.n6 10.6151
R1149 B.n695 B.n694 10.6151
R1150 B.n694 B.n693 10.6151
R1151 B.n693 B.n8 10.6151
R1152 B.n689 B.n8 10.6151
R1153 B.n689 B.n688 10.6151
R1154 B.n688 B.n687 10.6151
R1155 B.n687 B.n10 10.6151
R1156 B.n683 B.n10 10.6151
R1157 B.n683 B.n682 10.6151
R1158 B.n682 B.n681 10.6151
R1159 B.n681 B.n12 10.6151
R1160 B.n587 B.n586 9.36635
R1161 B.n569 B.n52 9.36635
R1162 B.n305 B.n144 9.36635
R1163 B.n323 B.n322 9.36635
R1164 B.n711 B.n0 2.81026
R1165 B.n711 B.n1 2.81026
R1166 B.n586 B.n585 1.24928
R1167 B.n572 B.n52 1.24928
R1168 B.n308 B.n144 1.24928
R1169 B.n322 B.n321 1.24928
C0 w_n1850_n4692# B 9.00586f
C1 VDD1 VDD2 0.736855f
C2 VN VTAIL 6.30745f
C3 VN VP 6.36969f
C4 VDD2 B 2.09588f
C5 VDD1 B 2.06527f
C6 w_n1850_n4692# VN 3.18059f
C7 VTAIL VP 6.322299f
C8 w_n1850_n4692# VTAIL 3.97236f
C9 VDD2 VN 6.86314f
C10 w_n1850_n4692# VP 3.41467f
C11 VDD1 VN 0.148416f
C12 VDD2 VTAIL 13.857f
C13 VN B 0.859128f
C14 VDD1 VTAIL 13.825701f
C15 VDD2 VP 0.304687f
C16 VDD1 VP 7.01276f
C17 B VTAIL 3.95081f
C18 w_n1850_n4692# VDD2 2.34065f
C19 B VP 1.24073f
C20 VDD1 w_n1850_n4692# 2.31432f
C21 VDD2 VSUBS 1.692355f
C22 VDD1 VSUBS 2.015116f
C23 VTAIL VSUBS 0.99217f
C24 VN VSUBS 5.01103f
C25 VP VSUBS 1.76959f
C26 B VSUBS 3.384403f
C27 w_n1850_n4692# VSUBS 0.106094p
C28 B.n0 VSUBS 0.005613f
C29 B.n1 VSUBS 0.005613f
C30 B.n2 VSUBS 0.008877f
C31 B.n3 VSUBS 0.008877f
C32 B.n4 VSUBS 0.008877f
C33 B.n5 VSUBS 0.008877f
C34 B.n6 VSUBS 0.008877f
C35 B.n7 VSUBS 0.008877f
C36 B.n8 VSUBS 0.008877f
C37 B.n9 VSUBS 0.008877f
C38 B.n10 VSUBS 0.008877f
C39 B.n11 VSUBS 0.008877f
C40 B.n12 VSUBS 0.019692f
C41 B.n13 VSUBS 0.008877f
C42 B.n14 VSUBS 0.008877f
C43 B.n15 VSUBS 0.008877f
C44 B.n16 VSUBS 0.008877f
C45 B.n17 VSUBS 0.008877f
C46 B.n18 VSUBS 0.008877f
C47 B.n19 VSUBS 0.008877f
C48 B.n20 VSUBS 0.008877f
C49 B.n21 VSUBS 0.008877f
C50 B.n22 VSUBS 0.008877f
C51 B.n23 VSUBS 0.008877f
C52 B.n24 VSUBS 0.008877f
C53 B.n25 VSUBS 0.008877f
C54 B.n26 VSUBS 0.008877f
C55 B.n27 VSUBS 0.008877f
C56 B.n28 VSUBS 0.008877f
C57 B.n29 VSUBS 0.008877f
C58 B.n30 VSUBS 0.008877f
C59 B.n31 VSUBS 0.008877f
C60 B.n32 VSUBS 0.008877f
C61 B.n33 VSUBS 0.008877f
C62 B.n34 VSUBS 0.008877f
C63 B.n35 VSUBS 0.008877f
C64 B.n36 VSUBS 0.008877f
C65 B.n37 VSUBS 0.008877f
C66 B.n38 VSUBS 0.008877f
C67 B.n39 VSUBS 0.008877f
C68 B.n40 VSUBS 0.008877f
C69 B.n41 VSUBS 0.008877f
C70 B.n42 VSUBS 0.008877f
C71 B.n43 VSUBS 0.008877f
C72 B.t5 VSUBS 0.799018f
C73 B.t4 VSUBS 0.810156f
C74 B.t3 VSUBS 0.735695f
C75 B.n44 VSUBS 0.253812f
C76 B.n45 VSUBS 0.081836f
C77 B.n46 VSUBS 0.008877f
C78 B.n47 VSUBS 0.008877f
C79 B.n48 VSUBS 0.008877f
C80 B.n49 VSUBS 0.008877f
C81 B.t11 VSUBS 0.798988f
C82 B.t10 VSUBS 0.810128f
C83 B.t9 VSUBS 0.735695f
C84 B.n50 VSUBS 0.253839f
C85 B.n51 VSUBS 0.081866f
C86 B.n52 VSUBS 0.020566f
C87 B.n53 VSUBS 0.008877f
C88 B.n54 VSUBS 0.008877f
C89 B.n55 VSUBS 0.008877f
C90 B.n56 VSUBS 0.008877f
C91 B.n57 VSUBS 0.008877f
C92 B.n58 VSUBS 0.008877f
C93 B.n59 VSUBS 0.008877f
C94 B.n60 VSUBS 0.008877f
C95 B.n61 VSUBS 0.008877f
C96 B.n62 VSUBS 0.008877f
C97 B.n63 VSUBS 0.008877f
C98 B.n64 VSUBS 0.008877f
C99 B.n65 VSUBS 0.008877f
C100 B.n66 VSUBS 0.008877f
C101 B.n67 VSUBS 0.008877f
C102 B.n68 VSUBS 0.008877f
C103 B.n69 VSUBS 0.008877f
C104 B.n70 VSUBS 0.008877f
C105 B.n71 VSUBS 0.008877f
C106 B.n72 VSUBS 0.008877f
C107 B.n73 VSUBS 0.008877f
C108 B.n74 VSUBS 0.008877f
C109 B.n75 VSUBS 0.008877f
C110 B.n76 VSUBS 0.008877f
C111 B.n77 VSUBS 0.008877f
C112 B.n78 VSUBS 0.008877f
C113 B.n79 VSUBS 0.008877f
C114 B.n80 VSUBS 0.008877f
C115 B.n81 VSUBS 0.008877f
C116 B.n82 VSUBS 0.008877f
C117 B.n83 VSUBS 0.019692f
C118 B.n84 VSUBS 0.008877f
C119 B.n85 VSUBS 0.008877f
C120 B.n86 VSUBS 0.008877f
C121 B.n87 VSUBS 0.008877f
C122 B.n88 VSUBS 0.008877f
C123 B.n89 VSUBS 0.008877f
C124 B.n90 VSUBS 0.008877f
C125 B.n91 VSUBS 0.008877f
C126 B.n92 VSUBS 0.008877f
C127 B.n93 VSUBS 0.008877f
C128 B.n94 VSUBS 0.008877f
C129 B.n95 VSUBS 0.008877f
C130 B.n96 VSUBS 0.008877f
C131 B.n97 VSUBS 0.008877f
C132 B.n98 VSUBS 0.008877f
C133 B.n99 VSUBS 0.008877f
C134 B.n100 VSUBS 0.008877f
C135 B.n101 VSUBS 0.008877f
C136 B.n102 VSUBS 0.008877f
C137 B.n103 VSUBS 0.008877f
C138 B.n104 VSUBS 0.019692f
C139 B.n105 VSUBS 0.008877f
C140 B.n106 VSUBS 0.008877f
C141 B.n107 VSUBS 0.008877f
C142 B.n108 VSUBS 0.008877f
C143 B.n109 VSUBS 0.008877f
C144 B.n110 VSUBS 0.008877f
C145 B.n111 VSUBS 0.008877f
C146 B.n112 VSUBS 0.008877f
C147 B.n113 VSUBS 0.008877f
C148 B.n114 VSUBS 0.008877f
C149 B.n115 VSUBS 0.008877f
C150 B.n116 VSUBS 0.008877f
C151 B.n117 VSUBS 0.008877f
C152 B.n118 VSUBS 0.008877f
C153 B.n119 VSUBS 0.008877f
C154 B.n120 VSUBS 0.008877f
C155 B.n121 VSUBS 0.008877f
C156 B.n122 VSUBS 0.008877f
C157 B.n123 VSUBS 0.008877f
C158 B.n124 VSUBS 0.008877f
C159 B.n125 VSUBS 0.008877f
C160 B.n126 VSUBS 0.008877f
C161 B.n127 VSUBS 0.008877f
C162 B.n128 VSUBS 0.008877f
C163 B.n129 VSUBS 0.008877f
C164 B.n130 VSUBS 0.008877f
C165 B.n131 VSUBS 0.008877f
C166 B.n132 VSUBS 0.008877f
C167 B.n133 VSUBS 0.008877f
C168 B.n134 VSUBS 0.008877f
C169 B.n135 VSUBS 0.008877f
C170 B.t7 VSUBS 0.798988f
C171 B.t8 VSUBS 0.810128f
C172 B.t6 VSUBS 0.735695f
C173 B.n136 VSUBS 0.253839f
C174 B.n137 VSUBS 0.081866f
C175 B.n138 VSUBS 0.008877f
C176 B.n139 VSUBS 0.008877f
C177 B.n140 VSUBS 0.008877f
C178 B.n141 VSUBS 0.008877f
C179 B.t1 VSUBS 0.799018f
C180 B.t2 VSUBS 0.810156f
C181 B.t0 VSUBS 0.735695f
C182 B.n142 VSUBS 0.253812f
C183 B.n143 VSUBS 0.081836f
C184 B.n144 VSUBS 0.020566f
C185 B.n145 VSUBS 0.008877f
C186 B.n146 VSUBS 0.008877f
C187 B.n147 VSUBS 0.008877f
C188 B.n148 VSUBS 0.008877f
C189 B.n149 VSUBS 0.008877f
C190 B.n150 VSUBS 0.008877f
C191 B.n151 VSUBS 0.008877f
C192 B.n152 VSUBS 0.008877f
C193 B.n153 VSUBS 0.008877f
C194 B.n154 VSUBS 0.008877f
C195 B.n155 VSUBS 0.008877f
C196 B.n156 VSUBS 0.008877f
C197 B.n157 VSUBS 0.008877f
C198 B.n158 VSUBS 0.008877f
C199 B.n159 VSUBS 0.008877f
C200 B.n160 VSUBS 0.008877f
C201 B.n161 VSUBS 0.008877f
C202 B.n162 VSUBS 0.008877f
C203 B.n163 VSUBS 0.008877f
C204 B.n164 VSUBS 0.008877f
C205 B.n165 VSUBS 0.008877f
C206 B.n166 VSUBS 0.008877f
C207 B.n167 VSUBS 0.008877f
C208 B.n168 VSUBS 0.008877f
C209 B.n169 VSUBS 0.008877f
C210 B.n170 VSUBS 0.008877f
C211 B.n171 VSUBS 0.008877f
C212 B.n172 VSUBS 0.008877f
C213 B.n173 VSUBS 0.008877f
C214 B.n174 VSUBS 0.008877f
C215 B.n175 VSUBS 0.019692f
C216 B.n176 VSUBS 0.008877f
C217 B.n177 VSUBS 0.008877f
C218 B.n178 VSUBS 0.008877f
C219 B.n179 VSUBS 0.008877f
C220 B.n180 VSUBS 0.008877f
C221 B.n181 VSUBS 0.008877f
C222 B.n182 VSUBS 0.008877f
C223 B.n183 VSUBS 0.008877f
C224 B.n184 VSUBS 0.008877f
C225 B.n185 VSUBS 0.008877f
C226 B.n186 VSUBS 0.008877f
C227 B.n187 VSUBS 0.008877f
C228 B.n188 VSUBS 0.008877f
C229 B.n189 VSUBS 0.008877f
C230 B.n190 VSUBS 0.008877f
C231 B.n191 VSUBS 0.008877f
C232 B.n192 VSUBS 0.008877f
C233 B.n193 VSUBS 0.008877f
C234 B.n194 VSUBS 0.008877f
C235 B.n195 VSUBS 0.008877f
C236 B.n196 VSUBS 0.008877f
C237 B.n197 VSUBS 0.008877f
C238 B.n198 VSUBS 0.008877f
C239 B.n199 VSUBS 0.008877f
C240 B.n200 VSUBS 0.008877f
C241 B.n201 VSUBS 0.008877f
C242 B.n202 VSUBS 0.008877f
C243 B.n203 VSUBS 0.008877f
C244 B.n204 VSUBS 0.008877f
C245 B.n205 VSUBS 0.008877f
C246 B.n206 VSUBS 0.008877f
C247 B.n207 VSUBS 0.008877f
C248 B.n208 VSUBS 0.008877f
C249 B.n209 VSUBS 0.008877f
C250 B.n210 VSUBS 0.008877f
C251 B.n211 VSUBS 0.008877f
C252 B.n212 VSUBS 0.008877f
C253 B.n213 VSUBS 0.008877f
C254 B.n214 VSUBS 0.019692f
C255 B.n215 VSUBS 0.021037f
C256 B.n216 VSUBS 0.021037f
C257 B.n217 VSUBS 0.008877f
C258 B.n218 VSUBS 0.008877f
C259 B.n219 VSUBS 0.008877f
C260 B.n220 VSUBS 0.008877f
C261 B.n221 VSUBS 0.008877f
C262 B.n222 VSUBS 0.008877f
C263 B.n223 VSUBS 0.008877f
C264 B.n224 VSUBS 0.008877f
C265 B.n225 VSUBS 0.008877f
C266 B.n226 VSUBS 0.008877f
C267 B.n227 VSUBS 0.008877f
C268 B.n228 VSUBS 0.008877f
C269 B.n229 VSUBS 0.008877f
C270 B.n230 VSUBS 0.008877f
C271 B.n231 VSUBS 0.008877f
C272 B.n232 VSUBS 0.008877f
C273 B.n233 VSUBS 0.008877f
C274 B.n234 VSUBS 0.008877f
C275 B.n235 VSUBS 0.008877f
C276 B.n236 VSUBS 0.008877f
C277 B.n237 VSUBS 0.008877f
C278 B.n238 VSUBS 0.008877f
C279 B.n239 VSUBS 0.008877f
C280 B.n240 VSUBS 0.008877f
C281 B.n241 VSUBS 0.008877f
C282 B.n242 VSUBS 0.008877f
C283 B.n243 VSUBS 0.008877f
C284 B.n244 VSUBS 0.008877f
C285 B.n245 VSUBS 0.008877f
C286 B.n246 VSUBS 0.008877f
C287 B.n247 VSUBS 0.008877f
C288 B.n248 VSUBS 0.008877f
C289 B.n249 VSUBS 0.008877f
C290 B.n250 VSUBS 0.008877f
C291 B.n251 VSUBS 0.008877f
C292 B.n252 VSUBS 0.008877f
C293 B.n253 VSUBS 0.008877f
C294 B.n254 VSUBS 0.008877f
C295 B.n255 VSUBS 0.008877f
C296 B.n256 VSUBS 0.008877f
C297 B.n257 VSUBS 0.008877f
C298 B.n258 VSUBS 0.008877f
C299 B.n259 VSUBS 0.008877f
C300 B.n260 VSUBS 0.008877f
C301 B.n261 VSUBS 0.008877f
C302 B.n262 VSUBS 0.008877f
C303 B.n263 VSUBS 0.008877f
C304 B.n264 VSUBS 0.008877f
C305 B.n265 VSUBS 0.008877f
C306 B.n266 VSUBS 0.008877f
C307 B.n267 VSUBS 0.008877f
C308 B.n268 VSUBS 0.008877f
C309 B.n269 VSUBS 0.008877f
C310 B.n270 VSUBS 0.008877f
C311 B.n271 VSUBS 0.008877f
C312 B.n272 VSUBS 0.008877f
C313 B.n273 VSUBS 0.008877f
C314 B.n274 VSUBS 0.008877f
C315 B.n275 VSUBS 0.008877f
C316 B.n276 VSUBS 0.008877f
C317 B.n277 VSUBS 0.008877f
C318 B.n278 VSUBS 0.008877f
C319 B.n279 VSUBS 0.008877f
C320 B.n280 VSUBS 0.008877f
C321 B.n281 VSUBS 0.008877f
C322 B.n282 VSUBS 0.008877f
C323 B.n283 VSUBS 0.008877f
C324 B.n284 VSUBS 0.008877f
C325 B.n285 VSUBS 0.008877f
C326 B.n286 VSUBS 0.008877f
C327 B.n287 VSUBS 0.008877f
C328 B.n288 VSUBS 0.008877f
C329 B.n289 VSUBS 0.008877f
C330 B.n290 VSUBS 0.008877f
C331 B.n291 VSUBS 0.008877f
C332 B.n292 VSUBS 0.008877f
C333 B.n293 VSUBS 0.008877f
C334 B.n294 VSUBS 0.008877f
C335 B.n295 VSUBS 0.008877f
C336 B.n296 VSUBS 0.008877f
C337 B.n297 VSUBS 0.008877f
C338 B.n298 VSUBS 0.008877f
C339 B.n299 VSUBS 0.008877f
C340 B.n300 VSUBS 0.008877f
C341 B.n301 VSUBS 0.008877f
C342 B.n302 VSUBS 0.008877f
C343 B.n303 VSUBS 0.008877f
C344 B.n304 VSUBS 0.008877f
C345 B.n305 VSUBS 0.008355f
C346 B.n306 VSUBS 0.008877f
C347 B.n307 VSUBS 0.008877f
C348 B.n308 VSUBS 0.004961f
C349 B.n309 VSUBS 0.008877f
C350 B.n310 VSUBS 0.008877f
C351 B.n311 VSUBS 0.008877f
C352 B.n312 VSUBS 0.008877f
C353 B.n313 VSUBS 0.008877f
C354 B.n314 VSUBS 0.008877f
C355 B.n315 VSUBS 0.008877f
C356 B.n316 VSUBS 0.008877f
C357 B.n317 VSUBS 0.008877f
C358 B.n318 VSUBS 0.008877f
C359 B.n319 VSUBS 0.008877f
C360 B.n320 VSUBS 0.008877f
C361 B.n321 VSUBS 0.004961f
C362 B.n322 VSUBS 0.020566f
C363 B.n323 VSUBS 0.008355f
C364 B.n324 VSUBS 0.008877f
C365 B.n325 VSUBS 0.008877f
C366 B.n326 VSUBS 0.008877f
C367 B.n327 VSUBS 0.008877f
C368 B.n328 VSUBS 0.008877f
C369 B.n329 VSUBS 0.008877f
C370 B.n330 VSUBS 0.008877f
C371 B.n331 VSUBS 0.008877f
C372 B.n332 VSUBS 0.008877f
C373 B.n333 VSUBS 0.008877f
C374 B.n334 VSUBS 0.008877f
C375 B.n335 VSUBS 0.008877f
C376 B.n336 VSUBS 0.008877f
C377 B.n337 VSUBS 0.008877f
C378 B.n338 VSUBS 0.008877f
C379 B.n339 VSUBS 0.008877f
C380 B.n340 VSUBS 0.008877f
C381 B.n341 VSUBS 0.008877f
C382 B.n342 VSUBS 0.008877f
C383 B.n343 VSUBS 0.008877f
C384 B.n344 VSUBS 0.008877f
C385 B.n345 VSUBS 0.008877f
C386 B.n346 VSUBS 0.008877f
C387 B.n347 VSUBS 0.008877f
C388 B.n348 VSUBS 0.008877f
C389 B.n349 VSUBS 0.008877f
C390 B.n350 VSUBS 0.008877f
C391 B.n351 VSUBS 0.008877f
C392 B.n352 VSUBS 0.008877f
C393 B.n353 VSUBS 0.008877f
C394 B.n354 VSUBS 0.008877f
C395 B.n355 VSUBS 0.008877f
C396 B.n356 VSUBS 0.008877f
C397 B.n357 VSUBS 0.008877f
C398 B.n358 VSUBS 0.008877f
C399 B.n359 VSUBS 0.008877f
C400 B.n360 VSUBS 0.008877f
C401 B.n361 VSUBS 0.008877f
C402 B.n362 VSUBS 0.008877f
C403 B.n363 VSUBS 0.008877f
C404 B.n364 VSUBS 0.008877f
C405 B.n365 VSUBS 0.008877f
C406 B.n366 VSUBS 0.008877f
C407 B.n367 VSUBS 0.008877f
C408 B.n368 VSUBS 0.008877f
C409 B.n369 VSUBS 0.008877f
C410 B.n370 VSUBS 0.008877f
C411 B.n371 VSUBS 0.008877f
C412 B.n372 VSUBS 0.008877f
C413 B.n373 VSUBS 0.008877f
C414 B.n374 VSUBS 0.008877f
C415 B.n375 VSUBS 0.008877f
C416 B.n376 VSUBS 0.008877f
C417 B.n377 VSUBS 0.008877f
C418 B.n378 VSUBS 0.008877f
C419 B.n379 VSUBS 0.008877f
C420 B.n380 VSUBS 0.008877f
C421 B.n381 VSUBS 0.008877f
C422 B.n382 VSUBS 0.008877f
C423 B.n383 VSUBS 0.008877f
C424 B.n384 VSUBS 0.008877f
C425 B.n385 VSUBS 0.008877f
C426 B.n386 VSUBS 0.008877f
C427 B.n387 VSUBS 0.008877f
C428 B.n388 VSUBS 0.008877f
C429 B.n389 VSUBS 0.008877f
C430 B.n390 VSUBS 0.008877f
C431 B.n391 VSUBS 0.008877f
C432 B.n392 VSUBS 0.008877f
C433 B.n393 VSUBS 0.008877f
C434 B.n394 VSUBS 0.008877f
C435 B.n395 VSUBS 0.008877f
C436 B.n396 VSUBS 0.008877f
C437 B.n397 VSUBS 0.008877f
C438 B.n398 VSUBS 0.008877f
C439 B.n399 VSUBS 0.008877f
C440 B.n400 VSUBS 0.008877f
C441 B.n401 VSUBS 0.008877f
C442 B.n402 VSUBS 0.008877f
C443 B.n403 VSUBS 0.008877f
C444 B.n404 VSUBS 0.008877f
C445 B.n405 VSUBS 0.008877f
C446 B.n406 VSUBS 0.008877f
C447 B.n407 VSUBS 0.008877f
C448 B.n408 VSUBS 0.008877f
C449 B.n409 VSUBS 0.008877f
C450 B.n410 VSUBS 0.008877f
C451 B.n411 VSUBS 0.008877f
C452 B.n412 VSUBS 0.008877f
C453 B.n413 VSUBS 0.021037f
C454 B.n414 VSUBS 0.021037f
C455 B.n415 VSUBS 0.019692f
C456 B.n416 VSUBS 0.008877f
C457 B.n417 VSUBS 0.008877f
C458 B.n418 VSUBS 0.008877f
C459 B.n419 VSUBS 0.008877f
C460 B.n420 VSUBS 0.008877f
C461 B.n421 VSUBS 0.008877f
C462 B.n422 VSUBS 0.008877f
C463 B.n423 VSUBS 0.008877f
C464 B.n424 VSUBS 0.008877f
C465 B.n425 VSUBS 0.008877f
C466 B.n426 VSUBS 0.008877f
C467 B.n427 VSUBS 0.008877f
C468 B.n428 VSUBS 0.008877f
C469 B.n429 VSUBS 0.008877f
C470 B.n430 VSUBS 0.008877f
C471 B.n431 VSUBS 0.008877f
C472 B.n432 VSUBS 0.008877f
C473 B.n433 VSUBS 0.008877f
C474 B.n434 VSUBS 0.008877f
C475 B.n435 VSUBS 0.008877f
C476 B.n436 VSUBS 0.008877f
C477 B.n437 VSUBS 0.008877f
C478 B.n438 VSUBS 0.008877f
C479 B.n439 VSUBS 0.008877f
C480 B.n440 VSUBS 0.008877f
C481 B.n441 VSUBS 0.008877f
C482 B.n442 VSUBS 0.008877f
C483 B.n443 VSUBS 0.008877f
C484 B.n444 VSUBS 0.008877f
C485 B.n445 VSUBS 0.008877f
C486 B.n446 VSUBS 0.008877f
C487 B.n447 VSUBS 0.008877f
C488 B.n448 VSUBS 0.008877f
C489 B.n449 VSUBS 0.008877f
C490 B.n450 VSUBS 0.008877f
C491 B.n451 VSUBS 0.008877f
C492 B.n452 VSUBS 0.008877f
C493 B.n453 VSUBS 0.008877f
C494 B.n454 VSUBS 0.008877f
C495 B.n455 VSUBS 0.008877f
C496 B.n456 VSUBS 0.008877f
C497 B.n457 VSUBS 0.008877f
C498 B.n458 VSUBS 0.008877f
C499 B.n459 VSUBS 0.008877f
C500 B.n460 VSUBS 0.008877f
C501 B.n461 VSUBS 0.008877f
C502 B.n462 VSUBS 0.008877f
C503 B.n463 VSUBS 0.008877f
C504 B.n464 VSUBS 0.008877f
C505 B.n465 VSUBS 0.008877f
C506 B.n466 VSUBS 0.008877f
C507 B.n467 VSUBS 0.008877f
C508 B.n468 VSUBS 0.008877f
C509 B.n469 VSUBS 0.008877f
C510 B.n470 VSUBS 0.008877f
C511 B.n471 VSUBS 0.008877f
C512 B.n472 VSUBS 0.008877f
C513 B.n473 VSUBS 0.008877f
C514 B.n474 VSUBS 0.008877f
C515 B.n475 VSUBS 0.008877f
C516 B.n476 VSUBS 0.008877f
C517 B.n477 VSUBS 0.008877f
C518 B.n478 VSUBS 0.020773f
C519 B.n479 VSUBS 0.019956f
C520 B.n480 VSUBS 0.021037f
C521 B.n481 VSUBS 0.008877f
C522 B.n482 VSUBS 0.008877f
C523 B.n483 VSUBS 0.008877f
C524 B.n484 VSUBS 0.008877f
C525 B.n485 VSUBS 0.008877f
C526 B.n486 VSUBS 0.008877f
C527 B.n487 VSUBS 0.008877f
C528 B.n488 VSUBS 0.008877f
C529 B.n489 VSUBS 0.008877f
C530 B.n490 VSUBS 0.008877f
C531 B.n491 VSUBS 0.008877f
C532 B.n492 VSUBS 0.008877f
C533 B.n493 VSUBS 0.008877f
C534 B.n494 VSUBS 0.008877f
C535 B.n495 VSUBS 0.008877f
C536 B.n496 VSUBS 0.008877f
C537 B.n497 VSUBS 0.008877f
C538 B.n498 VSUBS 0.008877f
C539 B.n499 VSUBS 0.008877f
C540 B.n500 VSUBS 0.008877f
C541 B.n501 VSUBS 0.008877f
C542 B.n502 VSUBS 0.008877f
C543 B.n503 VSUBS 0.008877f
C544 B.n504 VSUBS 0.008877f
C545 B.n505 VSUBS 0.008877f
C546 B.n506 VSUBS 0.008877f
C547 B.n507 VSUBS 0.008877f
C548 B.n508 VSUBS 0.008877f
C549 B.n509 VSUBS 0.008877f
C550 B.n510 VSUBS 0.008877f
C551 B.n511 VSUBS 0.008877f
C552 B.n512 VSUBS 0.008877f
C553 B.n513 VSUBS 0.008877f
C554 B.n514 VSUBS 0.008877f
C555 B.n515 VSUBS 0.008877f
C556 B.n516 VSUBS 0.008877f
C557 B.n517 VSUBS 0.008877f
C558 B.n518 VSUBS 0.008877f
C559 B.n519 VSUBS 0.008877f
C560 B.n520 VSUBS 0.008877f
C561 B.n521 VSUBS 0.008877f
C562 B.n522 VSUBS 0.008877f
C563 B.n523 VSUBS 0.008877f
C564 B.n524 VSUBS 0.008877f
C565 B.n525 VSUBS 0.008877f
C566 B.n526 VSUBS 0.008877f
C567 B.n527 VSUBS 0.008877f
C568 B.n528 VSUBS 0.008877f
C569 B.n529 VSUBS 0.008877f
C570 B.n530 VSUBS 0.008877f
C571 B.n531 VSUBS 0.008877f
C572 B.n532 VSUBS 0.008877f
C573 B.n533 VSUBS 0.008877f
C574 B.n534 VSUBS 0.008877f
C575 B.n535 VSUBS 0.008877f
C576 B.n536 VSUBS 0.008877f
C577 B.n537 VSUBS 0.008877f
C578 B.n538 VSUBS 0.008877f
C579 B.n539 VSUBS 0.008877f
C580 B.n540 VSUBS 0.008877f
C581 B.n541 VSUBS 0.008877f
C582 B.n542 VSUBS 0.008877f
C583 B.n543 VSUBS 0.008877f
C584 B.n544 VSUBS 0.008877f
C585 B.n545 VSUBS 0.008877f
C586 B.n546 VSUBS 0.008877f
C587 B.n547 VSUBS 0.008877f
C588 B.n548 VSUBS 0.008877f
C589 B.n549 VSUBS 0.008877f
C590 B.n550 VSUBS 0.008877f
C591 B.n551 VSUBS 0.008877f
C592 B.n552 VSUBS 0.008877f
C593 B.n553 VSUBS 0.008877f
C594 B.n554 VSUBS 0.008877f
C595 B.n555 VSUBS 0.008877f
C596 B.n556 VSUBS 0.008877f
C597 B.n557 VSUBS 0.008877f
C598 B.n558 VSUBS 0.008877f
C599 B.n559 VSUBS 0.008877f
C600 B.n560 VSUBS 0.008877f
C601 B.n561 VSUBS 0.008877f
C602 B.n562 VSUBS 0.008877f
C603 B.n563 VSUBS 0.008877f
C604 B.n564 VSUBS 0.008877f
C605 B.n565 VSUBS 0.008877f
C606 B.n566 VSUBS 0.008877f
C607 B.n567 VSUBS 0.008877f
C608 B.n568 VSUBS 0.008877f
C609 B.n569 VSUBS 0.008355f
C610 B.n570 VSUBS 0.008877f
C611 B.n571 VSUBS 0.008877f
C612 B.n572 VSUBS 0.004961f
C613 B.n573 VSUBS 0.008877f
C614 B.n574 VSUBS 0.008877f
C615 B.n575 VSUBS 0.008877f
C616 B.n576 VSUBS 0.008877f
C617 B.n577 VSUBS 0.008877f
C618 B.n578 VSUBS 0.008877f
C619 B.n579 VSUBS 0.008877f
C620 B.n580 VSUBS 0.008877f
C621 B.n581 VSUBS 0.008877f
C622 B.n582 VSUBS 0.008877f
C623 B.n583 VSUBS 0.008877f
C624 B.n584 VSUBS 0.008877f
C625 B.n585 VSUBS 0.004961f
C626 B.n586 VSUBS 0.020566f
C627 B.n587 VSUBS 0.008355f
C628 B.n588 VSUBS 0.008877f
C629 B.n589 VSUBS 0.008877f
C630 B.n590 VSUBS 0.008877f
C631 B.n591 VSUBS 0.008877f
C632 B.n592 VSUBS 0.008877f
C633 B.n593 VSUBS 0.008877f
C634 B.n594 VSUBS 0.008877f
C635 B.n595 VSUBS 0.008877f
C636 B.n596 VSUBS 0.008877f
C637 B.n597 VSUBS 0.008877f
C638 B.n598 VSUBS 0.008877f
C639 B.n599 VSUBS 0.008877f
C640 B.n600 VSUBS 0.008877f
C641 B.n601 VSUBS 0.008877f
C642 B.n602 VSUBS 0.008877f
C643 B.n603 VSUBS 0.008877f
C644 B.n604 VSUBS 0.008877f
C645 B.n605 VSUBS 0.008877f
C646 B.n606 VSUBS 0.008877f
C647 B.n607 VSUBS 0.008877f
C648 B.n608 VSUBS 0.008877f
C649 B.n609 VSUBS 0.008877f
C650 B.n610 VSUBS 0.008877f
C651 B.n611 VSUBS 0.008877f
C652 B.n612 VSUBS 0.008877f
C653 B.n613 VSUBS 0.008877f
C654 B.n614 VSUBS 0.008877f
C655 B.n615 VSUBS 0.008877f
C656 B.n616 VSUBS 0.008877f
C657 B.n617 VSUBS 0.008877f
C658 B.n618 VSUBS 0.008877f
C659 B.n619 VSUBS 0.008877f
C660 B.n620 VSUBS 0.008877f
C661 B.n621 VSUBS 0.008877f
C662 B.n622 VSUBS 0.008877f
C663 B.n623 VSUBS 0.008877f
C664 B.n624 VSUBS 0.008877f
C665 B.n625 VSUBS 0.008877f
C666 B.n626 VSUBS 0.008877f
C667 B.n627 VSUBS 0.008877f
C668 B.n628 VSUBS 0.008877f
C669 B.n629 VSUBS 0.008877f
C670 B.n630 VSUBS 0.008877f
C671 B.n631 VSUBS 0.008877f
C672 B.n632 VSUBS 0.008877f
C673 B.n633 VSUBS 0.008877f
C674 B.n634 VSUBS 0.008877f
C675 B.n635 VSUBS 0.008877f
C676 B.n636 VSUBS 0.008877f
C677 B.n637 VSUBS 0.008877f
C678 B.n638 VSUBS 0.008877f
C679 B.n639 VSUBS 0.008877f
C680 B.n640 VSUBS 0.008877f
C681 B.n641 VSUBS 0.008877f
C682 B.n642 VSUBS 0.008877f
C683 B.n643 VSUBS 0.008877f
C684 B.n644 VSUBS 0.008877f
C685 B.n645 VSUBS 0.008877f
C686 B.n646 VSUBS 0.008877f
C687 B.n647 VSUBS 0.008877f
C688 B.n648 VSUBS 0.008877f
C689 B.n649 VSUBS 0.008877f
C690 B.n650 VSUBS 0.008877f
C691 B.n651 VSUBS 0.008877f
C692 B.n652 VSUBS 0.008877f
C693 B.n653 VSUBS 0.008877f
C694 B.n654 VSUBS 0.008877f
C695 B.n655 VSUBS 0.008877f
C696 B.n656 VSUBS 0.008877f
C697 B.n657 VSUBS 0.008877f
C698 B.n658 VSUBS 0.008877f
C699 B.n659 VSUBS 0.008877f
C700 B.n660 VSUBS 0.008877f
C701 B.n661 VSUBS 0.008877f
C702 B.n662 VSUBS 0.008877f
C703 B.n663 VSUBS 0.008877f
C704 B.n664 VSUBS 0.008877f
C705 B.n665 VSUBS 0.008877f
C706 B.n666 VSUBS 0.008877f
C707 B.n667 VSUBS 0.008877f
C708 B.n668 VSUBS 0.008877f
C709 B.n669 VSUBS 0.008877f
C710 B.n670 VSUBS 0.008877f
C711 B.n671 VSUBS 0.008877f
C712 B.n672 VSUBS 0.008877f
C713 B.n673 VSUBS 0.008877f
C714 B.n674 VSUBS 0.008877f
C715 B.n675 VSUBS 0.008877f
C716 B.n676 VSUBS 0.008877f
C717 B.n677 VSUBS 0.021037f
C718 B.n678 VSUBS 0.021037f
C719 B.n679 VSUBS 0.019692f
C720 B.n680 VSUBS 0.008877f
C721 B.n681 VSUBS 0.008877f
C722 B.n682 VSUBS 0.008877f
C723 B.n683 VSUBS 0.008877f
C724 B.n684 VSUBS 0.008877f
C725 B.n685 VSUBS 0.008877f
C726 B.n686 VSUBS 0.008877f
C727 B.n687 VSUBS 0.008877f
C728 B.n688 VSUBS 0.008877f
C729 B.n689 VSUBS 0.008877f
C730 B.n690 VSUBS 0.008877f
C731 B.n691 VSUBS 0.008877f
C732 B.n692 VSUBS 0.008877f
C733 B.n693 VSUBS 0.008877f
C734 B.n694 VSUBS 0.008877f
C735 B.n695 VSUBS 0.008877f
C736 B.n696 VSUBS 0.008877f
C737 B.n697 VSUBS 0.008877f
C738 B.n698 VSUBS 0.008877f
C739 B.n699 VSUBS 0.008877f
C740 B.n700 VSUBS 0.008877f
C741 B.n701 VSUBS 0.008877f
C742 B.n702 VSUBS 0.008877f
C743 B.n703 VSUBS 0.008877f
C744 B.n704 VSUBS 0.008877f
C745 B.n705 VSUBS 0.008877f
C746 B.n706 VSUBS 0.008877f
C747 B.n707 VSUBS 0.008877f
C748 B.n708 VSUBS 0.008877f
C749 B.n709 VSUBS 0.008877f
C750 B.n710 VSUBS 0.008877f
C751 B.n711 VSUBS 0.0201f
C752 VDD1.t4 VSUBS 4.44914f
C753 VDD1.t5 VSUBS 4.44787f
C754 VDD1.t0 VSUBS 0.410384f
C755 VDD1.t2 VSUBS 0.410384f
C756 VDD1.n0 VSUBS 3.42584f
C757 VDD1.n1 VSUBS 3.57568f
C758 VDD1.t1 VSUBS 0.410384f
C759 VDD1.t3 VSUBS 0.410384f
C760 VDD1.n2 VSUBS 3.42408f
C761 VDD1.n3 VSUBS 3.42434f
C762 VP.n0 VSUBS 0.052175f
C763 VP.n1 VSUBS 0.01184f
C764 VP.n2 VSUBS 0.22271f
C765 VP.t2 VSUBS 2.12003f
C766 VP.t4 VSUBS 2.12003f
C767 VP.t1 VSUBS 2.14781f
C768 VP.n3 VSUBS 0.772602f
C769 VP.n4 VSUBS 0.798806f
C770 VP.n5 VSUBS 0.01184f
C771 VP.n6 VSUBS 0.792879f
C772 VP.n7 VSUBS 2.54309f
C773 VP.t0 VSUBS 2.12003f
C774 VP.n8 VSUBS 0.792879f
C775 VP.n9 VSUBS 2.58349f
C776 VP.n10 VSUBS 0.052175f
C777 VP.n11 VSUBS 0.052175f
C778 VP.t5 VSUBS 2.12003f
C779 VP.n12 VSUBS 0.793361f
C780 VP.n13 VSUBS 0.01184f
C781 VP.t3 VSUBS 2.12003f
C782 VP.n14 VSUBS 0.792879f
C783 VP.n15 VSUBS 0.040433f
C784 VTAIL.t6 VSUBS 0.412249f
C785 VTAIL.t10 VSUBS 0.412249f
C786 VTAIL.n0 VSUBS 3.26439f
C787 VTAIL.n1 VSUBS 0.803303f
C788 VTAIL.t2 VSUBS 4.26011f
C789 VTAIL.n2 VSUBS 0.99085f
C790 VTAIL.t3 VSUBS 0.412249f
C791 VTAIL.t4 VSUBS 0.412249f
C792 VTAIL.n3 VSUBS 3.26439f
C793 VTAIL.n4 VSUBS 2.77795f
C794 VTAIL.t9 VSUBS 0.412249f
C795 VTAIL.t8 VSUBS 0.412249f
C796 VTAIL.n5 VSUBS 3.2644f
C797 VTAIL.n6 VSUBS 2.77795f
C798 VTAIL.t5 VSUBS 4.26014f
C799 VTAIL.n7 VSUBS 0.990818f
C800 VTAIL.t0 VSUBS 0.412249f
C801 VTAIL.t1 VSUBS 0.412249f
C802 VTAIL.n8 VSUBS 3.2644f
C803 VTAIL.n9 VSUBS 0.862249f
C804 VTAIL.t11 VSUBS 4.26011f
C805 VTAIL.n10 VSUBS 2.82094f
C806 VTAIL.t7 VSUBS 4.26011f
C807 VTAIL.n11 VSUBS 2.79428f
C808 VDD2.t5 VSUBS 4.46613f
C809 VDD2.t2 VSUBS 0.412068f
C810 VDD2.t3 VSUBS 0.412068f
C811 VDD2.n0 VSUBS 3.4399f
C812 VDD2.n1 VSUBS 3.5001f
C813 VDD2.t4 VSUBS 4.45946f
C814 VDD2.n2 VSUBS 3.49542f
C815 VDD2.t1 VSUBS 0.412068f
C816 VDD2.t0 VSUBS 0.412068f
C817 VDD2.n3 VSUBS 3.43986f
C818 VN.n0 VSUBS 0.219122f
C819 VN.t4 VSUBS 2.11321f
C820 VN.n1 VSUBS 0.760155f
C821 VN.t0 VSUBS 2.08588f
C822 VN.n2 VSUBS 0.785937f
C823 VN.n3 VSUBS 0.011649f
C824 VN.t3 VSUBS 2.08588f
C825 VN.n4 VSUBS 0.780105f
C826 VN.n5 VSUBS 0.039782f
C827 VN.n6 VSUBS 0.219122f
C828 VN.t5 VSUBS 2.11321f
C829 VN.n7 VSUBS 0.760155f
C830 VN.t2 VSUBS 2.08588f
C831 VN.n8 VSUBS 0.785937f
C832 VN.n9 VSUBS 0.011649f
C833 VN.t1 VSUBS 2.08588f
C834 VN.n10 VSUBS 0.780105f
C835 VN.n11 VSUBS 2.53562f
.ends

