* NGSPICE file created from diff_pair_sample_0111.ext - technology: sky130A

.subckt diff_pair_sample_0111 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n2154_n4078# sky130_fd_pr__pfet_01v8 ad=6.0645 pd=31.88 as=6.0645 ps=31.88 w=15.55 l=2.63
X1 B.t11 B.t9 B.t10 w_n2154_n4078# sky130_fd_pr__pfet_01v8 ad=6.0645 pd=31.88 as=0 ps=0 w=15.55 l=2.63
X2 VDD1.t0 VP.t1 VTAIL.t3 w_n2154_n4078# sky130_fd_pr__pfet_01v8 ad=6.0645 pd=31.88 as=6.0645 ps=31.88 w=15.55 l=2.63
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n2154_n4078# sky130_fd_pr__pfet_01v8 ad=6.0645 pd=31.88 as=6.0645 ps=31.88 w=15.55 l=2.63
X4 B.t8 B.t6 B.t7 w_n2154_n4078# sky130_fd_pr__pfet_01v8 ad=6.0645 pd=31.88 as=0 ps=0 w=15.55 l=2.63
X5 VDD2.t0 VN.t1 VTAIL.t0 w_n2154_n4078# sky130_fd_pr__pfet_01v8 ad=6.0645 pd=31.88 as=6.0645 ps=31.88 w=15.55 l=2.63
X6 B.t5 B.t3 B.t4 w_n2154_n4078# sky130_fd_pr__pfet_01v8 ad=6.0645 pd=31.88 as=0 ps=0 w=15.55 l=2.63
X7 B.t2 B.t0 B.t1 w_n2154_n4078# sky130_fd_pr__pfet_01v8 ad=6.0645 pd=31.88 as=0 ps=0 w=15.55 l=2.63
R0 VP.n0 VP.t1 231.014
R1 VP.n0 VP.t0 183.589
R2 VP VP.n0 0.431811
R3 VTAIL.n338 VTAIL.n258 756.745
R4 VTAIL.n80 VTAIL.n0 756.745
R5 VTAIL.n252 VTAIL.n172 756.745
R6 VTAIL.n166 VTAIL.n86 756.745
R7 VTAIL.n287 VTAIL.n286 585
R8 VTAIL.n289 VTAIL.n288 585
R9 VTAIL.n282 VTAIL.n281 585
R10 VTAIL.n295 VTAIL.n294 585
R11 VTAIL.n297 VTAIL.n296 585
R12 VTAIL.n278 VTAIL.n277 585
R13 VTAIL.n303 VTAIL.n302 585
R14 VTAIL.n305 VTAIL.n304 585
R15 VTAIL.n274 VTAIL.n273 585
R16 VTAIL.n311 VTAIL.n310 585
R17 VTAIL.n313 VTAIL.n312 585
R18 VTAIL.n270 VTAIL.n269 585
R19 VTAIL.n319 VTAIL.n318 585
R20 VTAIL.n321 VTAIL.n320 585
R21 VTAIL.n266 VTAIL.n265 585
R22 VTAIL.n328 VTAIL.n327 585
R23 VTAIL.n329 VTAIL.n264 585
R24 VTAIL.n331 VTAIL.n330 585
R25 VTAIL.n262 VTAIL.n261 585
R26 VTAIL.n337 VTAIL.n336 585
R27 VTAIL.n339 VTAIL.n338 585
R28 VTAIL.n29 VTAIL.n28 585
R29 VTAIL.n31 VTAIL.n30 585
R30 VTAIL.n24 VTAIL.n23 585
R31 VTAIL.n37 VTAIL.n36 585
R32 VTAIL.n39 VTAIL.n38 585
R33 VTAIL.n20 VTAIL.n19 585
R34 VTAIL.n45 VTAIL.n44 585
R35 VTAIL.n47 VTAIL.n46 585
R36 VTAIL.n16 VTAIL.n15 585
R37 VTAIL.n53 VTAIL.n52 585
R38 VTAIL.n55 VTAIL.n54 585
R39 VTAIL.n12 VTAIL.n11 585
R40 VTAIL.n61 VTAIL.n60 585
R41 VTAIL.n63 VTAIL.n62 585
R42 VTAIL.n8 VTAIL.n7 585
R43 VTAIL.n70 VTAIL.n69 585
R44 VTAIL.n71 VTAIL.n6 585
R45 VTAIL.n73 VTAIL.n72 585
R46 VTAIL.n4 VTAIL.n3 585
R47 VTAIL.n79 VTAIL.n78 585
R48 VTAIL.n81 VTAIL.n80 585
R49 VTAIL.n253 VTAIL.n252 585
R50 VTAIL.n251 VTAIL.n250 585
R51 VTAIL.n176 VTAIL.n175 585
R52 VTAIL.n180 VTAIL.n178 585
R53 VTAIL.n245 VTAIL.n244 585
R54 VTAIL.n243 VTAIL.n242 585
R55 VTAIL.n182 VTAIL.n181 585
R56 VTAIL.n237 VTAIL.n236 585
R57 VTAIL.n235 VTAIL.n234 585
R58 VTAIL.n186 VTAIL.n185 585
R59 VTAIL.n229 VTAIL.n228 585
R60 VTAIL.n227 VTAIL.n226 585
R61 VTAIL.n190 VTAIL.n189 585
R62 VTAIL.n221 VTAIL.n220 585
R63 VTAIL.n219 VTAIL.n218 585
R64 VTAIL.n194 VTAIL.n193 585
R65 VTAIL.n213 VTAIL.n212 585
R66 VTAIL.n211 VTAIL.n210 585
R67 VTAIL.n198 VTAIL.n197 585
R68 VTAIL.n205 VTAIL.n204 585
R69 VTAIL.n203 VTAIL.n202 585
R70 VTAIL.n167 VTAIL.n166 585
R71 VTAIL.n165 VTAIL.n164 585
R72 VTAIL.n90 VTAIL.n89 585
R73 VTAIL.n94 VTAIL.n92 585
R74 VTAIL.n159 VTAIL.n158 585
R75 VTAIL.n157 VTAIL.n156 585
R76 VTAIL.n96 VTAIL.n95 585
R77 VTAIL.n151 VTAIL.n150 585
R78 VTAIL.n149 VTAIL.n148 585
R79 VTAIL.n100 VTAIL.n99 585
R80 VTAIL.n143 VTAIL.n142 585
R81 VTAIL.n141 VTAIL.n140 585
R82 VTAIL.n104 VTAIL.n103 585
R83 VTAIL.n135 VTAIL.n134 585
R84 VTAIL.n133 VTAIL.n132 585
R85 VTAIL.n108 VTAIL.n107 585
R86 VTAIL.n127 VTAIL.n126 585
R87 VTAIL.n125 VTAIL.n124 585
R88 VTAIL.n112 VTAIL.n111 585
R89 VTAIL.n119 VTAIL.n118 585
R90 VTAIL.n117 VTAIL.n116 585
R91 VTAIL.n285 VTAIL.t0 327.466
R92 VTAIL.n27 VTAIL.t2 327.466
R93 VTAIL.n201 VTAIL.t3 327.466
R94 VTAIL.n115 VTAIL.t1 327.466
R95 VTAIL.n288 VTAIL.n287 171.744
R96 VTAIL.n288 VTAIL.n281 171.744
R97 VTAIL.n295 VTAIL.n281 171.744
R98 VTAIL.n296 VTAIL.n295 171.744
R99 VTAIL.n296 VTAIL.n277 171.744
R100 VTAIL.n303 VTAIL.n277 171.744
R101 VTAIL.n304 VTAIL.n303 171.744
R102 VTAIL.n304 VTAIL.n273 171.744
R103 VTAIL.n311 VTAIL.n273 171.744
R104 VTAIL.n312 VTAIL.n311 171.744
R105 VTAIL.n312 VTAIL.n269 171.744
R106 VTAIL.n319 VTAIL.n269 171.744
R107 VTAIL.n320 VTAIL.n319 171.744
R108 VTAIL.n320 VTAIL.n265 171.744
R109 VTAIL.n328 VTAIL.n265 171.744
R110 VTAIL.n329 VTAIL.n328 171.744
R111 VTAIL.n330 VTAIL.n329 171.744
R112 VTAIL.n330 VTAIL.n261 171.744
R113 VTAIL.n337 VTAIL.n261 171.744
R114 VTAIL.n338 VTAIL.n337 171.744
R115 VTAIL.n30 VTAIL.n29 171.744
R116 VTAIL.n30 VTAIL.n23 171.744
R117 VTAIL.n37 VTAIL.n23 171.744
R118 VTAIL.n38 VTAIL.n37 171.744
R119 VTAIL.n38 VTAIL.n19 171.744
R120 VTAIL.n45 VTAIL.n19 171.744
R121 VTAIL.n46 VTAIL.n45 171.744
R122 VTAIL.n46 VTAIL.n15 171.744
R123 VTAIL.n53 VTAIL.n15 171.744
R124 VTAIL.n54 VTAIL.n53 171.744
R125 VTAIL.n54 VTAIL.n11 171.744
R126 VTAIL.n61 VTAIL.n11 171.744
R127 VTAIL.n62 VTAIL.n61 171.744
R128 VTAIL.n62 VTAIL.n7 171.744
R129 VTAIL.n70 VTAIL.n7 171.744
R130 VTAIL.n71 VTAIL.n70 171.744
R131 VTAIL.n72 VTAIL.n71 171.744
R132 VTAIL.n72 VTAIL.n3 171.744
R133 VTAIL.n79 VTAIL.n3 171.744
R134 VTAIL.n80 VTAIL.n79 171.744
R135 VTAIL.n252 VTAIL.n251 171.744
R136 VTAIL.n251 VTAIL.n175 171.744
R137 VTAIL.n180 VTAIL.n175 171.744
R138 VTAIL.n244 VTAIL.n180 171.744
R139 VTAIL.n244 VTAIL.n243 171.744
R140 VTAIL.n243 VTAIL.n181 171.744
R141 VTAIL.n236 VTAIL.n181 171.744
R142 VTAIL.n236 VTAIL.n235 171.744
R143 VTAIL.n235 VTAIL.n185 171.744
R144 VTAIL.n228 VTAIL.n185 171.744
R145 VTAIL.n228 VTAIL.n227 171.744
R146 VTAIL.n227 VTAIL.n189 171.744
R147 VTAIL.n220 VTAIL.n189 171.744
R148 VTAIL.n220 VTAIL.n219 171.744
R149 VTAIL.n219 VTAIL.n193 171.744
R150 VTAIL.n212 VTAIL.n193 171.744
R151 VTAIL.n212 VTAIL.n211 171.744
R152 VTAIL.n211 VTAIL.n197 171.744
R153 VTAIL.n204 VTAIL.n197 171.744
R154 VTAIL.n204 VTAIL.n203 171.744
R155 VTAIL.n166 VTAIL.n165 171.744
R156 VTAIL.n165 VTAIL.n89 171.744
R157 VTAIL.n94 VTAIL.n89 171.744
R158 VTAIL.n158 VTAIL.n94 171.744
R159 VTAIL.n158 VTAIL.n157 171.744
R160 VTAIL.n157 VTAIL.n95 171.744
R161 VTAIL.n150 VTAIL.n95 171.744
R162 VTAIL.n150 VTAIL.n149 171.744
R163 VTAIL.n149 VTAIL.n99 171.744
R164 VTAIL.n142 VTAIL.n99 171.744
R165 VTAIL.n142 VTAIL.n141 171.744
R166 VTAIL.n141 VTAIL.n103 171.744
R167 VTAIL.n134 VTAIL.n103 171.744
R168 VTAIL.n134 VTAIL.n133 171.744
R169 VTAIL.n133 VTAIL.n107 171.744
R170 VTAIL.n126 VTAIL.n107 171.744
R171 VTAIL.n126 VTAIL.n125 171.744
R172 VTAIL.n125 VTAIL.n111 171.744
R173 VTAIL.n118 VTAIL.n111 171.744
R174 VTAIL.n118 VTAIL.n117 171.744
R175 VTAIL.n287 VTAIL.t0 85.8723
R176 VTAIL.n29 VTAIL.t2 85.8723
R177 VTAIL.n203 VTAIL.t3 85.8723
R178 VTAIL.n117 VTAIL.t1 85.8723
R179 VTAIL.n343 VTAIL.n342 35.8702
R180 VTAIL.n85 VTAIL.n84 35.8702
R181 VTAIL.n257 VTAIL.n256 35.8702
R182 VTAIL.n171 VTAIL.n170 35.8702
R183 VTAIL.n171 VTAIL.n85 30.8755
R184 VTAIL.n343 VTAIL.n257 28.3238
R185 VTAIL.n286 VTAIL.n285 16.3895
R186 VTAIL.n28 VTAIL.n27 16.3895
R187 VTAIL.n202 VTAIL.n201 16.3895
R188 VTAIL.n116 VTAIL.n115 16.3895
R189 VTAIL.n331 VTAIL.n262 13.1884
R190 VTAIL.n73 VTAIL.n4 13.1884
R191 VTAIL.n178 VTAIL.n176 13.1884
R192 VTAIL.n92 VTAIL.n90 13.1884
R193 VTAIL.n289 VTAIL.n284 12.8005
R194 VTAIL.n332 VTAIL.n264 12.8005
R195 VTAIL.n336 VTAIL.n335 12.8005
R196 VTAIL.n31 VTAIL.n26 12.8005
R197 VTAIL.n74 VTAIL.n6 12.8005
R198 VTAIL.n78 VTAIL.n77 12.8005
R199 VTAIL.n250 VTAIL.n249 12.8005
R200 VTAIL.n246 VTAIL.n245 12.8005
R201 VTAIL.n205 VTAIL.n200 12.8005
R202 VTAIL.n164 VTAIL.n163 12.8005
R203 VTAIL.n160 VTAIL.n159 12.8005
R204 VTAIL.n119 VTAIL.n114 12.8005
R205 VTAIL.n290 VTAIL.n282 12.0247
R206 VTAIL.n327 VTAIL.n326 12.0247
R207 VTAIL.n339 VTAIL.n260 12.0247
R208 VTAIL.n32 VTAIL.n24 12.0247
R209 VTAIL.n69 VTAIL.n68 12.0247
R210 VTAIL.n81 VTAIL.n2 12.0247
R211 VTAIL.n253 VTAIL.n174 12.0247
R212 VTAIL.n242 VTAIL.n179 12.0247
R213 VTAIL.n206 VTAIL.n198 12.0247
R214 VTAIL.n167 VTAIL.n88 12.0247
R215 VTAIL.n156 VTAIL.n93 12.0247
R216 VTAIL.n120 VTAIL.n112 12.0247
R217 VTAIL.n294 VTAIL.n293 11.249
R218 VTAIL.n325 VTAIL.n266 11.249
R219 VTAIL.n340 VTAIL.n258 11.249
R220 VTAIL.n36 VTAIL.n35 11.249
R221 VTAIL.n67 VTAIL.n8 11.249
R222 VTAIL.n82 VTAIL.n0 11.249
R223 VTAIL.n254 VTAIL.n172 11.249
R224 VTAIL.n241 VTAIL.n182 11.249
R225 VTAIL.n210 VTAIL.n209 11.249
R226 VTAIL.n168 VTAIL.n86 11.249
R227 VTAIL.n155 VTAIL.n96 11.249
R228 VTAIL.n124 VTAIL.n123 11.249
R229 VTAIL.n297 VTAIL.n280 10.4732
R230 VTAIL.n322 VTAIL.n321 10.4732
R231 VTAIL.n39 VTAIL.n22 10.4732
R232 VTAIL.n64 VTAIL.n63 10.4732
R233 VTAIL.n238 VTAIL.n237 10.4732
R234 VTAIL.n213 VTAIL.n196 10.4732
R235 VTAIL.n152 VTAIL.n151 10.4732
R236 VTAIL.n127 VTAIL.n110 10.4732
R237 VTAIL.n298 VTAIL.n278 9.69747
R238 VTAIL.n318 VTAIL.n268 9.69747
R239 VTAIL.n40 VTAIL.n20 9.69747
R240 VTAIL.n60 VTAIL.n10 9.69747
R241 VTAIL.n234 VTAIL.n184 9.69747
R242 VTAIL.n214 VTAIL.n194 9.69747
R243 VTAIL.n148 VTAIL.n98 9.69747
R244 VTAIL.n128 VTAIL.n108 9.69747
R245 VTAIL.n342 VTAIL.n341 9.45567
R246 VTAIL.n84 VTAIL.n83 9.45567
R247 VTAIL.n256 VTAIL.n255 9.45567
R248 VTAIL.n170 VTAIL.n169 9.45567
R249 VTAIL.n341 VTAIL.n340 9.3005
R250 VTAIL.n260 VTAIL.n259 9.3005
R251 VTAIL.n335 VTAIL.n334 9.3005
R252 VTAIL.n307 VTAIL.n306 9.3005
R253 VTAIL.n276 VTAIL.n275 9.3005
R254 VTAIL.n301 VTAIL.n300 9.3005
R255 VTAIL.n299 VTAIL.n298 9.3005
R256 VTAIL.n280 VTAIL.n279 9.3005
R257 VTAIL.n293 VTAIL.n292 9.3005
R258 VTAIL.n291 VTAIL.n290 9.3005
R259 VTAIL.n284 VTAIL.n283 9.3005
R260 VTAIL.n309 VTAIL.n308 9.3005
R261 VTAIL.n272 VTAIL.n271 9.3005
R262 VTAIL.n315 VTAIL.n314 9.3005
R263 VTAIL.n317 VTAIL.n316 9.3005
R264 VTAIL.n268 VTAIL.n267 9.3005
R265 VTAIL.n323 VTAIL.n322 9.3005
R266 VTAIL.n325 VTAIL.n324 9.3005
R267 VTAIL.n326 VTAIL.n263 9.3005
R268 VTAIL.n333 VTAIL.n332 9.3005
R269 VTAIL.n83 VTAIL.n82 9.3005
R270 VTAIL.n2 VTAIL.n1 9.3005
R271 VTAIL.n77 VTAIL.n76 9.3005
R272 VTAIL.n49 VTAIL.n48 9.3005
R273 VTAIL.n18 VTAIL.n17 9.3005
R274 VTAIL.n43 VTAIL.n42 9.3005
R275 VTAIL.n41 VTAIL.n40 9.3005
R276 VTAIL.n22 VTAIL.n21 9.3005
R277 VTAIL.n35 VTAIL.n34 9.3005
R278 VTAIL.n33 VTAIL.n32 9.3005
R279 VTAIL.n26 VTAIL.n25 9.3005
R280 VTAIL.n51 VTAIL.n50 9.3005
R281 VTAIL.n14 VTAIL.n13 9.3005
R282 VTAIL.n57 VTAIL.n56 9.3005
R283 VTAIL.n59 VTAIL.n58 9.3005
R284 VTAIL.n10 VTAIL.n9 9.3005
R285 VTAIL.n65 VTAIL.n64 9.3005
R286 VTAIL.n67 VTAIL.n66 9.3005
R287 VTAIL.n68 VTAIL.n5 9.3005
R288 VTAIL.n75 VTAIL.n74 9.3005
R289 VTAIL.n188 VTAIL.n187 9.3005
R290 VTAIL.n231 VTAIL.n230 9.3005
R291 VTAIL.n233 VTAIL.n232 9.3005
R292 VTAIL.n184 VTAIL.n183 9.3005
R293 VTAIL.n239 VTAIL.n238 9.3005
R294 VTAIL.n241 VTAIL.n240 9.3005
R295 VTAIL.n179 VTAIL.n177 9.3005
R296 VTAIL.n247 VTAIL.n246 9.3005
R297 VTAIL.n255 VTAIL.n254 9.3005
R298 VTAIL.n174 VTAIL.n173 9.3005
R299 VTAIL.n249 VTAIL.n248 9.3005
R300 VTAIL.n225 VTAIL.n224 9.3005
R301 VTAIL.n223 VTAIL.n222 9.3005
R302 VTAIL.n192 VTAIL.n191 9.3005
R303 VTAIL.n217 VTAIL.n216 9.3005
R304 VTAIL.n215 VTAIL.n214 9.3005
R305 VTAIL.n196 VTAIL.n195 9.3005
R306 VTAIL.n209 VTAIL.n208 9.3005
R307 VTAIL.n207 VTAIL.n206 9.3005
R308 VTAIL.n200 VTAIL.n199 9.3005
R309 VTAIL.n102 VTAIL.n101 9.3005
R310 VTAIL.n145 VTAIL.n144 9.3005
R311 VTAIL.n147 VTAIL.n146 9.3005
R312 VTAIL.n98 VTAIL.n97 9.3005
R313 VTAIL.n153 VTAIL.n152 9.3005
R314 VTAIL.n155 VTAIL.n154 9.3005
R315 VTAIL.n93 VTAIL.n91 9.3005
R316 VTAIL.n161 VTAIL.n160 9.3005
R317 VTAIL.n169 VTAIL.n168 9.3005
R318 VTAIL.n88 VTAIL.n87 9.3005
R319 VTAIL.n163 VTAIL.n162 9.3005
R320 VTAIL.n139 VTAIL.n138 9.3005
R321 VTAIL.n137 VTAIL.n136 9.3005
R322 VTAIL.n106 VTAIL.n105 9.3005
R323 VTAIL.n131 VTAIL.n130 9.3005
R324 VTAIL.n129 VTAIL.n128 9.3005
R325 VTAIL.n110 VTAIL.n109 9.3005
R326 VTAIL.n123 VTAIL.n122 9.3005
R327 VTAIL.n121 VTAIL.n120 9.3005
R328 VTAIL.n114 VTAIL.n113 9.3005
R329 VTAIL.n302 VTAIL.n301 8.92171
R330 VTAIL.n317 VTAIL.n270 8.92171
R331 VTAIL.n44 VTAIL.n43 8.92171
R332 VTAIL.n59 VTAIL.n12 8.92171
R333 VTAIL.n233 VTAIL.n186 8.92171
R334 VTAIL.n218 VTAIL.n217 8.92171
R335 VTAIL.n147 VTAIL.n100 8.92171
R336 VTAIL.n132 VTAIL.n131 8.92171
R337 VTAIL.n305 VTAIL.n276 8.14595
R338 VTAIL.n314 VTAIL.n313 8.14595
R339 VTAIL.n47 VTAIL.n18 8.14595
R340 VTAIL.n56 VTAIL.n55 8.14595
R341 VTAIL.n230 VTAIL.n229 8.14595
R342 VTAIL.n221 VTAIL.n192 8.14595
R343 VTAIL.n144 VTAIL.n143 8.14595
R344 VTAIL.n135 VTAIL.n106 8.14595
R345 VTAIL.n306 VTAIL.n274 7.3702
R346 VTAIL.n310 VTAIL.n272 7.3702
R347 VTAIL.n48 VTAIL.n16 7.3702
R348 VTAIL.n52 VTAIL.n14 7.3702
R349 VTAIL.n226 VTAIL.n188 7.3702
R350 VTAIL.n222 VTAIL.n190 7.3702
R351 VTAIL.n140 VTAIL.n102 7.3702
R352 VTAIL.n136 VTAIL.n104 7.3702
R353 VTAIL.n309 VTAIL.n274 6.59444
R354 VTAIL.n310 VTAIL.n309 6.59444
R355 VTAIL.n51 VTAIL.n16 6.59444
R356 VTAIL.n52 VTAIL.n51 6.59444
R357 VTAIL.n226 VTAIL.n225 6.59444
R358 VTAIL.n225 VTAIL.n190 6.59444
R359 VTAIL.n140 VTAIL.n139 6.59444
R360 VTAIL.n139 VTAIL.n104 6.59444
R361 VTAIL.n306 VTAIL.n305 5.81868
R362 VTAIL.n313 VTAIL.n272 5.81868
R363 VTAIL.n48 VTAIL.n47 5.81868
R364 VTAIL.n55 VTAIL.n14 5.81868
R365 VTAIL.n229 VTAIL.n188 5.81868
R366 VTAIL.n222 VTAIL.n221 5.81868
R367 VTAIL.n143 VTAIL.n102 5.81868
R368 VTAIL.n136 VTAIL.n135 5.81868
R369 VTAIL.n302 VTAIL.n276 5.04292
R370 VTAIL.n314 VTAIL.n270 5.04292
R371 VTAIL.n44 VTAIL.n18 5.04292
R372 VTAIL.n56 VTAIL.n12 5.04292
R373 VTAIL.n230 VTAIL.n186 5.04292
R374 VTAIL.n218 VTAIL.n192 5.04292
R375 VTAIL.n144 VTAIL.n100 5.04292
R376 VTAIL.n132 VTAIL.n106 5.04292
R377 VTAIL.n301 VTAIL.n278 4.26717
R378 VTAIL.n318 VTAIL.n317 4.26717
R379 VTAIL.n43 VTAIL.n20 4.26717
R380 VTAIL.n60 VTAIL.n59 4.26717
R381 VTAIL.n234 VTAIL.n233 4.26717
R382 VTAIL.n217 VTAIL.n194 4.26717
R383 VTAIL.n148 VTAIL.n147 4.26717
R384 VTAIL.n131 VTAIL.n108 4.26717
R385 VTAIL.n285 VTAIL.n283 3.70982
R386 VTAIL.n27 VTAIL.n25 3.70982
R387 VTAIL.n201 VTAIL.n199 3.70982
R388 VTAIL.n115 VTAIL.n113 3.70982
R389 VTAIL.n298 VTAIL.n297 3.49141
R390 VTAIL.n321 VTAIL.n268 3.49141
R391 VTAIL.n40 VTAIL.n39 3.49141
R392 VTAIL.n63 VTAIL.n10 3.49141
R393 VTAIL.n237 VTAIL.n184 3.49141
R394 VTAIL.n214 VTAIL.n213 3.49141
R395 VTAIL.n151 VTAIL.n98 3.49141
R396 VTAIL.n128 VTAIL.n127 3.49141
R397 VTAIL.n294 VTAIL.n280 2.71565
R398 VTAIL.n322 VTAIL.n266 2.71565
R399 VTAIL.n342 VTAIL.n258 2.71565
R400 VTAIL.n36 VTAIL.n22 2.71565
R401 VTAIL.n64 VTAIL.n8 2.71565
R402 VTAIL.n84 VTAIL.n0 2.71565
R403 VTAIL.n256 VTAIL.n172 2.71565
R404 VTAIL.n238 VTAIL.n182 2.71565
R405 VTAIL.n210 VTAIL.n196 2.71565
R406 VTAIL.n170 VTAIL.n86 2.71565
R407 VTAIL.n152 VTAIL.n96 2.71565
R408 VTAIL.n124 VTAIL.n110 2.71565
R409 VTAIL.n293 VTAIL.n282 1.93989
R410 VTAIL.n327 VTAIL.n325 1.93989
R411 VTAIL.n340 VTAIL.n339 1.93989
R412 VTAIL.n35 VTAIL.n24 1.93989
R413 VTAIL.n69 VTAIL.n67 1.93989
R414 VTAIL.n82 VTAIL.n81 1.93989
R415 VTAIL.n254 VTAIL.n253 1.93989
R416 VTAIL.n242 VTAIL.n241 1.93989
R417 VTAIL.n209 VTAIL.n198 1.93989
R418 VTAIL.n168 VTAIL.n167 1.93989
R419 VTAIL.n156 VTAIL.n155 1.93989
R420 VTAIL.n123 VTAIL.n112 1.93989
R421 VTAIL.n257 VTAIL.n171 1.74619
R422 VTAIL VTAIL.n85 1.16645
R423 VTAIL.n290 VTAIL.n289 1.16414
R424 VTAIL.n326 VTAIL.n264 1.16414
R425 VTAIL.n336 VTAIL.n260 1.16414
R426 VTAIL.n32 VTAIL.n31 1.16414
R427 VTAIL.n68 VTAIL.n6 1.16414
R428 VTAIL.n78 VTAIL.n2 1.16414
R429 VTAIL.n250 VTAIL.n174 1.16414
R430 VTAIL.n245 VTAIL.n179 1.16414
R431 VTAIL.n206 VTAIL.n205 1.16414
R432 VTAIL.n164 VTAIL.n88 1.16414
R433 VTAIL.n159 VTAIL.n93 1.16414
R434 VTAIL.n120 VTAIL.n119 1.16414
R435 VTAIL VTAIL.n343 0.580241
R436 VTAIL.n286 VTAIL.n284 0.388379
R437 VTAIL.n332 VTAIL.n331 0.388379
R438 VTAIL.n335 VTAIL.n262 0.388379
R439 VTAIL.n28 VTAIL.n26 0.388379
R440 VTAIL.n74 VTAIL.n73 0.388379
R441 VTAIL.n77 VTAIL.n4 0.388379
R442 VTAIL.n249 VTAIL.n176 0.388379
R443 VTAIL.n246 VTAIL.n178 0.388379
R444 VTAIL.n202 VTAIL.n200 0.388379
R445 VTAIL.n163 VTAIL.n90 0.388379
R446 VTAIL.n160 VTAIL.n92 0.388379
R447 VTAIL.n116 VTAIL.n114 0.388379
R448 VTAIL.n291 VTAIL.n283 0.155672
R449 VTAIL.n292 VTAIL.n291 0.155672
R450 VTAIL.n292 VTAIL.n279 0.155672
R451 VTAIL.n299 VTAIL.n279 0.155672
R452 VTAIL.n300 VTAIL.n299 0.155672
R453 VTAIL.n300 VTAIL.n275 0.155672
R454 VTAIL.n307 VTAIL.n275 0.155672
R455 VTAIL.n308 VTAIL.n307 0.155672
R456 VTAIL.n308 VTAIL.n271 0.155672
R457 VTAIL.n315 VTAIL.n271 0.155672
R458 VTAIL.n316 VTAIL.n315 0.155672
R459 VTAIL.n316 VTAIL.n267 0.155672
R460 VTAIL.n323 VTAIL.n267 0.155672
R461 VTAIL.n324 VTAIL.n323 0.155672
R462 VTAIL.n324 VTAIL.n263 0.155672
R463 VTAIL.n333 VTAIL.n263 0.155672
R464 VTAIL.n334 VTAIL.n333 0.155672
R465 VTAIL.n334 VTAIL.n259 0.155672
R466 VTAIL.n341 VTAIL.n259 0.155672
R467 VTAIL.n33 VTAIL.n25 0.155672
R468 VTAIL.n34 VTAIL.n33 0.155672
R469 VTAIL.n34 VTAIL.n21 0.155672
R470 VTAIL.n41 VTAIL.n21 0.155672
R471 VTAIL.n42 VTAIL.n41 0.155672
R472 VTAIL.n42 VTAIL.n17 0.155672
R473 VTAIL.n49 VTAIL.n17 0.155672
R474 VTAIL.n50 VTAIL.n49 0.155672
R475 VTAIL.n50 VTAIL.n13 0.155672
R476 VTAIL.n57 VTAIL.n13 0.155672
R477 VTAIL.n58 VTAIL.n57 0.155672
R478 VTAIL.n58 VTAIL.n9 0.155672
R479 VTAIL.n65 VTAIL.n9 0.155672
R480 VTAIL.n66 VTAIL.n65 0.155672
R481 VTAIL.n66 VTAIL.n5 0.155672
R482 VTAIL.n75 VTAIL.n5 0.155672
R483 VTAIL.n76 VTAIL.n75 0.155672
R484 VTAIL.n76 VTAIL.n1 0.155672
R485 VTAIL.n83 VTAIL.n1 0.155672
R486 VTAIL.n255 VTAIL.n173 0.155672
R487 VTAIL.n248 VTAIL.n173 0.155672
R488 VTAIL.n248 VTAIL.n247 0.155672
R489 VTAIL.n247 VTAIL.n177 0.155672
R490 VTAIL.n240 VTAIL.n177 0.155672
R491 VTAIL.n240 VTAIL.n239 0.155672
R492 VTAIL.n239 VTAIL.n183 0.155672
R493 VTAIL.n232 VTAIL.n183 0.155672
R494 VTAIL.n232 VTAIL.n231 0.155672
R495 VTAIL.n231 VTAIL.n187 0.155672
R496 VTAIL.n224 VTAIL.n187 0.155672
R497 VTAIL.n224 VTAIL.n223 0.155672
R498 VTAIL.n223 VTAIL.n191 0.155672
R499 VTAIL.n216 VTAIL.n191 0.155672
R500 VTAIL.n216 VTAIL.n215 0.155672
R501 VTAIL.n215 VTAIL.n195 0.155672
R502 VTAIL.n208 VTAIL.n195 0.155672
R503 VTAIL.n208 VTAIL.n207 0.155672
R504 VTAIL.n207 VTAIL.n199 0.155672
R505 VTAIL.n169 VTAIL.n87 0.155672
R506 VTAIL.n162 VTAIL.n87 0.155672
R507 VTAIL.n162 VTAIL.n161 0.155672
R508 VTAIL.n161 VTAIL.n91 0.155672
R509 VTAIL.n154 VTAIL.n91 0.155672
R510 VTAIL.n154 VTAIL.n153 0.155672
R511 VTAIL.n153 VTAIL.n97 0.155672
R512 VTAIL.n146 VTAIL.n97 0.155672
R513 VTAIL.n146 VTAIL.n145 0.155672
R514 VTAIL.n145 VTAIL.n101 0.155672
R515 VTAIL.n138 VTAIL.n101 0.155672
R516 VTAIL.n138 VTAIL.n137 0.155672
R517 VTAIL.n137 VTAIL.n105 0.155672
R518 VTAIL.n130 VTAIL.n105 0.155672
R519 VTAIL.n130 VTAIL.n129 0.155672
R520 VTAIL.n129 VTAIL.n109 0.155672
R521 VTAIL.n122 VTAIL.n109 0.155672
R522 VTAIL.n122 VTAIL.n121 0.155672
R523 VTAIL.n121 VTAIL.n113 0.155672
R524 VDD1.n80 VDD1.n0 756.745
R525 VDD1.n165 VDD1.n85 756.745
R526 VDD1.n81 VDD1.n80 585
R527 VDD1.n79 VDD1.n78 585
R528 VDD1.n4 VDD1.n3 585
R529 VDD1.n8 VDD1.n6 585
R530 VDD1.n73 VDD1.n72 585
R531 VDD1.n71 VDD1.n70 585
R532 VDD1.n10 VDD1.n9 585
R533 VDD1.n65 VDD1.n64 585
R534 VDD1.n63 VDD1.n62 585
R535 VDD1.n14 VDD1.n13 585
R536 VDD1.n57 VDD1.n56 585
R537 VDD1.n55 VDD1.n54 585
R538 VDD1.n18 VDD1.n17 585
R539 VDD1.n49 VDD1.n48 585
R540 VDD1.n47 VDD1.n46 585
R541 VDD1.n22 VDD1.n21 585
R542 VDD1.n41 VDD1.n40 585
R543 VDD1.n39 VDD1.n38 585
R544 VDD1.n26 VDD1.n25 585
R545 VDD1.n33 VDD1.n32 585
R546 VDD1.n31 VDD1.n30 585
R547 VDD1.n114 VDD1.n113 585
R548 VDD1.n116 VDD1.n115 585
R549 VDD1.n109 VDD1.n108 585
R550 VDD1.n122 VDD1.n121 585
R551 VDD1.n124 VDD1.n123 585
R552 VDD1.n105 VDD1.n104 585
R553 VDD1.n130 VDD1.n129 585
R554 VDD1.n132 VDD1.n131 585
R555 VDD1.n101 VDD1.n100 585
R556 VDD1.n138 VDD1.n137 585
R557 VDD1.n140 VDD1.n139 585
R558 VDD1.n97 VDD1.n96 585
R559 VDD1.n146 VDD1.n145 585
R560 VDD1.n148 VDD1.n147 585
R561 VDD1.n93 VDD1.n92 585
R562 VDD1.n155 VDD1.n154 585
R563 VDD1.n156 VDD1.n91 585
R564 VDD1.n158 VDD1.n157 585
R565 VDD1.n89 VDD1.n88 585
R566 VDD1.n164 VDD1.n163 585
R567 VDD1.n166 VDD1.n165 585
R568 VDD1.n29 VDD1.t0 327.466
R569 VDD1.n112 VDD1.t1 327.466
R570 VDD1.n80 VDD1.n79 171.744
R571 VDD1.n79 VDD1.n3 171.744
R572 VDD1.n8 VDD1.n3 171.744
R573 VDD1.n72 VDD1.n8 171.744
R574 VDD1.n72 VDD1.n71 171.744
R575 VDD1.n71 VDD1.n9 171.744
R576 VDD1.n64 VDD1.n9 171.744
R577 VDD1.n64 VDD1.n63 171.744
R578 VDD1.n63 VDD1.n13 171.744
R579 VDD1.n56 VDD1.n13 171.744
R580 VDD1.n56 VDD1.n55 171.744
R581 VDD1.n55 VDD1.n17 171.744
R582 VDD1.n48 VDD1.n17 171.744
R583 VDD1.n48 VDD1.n47 171.744
R584 VDD1.n47 VDD1.n21 171.744
R585 VDD1.n40 VDD1.n21 171.744
R586 VDD1.n40 VDD1.n39 171.744
R587 VDD1.n39 VDD1.n25 171.744
R588 VDD1.n32 VDD1.n25 171.744
R589 VDD1.n32 VDD1.n31 171.744
R590 VDD1.n115 VDD1.n114 171.744
R591 VDD1.n115 VDD1.n108 171.744
R592 VDD1.n122 VDD1.n108 171.744
R593 VDD1.n123 VDD1.n122 171.744
R594 VDD1.n123 VDD1.n104 171.744
R595 VDD1.n130 VDD1.n104 171.744
R596 VDD1.n131 VDD1.n130 171.744
R597 VDD1.n131 VDD1.n100 171.744
R598 VDD1.n138 VDD1.n100 171.744
R599 VDD1.n139 VDD1.n138 171.744
R600 VDD1.n139 VDD1.n96 171.744
R601 VDD1.n146 VDD1.n96 171.744
R602 VDD1.n147 VDD1.n146 171.744
R603 VDD1.n147 VDD1.n92 171.744
R604 VDD1.n155 VDD1.n92 171.744
R605 VDD1.n156 VDD1.n155 171.744
R606 VDD1.n157 VDD1.n156 171.744
R607 VDD1.n157 VDD1.n88 171.744
R608 VDD1.n164 VDD1.n88 171.744
R609 VDD1.n165 VDD1.n164 171.744
R610 VDD1 VDD1.n169 95.8798
R611 VDD1.n31 VDD1.t0 85.8723
R612 VDD1.n114 VDD1.t1 85.8723
R613 VDD1 VDD1.n84 53.2451
R614 VDD1.n30 VDD1.n29 16.3895
R615 VDD1.n113 VDD1.n112 16.3895
R616 VDD1.n6 VDD1.n4 13.1884
R617 VDD1.n158 VDD1.n89 13.1884
R618 VDD1.n78 VDD1.n77 12.8005
R619 VDD1.n74 VDD1.n73 12.8005
R620 VDD1.n33 VDD1.n28 12.8005
R621 VDD1.n116 VDD1.n111 12.8005
R622 VDD1.n159 VDD1.n91 12.8005
R623 VDD1.n163 VDD1.n162 12.8005
R624 VDD1.n81 VDD1.n2 12.0247
R625 VDD1.n70 VDD1.n7 12.0247
R626 VDD1.n34 VDD1.n26 12.0247
R627 VDD1.n117 VDD1.n109 12.0247
R628 VDD1.n154 VDD1.n153 12.0247
R629 VDD1.n166 VDD1.n87 12.0247
R630 VDD1.n82 VDD1.n0 11.249
R631 VDD1.n69 VDD1.n10 11.249
R632 VDD1.n38 VDD1.n37 11.249
R633 VDD1.n121 VDD1.n120 11.249
R634 VDD1.n152 VDD1.n93 11.249
R635 VDD1.n167 VDD1.n85 11.249
R636 VDD1.n66 VDD1.n65 10.4732
R637 VDD1.n41 VDD1.n24 10.4732
R638 VDD1.n124 VDD1.n107 10.4732
R639 VDD1.n149 VDD1.n148 10.4732
R640 VDD1.n62 VDD1.n12 9.69747
R641 VDD1.n42 VDD1.n22 9.69747
R642 VDD1.n125 VDD1.n105 9.69747
R643 VDD1.n145 VDD1.n95 9.69747
R644 VDD1.n84 VDD1.n83 9.45567
R645 VDD1.n169 VDD1.n168 9.45567
R646 VDD1.n16 VDD1.n15 9.3005
R647 VDD1.n59 VDD1.n58 9.3005
R648 VDD1.n61 VDD1.n60 9.3005
R649 VDD1.n12 VDD1.n11 9.3005
R650 VDD1.n67 VDD1.n66 9.3005
R651 VDD1.n69 VDD1.n68 9.3005
R652 VDD1.n7 VDD1.n5 9.3005
R653 VDD1.n75 VDD1.n74 9.3005
R654 VDD1.n83 VDD1.n82 9.3005
R655 VDD1.n2 VDD1.n1 9.3005
R656 VDD1.n77 VDD1.n76 9.3005
R657 VDD1.n53 VDD1.n52 9.3005
R658 VDD1.n51 VDD1.n50 9.3005
R659 VDD1.n20 VDD1.n19 9.3005
R660 VDD1.n45 VDD1.n44 9.3005
R661 VDD1.n43 VDD1.n42 9.3005
R662 VDD1.n24 VDD1.n23 9.3005
R663 VDD1.n37 VDD1.n36 9.3005
R664 VDD1.n35 VDD1.n34 9.3005
R665 VDD1.n28 VDD1.n27 9.3005
R666 VDD1.n168 VDD1.n167 9.3005
R667 VDD1.n87 VDD1.n86 9.3005
R668 VDD1.n162 VDD1.n161 9.3005
R669 VDD1.n134 VDD1.n133 9.3005
R670 VDD1.n103 VDD1.n102 9.3005
R671 VDD1.n128 VDD1.n127 9.3005
R672 VDD1.n126 VDD1.n125 9.3005
R673 VDD1.n107 VDD1.n106 9.3005
R674 VDD1.n120 VDD1.n119 9.3005
R675 VDD1.n118 VDD1.n117 9.3005
R676 VDD1.n111 VDD1.n110 9.3005
R677 VDD1.n136 VDD1.n135 9.3005
R678 VDD1.n99 VDD1.n98 9.3005
R679 VDD1.n142 VDD1.n141 9.3005
R680 VDD1.n144 VDD1.n143 9.3005
R681 VDD1.n95 VDD1.n94 9.3005
R682 VDD1.n150 VDD1.n149 9.3005
R683 VDD1.n152 VDD1.n151 9.3005
R684 VDD1.n153 VDD1.n90 9.3005
R685 VDD1.n160 VDD1.n159 9.3005
R686 VDD1.n61 VDD1.n14 8.92171
R687 VDD1.n46 VDD1.n45 8.92171
R688 VDD1.n129 VDD1.n128 8.92171
R689 VDD1.n144 VDD1.n97 8.92171
R690 VDD1.n58 VDD1.n57 8.14595
R691 VDD1.n49 VDD1.n20 8.14595
R692 VDD1.n132 VDD1.n103 8.14595
R693 VDD1.n141 VDD1.n140 8.14595
R694 VDD1.n54 VDD1.n16 7.3702
R695 VDD1.n50 VDD1.n18 7.3702
R696 VDD1.n133 VDD1.n101 7.3702
R697 VDD1.n137 VDD1.n99 7.3702
R698 VDD1.n54 VDD1.n53 6.59444
R699 VDD1.n53 VDD1.n18 6.59444
R700 VDD1.n136 VDD1.n101 6.59444
R701 VDD1.n137 VDD1.n136 6.59444
R702 VDD1.n57 VDD1.n16 5.81868
R703 VDD1.n50 VDD1.n49 5.81868
R704 VDD1.n133 VDD1.n132 5.81868
R705 VDD1.n140 VDD1.n99 5.81868
R706 VDD1.n58 VDD1.n14 5.04292
R707 VDD1.n46 VDD1.n20 5.04292
R708 VDD1.n129 VDD1.n103 5.04292
R709 VDD1.n141 VDD1.n97 5.04292
R710 VDD1.n62 VDD1.n61 4.26717
R711 VDD1.n45 VDD1.n22 4.26717
R712 VDD1.n128 VDD1.n105 4.26717
R713 VDD1.n145 VDD1.n144 4.26717
R714 VDD1.n29 VDD1.n27 3.70982
R715 VDD1.n112 VDD1.n110 3.70982
R716 VDD1.n65 VDD1.n12 3.49141
R717 VDD1.n42 VDD1.n41 3.49141
R718 VDD1.n125 VDD1.n124 3.49141
R719 VDD1.n148 VDD1.n95 3.49141
R720 VDD1.n84 VDD1.n0 2.71565
R721 VDD1.n66 VDD1.n10 2.71565
R722 VDD1.n38 VDD1.n24 2.71565
R723 VDD1.n121 VDD1.n107 2.71565
R724 VDD1.n149 VDD1.n93 2.71565
R725 VDD1.n169 VDD1.n85 2.71565
R726 VDD1.n82 VDD1.n81 1.93989
R727 VDD1.n70 VDD1.n69 1.93989
R728 VDD1.n37 VDD1.n26 1.93989
R729 VDD1.n120 VDD1.n109 1.93989
R730 VDD1.n154 VDD1.n152 1.93989
R731 VDD1.n167 VDD1.n166 1.93989
R732 VDD1.n78 VDD1.n2 1.16414
R733 VDD1.n73 VDD1.n7 1.16414
R734 VDD1.n34 VDD1.n33 1.16414
R735 VDD1.n117 VDD1.n116 1.16414
R736 VDD1.n153 VDD1.n91 1.16414
R737 VDD1.n163 VDD1.n87 1.16414
R738 VDD1.n77 VDD1.n4 0.388379
R739 VDD1.n74 VDD1.n6 0.388379
R740 VDD1.n30 VDD1.n28 0.388379
R741 VDD1.n113 VDD1.n111 0.388379
R742 VDD1.n159 VDD1.n158 0.388379
R743 VDD1.n162 VDD1.n89 0.388379
R744 VDD1.n83 VDD1.n1 0.155672
R745 VDD1.n76 VDD1.n1 0.155672
R746 VDD1.n76 VDD1.n75 0.155672
R747 VDD1.n75 VDD1.n5 0.155672
R748 VDD1.n68 VDD1.n5 0.155672
R749 VDD1.n68 VDD1.n67 0.155672
R750 VDD1.n67 VDD1.n11 0.155672
R751 VDD1.n60 VDD1.n11 0.155672
R752 VDD1.n60 VDD1.n59 0.155672
R753 VDD1.n59 VDD1.n15 0.155672
R754 VDD1.n52 VDD1.n15 0.155672
R755 VDD1.n52 VDD1.n51 0.155672
R756 VDD1.n51 VDD1.n19 0.155672
R757 VDD1.n44 VDD1.n19 0.155672
R758 VDD1.n44 VDD1.n43 0.155672
R759 VDD1.n43 VDD1.n23 0.155672
R760 VDD1.n36 VDD1.n23 0.155672
R761 VDD1.n36 VDD1.n35 0.155672
R762 VDD1.n35 VDD1.n27 0.155672
R763 VDD1.n118 VDD1.n110 0.155672
R764 VDD1.n119 VDD1.n118 0.155672
R765 VDD1.n119 VDD1.n106 0.155672
R766 VDD1.n126 VDD1.n106 0.155672
R767 VDD1.n127 VDD1.n126 0.155672
R768 VDD1.n127 VDD1.n102 0.155672
R769 VDD1.n134 VDD1.n102 0.155672
R770 VDD1.n135 VDD1.n134 0.155672
R771 VDD1.n135 VDD1.n98 0.155672
R772 VDD1.n142 VDD1.n98 0.155672
R773 VDD1.n143 VDD1.n142 0.155672
R774 VDD1.n143 VDD1.n94 0.155672
R775 VDD1.n150 VDD1.n94 0.155672
R776 VDD1.n151 VDD1.n150 0.155672
R777 VDD1.n151 VDD1.n90 0.155672
R778 VDD1.n160 VDD1.n90 0.155672
R779 VDD1.n161 VDD1.n160 0.155672
R780 VDD1.n161 VDD1.n86 0.155672
R781 VDD1.n168 VDD1.n86 0.155672
R782 B.n384 B.n383 585
R783 B.n382 B.n103 585
R784 B.n381 B.n380 585
R785 B.n379 B.n104 585
R786 B.n378 B.n377 585
R787 B.n376 B.n105 585
R788 B.n375 B.n374 585
R789 B.n373 B.n106 585
R790 B.n372 B.n371 585
R791 B.n370 B.n107 585
R792 B.n369 B.n368 585
R793 B.n367 B.n108 585
R794 B.n366 B.n365 585
R795 B.n364 B.n109 585
R796 B.n363 B.n362 585
R797 B.n361 B.n110 585
R798 B.n360 B.n359 585
R799 B.n358 B.n111 585
R800 B.n357 B.n356 585
R801 B.n355 B.n112 585
R802 B.n354 B.n353 585
R803 B.n352 B.n113 585
R804 B.n351 B.n350 585
R805 B.n349 B.n114 585
R806 B.n348 B.n347 585
R807 B.n346 B.n115 585
R808 B.n345 B.n344 585
R809 B.n343 B.n116 585
R810 B.n342 B.n341 585
R811 B.n340 B.n117 585
R812 B.n339 B.n338 585
R813 B.n337 B.n118 585
R814 B.n336 B.n335 585
R815 B.n334 B.n119 585
R816 B.n333 B.n332 585
R817 B.n331 B.n120 585
R818 B.n330 B.n329 585
R819 B.n328 B.n121 585
R820 B.n327 B.n326 585
R821 B.n325 B.n122 585
R822 B.n324 B.n323 585
R823 B.n322 B.n123 585
R824 B.n321 B.n320 585
R825 B.n319 B.n124 585
R826 B.n318 B.n317 585
R827 B.n316 B.n125 585
R828 B.n315 B.n314 585
R829 B.n313 B.n126 585
R830 B.n312 B.n311 585
R831 B.n310 B.n127 585
R832 B.n309 B.n308 585
R833 B.n307 B.n128 585
R834 B.n305 B.n304 585
R835 B.n303 B.n131 585
R836 B.n302 B.n301 585
R837 B.n300 B.n132 585
R838 B.n299 B.n298 585
R839 B.n297 B.n133 585
R840 B.n296 B.n295 585
R841 B.n294 B.n134 585
R842 B.n293 B.n292 585
R843 B.n291 B.n135 585
R844 B.n290 B.n289 585
R845 B.n285 B.n136 585
R846 B.n284 B.n283 585
R847 B.n282 B.n137 585
R848 B.n281 B.n280 585
R849 B.n279 B.n138 585
R850 B.n278 B.n277 585
R851 B.n276 B.n139 585
R852 B.n275 B.n274 585
R853 B.n273 B.n140 585
R854 B.n272 B.n271 585
R855 B.n270 B.n141 585
R856 B.n269 B.n268 585
R857 B.n267 B.n142 585
R858 B.n266 B.n265 585
R859 B.n264 B.n143 585
R860 B.n263 B.n262 585
R861 B.n261 B.n144 585
R862 B.n260 B.n259 585
R863 B.n258 B.n145 585
R864 B.n257 B.n256 585
R865 B.n255 B.n146 585
R866 B.n254 B.n253 585
R867 B.n252 B.n147 585
R868 B.n251 B.n250 585
R869 B.n249 B.n148 585
R870 B.n248 B.n247 585
R871 B.n246 B.n149 585
R872 B.n245 B.n244 585
R873 B.n243 B.n150 585
R874 B.n242 B.n241 585
R875 B.n240 B.n151 585
R876 B.n239 B.n238 585
R877 B.n237 B.n152 585
R878 B.n236 B.n235 585
R879 B.n234 B.n153 585
R880 B.n233 B.n232 585
R881 B.n231 B.n154 585
R882 B.n230 B.n229 585
R883 B.n228 B.n155 585
R884 B.n227 B.n226 585
R885 B.n225 B.n156 585
R886 B.n224 B.n223 585
R887 B.n222 B.n157 585
R888 B.n221 B.n220 585
R889 B.n219 B.n158 585
R890 B.n218 B.n217 585
R891 B.n216 B.n159 585
R892 B.n215 B.n214 585
R893 B.n213 B.n160 585
R894 B.n212 B.n211 585
R895 B.n210 B.n161 585
R896 B.n385 B.n102 585
R897 B.n387 B.n386 585
R898 B.n388 B.n101 585
R899 B.n390 B.n389 585
R900 B.n391 B.n100 585
R901 B.n393 B.n392 585
R902 B.n394 B.n99 585
R903 B.n396 B.n395 585
R904 B.n397 B.n98 585
R905 B.n399 B.n398 585
R906 B.n400 B.n97 585
R907 B.n402 B.n401 585
R908 B.n403 B.n96 585
R909 B.n405 B.n404 585
R910 B.n406 B.n95 585
R911 B.n408 B.n407 585
R912 B.n409 B.n94 585
R913 B.n411 B.n410 585
R914 B.n412 B.n93 585
R915 B.n414 B.n413 585
R916 B.n415 B.n92 585
R917 B.n417 B.n416 585
R918 B.n418 B.n91 585
R919 B.n420 B.n419 585
R920 B.n421 B.n90 585
R921 B.n423 B.n422 585
R922 B.n424 B.n89 585
R923 B.n426 B.n425 585
R924 B.n427 B.n88 585
R925 B.n429 B.n428 585
R926 B.n430 B.n87 585
R927 B.n432 B.n431 585
R928 B.n433 B.n86 585
R929 B.n435 B.n434 585
R930 B.n436 B.n85 585
R931 B.n438 B.n437 585
R932 B.n439 B.n84 585
R933 B.n441 B.n440 585
R934 B.n442 B.n83 585
R935 B.n444 B.n443 585
R936 B.n445 B.n82 585
R937 B.n447 B.n446 585
R938 B.n448 B.n81 585
R939 B.n450 B.n449 585
R940 B.n451 B.n80 585
R941 B.n453 B.n452 585
R942 B.n454 B.n79 585
R943 B.n456 B.n455 585
R944 B.n457 B.n78 585
R945 B.n459 B.n458 585
R946 B.n460 B.n77 585
R947 B.n462 B.n461 585
R948 B.n634 B.n633 585
R949 B.n632 B.n15 585
R950 B.n631 B.n630 585
R951 B.n629 B.n16 585
R952 B.n628 B.n627 585
R953 B.n626 B.n17 585
R954 B.n625 B.n624 585
R955 B.n623 B.n18 585
R956 B.n622 B.n621 585
R957 B.n620 B.n19 585
R958 B.n619 B.n618 585
R959 B.n617 B.n20 585
R960 B.n616 B.n615 585
R961 B.n614 B.n21 585
R962 B.n613 B.n612 585
R963 B.n611 B.n22 585
R964 B.n610 B.n609 585
R965 B.n608 B.n23 585
R966 B.n607 B.n606 585
R967 B.n605 B.n24 585
R968 B.n604 B.n603 585
R969 B.n602 B.n25 585
R970 B.n601 B.n600 585
R971 B.n599 B.n26 585
R972 B.n598 B.n597 585
R973 B.n596 B.n27 585
R974 B.n595 B.n594 585
R975 B.n593 B.n28 585
R976 B.n592 B.n591 585
R977 B.n590 B.n29 585
R978 B.n589 B.n588 585
R979 B.n587 B.n30 585
R980 B.n586 B.n585 585
R981 B.n584 B.n31 585
R982 B.n583 B.n582 585
R983 B.n581 B.n32 585
R984 B.n580 B.n579 585
R985 B.n578 B.n33 585
R986 B.n577 B.n576 585
R987 B.n575 B.n34 585
R988 B.n574 B.n573 585
R989 B.n572 B.n35 585
R990 B.n571 B.n570 585
R991 B.n569 B.n36 585
R992 B.n568 B.n567 585
R993 B.n566 B.n37 585
R994 B.n565 B.n564 585
R995 B.n563 B.n38 585
R996 B.n562 B.n561 585
R997 B.n560 B.n39 585
R998 B.n559 B.n558 585
R999 B.n557 B.n40 585
R1000 B.n556 B.n555 585
R1001 B.n554 B.n41 585
R1002 B.n553 B.n552 585
R1003 B.n551 B.n45 585
R1004 B.n550 B.n549 585
R1005 B.n548 B.n46 585
R1006 B.n547 B.n546 585
R1007 B.n545 B.n47 585
R1008 B.n544 B.n543 585
R1009 B.n542 B.n48 585
R1010 B.n540 B.n539 585
R1011 B.n538 B.n51 585
R1012 B.n537 B.n536 585
R1013 B.n535 B.n52 585
R1014 B.n534 B.n533 585
R1015 B.n532 B.n53 585
R1016 B.n531 B.n530 585
R1017 B.n529 B.n54 585
R1018 B.n528 B.n527 585
R1019 B.n526 B.n55 585
R1020 B.n525 B.n524 585
R1021 B.n523 B.n56 585
R1022 B.n522 B.n521 585
R1023 B.n520 B.n57 585
R1024 B.n519 B.n518 585
R1025 B.n517 B.n58 585
R1026 B.n516 B.n515 585
R1027 B.n514 B.n59 585
R1028 B.n513 B.n512 585
R1029 B.n511 B.n60 585
R1030 B.n510 B.n509 585
R1031 B.n508 B.n61 585
R1032 B.n507 B.n506 585
R1033 B.n505 B.n62 585
R1034 B.n504 B.n503 585
R1035 B.n502 B.n63 585
R1036 B.n501 B.n500 585
R1037 B.n499 B.n64 585
R1038 B.n498 B.n497 585
R1039 B.n496 B.n65 585
R1040 B.n495 B.n494 585
R1041 B.n493 B.n66 585
R1042 B.n492 B.n491 585
R1043 B.n490 B.n67 585
R1044 B.n489 B.n488 585
R1045 B.n487 B.n68 585
R1046 B.n486 B.n485 585
R1047 B.n484 B.n69 585
R1048 B.n483 B.n482 585
R1049 B.n481 B.n70 585
R1050 B.n480 B.n479 585
R1051 B.n478 B.n71 585
R1052 B.n477 B.n476 585
R1053 B.n475 B.n72 585
R1054 B.n474 B.n473 585
R1055 B.n472 B.n73 585
R1056 B.n471 B.n470 585
R1057 B.n469 B.n74 585
R1058 B.n468 B.n467 585
R1059 B.n466 B.n75 585
R1060 B.n465 B.n464 585
R1061 B.n463 B.n76 585
R1062 B.n635 B.n14 585
R1063 B.n637 B.n636 585
R1064 B.n638 B.n13 585
R1065 B.n640 B.n639 585
R1066 B.n641 B.n12 585
R1067 B.n643 B.n642 585
R1068 B.n644 B.n11 585
R1069 B.n646 B.n645 585
R1070 B.n647 B.n10 585
R1071 B.n649 B.n648 585
R1072 B.n650 B.n9 585
R1073 B.n652 B.n651 585
R1074 B.n653 B.n8 585
R1075 B.n655 B.n654 585
R1076 B.n656 B.n7 585
R1077 B.n658 B.n657 585
R1078 B.n659 B.n6 585
R1079 B.n661 B.n660 585
R1080 B.n662 B.n5 585
R1081 B.n664 B.n663 585
R1082 B.n665 B.n4 585
R1083 B.n667 B.n666 585
R1084 B.n668 B.n3 585
R1085 B.n670 B.n669 585
R1086 B.n671 B.n0 585
R1087 B.n2 B.n1 585
R1088 B.n174 B.n173 585
R1089 B.n176 B.n175 585
R1090 B.n177 B.n172 585
R1091 B.n179 B.n178 585
R1092 B.n180 B.n171 585
R1093 B.n182 B.n181 585
R1094 B.n183 B.n170 585
R1095 B.n185 B.n184 585
R1096 B.n186 B.n169 585
R1097 B.n188 B.n187 585
R1098 B.n189 B.n168 585
R1099 B.n191 B.n190 585
R1100 B.n192 B.n167 585
R1101 B.n194 B.n193 585
R1102 B.n195 B.n166 585
R1103 B.n197 B.n196 585
R1104 B.n198 B.n165 585
R1105 B.n200 B.n199 585
R1106 B.n201 B.n164 585
R1107 B.n203 B.n202 585
R1108 B.n204 B.n163 585
R1109 B.n206 B.n205 585
R1110 B.n207 B.n162 585
R1111 B.n209 B.n208 585
R1112 B.n129 B.t7 497.084
R1113 B.n49 B.t11 497.084
R1114 B.n286 B.t4 497.084
R1115 B.n42 B.t2 497.084
R1116 B.n210 B.n209 478.086
R1117 B.n383 B.n102 478.086
R1118 B.n461 B.n76 478.086
R1119 B.n635 B.n634 478.086
R1120 B.n130 B.t8 439.678
R1121 B.n50 B.t10 439.678
R1122 B.n287 B.t5 439.678
R1123 B.n43 B.t1 439.678
R1124 B.n286 B.t3 350.584
R1125 B.n129 B.t6 350.584
R1126 B.n49 B.t9 350.584
R1127 B.n42 B.t0 350.584
R1128 B.n673 B.n672 256.663
R1129 B.n672 B.n671 235.042
R1130 B.n672 B.n2 235.042
R1131 B.n211 B.n210 163.367
R1132 B.n211 B.n160 163.367
R1133 B.n215 B.n160 163.367
R1134 B.n216 B.n215 163.367
R1135 B.n217 B.n216 163.367
R1136 B.n217 B.n158 163.367
R1137 B.n221 B.n158 163.367
R1138 B.n222 B.n221 163.367
R1139 B.n223 B.n222 163.367
R1140 B.n223 B.n156 163.367
R1141 B.n227 B.n156 163.367
R1142 B.n228 B.n227 163.367
R1143 B.n229 B.n228 163.367
R1144 B.n229 B.n154 163.367
R1145 B.n233 B.n154 163.367
R1146 B.n234 B.n233 163.367
R1147 B.n235 B.n234 163.367
R1148 B.n235 B.n152 163.367
R1149 B.n239 B.n152 163.367
R1150 B.n240 B.n239 163.367
R1151 B.n241 B.n240 163.367
R1152 B.n241 B.n150 163.367
R1153 B.n245 B.n150 163.367
R1154 B.n246 B.n245 163.367
R1155 B.n247 B.n246 163.367
R1156 B.n247 B.n148 163.367
R1157 B.n251 B.n148 163.367
R1158 B.n252 B.n251 163.367
R1159 B.n253 B.n252 163.367
R1160 B.n253 B.n146 163.367
R1161 B.n257 B.n146 163.367
R1162 B.n258 B.n257 163.367
R1163 B.n259 B.n258 163.367
R1164 B.n259 B.n144 163.367
R1165 B.n263 B.n144 163.367
R1166 B.n264 B.n263 163.367
R1167 B.n265 B.n264 163.367
R1168 B.n265 B.n142 163.367
R1169 B.n269 B.n142 163.367
R1170 B.n270 B.n269 163.367
R1171 B.n271 B.n270 163.367
R1172 B.n271 B.n140 163.367
R1173 B.n275 B.n140 163.367
R1174 B.n276 B.n275 163.367
R1175 B.n277 B.n276 163.367
R1176 B.n277 B.n138 163.367
R1177 B.n281 B.n138 163.367
R1178 B.n282 B.n281 163.367
R1179 B.n283 B.n282 163.367
R1180 B.n283 B.n136 163.367
R1181 B.n290 B.n136 163.367
R1182 B.n291 B.n290 163.367
R1183 B.n292 B.n291 163.367
R1184 B.n292 B.n134 163.367
R1185 B.n296 B.n134 163.367
R1186 B.n297 B.n296 163.367
R1187 B.n298 B.n297 163.367
R1188 B.n298 B.n132 163.367
R1189 B.n302 B.n132 163.367
R1190 B.n303 B.n302 163.367
R1191 B.n304 B.n303 163.367
R1192 B.n304 B.n128 163.367
R1193 B.n309 B.n128 163.367
R1194 B.n310 B.n309 163.367
R1195 B.n311 B.n310 163.367
R1196 B.n311 B.n126 163.367
R1197 B.n315 B.n126 163.367
R1198 B.n316 B.n315 163.367
R1199 B.n317 B.n316 163.367
R1200 B.n317 B.n124 163.367
R1201 B.n321 B.n124 163.367
R1202 B.n322 B.n321 163.367
R1203 B.n323 B.n322 163.367
R1204 B.n323 B.n122 163.367
R1205 B.n327 B.n122 163.367
R1206 B.n328 B.n327 163.367
R1207 B.n329 B.n328 163.367
R1208 B.n329 B.n120 163.367
R1209 B.n333 B.n120 163.367
R1210 B.n334 B.n333 163.367
R1211 B.n335 B.n334 163.367
R1212 B.n335 B.n118 163.367
R1213 B.n339 B.n118 163.367
R1214 B.n340 B.n339 163.367
R1215 B.n341 B.n340 163.367
R1216 B.n341 B.n116 163.367
R1217 B.n345 B.n116 163.367
R1218 B.n346 B.n345 163.367
R1219 B.n347 B.n346 163.367
R1220 B.n347 B.n114 163.367
R1221 B.n351 B.n114 163.367
R1222 B.n352 B.n351 163.367
R1223 B.n353 B.n352 163.367
R1224 B.n353 B.n112 163.367
R1225 B.n357 B.n112 163.367
R1226 B.n358 B.n357 163.367
R1227 B.n359 B.n358 163.367
R1228 B.n359 B.n110 163.367
R1229 B.n363 B.n110 163.367
R1230 B.n364 B.n363 163.367
R1231 B.n365 B.n364 163.367
R1232 B.n365 B.n108 163.367
R1233 B.n369 B.n108 163.367
R1234 B.n370 B.n369 163.367
R1235 B.n371 B.n370 163.367
R1236 B.n371 B.n106 163.367
R1237 B.n375 B.n106 163.367
R1238 B.n376 B.n375 163.367
R1239 B.n377 B.n376 163.367
R1240 B.n377 B.n104 163.367
R1241 B.n381 B.n104 163.367
R1242 B.n382 B.n381 163.367
R1243 B.n383 B.n382 163.367
R1244 B.n461 B.n460 163.367
R1245 B.n460 B.n459 163.367
R1246 B.n459 B.n78 163.367
R1247 B.n455 B.n78 163.367
R1248 B.n455 B.n454 163.367
R1249 B.n454 B.n453 163.367
R1250 B.n453 B.n80 163.367
R1251 B.n449 B.n80 163.367
R1252 B.n449 B.n448 163.367
R1253 B.n448 B.n447 163.367
R1254 B.n447 B.n82 163.367
R1255 B.n443 B.n82 163.367
R1256 B.n443 B.n442 163.367
R1257 B.n442 B.n441 163.367
R1258 B.n441 B.n84 163.367
R1259 B.n437 B.n84 163.367
R1260 B.n437 B.n436 163.367
R1261 B.n436 B.n435 163.367
R1262 B.n435 B.n86 163.367
R1263 B.n431 B.n86 163.367
R1264 B.n431 B.n430 163.367
R1265 B.n430 B.n429 163.367
R1266 B.n429 B.n88 163.367
R1267 B.n425 B.n88 163.367
R1268 B.n425 B.n424 163.367
R1269 B.n424 B.n423 163.367
R1270 B.n423 B.n90 163.367
R1271 B.n419 B.n90 163.367
R1272 B.n419 B.n418 163.367
R1273 B.n418 B.n417 163.367
R1274 B.n417 B.n92 163.367
R1275 B.n413 B.n92 163.367
R1276 B.n413 B.n412 163.367
R1277 B.n412 B.n411 163.367
R1278 B.n411 B.n94 163.367
R1279 B.n407 B.n94 163.367
R1280 B.n407 B.n406 163.367
R1281 B.n406 B.n405 163.367
R1282 B.n405 B.n96 163.367
R1283 B.n401 B.n96 163.367
R1284 B.n401 B.n400 163.367
R1285 B.n400 B.n399 163.367
R1286 B.n399 B.n98 163.367
R1287 B.n395 B.n98 163.367
R1288 B.n395 B.n394 163.367
R1289 B.n394 B.n393 163.367
R1290 B.n393 B.n100 163.367
R1291 B.n389 B.n100 163.367
R1292 B.n389 B.n388 163.367
R1293 B.n388 B.n387 163.367
R1294 B.n387 B.n102 163.367
R1295 B.n634 B.n15 163.367
R1296 B.n630 B.n15 163.367
R1297 B.n630 B.n629 163.367
R1298 B.n629 B.n628 163.367
R1299 B.n628 B.n17 163.367
R1300 B.n624 B.n17 163.367
R1301 B.n624 B.n623 163.367
R1302 B.n623 B.n622 163.367
R1303 B.n622 B.n19 163.367
R1304 B.n618 B.n19 163.367
R1305 B.n618 B.n617 163.367
R1306 B.n617 B.n616 163.367
R1307 B.n616 B.n21 163.367
R1308 B.n612 B.n21 163.367
R1309 B.n612 B.n611 163.367
R1310 B.n611 B.n610 163.367
R1311 B.n610 B.n23 163.367
R1312 B.n606 B.n23 163.367
R1313 B.n606 B.n605 163.367
R1314 B.n605 B.n604 163.367
R1315 B.n604 B.n25 163.367
R1316 B.n600 B.n25 163.367
R1317 B.n600 B.n599 163.367
R1318 B.n599 B.n598 163.367
R1319 B.n598 B.n27 163.367
R1320 B.n594 B.n27 163.367
R1321 B.n594 B.n593 163.367
R1322 B.n593 B.n592 163.367
R1323 B.n592 B.n29 163.367
R1324 B.n588 B.n29 163.367
R1325 B.n588 B.n587 163.367
R1326 B.n587 B.n586 163.367
R1327 B.n586 B.n31 163.367
R1328 B.n582 B.n31 163.367
R1329 B.n582 B.n581 163.367
R1330 B.n581 B.n580 163.367
R1331 B.n580 B.n33 163.367
R1332 B.n576 B.n33 163.367
R1333 B.n576 B.n575 163.367
R1334 B.n575 B.n574 163.367
R1335 B.n574 B.n35 163.367
R1336 B.n570 B.n35 163.367
R1337 B.n570 B.n569 163.367
R1338 B.n569 B.n568 163.367
R1339 B.n568 B.n37 163.367
R1340 B.n564 B.n37 163.367
R1341 B.n564 B.n563 163.367
R1342 B.n563 B.n562 163.367
R1343 B.n562 B.n39 163.367
R1344 B.n558 B.n39 163.367
R1345 B.n558 B.n557 163.367
R1346 B.n557 B.n556 163.367
R1347 B.n556 B.n41 163.367
R1348 B.n552 B.n41 163.367
R1349 B.n552 B.n551 163.367
R1350 B.n551 B.n550 163.367
R1351 B.n550 B.n46 163.367
R1352 B.n546 B.n46 163.367
R1353 B.n546 B.n545 163.367
R1354 B.n545 B.n544 163.367
R1355 B.n544 B.n48 163.367
R1356 B.n539 B.n48 163.367
R1357 B.n539 B.n538 163.367
R1358 B.n538 B.n537 163.367
R1359 B.n537 B.n52 163.367
R1360 B.n533 B.n52 163.367
R1361 B.n533 B.n532 163.367
R1362 B.n532 B.n531 163.367
R1363 B.n531 B.n54 163.367
R1364 B.n527 B.n54 163.367
R1365 B.n527 B.n526 163.367
R1366 B.n526 B.n525 163.367
R1367 B.n525 B.n56 163.367
R1368 B.n521 B.n56 163.367
R1369 B.n521 B.n520 163.367
R1370 B.n520 B.n519 163.367
R1371 B.n519 B.n58 163.367
R1372 B.n515 B.n58 163.367
R1373 B.n515 B.n514 163.367
R1374 B.n514 B.n513 163.367
R1375 B.n513 B.n60 163.367
R1376 B.n509 B.n60 163.367
R1377 B.n509 B.n508 163.367
R1378 B.n508 B.n507 163.367
R1379 B.n507 B.n62 163.367
R1380 B.n503 B.n62 163.367
R1381 B.n503 B.n502 163.367
R1382 B.n502 B.n501 163.367
R1383 B.n501 B.n64 163.367
R1384 B.n497 B.n64 163.367
R1385 B.n497 B.n496 163.367
R1386 B.n496 B.n495 163.367
R1387 B.n495 B.n66 163.367
R1388 B.n491 B.n66 163.367
R1389 B.n491 B.n490 163.367
R1390 B.n490 B.n489 163.367
R1391 B.n489 B.n68 163.367
R1392 B.n485 B.n68 163.367
R1393 B.n485 B.n484 163.367
R1394 B.n484 B.n483 163.367
R1395 B.n483 B.n70 163.367
R1396 B.n479 B.n70 163.367
R1397 B.n479 B.n478 163.367
R1398 B.n478 B.n477 163.367
R1399 B.n477 B.n72 163.367
R1400 B.n473 B.n72 163.367
R1401 B.n473 B.n472 163.367
R1402 B.n472 B.n471 163.367
R1403 B.n471 B.n74 163.367
R1404 B.n467 B.n74 163.367
R1405 B.n467 B.n466 163.367
R1406 B.n466 B.n465 163.367
R1407 B.n465 B.n76 163.367
R1408 B.n636 B.n635 163.367
R1409 B.n636 B.n13 163.367
R1410 B.n640 B.n13 163.367
R1411 B.n641 B.n640 163.367
R1412 B.n642 B.n641 163.367
R1413 B.n642 B.n11 163.367
R1414 B.n646 B.n11 163.367
R1415 B.n647 B.n646 163.367
R1416 B.n648 B.n647 163.367
R1417 B.n648 B.n9 163.367
R1418 B.n652 B.n9 163.367
R1419 B.n653 B.n652 163.367
R1420 B.n654 B.n653 163.367
R1421 B.n654 B.n7 163.367
R1422 B.n658 B.n7 163.367
R1423 B.n659 B.n658 163.367
R1424 B.n660 B.n659 163.367
R1425 B.n660 B.n5 163.367
R1426 B.n664 B.n5 163.367
R1427 B.n665 B.n664 163.367
R1428 B.n666 B.n665 163.367
R1429 B.n666 B.n3 163.367
R1430 B.n670 B.n3 163.367
R1431 B.n671 B.n670 163.367
R1432 B.n174 B.n2 163.367
R1433 B.n175 B.n174 163.367
R1434 B.n175 B.n172 163.367
R1435 B.n179 B.n172 163.367
R1436 B.n180 B.n179 163.367
R1437 B.n181 B.n180 163.367
R1438 B.n181 B.n170 163.367
R1439 B.n185 B.n170 163.367
R1440 B.n186 B.n185 163.367
R1441 B.n187 B.n186 163.367
R1442 B.n187 B.n168 163.367
R1443 B.n191 B.n168 163.367
R1444 B.n192 B.n191 163.367
R1445 B.n193 B.n192 163.367
R1446 B.n193 B.n166 163.367
R1447 B.n197 B.n166 163.367
R1448 B.n198 B.n197 163.367
R1449 B.n199 B.n198 163.367
R1450 B.n199 B.n164 163.367
R1451 B.n203 B.n164 163.367
R1452 B.n204 B.n203 163.367
R1453 B.n205 B.n204 163.367
R1454 B.n205 B.n162 163.367
R1455 B.n209 B.n162 163.367
R1456 B.n288 B.n287 59.5399
R1457 B.n306 B.n130 59.5399
R1458 B.n541 B.n50 59.5399
R1459 B.n44 B.n43 59.5399
R1460 B.n287 B.n286 57.4066
R1461 B.n130 B.n129 57.4066
R1462 B.n50 B.n49 57.4066
R1463 B.n43 B.n42 57.4066
R1464 B.n633 B.n14 31.0639
R1465 B.n463 B.n462 31.0639
R1466 B.n385 B.n384 31.0639
R1467 B.n208 B.n161 31.0639
R1468 B B.n673 18.0485
R1469 B.n637 B.n14 10.6151
R1470 B.n638 B.n637 10.6151
R1471 B.n639 B.n638 10.6151
R1472 B.n639 B.n12 10.6151
R1473 B.n643 B.n12 10.6151
R1474 B.n644 B.n643 10.6151
R1475 B.n645 B.n644 10.6151
R1476 B.n645 B.n10 10.6151
R1477 B.n649 B.n10 10.6151
R1478 B.n650 B.n649 10.6151
R1479 B.n651 B.n650 10.6151
R1480 B.n651 B.n8 10.6151
R1481 B.n655 B.n8 10.6151
R1482 B.n656 B.n655 10.6151
R1483 B.n657 B.n656 10.6151
R1484 B.n657 B.n6 10.6151
R1485 B.n661 B.n6 10.6151
R1486 B.n662 B.n661 10.6151
R1487 B.n663 B.n662 10.6151
R1488 B.n663 B.n4 10.6151
R1489 B.n667 B.n4 10.6151
R1490 B.n668 B.n667 10.6151
R1491 B.n669 B.n668 10.6151
R1492 B.n669 B.n0 10.6151
R1493 B.n633 B.n632 10.6151
R1494 B.n632 B.n631 10.6151
R1495 B.n631 B.n16 10.6151
R1496 B.n627 B.n16 10.6151
R1497 B.n627 B.n626 10.6151
R1498 B.n626 B.n625 10.6151
R1499 B.n625 B.n18 10.6151
R1500 B.n621 B.n18 10.6151
R1501 B.n621 B.n620 10.6151
R1502 B.n620 B.n619 10.6151
R1503 B.n619 B.n20 10.6151
R1504 B.n615 B.n20 10.6151
R1505 B.n615 B.n614 10.6151
R1506 B.n614 B.n613 10.6151
R1507 B.n613 B.n22 10.6151
R1508 B.n609 B.n22 10.6151
R1509 B.n609 B.n608 10.6151
R1510 B.n608 B.n607 10.6151
R1511 B.n607 B.n24 10.6151
R1512 B.n603 B.n24 10.6151
R1513 B.n603 B.n602 10.6151
R1514 B.n602 B.n601 10.6151
R1515 B.n601 B.n26 10.6151
R1516 B.n597 B.n26 10.6151
R1517 B.n597 B.n596 10.6151
R1518 B.n596 B.n595 10.6151
R1519 B.n595 B.n28 10.6151
R1520 B.n591 B.n28 10.6151
R1521 B.n591 B.n590 10.6151
R1522 B.n590 B.n589 10.6151
R1523 B.n589 B.n30 10.6151
R1524 B.n585 B.n30 10.6151
R1525 B.n585 B.n584 10.6151
R1526 B.n584 B.n583 10.6151
R1527 B.n583 B.n32 10.6151
R1528 B.n579 B.n32 10.6151
R1529 B.n579 B.n578 10.6151
R1530 B.n578 B.n577 10.6151
R1531 B.n577 B.n34 10.6151
R1532 B.n573 B.n34 10.6151
R1533 B.n573 B.n572 10.6151
R1534 B.n572 B.n571 10.6151
R1535 B.n571 B.n36 10.6151
R1536 B.n567 B.n36 10.6151
R1537 B.n567 B.n566 10.6151
R1538 B.n566 B.n565 10.6151
R1539 B.n565 B.n38 10.6151
R1540 B.n561 B.n38 10.6151
R1541 B.n561 B.n560 10.6151
R1542 B.n560 B.n559 10.6151
R1543 B.n559 B.n40 10.6151
R1544 B.n555 B.n554 10.6151
R1545 B.n554 B.n553 10.6151
R1546 B.n553 B.n45 10.6151
R1547 B.n549 B.n45 10.6151
R1548 B.n549 B.n548 10.6151
R1549 B.n548 B.n547 10.6151
R1550 B.n547 B.n47 10.6151
R1551 B.n543 B.n47 10.6151
R1552 B.n543 B.n542 10.6151
R1553 B.n540 B.n51 10.6151
R1554 B.n536 B.n51 10.6151
R1555 B.n536 B.n535 10.6151
R1556 B.n535 B.n534 10.6151
R1557 B.n534 B.n53 10.6151
R1558 B.n530 B.n53 10.6151
R1559 B.n530 B.n529 10.6151
R1560 B.n529 B.n528 10.6151
R1561 B.n528 B.n55 10.6151
R1562 B.n524 B.n55 10.6151
R1563 B.n524 B.n523 10.6151
R1564 B.n523 B.n522 10.6151
R1565 B.n522 B.n57 10.6151
R1566 B.n518 B.n57 10.6151
R1567 B.n518 B.n517 10.6151
R1568 B.n517 B.n516 10.6151
R1569 B.n516 B.n59 10.6151
R1570 B.n512 B.n59 10.6151
R1571 B.n512 B.n511 10.6151
R1572 B.n511 B.n510 10.6151
R1573 B.n510 B.n61 10.6151
R1574 B.n506 B.n61 10.6151
R1575 B.n506 B.n505 10.6151
R1576 B.n505 B.n504 10.6151
R1577 B.n504 B.n63 10.6151
R1578 B.n500 B.n63 10.6151
R1579 B.n500 B.n499 10.6151
R1580 B.n499 B.n498 10.6151
R1581 B.n498 B.n65 10.6151
R1582 B.n494 B.n65 10.6151
R1583 B.n494 B.n493 10.6151
R1584 B.n493 B.n492 10.6151
R1585 B.n492 B.n67 10.6151
R1586 B.n488 B.n67 10.6151
R1587 B.n488 B.n487 10.6151
R1588 B.n487 B.n486 10.6151
R1589 B.n486 B.n69 10.6151
R1590 B.n482 B.n69 10.6151
R1591 B.n482 B.n481 10.6151
R1592 B.n481 B.n480 10.6151
R1593 B.n480 B.n71 10.6151
R1594 B.n476 B.n71 10.6151
R1595 B.n476 B.n475 10.6151
R1596 B.n475 B.n474 10.6151
R1597 B.n474 B.n73 10.6151
R1598 B.n470 B.n73 10.6151
R1599 B.n470 B.n469 10.6151
R1600 B.n469 B.n468 10.6151
R1601 B.n468 B.n75 10.6151
R1602 B.n464 B.n75 10.6151
R1603 B.n464 B.n463 10.6151
R1604 B.n462 B.n77 10.6151
R1605 B.n458 B.n77 10.6151
R1606 B.n458 B.n457 10.6151
R1607 B.n457 B.n456 10.6151
R1608 B.n456 B.n79 10.6151
R1609 B.n452 B.n79 10.6151
R1610 B.n452 B.n451 10.6151
R1611 B.n451 B.n450 10.6151
R1612 B.n450 B.n81 10.6151
R1613 B.n446 B.n81 10.6151
R1614 B.n446 B.n445 10.6151
R1615 B.n445 B.n444 10.6151
R1616 B.n444 B.n83 10.6151
R1617 B.n440 B.n83 10.6151
R1618 B.n440 B.n439 10.6151
R1619 B.n439 B.n438 10.6151
R1620 B.n438 B.n85 10.6151
R1621 B.n434 B.n85 10.6151
R1622 B.n434 B.n433 10.6151
R1623 B.n433 B.n432 10.6151
R1624 B.n432 B.n87 10.6151
R1625 B.n428 B.n87 10.6151
R1626 B.n428 B.n427 10.6151
R1627 B.n427 B.n426 10.6151
R1628 B.n426 B.n89 10.6151
R1629 B.n422 B.n89 10.6151
R1630 B.n422 B.n421 10.6151
R1631 B.n421 B.n420 10.6151
R1632 B.n420 B.n91 10.6151
R1633 B.n416 B.n91 10.6151
R1634 B.n416 B.n415 10.6151
R1635 B.n415 B.n414 10.6151
R1636 B.n414 B.n93 10.6151
R1637 B.n410 B.n93 10.6151
R1638 B.n410 B.n409 10.6151
R1639 B.n409 B.n408 10.6151
R1640 B.n408 B.n95 10.6151
R1641 B.n404 B.n95 10.6151
R1642 B.n404 B.n403 10.6151
R1643 B.n403 B.n402 10.6151
R1644 B.n402 B.n97 10.6151
R1645 B.n398 B.n97 10.6151
R1646 B.n398 B.n397 10.6151
R1647 B.n397 B.n396 10.6151
R1648 B.n396 B.n99 10.6151
R1649 B.n392 B.n99 10.6151
R1650 B.n392 B.n391 10.6151
R1651 B.n391 B.n390 10.6151
R1652 B.n390 B.n101 10.6151
R1653 B.n386 B.n101 10.6151
R1654 B.n386 B.n385 10.6151
R1655 B.n173 B.n1 10.6151
R1656 B.n176 B.n173 10.6151
R1657 B.n177 B.n176 10.6151
R1658 B.n178 B.n177 10.6151
R1659 B.n178 B.n171 10.6151
R1660 B.n182 B.n171 10.6151
R1661 B.n183 B.n182 10.6151
R1662 B.n184 B.n183 10.6151
R1663 B.n184 B.n169 10.6151
R1664 B.n188 B.n169 10.6151
R1665 B.n189 B.n188 10.6151
R1666 B.n190 B.n189 10.6151
R1667 B.n190 B.n167 10.6151
R1668 B.n194 B.n167 10.6151
R1669 B.n195 B.n194 10.6151
R1670 B.n196 B.n195 10.6151
R1671 B.n196 B.n165 10.6151
R1672 B.n200 B.n165 10.6151
R1673 B.n201 B.n200 10.6151
R1674 B.n202 B.n201 10.6151
R1675 B.n202 B.n163 10.6151
R1676 B.n206 B.n163 10.6151
R1677 B.n207 B.n206 10.6151
R1678 B.n208 B.n207 10.6151
R1679 B.n212 B.n161 10.6151
R1680 B.n213 B.n212 10.6151
R1681 B.n214 B.n213 10.6151
R1682 B.n214 B.n159 10.6151
R1683 B.n218 B.n159 10.6151
R1684 B.n219 B.n218 10.6151
R1685 B.n220 B.n219 10.6151
R1686 B.n220 B.n157 10.6151
R1687 B.n224 B.n157 10.6151
R1688 B.n225 B.n224 10.6151
R1689 B.n226 B.n225 10.6151
R1690 B.n226 B.n155 10.6151
R1691 B.n230 B.n155 10.6151
R1692 B.n231 B.n230 10.6151
R1693 B.n232 B.n231 10.6151
R1694 B.n232 B.n153 10.6151
R1695 B.n236 B.n153 10.6151
R1696 B.n237 B.n236 10.6151
R1697 B.n238 B.n237 10.6151
R1698 B.n238 B.n151 10.6151
R1699 B.n242 B.n151 10.6151
R1700 B.n243 B.n242 10.6151
R1701 B.n244 B.n243 10.6151
R1702 B.n244 B.n149 10.6151
R1703 B.n248 B.n149 10.6151
R1704 B.n249 B.n248 10.6151
R1705 B.n250 B.n249 10.6151
R1706 B.n250 B.n147 10.6151
R1707 B.n254 B.n147 10.6151
R1708 B.n255 B.n254 10.6151
R1709 B.n256 B.n255 10.6151
R1710 B.n256 B.n145 10.6151
R1711 B.n260 B.n145 10.6151
R1712 B.n261 B.n260 10.6151
R1713 B.n262 B.n261 10.6151
R1714 B.n262 B.n143 10.6151
R1715 B.n266 B.n143 10.6151
R1716 B.n267 B.n266 10.6151
R1717 B.n268 B.n267 10.6151
R1718 B.n268 B.n141 10.6151
R1719 B.n272 B.n141 10.6151
R1720 B.n273 B.n272 10.6151
R1721 B.n274 B.n273 10.6151
R1722 B.n274 B.n139 10.6151
R1723 B.n278 B.n139 10.6151
R1724 B.n279 B.n278 10.6151
R1725 B.n280 B.n279 10.6151
R1726 B.n280 B.n137 10.6151
R1727 B.n284 B.n137 10.6151
R1728 B.n285 B.n284 10.6151
R1729 B.n289 B.n285 10.6151
R1730 B.n293 B.n135 10.6151
R1731 B.n294 B.n293 10.6151
R1732 B.n295 B.n294 10.6151
R1733 B.n295 B.n133 10.6151
R1734 B.n299 B.n133 10.6151
R1735 B.n300 B.n299 10.6151
R1736 B.n301 B.n300 10.6151
R1737 B.n301 B.n131 10.6151
R1738 B.n305 B.n131 10.6151
R1739 B.n308 B.n307 10.6151
R1740 B.n308 B.n127 10.6151
R1741 B.n312 B.n127 10.6151
R1742 B.n313 B.n312 10.6151
R1743 B.n314 B.n313 10.6151
R1744 B.n314 B.n125 10.6151
R1745 B.n318 B.n125 10.6151
R1746 B.n319 B.n318 10.6151
R1747 B.n320 B.n319 10.6151
R1748 B.n320 B.n123 10.6151
R1749 B.n324 B.n123 10.6151
R1750 B.n325 B.n324 10.6151
R1751 B.n326 B.n325 10.6151
R1752 B.n326 B.n121 10.6151
R1753 B.n330 B.n121 10.6151
R1754 B.n331 B.n330 10.6151
R1755 B.n332 B.n331 10.6151
R1756 B.n332 B.n119 10.6151
R1757 B.n336 B.n119 10.6151
R1758 B.n337 B.n336 10.6151
R1759 B.n338 B.n337 10.6151
R1760 B.n338 B.n117 10.6151
R1761 B.n342 B.n117 10.6151
R1762 B.n343 B.n342 10.6151
R1763 B.n344 B.n343 10.6151
R1764 B.n344 B.n115 10.6151
R1765 B.n348 B.n115 10.6151
R1766 B.n349 B.n348 10.6151
R1767 B.n350 B.n349 10.6151
R1768 B.n350 B.n113 10.6151
R1769 B.n354 B.n113 10.6151
R1770 B.n355 B.n354 10.6151
R1771 B.n356 B.n355 10.6151
R1772 B.n356 B.n111 10.6151
R1773 B.n360 B.n111 10.6151
R1774 B.n361 B.n360 10.6151
R1775 B.n362 B.n361 10.6151
R1776 B.n362 B.n109 10.6151
R1777 B.n366 B.n109 10.6151
R1778 B.n367 B.n366 10.6151
R1779 B.n368 B.n367 10.6151
R1780 B.n368 B.n107 10.6151
R1781 B.n372 B.n107 10.6151
R1782 B.n373 B.n372 10.6151
R1783 B.n374 B.n373 10.6151
R1784 B.n374 B.n105 10.6151
R1785 B.n378 B.n105 10.6151
R1786 B.n379 B.n378 10.6151
R1787 B.n380 B.n379 10.6151
R1788 B.n380 B.n103 10.6151
R1789 B.n384 B.n103 10.6151
R1790 B.n44 B.n40 9.36635
R1791 B.n541 B.n540 9.36635
R1792 B.n289 B.n288 9.36635
R1793 B.n307 B.n306 9.36635
R1794 B.n673 B.n0 8.11757
R1795 B.n673 B.n1 8.11757
R1796 B.n555 B.n44 1.24928
R1797 B.n542 B.n541 1.24928
R1798 B.n288 B.n135 1.24928
R1799 B.n306 B.n305 1.24928
R1800 VN VN.t0 231.017
R1801 VN VN.t1 184.019
R1802 VDD2.n165 VDD2.n85 756.745
R1803 VDD2.n80 VDD2.n0 756.745
R1804 VDD2.n166 VDD2.n165 585
R1805 VDD2.n164 VDD2.n163 585
R1806 VDD2.n89 VDD2.n88 585
R1807 VDD2.n93 VDD2.n91 585
R1808 VDD2.n158 VDD2.n157 585
R1809 VDD2.n156 VDD2.n155 585
R1810 VDD2.n95 VDD2.n94 585
R1811 VDD2.n150 VDD2.n149 585
R1812 VDD2.n148 VDD2.n147 585
R1813 VDD2.n99 VDD2.n98 585
R1814 VDD2.n142 VDD2.n141 585
R1815 VDD2.n140 VDD2.n139 585
R1816 VDD2.n103 VDD2.n102 585
R1817 VDD2.n134 VDD2.n133 585
R1818 VDD2.n132 VDD2.n131 585
R1819 VDD2.n107 VDD2.n106 585
R1820 VDD2.n126 VDD2.n125 585
R1821 VDD2.n124 VDD2.n123 585
R1822 VDD2.n111 VDD2.n110 585
R1823 VDD2.n118 VDD2.n117 585
R1824 VDD2.n116 VDD2.n115 585
R1825 VDD2.n29 VDD2.n28 585
R1826 VDD2.n31 VDD2.n30 585
R1827 VDD2.n24 VDD2.n23 585
R1828 VDD2.n37 VDD2.n36 585
R1829 VDD2.n39 VDD2.n38 585
R1830 VDD2.n20 VDD2.n19 585
R1831 VDD2.n45 VDD2.n44 585
R1832 VDD2.n47 VDD2.n46 585
R1833 VDD2.n16 VDD2.n15 585
R1834 VDD2.n53 VDD2.n52 585
R1835 VDD2.n55 VDD2.n54 585
R1836 VDD2.n12 VDD2.n11 585
R1837 VDD2.n61 VDD2.n60 585
R1838 VDD2.n63 VDD2.n62 585
R1839 VDD2.n8 VDD2.n7 585
R1840 VDD2.n70 VDD2.n69 585
R1841 VDD2.n71 VDD2.n6 585
R1842 VDD2.n73 VDD2.n72 585
R1843 VDD2.n4 VDD2.n3 585
R1844 VDD2.n79 VDD2.n78 585
R1845 VDD2.n81 VDD2.n80 585
R1846 VDD2.n114 VDD2.t1 327.466
R1847 VDD2.n27 VDD2.t0 327.466
R1848 VDD2.n165 VDD2.n164 171.744
R1849 VDD2.n164 VDD2.n88 171.744
R1850 VDD2.n93 VDD2.n88 171.744
R1851 VDD2.n157 VDD2.n93 171.744
R1852 VDD2.n157 VDD2.n156 171.744
R1853 VDD2.n156 VDD2.n94 171.744
R1854 VDD2.n149 VDD2.n94 171.744
R1855 VDD2.n149 VDD2.n148 171.744
R1856 VDD2.n148 VDD2.n98 171.744
R1857 VDD2.n141 VDD2.n98 171.744
R1858 VDD2.n141 VDD2.n140 171.744
R1859 VDD2.n140 VDD2.n102 171.744
R1860 VDD2.n133 VDD2.n102 171.744
R1861 VDD2.n133 VDD2.n132 171.744
R1862 VDD2.n132 VDD2.n106 171.744
R1863 VDD2.n125 VDD2.n106 171.744
R1864 VDD2.n125 VDD2.n124 171.744
R1865 VDD2.n124 VDD2.n110 171.744
R1866 VDD2.n117 VDD2.n110 171.744
R1867 VDD2.n117 VDD2.n116 171.744
R1868 VDD2.n30 VDD2.n29 171.744
R1869 VDD2.n30 VDD2.n23 171.744
R1870 VDD2.n37 VDD2.n23 171.744
R1871 VDD2.n38 VDD2.n37 171.744
R1872 VDD2.n38 VDD2.n19 171.744
R1873 VDD2.n45 VDD2.n19 171.744
R1874 VDD2.n46 VDD2.n45 171.744
R1875 VDD2.n46 VDD2.n15 171.744
R1876 VDD2.n53 VDD2.n15 171.744
R1877 VDD2.n54 VDD2.n53 171.744
R1878 VDD2.n54 VDD2.n11 171.744
R1879 VDD2.n61 VDD2.n11 171.744
R1880 VDD2.n62 VDD2.n61 171.744
R1881 VDD2.n62 VDD2.n7 171.744
R1882 VDD2.n70 VDD2.n7 171.744
R1883 VDD2.n71 VDD2.n70 171.744
R1884 VDD2.n72 VDD2.n71 171.744
R1885 VDD2.n72 VDD2.n3 171.744
R1886 VDD2.n79 VDD2.n3 171.744
R1887 VDD2.n80 VDD2.n79 171.744
R1888 VDD2.n170 VDD2.n84 94.7171
R1889 VDD2.n116 VDD2.t1 85.8723
R1890 VDD2.n29 VDD2.t0 85.8723
R1891 VDD2.n170 VDD2.n169 52.549
R1892 VDD2.n115 VDD2.n114 16.3895
R1893 VDD2.n28 VDD2.n27 16.3895
R1894 VDD2.n91 VDD2.n89 13.1884
R1895 VDD2.n73 VDD2.n4 13.1884
R1896 VDD2.n163 VDD2.n162 12.8005
R1897 VDD2.n159 VDD2.n158 12.8005
R1898 VDD2.n118 VDD2.n113 12.8005
R1899 VDD2.n31 VDD2.n26 12.8005
R1900 VDD2.n74 VDD2.n6 12.8005
R1901 VDD2.n78 VDD2.n77 12.8005
R1902 VDD2.n166 VDD2.n87 12.0247
R1903 VDD2.n155 VDD2.n92 12.0247
R1904 VDD2.n119 VDD2.n111 12.0247
R1905 VDD2.n32 VDD2.n24 12.0247
R1906 VDD2.n69 VDD2.n68 12.0247
R1907 VDD2.n81 VDD2.n2 12.0247
R1908 VDD2.n167 VDD2.n85 11.249
R1909 VDD2.n154 VDD2.n95 11.249
R1910 VDD2.n123 VDD2.n122 11.249
R1911 VDD2.n36 VDD2.n35 11.249
R1912 VDD2.n67 VDD2.n8 11.249
R1913 VDD2.n82 VDD2.n0 11.249
R1914 VDD2.n151 VDD2.n150 10.4732
R1915 VDD2.n126 VDD2.n109 10.4732
R1916 VDD2.n39 VDD2.n22 10.4732
R1917 VDD2.n64 VDD2.n63 10.4732
R1918 VDD2.n147 VDD2.n97 9.69747
R1919 VDD2.n127 VDD2.n107 9.69747
R1920 VDD2.n40 VDD2.n20 9.69747
R1921 VDD2.n60 VDD2.n10 9.69747
R1922 VDD2.n169 VDD2.n168 9.45567
R1923 VDD2.n84 VDD2.n83 9.45567
R1924 VDD2.n101 VDD2.n100 9.3005
R1925 VDD2.n144 VDD2.n143 9.3005
R1926 VDD2.n146 VDD2.n145 9.3005
R1927 VDD2.n97 VDD2.n96 9.3005
R1928 VDD2.n152 VDD2.n151 9.3005
R1929 VDD2.n154 VDD2.n153 9.3005
R1930 VDD2.n92 VDD2.n90 9.3005
R1931 VDD2.n160 VDD2.n159 9.3005
R1932 VDD2.n168 VDD2.n167 9.3005
R1933 VDD2.n87 VDD2.n86 9.3005
R1934 VDD2.n162 VDD2.n161 9.3005
R1935 VDD2.n138 VDD2.n137 9.3005
R1936 VDD2.n136 VDD2.n135 9.3005
R1937 VDD2.n105 VDD2.n104 9.3005
R1938 VDD2.n130 VDD2.n129 9.3005
R1939 VDD2.n128 VDD2.n127 9.3005
R1940 VDD2.n109 VDD2.n108 9.3005
R1941 VDD2.n122 VDD2.n121 9.3005
R1942 VDD2.n120 VDD2.n119 9.3005
R1943 VDD2.n113 VDD2.n112 9.3005
R1944 VDD2.n83 VDD2.n82 9.3005
R1945 VDD2.n2 VDD2.n1 9.3005
R1946 VDD2.n77 VDD2.n76 9.3005
R1947 VDD2.n49 VDD2.n48 9.3005
R1948 VDD2.n18 VDD2.n17 9.3005
R1949 VDD2.n43 VDD2.n42 9.3005
R1950 VDD2.n41 VDD2.n40 9.3005
R1951 VDD2.n22 VDD2.n21 9.3005
R1952 VDD2.n35 VDD2.n34 9.3005
R1953 VDD2.n33 VDD2.n32 9.3005
R1954 VDD2.n26 VDD2.n25 9.3005
R1955 VDD2.n51 VDD2.n50 9.3005
R1956 VDD2.n14 VDD2.n13 9.3005
R1957 VDD2.n57 VDD2.n56 9.3005
R1958 VDD2.n59 VDD2.n58 9.3005
R1959 VDD2.n10 VDD2.n9 9.3005
R1960 VDD2.n65 VDD2.n64 9.3005
R1961 VDD2.n67 VDD2.n66 9.3005
R1962 VDD2.n68 VDD2.n5 9.3005
R1963 VDD2.n75 VDD2.n74 9.3005
R1964 VDD2.n146 VDD2.n99 8.92171
R1965 VDD2.n131 VDD2.n130 8.92171
R1966 VDD2.n44 VDD2.n43 8.92171
R1967 VDD2.n59 VDD2.n12 8.92171
R1968 VDD2.n143 VDD2.n142 8.14595
R1969 VDD2.n134 VDD2.n105 8.14595
R1970 VDD2.n47 VDD2.n18 8.14595
R1971 VDD2.n56 VDD2.n55 8.14595
R1972 VDD2.n139 VDD2.n101 7.3702
R1973 VDD2.n135 VDD2.n103 7.3702
R1974 VDD2.n48 VDD2.n16 7.3702
R1975 VDD2.n52 VDD2.n14 7.3702
R1976 VDD2.n139 VDD2.n138 6.59444
R1977 VDD2.n138 VDD2.n103 6.59444
R1978 VDD2.n51 VDD2.n16 6.59444
R1979 VDD2.n52 VDD2.n51 6.59444
R1980 VDD2.n142 VDD2.n101 5.81868
R1981 VDD2.n135 VDD2.n134 5.81868
R1982 VDD2.n48 VDD2.n47 5.81868
R1983 VDD2.n55 VDD2.n14 5.81868
R1984 VDD2.n143 VDD2.n99 5.04292
R1985 VDD2.n131 VDD2.n105 5.04292
R1986 VDD2.n44 VDD2.n18 5.04292
R1987 VDD2.n56 VDD2.n12 5.04292
R1988 VDD2.n147 VDD2.n146 4.26717
R1989 VDD2.n130 VDD2.n107 4.26717
R1990 VDD2.n43 VDD2.n20 4.26717
R1991 VDD2.n60 VDD2.n59 4.26717
R1992 VDD2.n114 VDD2.n112 3.70982
R1993 VDD2.n27 VDD2.n25 3.70982
R1994 VDD2.n150 VDD2.n97 3.49141
R1995 VDD2.n127 VDD2.n126 3.49141
R1996 VDD2.n40 VDD2.n39 3.49141
R1997 VDD2.n63 VDD2.n10 3.49141
R1998 VDD2.n169 VDD2.n85 2.71565
R1999 VDD2.n151 VDD2.n95 2.71565
R2000 VDD2.n123 VDD2.n109 2.71565
R2001 VDD2.n36 VDD2.n22 2.71565
R2002 VDD2.n64 VDD2.n8 2.71565
R2003 VDD2.n84 VDD2.n0 2.71565
R2004 VDD2.n167 VDD2.n166 1.93989
R2005 VDD2.n155 VDD2.n154 1.93989
R2006 VDD2.n122 VDD2.n111 1.93989
R2007 VDD2.n35 VDD2.n24 1.93989
R2008 VDD2.n69 VDD2.n67 1.93989
R2009 VDD2.n82 VDD2.n81 1.93989
R2010 VDD2.n163 VDD2.n87 1.16414
R2011 VDD2.n158 VDD2.n92 1.16414
R2012 VDD2.n119 VDD2.n118 1.16414
R2013 VDD2.n32 VDD2.n31 1.16414
R2014 VDD2.n68 VDD2.n6 1.16414
R2015 VDD2.n78 VDD2.n2 1.16414
R2016 VDD2 VDD2.n170 0.696621
R2017 VDD2.n162 VDD2.n89 0.388379
R2018 VDD2.n159 VDD2.n91 0.388379
R2019 VDD2.n115 VDD2.n113 0.388379
R2020 VDD2.n28 VDD2.n26 0.388379
R2021 VDD2.n74 VDD2.n73 0.388379
R2022 VDD2.n77 VDD2.n4 0.388379
R2023 VDD2.n168 VDD2.n86 0.155672
R2024 VDD2.n161 VDD2.n86 0.155672
R2025 VDD2.n161 VDD2.n160 0.155672
R2026 VDD2.n160 VDD2.n90 0.155672
R2027 VDD2.n153 VDD2.n90 0.155672
R2028 VDD2.n153 VDD2.n152 0.155672
R2029 VDD2.n152 VDD2.n96 0.155672
R2030 VDD2.n145 VDD2.n96 0.155672
R2031 VDD2.n145 VDD2.n144 0.155672
R2032 VDD2.n144 VDD2.n100 0.155672
R2033 VDD2.n137 VDD2.n100 0.155672
R2034 VDD2.n137 VDD2.n136 0.155672
R2035 VDD2.n136 VDD2.n104 0.155672
R2036 VDD2.n129 VDD2.n104 0.155672
R2037 VDD2.n129 VDD2.n128 0.155672
R2038 VDD2.n128 VDD2.n108 0.155672
R2039 VDD2.n121 VDD2.n108 0.155672
R2040 VDD2.n121 VDD2.n120 0.155672
R2041 VDD2.n120 VDD2.n112 0.155672
R2042 VDD2.n33 VDD2.n25 0.155672
R2043 VDD2.n34 VDD2.n33 0.155672
R2044 VDD2.n34 VDD2.n21 0.155672
R2045 VDD2.n41 VDD2.n21 0.155672
R2046 VDD2.n42 VDD2.n41 0.155672
R2047 VDD2.n42 VDD2.n17 0.155672
R2048 VDD2.n49 VDD2.n17 0.155672
R2049 VDD2.n50 VDD2.n49 0.155672
R2050 VDD2.n50 VDD2.n13 0.155672
R2051 VDD2.n57 VDD2.n13 0.155672
R2052 VDD2.n58 VDD2.n57 0.155672
R2053 VDD2.n58 VDD2.n9 0.155672
R2054 VDD2.n65 VDD2.n9 0.155672
R2055 VDD2.n66 VDD2.n65 0.155672
R2056 VDD2.n66 VDD2.n5 0.155672
R2057 VDD2.n75 VDD2.n5 0.155672
R2058 VDD2.n76 VDD2.n75 0.155672
R2059 VDD2.n76 VDD2.n1 0.155672
R2060 VDD2.n83 VDD2.n1 0.155672
C0 B VN 1.09664f
C1 VN w_n2154_n4078# 3.05948f
C2 VN VP 6.13145f
C3 VTAIL B 4.46651f
C4 VTAIL w_n2154_n4078# 3.24504f
C5 VTAIL VP 3.05785f
C6 B w_n2154_n4078# 9.83662f
C7 B VP 1.54796f
C8 VP w_n2154_n4078# 3.33392f
C9 VN VDD2 3.5352f
C10 VN VDD1 0.148136f
C11 VTAIL VDD2 6.05729f
C12 VTAIL VDD1 6.00726f
C13 B VDD2 2.02065f
C14 B VDD1 1.9903f
C15 VDD2 w_n2154_n4078# 2.05709f
C16 VP VDD2 0.334606f
C17 w_n2154_n4078# VDD1 2.03084f
C18 VP VDD1 3.71854f
C19 VDD2 VDD1 0.678631f
C20 VTAIL VN 3.04351f
C21 VDD2 VSUBS 1.055002f
C22 VDD1 VSUBS 4.68326f
C23 VTAIL VSUBS 1.144152f
C24 VN VSUBS 8.61801f
C25 VP VSUBS 1.827816f
C26 B VSUBS 4.231579f
C27 w_n2154_n4078# VSUBS 0.107657p
C28 VDD2.n0 VSUBS 0.031696f
C29 VDD2.n1 VSUBS 0.028624f
C30 VDD2.n2 VSUBS 0.015381f
C31 VDD2.n3 VSUBS 0.036356f
C32 VDD2.n4 VSUBS 0.015834f
C33 VDD2.n5 VSUBS 0.028624f
C34 VDD2.n6 VSUBS 0.016286f
C35 VDD2.n7 VSUBS 0.036356f
C36 VDD2.n8 VSUBS 0.016286f
C37 VDD2.n9 VSUBS 0.028624f
C38 VDD2.n10 VSUBS 0.015381f
C39 VDD2.n11 VSUBS 0.036356f
C40 VDD2.n12 VSUBS 0.016286f
C41 VDD2.n13 VSUBS 0.028624f
C42 VDD2.n14 VSUBS 0.015381f
C43 VDD2.n15 VSUBS 0.036356f
C44 VDD2.n16 VSUBS 0.016286f
C45 VDD2.n17 VSUBS 0.028624f
C46 VDD2.n18 VSUBS 0.015381f
C47 VDD2.n19 VSUBS 0.036356f
C48 VDD2.n20 VSUBS 0.016286f
C49 VDD2.n21 VSUBS 0.028624f
C50 VDD2.n22 VSUBS 0.015381f
C51 VDD2.n23 VSUBS 0.036356f
C52 VDD2.n24 VSUBS 0.016286f
C53 VDD2.n25 VSUBS 1.89917f
C54 VDD2.n26 VSUBS 0.015381f
C55 VDD2.t0 VSUBS 0.07787f
C56 VDD2.n27 VSUBS 0.206419f
C57 VDD2.n28 VSUBS 0.023128f
C58 VDD2.n29 VSUBS 0.027267f
C59 VDD2.n30 VSUBS 0.036356f
C60 VDD2.n31 VSUBS 0.016286f
C61 VDD2.n32 VSUBS 0.015381f
C62 VDD2.n33 VSUBS 0.028624f
C63 VDD2.n34 VSUBS 0.028624f
C64 VDD2.n35 VSUBS 0.015381f
C65 VDD2.n36 VSUBS 0.016286f
C66 VDD2.n37 VSUBS 0.036356f
C67 VDD2.n38 VSUBS 0.036356f
C68 VDD2.n39 VSUBS 0.016286f
C69 VDD2.n40 VSUBS 0.015381f
C70 VDD2.n41 VSUBS 0.028624f
C71 VDD2.n42 VSUBS 0.028624f
C72 VDD2.n43 VSUBS 0.015381f
C73 VDD2.n44 VSUBS 0.016286f
C74 VDD2.n45 VSUBS 0.036356f
C75 VDD2.n46 VSUBS 0.036356f
C76 VDD2.n47 VSUBS 0.016286f
C77 VDD2.n48 VSUBS 0.015381f
C78 VDD2.n49 VSUBS 0.028624f
C79 VDD2.n50 VSUBS 0.028624f
C80 VDD2.n51 VSUBS 0.015381f
C81 VDD2.n52 VSUBS 0.016286f
C82 VDD2.n53 VSUBS 0.036356f
C83 VDD2.n54 VSUBS 0.036356f
C84 VDD2.n55 VSUBS 0.016286f
C85 VDD2.n56 VSUBS 0.015381f
C86 VDD2.n57 VSUBS 0.028624f
C87 VDD2.n58 VSUBS 0.028624f
C88 VDD2.n59 VSUBS 0.015381f
C89 VDD2.n60 VSUBS 0.016286f
C90 VDD2.n61 VSUBS 0.036356f
C91 VDD2.n62 VSUBS 0.036356f
C92 VDD2.n63 VSUBS 0.016286f
C93 VDD2.n64 VSUBS 0.015381f
C94 VDD2.n65 VSUBS 0.028624f
C95 VDD2.n66 VSUBS 0.028624f
C96 VDD2.n67 VSUBS 0.015381f
C97 VDD2.n68 VSUBS 0.015381f
C98 VDD2.n69 VSUBS 0.016286f
C99 VDD2.n70 VSUBS 0.036356f
C100 VDD2.n71 VSUBS 0.036356f
C101 VDD2.n72 VSUBS 0.036356f
C102 VDD2.n73 VSUBS 0.015834f
C103 VDD2.n74 VSUBS 0.015381f
C104 VDD2.n75 VSUBS 0.028624f
C105 VDD2.n76 VSUBS 0.028624f
C106 VDD2.n77 VSUBS 0.015381f
C107 VDD2.n78 VSUBS 0.016286f
C108 VDD2.n79 VSUBS 0.036356f
C109 VDD2.n80 VSUBS 0.088846f
C110 VDD2.n81 VSUBS 0.016286f
C111 VDD2.n82 VSUBS 0.015381f
C112 VDD2.n83 VSUBS 0.073593f
C113 VDD2.n84 VSUBS 0.959327f
C114 VDD2.n85 VSUBS 0.031696f
C115 VDD2.n86 VSUBS 0.028624f
C116 VDD2.n87 VSUBS 0.015381f
C117 VDD2.n88 VSUBS 0.036356f
C118 VDD2.n89 VSUBS 0.015834f
C119 VDD2.n90 VSUBS 0.028624f
C120 VDD2.n91 VSUBS 0.015834f
C121 VDD2.n92 VSUBS 0.015381f
C122 VDD2.n93 VSUBS 0.036356f
C123 VDD2.n94 VSUBS 0.036356f
C124 VDD2.n95 VSUBS 0.016286f
C125 VDD2.n96 VSUBS 0.028624f
C126 VDD2.n97 VSUBS 0.015381f
C127 VDD2.n98 VSUBS 0.036356f
C128 VDD2.n99 VSUBS 0.016286f
C129 VDD2.n100 VSUBS 0.028624f
C130 VDD2.n101 VSUBS 0.015381f
C131 VDD2.n102 VSUBS 0.036356f
C132 VDD2.n103 VSUBS 0.016286f
C133 VDD2.n104 VSUBS 0.028624f
C134 VDD2.n105 VSUBS 0.015381f
C135 VDD2.n106 VSUBS 0.036356f
C136 VDD2.n107 VSUBS 0.016286f
C137 VDD2.n108 VSUBS 0.028624f
C138 VDD2.n109 VSUBS 0.015381f
C139 VDD2.n110 VSUBS 0.036356f
C140 VDD2.n111 VSUBS 0.016286f
C141 VDD2.n112 VSUBS 1.89918f
C142 VDD2.n113 VSUBS 0.015381f
C143 VDD2.t1 VSUBS 0.07787f
C144 VDD2.n114 VSUBS 0.206419f
C145 VDD2.n115 VSUBS 0.023128f
C146 VDD2.n116 VSUBS 0.027267f
C147 VDD2.n117 VSUBS 0.036356f
C148 VDD2.n118 VSUBS 0.016286f
C149 VDD2.n119 VSUBS 0.015381f
C150 VDD2.n120 VSUBS 0.028624f
C151 VDD2.n121 VSUBS 0.028624f
C152 VDD2.n122 VSUBS 0.015381f
C153 VDD2.n123 VSUBS 0.016286f
C154 VDD2.n124 VSUBS 0.036356f
C155 VDD2.n125 VSUBS 0.036356f
C156 VDD2.n126 VSUBS 0.016286f
C157 VDD2.n127 VSUBS 0.015381f
C158 VDD2.n128 VSUBS 0.028624f
C159 VDD2.n129 VSUBS 0.028624f
C160 VDD2.n130 VSUBS 0.015381f
C161 VDD2.n131 VSUBS 0.016286f
C162 VDD2.n132 VSUBS 0.036356f
C163 VDD2.n133 VSUBS 0.036356f
C164 VDD2.n134 VSUBS 0.016286f
C165 VDD2.n135 VSUBS 0.015381f
C166 VDD2.n136 VSUBS 0.028624f
C167 VDD2.n137 VSUBS 0.028624f
C168 VDD2.n138 VSUBS 0.015381f
C169 VDD2.n139 VSUBS 0.016286f
C170 VDD2.n140 VSUBS 0.036356f
C171 VDD2.n141 VSUBS 0.036356f
C172 VDD2.n142 VSUBS 0.016286f
C173 VDD2.n143 VSUBS 0.015381f
C174 VDD2.n144 VSUBS 0.028624f
C175 VDD2.n145 VSUBS 0.028624f
C176 VDD2.n146 VSUBS 0.015381f
C177 VDD2.n147 VSUBS 0.016286f
C178 VDD2.n148 VSUBS 0.036356f
C179 VDD2.n149 VSUBS 0.036356f
C180 VDD2.n150 VSUBS 0.016286f
C181 VDD2.n151 VSUBS 0.015381f
C182 VDD2.n152 VSUBS 0.028624f
C183 VDD2.n153 VSUBS 0.028624f
C184 VDD2.n154 VSUBS 0.015381f
C185 VDD2.n155 VSUBS 0.016286f
C186 VDD2.n156 VSUBS 0.036356f
C187 VDD2.n157 VSUBS 0.036356f
C188 VDD2.n158 VSUBS 0.016286f
C189 VDD2.n159 VSUBS 0.015381f
C190 VDD2.n160 VSUBS 0.028624f
C191 VDD2.n161 VSUBS 0.028624f
C192 VDD2.n162 VSUBS 0.015381f
C193 VDD2.n163 VSUBS 0.016286f
C194 VDD2.n164 VSUBS 0.036356f
C195 VDD2.n165 VSUBS 0.088846f
C196 VDD2.n166 VSUBS 0.016286f
C197 VDD2.n167 VSUBS 0.015381f
C198 VDD2.n168 VSUBS 0.073593f
C199 VDD2.n169 VSUBS 0.064647f
C200 VDD2.n170 VSUBS 3.96048f
C201 VN.t1 VSUBS 4.48872f
C202 VN.t0 VSUBS 5.16967f
C203 B.n0 VSUBS 0.005631f
C204 B.n1 VSUBS 0.005631f
C205 B.n2 VSUBS 0.008328f
C206 B.n3 VSUBS 0.006382f
C207 B.n4 VSUBS 0.006382f
C208 B.n5 VSUBS 0.006382f
C209 B.n6 VSUBS 0.006382f
C210 B.n7 VSUBS 0.006382f
C211 B.n8 VSUBS 0.006382f
C212 B.n9 VSUBS 0.006382f
C213 B.n10 VSUBS 0.006382f
C214 B.n11 VSUBS 0.006382f
C215 B.n12 VSUBS 0.006382f
C216 B.n13 VSUBS 0.006382f
C217 B.n14 VSUBS 0.01396f
C218 B.n15 VSUBS 0.006382f
C219 B.n16 VSUBS 0.006382f
C220 B.n17 VSUBS 0.006382f
C221 B.n18 VSUBS 0.006382f
C222 B.n19 VSUBS 0.006382f
C223 B.n20 VSUBS 0.006382f
C224 B.n21 VSUBS 0.006382f
C225 B.n22 VSUBS 0.006382f
C226 B.n23 VSUBS 0.006382f
C227 B.n24 VSUBS 0.006382f
C228 B.n25 VSUBS 0.006382f
C229 B.n26 VSUBS 0.006382f
C230 B.n27 VSUBS 0.006382f
C231 B.n28 VSUBS 0.006382f
C232 B.n29 VSUBS 0.006382f
C233 B.n30 VSUBS 0.006382f
C234 B.n31 VSUBS 0.006382f
C235 B.n32 VSUBS 0.006382f
C236 B.n33 VSUBS 0.006382f
C237 B.n34 VSUBS 0.006382f
C238 B.n35 VSUBS 0.006382f
C239 B.n36 VSUBS 0.006382f
C240 B.n37 VSUBS 0.006382f
C241 B.n38 VSUBS 0.006382f
C242 B.n39 VSUBS 0.006382f
C243 B.n40 VSUBS 0.006007f
C244 B.n41 VSUBS 0.006382f
C245 B.t1 VSUBS 0.266822f
C246 B.t2 VSUBS 0.297219f
C247 B.t0 VSUBS 1.67168f
C248 B.n42 VSUBS 0.46081f
C249 B.n43 VSUBS 0.272308f
C250 B.n44 VSUBS 0.014787f
C251 B.n45 VSUBS 0.006382f
C252 B.n46 VSUBS 0.006382f
C253 B.n47 VSUBS 0.006382f
C254 B.n48 VSUBS 0.006382f
C255 B.t10 VSUBS 0.266825f
C256 B.t11 VSUBS 0.297221f
C257 B.t9 VSUBS 1.67168f
C258 B.n49 VSUBS 0.460807f
C259 B.n50 VSUBS 0.272305f
C260 B.n51 VSUBS 0.006382f
C261 B.n52 VSUBS 0.006382f
C262 B.n53 VSUBS 0.006382f
C263 B.n54 VSUBS 0.006382f
C264 B.n55 VSUBS 0.006382f
C265 B.n56 VSUBS 0.006382f
C266 B.n57 VSUBS 0.006382f
C267 B.n58 VSUBS 0.006382f
C268 B.n59 VSUBS 0.006382f
C269 B.n60 VSUBS 0.006382f
C270 B.n61 VSUBS 0.006382f
C271 B.n62 VSUBS 0.006382f
C272 B.n63 VSUBS 0.006382f
C273 B.n64 VSUBS 0.006382f
C274 B.n65 VSUBS 0.006382f
C275 B.n66 VSUBS 0.006382f
C276 B.n67 VSUBS 0.006382f
C277 B.n68 VSUBS 0.006382f
C278 B.n69 VSUBS 0.006382f
C279 B.n70 VSUBS 0.006382f
C280 B.n71 VSUBS 0.006382f
C281 B.n72 VSUBS 0.006382f
C282 B.n73 VSUBS 0.006382f
C283 B.n74 VSUBS 0.006382f
C284 B.n75 VSUBS 0.006382f
C285 B.n76 VSUBS 0.014946f
C286 B.n77 VSUBS 0.006382f
C287 B.n78 VSUBS 0.006382f
C288 B.n79 VSUBS 0.006382f
C289 B.n80 VSUBS 0.006382f
C290 B.n81 VSUBS 0.006382f
C291 B.n82 VSUBS 0.006382f
C292 B.n83 VSUBS 0.006382f
C293 B.n84 VSUBS 0.006382f
C294 B.n85 VSUBS 0.006382f
C295 B.n86 VSUBS 0.006382f
C296 B.n87 VSUBS 0.006382f
C297 B.n88 VSUBS 0.006382f
C298 B.n89 VSUBS 0.006382f
C299 B.n90 VSUBS 0.006382f
C300 B.n91 VSUBS 0.006382f
C301 B.n92 VSUBS 0.006382f
C302 B.n93 VSUBS 0.006382f
C303 B.n94 VSUBS 0.006382f
C304 B.n95 VSUBS 0.006382f
C305 B.n96 VSUBS 0.006382f
C306 B.n97 VSUBS 0.006382f
C307 B.n98 VSUBS 0.006382f
C308 B.n99 VSUBS 0.006382f
C309 B.n100 VSUBS 0.006382f
C310 B.n101 VSUBS 0.006382f
C311 B.n102 VSUBS 0.01396f
C312 B.n103 VSUBS 0.006382f
C313 B.n104 VSUBS 0.006382f
C314 B.n105 VSUBS 0.006382f
C315 B.n106 VSUBS 0.006382f
C316 B.n107 VSUBS 0.006382f
C317 B.n108 VSUBS 0.006382f
C318 B.n109 VSUBS 0.006382f
C319 B.n110 VSUBS 0.006382f
C320 B.n111 VSUBS 0.006382f
C321 B.n112 VSUBS 0.006382f
C322 B.n113 VSUBS 0.006382f
C323 B.n114 VSUBS 0.006382f
C324 B.n115 VSUBS 0.006382f
C325 B.n116 VSUBS 0.006382f
C326 B.n117 VSUBS 0.006382f
C327 B.n118 VSUBS 0.006382f
C328 B.n119 VSUBS 0.006382f
C329 B.n120 VSUBS 0.006382f
C330 B.n121 VSUBS 0.006382f
C331 B.n122 VSUBS 0.006382f
C332 B.n123 VSUBS 0.006382f
C333 B.n124 VSUBS 0.006382f
C334 B.n125 VSUBS 0.006382f
C335 B.n126 VSUBS 0.006382f
C336 B.n127 VSUBS 0.006382f
C337 B.n128 VSUBS 0.006382f
C338 B.t8 VSUBS 0.266825f
C339 B.t7 VSUBS 0.297221f
C340 B.t6 VSUBS 1.67168f
C341 B.n129 VSUBS 0.460807f
C342 B.n130 VSUBS 0.272305f
C343 B.n131 VSUBS 0.006382f
C344 B.n132 VSUBS 0.006382f
C345 B.n133 VSUBS 0.006382f
C346 B.n134 VSUBS 0.006382f
C347 B.n135 VSUBS 0.003566f
C348 B.n136 VSUBS 0.006382f
C349 B.n137 VSUBS 0.006382f
C350 B.n138 VSUBS 0.006382f
C351 B.n139 VSUBS 0.006382f
C352 B.n140 VSUBS 0.006382f
C353 B.n141 VSUBS 0.006382f
C354 B.n142 VSUBS 0.006382f
C355 B.n143 VSUBS 0.006382f
C356 B.n144 VSUBS 0.006382f
C357 B.n145 VSUBS 0.006382f
C358 B.n146 VSUBS 0.006382f
C359 B.n147 VSUBS 0.006382f
C360 B.n148 VSUBS 0.006382f
C361 B.n149 VSUBS 0.006382f
C362 B.n150 VSUBS 0.006382f
C363 B.n151 VSUBS 0.006382f
C364 B.n152 VSUBS 0.006382f
C365 B.n153 VSUBS 0.006382f
C366 B.n154 VSUBS 0.006382f
C367 B.n155 VSUBS 0.006382f
C368 B.n156 VSUBS 0.006382f
C369 B.n157 VSUBS 0.006382f
C370 B.n158 VSUBS 0.006382f
C371 B.n159 VSUBS 0.006382f
C372 B.n160 VSUBS 0.006382f
C373 B.n161 VSUBS 0.014946f
C374 B.n162 VSUBS 0.006382f
C375 B.n163 VSUBS 0.006382f
C376 B.n164 VSUBS 0.006382f
C377 B.n165 VSUBS 0.006382f
C378 B.n166 VSUBS 0.006382f
C379 B.n167 VSUBS 0.006382f
C380 B.n168 VSUBS 0.006382f
C381 B.n169 VSUBS 0.006382f
C382 B.n170 VSUBS 0.006382f
C383 B.n171 VSUBS 0.006382f
C384 B.n172 VSUBS 0.006382f
C385 B.n173 VSUBS 0.006382f
C386 B.n174 VSUBS 0.006382f
C387 B.n175 VSUBS 0.006382f
C388 B.n176 VSUBS 0.006382f
C389 B.n177 VSUBS 0.006382f
C390 B.n178 VSUBS 0.006382f
C391 B.n179 VSUBS 0.006382f
C392 B.n180 VSUBS 0.006382f
C393 B.n181 VSUBS 0.006382f
C394 B.n182 VSUBS 0.006382f
C395 B.n183 VSUBS 0.006382f
C396 B.n184 VSUBS 0.006382f
C397 B.n185 VSUBS 0.006382f
C398 B.n186 VSUBS 0.006382f
C399 B.n187 VSUBS 0.006382f
C400 B.n188 VSUBS 0.006382f
C401 B.n189 VSUBS 0.006382f
C402 B.n190 VSUBS 0.006382f
C403 B.n191 VSUBS 0.006382f
C404 B.n192 VSUBS 0.006382f
C405 B.n193 VSUBS 0.006382f
C406 B.n194 VSUBS 0.006382f
C407 B.n195 VSUBS 0.006382f
C408 B.n196 VSUBS 0.006382f
C409 B.n197 VSUBS 0.006382f
C410 B.n198 VSUBS 0.006382f
C411 B.n199 VSUBS 0.006382f
C412 B.n200 VSUBS 0.006382f
C413 B.n201 VSUBS 0.006382f
C414 B.n202 VSUBS 0.006382f
C415 B.n203 VSUBS 0.006382f
C416 B.n204 VSUBS 0.006382f
C417 B.n205 VSUBS 0.006382f
C418 B.n206 VSUBS 0.006382f
C419 B.n207 VSUBS 0.006382f
C420 B.n208 VSUBS 0.01396f
C421 B.n209 VSUBS 0.01396f
C422 B.n210 VSUBS 0.014946f
C423 B.n211 VSUBS 0.006382f
C424 B.n212 VSUBS 0.006382f
C425 B.n213 VSUBS 0.006382f
C426 B.n214 VSUBS 0.006382f
C427 B.n215 VSUBS 0.006382f
C428 B.n216 VSUBS 0.006382f
C429 B.n217 VSUBS 0.006382f
C430 B.n218 VSUBS 0.006382f
C431 B.n219 VSUBS 0.006382f
C432 B.n220 VSUBS 0.006382f
C433 B.n221 VSUBS 0.006382f
C434 B.n222 VSUBS 0.006382f
C435 B.n223 VSUBS 0.006382f
C436 B.n224 VSUBS 0.006382f
C437 B.n225 VSUBS 0.006382f
C438 B.n226 VSUBS 0.006382f
C439 B.n227 VSUBS 0.006382f
C440 B.n228 VSUBS 0.006382f
C441 B.n229 VSUBS 0.006382f
C442 B.n230 VSUBS 0.006382f
C443 B.n231 VSUBS 0.006382f
C444 B.n232 VSUBS 0.006382f
C445 B.n233 VSUBS 0.006382f
C446 B.n234 VSUBS 0.006382f
C447 B.n235 VSUBS 0.006382f
C448 B.n236 VSUBS 0.006382f
C449 B.n237 VSUBS 0.006382f
C450 B.n238 VSUBS 0.006382f
C451 B.n239 VSUBS 0.006382f
C452 B.n240 VSUBS 0.006382f
C453 B.n241 VSUBS 0.006382f
C454 B.n242 VSUBS 0.006382f
C455 B.n243 VSUBS 0.006382f
C456 B.n244 VSUBS 0.006382f
C457 B.n245 VSUBS 0.006382f
C458 B.n246 VSUBS 0.006382f
C459 B.n247 VSUBS 0.006382f
C460 B.n248 VSUBS 0.006382f
C461 B.n249 VSUBS 0.006382f
C462 B.n250 VSUBS 0.006382f
C463 B.n251 VSUBS 0.006382f
C464 B.n252 VSUBS 0.006382f
C465 B.n253 VSUBS 0.006382f
C466 B.n254 VSUBS 0.006382f
C467 B.n255 VSUBS 0.006382f
C468 B.n256 VSUBS 0.006382f
C469 B.n257 VSUBS 0.006382f
C470 B.n258 VSUBS 0.006382f
C471 B.n259 VSUBS 0.006382f
C472 B.n260 VSUBS 0.006382f
C473 B.n261 VSUBS 0.006382f
C474 B.n262 VSUBS 0.006382f
C475 B.n263 VSUBS 0.006382f
C476 B.n264 VSUBS 0.006382f
C477 B.n265 VSUBS 0.006382f
C478 B.n266 VSUBS 0.006382f
C479 B.n267 VSUBS 0.006382f
C480 B.n268 VSUBS 0.006382f
C481 B.n269 VSUBS 0.006382f
C482 B.n270 VSUBS 0.006382f
C483 B.n271 VSUBS 0.006382f
C484 B.n272 VSUBS 0.006382f
C485 B.n273 VSUBS 0.006382f
C486 B.n274 VSUBS 0.006382f
C487 B.n275 VSUBS 0.006382f
C488 B.n276 VSUBS 0.006382f
C489 B.n277 VSUBS 0.006382f
C490 B.n278 VSUBS 0.006382f
C491 B.n279 VSUBS 0.006382f
C492 B.n280 VSUBS 0.006382f
C493 B.n281 VSUBS 0.006382f
C494 B.n282 VSUBS 0.006382f
C495 B.n283 VSUBS 0.006382f
C496 B.n284 VSUBS 0.006382f
C497 B.n285 VSUBS 0.006382f
C498 B.t5 VSUBS 0.266822f
C499 B.t4 VSUBS 0.297219f
C500 B.t3 VSUBS 1.67168f
C501 B.n286 VSUBS 0.46081f
C502 B.n287 VSUBS 0.272308f
C503 B.n288 VSUBS 0.014787f
C504 B.n289 VSUBS 0.006007f
C505 B.n290 VSUBS 0.006382f
C506 B.n291 VSUBS 0.006382f
C507 B.n292 VSUBS 0.006382f
C508 B.n293 VSUBS 0.006382f
C509 B.n294 VSUBS 0.006382f
C510 B.n295 VSUBS 0.006382f
C511 B.n296 VSUBS 0.006382f
C512 B.n297 VSUBS 0.006382f
C513 B.n298 VSUBS 0.006382f
C514 B.n299 VSUBS 0.006382f
C515 B.n300 VSUBS 0.006382f
C516 B.n301 VSUBS 0.006382f
C517 B.n302 VSUBS 0.006382f
C518 B.n303 VSUBS 0.006382f
C519 B.n304 VSUBS 0.006382f
C520 B.n305 VSUBS 0.003566f
C521 B.n306 VSUBS 0.014787f
C522 B.n307 VSUBS 0.006007f
C523 B.n308 VSUBS 0.006382f
C524 B.n309 VSUBS 0.006382f
C525 B.n310 VSUBS 0.006382f
C526 B.n311 VSUBS 0.006382f
C527 B.n312 VSUBS 0.006382f
C528 B.n313 VSUBS 0.006382f
C529 B.n314 VSUBS 0.006382f
C530 B.n315 VSUBS 0.006382f
C531 B.n316 VSUBS 0.006382f
C532 B.n317 VSUBS 0.006382f
C533 B.n318 VSUBS 0.006382f
C534 B.n319 VSUBS 0.006382f
C535 B.n320 VSUBS 0.006382f
C536 B.n321 VSUBS 0.006382f
C537 B.n322 VSUBS 0.006382f
C538 B.n323 VSUBS 0.006382f
C539 B.n324 VSUBS 0.006382f
C540 B.n325 VSUBS 0.006382f
C541 B.n326 VSUBS 0.006382f
C542 B.n327 VSUBS 0.006382f
C543 B.n328 VSUBS 0.006382f
C544 B.n329 VSUBS 0.006382f
C545 B.n330 VSUBS 0.006382f
C546 B.n331 VSUBS 0.006382f
C547 B.n332 VSUBS 0.006382f
C548 B.n333 VSUBS 0.006382f
C549 B.n334 VSUBS 0.006382f
C550 B.n335 VSUBS 0.006382f
C551 B.n336 VSUBS 0.006382f
C552 B.n337 VSUBS 0.006382f
C553 B.n338 VSUBS 0.006382f
C554 B.n339 VSUBS 0.006382f
C555 B.n340 VSUBS 0.006382f
C556 B.n341 VSUBS 0.006382f
C557 B.n342 VSUBS 0.006382f
C558 B.n343 VSUBS 0.006382f
C559 B.n344 VSUBS 0.006382f
C560 B.n345 VSUBS 0.006382f
C561 B.n346 VSUBS 0.006382f
C562 B.n347 VSUBS 0.006382f
C563 B.n348 VSUBS 0.006382f
C564 B.n349 VSUBS 0.006382f
C565 B.n350 VSUBS 0.006382f
C566 B.n351 VSUBS 0.006382f
C567 B.n352 VSUBS 0.006382f
C568 B.n353 VSUBS 0.006382f
C569 B.n354 VSUBS 0.006382f
C570 B.n355 VSUBS 0.006382f
C571 B.n356 VSUBS 0.006382f
C572 B.n357 VSUBS 0.006382f
C573 B.n358 VSUBS 0.006382f
C574 B.n359 VSUBS 0.006382f
C575 B.n360 VSUBS 0.006382f
C576 B.n361 VSUBS 0.006382f
C577 B.n362 VSUBS 0.006382f
C578 B.n363 VSUBS 0.006382f
C579 B.n364 VSUBS 0.006382f
C580 B.n365 VSUBS 0.006382f
C581 B.n366 VSUBS 0.006382f
C582 B.n367 VSUBS 0.006382f
C583 B.n368 VSUBS 0.006382f
C584 B.n369 VSUBS 0.006382f
C585 B.n370 VSUBS 0.006382f
C586 B.n371 VSUBS 0.006382f
C587 B.n372 VSUBS 0.006382f
C588 B.n373 VSUBS 0.006382f
C589 B.n374 VSUBS 0.006382f
C590 B.n375 VSUBS 0.006382f
C591 B.n376 VSUBS 0.006382f
C592 B.n377 VSUBS 0.006382f
C593 B.n378 VSUBS 0.006382f
C594 B.n379 VSUBS 0.006382f
C595 B.n380 VSUBS 0.006382f
C596 B.n381 VSUBS 0.006382f
C597 B.n382 VSUBS 0.006382f
C598 B.n383 VSUBS 0.014946f
C599 B.n384 VSUBS 0.014154f
C600 B.n385 VSUBS 0.014753f
C601 B.n386 VSUBS 0.006382f
C602 B.n387 VSUBS 0.006382f
C603 B.n388 VSUBS 0.006382f
C604 B.n389 VSUBS 0.006382f
C605 B.n390 VSUBS 0.006382f
C606 B.n391 VSUBS 0.006382f
C607 B.n392 VSUBS 0.006382f
C608 B.n393 VSUBS 0.006382f
C609 B.n394 VSUBS 0.006382f
C610 B.n395 VSUBS 0.006382f
C611 B.n396 VSUBS 0.006382f
C612 B.n397 VSUBS 0.006382f
C613 B.n398 VSUBS 0.006382f
C614 B.n399 VSUBS 0.006382f
C615 B.n400 VSUBS 0.006382f
C616 B.n401 VSUBS 0.006382f
C617 B.n402 VSUBS 0.006382f
C618 B.n403 VSUBS 0.006382f
C619 B.n404 VSUBS 0.006382f
C620 B.n405 VSUBS 0.006382f
C621 B.n406 VSUBS 0.006382f
C622 B.n407 VSUBS 0.006382f
C623 B.n408 VSUBS 0.006382f
C624 B.n409 VSUBS 0.006382f
C625 B.n410 VSUBS 0.006382f
C626 B.n411 VSUBS 0.006382f
C627 B.n412 VSUBS 0.006382f
C628 B.n413 VSUBS 0.006382f
C629 B.n414 VSUBS 0.006382f
C630 B.n415 VSUBS 0.006382f
C631 B.n416 VSUBS 0.006382f
C632 B.n417 VSUBS 0.006382f
C633 B.n418 VSUBS 0.006382f
C634 B.n419 VSUBS 0.006382f
C635 B.n420 VSUBS 0.006382f
C636 B.n421 VSUBS 0.006382f
C637 B.n422 VSUBS 0.006382f
C638 B.n423 VSUBS 0.006382f
C639 B.n424 VSUBS 0.006382f
C640 B.n425 VSUBS 0.006382f
C641 B.n426 VSUBS 0.006382f
C642 B.n427 VSUBS 0.006382f
C643 B.n428 VSUBS 0.006382f
C644 B.n429 VSUBS 0.006382f
C645 B.n430 VSUBS 0.006382f
C646 B.n431 VSUBS 0.006382f
C647 B.n432 VSUBS 0.006382f
C648 B.n433 VSUBS 0.006382f
C649 B.n434 VSUBS 0.006382f
C650 B.n435 VSUBS 0.006382f
C651 B.n436 VSUBS 0.006382f
C652 B.n437 VSUBS 0.006382f
C653 B.n438 VSUBS 0.006382f
C654 B.n439 VSUBS 0.006382f
C655 B.n440 VSUBS 0.006382f
C656 B.n441 VSUBS 0.006382f
C657 B.n442 VSUBS 0.006382f
C658 B.n443 VSUBS 0.006382f
C659 B.n444 VSUBS 0.006382f
C660 B.n445 VSUBS 0.006382f
C661 B.n446 VSUBS 0.006382f
C662 B.n447 VSUBS 0.006382f
C663 B.n448 VSUBS 0.006382f
C664 B.n449 VSUBS 0.006382f
C665 B.n450 VSUBS 0.006382f
C666 B.n451 VSUBS 0.006382f
C667 B.n452 VSUBS 0.006382f
C668 B.n453 VSUBS 0.006382f
C669 B.n454 VSUBS 0.006382f
C670 B.n455 VSUBS 0.006382f
C671 B.n456 VSUBS 0.006382f
C672 B.n457 VSUBS 0.006382f
C673 B.n458 VSUBS 0.006382f
C674 B.n459 VSUBS 0.006382f
C675 B.n460 VSUBS 0.006382f
C676 B.n461 VSUBS 0.01396f
C677 B.n462 VSUBS 0.01396f
C678 B.n463 VSUBS 0.014946f
C679 B.n464 VSUBS 0.006382f
C680 B.n465 VSUBS 0.006382f
C681 B.n466 VSUBS 0.006382f
C682 B.n467 VSUBS 0.006382f
C683 B.n468 VSUBS 0.006382f
C684 B.n469 VSUBS 0.006382f
C685 B.n470 VSUBS 0.006382f
C686 B.n471 VSUBS 0.006382f
C687 B.n472 VSUBS 0.006382f
C688 B.n473 VSUBS 0.006382f
C689 B.n474 VSUBS 0.006382f
C690 B.n475 VSUBS 0.006382f
C691 B.n476 VSUBS 0.006382f
C692 B.n477 VSUBS 0.006382f
C693 B.n478 VSUBS 0.006382f
C694 B.n479 VSUBS 0.006382f
C695 B.n480 VSUBS 0.006382f
C696 B.n481 VSUBS 0.006382f
C697 B.n482 VSUBS 0.006382f
C698 B.n483 VSUBS 0.006382f
C699 B.n484 VSUBS 0.006382f
C700 B.n485 VSUBS 0.006382f
C701 B.n486 VSUBS 0.006382f
C702 B.n487 VSUBS 0.006382f
C703 B.n488 VSUBS 0.006382f
C704 B.n489 VSUBS 0.006382f
C705 B.n490 VSUBS 0.006382f
C706 B.n491 VSUBS 0.006382f
C707 B.n492 VSUBS 0.006382f
C708 B.n493 VSUBS 0.006382f
C709 B.n494 VSUBS 0.006382f
C710 B.n495 VSUBS 0.006382f
C711 B.n496 VSUBS 0.006382f
C712 B.n497 VSUBS 0.006382f
C713 B.n498 VSUBS 0.006382f
C714 B.n499 VSUBS 0.006382f
C715 B.n500 VSUBS 0.006382f
C716 B.n501 VSUBS 0.006382f
C717 B.n502 VSUBS 0.006382f
C718 B.n503 VSUBS 0.006382f
C719 B.n504 VSUBS 0.006382f
C720 B.n505 VSUBS 0.006382f
C721 B.n506 VSUBS 0.006382f
C722 B.n507 VSUBS 0.006382f
C723 B.n508 VSUBS 0.006382f
C724 B.n509 VSUBS 0.006382f
C725 B.n510 VSUBS 0.006382f
C726 B.n511 VSUBS 0.006382f
C727 B.n512 VSUBS 0.006382f
C728 B.n513 VSUBS 0.006382f
C729 B.n514 VSUBS 0.006382f
C730 B.n515 VSUBS 0.006382f
C731 B.n516 VSUBS 0.006382f
C732 B.n517 VSUBS 0.006382f
C733 B.n518 VSUBS 0.006382f
C734 B.n519 VSUBS 0.006382f
C735 B.n520 VSUBS 0.006382f
C736 B.n521 VSUBS 0.006382f
C737 B.n522 VSUBS 0.006382f
C738 B.n523 VSUBS 0.006382f
C739 B.n524 VSUBS 0.006382f
C740 B.n525 VSUBS 0.006382f
C741 B.n526 VSUBS 0.006382f
C742 B.n527 VSUBS 0.006382f
C743 B.n528 VSUBS 0.006382f
C744 B.n529 VSUBS 0.006382f
C745 B.n530 VSUBS 0.006382f
C746 B.n531 VSUBS 0.006382f
C747 B.n532 VSUBS 0.006382f
C748 B.n533 VSUBS 0.006382f
C749 B.n534 VSUBS 0.006382f
C750 B.n535 VSUBS 0.006382f
C751 B.n536 VSUBS 0.006382f
C752 B.n537 VSUBS 0.006382f
C753 B.n538 VSUBS 0.006382f
C754 B.n539 VSUBS 0.006382f
C755 B.n540 VSUBS 0.006007f
C756 B.n541 VSUBS 0.014787f
C757 B.n542 VSUBS 0.003566f
C758 B.n543 VSUBS 0.006382f
C759 B.n544 VSUBS 0.006382f
C760 B.n545 VSUBS 0.006382f
C761 B.n546 VSUBS 0.006382f
C762 B.n547 VSUBS 0.006382f
C763 B.n548 VSUBS 0.006382f
C764 B.n549 VSUBS 0.006382f
C765 B.n550 VSUBS 0.006382f
C766 B.n551 VSUBS 0.006382f
C767 B.n552 VSUBS 0.006382f
C768 B.n553 VSUBS 0.006382f
C769 B.n554 VSUBS 0.006382f
C770 B.n555 VSUBS 0.003566f
C771 B.n556 VSUBS 0.006382f
C772 B.n557 VSUBS 0.006382f
C773 B.n558 VSUBS 0.006382f
C774 B.n559 VSUBS 0.006382f
C775 B.n560 VSUBS 0.006382f
C776 B.n561 VSUBS 0.006382f
C777 B.n562 VSUBS 0.006382f
C778 B.n563 VSUBS 0.006382f
C779 B.n564 VSUBS 0.006382f
C780 B.n565 VSUBS 0.006382f
C781 B.n566 VSUBS 0.006382f
C782 B.n567 VSUBS 0.006382f
C783 B.n568 VSUBS 0.006382f
C784 B.n569 VSUBS 0.006382f
C785 B.n570 VSUBS 0.006382f
C786 B.n571 VSUBS 0.006382f
C787 B.n572 VSUBS 0.006382f
C788 B.n573 VSUBS 0.006382f
C789 B.n574 VSUBS 0.006382f
C790 B.n575 VSUBS 0.006382f
C791 B.n576 VSUBS 0.006382f
C792 B.n577 VSUBS 0.006382f
C793 B.n578 VSUBS 0.006382f
C794 B.n579 VSUBS 0.006382f
C795 B.n580 VSUBS 0.006382f
C796 B.n581 VSUBS 0.006382f
C797 B.n582 VSUBS 0.006382f
C798 B.n583 VSUBS 0.006382f
C799 B.n584 VSUBS 0.006382f
C800 B.n585 VSUBS 0.006382f
C801 B.n586 VSUBS 0.006382f
C802 B.n587 VSUBS 0.006382f
C803 B.n588 VSUBS 0.006382f
C804 B.n589 VSUBS 0.006382f
C805 B.n590 VSUBS 0.006382f
C806 B.n591 VSUBS 0.006382f
C807 B.n592 VSUBS 0.006382f
C808 B.n593 VSUBS 0.006382f
C809 B.n594 VSUBS 0.006382f
C810 B.n595 VSUBS 0.006382f
C811 B.n596 VSUBS 0.006382f
C812 B.n597 VSUBS 0.006382f
C813 B.n598 VSUBS 0.006382f
C814 B.n599 VSUBS 0.006382f
C815 B.n600 VSUBS 0.006382f
C816 B.n601 VSUBS 0.006382f
C817 B.n602 VSUBS 0.006382f
C818 B.n603 VSUBS 0.006382f
C819 B.n604 VSUBS 0.006382f
C820 B.n605 VSUBS 0.006382f
C821 B.n606 VSUBS 0.006382f
C822 B.n607 VSUBS 0.006382f
C823 B.n608 VSUBS 0.006382f
C824 B.n609 VSUBS 0.006382f
C825 B.n610 VSUBS 0.006382f
C826 B.n611 VSUBS 0.006382f
C827 B.n612 VSUBS 0.006382f
C828 B.n613 VSUBS 0.006382f
C829 B.n614 VSUBS 0.006382f
C830 B.n615 VSUBS 0.006382f
C831 B.n616 VSUBS 0.006382f
C832 B.n617 VSUBS 0.006382f
C833 B.n618 VSUBS 0.006382f
C834 B.n619 VSUBS 0.006382f
C835 B.n620 VSUBS 0.006382f
C836 B.n621 VSUBS 0.006382f
C837 B.n622 VSUBS 0.006382f
C838 B.n623 VSUBS 0.006382f
C839 B.n624 VSUBS 0.006382f
C840 B.n625 VSUBS 0.006382f
C841 B.n626 VSUBS 0.006382f
C842 B.n627 VSUBS 0.006382f
C843 B.n628 VSUBS 0.006382f
C844 B.n629 VSUBS 0.006382f
C845 B.n630 VSUBS 0.006382f
C846 B.n631 VSUBS 0.006382f
C847 B.n632 VSUBS 0.006382f
C848 B.n633 VSUBS 0.014946f
C849 B.n634 VSUBS 0.014946f
C850 B.n635 VSUBS 0.01396f
C851 B.n636 VSUBS 0.006382f
C852 B.n637 VSUBS 0.006382f
C853 B.n638 VSUBS 0.006382f
C854 B.n639 VSUBS 0.006382f
C855 B.n640 VSUBS 0.006382f
C856 B.n641 VSUBS 0.006382f
C857 B.n642 VSUBS 0.006382f
C858 B.n643 VSUBS 0.006382f
C859 B.n644 VSUBS 0.006382f
C860 B.n645 VSUBS 0.006382f
C861 B.n646 VSUBS 0.006382f
C862 B.n647 VSUBS 0.006382f
C863 B.n648 VSUBS 0.006382f
C864 B.n649 VSUBS 0.006382f
C865 B.n650 VSUBS 0.006382f
C866 B.n651 VSUBS 0.006382f
C867 B.n652 VSUBS 0.006382f
C868 B.n653 VSUBS 0.006382f
C869 B.n654 VSUBS 0.006382f
C870 B.n655 VSUBS 0.006382f
C871 B.n656 VSUBS 0.006382f
C872 B.n657 VSUBS 0.006382f
C873 B.n658 VSUBS 0.006382f
C874 B.n659 VSUBS 0.006382f
C875 B.n660 VSUBS 0.006382f
C876 B.n661 VSUBS 0.006382f
C877 B.n662 VSUBS 0.006382f
C878 B.n663 VSUBS 0.006382f
C879 B.n664 VSUBS 0.006382f
C880 B.n665 VSUBS 0.006382f
C881 B.n666 VSUBS 0.006382f
C882 B.n667 VSUBS 0.006382f
C883 B.n668 VSUBS 0.006382f
C884 B.n669 VSUBS 0.006382f
C885 B.n670 VSUBS 0.006382f
C886 B.n671 VSUBS 0.008328f
C887 B.n672 VSUBS 0.008872f
C888 B.n673 VSUBS 0.017642f
C889 VDD1.n0 VSUBS 0.026862f
C890 VDD1.n1 VSUBS 0.024258f
C891 VDD1.n2 VSUBS 0.013035f
C892 VDD1.n3 VSUBS 0.030811f
C893 VDD1.n4 VSUBS 0.013419f
C894 VDD1.n5 VSUBS 0.024258f
C895 VDD1.n6 VSUBS 0.013419f
C896 VDD1.n7 VSUBS 0.013035f
C897 VDD1.n8 VSUBS 0.030811f
C898 VDD1.n9 VSUBS 0.030811f
C899 VDD1.n10 VSUBS 0.013802f
C900 VDD1.n11 VSUBS 0.024258f
C901 VDD1.n12 VSUBS 0.013035f
C902 VDD1.n13 VSUBS 0.030811f
C903 VDD1.n14 VSUBS 0.013802f
C904 VDD1.n15 VSUBS 0.024258f
C905 VDD1.n16 VSUBS 0.013035f
C906 VDD1.n17 VSUBS 0.030811f
C907 VDD1.n18 VSUBS 0.013802f
C908 VDD1.n19 VSUBS 0.024258f
C909 VDD1.n20 VSUBS 0.013035f
C910 VDD1.n21 VSUBS 0.030811f
C911 VDD1.n22 VSUBS 0.013802f
C912 VDD1.n23 VSUBS 0.024258f
C913 VDD1.n24 VSUBS 0.013035f
C914 VDD1.n25 VSUBS 0.030811f
C915 VDD1.n26 VSUBS 0.013802f
C916 VDD1.n27 VSUBS 1.6095f
C917 VDD1.n28 VSUBS 0.013035f
C918 VDD1.t0 VSUBS 0.065993f
C919 VDD1.n29 VSUBS 0.174935f
C920 VDD1.n30 VSUBS 0.0196f
C921 VDD1.n31 VSUBS 0.023108f
C922 VDD1.n32 VSUBS 0.030811f
C923 VDD1.n33 VSUBS 0.013802f
C924 VDD1.n34 VSUBS 0.013035f
C925 VDD1.n35 VSUBS 0.024258f
C926 VDD1.n36 VSUBS 0.024258f
C927 VDD1.n37 VSUBS 0.013035f
C928 VDD1.n38 VSUBS 0.013802f
C929 VDD1.n39 VSUBS 0.030811f
C930 VDD1.n40 VSUBS 0.030811f
C931 VDD1.n41 VSUBS 0.013802f
C932 VDD1.n42 VSUBS 0.013035f
C933 VDD1.n43 VSUBS 0.024258f
C934 VDD1.n44 VSUBS 0.024258f
C935 VDD1.n45 VSUBS 0.013035f
C936 VDD1.n46 VSUBS 0.013802f
C937 VDD1.n47 VSUBS 0.030811f
C938 VDD1.n48 VSUBS 0.030811f
C939 VDD1.n49 VSUBS 0.013802f
C940 VDD1.n50 VSUBS 0.013035f
C941 VDD1.n51 VSUBS 0.024258f
C942 VDD1.n52 VSUBS 0.024258f
C943 VDD1.n53 VSUBS 0.013035f
C944 VDD1.n54 VSUBS 0.013802f
C945 VDD1.n55 VSUBS 0.030811f
C946 VDD1.n56 VSUBS 0.030811f
C947 VDD1.n57 VSUBS 0.013802f
C948 VDD1.n58 VSUBS 0.013035f
C949 VDD1.n59 VSUBS 0.024258f
C950 VDD1.n60 VSUBS 0.024258f
C951 VDD1.n61 VSUBS 0.013035f
C952 VDD1.n62 VSUBS 0.013802f
C953 VDD1.n63 VSUBS 0.030811f
C954 VDD1.n64 VSUBS 0.030811f
C955 VDD1.n65 VSUBS 0.013802f
C956 VDD1.n66 VSUBS 0.013035f
C957 VDD1.n67 VSUBS 0.024258f
C958 VDD1.n68 VSUBS 0.024258f
C959 VDD1.n69 VSUBS 0.013035f
C960 VDD1.n70 VSUBS 0.013802f
C961 VDD1.n71 VSUBS 0.030811f
C962 VDD1.n72 VSUBS 0.030811f
C963 VDD1.n73 VSUBS 0.013802f
C964 VDD1.n74 VSUBS 0.013035f
C965 VDD1.n75 VSUBS 0.024258f
C966 VDD1.n76 VSUBS 0.024258f
C967 VDD1.n77 VSUBS 0.013035f
C968 VDD1.n78 VSUBS 0.013802f
C969 VDD1.n79 VSUBS 0.030811f
C970 VDD1.n80 VSUBS 0.075295f
C971 VDD1.n81 VSUBS 0.013802f
C972 VDD1.n82 VSUBS 0.013035f
C973 VDD1.n83 VSUBS 0.062368f
C974 VDD1.n84 VSUBS 0.056156f
C975 VDD1.n85 VSUBS 0.026862f
C976 VDD1.n86 VSUBS 0.024258f
C977 VDD1.n87 VSUBS 0.013035f
C978 VDD1.n88 VSUBS 0.030811f
C979 VDD1.n89 VSUBS 0.013419f
C980 VDD1.n90 VSUBS 0.024258f
C981 VDD1.n91 VSUBS 0.013802f
C982 VDD1.n92 VSUBS 0.030811f
C983 VDD1.n93 VSUBS 0.013802f
C984 VDD1.n94 VSUBS 0.024258f
C985 VDD1.n95 VSUBS 0.013035f
C986 VDD1.n96 VSUBS 0.030811f
C987 VDD1.n97 VSUBS 0.013802f
C988 VDD1.n98 VSUBS 0.024258f
C989 VDD1.n99 VSUBS 0.013035f
C990 VDD1.n100 VSUBS 0.030811f
C991 VDD1.n101 VSUBS 0.013802f
C992 VDD1.n102 VSUBS 0.024258f
C993 VDD1.n103 VSUBS 0.013035f
C994 VDD1.n104 VSUBS 0.030811f
C995 VDD1.n105 VSUBS 0.013802f
C996 VDD1.n106 VSUBS 0.024258f
C997 VDD1.n107 VSUBS 0.013035f
C998 VDD1.n108 VSUBS 0.030811f
C999 VDD1.n109 VSUBS 0.013802f
C1000 VDD1.n110 VSUBS 1.6095f
C1001 VDD1.n111 VSUBS 0.013035f
C1002 VDD1.t1 VSUBS 0.065993f
C1003 VDD1.n112 VSUBS 0.174935f
C1004 VDD1.n113 VSUBS 0.0196f
C1005 VDD1.n114 VSUBS 0.023108f
C1006 VDD1.n115 VSUBS 0.030811f
C1007 VDD1.n116 VSUBS 0.013802f
C1008 VDD1.n117 VSUBS 0.013035f
C1009 VDD1.n118 VSUBS 0.024258f
C1010 VDD1.n119 VSUBS 0.024258f
C1011 VDD1.n120 VSUBS 0.013035f
C1012 VDD1.n121 VSUBS 0.013802f
C1013 VDD1.n122 VSUBS 0.030811f
C1014 VDD1.n123 VSUBS 0.030811f
C1015 VDD1.n124 VSUBS 0.013802f
C1016 VDD1.n125 VSUBS 0.013035f
C1017 VDD1.n126 VSUBS 0.024258f
C1018 VDD1.n127 VSUBS 0.024258f
C1019 VDD1.n128 VSUBS 0.013035f
C1020 VDD1.n129 VSUBS 0.013802f
C1021 VDD1.n130 VSUBS 0.030811f
C1022 VDD1.n131 VSUBS 0.030811f
C1023 VDD1.n132 VSUBS 0.013802f
C1024 VDD1.n133 VSUBS 0.013035f
C1025 VDD1.n134 VSUBS 0.024258f
C1026 VDD1.n135 VSUBS 0.024258f
C1027 VDD1.n136 VSUBS 0.013035f
C1028 VDD1.n137 VSUBS 0.013802f
C1029 VDD1.n138 VSUBS 0.030811f
C1030 VDD1.n139 VSUBS 0.030811f
C1031 VDD1.n140 VSUBS 0.013802f
C1032 VDD1.n141 VSUBS 0.013035f
C1033 VDD1.n142 VSUBS 0.024258f
C1034 VDD1.n143 VSUBS 0.024258f
C1035 VDD1.n144 VSUBS 0.013035f
C1036 VDD1.n145 VSUBS 0.013802f
C1037 VDD1.n146 VSUBS 0.030811f
C1038 VDD1.n147 VSUBS 0.030811f
C1039 VDD1.n148 VSUBS 0.013802f
C1040 VDD1.n149 VSUBS 0.013035f
C1041 VDD1.n150 VSUBS 0.024258f
C1042 VDD1.n151 VSUBS 0.024258f
C1043 VDD1.n152 VSUBS 0.013035f
C1044 VDD1.n153 VSUBS 0.013035f
C1045 VDD1.n154 VSUBS 0.013802f
C1046 VDD1.n155 VSUBS 0.030811f
C1047 VDD1.n156 VSUBS 0.030811f
C1048 VDD1.n157 VSUBS 0.030811f
C1049 VDD1.n158 VSUBS 0.013419f
C1050 VDD1.n159 VSUBS 0.013035f
C1051 VDD1.n160 VSUBS 0.024258f
C1052 VDD1.n161 VSUBS 0.024258f
C1053 VDD1.n162 VSUBS 0.013035f
C1054 VDD1.n163 VSUBS 0.013802f
C1055 VDD1.n164 VSUBS 0.030811f
C1056 VDD1.n165 VSUBS 0.075295f
C1057 VDD1.n166 VSUBS 0.013802f
C1058 VDD1.n167 VSUBS 0.013035f
C1059 VDD1.n168 VSUBS 0.062368f
C1060 VDD1.n169 VSUBS 0.862117f
C1061 VTAIL.n0 VSUBS 0.031675f
C1062 VTAIL.n1 VSUBS 0.028605f
C1063 VTAIL.n2 VSUBS 0.015371f
C1064 VTAIL.n3 VSUBS 0.036332f
C1065 VTAIL.n4 VSUBS 0.015823f
C1066 VTAIL.n5 VSUBS 0.028605f
C1067 VTAIL.n6 VSUBS 0.016275f
C1068 VTAIL.n7 VSUBS 0.036332f
C1069 VTAIL.n8 VSUBS 0.016275f
C1070 VTAIL.n9 VSUBS 0.028605f
C1071 VTAIL.n10 VSUBS 0.015371f
C1072 VTAIL.n11 VSUBS 0.036332f
C1073 VTAIL.n12 VSUBS 0.016275f
C1074 VTAIL.n13 VSUBS 0.028605f
C1075 VTAIL.n14 VSUBS 0.015371f
C1076 VTAIL.n15 VSUBS 0.036332f
C1077 VTAIL.n16 VSUBS 0.016275f
C1078 VTAIL.n17 VSUBS 0.028605f
C1079 VTAIL.n18 VSUBS 0.015371f
C1080 VTAIL.n19 VSUBS 0.036332f
C1081 VTAIL.n20 VSUBS 0.016275f
C1082 VTAIL.n21 VSUBS 0.028605f
C1083 VTAIL.n22 VSUBS 0.015371f
C1084 VTAIL.n23 VSUBS 0.036332f
C1085 VTAIL.n24 VSUBS 0.016275f
C1086 VTAIL.n25 VSUBS 1.89792f
C1087 VTAIL.n26 VSUBS 0.015371f
C1088 VTAIL.t2 VSUBS 0.077818f
C1089 VTAIL.n27 VSUBS 0.206282f
C1090 VTAIL.n28 VSUBS 0.023113f
C1091 VTAIL.n29 VSUBS 0.027249f
C1092 VTAIL.n30 VSUBS 0.036332f
C1093 VTAIL.n31 VSUBS 0.016275f
C1094 VTAIL.n32 VSUBS 0.015371f
C1095 VTAIL.n33 VSUBS 0.028605f
C1096 VTAIL.n34 VSUBS 0.028605f
C1097 VTAIL.n35 VSUBS 0.015371f
C1098 VTAIL.n36 VSUBS 0.016275f
C1099 VTAIL.n37 VSUBS 0.036332f
C1100 VTAIL.n38 VSUBS 0.036332f
C1101 VTAIL.n39 VSUBS 0.016275f
C1102 VTAIL.n40 VSUBS 0.015371f
C1103 VTAIL.n41 VSUBS 0.028605f
C1104 VTAIL.n42 VSUBS 0.028605f
C1105 VTAIL.n43 VSUBS 0.015371f
C1106 VTAIL.n44 VSUBS 0.016275f
C1107 VTAIL.n45 VSUBS 0.036332f
C1108 VTAIL.n46 VSUBS 0.036332f
C1109 VTAIL.n47 VSUBS 0.016275f
C1110 VTAIL.n48 VSUBS 0.015371f
C1111 VTAIL.n49 VSUBS 0.028605f
C1112 VTAIL.n50 VSUBS 0.028605f
C1113 VTAIL.n51 VSUBS 0.015371f
C1114 VTAIL.n52 VSUBS 0.016275f
C1115 VTAIL.n53 VSUBS 0.036332f
C1116 VTAIL.n54 VSUBS 0.036332f
C1117 VTAIL.n55 VSUBS 0.016275f
C1118 VTAIL.n56 VSUBS 0.015371f
C1119 VTAIL.n57 VSUBS 0.028605f
C1120 VTAIL.n58 VSUBS 0.028605f
C1121 VTAIL.n59 VSUBS 0.015371f
C1122 VTAIL.n60 VSUBS 0.016275f
C1123 VTAIL.n61 VSUBS 0.036332f
C1124 VTAIL.n62 VSUBS 0.036332f
C1125 VTAIL.n63 VSUBS 0.016275f
C1126 VTAIL.n64 VSUBS 0.015371f
C1127 VTAIL.n65 VSUBS 0.028605f
C1128 VTAIL.n66 VSUBS 0.028605f
C1129 VTAIL.n67 VSUBS 0.015371f
C1130 VTAIL.n68 VSUBS 0.015371f
C1131 VTAIL.n69 VSUBS 0.016275f
C1132 VTAIL.n70 VSUBS 0.036332f
C1133 VTAIL.n71 VSUBS 0.036332f
C1134 VTAIL.n72 VSUBS 0.036332f
C1135 VTAIL.n73 VSUBS 0.015823f
C1136 VTAIL.n74 VSUBS 0.015371f
C1137 VTAIL.n75 VSUBS 0.028605f
C1138 VTAIL.n76 VSUBS 0.028605f
C1139 VTAIL.n77 VSUBS 0.015371f
C1140 VTAIL.n78 VSUBS 0.016275f
C1141 VTAIL.n79 VSUBS 0.036332f
C1142 VTAIL.n80 VSUBS 0.088787f
C1143 VTAIL.n81 VSUBS 0.016275f
C1144 VTAIL.n82 VSUBS 0.015371f
C1145 VTAIL.n83 VSUBS 0.073544f
C1146 VTAIL.n84 VSUBS 0.044905f
C1147 VTAIL.n85 VSUBS 2.23065f
C1148 VTAIL.n86 VSUBS 0.031675f
C1149 VTAIL.n87 VSUBS 0.028605f
C1150 VTAIL.n88 VSUBS 0.015371f
C1151 VTAIL.n89 VSUBS 0.036332f
C1152 VTAIL.n90 VSUBS 0.015823f
C1153 VTAIL.n91 VSUBS 0.028605f
C1154 VTAIL.n92 VSUBS 0.015823f
C1155 VTAIL.n93 VSUBS 0.015371f
C1156 VTAIL.n94 VSUBS 0.036332f
C1157 VTAIL.n95 VSUBS 0.036332f
C1158 VTAIL.n96 VSUBS 0.016275f
C1159 VTAIL.n97 VSUBS 0.028605f
C1160 VTAIL.n98 VSUBS 0.015371f
C1161 VTAIL.n99 VSUBS 0.036332f
C1162 VTAIL.n100 VSUBS 0.016275f
C1163 VTAIL.n101 VSUBS 0.028605f
C1164 VTAIL.n102 VSUBS 0.015371f
C1165 VTAIL.n103 VSUBS 0.036332f
C1166 VTAIL.n104 VSUBS 0.016275f
C1167 VTAIL.n105 VSUBS 0.028605f
C1168 VTAIL.n106 VSUBS 0.015371f
C1169 VTAIL.n107 VSUBS 0.036332f
C1170 VTAIL.n108 VSUBS 0.016275f
C1171 VTAIL.n109 VSUBS 0.028605f
C1172 VTAIL.n110 VSUBS 0.015371f
C1173 VTAIL.n111 VSUBS 0.036332f
C1174 VTAIL.n112 VSUBS 0.016275f
C1175 VTAIL.n113 VSUBS 1.89792f
C1176 VTAIL.n114 VSUBS 0.015371f
C1177 VTAIL.t1 VSUBS 0.077818f
C1178 VTAIL.n115 VSUBS 0.206282f
C1179 VTAIL.n116 VSUBS 0.023113f
C1180 VTAIL.n117 VSUBS 0.027249f
C1181 VTAIL.n118 VSUBS 0.036332f
C1182 VTAIL.n119 VSUBS 0.016275f
C1183 VTAIL.n120 VSUBS 0.015371f
C1184 VTAIL.n121 VSUBS 0.028605f
C1185 VTAIL.n122 VSUBS 0.028605f
C1186 VTAIL.n123 VSUBS 0.015371f
C1187 VTAIL.n124 VSUBS 0.016275f
C1188 VTAIL.n125 VSUBS 0.036332f
C1189 VTAIL.n126 VSUBS 0.036332f
C1190 VTAIL.n127 VSUBS 0.016275f
C1191 VTAIL.n128 VSUBS 0.015371f
C1192 VTAIL.n129 VSUBS 0.028605f
C1193 VTAIL.n130 VSUBS 0.028605f
C1194 VTAIL.n131 VSUBS 0.015371f
C1195 VTAIL.n132 VSUBS 0.016275f
C1196 VTAIL.n133 VSUBS 0.036332f
C1197 VTAIL.n134 VSUBS 0.036332f
C1198 VTAIL.n135 VSUBS 0.016275f
C1199 VTAIL.n136 VSUBS 0.015371f
C1200 VTAIL.n137 VSUBS 0.028605f
C1201 VTAIL.n138 VSUBS 0.028605f
C1202 VTAIL.n139 VSUBS 0.015371f
C1203 VTAIL.n140 VSUBS 0.016275f
C1204 VTAIL.n141 VSUBS 0.036332f
C1205 VTAIL.n142 VSUBS 0.036332f
C1206 VTAIL.n143 VSUBS 0.016275f
C1207 VTAIL.n144 VSUBS 0.015371f
C1208 VTAIL.n145 VSUBS 0.028605f
C1209 VTAIL.n146 VSUBS 0.028605f
C1210 VTAIL.n147 VSUBS 0.015371f
C1211 VTAIL.n148 VSUBS 0.016275f
C1212 VTAIL.n149 VSUBS 0.036332f
C1213 VTAIL.n150 VSUBS 0.036332f
C1214 VTAIL.n151 VSUBS 0.016275f
C1215 VTAIL.n152 VSUBS 0.015371f
C1216 VTAIL.n153 VSUBS 0.028605f
C1217 VTAIL.n154 VSUBS 0.028605f
C1218 VTAIL.n155 VSUBS 0.015371f
C1219 VTAIL.n156 VSUBS 0.016275f
C1220 VTAIL.n157 VSUBS 0.036332f
C1221 VTAIL.n158 VSUBS 0.036332f
C1222 VTAIL.n159 VSUBS 0.016275f
C1223 VTAIL.n160 VSUBS 0.015371f
C1224 VTAIL.n161 VSUBS 0.028605f
C1225 VTAIL.n162 VSUBS 0.028605f
C1226 VTAIL.n163 VSUBS 0.015371f
C1227 VTAIL.n164 VSUBS 0.016275f
C1228 VTAIL.n165 VSUBS 0.036332f
C1229 VTAIL.n166 VSUBS 0.088787f
C1230 VTAIL.n167 VSUBS 0.016275f
C1231 VTAIL.n168 VSUBS 0.015371f
C1232 VTAIL.n169 VSUBS 0.073544f
C1233 VTAIL.n170 VSUBS 0.044905f
C1234 VTAIL.n171 VSUBS 2.28408f
C1235 VTAIL.n172 VSUBS 0.031675f
C1236 VTAIL.n173 VSUBS 0.028605f
C1237 VTAIL.n174 VSUBS 0.015371f
C1238 VTAIL.n175 VSUBS 0.036332f
C1239 VTAIL.n176 VSUBS 0.015823f
C1240 VTAIL.n177 VSUBS 0.028605f
C1241 VTAIL.n178 VSUBS 0.015823f
C1242 VTAIL.n179 VSUBS 0.015371f
C1243 VTAIL.n180 VSUBS 0.036332f
C1244 VTAIL.n181 VSUBS 0.036332f
C1245 VTAIL.n182 VSUBS 0.016275f
C1246 VTAIL.n183 VSUBS 0.028605f
C1247 VTAIL.n184 VSUBS 0.015371f
C1248 VTAIL.n185 VSUBS 0.036332f
C1249 VTAIL.n186 VSUBS 0.016275f
C1250 VTAIL.n187 VSUBS 0.028605f
C1251 VTAIL.n188 VSUBS 0.015371f
C1252 VTAIL.n189 VSUBS 0.036332f
C1253 VTAIL.n190 VSUBS 0.016275f
C1254 VTAIL.n191 VSUBS 0.028605f
C1255 VTAIL.n192 VSUBS 0.015371f
C1256 VTAIL.n193 VSUBS 0.036332f
C1257 VTAIL.n194 VSUBS 0.016275f
C1258 VTAIL.n195 VSUBS 0.028605f
C1259 VTAIL.n196 VSUBS 0.015371f
C1260 VTAIL.n197 VSUBS 0.036332f
C1261 VTAIL.n198 VSUBS 0.016275f
C1262 VTAIL.n199 VSUBS 1.89792f
C1263 VTAIL.n200 VSUBS 0.015371f
C1264 VTAIL.t3 VSUBS 0.077818f
C1265 VTAIL.n201 VSUBS 0.206282f
C1266 VTAIL.n202 VSUBS 0.023113f
C1267 VTAIL.n203 VSUBS 0.027249f
C1268 VTAIL.n204 VSUBS 0.036332f
C1269 VTAIL.n205 VSUBS 0.016275f
C1270 VTAIL.n206 VSUBS 0.015371f
C1271 VTAIL.n207 VSUBS 0.028605f
C1272 VTAIL.n208 VSUBS 0.028605f
C1273 VTAIL.n209 VSUBS 0.015371f
C1274 VTAIL.n210 VSUBS 0.016275f
C1275 VTAIL.n211 VSUBS 0.036332f
C1276 VTAIL.n212 VSUBS 0.036332f
C1277 VTAIL.n213 VSUBS 0.016275f
C1278 VTAIL.n214 VSUBS 0.015371f
C1279 VTAIL.n215 VSUBS 0.028605f
C1280 VTAIL.n216 VSUBS 0.028605f
C1281 VTAIL.n217 VSUBS 0.015371f
C1282 VTAIL.n218 VSUBS 0.016275f
C1283 VTAIL.n219 VSUBS 0.036332f
C1284 VTAIL.n220 VSUBS 0.036332f
C1285 VTAIL.n221 VSUBS 0.016275f
C1286 VTAIL.n222 VSUBS 0.015371f
C1287 VTAIL.n223 VSUBS 0.028605f
C1288 VTAIL.n224 VSUBS 0.028605f
C1289 VTAIL.n225 VSUBS 0.015371f
C1290 VTAIL.n226 VSUBS 0.016275f
C1291 VTAIL.n227 VSUBS 0.036332f
C1292 VTAIL.n228 VSUBS 0.036332f
C1293 VTAIL.n229 VSUBS 0.016275f
C1294 VTAIL.n230 VSUBS 0.015371f
C1295 VTAIL.n231 VSUBS 0.028605f
C1296 VTAIL.n232 VSUBS 0.028605f
C1297 VTAIL.n233 VSUBS 0.015371f
C1298 VTAIL.n234 VSUBS 0.016275f
C1299 VTAIL.n235 VSUBS 0.036332f
C1300 VTAIL.n236 VSUBS 0.036332f
C1301 VTAIL.n237 VSUBS 0.016275f
C1302 VTAIL.n238 VSUBS 0.015371f
C1303 VTAIL.n239 VSUBS 0.028605f
C1304 VTAIL.n240 VSUBS 0.028605f
C1305 VTAIL.n241 VSUBS 0.015371f
C1306 VTAIL.n242 VSUBS 0.016275f
C1307 VTAIL.n243 VSUBS 0.036332f
C1308 VTAIL.n244 VSUBS 0.036332f
C1309 VTAIL.n245 VSUBS 0.016275f
C1310 VTAIL.n246 VSUBS 0.015371f
C1311 VTAIL.n247 VSUBS 0.028605f
C1312 VTAIL.n248 VSUBS 0.028605f
C1313 VTAIL.n249 VSUBS 0.015371f
C1314 VTAIL.n250 VSUBS 0.016275f
C1315 VTAIL.n251 VSUBS 0.036332f
C1316 VTAIL.n252 VSUBS 0.088787f
C1317 VTAIL.n253 VSUBS 0.016275f
C1318 VTAIL.n254 VSUBS 0.015371f
C1319 VTAIL.n255 VSUBS 0.073544f
C1320 VTAIL.n256 VSUBS 0.044905f
C1321 VTAIL.n257 VSUBS 2.04889f
C1322 VTAIL.n258 VSUBS 0.031675f
C1323 VTAIL.n259 VSUBS 0.028605f
C1324 VTAIL.n260 VSUBS 0.015371f
C1325 VTAIL.n261 VSUBS 0.036332f
C1326 VTAIL.n262 VSUBS 0.015823f
C1327 VTAIL.n263 VSUBS 0.028605f
C1328 VTAIL.n264 VSUBS 0.016275f
C1329 VTAIL.n265 VSUBS 0.036332f
C1330 VTAIL.n266 VSUBS 0.016275f
C1331 VTAIL.n267 VSUBS 0.028605f
C1332 VTAIL.n268 VSUBS 0.015371f
C1333 VTAIL.n269 VSUBS 0.036332f
C1334 VTAIL.n270 VSUBS 0.016275f
C1335 VTAIL.n271 VSUBS 0.028605f
C1336 VTAIL.n272 VSUBS 0.015371f
C1337 VTAIL.n273 VSUBS 0.036332f
C1338 VTAIL.n274 VSUBS 0.016275f
C1339 VTAIL.n275 VSUBS 0.028605f
C1340 VTAIL.n276 VSUBS 0.015371f
C1341 VTAIL.n277 VSUBS 0.036332f
C1342 VTAIL.n278 VSUBS 0.016275f
C1343 VTAIL.n279 VSUBS 0.028605f
C1344 VTAIL.n280 VSUBS 0.015371f
C1345 VTAIL.n281 VSUBS 0.036332f
C1346 VTAIL.n282 VSUBS 0.016275f
C1347 VTAIL.n283 VSUBS 1.89792f
C1348 VTAIL.n284 VSUBS 0.015371f
C1349 VTAIL.t0 VSUBS 0.077818f
C1350 VTAIL.n285 VSUBS 0.206282f
C1351 VTAIL.n286 VSUBS 0.023113f
C1352 VTAIL.n287 VSUBS 0.027249f
C1353 VTAIL.n288 VSUBS 0.036332f
C1354 VTAIL.n289 VSUBS 0.016275f
C1355 VTAIL.n290 VSUBS 0.015371f
C1356 VTAIL.n291 VSUBS 0.028605f
C1357 VTAIL.n292 VSUBS 0.028605f
C1358 VTAIL.n293 VSUBS 0.015371f
C1359 VTAIL.n294 VSUBS 0.016275f
C1360 VTAIL.n295 VSUBS 0.036332f
C1361 VTAIL.n296 VSUBS 0.036332f
C1362 VTAIL.n297 VSUBS 0.016275f
C1363 VTAIL.n298 VSUBS 0.015371f
C1364 VTAIL.n299 VSUBS 0.028605f
C1365 VTAIL.n300 VSUBS 0.028605f
C1366 VTAIL.n301 VSUBS 0.015371f
C1367 VTAIL.n302 VSUBS 0.016275f
C1368 VTAIL.n303 VSUBS 0.036332f
C1369 VTAIL.n304 VSUBS 0.036332f
C1370 VTAIL.n305 VSUBS 0.016275f
C1371 VTAIL.n306 VSUBS 0.015371f
C1372 VTAIL.n307 VSUBS 0.028605f
C1373 VTAIL.n308 VSUBS 0.028605f
C1374 VTAIL.n309 VSUBS 0.015371f
C1375 VTAIL.n310 VSUBS 0.016275f
C1376 VTAIL.n311 VSUBS 0.036332f
C1377 VTAIL.n312 VSUBS 0.036332f
C1378 VTAIL.n313 VSUBS 0.016275f
C1379 VTAIL.n314 VSUBS 0.015371f
C1380 VTAIL.n315 VSUBS 0.028605f
C1381 VTAIL.n316 VSUBS 0.028605f
C1382 VTAIL.n317 VSUBS 0.015371f
C1383 VTAIL.n318 VSUBS 0.016275f
C1384 VTAIL.n319 VSUBS 0.036332f
C1385 VTAIL.n320 VSUBS 0.036332f
C1386 VTAIL.n321 VSUBS 0.016275f
C1387 VTAIL.n322 VSUBS 0.015371f
C1388 VTAIL.n323 VSUBS 0.028605f
C1389 VTAIL.n324 VSUBS 0.028605f
C1390 VTAIL.n325 VSUBS 0.015371f
C1391 VTAIL.n326 VSUBS 0.015371f
C1392 VTAIL.n327 VSUBS 0.016275f
C1393 VTAIL.n328 VSUBS 0.036332f
C1394 VTAIL.n329 VSUBS 0.036332f
C1395 VTAIL.n330 VSUBS 0.036332f
C1396 VTAIL.n331 VSUBS 0.015823f
C1397 VTAIL.n332 VSUBS 0.015371f
C1398 VTAIL.n333 VSUBS 0.028605f
C1399 VTAIL.n334 VSUBS 0.028605f
C1400 VTAIL.n335 VSUBS 0.015371f
C1401 VTAIL.n336 VSUBS 0.016275f
C1402 VTAIL.n337 VSUBS 0.036332f
C1403 VTAIL.n338 VSUBS 0.088787f
C1404 VTAIL.n339 VSUBS 0.016275f
C1405 VTAIL.n340 VSUBS 0.015371f
C1406 VTAIL.n341 VSUBS 0.073544f
C1407 VTAIL.n342 VSUBS 0.044905f
C1408 VTAIL.n343 VSUBS 1.94142f
C1409 VP.t0 VSUBS 4.64333f
C1410 VP.t1 VSUBS 5.35002f
C1411 VP.n0 VSUBS 6.10837f
.ends

