* NGSPICE file created from diff_pair_sample_0139.ext - technology: sky130A

.subckt diff_pair_sample_0139 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2210_n4966# sky130_fd_pr__pfet_01v8 ad=7.7961 pd=40.76 as=0 ps=0 w=19.99 l=2.77
X1 VDD1.t1 VP.t0 VTAIL.t2 w_n2210_n4966# sky130_fd_pr__pfet_01v8 ad=7.7961 pd=40.76 as=7.7961 ps=40.76 w=19.99 l=2.77
X2 VDD1.t0 VP.t1 VTAIL.t3 w_n2210_n4966# sky130_fd_pr__pfet_01v8 ad=7.7961 pd=40.76 as=7.7961 ps=40.76 w=19.99 l=2.77
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n2210_n4966# sky130_fd_pr__pfet_01v8 ad=7.7961 pd=40.76 as=7.7961 ps=40.76 w=19.99 l=2.77
X4 VDD2.t0 VN.t1 VTAIL.t0 w_n2210_n4966# sky130_fd_pr__pfet_01v8 ad=7.7961 pd=40.76 as=7.7961 ps=40.76 w=19.99 l=2.77
X5 B.t8 B.t6 B.t7 w_n2210_n4966# sky130_fd_pr__pfet_01v8 ad=7.7961 pd=40.76 as=0 ps=0 w=19.99 l=2.77
X6 B.t5 B.t3 B.t4 w_n2210_n4966# sky130_fd_pr__pfet_01v8 ad=7.7961 pd=40.76 as=0 ps=0 w=19.99 l=2.77
X7 B.t2 B.t0 B.t1 w_n2210_n4966# sky130_fd_pr__pfet_01v8 ad=7.7961 pd=40.76 as=0 ps=0 w=19.99 l=2.77
R0 B.n452 B.n117 585
R1 B.n451 B.n450 585
R2 B.n449 B.n118 585
R3 B.n448 B.n447 585
R4 B.n446 B.n119 585
R5 B.n445 B.n444 585
R6 B.n443 B.n120 585
R7 B.n442 B.n441 585
R8 B.n440 B.n121 585
R9 B.n439 B.n438 585
R10 B.n437 B.n122 585
R11 B.n436 B.n435 585
R12 B.n434 B.n123 585
R13 B.n433 B.n432 585
R14 B.n431 B.n124 585
R15 B.n430 B.n429 585
R16 B.n428 B.n125 585
R17 B.n427 B.n426 585
R18 B.n425 B.n126 585
R19 B.n424 B.n423 585
R20 B.n422 B.n127 585
R21 B.n421 B.n420 585
R22 B.n419 B.n128 585
R23 B.n418 B.n417 585
R24 B.n416 B.n129 585
R25 B.n415 B.n414 585
R26 B.n413 B.n130 585
R27 B.n412 B.n411 585
R28 B.n410 B.n131 585
R29 B.n409 B.n408 585
R30 B.n407 B.n132 585
R31 B.n406 B.n405 585
R32 B.n404 B.n133 585
R33 B.n403 B.n402 585
R34 B.n401 B.n134 585
R35 B.n400 B.n399 585
R36 B.n398 B.n135 585
R37 B.n397 B.n396 585
R38 B.n395 B.n136 585
R39 B.n394 B.n393 585
R40 B.n392 B.n137 585
R41 B.n391 B.n390 585
R42 B.n389 B.n138 585
R43 B.n388 B.n387 585
R44 B.n386 B.n139 585
R45 B.n385 B.n384 585
R46 B.n383 B.n140 585
R47 B.n382 B.n381 585
R48 B.n380 B.n141 585
R49 B.n379 B.n378 585
R50 B.n377 B.n142 585
R51 B.n376 B.n375 585
R52 B.n374 B.n143 585
R53 B.n373 B.n372 585
R54 B.n371 B.n144 585
R55 B.n370 B.n369 585
R56 B.n368 B.n145 585
R57 B.n367 B.n366 585
R58 B.n365 B.n146 585
R59 B.n364 B.n363 585
R60 B.n362 B.n147 585
R61 B.n361 B.n360 585
R62 B.n359 B.n148 585
R63 B.n358 B.n357 585
R64 B.n356 B.n149 585
R65 B.n355 B.n354 585
R66 B.n350 B.n150 585
R67 B.n349 B.n348 585
R68 B.n347 B.n151 585
R69 B.n346 B.n345 585
R70 B.n344 B.n152 585
R71 B.n343 B.n342 585
R72 B.n341 B.n153 585
R73 B.n340 B.n339 585
R74 B.n338 B.n154 585
R75 B.n336 B.n335 585
R76 B.n334 B.n157 585
R77 B.n333 B.n332 585
R78 B.n331 B.n158 585
R79 B.n330 B.n329 585
R80 B.n328 B.n159 585
R81 B.n327 B.n326 585
R82 B.n325 B.n160 585
R83 B.n324 B.n323 585
R84 B.n322 B.n161 585
R85 B.n321 B.n320 585
R86 B.n319 B.n162 585
R87 B.n318 B.n317 585
R88 B.n316 B.n163 585
R89 B.n315 B.n314 585
R90 B.n313 B.n164 585
R91 B.n312 B.n311 585
R92 B.n310 B.n165 585
R93 B.n309 B.n308 585
R94 B.n307 B.n166 585
R95 B.n306 B.n305 585
R96 B.n304 B.n167 585
R97 B.n303 B.n302 585
R98 B.n301 B.n168 585
R99 B.n300 B.n299 585
R100 B.n298 B.n169 585
R101 B.n297 B.n296 585
R102 B.n295 B.n170 585
R103 B.n294 B.n293 585
R104 B.n292 B.n171 585
R105 B.n291 B.n290 585
R106 B.n289 B.n172 585
R107 B.n288 B.n287 585
R108 B.n286 B.n173 585
R109 B.n285 B.n284 585
R110 B.n283 B.n174 585
R111 B.n282 B.n281 585
R112 B.n280 B.n175 585
R113 B.n279 B.n278 585
R114 B.n277 B.n176 585
R115 B.n276 B.n275 585
R116 B.n274 B.n177 585
R117 B.n273 B.n272 585
R118 B.n271 B.n178 585
R119 B.n270 B.n269 585
R120 B.n268 B.n179 585
R121 B.n267 B.n266 585
R122 B.n265 B.n180 585
R123 B.n264 B.n263 585
R124 B.n262 B.n181 585
R125 B.n261 B.n260 585
R126 B.n259 B.n182 585
R127 B.n258 B.n257 585
R128 B.n256 B.n183 585
R129 B.n255 B.n254 585
R130 B.n253 B.n184 585
R131 B.n252 B.n251 585
R132 B.n250 B.n185 585
R133 B.n249 B.n248 585
R134 B.n247 B.n186 585
R135 B.n246 B.n245 585
R136 B.n244 B.n187 585
R137 B.n243 B.n242 585
R138 B.n241 B.n188 585
R139 B.n240 B.n239 585
R140 B.n454 B.n453 585
R141 B.n455 B.n116 585
R142 B.n457 B.n456 585
R143 B.n458 B.n115 585
R144 B.n460 B.n459 585
R145 B.n461 B.n114 585
R146 B.n463 B.n462 585
R147 B.n464 B.n113 585
R148 B.n466 B.n465 585
R149 B.n467 B.n112 585
R150 B.n469 B.n468 585
R151 B.n470 B.n111 585
R152 B.n472 B.n471 585
R153 B.n473 B.n110 585
R154 B.n475 B.n474 585
R155 B.n476 B.n109 585
R156 B.n478 B.n477 585
R157 B.n479 B.n108 585
R158 B.n481 B.n480 585
R159 B.n482 B.n107 585
R160 B.n484 B.n483 585
R161 B.n485 B.n106 585
R162 B.n487 B.n486 585
R163 B.n488 B.n105 585
R164 B.n490 B.n489 585
R165 B.n491 B.n104 585
R166 B.n493 B.n492 585
R167 B.n494 B.n103 585
R168 B.n496 B.n495 585
R169 B.n497 B.n102 585
R170 B.n499 B.n498 585
R171 B.n500 B.n101 585
R172 B.n502 B.n501 585
R173 B.n503 B.n100 585
R174 B.n505 B.n504 585
R175 B.n506 B.n99 585
R176 B.n508 B.n507 585
R177 B.n509 B.n98 585
R178 B.n511 B.n510 585
R179 B.n512 B.n97 585
R180 B.n514 B.n513 585
R181 B.n515 B.n96 585
R182 B.n517 B.n516 585
R183 B.n518 B.n95 585
R184 B.n520 B.n519 585
R185 B.n521 B.n94 585
R186 B.n523 B.n522 585
R187 B.n524 B.n93 585
R188 B.n526 B.n525 585
R189 B.n527 B.n92 585
R190 B.n529 B.n528 585
R191 B.n530 B.n91 585
R192 B.n532 B.n531 585
R193 B.n533 B.n90 585
R194 B.n744 B.n15 585
R195 B.n743 B.n742 585
R196 B.n741 B.n16 585
R197 B.n740 B.n739 585
R198 B.n738 B.n17 585
R199 B.n737 B.n736 585
R200 B.n735 B.n18 585
R201 B.n734 B.n733 585
R202 B.n732 B.n19 585
R203 B.n731 B.n730 585
R204 B.n729 B.n20 585
R205 B.n728 B.n727 585
R206 B.n726 B.n21 585
R207 B.n725 B.n724 585
R208 B.n723 B.n22 585
R209 B.n722 B.n721 585
R210 B.n720 B.n23 585
R211 B.n719 B.n718 585
R212 B.n717 B.n24 585
R213 B.n716 B.n715 585
R214 B.n714 B.n25 585
R215 B.n713 B.n712 585
R216 B.n711 B.n26 585
R217 B.n710 B.n709 585
R218 B.n708 B.n27 585
R219 B.n707 B.n706 585
R220 B.n705 B.n28 585
R221 B.n704 B.n703 585
R222 B.n702 B.n29 585
R223 B.n701 B.n700 585
R224 B.n699 B.n30 585
R225 B.n698 B.n697 585
R226 B.n696 B.n31 585
R227 B.n695 B.n694 585
R228 B.n693 B.n32 585
R229 B.n692 B.n691 585
R230 B.n690 B.n33 585
R231 B.n689 B.n688 585
R232 B.n687 B.n34 585
R233 B.n686 B.n685 585
R234 B.n684 B.n35 585
R235 B.n683 B.n682 585
R236 B.n681 B.n36 585
R237 B.n680 B.n679 585
R238 B.n678 B.n37 585
R239 B.n677 B.n676 585
R240 B.n675 B.n38 585
R241 B.n674 B.n673 585
R242 B.n672 B.n39 585
R243 B.n671 B.n670 585
R244 B.n669 B.n40 585
R245 B.n668 B.n667 585
R246 B.n666 B.n41 585
R247 B.n665 B.n664 585
R248 B.n663 B.n42 585
R249 B.n662 B.n661 585
R250 B.n660 B.n43 585
R251 B.n659 B.n658 585
R252 B.n657 B.n44 585
R253 B.n656 B.n655 585
R254 B.n654 B.n45 585
R255 B.n653 B.n652 585
R256 B.n651 B.n46 585
R257 B.n650 B.n649 585
R258 B.n648 B.n47 585
R259 B.n646 B.n645 585
R260 B.n644 B.n50 585
R261 B.n643 B.n642 585
R262 B.n641 B.n51 585
R263 B.n640 B.n639 585
R264 B.n638 B.n52 585
R265 B.n637 B.n636 585
R266 B.n635 B.n53 585
R267 B.n634 B.n633 585
R268 B.n632 B.n54 585
R269 B.n631 B.n630 585
R270 B.n629 B.n55 585
R271 B.n628 B.n627 585
R272 B.n626 B.n59 585
R273 B.n625 B.n624 585
R274 B.n623 B.n60 585
R275 B.n622 B.n621 585
R276 B.n620 B.n61 585
R277 B.n619 B.n618 585
R278 B.n617 B.n62 585
R279 B.n616 B.n615 585
R280 B.n614 B.n63 585
R281 B.n613 B.n612 585
R282 B.n611 B.n64 585
R283 B.n610 B.n609 585
R284 B.n608 B.n65 585
R285 B.n607 B.n606 585
R286 B.n605 B.n66 585
R287 B.n604 B.n603 585
R288 B.n602 B.n67 585
R289 B.n601 B.n600 585
R290 B.n599 B.n68 585
R291 B.n598 B.n597 585
R292 B.n596 B.n69 585
R293 B.n595 B.n594 585
R294 B.n593 B.n70 585
R295 B.n592 B.n591 585
R296 B.n590 B.n71 585
R297 B.n589 B.n588 585
R298 B.n587 B.n72 585
R299 B.n586 B.n585 585
R300 B.n584 B.n73 585
R301 B.n583 B.n582 585
R302 B.n581 B.n74 585
R303 B.n580 B.n579 585
R304 B.n578 B.n75 585
R305 B.n577 B.n576 585
R306 B.n575 B.n76 585
R307 B.n574 B.n573 585
R308 B.n572 B.n77 585
R309 B.n571 B.n570 585
R310 B.n569 B.n78 585
R311 B.n568 B.n567 585
R312 B.n566 B.n79 585
R313 B.n565 B.n564 585
R314 B.n563 B.n80 585
R315 B.n562 B.n561 585
R316 B.n560 B.n81 585
R317 B.n559 B.n558 585
R318 B.n557 B.n82 585
R319 B.n556 B.n555 585
R320 B.n554 B.n83 585
R321 B.n553 B.n552 585
R322 B.n551 B.n84 585
R323 B.n550 B.n549 585
R324 B.n548 B.n85 585
R325 B.n547 B.n546 585
R326 B.n545 B.n86 585
R327 B.n544 B.n543 585
R328 B.n542 B.n87 585
R329 B.n541 B.n540 585
R330 B.n539 B.n88 585
R331 B.n538 B.n537 585
R332 B.n536 B.n89 585
R333 B.n535 B.n534 585
R334 B.n746 B.n745 585
R335 B.n747 B.n14 585
R336 B.n749 B.n748 585
R337 B.n750 B.n13 585
R338 B.n752 B.n751 585
R339 B.n753 B.n12 585
R340 B.n755 B.n754 585
R341 B.n756 B.n11 585
R342 B.n758 B.n757 585
R343 B.n759 B.n10 585
R344 B.n761 B.n760 585
R345 B.n762 B.n9 585
R346 B.n764 B.n763 585
R347 B.n765 B.n8 585
R348 B.n767 B.n766 585
R349 B.n768 B.n7 585
R350 B.n770 B.n769 585
R351 B.n771 B.n6 585
R352 B.n773 B.n772 585
R353 B.n774 B.n5 585
R354 B.n776 B.n775 585
R355 B.n777 B.n4 585
R356 B.n779 B.n778 585
R357 B.n780 B.n3 585
R358 B.n782 B.n781 585
R359 B.n783 B.n0 585
R360 B.n2 B.n1 585
R361 B.n202 B.n201 585
R362 B.n204 B.n203 585
R363 B.n205 B.n200 585
R364 B.n207 B.n206 585
R365 B.n208 B.n199 585
R366 B.n210 B.n209 585
R367 B.n211 B.n198 585
R368 B.n213 B.n212 585
R369 B.n214 B.n197 585
R370 B.n216 B.n215 585
R371 B.n217 B.n196 585
R372 B.n219 B.n218 585
R373 B.n220 B.n195 585
R374 B.n222 B.n221 585
R375 B.n223 B.n194 585
R376 B.n225 B.n224 585
R377 B.n226 B.n193 585
R378 B.n228 B.n227 585
R379 B.n229 B.n192 585
R380 B.n231 B.n230 585
R381 B.n232 B.n191 585
R382 B.n234 B.n233 585
R383 B.n235 B.n190 585
R384 B.n237 B.n236 585
R385 B.n238 B.n189 585
R386 B.n239 B.n238 458.866
R387 B.n453 B.n452 458.866
R388 B.n535 B.n90 458.866
R389 B.n746 B.n15 458.866
R390 B.n155 B.t6 382.211
R391 B.n351 B.t0 382.211
R392 B.n56 B.t9 382.211
R393 B.n48 B.t3 382.211
R394 B.n785 B.n784 256.663
R395 B.n784 B.n783 235.042
R396 B.n784 B.n2 235.042
R397 B.n351 B.t1 171.385
R398 B.n56 B.t11 171.385
R399 B.n155 B.t7 171.358
R400 B.n48 B.t5 171.358
R401 B.n239 B.n188 163.367
R402 B.n243 B.n188 163.367
R403 B.n244 B.n243 163.367
R404 B.n245 B.n244 163.367
R405 B.n245 B.n186 163.367
R406 B.n249 B.n186 163.367
R407 B.n250 B.n249 163.367
R408 B.n251 B.n250 163.367
R409 B.n251 B.n184 163.367
R410 B.n255 B.n184 163.367
R411 B.n256 B.n255 163.367
R412 B.n257 B.n256 163.367
R413 B.n257 B.n182 163.367
R414 B.n261 B.n182 163.367
R415 B.n262 B.n261 163.367
R416 B.n263 B.n262 163.367
R417 B.n263 B.n180 163.367
R418 B.n267 B.n180 163.367
R419 B.n268 B.n267 163.367
R420 B.n269 B.n268 163.367
R421 B.n269 B.n178 163.367
R422 B.n273 B.n178 163.367
R423 B.n274 B.n273 163.367
R424 B.n275 B.n274 163.367
R425 B.n275 B.n176 163.367
R426 B.n279 B.n176 163.367
R427 B.n280 B.n279 163.367
R428 B.n281 B.n280 163.367
R429 B.n281 B.n174 163.367
R430 B.n285 B.n174 163.367
R431 B.n286 B.n285 163.367
R432 B.n287 B.n286 163.367
R433 B.n287 B.n172 163.367
R434 B.n291 B.n172 163.367
R435 B.n292 B.n291 163.367
R436 B.n293 B.n292 163.367
R437 B.n293 B.n170 163.367
R438 B.n297 B.n170 163.367
R439 B.n298 B.n297 163.367
R440 B.n299 B.n298 163.367
R441 B.n299 B.n168 163.367
R442 B.n303 B.n168 163.367
R443 B.n304 B.n303 163.367
R444 B.n305 B.n304 163.367
R445 B.n305 B.n166 163.367
R446 B.n309 B.n166 163.367
R447 B.n310 B.n309 163.367
R448 B.n311 B.n310 163.367
R449 B.n311 B.n164 163.367
R450 B.n315 B.n164 163.367
R451 B.n316 B.n315 163.367
R452 B.n317 B.n316 163.367
R453 B.n317 B.n162 163.367
R454 B.n321 B.n162 163.367
R455 B.n322 B.n321 163.367
R456 B.n323 B.n322 163.367
R457 B.n323 B.n160 163.367
R458 B.n327 B.n160 163.367
R459 B.n328 B.n327 163.367
R460 B.n329 B.n328 163.367
R461 B.n329 B.n158 163.367
R462 B.n333 B.n158 163.367
R463 B.n334 B.n333 163.367
R464 B.n335 B.n334 163.367
R465 B.n335 B.n154 163.367
R466 B.n340 B.n154 163.367
R467 B.n341 B.n340 163.367
R468 B.n342 B.n341 163.367
R469 B.n342 B.n152 163.367
R470 B.n346 B.n152 163.367
R471 B.n347 B.n346 163.367
R472 B.n348 B.n347 163.367
R473 B.n348 B.n150 163.367
R474 B.n355 B.n150 163.367
R475 B.n356 B.n355 163.367
R476 B.n357 B.n356 163.367
R477 B.n357 B.n148 163.367
R478 B.n361 B.n148 163.367
R479 B.n362 B.n361 163.367
R480 B.n363 B.n362 163.367
R481 B.n363 B.n146 163.367
R482 B.n367 B.n146 163.367
R483 B.n368 B.n367 163.367
R484 B.n369 B.n368 163.367
R485 B.n369 B.n144 163.367
R486 B.n373 B.n144 163.367
R487 B.n374 B.n373 163.367
R488 B.n375 B.n374 163.367
R489 B.n375 B.n142 163.367
R490 B.n379 B.n142 163.367
R491 B.n380 B.n379 163.367
R492 B.n381 B.n380 163.367
R493 B.n381 B.n140 163.367
R494 B.n385 B.n140 163.367
R495 B.n386 B.n385 163.367
R496 B.n387 B.n386 163.367
R497 B.n387 B.n138 163.367
R498 B.n391 B.n138 163.367
R499 B.n392 B.n391 163.367
R500 B.n393 B.n392 163.367
R501 B.n393 B.n136 163.367
R502 B.n397 B.n136 163.367
R503 B.n398 B.n397 163.367
R504 B.n399 B.n398 163.367
R505 B.n399 B.n134 163.367
R506 B.n403 B.n134 163.367
R507 B.n404 B.n403 163.367
R508 B.n405 B.n404 163.367
R509 B.n405 B.n132 163.367
R510 B.n409 B.n132 163.367
R511 B.n410 B.n409 163.367
R512 B.n411 B.n410 163.367
R513 B.n411 B.n130 163.367
R514 B.n415 B.n130 163.367
R515 B.n416 B.n415 163.367
R516 B.n417 B.n416 163.367
R517 B.n417 B.n128 163.367
R518 B.n421 B.n128 163.367
R519 B.n422 B.n421 163.367
R520 B.n423 B.n422 163.367
R521 B.n423 B.n126 163.367
R522 B.n427 B.n126 163.367
R523 B.n428 B.n427 163.367
R524 B.n429 B.n428 163.367
R525 B.n429 B.n124 163.367
R526 B.n433 B.n124 163.367
R527 B.n434 B.n433 163.367
R528 B.n435 B.n434 163.367
R529 B.n435 B.n122 163.367
R530 B.n439 B.n122 163.367
R531 B.n440 B.n439 163.367
R532 B.n441 B.n440 163.367
R533 B.n441 B.n120 163.367
R534 B.n445 B.n120 163.367
R535 B.n446 B.n445 163.367
R536 B.n447 B.n446 163.367
R537 B.n447 B.n118 163.367
R538 B.n451 B.n118 163.367
R539 B.n452 B.n451 163.367
R540 B.n531 B.n90 163.367
R541 B.n531 B.n530 163.367
R542 B.n530 B.n529 163.367
R543 B.n529 B.n92 163.367
R544 B.n525 B.n92 163.367
R545 B.n525 B.n524 163.367
R546 B.n524 B.n523 163.367
R547 B.n523 B.n94 163.367
R548 B.n519 B.n94 163.367
R549 B.n519 B.n518 163.367
R550 B.n518 B.n517 163.367
R551 B.n517 B.n96 163.367
R552 B.n513 B.n96 163.367
R553 B.n513 B.n512 163.367
R554 B.n512 B.n511 163.367
R555 B.n511 B.n98 163.367
R556 B.n507 B.n98 163.367
R557 B.n507 B.n506 163.367
R558 B.n506 B.n505 163.367
R559 B.n505 B.n100 163.367
R560 B.n501 B.n100 163.367
R561 B.n501 B.n500 163.367
R562 B.n500 B.n499 163.367
R563 B.n499 B.n102 163.367
R564 B.n495 B.n102 163.367
R565 B.n495 B.n494 163.367
R566 B.n494 B.n493 163.367
R567 B.n493 B.n104 163.367
R568 B.n489 B.n104 163.367
R569 B.n489 B.n488 163.367
R570 B.n488 B.n487 163.367
R571 B.n487 B.n106 163.367
R572 B.n483 B.n106 163.367
R573 B.n483 B.n482 163.367
R574 B.n482 B.n481 163.367
R575 B.n481 B.n108 163.367
R576 B.n477 B.n108 163.367
R577 B.n477 B.n476 163.367
R578 B.n476 B.n475 163.367
R579 B.n475 B.n110 163.367
R580 B.n471 B.n110 163.367
R581 B.n471 B.n470 163.367
R582 B.n470 B.n469 163.367
R583 B.n469 B.n112 163.367
R584 B.n465 B.n112 163.367
R585 B.n465 B.n464 163.367
R586 B.n464 B.n463 163.367
R587 B.n463 B.n114 163.367
R588 B.n459 B.n114 163.367
R589 B.n459 B.n458 163.367
R590 B.n458 B.n457 163.367
R591 B.n457 B.n116 163.367
R592 B.n453 B.n116 163.367
R593 B.n742 B.n15 163.367
R594 B.n742 B.n741 163.367
R595 B.n741 B.n740 163.367
R596 B.n740 B.n17 163.367
R597 B.n736 B.n17 163.367
R598 B.n736 B.n735 163.367
R599 B.n735 B.n734 163.367
R600 B.n734 B.n19 163.367
R601 B.n730 B.n19 163.367
R602 B.n730 B.n729 163.367
R603 B.n729 B.n728 163.367
R604 B.n728 B.n21 163.367
R605 B.n724 B.n21 163.367
R606 B.n724 B.n723 163.367
R607 B.n723 B.n722 163.367
R608 B.n722 B.n23 163.367
R609 B.n718 B.n23 163.367
R610 B.n718 B.n717 163.367
R611 B.n717 B.n716 163.367
R612 B.n716 B.n25 163.367
R613 B.n712 B.n25 163.367
R614 B.n712 B.n711 163.367
R615 B.n711 B.n710 163.367
R616 B.n710 B.n27 163.367
R617 B.n706 B.n27 163.367
R618 B.n706 B.n705 163.367
R619 B.n705 B.n704 163.367
R620 B.n704 B.n29 163.367
R621 B.n700 B.n29 163.367
R622 B.n700 B.n699 163.367
R623 B.n699 B.n698 163.367
R624 B.n698 B.n31 163.367
R625 B.n694 B.n31 163.367
R626 B.n694 B.n693 163.367
R627 B.n693 B.n692 163.367
R628 B.n692 B.n33 163.367
R629 B.n688 B.n33 163.367
R630 B.n688 B.n687 163.367
R631 B.n687 B.n686 163.367
R632 B.n686 B.n35 163.367
R633 B.n682 B.n35 163.367
R634 B.n682 B.n681 163.367
R635 B.n681 B.n680 163.367
R636 B.n680 B.n37 163.367
R637 B.n676 B.n37 163.367
R638 B.n676 B.n675 163.367
R639 B.n675 B.n674 163.367
R640 B.n674 B.n39 163.367
R641 B.n670 B.n39 163.367
R642 B.n670 B.n669 163.367
R643 B.n669 B.n668 163.367
R644 B.n668 B.n41 163.367
R645 B.n664 B.n41 163.367
R646 B.n664 B.n663 163.367
R647 B.n663 B.n662 163.367
R648 B.n662 B.n43 163.367
R649 B.n658 B.n43 163.367
R650 B.n658 B.n657 163.367
R651 B.n657 B.n656 163.367
R652 B.n656 B.n45 163.367
R653 B.n652 B.n45 163.367
R654 B.n652 B.n651 163.367
R655 B.n651 B.n650 163.367
R656 B.n650 B.n47 163.367
R657 B.n645 B.n47 163.367
R658 B.n645 B.n644 163.367
R659 B.n644 B.n643 163.367
R660 B.n643 B.n51 163.367
R661 B.n639 B.n51 163.367
R662 B.n639 B.n638 163.367
R663 B.n638 B.n637 163.367
R664 B.n637 B.n53 163.367
R665 B.n633 B.n53 163.367
R666 B.n633 B.n632 163.367
R667 B.n632 B.n631 163.367
R668 B.n631 B.n55 163.367
R669 B.n627 B.n55 163.367
R670 B.n627 B.n626 163.367
R671 B.n626 B.n625 163.367
R672 B.n625 B.n60 163.367
R673 B.n621 B.n60 163.367
R674 B.n621 B.n620 163.367
R675 B.n620 B.n619 163.367
R676 B.n619 B.n62 163.367
R677 B.n615 B.n62 163.367
R678 B.n615 B.n614 163.367
R679 B.n614 B.n613 163.367
R680 B.n613 B.n64 163.367
R681 B.n609 B.n64 163.367
R682 B.n609 B.n608 163.367
R683 B.n608 B.n607 163.367
R684 B.n607 B.n66 163.367
R685 B.n603 B.n66 163.367
R686 B.n603 B.n602 163.367
R687 B.n602 B.n601 163.367
R688 B.n601 B.n68 163.367
R689 B.n597 B.n68 163.367
R690 B.n597 B.n596 163.367
R691 B.n596 B.n595 163.367
R692 B.n595 B.n70 163.367
R693 B.n591 B.n70 163.367
R694 B.n591 B.n590 163.367
R695 B.n590 B.n589 163.367
R696 B.n589 B.n72 163.367
R697 B.n585 B.n72 163.367
R698 B.n585 B.n584 163.367
R699 B.n584 B.n583 163.367
R700 B.n583 B.n74 163.367
R701 B.n579 B.n74 163.367
R702 B.n579 B.n578 163.367
R703 B.n578 B.n577 163.367
R704 B.n577 B.n76 163.367
R705 B.n573 B.n76 163.367
R706 B.n573 B.n572 163.367
R707 B.n572 B.n571 163.367
R708 B.n571 B.n78 163.367
R709 B.n567 B.n78 163.367
R710 B.n567 B.n566 163.367
R711 B.n566 B.n565 163.367
R712 B.n565 B.n80 163.367
R713 B.n561 B.n80 163.367
R714 B.n561 B.n560 163.367
R715 B.n560 B.n559 163.367
R716 B.n559 B.n82 163.367
R717 B.n555 B.n82 163.367
R718 B.n555 B.n554 163.367
R719 B.n554 B.n553 163.367
R720 B.n553 B.n84 163.367
R721 B.n549 B.n84 163.367
R722 B.n549 B.n548 163.367
R723 B.n548 B.n547 163.367
R724 B.n547 B.n86 163.367
R725 B.n543 B.n86 163.367
R726 B.n543 B.n542 163.367
R727 B.n542 B.n541 163.367
R728 B.n541 B.n88 163.367
R729 B.n537 B.n88 163.367
R730 B.n537 B.n536 163.367
R731 B.n536 B.n535 163.367
R732 B.n747 B.n746 163.367
R733 B.n748 B.n747 163.367
R734 B.n748 B.n13 163.367
R735 B.n752 B.n13 163.367
R736 B.n753 B.n752 163.367
R737 B.n754 B.n753 163.367
R738 B.n754 B.n11 163.367
R739 B.n758 B.n11 163.367
R740 B.n759 B.n758 163.367
R741 B.n760 B.n759 163.367
R742 B.n760 B.n9 163.367
R743 B.n764 B.n9 163.367
R744 B.n765 B.n764 163.367
R745 B.n766 B.n765 163.367
R746 B.n766 B.n7 163.367
R747 B.n770 B.n7 163.367
R748 B.n771 B.n770 163.367
R749 B.n772 B.n771 163.367
R750 B.n772 B.n5 163.367
R751 B.n776 B.n5 163.367
R752 B.n777 B.n776 163.367
R753 B.n778 B.n777 163.367
R754 B.n778 B.n3 163.367
R755 B.n782 B.n3 163.367
R756 B.n783 B.n782 163.367
R757 B.n202 B.n2 163.367
R758 B.n203 B.n202 163.367
R759 B.n203 B.n200 163.367
R760 B.n207 B.n200 163.367
R761 B.n208 B.n207 163.367
R762 B.n209 B.n208 163.367
R763 B.n209 B.n198 163.367
R764 B.n213 B.n198 163.367
R765 B.n214 B.n213 163.367
R766 B.n215 B.n214 163.367
R767 B.n215 B.n196 163.367
R768 B.n219 B.n196 163.367
R769 B.n220 B.n219 163.367
R770 B.n221 B.n220 163.367
R771 B.n221 B.n194 163.367
R772 B.n225 B.n194 163.367
R773 B.n226 B.n225 163.367
R774 B.n227 B.n226 163.367
R775 B.n227 B.n192 163.367
R776 B.n231 B.n192 163.367
R777 B.n232 B.n231 163.367
R778 B.n233 B.n232 163.367
R779 B.n233 B.n190 163.367
R780 B.n237 B.n190 163.367
R781 B.n238 B.n237 163.367
R782 B.n352 B.t2 111.263
R783 B.n57 B.t10 111.263
R784 B.n156 B.t8 111.237
R785 B.n49 B.t4 111.237
R786 B.n156 B.n155 60.1217
R787 B.n352 B.n351 60.1217
R788 B.n57 B.n56 60.1217
R789 B.n49 B.n48 60.1217
R790 B.n337 B.n156 59.5399
R791 B.n353 B.n352 59.5399
R792 B.n58 B.n57 59.5399
R793 B.n647 B.n49 59.5399
R794 B.n745 B.n744 29.8151
R795 B.n534 B.n533 29.8151
R796 B.n454 B.n117 29.8151
R797 B.n240 B.n189 29.8151
R798 B B.n785 18.0485
R799 B.n745 B.n14 10.6151
R800 B.n749 B.n14 10.6151
R801 B.n750 B.n749 10.6151
R802 B.n751 B.n750 10.6151
R803 B.n751 B.n12 10.6151
R804 B.n755 B.n12 10.6151
R805 B.n756 B.n755 10.6151
R806 B.n757 B.n756 10.6151
R807 B.n757 B.n10 10.6151
R808 B.n761 B.n10 10.6151
R809 B.n762 B.n761 10.6151
R810 B.n763 B.n762 10.6151
R811 B.n763 B.n8 10.6151
R812 B.n767 B.n8 10.6151
R813 B.n768 B.n767 10.6151
R814 B.n769 B.n768 10.6151
R815 B.n769 B.n6 10.6151
R816 B.n773 B.n6 10.6151
R817 B.n774 B.n773 10.6151
R818 B.n775 B.n774 10.6151
R819 B.n775 B.n4 10.6151
R820 B.n779 B.n4 10.6151
R821 B.n780 B.n779 10.6151
R822 B.n781 B.n780 10.6151
R823 B.n781 B.n0 10.6151
R824 B.n744 B.n743 10.6151
R825 B.n743 B.n16 10.6151
R826 B.n739 B.n16 10.6151
R827 B.n739 B.n738 10.6151
R828 B.n738 B.n737 10.6151
R829 B.n737 B.n18 10.6151
R830 B.n733 B.n18 10.6151
R831 B.n733 B.n732 10.6151
R832 B.n732 B.n731 10.6151
R833 B.n731 B.n20 10.6151
R834 B.n727 B.n20 10.6151
R835 B.n727 B.n726 10.6151
R836 B.n726 B.n725 10.6151
R837 B.n725 B.n22 10.6151
R838 B.n721 B.n22 10.6151
R839 B.n721 B.n720 10.6151
R840 B.n720 B.n719 10.6151
R841 B.n719 B.n24 10.6151
R842 B.n715 B.n24 10.6151
R843 B.n715 B.n714 10.6151
R844 B.n714 B.n713 10.6151
R845 B.n713 B.n26 10.6151
R846 B.n709 B.n26 10.6151
R847 B.n709 B.n708 10.6151
R848 B.n708 B.n707 10.6151
R849 B.n707 B.n28 10.6151
R850 B.n703 B.n28 10.6151
R851 B.n703 B.n702 10.6151
R852 B.n702 B.n701 10.6151
R853 B.n701 B.n30 10.6151
R854 B.n697 B.n30 10.6151
R855 B.n697 B.n696 10.6151
R856 B.n696 B.n695 10.6151
R857 B.n695 B.n32 10.6151
R858 B.n691 B.n32 10.6151
R859 B.n691 B.n690 10.6151
R860 B.n690 B.n689 10.6151
R861 B.n689 B.n34 10.6151
R862 B.n685 B.n34 10.6151
R863 B.n685 B.n684 10.6151
R864 B.n684 B.n683 10.6151
R865 B.n683 B.n36 10.6151
R866 B.n679 B.n36 10.6151
R867 B.n679 B.n678 10.6151
R868 B.n678 B.n677 10.6151
R869 B.n677 B.n38 10.6151
R870 B.n673 B.n38 10.6151
R871 B.n673 B.n672 10.6151
R872 B.n672 B.n671 10.6151
R873 B.n671 B.n40 10.6151
R874 B.n667 B.n40 10.6151
R875 B.n667 B.n666 10.6151
R876 B.n666 B.n665 10.6151
R877 B.n665 B.n42 10.6151
R878 B.n661 B.n42 10.6151
R879 B.n661 B.n660 10.6151
R880 B.n660 B.n659 10.6151
R881 B.n659 B.n44 10.6151
R882 B.n655 B.n44 10.6151
R883 B.n655 B.n654 10.6151
R884 B.n654 B.n653 10.6151
R885 B.n653 B.n46 10.6151
R886 B.n649 B.n46 10.6151
R887 B.n649 B.n648 10.6151
R888 B.n646 B.n50 10.6151
R889 B.n642 B.n50 10.6151
R890 B.n642 B.n641 10.6151
R891 B.n641 B.n640 10.6151
R892 B.n640 B.n52 10.6151
R893 B.n636 B.n52 10.6151
R894 B.n636 B.n635 10.6151
R895 B.n635 B.n634 10.6151
R896 B.n634 B.n54 10.6151
R897 B.n630 B.n629 10.6151
R898 B.n629 B.n628 10.6151
R899 B.n628 B.n59 10.6151
R900 B.n624 B.n59 10.6151
R901 B.n624 B.n623 10.6151
R902 B.n623 B.n622 10.6151
R903 B.n622 B.n61 10.6151
R904 B.n618 B.n61 10.6151
R905 B.n618 B.n617 10.6151
R906 B.n617 B.n616 10.6151
R907 B.n616 B.n63 10.6151
R908 B.n612 B.n63 10.6151
R909 B.n612 B.n611 10.6151
R910 B.n611 B.n610 10.6151
R911 B.n610 B.n65 10.6151
R912 B.n606 B.n65 10.6151
R913 B.n606 B.n605 10.6151
R914 B.n605 B.n604 10.6151
R915 B.n604 B.n67 10.6151
R916 B.n600 B.n67 10.6151
R917 B.n600 B.n599 10.6151
R918 B.n599 B.n598 10.6151
R919 B.n598 B.n69 10.6151
R920 B.n594 B.n69 10.6151
R921 B.n594 B.n593 10.6151
R922 B.n593 B.n592 10.6151
R923 B.n592 B.n71 10.6151
R924 B.n588 B.n71 10.6151
R925 B.n588 B.n587 10.6151
R926 B.n587 B.n586 10.6151
R927 B.n586 B.n73 10.6151
R928 B.n582 B.n73 10.6151
R929 B.n582 B.n581 10.6151
R930 B.n581 B.n580 10.6151
R931 B.n580 B.n75 10.6151
R932 B.n576 B.n75 10.6151
R933 B.n576 B.n575 10.6151
R934 B.n575 B.n574 10.6151
R935 B.n574 B.n77 10.6151
R936 B.n570 B.n77 10.6151
R937 B.n570 B.n569 10.6151
R938 B.n569 B.n568 10.6151
R939 B.n568 B.n79 10.6151
R940 B.n564 B.n79 10.6151
R941 B.n564 B.n563 10.6151
R942 B.n563 B.n562 10.6151
R943 B.n562 B.n81 10.6151
R944 B.n558 B.n81 10.6151
R945 B.n558 B.n557 10.6151
R946 B.n557 B.n556 10.6151
R947 B.n556 B.n83 10.6151
R948 B.n552 B.n83 10.6151
R949 B.n552 B.n551 10.6151
R950 B.n551 B.n550 10.6151
R951 B.n550 B.n85 10.6151
R952 B.n546 B.n85 10.6151
R953 B.n546 B.n545 10.6151
R954 B.n545 B.n544 10.6151
R955 B.n544 B.n87 10.6151
R956 B.n540 B.n87 10.6151
R957 B.n540 B.n539 10.6151
R958 B.n539 B.n538 10.6151
R959 B.n538 B.n89 10.6151
R960 B.n534 B.n89 10.6151
R961 B.n533 B.n532 10.6151
R962 B.n532 B.n91 10.6151
R963 B.n528 B.n91 10.6151
R964 B.n528 B.n527 10.6151
R965 B.n527 B.n526 10.6151
R966 B.n526 B.n93 10.6151
R967 B.n522 B.n93 10.6151
R968 B.n522 B.n521 10.6151
R969 B.n521 B.n520 10.6151
R970 B.n520 B.n95 10.6151
R971 B.n516 B.n95 10.6151
R972 B.n516 B.n515 10.6151
R973 B.n515 B.n514 10.6151
R974 B.n514 B.n97 10.6151
R975 B.n510 B.n97 10.6151
R976 B.n510 B.n509 10.6151
R977 B.n509 B.n508 10.6151
R978 B.n508 B.n99 10.6151
R979 B.n504 B.n99 10.6151
R980 B.n504 B.n503 10.6151
R981 B.n503 B.n502 10.6151
R982 B.n502 B.n101 10.6151
R983 B.n498 B.n101 10.6151
R984 B.n498 B.n497 10.6151
R985 B.n497 B.n496 10.6151
R986 B.n496 B.n103 10.6151
R987 B.n492 B.n103 10.6151
R988 B.n492 B.n491 10.6151
R989 B.n491 B.n490 10.6151
R990 B.n490 B.n105 10.6151
R991 B.n486 B.n105 10.6151
R992 B.n486 B.n485 10.6151
R993 B.n485 B.n484 10.6151
R994 B.n484 B.n107 10.6151
R995 B.n480 B.n107 10.6151
R996 B.n480 B.n479 10.6151
R997 B.n479 B.n478 10.6151
R998 B.n478 B.n109 10.6151
R999 B.n474 B.n109 10.6151
R1000 B.n474 B.n473 10.6151
R1001 B.n473 B.n472 10.6151
R1002 B.n472 B.n111 10.6151
R1003 B.n468 B.n111 10.6151
R1004 B.n468 B.n467 10.6151
R1005 B.n467 B.n466 10.6151
R1006 B.n466 B.n113 10.6151
R1007 B.n462 B.n113 10.6151
R1008 B.n462 B.n461 10.6151
R1009 B.n461 B.n460 10.6151
R1010 B.n460 B.n115 10.6151
R1011 B.n456 B.n115 10.6151
R1012 B.n456 B.n455 10.6151
R1013 B.n455 B.n454 10.6151
R1014 B.n201 B.n1 10.6151
R1015 B.n204 B.n201 10.6151
R1016 B.n205 B.n204 10.6151
R1017 B.n206 B.n205 10.6151
R1018 B.n206 B.n199 10.6151
R1019 B.n210 B.n199 10.6151
R1020 B.n211 B.n210 10.6151
R1021 B.n212 B.n211 10.6151
R1022 B.n212 B.n197 10.6151
R1023 B.n216 B.n197 10.6151
R1024 B.n217 B.n216 10.6151
R1025 B.n218 B.n217 10.6151
R1026 B.n218 B.n195 10.6151
R1027 B.n222 B.n195 10.6151
R1028 B.n223 B.n222 10.6151
R1029 B.n224 B.n223 10.6151
R1030 B.n224 B.n193 10.6151
R1031 B.n228 B.n193 10.6151
R1032 B.n229 B.n228 10.6151
R1033 B.n230 B.n229 10.6151
R1034 B.n230 B.n191 10.6151
R1035 B.n234 B.n191 10.6151
R1036 B.n235 B.n234 10.6151
R1037 B.n236 B.n235 10.6151
R1038 B.n236 B.n189 10.6151
R1039 B.n241 B.n240 10.6151
R1040 B.n242 B.n241 10.6151
R1041 B.n242 B.n187 10.6151
R1042 B.n246 B.n187 10.6151
R1043 B.n247 B.n246 10.6151
R1044 B.n248 B.n247 10.6151
R1045 B.n248 B.n185 10.6151
R1046 B.n252 B.n185 10.6151
R1047 B.n253 B.n252 10.6151
R1048 B.n254 B.n253 10.6151
R1049 B.n254 B.n183 10.6151
R1050 B.n258 B.n183 10.6151
R1051 B.n259 B.n258 10.6151
R1052 B.n260 B.n259 10.6151
R1053 B.n260 B.n181 10.6151
R1054 B.n264 B.n181 10.6151
R1055 B.n265 B.n264 10.6151
R1056 B.n266 B.n265 10.6151
R1057 B.n266 B.n179 10.6151
R1058 B.n270 B.n179 10.6151
R1059 B.n271 B.n270 10.6151
R1060 B.n272 B.n271 10.6151
R1061 B.n272 B.n177 10.6151
R1062 B.n276 B.n177 10.6151
R1063 B.n277 B.n276 10.6151
R1064 B.n278 B.n277 10.6151
R1065 B.n278 B.n175 10.6151
R1066 B.n282 B.n175 10.6151
R1067 B.n283 B.n282 10.6151
R1068 B.n284 B.n283 10.6151
R1069 B.n284 B.n173 10.6151
R1070 B.n288 B.n173 10.6151
R1071 B.n289 B.n288 10.6151
R1072 B.n290 B.n289 10.6151
R1073 B.n290 B.n171 10.6151
R1074 B.n294 B.n171 10.6151
R1075 B.n295 B.n294 10.6151
R1076 B.n296 B.n295 10.6151
R1077 B.n296 B.n169 10.6151
R1078 B.n300 B.n169 10.6151
R1079 B.n301 B.n300 10.6151
R1080 B.n302 B.n301 10.6151
R1081 B.n302 B.n167 10.6151
R1082 B.n306 B.n167 10.6151
R1083 B.n307 B.n306 10.6151
R1084 B.n308 B.n307 10.6151
R1085 B.n308 B.n165 10.6151
R1086 B.n312 B.n165 10.6151
R1087 B.n313 B.n312 10.6151
R1088 B.n314 B.n313 10.6151
R1089 B.n314 B.n163 10.6151
R1090 B.n318 B.n163 10.6151
R1091 B.n319 B.n318 10.6151
R1092 B.n320 B.n319 10.6151
R1093 B.n320 B.n161 10.6151
R1094 B.n324 B.n161 10.6151
R1095 B.n325 B.n324 10.6151
R1096 B.n326 B.n325 10.6151
R1097 B.n326 B.n159 10.6151
R1098 B.n330 B.n159 10.6151
R1099 B.n331 B.n330 10.6151
R1100 B.n332 B.n331 10.6151
R1101 B.n332 B.n157 10.6151
R1102 B.n336 B.n157 10.6151
R1103 B.n339 B.n338 10.6151
R1104 B.n339 B.n153 10.6151
R1105 B.n343 B.n153 10.6151
R1106 B.n344 B.n343 10.6151
R1107 B.n345 B.n344 10.6151
R1108 B.n345 B.n151 10.6151
R1109 B.n349 B.n151 10.6151
R1110 B.n350 B.n349 10.6151
R1111 B.n354 B.n350 10.6151
R1112 B.n358 B.n149 10.6151
R1113 B.n359 B.n358 10.6151
R1114 B.n360 B.n359 10.6151
R1115 B.n360 B.n147 10.6151
R1116 B.n364 B.n147 10.6151
R1117 B.n365 B.n364 10.6151
R1118 B.n366 B.n365 10.6151
R1119 B.n366 B.n145 10.6151
R1120 B.n370 B.n145 10.6151
R1121 B.n371 B.n370 10.6151
R1122 B.n372 B.n371 10.6151
R1123 B.n372 B.n143 10.6151
R1124 B.n376 B.n143 10.6151
R1125 B.n377 B.n376 10.6151
R1126 B.n378 B.n377 10.6151
R1127 B.n378 B.n141 10.6151
R1128 B.n382 B.n141 10.6151
R1129 B.n383 B.n382 10.6151
R1130 B.n384 B.n383 10.6151
R1131 B.n384 B.n139 10.6151
R1132 B.n388 B.n139 10.6151
R1133 B.n389 B.n388 10.6151
R1134 B.n390 B.n389 10.6151
R1135 B.n390 B.n137 10.6151
R1136 B.n394 B.n137 10.6151
R1137 B.n395 B.n394 10.6151
R1138 B.n396 B.n395 10.6151
R1139 B.n396 B.n135 10.6151
R1140 B.n400 B.n135 10.6151
R1141 B.n401 B.n400 10.6151
R1142 B.n402 B.n401 10.6151
R1143 B.n402 B.n133 10.6151
R1144 B.n406 B.n133 10.6151
R1145 B.n407 B.n406 10.6151
R1146 B.n408 B.n407 10.6151
R1147 B.n408 B.n131 10.6151
R1148 B.n412 B.n131 10.6151
R1149 B.n413 B.n412 10.6151
R1150 B.n414 B.n413 10.6151
R1151 B.n414 B.n129 10.6151
R1152 B.n418 B.n129 10.6151
R1153 B.n419 B.n418 10.6151
R1154 B.n420 B.n419 10.6151
R1155 B.n420 B.n127 10.6151
R1156 B.n424 B.n127 10.6151
R1157 B.n425 B.n424 10.6151
R1158 B.n426 B.n425 10.6151
R1159 B.n426 B.n125 10.6151
R1160 B.n430 B.n125 10.6151
R1161 B.n431 B.n430 10.6151
R1162 B.n432 B.n431 10.6151
R1163 B.n432 B.n123 10.6151
R1164 B.n436 B.n123 10.6151
R1165 B.n437 B.n436 10.6151
R1166 B.n438 B.n437 10.6151
R1167 B.n438 B.n121 10.6151
R1168 B.n442 B.n121 10.6151
R1169 B.n443 B.n442 10.6151
R1170 B.n444 B.n443 10.6151
R1171 B.n444 B.n119 10.6151
R1172 B.n448 B.n119 10.6151
R1173 B.n449 B.n448 10.6151
R1174 B.n450 B.n449 10.6151
R1175 B.n450 B.n117 10.6151
R1176 B.n648 B.n647 9.36635
R1177 B.n630 B.n58 9.36635
R1178 B.n337 B.n336 9.36635
R1179 B.n353 B.n149 9.36635
R1180 B.n785 B.n0 8.11757
R1181 B.n785 B.n1 8.11757
R1182 B.n647 B.n646 1.24928
R1183 B.n58 B.n54 1.24928
R1184 B.n338 B.n337 1.24928
R1185 B.n354 B.n353 1.24928
R1186 VP.n0 VP.t1 266.178
R1187 VP.n0 VP.t0 215.017
R1188 VP VP.n0 0.431811
R1189 VTAIL.n2 VTAIL.t3 51.9591
R1190 VTAIL.n1 VTAIL.t1 51.959
R1191 VTAIL.n3 VTAIL.t0 51.9589
R1192 VTAIL.n0 VTAIL.t2 51.9589
R1193 VTAIL.n1 VTAIL.n0 34.9445
R1194 VTAIL.n3 VTAIL.n2 32.2721
R1195 VTAIL.n2 VTAIL.n1 1.80653
R1196 VTAIL VTAIL.n0 1.19662
R1197 VTAIL VTAIL.n3 0.610414
R1198 VDD1 VDD1.t1 116.067
R1199 VDD1 VDD1.t0 69.3642
R1200 VN VN.t0 266.178
R1201 VN VN.t1 215.447
R1202 VDD2.n0 VDD2.t0 114.874
R1203 VDD2.n0 VDD2.t1 68.6379
R1204 VDD2 VDD2.n0 0.726793
C0 w_n2210_n4966# B 11.232401f
C1 B VTAIL 5.53507f
C2 VDD2 VN 4.509f
C3 VP VN 7.0172f
C4 VDD1 VN 0.1482f
C5 w_n2210_n4966# VN 3.22669f
C6 VN VTAIL 3.82911f
C7 VDD2 VP 0.340811f
C8 VDD2 VDD1 0.696022f
C9 VDD1 VP 4.69783f
C10 VDD2 w_n2210_n4966# 2.38127f
C11 w_n2210_n4966# VP 3.50857f
C12 VDD1 w_n2210_n4966# 2.35329f
C13 VN B 1.17238f
C14 VDD2 VTAIL 7.22988f
C15 VP VTAIL 3.84349f
C16 VDD1 VTAIL 7.17969f
C17 w_n2210_n4966# VTAIL 3.85048f
C18 VDD2 B 2.39399f
C19 VP B 1.63648f
C20 VDD1 B 2.3624f
C21 VDD2 VSUBS 1.201377f
C22 VDD1 VSUBS 7.080801f
C23 VTAIL VSUBS 1.334253f
C24 VN VSUBS 9.5472f
C25 VP VSUBS 2.026141f
C26 B VSUBS 4.710275f
C27 w_n2210_n4966# VSUBS 0.134006p
C28 VDD2.t0 VSUBS 5.97247f
C29 VDD2.t1 VSUBS 4.79975f
C30 VDD2.n0 VSUBS 5.54144f
C31 VN.t1 VSUBS 5.52234f
C32 VN.t0 VSUBS 6.23052f
C33 VDD1.t0 VSUBS 4.83563f
C34 VDD1.t1 VSUBS 6.06613f
C35 VTAIL.t2 VSUBS 4.56529f
C36 VTAIL.n0 VSUBS 3.34976f
C37 VTAIL.t1 VSUBS 4.56532f
C38 VTAIL.n1 VSUBS 3.40435f
C39 VTAIL.t3 VSUBS 4.56531f
C40 VTAIL.n2 VSUBS 3.16501f
C41 VTAIL.t0 VSUBS 4.56529f
C42 VTAIL.n3 VSUBS 3.05791f
C43 VP.t0 VSUBS 5.68244f
C44 VP.t1 VSUBS 6.41386f
C45 VP.n0 VSUBS 6.8088f
C46 B.n0 VSUBS 0.00581f
C47 B.n1 VSUBS 0.00581f
C48 B.n2 VSUBS 0.008592f
C49 B.n3 VSUBS 0.006584f
C50 B.n4 VSUBS 0.006584f
C51 B.n5 VSUBS 0.006584f
C52 B.n6 VSUBS 0.006584f
C53 B.n7 VSUBS 0.006584f
C54 B.n8 VSUBS 0.006584f
C55 B.n9 VSUBS 0.006584f
C56 B.n10 VSUBS 0.006584f
C57 B.n11 VSUBS 0.006584f
C58 B.n12 VSUBS 0.006584f
C59 B.n13 VSUBS 0.006584f
C60 B.n14 VSUBS 0.006584f
C61 B.n15 VSUBS 0.014888f
C62 B.n16 VSUBS 0.006584f
C63 B.n17 VSUBS 0.006584f
C64 B.n18 VSUBS 0.006584f
C65 B.n19 VSUBS 0.006584f
C66 B.n20 VSUBS 0.006584f
C67 B.n21 VSUBS 0.006584f
C68 B.n22 VSUBS 0.006584f
C69 B.n23 VSUBS 0.006584f
C70 B.n24 VSUBS 0.006584f
C71 B.n25 VSUBS 0.006584f
C72 B.n26 VSUBS 0.006584f
C73 B.n27 VSUBS 0.006584f
C74 B.n28 VSUBS 0.006584f
C75 B.n29 VSUBS 0.006584f
C76 B.n30 VSUBS 0.006584f
C77 B.n31 VSUBS 0.006584f
C78 B.n32 VSUBS 0.006584f
C79 B.n33 VSUBS 0.006584f
C80 B.n34 VSUBS 0.006584f
C81 B.n35 VSUBS 0.006584f
C82 B.n36 VSUBS 0.006584f
C83 B.n37 VSUBS 0.006584f
C84 B.n38 VSUBS 0.006584f
C85 B.n39 VSUBS 0.006584f
C86 B.n40 VSUBS 0.006584f
C87 B.n41 VSUBS 0.006584f
C88 B.n42 VSUBS 0.006584f
C89 B.n43 VSUBS 0.006584f
C90 B.n44 VSUBS 0.006584f
C91 B.n45 VSUBS 0.006584f
C92 B.n46 VSUBS 0.006584f
C93 B.n47 VSUBS 0.006584f
C94 B.t4 VSUBS 0.639236f
C95 B.t5 VSUBS 0.659988f
C96 B.t3 VSUBS 2.30477f
C97 B.n48 VSUBS 0.378408f
C98 B.n49 VSUBS 0.068538f
C99 B.n50 VSUBS 0.006584f
C100 B.n51 VSUBS 0.006584f
C101 B.n52 VSUBS 0.006584f
C102 B.n53 VSUBS 0.006584f
C103 B.n54 VSUBS 0.00368f
C104 B.n55 VSUBS 0.006584f
C105 B.t10 VSUBS 0.63921f
C106 B.t11 VSUBS 0.659968f
C107 B.t9 VSUBS 2.30477f
C108 B.n56 VSUBS 0.378429f
C109 B.n57 VSUBS 0.068565f
C110 B.n58 VSUBS 0.015256f
C111 B.n59 VSUBS 0.006584f
C112 B.n60 VSUBS 0.006584f
C113 B.n61 VSUBS 0.006584f
C114 B.n62 VSUBS 0.006584f
C115 B.n63 VSUBS 0.006584f
C116 B.n64 VSUBS 0.006584f
C117 B.n65 VSUBS 0.006584f
C118 B.n66 VSUBS 0.006584f
C119 B.n67 VSUBS 0.006584f
C120 B.n68 VSUBS 0.006584f
C121 B.n69 VSUBS 0.006584f
C122 B.n70 VSUBS 0.006584f
C123 B.n71 VSUBS 0.006584f
C124 B.n72 VSUBS 0.006584f
C125 B.n73 VSUBS 0.006584f
C126 B.n74 VSUBS 0.006584f
C127 B.n75 VSUBS 0.006584f
C128 B.n76 VSUBS 0.006584f
C129 B.n77 VSUBS 0.006584f
C130 B.n78 VSUBS 0.006584f
C131 B.n79 VSUBS 0.006584f
C132 B.n80 VSUBS 0.006584f
C133 B.n81 VSUBS 0.006584f
C134 B.n82 VSUBS 0.006584f
C135 B.n83 VSUBS 0.006584f
C136 B.n84 VSUBS 0.006584f
C137 B.n85 VSUBS 0.006584f
C138 B.n86 VSUBS 0.006584f
C139 B.n87 VSUBS 0.006584f
C140 B.n88 VSUBS 0.006584f
C141 B.n89 VSUBS 0.006584f
C142 B.n90 VSUBS 0.014161f
C143 B.n91 VSUBS 0.006584f
C144 B.n92 VSUBS 0.006584f
C145 B.n93 VSUBS 0.006584f
C146 B.n94 VSUBS 0.006584f
C147 B.n95 VSUBS 0.006584f
C148 B.n96 VSUBS 0.006584f
C149 B.n97 VSUBS 0.006584f
C150 B.n98 VSUBS 0.006584f
C151 B.n99 VSUBS 0.006584f
C152 B.n100 VSUBS 0.006584f
C153 B.n101 VSUBS 0.006584f
C154 B.n102 VSUBS 0.006584f
C155 B.n103 VSUBS 0.006584f
C156 B.n104 VSUBS 0.006584f
C157 B.n105 VSUBS 0.006584f
C158 B.n106 VSUBS 0.006584f
C159 B.n107 VSUBS 0.006584f
C160 B.n108 VSUBS 0.006584f
C161 B.n109 VSUBS 0.006584f
C162 B.n110 VSUBS 0.006584f
C163 B.n111 VSUBS 0.006584f
C164 B.n112 VSUBS 0.006584f
C165 B.n113 VSUBS 0.006584f
C166 B.n114 VSUBS 0.006584f
C167 B.n115 VSUBS 0.006584f
C168 B.n116 VSUBS 0.006584f
C169 B.n117 VSUBS 0.014036f
C170 B.n118 VSUBS 0.006584f
C171 B.n119 VSUBS 0.006584f
C172 B.n120 VSUBS 0.006584f
C173 B.n121 VSUBS 0.006584f
C174 B.n122 VSUBS 0.006584f
C175 B.n123 VSUBS 0.006584f
C176 B.n124 VSUBS 0.006584f
C177 B.n125 VSUBS 0.006584f
C178 B.n126 VSUBS 0.006584f
C179 B.n127 VSUBS 0.006584f
C180 B.n128 VSUBS 0.006584f
C181 B.n129 VSUBS 0.006584f
C182 B.n130 VSUBS 0.006584f
C183 B.n131 VSUBS 0.006584f
C184 B.n132 VSUBS 0.006584f
C185 B.n133 VSUBS 0.006584f
C186 B.n134 VSUBS 0.006584f
C187 B.n135 VSUBS 0.006584f
C188 B.n136 VSUBS 0.006584f
C189 B.n137 VSUBS 0.006584f
C190 B.n138 VSUBS 0.006584f
C191 B.n139 VSUBS 0.006584f
C192 B.n140 VSUBS 0.006584f
C193 B.n141 VSUBS 0.006584f
C194 B.n142 VSUBS 0.006584f
C195 B.n143 VSUBS 0.006584f
C196 B.n144 VSUBS 0.006584f
C197 B.n145 VSUBS 0.006584f
C198 B.n146 VSUBS 0.006584f
C199 B.n147 VSUBS 0.006584f
C200 B.n148 VSUBS 0.006584f
C201 B.n149 VSUBS 0.006197f
C202 B.n150 VSUBS 0.006584f
C203 B.n151 VSUBS 0.006584f
C204 B.n152 VSUBS 0.006584f
C205 B.n153 VSUBS 0.006584f
C206 B.n154 VSUBS 0.006584f
C207 B.t8 VSUBS 0.639236f
C208 B.t7 VSUBS 0.659988f
C209 B.t6 VSUBS 2.30477f
C210 B.n155 VSUBS 0.378408f
C211 B.n156 VSUBS 0.068538f
C212 B.n157 VSUBS 0.006584f
C213 B.n158 VSUBS 0.006584f
C214 B.n159 VSUBS 0.006584f
C215 B.n160 VSUBS 0.006584f
C216 B.n161 VSUBS 0.006584f
C217 B.n162 VSUBS 0.006584f
C218 B.n163 VSUBS 0.006584f
C219 B.n164 VSUBS 0.006584f
C220 B.n165 VSUBS 0.006584f
C221 B.n166 VSUBS 0.006584f
C222 B.n167 VSUBS 0.006584f
C223 B.n168 VSUBS 0.006584f
C224 B.n169 VSUBS 0.006584f
C225 B.n170 VSUBS 0.006584f
C226 B.n171 VSUBS 0.006584f
C227 B.n172 VSUBS 0.006584f
C228 B.n173 VSUBS 0.006584f
C229 B.n174 VSUBS 0.006584f
C230 B.n175 VSUBS 0.006584f
C231 B.n176 VSUBS 0.006584f
C232 B.n177 VSUBS 0.006584f
C233 B.n178 VSUBS 0.006584f
C234 B.n179 VSUBS 0.006584f
C235 B.n180 VSUBS 0.006584f
C236 B.n181 VSUBS 0.006584f
C237 B.n182 VSUBS 0.006584f
C238 B.n183 VSUBS 0.006584f
C239 B.n184 VSUBS 0.006584f
C240 B.n185 VSUBS 0.006584f
C241 B.n186 VSUBS 0.006584f
C242 B.n187 VSUBS 0.006584f
C243 B.n188 VSUBS 0.006584f
C244 B.n189 VSUBS 0.014161f
C245 B.n190 VSUBS 0.006584f
C246 B.n191 VSUBS 0.006584f
C247 B.n192 VSUBS 0.006584f
C248 B.n193 VSUBS 0.006584f
C249 B.n194 VSUBS 0.006584f
C250 B.n195 VSUBS 0.006584f
C251 B.n196 VSUBS 0.006584f
C252 B.n197 VSUBS 0.006584f
C253 B.n198 VSUBS 0.006584f
C254 B.n199 VSUBS 0.006584f
C255 B.n200 VSUBS 0.006584f
C256 B.n201 VSUBS 0.006584f
C257 B.n202 VSUBS 0.006584f
C258 B.n203 VSUBS 0.006584f
C259 B.n204 VSUBS 0.006584f
C260 B.n205 VSUBS 0.006584f
C261 B.n206 VSUBS 0.006584f
C262 B.n207 VSUBS 0.006584f
C263 B.n208 VSUBS 0.006584f
C264 B.n209 VSUBS 0.006584f
C265 B.n210 VSUBS 0.006584f
C266 B.n211 VSUBS 0.006584f
C267 B.n212 VSUBS 0.006584f
C268 B.n213 VSUBS 0.006584f
C269 B.n214 VSUBS 0.006584f
C270 B.n215 VSUBS 0.006584f
C271 B.n216 VSUBS 0.006584f
C272 B.n217 VSUBS 0.006584f
C273 B.n218 VSUBS 0.006584f
C274 B.n219 VSUBS 0.006584f
C275 B.n220 VSUBS 0.006584f
C276 B.n221 VSUBS 0.006584f
C277 B.n222 VSUBS 0.006584f
C278 B.n223 VSUBS 0.006584f
C279 B.n224 VSUBS 0.006584f
C280 B.n225 VSUBS 0.006584f
C281 B.n226 VSUBS 0.006584f
C282 B.n227 VSUBS 0.006584f
C283 B.n228 VSUBS 0.006584f
C284 B.n229 VSUBS 0.006584f
C285 B.n230 VSUBS 0.006584f
C286 B.n231 VSUBS 0.006584f
C287 B.n232 VSUBS 0.006584f
C288 B.n233 VSUBS 0.006584f
C289 B.n234 VSUBS 0.006584f
C290 B.n235 VSUBS 0.006584f
C291 B.n236 VSUBS 0.006584f
C292 B.n237 VSUBS 0.006584f
C293 B.n238 VSUBS 0.014161f
C294 B.n239 VSUBS 0.014888f
C295 B.n240 VSUBS 0.014888f
C296 B.n241 VSUBS 0.006584f
C297 B.n242 VSUBS 0.006584f
C298 B.n243 VSUBS 0.006584f
C299 B.n244 VSUBS 0.006584f
C300 B.n245 VSUBS 0.006584f
C301 B.n246 VSUBS 0.006584f
C302 B.n247 VSUBS 0.006584f
C303 B.n248 VSUBS 0.006584f
C304 B.n249 VSUBS 0.006584f
C305 B.n250 VSUBS 0.006584f
C306 B.n251 VSUBS 0.006584f
C307 B.n252 VSUBS 0.006584f
C308 B.n253 VSUBS 0.006584f
C309 B.n254 VSUBS 0.006584f
C310 B.n255 VSUBS 0.006584f
C311 B.n256 VSUBS 0.006584f
C312 B.n257 VSUBS 0.006584f
C313 B.n258 VSUBS 0.006584f
C314 B.n259 VSUBS 0.006584f
C315 B.n260 VSUBS 0.006584f
C316 B.n261 VSUBS 0.006584f
C317 B.n262 VSUBS 0.006584f
C318 B.n263 VSUBS 0.006584f
C319 B.n264 VSUBS 0.006584f
C320 B.n265 VSUBS 0.006584f
C321 B.n266 VSUBS 0.006584f
C322 B.n267 VSUBS 0.006584f
C323 B.n268 VSUBS 0.006584f
C324 B.n269 VSUBS 0.006584f
C325 B.n270 VSUBS 0.006584f
C326 B.n271 VSUBS 0.006584f
C327 B.n272 VSUBS 0.006584f
C328 B.n273 VSUBS 0.006584f
C329 B.n274 VSUBS 0.006584f
C330 B.n275 VSUBS 0.006584f
C331 B.n276 VSUBS 0.006584f
C332 B.n277 VSUBS 0.006584f
C333 B.n278 VSUBS 0.006584f
C334 B.n279 VSUBS 0.006584f
C335 B.n280 VSUBS 0.006584f
C336 B.n281 VSUBS 0.006584f
C337 B.n282 VSUBS 0.006584f
C338 B.n283 VSUBS 0.006584f
C339 B.n284 VSUBS 0.006584f
C340 B.n285 VSUBS 0.006584f
C341 B.n286 VSUBS 0.006584f
C342 B.n287 VSUBS 0.006584f
C343 B.n288 VSUBS 0.006584f
C344 B.n289 VSUBS 0.006584f
C345 B.n290 VSUBS 0.006584f
C346 B.n291 VSUBS 0.006584f
C347 B.n292 VSUBS 0.006584f
C348 B.n293 VSUBS 0.006584f
C349 B.n294 VSUBS 0.006584f
C350 B.n295 VSUBS 0.006584f
C351 B.n296 VSUBS 0.006584f
C352 B.n297 VSUBS 0.006584f
C353 B.n298 VSUBS 0.006584f
C354 B.n299 VSUBS 0.006584f
C355 B.n300 VSUBS 0.006584f
C356 B.n301 VSUBS 0.006584f
C357 B.n302 VSUBS 0.006584f
C358 B.n303 VSUBS 0.006584f
C359 B.n304 VSUBS 0.006584f
C360 B.n305 VSUBS 0.006584f
C361 B.n306 VSUBS 0.006584f
C362 B.n307 VSUBS 0.006584f
C363 B.n308 VSUBS 0.006584f
C364 B.n309 VSUBS 0.006584f
C365 B.n310 VSUBS 0.006584f
C366 B.n311 VSUBS 0.006584f
C367 B.n312 VSUBS 0.006584f
C368 B.n313 VSUBS 0.006584f
C369 B.n314 VSUBS 0.006584f
C370 B.n315 VSUBS 0.006584f
C371 B.n316 VSUBS 0.006584f
C372 B.n317 VSUBS 0.006584f
C373 B.n318 VSUBS 0.006584f
C374 B.n319 VSUBS 0.006584f
C375 B.n320 VSUBS 0.006584f
C376 B.n321 VSUBS 0.006584f
C377 B.n322 VSUBS 0.006584f
C378 B.n323 VSUBS 0.006584f
C379 B.n324 VSUBS 0.006584f
C380 B.n325 VSUBS 0.006584f
C381 B.n326 VSUBS 0.006584f
C382 B.n327 VSUBS 0.006584f
C383 B.n328 VSUBS 0.006584f
C384 B.n329 VSUBS 0.006584f
C385 B.n330 VSUBS 0.006584f
C386 B.n331 VSUBS 0.006584f
C387 B.n332 VSUBS 0.006584f
C388 B.n333 VSUBS 0.006584f
C389 B.n334 VSUBS 0.006584f
C390 B.n335 VSUBS 0.006584f
C391 B.n336 VSUBS 0.006197f
C392 B.n337 VSUBS 0.015256f
C393 B.n338 VSUBS 0.00368f
C394 B.n339 VSUBS 0.006584f
C395 B.n340 VSUBS 0.006584f
C396 B.n341 VSUBS 0.006584f
C397 B.n342 VSUBS 0.006584f
C398 B.n343 VSUBS 0.006584f
C399 B.n344 VSUBS 0.006584f
C400 B.n345 VSUBS 0.006584f
C401 B.n346 VSUBS 0.006584f
C402 B.n347 VSUBS 0.006584f
C403 B.n348 VSUBS 0.006584f
C404 B.n349 VSUBS 0.006584f
C405 B.n350 VSUBS 0.006584f
C406 B.t2 VSUBS 0.63921f
C407 B.t1 VSUBS 0.659968f
C408 B.t0 VSUBS 2.30477f
C409 B.n351 VSUBS 0.378429f
C410 B.n352 VSUBS 0.068565f
C411 B.n353 VSUBS 0.015256f
C412 B.n354 VSUBS 0.00368f
C413 B.n355 VSUBS 0.006584f
C414 B.n356 VSUBS 0.006584f
C415 B.n357 VSUBS 0.006584f
C416 B.n358 VSUBS 0.006584f
C417 B.n359 VSUBS 0.006584f
C418 B.n360 VSUBS 0.006584f
C419 B.n361 VSUBS 0.006584f
C420 B.n362 VSUBS 0.006584f
C421 B.n363 VSUBS 0.006584f
C422 B.n364 VSUBS 0.006584f
C423 B.n365 VSUBS 0.006584f
C424 B.n366 VSUBS 0.006584f
C425 B.n367 VSUBS 0.006584f
C426 B.n368 VSUBS 0.006584f
C427 B.n369 VSUBS 0.006584f
C428 B.n370 VSUBS 0.006584f
C429 B.n371 VSUBS 0.006584f
C430 B.n372 VSUBS 0.006584f
C431 B.n373 VSUBS 0.006584f
C432 B.n374 VSUBS 0.006584f
C433 B.n375 VSUBS 0.006584f
C434 B.n376 VSUBS 0.006584f
C435 B.n377 VSUBS 0.006584f
C436 B.n378 VSUBS 0.006584f
C437 B.n379 VSUBS 0.006584f
C438 B.n380 VSUBS 0.006584f
C439 B.n381 VSUBS 0.006584f
C440 B.n382 VSUBS 0.006584f
C441 B.n383 VSUBS 0.006584f
C442 B.n384 VSUBS 0.006584f
C443 B.n385 VSUBS 0.006584f
C444 B.n386 VSUBS 0.006584f
C445 B.n387 VSUBS 0.006584f
C446 B.n388 VSUBS 0.006584f
C447 B.n389 VSUBS 0.006584f
C448 B.n390 VSUBS 0.006584f
C449 B.n391 VSUBS 0.006584f
C450 B.n392 VSUBS 0.006584f
C451 B.n393 VSUBS 0.006584f
C452 B.n394 VSUBS 0.006584f
C453 B.n395 VSUBS 0.006584f
C454 B.n396 VSUBS 0.006584f
C455 B.n397 VSUBS 0.006584f
C456 B.n398 VSUBS 0.006584f
C457 B.n399 VSUBS 0.006584f
C458 B.n400 VSUBS 0.006584f
C459 B.n401 VSUBS 0.006584f
C460 B.n402 VSUBS 0.006584f
C461 B.n403 VSUBS 0.006584f
C462 B.n404 VSUBS 0.006584f
C463 B.n405 VSUBS 0.006584f
C464 B.n406 VSUBS 0.006584f
C465 B.n407 VSUBS 0.006584f
C466 B.n408 VSUBS 0.006584f
C467 B.n409 VSUBS 0.006584f
C468 B.n410 VSUBS 0.006584f
C469 B.n411 VSUBS 0.006584f
C470 B.n412 VSUBS 0.006584f
C471 B.n413 VSUBS 0.006584f
C472 B.n414 VSUBS 0.006584f
C473 B.n415 VSUBS 0.006584f
C474 B.n416 VSUBS 0.006584f
C475 B.n417 VSUBS 0.006584f
C476 B.n418 VSUBS 0.006584f
C477 B.n419 VSUBS 0.006584f
C478 B.n420 VSUBS 0.006584f
C479 B.n421 VSUBS 0.006584f
C480 B.n422 VSUBS 0.006584f
C481 B.n423 VSUBS 0.006584f
C482 B.n424 VSUBS 0.006584f
C483 B.n425 VSUBS 0.006584f
C484 B.n426 VSUBS 0.006584f
C485 B.n427 VSUBS 0.006584f
C486 B.n428 VSUBS 0.006584f
C487 B.n429 VSUBS 0.006584f
C488 B.n430 VSUBS 0.006584f
C489 B.n431 VSUBS 0.006584f
C490 B.n432 VSUBS 0.006584f
C491 B.n433 VSUBS 0.006584f
C492 B.n434 VSUBS 0.006584f
C493 B.n435 VSUBS 0.006584f
C494 B.n436 VSUBS 0.006584f
C495 B.n437 VSUBS 0.006584f
C496 B.n438 VSUBS 0.006584f
C497 B.n439 VSUBS 0.006584f
C498 B.n440 VSUBS 0.006584f
C499 B.n441 VSUBS 0.006584f
C500 B.n442 VSUBS 0.006584f
C501 B.n443 VSUBS 0.006584f
C502 B.n444 VSUBS 0.006584f
C503 B.n445 VSUBS 0.006584f
C504 B.n446 VSUBS 0.006584f
C505 B.n447 VSUBS 0.006584f
C506 B.n448 VSUBS 0.006584f
C507 B.n449 VSUBS 0.006584f
C508 B.n450 VSUBS 0.006584f
C509 B.n451 VSUBS 0.006584f
C510 B.n452 VSUBS 0.014888f
C511 B.n453 VSUBS 0.014161f
C512 B.n454 VSUBS 0.015013f
C513 B.n455 VSUBS 0.006584f
C514 B.n456 VSUBS 0.006584f
C515 B.n457 VSUBS 0.006584f
C516 B.n458 VSUBS 0.006584f
C517 B.n459 VSUBS 0.006584f
C518 B.n460 VSUBS 0.006584f
C519 B.n461 VSUBS 0.006584f
C520 B.n462 VSUBS 0.006584f
C521 B.n463 VSUBS 0.006584f
C522 B.n464 VSUBS 0.006584f
C523 B.n465 VSUBS 0.006584f
C524 B.n466 VSUBS 0.006584f
C525 B.n467 VSUBS 0.006584f
C526 B.n468 VSUBS 0.006584f
C527 B.n469 VSUBS 0.006584f
C528 B.n470 VSUBS 0.006584f
C529 B.n471 VSUBS 0.006584f
C530 B.n472 VSUBS 0.006584f
C531 B.n473 VSUBS 0.006584f
C532 B.n474 VSUBS 0.006584f
C533 B.n475 VSUBS 0.006584f
C534 B.n476 VSUBS 0.006584f
C535 B.n477 VSUBS 0.006584f
C536 B.n478 VSUBS 0.006584f
C537 B.n479 VSUBS 0.006584f
C538 B.n480 VSUBS 0.006584f
C539 B.n481 VSUBS 0.006584f
C540 B.n482 VSUBS 0.006584f
C541 B.n483 VSUBS 0.006584f
C542 B.n484 VSUBS 0.006584f
C543 B.n485 VSUBS 0.006584f
C544 B.n486 VSUBS 0.006584f
C545 B.n487 VSUBS 0.006584f
C546 B.n488 VSUBS 0.006584f
C547 B.n489 VSUBS 0.006584f
C548 B.n490 VSUBS 0.006584f
C549 B.n491 VSUBS 0.006584f
C550 B.n492 VSUBS 0.006584f
C551 B.n493 VSUBS 0.006584f
C552 B.n494 VSUBS 0.006584f
C553 B.n495 VSUBS 0.006584f
C554 B.n496 VSUBS 0.006584f
C555 B.n497 VSUBS 0.006584f
C556 B.n498 VSUBS 0.006584f
C557 B.n499 VSUBS 0.006584f
C558 B.n500 VSUBS 0.006584f
C559 B.n501 VSUBS 0.006584f
C560 B.n502 VSUBS 0.006584f
C561 B.n503 VSUBS 0.006584f
C562 B.n504 VSUBS 0.006584f
C563 B.n505 VSUBS 0.006584f
C564 B.n506 VSUBS 0.006584f
C565 B.n507 VSUBS 0.006584f
C566 B.n508 VSUBS 0.006584f
C567 B.n509 VSUBS 0.006584f
C568 B.n510 VSUBS 0.006584f
C569 B.n511 VSUBS 0.006584f
C570 B.n512 VSUBS 0.006584f
C571 B.n513 VSUBS 0.006584f
C572 B.n514 VSUBS 0.006584f
C573 B.n515 VSUBS 0.006584f
C574 B.n516 VSUBS 0.006584f
C575 B.n517 VSUBS 0.006584f
C576 B.n518 VSUBS 0.006584f
C577 B.n519 VSUBS 0.006584f
C578 B.n520 VSUBS 0.006584f
C579 B.n521 VSUBS 0.006584f
C580 B.n522 VSUBS 0.006584f
C581 B.n523 VSUBS 0.006584f
C582 B.n524 VSUBS 0.006584f
C583 B.n525 VSUBS 0.006584f
C584 B.n526 VSUBS 0.006584f
C585 B.n527 VSUBS 0.006584f
C586 B.n528 VSUBS 0.006584f
C587 B.n529 VSUBS 0.006584f
C588 B.n530 VSUBS 0.006584f
C589 B.n531 VSUBS 0.006584f
C590 B.n532 VSUBS 0.006584f
C591 B.n533 VSUBS 0.014161f
C592 B.n534 VSUBS 0.014888f
C593 B.n535 VSUBS 0.014888f
C594 B.n536 VSUBS 0.006584f
C595 B.n537 VSUBS 0.006584f
C596 B.n538 VSUBS 0.006584f
C597 B.n539 VSUBS 0.006584f
C598 B.n540 VSUBS 0.006584f
C599 B.n541 VSUBS 0.006584f
C600 B.n542 VSUBS 0.006584f
C601 B.n543 VSUBS 0.006584f
C602 B.n544 VSUBS 0.006584f
C603 B.n545 VSUBS 0.006584f
C604 B.n546 VSUBS 0.006584f
C605 B.n547 VSUBS 0.006584f
C606 B.n548 VSUBS 0.006584f
C607 B.n549 VSUBS 0.006584f
C608 B.n550 VSUBS 0.006584f
C609 B.n551 VSUBS 0.006584f
C610 B.n552 VSUBS 0.006584f
C611 B.n553 VSUBS 0.006584f
C612 B.n554 VSUBS 0.006584f
C613 B.n555 VSUBS 0.006584f
C614 B.n556 VSUBS 0.006584f
C615 B.n557 VSUBS 0.006584f
C616 B.n558 VSUBS 0.006584f
C617 B.n559 VSUBS 0.006584f
C618 B.n560 VSUBS 0.006584f
C619 B.n561 VSUBS 0.006584f
C620 B.n562 VSUBS 0.006584f
C621 B.n563 VSUBS 0.006584f
C622 B.n564 VSUBS 0.006584f
C623 B.n565 VSUBS 0.006584f
C624 B.n566 VSUBS 0.006584f
C625 B.n567 VSUBS 0.006584f
C626 B.n568 VSUBS 0.006584f
C627 B.n569 VSUBS 0.006584f
C628 B.n570 VSUBS 0.006584f
C629 B.n571 VSUBS 0.006584f
C630 B.n572 VSUBS 0.006584f
C631 B.n573 VSUBS 0.006584f
C632 B.n574 VSUBS 0.006584f
C633 B.n575 VSUBS 0.006584f
C634 B.n576 VSUBS 0.006584f
C635 B.n577 VSUBS 0.006584f
C636 B.n578 VSUBS 0.006584f
C637 B.n579 VSUBS 0.006584f
C638 B.n580 VSUBS 0.006584f
C639 B.n581 VSUBS 0.006584f
C640 B.n582 VSUBS 0.006584f
C641 B.n583 VSUBS 0.006584f
C642 B.n584 VSUBS 0.006584f
C643 B.n585 VSUBS 0.006584f
C644 B.n586 VSUBS 0.006584f
C645 B.n587 VSUBS 0.006584f
C646 B.n588 VSUBS 0.006584f
C647 B.n589 VSUBS 0.006584f
C648 B.n590 VSUBS 0.006584f
C649 B.n591 VSUBS 0.006584f
C650 B.n592 VSUBS 0.006584f
C651 B.n593 VSUBS 0.006584f
C652 B.n594 VSUBS 0.006584f
C653 B.n595 VSUBS 0.006584f
C654 B.n596 VSUBS 0.006584f
C655 B.n597 VSUBS 0.006584f
C656 B.n598 VSUBS 0.006584f
C657 B.n599 VSUBS 0.006584f
C658 B.n600 VSUBS 0.006584f
C659 B.n601 VSUBS 0.006584f
C660 B.n602 VSUBS 0.006584f
C661 B.n603 VSUBS 0.006584f
C662 B.n604 VSUBS 0.006584f
C663 B.n605 VSUBS 0.006584f
C664 B.n606 VSUBS 0.006584f
C665 B.n607 VSUBS 0.006584f
C666 B.n608 VSUBS 0.006584f
C667 B.n609 VSUBS 0.006584f
C668 B.n610 VSUBS 0.006584f
C669 B.n611 VSUBS 0.006584f
C670 B.n612 VSUBS 0.006584f
C671 B.n613 VSUBS 0.006584f
C672 B.n614 VSUBS 0.006584f
C673 B.n615 VSUBS 0.006584f
C674 B.n616 VSUBS 0.006584f
C675 B.n617 VSUBS 0.006584f
C676 B.n618 VSUBS 0.006584f
C677 B.n619 VSUBS 0.006584f
C678 B.n620 VSUBS 0.006584f
C679 B.n621 VSUBS 0.006584f
C680 B.n622 VSUBS 0.006584f
C681 B.n623 VSUBS 0.006584f
C682 B.n624 VSUBS 0.006584f
C683 B.n625 VSUBS 0.006584f
C684 B.n626 VSUBS 0.006584f
C685 B.n627 VSUBS 0.006584f
C686 B.n628 VSUBS 0.006584f
C687 B.n629 VSUBS 0.006584f
C688 B.n630 VSUBS 0.006197f
C689 B.n631 VSUBS 0.006584f
C690 B.n632 VSUBS 0.006584f
C691 B.n633 VSUBS 0.006584f
C692 B.n634 VSUBS 0.006584f
C693 B.n635 VSUBS 0.006584f
C694 B.n636 VSUBS 0.006584f
C695 B.n637 VSUBS 0.006584f
C696 B.n638 VSUBS 0.006584f
C697 B.n639 VSUBS 0.006584f
C698 B.n640 VSUBS 0.006584f
C699 B.n641 VSUBS 0.006584f
C700 B.n642 VSUBS 0.006584f
C701 B.n643 VSUBS 0.006584f
C702 B.n644 VSUBS 0.006584f
C703 B.n645 VSUBS 0.006584f
C704 B.n646 VSUBS 0.00368f
C705 B.n647 VSUBS 0.015256f
C706 B.n648 VSUBS 0.006197f
C707 B.n649 VSUBS 0.006584f
C708 B.n650 VSUBS 0.006584f
C709 B.n651 VSUBS 0.006584f
C710 B.n652 VSUBS 0.006584f
C711 B.n653 VSUBS 0.006584f
C712 B.n654 VSUBS 0.006584f
C713 B.n655 VSUBS 0.006584f
C714 B.n656 VSUBS 0.006584f
C715 B.n657 VSUBS 0.006584f
C716 B.n658 VSUBS 0.006584f
C717 B.n659 VSUBS 0.006584f
C718 B.n660 VSUBS 0.006584f
C719 B.n661 VSUBS 0.006584f
C720 B.n662 VSUBS 0.006584f
C721 B.n663 VSUBS 0.006584f
C722 B.n664 VSUBS 0.006584f
C723 B.n665 VSUBS 0.006584f
C724 B.n666 VSUBS 0.006584f
C725 B.n667 VSUBS 0.006584f
C726 B.n668 VSUBS 0.006584f
C727 B.n669 VSUBS 0.006584f
C728 B.n670 VSUBS 0.006584f
C729 B.n671 VSUBS 0.006584f
C730 B.n672 VSUBS 0.006584f
C731 B.n673 VSUBS 0.006584f
C732 B.n674 VSUBS 0.006584f
C733 B.n675 VSUBS 0.006584f
C734 B.n676 VSUBS 0.006584f
C735 B.n677 VSUBS 0.006584f
C736 B.n678 VSUBS 0.006584f
C737 B.n679 VSUBS 0.006584f
C738 B.n680 VSUBS 0.006584f
C739 B.n681 VSUBS 0.006584f
C740 B.n682 VSUBS 0.006584f
C741 B.n683 VSUBS 0.006584f
C742 B.n684 VSUBS 0.006584f
C743 B.n685 VSUBS 0.006584f
C744 B.n686 VSUBS 0.006584f
C745 B.n687 VSUBS 0.006584f
C746 B.n688 VSUBS 0.006584f
C747 B.n689 VSUBS 0.006584f
C748 B.n690 VSUBS 0.006584f
C749 B.n691 VSUBS 0.006584f
C750 B.n692 VSUBS 0.006584f
C751 B.n693 VSUBS 0.006584f
C752 B.n694 VSUBS 0.006584f
C753 B.n695 VSUBS 0.006584f
C754 B.n696 VSUBS 0.006584f
C755 B.n697 VSUBS 0.006584f
C756 B.n698 VSUBS 0.006584f
C757 B.n699 VSUBS 0.006584f
C758 B.n700 VSUBS 0.006584f
C759 B.n701 VSUBS 0.006584f
C760 B.n702 VSUBS 0.006584f
C761 B.n703 VSUBS 0.006584f
C762 B.n704 VSUBS 0.006584f
C763 B.n705 VSUBS 0.006584f
C764 B.n706 VSUBS 0.006584f
C765 B.n707 VSUBS 0.006584f
C766 B.n708 VSUBS 0.006584f
C767 B.n709 VSUBS 0.006584f
C768 B.n710 VSUBS 0.006584f
C769 B.n711 VSUBS 0.006584f
C770 B.n712 VSUBS 0.006584f
C771 B.n713 VSUBS 0.006584f
C772 B.n714 VSUBS 0.006584f
C773 B.n715 VSUBS 0.006584f
C774 B.n716 VSUBS 0.006584f
C775 B.n717 VSUBS 0.006584f
C776 B.n718 VSUBS 0.006584f
C777 B.n719 VSUBS 0.006584f
C778 B.n720 VSUBS 0.006584f
C779 B.n721 VSUBS 0.006584f
C780 B.n722 VSUBS 0.006584f
C781 B.n723 VSUBS 0.006584f
C782 B.n724 VSUBS 0.006584f
C783 B.n725 VSUBS 0.006584f
C784 B.n726 VSUBS 0.006584f
C785 B.n727 VSUBS 0.006584f
C786 B.n728 VSUBS 0.006584f
C787 B.n729 VSUBS 0.006584f
C788 B.n730 VSUBS 0.006584f
C789 B.n731 VSUBS 0.006584f
C790 B.n732 VSUBS 0.006584f
C791 B.n733 VSUBS 0.006584f
C792 B.n734 VSUBS 0.006584f
C793 B.n735 VSUBS 0.006584f
C794 B.n736 VSUBS 0.006584f
C795 B.n737 VSUBS 0.006584f
C796 B.n738 VSUBS 0.006584f
C797 B.n739 VSUBS 0.006584f
C798 B.n740 VSUBS 0.006584f
C799 B.n741 VSUBS 0.006584f
C800 B.n742 VSUBS 0.006584f
C801 B.n743 VSUBS 0.006584f
C802 B.n744 VSUBS 0.014888f
C803 B.n745 VSUBS 0.014161f
C804 B.n746 VSUBS 0.014161f
C805 B.n747 VSUBS 0.006584f
C806 B.n748 VSUBS 0.006584f
C807 B.n749 VSUBS 0.006584f
C808 B.n750 VSUBS 0.006584f
C809 B.n751 VSUBS 0.006584f
C810 B.n752 VSUBS 0.006584f
C811 B.n753 VSUBS 0.006584f
C812 B.n754 VSUBS 0.006584f
C813 B.n755 VSUBS 0.006584f
C814 B.n756 VSUBS 0.006584f
C815 B.n757 VSUBS 0.006584f
C816 B.n758 VSUBS 0.006584f
C817 B.n759 VSUBS 0.006584f
C818 B.n760 VSUBS 0.006584f
C819 B.n761 VSUBS 0.006584f
C820 B.n762 VSUBS 0.006584f
C821 B.n763 VSUBS 0.006584f
C822 B.n764 VSUBS 0.006584f
C823 B.n765 VSUBS 0.006584f
C824 B.n766 VSUBS 0.006584f
C825 B.n767 VSUBS 0.006584f
C826 B.n768 VSUBS 0.006584f
C827 B.n769 VSUBS 0.006584f
C828 B.n770 VSUBS 0.006584f
C829 B.n771 VSUBS 0.006584f
C830 B.n772 VSUBS 0.006584f
C831 B.n773 VSUBS 0.006584f
C832 B.n774 VSUBS 0.006584f
C833 B.n775 VSUBS 0.006584f
C834 B.n776 VSUBS 0.006584f
C835 B.n777 VSUBS 0.006584f
C836 B.n778 VSUBS 0.006584f
C837 B.n779 VSUBS 0.006584f
C838 B.n780 VSUBS 0.006584f
C839 B.n781 VSUBS 0.006584f
C840 B.n782 VSUBS 0.006584f
C841 B.n783 VSUBS 0.008592f
C842 B.n784 VSUBS 0.009153f
C843 B.n785 VSUBS 0.018202f
.ends

