* NGSPICE file created from diff_pair_sample_0892.ext - technology: sky130A

.subckt diff_pair_sample_0892 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t3 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
X1 VTAIL.t3 VP.t0 VDD1.t9 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
X2 B.t11 B.t9 B.t10 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=3.3111 pd=17.76 as=0 ps=0 w=8.49 l=2.09
X3 B.t8 B.t6 B.t7 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=3.3111 pd=17.76 as=0 ps=0 w=8.49 l=2.09
X4 VDD1.t8 VP.t1 VTAIL.t1 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=3.3111 ps=17.76 w=8.49 l=2.09
X5 VTAIL.t18 VN.t1 VDD2.t2 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
X6 VDD1.t7 VP.t2 VTAIL.t2 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=3.3111 pd=17.76 as=1.40085 ps=8.82 w=8.49 l=2.09
X7 VTAIL.t17 VN.t2 VDD2.t8 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
X8 VDD1.t6 VP.t3 VTAIL.t5 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
X9 VDD2.t7 VN.t3 VTAIL.t16 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=3.3111 ps=17.76 w=8.49 l=2.09
X10 VTAIL.t15 VN.t4 VDD2.t6 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
X11 B.t5 B.t3 B.t4 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=3.3111 pd=17.76 as=0 ps=0 w=8.49 l=2.09
X12 VDD2.t9 VN.t5 VTAIL.t14 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=3.3111 pd=17.76 as=1.40085 ps=8.82 w=8.49 l=2.09
X13 VDD1.t5 VP.t4 VTAIL.t0 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=3.3111 ps=17.76 w=8.49 l=2.09
X14 B.t2 B.t0 B.t1 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=3.3111 pd=17.76 as=0 ps=0 w=8.49 l=2.09
X15 VDD1.t4 VP.t5 VTAIL.t4 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=3.3111 pd=17.76 as=1.40085 ps=8.82 w=8.49 l=2.09
X16 VDD1.t3 VP.t6 VTAIL.t8 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
X17 VDD2.t4 VN.t6 VTAIL.t13 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=3.3111 ps=17.76 w=8.49 l=2.09
X18 VDD2.t5 VN.t7 VTAIL.t12 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
X19 VDD2.t0 VN.t8 VTAIL.t11 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=3.3111 pd=17.76 as=1.40085 ps=8.82 w=8.49 l=2.09
X20 VTAIL.t7 VP.t7 VDD1.t2 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
X21 VTAIL.t6 VP.t8 VDD1.t1 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
X22 VDD2.t1 VN.t9 VTAIL.t10 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
X23 VTAIL.t9 VP.t9 VDD1.t0 w_n3874_n2666# sky130_fd_pr__pfet_01v8 ad=1.40085 pd=8.82 as=1.40085 ps=8.82 w=8.49 l=2.09
R0 VN.n63 VN.n33 161.3
R1 VN.n62 VN.n61 161.3
R2 VN.n60 VN.n34 161.3
R3 VN.n59 VN.n58 161.3
R4 VN.n57 VN.n35 161.3
R5 VN.n55 VN.n54 161.3
R6 VN.n53 VN.n36 161.3
R7 VN.n52 VN.n51 161.3
R8 VN.n50 VN.n37 161.3
R9 VN.n49 VN.n48 161.3
R10 VN.n47 VN.n38 161.3
R11 VN.n46 VN.n45 161.3
R12 VN.n44 VN.n39 161.3
R13 VN.n43 VN.n42 161.3
R14 VN.n30 VN.n0 161.3
R15 VN.n29 VN.n28 161.3
R16 VN.n27 VN.n1 161.3
R17 VN.n26 VN.n25 161.3
R18 VN.n24 VN.n2 161.3
R19 VN.n22 VN.n21 161.3
R20 VN.n20 VN.n3 161.3
R21 VN.n19 VN.n18 161.3
R22 VN.n17 VN.n4 161.3
R23 VN.n16 VN.n15 161.3
R24 VN.n14 VN.n5 161.3
R25 VN.n13 VN.n12 161.3
R26 VN.n11 VN.n6 161.3
R27 VN.n10 VN.n9 161.3
R28 VN.n8 VN.t5 131.347
R29 VN.n41 VN.t3 131.347
R30 VN.n16 VN.t7 97.8995
R31 VN.n7 VN.t0 97.8995
R32 VN.n23 VN.t2 97.8995
R33 VN.n31 VN.t6 97.8995
R34 VN.n49 VN.t9 97.8995
R35 VN.n40 VN.t1 97.8995
R36 VN.n56 VN.t4 97.8995
R37 VN.n64 VN.t8 97.8995
R38 VN.n32 VN.n31 94.1189
R39 VN.n65 VN.n64 94.1189
R40 VN.n12 VN.n11 56.5193
R41 VN.n18 VN.n3 56.5193
R42 VN.n45 VN.n44 56.5193
R43 VN.n51 VN.n36 56.5193
R44 VN.n29 VN.n1 53.1199
R45 VN.n62 VN.n34 53.1199
R46 VN.n8 VN.n7 50.0611
R47 VN.n41 VN.n40 50.0611
R48 VN VN.n65 47.9603
R49 VN.n25 VN.n1 27.8669
R50 VN.n58 VN.n34 27.8669
R51 VN.n11 VN.n10 24.4675
R52 VN.n12 VN.n5 24.4675
R53 VN.n16 VN.n5 24.4675
R54 VN.n17 VN.n16 24.4675
R55 VN.n18 VN.n17 24.4675
R56 VN.n22 VN.n3 24.4675
R57 VN.n25 VN.n24 24.4675
R58 VN.n30 VN.n29 24.4675
R59 VN.n44 VN.n43 24.4675
R60 VN.n51 VN.n50 24.4675
R61 VN.n50 VN.n49 24.4675
R62 VN.n49 VN.n38 24.4675
R63 VN.n45 VN.n38 24.4675
R64 VN.n58 VN.n57 24.4675
R65 VN.n55 VN.n36 24.4675
R66 VN.n63 VN.n62 24.4675
R67 VN.n10 VN.n7 20.5528
R68 VN.n23 VN.n22 20.5528
R69 VN.n43 VN.n40 20.5528
R70 VN.n56 VN.n55 20.5528
R71 VN.n31 VN.n30 16.6381
R72 VN.n64 VN.n63 16.6381
R73 VN.n42 VN.n41 9.28282
R74 VN.n9 VN.n8 9.28282
R75 VN.n24 VN.n23 3.91522
R76 VN.n57 VN.n56 3.91522
R77 VN.n65 VN.n33 0.278367
R78 VN.n32 VN.n0 0.278367
R79 VN.n61 VN.n33 0.189894
R80 VN.n61 VN.n60 0.189894
R81 VN.n60 VN.n59 0.189894
R82 VN.n59 VN.n35 0.189894
R83 VN.n54 VN.n35 0.189894
R84 VN.n54 VN.n53 0.189894
R85 VN.n53 VN.n52 0.189894
R86 VN.n52 VN.n37 0.189894
R87 VN.n48 VN.n37 0.189894
R88 VN.n48 VN.n47 0.189894
R89 VN.n47 VN.n46 0.189894
R90 VN.n46 VN.n39 0.189894
R91 VN.n42 VN.n39 0.189894
R92 VN.n9 VN.n6 0.189894
R93 VN.n13 VN.n6 0.189894
R94 VN.n14 VN.n13 0.189894
R95 VN.n15 VN.n14 0.189894
R96 VN.n15 VN.n4 0.189894
R97 VN.n19 VN.n4 0.189894
R98 VN.n20 VN.n19 0.189894
R99 VN.n21 VN.n20 0.189894
R100 VN.n21 VN.n2 0.189894
R101 VN.n26 VN.n2 0.189894
R102 VN.n27 VN.n26 0.189894
R103 VN.n28 VN.n27 0.189894
R104 VN.n28 VN.n0 0.189894
R105 VN VN.n32 0.153454
R106 VDD2.n1 VDD2.t9 87.032
R107 VDD2.n4 VDD2.t0 84.946
R108 VDD2.n3 VDD2.n2 82.6267
R109 VDD2 VDD2.n7 82.6239
R110 VDD2.n6 VDD2.n5 81.1174
R111 VDD2.n1 VDD2.n0 81.1174
R112 VDD2.n4 VDD2.n3 40.9437
R113 VDD2.n7 VDD2.t2 3.82912
R114 VDD2.n7 VDD2.t7 3.82912
R115 VDD2.n5 VDD2.t6 3.82912
R116 VDD2.n5 VDD2.t1 3.82912
R117 VDD2.n2 VDD2.t8 3.82912
R118 VDD2.n2 VDD2.t4 3.82912
R119 VDD2.n0 VDD2.t3 3.82912
R120 VDD2.n0 VDD2.t5 3.82912
R121 VDD2.n6 VDD2.n4 2.08671
R122 VDD2 VDD2.n6 0.580241
R123 VDD2.n3 VDD2.n1 0.466706
R124 VTAIL.n11 VTAIL.t16 68.2672
R125 VTAIL.n16 VTAIL.t0 68.2672
R126 VTAIL.n17 VTAIL.t13 68.267
R127 VTAIL.n2 VTAIL.t1 68.267
R128 VTAIL.n15 VTAIL.n14 64.4386
R129 VTAIL.n13 VTAIL.n12 64.4386
R130 VTAIL.n10 VTAIL.n9 64.4386
R131 VTAIL.n8 VTAIL.n7 64.4386
R132 VTAIL.n19 VTAIL.n18 64.4386
R133 VTAIL.n1 VTAIL.n0 64.4386
R134 VTAIL.n4 VTAIL.n3 64.4386
R135 VTAIL.n6 VTAIL.n5 64.4386
R136 VTAIL.n8 VTAIL.n6 23.8583
R137 VTAIL.n17 VTAIL.n16 21.7721
R138 VTAIL.n18 VTAIL.t12 3.82912
R139 VTAIL.n18 VTAIL.t17 3.82912
R140 VTAIL.n0 VTAIL.t14 3.82912
R141 VTAIL.n0 VTAIL.t19 3.82912
R142 VTAIL.n3 VTAIL.t5 3.82912
R143 VTAIL.n3 VTAIL.t9 3.82912
R144 VTAIL.n5 VTAIL.t4 3.82912
R145 VTAIL.n5 VTAIL.t7 3.82912
R146 VTAIL.n14 VTAIL.t8 3.82912
R147 VTAIL.n14 VTAIL.t3 3.82912
R148 VTAIL.n12 VTAIL.t2 3.82912
R149 VTAIL.n12 VTAIL.t6 3.82912
R150 VTAIL.n9 VTAIL.t10 3.82912
R151 VTAIL.n9 VTAIL.t18 3.82912
R152 VTAIL.n7 VTAIL.t11 3.82912
R153 VTAIL.n7 VTAIL.t15 3.82912
R154 VTAIL.n10 VTAIL.n8 2.08671
R155 VTAIL.n11 VTAIL.n10 2.08671
R156 VTAIL.n15 VTAIL.n13 2.08671
R157 VTAIL.n16 VTAIL.n15 2.08671
R158 VTAIL.n6 VTAIL.n4 2.08671
R159 VTAIL.n4 VTAIL.n2 2.08671
R160 VTAIL.n19 VTAIL.n17 2.08671
R161 VTAIL VTAIL.n1 1.62334
R162 VTAIL.n13 VTAIL.n11 1.51343
R163 VTAIL.n2 VTAIL.n1 1.51343
R164 VTAIL VTAIL.n19 0.463862
R165 VP.n20 VP.n19 161.3
R166 VP.n21 VP.n16 161.3
R167 VP.n23 VP.n22 161.3
R168 VP.n24 VP.n15 161.3
R169 VP.n26 VP.n25 161.3
R170 VP.n27 VP.n14 161.3
R171 VP.n29 VP.n28 161.3
R172 VP.n30 VP.n13 161.3
R173 VP.n32 VP.n31 161.3
R174 VP.n34 VP.n12 161.3
R175 VP.n36 VP.n35 161.3
R176 VP.n37 VP.n11 161.3
R177 VP.n39 VP.n38 161.3
R178 VP.n40 VP.n10 161.3
R179 VP.n74 VP.n0 161.3
R180 VP.n73 VP.n72 161.3
R181 VP.n71 VP.n1 161.3
R182 VP.n70 VP.n69 161.3
R183 VP.n68 VP.n2 161.3
R184 VP.n66 VP.n65 161.3
R185 VP.n64 VP.n3 161.3
R186 VP.n63 VP.n62 161.3
R187 VP.n61 VP.n4 161.3
R188 VP.n60 VP.n59 161.3
R189 VP.n58 VP.n5 161.3
R190 VP.n57 VP.n56 161.3
R191 VP.n55 VP.n6 161.3
R192 VP.n54 VP.n53 161.3
R193 VP.n52 VP.n51 161.3
R194 VP.n50 VP.n8 161.3
R195 VP.n49 VP.n48 161.3
R196 VP.n47 VP.n9 161.3
R197 VP.n46 VP.n45 161.3
R198 VP.n18 VP.t2 131.347
R199 VP.n60 VP.t3 97.8995
R200 VP.n44 VP.t5 97.8995
R201 VP.n7 VP.t7 97.8995
R202 VP.n67 VP.t9 97.8995
R203 VP.n75 VP.t1 97.8995
R204 VP.n26 VP.t6 97.8995
R205 VP.n41 VP.t4 97.8995
R206 VP.n33 VP.t0 97.8995
R207 VP.n17 VP.t8 97.8995
R208 VP.n44 VP.n43 94.1189
R209 VP.n76 VP.n75 94.1189
R210 VP.n42 VP.n41 94.1189
R211 VP.n56 VP.n55 56.5193
R212 VP.n62 VP.n3 56.5193
R213 VP.n28 VP.n13 56.5193
R214 VP.n22 VP.n21 56.5193
R215 VP.n49 VP.n9 53.1199
R216 VP.n73 VP.n1 53.1199
R217 VP.n39 VP.n11 53.1199
R218 VP.n18 VP.n17 50.0611
R219 VP.n43 VP.n42 47.6814
R220 VP.n50 VP.n49 27.8669
R221 VP.n69 VP.n1 27.8669
R222 VP.n35 VP.n11 27.8669
R223 VP.n45 VP.n9 24.4675
R224 VP.n51 VP.n50 24.4675
R225 VP.n55 VP.n54 24.4675
R226 VP.n56 VP.n5 24.4675
R227 VP.n60 VP.n5 24.4675
R228 VP.n61 VP.n60 24.4675
R229 VP.n62 VP.n61 24.4675
R230 VP.n66 VP.n3 24.4675
R231 VP.n69 VP.n68 24.4675
R232 VP.n74 VP.n73 24.4675
R233 VP.n40 VP.n39 24.4675
R234 VP.n32 VP.n13 24.4675
R235 VP.n35 VP.n34 24.4675
R236 VP.n22 VP.n15 24.4675
R237 VP.n26 VP.n15 24.4675
R238 VP.n27 VP.n26 24.4675
R239 VP.n28 VP.n27 24.4675
R240 VP.n21 VP.n20 24.4675
R241 VP.n54 VP.n7 20.5528
R242 VP.n67 VP.n66 20.5528
R243 VP.n33 VP.n32 20.5528
R244 VP.n20 VP.n17 20.5528
R245 VP.n45 VP.n44 16.6381
R246 VP.n75 VP.n74 16.6381
R247 VP.n41 VP.n40 16.6381
R248 VP.n19 VP.n18 9.28282
R249 VP.n51 VP.n7 3.91522
R250 VP.n68 VP.n67 3.91522
R251 VP.n34 VP.n33 3.91522
R252 VP.n42 VP.n10 0.278367
R253 VP.n46 VP.n43 0.278367
R254 VP.n76 VP.n0 0.278367
R255 VP.n19 VP.n16 0.189894
R256 VP.n23 VP.n16 0.189894
R257 VP.n24 VP.n23 0.189894
R258 VP.n25 VP.n24 0.189894
R259 VP.n25 VP.n14 0.189894
R260 VP.n29 VP.n14 0.189894
R261 VP.n30 VP.n29 0.189894
R262 VP.n31 VP.n30 0.189894
R263 VP.n31 VP.n12 0.189894
R264 VP.n36 VP.n12 0.189894
R265 VP.n37 VP.n36 0.189894
R266 VP.n38 VP.n37 0.189894
R267 VP.n38 VP.n10 0.189894
R268 VP.n47 VP.n46 0.189894
R269 VP.n48 VP.n47 0.189894
R270 VP.n48 VP.n8 0.189894
R271 VP.n52 VP.n8 0.189894
R272 VP.n53 VP.n52 0.189894
R273 VP.n53 VP.n6 0.189894
R274 VP.n57 VP.n6 0.189894
R275 VP.n58 VP.n57 0.189894
R276 VP.n59 VP.n58 0.189894
R277 VP.n59 VP.n4 0.189894
R278 VP.n63 VP.n4 0.189894
R279 VP.n64 VP.n63 0.189894
R280 VP.n65 VP.n64 0.189894
R281 VP.n65 VP.n2 0.189894
R282 VP.n70 VP.n2 0.189894
R283 VP.n71 VP.n70 0.189894
R284 VP.n72 VP.n71 0.189894
R285 VP.n72 VP.n0 0.189894
R286 VP VP.n76 0.153454
R287 VDD1.n1 VDD1.t7 87.0322
R288 VDD1.n3 VDD1.t4 87.032
R289 VDD1.n5 VDD1.n4 82.6267
R290 VDD1.n7 VDD1.n6 81.1174
R291 VDD1.n1 VDD1.n0 81.1174
R292 VDD1.n3 VDD1.n2 81.1174
R293 VDD1.n7 VDD1.n5 42.5699
R294 VDD1.n6 VDD1.t9 3.82912
R295 VDD1.n6 VDD1.t5 3.82912
R296 VDD1.n0 VDD1.t1 3.82912
R297 VDD1.n0 VDD1.t3 3.82912
R298 VDD1.n4 VDD1.t0 3.82912
R299 VDD1.n4 VDD1.t8 3.82912
R300 VDD1.n2 VDD1.t2 3.82912
R301 VDD1.n2 VDD1.t6 3.82912
R302 VDD1 VDD1.n7 1.50697
R303 VDD1 VDD1.n1 0.580241
R304 VDD1.n5 VDD1.n3 0.466706
R305 B.n525 B.n524 585
R306 B.n526 B.n67 585
R307 B.n528 B.n527 585
R308 B.n529 B.n66 585
R309 B.n531 B.n530 585
R310 B.n532 B.n65 585
R311 B.n534 B.n533 585
R312 B.n535 B.n64 585
R313 B.n537 B.n536 585
R314 B.n538 B.n63 585
R315 B.n540 B.n539 585
R316 B.n541 B.n62 585
R317 B.n543 B.n542 585
R318 B.n544 B.n61 585
R319 B.n546 B.n545 585
R320 B.n547 B.n60 585
R321 B.n549 B.n548 585
R322 B.n550 B.n59 585
R323 B.n552 B.n551 585
R324 B.n553 B.n58 585
R325 B.n555 B.n554 585
R326 B.n556 B.n57 585
R327 B.n558 B.n557 585
R328 B.n559 B.n56 585
R329 B.n561 B.n560 585
R330 B.n562 B.n55 585
R331 B.n564 B.n563 585
R332 B.n565 B.n54 585
R333 B.n567 B.n566 585
R334 B.n568 B.n53 585
R335 B.n570 B.n569 585
R336 B.n572 B.n571 585
R337 B.n573 B.n49 585
R338 B.n575 B.n574 585
R339 B.n576 B.n48 585
R340 B.n578 B.n577 585
R341 B.n579 B.n47 585
R342 B.n581 B.n580 585
R343 B.n582 B.n46 585
R344 B.n584 B.n583 585
R345 B.n585 B.n43 585
R346 B.n588 B.n587 585
R347 B.n589 B.n42 585
R348 B.n591 B.n590 585
R349 B.n592 B.n41 585
R350 B.n594 B.n593 585
R351 B.n595 B.n40 585
R352 B.n597 B.n596 585
R353 B.n598 B.n39 585
R354 B.n600 B.n599 585
R355 B.n601 B.n38 585
R356 B.n603 B.n602 585
R357 B.n604 B.n37 585
R358 B.n606 B.n605 585
R359 B.n607 B.n36 585
R360 B.n609 B.n608 585
R361 B.n610 B.n35 585
R362 B.n612 B.n611 585
R363 B.n613 B.n34 585
R364 B.n615 B.n614 585
R365 B.n616 B.n33 585
R366 B.n618 B.n617 585
R367 B.n619 B.n32 585
R368 B.n621 B.n620 585
R369 B.n622 B.n31 585
R370 B.n624 B.n623 585
R371 B.n625 B.n30 585
R372 B.n627 B.n626 585
R373 B.n628 B.n29 585
R374 B.n630 B.n629 585
R375 B.n631 B.n28 585
R376 B.n633 B.n632 585
R377 B.n523 B.n68 585
R378 B.n522 B.n521 585
R379 B.n520 B.n69 585
R380 B.n519 B.n518 585
R381 B.n517 B.n70 585
R382 B.n516 B.n515 585
R383 B.n514 B.n71 585
R384 B.n513 B.n512 585
R385 B.n511 B.n72 585
R386 B.n510 B.n509 585
R387 B.n508 B.n73 585
R388 B.n507 B.n506 585
R389 B.n505 B.n74 585
R390 B.n504 B.n503 585
R391 B.n502 B.n75 585
R392 B.n501 B.n500 585
R393 B.n499 B.n76 585
R394 B.n498 B.n497 585
R395 B.n496 B.n77 585
R396 B.n495 B.n494 585
R397 B.n493 B.n78 585
R398 B.n492 B.n491 585
R399 B.n490 B.n79 585
R400 B.n489 B.n488 585
R401 B.n487 B.n80 585
R402 B.n486 B.n485 585
R403 B.n484 B.n81 585
R404 B.n483 B.n482 585
R405 B.n481 B.n82 585
R406 B.n480 B.n479 585
R407 B.n478 B.n83 585
R408 B.n477 B.n476 585
R409 B.n475 B.n84 585
R410 B.n474 B.n473 585
R411 B.n472 B.n85 585
R412 B.n471 B.n470 585
R413 B.n469 B.n86 585
R414 B.n468 B.n467 585
R415 B.n466 B.n87 585
R416 B.n465 B.n464 585
R417 B.n463 B.n88 585
R418 B.n462 B.n461 585
R419 B.n460 B.n89 585
R420 B.n459 B.n458 585
R421 B.n457 B.n90 585
R422 B.n456 B.n455 585
R423 B.n454 B.n91 585
R424 B.n453 B.n452 585
R425 B.n451 B.n92 585
R426 B.n450 B.n449 585
R427 B.n448 B.n93 585
R428 B.n447 B.n446 585
R429 B.n445 B.n94 585
R430 B.n444 B.n443 585
R431 B.n442 B.n95 585
R432 B.n441 B.n440 585
R433 B.n439 B.n96 585
R434 B.n438 B.n437 585
R435 B.n436 B.n97 585
R436 B.n435 B.n434 585
R437 B.n433 B.n98 585
R438 B.n432 B.n431 585
R439 B.n430 B.n99 585
R440 B.n429 B.n428 585
R441 B.n427 B.n100 585
R442 B.n426 B.n425 585
R443 B.n424 B.n101 585
R444 B.n423 B.n422 585
R445 B.n421 B.n102 585
R446 B.n420 B.n419 585
R447 B.n418 B.n103 585
R448 B.n417 B.n416 585
R449 B.n415 B.n104 585
R450 B.n414 B.n413 585
R451 B.n412 B.n105 585
R452 B.n411 B.n410 585
R453 B.n409 B.n106 585
R454 B.n408 B.n407 585
R455 B.n406 B.n107 585
R456 B.n405 B.n404 585
R457 B.n403 B.n108 585
R458 B.n402 B.n401 585
R459 B.n400 B.n109 585
R460 B.n399 B.n398 585
R461 B.n397 B.n110 585
R462 B.n396 B.n395 585
R463 B.n394 B.n111 585
R464 B.n393 B.n392 585
R465 B.n391 B.n112 585
R466 B.n390 B.n389 585
R467 B.n388 B.n113 585
R468 B.n387 B.n386 585
R469 B.n385 B.n114 585
R470 B.n384 B.n383 585
R471 B.n382 B.n115 585
R472 B.n381 B.n380 585
R473 B.n379 B.n116 585
R474 B.n378 B.n377 585
R475 B.n376 B.n117 585
R476 B.n375 B.n374 585
R477 B.n373 B.n118 585
R478 B.n372 B.n371 585
R479 B.n370 B.n119 585
R480 B.n261 B.n260 585
R481 B.n262 B.n159 585
R482 B.n264 B.n263 585
R483 B.n265 B.n158 585
R484 B.n267 B.n266 585
R485 B.n268 B.n157 585
R486 B.n270 B.n269 585
R487 B.n271 B.n156 585
R488 B.n273 B.n272 585
R489 B.n274 B.n155 585
R490 B.n276 B.n275 585
R491 B.n277 B.n154 585
R492 B.n279 B.n278 585
R493 B.n280 B.n153 585
R494 B.n282 B.n281 585
R495 B.n283 B.n152 585
R496 B.n285 B.n284 585
R497 B.n286 B.n151 585
R498 B.n288 B.n287 585
R499 B.n289 B.n150 585
R500 B.n291 B.n290 585
R501 B.n292 B.n149 585
R502 B.n294 B.n293 585
R503 B.n295 B.n148 585
R504 B.n297 B.n296 585
R505 B.n298 B.n147 585
R506 B.n300 B.n299 585
R507 B.n301 B.n146 585
R508 B.n303 B.n302 585
R509 B.n304 B.n145 585
R510 B.n306 B.n305 585
R511 B.n308 B.n307 585
R512 B.n309 B.n141 585
R513 B.n311 B.n310 585
R514 B.n312 B.n140 585
R515 B.n314 B.n313 585
R516 B.n315 B.n139 585
R517 B.n317 B.n316 585
R518 B.n318 B.n138 585
R519 B.n320 B.n319 585
R520 B.n321 B.n135 585
R521 B.n324 B.n323 585
R522 B.n325 B.n134 585
R523 B.n327 B.n326 585
R524 B.n328 B.n133 585
R525 B.n330 B.n329 585
R526 B.n331 B.n132 585
R527 B.n333 B.n332 585
R528 B.n334 B.n131 585
R529 B.n336 B.n335 585
R530 B.n337 B.n130 585
R531 B.n339 B.n338 585
R532 B.n340 B.n129 585
R533 B.n342 B.n341 585
R534 B.n343 B.n128 585
R535 B.n345 B.n344 585
R536 B.n346 B.n127 585
R537 B.n348 B.n347 585
R538 B.n349 B.n126 585
R539 B.n351 B.n350 585
R540 B.n352 B.n125 585
R541 B.n354 B.n353 585
R542 B.n355 B.n124 585
R543 B.n357 B.n356 585
R544 B.n358 B.n123 585
R545 B.n360 B.n359 585
R546 B.n361 B.n122 585
R547 B.n363 B.n362 585
R548 B.n364 B.n121 585
R549 B.n366 B.n365 585
R550 B.n367 B.n120 585
R551 B.n369 B.n368 585
R552 B.n259 B.n160 585
R553 B.n258 B.n257 585
R554 B.n256 B.n161 585
R555 B.n255 B.n254 585
R556 B.n253 B.n162 585
R557 B.n252 B.n251 585
R558 B.n250 B.n163 585
R559 B.n249 B.n248 585
R560 B.n247 B.n164 585
R561 B.n246 B.n245 585
R562 B.n244 B.n165 585
R563 B.n243 B.n242 585
R564 B.n241 B.n166 585
R565 B.n240 B.n239 585
R566 B.n238 B.n167 585
R567 B.n237 B.n236 585
R568 B.n235 B.n168 585
R569 B.n234 B.n233 585
R570 B.n232 B.n169 585
R571 B.n231 B.n230 585
R572 B.n229 B.n170 585
R573 B.n228 B.n227 585
R574 B.n226 B.n171 585
R575 B.n225 B.n224 585
R576 B.n223 B.n172 585
R577 B.n222 B.n221 585
R578 B.n220 B.n173 585
R579 B.n219 B.n218 585
R580 B.n217 B.n174 585
R581 B.n216 B.n215 585
R582 B.n214 B.n175 585
R583 B.n213 B.n212 585
R584 B.n211 B.n176 585
R585 B.n210 B.n209 585
R586 B.n208 B.n177 585
R587 B.n207 B.n206 585
R588 B.n205 B.n178 585
R589 B.n204 B.n203 585
R590 B.n202 B.n179 585
R591 B.n201 B.n200 585
R592 B.n199 B.n180 585
R593 B.n198 B.n197 585
R594 B.n196 B.n181 585
R595 B.n195 B.n194 585
R596 B.n193 B.n182 585
R597 B.n192 B.n191 585
R598 B.n190 B.n183 585
R599 B.n189 B.n188 585
R600 B.n187 B.n184 585
R601 B.n186 B.n185 585
R602 B.n2 B.n0 585
R603 B.n709 B.n1 585
R604 B.n708 B.n707 585
R605 B.n706 B.n3 585
R606 B.n705 B.n704 585
R607 B.n703 B.n4 585
R608 B.n702 B.n701 585
R609 B.n700 B.n5 585
R610 B.n699 B.n698 585
R611 B.n697 B.n6 585
R612 B.n696 B.n695 585
R613 B.n694 B.n7 585
R614 B.n693 B.n692 585
R615 B.n691 B.n8 585
R616 B.n690 B.n689 585
R617 B.n688 B.n9 585
R618 B.n687 B.n686 585
R619 B.n685 B.n10 585
R620 B.n684 B.n683 585
R621 B.n682 B.n11 585
R622 B.n681 B.n680 585
R623 B.n679 B.n12 585
R624 B.n678 B.n677 585
R625 B.n676 B.n13 585
R626 B.n675 B.n674 585
R627 B.n673 B.n14 585
R628 B.n672 B.n671 585
R629 B.n670 B.n15 585
R630 B.n669 B.n668 585
R631 B.n667 B.n16 585
R632 B.n666 B.n665 585
R633 B.n664 B.n17 585
R634 B.n663 B.n662 585
R635 B.n661 B.n18 585
R636 B.n660 B.n659 585
R637 B.n658 B.n19 585
R638 B.n657 B.n656 585
R639 B.n655 B.n20 585
R640 B.n654 B.n653 585
R641 B.n652 B.n21 585
R642 B.n651 B.n650 585
R643 B.n649 B.n22 585
R644 B.n648 B.n647 585
R645 B.n646 B.n23 585
R646 B.n645 B.n644 585
R647 B.n643 B.n24 585
R648 B.n642 B.n641 585
R649 B.n640 B.n25 585
R650 B.n639 B.n638 585
R651 B.n637 B.n26 585
R652 B.n636 B.n635 585
R653 B.n634 B.n27 585
R654 B.n711 B.n710 585
R655 B.n260 B.n259 482.89
R656 B.n632 B.n27 482.89
R657 B.n368 B.n119 482.89
R658 B.n524 B.n523 482.89
R659 B.n136 B.t6 305.021
R660 B.n142 B.t9 305.021
R661 B.n44 B.t0 305.021
R662 B.n50 B.t3 305.021
R663 B.n259 B.n258 163.367
R664 B.n258 B.n161 163.367
R665 B.n254 B.n161 163.367
R666 B.n254 B.n253 163.367
R667 B.n253 B.n252 163.367
R668 B.n252 B.n163 163.367
R669 B.n248 B.n163 163.367
R670 B.n248 B.n247 163.367
R671 B.n247 B.n246 163.367
R672 B.n246 B.n165 163.367
R673 B.n242 B.n165 163.367
R674 B.n242 B.n241 163.367
R675 B.n241 B.n240 163.367
R676 B.n240 B.n167 163.367
R677 B.n236 B.n167 163.367
R678 B.n236 B.n235 163.367
R679 B.n235 B.n234 163.367
R680 B.n234 B.n169 163.367
R681 B.n230 B.n169 163.367
R682 B.n230 B.n229 163.367
R683 B.n229 B.n228 163.367
R684 B.n228 B.n171 163.367
R685 B.n224 B.n171 163.367
R686 B.n224 B.n223 163.367
R687 B.n223 B.n222 163.367
R688 B.n222 B.n173 163.367
R689 B.n218 B.n173 163.367
R690 B.n218 B.n217 163.367
R691 B.n217 B.n216 163.367
R692 B.n216 B.n175 163.367
R693 B.n212 B.n175 163.367
R694 B.n212 B.n211 163.367
R695 B.n211 B.n210 163.367
R696 B.n210 B.n177 163.367
R697 B.n206 B.n177 163.367
R698 B.n206 B.n205 163.367
R699 B.n205 B.n204 163.367
R700 B.n204 B.n179 163.367
R701 B.n200 B.n179 163.367
R702 B.n200 B.n199 163.367
R703 B.n199 B.n198 163.367
R704 B.n198 B.n181 163.367
R705 B.n194 B.n181 163.367
R706 B.n194 B.n193 163.367
R707 B.n193 B.n192 163.367
R708 B.n192 B.n183 163.367
R709 B.n188 B.n183 163.367
R710 B.n188 B.n187 163.367
R711 B.n187 B.n186 163.367
R712 B.n186 B.n2 163.367
R713 B.n710 B.n2 163.367
R714 B.n710 B.n709 163.367
R715 B.n709 B.n708 163.367
R716 B.n708 B.n3 163.367
R717 B.n704 B.n3 163.367
R718 B.n704 B.n703 163.367
R719 B.n703 B.n702 163.367
R720 B.n702 B.n5 163.367
R721 B.n698 B.n5 163.367
R722 B.n698 B.n697 163.367
R723 B.n697 B.n696 163.367
R724 B.n696 B.n7 163.367
R725 B.n692 B.n7 163.367
R726 B.n692 B.n691 163.367
R727 B.n691 B.n690 163.367
R728 B.n690 B.n9 163.367
R729 B.n686 B.n9 163.367
R730 B.n686 B.n685 163.367
R731 B.n685 B.n684 163.367
R732 B.n684 B.n11 163.367
R733 B.n680 B.n11 163.367
R734 B.n680 B.n679 163.367
R735 B.n679 B.n678 163.367
R736 B.n678 B.n13 163.367
R737 B.n674 B.n13 163.367
R738 B.n674 B.n673 163.367
R739 B.n673 B.n672 163.367
R740 B.n672 B.n15 163.367
R741 B.n668 B.n15 163.367
R742 B.n668 B.n667 163.367
R743 B.n667 B.n666 163.367
R744 B.n666 B.n17 163.367
R745 B.n662 B.n17 163.367
R746 B.n662 B.n661 163.367
R747 B.n661 B.n660 163.367
R748 B.n660 B.n19 163.367
R749 B.n656 B.n19 163.367
R750 B.n656 B.n655 163.367
R751 B.n655 B.n654 163.367
R752 B.n654 B.n21 163.367
R753 B.n650 B.n21 163.367
R754 B.n650 B.n649 163.367
R755 B.n649 B.n648 163.367
R756 B.n648 B.n23 163.367
R757 B.n644 B.n23 163.367
R758 B.n644 B.n643 163.367
R759 B.n643 B.n642 163.367
R760 B.n642 B.n25 163.367
R761 B.n638 B.n25 163.367
R762 B.n638 B.n637 163.367
R763 B.n637 B.n636 163.367
R764 B.n636 B.n27 163.367
R765 B.n260 B.n159 163.367
R766 B.n264 B.n159 163.367
R767 B.n265 B.n264 163.367
R768 B.n266 B.n265 163.367
R769 B.n266 B.n157 163.367
R770 B.n270 B.n157 163.367
R771 B.n271 B.n270 163.367
R772 B.n272 B.n271 163.367
R773 B.n272 B.n155 163.367
R774 B.n276 B.n155 163.367
R775 B.n277 B.n276 163.367
R776 B.n278 B.n277 163.367
R777 B.n278 B.n153 163.367
R778 B.n282 B.n153 163.367
R779 B.n283 B.n282 163.367
R780 B.n284 B.n283 163.367
R781 B.n284 B.n151 163.367
R782 B.n288 B.n151 163.367
R783 B.n289 B.n288 163.367
R784 B.n290 B.n289 163.367
R785 B.n290 B.n149 163.367
R786 B.n294 B.n149 163.367
R787 B.n295 B.n294 163.367
R788 B.n296 B.n295 163.367
R789 B.n296 B.n147 163.367
R790 B.n300 B.n147 163.367
R791 B.n301 B.n300 163.367
R792 B.n302 B.n301 163.367
R793 B.n302 B.n145 163.367
R794 B.n306 B.n145 163.367
R795 B.n307 B.n306 163.367
R796 B.n307 B.n141 163.367
R797 B.n311 B.n141 163.367
R798 B.n312 B.n311 163.367
R799 B.n313 B.n312 163.367
R800 B.n313 B.n139 163.367
R801 B.n317 B.n139 163.367
R802 B.n318 B.n317 163.367
R803 B.n319 B.n318 163.367
R804 B.n319 B.n135 163.367
R805 B.n324 B.n135 163.367
R806 B.n325 B.n324 163.367
R807 B.n326 B.n325 163.367
R808 B.n326 B.n133 163.367
R809 B.n330 B.n133 163.367
R810 B.n331 B.n330 163.367
R811 B.n332 B.n331 163.367
R812 B.n332 B.n131 163.367
R813 B.n336 B.n131 163.367
R814 B.n337 B.n336 163.367
R815 B.n338 B.n337 163.367
R816 B.n338 B.n129 163.367
R817 B.n342 B.n129 163.367
R818 B.n343 B.n342 163.367
R819 B.n344 B.n343 163.367
R820 B.n344 B.n127 163.367
R821 B.n348 B.n127 163.367
R822 B.n349 B.n348 163.367
R823 B.n350 B.n349 163.367
R824 B.n350 B.n125 163.367
R825 B.n354 B.n125 163.367
R826 B.n355 B.n354 163.367
R827 B.n356 B.n355 163.367
R828 B.n356 B.n123 163.367
R829 B.n360 B.n123 163.367
R830 B.n361 B.n360 163.367
R831 B.n362 B.n361 163.367
R832 B.n362 B.n121 163.367
R833 B.n366 B.n121 163.367
R834 B.n367 B.n366 163.367
R835 B.n368 B.n367 163.367
R836 B.n372 B.n119 163.367
R837 B.n373 B.n372 163.367
R838 B.n374 B.n373 163.367
R839 B.n374 B.n117 163.367
R840 B.n378 B.n117 163.367
R841 B.n379 B.n378 163.367
R842 B.n380 B.n379 163.367
R843 B.n380 B.n115 163.367
R844 B.n384 B.n115 163.367
R845 B.n385 B.n384 163.367
R846 B.n386 B.n385 163.367
R847 B.n386 B.n113 163.367
R848 B.n390 B.n113 163.367
R849 B.n391 B.n390 163.367
R850 B.n392 B.n391 163.367
R851 B.n392 B.n111 163.367
R852 B.n396 B.n111 163.367
R853 B.n397 B.n396 163.367
R854 B.n398 B.n397 163.367
R855 B.n398 B.n109 163.367
R856 B.n402 B.n109 163.367
R857 B.n403 B.n402 163.367
R858 B.n404 B.n403 163.367
R859 B.n404 B.n107 163.367
R860 B.n408 B.n107 163.367
R861 B.n409 B.n408 163.367
R862 B.n410 B.n409 163.367
R863 B.n410 B.n105 163.367
R864 B.n414 B.n105 163.367
R865 B.n415 B.n414 163.367
R866 B.n416 B.n415 163.367
R867 B.n416 B.n103 163.367
R868 B.n420 B.n103 163.367
R869 B.n421 B.n420 163.367
R870 B.n422 B.n421 163.367
R871 B.n422 B.n101 163.367
R872 B.n426 B.n101 163.367
R873 B.n427 B.n426 163.367
R874 B.n428 B.n427 163.367
R875 B.n428 B.n99 163.367
R876 B.n432 B.n99 163.367
R877 B.n433 B.n432 163.367
R878 B.n434 B.n433 163.367
R879 B.n434 B.n97 163.367
R880 B.n438 B.n97 163.367
R881 B.n439 B.n438 163.367
R882 B.n440 B.n439 163.367
R883 B.n440 B.n95 163.367
R884 B.n444 B.n95 163.367
R885 B.n445 B.n444 163.367
R886 B.n446 B.n445 163.367
R887 B.n446 B.n93 163.367
R888 B.n450 B.n93 163.367
R889 B.n451 B.n450 163.367
R890 B.n452 B.n451 163.367
R891 B.n452 B.n91 163.367
R892 B.n456 B.n91 163.367
R893 B.n457 B.n456 163.367
R894 B.n458 B.n457 163.367
R895 B.n458 B.n89 163.367
R896 B.n462 B.n89 163.367
R897 B.n463 B.n462 163.367
R898 B.n464 B.n463 163.367
R899 B.n464 B.n87 163.367
R900 B.n468 B.n87 163.367
R901 B.n469 B.n468 163.367
R902 B.n470 B.n469 163.367
R903 B.n470 B.n85 163.367
R904 B.n474 B.n85 163.367
R905 B.n475 B.n474 163.367
R906 B.n476 B.n475 163.367
R907 B.n476 B.n83 163.367
R908 B.n480 B.n83 163.367
R909 B.n481 B.n480 163.367
R910 B.n482 B.n481 163.367
R911 B.n482 B.n81 163.367
R912 B.n486 B.n81 163.367
R913 B.n487 B.n486 163.367
R914 B.n488 B.n487 163.367
R915 B.n488 B.n79 163.367
R916 B.n492 B.n79 163.367
R917 B.n493 B.n492 163.367
R918 B.n494 B.n493 163.367
R919 B.n494 B.n77 163.367
R920 B.n498 B.n77 163.367
R921 B.n499 B.n498 163.367
R922 B.n500 B.n499 163.367
R923 B.n500 B.n75 163.367
R924 B.n504 B.n75 163.367
R925 B.n505 B.n504 163.367
R926 B.n506 B.n505 163.367
R927 B.n506 B.n73 163.367
R928 B.n510 B.n73 163.367
R929 B.n511 B.n510 163.367
R930 B.n512 B.n511 163.367
R931 B.n512 B.n71 163.367
R932 B.n516 B.n71 163.367
R933 B.n517 B.n516 163.367
R934 B.n518 B.n517 163.367
R935 B.n518 B.n69 163.367
R936 B.n522 B.n69 163.367
R937 B.n523 B.n522 163.367
R938 B.n632 B.n631 163.367
R939 B.n631 B.n630 163.367
R940 B.n630 B.n29 163.367
R941 B.n626 B.n29 163.367
R942 B.n626 B.n625 163.367
R943 B.n625 B.n624 163.367
R944 B.n624 B.n31 163.367
R945 B.n620 B.n31 163.367
R946 B.n620 B.n619 163.367
R947 B.n619 B.n618 163.367
R948 B.n618 B.n33 163.367
R949 B.n614 B.n33 163.367
R950 B.n614 B.n613 163.367
R951 B.n613 B.n612 163.367
R952 B.n612 B.n35 163.367
R953 B.n608 B.n35 163.367
R954 B.n608 B.n607 163.367
R955 B.n607 B.n606 163.367
R956 B.n606 B.n37 163.367
R957 B.n602 B.n37 163.367
R958 B.n602 B.n601 163.367
R959 B.n601 B.n600 163.367
R960 B.n600 B.n39 163.367
R961 B.n596 B.n39 163.367
R962 B.n596 B.n595 163.367
R963 B.n595 B.n594 163.367
R964 B.n594 B.n41 163.367
R965 B.n590 B.n41 163.367
R966 B.n590 B.n589 163.367
R967 B.n589 B.n588 163.367
R968 B.n588 B.n43 163.367
R969 B.n583 B.n43 163.367
R970 B.n583 B.n582 163.367
R971 B.n582 B.n581 163.367
R972 B.n581 B.n47 163.367
R973 B.n577 B.n47 163.367
R974 B.n577 B.n576 163.367
R975 B.n576 B.n575 163.367
R976 B.n575 B.n49 163.367
R977 B.n571 B.n49 163.367
R978 B.n571 B.n570 163.367
R979 B.n570 B.n53 163.367
R980 B.n566 B.n53 163.367
R981 B.n566 B.n565 163.367
R982 B.n565 B.n564 163.367
R983 B.n564 B.n55 163.367
R984 B.n560 B.n55 163.367
R985 B.n560 B.n559 163.367
R986 B.n559 B.n558 163.367
R987 B.n558 B.n57 163.367
R988 B.n554 B.n57 163.367
R989 B.n554 B.n553 163.367
R990 B.n553 B.n552 163.367
R991 B.n552 B.n59 163.367
R992 B.n548 B.n59 163.367
R993 B.n548 B.n547 163.367
R994 B.n547 B.n546 163.367
R995 B.n546 B.n61 163.367
R996 B.n542 B.n61 163.367
R997 B.n542 B.n541 163.367
R998 B.n541 B.n540 163.367
R999 B.n540 B.n63 163.367
R1000 B.n536 B.n63 163.367
R1001 B.n536 B.n535 163.367
R1002 B.n535 B.n534 163.367
R1003 B.n534 B.n65 163.367
R1004 B.n530 B.n65 163.367
R1005 B.n530 B.n529 163.367
R1006 B.n529 B.n528 163.367
R1007 B.n528 B.n67 163.367
R1008 B.n524 B.n67 163.367
R1009 B.n136 B.t8 161.724
R1010 B.n50 B.t4 161.724
R1011 B.n142 B.t11 161.714
R1012 B.n44 B.t1 161.714
R1013 B.n137 B.t7 114.79
R1014 B.n51 B.t5 114.79
R1015 B.n143 B.t10 114.781
R1016 B.n45 B.t2 114.781
R1017 B.n322 B.n137 59.5399
R1018 B.n144 B.n143 59.5399
R1019 B.n586 B.n45 59.5399
R1020 B.n52 B.n51 59.5399
R1021 B.n137 B.n136 46.9338
R1022 B.n143 B.n142 46.9338
R1023 B.n45 B.n44 46.9338
R1024 B.n51 B.n50 46.9338
R1025 B.n634 B.n633 31.3761
R1026 B.n525 B.n68 31.3761
R1027 B.n370 B.n369 31.3761
R1028 B.n261 B.n160 31.3761
R1029 B B.n711 18.0485
R1030 B.n633 B.n28 10.6151
R1031 B.n629 B.n28 10.6151
R1032 B.n629 B.n628 10.6151
R1033 B.n628 B.n627 10.6151
R1034 B.n627 B.n30 10.6151
R1035 B.n623 B.n30 10.6151
R1036 B.n623 B.n622 10.6151
R1037 B.n622 B.n621 10.6151
R1038 B.n621 B.n32 10.6151
R1039 B.n617 B.n32 10.6151
R1040 B.n617 B.n616 10.6151
R1041 B.n616 B.n615 10.6151
R1042 B.n615 B.n34 10.6151
R1043 B.n611 B.n34 10.6151
R1044 B.n611 B.n610 10.6151
R1045 B.n610 B.n609 10.6151
R1046 B.n609 B.n36 10.6151
R1047 B.n605 B.n36 10.6151
R1048 B.n605 B.n604 10.6151
R1049 B.n604 B.n603 10.6151
R1050 B.n603 B.n38 10.6151
R1051 B.n599 B.n38 10.6151
R1052 B.n599 B.n598 10.6151
R1053 B.n598 B.n597 10.6151
R1054 B.n597 B.n40 10.6151
R1055 B.n593 B.n40 10.6151
R1056 B.n593 B.n592 10.6151
R1057 B.n592 B.n591 10.6151
R1058 B.n591 B.n42 10.6151
R1059 B.n587 B.n42 10.6151
R1060 B.n585 B.n584 10.6151
R1061 B.n584 B.n46 10.6151
R1062 B.n580 B.n46 10.6151
R1063 B.n580 B.n579 10.6151
R1064 B.n579 B.n578 10.6151
R1065 B.n578 B.n48 10.6151
R1066 B.n574 B.n48 10.6151
R1067 B.n574 B.n573 10.6151
R1068 B.n573 B.n572 10.6151
R1069 B.n569 B.n568 10.6151
R1070 B.n568 B.n567 10.6151
R1071 B.n567 B.n54 10.6151
R1072 B.n563 B.n54 10.6151
R1073 B.n563 B.n562 10.6151
R1074 B.n562 B.n561 10.6151
R1075 B.n561 B.n56 10.6151
R1076 B.n557 B.n56 10.6151
R1077 B.n557 B.n556 10.6151
R1078 B.n556 B.n555 10.6151
R1079 B.n555 B.n58 10.6151
R1080 B.n551 B.n58 10.6151
R1081 B.n551 B.n550 10.6151
R1082 B.n550 B.n549 10.6151
R1083 B.n549 B.n60 10.6151
R1084 B.n545 B.n60 10.6151
R1085 B.n545 B.n544 10.6151
R1086 B.n544 B.n543 10.6151
R1087 B.n543 B.n62 10.6151
R1088 B.n539 B.n62 10.6151
R1089 B.n539 B.n538 10.6151
R1090 B.n538 B.n537 10.6151
R1091 B.n537 B.n64 10.6151
R1092 B.n533 B.n64 10.6151
R1093 B.n533 B.n532 10.6151
R1094 B.n532 B.n531 10.6151
R1095 B.n531 B.n66 10.6151
R1096 B.n527 B.n66 10.6151
R1097 B.n527 B.n526 10.6151
R1098 B.n526 B.n525 10.6151
R1099 B.n371 B.n370 10.6151
R1100 B.n371 B.n118 10.6151
R1101 B.n375 B.n118 10.6151
R1102 B.n376 B.n375 10.6151
R1103 B.n377 B.n376 10.6151
R1104 B.n377 B.n116 10.6151
R1105 B.n381 B.n116 10.6151
R1106 B.n382 B.n381 10.6151
R1107 B.n383 B.n382 10.6151
R1108 B.n383 B.n114 10.6151
R1109 B.n387 B.n114 10.6151
R1110 B.n388 B.n387 10.6151
R1111 B.n389 B.n388 10.6151
R1112 B.n389 B.n112 10.6151
R1113 B.n393 B.n112 10.6151
R1114 B.n394 B.n393 10.6151
R1115 B.n395 B.n394 10.6151
R1116 B.n395 B.n110 10.6151
R1117 B.n399 B.n110 10.6151
R1118 B.n400 B.n399 10.6151
R1119 B.n401 B.n400 10.6151
R1120 B.n401 B.n108 10.6151
R1121 B.n405 B.n108 10.6151
R1122 B.n406 B.n405 10.6151
R1123 B.n407 B.n406 10.6151
R1124 B.n407 B.n106 10.6151
R1125 B.n411 B.n106 10.6151
R1126 B.n412 B.n411 10.6151
R1127 B.n413 B.n412 10.6151
R1128 B.n413 B.n104 10.6151
R1129 B.n417 B.n104 10.6151
R1130 B.n418 B.n417 10.6151
R1131 B.n419 B.n418 10.6151
R1132 B.n419 B.n102 10.6151
R1133 B.n423 B.n102 10.6151
R1134 B.n424 B.n423 10.6151
R1135 B.n425 B.n424 10.6151
R1136 B.n425 B.n100 10.6151
R1137 B.n429 B.n100 10.6151
R1138 B.n430 B.n429 10.6151
R1139 B.n431 B.n430 10.6151
R1140 B.n431 B.n98 10.6151
R1141 B.n435 B.n98 10.6151
R1142 B.n436 B.n435 10.6151
R1143 B.n437 B.n436 10.6151
R1144 B.n437 B.n96 10.6151
R1145 B.n441 B.n96 10.6151
R1146 B.n442 B.n441 10.6151
R1147 B.n443 B.n442 10.6151
R1148 B.n443 B.n94 10.6151
R1149 B.n447 B.n94 10.6151
R1150 B.n448 B.n447 10.6151
R1151 B.n449 B.n448 10.6151
R1152 B.n449 B.n92 10.6151
R1153 B.n453 B.n92 10.6151
R1154 B.n454 B.n453 10.6151
R1155 B.n455 B.n454 10.6151
R1156 B.n455 B.n90 10.6151
R1157 B.n459 B.n90 10.6151
R1158 B.n460 B.n459 10.6151
R1159 B.n461 B.n460 10.6151
R1160 B.n461 B.n88 10.6151
R1161 B.n465 B.n88 10.6151
R1162 B.n466 B.n465 10.6151
R1163 B.n467 B.n466 10.6151
R1164 B.n467 B.n86 10.6151
R1165 B.n471 B.n86 10.6151
R1166 B.n472 B.n471 10.6151
R1167 B.n473 B.n472 10.6151
R1168 B.n473 B.n84 10.6151
R1169 B.n477 B.n84 10.6151
R1170 B.n478 B.n477 10.6151
R1171 B.n479 B.n478 10.6151
R1172 B.n479 B.n82 10.6151
R1173 B.n483 B.n82 10.6151
R1174 B.n484 B.n483 10.6151
R1175 B.n485 B.n484 10.6151
R1176 B.n485 B.n80 10.6151
R1177 B.n489 B.n80 10.6151
R1178 B.n490 B.n489 10.6151
R1179 B.n491 B.n490 10.6151
R1180 B.n491 B.n78 10.6151
R1181 B.n495 B.n78 10.6151
R1182 B.n496 B.n495 10.6151
R1183 B.n497 B.n496 10.6151
R1184 B.n497 B.n76 10.6151
R1185 B.n501 B.n76 10.6151
R1186 B.n502 B.n501 10.6151
R1187 B.n503 B.n502 10.6151
R1188 B.n503 B.n74 10.6151
R1189 B.n507 B.n74 10.6151
R1190 B.n508 B.n507 10.6151
R1191 B.n509 B.n508 10.6151
R1192 B.n509 B.n72 10.6151
R1193 B.n513 B.n72 10.6151
R1194 B.n514 B.n513 10.6151
R1195 B.n515 B.n514 10.6151
R1196 B.n515 B.n70 10.6151
R1197 B.n519 B.n70 10.6151
R1198 B.n520 B.n519 10.6151
R1199 B.n521 B.n520 10.6151
R1200 B.n521 B.n68 10.6151
R1201 B.n262 B.n261 10.6151
R1202 B.n263 B.n262 10.6151
R1203 B.n263 B.n158 10.6151
R1204 B.n267 B.n158 10.6151
R1205 B.n268 B.n267 10.6151
R1206 B.n269 B.n268 10.6151
R1207 B.n269 B.n156 10.6151
R1208 B.n273 B.n156 10.6151
R1209 B.n274 B.n273 10.6151
R1210 B.n275 B.n274 10.6151
R1211 B.n275 B.n154 10.6151
R1212 B.n279 B.n154 10.6151
R1213 B.n280 B.n279 10.6151
R1214 B.n281 B.n280 10.6151
R1215 B.n281 B.n152 10.6151
R1216 B.n285 B.n152 10.6151
R1217 B.n286 B.n285 10.6151
R1218 B.n287 B.n286 10.6151
R1219 B.n287 B.n150 10.6151
R1220 B.n291 B.n150 10.6151
R1221 B.n292 B.n291 10.6151
R1222 B.n293 B.n292 10.6151
R1223 B.n293 B.n148 10.6151
R1224 B.n297 B.n148 10.6151
R1225 B.n298 B.n297 10.6151
R1226 B.n299 B.n298 10.6151
R1227 B.n299 B.n146 10.6151
R1228 B.n303 B.n146 10.6151
R1229 B.n304 B.n303 10.6151
R1230 B.n305 B.n304 10.6151
R1231 B.n309 B.n308 10.6151
R1232 B.n310 B.n309 10.6151
R1233 B.n310 B.n140 10.6151
R1234 B.n314 B.n140 10.6151
R1235 B.n315 B.n314 10.6151
R1236 B.n316 B.n315 10.6151
R1237 B.n316 B.n138 10.6151
R1238 B.n320 B.n138 10.6151
R1239 B.n321 B.n320 10.6151
R1240 B.n323 B.n134 10.6151
R1241 B.n327 B.n134 10.6151
R1242 B.n328 B.n327 10.6151
R1243 B.n329 B.n328 10.6151
R1244 B.n329 B.n132 10.6151
R1245 B.n333 B.n132 10.6151
R1246 B.n334 B.n333 10.6151
R1247 B.n335 B.n334 10.6151
R1248 B.n335 B.n130 10.6151
R1249 B.n339 B.n130 10.6151
R1250 B.n340 B.n339 10.6151
R1251 B.n341 B.n340 10.6151
R1252 B.n341 B.n128 10.6151
R1253 B.n345 B.n128 10.6151
R1254 B.n346 B.n345 10.6151
R1255 B.n347 B.n346 10.6151
R1256 B.n347 B.n126 10.6151
R1257 B.n351 B.n126 10.6151
R1258 B.n352 B.n351 10.6151
R1259 B.n353 B.n352 10.6151
R1260 B.n353 B.n124 10.6151
R1261 B.n357 B.n124 10.6151
R1262 B.n358 B.n357 10.6151
R1263 B.n359 B.n358 10.6151
R1264 B.n359 B.n122 10.6151
R1265 B.n363 B.n122 10.6151
R1266 B.n364 B.n363 10.6151
R1267 B.n365 B.n364 10.6151
R1268 B.n365 B.n120 10.6151
R1269 B.n369 B.n120 10.6151
R1270 B.n257 B.n160 10.6151
R1271 B.n257 B.n256 10.6151
R1272 B.n256 B.n255 10.6151
R1273 B.n255 B.n162 10.6151
R1274 B.n251 B.n162 10.6151
R1275 B.n251 B.n250 10.6151
R1276 B.n250 B.n249 10.6151
R1277 B.n249 B.n164 10.6151
R1278 B.n245 B.n164 10.6151
R1279 B.n245 B.n244 10.6151
R1280 B.n244 B.n243 10.6151
R1281 B.n243 B.n166 10.6151
R1282 B.n239 B.n166 10.6151
R1283 B.n239 B.n238 10.6151
R1284 B.n238 B.n237 10.6151
R1285 B.n237 B.n168 10.6151
R1286 B.n233 B.n168 10.6151
R1287 B.n233 B.n232 10.6151
R1288 B.n232 B.n231 10.6151
R1289 B.n231 B.n170 10.6151
R1290 B.n227 B.n170 10.6151
R1291 B.n227 B.n226 10.6151
R1292 B.n226 B.n225 10.6151
R1293 B.n225 B.n172 10.6151
R1294 B.n221 B.n172 10.6151
R1295 B.n221 B.n220 10.6151
R1296 B.n220 B.n219 10.6151
R1297 B.n219 B.n174 10.6151
R1298 B.n215 B.n174 10.6151
R1299 B.n215 B.n214 10.6151
R1300 B.n214 B.n213 10.6151
R1301 B.n213 B.n176 10.6151
R1302 B.n209 B.n176 10.6151
R1303 B.n209 B.n208 10.6151
R1304 B.n208 B.n207 10.6151
R1305 B.n207 B.n178 10.6151
R1306 B.n203 B.n178 10.6151
R1307 B.n203 B.n202 10.6151
R1308 B.n202 B.n201 10.6151
R1309 B.n201 B.n180 10.6151
R1310 B.n197 B.n180 10.6151
R1311 B.n197 B.n196 10.6151
R1312 B.n196 B.n195 10.6151
R1313 B.n195 B.n182 10.6151
R1314 B.n191 B.n182 10.6151
R1315 B.n191 B.n190 10.6151
R1316 B.n190 B.n189 10.6151
R1317 B.n189 B.n184 10.6151
R1318 B.n185 B.n184 10.6151
R1319 B.n185 B.n0 10.6151
R1320 B.n707 B.n1 10.6151
R1321 B.n707 B.n706 10.6151
R1322 B.n706 B.n705 10.6151
R1323 B.n705 B.n4 10.6151
R1324 B.n701 B.n4 10.6151
R1325 B.n701 B.n700 10.6151
R1326 B.n700 B.n699 10.6151
R1327 B.n699 B.n6 10.6151
R1328 B.n695 B.n6 10.6151
R1329 B.n695 B.n694 10.6151
R1330 B.n694 B.n693 10.6151
R1331 B.n693 B.n8 10.6151
R1332 B.n689 B.n8 10.6151
R1333 B.n689 B.n688 10.6151
R1334 B.n688 B.n687 10.6151
R1335 B.n687 B.n10 10.6151
R1336 B.n683 B.n10 10.6151
R1337 B.n683 B.n682 10.6151
R1338 B.n682 B.n681 10.6151
R1339 B.n681 B.n12 10.6151
R1340 B.n677 B.n12 10.6151
R1341 B.n677 B.n676 10.6151
R1342 B.n676 B.n675 10.6151
R1343 B.n675 B.n14 10.6151
R1344 B.n671 B.n14 10.6151
R1345 B.n671 B.n670 10.6151
R1346 B.n670 B.n669 10.6151
R1347 B.n669 B.n16 10.6151
R1348 B.n665 B.n16 10.6151
R1349 B.n665 B.n664 10.6151
R1350 B.n664 B.n663 10.6151
R1351 B.n663 B.n18 10.6151
R1352 B.n659 B.n18 10.6151
R1353 B.n659 B.n658 10.6151
R1354 B.n658 B.n657 10.6151
R1355 B.n657 B.n20 10.6151
R1356 B.n653 B.n20 10.6151
R1357 B.n653 B.n652 10.6151
R1358 B.n652 B.n651 10.6151
R1359 B.n651 B.n22 10.6151
R1360 B.n647 B.n22 10.6151
R1361 B.n647 B.n646 10.6151
R1362 B.n646 B.n645 10.6151
R1363 B.n645 B.n24 10.6151
R1364 B.n641 B.n24 10.6151
R1365 B.n641 B.n640 10.6151
R1366 B.n640 B.n639 10.6151
R1367 B.n639 B.n26 10.6151
R1368 B.n635 B.n26 10.6151
R1369 B.n635 B.n634 10.6151
R1370 B.n587 B.n586 9.36635
R1371 B.n569 B.n52 9.36635
R1372 B.n305 B.n144 9.36635
R1373 B.n323 B.n322 9.36635
R1374 B.n711 B.n0 2.81026
R1375 B.n711 B.n1 2.81026
R1376 B.n586 B.n585 1.24928
R1377 B.n572 B.n52 1.24928
R1378 B.n308 B.n144 1.24928
R1379 B.n322 B.n321 1.24928
C0 VDD1 VTAIL 8.60097f
C1 VDD2 VTAIL 8.648849f
C2 w_n3874_n2666# VTAIL 2.64876f
C3 VP VTAIL 7.92701f
C4 B VN 1.11243f
C5 VDD1 VN 0.152274f
C6 VDD2 VN 7.33348f
C7 w_n3874_n2666# VN 8.06795f
C8 VP VN 6.99902f
C9 B VDD1 2.00619f
C10 B VDD2 2.10424f
C11 B w_n3874_n2666# 8.70504f
C12 B VP 1.95511f
C13 VN VTAIL 7.91274f
C14 B VTAIL 2.75238f
C15 VDD2 VDD1 1.84265f
C16 w_n3874_n2666# VDD1 2.34996f
C17 VP VDD1 7.69634f
C18 w_n3874_n2666# VDD2 2.4671f
C19 VP VDD2 0.5183f
C20 w_n3874_n2666# VP 8.57076f
C21 VDD2 VSUBS 1.838412f
C22 VDD1 VSUBS 1.640555f
C23 VTAIL VSUBS 1.062329f
C24 VN VSUBS 6.746f
C25 VP VSUBS 3.463377f
C26 B VSUBS 4.436697f
C27 w_n3874_n2666# VSUBS 0.127981p
C28 B.n0 VSUBS 0.006055f
C29 B.n1 VSUBS 0.006055f
C30 B.n2 VSUBS 0.009576f
C31 B.n3 VSUBS 0.009576f
C32 B.n4 VSUBS 0.009576f
C33 B.n5 VSUBS 0.009576f
C34 B.n6 VSUBS 0.009576f
C35 B.n7 VSUBS 0.009576f
C36 B.n8 VSUBS 0.009576f
C37 B.n9 VSUBS 0.009576f
C38 B.n10 VSUBS 0.009576f
C39 B.n11 VSUBS 0.009576f
C40 B.n12 VSUBS 0.009576f
C41 B.n13 VSUBS 0.009576f
C42 B.n14 VSUBS 0.009576f
C43 B.n15 VSUBS 0.009576f
C44 B.n16 VSUBS 0.009576f
C45 B.n17 VSUBS 0.009576f
C46 B.n18 VSUBS 0.009576f
C47 B.n19 VSUBS 0.009576f
C48 B.n20 VSUBS 0.009576f
C49 B.n21 VSUBS 0.009576f
C50 B.n22 VSUBS 0.009576f
C51 B.n23 VSUBS 0.009576f
C52 B.n24 VSUBS 0.009576f
C53 B.n25 VSUBS 0.009576f
C54 B.n26 VSUBS 0.009576f
C55 B.n27 VSUBS 0.021526f
C56 B.n28 VSUBS 0.009576f
C57 B.n29 VSUBS 0.009576f
C58 B.n30 VSUBS 0.009576f
C59 B.n31 VSUBS 0.009576f
C60 B.n32 VSUBS 0.009576f
C61 B.n33 VSUBS 0.009576f
C62 B.n34 VSUBS 0.009576f
C63 B.n35 VSUBS 0.009576f
C64 B.n36 VSUBS 0.009576f
C65 B.n37 VSUBS 0.009576f
C66 B.n38 VSUBS 0.009576f
C67 B.n39 VSUBS 0.009576f
C68 B.n40 VSUBS 0.009576f
C69 B.n41 VSUBS 0.009576f
C70 B.n42 VSUBS 0.009576f
C71 B.n43 VSUBS 0.009576f
C72 B.t2 VSUBS 0.361714f
C73 B.t1 VSUBS 0.385314f
C74 B.t0 VSUBS 1.11287f
C75 B.n44 VSUBS 0.198654f
C76 B.n45 VSUBS 0.094975f
C77 B.n46 VSUBS 0.009576f
C78 B.n47 VSUBS 0.009576f
C79 B.n48 VSUBS 0.009576f
C80 B.n49 VSUBS 0.009576f
C81 B.t5 VSUBS 0.36171f
C82 B.t4 VSUBS 0.38531f
C83 B.t3 VSUBS 1.11287f
C84 B.n50 VSUBS 0.198658f
C85 B.n51 VSUBS 0.094978f
C86 B.n52 VSUBS 0.022186f
C87 B.n53 VSUBS 0.009576f
C88 B.n54 VSUBS 0.009576f
C89 B.n55 VSUBS 0.009576f
C90 B.n56 VSUBS 0.009576f
C91 B.n57 VSUBS 0.009576f
C92 B.n58 VSUBS 0.009576f
C93 B.n59 VSUBS 0.009576f
C94 B.n60 VSUBS 0.009576f
C95 B.n61 VSUBS 0.009576f
C96 B.n62 VSUBS 0.009576f
C97 B.n63 VSUBS 0.009576f
C98 B.n64 VSUBS 0.009576f
C99 B.n65 VSUBS 0.009576f
C100 B.n66 VSUBS 0.009576f
C101 B.n67 VSUBS 0.009576f
C102 B.n68 VSUBS 0.022703f
C103 B.n69 VSUBS 0.009576f
C104 B.n70 VSUBS 0.009576f
C105 B.n71 VSUBS 0.009576f
C106 B.n72 VSUBS 0.009576f
C107 B.n73 VSUBS 0.009576f
C108 B.n74 VSUBS 0.009576f
C109 B.n75 VSUBS 0.009576f
C110 B.n76 VSUBS 0.009576f
C111 B.n77 VSUBS 0.009576f
C112 B.n78 VSUBS 0.009576f
C113 B.n79 VSUBS 0.009576f
C114 B.n80 VSUBS 0.009576f
C115 B.n81 VSUBS 0.009576f
C116 B.n82 VSUBS 0.009576f
C117 B.n83 VSUBS 0.009576f
C118 B.n84 VSUBS 0.009576f
C119 B.n85 VSUBS 0.009576f
C120 B.n86 VSUBS 0.009576f
C121 B.n87 VSUBS 0.009576f
C122 B.n88 VSUBS 0.009576f
C123 B.n89 VSUBS 0.009576f
C124 B.n90 VSUBS 0.009576f
C125 B.n91 VSUBS 0.009576f
C126 B.n92 VSUBS 0.009576f
C127 B.n93 VSUBS 0.009576f
C128 B.n94 VSUBS 0.009576f
C129 B.n95 VSUBS 0.009576f
C130 B.n96 VSUBS 0.009576f
C131 B.n97 VSUBS 0.009576f
C132 B.n98 VSUBS 0.009576f
C133 B.n99 VSUBS 0.009576f
C134 B.n100 VSUBS 0.009576f
C135 B.n101 VSUBS 0.009576f
C136 B.n102 VSUBS 0.009576f
C137 B.n103 VSUBS 0.009576f
C138 B.n104 VSUBS 0.009576f
C139 B.n105 VSUBS 0.009576f
C140 B.n106 VSUBS 0.009576f
C141 B.n107 VSUBS 0.009576f
C142 B.n108 VSUBS 0.009576f
C143 B.n109 VSUBS 0.009576f
C144 B.n110 VSUBS 0.009576f
C145 B.n111 VSUBS 0.009576f
C146 B.n112 VSUBS 0.009576f
C147 B.n113 VSUBS 0.009576f
C148 B.n114 VSUBS 0.009576f
C149 B.n115 VSUBS 0.009576f
C150 B.n116 VSUBS 0.009576f
C151 B.n117 VSUBS 0.009576f
C152 B.n118 VSUBS 0.009576f
C153 B.n119 VSUBS 0.021526f
C154 B.n120 VSUBS 0.009576f
C155 B.n121 VSUBS 0.009576f
C156 B.n122 VSUBS 0.009576f
C157 B.n123 VSUBS 0.009576f
C158 B.n124 VSUBS 0.009576f
C159 B.n125 VSUBS 0.009576f
C160 B.n126 VSUBS 0.009576f
C161 B.n127 VSUBS 0.009576f
C162 B.n128 VSUBS 0.009576f
C163 B.n129 VSUBS 0.009576f
C164 B.n130 VSUBS 0.009576f
C165 B.n131 VSUBS 0.009576f
C166 B.n132 VSUBS 0.009576f
C167 B.n133 VSUBS 0.009576f
C168 B.n134 VSUBS 0.009576f
C169 B.n135 VSUBS 0.009576f
C170 B.t7 VSUBS 0.36171f
C171 B.t8 VSUBS 0.38531f
C172 B.t6 VSUBS 1.11287f
C173 B.n136 VSUBS 0.198658f
C174 B.n137 VSUBS 0.094978f
C175 B.n138 VSUBS 0.009576f
C176 B.n139 VSUBS 0.009576f
C177 B.n140 VSUBS 0.009576f
C178 B.n141 VSUBS 0.009576f
C179 B.t10 VSUBS 0.361714f
C180 B.t11 VSUBS 0.385314f
C181 B.t9 VSUBS 1.11287f
C182 B.n142 VSUBS 0.198654f
C183 B.n143 VSUBS 0.094975f
C184 B.n144 VSUBS 0.022186f
C185 B.n145 VSUBS 0.009576f
C186 B.n146 VSUBS 0.009576f
C187 B.n147 VSUBS 0.009576f
C188 B.n148 VSUBS 0.009576f
C189 B.n149 VSUBS 0.009576f
C190 B.n150 VSUBS 0.009576f
C191 B.n151 VSUBS 0.009576f
C192 B.n152 VSUBS 0.009576f
C193 B.n153 VSUBS 0.009576f
C194 B.n154 VSUBS 0.009576f
C195 B.n155 VSUBS 0.009576f
C196 B.n156 VSUBS 0.009576f
C197 B.n157 VSUBS 0.009576f
C198 B.n158 VSUBS 0.009576f
C199 B.n159 VSUBS 0.009576f
C200 B.n160 VSUBS 0.021526f
C201 B.n161 VSUBS 0.009576f
C202 B.n162 VSUBS 0.009576f
C203 B.n163 VSUBS 0.009576f
C204 B.n164 VSUBS 0.009576f
C205 B.n165 VSUBS 0.009576f
C206 B.n166 VSUBS 0.009576f
C207 B.n167 VSUBS 0.009576f
C208 B.n168 VSUBS 0.009576f
C209 B.n169 VSUBS 0.009576f
C210 B.n170 VSUBS 0.009576f
C211 B.n171 VSUBS 0.009576f
C212 B.n172 VSUBS 0.009576f
C213 B.n173 VSUBS 0.009576f
C214 B.n174 VSUBS 0.009576f
C215 B.n175 VSUBS 0.009576f
C216 B.n176 VSUBS 0.009576f
C217 B.n177 VSUBS 0.009576f
C218 B.n178 VSUBS 0.009576f
C219 B.n179 VSUBS 0.009576f
C220 B.n180 VSUBS 0.009576f
C221 B.n181 VSUBS 0.009576f
C222 B.n182 VSUBS 0.009576f
C223 B.n183 VSUBS 0.009576f
C224 B.n184 VSUBS 0.009576f
C225 B.n185 VSUBS 0.009576f
C226 B.n186 VSUBS 0.009576f
C227 B.n187 VSUBS 0.009576f
C228 B.n188 VSUBS 0.009576f
C229 B.n189 VSUBS 0.009576f
C230 B.n190 VSUBS 0.009576f
C231 B.n191 VSUBS 0.009576f
C232 B.n192 VSUBS 0.009576f
C233 B.n193 VSUBS 0.009576f
C234 B.n194 VSUBS 0.009576f
C235 B.n195 VSUBS 0.009576f
C236 B.n196 VSUBS 0.009576f
C237 B.n197 VSUBS 0.009576f
C238 B.n198 VSUBS 0.009576f
C239 B.n199 VSUBS 0.009576f
C240 B.n200 VSUBS 0.009576f
C241 B.n201 VSUBS 0.009576f
C242 B.n202 VSUBS 0.009576f
C243 B.n203 VSUBS 0.009576f
C244 B.n204 VSUBS 0.009576f
C245 B.n205 VSUBS 0.009576f
C246 B.n206 VSUBS 0.009576f
C247 B.n207 VSUBS 0.009576f
C248 B.n208 VSUBS 0.009576f
C249 B.n209 VSUBS 0.009576f
C250 B.n210 VSUBS 0.009576f
C251 B.n211 VSUBS 0.009576f
C252 B.n212 VSUBS 0.009576f
C253 B.n213 VSUBS 0.009576f
C254 B.n214 VSUBS 0.009576f
C255 B.n215 VSUBS 0.009576f
C256 B.n216 VSUBS 0.009576f
C257 B.n217 VSUBS 0.009576f
C258 B.n218 VSUBS 0.009576f
C259 B.n219 VSUBS 0.009576f
C260 B.n220 VSUBS 0.009576f
C261 B.n221 VSUBS 0.009576f
C262 B.n222 VSUBS 0.009576f
C263 B.n223 VSUBS 0.009576f
C264 B.n224 VSUBS 0.009576f
C265 B.n225 VSUBS 0.009576f
C266 B.n226 VSUBS 0.009576f
C267 B.n227 VSUBS 0.009576f
C268 B.n228 VSUBS 0.009576f
C269 B.n229 VSUBS 0.009576f
C270 B.n230 VSUBS 0.009576f
C271 B.n231 VSUBS 0.009576f
C272 B.n232 VSUBS 0.009576f
C273 B.n233 VSUBS 0.009576f
C274 B.n234 VSUBS 0.009576f
C275 B.n235 VSUBS 0.009576f
C276 B.n236 VSUBS 0.009576f
C277 B.n237 VSUBS 0.009576f
C278 B.n238 VSUBS 0.009576f
C279 B.n239 VSUBS 0.009576f
C280 B.n240 VSUBS 0.009576f
C281 B.n241 VSUBS 0.009576f
C282 B.n242 VSUBS 0.009576f
C283 B.n243 VSUBS 0.009576f
C284 B.n244 VSUBS 0.009576f
C285 B.n245 VSUBS 0.009576f
C286 B.n246 VSUBS 0.009576f
C287 B.n247 VSUBS 0.009576f
C288 B.n248 VSUBS 0.009576f
C289 B.n249 VSUBS 0.009576f
C290 B.n250 VSUBS 0.009576f
C291 B.n251 VSUBS 0.009576f
C292 B.n252 VSUBS 0.009576f
C293 B.n253 VSUBS 0.009576f
C294 B.n254 VSUBS 0.009576f
C295 B.n255 VSUBS 0.009576f
C296 B.n256 VSUBS 0.009576f
C297 B.n257 VSUBS 0.009576f
C298 B.n258 VSUBS 0.009576f
C299 B.n259 VSUBS 0.021526f
C300 B.n260 VSUBS 0.022129f
C301 B.n261 VSUBS 0.022129f
C302 B.n262 VSUBS 0.009576f
C303 B.n263 VSUBS 0.009576f
C304 B.n264 VSUBS 0.009576f
C305 B.n265 VSUBS 0.009576f
C306 B.n266 VSUBS 0.009576f
C307 B.n267 VSUBS 0.009576f
C308 B.n268 VSUBS 0.009576f
C309 B.n269 VSUBS 0.009576f
C310 B.n270 VSUBS 0.009576f
C311 B.n271 VSUBS 0.009576f
C312 B.n272 VSUBS 0.009576f
C313 B.n273 VSUBS 0.009576f
C314 B.n274 VSUBS 0.009576f
C315 B.n275 VSUBS 0.009576f
C316 B.n276 VSUBS 0.009576f
C317 B.n277 VSUBS 0.009576f
C318 B.n278 VSUBS 0.009576f
C319 B.n279 VSUBS 0.009576f
C320 B.n280 VSUBS 0.009576f
C321 B.n281 VSUBS 0.009576f
C322 B.n282 VSUBS 0.009576f
C323 B.n283 VSUBS 0.009576f
C324 B.n284 VSUBS 0.009576f
C325 B.n285 VSUBS 0.009576f
C326 B.n286 VSUBS 0.009576f
C327 B.n287 VSUBS 0.009576f
C328 B.n288 VSUBS 0.009576f
C329 B.n289 VSUBS 0.009576f
C330 B.n290 VSUBS 0.009576f
C331 B.n291 VSUBS 0.009576f
C332 B.n292 VSUBS 0.009576f
C333 B.n293 VSUBS 0.009576f
C334 B.n294 VSUBS 0.009576f
C335 B.n295 VSUBS 0.009576f
C336 B.n296 VSUBS 0.009576f
C337 B.n297 VSUBS 0.009576f
C338 B.n298 VSUBS 0.009576f
C339 B.n299 VSUBS 0.009576f
C340 B.n300 VSUBS 0.009576f
C341 B.n301 VSUBS 0.009576f
C342 B.n302 VSUBS 0.009576f
C343 B.n303 VSUBS 0.009576f
C344 B.n304 VSUBS 0.009576f
C345 B.n305 VSUBS 0.009013f
C346 B.n306 VSUBS 0.009576f
C347 B.n307 VSUBS 0.009576f
C348 B.n308 VSUBS 0.005351f
C349 B.n309 VSUBS 0.009576f
C350 B.n310 VSUBS 0.009576f
C351 B.n311 VSUBS 0.009576f
C352 B.n312 VSUBS 0.009576f
C353 B.n313 VSUBS 0.009576f
C354 B.n314 VSUBS 0.009576f
C355 B.n315 VSUBS 0.009576f
C356 B.n316 VSUBS 0.009576f
C357 B.n317 VSUBS 0.009576f
C358 B.n318 VSUBS 0.009576f
C359 B.n319 VSUBS 0.009576f
C360 B.n320 VSUBS 0.009576f
C361 B.n321 VSUBS 0.005351f
C362 B.n322 VSUBS 0.022186f
C363 B.n323 VSUBS 0.009013f
C364 B.n324 VSUBS 0.009576f
C365 B.n325 VSUBS 0.009576f
C366 B.n326 VSUBS 0.009576f
C367 B.n327 VSUBS 0.009576f
C368 B.n328 VSUBS 0.009576f
C369 B.n329 VSUBS 0.009576f
C370 B.n330 VSUBS 0.009576f
C371 B.n331 VSUBS 0.009576f
C372 B.n332 VSUBS 0.009576f
C373 B.n333 VSUBS 0.009576f
C374 B.n334 VSUBS 0.009576f
C375 B.n335 VSUBS 0.009576f
C376 B.n336 VSUBS 0.009576f
C377 B.n337 VSUBS 0.009576f
C378 B.n338 VSUBS 0.009576f
C379 B.n339 VSUBS 0.009576f
C380 B.n340 VSUBS 0.009576f
C381 B.n341 VSUBS 0.009576f
C382 B.n342 VSUBS 0.009576f
C383 B.n343 VSUBS 0.009576f
C384 B.n344 VSUBS 0.009576f
C385 B.n345 VSUBS 0.009576f
C386 B.n346 VSUBS 0.009576f
C387 B.n347 VSUBS 0.009576f
C388 B.n348 VSUBS 0.009576f
C389 B.n349 VSUBS 0.009576f
C390 B.n350 VSUBS 0.009576f
C391 B.n351 VSUBS 0.009576f
C392 B.n352 VSUBS 0.009576f
C393 B.n353 VSUBS 0.009576f
C394 B.n354 VSUBS 0.009576f
C395 B.n355 VSUBS 0.009576f
C396 B.n356 VSUBS 0.009576f
C397 B.n357 VSUBS 0.009576f
C398 B.n358 VSUBS 0.009576f
C399 B.n359 VSUBS 0.009576f
C400 B.n360 VSUBS 0.009576f
C401 B.n361 VSUBS 0.009576f
C402 B.n362 VSUBS 0.009576f
C403 B.n363 VSUBS 0.009576f
C404 B.n364 VSUBS 0.009576f
C405 B.n365 VSUBS 0.009576f
C406 B.n366 VSUBS 0.009576f
C407 B.n367 VSUBS 0.009576f
C408 B.n368 VSUBS 0.022129f
C409 B.n369 VSUBS 0.022129f
C410 B.n370 VSUBS 0.021526f
C411 B.n371 VSUBS 0.009576f
C412 B.n372 VSUBS 0.009576f
C413 B.n373 VSUBS 0.009576f
C414 B.n374 VSUBS 0.009576f
C415 B.n375 VSUBS 0.009576f
C416 B.n376 VSUBS 0.009576f
C417 B.n377 VSUBS 0.009576f
C418 B.n378 VSUBS 0.009576f
C419 B.n379 VSUBS 0.009576f
C420 B.n380 VSUBS 0.009576f
C421 B.n381 VSUBS 0.009576f
C422 B.n382 VSUBS 0.009576f
C423 B.n383 VSUBS 0.009576f
C424 B.n384 VSUBS 0.009576f
C425 B.n385 VSUBS 0.009576f
C426 B.n386 VSUBS 0.009576f
C427 B.n387 VSUBS 0.009576f
C428 B.n388 VSUBS 0.009576f
C429 B.n389 VSUBS 0.009576f
C430 B.n390 VSUBS 0.009576f
C431 B.n391 VSUBS 0.009576f
C432 B.n392 VSUBS 0.009576f
C433 B.n393 VSUBS 0.009576f
C434 B.n394 VSUBS 0.009576f
C435 B.n395 VSUBS 0.009576f
C436 B.n396 VSUBS 0.009576f
C437 B.n397 VSUBS 0.009576f
C438 B.n398 VSUBS 0.009576f
C439 B.n399 VSUBS 0.009576f
C440 B.n400 VSUBS 0.009576f
C441 B.n401 VSUBS 0.009576f
C442 B.n402 VSUBS 0.009576f
C443 B.n403 VSUBS 0.009576f
C444 B.n404 VSUBS 0.009576f
C445 B.n405 VSUBS 0.009576f
C446 B.n406 VSUBS 0.009576f
C447 B.n407 VSUBS 0.009576f
C448 B.n408 VSUBS 0.009576f
C449 B.n409 VSUBS 0.009576f
C450 B.n410 VSUBS 0.009576f
C451 B.n411 VSUBS 0.009576f
C452 B.n412 VSUBS 0.009576f
C453 B.n413 VSUBS 0.009576f
C454 B.n414 VSUBS 0.009576f
C455 B.n415 VSUBS 0.009576f
C456 B.n416 VSUBS 0.009576f
C457 B.n417 VSUBS 0.009576f
C458 B.n418 VSUBS 0.009576f
C459 B.n419 VSUBS 0.009576f
C460 B.n420 VSUBS 0.009576f
C461 B.n421 VSUBS 0.009576f
C462 B.n422 VSUBS 0.009576f
C463 B.n423 VSUBS 0.009576f
C464 B.n424 VSUBS 0.009576f
C465 B.n425 VSUBS 0.009576f
C466 B.n426 VSUBS 0.009576f
C467 B.n427 VSUBS 0.009576f
C468 B.n428 VSUBS 0.009576f
C469 B.n429 VSUBS 0.009576f
C470 B.n430 VSUBS 0.009576f
C471 B.n431 VSUBS 0.009576f
C472 B.n432 VSUBS 0.009576f
C473 B.n433 VSUBS 0.009576f
C474 B.n434 VSUBS 0.009576f
C475 B.n435 VSUBS 0.009576f
C476 B.n436 VSUBS 0.009576f
C477 B.n437 VSUBS 0.009576f
C478 B.n438 VSUBS 0.009576f
C479 B.n439 VSUBS 0.009576f
C480 B.n440 VSUBS 0.009576f
C481 B.n441 VSUBS 0.009576f
C482 B.n442 VSUBS 0.009576f
C483 B.n443 VSUBS 0.009576f
C484 B.n444 VSUBS 0.009576f
C485 B.n445 VSUBS 0.009576f
C486 B.n446 VSUBS 0.009576f
C487 B.n447 VSUBS 0.009576f
C488 B.n448 VSUBS 0.009576f
C489 B.n449 VSUBS 0.009576f
C490 B.n450 VSUBS 0.009576f
C491 B.n451 VSUBS 0.009576f
C492 B.n452 VSUBS 0.009576f
C493 B.n453 VSUBS 0.009576f
C494 B.n454 VSUBS 0.009576f
C495 B.n455 VSUBS 0.009576f
C496 B.n456 VSUBS 0.009576f
C497 B.n457 VSUBS 0.009576f
C498 B.n458 VSUBS 0.009576f
C499 B.n459 VSUBS 0.009576f
C500 B.n460 VSUBS 0.009576f
C501 B.n461 VSUBS 0.009576f
C502 B.n462 VSUBS 0.009576f
C503 B.n463 VSUBS 0.009576f
C504 B.n464 VSUBS 0.009576f
C505 B.n465 VSUBS 0.009576f
C506 B.n466 VSUBS 0.009576f
C507 B.n467 VSUBS 0.009576f
C508 B.n468 VSUBS 0.009576f
C509 B.n469 VSUBS 0.009576f
C510 B.n470 VSUBS 0.009576f
C511 B.n471 VSUBS 0.009576f
C512 B.n472 VSUBS 0.009576f
C513 B.n473 VSUBS 0.009576f
C514 B.n474 VSUBS 0.009576f
C515 B.n475 VSUBS 0.009576f
C516 B.n476 VSUBS 0.009576f
C517 B.n477 VSUBS 0.009576f
C518 B.n478 VSUBS 0.009576f
C519 B.n479 VSUBS 0.009576f
C520 B.n480 VSUBS 0.009576f
C521 B.n481 VSUBS 0.009576f
C522 B.n482 VSUBS 0.009576f
C523 B.n483 VSUBS 0.009576f
C524 B.n484 VSUBS 0.009576f
C525 B.n485 VSUBS 0.009576f
C526 B.n486 VSUBS 0.009576f
C527 B.n487 VSUBS 0.009576f
C528 B.n488 VSUBS 0.009576f
C529 B.n489 VSUBS 0.009576f
C530 B.n490 VSUBS 0.009576f
C531 B.n491 VSUBS 0.009576f
C532 B.n492 VSUBS 0.009576f
C533 B.n493 VSUBS 0.009576f
C534 B.n494 VSUBS 0.009576f
C535 B.n495 VSUBS 0.009576f
C536 B.n496 VSUBS 0.009576f
C537 B.n497 VSUBS 0.009576f
C538 B.n498 VSUBS 0.009576f
C539 B.n499 VSUBS 0.009576f
C540 B.n500 VSUBS 0.009576f
C541 B.n501 VSUBS 0.009576f
C542 B.n502 VSUBS 0.009576f
C543 B.n503 VSUBS 0.009576f
C544 B.n504 VSUBS 0.009576f
C545 B.n505 VSUBS 0.009576f
C546 B.n506 VSUBS 0.009576f
C547 B.n507 VSUBS 0.009576f
C548 B.n508 VSUBS 0.009576f
C549 B.n509 VSUBS 0.009576f
C550 B.n510 VSUBS 0.009576f
C551 B.n511 VSUBS 0.009576f
C552 B.n512 VSUBS 0.009576f
C553 B.n513 VSUBS 0.009576f
C554 B.n514 VSUBS 0.009576f
C555 B.n515 VSUBS 0.009576f
C556 B.n516 VSUBS 0.009576f
C557 B.n517 VSUBS 0.009576f
C558 B.n518 VSUBS 0.009576f
C559 B.n519 VSUBS 0.009576f
C560 B.n520 VSUBS 0.009576f
C561 B.n521 VSUBS 0.009576f
C562 B.n522 VSUBS 0.009576f
C563 B.n523 VSUBS 0.021526f
C564 B.n524 VSUBS 0.022129f
C565 B.n525 VSUBS 0.020951f
C566 B.n526 VSUBS 0.009576f
C567 B.n527 VSUBS 0.009576f
C568 B.n528 VSUBS 0.009576f
C569 B.n529 VSUBS 0.009576f
C570 B.n530 VSUBS 0.009576f
C571 B.n531 VSUBS 0.009576f
C572 B.n532 VSUBS 0.009576f
C573 B.n533 VSUBS 0.009576f
C574 B.n534 VSUBS 0.009576f
C575 B.n535 VSUBS 0.009576f
C576 B.n536 VSUBS 0.009576f
C577 B.n537 VSUBS 0.009576f
C578 B.n538 VSUBS 0.009576f
C579 B.n539 VSUBS 0.009576f
C580 B.n540 VSUBS 0.009576f
C581 B.n541 VSUBS 0.009576f
C582 B.n542 VSUBS 0.009576f
C583 B.n543 VSUBS 0.009576f
C584 B.n544 VSUBS 0.009576f
C585 B.n545 VSUBS 0.009576f
C586 B.n546 VSUBS 0.009576f
C587 B.n547 VSUBS 0.009576f
C588 B.n548 VSUBS 0.009576f
C589 B.n549 VSUBS 0.009576f
C590 B.n550 VSUBS 0.009576f
C591 B.n551 VSUBS 0.009576f
C592 B.n552 VSUBS 0.009576f
C593 B.n553 VSUBS 0.009576f
C594 B.n554 VSUBS 0.009576f
C595 B.n555 VSUBS 0.009576f
C596 B.n556 VSUBS 0.009576f
C597 B.n557 VSUBS 0.009576f
C598 B.n558 VSUBS 0.009576f
C599 B.n559 VSUBS 0.009576f
C600 B.n560 VSUBS 0.009576f
C601 B.n561 VSUBS 0.009576f
C602 B.n562 VSUBS 0.009576f
C603 B.n563 VSUBS 0.009576f
C604 B.n564 VSUBS 0.009576f
C605 B.n565 VSUBS 0.009576f
C606 B.n566 VSUBS 0.009576f
C607 B.n567 VSUBS 0.009576f
C608 B.n568 VSUBS 0.009576f
C609 B.n569 VSUBS 0.009013f
C610 B.n570 VSUBS 0.009576f
C611 B.n571 VSUBS 0.009576f
C612 B.n572 VSUBS 0.005351f
C613 B.n573 VSUBS 0.009576f
C614 B.n574 VSUBS 0.009576f
C615 B.n575 VSUBS 0.009576f
C616 B.n576 VSUBS 0.009576f
C617 B.n577 VSUBS 0.009576f
C618 B.n578 VSUBS 0.009576f
C619 B.n579 VSUBS 0.009576f
C620 B.n580 VSUBS 0.009576f
C621 B.n581 VSUBS 0.009576f
C622 B.n582 VSUBS 0.009576f
C623 B.n583 VSUBS 0.009576f
C624 B.n584 VSUBS 0.009576f
C625 B.n585 VSUBS 0.005351f
C626 B.n586 VSUBS 0.022186f
C627 B.n587 VSUBS 0.009013f
C628 B.n588 VSUBS 0.009576f
C629 B.n589 VSUBS 0.009576f
C630 B.n590 VSUBS 0.009576f
C631 B.n591 VSUBS 0.009576f
C632 B.n592 VSUBS 0.009576f
C633 B.n593 VSUBS 0.009576f
C634 B.n594 VSUBS 0.009576f
C635 B.n595 VSUBS 0.009576f
C636 B.n596 VSUBS 0.009576f
C637 B.n597 VSUBS 0.009576f
C638 B.n598 VSUBS 0.009576f
C639 B.n599 VSUBS 0.009576f
C640 B.n600 VSUBS 0.009576f
C641 B.n601 VSUBS 0.009576f
C642 B.n602 VSUBS 0.009576f
C643 B.n603 VSUBS 0.009576f
C644 B.n604 VSUBS 0.009576f
C645 B.n605 VSUBS 0.009576f
C646 B.n606 VSUBS 0.009576f
C647 B.n607 VSUBS 0.009576f
C648 B.n608 VSUBS 0.009576f
C649 B.n609 VSUBS 0.009576f
C650 B.n610 VSUBS 0.009576f
C651 B.n611 VSUBS 0.009576f
C652 B.n612 VSUBS 0.009576f
C653 B.n613 VSUBS 0.009576f
C654 B.n614 VSUBS 0.009576f
C655 B.n615 VSUBS 0.009576f
C656 B.n616 VSUBS 0.009576f
C657 B.n617 VSUBS 0.009576f
C658 B.n618 VSUBS 0.009576f
C659 B.n619 VSUBS 0.009576f
C660 B.n620 VSUBS 0.009576f
C661 B.n621 VSUBS 0.009576f
C662 B.n622 VSUBS 0.009576f
C663 B.n623 VSUBS 0.009576f
C664 B.n624 VSUBS 0.009576f
C665 B.n625 VSUBS 0.009576f
C666 B.n626 VSUBS 0.009576f
C667 B.n627 VSUBS 0.009576f
C668 B.n628 VSUBS 0.009576f
C669 B.n629 VSUBS 0.009576f
C670 B.n630 VSUBS 0.009576f
C671 B.n631 VSUBS 0.009576f
C672 B.n632 VSUBS 0.022129f
C673 B.n633 VSUBS 0.022129f
C674 B.n634 VSUBS 0.021526f
C675 B.n635 VSUBS 0.009576f
C676 B.n636 VSUBS 0.009576f
C677 B.n637 VSUBS 0.009576f
C678 B.n638 VSUBS 0.009576f
C679 B.n639 VSUBS 0.009576f
C680 B.n640 VSUBS 0.009576f
C681 B.n641 VSUBS 0.009576f
C682 B.n642 VSUBS 0.009576f
C683 B.n643 VSUBS 0.009576f
C684 B.n644 VSUBS 0.009576f
C685 B.n645 VSUBS 0.009576f
C686 B.n646 VSUBS 0.009576f
C687 B.n647 VSUBS 0.009576f
C688 B.n648 VSUBS 0.009576f
C689 B.n649 VSUBS 0.009576f
C690 B.n650 VSUBS 0.009576f
C691 B.n651 VSUBS 0.009576f
C692 B.n652 VSUBS 0.009576f
C693 B.n653 VSUBS 0.009576f
C694 B.n654 VSUBS 0.009576f
C695 B.n655 VSUBS 0.009576f
C696 B.n656 VSUBS 0.009576f
C697 B.n657 VSUBS 0.009576f
C698 B.n658 VSUBS 0.009576f
C699 B.n659 VSUBS 0.009576f
C700 B.n660 VSUBS 0.009576f
C701 B.n661 VSUBS 0.009576f
C702 B.n662 VSUBS 0.009576f
C703 B.n663 VSUBS 0.009576f
C704 B.n664 VSUBS 0.009576f
C705 B.n665 VSUBS 0.009576f
C706 B.n666 VSUBS 0.009576f
C707 B.n667 VSUBS 0.009576f
C708 B.n668 VSUBS 0.009576f
C709 B.n669 VSUBS 0.009576f
C710 B.n670 VSUBS 0.009576f
C711 B.n671 VSUBS 0.009576f
C712 B.n672 VSUBS 0.009576f
C713 B.n673 VSUBS 0.009576f
C714 B.n674 VSUBS 0.009576f
C715 B.n675 VSUBS 0.009576f
C716 B.n676 VSUBS 0.009576f
C717 B.n677 VSUBS 0.009576f
C718 B.n678 VSUBS 0.009576f
C719 B.n679 VSUBS 0.009576f
C720 B.n680 VSUBS 0.009576f
C721 B.n681 VSUBS 0.009576f
C722 B.n682 VSUBS 0.009576f
C723 B.n683 VSUBS 0.009576f
C724 B.n684 VSUBS 0.009576f
C725 B.n685 VSUBS 0.009576f
C726 B.n686 VSUBS 0.009576f
C727 B.n687 VSUBS 0.009576f
C728 B.n688 VSUBS 0.009576f
C729 B.n689 VSUBS 0.009576f
C730 B.n690 VSUBS 0.009576f
C731 B.n691 VSUBS 0.009576f
C732 B.n692 VSUBS 0.009576f
C733 B.n693 VSUBS 0.009576f
C734 B.n694 VSUBS 0.009576f
C735 B.n695 VSUBS 0.009576f
C736 B.n696 VSUBS 0.009576f
C737 B.n697 VSUBS 0.009576f
C738 B.n698 VSUBS 0.009576f
C739 B.n699 VSUBS 0.009576f
C740 B.n700 VSUBS 0.009576f
C741 B.n701 VSUBS 0.009576f
C742 B.n702 VSUBS 0.009576f
C743 B.n703 VSUBS 0.009576f
C744 B.n704 VSUBS 0.009576f
C745 B.n705 VSUBS 0.009576f
C746 B.n706 VSUBS 0.009576f
C747 B.n707 VSUBS 0.009576f
C748 B.n708 VSUBS 0.009576f
C749 B.n709 VSUBS 0.009576f
C750 B.n710 VSUBS 0.009576f
C751 B.n711 VSUBS 0.021683f
C752 VDD1.t7 VSUBS 1.85291f
C753 VDD1.t1 VSUBS 0.192118f
C754 VDD1.t3 VSUBS 0.192118f
C755 VDD1.n0 VSUBS 1.38738f
C756 VDD1.n1 VSUBS 1.53547f
C757 VDD1.t4 VSUBS 1.85291f
C758 VDD1.t2 VSUBS 0.192118f
C759 VDD1.t6 VSUBS 0.192118f
C760 VDD1.n2 VSUBS 1.38738f
C761 VDD1.n3 VSUBS 1.52643f
C762 VDD1.t0 VSUBS 0.192118f
C763 VDD1.t8 VSUBS 0.192118f
C764 VDD1.n4 VSUBS 1.40304f
C765 VDD1.n5 VSUBS 3.17758f
C766 VDD1.t9 VSUBS 0.192118f
C767 VDD1.t5 VSUBS 0.192118f
C768 VDD1.n6 VSUBS 1.38738f
C769 VDD1.n7 VSUBS 3.36007f
C770 VP.n0 VSUBS 0.047262f
C771 VP.t1 VSUBS 1.71264f
C772 VP.n1 VSUBS 0.037599f
C773 VP.n2 VSUBS 0.035848f
C774 VP.t9 VSUBS 1.71264f
C775 VP.n3 VSUBS 0.056328f
C776 VP.n4 VSUBS 0.035848f
C777 VP.t3 VSUBS 1.71264f
C778 VP.n5 VSUBS 0.066812f
C779 VP.n6 VSUBS 0.035848f
C780 VP.t7 VSUBS 1.71264f
C781 VP.n7 VSUBS 0.627195f
C782 VP.n8 VSUBS 0.035848f
C783 VP.n9 VSUBS 0.063606f
C784 VP.n10 VSUBS 0.047262f
C785 VP.t4 VSUBS 1.71264f
C786 VP.n11 VSUBS 0.037599f
C787 VP.n12 VSUBS 0.035848f
C788 VP.t0 VSUBS 1.71264f
C789 VP.n13 VSUBS 0.056328f
C790 VP.n14 VSUBS 0.035848f
C791 VP.t6 VSUBS 1.71264f
C792 VP.n15 VSUBS 0.066812f
C793 VP.n16 VSUBS 0.035848f
C794 VP.t8 VSUBS 1.71264f
C795 VP.n17 VSUBS 0.727929f
C796 VP.t2 VSUBS 1.92039f
C797 VP.n18 VSUBS 0.705794f
C798 VP.n19 VSUBS 0.301507f
C799 VP.n20 VSUBS 0.061534f
C800 VP.n21 VSUBS 0.056328f
C801 VP.n22 VSUBS 0.048336f
C802 VP.n23 VSUBS 0.035848f
C803 VP.n24 VSUBS 0.035848f
C804 VP.n25 VSUBS 0.035848f
C805 VP.n26 VSUBS 0.661022f
C806 VP.n27 VSUBS 0.066812f
C807 VP.n28 VSUBS 0.048336f
C808 VP.n29 VSUBS 0.035848f
C809 VP.n30 VSUBS 0.035848f
C810 VP.n31 VSUBS 0.035848f
C811 VP.n32 VSUBS 0.061534f
C812 VP.n33 VSUBS 0.627195f
C813 VP.n34 VSUBS 0.039104f
C814 VP.n35 VSUBS 0.070271f
C815 VP.n36 VSUBS 0.035848f
C816 VP.n37 VSUBS 0.035848f
C817 VP.n38 VSUBS 0.035848f
C818 VP.n39 VSUBS 0.063606f
C819 VP.n40 VSUBS 0.056257f
C820 VP.n41 VSUBS 0.735251f
C821 VP.n42 VSUBS 1.84653f
C822 VP.n43 VSUBS 1.87356f
C823 VP.t5 VSUBS 1.71264f
C824 VP.n44 VSUBS 0.735251f
C825 VP.n45 VSUBS 0.056257f
C826 VP.n46 VSUBS 0.047262f
C827 VP.n47 VSUBS 0.035848f
C828 VP.n48 VSUBS 0.035848f
C829 VP.n49 VSUBS 0.037599f
C830 VP.n50 VSUBS 0.070271f
C831 VP.n51 VSUBS 0.039104f
C832 VP.n52 VSUBS 0.035848f
C833 VP.n53 VSUBS 0.035848f
C834 VP.n54 VSUBS 0.061534f
C835 VP.n55 VSUBS 0.056328f
C836 VP.n56 VSUBS 0.048336f
C837 VP.n57 VSUBS 0.035848f
C838 VP.n58 VSUBS 0.035848f
C839 VP.n59 VSUBS 0.035848f
C840 VP.n60 VSUBS 0.661022f
C841 VP.n61 VSUBS 0.066812f
C842 VP.n62 VSUBS 0.048336f
C843 VP.n63 VSUBS 0.035848f
C844 VP.n64 VSUBS 0.035848f
C845 VP.n65 VSUBS 0.035848f
C846 VP.n66 VSUBS 0.061534f
C847 VP.n67 VSUBS 0.627195f
C848 VP.n68 VSUBS 0.039104f
C849 VP.n69 VSUBS 0.070271f
C850 VP.n70 VSUBS 0.035848f
C851 VP.n71 VSUBS 0.035848f
C852 VP.n72 VSUBS 0.035848f
C853 VP.n73 VSUBS 0.063606f
C854 VP.n74 VSUBS 0.056257f
C855 VP.n75 VSUBS 0.735251f
C856 VP.n76 VSUBS 0.047253f
C857 VTAIL.t14 VSUBS 0.201765f
C858 VTAIL.t19 VSUBS 0.201765f
C859 VTAIL.n0 VSUBS 1.31894f
C860 VTAIL.n1 VSUBS 0.940405f
C861 VTAIL.t1 VSUBS 1.77569f
C862 VTAIL.n2 VSUBS 1.07882f
C863 VTAIL.t5 VSUBS 0.201765f
C864 VTAIL.t9 VSUBS 0.201765f
C865 VTAIL.n3 VSUBS 1.31894f
C866 VTAIL.n4 VSUBS 1.04086f
C867 VTAIL.t4 VSUBS 0.201765f
C868 VTAIL.t7 VSUBS 0.201765f
C869 VTAIL.n5 VSUBS 1.31894f
C870 VTAIL.n6 VSUBS 2.36077f
C871 VTAIL.t11 VSUBS 0.201765f
C872 VTAIL.t15 VSUBS 0.201765f
C873 VTAIL.n7 VSUBS 1.31894f
C874 VTAIL.n8 VSUBS 2.36076f
C875 VTAIL.t10 VSUBS 0.201765f
C876 VTAIL.t18 VSUBS 0.201765f
C877 VTAIL.n9 VSUBS 1.31894f
C878 VTAIL.n10 VSUBS 1.04085f
C879 VTAIL.t16 VSUBS 1.7757f
C880 VTAIL.n11 VSUBS 1.07882f
C881 VTAIL.t2 VSUBS 0.201765f
C882 VTAIL.t6 VSUBS 0.201765f
C883 VTAIL.n12 VSUBS 1.31894f
C884 VTAIL.n13 VSUBS 0.9853f
C885 VTAIL.t8 VSUBS 0.201765f
C886 VTAIL.t3 VSUBS 0.201765f
C887 VTAIL.n14 VSUBS 1.31894f
C888 VTAIL.n15 VSUBS 1.04085f
C889 VTAIL.t0 VSUBS 1.7757f
C890 VTAIL.n16 VSUBS 2.25212f
C891 VTAIL.t13 VSUBS 1.77569f
C892 VTAIL.n17 VSUBS 2.25213f
C893 VTAIL.t12 VSUBS 0.201765f
C894 VTAIL.t17 VSUBS 0.201765f
C895 VTAIL.n18 VSUBS 1.31894f
C896 VTAIL.n19 VSUBS 0.8836f
C897 VDD2.t9 VSUBS 1.85343f
C898 VDD2.t3 VSUBS 0.192172f
C899 VDD2.t5 VSUBS 0.192172f
C900 VDD2.n0 VSUBS 1.38777f
C901 VDD2.n1 VSUBS 1.52686f
C902 VDD2.t8 VSUBS 0.192172f
C903 VDD2.t4 VSUBS 0.192172f
C904 VDD2.n2 VSUBS 1.40343f
C905 VDD2.n3 VSUBS 3.05341f
C906 VDD2.t0 VSUBS 1.83437f
C907 VDD2.n4 VSUBS 3.31876f
C908 VDD2.t6 VSUBS 0.192172f
C909 VDD2.t1 VSUBS 0.192172f
C910 VDD2.n5 VSUBS 1.38777f
C911 VDD2.n6 VSUBS 0.759715f
C912 VDD2.t2 VSUBS 0.192172f
C913 VDD2.t7 VSUBS 0.192172f
C914 VDD2.n7 VSUBS 1.4034f
C915 VN.n0 VSUBS 0.045825f
C916 VN.t6 VSUBS 1.66056f
C917 VN.n1 VSUBS 0.036455f
C918 VN.n2 VSUBS 0.034758f
C919 VN.t2 VSUBS 1.66056f
C920 VN.n3 VSUBS 0.054615f
C921 VN.n4 VSUBS 0.034758f
C922 VN.t7 VSUBS 1.66056f
C923 VN.n5 VSUBS 0.06478f
C924 VN.n6 VSUBS 0.034758f
C925 VN.t0 VSUBS 1.66056f
C926 VN.n7 VSUBS 0.705791f
C927 VN.t5 VSUBS 1.86199f
C928 VN.n8 VSUBS 0.68433f
C929 VN.n9 VSUBS 0.292337f
C930 VN.n10 VSUBS 0.059663f
C931 VN.n11 VSUBS 0.054615f
C932 VN.n12 VSUBS 0.046866f
C933 VN.n13 VSUBS 0.034758f
C934 VN.n14 VSUBS 0.034758f
C935 VN.n15 VSUBS 0.034758f
C936 VN.n16 VSUBS 0.640919f
C937 VN.n17 VSUBS 0.06478f
C938 VN.n18 VSUBS 0.046866f
C939 VN.n19 VSUBS 0.034758f
C940 VN.n20 VSUBS 0.034758f
C941 VN.n21 VSUBS 0.034758f
C942 VN.n22 VSUBS 0.059663f
C943 VN.n23 VSUBS 0.608121f
C944 VN.n24 VSUBS 0.037915f
C945 VN.n25 VSUBS 0.068133f
C946 VN.n26 VSUBS 0.034758f
C947 VN.n27 VSUBS 0.034758f
C948 VN.n28 VSUBS 0.034758f
C949 VN.n29 VSUBS 0.061672f
C950 VN.n30 VSUBS 0.054546f
C951 VN.n31 VSUBS 0.712891f
C952 VN.n32 VSUBS 0.045816f
C953 VN.n33 VSUBS 0.045825f
C954 VN.t8 VSUBS 1.66056f
C955 VN.n34 VSUBS 0.036455f
C956 VN.n35 VSUBS 0.034758f
C957 VN.t4 VSUBS 1.66056f
C958 VN.n36 VSUBS 0.054615f
C959 VN.n37 VSUBS 0.034758f
C960 VN.t9 VSUBS 1.66056f
C961 VN.n38 VSUBS 0.06478f
C962 VN.n39 VSUBS 0.034758f
C963 VN.t1 VSUBS 1.66056f
C964 VN.n40 VSUBS 0.705791f
C965 VN.t3 VSUBS 1.86199f
C966 VN.n41 VSUBS 0.68433f
C967 VN.n42 VSUBS 0.292337f
C968 VN.n43 VSUBS 0.059663f
C969 VN.n44 VSUBS 0.054615f
C970 VN.n45 VSUBS 0.046866f
C971 VN.n46 VSUBS 0.034758f
C972 VN.n47 VSUBS 0.034758f
C973 VN.n48 VSUBS 0.034758f
C974 VN.n49 VSUBS 0.640919f
C975 VN.n50 VSUBS 0.06478f
C976 VN.n51 VSUBS 0.046866f
C977 VN.n52 VSUBS 0.034758f
C978 VN.n53 VSUBS 0.034758f
C979 VN.n54 VSUBS 0.034758f
C980 VN.n55 VSUBS 0.059663f
C981 VN.n56 VSUBS 0.608121f
C982 VN.n57 VSUBS 0.037915f
C983 VN.n58 VSUBS 0.068133f
C984 VN.n59 VSUBS 0.034758f
C985 VN.n60 VSUBS 0.034758f
C986 VN.n61 VSUBS 0.034758f
C987 VN.n62 VSUBS 0.061672f
C988 VN.n63 VSUBS 0.054546f
C989 VN.n64 VSUBS 0.712891f
C990 VN.n65 VSUBS 1.8092f
.ends

