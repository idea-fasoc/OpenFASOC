* NGSPICE file created from diff_pair_sample_0469.ext - technology: sky130A

.subckt diff_pair_sample_0469 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X1 VDD1.t8 VP.t1 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=2.6247 ps=14.24 w=6.73 l=3.37
X2 VDD1.t7 VP.t2 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=2.6247 ps=14.24 w=6.73 l=3.37
X3 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=2.6247 pd=14.24 as=0 ps=0 w=6.73 l=3.37
X4 VTAIL.t17 VP.t3 VDD1.t6 B.t8 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X5 VDD2.t9 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.6247 pd=14.24 as=1.11045 ps=7.06 w=6.73 l=3.37
X6 VDD2.t8 VN.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.6247 pd=14.24 as=1.11045 ps=7.06 w=6.73 l=3.37
X7 VTAIL.t12 VP.t4 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X8 VDD1.t4 VP.t5 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X9 VTAIL.t4 VN.t2 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X10 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=2.6247 pd=14.24 as=0 ps=0 w=6.73 l=3.37
X11 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=2.6247 pd=14.24 as=0 ps=0 w=6.73 l=3.37
X12 VTAIL.t19 VP.t6 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X13 VTAIL.t3 VN.t3 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X14 VTAIL.t8 VN.t4 VDD2.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X15 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.6247 pd=14.24 as=0 ps=0 w=6.73 l=3.37
X16 VDD2.t4 VN.t5 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=2.6247 ps=14.24 w=6.73 l=3.37
X17 VTAIL.t7 VN.t6 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X18 VTAIL.t11 VP.t7 VDD1.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X19 VDD2.t2 VN.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X20 VDD1.t1 VP.t8 VTAIL.t18 B.t6 sky130_fd_pr__nfet_01v8 ad=2.6247 pd=14.24 as=1.11045 ps=7.06 w=6.73 l=3.37
X21 VDD2.t1 VN.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=2.6247 ps=14.24 w=6.73 l=3.37
X22 VDD2.t0 VN.t9 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.11045 pd=7.06 as=1.11045 ps=7.06 w=6.73 l=3.37
X23 VDD1.t0 VP.t9 VTAIL.t16 B.t2 sky130_fd_pr__nfet_01v8 ad=2.6247 pd=14.24 as=1.11045 ps=7.06 w=6.73 l=3.37
R0 VP.n32 VP.n31 161.3
R1 VP.n33 VP.n28 161.3
R2 VP.n35 VP.n34 161.3
R3 VP.n36 VP.n27 161.3
R4 VP.n38 VP.n37 161.3
R5 VP.n39 VP.n26 161.3
R6 VP.n41 VP.n40 161.3
R7 VP.n43 VP.n42 161.3
R8 VP.n44 VP.n24 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n47 VP.n23 161.3
R11 VP.n49 VP.n48 161.3
R12 VP.n50 VP.n22 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n21 161.3
R15 VP.n56 VP.n55 161.3
R16 VP.n57 VP.n20 161.3
R17 VP.n59 VP.n58 161.3
R18 VP.n60 VP.n19 161.3
R19 VP.n62 VP.n61 161.3
R20 VP.n63 VP.n18 161.3
R21 VP.n65 VP.n64 161.3
R22 VP.n115 VP.n114 161.3
R23 VP.n113 VP.n1 161.3
R24 VP.n112 VP.n111 161.3
R25 VP.n110 VP.n2 161.3
R26 VP.n109 VP.n108 161.3
R27 VP.n107 VP.n3 161.3
R28 VP.n106 VP.n105 161.3
R29 VP.n104 VP.n4 161.3
R30 VP.n103 VP.n102 161.3
R31 VP.n100 VP.n5 161.3
R32 VP.n99 VP.n98 161.3
R33 VP.n97 VP.n6 161.3
R34 VP.n96 VP.n95 161.3
R35 VP.n94 VP.n7 161.3
R36 VP.n93 VP.n92 161.3
R37 VP.n91 VP.n90 161.3
R38 VP.n89 VP.n9 161.3
R39 VP.n88 VP.n87 161.3
R40 VP.n86 VP.n10 161.3
R41 VP.n85 VP.n84 161.3
R42 VP.n83 VP.n11 161.3
R43 VP.n82 VP.n81 161.3
R44 VP.n80 VP.n79 161.3
R45 VP.n78 VP.n13 161.3
R46 VP.n77 VP.n76 161.3
R47 VP.n75 VP.n14 161.3
R48 VP.n74 VP.n73 161.3
R49 VP.n72 VP.n15 161.3
R50 VP.n71 VP.n70 161.3
R51 VP.n69 VP.n16 161.3
R52 VP.n68 VP.n67 82.7273
R53 VP.n116 VP.n0 82.7273
R54 VP.n66 VP.n17 82.7273
R55 VP.n30 VP.t8 81.0578
R56 VP.n73 VP.n14 56.5193
R57 VP.n108 VP.n2 56.5193
R58 VP.n58 VP.n19 56.5193
R59 VP.n68 VP.n66 53.3251
R60 VP.n30 VP.n29 52.4975
R61 VP.n84 VP.n10 50.2061
R62 VP.n99 VP.n6 50.2061
R63 VP.n49 VP.n23 50.2061
R64 VP.n34 VP.n27 50.2061
R65 VP.n67 VP.t9 48.129
R66 VP.n12 VP.t4 48.129
R67 VP.n8 VP.t0 48.129
R68 VP.n101 VP.t6 48.129
R69 VP.n0 VP.t1 48.129
R70 VP.n17 VP.t2 48.129
R71 VP.n51 VP.t3 48.129
R72 VP.n25 VP.t5 48.129
R73 VP.n29 VP.t7 48.129
R74 VP.n88 VP.n10 30.7807
R75 VP.n95 VP.n6 30.7807
R76 VP.n45 VP.n23 30.7807
R77 VP.n38 VP.n27 30.7807
R78 VP.n71 VP.n16 24.4675
R79 VP.n72 VP.n71 24.4675
R80 VP.n73 VP.n72 24.4675
R81 VP.n77 VP.n14 24.4675
R82 VP.n78 VP.n77 24.4675
R83 VP.n79 VP.n78 24.4675
R84 VP.n83 VP.n82 24.4675
R85 VP.n84 VP.n83 24.4675
R86 VP.n89 VP.n88 24.4675
R87 VP.n90 VP.n89 24.4675
R88 VP.n94 VP.n93 24.4675
R89 VP.n95 VP.n94 24.4675
R90 VP.n100 VP.n99 24.4675
R91 VP.n102 VP.n100 24.4675
R92 VP.n106 VP.n4 24.4675
R93 VP.n107 VP.n106 24.4675
R94 VP.n108 VP.n107 24.4675
R95 VP.n112 VP.n2 24.4675
R96 VP.n113 VP.n112 24.4675
R97 VP.n114 VP.n113 24.4675
R98 VP.n62 VP.n19 24.4675
R99 VP.n63 VP.n62 24.4675
R100 VP.n64 VP.n63 24.4675
R101 VP.n50 VP.n49 24.4675
R102 VP.n52 VP.n50 24.4675
R103 VP.n56 VP.n21 24.4675
R104 VP.n57 VP.n56 24.4675
R105 VP.n58 VP.n57 24.4675
R106 VP.n39 VP.n38 24.4675
R107 VP.n40 VP.n39 24.4675
R108 VP.n44 VP.n43 24.4675
R109 VP.n45 VP.n44 24.4675
R110 VP.n33 VP.n32 24.4675
R111 VP.n34 VP.n33 24.4675
R112 VP.n82 VP.n12 22.0208
R113 VP.n102 VP.n101 22.0208
R114 VP.n52 VP.n51 22.0208
R115 VP.n32 VP.n29 22.0208
R116 VP.n90 VP.n8 12.234
R117 VP.n93 VP.n8 12.234
R118 VP.n40 VP.n25 12.234
R119 VP.n43 VP.n25 12.234
R120 VP.n67 VP.n16 7.3406
R121 VP.n114 VP.n0 7.3406
R122 VP.n64 VP.n17 7.3406
R123 VP.n31 VP.n30 3.24374
R124 VP.n79 VP.n12 2.4472
R125 VP.n101 VP.n4 2.4472
R126 VP.n51 VP.n21 2.4472
R127 VP.n66 VP.n65 0.354971
R128 VP.n69 VP.n68 0.354971
R129 VP.n116 VP.n115 0.354971
R130 VP VP.n116 0.26696
R131 VP.n31 VP.n28 0.189894
R132 VP.n35 VP.n28 0.189894
R133 VP.n36 VP.n35 0.189894
R134 VP.n37 VP.n36 0.189894
R135 VP.n37 VP.n26 0.189894
R136 VP.n41 VP.n26 0.189894
R137 VP.n42 VP.n41 0.189894
R138 VP.n42 VP.n24 0.189894
R139 VP.n46 VP.n24 0.189894
R140 VP.n47 VP.n46 0.189894
R141 VP.n48 VP.n47 0.189894
R142 VP.n48 VP.n22 0.189894
R143 VP.n53 VP.n22 0.189894
R144 VP.n54 VP.n53 0.189894
R145 VP.n55 VP.n54 0.189894
R146 VP.n55 VP.n20 0.189894
R147 VP.n59 VP.n20 0.189894
R148 VP.n60 VP.n59 0.189894
R149 VP.n61 VP.n60 0.189894
R150 VP.n61 VP.n18 0.189894
R151 VP.n65 VP.n18 0.189894
R152 VP.n70 VP.n69 0.189894
R153 VP.n70 VP.n15 0.189894
R154 VP.n74 VP.n15 0.189894
R155 VP.n75 VP.n74 0.189894
R156 VP.n76 VP.n75 0.189894
R157 VP.n76 VP.n13 0.189894
R158 VP.n80 VP.n13 0.189894
R159 VP.n81 VP.n80 0.189894
R160 VP.n81 VP.n11 0.189894
R161 VP.n85 VP.n11 0.189894
R162 VP.n86 VP.n85 0.189894
R163 VP.n87 VP.n86 0.189894
R164 VP.n87 VP.n9 0.189894
R165 VP.n91 VP.n9 0.189894
R166 VP.n92 VP.n91 0.189894
R167 VP.n92 VP.n7 0.189894
R168 VP.n96 VP.n7 0.189894
R169 VP.n97 VP.n96 0.189894
R170 VP.n98 VP.n97 0.189894
R171 VP.n98 VP.n5 0.189894
R172 VP.n103 VP.n5 0.189894
R173 VP.n104 VP.n103 0.189894
R174 VP.n105 VP.n104 0.189894
R175 VP.n105 VP.n3 0.189894
R176 VP.n109 VP.n3 0.189894
R177 VP.n110 VP.n109 0.189894
R178 VP.n111 VP.n110 0.189894
R179 VP.n111 VP.n1 0.189894
R180 VP.n115 VP.n1 0.189894
R181 VTAIL.n152 VTAIL.n122 289.615
R182 VTAIL.n32 VTAIL.n2 289.615
R183 VTAIL.n116 VTAIL.n86 289.615
R184 VTAIL.n76 VTAIL.n46 289.615
R185 VTAIL.n135 VTAIL.n134 185
R186 VTAIL.n137 VTAIL.n136 185
R187 VTAIL.n130 VTAIL.n129 185
R188 VTAIL.n143 VTAIL.n142 185
R189 VTAIL.n145 VTAIL.n144 185
R190 VTAIL.n126 VTAIL.n125 185
R191 VTAIL.n151 VTAIL.n150 185
R192 VTAIL.n153 VTAIL.n152 185
R193 VTAIL.n15 VTAIL.n14 185
R194 VTAIL.n17 VTAIL.n16 185
R195 VTAIL.n10 VTAIL.n9 185
R196 VTAIL.n23 VTAIL.n22 185
R197 VTAIL.n25 VTAIL.n24 185
R198 VTAIL.n6 VTAIL.n5 185
R199 VTAIL.n31 VTAIL.n30 185
R200 VTAIL.n33 VTAIL.n32 185
R201 VTAIL.n117 VTAIL.n116 185
R202 VTAIL.n115 VTAIL.n114 185
R203 VTAIL.n90 VTAIL.n89 185
R204 VTAIL.n109 VTAIL.n108 185
R205 VTAIL.n107 VTAIL.n106 185
R206 VTAIL.n94 VTAIL.n93 185
R207 VTAIL.n101 VTAIL.n100 185
R208 VTAIL.n99 VTAIL.n98 185
R209 VTAIL.n77 VTAIL.n76 185
R210 VTAIL.n75 VTAIL.n74 185
R211 VTAIL.n50 VTAIL.n49 185
R212 VTAIL.n69 VTAIL.n68 185
R213 VTAIL.n67 VTAIL.n66 185
R214 VTAIL.n54 VTAIL.n53 185
R215 VTAIL.n61 VTAIL.n60 185
R216 VTAIL.n59 VTAIL.n58 185
R217 VTAIL.n133 VTAIL.t5 147.659
R218 VTAIL.n13 VTAIL.t15 147.659
R219 VTAIL.n97 VTAIL.t10 147.659
R220 VTAIL.n57 VTAIL.t9 147.659
R221 VTAIL.n136 VTAIL.n135 104.615
R222 VTAIL.n136 VTAIL.n129 104.615
R223 VTAIL.n143 VTAIL.n129 104.615
R224 VTAIL.n144 VTAIL.n143 104.615
R225 VTAIL.n144 VTAIL.n125 104.615
R226 VTAIL.n151 VTAIL.n125 104.615
R227 VTAIL.n152 VTAIL.n151 104.615
R228 VTAIL.n16 VTAIL.n15 104.615
R229 VTAIL.n16 VTAIL.n9 104.615
R230 VTAIL.n23 VTAIL.n9 104.615
R231 VTAIL.n24 VTAIL.n23 104.615
R232 VTAIL.n24 VTAIL.n5 104.615
R233 VTAIL.n31 VTAIL.n5 104.615
R234 VTAIL.n32 VTAIL.n31 104.615
R235 VTAIL.n116 VTAIL.n115 104.615
R236 VTAIL.n115 VTAIL.n89 104.615
R237 VTAIL.n108 VTAIL.n89 104.615
R238 VTAIL.n108 VTAIL.n107 104.615
R239 VTAIL.n107 VTAIL.n93 104.615
R240 VTAIL.n100 VTAIL.n93 104.615
R241 VTAIL.n100 VTAIL.n99 104.615
R242 VTAIL.n76 VTAIL.n75 104.615
R243 VTAIL.n75 VTAIL.n49 104.615
R244 VTAIL.n68 VTAIL.n49 104.615
R245 VTAIL.n68 VTAIL.n67 104.615
R246 VTAIL.n67 VTAIL.n53 104.615
R247 VTAIL.n60 VTAIL.n53 104.615
R248 VTAIL.n60 VTAIL.n59 104.615
R249 VTAIL.n135 VTAIL.t5 52.3082
R250 VTAIL.n15 VTAIL.t15 52.3082
R251 VTAIL.n99 VTAIL.t10 52.3082
R252 VTAIL.n59 VTAIL.t9 52.3082
R253 VTAIL.n85 VTAIL.n84 49.5893
R254 VTAIL.n83 VTAIL.n82 49.5893
R255 VTAIL.n45 VTAIL.n44 49.5893
R256 VTAIL.n43 VTAIL.n42 49.5893
R257 VTAIL.n159 VTAIL.n158 49.5891
R258 VTAIL.n1 VTAIL.n0 49.5891
R259 VTAIL.n39 VTAIL.n38 49.5891
R260 VTAIL.n41 VTAIL.n40 49.5891
R261 VTAIL.n157 VTAIL.n156 32.3793
R262 VTAIL.n37 VTAIL.n36 32.3793
R263 VTAIL.n121 VTAIL.n120 32.3793
R264 VTAIL.n81 VTAIL.n80 32.3793
R265 VTAIL.n43 VTAIL.n41 24.5479
R266 VTAIL.n157 VTAIL.n121 21.3583
R267 VTAIL.n134 VTAIL.n133 15.6676
R268 VTAIL.n14 VTAIL.n13 15.6676
R269 VTAIL.n98 VTAIL.n97 15.6676
R270 VTAIL.n58 VTAIL.n57 15.6676
R271 VTAIL.n137 VTAIL.n132 12.8005
R272 VTAIL.n17 VTAIL.n12 12.8005
R273 VTAIL.n101 VTAIL.n96 12.8005
R274 VTAIL.n61 VTAIL.n56 12.8005
R275 VTAIL.n138 VTAIL.n130 12.0247
R276 VTAIL.n18 VTAIL.n10 12.0247
R277 VTAIL.n102 VTAIL.n94 12.0247
R278 VTAIL.n62 VTAIL.n54 12.0247
R279 VTAIL.n142 VTAIL.n141 11.249
R280 VTAIL.n22 VTAIL.n21 11.249
R281 VTAIL.n106 VTAIL.n105 11.249
R282 VTAIL.n66 VTAIL.n65 11.249
R283 VTAIL.n145 VTAIL.n128 10.4732
R284 VTAIL.n25 VTAIL.n8 10.4732
R285 VTAIL.n109 VTAIL.n92 10.4732
R286 VTAIL.n69 VTAIL.n52 10.4732
R287 VTAIL.n146 VTAIL.n126 9.69747
R288 VTAIL.n26 VTAIL.n6 9.69747
R289 VTAIL.n110 VTAIL.n90 9.69747
R290 VTAIL.n70 VTAIL.n50 9.69747
R291 VTAIL.n156 VTAIL.n155 9.45567
R292 VTAIL.n36 VTAIL.n35 9.45567
R293 VTAIL.n120 VTAIL.n119 9.45567
R294 VTAIL.n80 VTAIL.n79 9.45567
R295 VTAIL.n124 VTAIL.n123 9.3005
R296 VTAIL.n149 VTAIL.n148 9.3005
R297 VTAIL.n147 VTAIL.n146 9.3005
R298 VTAIL.n128 VTAIL.n127 9.3005
R299 VTAIL.n141 VTAIL.n140 9.3005
R300 VTAIL.n139 VTAIL.n138 9.3005
R301 VTAIL.n132 VTAIL.n131 9.3005
R302 VTAIL.n155 VTAIL.n154 9.3005
R303 VTAIL.n4 VTAIL.n3 9.3005
R304 VTAIL.n29 VTAIL.n28 9.3005
R305 VTAIL.n27 VTAIL.n26 9.3005
R306 VTAIL.n8 VTAIL.n7 9.3005
R307 VTAIL.n21 VTAIL.n20 9.3005
R308 VTAIL.n19 VTAIL.n18 9.3005
R309 VTAIL.n12 VTAIL.n11 9.3005
R310 VTAIL.n35 VTAIL.n34 9.3005
R311 VTAIL.n119 VTAIL.n118 9.3005
R312 VTAIL.n88 VTAIL.n87 9.3005
R313 VTAIL.n113 VTAIL.n112 9.3005
R314 VTAIL.n111 VTAIL.n110 9.3005
R315 VTAIL.n92 VTAIL.n91 9.3005
R316 VTAIL.n105 VTAIL.n104 9.3005
R317 VTAIL.n103 VTAIL.n102 9.3005
R318 VTAIL.n96 VTAIL.n95 9.3005
R319 VTAIL.n79 VTAIL.n78 9.3005
R320 VTAIL.n48 VTAIL.n47 9.3005
R321 VTAIL.n73 VTAIL.n72 9.3005
R322 VTAIL.n71 VTAIL.n70 9.3005
R323 VTAIL.n52 VTAIL.n51 9.3005
R324 VTAIL.n65 VTAIL.n64 9.3005
R325 VTAIL.n63 VTAIL.n62 9.3005
R326 VTAIL.n56 VTAIL.n55 9.3005
R327 VTAIL.n150 VTAIL.n149 8.92171
R328 VTAIL.n30 VTAIL.n29 8.92171
R329 VTAIL.n114 VTAIL.n113 8.92171
R330 VTAIL.n74 VTAIL.n73 8.92171
R331 VTAIL.n153 VTAIL.n124 8.14595
R332 VTAIL.n33 VTAIL.n4 8.14595
R333 VTAIL.n117 VTAIL.n88 8.14595
R334 VTAIL.n77 VTAIL.n48 8.14595
R335 VTAIL.n154 VTAIL.n122 7.3702
R336 VTAIL.n34 VTAIL.n2 7.3702
R337 VTAIL.n118 VTAIL.n86 7.3702
R338 VTAIL.n78 VTAIL.n46 7.3702
R339 VTAIL.n156 VTAIL.n122 6.59444
R340 VTAIL.n36 VTAIL.n2 6.59444
R341 VTAIL.n120 VTAIL.n86 6.59444
R342 VTAIL.n80 VTAIL.n46 6.59444
R343 VTAIL.n154 VTAIL.n153 5.81868
R344 VTAIL.n34 VTAIL.n33 5.81868
R345 VTAIL.n118 VTAIL.n117 5.81868
R346 VTAIL.n78 VTAIL.n77 5.81868
R347 VTAIL.n150 VTAIL.n124 5.04292
R348 VTAIL.n30 VTAIL.n4 5.04292
R349 VTAIL.n114 VTAIL.n88 5.04292
R350 VTAIL.n74 VTAIL.n48 5.04292
R351 VTAIL.n133 VTAIL.n131 4.38571
R352 VTAIL.n13 VTAIL.n11 4.38571
R353 VTAIL.n97 VTAIL.n95 4.38571
R354 VTAIL.n57 VTAIL.n55 4.38571
R355 VTAIL.n149 VTAIL.n126 4.26717
R356 VTAIL.n29 VTAIL.n6 4.26717
R357 VTAIL.n113 VTAIL.n90 4.26717
R358 VTAIL.n73 VTAIL.n50 4.26717
R359 VTAIL.n146 VTAIL.n145 3.49141
R360 VTAIL.n26 VTAIL.n25 3.49141
R361 VTAIL.n110 VTAIL.n109 3.49141
R362 VTAIL.n70 VTAIL.n69 3.49141
R363 VTAIL.n45 VTAIL.n43 3.19016
R364 VTAIL.n81 VTAIL.n45 3.19016
R365 VTAIL.n85 VTAIL.n83 3.19016
R366 VTAIL.n121 VTAIL.n85 3.19016
R367 VTAIL.n41 VTAIL.n39 3.19016
R368 VTAIL.n39 VTAIL.n37 3.19016
R369 VTAIL.n159 VTAIL.n157 3.19016
R370 VTAIL.n158 VTAIL.t0 2.94255
R371 VTAIL.n158 VTAIL.t8 2.94255
R372 VTAIL.n0 VTAIL.t6 2.94255
R373 VTAIL.n0 VTAIL.t7 2.94255
R374 VTAIL.n38 VTAIL.t13 2.94255
R375 VTAIL.n38 VTAIL.t19 2.94255
R376 VTAIL.n40 VTAIL.t16 2.94255
R377 VTAIL.n40 VTAIL.t12 2.94255
R378 VTAIL.n84 VTAIL.t14 2.94255
R379 VTAIL.n84 VTAIL.t17 2.94255
R380 VTAIL.n82 VTAIL.t18 2.94255
R381 VTAIL.n82 VTAIL.t11 2.94255
R382 VTAIL.n44 VTAIL.t1 2.94255
R383 VTAIL.n44 VTAIL.t3 2.94255
R384 VTAIL.n42 VTAIL.t2 2.94255
R385 VTAIL.n42 VTAIL.t4 2.94255
R386 VTAIL.n142 VTAIL.n128 2.71565
R387 VTAIL.n22 VTAIL.n8 2.71565
R388 VTAIL.n106 VTAIL.n92 2.71565
R389 VTAIL.n66 VTAIL.n52 2.71565
R390 VTAIL VTAIL.n1 2.45093
R391 VTAIL.n83 VTAIL.n81 2.06516
R392 VTAIL.n37 VTAIL.n1 2.06516
R393 VTAIL.n141 VTAIL.n130 1.93989
R394 VTAIL.n21 VTAIL.n10 1.93989
R395 VTAIL.n105 VTAIL.n94 1.93989
R396 VTAIL.n65 VTAIL.n54 1.93989
R397 VTAIL.n138 VTAIL.n137 1.16414
R398 VTAIL.n18 VTAIL.n17 1.16414
R399 VTAIL.n102 VTAIL.n101 1.16414
R400 VTAIL.n62 VTAIL.n61 1.16414
R401 VTAIL VTAIL.n159 0.739724
R402 VTAIL.n134 VTAIL.n132 0.388379
R403 VTAIL.n14 VTAIL.n12 0.388379
R404 VTAIL.n98 VTAIL.n96 0.388379
R405 VTAIL.n58 VTAIL.n56 0.388379
R406 VTAIL.n139 VTAIL.n131 0.155672
R407 VTAIL.n140 VTAIL.n139 0.155672
R408 VTAIL.n140 VTAIL.n127 0.155672
R409 VTAIL.n147 VTAIL.n127 0.155672
R410 VTAIL.n148 VTAIL.n147 0.155672
R411 VTAIL.n148 VTAIL.n123 0.155672
R412 VTAIL.n155 VTAIL.n123 0.155672
R413 VTAIL.n19 VTAIL.n11 0.155672
R414 VTAIL.n20 VTAIL.n19 0.155672
R415 VTAIL.n20 VTAIL.n7 0.155672
R416 VTAIL.n27 VTAIL.n7 0.155672
R417 VTAIL.n28 VTAIL.n27 0.155672
R418 VTAIL.n28 VTAIL.n3 0.155672
R419 VTAIL.n35 VTAIL.n3 0.155672
R420 VTAIL.n119 VTAIL.n87 0.155672
R421 VTAIL.n112 VTAIL.n87 0.155672
R422 VTAIL.n112 VTAIL.n111 0.155672
R423 VTAIL.n111 VTAIL.n91 0.155672
R424 VTAIL.n104 VTAIL.n91 0.155672
R425 VTAIL.n104 VTAIL.n103 0.155672
R426 VTAIL.n103 VTAIL.n95 0.155672
R427 VTAIL.n79 VTAIL.n47 0.155672
R428 VTAIL.n72 VTAIL.n47 0.155672
R429 VTAIL.n72 VTAIL.n71 0.155672
R430 VTAIL.n71 VTAIL.n51 0.155672
R431 VTAIL.n64 VTAIL.n51 0.155672
R432 VTAIL.n64 VTAIL.n63 0.155672
R433 VTAIL.n63 VTAIL.n55 0.155672
R434 VDD1.n30 VDD1.n0 289.615
R435 VDD1.n67 VDD1.n37 289.615
R436 VDD1.n31 VDD1.n30 185
R437 VDD1.n29 VDD1.n28 185
R438 VDD1.n4 VDD1.n3 185
R439 VDD1.n23 VDD1.n22 185
R440 VDD1.n21 VDD1.n20 185
R441 VDD1.n8 VDD1.n7 185
R442 VDD1.n15 VDD1.n14 185
R443 VDD1.n13 VDD1.n12 185
R444 VDD1.n50 VDD1.n49 185
R445 VDD1.n52 VDD1.n51 185
R446 VDD1.n45 VDD1.n44 185
R447 VDD1.n58 VDD1.n57 185
R448 VDD1.n60 VDD1.n59 185
R449 VDD1.n41 VDD1.n40 185
R450 VDD1.n66 VDD1.n65 185
R451 VDD1.n68 VDD1.n67 185
R452 VDD1.n11 VDD1.t1 147.659
R453 VDD1.n48 VDD1.t0 147.659
R454 VDD1.n30 VDD1.n29 104.615
R455 VDD1.n29 VDD1.n3 104.615
R456 VDD1.n22 VDD1.n3 104.615
R457 VDD1.n22 VDD1.n21 104.615
R458 VDD1.n21 VDD1.n7 104.615
R459 VDD1.n14 VDD1.n7 104.615
R460 VDD1.n14 VDD1.n13 104.615
R461 VDD1.n51 VDD1.n50 104.615
R462 VDD1.n51 VDD1.n44 104.615
R463 VDD1.n58 VDD1.n44 104.615
R464 VDD1.n59 VDD1.n58 104.615
R465 VDD1.n59 VDD1.n40 104.615
R466 VDD1.n66 VDD1.n40 104.615
R467 VDD1.n67 VDD1.n66 104.615
R468 VDD1.n75 VDD1.n74 68.6048
R469 VDD1.n36 VDD1.n35 66.2681
R470 VDD1.n77 VDD1.n76 66.2679
R471 VDD1.n73 VDD1.n72 66.2679
R472 VDD1.n13 VDD1.t1 52.3082
R473 VDD1.n50 VDD1.t0 52.3082
R474 VDD1.n36 VDD1.n34 52.2477
R475 VDD1.n73 VDD1.n71 52.2477
R476 VDD1.n77 VDD1.n75 46.8457
R477 VDD1.n12 VDD1.n11 15.6676
R478 VDD1.n49 VDD1.n48 15.6676
R479 VDD1.n15 VDD1.n10 12.8005
R480 VDD1.n52 VDD1.n47 12.8005
R481 VDD1.n16 VDD1.n8 12.0247
R482 VDD1.n53 VDD1.n45 12.0247
R483 VDD1.n20 VDD1.n19 11.249
R484 VDD1.n57 VDD1.n56 11.249
R485 VDD1.n23 VDD1.n6 10.4732
R486 VDD1.n60 VDD1.n43 10.4732
R487 VDD1.n24 VDD1.n4 9.69747
R488 VDD1.n61 VDD1.n41 9.69747
R489 VDD1.n34 VDD1.n33 9.45567
R490 VDD1.n71 VDD1.n70 9.45567
R491 VDD1.n33 VDD1.n32 9.3005
R492 VDD1.n2 VDD1.n1 9.3005
R493 VDD1.n27 VDD1.n26 9.3005
R494 VDD1.n25 VDD1.n24 9.3005
R495 VDD1.n6 VDD1.n5 9.3005
R496 VDD1.n19 VDD1.n18 9.3005
R497 VDD1.n17 VDD1.n16 9.3005
R498 VDD1.n10 VDD1.n9 9.3005
R499 VDD1.n39 VDD1.n38 9.3005
R500 VDD1.n64 VDD1.n63 9.3005
R501 VDD1.n62 VDD1.n61 9.3005
R502 VDD1.n43 VDD1.n42 9.3005
R503 VDD1.n56 VDD1.n55 9.3005
R504 VDD1.n54 VDD1.n53 9.3005
R505 VDD1.n47 VDD1.n46 9.3005
R506 VDD1.n70 VDD1.n69 9.3005
R507 VDD1.n28 VDD1.n27 8.92171
R508 VDD1.n65 VDD1.n64 8.92171
R509 VDD1.n31 VDD1.n2 8.14595
R510 VDD1.n68 VDD1.n39 8.14595
R511 VDD1.n32 VDD1.n0 7.3702
R512 VDD1.n69 VDD1.n37 7.3702
R513 VDD1.n34 VDD1.n0 6.59444
R514 VDD1.n71 VDD1.n37 6.59444
R515 VDD1.n32 VDD1.n31 5.81868
R516 VDD1.n69 VDD1.n68 5.81868
R517 VDD1.n28 VDD1.n2 5.04292
R518 VDD1.n65 VDD1.n39 5.04292
R519 VDD1.n11 VDD1.n9 4.38571
R520 VDD1.n48 VDD1.n46 4.38571
R521 VDD1.n27 VDD1.n4 4.26717
R522 VDD1.n64 VDD1.n41 4.26717
R523 VDD1.n24 VDD1.n23 3.49141
R524 VDD1.n61 VDD1.n60 3.49141
R525 VDD1.n76 VDD1.t6 2.94255
R526 VDD1.n76 VDD1.t7 2.94255
R527 VDD1.n35 VDD1.t2 2.94255
R528 VDD1.n35 VDD1.t4 2.94255
R529 VDD1.n74 VDD1.t3 2.94255
R530 VDD1.n74 VDD1.t8 2.94255
R531 VDD1.n72 VDD1.t5 2.94255
R532 VDD1.n72 VDD1.t9 2.94255
R533 VDD1.n20 VDD1.n6 2.71565
R534 VDD1.n57 VDD1.n43 2.71565
R535 VDD1 VDD1.n77 2.33455
R536 VDD1.n19 VDD1.n8 1.93989
R537 VDD1.n56 VDD1.n45 1.93989
R538 VDD1.n16 VDD1.n15 1.16414
R539 VDD1.n53 VDD1.n52 1.16414
R540 VDD1 VDD1.n36 0.856103
R541 VDD1.n75 VDD1.n73 0.742568
R542 VDD1.n12 VDD1.n10 0.388379
R543 VDD1.n49 VDD1.n47 0.388379
R544 VDD1.n33 VDD1.n1 0.155672
R545 VDD1.n26 VDD1.n1 0.155672
R546 VDD1.n26 VDD1.n25 0.155672
R547 VDD1.n25 VDD1.n5 0.155672
R548 VDD1.n18 VDD1.n5 0.155672
R549 VDD1.n18 VDD1.n17 0.155672
R550 VDD1.n17 VDD1.n9 0.155672
R551 VDD1.n54 VDD1.n46 0.155672
R552 VDD1.n55 VDD1.n54 0.155672
R553 VDD1.n55 VDD1.n42 0.155672
R554 VDD1.n62 VDD1.n42 0.155672
R555 VDD1.n63 VDD1.n62 0.155672
R556 VDD1.n63 VDD1.n38 0.155672
R557 VDD1.n70 VDD1.n38 0.155672
R558 B.n910 B.n909 585
R559 B.n291 B.n164 585
R560 B.n290 B.n289 585
R561 B.n288 B.n287 585
R562 B.n286 B.n285 585
R563 B.n284 B.n283 585
R564 B.n282 B.n281 585
R565 B.n280 B.n279 585
R566 B.n278 B.n277 585
R567 B.n276 B.n275 585
R568 B.n274 B.n273 585
R569 B.n272 B.n271 585
R570 B.n270 B.n269 585
R571 B.n268 B.n267 585
R572 B.n266 B.n265 585
R573 B.n264 B.n263 585
R574 B.n262 B.n261 585
R575 B.n260 B.n259 585
R576 B.n258 B.n257 585
R577 B.n256 B.n255 585
R578 B.n254 B.n253 585
R579 B.n252 B.n251 585
R580 B.n250 B.n249 585
R581 B.n248 B.n247 585
R582 B.n246 B.n245 585
R583 B.n244 B.n243 585
R584 B.n242 B.n241 585
R585 B.n240 B.n239 585
R586 B.n238 B.n237 585
R587 B.n236 B.n235 585
R588 B.n234 B.n233 585
R589 B.n232 B.n231 585
R590 B.n230 B.n229 585
R591 B.n228 B.n227 585
R592 B.n226 B.n225 585
R593 B.n224 B.n223 585
R594 B.n222 B.n221 585
R595 B.n220 B.n219 585
R596 B.n218 B.n217 585
R597 B.n216 B.n215 585
R598 B.n214 B.n213 585
R599 B.n212 B.n211 585
R600 B.n210 B.n209 585
R601 B.n208 B.n207 585
R602 B.n206 B.n205 585
R603 B.n204 B.n203 585
R604 B.n202 B.n201 585
R605 B.n200 B.n199 585
R606 B.n198 B.n197 585
R607 B.n196 B.n195 585
R608 B.n194 B.n193 585
R609 B.n192 B.n191 585
R610 B.n190 B.n189 585
R611 B.n188 B.n187 585
R612 B.n186 B.n185 585
R613 B.n184 B.n183 585
R614 B.n182 B.n181 585
R615 B.n180 B.n179 585
R616 B.n178 B.n177 585
R617 B.n176 B.n175 585
R618 B.n174 B.n173 585
R619 B.n172 B.n171 585
R620 B.n908 B.n133 585
R621 B.n913 B.n133 585
R622 B.n907 B.n132 585
R623 B.n914 B.n132 585
R624 B.n906 B.n905 585
R625 B.n905 B.n128 585
R626 B.n904 B.n127 585
R627 B.n920 B.n127 585
R628 B.n903 B.n126 585
R629 B.n921 B.n126 585
R630 B.n902 B.n125 585
R631 B.n922 B.n125 585
R632 B.n901 B.n900 585
R633 B.n900 B.n121 585
R634 B.n899 B.n120 585
R635 B.n928 B.n120 585
R636 B.n898 B.n119 585
R637 B.n929 B.n119 585
R638 B.n897 B.n118 585
R639 B.n930 B.n118 585
R640 B.n896 B.n895 585
R641 B.n895 B.n114 585
R642 B.n894 B.n113 585
R643 B.n936 B.n113 585
R644 B.n893 B.n112 585
R645 B.n937 B.n112 585
R646 B.n892 B.n111 585
R647 B.n938 B.n111 585
R648 B.n891 B.n890 585
R649 B.n890 B.n107 585
R650 B.n889 B.n106 585
R651 B.n944 B.n106 585
R652 B.n888 B.n105 585
R653 B.n945 B.n105 585
R654 B.n887 B.n104 585
R655 B.n946 B.n104 585
R656 B.n886 B.n885 585
R657 B.n885 B.n100 585
R658 B.n884 B.n99 585
R659 B.n952 B.n99 585
R660 B.n883 B.n98 585
R661 B.n953 B.n98 585
R662 B.n882 B.n97 585
R663 B.n954 B.n97 585
R664 B.n881 B.n880 585
R665 B.n880 B.n96 585
R666 B.n879 B.n92 585
R667 B.n960 B.n92 585
R668 B.n878 B.n91 585
R669 B.n961 B.n91 585
R670 B.n877 B.n90 585
R671 B.n962 B.n90 585
R672 B.n876 B.n875 585
R673 B.n875 B.n86 585
R674 B.n874 B.n85 585
R675 B.n968 B.n85 585
R676 B.n873 B.n84 585
R677 B.n969 B.n84 585
R678 B.n872 B.n83 585
R679 B.n970 B.n83 585
R680 B.n871 B.n870 585
R681 B.n870 B.n79 585
R682 B.n869 B.n78 585
R683 B.n976 B.n78 585
R684 B.n868 B.n77 585
R685 B.n977 B.n77 585
R686 B.n867 B.n76 585
R687 B.n978 B.n76 585
R688 B.n866 B.n865 585
R689 B.n865 B.n72 585
R690 B.n864 B.n71 585
R691 B.n984 B.n71 585
R692 B.n863 B.n70 585
R693 B.n985 B.n70 585
R694 B.n862 B.n69 585
R695 B.n986 B.n69 585
R696 B.n861 B.n860 585
R697 B.n860 B.n65 585
R698 B.n859 B.n64 585
R699 B.n992 B.n64 585
R700 B.n858 B.n63 585
R701 B.n993 B.n63 585
R702 B.n857 B.n62 585
R703 B.n994 B.n62 585
R704 B.n856 B.n855 585
R705 B.n855 B.n58 585
R706 B.n854 B.n57 585
R707 B.n1000 B.n57 585
R708 B.n853 B.n56 585
R709 B.n1001 B.n56 585
R710 B.n852 B.n55 585
R711 B.n1002 B.n55 585
R712 B.n851 B.n850 585
R713 B.n850 B.n51 585
R714 B.n849 B.n50 585
R715 B.n1008 B.n50 585
R716 B.n848 B.n49 585
R717 B.n1009 B.n49 585
R718 B.n847 B.n48 585
R719 B.n1010 B.n48 585
R720 B.n846 B.n845 585
R721 B.n845 B.n44 585
R722 B.n844 B.n43 585
R723 B.n1016 B.n43 585
R724 B.n843 B.n42 585
R725 B.n1017 B.n42 585
R726 B.n842 B.n41 585
R727 B.n1018 B.n41 585
R728 B.n841 B.n840 585
R729 B.n840 B.n37 585
R730 B.n839 B.n36 585
R731 B.n1024 B.n36 585
R732 B.n838 B.n35 585
R733 B.n1025 B.n35 585
R734 B.n837 B.n34 585
R735 B.n1026 B.n34 585
R736 B.n836 B.n835 585
R737 B.n835 B.n30 585
R738 B.n834 B.n29 585
R739 B.n1032 B.n29 585
R740 B.n833 B.n28 585
R741 B.n1033 B.n28 585
R742 B.n832 B.n27 585
R743 B.n1034 B.n27 585
R744 B.n831 B.n830 585
R745 B.n830 B.n23 585
R746 B.n829 B.n22 585
R747 B.n1040 B.n22 585
R748 B.n828 B.n21 585
R749 B.n1041 B.n21 585
R750 B.n827 B.n20 585
R751 B.n1042 B.n20 585
R752 B.n826 B.n825 585
R753 B.n825 B.n19 585
R754 B.n824 B.n15 585
R755 B.n1048 B.n15 585
R756 B.n823 B.n14 585
R757 B.n1049 B.n14 585
R758 B.n822 B.n13 585
R759 B.n1050 B.n13 585
R760 B.n821 B.n820 585
R761 B.n820 B.n12 585
R762 B.n819 B.n818 585
R763 B.n819 B.n8 585
R764 B.n817 B.n7 585
R765 B.n1057 B.n7 585
R766 B.n816 B.n6 585
R767 B.n1058 B.n6 585
R768 B.n815 B.n5 585
R769 B.n1059 B.n5 585
R770 B.n814 B.n813 585
R771 B.n813 B.n4 585
R772 B.n812 B.n292 585
R773 B.n812 B.n811 585
R774 B.n802 B.n293 585
R775 B.n294 B.n293 585
R776 B.n804 B.n803 585
R777 B.n805 B.n804 585
R778 B.n801 B.n299 585
R779 B.n299 B.n298 585
R780 B.n800 B.n799 585
R781 B.n799 B.n798 585
R782 B.n301 B.n300 585
R783 B.n791 B.n301 585
R784 B.n790 B.n789 585
R785 B.n792 B.n790 585
R786 B.n788 B.n306 585
R787 B.n306 B.n305 585
R788 B.n787 B.n786 585
R789 B.n786 B.n785 585
R790 B.n308 B.n307 585
R791 B.n309 B.n308 585
R792 B.n778 B.n777 585
R793 B.n779 B.n778 585
R794 B.n776 B.n314 585
R795 B.n314 B.n313 585
R796 B.n775 B.n774 585
R797 B.n774 B.n773 585
R798 B.n316 B.n315 585
R799 B.n317 B.n316 585
R800 B.n766 B.n765 585
R801 B.n767 B.n766 585
R802 B.n764 B.n322 585
R803 B.n322 B.n321 585
R804 B.n763 B.n762 585
R805 B.n762 B.n761 585
R806 B.n324 B.n323 585
R807 B.n325 B.n324 585
R808 B.n754 B.n753 585
R809 B.n755 B.n754 585
R810 B.n752 B.n330 585
R811 B.n330 B.n329 585
R812 B.n751 B.n750 585
R813 B.n750 B.n749 585
R814 B.n332 B.n331 585
R815 B.n333 B.n332 585
R816 B.n742 B.n741 585
R817 B.n743 B.n742 585
R818 B.n740 B.n338 585
R819 B.n338 B.n337 585
R820 B.n739 B.n738 585
R821 B.n738 B.n737 585
R822 B.n340 B.n339 585
R823 B.n341 B.n340 585
R824 B.n730 B.n729 585
R825 B.n731 B.n730 585
R826 B.n728 B.n345 585
R827 B.n349 B.n345 585
R828 B.n727 B.n726 585
R829 B.n726 B.n725 585
R830 B.n347 B.n346 585
R831 B.n348 B.n347 585
R832 B.n718 B.n717 585
R833 B.n719 B.n718 585
R834 B.n716 B.n354 585
R835 B.n354 B.n353 585
R836 B.n715 B.n714 585
R837 B.n714 B.n713 585
R838 B.n356 B.n355 585
R839 B.n357 B.n356 585
R840 B.n706 B.n705 585
R841 B.n707 B.n706 585
R842 B.n704 B.n362 585
R843 B.n362 B.n361 585
R844 B.n703 B.n702 585
R845 B.n702 B.n701 585
R846 B.n364 B.n363 585
R847 B.n365 B.n364 585
R848 B.n694 B.n693 585
R849 B.n695 B.n694 585
R850 B.n692 B.n370 585
R851 B.n370 B.n369 585
R852 B.n691 B.n690 585
R853 B.n690 B.n689 585
R854 B.n372 B.n371 585
R855 B.n373 B.n372 585
R856 B.n682 B.n681 585
R857 B.n683 B.n682 585
R858 B.n680 B.n378 585
R859 B.n378 B.n377 585
R860 B.n679 B.n678 585
R861 B.n678 B.n677 585
R862 B.n380 B.n379 585
R863 B.n381 B.n380 585
R864 B.n670 B.n669 585
R865 B.n671 B.n670 585
R866 B.n668 B.n386 585
R867 B.n386 B.n385 585
R868 B.n667 B.n666 585
R869 B.n666 B.n665 585
R870 B.n388 B.n387 585
R871 B.n658 B.n388 585
R872 B.n657 B.n656 585
R873 B.n659 B.n657 585
R874 B.n655 B.n393 585
R875 B.n393 B.n392 585
R876 B.n654 B.n653 585
R877 B.n653 B.n652 585
R878 B.n395 B.n394 585
R879 B.n396 B.n395 585
R880 B.n645 B.n644 585
R881 B.n646 B.n645 585
R882 B.n643 B.n401 585
R883 B.n401 B.n400 585
R884 B.n642 B.n641 585
R885 B.n641 B.n640 585
R886 B.n403 B.n402 585
R887 B.n404 B.n403 585
R888 B.n633 B.n632 585
R889 B.n634 B.n633 585
R890 B.n631 B.n409 585
R891 B.n409 B.n408 585
R892 B.n630 B.n629 585
R893 B.n629 B.n628 585
R894 B.n411 B.n410 585
R895 B.n412 B.n411 585
R896 B.n621 B.n620 585
R897 B.n622 B.n621 585
R898 B.n619 B.n416 585
R899 B.n420 B.n416 585
R900 B.n618 B.n617 585
R901 B.n617 B.n616 585
R902 B.n418 B.n417 585
R903 B.n419 B.n418 585
R904 B.n609 B.n608 585
R905 B.n610 B.n609 585
R906 B.n607 B.n425 585
R907 B.n425 B.n424 585
R908 B.n606 B.n605 585
R909 B.n605 B.n604 585
R910 B.n427 B.n426 585
R911 B.n428 B.n427 585
R912 B.n597 B.n596 585
R913 B.n598 B.n597 585
R914 B.n595 B.n433 585
R915 B.n433 B.n432 585
R916 B.n590 B.n589 585
R917 B.n588 B.n466 585
R918 B.n587 B.n465 585
R919 B.n592 B.n465 585
R920 B.n586 B.n585 585
R921 B.n584 B.n583 585
R922 B.n582 B.n581 585
R923 B.n580 B.n579 585
R924 B.n578 B.n577 585
R925 B.n576 B.n575 585
R926 B.n574 B.n573 585
R927 B.n572 B.n571 585
R928 B.n570 B.n569 585
R929 B.n568 B.n567 585
R930 B.n566 B.n565 585
R931 B.n564 B.n563 585
R932 B.n562 B.n561 585
R933 B.n560 B.n559 585
R934 B.n558 B.n557 585
R935 B.n556 B.n555 585
R936 B.n554 B.n553 585
R937 B.n552 B.n551 585
R938 B.n550 B.n549 585
R939 B.n548 B.n547 585
R940 B.n546 B.n545 585
R941 B.n544 B.n543 585
R942 B.n542 B.n541 585
R943 B.n539 B.n538 585
R944 B.n537 B.n536 585
R945 B.n535 B.n534 585
R946 B.n533 B.n532 585
R947 B.n531 B.n530 585
R948 B.n529 B.n528 585
R949 B.n527 B.n526 585
R950 B.n525 B.n524 585
R951 B.n523 B.n522 585
R952 B.n521 B.n520 585
R953 B.n518 B.n517 585
R954 B.n516 B.n515 585
R955 B.n514 B.n513 585
R956 B.n512 B.n511 585
R957 B.n510 B.n509 585
R958 B.n508 B.n507 585
R959 B.n506 B.n505 585
R960 B.n504 B.n503 585
R961 B.n502 B.n501 585
R962 B.n500 B.n499 585
R963 B.n498 B.n497 585
R964 B.n496 B.n495 585
R965 B.n494 B.n493 585
R966 B.n492 B.n491 585
R967 B.n490 B.n489 585
R968 B.n488 B.n487 585
R969 B.n486 B.n485 585
R970 B.n484 B.n483 585
R971 B.n482 B.n481 585
R972 B.n480 B.n479 585
R973 B.n478 B.n477 585
R974 B.n476 B.n475 585
R975 B.n474 B.n473 585
R976 B.n472 B.n471 585
R977 B.n435 B.n434 585
R978 B.n594 B.n593 585
R979 B.n593 B.n592 585
R980 B.n431 B.n430 585
R981 B.n432 B.n431 585
R982 B.n600 B.n599 585
R983 B.n599 B.n598 585
R984 B.n601 B.n429 585
R985 B.n429 B.n428 585
R986 B.n603 B.n602 585
R987 B.n604 B.n603 585
R988 B.n423 B.n422 585
R989 B.n424 B.n423 585
R990 B.n612 B.n611 585
R991 B.n611 B.n610 585
R992 B.n613 B.n421 585
R993 B.n421 B.n419 585
R994 B.n615 B.n614 585
R995 B.n616 B.n615 585
R996 B.n415 B.n414 585
R997 B.n420 B.n415 585
R998 B.n624 B.n623 585
R999 B.n623 B.n622 585
R1000 B.n625 B.n413 585
R1001 B.n413 B.n412 585
R1002 B.n627 B.n626 585
R1003 B.n628 B.n627 585
R1004 B.n407 B.n406 585
R1005 B.n408 B.n407 585
R1006 B.n636 B.n635 585
R1007 B.n635 B.n634 585
R1008 B.n637 B.n405 585
R1009 B.n405 B.n404 585
R1010 B.n639 B.n638 585
R1011 B.n640 B.n639 585
R1012 B.n399 B.n398 585
R1013 B.n400 B.n399 585
R1014 B.n648 B.n647 585
R1015 B.n647 B.n646 585
R1016 B.n649 B.n397 585
R1017 B.n397 B.n396 585
R1018 B.n651 B.n650 585
R1019 B.n652 B.n651 585
R1020 B.n391 B.n390 585
R1021 B.n392 B.n391 585
R1022 B.n661 B.n660 585
R1023 B.n660 B.n659 585
R1024 B.n662 B.n389 585
R1025 B.n658 B.n389 585
R1026 B.n664 B.n663 585
R1027 B.n665 B.n664 585
R1028 B.n384 B.n383 585
R1029 B.n385 B.n384 585
R1030 B.n673 B.n672 585
R1031 B.n672 B.n671 585
R1032 B.n674 B.n382 585
R1033 B.n382 B.n381 585
R1034 B.n676 B.n675 585
R1035 B.n677 B.n676 585
R1036 B.n376 B.n375 585
R1037 B.n377 B.n376 585
R1038 B.n685 B.n684 585
R1039 B.n684 B.n683 585
R1040 B.n686 B.n374 585
R1041 B.n374 B.n373 585
R1042 B.n688 B.n687 585
R1043 B.n689 B.n688 585
R1044 B.n368 B.n367 585
R1045 B.n369 B.n368 585
R1046 B.n697 B.n696 585
R1047 B.n696 B.n695 585
R1048 B.n698 B.n366 585
R1049 B.n366 B.n365 585
R1050 B.n700 B.n699 585
R1051 B.n701 B.n700 585
R1052 B.n360 B.n359 585
R1053 B.n361 B.n360 585
R1054 B.n709 B.n708 585
R1055 B.n708 B.n707 585
R1056 B.n710 B.n358 585
R1057 B.n358 B.n357 585
R1058 B.n712 B.n711 585
R1059 B.n713 B.n712 585
R1060 B.n352 B.n351 585
R1061 B.n353 B.n352 585
R1062 B.n721 B.n720 585
R1063 B.n720 B.n719 585
R1064 B.n722 B.n350 585
R1065 B.n350 B.n348 585
R1066 B.n724 B.n723 585
R1067 B.n725 B.n724 585
R1068 B.n344 B.n343 585
R1069 B.n349 B.n344 585
R1070 B.n733 B.n732 585
R1071 B.n732 B.n731 585
R1072 B.n734 B.n342 585
R1073 B.n342 B.n341 585
R1074 B.n736 B.n735 585
R1075 B.n737 B.n736 585
R1076 B.n336 B.n335 585
R1077 B.n337 B.n336 585
R1078 B.n745 B.n744 585
R1079 B.n744 B.n743 585
R1080 B.n746 B.n334 585
R1081 B.n334 B.n333 585
R1082 B.n748 B.n747 585
R1083 B.n749 B.n748 585
R1084 B.n328 B.n327 585
R1085 B.n329 B.n328 585
R1086 B.n757 B.n756 585
R1087 B.n756 B.n755 585
R1088 B.n758 B.n326 585
R1089 B.n326 B.n325 585
R1090 B.n760 B.n759 585
R1091 B.n761 B.n760 585
R1092 B.n320 B.n319 585
R1093 B.n321 B.n320 585
R1094 B.n769 B.n768 585
R1095 B.n768 B.n767 585
R1096 B.n770 B.n318 585
R1097 B.n318 B.n317 585
R1098 B.n772 B.n771 585
R1099 B.n773 B.n772 585
R1100 B.n312 B.n311 585
R1101 B.n313 B.n312 585
R1102 B.n781 B.n780 585
R1103 B.n780 B.n779 585
R1104 B.n782 B.n310 585
R1105 B.n310 B.n309 585
R1106 B.n784 B.n783 585
R1107 B.n785 B.n784 585
R1108 B.n304 B.n303 585
R1109 B.n305 B.n304 585
R1110 B.n794 B.n793 585
R1111 B.n793 B.n792 585
R1112 B.n795 B.n302 585
R1113 B.n791 B.n302 585
R1114 B.n797 B.n796 585
R1115 B.n798 B.n797 585
R1116 B.n297 B.n296 585
R1117 B.n298 B.n297 585
R1118 B.n807 B.n806 585
R1119 B.n806 B.n805 585
R1120 B.n808 B.n295 585
R1121 B.n295 B.n294 585
R1122 B.n810 B.n809 585
R1123 B.n811 B.n810 585
R1124 B.n3 B.n0 585
R1125 B.n4 B.n3 585
R1126 B.n1056 B.n1 585
R1127 B.n1057 B.n1056 585
R1128 B.n1055 B.n1054 585
R1129 B.n1055 B.n8 585
R1130 B.n1053 B.n9 585
R1131 B.n12 B.n9 585
R1132 B.n1052 B.n1051 585
R1133 B.n1051 B.n1050 585
R1134 B.n11 B.n10 585
R1135 B.n1049 B.n11 585
R1136 B.n1047 B.n1046 585
R1137 B.n1048 B.n1047 585
R1138 B.n1045 B.n16 585
R1139 B.n19 B.n16 585
R1140 B.n1044 B.n1043 585
R1141 B.n1043 B.n1042 585
R1142 B.n18 B.n17 585
R1143 B.n1041 B.n18 585
R1144 B.n1039 B.n1038 585
R1145 B.n1040 B.n1039 585
R1146 B.n1037 B.n24 585
R1147 B.n24 B.n23 585
R1148 B.n1036 B.n1035 585
R1149 B.n1035 B.n1034 585
R1150 B.n26 B.n25 585
R1151 B.n1033 B.n26 585
R1152 B.n1031 B.n1030 585
R1153 B.n1032 B.n1031 585
R1154 B.n1029 B.n31 585
R1155 B.n31 B.n30 585
R1156 B.n1028 B.n1027 585
R1157 B.n1027 B.n1026 585
R1158 B.n33 B.n32 585
R1159 B.n1025 B.n33 585
R1160 B.n1023 B.n1022 585
R1161 B.n1024 B.n1023 585
R1162 B.n1021 B.n38 585
R1163 B.n38 B.n37 585
R1164 B.n1020 B.n1019 585
R1165 B.n1019 B.n1018 585
R1166 B.n40 B.n39 585
R1167 B.n1017 B.n40 585
R1168 B.n1015 B.n1014 585
R1169 B.n1016 B.n1015 585
R1170 B.n1013 B.n45 585
R1171 B.n45 B.n44 585
R1172 B.n1012 B.n1011 585
R1173 B.n1011 B.n1010 585
R1174 B.n47 B.n46 585
R1175 B.n1009 B.n47 585
R1176 B.n1007 B.n1006 585
R1177 B.n1008 B.n1007 585
R1178 B.n1005 B.n52 585
R1179 B.n52 B.n51 585
R1180 B.n1004 B.n1003 585
R1181 B.n1003 B.n1002 585
R1182 B.n54 B.n53 585
R1183 B.n1001 B.n54 585
R1184 B.n999 B.n998 585
R1185 B.n1000 B.n999 585
R1186 B.n997 B.n59 585
R1187 B.n59 B.n58 585
R1188 B.n996 B.n995 585
R1189 B.n995 B.n994 585
R1190 B.n61 B.n60 585
R1191 B.n993 B.n61 585
R1192 B.n991 B.n990 585
R1193 B.n992 B.n991 585
R1194 B.n989 B.n66 585
R1195 B.n66 B.n65 585
R1196 B.n988 B.n987 585
R1197 B.n987 B.n986 585
R1198 B.n68 B.n67 585
R1199 B.n985 B.n68 585
R1200 B.n983 B.n982 585
R1201 B.n984 B.n983 585
R1202 B.n981 B.n73 585
R1203 B.n73 B.n72 585
R1204 B.n980 B.n979 585
R1205 B.n979 B.n978 585
R1206 B.n75 B.n74 585
R1207 B.n977 B.n75 585
R1208 B.n975 B.n974 585
R1209 B.n976 B.n975 585
R1210 B.n973 B.n80 585
R1211 B.n80 B.n79 585
R1212 B.n972 B.n971 585
R1213 B.n971 B.n970 585
R1214 B.n82 B.n81 585
R1215 B.n969 B.n82 585
R1216 B.n967 B.n966 585
R1217 B.n968 B.n967 585
R1218 B.n965 B.n87 585
R1219 B.n87 B.n86 585
R1220 B.n964 B.n963 585
R1221 B.n963 B.n962 585
R1222 B.n89 B.n88 585
R1223 B.n961 B.n89 585
R1224 B.n959 B.n958 585
R1225 B.n960 B.n959 585
R1226 B.n957 B.n93 585
R1227 B.n96 B.n93 585
R1228 B.n956 B.n955 585
R1229 B.n955 B.n954 585
R1230 B.n95 B.n94 585
R1231 B.n953 B.n95 585
R1232 B.n951 B.n950 585
R1233 B.n952 B.n951 585
R1234 B.n949 B.n101 585
R1235 B.n101 B.n100 585
R1236 B.n948 B.n947 585
R1237 B.n947 B.n946 585
R1238 B.n103 B.n102 585
R1239 B.n945 B.n103 585
R1240 B.n943 B.n942 585
R1241 B.n944 B.n943 585
R1242 B.n941 B.n108 585
R1243 B.n108 B.n107 585
R1244 B.n940 B.n939 585
R1245 B.n939 B.n938 585
R1246 B.n110 B.n109 585
R1247 B.n937 B.n110 585
R1248 B.n935 B.n934 585
R1249 B.n936 B.n935 585
R1250 B.n933 B.n115 585
R1251 B.n115 B.n114 585
R1252 B.n932 B.n931 585
R1253 B.n931 B.n930 585
R1254 B.n117 B.n116 585
R1255 B.n929 B.n117 585
R1256 B.n927 B.n926 585
R1257 B.n928 B.n927 585
R1258 B.n925 B.n122 585
R1259 B.n122 B.n121 585
R1260 B.n924 B.n923 585
R1261 B.n923 B.n922 585
R1262 B.n124 B.n123 585
R1263 B.n921 B.n124 585
R1264 B.n919 B.n918 585
R1265 B.n920 B.n919 585
R1266 B.n917 B.n129 585
R1267 B.n129 B.n128 585
R1268 B.n916 B.n915 585
R1269 B.n915 B.n914 585
R1270 B.n131 B.n130 585
R1271 B.n913 B.n131 585
R1272 B.n1060 B.n1059 585
R1273 B.n1058 B.n2 585
R1274 B.n171 B.n131 468.476
R1275 B.n910 B.n133 468.476
R1276 B.n593 B.n433 468.476
R1277 B.n590 B.n431 468.476
R1278 B.n165 B.t15 263.392
R1279 B.n469 B.t23 263.392
R1280 B.n168 B.t12 263.392
R1281 B.n467 B.t20 263.392
R1282 B.n168 B.t10 257.101
R1283 B.n165 B.t14 257.101
R1284 B.n469 B.t21 257.101
R1285 B.n467 B.t17 257.101
R1286 B.n912 B.n911 256.663
R1287 B.n912 B.n163 256.663
R1288 B.n912 B.n162 256.663
R1289 B.n912 B.n161 256.663
R1290 B.n912 B.n160 256.663
R1291 B.n912 B.n159 256.663
R1292 B.n912 B.n158 256.663
R1293 B.n912 B.n157 256.663
R1294 B.n912 B.n156 256.663
R1295 B.n912 B.n155 256.663
R1296 B.n912 B.n154 256.663
R1297 B.n912 B.n153 256.663
R1298 B.n912 B.n152 256.663
R1299 B.n912 B.n151 256.663
R1300 B.n912 B.n150 256.663
R1301 B.n912 B.n149 256.663
R1302 B.n912 B.n148 256.663
R1303 B.n912 B.n147 256.663
R1304 B.n912 B.n146 256.663
R1305 B.n912 B.n145 256.663
R1306 B.n912 B.n144 256.663
R1307 B.n912 B.n143 256.663
R1308 B.n912 B.n142 256.663
R1309 B.n912 B.n141 256.663
R1310 B.n912 B.n140 256.663
R1311 B.n912 B.n139 256.663
R1312 B.n912 B.n138 256.663
R1313 B.n912 B.n137 256.663
R1314 B.n912 B.n136 256.663
R1315 B.n912 B.n135 256.663
R1316 B.n912 B.n134 256.663
R1317 B.n592 B.n591 256.663
R1318 B.n592 B.n436 256.663
R1319 B.n592 B.n437 256.663
R1320 B.n592 B.n438 256.663
R1321 B.n592 B.n439 256.663
R1322 B.n592 B.n440 256.663
R1323 B.n592 B.n441 256.663
R1324 B.n592 B.n442 256.663
R1325 B.n592 B.n443 256.663
R1326 B.n592 B.n444 256.663
R1327 B.n592 B.n445 256.663
R1328 B.n592 B.n446 256.663
R1329 B.n592 B.n447 256.663
R1330 B.n592 B.n448 256.663
R1331 B.n592 B.n449 256.663
R1332 B.n592 B.n450 256.663
R1333 B.n592 B.n451 256.663
R1334 B.n592 B.n452 256.663
R1335 B.n592 B.n453 256.663
R1336 B.n592 B.n454 256.663
R1337 B.n592 B.n455 256.663
R1338 B.n592 B.n456 256.663
R1339 B.n592 B.n457 256.663
R1340 B.n592 B.n458 256.663
R1341 B.n592 B.n459 256.663
R1342 B.n592 B.n460 256.663
R1343 B.n592 B.n461 256.663
R1344 B.n592 B.n462 256.663
R1345 B.n592 B.n463 256.663
R1346 B.n592 B.n464 256.663
R1347 B.n1062 B.n1061 256.663
R1348 B.n166 B.t16 191.635
R1349 B.n470 B.t22 191.635
R1350 B.n169 B.t13 191.635
R1351 B.n468 B.t19 191.635
R1352 B.n175 B.n174 163.367
R1353 B.n179 B.n178 163.367
R1354 B.n183 B.n182 163.367
R1355 B.n187 B.n186 163.367
R1356 B.n191 B.n190 163.367
R1357 B.n195 B.n194 163.367
R1358 B.n199 B.n198 163.367
R1359 B.n203 B.n202 163.367
R1360 B.n207 B.n206 163.367
R1361 B.n211 B.n210 163.367
R1362 B.n215 B.n214 163.367
R1363 B.n219 B.n218 163.367
R1364 B.n223 B.n222 163.367
R1365 B.n227 B.n226 163.367
R1366 B.n231 B.n230 163.367
R1367 B.n235 B.n234 163.367
R1368 B.n239 B.n238 163.367
R1369 B.n243 B.n242 163.367
R1370 B.n247 B.n246 163.367
R1371 B.n251 B.n250 163.367
R1372 B.n255 B.n254 163.367
R1373 B.n259 B.n258 163.367
R1374 B.n263 B.n262 163.367
R1375 B.n267 B.n266 163.367
R1376 B.n271 B.n270 163.367
R1377 B.n275 B.n274 163.367
R1378 B.n279 B.n278 163.367
R1379 B.n283 B.n282 163.367
R1380 B.n287 B.n286 163.367
R1381 B.n289 B.n164 163.367
R1382 B.n597 B.n433 163.367
R1383 B.n597 B.n427 163.367
R1384 B.n605 B.n427 163.367
R1385 B.n605 B.n425 163.367
R1386 B.n609 B.n425 163.367
R1387 B.n609 B.n418 163.367
R1388 B.n617 B.n418 163.367
R1389 B.n617 B.n416 163.367
R1390 B.n621 B.n416 163.367
R1391 B.n621 B.n411 163.367
R1392 B.n629 B.n411 163.367
R1393 B.n629 B.n409 163.367
R1394 B.n633 B.n409 163.367
R1395 B.n633 B.n403 163.367
R1396 B.n641 B.n403 163.367
R1397 B.n641 B.n401 163.367
R1398 B.n645 B.n401 163.367
R1399 B.n645 B.n395 163.367
R1400 B.n653 B.n395 163.367
R1401 B.n653 B.n393 163.367
R1402 B.n657 B.n393 163.367
R1403 B.n657 B.n388 163.367
R1404 B.n666 B.n388 163.367
R1405 B.n666 B.n386 163.367
R1406 B.n670 B.n386 163.367
R1407 B.n670 B.n380 163.367
R1408 B.n678 B.n380 163.367
R1409 B.n678 B.n378 163.367
R1410 B.n682 B.n378 163.367
R1411 B.n682 B.n372 163.367
R1412 B.n690 B.n372 163.367
R1413 B.n690 B.n370 163.367
R1414 B.n694 B.n370 163.367
R1415 B.n694 B.n364 163.367
R1416 B.n702 B.n364 163.367
R1417 B.n702 B.n362 163.367
R1418 B.n706 B.n362 163.367
R1419 B.n706 B.n356 163.367
R1420 B.n714 B.n356 163.367
R1421 B.n714 B.n354 163.367
R1422 B.n718 B.n354 163.367
R1423 B.n718 B.n347 163.367
R1424 B.n726 B.n347 163.367
R1425 B.n726 B.n345 163.367
R1426 B.n730 B.n345 163.367
R1427 B.n730 B.n340 163.367
R1428 B.n738 B.n340 163.367
R1429 B.n738 B.n338 163.367
R1430 B.n742 B.n338 163.367
R1431 B.n742 B.n332 163.367
R1432 B.n750 B.n332 163.367
R1433 B.n750 B.n330 163.367
R1434 B.n754 B.n330 163.367
R1435 B.n754 B.n324 163.367
R1436 B.n762 B.n324 163.367
R1437 B.n762 B.n322 163.367
R1438 B.n766 B.n322 163.367
R1439 B.n766 B.n316 163.367
R1440 B.n774 B.n316 163.367
R1441 B.n774 B.n314 163.367
R1442 B.n778 B.n314 163.367
R1443 B.n778 B.n308 163.367
R1444 B.n786 B.n308 163.367
R1445 B.n786 B.n306 163.367
R1446 B.n790 B.n306 163.367
R1447 B.n790 B.n301 163.367
R1448 B.n799 B.n301 163.367
R1449 B.n799 B.n299 163.367
R1450 B.n804 B.n299 163.367
R1451 B.n804 B.n293 163.367
R1452 B.n812 B.n293 163.367
R1453 B.n813 B.n812 163.367
R1454 B.n813 B.n5 163.367
R1455 B.n6 B.n5 163.367
R1456 B.n7 B.n6 163.367
R1457 B.n819 B.n7 163.367
R1458 B.n820 B.n819 163.367
R1459 B.n820 B.n13 163.367
R1460 B.n14 B.n13 163.367
R1461 B.n15 B.n14 163.367
R1462 B.n825 B.n15 163.367
R1463 B.n825 B.n20 163.367
R1464 B.n21 B.n20 163.367
R1465 B.n22 B.n21 163.367
R1466 B.n830 B.n22 163.367
R1467 B.n830 B.n27 163.367
R1468 B.n28 B.n27 163.367
R1469 B.n29 B.n28 163.367
R1470 B.n835 B.n29 163.367
R1471 B.n835 B.n34 163.367
R1472 B.n35 B.n34 163.367
R1473 B.n36 B.n35 163.367
R1474 B.n840 B.n36 163.367
R1475 B.n840 B.n41 163.367
R1476 B.n42 B.n41 163.367
R1477 B.n43 B.n42 163.367
R1478 B.n845 B.n43 163.367
R1479 B.n845 B.n48 163.367
R1480 B.n49 B.n48 163.367
R1481 B.n50 B.n49 163.367
R1482 B.n850 B.n50 163.367
R1483 B.n850 B.n55 163.367
R1484 B.n56 B.n55 163.367
R1485 B.n57 B.n56 163.367
R1486 B.n855 B.n57 163.367
R1487 B.n855 B.n62 163.367
R1488 B.n63 B.n62 163.367
R1489 B.n64 B.n63 163.367
R1490 B.n860 B.n64 163.367
R1491 B.n860 B.n69 163.367
R1492 B.n70 B.n69 163.367
R1493 B.n71 B.n70 163.367
R1494 B.n865 B.n71 163.367
R1495 B.n865 B.n76 163.367
R1496 B.n77 B.n76 163.367
R1497 B.n78 B.n77 163.367
R1498 B.n870 B.n78 163.367
R1499 B.n870 B.n83 163.367
R1500 B.n84 B.n83 163.367
R1501 B.n85 B.n84 163.367
R1502 B.n875 B.n85 163.367
R1503 B.n875 B.n90 163.367
R1504 B.n91 B.n90 163.367
R1505 B.n92 B.n91 163.367
R1506 B.n880 B.n92 163.367
R1507 B.n880 B.n97 163.367
R1508 B.n98 B.n97 163.367
R1509 B.n99 B.n98 163.367
R1510 B.n885 B.n99 163.367
R1511 B.n885 B.n104 163.367
R1512 B.n105 B.n104 163.367
R1513 B.n106 B.n105 163.367
R1514 B.n890 B.n106 163.367
R1515 B.n890 B.n111 163.367
R1516 B.n112 B.n111 163.367
R1517 B.n113 B.n112 163.367
R1518 B.n895 B.n113 163.367
R1519 B.n895 B.n118 163.367
R1520 B.n119 B.n118 163.367
R1521 B.n120 B.n119 163.367
R1522 B.n900 B.n120 163.367
R1523 B.n900 B.n125 163.367
R1524 B.n126 B.n125 163.367
R1525 B.n127 B.n126 163.367
R1526 B.n905 B.n127 163.367
R1527 B.n905 B.n132 163.367
R1528 B.n133 B.n132 163.367
R1529 B.n466 B.n465 163.367
R1530 B.n585 B.n465 163.367
R1531 B.n583 B.n582 163.367
R1532 B.n579 B.n578 163.367
R1533 B.n575 B.n574 163.367
R1534 B.n571 B.n570 163.367
R1535 B.n567 B.n566 163.367
R1536 B.n563 B.n562 163.367
R1537 B.n559 B.n558 163.367
R1538 B.n555 B.n554 163.367
R1539 B.n551 B.n550 163.367
R1540 B.n547 B.n546 163.367
R1541 B.n543 B.n542 163.367
R1542 B.n538 B.n537 163.367
R1543 B.n534 B.n533 163.367
R1544 B.n530 B.n529 163.367
R1545 B.n526 B.n525 163.367
R1546 B.n522 B.n521 163.367
R1547 B.n517 B.n516 163.367
R1548 B.n513 B.n512 163.367
R1549 B.n509 B.n508 163.367
R1550 B.n505 B.n504 163.367
R1551 B.n501 B.n500 163.367
R1552 B.n497 B.n496 163.367
R1553 B.n493 B.n492 163.367
R1554 B.n489 B.n488 163.367
R1555 B.n485 B.n484 163.367
R1556 B.n481 B.n480 163.367
R1557 B.n477 B.n476 163.367
R1558 B.n473 B.n472 163.367
R1559 B.n593 B.n435 163.367
R1560 B.n599 B.n431 163.367
R1561 B.n599 B.n429 163.367
R1562 B.n603 B.n429 163.367
R1563 B.n603 B.n423 163.367
R1564 B.n611 B.n423 163.367
R1565 B.n611 B.n421 163.367
R1566 B.n615 B.n421 163.367
R1567 B.n615 B.n415 163.367
R1568 B.n623 B.n415 163.367
R1569 B.n623 B.n413 163.367
R1570 B.n627 B.n413 163.367
R1571 B.n627 B.n407 163.367
R1572 B.n635 B.n407 163.367
R1573 B.n635 B.n405 163.367
R1574 B.n639 B.n405 163.367
R1575 B.n639 B.n399 163.367
R1576 B.n647 B.n399 163.367
R1577 B.n647 B.n397 163.367
R1578 B.n651 B.n397 163.367
R1579 B.n651 B.n391 163.367
R1580 B.n660 B.n391 163.367
R1581 B.n660 B.n389 163.367
R1582 B.n664 B.n389 163.367
R1583 B.n664 B.n384 163.367
R1584 B.n672 B.n384 163.367
R1585 B.n672 B.n382 163.367
R1586 B.n676 B.n382 163.367
R1587 B.n676 B.n376 163.367
R1588 B.n684 B.n376 163.367
R1589 B.n684 B.n374 163.367
R1590 B.n688 B.n374 163.367
R1591 B.n688 B.n368 163.367
R1592 B.n696 B.n368 163.367
R1593 B.n696 B.n366 163.367
R1594 B.n700 B.n366 163.367
R1595 B.n700 B.n360 163.367
R1596 B.n708 B.n360 163.367
R1597 B.n708 B.n358 163.367
R1598 B.n712 B.n358 163.367
R1599 B.n712 B.n352 163.367
R1600 B.n720 B.n352 163.367
R1601 B.n720 B.n350 163.367
R1602 B.n724 B.n350 163.367
R1603 B.n724 B.n344 163.367
R1604 B.n732 B.n344 163.367
R1605 B.n732 B.n342 163.367
R1606 B.n736 B.n342 163.367
R1607 B.n736 B.n336 163.367
R1608 B.n744 B.n336 163.367
R1609 B.n744 B.n334 163.367
R1610 B.n748 B.n334 163.367
R1611 B.n748 B.n328 163.367
R1612 B.n756 B.n328 163.367
R1613 B.n756 B.n326 163.367
R1614 B.n760 B.n326 163.367
R1615 B.n760 B.n320 163.367
R1616 B.n768 B.n320 163.367
R1617 B.n768 B.n318 163.367
R1618 B.n772 B.n318 163.367
R1619 B.n772 B.n312 163.367
R1620 B.n780 B.n312 163.367
R1621 B.n780 B.n310 163.367
R1622 B.n784 B.n310 163.367
R1623 B.n784 B.n304 163.367
R1624 B.n793 B.n304 163.367
R1625 B.n793 B.n302 163.367
R1626 B.n797 B.n302 163.367
R1627 B.n797 B.n297 163.367
R1628 B.n806 B.n297 163.367
R1629 B.n806 B.n295 163.367
R1630 B.n810 B.n295 163.367
R1631 B.n810 B.n3 163.367
R1632 B.n1060 B.n3 163.367
R1633 B.n1056 B.n2 163.367
R1634 B.n1056 B.n1055 163.367
R1635 B.n1055 B.n9 163.367
R1636 B.n1051 B.n9 163.367
R1637 B.n1051 B.n11 163.367
R1638 B.n1047 B.n11 163.367
R1639 B.n1047 B.n16 163.367
R1640 B.n1043 B.n16 163.367
R1641 B.n1043 B.n18 163.367
R1642 B.n1039 B.n18 163.367
R1643 B.n1039 B.n24 163.367
R1644 B.n1035 B.n24 163.367
R1645 B.n1035 B.n26 163.367
R1646 B.n1031 B.n26 163.367
R1647 B.n1031 B.n31 163.367
R1648 B.n1027 B.n31 163.367
R1649 B.n1027 B.n33 163.367
R1650 B.n1023 B.n33 163.367
R1651 B.n1023 B.n38 163.367
R1652 B.n1019 B.n38 163.367
R1653 B.n1019 B.n40 163.367
R1654 B.n1015 B.n40 163.367
R1655 B.n1015 B.n45 163.367
R1656 B.n1011 B.n45 163.367
R1657 B.n1011 B.n47 163.367
R1658 B.n1007 B.n47 163.367
R1659 B.n1007 B.n52 163.367
R1660 B.n1003 B.n52 163.367
R1661 B.n1003 B.n54 163.367
R1662 B.n999 B.n54 163.367
R1663 B.n999 B.n59 163.367
R1664 B.n995 B.n59 163.367
R1665 B.n995 B.n61 163.367
R1666 B.n991 B.n61 163.367
R1667 B.n991 B.n66 163.367
R1668 B.n987 B.n66 163.367
R1669 B.n987 B.n68 163.367
R1670 B.n983 B.n68 163.367
R1671 B.n983 B.n73 163.367
R1672 B.n979 B.n73 163.367
R1673 B.n979 B.n75 163.367
R1674 B.n975 B.n75 163.367
R1675 B.n975 B.n80 163.367
R1676 B.n971 B.n80 163.367
R1677 B.n971 B.n82 163.367
R1678 B.n967 B.n82 163.367
R1679 B.n967 B.n87 163.367
R1680 B.n963 B.n87 163.367
R1681 B.n963 B.n89 163.367
R1682 B.n959 B.n89 163.367
R1683 B.n959 B.n93 163.367
R1684 B.n955 B.n93 163.367
R1685 B.n955 B.n95 163.367
R1686 B.n951 B.n95 163.367
R1687 B.n951 B.n101 163.367
R1688 B.n947 B.n101 163.367
R1689 B.n947 B.n103 163.367
R1690 B.n943 B.n103 163.367
R1691 B.n943 B.n108 163.367
R1692 B.n939 B.n108 163.367
R1693 B.n939 B.n110 163.367
R1694 B.n935 B.n110 163.367
R1695 B.n935 B.n115 163.367
R1696 B.n931 B.n115 163.367
R1697 B.n931 B.n117 163.367
R1698 B.n927 B.n117 163.367
R1699 B.n927 B.n122 163.367
R1700 B.n923 B.n122 163.367
R1701 B.n923 B.n124 163.367
R1702 B.n919 B.n124 163.367
R1703 B.n919 B.n129 163.367
R1704 B.n915 B.n129 163.367
R1705 B.n915 B.n131 163.367
R1706 B.n592 B.n432 107.206
R1707 B.n913 B.n912 107.206
R1708 B.n169 B.n168 71.7581
R1709 B.n166 B.n165 71.7581
R1710 B.n470 B.n469 71.7581
R1711 B.n468 B.n467 71.7581
R1712 B.n171 B.n134 71.676
R1713 B.n175 B.n135 71.676
R1714 B.n179 B.n136 71.676
R1715 B.n183 B.n137 71.676
R1716 B.n187 B.n138 71.676
R1717 B.n191 B.n139 71.676
R1718 B.n195 B.n140 71.676
R1719 B.n199 B.n141 71.676
R1720 B.n203 B.n142 71.676
R1721 B.n207 B.n143 71.676
R1722 B.n211 B.n144 71.676
R1723 B.n215 B.n145 71.676
R1724 B.n219 B.n146 71.676
R1725 B.n223 B.n147 71.676
R1726 B.n227 B.n148 71.676
R1727 B.n231 B.n149 71.676
R1728 B.n235 B.n150 71.676
R1729 B.n239 B.n151 71.676
R1730 B.n243 B.n152 71.676
R1731 B.n247 B.n153 71.676
R1732 B.n251 B.n154 71.676
R1733 B.n255 B.n155 71.676
R1734 B.n259 B.n156 71.676
R1735 B.n263 B.n157 71.676
R1736 B.n267 B.n158 71.676
R1737 B.n271 B.n159 71.676
R1738 B.n275 B.n160 71.676
R1739 B.n279 B.n161 71.676
R1740 B.n283 B.n162 71.676
R1741 B.n287 B.n163 71.676
R1742 B.n911 B.n164 71.676
R1743 B.n911 B.n910 71.676
R1744 B.n289 B.n163 71.676
R1745 B.n286 B.n162 71.676
R1746 B.n282 B.n161 71.676
R1747 B.n278 B.n160 71.676
R1748 B.n274 B.n159 71.676
R1749 B.n270 B.n158 71.676
R1750 B.n266 B.n157 71.676
R1751 B.n262 B.n156 71.676
R1752 B.n258 B.n155 71.676
R1753 B.n254 B.n154 71.676
R1754 B.n250 B.n153 71.676
R1755 B.n246 B.n152 71.676
R1756 B.n242 B.n151 71.676
R1757 B.n238 B.n150 71.676
R1758 B.n234 B.n149 71.676
R1759 B.n230 B.n148 71.676
R1760 B.n226 B.n147 71.676
R1761 B.n222 B.n146 71.676
R1762 B.n218 B.n145 71.676
R1763 B.n214 B.n144 71.676
R1764 B.n210 B.n143 71.676
R1765 B.n206 B.n142 71.676
R1766 B.n202 B.n141 71.676
R1767 B.n198 B.n140 71.676
R1768 B.n194 B.n139 71.676
R1769 B.n190 B.n138 71.676
R1770 B.n186 B.n137 71.676
R1771 B.n182 B.n136 71.676
R1772 B.n178 B.n135 71.676
R1773 B.n174 B.n134 71.676
R1774 B.n591 B.n590 71.676
R1775 B.n585 B.n436 71.676
R1776 B.n582 B.n437 71.676
R1777 B.n578 B.n438 71.676
R1778 B.n574 B.n439 71.676
R1779 B.n570 B.n440 71.676
R1780 B.n566 B.n441 71.676
R1781 B.n562 B.n442 71.676
R1782 B.n558 B.n443 71.676
R1783 B.n554 B.n444 71.676
R1784 B.n550 B.n445 71.676
R1785 B.n546 B.n446 71.676
R1786 B.n542 B.n447 71.676
R1787 B.n537 B.n448 71.676
R1788 B.n533 B.n449 71.676
R1789 B.n529 B.n450 71.676
R1790 B.n525 B.n451 71.676
R1791 B.n521 B.n452 71.676
R1792 B.n516 B.n453 71.676
R1793 B.n512 B.n454 71.676
R1794 B.n508 B.n455 71.676
R1795 B.n504 B.n456 71.676
R1796 B.n500 B.n457 71.676
R1797 B.n496 B.n458 71.676
R1798 B.n492 B.n459 71.676
R1799 B.n488 B.n460 71.676
R1800 B.n484 B.n461 71.676
R1801 B.n480 B.n462 71.676
R1802 B.n476 B.n463 71.676
R1803 B.n472 B.n464 71.676
R1804 B.n591 B.n466 71.676
R1805 B.n583 B.n436 71.676
R1806 B.n579 B.n437 71.676
R1807 B.n575 B.n438 71.676
R1808 B.n571 B.n439 71.676
R1809 B.n567 B.n440 71.676
R1810 B.n563 B.n441 71.676
R1811 B.n559 B.n442 71.676
R1812 B.n555 B.n443 71.676
R1813 B.n551 B.n444 71.676
R1814 B.n547 B.n445 71.676
R1815 B.n543 B.n446 71.676
R1816 B.n538 B.n447 71.676
R1817 B.n534 B.n448 71.676
R1818 B.n530 B.n449 71.676
R1819 B.n526 B.n450 71.676
R1820 B.n522 B.n451 71.676
R1821 B.n517 B.n452 71.676
R1822 B.n513 B.n453 71.676
R1823 B.n509 B.n454 71.676
R1824 B.n505 B.n455 71.676
R1825 B.n501 B.n456 71.676
R1826 B.n497 B.n457 71.676
R1827 B.n493 B.n458 71.676
R1828 B.n489 B.n459 71.676
R1829 B.n485 B.n460 71.676
R1830 B.n481 B.n461 71.676
R1831 B.n477 B.n462 71.676
R1832 B.n473 B.n463 71.676
R1833 B.n464 B.n435 71.676
R1834 B.n1061 B.n1060 71.676
R1835 B.n1061 B.n2 71.676
R1836 B.n598 B.n432 62.3079
R1837 B.n598 B.n428 62.3079
R1838 B.n604 B.n428 62.3079
R1839 B.n604 B.n424 62.3079
R1840 B.n610 B.n424 62.3079
R1841 B.n610 B.n419 62.3079
R1842 B.n616 B.n419 62.3079
R1843 B.n616 B.n420 62.3079
R1844 B.n622 B.n412 62.3079
R1845 B.n628 B.n412 62.3079
R1846 B.n628 B.n408 62.3079
R1847 B.n634 B.n408 62.3079
R1848 B.n634 B.n404 62.3079
R1849 B.n640 B.n404 62.3079
R1850 B.n640 B.n400 62.3079
R1851 B.n646 B.n400 62.3079
R1852 B.n646 B.n396 62.3079
R1853 B.n652 B.n396 62.3079
R1854 B.n652 B.n392 62.3079
R1855 B.n659 B.n392 62.3079
R1856 B.n659 B.n658 62.3079
R1857 B.n665 B.n385 62.3079
R1858 B.n671 B.n385 62.3079
R1859 B.n671 B.n381 62.3079
R1860 B.n677 B.n381 62.3079
R1861 B.n677 B.n377 62.3079
R1862 B.n683 B.n377 62.3079
R1863 B.n683 B.n373 62.3079
R1864 B.n689 B.n373 62.3079
R1865 B.n689 B.n369 62.3079
R1866 B.n695 B.n369 62.3079
R1867 B.n701 B.n365 62.3079
R1868 B.n701 B.n361 62.3079
R1869 B.n707 B.n361 62.3079
R1870 B.n707 B.n357 62.3079
R1871 B.n713 B.n357 62.3079
R1872 B.n713 B.n353 62.3079
R1873 B.n719 B.n353 62.3079
R1874 B.n719 B.n348 62.3079
R1875 B.n725 B.n348 62.3079
R1876 B.n725 B.n349 62.3079
R1877 B.n731 B.n341 62.3079
R1878 B.n737 B.n341 62.3079
R1879 B.n737 B.n337 62.3079
R1880 B.n743 B.n337 62.3079
R1881 B.n743 B.n333 62.3079
R1882 B.n749 B.n333 62.3079
R1883 B.n749 B.n329 62.3079
R1884 B.n755 B.n329 62.3079
R1885 B.n755 B.n325 62.3079
R1886 B.n761 B.n325 62.3079
R1887 B.n767 B.n321 62.3079
R1888 B.n767 B.n317 62.3079
R1889 B.n773 B.n317 62.3079
R1890 B.n773 B.n313 62.3079
R1891 B.n779 B.n313 62.3079
R1892 B.n779 B.n309 62.3079
R1893 B.n785 B.n309 62.3079
R1894 B.n785 B.n305 62.3079
R1895 B.n792 B.n305 62.3079
R1896 B.n792 B.n791 62.3079
R1897 B.n798 B.n298 62.3079
R1898 B.n805 B.n298 62.3079
R1899 B.n805 B.n294 62.3079
R1900 B.n811 B.n294 62.3079
R1901 B.n811 B.n4 62.3079
R1902 B.n1059 B.n4 62.3079
R1903 B.n1059 B.n1058 62.3079
R1904 B.n1058 B.n1057 62.3079
R1905 B.n1057 B.n8 62.3079
R1906 B.n12 B.n8 62.3079
R1907 B.n1050 B.n12 62.3079
R1908 B.n1050 B.n1049 62.3079
R1909 B.n1049 B.n1048 62.3079
R1910 B.n1042 B.n19 62.3079
R1911 B.n1042 B.n1041 62.3079
R1912 B.n1041 B.n1040 62.3079
R1913 B.n1040 B.n23 62.3079
R1914 B.n1034 B.n23 62.3079
R1915 B.n1034 B.n1033 62.3079
R1916 B.n1033 B.n1032 62.3079
R1917 B.n1032 B.n30 62.3079
R1918 B.n1026 B.n30 62.3079
R1919 B.n1026 B.n1025 62.3079
R1920 B.n1024 B.n37 62.3079
R1921 B.n1018 B.n37 62.3079
R1922 B.n1018 B.n1017 62.3079
R1923 B.n1017 B.n1016 62.3079
R1924 B.n1016 B.n44 62.3079
R1925 B.n1010 B.n44 62.3079
R1926 B.n1010 B.n1009 62.3079
R1927 B.n1009 B.n1008 62.3079
R1928 B.n1008 B.n51 62.3079
R1929 B.n1002 B.n51 62.3079
R1930 B.n1001 B.n1000 62.3079
R1931 B.n1000 B.n58 62.3079
R1932 B.n994 B.n58 62.3079
R1933 B.n994 B.n993 62.3079
R1934 B.n993 B.n992 62.3079
R1935 B.n992 B.n65 62.3079
R1936 B.n986 B.n65 62.3079
R1937 B.n986 B.n985 62.3079
R1938 B.n985 B.n984 62.3079
R1939 B.n984 B.n72 62.3079
R1940 B.n978 B.n977 62.3079
R1941 B.n977 B.n976 62.3079
R1942 B.n976 B.n79 62.3079
R1943 B.n970 B.n79 62.3079
R1944 B.n970 B.n969 62.3079
R1945 B.n969 B.n968 62.3079
R1946 B.n968 B.n86 62.3079
R1947 B.n962 B.n86 62.3079
R1948 B.n962 B.n961 62.3079
R1949 B.n961 B.n960 62.3079
R1950 B.n954 B.n96 62.3079
R1951 B.n954 B.n953 62.3079
R1952 B.n953 B.n952 62.3079
R1953 B.n952 B.n100 62.3079
R1954 B.n946 B.n100 62.3079
R1955 B.n946 B.n945 62.3079
R1956 B.n945 B.n944 62.3079
R1957 B.n944 B.n107 62.3079
R1958 B.n938 B.n107 62.3079
R1959 B.n938 B.n937 62.3079
R1960 B.n937 B.n936 62.3079
R1961 B.n936 B.n114 62.3079
R1962 B.n930 B.n114 62.3079
R1963 B.n929 B.n928 62.3079
R1964 B.n928 B.n121 62.3079
R1965 B.n922 B.n121 62.3079
R1966 B.n922 B.n921 62.3079
R1967 B.n921 B.n920 62.3079
R1968 B.n920 B.n128 62.3079
R1969 B.n914 B.n128 62.3079
R1970 B.n914 B.n913 62.3079
R1971 B.n170 B.n169 59.5399
R1972 B.n167 B.n166 59.5399
R1973 B.n519 B.n470 59.5399
R1974 B.n540 B.n468 59.5399
R1975 B.n658 B.t2 57.7264
R1976 B.n96 B.t5 57.7264
R1977 B.n420 B.t18 52.2287
R1978 B.t11 B.n929 52.2287
R1979 B.n695 B.t4 50.3962
R1980 B.n978 B.t8 50.3962
R1981 B.n349 B.t1 43.0659
R1982 B.t0 B.n1001 43.0659
R1983 B.n761 B.t3 35.7356
R1984 B.t7 B.n1024 35.7356
R1985 B.n798 B.t9 33.903
R1986 B.n1048 B.t6 33.903
R1987 B.n589 B.n430 30.4395
R1988 B.n595 B.n594 30.4395
R1989 B.n909 B.n908 30.4395
R1990 B.n172 B.n130 30.4395
R1991 B.n791 B.t9 28.4053
R1992 B.n19 B.t6 28.4053
R1993 B.t3 B.n321 26.5728
R1994 B.n1025 B.t7 26.5728
R1995 B.n731 B.t1 19.2425
R1996 B.n1002 B.t0 19.2425
R1997 B B.n1062 18.0485
R1998 B.t4 B.n365 11.9122
R1999 B.t8 B.n72 11.9122
R2000 B.n600 B.n430 10.6151
R2001 B.n601 B.n600 10.6151
R2002 B.n602 B.n601 10.6151
R2003 B.n602 B.n422 10.6151
R2004 B.n612 B.n422 10.6151
R2005 B.n613 B.n612 10.6151
R2006 B.n614 B.n613 10.6151
R2007 B.n614 B.n414 10.6151
R2008 B.n624 B.n414 10.6151
R2009 B.n625 B.n624 10.6151
R2010 B.n626 B.n625 10.6151
R2011 B.n626 B.n406 10.6151
R2012 B.n636 B.n406 10.6151
R2013 B.n637 B.n636 10.6151
R2014 B.n638 B.n637 10.6151
R2015 B.n638 B.n398 10.6151
R2016 B.n648 B.n398 10.6151
R2017 B.n649 B.n648 10.6151
R2018 B.n650 B.n649 10.6151
R2019 B.n650 B.n390 10.6151
R2020 B.n661 B.n390 10.6151
R2021 B.n662 B.n661 10.6151
R2022 B.n663 B.n662 10.6151
R2023 B.n663 B.n383 10.6151
R2024 B.n673 B.n383 10.6151
R2025 B.n674 B.n673 10.6151
R2026 B.n675 B.n674 10.6151
R2027 B.n675 B.n375 10.6151
R2028 B.n685 B.n375 10.6151
R2029 B.n686 B.n685 10.6151
R2030 B.n687 B.n686 10.6151
R2031 B.n687 B.n367 10.6151
R2032 B.n697 B.n367 10.6151
R2033 B.n698 B.n697 10.6151
R2034 B.n699 B.n698 10.6151
R2035 B.n699 B.n359 10.6151
R2036 B.n709 B.n359 10.6151
R2037 B.n710 B.n709 10.6151
R2038 B.n711 B.n710 10.6151
R2039 B.n711 B.n351 10.6151
R2040 B.n721 B.n351 10.6151
R2041 B.n722 B.n721 10.6151
R2042 B.n723 B.n722 10.6151
R2043 B.n723 B.n343 10.6151
R2044 B.n733 B.n343 10.6151
R2045 B.n734 B.n733 10.6151
R2046 B.n735 B.n734 10.6151
R2047 B.n735 B.n335 10.6151
R2048 B.n745 B.n335 10.6151
R2049 B.n746 B.n745 10.6151
R2050 B.n747 B.n746 10.6151
R2051 B.n747 B.n327 10.6151
R2052 B.n757 B.n327 10.6151
R2053 B.n758 B.n757 10.6151
R2054 B.n759 B.n758 10.6151
R2055 B.n759 B.n319 10.6151
R2056 B.n769 B.n319 10.6151
R2057 B.n770 B.n769 10.6151
R2058 B.n771 B.n770 10.6151
R2059 B.n771 B.n311 10.6151
R2060 B.n781 B.n311 10.6151
R2061 B.n782 B.n781 10.6151
R2062 B.n783 B.n782 10.6151
R2063 B.n783 B.n303 10.6151
R2064 B.n794 B.n303 10.6151
R2065 B.n795 B.n794 10.6151
R2066 B.n796 B.n795 10.6151
R2067 B.n796 B.n296 10.6151
R2068 B.n807 B.n296 10.6151
R2069 B.n808 B.n807 10.6151
R2070 B.n809 B.n808 10.6151
R2071 B.n809 B.n0 10.6151
R2072 B.n589 B.n588 10.6151
R2073 B.n588 B.n587 10.6151
R2074 B.n587 B.n586 10.6151
R2075 B.n586 B.n584 10.6151
R2076 B.n584 B.n581 10.6151
R2077 B.n581 B.n580 10.6151
R2078 B.n580 B.n577 10.6151
R2079 B.n577 B.n576 10.6151
R2080 B.n576 B.n573 10.6151
R2081 B.n573 B.n572 10.6151
R2082 B.n572 B.n569 10.6151
R2083 B.n569 B.n568 10.6151
R2084 B.n568 B.n565 10.6151
R2085 B.n565 B.n564 10.6151
R2086 B.n564 B.n561 10.6151
R2087 B.n561 B.n560 10.6151
R2088 B.n560 B.n557 10.6151
R2089 B.n557 B.n556 10.6151
R2090 B.n556 B.n553 10.6151
R2091 B.n553 B.n552 10.6151
R2092 B.n552 B.n549 10.6151
R2093 B.n549 B.n548 10.6151
R2094 B.n548 B.n545 10.6151
R2095 B.n545 B.n544 10.6151
R2096 B.n544 B.n541 10.6151
R2097 B.n539 B.n536 10.6151
R2098 B.n536 B.n535 10.6151
R2099 B.n535 B.n532 10.6151
R2100 B.n532 B.n531 10.6151
R2101 B.n531 B.n528 10.6151
R2102 B.n528 B.n527 10.6151
R2103 B.n527 B.n524 10.6151
R2104 B.n524 B.n523 10.6151
R2105 B.n523 B.n520 10.6151
R2106 B.n518 B.n515 10.6151
R2107 B.n515 B.n514 10.6151
R2108 B.n514 B.n511 10.6151
R2109 B.n511 B.n510 10.6151
R2110 B.n510 B.n507 10.6151
R2111 B.n507 B.n506 10.6151
R2112 B.n506 B.n503 10.6151
R2113 B.n503 B.n502 10.6151
R2114 B.n502 B.n499 10.6151
R2115 B.n499 B.n498 10.6151
R2116 B.n498 B.n495 10.6151
R2117 B.n495 B.n494 10.6151
R2118 B.n494 B.n491 10.6151
R2119 B.n491 B.n490 10.6151
R2120 B.n490 B.n487 10.6151
R2121 B.n487 B.n486 10.6151
R2122 B.n486 B.n483 10.6151
R2123 B.n483 B.n482 10.6151
R2124 B.n482 B.n479 10.6151
R2125 B.n479 B.n478 10.6151
R2126 B.n478 B.n475 10.6151
R2127 B.n475 B.n474 10.6151
R2128 B.n474 B.n471 10.6151
R2129 B.n471 B.n434 10.6151
R2130 B.n594 B.n434 10.6151
R2131 B.n596 B.n595 10.6151
R2132 B.n596 B.n426 10.6151
R2133 B.n606 B.n426 10.6151
R2134 B.n607 B.n606 10.6151
R2135 B.n608 B.n607 10.6151
R2136 B.n608 B.n417 10.6151
R2137 B.n618 B.n417 10.6151
R2138 B.n619 B.n618 10.6151
R2139 B.n620 B.n619 10.6151
R2140 B.n620 B.n410 10.6151
R2141 B.n630 B.n410 10.6151
R2142 B.n631 B.n630 10.6151
R2143 B.n632 B.n631 10.6151
R2144 B.n632 B.n402 10.6151
R2145 B.n642 B.n402 10.6151
R2146 B.n643 B.n642 10.6151
R2147 B.n644 B.n643 10.6151
R2148 B.n644 B.n394 10.6151
R2149 B.n654 B.n394 10.6151
R2150 B.n655 B.n654 10.6151
R2151 B.n656 B.n655 10.6151
R2152 B.n656 B.n387 10.6151
R2153 B.n667 B.n387 10.6151
R2154 B.n668 B.n667 10.6151
R2155 B.n669 B.n668 10.6151
R2156 B.n669 B.n379 10.6151
R2157 B.n679 B.n379 10.6151
R2158 B.n680 B.n679 10.6151
R2159 B.n681 B.n680 10.6151
R2160 B.n681 B.n371 10.6151
R2161 B.n691 B.n371 10.6151
R2162 B.n692 B.n691 10.6151
R2163 B.n693 B.n692 10.6151
R2164 B.n693 B.n363 10.6151
R2165 B.n703 B.n363 10.6151
R2166 B.n704 B.n703 10.6151
R2167 B.n705 B.n704 10.6151
R2168 B.n705 B.n355 10.6151
R2169 B.n715 B.n355 10.6151
R2170 B.n716 B.n715 10.6151
R2171 B.n717 B.n716 10.6151
R2172 B.n717 B.n346 10.6151
R2173 B.n727 B.n346 10.6151
R2174 B.n728 B.n727 10.6151
R2175 B.n729 B.n728 10.6151
R2176 B.n729 B.n339 10.6151
R2177 B.n739 B.n339 10.6151
R2178 B.n740 B.n739 10.6151
R2179 B.n741 B.n740 10.6151
R2180 B.n741 B.n331 10.6151
R2181 B.n751 B.n331 10.6151
R2182 B.n752 B.n751 10.6151
R2183 B.n753 B.n752 10.6151
R2184 B.n753 B.n323 10.6151
R2185 B.n763 B.n323 10.6151
R2186 B.n764 B.n763 10.6151
R2187 B.n765 B.n764 10.6151
R2188 B.n765 B.n315 10.6151
R2189 B.n775 B.n315 10.6151
R2190 B.n776 B.n775 10.6151
R2191 B.n777 B.n776 10.6151
R2192 B.n777 B.n307 10.6151
R2193 B.n787 B.n307 10.6151
R2194 B.n788 B.n787 10.6151
R2195 B.n789 B.n788 10.6151
R2196 B.n789 B.n300 10.6151
R2197 B.n800 B.n300 10.6151
R2198 B.n801 B.n800 10.6151
R2199 B.n803 B.n801 10.6151
R2200 B.n803 B.n802 10.6151
R2201 B.n802 B.n292 10.6151
R2202 B.n814 B.n292 10.6151
R2203 B.n815 B.n814 10.6151
R2204 B.n816 B.n815 10.6151
R2205 B.n817 B.n816 10.6151
R2206 B.n818 B.n817 10.6151
R2207 B.n821 B.n818 10.6151
R2208 B.n822 B.n821 10.6151
R2209 B.n823 B.n822 10.6151
R2210 B.n824 B.n823 10.6151
R2211 B.n826 B.n824 10.6151
R2212 B.n827 B.n826 10.6151
R2213 B.n828 B.n827 10.6151
R2214 B.n829 B.n828 10.6151
R2215 B.n831 B.n829 10.6151
R2216 B.n832 B.n831 10.6151
R2217 B.n833 B.n832 10.6151
R2218 B.n834 B.n833 10.6151
R2219 B.n836 B.n834 10.6151
R2220 B.n837 B.n836 10.6151
R2221 B.n838 B.n837 10.6151
R2222 B.n839 B.n838 10.6151
R2223 B.n841 B.n839 10.6151
R2224 B.n842 B.n841 10.6151
R2225 B.n843 B.n842 10.6151
R2226 B.n844 B.n843 10.6151
R2227 B.n846 B.n844 10.6151
R2228 B.n847 B.n846 10.6151
R2229 B.n848 B.n847 10.6151
R2230 B.n849 B.n848 10.6151
R2231 B.n851 B.n849 10.6151
R2232 B.n852 B.n851 10.6151
R2233 B.n853 B.n852 10.6151
R2234 B.n854 B.n853 10.6151
R2235 B.n856 B.n854 10.6151
R2236 B.n857 B.n856 10.6151
R2237 B.n858 B.n857 10.6151
R2238 B.n859 B.n858 10.6151
R2239 B.n861 B.n859 10.6151
R2240 B.n862 B.n861 10.6151
R2241 B.n863 B.n862 10.6151
R2242 B.n864 B.n863 10.6151
R2243 B.n866 B.n864 10.6151
R2244 B.n867 B.n866 10.6151
R2245 B.n868 B.n867 10.6151
R2246 B.n869 B.n868 10.6151
R2247 B.n871 B.n869 10.6151
R2248 B.n872 B.n871 10.6151
R2249 B.n873 B.n872 10.6151
R2250 B.n874 B.n873 10.6151
R2251 B.n876 B.n874 10.6151
R2252 B.n877 B.n876 10.6151
R2253 B.n878 B.n877 10.6151
R2254 B.n879 B.n878 10.6151
R2255 B.n881 B.n879 10.6151
R2256 B.n882 B.n881 10.6151
R2257 B.n883 B.n882 10.6151
R2258 B.n884 B.n883 10.6151
R2259 B.n886 B.n884 10.6151
R2260 B.n887 B.n886 10.6151
R2261 B.n888 B.n887 10.6151
R2262 B.n889 B.n888 10.6151
R2263 B.n891 B.n889 10.6151
R2264 B.n892 B.n891 10.6151
R2265 B.n893 B.n892 10.6151
R2266 B.n894 B.n893 10.6151
R2267 B.n896 B.n894 10.6151
R2268 B.n897 B.n896 10.6151
R2269 B.n898 B.n897 10.6151
R2270 B.n899 B.n898 10.6151
R2271 B.n901 B.n899 10.6151
R2272 B.n902 B.n901 10.6151
R2273 B.n903 B.n902 10.6151
R2274 B.n904 B.n903 10.6151
R2275 B.n906 B.n904 10.6151
R2276 B.n907 B.n906 10.6151
R2277 B.n908 B.n907 10.6151
R2278 B.n1054 B.n1 10.6151
R2279 B.n1054 B.n1053 10.6151
R2280 B.n1053 B.n1052 10.6151
R2281 B.n1052 B.n10 10.6151
R2282 B.n1046 B.n10 10.6151
R2283 B.n1046 B.n1045 10.6151
R2284 B.n1045 B.n1044 10.6151
R2285 B.n1044 B.n17 10.6151
R2286 B.n1038 B.n17 10.6151
R2287 B.n1038 B.n1037 10.6151
R2288 B.n1037 B.n1036 10.6151
R2289 B.n1036 B.n25 10.6151
R2290 B.n1030 B.n25 10.6151
R2291 B.n1030 B.n1029 10.6151
R2292 B.n1029 B.n1028 10.6151
R2293 B.n1028 B.n32 10.6151
R2294 B.n1022 B.n32 10.6151
R2295 B.n1022 B.n1021 10.6151
R2296 B.n1021 B.n1020 10.6151
R2297 B.n1020 B.n39 10.6151
R2298 B.n1014 B.n39 10.6151
R2299 B.n1014 B.n1013 10.6151
R2300 B.n1013 B.n1012 10.6151
R2301 B.n1012 B.n46 10.6151
R2302 B.n1006 B.n46 10.6151
R2303 B.n1006 B.n1005 10.6151
R2304 B.n1005 B.n1004 10.6151
R2305 B.n1004 B.n53 10.6151
R2306 B.n998 B.n53 10.6151
R2307 B.n998 B.n997 10.6151
R2308 B.n997 B.n996 10.6151
R2309 B.n996 B.n60 10.6151
R2310 B.n990 B.n60 10.6151
R2311 B.n990 B.n989 10.6151
R2312 B.n989 B.n988 10.6151
R2313 B.n988 B.n67 10.6151
R2314 B.n982 B.n67 10.6151
R2315 B.n982 B.n981 10.6151
R2316 B.n981 B.n980 10.6151
R2317 B.n980 B.n74 10.6151
R2318 B.n974 B.n74 10.6151
R2319 B.n974 B.n973 10.6151
R2320 B.n973 B.n972 10.6151
R2321 B.n972 B.n81 10.6151
R2322 B.n966 B.n81 10.6151
R2323 B.n966 B.n965 10.6151
R2324 B.n965 B.n964 10.6151
R2325 B.n964 B.n88 10.6151
R2326 B.n958 B.n88 10.6151
R2327 B.n958 B.n957 10.6151
R2328 B.n957 B.n956 10.6151
R2329 B.n956 B.n94 10.6151
R2330 B.n950 B.n94 10.6151
R2331 B.n950 B.n949 10.6151
R2332 B.n949 B.n948 10.6151
R2333 B.n948 B.n102 10.6151
R2334 B.n942 B.n102 10.6151
R2335 B.n942 B.n941 10.6151
R2336 B.n941 B.n940 10.6151
R2337 B.n940 B.n109 10.6151
R2338 B.n934 B.n109 10.6151
R2339 B.n934 B.n933 10.6151
R2340 B.n933 B.n932 10.6151
R2341 B.n932 B.n116 10.6151
R2342 B.n926 B.n116 10.6151
R2343 B.n926 B.n925 10.6151
R2344 B.n925 B.n924 10.6151
R2345 B.n924 B.n123 10.6151
R2346 B.n918 B.n123 10.6151
R2347 B.n918 B.n917 10.6151
R2348 B.n917 B.n916 10.6151
R2349 B.n916 B.n130 10.6151
R2350 B.n173 B.n172 10.6151
R2351 B.n176 B.n173 10.6151
R2352 B.n177 B.n176 10.6151
R2353 B.n180 B.n177 10.6151
R2354 B.n181 B.n180 10.6151
R2355 B.n184 B.n181 10.6151
R2356 B.n185 B.n184 10.6151
R2357 B.n188 B.n185 10.6151
R2358 B.n189 B.n188 10.6151
R2359 B.n192 B.n189 10.6151
R2360 B.n193 B.n192 10.6151
R2361 B.n196 B.n193 10.6151
R2362 B.n197 B.n196 10.6151
R2363 B.n200 B.n197 10.6151
R2364 B.n201 B.n200 10.6151
R2365 B.n204 B.n201 10.6151
R2366 B.n205 B.n204 10.6151
R2367 B.n208 B.n205 10.6151
R2368 B.n209 B.n208 10.6151
R2369 B.n212 B.n209 10.6151
R2370 B.n213 B.n212 10.6151
R2371 B.n216 B.n213 10.6151
R2372 B.n217 B.n216 10.6151
R2373 B.n220 B.n217 10.6151
R2374 B.n221 B.n220 10.6151
R2375 B.n225 B.n224 10.6151
R2376 B.n228 B.n225 10.6151
R2377 B.n229 B.n228 10.6151
R2378 B.n232 B.n229 10.6151
R2379 B.n233 B.n232 10.6151
R2380 B.n236 B.n233 10.6151
R2381 B.n237 B.n236 10.6151
R2382 B.n240 B.n237 10.6151
R2383 B.n241 B.n240 10.6151
R2384 B.n245 B.n244 10.6151
R2385 B.n248 B.n245 10.6151
R2386 B.n249 B.n248 10.6151
R2387 B.n252 B.n249 10.6151
R2388 B.n253 B.n252 10.6151
R2389 B.n256 B.n253 10.6151
R2390 B.n257 B.n256 10.6151
R2391 B.n260 B.n257 10.6151
R2392 B.n261 B.n260 10.6151
R2393 B.n264 B.n261 10.6151
R2394 B.n265 B.n264 10.6151
R2395 B.n268 B.n265 10.6151
R2396 B.n269 B.n268 10.6151
R2397 B.n272 B.n269 10.6151
R2398 B.n273 B.n272 10.6151
R2399 B.n276 B.n273 10.6151
R2400 B.n277 B.n276 10.6151
R2401 B.n280 B.n277 10.6151
R2402 B.n281 B.n280 10.6151
R2403 B.n284 B.n281 10.6151
R2404 B.n285 B.n284 10.6151
R2405 B.n288 B.n285 10.6151
R2406 B.n290 B.n288 10.6151
R2407 B.n291 B.n290 10.6151
R2408 B.n909 B.n291 10.6151
R2409 B.n622 B.t18 10.0796
R2410 B.n930 B.t11 10.0796
R2411 B.n541 B.n540 9.36635
R2412 B.n519 B.n518 9.36635
R2413 B.n221 B.n170 9.36635
R2414 B.n244 B.n167 9.36635
R2415 B.n1062 B.n0 8.11757
R2416 B.n1062 B.n1 8.11757
R2417 B.n665 B.t2 4.58192
R2418 B.n960 B.t5 4.58192
R2419 B.n540 B.n539 1.24928
R2420 B.n520 B.n519 1.24928
R2421 B.n224 B.n170 1.24928
R2422 B.n241 B.n167 1.24928
R2423 VN.n98 VN.n97 161.3
R2424 VN.n96 VN.n51 161.3
R2425 VN.n95 VN.n94 161.3
R2426 VN.n93 VN.n52 161.3
R2427 VN.n92 VN.n91 161.3
R2428 VN.n90 VN.n53 161.3
R2429 VN.n89 VN.n88 161.3
R2430 VN.n87 VN.n54 161.3
R2431 VN.n86 VN.n85 161.3
R2432 VN.n84 VN.n55 161.3
R2433 VN.n83 VN.n82 161.3
R2434 VN.n81 VN.n57 161.3
R2435 VN.n80 VN.n79 161.3
R2436 VN.n78 VN.n58 161.3
R2437 VN.n77 VN.n76 161.3
R2438 VN.n75 VN.n74 161.3
R2439 VN.n73 VN.n60 161.3
R2440 VN.n72 VN.n71 161.3
R2441 VN.n70 VN.n61 161.3
R2442 VN.n69 VN.n68 161.3
R2443 VN.n67 VN.n62 161.3
R2444 VN.n66 VN.n65 161.3
R2445 VN.n48 VN.n47 161.3
R2446 VN.n46 VN.n1 161.3
R2447 VN.n45 VN.n44 161.3
R2448 VN.n43 VN.n2 161.3
R2449 VN.n42 VN.n41 161.3
R2450 VN.n40 VN.n3 161.3
R2451 VN.n39 VN.n38 161.3
R2452 VN.n37 VN.n4 161.3
R2453 VN.n36 VN.n35 161.3
R2454 VN.n33 VN.n5 161.3
R2455 VN.n32 VN.n31 161.3
R2456 VN.n30 VN.n6 161.3
R2457 VN.n29 VN.n28 161.3
R2458 VN.n27 VN.n7 161.3
R2459 VN.n26 VN.n25 161.3
R2460 VN.n24 VN.n23 161.3
R2461 VN.n22 VN.n9 161.3
R2462 VN.n21 VN.n20 161.3
R2463 VN.n19 VN.n10 161.3
R2464 VN.n18 VN.n17 161.3
R2465 VN.n16 VN.n11 161.3
R2466 VN.n15 VN.n14 161.3
R2467 VN.n49 VN.n0 82.7273
R2468 VN.n99 VN.n50 82.7273
R2469 VN.n13 VN.t1 81.058
R2470 VN.n64 VN.t5 81.058
R2471 VN.n41 VN.n2 56.5193
R2472 VN.n91 VN.n52 56.5193
R2473 VN VN.n99 53.4904
R2474 VN.n64 VN.n63 52.4975
R2475 VN.n13 VN.n12 52.4975
R2476 VN.n17 VN.n10 50.2061
R2477 VN.n32 VN.n6 50.2061
R2478 VN.n68 VN.n61 50.2061
R2479 VN.n83 VN.n57 50.2061
R2480 VN.n12 VN.t6 48.129
R2481 VN.n8 VN.t9 48.129
R2482 VN.n34 VN.t4 48.129
R2483 VN.n0 VN.t8 48.129
R2484 VN.n63 VN.t3 48.129
R2485 VN.n59 VN.t7 48.129
R2486 VN.n56 VN.t2 48.129
R2487 VN.n50 VN.t0 48.129
R2488 VN.n21 VN.n10 30.7807
R2489 VN.n28 VN.n6 30.7807
R2490 VN.n72 VN.n61 30.7807
R2491 VN.n79 VN.n57 30.7807
R2492 VN.n16 VN.n15 24.4675
R2493 VN.n17 VN.n16 24.4675
R2494 VN.n22 VN.n21 24.4675
R2495 VN.n23 VN.n22 24.4675
R2496 VN.n27 VN.n26 24.4675
R2497 VN.n28 VN.n27 24.4675
R2498 VN.n33 VN.n32 24.4675
R2499 VN.n35 VN.n33 24.4675
R2500 VN.n39 VN.n4 24.4675
R2501 VN.n40 VN.n39 24.4675
R2502 VN.n41 VN.n40 24.4675
R2503 VN.n45 VN.n2 24.4675
R2504 VN.n46 VN.n45 24.4675
R2505 VN.n47 VN.n46 24.4675
R2506 VN.n68 VN.n67 24.4675
R2507 VN.n67 VN.n66 24.4675
R2508 VN.n79 VN.n78 24.4675
R2509 VN.n78 VN.n77 24.4675
R2510 VN.n74 VN.n73 24.4675
R2511 VN.n73 VN.n72 24.4675
R2512 VN.n91 VN.n90 24.4675
R2513 VN.n90 VN.n89 24.4675
R2514 VN.n89 VN.n54 24.4675
R2515 VN.n85 VN.n84 24.4675
R2516 VN.n84 VN.n83 24.4675
R2517 VN.n97 VN.n96 24.4675
R2518 VN.n96 VN.n95 24.4675
R2519 VN.n95 VN.n52 24.4675
R2520 VN.n15 VN.n12 22.0208
R2521 VN.n35 VN.n34 22.0208
R2522 VN.n66 VN.n63 22.0208
R2523 VN.n85 VN.n56 22.0208
R2524 VN.n23 VN.n8 12.234
R2525 VN.n26 VN.n8 12.234
R2526 VN.n77 VN.n59 12.234
R2527 VN.n74 VN.n59 12.234
R2528 VN.n47 VN.n0 7.3406
R2529 VN.n97 VN.n50 7.3406
R2530 VN.n65 VN.n64 3.24375
R2531 VN.n14 VN.n13 3.24375
R2532 VN.n34 VN.n4 2.4472
R2533 VN.n56 VN.n54 2.4472
R2534 VN.n99 VN.n98 0.354971
R2535 VN.n49 VN.n48 0.354971
R2536 VN VN.n49 0.26696
R2537 VN.n98 VN.n51 0.189894
R2538 VN.n94 VN.n51 0.189894
R2539 VN.n94 VN.n93 0.189894
R2540 VN.n93 VN.n92 0.189894
R2541 VN.n92 VN.n53 0.189894
R2542 VN.n88 VN.n53 0.189894
R2543 VN.n88 VN.n87 0.189894
R2544 VN.n87 VN.n86 0.189894
R2545 VN.n86 VN.n55 0.189894
R2546 VN.n82 VN.n55 0.189894
R2547 VN.n82 VN.n81 0.189894
R2548 VN.n81 VN.n80 0.189894
R2549 VN.n80 VN.n58 0.189894
R2550 VN.n76 VN.n58 0.189894
R2551 VN.n76 VN.n75 0.189894
R2552 VN.n75 VN.n60 0.189894
R2553 VN.n71 VN.n60 0.189894
R2554 VN.n71 VN.n70 0.189894
R2555 VN.n70 VN.n69 0.189894
R2556 VN.n69 VN.n62 0.189894
R2557 VN.n65 VN.n62 0.189894
R2558 VN.n14 VN.n11 0.189894
R2559 VN.n18 VN.n11 0.189894
R2560 VN.n19 VN.n18 0.189894
R2561 VN.n20 VN.n19 0.189894
R2562 VN.n20 VN.n9 0.189894
R2563 VN.n24 VN.n9 0.189894
R2564 VN.n25 VN.n24 0.189894
R2565 VN.n25 VN.n7 0.189894
R2566 VN.n29 VN.n7 0.189894
R2567 VN.n30 VN.n29 0.189894
R2568 VN.n31 VN.n30 0.189894
R2569 VN.n31 VN.n5 0.189894
R2570 VN.n36 VN.n5 0.189894
R2571 VN.n37 VN.n36 0.189894
R2572 VN.n38 VN.n37 0.189894
R2573 VN.n38 VN.n3 0.189894
R2574 VN.n42 VN.n3 0.189894
R2575 VN.n43 VN.n42 0.189894
R2576 VN.n44 VN.n43 0.189894
R2577 VN.n44 VN.n1 0.189894
R2578 VN.n48 VN.n1 0.189894
R2579 VDD2.n69 VDD2.n39 289.615
R2580 VDD2.n30 VDD2.n0 289.615
R2581 VDD2.n70 VDD2.n69 185
R2582 VDD2.n68 VDD2.n67 185
R2583 VDD2.n43 VDD2.n42 185
R2584 VDD2.n62 VDD2.n61 185
R2585 VDD2.n60 VDD2.n59 185
R2586 VDD2.n47 VDD2.n46 185
R2587 VDD2.n54 VDD2.n53 185
R2588 VDD2.n52 VDD2.n51 185
R2589 VDD2.n13 VDD2.n12 185
R2590 VDD2.n15 VDD2.n14 185
R2591 VDD2.n8 VDD2.n7 185
R2592 VDD2.n21 VDD2.n20 185
R2593 VDD2.n23 VDD2.n22 185
R2594 VDD2.n4 VDD2.n3 185
R2595 VDD2.n29 VDD2.n28 185
R2596 VDD2.n31 VDD2.n30 185
R2597 VDD2.n50 VDD2.t9 147.659
R2598 VDD2.n11 VDD2.t8 147.659
R2599 VDD2.n69 VDD2.n68 104.615
R2600 VDD2.n68 VDD2.n42 104.615
R2601 VDD2.n61 VDD2.n42 104.615
R2602 VDD2.n61 VDD2.n60 104.615
R2603 VDD2.n60 VDD2.n46 104.615
R2604 VDD2.n53 VDD2.n46 104.615
R2605 VDD2.n53 VDD2.n52 104.615
R2606 VDD2.n14 VDD2.n13 104.615
R2607 VDD2.n14 VDD2.n7 104.615
R2608 VDD2.n21 VDD2.n7 104.615
R2609 VDD2.n22 VDD2.n21 104.615
R2610 VDD2.n22 VDD2.n3 104.615
R2611 VDD2.n29 VDD2.n3 104.615
R2612 VDD2.n30 VDD2.n29 104.615
R2613 VDD2.n38 VDD2.n37 68.6048
R2614 VDD2 VDD2.n77 68.6019
R2615 VDD2.n76 VDD2.n75 66.2681
R2616 VDD2.n36 VDD2.n35 66.2679
R2617 VDD2.n52 VDD2.t9 52.3082
R2618 VDD2.n13 VDD2.t8 52.3082
R2619 VDD2.n36 VDD2.n34 52.2477
R2620 VDD2.n74 VDD2.n73 49.0581
R2621 VDD2.n74 VDD2.n38 44.6679
R2622 VDD2.n51 VDD2.n50 15.6676
R2623 VDD2.n12 VDD2.n11 15.6676
R2624 VDD2.n54 VDD2.n49 12.8005
R2625 VDD2.n15 VDD2.n10 12.8005
R2626 VDD2.n55 VDD2.n47 12.0247
R2627 VDD2.n16 VDD2.n8 12.0247
R2628 VDD2.n59 VDD2.n58 11.249
R2629 VDD2.n20 VDD2.n19 11.249
R2630 VDD2.n62 VDD2.n45 10.4732
R2631 VDD2.n23 VDD2.n6 10.4732
R2632 VDD2.n63 VDD2.n43 9.69747
R2633 VDD2.n24 VDD2.n4 9.69747
R2634 VDD2.n73 VDD2.n72 9.45567
R2635 VDD2.n34 VDD2.n33 9.45567
R2636 VDD2.n72 VDD2.n71 9.3005
R2637 VDD2.n41 VDD2.n40 9.3005
R2638 VDD2.n66 VDD2.n65 9.3005
R2639 VDD2.n64 VDD2.n63 9.3005
R2640 VDD2.n45 VDD2.n44 9.3005
R2641 VDD2.n58 VDD2.n57 9.3005
R2642 VDD2.n56 VDD2.n55 9.3005
R2643 VDD2.n49 VDD2.n48 9.3005
R2644 VDD2.n2 VDD2.n1 9.3005
R2645 VDD2.n27 VDD2.n26 9.3005
R2646 VDD2.n25 VDD2.n24 9.3005
R2647 VDD2.n6 VDD2.n5 9.3005
R2648 VDD2.n19 VDD2.n18 9.3005
R2649 VDD2.n17 VDD2.n16 9.3005
R2650 VDD2.n10 VDD2.n9 9.3005
R2651 VDD2.n33 VDD2.n32 9.3005
R2652 VDD2.n67 VDD2.n66 8.92171
R2653 VDD2.n28 VDD2.n27 8.92171
R2654 VDD2.n70 VDD2.n41 8.14595
R2655 VDD2.n31 VDD2.n2 8.14595
R2656 VDD2.n71 VDD2.n39 7.3702
R2657 VDD2.n32 VDD2.n0 7.3702
R2658 VDD2.n73 VDD2.n39 6.59444
R2659 VDD2.n34 VDD2.n0 6.59444
R2660 VDD2.n71 VDD2.n70 5.81868
R2661 VDD2.n32 VDD2.n31 5.81868
R2662 VDD2.n67 VDD2.n41 5.04292
R2663 VDD2.n28 VDD2.n2 5.04292
R2664 VDD2.n50 VDD2.n48 4.38571
R2665 VDD2.n11 VDD2.n9 4.38571
R2666 VDD2.n66 VDD2.n43 4.26717
R2667 VDD2.n27 VDD2.n4 4.26717
R2668 VDD2.n63 VDD2.n62 3.49141
R2669 VDD2.n24 VDD2.n23 3.49141
R2670 VDD2.n76 VDD2.n74 3.19016
R2671 VDD2.n77 VDD2.t6 2.94255
R2672 VDD2.n77 VDD2.t4 2.94255
R2673 VDD2.n75 VDD2.t7 2.94255
R2674 VDD2.n75 VDD2.t2 2.94255
R2675 VDD2.n37 VDD2.t5 2.94255
R2676 VDD2.n37 VDD2.t1 2.94255
R2677 VDD2.n35 VDD2.t3 2.94255
R2678 VDD2.n35 VDD2.t0 2.94255
R2679 VDD2.n59 VDD2.n45 2.71565
R2680 VDD2.n20 VDD2.n6 2.71565
R2681 VDD2.n58 VDD2.n47 1.93989
R2682 VDD2.n19 VDD2.n8 1.93989
R2683 VDD2.n55 VDD2.n54 1.16414
R2684 VDD2.n16 VDD2.n15 1.16414
R2685 VDD2 VDD2.n76 0.856103
R2686 VDD2.n38 VDD2.n36 0.742568
R2687 VDD2.n51 VDD2.n49 0.388379
R2688 VDD2.n12 VDD2.n10 0.388379
R2689 VDD2.n72 VDD2.n40 0.155672
R2690 VDD2.n65 VDD2.n40 0.155672
R2691 VDD2.n65 VDD2.n64 0.155672
R2692 VDD2.n64 VDD2.n44 0.155672
R2693 VDD2.n57 VDD2.n44 0.155672
R2694 VDD2.n57 VDD2.n56 0.155672
R2695 VDD2.n56 VDD2.n48 0.155672
R2696 VDD2.n17 VDD2.n9 0.155672
R2697 VDD2.n18 VDD2.n17 0.155672
R2698 VDD2.n18 VDD2.n5 0.155672
R2699 VDD2.n25 VDD2.n5 0.155672
R2700 VDD2.n26 VDD2.n25 0.155672
R2701 VDD2.n26 VDD2.n1 0.155672
R2702 VDD2.n33 VDD2.n1 0.155672
C0 VDD1 VDD2 2.67584f
C1 VN VP 8.562611f
C2 VN VTAIL 7.96589f
C3 VDD1 VP 7.02562f
C4 VDD2 VP 0.681531f
C5 VDD1 VTAIL 8.570331f
C6 VDD2 VTAIL 8.628059f
C7 VDD1 VN 0.155169f
C8 VDD2 VN 6.50244f
C9 VTAIL VP 7.98007f
C10 VDD2 B 7.233233f
C11 VDD1 B 7.160848f
C12 VTAIL B 6.124303f
C13 VN B 21.202488f
C14 VP B 19.764212f
C15 VDD2.n0 B 0.037836f
C16 VDD2.n1 B 0.026287f
C17 VDD2.n2 B 0.014126f
C18 VDD2.n3 B 0.033388f
C19 VDD2.n4 B 0.014957f
C20 VDD2.n5 B 0.026287f
C21 VDD2.n6 B 0.014126f
C22 VDD2.n7 B 0.033388f
C23 VDD2.n8 B 0.014957f
C24 VDD2.n9 B 0.71367f
C25 VDD2.n10 B 0.014126f
C26 VDD2.t8 B 0.054403f
C27 VDD2.n11 B 0.117143f
C28 VDD2.n12 B 0.019723f
C29 VDD2.n13 B 0.025041f
C30 VDD2.n14 B 0.033388f
C31 VDD2.n15 B 0.014957f
C32 VDD2.n16 B 0.014126f
C33 VDD2.n17 B 0.026287f
C34 VDD2.n18 B 0.026287f
C35 VDD2.n19 B 0.014126f
C36 VDD2.n20 B 0.014957f
C37 VDD2.n21 B 0.033388f
C38 VDD2.n22 B 0.033388f
C39 VDD2.n23 B 0.014957f
C40 VDD2.n24 B 0.014126f
C41 VDD2.n25 B 0.026287f
C42 VDD2.n26 B 0.026287f
C43 VDD2.n27 B 0.014126f
C44 VDD2.n28 B 0.014957f
C45 VDD2.n29 B 0.033388f
C46 VDD2.n30 B 0.073848f
C47 VDD2.n31 B 0.014957f
C48 VDD2.n32 B 0.014126f
C49 VDD2.n33 B 0.061121f
C50 VDD2.n34 B 0.079238f
C51 VDD2.t3 B 0.139803f
C52 VDD2.t0 B 0.139803f
C53 VDD2.n35 B 1.1816f
C54 VDD2.n36 B 0.850789f
C55 VDD2.t5 B 0.139803f
C56 VDD2.t1 B 0.139803f
C57 VDD2.n37 B 1.20526f
C58 VDD2.n38 B 3.13638f
C59 VDD2.n39 B 0.037836f
C60 VDD2.n40 B 0.026287f
C61 VDD2.n41 B 0.014126f
C62 VDD2.n42 B 0.033388f
C63 VDD2.n43 B 0.014957f
C64 VDD2.n44 B 0.026287f
C65 VDD2.n45 B 0.014126f
C66 VDD2.n46 B 0.033388f
C67 VDD2.n47 B 0.014957f
C68 VDD2.n48 B 0.71367f
C69 VDD2.n49 B 0.014126f
C70 VDD2.t9 B 0.054403f
C71 VDD2.n50 B 0.117143f
C72 VDD2.n51 B 0.019723f
C73 VDD2.n52 B 0.025041f
C74 VDD2.n53 B 0.033388f
C75 VDD2.n54 B 0.014957f
C76 VDD2.n55 B 0.014126f
C77 VDD2.n56 B 0.026287f
C78 VDD2.n57 B 0.026287f
C79 VDD2.n58 B 0.014126f
C80 VDD2.n59 B 0.014957f
C81 VDD2.n60 B 0.033388f
C82 VDD2.n61 B 0.033388f
C83 VDD2.n62 B 0.014957f
C84 VDD2.n63 B 0.014126f
C85 VDD2.n64 B 0.026287f
C86 VDD2.n65 B 0.026287f
C87 VDD2.n66 B 0.014126f
C88 VDD2.n67 B 0.014957f
C89 VDD2.n68 B 0.033388f
C90 VDD2.n69 B 0.073848f
C91 VDD2.n70 B 0.014957f
C92 VDD2.n71 B 0.014126f
C93 VDD2.n72 B 0.061121f
C94 VDD2.n73 B 0.059641f
C95 VDD2.n74 B 2.92602f
C96 VDD2.t7 B 0.139803f
C97 VDD2.t2 B 0.139803f
C98 VDD2.n75 B 1.18161f
C99 VDD2.n76 B 0.558176f
C100 VDD2.t6 B 0.139803f
C101 VDD2.t4 B 0.139803f
C102 VDD2.n77 B 1.20521f
C103 VN.t8 B 1.22904f
C104 VN.n0 B 0.522539f
C105 VN.n1 B 0.020344f
C106 VN.n2 B 0.026864f
C107 VN.n3 B 0.020344f
C108 VN.n4 B 0.021069f
C109 VN.n5 B 0.020344f
C110 VN.n6 B 0.019219f
C111 VN.n7 B 0.020344f
C112 VN.t9 B 1.22904f
C113 VN.n8 B 0.449747f
C114 VN.n9 B 0.020344f
C115 VN.n10 B 0.019219f
C116 VN.n11 B 0.020344f
C117 VN.t6 B 1.22904f
C118 VN.n12 B 0.527141f
C119 VN.t1 B 1.47186f
C120 VN.n13 B 0.498236f
C121 VN.n14 B 0.249004f
C122 VN.n15 B 0.036045f
C123 VN.n16 B 0.037917f
C124 VN.n17 B 0.037339f
C125 VN.n18 B 0.020344f
C126 VN.n19 B 0.020344f
C127 VN.n20 B 0.020344f
C128 VN.n21 B 0.040756f
C129 VN.n22 B 0.037917f
C130 VN.n23 B 0.028557f
C131 VN.n24 B 0.020344f
C132 VN.n25 B 0.020344f
C133 VN.n26 B 0.028557f
C134 VN.n27 B 0.037917f
C135 VN.n28 B 0.040756f
C136 VN.n29 B 0.020344f
C137 VN.n30 B 0.020344f
C138 VN.n31 B 0.020344f
C139 VN.n32 B 0.037339f
C140 VN.n33 B 0.037917f
C141 VN.t4 B 1.22904f
C142 VN.n34 B 0.449747f
C143 VN.n35 B 0.036045f
C144 VN.n36 B 0.020344f
C145 VN.n37 B 0.020344f
C146 VN.n38 B 0.020344f
C147 VN.n39 B 0.037917f
C148 VN.n40 B 0.037917f
C149 VN.n41 B 0.032534f
C150 VN.n42 B 0.020344f
C151 VN.n43 B 0.020344f
C152 VN.n44 B 0.020344f
C153 VN.n45 B 0.037917f
C154 VN.n46 B 0.037917f
C155 VN.n47 B 0.024813f
C156 VN.n48 B 0.032835f
C157 VN.n49 B 0.055124f
C158 VN.t0 B 1.22904f
C159 VN.n50 B 0.522539f
C160 VN.n51 B 0.020344f
C161 VN.n52 B 0.026864f
C162 VN.n53 B 0.020344f
C163 VN.n54 B 0.021069f
C164 VN.n55 B 0.020344f
C165 VN.t2 B 1.22904f
C166 VN.n56 B 0.449747f
C167 VN.n57 B 0.019219f
C168 VN.n58 B 0.020344f
C169 VN.t7 B 1.22904f
C170 VN.n59 B 0.449747f
C171 VN.n60 B 0.020344f
C172 VN.n61 B 0.019219f
C173 VN.n62 B 0.020344f
C174 VN.t3 B 1.22904f
C175 VN.n63 B 0.527141f
C176 VN.t5 B 1.47186f
C177 VN.n64 B 0.498237f
C178 VN.n65 B 0.249004f
C179 VN.n66 B 0.036045f
C180 VN.n67 B 0.037917f
C181 VN.n68 B 0.037339f
C182 VN.n69 B 0.020344f
C183 VN.n70 B 0.020344f
C184 VN.n71 B 0.020344f
C185 VN.n72 B 0.040756f
C186 VN.n73 B 0.037917f
C187 VN.n74 B 0.028557f
C188 VN.n75 B 0.020344f
C189 VN.n76 B 0.020344f
C190 VN.n77 B 0.028557f
C191 VN.n78 B 0.037917f
C192 VN.n79 B 0.040756f
C193 VN.n80 B 0.020344f
C194 VN.n81 B 0.020344f
C195 VN.n82 B 0.020344f
C196 VN.n83 B 0.037339f
C197 VN.n84 B 0.037917f
C198 VN.n85 B 0.036045f
C199 VN.n86 B 0.020344f
C200 VN.n87 B 0.020344f
C201 VN.n88 B 0.020344f
C202 VN.n89 B 0.037917f
C203 VN.n90 B 0.037917f
C204 VN.n91 B 0.032534f
C205 VN.n92 B 0.020344f
C206 VN.n93 B 0.020344f
C207 VN.n94 B 0.020344f
C208 VN.n95 B 0.037917f
C209 VN.n96 B 0.037917f
C210 VN.n97 B 0.024813f
C211 VN.n98 B 0.032835f
C212 VN.n99 B 1.28041f
C213 VDD1.n0 B 0.038688f
C214 VDD1.n1 B 0.026879f
C215 VDD1.n2 B 0.014444f
C216 VDD1.n3 B 0.03414f
C217 VDD1.n4 B 0.015293f
C218 VDD1.n5 B 0.026879f
C219 VDD1.n6 B 0.014444f
C220 VDD1.n7 B 0.03414f
C221 VDD1.n8 B 0.015293f
C222 VDD1.n9 B 0.729737f
C223 VDD1.n10 B 0.014444f
C224 VDD1.t1 B 0.055628f
C225 VDD1.n11 B 0.11978f
C226 VDD1.n12 B 0.020167f
C227 VDD1.n13 B 0.025605f
C228 VDD1.n14 B 0.03414f
C229 VDD1.n15 B 0.015293f
C230 VDD1.n16 B 0.014444f
C231 VDD1.n17 B 0.026879f
C232 VDD1.n18 B 0.026879f
C233 VDD1.n19 B 0.014444f
C234 VDD1.n20 B 0.015293f
C235 VDD1.n21 B 0.03414f
C236 VDD1.n22 B 0.03414f
C237 VDD1.n23 B 0.015293f
C238 VDD1.n24 B 0.014444f
C239 VDD1.n25 B 0.026879f
C240 VDD1.n26 B 0.026879f
C241 VDD1.n27 B 0.014444f
C242 VDD1.n28 B 0.015293f
C243 VDD1.n29 B 0.03414f
C244 VDD1.n30 B 0.07551f
C245 VDD1.n31 B 0.015293f
C246 VDD1.n32 B 0.014444f
C247 VDD1.n33 B 0.062497f
C248 VDD1.n34 B 0.081021f
C249 VDD1.t2 B 0.14295f
C250 VDD1.t4 B 0.14295f
C251 VDD1.n35 B 1.20821f
C252 VDD1.n36 B 0.878931f
C253 VDD1.n37 B 0.038688f
C254 VDD1.n38 B 0.026879f
C255 VDD1.n39 B 0.014444f
C256 VDD1.n40 B 0.03414f
C257 VDD1.n41 B 0.015293f
C258 VDD1.n42 B 0.026879f
C259 VDD1.n43 B 0.014444f
C260 VDD1.n44 B 0.03414f
C261 VDD1.n45 B 0.015293f
C262 VDD1.n46 B 0.729737f
C263 VDD1.n47 B 0.014444f
C264 VDD1.t0 B 0.055628f
C265 VDD1.n48 B 0.11978f
C266 VDD1.n49 B 0.020167f
C267 VDD1.n50 B 0.025605f
C268 VDD1.n51 B 0.03414f
C269 VDD1.n52 B 0.015293f
C270 VDD1.n53 B 0.014444f
C271 VDD1.n54 B 0.026879f
C272 VDD1.n55 B 0.026879f
C273 VDD1.n56 B 0.014444f
C274 VDD1.n57 B 0.015293f
C275 VDD1.n58 B 0.03414f
C276 VDD1.n59 B 0.03414f
C277 VDD1.n60 B 0.015293f
C278 VDD1.n61 B 0.014444f
C279 VDD1.n62 B 0.026879f
C280 VDD1.n63 B 0.026879f
C281 VDD1.n64 B 0.014444f
C282 VDD1.n65 B 0.015293f
C283 VDD1.n66 B 0.03414f
C284 VDD1.n67 B 0.07551f
C285 VDD1.n68 B 0.015293f
C286 VDD1.n69 B 0.014444f
C287 VDD1.n70 B 0.062497f
C288 VDD1.n71 B 0.081021f
C289 VDD1.t5 B 0.14295f
C290 VDD1.t9 B 0.14295f
C291 VDD1.n72 B 1.2082f
C292 VDD1.n73 B 0.869943f
C293 VDD1.t3 B 0.14295f
C294 VDD1.t8 B 0.14295f
C295 VDD1.n74 B 1.23239f
C296 VDD1.n75 B 3.35912f
C297 VDD1.t6 B 0.14295f
C298 VDD1.t7 B 0.14295f
C299 VDD1.n76 B 1.2082f
C300 VDD1.n77 B 3.32043f
C301 VTAIL.t6 B 0.154016f
C302 VTAIL.t7 B 0.154016f
C303 VTAIL.n0 B 1.22372f
C304 VTAIL.n1 B 0.697416f
C305 VTAIL.n2 B 0.041683f
C306 VTAIL.n3 B 0.02896f
C307 VTAIL.n4 B 0.015562f
C308 VTAIL.n5 B 0.036782f
C309 VTAIL.n6 B 0.016477f
C310 VTAIL.n7 B 0.02896f
C311 VTAIL.n8 B 0.015562f
C312 VTAIL.n9 B 0.036782f
C313 VTAIL.n10 B 0.016477f
C314 VTAIL.n11 B 0.786223f
C315 VTAIL.n12 B 0.015562f
C316 VTAIL.t15 B 0.059934f
C317 VTAIL.n13 B 0.129052f
C318 VTAIL.n14 B 0.021728f
C319 VTAIL.n15 B 0.027587f
C320 VTAIL.n16 B 0.036782f
C321 VTAIL.n17 B 0.016477f
C322 VTAIL.n18 B 0.015562f
C323 VTAIL.n19 B 0.02896f
C324 VTAIL.n20 B 0.02896f
C325 VTAIL.n21 B 0.015562f
C326 VTAIL.n22 B 0.016477f
C327 VTAIL.n23 B 0.036782f
C328 VTAIL.n24 B 0.036782f
C329 VTAIL.n25 B 0.016477f
C330 VTAIL.n26 B 0.015562f
C331 VTAIL.n27 B 0.02896f
C332 VTAIL.n28 B 0.02896f
C333 VTAIL.n29 B 0.015562f
C334 VTAIL.n30 B 0.016477f
C335 VTAIL.n31 B 0.036782f
C336 VTAIL.n32 B 0.081355f
C337 VTAIL.n33 B 0.016477f
C338 VTAIL.n34 B 0.015562f
C339 VTAIL.n35 B 0.067335f
C340 VTAIL.n36 B 0.045711f
C341 VTAIL.n37 B 0.515263f
C342 VTAIL.t13 B 0.154016f
C343 VTAIL.t19 B 0.154016f
C344 VTAIL.n38 B 1.22372f
C345 VTAIL.n39 B 0.871376f
C346 VTAIL.t16 B 0.154016f
C347 VTAIL.t12 B 0.154016f
C348 VTAIL.n40 B 1.22372f
C349 VTAIL.n41 B 2.10379f
C350 VTAIL.t2 B 0.154016f
C351 VTAIL.t4 B 0.154016f
C352 VTAIL.n42 B 1.22373f
C353 VTAIL.n43 B 2.10378f
C354 VTAIL.t1 B 0.154016f
C355 VTAIL.t3 B 0.154016f
C356 VTAIL.n44 B 1.22373f
C357 VTAIL.n45 B 0.871368f
C358 VTAIL.n46 B 0.041683f
C359 VTAIL.n47 B 0.02896f
C360 VTAIL.n48 B 0.015562f
C361 VTAIL.n49 B 0.036782f
C362 VTAIL.n50 B 0.016477f
C363 VTAIL.n51 B 0.02896f
C364 VTAIL.n52 B 0.015562f
C365 VTAIL.n53 B 0.036782f
C366 VTAIL.n54 B 0.016477f
C367 VTAIL.n55 B 0.786223f
C368 VTAIL.n56 B 0.015562f
C369 VTAIL.t9 B 0.059934f
C370 VTAIL.n57 B 0.129052f
C371 VTAIL.n58 B 0.021728f
C372 VTAIL.n59 B 0.027587f
C373 VTAIL.n60 B 0.036782f
C374 VTAIL.n61 B 0.016477f
C375 VTAIL.n62 B 0.015562f
C376 VTAIL.n63 B 0.02896f
C377 VTAIL.n64 B 0.02896f
C378 VTAIL.n65 B 0.015562f
C379 VTAIL.n66 B 0.016477f
C380 VTAIL.n67 B 0.036782f
C381 VTAIL.n68 B 0.036782f
C382 VTAIL.n69 B 0.016477f
C383 VTAIL.n70 B 0.015562f
C384 VTAIL.n71 B 0.02896f
C385 VTAIL.n72 B 0.02896f
C386 VTAIL.n73 B 0.015562f
C387 VTAIL.n74 B 0.016477f
C388 VTAIL.n75 B 0.036782f
C389 VTAIL.n76 B 0.081355f
C390 VTAIL.n77 B 0.016477f
C391 VTAIL.n78 B 0.015562f
C392 VTAIL.n79 B 0.067335f
C393 VTAIL.n80 B 0.045711f
C394 VTAIL.n81 B 0.515263f
C395 VTAIL.t18 B 0.154016f
C396 VTAIL.t11 B 0.154016f
C397 VTAIL.n82 B 1.22373f
C398 VTAIL.n83 B 0.766388f
C399 VTAIL.t14 B 0.154016f
C400 VTAIL.t17 B 0.154016f
C401 VTAIL.n84 B 1.22373f
C402 VTAIL.n85 B 0.871368f
C403 VTAIL.n86 B 0.041683f
C404 VTAIL.n87 B 0.02896f
C405 VTAIL.n88 B 0.015562f
C406 VTAIL.n89 B 0.036782f
C407 VTAIL.n90 B 0.016477f
C408 VTAIL.n91 B 0.02896f
C409 VTAIL.n92 B 0.015562f
C410 VTAIL.n93 B 0.036782f
C411 VTAIL.n94 B 0.016477f
C412 VTAIL.n95 B 0.786223f
C413 VTAIL.n96 B 0.015562f
C414 VTAIL.t10 B 0.059934f
C415 VTAIL.n97 B 0.129052f
C416 VTAIL.n98 B 0.021728f
C417 VTAIL.n99 B 0.027587f
C418 VTAIL.n100 B 0.036782f
C419 VTAIL.n101 B 0.016477f
C420 VTAIL.n102 B 0.015562f
C421 VTAIL.n103 B 0.02896f
C422 VTAIL.n104 B 0.02896f
C423 VTAIL.n105 B 0.015562f
C424 VTAIL.n106 B 0.016477f
C425 VTAIL.n107 B 0.036782f
C426 VTAIL.n108 B 0.036782f
C427 VTAIL.n109 B 0.016477f
C428 VTAIL.n110 B 0.015562f
C429 VTAIL.n111 B 0.02896f
C430 VTAIL.n112 B 0.02896f
C431 VTAIL.n113 B 0.015562f
C432 VTAIL.n114 B 0.016477f
C433 VTAIL.n115 B 0.036782f
C434 VTAIL.n116 B 0.081355f
C435 VTAIL.n117 B 0.016477f
C436 VTAIL.n118 B 0.015562f
C437 VTAIL.n119 B 0.067335f
C438 VTAIL.n120 B 0.045711f
C439 VTAIL.n121 B 1.55502f
C440 VTAIL.n122 B 0.041683f
C441 VTAIL.n123 B 0.02896f
C442 VTAIL.n124 B 0.015562f
C443 VTAIL.n125 B 0.036782f
C444 VTAIL.n126 B 0.016477f
C445 VTAIL.n127 B 0.02896f
C446 VTAIL.n128 B 0.015562f
C447 VTAIL.n129 B 0.036782f
C448 VTAIL.n130 B 0.016477f
C449 VTAIL.n131 B 0.786223f
C450 VTAIL.n132 B 0.015562f
C451 VTAIL.t5 B 0.059934f
C452 VTAIL.n133 B 0.129052f
C453 VTAIL.n134 B 0.021728f
C454 VTAIL.n135 B 0.027587f
C455 VTAIL.n136 B 0.036782f
C456 VTAIL.n137 B 0.016477f
C457 VTAIL.n138 B 0.015562f
C458 VTAIL.n139 B 0.02896f
C459 VTAIL.n140 B 0.02896f
C460 VTAIL.n141 B 0.015562f
C461 VTAIL.n142 B 0.016477f
C462 VTAIL.n143 B 0.036782f
C463 VTAIL.n144 B 0.036782f
C464 VTAIL.n145 B 0.016477f
C465 VTAIL.n146 B 0.015562f
C466 VTAIL.n147 B 0.02896f
C467 VTAIL.n148 B 0.02896f
C468 VTAIL.n149 B 0.015562f
C469 VTAIL.n150 B 0.016477f
C470 VTAIL.n151 B 0.036782f
C471 VTAIL.n152 B 0.081355f
C472 VTAIL.n153 B 0.016477f
C473 VTAIL.n154 B 0.015562f
C474 VTAIL.n155 B 0.067335f
C475 VTAIL.n156 B 0.045711f
C476 VTAIL.n157 B 1.55502f
C477 VTAIL.t0 B 0.154016f
C478 VTAIL.t8 B 0.154016f
C479 VTAIL.n158 B 1.22372f
C480 VTAIL.n159 B 0.642714f
C481 VP.t1 B 1.2572f
C482 VP.n0 B 0.534511f
C483 VP.n1 B 0.02081f
C484 VP.n2 B 0.02748f
C485 VP.n3 B 0.02081f
C486 VP.n4 B 0.021552f
C487 VP.n5 B 0.02081f
C488 VP.n6 B 0.019659f
C489 VP.n7 B 0.02081f
C490 VP.t0 B 1.2572f
C491 VP.n8 B 0.460052f
C492 VP.n9 B 0.02081f
C493 VP.n10 B 0.019659f
C494 VP.n11 B 0.02081f
C495 VP.t4 B 1.2572f
C496 VP.n12 B 0.460052f
C497 VP.n13 B 0.02081f
C498 VP.n14 B 0.033279f
C499 VP.n15 B 0.02081f
C500 VP.n16 B 0.025381f
C501 VP.t2 B 1.2572f
C502 VP.n17 B 0.534511f
C503 VP.n18 B 0.02081f
C504 VP.n19 B 0.02748f
C505 VP.n20 B 0.02081f
C506 VP.n21 B 0.021552f
C507 VP.n22 B 0.02081f
C508 VP.n23 B 0.019659f
C509 VP.n24 B 0.02081f
C510 VP.t5 B 1.2572f
C511 VP.n25 B 0.460052f
C512 VP.n26 B 0.02081f
C513 VP.n27 B 0.019659f
C514 VP.n28 B 0.02081f
C515 VP.t7 B 1.2572f
C516 VP.n29 B 0.539219f
C517 VP.t8 B 1.50558f
C518 VP.n30 B 0.509652f
C519 VP.n31 B 0.254709f
C520 VP.n32 B 0.03687f
C521 VP.n33 B 0.038785f
C522 VP.n34 B 0.038194f
C523 VP.n35 B 0.02081f
C524 VP.n36 B 0.02081f
C525 VP.n37 B 0.02081f
C526 VP.n38 B 0.04169f
C527 VP.n39 B 0.038785f
C528 VP.n40 B 0.029211f
C529 VP.n41 B 0.02081f
C530 VP.n42 B 0.02081f
C531 VP.n43 B 0.029211f
C532 VP.n44 B 0.038785f
C533 VP.n45 B 0.04169f
C534 VP.n46 B 0.02081f
C535 VP.n47 B 0.02081f
C536 VP.n48 B 0.02081f
C537 VP.n49 B 0.038194f
C538 VP.n50 B 0.038785f
C539 VP.t3 B 1.2572f
C540 VP.n51 B 0.460052f
C541 VP.n52 B 0.03687f
C542 VP.n53 B 0.02081f
C543 VP.n54 B 0.02081f
C544 VP.n55 B 0.02081f
C545 VP.n56 B 0.038785f
C546 VP.n57 B 0.038785f
C547 VP.n58 B 0.033279f
C548 VP.n59 B 0.02081f
C549 VP.n60 B 0.02081f
C550 VP.n61 B 0.02081f
C551 VP.n62 B 0.038785f
C552 VP.n63 B 0.038785f
C553 VP.n64 B 0.025381f
C554 VP.n65 B 0.033587f
C555 VP.n66 B 1.3014f
C556 VP.t9 B 1.2572f
C557 VP.n67 B 0.534511f
C558 VP.n68 B 1.31543f
C559 VP.n69 B 0.033587f
C560 VP.n70 B 0.02081f
C561 VP.n71 B 0.038785f
C562 VP.n72 B 0.038785f
C563 VP.n73 B 0.02748f
C564 VP.n74 B 0.02081f
C565 VP.n75 B 0.02081f
C566 VP.n76 B 0.02081f
C567 VP.n77 B 0.038785f
C568 VP.n78 B 0.038785f
C569 VP.n79 B 0.021552f
C570 VP.n80 B 0.02081f
C571 VP.n81 B 0.02081f
C572 VP.n82 B 0.03687f
C573 VP.n83 B 0.038785f
C574 VP.n84 B 0.038194f
C575 VP.n85 B 0.02081f
C576 VP.n86 B 0.02081f
C577 VP.n87 B 0.02081f
C578 VP.n88 B 0.04169f
C579 VP.n89 B 0.038785f
C580 VP.n90 B 0.029211f
C581 VP.n91 B 0.02081f
C582 VP.n92 B 0.02081f
C583 VP.n93 B 0.029211f
C584 VP.n94 B 0.038785f
C585 VP.n95 B 0.04169f
C586 VP.n96 B 0.02081f
C587 VP.n97 B 0.02081f
C588 VP.n98 B 0.02081f
C589 VP.n99 B 0.038194f
C590 VP.n100 B 0.038785f
C591 VP.t6 B 1.2572f
C592 VP.n101 B 0.460052f
C593 VP.n102 B 0.03687f
C594 VP.n103 B 0.02081f
C595 VP.n104 B 0.02081f
C596 VP.n105 B 0.02081f
C597 VP.n106 B 0.038785f
C598 VP.n107 B 0.038785f
C599 VP.n108 B 0.033279f
C600 VP.n109 B 0.02081f
C601 VP.n110 B 0.02081f
C602 VP.n111 B 0.02081f
C603 VP.n112 B 0.038785f
C604 VP.n113 B 0.038785f
C605 VP.n114 B 0.025381f
C606 VP.n115 B 0.033587f
C607 VP.n116 B 0.056387f
.ends

