* NGSPICE file created from diff_pair_sample_0245.ext - technology: sky130A

.subckt diff_pair_sample_0245 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t13 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.69
X1 B.t11 B.t9 B.t10 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.69
X2 VTAIL.t6 VP.t0 VDD1.t9 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X3 VDD2.t8 VN.t1 VTAIL.t10 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X4 VDD1.t8 VP.t1 VTAIL.t19 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X5 VDD1.t7 VP.t2 VTAIL.t3 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.69
X6 VTAIL.t2 VP.t3 VDD1.t6 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X7 VTAIL.t12 VN.t2 VDD2.t7 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X8 VTAIL.t0 VP.t4 VDD1.t5 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X9 VDD1.t4 VP.t5 VTAIL.t1 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.69
X10 VDD2.t6 VN.t3 VTAIL.t9 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.69
X11 VDD1.t3 VP.t6 VTAIL.t4 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X12 VDD2.t5 VN.t4 VTAIL.t18 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.69
X13 VDD2.t4 VN.t5 VTAIL.t11 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.69
X14 VTAIL.t17 VN.t6 VDD2.t3 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X15 VDD1.t2 VP.t7 VTAIL.t7 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=2.0709 ps=11.4 w=5.31 l=3.69
X16 VTAIL.t5 VP.t8 VDD1.t1 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X17 B.t8 B.t6 B.t7 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.69
X18 VTAIL.t16 VN.t7 VDD2.t2 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X19 B.t5 B.t3 B.t4 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.69
X20 VDD2.t1 VN.t8 VTAIL.t15 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X21 B.t2 B.t0 B.t1 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0 ps=0 w=5.31 l=3.69
X22 VTAIL.t14 VN.t9 VDD2.t0 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=0.87615 pd=5.64 as=0.87615 ps=5.64 w=5.31 l=3.69
X23 VDD1.t0 VP.t9 VTAIL.t8 w_n5794_n2030# sky130_fd_pr__pfet_01v8 ad=2.0709 pd=11.4 as=0.87615 ps=5.64 w=5.31 l=3.69
R0 VN.n108 VN.n107 161.3
R1 VN.n106 VN.n56 161.3
R2 VN.n105 VN.n104 161.3
R3 VN.n103 VN.n57 161.3
R4 VN.n102 VN.n101 161.3
R5 VN.n100 VN.n58 161.3
R6 VN.n99 VN.n98 161.3
R7 VN.n97 VN.n59 161.3
R8 VN.n96 VN.n95 161.3
R9 VN.n94 VN.n60 161.3
R10 VN.n93 VN.n92 161.3
R11 VN.n91 VN.n62 161.3
R12 VN.n90 VN.n89 161.3
R13 VN.n88 VN.n63 161.3
R14 VN.n87 VN.n86 161.3
R15 VN.n85 VN.n64 161.3
R16 VN.n84 VN.n83 161.3
R17 VN.n82 VN.n65 161.3
R18 VN.n81 VN.n80 161.3
R19 VN.n79 VN.n66 161.3
R20 VN.n78 VN.n77 161.3
R21 VN.n76 VN.n67 161.3
R22 VN.n75 VN.n74 161.3
R23 VN.n73 VN.n68 161.3
R24 VN.n72 VN.n71 161.3
R25 VN.n53 VN.n52 161.3
R26 VN.n51 VN.n1 161.3
R27 VN.n50 VN.n49 161.3
R28 VN.n48 VN.n2 161.3
R29 VN.n47 VN.n46 161.3
R30 VN.n45 VN.n3 161.3
R31 VN.n44 VN.n43 161.3
R32 VN.n42 VN.n4 161.3
R33 VN.n41 VN.n40 161.3
R34 VN.n38 VN.n5 161.3
R35 VN.n37 VN.n36 161.3
R36 VN.n35 VN.n6 161.3
R37 VN.n34 VN.n33 161.3
R38 VN.n32 VN.n7 161.3
R39 VN.n31 VN.n30 161.3
R40 VN.n29 VN.n8 161.3
R41 VN.n28 VN.n27 161.3
R42 VN.n26 VN.n9 161.3
R43 VN.n25 VN.n24 161.3
R44 VN.n23 VN.n10 161.3
R45 VN.n22 VN.n21 161.3
R46 VN.n20 VN.n11 161.3
R47 VN.n19 VN.n18 161.3
R48 VN.n17 VN.n12 161.3
R49 VN.n16 VN.n15 161.3
R50 VN.n54 VN.n0 88.1101
R51 VN.n109 VN.n55 88.1101
R52 VN.n14 VN.n13 74.0089
R53 VN.n70 VN.n69 74.0089
R54 VN.n69 VN.t4 66.2847
R55 VN.n13 VN.t0 66.2847
R56 VN VN.n109 54.1495
R57 VN.n46 VN.n2 43.4072
R58 VN.n101 VN.n57 43.4072
R59 VN.n21 VN.n20 41.4647
R60 VN.n33 VN.n6 41.4647
R61 VN.n77 VN.n76 41.4647
R62 VN.n89 VN.n62 41.4647
R63 VN.n21 VN.n10 39.5221
R64 VN.n33 VN.n32 39.5221
R65 VN.n77 VN.n66 39.5221
R66 VN.n89 VN.n88 39.5221
R67 VN.n46 VN.n45 37.5796
R68 VN.n101 VN.n100 37.5796
R69 VN.n27 VN.t8 34.681
R70 VN.n14 VN.t9 34.681
R71 VN.n39 VN.t6 34.681
R72 VN.n0 VN.t5 34.681
R73 VN.n83 VN.t1 34.681
R74 VN.n70 VN.t7 34.681
R75 VN.n61 VN.t2 34.681
R76 VN.n55 VN.t3 34.681
R77 VN.n15 VN.n12 24.4675
R78 VN.n19 VN.n12 24.4675
R79 VN.n20 VN.n19 24.4675
R80 VN.n25 VN.n10 24.4675
R81 VN.n26 VN.n25 24.4675
R82 VN.n27 VN.n26 24.4675
R83 VN.n27 VN.n8 24.4675
R84 VN.n31 VN.n8 24.4675
R85 VN.n32 VN.n31 24.4675
R86 VN.n37 VN.n6 24.4675
R87 VN.n38 VN.n37 24.4675
R88 VN.n40 VN.n38 24.4675
R89 VN.n44 VN.n4 24.4675
R90 VN.n45 VN.n44 24.4675
R91 VN.n50 VN.n2 24.4675
R92 VN.n51 VN.n50 24.4675
R93 VN.n52 VN.n51 24.4675
R94 VN.n76 VN.n75 24.4675
R95 VN.n75 VN.n68 24.4675
R96 VN.n71 VN.n68 24.4675
R97 VN.n88 VN.n87 24.4675
R98 VN.n87 VN.n64 24.4675
R99 VN.n83 VN.n64 24.4675
R100 VN.n83 VN.n82 24.4675
R101 VN.n82 VN.n81 24.4675
R102 VN.n81 VN.n66 24.4675
R103 VN.n100 VN.n99 24.4675
R104 VN.n99 VN.n59 24.4675
R105 VN.n95 VN.n94 24.4675
R106 VN.n94 VN.n93 24.4675
R107 VN.n93 VN.n62 24.4675
R108 VN.n107 VN.n106 24.4675
R109 VN.n106 VN.n105 24.4675
R110 VN.n105 VN.n57 24.4675
R111 VN.n39 VN.n4 23.4888
R112 VN.n61 VN.n59 23.4888
R113 VN.n72 VN.n69 3.40897
R114 VN.n16 VN.n13 3.40897
R115 VN.n52 VN.n0 1.95786
R116 VN.n107 VN.n55 1.95786
R117 VN.n15 VN.n14 0.97918
R118 VN.n40 VN.n39 0.97918
R119 VN.n71 VN.n70 0.97918
R120 VN.n95 VN.n61 0.97918
R121 VN.n109 VN.n108 0.354971
R122 VN.n54 VN.n53 0.354971
R123 VN VN.n54 0.26696
R124 VN.n108 VN.n56 0.189894
R125 VN.n104 VN.n56 0.189894
R126 VN.n104 VN.n103 0.189894
R127 VN.n103 VN.n102 0.189894
R128 VN.n102 VN.n58 0.189894
R129 VN.n98 VN.n58 0.189894
R130 VN.n98 VN.n97 0.189894
R131 VN.n97 VN.n96 0.189894
R132 VN.n96 VN.n60 0.189894
R133 VN.n92 VN.n60 0.189894
R134 VN.n92 VN.n91 0.189894
R135 VN.n91 VN.n90 0.189894
R136 VN.n90 VN.n63 0.189894
R137 VN.n86 VN.n63 0.189894
R138 VN.n86 VN.n85 0.189894
R139 VN.n85 VN.n84 0.189894
R140 VN.n84 VN.n65 0.189894
R141 VN.n80 VN.n65 0.189894
R142 VN.n80 VN.n79 0.189894
R143 VN.n79 VN.n78 0.189894
R144 VN.n78 VN.n67 0.189894
R145 VN.n74 VN.n67 0.189894
R146 VN.n74 VN.n73 0.189894
R147 VN.n73 VN.n72 0.189894
R148 VN.n17 VN.n16 0.189894
R149 VN.n18 VN.n17 0.189894
R150 VN.n18 VN.n11 0.189894
R151 VN.n22 VN.n11 0.189894
R152 VN.n23 VN.n22 0.189894
R153 VN.n24 VN.n23 0.189894
R154 VN.n24 VN.n9 0.189894
R155 VN.n28 VN.n9 0.189894
R156 VN.n29 VN.n28 0.189894
R157 VN.n30 VN.n29 0.189894
R158 VN.n30 VN.n7 0.189894
R159 VN.n34 VN.n7 0.189894
R160 VN.n35 VN.n34 0.189894
R161 VN.n36 VN.n35 0.189894
R162 VN.n36 VN.n5 0.189894
R163 VN.n41 VN.n5 0.189894
R164 VN.n42 VN.n41 0.189894
R165 VN.n43 VN.n42 0.189894
R166 VN.n43 VN.n3 0.189894
R167 VN.n47 VN.n3 0.189894
R168 VN.n48 VN.n47 0.189894
R169 VN.n49 VN.n48 0.189894
R170 VN.n49 VN.n1 0.189894
R171 VN.n53 VN.n1 0.189894
R172 VTAIL.n120 VTAIL.n98 756.745
R173 VTAIL.n24 VTAIL.n2 756.745
R174 VTAIL.n92 VTAIL.n70 756.745
R175 VTAIL.n60 VTAIL.n38 756.745
R176 VTAIL.n106 VTAIL.n105 585
R177 VTAIL.n111 VTAIL.n110 585
R178 VTAIL.n113 VTAIL.n112 585
R179 VTAIL.n102 VTAIL.n101 585
R180 VTAIL.n119 VTAIL.n118 585
R181 VTAIL.n121 VTAIL.n120 585
R182 VTAIL.n10 VTAIL.n9 585
R183 VTAIL.n15 VTAIL.n14 585
R184 VTAIL.n17 VTAIL.n16 585
R185 VTAIL.n6 VTAIL.n5 585
R186 VTAIL.n23 VTAIL.n22 585
R187 VTAIL.n25 VTAIL.n24 585
R188 VTAIL.n93 VTAIL.n92 585
R189 VTAIL.n91 VTAIL.n90 585
R190 VTAIL.n74 VTAIL.n73 585
R191 VTAIL.n85 VTAIL.n84 585
R192 VTAIL.n83 VTAIL.n82 585
R193 VTAIL.n78 VTAIL.n77 585
R194 VTAIL.n61 VTAIL.n60 585
R195 VTAIL.n59 VTAIL.n58 585
R196 VTAIL.n42 VTAIL.n41 585
R197 VTAIL.n53 VTAIL.n52 585
R198 VTAIL.n51 VTAIL.n50 585
R199 VTAIL.n46 VTAIL.n45 585
R200 VTAIL.n107 VTAIL.t11 327.856
R201 VTAIL.n11 VTAIL.t7 327.856
R202 VTAIL.n79 VTAIL.t1 327.856
R203 VTAIL.n47 VTAIL.t18 327.856
R204 VTAIL.n111 VTAIL.n105 171.744
R205 VTAIL.n112 VTAIL.n111 171.744
R206 VTAIL.n112 VTAIL.n101 171.744
R207 VTAIL.n119 VTAIL.n101 171.744
R208 VTAIL.n120 VTAIL.n119 171.744
R209 VTAIL.n15 VTAIL.n9 171.744
R210 VTAIL.n16 VTAIL.n15 171.744
R211 VTAIL.n16 VTAIL.n5 171.744
R212 VTAIL.n23 VTAIL.n5 171.744
R213 VTAIL.n24 VTAIL.n23 171.744
R214 VTAIL.n92 VTAIL.n91 171.744
R215 VTAIL.n91 VTAIL.n73 171.744
R216 VTAIL.n84 VTAIL.n73 171.744
R217 VTAIL.n84 VTAIL.n83 171.744
R218 VTAIL.n83 VTAIL.n77 171.744
R219 VTAIL.n60 VTAIL.n59 171.744
R220 VTAIL.n59 VTAIL.n41 171.744
R221 VTAIL.n52 VTAIL.n41 171.744
R222 VTAIL.n52 VTAIL.n51 171.744
R223 VTAIL.n51 VTAIL.n45 171.744
R224 VTAIL.t11 VTAIL.n105 85.8723
R225 VTAIL.t7 VTAIL.n9 85.8723
R226 VTAIL.t1 VTAIL.n77 85.8723
R227 VTAIL.t18 VTAIL.n45 85.8723
R228 VTAIL.n69 VTAIL.n68 81.234
R229 VTAIL.n67 VTAIL.n66 81.234
R230 VTAIL.n37 VTAIL.n36 81.234
R231 VTAIL.n35 VTAIL.n34 81.234
R232 VTAIL.n127 VTAIL.n126 81.2338
R233 VTAIL.n1 VTAIL.n0 81.2338
R234 VTAIL.n31 VTAIL.n30 81.2338
R235 VTAIL.n33 VTAIL.n32 81.2338
R236 VTAIL.n125 VTAIL.n124 32.7672
R237 VTAIL.n29 VTAIL.n28 32.7672
R238 VTAIL.n97 VTAIL.n96 32.7672
R239 VTAIL.n65 VTAIL.n64 32.7672
R240 VTAIL.n35 VTAIL.n33 23.8755
R241 VTAIL.n125 VTAIL.n97 20.41
R242 VTAIL.n107 VTAIL.n106 16.381
R243 VTAIL.n11 VTAIL.n10 16.381
R244 VTAIL.n79 VTAIL.n78 16.381
R245 VTAIL.n47 VTAIL.n46 16.381
R246 VTAIL.n110 VTAIL.n109 12.8005
R247 VTAIL.n14 VTAIL.n13 12.8005
R248 VTAIL.n82 VTAIL.n81 12.8005
R249 VTAIL.n50 VTAIL.n49 12.8005
R250 VTAIL.n113 VTAIL.n104 12.0247
R251 VTAIL.n17 VTAIL.n8 12.0247
R252 VTAIL.n85 VTAIL.n76 12.0247
R253 VTAIL.n53 VTAIL.n44 12.0247
R254 VTAIL.n114 VTAIL.n102 11.249
R255 VTAIL.n18 VTAIL.n6 11.249
R256 VTAIL.n86 VTAIL.n74 11.249
R257 VTAIL.n54 VTAIL.n42 11.249
R258 VTAIL.n118 VTAIL.n117 10.4732
R259 VTAIL.n22 VTAIL.n21 10.4732
R260 VTAIL.n90 VTAIL.n89 10.4732
R261 VTAIL.n58 VTAIL.n57 10.4732
R262 VTAIL.n121 VTAIL.n100 9.69747
R263 VTAIL.n25 VTAIL.n4 9.69747
R264 VTAIL.n93 VTAIL.n72 9.69747
R265 VTAIL.n61 VTAIL.n40 9.69747
R266 VTAIL.n124 VTAIL.n123 9.45567
R267 VTAIL.n28 VTAIL.n27 9.45567
R268 VTAIL.n96 VTAIL.n95 9.45567
R269 VTAIL.n64 VTAIL.n63 9.45567
R270 VTAIL.n123 VTAIL.n122 9.3005
R271 VTAIL.n100 VTAIL.n99 9.3005
R272 VTAIL.n117 VTAIL.n116 9.3005
R273 VTAIL.n115 VTAIL.n114 9.3005
R274 VTAIL.n104 VTAIL.n103 9.3005
R275 VTAIL.n109 VTAIL.n108 9.3005
R276 VTAIL.n27 VTAIL.n26 9.3005
R277 VTAIL.n4 VTAIL.n3 9.3005
R278 VTAIL.n21 VTAIL.n20 9.3005
R279 VTAIL.n19 VTAIL.n18 9.3005
R280 VTAIL.n8 VTAIL.n7 9.3005
R281 VTAIL.n13 VTAIL.n12 9.3005
R282 VTAIL.n95 VTAIL.n94 9.3005
R283 VTAIL.n72 VTAIL.n71 9.3005
R284 VTAIL.n89 VTAIL.n88 9.3005
R285 VTAIL.n87 VTAIL.n86 9.3005
R286 VTAIL.n76 VTAIL.n75 9.3005
R287 VTAIL.n81 VTAIL.n80 9.3005
R288 VTAIL.n63 VTAIL.n62 9.3005
R289 VTAIL.n40 VTAIL.n39 9.3005
R290 VTAIL.n57 VTAIL.n56 9.3005
R291 VTAIL.n55 VTAIL.n54 9.3005
R292 VTAIL.n44 VTAIL.n43 9.3005
R293 VTAIL.n49 VTAIL.n48 9.3005
R294 VTAIL.n122 VTAIL.n98 8.92171
R295 VTAIL.n26 VTAIL.n2 8.92171
R296 VTAIL.n94 VTAIL.n70 8.92171
R297 VTAIL.n62 VTAIL.n38 8.92171
R298 VTAIL.n126 VTAIL.t15 6.12197
R299 VTAIL.n126 VTAIL.t17 6.12197
R300 VTAIL.n0 VTAIL.t13 6.12197
R301 VTAIL.n0 VTAIL.t14 6.12197
R302 VTAIL.n30 VTAIL.t4 6.12197
R303 VTAIL.n30 VTAIL.t5 6.12197
R304 VTAIL.n32 VTAIL.t3 6.12197
R305 VTAIL.n32 VTAIL.t0 6.12197
R306 VTAIL.n68 VTAIL.t19 6.12197
R307 VTAIL.n68 VTAIL.t2 6.12197
R308 VTAIL.n66 VTAIL.t8 6.12197
R309 VTAIL.n66 VTAIL.t6 6.12197
R310 VTAIL.n36 VTAIL.t10 6.12197
R311 VTAIL.n36 VTAIL.t16 6.12197
R312 VTAIL.n34 VTAIL.t9 6.12197
R313 VTAIL.n34 VTAIL.t12 6.12197
R314 VTAIL.n124 VTAIL.n98 5.04292
R315 VTAIL.n28 VTAIL.n2 5.04292
R316 VTAIL.n96 VTAIL.n70 5.04292
R317 VTAIL.n64 VTAIL.n38 5.04292
R318 VTAIL.n122 VTAIL.n121 4.26717
R319 VTAIL.n26 VTAIL.n25 4.26717
R320 VTAIL.n94 VTAIL.n93 4.26717
R321 VTAIL.n62 VTAIL.n61 4.26717
R322 VTAIL.n80 VTAIL.n79 3.71853
R323 VTAIL.n48 VTAIL.n47 3.71853
R324 VTAIL.n108 VTAIL.n107 3.71853
R325 VTAIL.n12 VTAIL.n11 3.71853
R326 VTAIL.n118 VTAIL.n100 3.49141
R327 VTAIL.n22 VTAIL.n4 3.49141
R328 VTAIL.n90 VTAIL.n72 3.49141
R329 VTAIL.n58 VTAIL.n40 3.49141
R330 VTAIL.n37 VTAIL.n35 3.46602
R331 VTAIL.n65 VTAIL.n37 3.46602
R332 VTAIL.n69 VTAIL.n67 3.46602
R333 VTAIL.n97 VTAIL.n69 3.46602
R334 VTAIL.n33 VTAIL.n31 3.46602
R335 VTAIL.n31 VTAIL.n29 3.46602
R336 VTAIL.n127 VTAIL.n125 3.46602
R337 VTAIL.n117 VTAIL.n102 2.71565
R338 VTAIL.n21 VTAIL.n6 2.71565
R339 VTAIL.n89 VTAIL.n74 2.71565
R340 VTAIL.n57 VTAIL.n42 2.71565
R341 VTAIL VTAIL.n1 2.65783
R342 VTAIL.n67 VTAIL.n65 2.20309
R343 VTAIL.n29 VTAIL.n1 2.20309
R344 VTAIL.n114 VTAIL.n113 1.93989
R345 VTAIL.n18 VTAIL.n17 1.93989
R346 VTAIL.n86 VTAIL.n85 1.93989
R347 VTAIL.n54 VTAIL.n53 1.93989
R348 VTAIL.n110 VTAIL.n104 1.16414
R349 VTAIL.n14 VTAIL.n8 1.16414
R350 VTAIL.n82 VTAIL.n76 1.16414
R351 VTAIL.n50 VTAIL.n44 1.16414
R352 VTAIL VTAIL.n127 0.80869
R353 VTAIL.n109 VTAIL.n106 0.388379
R354 VTAIL.n13 VTAIL.n10 0.388379
R355 VTAIL.n81 VTAIL.n78 0.388379
R356 VTAIL.n49 VTAIL.n46 0.388379
R357 VTAIL.n108 VTAIL.n103 0.155672
R358 VTAIL.n115 VTAIL.n103 0.155672
R359 VTAIL.n116 VTAIL.n115 0.155672
R360 VTAIL.n116 VTAIL.n99 0.155672
R361 VTAIL.n123 VTAIL.n99 0.155672
R362 VTAIL.n12 VTAIL.n7 0.155672
R363 VTAIL.n19 VTAIL.n7 0.155672
R364 VTAIL.n20 VTAIL.n19 0.155672
R365 VTAIL.n20 VTAIL.n3 0.155672
R366 VTAIL.n27 VTAIL.n3 0.155672
R367 VTAIL.n95 VTAIL.n71 0.155672
R368 VTAIL.n88 VTAIL.n71 0.155672
R369 VTAIL.n88 VTAIL.n87 0.155672
R370 VTAIL.n87 VTAIL.n75 0.155672
R371 VTAIL.n80 VTAIL.n75 0.155672
R372 VTAIL.n63 VTAIL.n39 0.155672
R373 VTAIL.n56 VTAIL.n39 0.155672
R374 VTAIL.n56 VTAIL.n55 0.155672
R375 VTAIL.n55 VTAIL.n43 0.155672
R376 VTAIL.n48 VTAIL.n43 0.155672
R377 VDD2.n53 VDD2.n31 756.745
R378 VDD2.n22 VDD2.n0 756.745
R379 VDD2.n54 VDD2.n53 585
R380 VDD2.n52 VDD2.n51 585
R381 VDD2.n35 VDD2.n34 585
R382 VDD2.n46 VDD2.n45 585
R383 VDD2.n44 VDD2.n43 585
R384 VDD2.n39 VDD2.n38 585
R385 VDD2.n8 VDD2.n7 585
R386 VDD2.n13 VDD2.n12 585
R387 VDD2.n15 VDD2.n14 585
R388 VDD2.n4 VDD2.n3 585
R389 VDD2.n21 VDD2.n20 585
R390 VDD2.n23 VDD2.n22 585
R391 VDD2.n40 VDD2.t6 327.856
R392 VDD2.n9 VDD2.t9 327.856
R393 VDD2.n53 VDD2.n52 171.744
R394 VDD2.n52 VDD2.n34 171.744
R395 VDD2.n45 VDD2.n34 171.744
R396 VDD2.n45 VDD2.n44 171.744
R397 VDD2.n44 VDD2.n38 171.744
R398 VDD2.n13 VDD2.n7 171.744
R399 VDD2.n14 VDD2.n13 171.744
R400 VDD2.n14 VDD2.n3 171.744
R401 VDD2.n21 VDD2.n3 171.744
R402 VDD2.n22 VDD2.n21 171.744
R403 VDD2.n30 VDD2.n29 100.457
R404 VDD2 VDD2.n61 100.454
R405 VDD2.n60 VDD2.n59 97.9127
R406 VDD2.n28 VDD2.n27 97.9126
R407 VDD2.t6 VDD2.n38 85.8723
R408 VDD2.t9 VDD2.n7 85.8723
R409 VDD2.n28 VDD2.n26 52.9115
R410 VDD2.n58 VDD2.n57 49.446
R411 VDD2.n58 VDD2.n30 44.7541
R412 VDD2.n40 VDD2.n39 16.381
R413 VDD2.n9 VDD2.n8 16.381
R414 VDD2.n43 VDD2.n42 12.8005
R415 VDD2.n12 VDD2.n11 12.8005
R416 VDD2.n46 VDD2.n37 12.0247
R417 VDD2.n15 VDD2.n6 12.0247
R418 VDD2.n47 VDD2.n35 11.249
R419 VDD2.n16 VDD2.n4 11.249
R420 VDD2.n51 VDD2.n50 10.4732
R421 VDD2.n20 VDD2.n19 10.4732
R422 VDD2.n54 VDD2.n33 9.69747
R423 VDD2.n23 VDD2.n2 9.69747
R424 VDD2.n57 VDD2.n56 9.45567
R425 VDD2.n26 VDD2.n25 9.45567
R426 VDD2.n56 VDD2.n55 9.3005
R427 VDD2.n33 VDD2.n32 9.3005
R428 VDD2.n50 VDD2.n49 9.3005
R429 VDD2.n48 VDD2.n47 9.3005
R430 VDD2.n37 VDD2.n36 9.3005
R431 VDD2.n42 VDD2.n41 9.3005
R432 VDD2.n25 VDD2.n24 9.3005
R433 VDD2.n2 VDD2.n1 9.3005
R434 VDD2.n19 VDD2.n18 9.3005
R435 VDD2.n17 VDD2.n16 9.3005
R436 VDD2.n6 VDD2.n5 9.3005
R437 VDD2.n11 VDD2.n10 9.3005
R438 VDD2.n55 VDD2.n31 8.92171
R439 VDD2.n24 VDD2.n0 8.92171
R440 VDD2.n61 VDD2.t2 6.12197
R441 VDD2.n61 VDD2.t5 6.12197
R442 VDD2.n59 VDD2.t7 6.12197
R443 VDD2.n59 VDD2.t8 6.12197
R444 VDD2.n29 VDD2.t3 6.12197
R445 VDD2.n29 VDD2.t4 6.12197
R446 VDD2.n27 VDD2.t0 6.12197
R447 VDD2.n27 VDD2.t1 6.12197
R448 VDD2.n57 VDD2.n31 5.04292
R449 VDD2.n26 VDD2.n0 5.04292
R450 VDD2.n55 VDD2.n54 4.26717
R451 VDD2.n24 VDD2.n23 4.26717
R452 VDD2.n41 VDD2.n40 3.71853
R453 VDD2.n10 VDD2.n9 3.71853
R454 VDD2.n51 VDD2.n33 3.49141
R455 VDD2.n20 VDD2.n2 3.49141
R456 VDD2.n60 VDD2.n58 3.46602
R457 VDD2.n50 VDD2.n35 2.71565
R458 VDD2.n19 VDD2.n4 2.71565
R459 VDD2.n47 VDD2.n46 1.93989
R460 VDD2.n16 VDD2.n15 1.93989
R461 VDD2.n43 VDD2.n37 1.16414
R462 VDD2.n12 VDD2.n6 1.16414
R463 VDD2 VDD2.n60 0.925069
R464 VDD2.n30 VDD2.n28 0.811533
R465 VDD2.n42 VDD2.n39 0.388379
R466 VDD2.n11 VDD2.n8 0.388379
R467 VDD2.n56 VDD2.n32 0.155672
R468 VDD2.n49 VDD2.n32 0.155672
R469 VDD2.n49 VDD2.n48 0.155672
R470 VDD2.n48 VDD2.n36 0.155672
R471 VDD2.n41 VDD2.n36 0.155672
R472 VDD2.n10 VDD2.n5 0.155672
R473 VDD2.n17 VDD2.n5 0.155672
R474 VDD2.n18 VDD2.n17 0.155672
R475 VDD2.n18 VDD2.n1 0.155672
R476 VDD2.n25 VDD2.n1 0.155672
R477 B.n660 B.n659 585
R478 B.n661 B.n72 585
R479 B.n663 B.n662 585
R480 B.n664 B.n71 585
R481 B.n666 B.n665 585
R482 B.n667 B.n70 585
R483 B.n669 B.n668 585
R484 B.n670 B.n69 585
R485 B.n672 B.n671 585
R486 B.n673 B.n68 585
R487 B.n675 B.n674 585
R488 B.n676 B.n67 585
R489 B.n678 B.n677 585
R490 B.n679 B.n66 585
R491 B.n681 B.n680 585
R492 B.n682 B.n65 585
R493 B.n684 B.n683 585
R494 B.n685 B.n64 585
R495 B.n687 B.n686 585
R496 B.n688 B.n63 585
R497 B.n690 B.n689 585
R498 B.n691 B.n60 585
R499 B.n694 B.n693 585
R500 B.n695 B.n59 585
R501 B.n697 B.n696 585
R502 B.n698 B.n58 585
R503 B.n700 B.n699 585
R504 B.n701 B.n57 585
R505 B.n703 B.n702 585
R506 B.n704 B.n53 585
R507 B.n706 B.n705 585
R508 B.n707 B.n52 585
R509 B.n709 B.n708 585
R510 B.n710 B.n51 585
R511 B.n712 B.n711 585
R512 B.n713 B.n50 585
R513 B.n715 B.n714 585
R514 B.n716 B.n49 585
R515 B.n718 B.n717 585
R516 B.n719 B.n48 585
R517 B.n721 B.n720 585
R518 B.n722 B.n47 585
R519 B.n724 B.n723 585
R520 B.n725 B.n46 585
R521 B.n727 B.n726 585
R522 B.n728 B.n45 585
R523 B.n730 B.n729 585
R524 B.n731 B.n44 585
R525 B.n733 B.n732 585
R526 B.n734 B.n43 585
R527 B.n736 B.n735 585
R528 B.n737 B.n42 585
R529 B.n739 B.n738 585
R530 B.n658 B.n73 585
R531 B.n657 B.n656 585
R532 B.n655 B.n74 585
R533 B.n654 B.n653 585
R534 B.n652 B.n75 585
R535 B.n651 B.n650 585
R536 B.n649 B.n76 585
R537 B.n648 B.n647 585
R538 B.n646 B.n77 585
R539 B.n645 B.n644 585
R540 B.n643 B.n78 585
R541 B.n642 B.n641 585
R542 B.n640 B.n79 585
R543 B.n639 B.n638 585
R544 B.n637 B.n80 585
R545 B.n636 B.n635 585
R546 B.n634 B.n81 585
R547 B.n633 B.n632 585
R548 B.n631 B.n82 585
R549 B.n630 B.n629 585
R550 B.n628 B.n83 585
R551 B.n627 B.n626 585
R552 B.n625 B.n84 585
R553 B.n624 B.n623 585
R554 B.n622 B.n85 585
R555 B.n621 B.n620 585
R556 B.n619 B.n86 585
R557 B.n618 B.n617 585
R558 B.n616 B.n87 585
R559 B.n615 B.n614 585
R560 B.n613 B.n88 585
R561 B.n612 B.n611 585
R562 B.n610 B.n89 585
R563 B.n609 B.n608 585
R564 B.n607 B.n90 585
R565 B.n606 B.n605 585
R566 B.n604 B.n91 585
R567 B.n603 B.n602 585
R568 B.n601 B.n92 585
R569 B.n600 B.n599 585
R570 B.n598 B.n93 585
R571 B.n597 B.n596 585
R572 B.n595 B.n94 585
R573 B.n594 B.n593 585
R574 B.n592 B.n95 585
R575 B.n591 B.n590 585
R576 B.n589 B.n96 585
R577 B.n588 B.n587 585
R578 B.n586 B.n97 585
R579 B.n585 B.n584 585
R580 B.n583 B.n98 585
R581 B.n582 B.n581 585
R582 B.n580 B.n99 585
R583 B.n579 B.n578 585
R584 B.n577 B.n100 585
R585 B.n576 B.n575 585
R586 B.n574 B.n101 585
R587 B.n573 B.n572 585
R588 B.n571 B.n102 585
R589 B.n570 B.n569 585
R590 B.n568 B.n103 585
R591 B.n567 B.n566 585
R592 B.n565 B.n104 585
R593 B.n564 B.n563 585
R594 B.n562 B.n105 585
R595 B.n561 B.n560 585
R596 B.n559 B.n106 585
R597 B.n558 B.n557 585
R598 B.n556 B.n107 585
R599 B.n555 B.n554 585
R600 B.n553 B.n108 585
R601 B.n552 B.n551 585
R602 B.n550 B.n109 585
R603 B.n549 B.n548 585
R604 B.n547 B.n110 585
R605 B.n546 B.n545 585
R606 B.n544 B.n111 585
R607 B.n543 B.n542 585
R608 B.n541 B.n112 585
R609 B.n540 B.n539 585
R610 B.n538 B.n113 585
R611 B.n537 B.n536 585
R612 B.n535 B.n114 585
R613 B.n534 B.n533 585
R614 B.n532 B.n115 585
R615 B.n531 B.n530 585
R616 B.n529 B.n116 585
R617 B.n528 B.n527 585
R618 B.n526 B.n117 585
R619 B.n525 B.n524 585
R620 B.n523 B.n118 585
R621 B.n522 B.n521 585
R622 B.n520 B.n119 585
R623 B.n519 B.n518 585
R624 B.n517 B.n120 585
R625 B.n516 B.n515 585
R626 B.n514 B.n121 585
R627 B.n513 B.n512 585
R628 B.n511 B.n122 585
R629 B.n510 B.n509 585
R630 B.n508 B.n123 585
R631 B.n507 B.n506 585
R632 B.n505 B.n124 585
R633 B.n504 B.n503 585
R634 B.n502 B.n125 585
R635 B.n501 B.n500 585
R636 B.n499 B.n126 585
R637 B.n498 B.n497 585
R638 B.n496 B.n127 585
R639 B.n495 B.n494 585
R640 B.n493 B.n128 585
R641 B.n492 B.n491 585
R642 B.n490 B.n129 585
R643 B.n489 B.n488 585
R644 B.n487 B.n130 585
R645 B.n486 B.n485 585
R646 B.n484 B.n131 585
R647 B.n483 B.n482 585
R648 B.n481 B.n132 585
R649 B.n480 B.n479 585
R650 B.n478 B.n133 585
R651 B.n477 B.n476 585
R652 B.n475 B.n134 585
R653 B.n474 B.n473 585
R654 B.n472 B.n135 585
R655 B.n471 B.n470 585
R656 B.n469 B.n136 585
R657 B.n468 B.n467 585
R658 B.n466 B.n137 585
R659 B.n465 B.n464 585
R660 B.n463 B.n138 585
R661 B.n462 B.n461 585
R662 B.n460 B.n139 585
R663 B.n459 B.n458 585
R664 B.n457 B.n140 585
R665 B.n456 B.n455 585
R666 B.n454 B.n141 585
R667 B.n453 B.n452 585
R668 B.n451 B.n142 585
R669 B.n450 B.n449 585
R670 B.n448 B.n143 585
R671 B.n447 B.n446 585
R672 B.n445 B.n144 585
R673 B.n444 B.n443 585
R674 B.n442 B.n145 585
R675 B.n441 B.n440 585
R676 B.n439 B.n146 585
R677 B.n438 B.n437 585
R678 B.n436 B.n147 585
R679 B.n435 B.n434 585
R680 B.n433 B.n148 585
R681 B.n432 B.n431 585
R682 B.n430 B.n149 585
R683 B.n429 B.n428 585
R684 B.n427 B.n150 585
R685 B.n426 B.n425 585
R686 B.n424 B.n151 585
R687 B.n423 B.n422 585
R688 B.n421 B.n152 585
R689 B.n338 B.n337 585
R690 B.n339 B.n180 585
R691 B.n341 B.n340 585
R692 B.n342 B.n179 585
R693 B.n344 B.n343 585
R694 B.n345 B.n178 585
R695 B.n347 B.n346 585
R696 B.n348 B.n177 585
R697 B.n350 B.n349 585
R698 B.n351 B.n176 585
R699 B.n353 B.n352 585
R700 B.n354 B.n175 585
R701 B.n356 B.n355 585
R702 B.n357 B.n174 585
R703 B.n359 B.n358 585
R704 B.n360 B.n173 585
R705 B.n362 B.n361 585
R706 B.n363 B.n172 585
R707 B.n365 B.n364 585
R708 B.n366 B.n171 585
R709 B.n368 B.n367 585
R710 B.n369 B.n168 585
R711 B.n372 B.n371 585
R712 B.n373 B.n167 585
R713 B.n375 B.n374 585
R714 B.n376 B.n166 585
R715 B.n378 B.n377 585
R716 B.n379 B.n165 585
R717 B.n381 B.n380 585
R718 B.n382 B.n164 585
R719 B.n387 B.n386 585
R720 B.n388 B.n163 585
R721 B.n390 B.n389 585
R722 B.n391 B.n162 585
R723 B.n393 B.n392 585
R724 B.n394 B.n161 585
R725 B.n396 B.n395 585
R726 B.n397 B.n160 585
R727 B.n399 B.n398 585
R728 B.n400 B.n159 585
R729 B.n402 B.n401 585
R730 B.n403 B.n158 585
R731 B.n405 B.n404 585
R732 B.n406 B.n157 585
R733 B.n408 B.n407 585
R734 B.n409 B.n156 585
R735 B.n411 B.n410 585
R736 B.n412 B.n155 585
R737 B.n414 B.n413 585
R738 B.n415 B.n154 585
R739 B.n417 B.n416 585
R740 B.n418 B.n153 585
R741 B.n420 B.n419 585
R742 B.n336 B.n181 585
R743 B.n335 B.n334 585
R744 B.n333 B.n182 585
R745 B.n332 B.n331 585
R746 B.n330 B.n183 585
R747 B.n329 B.n328 585
R748 B.n327 B.n184 585
R749 B.n326 B.n325 585
R750 B.n324 B.n185 585
R751 B.n323 B.n322 585
R752 B.n321 B.n186 585
R753 B.n320 B.n319 585
R754 B.n318 B.n187 585
R755 B.n317 B.n316 585
R756 B.n315 B.n188 585
R757 B.n314 B.n313 585
R758 B.n312 B.n189 585
R759 B.n311 B.n310 585
R760 B.n309 B.n190 585
R761 B.n308 B.n307 585
R762 B.n306 B.n191 585
R763 B.n305 B.n304 585
R764 B.n303 B.n192 585
R765 B.n302 B.n301 585
R766 B.n300 B.n193 585
R767 B.n299 B.n298 585
R768 B.n297 B.n194 585
R769 B.n296 B.n295 585
R770 B.n294 B.n195 585
R771 B.n293 B.n292 585
R772 B.n291 B.n196 585
R773 B.n290 B.n289 585
R774 B.n288 B.n197 585
R775 B.n287 B.n286 585
R776 B.n285 B.n198 585
R777 B.n284 B.n283 585
R778 B.n282 B.n199 585
R779 B.n281 B.n280 585
R780 B.n279 B.n200 585
R781 B.n278 B.n277 585
R782 B.n276 B.n201 585
R783 B.n275 B.n274 585
R784 B.n273 B.n202 585
R785 B.n272 B.n271 585
R786 B.n270 B.n203 585
R787 B.n269 B.n268 585
R788 B.n267 B.n204 585
R789 B.n266 B.n265 585
R790 B.n264 B.n205 585
R791 B.n263 B.n262 585
R792 B.n261 B.n206 585
R793 B.n260 B.n259 585
R794 B.n258 B.n207 585
R795 B.n257 B.n256 585
R796 B.n255 B.n208 585
R797 B.n254 B.n253 585
R798 B.n252 B.n209 585
R799 B.n251 B.n250 585
R800 B.n249 B.n210 585
R801 B.n248 B.n247 585
R802 B.n246 B.n211 585
R803 B.n245 B.n244 585
R804 B.n243 B.n212 585
R805 B.n242 B.n241 585
R806 B.n240 B.n213 585
R807 B.n239 B.n238 585
R808 B.n237 B.n214 585
R809 B.n236 B.n235 585
R810 B.n234 B.n215 585
R811 B.n233 B.n232 585
R812 B.n231 B.n216 585
R813 B.n230 B.n229 585
R814 B.n228 B.n217 585
R815 B.n227 B.n226 585
R816 B.n225 B.n218 585
R817 B.n224 B.n223 585
R818 B.n222 B.n219 585
R819 B.n221 B.n220 585
R820 B.n2 B.n0 585
R821 B.n857 B.n1 585
R822 B.n856 B.n855 585
R823 B.n854 B.n3 585
R824 B.n853 B.n852 585
R825 B.n851 B.n4 585
R826 B.n850 B.n849 585
R827 B.n848 B.n5 585
R828 B.n847 B.n846 585
R829 B.n845 B.n6 585
R830 B.n844 B.n843 585
R831 B.n842 B.n7 585
R832 B.n841 B.n840 585
R833 B.n839 B.n8 585
R834 B.n838 B.n837 585
R835 B.n836 B.n9 585
R836 B.n835 B.n834 585
R837 B.n833 B.n10 585
R838 B.n832 B.n831 585
R839 B.n830 B.n11 585
R840 B.n829 B.n828 585
R841 B.n827 B.n12 585
R842 B.n826 B.n825 585
R843 B.n824 B.n13 585
R844 B.n823 B.n822 585
R845 B.n821 B.n14 585
R846 B.n820 B.n819 585
R847 B.n818 B.n15 585
R848 B.n817 B.n816 585
R849 B.n815 B.n16 585
R850 B.n814 B.n813 585
R851 B.n812 B.n17 585
R852 B.n811 B.n810 585
R853 B.n809 B.n18 585
R854 B.n808 B.n807 585
R855 B.n806 B.n19 585
R856 B.n805 B.n804 585
R857 B.n803 B.n20 585
R858 B.n802 B.n801 585
R859 B.n800 B.n21 585
R860 B.n799 B.n798 585
R861 B.n797 B.n22 585
R862 B.n796 B.n795 585
R863 B.n794 B.n23 585
R864 B.n793 B.n792 585
R865 B.n791 B.n24 585
R866 B.n790 B.n789 585
R867 B.n788 B.n25 585
R868 B.n787 B.n786 585
R869 B.n785 B.n26 585
R870 B.n784 B.n783 585
R871 B.n782 B.n27 585
R872 B.n781 B.n780 585
R873 B.n779 B.n28 585
R874 B.n778 B.n777 585
R875 B.n776 B.n29 585
R876 B.n775 B.n774 585
R877 B.n773 B.n30 585
R878 B.n772 B.n771 585
R879 B.n770 B.n31 585
R880 B.n769 B.n768 585
R881 B.n767 B.n32 585
R882 B.n766 B.n765 585
R883 B.n764 B.n33 585
R884 B.n763 B.n762 585
R885 B.n761 B.n34 585
R886 B.n760 B.n759 585
R887 B.n758 B.n35 585
R888 B.n757 B.n756 585
R889 B.n755 B.n36 585
R890 B.n754 B.n753 585
R891 B.n752 B.n37 585
R892 B.n751 B.n750 585
R893 B.n749 B.n38 585
R894 B.n748 B.n747 585
R895 B.n746 B.n39 585
R896 B.n745 B.n744 585
R897 B.n743 B.n40 585
R898 B.n742 B.n741 585
R899 B.n740 B.n41 585
R900 B.n859 B.n858 585
R901 B.n337 B.n336 545.355
R902 B.n738 B.n41 545.355
R903 B.n419 B.n152 545.355
R904 B.n659 B.n658 545.355
R905 B.n383 B.t2 334.193
R906 B.n61 B.t7 334.193
R907 B.n169 B.t5 334.193
R908 B.n54 B.t10 334.193
R909 B.n384 B.t1 256.231
R910 B.n62 B.t8 256.231
R911 B.n170 B.t4 256.231
R912 B.n55 B.t11 256.231
R913 B.n383 B.t0 243.936
R914 B.n169 B.t3 243.936
R915 B.n54 B.t9 243.936
R916 B.n61 B.t6 243.936
R917 B.n336 B.n335 163.367
R918 B.n335 B.n182 163.367
R919 B.n331 B.n182 163.367
R920 B.n331 B.n330 163.367
R921 B.n330 B.n329 163.367
R922 B.n329 B.n184 163.367
R923 B.n325 B.n184 163.367
R924 B.n325 B.n324 163.367
R925 B.n324 B.n323 163.367
R926 B.n323 B.n186 163.367
R927 B.n319 B.n186 163.367
R928 B.n319 B.n318 163.367
R929 B.n318 B.n317 163.367
R930 B.n317 B.n188 163.367
R931 B.n313 B.n188 163.367
R932 B.n313 B.n312 163.367
R933 B.n312 B.n311 163.367
R934 B.n311 B.n190 163.367
R935 B.n307 B.n190 163.367
R936 B.n307 B.n306 163.367
R937 B.n306 B.n305 163.367
R938 B.n305 B.n192 163.367
R939 B.n301 B.n192 163.367
R940 B.n301 B.n300 163.367
R941 B.n300 B.n299 163.367
R942 B.n299 B.n194 163.367
R943 B.n295 B.n194 163.367
R944 B.n295 B.n294 163.367
R945 B.n294 B.n293 163.367
R946 B.n293 B.n196 163.367
R947 B.n289 B.n196 163.367
R948 B.n289 B.n288 163.367
R949 B.n288 B.n287 163.367
R950 B.n287 B.n198 163.367
R951 B.n283 B.n198 163.367
R952 B.n283 B.n282 163.367
R953 B.n282 B.n281 163.367
R954 B.n281 B.n200 163.367
R955 B.n277 B.n200 163.367
R956 B.n277 B.n276 163.367
R957 B.n276 B.n275 163.367
R958 B.n275 B.n202 163.367
R959 B.n271 B.n202 163.367
R960 B.n271 B.n270 163.367
R961 B.n270 B.n269 163.367
R962 B.n269 B.n204 163.367
R963 B.n265 B.n204 163.367
R964 B.n265 B.n264 163.367
R965 B.n264 B.n263 163.367
R966 B.n263 B.n206 163.367
R967 B.n259 B.n206 163.367
R968 B.n259 B.n258 163.367
R969 B.n258 B.n257 163.367
R970 B.n257 B.n208 163.367
R971 B.n253 B.n208 163.367
R972 B.n253 B.n252 163.367
R973 B.n252 B.n251 163.367
R974 B.n251 B.n210 163.367
R975 B.n247 B.n210 163.367
R976 B.n247 B.n246 163.367
R977 B.n246 B.n245 163.367
R978 B.n245 B.n212 163.367
R979 B.n241 B.n212 163.367
R980 B.n241 B.n240 163.367
R981 B.n240 B.n239 163.367
R982 B.n239 B.n214 163.367
R983 B.n235 B.n214 163.367
R984 B.n235 B.n234 163.367
R985 B.n234 B.n233 163.367
R986 B.n233 B.n216 163.367
R987 B.n229 B.n216 163.367
R988 B.n229 B.n228 163.367
R989 B.n228 B.n227 163.367
R990 B.n227 B.n218 163.367
R991 B.n223 B.n218 163.367
R992 B.n223 B.n222 163.367
R993 B.n222 B.n221 163.367
R994 B.n221 B.n2 163.367
R995 B.n858 B.n2 163.367
R996 B.n858 B.n857 163.367
R997 B.n857 B.n856 163.367
R998 B.n856 B.n3 163.367
R999 B.n852 B.n3 163.367
R1000 B.n852 B.n851 163.367
R1001 B.n851 B.n850 163.367
R1002 B.n850 B.n5 163.367
R1003 B.n846 B.n5 163.367
R1004 B.n846 B.n845 163.367
R1005 B.n845 B.n844 163.367
R1006 B.n844 B.n7 163.367
R1007 B.n840 B.n7 163.367
R1008 B.n840 B.n839 163.367
R1009 B.n839 B.n838 163.367
R1010 B.n838 B.n9 163.367
R1011 B.n834 B.n9 163.367
R1012 B.n834 B.n833 163.367
R1013 B.n833 B.n832 163.367
R1014 B.n832 B.n11 163.367
R1015 B.n828 B.n11 163.367
R1016 B.n828 B.n827 163.367
R1017 B.n827 B.n826 163.367
R1018 B.n826 B.n13 163.367
R1019 B.n822 B.n13 163.367
R1020 B.n822 B.n821 163.367
R1021 B.n821 B.n820 163.367
R1022 B.n820 B.n15 163.367
R1023 B.n816 B.n15 163.367
R1024 B.n816 B.n815 163.367
R1025 B.n815 B.n814 163.367
R1026 B.n814 B.n17 163.367
R1027 B.n810 B.n17 163.367
R1028 B.n810 B.n809 163.367
R1029 B.n809 B.n808 163.367
R1030 B.n808 B.n19 163.367
R1031 B.n804 B.n19 163.367
R1032 B.n804 B.n803 163.367
R1033 B.n803 B.n802 163.367
R1034 B.n802 B.n21 163.367
R1035 B.n798 B.n21 163.367
R1036 B.n798 B.n797 163.367
R1037 B.n797 B.n796 163.367
R1038 B.n796 B.n23 163.367
R1039 B.n792 B.n23 163.367
R1040 B.n792 B.n791 163.367
R1041 B.n791 B.n790 163.367
R1042 B.n790 B.n25 163.367
R1043 B.n786 B.n25 163.367
R1044 B.n786 B.n785 163.367
R1045 B.n785 B.n784 163.367
R1046 B.n784 B.n27 163.367
R1047 B.n780 B.n27 163.367
R1048 B.n780 B.n779 163.367
R1049 B.n779 B.n778 163.367
R1050 B.n778 B.n29 163.367
R1051 B.n774 B.n29 163.367
R1052 B.n774 B.n773 163.367
R1053 B.n773 B.n772 163.367
R1054 B.n772 B.n31 163.367
R1055 B.n768 B.n31 163.367
R1056 B.n768 B.n767 163.367
R1057 B.n767 B.n766 163.367
R1058 B.n766 B.n33 163.367
R1059 B.n762 B.n33 163.367
R1060 B.n762 B.n761 163.367
R1061 B.n761 B.n760 163.367
R1062 B.n760 B.n35 163.367
R1063 B.n756 B.n35 163.367
R1064 B.n756 B.n755 163.367
R1065 B.n755 B.n754 163.367
R1066 B.n754 B.n37 163.367
R1067 B.n750 B.n37 163.367
R1068 B.n750 B.n749 163.367
R1069 B.n749 B.n748 163.367
R1070 B.n748 B.n39 163.367
R1071 B.n744 B.n39 163.367
R1072 B.n744 B.n743 163.367
R1073 B.n743 B.n742 163.367
R1074 B.n742 B.n41 163.367
R1075 B.n337 B.n180 163.367
R1076 B.n341 B.n180 163.367
R1077 B.n342 B.n341 163.367
R1078 B.n343 B.n342 163.367
R1079 B.n343 B.n178 163.367
R1080 B.n347 B.n178 163.367
R1081 B.n348 B.n347 163.367
R1082 B.n349 B.n348 163.367
R1083 B.n349 B.n176 163.367
R1084 B.n353 B.n176 163.367
R1085 B.n354 B.n353 163.367
R1086 B.n355 B.n354 163.367
R1087 B.n355 B.n174 163.367
R1088 B.n359 B.n174 163.367
R1089 B.n360 B.n359 163.367
R1090 B.n361 B.n360 163.367
R1091 B.n361 B.n172 163.367
R1092 B.n365 B.n172 163.367
R1093 B.n366 B.n365 163.367
R1094 B.n367 B.n366 163.367
R1095 B.n367 B.n168 163.367
R1096 B.n372 B.n168 163.367
R1097 B.n373 B.n372 163.367
R1098 B.n374 B.n373 163.367
R1099 B.n374 B.n166 163.367
R1100 B.n378 B.n166 163.367
R1101 B.n379 B.n378 163.367
R1102 B.n380 B.n379 163.367
R1103 B.n380 B.n164 163.367
R1104 B.n387 B.n164 163.367
R1105 B.n388 B.n387 163.367
R1106 B.n389 B.n388 163.367
R1107 B.n389 B.n162 163.367
R1108 B.n393 B.n162 163.367
R1109 B.n394 B.n393 163.367
R1110 B.n395 B.n394 163.367
R1111 B.n395 B.n160 163.367
R1112 B.n399 B.n160 163.367
R1113 B.n400 B.n399 163.367
R1114 B.n401 B.n400 163.367
R1115 B.n401 B.n158 163.367
R1116 B.n405 B.n158 163.367
R1117 B.n406 B.n405 163.367
R1118 B.n407 B.n406 163.367
R1119 B.n407 B.n156 163.367
R1120 B.n411 B.n156 163.367
R1121 B.n412 B.n411 163.367
R1122 B.n413 B.n412 163.367
R1123 B.n413 B.n154 163.367
R1124 B.n417 B.n154 163.367
R1125 B.n418 B.n417 163.367
R1126 B.n419 B.n418 163.367
R1127 B.n423 B.n152 163.367
R1128 B.n424 B.n423 163.367
R1129 B.n425 B.n424 163.367
R1130 B.n425 B.n150 163.367
R1131 B.n429 B.n150 163.367
R1132 B.n430 B.n429 163.367
R1133 B.n431 B.n430 163.367
R1134 B.n431 B.n148 163.367
R1135 B.n435 B.n148 163.367
R1136 B.n436 B.n435 163.367
R1137 B.n437 B.n436 163.367
R1138 B.n437 B.n146 163.367
R1139 B.n441 B.n146 163.367
R1140 B.n442 B.n441 163.367
R1141 B.n443 B.n442 163.367
R1142 B.n443 B.n144 163.367
R1143 B.n447 B.n144 163.367
R1144 B.n448 B.n447 163.367
R1145 B.n449 B.n448 163.367
R1146 B.n449 B.n142 163.367
R1147 B.n453 B.n142 163.367
R1148 B.n454 B.n453 163.367
R1149 B.n455 B.n454 163.367
R1150 B.n455 B.n140 163.367
R1151 B.n459 B.n140 163.367
R1152 B.n460 B.n459 163.367
R1153 B.n461 B.n460 163.367
R1154 B.n461 B.n138 163.367
R1155 B.n465 B.n138 163.367
R1156 B.n466 B.n465 163.367
R1157 B.n467 B.n466 163.367
R1158 B.n467 B.n136 163.367
R1159 B.n471 B.n136 163.367
R1160 B.n472 B.n471 163.367
R1161 B.n473 B.n472 163.367
R1162 B.n473 B.n134 163.367
R1163 B.n477 B.n134 163.367
R1164 B.n478 B.n477 163.367
R1165 B.n479 B.n478 163.367
R1166 B.n479 B.n132 163.367
R1167 B.n483 B.n132 163.367
R1168 B.n484 B.n483 163.367
R1169 B.n485 B.n484 163.367
R1170 B.n485 B.n130 163.367
R1171 B.n489 B.n130 163.367
R1172 B.n490 B.n489 163.367
R1173 B.n491 B.n490 163.367
R1174 B.n491 B.n128 163.367
R1175 B.n495 B.n128 163.367
R1176 B.n496 B.n495 163.367
R1177 B.n497 B.n496 163.367
R1178 B.n497 B.n126 163.367
R1179 B.n501 B.n126 163.367
R1180 B.n502 B.n501 163.367
R1181 B.n503 B.n502 163.367
R1182 B.n503 B.n124 163.367
R1183 B.n507 B.n124 163.367
R1184 B.n508 B.n507 163.367
R1185 B.n509 B.n508 163.367
R1186 B.n509 B.n122 163.367
R1187 B.n513 B.n122 163.367
R1188 B.n514 B.n513 163.367
R1189 B.n515 B.n514 163.367
R1190 B.n515 B.n120 163.367
R1191 B.n519 B.n120 163.367
R1192 B.n520 B.n519 163.367
R1193 B.n521 B.n520 163.367
R1194 B.n521 B.n118 163.367
R1195 B.n525 B.n118 163.367
R1196 B.n526 B.n525 163.367
R1197 B.n527 B.n526 163.367
R1198 B.n527 B.n116 163.367
R1199 B.n531 B.n116 163.367
R1200 B.n532 B.n531 163.367
R1201 B.n533 B.n532 163.367
R1202 B.n533 B.n114 163.367
R1203 B.n537 B.n114 163.367
R1204 B.n538 B.n537 163.367
R1205 B.n539 B.n538 163.367
R1206 B.n539 B.n112 163.367
R1207 B.n543 B.n112 163.367
R1208 B.n544 B.n543 163.367
R1209 B.n545 B.n544 163.367
R1210 B.n545 B.n110 163.367
R1211 B.n549 B.n110 163.367
R1212 B.n550 B.n549 163.367
R1213 B.n551 B.n550 163.367
R1214 B.n551 B.n108 163.367
R1215 B.n555 B.n108 163.367
R1216 B.n556 B.n555 163.367
R1217 B.n557 B.n556 163.367
R1218 B.n557 B.n106 163.367
R1219 B.n561 B.n106 163.367
R1220 B.n562 B.n561 163.367
R1221 B.n563 B.n562 163.367
R1222 B.n563 B.n104 163.367
R1223 B.n567 B.n104 163.367
R1224 B.n568 B.n567 163.367
R1225 B.n569 B.n568 163.367
R1226 B.n569 B.n102 163.367
R1227 B.n573 B.n102 163.367
R1228 B.n574 B.n573 163.367
R1229 B.n575 B.n574 163.367
R1230 B.n575 B.n100 163.367
R1231 B.n579 B.n100 163.367
R1232 B.n580 B.n579 163.367
R1233 B.n581 B.n580 163.367
R1234 B.n581 B.n98 163.367
R1235 B.n585 B.n98 163.367
R1236 B.n586 B.n585 163.367
R1237 B.n587 B.n586 163.367
R1238 B.n587 B.n96 163.367
R1239 B.n591 B.n96 163.367
R1240 B.n592 B.n591 163.367
R1241 B.n593 B.n592 163.367
R1242 B.n593 B.n94 163.367
R1243 B.n597 B.n94 163.367
R1244 B.n598 B.n597 163.367
R1245 B.n599 B.n598 163.367
R1246 B.n599 B.n92 163.367
R1247 B.n603 B.n92 163.367
R1248 B.n604 B.n603 163.367
R1249 B.n605 B.n604 163.367
R1250 B.n605 B.n90 163.367
R1251 B.n609 B.n90 163.367
R1252 B.n610 B.n609 163.367
R1253 B.n611 B.n610 163.367
R1254 B.n611 B.n88 163.367
R1255 B.n615 B.n88 163.367
R1256 B.n616 B.n615 163.367
R1257 B.n617 B.n616 163.367
R1258 B.n617 B.n86 163.367
R1259 B.n621 B.n86 163.367
R1260 B.n622 B.n621 163.367
R1261 B.n623 B.n622 163.367
R1262 B.n623 B.n84 163.367
R1263 B.n627 B.n84 163.367
R1264 B.n628 B.n627 163.367
R1265 B.n629 B.n628 163.367
R1266 B.n629 B.n82 163.367
R1267 B.n633 B.n82 163.367
R1268 B.n634 B.n633 163.367
R1269 B.n635 B.n634 163.367
R1270 B.n635 B.n80 163.367
R1271 B.n639 B.n80 163.367
R1272 B.n640 B.n639 163.367
R1273 B.n641 B.n640 163.367
R1274 B.n641 B.n78 163.367
R1275 B.n645 B.n78 163.367
R1276 B.n646 B.n645 163.367
R1277 B.n647 B.n646 163.367
R1278 B.n647 B.n76 163.367
R1279 B.n651 B.n76 163.367
R1280 B.n652 B.n651 163.367
R1281 B.n653 B.n652 163.367
R1282 B.n653 B.n74 163.367
R1283 B.n657 B.n74 163.367
R1284 B.n658 B.n657 163.367
R1285 B.n738 B.n737 163.367
R1286 B.n737 B.n736 163.367
R1287 B.n736 B.n43 163.367
R1288 B.n732 B.n43 163.367
R1289 B.n732 B.n731 163.367
R1290 B.n731 B.n730 163.367
R1291 B.n730 B.n45 163.367
R1292 B.n726 B.n45 163.367
R1293 B.n726 B.n725 163.367
R1294 B.n725 B.n724 163.367
R1295 B.n724 B.n47 163.367
R1296 B.n720 B.n47 163.367
R1297 B.n720 B.n719 163.367
R1298 B.n719 B.n718 163.367
R1299 B.n718 B.n49 163.367
R1300 B.n714 B.n49 163.367
R1301 B.n714 B.n713 163.367
R1302 B.n713 B.n712 163.367
R1303 B.n712 B.n51 163.367
R1304 B.n708 B.n51 163.367
R1305 B.n708 B.n707 163.367
R1306 B.n707 B.n706 163.367
R1307 B.n706 B.n53 163.367
R1308 B.n702 B.n53 163.367
R1309 B.n702 B.n701 163.367
R1310 B.n701 B.n700 163.367
R1311 B.n700 B.n58 163.367
R1312 B.n696 B.n58 163.367
R1313 B.n696 B.n695 163.367
R1314 B.n695 B.n694 163.367
R1315 B.n694 B.n60 163.367
R1316 B.n689 B.n60 163.367
R1317 B.n689 B.n688 163.367
R1318 B.n688 B.n687 163.367
R1319 B.n687 B.n64 163.367
R1320 B.n683 B.n64 163.367
R1321 B.n683 B.n682 163.367
R1322 B.n682 B.n681 163.367
R1323 B.n681 B.n66 163.367
R1324 B.n677 B.n66 163.367
R1325 B.n677 B.n676 163.367
R1326 B.n676 B.n675 163.367
R1327 B.n675 B.n68 163.367
R1328 B.n671 B.n68 163.367
R1329 B.n671 B.n670 163.367
R1330 B.n670 B.n669 163.367
R1331 B.n669 B.n70 163.367
R1332 B.n665 B.n70 163.367
R1333 B.n665 B.n664 163.367
R1334 B.n664 B.n663 163.367
R1335 B.n663 B.n72 163.367
R1336 B.n659 B.n72 163.367
R1337 B.n384 B.n383 77.9641
R1338 B.n170 B.n169 77.9641
R1339 B.n55 B.n54 77.9641
R1340 B.n62 B.n61 77.9641
R1341 B.n385 B.n384 59.5399
R1342 B.n370 B.n170 59.5399
R1343 B.n56 B.n55 59.5399
R1344 B.n692 B.n62 59.5399
R1345 B.n740 B.n739 35.4346
R1346 B.n660 B.n73 35.4346
R1347 B.n421 B.n420 35.4346
R1348 B.n338 B.n181 35.4346
R1349 B B.n859 18.0485
R1350 B.n739 B.n42 10.6151
R1351 B.n735 B.n42 10.6151
R1352 B.n735 B.n734 10.6151
R1353 B.n734 B.n733 10.6151
R1354 B.n733 B.n44 10.6151
R1355 B.n729 B.n44 10.6151
R1356 B.n729 B.n728 10.6151
R1357 B.n728 B.n727 10.6151
R1358 B.n727 B.n46 10.6151
R1359 B.n723 B.n46 10.6151
R1360 B.n723 B.n722 10.6151
R1361 B.n722 B.n721 10.6151
R1362 B.n721 B.n48 10.6151
R1363 B.n717 B.n48 10.6151
R1364 B.n717 B.n716 10.6151
R1365 B.n716 B.n715 10.6151
R1366 B.n715 B.n50 10.6151
R1367 B.n711 B.n50 10.6151
R1368 B.n711 B.n710 10.6151
R1369 B.n710 B.n709 10.6151
R1370 B.n709 B.n52 10.6151
R1371 B.n705 B.n704 10.6151
R1372 B.n704 B.n703 10.6151
R1373 B.n703 B.n57 10.6151
R1374 B.n699 B.n57 10.6151
R1375 B.n699 B.n698 10.6151
R1376 B.n698 B.n697 10.6151
R1377 B.n697 B.n59 10.6151
R1378 B.n693 B.n59 10.6151
R1379 B.n691 B.n690 10.6151
R1380 B.n690 B.n63 10.6151
R1381 B.n686 B.n63 10.6151
R1382 B.n686 B.n685 10.6151
R1383 B.n685 B.n684 10.6151
R1384 B.n684 B.n65 10.6151
R1385 B.n680 B.n65 10.6151
R1386 B.n680 B.n679 10.6151
R1387 B.n679 B.n678 10.6151
R1388 B.n678 B.n67 10.6151
R1389 B.n674 B.n67 10.6151
R1390 B.n674 B.n673 10.6151
R1391 B.n673 B.n672 10.6151
R1392 B.n672 B.n69 10.6151
R1393 B.n668 B.n69 10.6151
R1394 B.n668 B.n667 10.6151
R1395 B.n667 B.n666 10.6151
R1396 B.n666 B.n71 10.6151
R1397 B.n662 B.n71 10.6151
R1398 B.n662 B.n661 10.6151
R1399 B.n661 B.n660 10.6151
R1400 B.n422 B.n421 10.6151
R1401 B.n422 B.n151 10.6151
R1402 B.n426 B.n151 10.6151
R1403 B.n427 B.n426 10.6151
R1404 B.n428 B.n427 10.6151
R1405 B.n428 B.n149 10.6151
R1406 B.n432 B.n149 10.6151
R1407 B.n433 B.n432 10.6151
R1408 B.n434 B.n433 10.6151
R1409 B.n434 B.n147 10.6151
R1410 B.n438 B.n147 10.6151
R1411 B.n439 B.n438 10.6151
R1412 B.n440 B.n439 10.6151
R1413 B.n440 B.n145 10.6151
R1414 B.n444 B.n145 10.6151
R1415 B.n445 B.n444 10.6151
R1416 B.n446 B.n445 10.6151
R1417 B.n446 B.n143 10.6151
R1418 B.n450 B.n143 10.6151
R1419 B.n451 B.n450 10.6151
R1420 B.n452 B.n451 10.6151
R1421 B.n452 B.n141 10.6151
R1422 B.n456 B.n141 10.6151
R1423 B.n457 B.n456 10.6151
R1424 B.n458 B.n457 10.6151
R1425 B.n458 B.n139 10.6151
R1426 B.n462 B.n139 10.6151
R1427 B.n463 B.n462 10.6151
R1428 B.n464 B.n463 10.6151
R1429 B.n464 B.n137 10.6151
R1430 B.n468 B.n137 10.6151
R1431 B.n469 B.n468 10.6151
R1432 B.n470 B.n469 10.6151
R1433 B.n470 B.n135 10.6151
R1434 B.n474 B.n135 10.6151
R1435 B.n475 B.n474 10.6151
R1436 B.n476 B.n475 10.6151
R1437 B.n476 B.n133 10.6151
R1438 B.n480 B.n133 10.6151
R1439 B.n481 B.n480 10.6151
R1440 B.n482 B.n481 10.6151
R1441 B.n482 B.n131 10.6151
R1442 B.n486 B.n131 10.6151
R1443 B.n487 B.n486 10.6151
R1444 B.n488 B.n487 10.6151
R1445 B.n488 B.n129 10.6151
R1446 B.n492 B.n129 10.6151
R1447 B.n493 B.n492 10.6151
R1448 B.n494 B.n493 10.6151
R1449 B.n494 B.n127 10.6151
R1450 B.n498 B.n127 10.6151
R1451 B.n499 B.n498 10.6151
R1452 B.n500 B.n499 10.6151
R1453 B.n500 B.n125 10.6151
R1454 B.n504 B.n125 10.6151
R1455 B.n505 B.n504 10.6151
R1456 B.n506 B.n505 10.6151
R1457 B.n506 B.n123 10.6151
R1458 B.n510 B.n123 10.6151
R1459 B.n511 B.n510 10.6151
R1460 B.n512 B.n511 10.6151
R1461 B.n512 B.n121 10.6151
R1462 B.n516 B.n121 10.6151
R1463 B.n517 B.n516 10.6151
R1464 B.n518 B.n517 10.6151
R1465 B.n518 B.n119 10.6151
R1466 B.n522 B.n119 10.6151
R1467 B.n523 B.n522 10.6151
R1468 B.n524 B.n523 10.6151
R1469 B.n524 B.n117 10.6151
R1470 B.n528 B.n117 10.6151
R1471 B.n529 B.n528 10.6151
R1472 B.n530 B.n529 10.6151
R1473 B.n530 B.n115 10.6151
R1474 B.n534 B.n115 10.6151
R1475 B.n535 B.n534 10.6151
R1476 B.n536 B.n535 10.6151
R1477 B.n536 B.n113 10.6151
R1478 B.n540 B.n113 10.6151
R1479 B.n541 B.n540 10.6151
R1480 B.n542 B.n541 10.6151
R1481 B.n542 B.n111 10.6151
R1482 B.n546 B.n111 10.6151
R1483 B.n547 B.n546 10.6151
R1484 B.n548 B.n547 10.6151
R1485 B.n548 B.n109 10.6151
R1486 B.n552 B.n109 10.6151
R1487 B.n553 B.n552 10.6151
R1488 B.n554 B.n553 10.6151
R1489 B.n554 B.n107 10.6151
R1490 B.n558 B.n107 10.6151
R1491 B.n559 B.n558 10.6151
R1492 B.n560 B.n559 10.6151
R1493 B.n560 B.n105 10.6151
R1494 B.n564 B.n105 10.6151
R1495 B.n565 B.n564 10.6151
R1496 B.n566 B.n565 10.6151
R1497 B.n566 B.n103 10.6151
R1498 B.n570 B.n103 10.6151
R1499 B.n571 B.n570 10.6151
R1500 B.n572 B.n571 10.6151
R1501 B.n572 B.n101 10.6151
R1502 B.n576 B.n101 10.6151
R1503 B.n577 B.n576 10.6151
R1504 B.n578 B.n577 10.6151
R1505 B.n578 B.n99 10.6151
R1506 B.n582 B.n99 10.6151
R1507 B.n583 B.n582 10.6151
R1508 B.n584 B.n583 10.6151
R1509 B.n584 B.n97 10.6151
R1510 B.n588 B.n97 10.6151
R1511 B.n589 B.n588 10.6151
R1512 B.n590 B.n589 10.6151
R1513 B.n590 B.n95 10.6151
R1514 B.n594 B.n95 10.6151
R1515 B.n595 B.n594 10.6151
R1516 B.n596 B.n595 10.6151
R1517 B.n596 B.n93 10.6151
R1518 B.n600 B.n93 10.6151
R1519 B.n601 B.n600 10.6151
R1520 B.n602 B.n601 10.6151
R1521 B.n602 B.n91 10.6151
R1522 B.n606 B.n91 10.6151
R1523 B.n607 B.n606 10.6151
R1524 B.n608 B.n607 10.6151
R1525 B.n608 B.n89 10.6151
R1526 B.n612 B.n89 10.6151
R1527 B.n613 B.n612 10.6151
R1528 B.n614 B.n613 10.6151
R1529 B.n614 B.n87 10.6151
R1530 B.n618 B.n87 10.6151
R1531 B.n619 B.n618 10.6151
R1532 B.n620 B.n619 10.6151
R1533 B.n620 B.n85 10.6151
R1534 B.n624 B.n85 10.6151
R1535 B.n625 B.n624 10.6151
R1536 B.n626 B.n625 10.6151
R1537 B.n626 B.n83 10.6151
R1538 B.n630 B.n83 10.6151
R1539 B.n631 B.n630 10.6151
R1540 B.n632 B.n631 10.6151
R1541 B.n632 B.n81 10.6151
R1542 B.n636 B.n81 10.6151
R1543 B.n637 B.n636 10.6151
R1544 B.n638 B.n637 10.6151
R1545 B.n638 B.n79 10.6151
R1546 B.n642 B.n79 10.6151
R1547 B.n643 B.n642 10.6151
R1548 B.n644 B.n643 10.6151
R1549 B.n644 B.n77 10.6151
R1550 B.n648 B.n77 10.6151
R1551 B.n649 B.n648 10.6151
R1552 B.n650 B.n649 10.6151
R1553 B.n650 B.n75 10.6151
R1554 B.n654 B.n75 10.6151
R1555 B.n655 B.n654 10.6151
R1556 B.n656 B.n655 10.6151
R1557 B.n656 B.n73 10.6151
R1558 B.n339 B.n338 10.6151
R1559 B.n340 B.n339 10.6151
R1560 B.n340 B.n179 10.6151
R1561 B.n344 B.n179 10.6151
R1562 B.n345 B.n344 10.6151
R1563 B.n346 B.n345 10.6151
R1564 B.n346 B.n177 10.6151
R1565 B.n350 B.n177 10.6151
R1566 B.n351 B.n350 10.6151
R1567 B.n352 B.n351 10.6151
R1568 B.n352 B.n175 10.6151
R1569 B.n356 B.n175 10.6151
R1570 B.n357 B.n356 10.6151
R1571 B.n358 B.n357 10.6151
R1572 B.n358 B.n173 10.6151
R1573 B.n362 B.n173 10.6151
R1574 B.n363 B.n362 10.6151
R1575 B.n364 B.n363 10.6151
R1576 B.n364 B.n171 10.6151
R1577 B.n368 B.n171 10.6151
R1578 B.n369 B.n368 10.6151
R1579 B.n371 B.n167 10.6151
R1580 B.n375 B.n167 10.6151
R1581 B.n376 B.n375 10.6151
R1582 B.n377 B.n376 10.6151
R1583 B.n377 B.n165 10.6151
R1584 B.n381 B.n165 10.6151
R1585 B.n382 B.n381 10.6151
R1586 B.n386 B.n382 10.6151
R1587 B.n390 B.n163 10.6151
R1588 B.n391 B.n390 10.6151
R1589 B.n392 B.n391 10.6151
R1590 B.n392 B.n161 10.6151
R1591 B.n396 B.n161 10.6151
R1592 B.n397 B.n396 10.6151
R1593 B.n398 B.n397 10.6151
R1594 B.n398 B.n159 10.6151
R1595 B.n402 B.n159 10.6151
R1596 B.n403 B.n402 10.6151
R1597 B.n404 B.n403 10.6151
R1598 B.n404 B.n157 10.6151
R1599 B.n408 B.n157 10.6151
R1600 B.n409 B.n408 10.6151
R1601 B.n410 B.n409 10.6151
R1602 B.n410 B.n155 10.6151
R1603 B.n414 B.n155 10.6151
R1604 B.n415 B.n414 10.6151
R1605 B.n416 B.n415 10.6151
R1606 B.n416 B.n153 10.6151
R1607 B.n420 B.n153 10.6151
R1608 B.n334 B.n181 10.6151
R1609 B.n334 B.n333 10.6151
R1610 B.n333 B.n332 10.6151
R1611 B.n332 B.n183 10.6151
R1612 B.n328 B.n183 10.6151
R1613 B.n328 B.n327 10.6151
R1614 B.n327 B.n326 10.6151
R1615 B.n326 B.n185 10.6151
R1616 B.n322 B.n185 10.6151
R1617 B.n322 B.n321 10.6151
R1618 B.n321 B.n320 10.6151
R1619 B.n320 B.n187 10.6151
R1620 B.n316 B.n187 10.6151
R1621 B.n316 B.n315 10.6151
R1622 B.n315 B.n314 10.6151
R1623 B.n314 B.n189 10.6151
R1624 B.n310 B.n189 10.6151
R1625 B.n310 B.n309 10.6151
R1626 B.n309 B.n308 10.6151
R1627 B.n308 B.n191 10.6151
R1628 B.n304 B.n191 10.6151
R1629 B.n304 B.n303 10.6151
R1630 B.n303 B.n302 10.6151
R1631 B.n302 B.n193 10.6151
R1632 B.n298 B.n193 10.6151
R1633 B.n298 B.n297 10.6151
R1634 B.n297 B.n296 10.6151
R1635 B.n296 B.n195 10.6151
R1636 B.n292 B.n195 10.6151
R1637 B.n292 B.n291 10.6151
R1638 B.n291 B.n290 10.6151
R1639 B.n290 B.n197 10.6151
R1640 B.n286 B.n197 10.6151
R1641 B.n286 B.n285 10.6151
R1642 B.n285 B.n284 10.6151
R1643 B.n284 B.n199 10.6151
R1644 B.n280 B.n199 10.6151
R1645 B.n280 B.n279 10.6151
R1646 B.n279 B.n278 10.6151
R1647 B.n278 B.n201 10.6151
R1648 B.n274 B.n201 10.6151
R1649 B.n274 B.n273 10.6151
R1650 B.n273 B.n272 10.6151
R1651 B.n272 B.n203 10.6151
R1652 B.n268 B.n203 10.6151
R1653 B.n268 B.n267 10.6151
R1654 B.n267 B.n266 10.6151
R1655 B.n266 B.n205 10.6151
R1656 B.n262 B.n205 10.6151
R1657 B.n262 B.n261 10.6151
R1658 B.n261 B.n260 10.6151
R1659 B.n260 B.n207 10.6151
R1660 B.n256 B.n207 10.6151
R1661 B.n256 B.n255 10.6151
R1662 B.n255 B.n254 10.6151
R1663 B.n254 B.n209 10.6151
R1664 B.n250 B.n209 10.6151
R1665 B.n250 B.n249 10.6151
R1666 B.n249 B.n248 10.6151
R1667 B.n248 B.n211 10.6151
R1668 B.n244 B.n211 10.6151
R1669 B.n244 B.n243 10.6151
R1670 B.n243 B.n242 10.6151
R1671 B.n242 B.n213 10.6151
R1672 B.n238 B.n213 10.6151
R1673 B.n238 B.n237 10.6151
R1674 B.n237 B.n236 10.6151
R1675 B.n236 B.n215 10.6151
R1676 B.n232 B.n215 10.6151
R1677 B.n232 B.n231 10.6151
R1678 B.n231 B.n230 10.6151
R1679 B.n230 B.n217 10.6151
R1680 B.n226 B.n217 10.6151
R1681 B.n226 B.n225 10.6151
R1682 B.n225 B.n224 10.6151
R1683 B.n224 B.n219 10.6151
R1684 B.n220 B.n219 10.6151
R1685 B.n220 B.n0 10.6151
R1686 B.n855 B.n1 10.6151
R1687 B.n855 B.n854 10.6151
R1688 B.n854 B.n853 10.6151
R1689 B.n853 B.n4 10.6151
R1690 B.n849 B.n4 10.6151
R1691 B.n849 B.n848 10.6151
R1692 B.n848 B.n847 10.6151
R1693 B.n847 B.n6 10.6151
R1694 B.n843 B.n6 10.6151
R1695 B.n843 B.n842 10.6151
R1696 B.n842 B.n841 10.6151
R1697 B.n841 B.n8 10.6151
R1698 B.n837 B.n8 10.6151
R1699 B.n837 B.n836 10.6151
R1700 B.n836 B.n835 10.6151
R1701 B.n835 B.n10 10.6151
R1702 B.n831 B.n10 10.6151
R1703 B.n831 B.n830 10.6151
R1704 B.n830 B.n829 10.6151
R1705 B.n829 B.n12 10.6151
R1706 B.n825 B.n12 10.6151
R1707 B.n825 B.n824 10.6151
R1708 B.n824 B.n823 10.6151
R1709 B.n823 B.n14 10.6151
R1710 B.n819 B.n14 10.6151
R1711 B.n819 B.n818 10.6151
R1712 B.n818 B.n817 10.6151
R1713 B.n817 B.n16 10.6151
R1714 B.n813 B.n16 10.6151
R1715 B.n813 B.n812 10.6151
R1716 B.n812 B.n811 10.6151
R1717 B.n811 B.n18 10.6151
R1718 B.n807 B.n18 10.6151
R1719 B.n807 B.n806 10.6151
R1720 B.n806 B.n805 10.6151
R1721 B.n805 B.n20 10.6151
R1722 B.n801 B.n20 10.6151
R1723 B.n801 B.n800 10.6151
R1724 B.n800 B.n799 10.6151
R1725 B.n799 B.n22 10.6151
R1726 B.n795 B.n22 10.6151
R1727 B.n795 B.n794 10.6151
R1728 B.n794 B.n793 10.6151
R1729 B.n793 B.n24 10.6151
R1730 B.n789 B.n24 10.6151
R1731 B.n789 B.n788 10.6151
R1732 B.n788 B.n787 10.6151
R1733 B.n787 B.n26 10.6151
R1734 B.n783 B.n26 10.6151
R1735 B.n783 B.n782 10.6151
R1736 B.n782 B.n781 10.6151
R1737 B.n781 B.n28 10.6151
R1738 B.n777 B.n28 10.6151
R1739 B.n777 B.n776 10.6151
R1740 B.n776 B.n775 10.6151
R1741 B.n775 B.n30 10.6151
R1742 B.n771 B.n30 10.6151
R1743 B.n771 B.n770 10.6151
R1744 B.n770 B.n769 10.6151
R1745 B.n769 B.n32 10.6151
R1746 B.n765 B.n32 10.6151
R1747 B.n765 B.n764 10.6151
R1748 B.n764 B.n763 10.6151
R1749 B.n763 B.n34 10.6151
R1750 B.n759 B.n34 10.6151
R1751 B.n759 B.n758 10.6151
R1752 B.n758 B.n757 10.6151
R1753 B.n757 B.n36 10.6151
R1754 B.n753 B.n36 10.6151
R1755 B.n753 B.n752 10.6151
R1756 B.n752 B.n751 10.6151
R1757 B.n751 B.n38 10.6151
R1758 B.n747 B.n38 10.6151
R1759 B.n747 B.n746 10.6151
R1760 B.n746 B.n745 10.6151
R1761 B.n745 B.n40 10.6151
R1762 B.n741 B.n40 10.6151
R1763 B.n741 B.n740 10.6151
R1764 B.n705 B.n56 6.5566
R1765 B.n693 B.n692 6.5566
R1766 B.n371 B.n370 6.5566
R1767 B.n386 B.n385 6.5566
R1768 B.n56 B.n52 4.05904
R1769 B.n692 B.n691 4.05904
R1770 B.n370 B.n369 4.05904
R1771 B.n385 B.n163 4.05904
R1772 B.n859 B.n0 2.81026
R1773 B.n859 B.n1 2.81026
R1774 VP.n33 VP.n32 161.3
R1775 VP.n34 VP.n29 161.3
R1776 VP.n36 VP.n35 161.3
R1777 VP.n37 VP.n28 161.3
R1778 VP.n39 VP.n38 161.3
R1779 VP.n40 VP.n27 161.3
R1780 VP.n42 VP.n41 161.3
R1781 VP.n43 VP.n26 161.3
R1782 VP.n45 VP.n44 161.3
R1783 VP.n46 VP.n25 161.3
R1784 VP.n48 VP.n47 161.3
R1785 VP.n49 VP.n24 161.3
R1786 VP.n51 VP.n50 161.3
R1787 VP.n52 VP.n23 161.3
R1788 VP.n54 VP.n53 161.3
R1789 VP.n55 VP.n22 161.3
R1790 VP.n58 VP.n57 161.3
R1791 VP.n59 VP.n21 161.3
R1792 VP.n61 VP.n60 161.3
R1793 VP.n62 VP.n20 161.3
R1794 VP.n64 VP.n63 161.3
R1795 VP.n65 VP.n19 161.3
R1796 VP.n67 VP.n66 161.3
R1797 VP.n68 VP.n18 161.3
R1798 VP.n70 VP.n69 161.3
R1799 VP.n125 VP.n124 161.3
R1800 VP.n123 VP.n1 161.3
R1801 VP.n122 VP.n121 161.3
R1802 VP.n120 VP.n2 161.3
R1803 VP.n119 VP.n118 161.3
R1804 VP.n117 VP.n3 161.3
R1805 VP.n116 VP.n115 161.3
R1806 VP.n114 VP.n4 161.3
R1807 VP.n113 VP.n112 161.3
R1808 VP.n110 VP.n5 161.3
R1809 VP.n109 VP.n108 161.3
R1810 VP.n107 VP.n6 161.3
R1811 VP.n106 VP.n105 161.3
R1812 VP.n104 VP.n7 161.3
R1813 VP.n103 VP.n102 161.3
R1814 VP.n101 VP.n8 161.3
R1815 VP.n100 VP.n99 161.3
R1816 VP.n98 VP.n9 161.3
R1817 VP.n97 VP.n96 161.3
R1818 VP.n95 VP.n10 161.3
R1819 VP.n94 VP.n93 161.3
R1820 VP.n92 VP.n11 161.3
R1821 VP.n91 VP.n90 161.3
R1822 VP.n89 VP.n12 161.3
R1823 VP.n88 VP.n87 161.3
R1824 VP.n85 VP.n13 161.3
R1825 VP.n84 VP.n83 161.3
R1826 VP.n82 VP.n14 161.3
R1827 VP.n81 VP.n80 161.3
R1828 VP.n79 VP.n15 161.3
R1829 VP.n78 VP.n77 161.3
R1830 VP.n76 VP.n16 161.3
R1831 VP.n75 VP.n74 161.3
R1832 VP.n73 VP.n72 88.1101
R1833 VP.n126 VP.n0 88.1101
R1834 VP.n71 VP.n17 88.1101
R1835 VP.n31 VP.n30 74.0089
R1836 VP.n30 VP.t9 66.2846
R1837 VP.n72 VP.n71 53.9842
R1838 VP.n80 VP.n79 43.4072
R1839 VP.n118 VP.n2 43.4072
R1840 VP.n63 VP.n19 43.4072
R1841 VP.n93 VP.n92 41.4647
R1842 VP.n105 VP.n6 41.4647
R1843 VP.n50 VP.n23 41.4647
R1844 VP.n38 VP.n37 41.4647
R1845 VP.n93 VP.n10 39.5221
R1846 VP.n105 VP.n104 39.5221
R1847 VP.n50 VP.n49 39.5221
R1848 VP.n38 VP.n27 39.5221
R1849 VP.n80 VP.n14 37.5796
R1850 VP.n118 VP.n117 37.5796
R1851 VP.n63 VP.n62 37.5796
R1852 VP.n99 VP.t6 34.681
R1853 VP.n73 VP.t2 34.681
R1854 VP.n86 VP.t4 34.681
R1855 VP.n111 VP.t8 34.681
R1856 VP.n0 VP.t7 34.681
R1857 VP.n44 VP.t1 34.681
R1858 VP.n17 VP.t5 34.681
R1859 VP.n56 VP.t3 34.681
R1860 VP.n31 VP.t0 34.681
R1861 VP.n74 VP.n16 24.4675
R1862 VP.n78 VP.n16 24.4675
R1863 VP.n79 VP.n78 24.4675
R1864 VP.n84 VP.n14 24.4675
R1865 VP.n85 VP.n84 24.4675
R1866 VP.n87 VP.n12 24.4675
R1867 VP.n91 VP.n12 24.4675
R1868 VP.n92 VP.n91 24.4675
R1869 VP.n97 VP.n10 24.4675
R1870 VP.n98 VP.n97 24.4675
R1871 VP.n99 VP.n98 24.4675
R1872 VP.n99 VP.n8 24.4675
R1873 VP.n103 VP.n8 24.4675
R1874 VP.n104 VP.n103 24.4675
R1875 VP.n109 VP.n6 24.4675
R1876 VP.n110 VP.n109 24.4675
R1877 VP.n112 VP.n110 24.4675
R1878 VP.n116 VP.n4 24.4675
R1879 VP.n117 VP.n116 24.4675
R1880 VP.n122 VP.n2 24.4675
R1881 VP.n123 VP.n122 24.4675
R1882 VP.n124 VP.n123 24.4675
R1883 VP.n67 VP.n19 24.4675
R1884 VP.n68 VP.n67 24.4675
R1885 VP.n69 VP.n68 24.4675
R1886 VP.n54 VP.n23 24.4675
R1887 VP.n55 VP.n54 24.4675
R1888 VP.n57 VP.n55 24.4675
R1889 VP.n61 VP.n21 24.4675
R1890 VP.n62 VP.n61 24.4675
R1891 VP.n42 VP.n27 24.4675
R1892 VP.n43 VP.n42 24.4675
R1893 VP.n44 VP.n43 24.4675
R1894 VP.n44 VP.n25 24.4675
R1895 VP.n48 VP.n25 24.4675
R1896 VP.n49 VP.n48 24.4675
R1897 VP.n32 VP.n29 24.4675
R1898 VP.n36 VP.n29 24.4675
R1899 VP.n37 VP.n36 24.4675
R1900 VP.n86 VP.n85 23.4888
R1901 VP.n111 VP.n4 23.4888
R1902 VP.n56 VP.n21 23.4888
R1903 VP.n33 VP.n30 3.40896
R1904 VP.n74 VP.n73 1.95786
R1905 VP.n124 VP.n0 1.95786
R1906 VP.n69 VP.n17 1.95786
R1907 VP.n87 VP.n86 0.97918
R1908 VP.n112 VP.n111 0.97918
R1909 VP.n57 VP.n56 0.97918
R1910 VP.n32 VP.n31 0.97918
R1911 VP.n71 VP.n70 0.354971
R1912 VP.n75 VP.n72 0.354971
R1913 VP.n126 VP.n125 0.354971
R1914 VP VP.n126 0.26696
R1915 VP.n34 VP.n33 0.189894
R1916 VP.n35 VP.n34 0.189894
R1917 VP.n35 VP.n28 0.189894
R1918 VP.n39 VP.n28 0.189894
R1919 VP.n40 VP.n39 0.189894
R1920 VP.n41 VP.n40 0.189894
R1921 VP.n41 VP.n26 0.189894
R1922 VP.n45 VP.n26 0.189894
R1923 VP.n46 VP.n45 0.189894
R1924 VP.n47 VP.n46 0.189894
R1925 VP.n47 VP.n24 0.189894
R1926 VP.n51 VP.n24 0.189894
R1927 VP.n52 VP.n51 0.189894
R1928 VP.n53 VP.n52 0.189894
R1929 VP.n53 VP.n22 0.189894
R1930 VP.n58 VP.n22 0.189894
R1931 VP.n59 VP.n58 0.189894
R1932 VP.n60 VP.n59 0.189894
R1933 VP.n60 VP.n20 0.189894
R1934 VP.n64 VP.n20 0.189894
R1935 VP.n65 VP.n64 0.189894
R1936 VP.n66 VP.n65 0.189894
R1937 VP.n66 VP.n18 0.189894
R1938 VP.n70 VP.n18 0.189894
R1939 VP.n76 VP.n75 0.189894
R1940 VP.n77 VP.n76 0.189894
R1941 VP.n77 VP.n15 0.189894
R1942 VP.n81 VP.n15 0.189894
R1943 VP.n82 VP.n81 0.189894
R1944 VP.n83 VP.n82 0.189894
R1945 VP.n83 VP.n13 0.189894
R1946 VP.n88 VP.n13 0.189894
R1947 VP.n89 VP.n88 0.189894
R1948 VP.n90 VP.n89 0.189894
R1949 VP.n90 VP.n11 0.189894
R1950 VP.n94 VP.n11 0.189894
R1951 VP.n95 VP.n94 0.189894
R1952 VP.n96 VP.n95 0.189894
R1953 VP.n96 VP.n9 0.189894
R1954 VP.n100 VP.n9 0.189894
R1955 VP.n101 VP.n100 0.189894
R1956 VP.n102 VP.n101 0.189894
R1957 VP.n102 VP.n7 0.189894
R1958 VP.n106 VP.n7 0.189894
R1959 VP.n107 VP.n106 0.189894
R1960 VP.n108 VP.n107 0.189894
R1961 VP.n108 VP.n5 0.189894
R1962 VP.n113 VP.n5 0.189894
R1963 VP.n114 VP.n113 0.189894
R1964 VP.n115 VP.n114 0.189894
R1965 VP.n115 VP.n3 0.189894
R1966 VP.n119 VP.n3 0.189894
R1967 VP.n120 VP.n119 0.189894
R1968 VP.n121 VP.n120 0.189894
R1969 VP.n121 VP.n1 0.189894
R1970 VP.n125 VP.n1 0.189894
R1971 VDD1.n22 VDD1.n0 756.745
R1972 VDD1.n51 VDD1.n29 756.745
R1973 VDD1.n23 VDD1.n22 585
R1974 VDD1.n21 VDD1.n20 585
R1975 VDD1.n4 VDD1.n3 585
R1976 VDD1.n15 VDD1.n14 585
R1977 VDD1.n13 VDD1.n12 585
R1978 VDD1.n8 VDD1.n7 585
R1979 VDD1.n37 VDD1.n36 585
R1980 VDD1.n42 VDD1.n41 585
R1981 VDD1.n44 VDD1.n43 585
R1982 VDD1.n33 VDD1.n32 585
R1983 VDD1.n50 VDD1.n49 585
R1984 VDD1.n52 VDD1.n51 585
R1985 VDD1.n9 VDD1.t0 327.856
R1986 VDD1.n38 VDD1.t7 327.856
R1987 VDD1.n22 VDD1.n21 171.744
R1988 VDD1.n21 VDD1.n3 171.744
R1989 VDD1.n14 VDD1.n3 171.744
R1990 VDD1.n14 VDD1.n13 171.744
R1991 VDD1.n13 VDD1.n7 171.744
R1992 VDD1.n42 VDD1.n36 171.744
R1993 VDD1.n43 VDD1.n42 171.744
R1994 VDD1.n43 VDD1.n32 171.744
R1995 VDD1.n50 VDD1.n32 171.744
R1996 VDD1.n51 VDD1.n50 171.744
R1997 VDD1.n59 VDD1.n58 100.457
R1998 VDD1.n28 VDD1.n27 97.9127
R1999 VDD1.n57 VDD1.n56 97.9126
R2000 VDD1.n61 VDD1.n60 97.9126
R2001 VDD1.t0 VDD1.n7 85.8723
R2002 VDD1.t7 VDD1.n36 85.8723
R2003 VDD1.n28 VDD1.n26 52.9115
R2004 VDD1.n57 VDD1.n55 52.9115
R2005 VDD1.n61 VDD1.n59 47.0699
R2006 VDD1.n9 VDD1.n8 16.381
R2007 VDD1.n38 VDD1.n37 16.381
R2008 VDD1.n12 VDD1.n11 12.8005
R2009 VDD1.n41 VDD1.n40 12.8005
R2010 VDD1.n15 VDD1.n6 12.0247
R2011 VDD1.n44 VDD1.n35 12.0247
R2012 VDD1.n16 VDD1.n4 11.249
R2013 VDD1.n45 VDD1.n33 11.249
R2014 VDD1.n20 VDD1.n19 10.4732
R2015 VDD1.n49 VDD1.n48 10.4732
R2016 VDD1.n23 VDD1.n2 9.69747
R2017 VDD1.n52 VDD1.n31 9.69747
R2018 VDD1.n26 VDD1.n25 9.45567
R2019 VDD1.n55 VDD1.n54 9.45567
R2020 VDD1.n25 VDD1.n24 9.3005
R2021 VDD1.n2 VDD1.n1 9.3005
R2022 VDD1.n19 VDD1.n18 9.3005
R2023 VDD1.n17 VDD1.n16 9.3005
R2024 VDD1.n6 VDD1.n5 9.3005
R2025 VDD1.n11 VDD1.n10 9.3005
R2026 VDD1.n54 VDD1.n53 9.3005
R2027 VDD1.n31 VDD1.n30 9.3005
R2028 VDD1.n48 VDD1.n47 9.3005
R2029 VDD1.n46 VDD1.n45 9.3005
R2030 VDD1.n35 VDD1.n34 9.3005
R2031 VDD1.n40 VDD1.n39 9.3005
R2032 VDD1.n24 VDD1.n0 8.92171
R2033 VDD1.n53 VDD1.n29 8.92171
R2034 VDD1.n60 VDD1.t6 6.12197
R2035 VDD1.n60 VDD1.t4 6.12197
R2036 VDD1.n27 VDD1.t9 6.12197
R2037 VDD1.n27 VDD1.t8 6.12197
R2038 VDD1.n58 VDD1.t1 6.12197
R2039 VDD1.n58 VDD1.t2 6.12197
R2040 VDD1.n56 VDD1.t5 6.12197
R2041 VDD1.n56 VDD1.t3 6.12197
R2042 VDD1.n26 VDD1.n0 5.04292
R2043 VDD1.n55 VDD1.n29 5.04292
R2044 VDD1.n24 VDD1.n23 4.26717
R2045 VDD1.n53 VDD1.n52 4.26717
R2046 VDD1.n10 VDD1.n9 3.71853
R2047 VDD1.n39 VDD1.n38 3.71853
R2048 VDD1.n20 VDD1.n2 3.49141
R2049 VDD1.n49 VDD1.n31 3.49141
R2050 VDD1.n19 VDD1.n4 2.71565
R2051 VDD1.n48 VDD1.n33 2.71565
R2052 VDD1 VDD1.n61 2.54145
R2053 VDD1.n16 VDD1.n15 1.93989
R2054 VDD1.n45 VDD1.n44 1.93989
R2055 VDD1.n12 VDD1.n6 1.16414
R2056 VDD1.n41 VDD1.n35 1.16414
R2057 VDD1 VDD1.n28 0.925069
R2058 VDD1.n59 VDD1.n57 0.811533
R2059 VDD1.n11 VDD1.n8 0.388379
R2060 VDD1.n40 VDD1.n37 0.388379
R2061 VDD1.n25 VDD1.n1 0.155672
R2062 VDD1.n18 VDD1.n1 0.155672
R2063 VDD1.n18 VDD1.n17 0.155672
R2064 VDD1.n17 VDD1.n5 0.155672
R2065 VDD1.n10 VDD1.n5 0.155672
R2066 VDD1.n39 VDD1.n34 0.155672
R2067 VDD1.n46 VDD1.n34 0.155672
R2068 VDD1.n47 VDD1.n46 0.155672
R2069 VDD1.n47 VDD1.n30 0.155672
R2070 VDD1.n54 VDD1.n30 0.155672
C0 VDD2 VN 5.3289f
C1 w_n5794_n2030# B 10.522099f
C2 w_n5794_n2030# VDD2 2.93809f
C3 VN VP 8.76997f
C4 B VTAIL 2.52919f
C5 w_n5794_n2030# VP 13.3952f
C6 VDD2 VTAIL 8.368259f
C7 B VDD1 2.3642f
C8 w_n5794_n2030# VN 12.637599f
C9 VTAIL VP 7.06016f
C10 VDD2 VDD1 2.88153f
C11 VN VTAIL 7.04588f
C12 VDD1 VP 5.89202f
C13 w_n5794_n2030# VTAIL 2.44542f
C14 VDD2 B 2.52477f
C15 VN VDD1 0.1555f
C16 B VP 2.7516f
C17 w_n5794_n2030# VDD1 2.73815f
C18 VDD2 VP 0.726029f
C19 B VN 1.47146f
C20 VTAIL VDD1 8.30804f
C21 VDD2 VSUBS 2.526222f
C22 VDD1 VSUBS 2.276457f
C23 VTAIL VSUBS 0.782279f
C24 VN VSUBS 9.32371f
C25 VP VSUBS 5.080829f
C26 B VSUBS 5.979703f
C27 w_n5794_n2030# VSUBS 0.147191p
C28 VDD1.n0 VSUBS 0.03961f
C29 VDD1.n1 VSUBS 0.036327f
C30 VDD1.n2 VSUBS 0.019521f
C31 VDD1.n3 VSUBS 0.04614f
C32 VDD1.n4 VSUBS 0.020669f
C33 VDD1.n5 VSUBS 0.036327f
C34 VDD1.n6 VSUBS 0.019521f
C35 VDD1.n7 VSUBS 0.034605f
C36 VDD1.n8 VSUBS 0.029308f
C37 VDD1.t0 VSUBS 0.099594f
C38 VDD1.n9 VSUBS 0.153778f
C39 VDD1.n10 VSUBS 0.718361f
C40 VDD1.n11 VSUBS 0.019521f
C41 VDD1.n12 VSUBS 0.020669f
C42 VDD1.n13 VSUBS 0.04614f
C43 VDD1.n14 VSUBS 0.04614f
C44 VDD1.n15 VSUBS 0.020669f
C45 VDD1.n16 VSUBS 0.019521f
C46 VDD1.n17 VSUBS 0.036327f
C47 VDD1.n18 VSUBS 0.036327f
C48 VDD1.n19 VSUBS 0.019521f
C49 VDD1.n20 VSUBS 0.020669f
C50 VDD1.n21 VSUBS 0.04614f
C51 VDD1.n22 VSUBS 0.110658f
C52 VDD1.n23 VSUBS 0.020669f
C53 VDD1.n24 VSUBS 0.019521f
C54 VDD1.n25 VSUBS 0.085458f
C55 VDD1.n26 VSUBS 0.111927f
C56 VDD1.t9 VSUBS 0.152435f
C57 VDD1.t8 VSUBS 0.152435f
C58 VDD1.n27 VSUBS 0.975638f
C59 VDD1.n28 VSUBS 1.52637f
C60 VDD1.n29 VSUBS 0.03961f
C61 VDD1.n30 VSUBS 0.036327f
C62 VDD1.n31 VSUBS 0.019521f
C63 VDD1.n32 VSUBS 0.04614f
C64 VDD1.n33 VSUBS 0.020669f
C65 VDD1.n34 VSUBS 0.036327f
C66 VDD1.n35 VSUBS 0.019521f
C67 VDD1.n36 VSUBS 0.034605f
C68 VDD1.n37 VSUBS 0.029308f
C69 VDD1.t7 VSUBS 0.099594f
C70 VDD1.n38 VSUBS 0.153778f
C71 VDD1.n39 VSUBS 0.718361f
C72 VDD1.n40 VSUBS 0.019521f
C73 VDD1.n41 VSUBS 0.020669f
C74 VDD1.n42 VSUBS 0.04614f
C75 VDD1.n43 VSUBS 0.04614f
C76 VDD1.n44 VSUBS 0.020669f
C77 VDD1.n45 VSUBS 0.019521f
C78 VDD1.n46 VSUBS 0.036327f
C79 VDD1.n47 VSUBS 0.036327f
C80 VDD1.n48 VSUBS 0.019521f
C81 VDD1.n49 VSUBS 0.020669f
C82 VDD1.n50 VSUBS 0.04614f
C83 VDD1.n51 VSUBS 0.110658f
C84 VDD1.n52 VSUBS 0.020669f
C85 VDD1.n53 VSUBS 0.019521f
C86 VDD1.n54 VSUBS 0.085458f
C87 VDD1.n55 VSUBS 0.111927f
C88 VDD1.t5 VSUBS 0.152435f
C89 VDD1.t3 VSUBS 0.152435f
C90 VDD1.n56 VSUBS 0.975633f
C91 VDD1.n57 VSUBS 1.51413f
C92 VDD1.t1 VSUBS 0.152435f
C93 VDD1.t2 VSUBS 0.152435f
C94 VDD1.n58 VSUBS 1.00819f
C95 VDD1.n59 VSUBS 4.93981f
C96 VDD1.t6 VSUBS 0.152435f
C97 VDD1.t4 VSUBS 0.152435f
C98 VDD1.n60 VSUBS 0.975633f
C99 VDD1.n61 VSUBS 4.79219f
C100 VP.t7 VSUBS 1.88781f
C101 VP.n0 VSUBS 0.83733f
C102 VP.n1 VSUBS 0.036682f
C103 VP.n2 VSUBS 0.071603f
C104 VP.n3 VSUBS 0.036682f
C105 VP.n4 VSUBS 0.067016f
C106 VP.n5 VSUBS 0.036682f
C107 VP.n6 VSUBS 0.072514f
C108 VP.n7 VSUBS 0.036682f
C109 VP.n8 VSUBS 0.068366f
C110 VP.n9 VSUBS 0.036682f
C111 VP.t6 VSUBS 1.88781f
C112 VP.n10 VSUBS 0.073249f
C113 VP.n11 VSUBS 0.036682f
C114 VP.n12 VSUBS 0.068366f
C115 VP.n13 VSUBS 0.036682f
C116 VP.t4 VSUBS 1.88781f
C117 VP.n14 VSUBS 0.073781f
C118 VP.n15 VSUBS 0.036682f
C119 VP.n16 VSUBS 0.068366f
C120 VP.t5 VSUBS 1.88781f
C121 VP.n17 VSUBS 0.83733f
C122 VP.n18 VSUBS 0.036682f
C123 VP.n19 VSUBS 0.071603f
C124 VP.n20 VSUBS 0.036682f
C125 VP.n21 VSUBS 0.067016f
C126 VP.n22 VSUBS 0.036682f
C127 VP.n23 VSUBS 0.072514f
C128 VP.n24 VSUBS 0.036682f
C129 VP.n25 VSUBS 0.068366f
C130 VP.n26 VSUBS 0.036682f
C131 VP.t1 VSUBS 1.88781f
C132 VP.n27 VSUBS 0.073249f
C133 VP.n28 VSUBS 0.036682f
C134 VP.n29 VSUBS 0.068366f
C135 VP.t9 VSUBS 2.35674f
C136 VP.n30 VSUBS 0.805773f
C137 VP.t0 VSUBS 1.88781f
C138 VP.n31 VSUBS 0.821395f
C139 VP.n32 VSUBS 0.035963f
C140 VP.n33 VSUBS 0.466048f
C141 VP.n34 VSUBS 0.036682f
C142 VP.n35 VSUBS 0.036682f
C143 VP.n36 VSUBS 0.068366f
C144 VP.n37 VSUBS 0.072514f
C145 VP.n38 VSUBS 0.029701f
C146 VP.n39 VSUBS 0.036682f
C147 VP.n40 VSUBS 0.036682f
C148 VP.n41 VSUBS 0.036682f
C149 VP.n42 VSUBS 0.068366f
C150 VP.n43 VSUBS 0.068366f
C151 VP.n44 VSUBS 0.739784f
C152 VP.n45 VSUBS 0.036682f
C153 VP.n46 VSUBS 0.036682f
C154 VP.n47 VSUBS 0.036682f
C155 VP.n48 VSUBS 0.068366f
C156 VP.n49 VSUBS 0.073249f
C157 VP.n50 VSUBS 0.029701f
C158 VP.n51 VSUBS 0.036682f
C159 VP.n52 VSUBS 0.036682f
C160 VP.n53 VSUBS 0.036682f
C161 VP.n54 VSUBS 0.068366f
C162 VP.n55 VSUBS 0.068366f
C163 VP.t3 VSUBS 1.88781f
C164 VP.n56 VSUBS 0.705171f
C165 VP.n57 VSUBS 0.035963f
C166 VP.n58 VSUBS 0.036682f
C167 VP.n59 VSUBS 0.036682f
C168 VP.n60 VSUBS 0.036682f
C169 VP.n61 VSUBS 0.068366f
C170 VP.n62 VSUBS 0.073781f
C171 VP.n63 VSUBS 0.03008f
C172 VP.n64 VSUBS 0.036682f
C173 VP.n65 VSUBS 0.036682f
C174 VP.n66 VSUBS 0.036682f
C175 VP.n67 VSUBS 0.068366f
C176 VP.n68 VSUBS 0.068366f
C177 VP.n69 VSUBS 0.037313f
C178 VP.n70 VSUBS 0.059204f
C179 VP.n71 VSUBS 2.34673f
C180 VP.n72 VSUBS 2.37116f
C181 VP.t2 VSUBS 1.88781f
C182 VP.n73 VSUBS 0.83733f
C183 VP.n74 VSUBS 0.037313f
C184 VP.n75 VSUBS 0.059204f
C185 VP.n76 VSUBS 0.036682f
C186 VP.n77 VSUBS 0.036682f
C187 VP.n78 VSUBS 0.068366f
C188 VP.n79 VSUBS 0.071603f
C189 VP.n80 VSUBS 0.03008f
C190 VP.n81 VSUBS 0.036682f
C191 VP.n82 VSUBS 0.036682f
C192 VP.n83 VSUBS 0.036682f
C193 VP.n84 VSUBS 0.068366f
C194 VP.n85 VSUBS 0.067016f
C195 VP.n86 VSUBS 0.705171f
C196 VP.n87 VSUBS 0.035963f
C197 VP.n88 VSUBS 0.036682f
C198 VP.n89 VSUBS 0.036682f
C199 VP.n90 VSUBS 0.036682f
C200 VP.n91 VSUBS 0.068366f
C201 VP.n92 VSUBS 0.072514f
C202 VP.n93 VSUBS 0.029701f
C203 VP.n94 VSUBS 0.036682f
C204 VP.n95 VSUBS 0.036682f
C205 VP.n96 VSUBS 0.036682f
C206 VP.n97 VSUBS 0.068366f
C207 VP.n98 VSUBS 0.068366f
C208 VP.n99 VSUBS 0.739784f
C209 VP.n100 VSUBS 0.036682f
C210 VP.n101 VSUBS 0.036682f
C211 VP.n102 VSUBS 0.036682f
C212 VP.n103 VSUBS 0.068366f
C213 VP.n104 VSUBS 0.073249f
C214 VP.n105 VSUBS 0.029701f
C215 VP.n106 VSUBS 0.036682f
C216 VP.n107 VSUBS 0.036682f
C217 VP.n108 VSUBS 0.036682f
C218 VP.n109 VSUBS 0.068366f
C219 VP.n110 VSUBS 0.068366f
C220 VP.t8 VSUBS 1.88781f
C221 VP.n111 VSUBS 0.705171f
C222 VP.n112 VSUBS 0.035963f
C223 VP.n113 VSUBS 0.036682f
C224 VP.n114 VSUBS 0.036682f
C225 VP.n115 VSUBS 0.036682f
C226 VP.n116 VSUBS 0.068366f
C227 VP.n117 VSUBS 0.073781f
C228 VP.n118 VSUBS 0.03008f
C229 VP.n119 VSUBS 0.036682f
C230 VP.n120 VSUBS 0.036682f
C231 VP.n121 VSUBS 0.036682f
C232 VP.n122 VSUBS 0.068366f
C233 VP.n123 VSUBS 0.068366f
C234 VP.n124 VSUBS 0.037313f
C235 VP.n125 VSUBS 0.059204f
C236 VP.n126 VSUBS 0.111388f
C237 B.n0 VSUBS 0.007624f
C238 B.n1 VSUBS 0.007624f
C239 B.n2 VSUBS 0.012056f
C240 B.n3 VSUBS 0.012056f
C241 B.n4 VSUBS 0.012056f
C242 B.n5 VSUBS 0.012056f
C243 B.n6 VSUBS 0.012056f
C244 B.n7 VSUBS 0.012056f
C245 B.n8 VSUBS 0.012056f
C246 B.n9 VSUBS 0.012056f
C247 B.n10 VSUBS 0.012056f
C248 B.n11 VSUBS 0.012056f
C249 B.n12 VSUBS 0.012056f
C250 B.n13 VSUBS 0.012056f
C251 B.n14 VSUBS 0.012056f
C252 B.n15 VSUBS 0.012056f
C253 B.n16 VSUBS 0.012056f
C254 B.n17 VSUBS 0.012056f
C255 B.n18 VSUBS 0.012056f
C256 B.n19 VSUBS 0.012056f
C257 B.n20 VSUBS 0.012056f
C258 B.n21 VSUBS 0.012056f
C259 B.n22 VSUBS 0.012056f
C260 B.n23 VSUBS 0.012056f
C261 B.n24 VSUBS 0.012056f
C262 B.n25 VSUBS 0.012056f
C263 B.n26 VSUBS 0.012056f
C264 B.n27 VSUBS 0.012056f
C265 B.n28 VSUBS 0.012056f
C266 B.n29 VSUBS 0.012056f
C267 B.n30 VSUBS 0.012056f
C268 B.n31 VSUBS 0.012056f
C269 B.n32 VSUBS 0.012056f
C270 B.n33 VSUBS 0.012056f
C271 B.n34 VSUBS 0.012056f
C272 B.n35 VSUBS 0.012056f
C273 B.n36 VSUBS 0.012056f
C274 B.n37 VSUBS 0.012056f
C275 B.n38 VSUBS 0.012056f
C276 B.n39 VSUBS 0.012056f
C277 B.n40 VSUBS 0.012056f
C278 B.n41 VSUBS 0.029353f
C279 B.n42 VSUBS 0.012056f
C280 B.n43 VSUBS 0.012056f
C281 B.n44 VSUBS 0.012056f
C282 B.n45 VSUBS 0.012056f
C283 B.n46 VSUBS 0.012056f
C284 B.n47 VSUBS 0.012056f
C285 B.n48 VSUBS 0.012056f
C286 B.n49 VSUBS 0.012056f
C287 B.n50 VSUBS 0.012056f
C288 B.n51 VSUBS 0.012056f
C289 B.n52 VSUBS 0.008333f
C290 B.n53 VSUBS 0.012056f
C291 B.t11 VSUBS 0.134014f
C292 B.t10 VSUBS 0.189341f
C293 B.t9 VSUBS 1.62753f
C294 B.n54 VSUBS 0.315658f
C295 B.n55 VSUBS 0.254357f
C296 B.n56 VSUBS 0.027932f
C297 B.n57 VSUBS 0.012056f
C298 B.n58 VSUBS 0.012056f
C299 B.n59 VSUBS 0.012056f
C300 B.n60 VSUBS 0.012056f
C301 B.t8 VSUBS 0.134017f
C302 B.t7 VSUBS 0.189343f
C303 B.t6 VSUBS 1.62753f
C304 B.n61 VSUBS 0.315656f
C305 B.n62 VSUBS 0.254354f
C306 B.n63 VSUBS 0.012056f
C307 B.n64 VSUBS 0.012056f
C308 B.n65 VSUBS 0.012056f
C309 B.n66 VSUBS 0.012056f
C310 B.n67 VSUBS 0.012056f
C311 B.n68 VSUBS 0.012056f
C312 B.n69 VSUBS 0.012056f
C313 B.n70 VSUBS 0.012056f
C314 B.n71 VSUBS 0.012056f
C315 B.n72 VSUBS 0.012056f
C316 B.n73 VSUBS 0.030666f
C317 B.n74 VSUBS 0.012056f
C318 B.n75 VSUBS 0.012056f
C319 B.n76 VSUBS 0.012056f
C320 B.n77 VSUBS 0.012056f
C321 B.n78 VSUBS 0.012056f
C322 B.n79 VSUBS 0.012056f
C323 B.n80 VSUBS 0.012056f
C324 B.n81 VSUBS 0.012056f
C325 B.n82 VSUBS 0.012056f
C326 B.n83 VSUBS 0.012056f
C327 B.n84 VSUBS 0.012056f
C328 B.n85 VSUBS 0.012056f
C329 B.n86 VSUBS 0.012056f
C330 B.n87 VSUBS 0.012056f
C331 B.n88 VSUBS 0.012056f
C332 B.n89 VSUBS 0.012056f
C333 B.n90 VSUBS 0.012056f
C334 B.n91 VSUBS 0.012056f
C335 B.n92 VSUBS 0.012056f
C336 B.n93 VSUBS 0.012056f
C337 B.n94 VSUBS 0.012056f
C338 B.n95 VSUBS 0.012056f
C339 B.n96 VSUBS 0.012056f
C340 B.n97 VSUBS 0.012056f
C341 B.n98 VSUBS 0.012056f
C342 B.n99 VSUBS 0.012056f
C343 B.n100 VSUBS 0.012056f
C344 B.n101 VSUBS 0.012056f
C345 B.n102 VSUBS 0.012056f
C346 B.n103 VSUBS 0.012056f
C347 B.n104 VSUBS 0.012056f
C348 B.n105 VSUBS 0.012056f
C349 B.n106 VSUBS 0.012056f
C350 B.n107 VSUBS 0.012056f
C351 B.n108 VSUBS 0.012056f
C352 B.n109 VSUBS 0.012056f
C353 B.n110 VSUBS 0.012056f
C354 B.n111 VSUBS 0.012056f
C355 B.n112 VSUBS 0.012056f
C356 B.n113 VSUBS 0.012056f
C357 B.n114 VSUBS 0.012056f
C358 B.n115 VSUBS 0.012056f
C359 B.n116 VSUBS 0.012056f
C360 B.n117 VSUBS 0.012056f
C361 B.n118 VSUBS 0.012056f
C362 B.n119 VSUBS 0.012056f
C363 B.n120 VSUBS 0.012056f
C364 B.n121 VSUBS 0.012056f
C365 B.n122 VSUBS 0.012056f
C366 B.n123 VSUBS 0.012056f
C367 B.n124 VSUBS 0.012056f
C368 B.n125 VSUBS 0.012056f
C369 B.n126 VSUBS 0.012056f
C370 B.n127 VSUBS 0.012056f
C371 B.n128 VSUBS 0.012056f
C372 B.n129 VSUBS 0.012056f
C373 B.n130 VSUBS 0.012056f
C374 B.n131 VSUBS 0.012056f
C375 B.n132 VSUBS 0.012056f
C376 B.n133 VSUBS 0.012056f
C377 B.n134 VSUBS 0.012056f
C378 B.n135 VSUBS 0.012056f
C379 B.n136 VSUBS 0.012056f
C380 B.n137 VSUBS 0.012056f
C381 B.n138 VSUBS 0.012056f
C382 B.n139 VSUBS 0.012056f
C383 B.n140 VSUBS 0.012056f
C384 B.n141 VSUBS 0.012056f
C385 B.n142 VSUBS 0.012056f
C386 B.n143 VSUBS 0.012056f
C387 B.n144 VSUBS 0.012056f
C388 B.n145 VSUBS 0.012056f
C389 B.n146 VSUBS 0.012056f
C390 B.n147 VSUBS 0.012056f
C391 B.n148 VSUBS 0.012056f
C392 B.n149 VSUBS 0.012056f
C393 B.n150 VSUBS 0.012056f
C394 B.n151 VSUBS 0.012056f
C395 B.n152 VSUBS 0.029353f
C396 B.n153 VSUBS 0.012056f
C397 B.n154 VSUBS 0.012056f
C398 B.n155 VSUBS 0.012056f
C399 B.n156 VSUBS 0.012056f
C400 B.n157 VSUBS 0.012056f
C401 B.n158 VSUBS 0.012056f
C402 B.n159 VSUBS 0.012056f
C403 B.n160 VSUBS 0.012056f
C404 B.n161 VSUBS 0.012056f
C405 B.n162 VSUBS 0.012056f
C406 B.n163 VSUBS 0.008333f
C407 B.n164 VSUBS 0.012056f
C408 B.n165 VSUBS 0.012056f
C409 B.n166 VSUBS 0.012056f
C410 B.n167 VSUBS 0.012056f
C411 B.n168 VSUBS 0.012056f
C412 B.t4 VSUBS 0.134014f
C413 B.t5 VSUBS 0.189341f
C414 B.t3 VSUBS 1.62753f
C415 B.n169 VSUBS 0.315658f
C416 B.n170 VSUBS 0.254357f
C417 B.n171 VSUBS 0.012056f
C418 B.n172 VSUBS 0.012056f
C419 B.n173 VSUBS 0.012056f
C420 B.n174 VSUBS 0.012056f
C421 B.n175 VSUBS 0.012056f
C422 B.n176 VSUBS 0.012056f
C423 B.n177 VSUBS 0.012056f
C424 B.n178 VSUBS 0.012056f
C425 B.n179 VSUBS 0.012056f
C426 B.n180 VSUBS 0.012056f
C427 B.n181 VSUBS 0.029353f
C428 B.n182 VSUBS 0.012056f
C429 B.n183 VSUBS 0.012056f
C430 B.n184 VSUBS 0.012056f
C431 B.n185 VSUBS 0.012056f
C432 B.n186 VSUBS 0.012056f
C433 B.n187 VSUBS 0.012056f
C434 B.n188 VSUBS 0.012056f
C435 B.n189 VSUBS 0.012056f
C436 B.n190 VSUBS 0.012056f
C437 B.n191 VSUBS 0.012056f
C438 B.n192 VSUBS 0.012056f
C439 B.n193 VSUBS 0.012056f
C440 B.n194 VSUBS 0.012056f
C441 B.n195 VSUBS 0.012056f
C442 B.n196 VSUBS 0.012056f
C443 B.n197 VSUBS 0.012056f
C444 B.n198 VSUBS 0.012056f
C445 B.n199 VSUBS 0.012056f
C446 B.n200 VSUBS 0.012056f
C447 B.n201 VSUBS 0.012056f
C448 B.n202 VSUBS 0.012056f
C449 B.n203 VSUBS 0.012056f
C450 B.n204 VSUBS 0.012056f
C451 B.n205 VSUBS 0.012056f
C452 B.n206 VSUBS 0.012056f
C453 B.n207 VSUBS 0.012056f
C454 B.n208 VSUBS 0.012056f
C455 B.n209 VSUBS 0.012056f
C456 B.n210 VSUBS 0.012056f
C457 B.n211 VSUBS 0.012056f
C458 B.n212 VSUBS 0.012056f
C459 B.n213 VSUBS 0.012056f
C460 B.n214 VSUBS 0.012056f
C461 B.n215 VSUBS 0.012056f
C462 B.n216 VSUBS 0.012056f
C463 B.n217 VSUBS 0.012056f
C464 B.n218 VSUBS 0.012056f
C465 B.n219 VSUBS 0.012056f
C466 B.n220 VSUBS 0.012056f
C467 B.n221 VSUBS 0.012056f
C468 B.n222 VSUBS 0.012056f
C469 B.n223 VSUBS 0.012056f
C470 B.n224 VSUBS 0.012056f
C471 B.n225 VSUBS 0.012056f
C472 B.n226 VSUBS 0.012056f
C473 B.n227 VSUBS 0.012056f
C474 B.n228 VSUBS 0.012056f
C475 B.n229 VSUBS 0.012056f
C476 B.n230 VSUBS 0.012056f
C477 B.n231 VSUBS 0.012056f
C478 B.n232 VSUBS 0.012056f
C479 B.n233 VSUBS 0.012056f
C480 B.n234 VSUBS 0.012056f
C481 B.n235 VSUBS 0.012056f
C482 B.n236 VSUBS 0.012056f
C483 B.n237 VSUBS 0.012056f
C484 B.n238 VSUBS 0.012056f
C485 B.n239 VSUBS 0.012056f
C486 B.n240 VSUBS 0.012056f
C487 B.n241 VSUBS 0.012056f
C488 B.n242 VSUBS 0.012056f
C489 B.n243 VSUBS 0.012056f
C490 B.n244 VSUBS 0.012056f
C491 B.n245 VSUBS 0.012056f
C492 B.n246 VSUBS 0.012056f
C493 B.n247 VSUBS 0.012056f
C494 B.n248 VSUBS 0.012056f
C495 B.n249 VSUBS 0.012056f
C496 B.n250 VSUBS 0.012056f
C497 B.n251 VSUBS 0.012056f
C498 B.n252 VSUBS 0.012056f
C499 B.n253 VSUBS 0.012056f
C500 B.n254 VSUBS 0.012056f
C501 B.n255 VSUBS 0.012056f
C502 B.n256 VSUBS 0.012056f
C503 B.n257 VSUBS 0.012056f
C504 B.n258 VSUBS 0.012056f
C505 B.n259 VSUBS 0.012056f
C506 B.n260 VSUBS 0.012056f
C507 B.n261 VSUBS 0.012056f
C508 B.n262 VSUBS 0.012056f
C509 B.n263 VSUBS 0.012056f
C510 B.n264 VSUBS 0.012056f
C511 B.n265 VSUBS 0.012056f
C512 B.n266 VSUBS 0.012056f
C513 B.n267 VSUBS 0.012056f
C514 B.n268 VSUBS 0.012056f
C515 B.n269 VSUBS 0.012056f
C516 B.n270 VSUBS 0.012056f
C517 B.n271 VSUBS 0.012056f
C518 B.n272 VSUBS 0.012056f
C519 B.n273 VSUBS 0.012056f
C520 B.n274 VSUBS 0.012056f
C521 B.n275 VSUBS 0.012056f
C522 B.n276 VSUBS 0.012056f
C523 B.n277 VSUBS 0.012056f
C524 B.n278 VSUBS 0.012056f
C525 B.n279 VSUBS 0.012056f
C526 B.n280 VSUBS 0.012056f
C527 B.n281 VSUBS 0.012056f
C528 B.n282 VSUBS 0.012056f
C529 B.n283 VSUBS 0.012056f
C530 B.n284 VSUBS 0.012056f
C531 B.n285 VSUBS 0.012056f
C532 B.n286 VSUBS 0.012056f
C533 B.n287 VSUBS 0.012056f
C534 B.n288 VSUBS 0.012056f
C535 B.n289 VSUBS 0.012056f
C536 B.n290 VSUBS 0.012056f
C537 B.n291 VSUBS 0.012056f
C538 B.n292 VSUBS 0.012056f
C539 B.n293 VSUBS 0.012056f
C540 B.n294 VSUBS 0.012056f
C541 B.n295 VSUBS 0.012056f
C542 B.n296 VSUBS 0.012056f
C543 B.n297 VSUBS 0.012056f
C544 B.n298 VSUBS 0.012056f
C545 B.n299 VSUBS 0.012056f
C546 B.n300 VSUBS 0.012056f
C547 B.n301 VSUBS 0.012056f
C548 B.n302 VSUBS 0.012056f
C549 B.n303 VSUBS 0.012056f
C550 B.n304 VSUBS 0.012056f
C551 B.n305 VSUBS 0.012056f
C552 B.n306 VSUBS 0.012056f
C553 B.n307 VSUBS 0.012056f
C554 B.n308 VSUBS 0.012056f
C555 B.n309 VSUBS 0.012056f
C556 B.n310 VSUBS 0.012056f
C557 B.n311 VSUBS 0.012056f
C558 B.n312 VSUBS 0.012056f
C559 B.n313 VSUBS 0.012056f
C560 B.n314 VSUBS 0.012056f
C561 B.n315 VSUBS 0.012056f
C562 B.n316 VSUBS 0.012056f
C563 B.n317 VSUBS 0.012056f
C564 B.n318 VSUBS 0.012056f
C565 B.n319 VSUBS 0.012056f
C566 B.n320 VSUBS 0.012056f
C567 B.n321 VSUBS 0.012056f
C568 B.n322 VSUBS 0.012056f
C569 B.n323 VSUBS 0.012056f
C570 B.n324 VSUBS 0.012056f
C571 B.n325 VSUBS 0.012056f
C572 B.n326 VSUBS 0.012056f
C573 B.n327 VSUBS 0.012056f
C574 B.n328 VSUBS 0.012056f
C575 B.n329 VSUBS 0.012056f
C576 B.n330 VSUBS 0.012056f
C577 B.n331 VSUBS 0.012056f
C578 B.n332 VSUBS 0.012056f
C579 B.n333 VSUBS 0.012056f
C580 B.n334 VSUBS 0.012056f
C581 B.n335 VSUBS 0.012056f
C582 B.n336 VSUBS 0.029353f
C583 B.n337 VSUBS 0.030218f
C584 B.n338 VSUBS 0.030218f
C585 B.n339 VSUBS 0.012056f
C586 B.n340 VSUBS 0.012056f
C587 B.n341 VSUBS 0.012056f
C588 B.n342 VSUBS 0.012056f
C589 B.n343 VSUBS 0.012056f
C590 B.n344 VSUBS 0.012056f
C591 B.n345 VSUBS 0.012056f
C592 B.n346 VSUBS 0.012056f
C593 B.n347 VSUBS 0.012056f
C594 B.n348 VSUBS 0.012056f
C595 B.n349 VSUBS 0.012056f
C596 B.n350 VSUBS 0.012056f
C597 B.n351 VSUBS 0.012056f
C598 B.n352 VSUBS 0.012056f
C599 B.n353 VSUBS 0.012056f
C600 B.n354 VSUBS 0.012056f
C601 B.n355 VSUBS 0.012056f
C602 B.n356 VSUBS 0.012056f
C603 B.n357 VSUBS 0.012056f
C604 B.n358 VSUBS 0.012056f
C605 B.n359 VSUBS 0.012056f
C606 B.n360 VSUBS 0.012056f
C607 B.n361 VSUBS 0.012056f
C608 B.n362 VSUBS 0.012056f
C609 B.n363 VSUBS 0.012056f
C610 B.n364 VSUBS 0.012056f
C611 B.n365 VSUBS 0.012056f
C612 B.n366 VSUBS 0.012056f
C613 B.n367 VSUBS 0.012056f
C614 B.n368 VSUBS 0.012056f
C615 B.n369 VSUBS 0.008333f
C616 B.n370 VSUBS 0.027932f
C617 B.n371 VSUBS 0.009751f
C618 B.n372 VSUBS 0.012056f
C619 B.n373 VSUBS 0.012056f
C620 B.n374 VSUBS 0.012056f
C621 B.n375 VSUBS 0.012056f
C622 B.n376 VSUBS 0.012056f
C623 B.n377 VSUBS 0.012056f
C624 B.n378 VSUBS 0.012056f
C625 B.n379 VSUBS 0.012056f
C626 B.n380 VSUBS 0.012056f
C627 B.n381 VSUBS 0.012056f
C628 B.n382 VSUBS 0.012056f
C629 B.t1 VSUBS 0.134017f
C630 B.t2 VSUBS 0.189343f
C631 B.t0 VSUBS 1.62753f
C632 B.n383 VSUBS 0.315656f
C633 B.n384 VSUBS 0.254354f
C634 B.n385 VSUBS 0.027932f
C635 B.n386 VSUBS 0.009751f
C636 B.n387 VSUBS 0.012056f
C637 B.n388 VSUBS 0.012056f
C638 B.n389 VSUBS 0.012056f
C639 B.n390 VSUBS 0.012056f
C640 B.n391 VSUBS 0.012056f
C641 B.n392 VSUBS 0.012056f
C642 B.n393 VSUBS 0.012056f
C643 B.n394 VSUBS 0.012056f
C644 B.n395 VSUBS 0.012056f
C645 B.n396 VSUBS 0.012056f
C646 B.n397 VSUBS 0.012056f
C647 B.n398 VSUBS 0.012056f
C648 B.n399 VSUBS 0.012056f
C649 B.n400 VSUBS 0.012056f
C650 B.n401 VSUBS 0.012056f
C651 B.n402 VSUBS 0.012056f
C652 B.n403 VSUBS 0.012056f
C653 B.n404 VSUBS 0.012056f
C654 B.n405 VSUBS 0.012056f
C655 B.n406 VSUBS 0.012056f
C656 B.n407 VSUBS 0.012056f
C657 B.n408 VSUBS 0.012056f
C658 B.n409 VSUBS 0.012056f
C659 B.n410 VSUBS 0.012056f
C660 B.n411 VSUBS 0.012056f
C661 B.n412 VSUBS 0.012056f
C662 B.n413 VSUBS 0.012056f
C663 B.n414 VSUBS 0.012056f
C664 B.n415 VSUBS 0.012056f
C665 B.n416 VSUBS 0.012056f
C666 B.n417 VSUBS 0.012056f
C667 B.n418 VSUBS 0.012056f
C668 B.n419 VSUBS 0.030218f
C669 B.n420 VSUBS 0.030218f
C670 B.n421 VSUBS 0.029353f
C671 B.n422 VSUBS 0.012056f
C672 B.n423 VSUBS 0.012056f
C673 B.n424 VSUBS 0.012056f
C674 B.n425 VSUBS 0.012056f
C675 B.n426 VSUBS 0.012056f
C676 B.n427 VSUBS 0.012056f
C677 B.n428 VSUBS 0.012056f
C678 B.n429 VSUBS 0.012056f
C679 B.n430 VSUBS 0.012056f
C680 B.n431 VSUBS 0.012056f
C681 B.n432 VSUBS 0.012056f
C682 B.n433 VSUBS 0.012056f
C683 B.n434 VSUBS 0.012056f
C684 B.n435 VSUBS 0.012056f
C685 B.n436 VSUBS 0.012056f
C686 B.n437 VSUBS 0.012056f
C687 B.n438 VSUBS 0.012056f
C688 B.n439 VSUBS 0.012056f
C689 B.n440 VSUBS 0.012056f
C690 B.n441 VSUBS 0.012056f
C691 B.n442 VSUBS 0.012056f
C692 B.n443 VSUBS 0.012056f
C693 B.n444 VSUBS 0.012056f
C694 B.n445 VSUBS 0.012056f
C695 B.n446 VSUBS 0.012056f
C696 B.n447 VSUBS 0.012056f
C697 B.n448 VSUBS 0.012056f
C698 B.n449 VSUBS 0.012056f
C699 B.n450 VSUBS 0.012056f
C700 B.n451 VSUBS 0.012056f
C701 B.n452 VSUBS 0.012056f
C702 B.n453 VSUBS 0.012056f
C703 B.n454 VSUBS 0.012056f
C704 B.n455 VSUBS 0.012056f
C705 B.n456 VSUBS 0.012056f
C706 B.n457 VSUBS 0.012056f
C707 B.n458 VSUBS 0.012056f
C708 B.n459 VSUBS 0.012056f
C709 B.n460 VSUBS 0.012056f
C710 B.n461 VSUBS 0.012056f
C711 B.n462 VSUBS 0.012056f
C712 B.n463 VSUBS 0.012056f
C713 B.n464 VSUBS 0.012056f
C714 B.n465 VSUBS 0.012056f
C715 B.n466 VSUBS 0.012056f
C716 B.n467 VSUBS 0.012056f
C717 B.n468 VSUBS 0.012056f
C718 B.n469 VSUBS 0.012056f
C719 B.n470 VSUBS 0.012056f
C720 B.n471 VSUBS 0.012056f
C721 B.n472 VSUBS 0.012056f
C722 B.n473 VSUBS 0.012056f
C723 B.n474 VSUBS 0.012056f
C724 B.n475 VSUBS 0.012056f
C725 B.n476 VSUBS 0.012056f
C726 B.n477 VSUBS 0.012056f
C727 B.n478 VSUBS 0.012056f
C728 B.n479 VSUBS 0.012056f
C729 B.n480 VSUBS 0.012056f
C730 B.n481 VSUBS 0.012056f
C731 B.n482 VSUBS 0.012056f
C732 B.n483 VSUBS 0.012056f
C733 B.n484 VSUBS 0.012056f
C734 B.n485 VSUBS 0.012056f
C735 B.n486 VSUBS 0.012056f
C736 B.n487 VSUBS 0.012056f
C737 B.n488 VSUBS 0.012056f
C738 B.n489 VSUBS 0.012056f
C739 B.n490 VSUBS 0.012056f
C740 B.n491 VSUBS 0.012056f
C741 B.n492 VSUBS 0.012056f
C742 B.n493 VSUBS 0.012056f
C743 B.n494 VSUBS 0.012056f
C744 B.n495 VSUBS 0.012056f
C745 B.n496 VSUBS 0.012056f
C746 B.n497 VSUBS 0.012056f
C747 B.n498 VSUBS 0.012056f
C748 B.n499 VSUBS 0.012056f
C749 B.n500 VSUBS 0.012056f
C750 B.n501 VSUBS 0.012056f
C751 B.n502 VSUBS 0.012056f
C752 B.n503 VSUBS 0.012056f
C753 B.n504 VSUBS 0.012056f
C754 B.n505 VSUBS 0.012056f
C755 B.n506 VSUBS 0.012056f
C756 B.n507 VSUBS 0.012056f
C757 B.n508 VSUBS 0.012056f
C758 B.n509 VSUBS 0.012056f
C759 B.n510 VSUBS 0.012056f
C760 B.n511 VSUBS 0.012056f
C761 B.n512 VSUBS 0.012056f
C762 B.n513 VSUBS 0.012056f
C763 B.n514 VSUBS 0.012056f
C764 B.n515 VSUBS 0.012056f
C765 B.n516 VSUBS 0.012056f
C766 B.n517 VSUBS 0.012056f
C767 B.n518 VSUBS 0.012056f
C768 B.n519 VSUBS 0.012056f
C769 B.n520 VSUBS 0.012056f
C770 B.n521 VSUBS 0.012056f
C771 B.n522 VSUBS 0.012056f
C772 B.n523 VSUBS 0.012056f
C773 B.n524 VSUBS 0.012056f
C774 B.n525 VSUBS 0.012056f
C775 B.n526 VSUBS 0.012056f
C776 B.n527 VSUBS 0.012056f
C777 B.n528 VSUBS 0.012056f
C778 B.n529 VSUBS 0.012056f
C779 B.n530 VSUBS 0.012056f
C780 B.n531 VSUBS 0.012056f
C781 B.n532 VSUBS 0.012056f
C782 B.n533 VSUBS 0.012056f
C783 B.n534 VSUBS 0.012056f
C784 B.n535 VSUBS 0.012056f
C785 B.n536 VSUBS 0.012056f
C786 B.n537 VSUBS 0.012056f
C787 B.n538 VSUBS 0.012056f
C788 B.n539 VSUBS 0.012056f
C789 B.n540 VSUBS 0.012056f
C790 B.n541 VSUBS 0.012056f
C791 B.n542 VSUBS 0.012056f
C792 B.n543 VSUBS 0.012056f
C793 B.n544 VSUBS 0.012056f
C794 B.n545 VSUBS 0.012056f
C795 B.n546 VSUBS 0.012056f
C796 B.n547 VSUBS 0.012056f
C797 B.n548 VSUBS 0.012056f
C798 B.n549 VSUBS 0.012056f
C799 B.n550 VSUBS 0.012056f
C800 B.n551 VSUBS 0.012056f
C801 B.n552 VSUBS 0.012056f
C802 B.n553 VSUBS 0.012056f
C803 B.n554 VSUBS 0.012056f
C804 B.n555 VSUBS 0.012056f
C805 B.n556 VSUBS 0.012056f
C806 B.n557 VSUBS 0.012056f
C807 B.n558 VSUBS 0.012056f
C808 B.n559 VSUBS 0.012056f
C809 B.n560 VSUBS 0.012056f
C810 B.n561 VSUBS 0.012056f
C811 B.n562 VSUBS 0.012056f
C812 B.n563 VSUBS 0.012056f
C813 B.n564 VSUBS 0.012056f
C814 B.n565 VSUBS 0.012056f
C815 B.n566 VSUBS 0.012056f
C816 B.n567 VSUBS 0.012056f
C817 B.n568 VSUBS 0.012056f
C818 B.n569 VSUBS 0.012056f
C819 B.n570 VSUBS 0.012056f
C820 B.n571 VSUBS 0.012056f
C821 B.n572 VSUBS 0.012056f
C822 B.n573 VSUBS 0.012056f
C823 B.n574 VSUBS 0.012056f
C824 B.n575 VSUBS 0.012056f
C825 B.n576 VSUBS 0.012056f
C826 B.n577 VSUBS 0.012056f
C827 B.n578 VSUBS 0.012056f
C828 B.n579 VSUBS 0.012056f
C829 B.n580 VSUBS 0.012056f
C830 B.n581 VSUBS 0.012056f
C831 B.n582 VSUBS 0.012056f
C832 B.n583 VSUBS 0.012056f
C833 B.n584 VSUBS 0.012056f
C834 B.n585 VSUBS 0.012056f
C835 B.n586 VSUBS 0.012056f
C836 B.n587 VSUBS 0.012056f
C837 B.n588 VSUBS 0.012056f
C838 B.n589 VSUBS 0.012056f
C839 B.n590 VSUBS 0.012056f
C840 B.n591 VSUBS 0.012056f
C841 B.n592 VSUBS 0.012056f
C842 B.n593 VSUBS 0.012056f
C843 B.n594 VSUBS 0.012056f
C844 B.n595 VSUBS 0.012056f
C845 B.n596 VSUBS 0.012056f
C846 B.n597 VSUBS 0.012056f
C847 B.n598 VSUBS 0.012056f
C848 B.n599 VSUBS 0.012056f
C849 B.n600 VSUBS 0.012056f
C850 B.n601 VSUBS 0.012056f
C851 B.n602 VSUBS 0.012056f
C852 B.n603 VSUBS 0.012056f
C853 B.n604 VSUBS 0.012056f
C854 B.n605 VSUBS 0.012056f
C855 B.n606 VSUBS 0.012056f
C856 B.n607 VSUBS 0.012056f
C857 B.n608 VSUBS 0.012056f
C858 B.n609 VSUBS 0.012056f
C859 B.n610 VSUBS 0.012056f
C860 B.n611 VSUBS 0.012056f
C861 B.n612 VSUBS 0.012056f
C862 B.n613 VSUBS 0.012056f
C863 B.n614 VSUBS 0.012056f
C864 B.n615 VSUBS 0.012056f
C865 B.n616 VSUBS 0.012056f
C866 B.n617 VSUBS 0.012056f
C867 B.n618 VSUBS 0.012056f
C868 B.n619 VSUBS 0.012056f
C869 B.n620 VSUBS 0.012056f
C870 B.n621 VSUBS 0.012056f
C871 B.n622 VSUBS 0.012056f
C872 B.n623 VSUBS 0.012056f
C873 B.n624 VSUBS 0.012056f
C874 B.n625 VSUBS 0.012056f
C875 B.n626 VSUBS 0.012056f
C876 B.n627 VSUBS 0.012056f
C877 B.n628 VSUBS 0.012056f
C878 B.n629 VSUBS 0.012056f
C879 B.n630 VSUBS 0.012056f
C880 B.n631 VSUBS 0.012056f
C881 B.n632 VSUBS 0.012056f
C882 B.n633 VSUBS 0.012056f
C883 B.n634 VSUBS 0.012056f
C884 B.n635 VSUBS 0.012056f
C885 B.n636 VSUBS 0.012056f
C886 B.n637 VSUBS 0.012056f
C887 B.n638 VSUBS 0.012056f
C888 B.n639 VSUBS 0.012056f
C889 B.n640 VSUBS 0.012056f
C890 B.n641 VSUBS 0.012056f
C891 B.n642 VSUBS 0.012056f
C892 B.n643 VSUBS 0.012056f
C893 B.n644 VSUBS 0.012056f
C894 B.n645 VSUBS 0.012056f
C895 B.n646 VSUBS 0.012056f
C896 B.n647 VSUBS 0.012056f
C897 B.n648 VSUBS 0.012056f
C898 B.n649 VSUBS 0.012056f
C899 B.n650 VSUBS 0.012056f
C900 B.n651 VSUBS 0.012056f
C901 B.n652 VSUBS 0.012056f
C902 B.n653 VSUBS 0.012056f
C903 B.n654 VSUBS 0.012056f
C904 B.n655 VSUBS 0.012056f
C905 B.n656 VSUBS 0.012056f
C906 B.n657 VSUBS 0.012056f
C907 B.n658 VSUBS 0.029353f
C908 B.n659 VSUBS 0.030218f
C909 B.n660 VSUBS 0.028905f
C910 B.n661 VSUBS 0.012056f
C911 B.n662 VSUBS 0.012056f
C912 B.n663 VSUBS 0.012056f
C913 B.n664 VSUBS 0.012056f
C914 B.n665 VSUBS 0.012056f
C915 B.n666 VSUBS 0.012056f
C916 B.n667 VSUBS 0.012056f
C917 B.n668 VSUBS 0.012056f
C918 B.n669 VSUBS 0.012056f
C919 B.n670 VSUBS 0.012056f
C920 B.n671 VSUBS 0.012056f
C921 B.n672 VSUBS 0.012056f
C922 B.n673 VSUBS 0.012056f
C923 B.n674 VSUBS 0.012056f
C924 B.n675 VSUBS 0.012056f
C925 B.n676 VSUBS 0.012056f
C926 B.n677 VSUBS 0.012056f
C927 B.n678 VSUBS 0.012056f
C928 B.n679 VSUBS 0.012056f
C929 B.n680 VSUBS 0.012056f
C930 B.n681 VSUBS 0.012056f
C931 B.n682 VSUBS 0.012056f
C932 B.n683 VSUBS 0.012056f
C933 B.n684 VSUBS 0.012056f
C934 B.n685 VSUBS 0.012056f
C935 B.n686 VSUBS 0.012056f
C936 B.n687 VSUBS 0.012056f
C937 B.n688 VSUBS 0.012056f
C938 B.n689 VSUBS 0.012056f
C939 B.n690 VSUBS 0.012056f
C940 B.n691 VSUBS 0.008333f
C941 B.n692 VSUBS 0.027932f
C942 B.n693 VSUBS 0.009751f
C943 B.n694 VSUBS 0.012056f
C944 B.n695 VSUBS 0.012056f
C945 B.n696 VSUBS 0.012056f
C946 B.n697 VSUBS 0.012056f
C947 B.n698 VSUBS 0.012056f
C948 B.n699 VSUBS 0.012056f
C949 B.n700 VSUBS 0.012056f
C950 B.n701 VSUBS 0.012056f
C951 B.n702 VSUBS 0.012056f
C952 B.n703 VSUBS 0.012056f
C953 B.n704 VSUBS 0.012056f
C954 B.n705 VSUBS 0.009751f
C955 B.n706 VSUBS 0.012056f
C956 B.n707 VSUBS 0.012056f
C957 B.n708 VSUBS 0.012056f
C958 B.n709 VSUBS 0.012056f
C959 B.n710 VSUBS 0.012056f
C960 B.n711 VSUBS 0.012056f
C961 B.n712 VSUBS 0.012056f
C962 B.n713 VSUBS 0.012056f
C963 B.n714 VSUBS 0.012056f
C964 B.n715 VSUBS 0.012056f
C965 B.n716 VSUBS 0.012056f
C966 B.n717 VSUBS 0.012056f
C967 B.n718 VSUBS 0.012056f
C968 B.n719 VSUBS 0.012056f
C969 B.n720 VSUBS 0.012056f
C970 B.n721 VSUBS 0.012056f
C971 B.n722 VSUBS 0.012056f
C972 B.n723 VSUBS 0.012056f
C973 B.n724 VSUBS 0.012056f
C974 B.n725 VSUBS 0.012056f
C975 B.n726 VSUBS 0.012056f
C976 B.n727 VSUBS 0.012056f
C977 B.n728 VSUBS 0.012056f
C978 B.n729 VSUBS 0.012056f
C979 B.n730 VSUBS 0.012056f
C980 B.n731 VSUBS 0.012056f
C981 B.n732 VSUBS 0.012056f
C982 B.n733 VSUBS 0.012056f
C983 B.n734 VSUBS 0.012056f
C984 B.n735 VSUBS 0.012056f
C985 B.n736 VSUBS 0.012056f
C986 B.n737 VSUBS 0.012056f
C987 B.n738 VSUBS 0.030218f
C988 B.n739 VSUBS 0.030218f
C989 B.n740 VSUBS 0.029353f
C990 B.n741 VSUBS 0.012056f
C991 B.n742 VSUBS 0.012056f
C992 B.n743 VSUBS 0.012056f
C993 B.n744 VSUBS 0.012056f
C994 B.n745 VSUBS 0.012056f
C995 B.n746 VSUBS 0.012056f
C996 B.n747 VSUBS 0.012056f
C997 B.n748 VSUBS 0.012056f
C998 B.n749 VSUBS 0.012056f
C999 B.n750 VSUBS 0.012056f
C1000 B.n751 VSUBS 0.012056f
C1001 B.n752 VSUBS 0.012056f
C1002 B.n753 VSUBS 0.012056f
C1003 B.n754 VSUBS 0.012056f
C1004 B.n755 VSUBS 0.012056f
C1005 B.n756 VSUBS 0.012056f
C1006 B.n757 VSUBS 0.012056f
C1007 B.n758 VSUBS 0.012056f
C1008 B.n759 VSUBS 0.012056f
C1009 B.n760 VSUBS 0.012056f
C1010 B.n761 VSUBS 0.012056f
C1011 B.n762 VSUBS 0.012056f
C1012 B.n763 VSUBS 0.012056f
C1013 B.n764 VSUBS 0.012056f
C1014 B.n765 VSUBS 0.012056f
C1015 B.n766 VSUBS 0.012056f
C1016 B.n767 VSUBS 0.012056f
C1017 B.n768 VSUBS 0.012056f
C1018 B.n769 VSUBS 0.012056f
C1019 B.n770 VSUBS 0.012056f
C1020 B.n771 VSUBS 0.012056f
C1021 B.n772 VSUBS 0.012056f
C1022 B.n773 VSUBS 0.012056f
C1023 B.n774 VSUBS 0.012056f
C1024 B.n775 VSUBS 0.012056f
C1025 B.n776 VSUBS 0.012056f
C1026 B.n777 VSUBS 0.012056f
C1027 B.n778 VSUBS 0.012056f
C1028 B.n779 VSUBS 0.012056f
C1029 B.n780 VSUBS 0.012056f
C1030 B.n781 VSUBS 0.012056f
C1031 B.n782 VSUBS 0.012056f
C1032 B.n783 VSUBS 0.012056f
C1033 B.n784 VSUBS 0.012056f
C1034 B.n785 VSUBS 0.012056f
C1035 B.n786 VSUBS 0.012056f
C1036 B.n787 VSUBS 0.012056f
C1037 B.n788 VSUBS 0.012056f
C1038 B.n789 VSUBS 0.012056f
C1039 B.n790 VSUBS 0.012056f
C1040 B.n791 VSUBS 0.012056f
C1041 B.n792 VSUBS 0.012056f
C1042 B.n793 VSUBS 0.012056f
C1043 B.n794 VSUBS 0.012056f
C1044 B.n795 VSUBS 0.012056f
C1045 B.n796 VSUBS 0.012056f
C1046 B.n797 VSUBS 0.012056f
C1047 B.n798 VSUBS 0.012056f
C1048 B.n799 VSUBS 0.012056f
C1049 B.n800 VSUBS 0.012056f
C1050 B.n801 VSUBS 0.012056f
C1051 B.n802 VSUBS 0.012056f
C1052 B.n803 VSUBS 0.012056f
C1053 B.n804 VSUBS 0.012056f
C1054 B.n805 VSUBS 0.012056f
C1055 B.n806 VSUBS 0.012056f
C1056 B.n807 VSUBS 0.012056f
C1057 B.n808 VSUBS 0.012056f
C1058 B.n809 VSUBS 0.012056f
C1059 B.n810 VSUBS 0.012056f
C1060 B.n811 VSUBS 0.012056f
C1061 B.n812 VSUBS 0.012056f
C1062 B.n813 VSUBS 0.012056f
C1063 B.n814 VSUBS 0.012056f
C1064 B.n815 VSUBS 0.012056f
C1065 B.n816 VSUBS 0.012056f
C1066 B.n817 VSUBS 0.012056f
C1067 B.n818 VSUBS 0.012056f
C1068 B.n819 VSUBS 0.012056f
C1069 B.n820 VSUBS 0.012056f
C1070 B.n821 VSUBS 0.012056f
C1071 B.n822 VSUBS 0.012056f
C1072 B.n823 VSUBS 0.012056f
C1073 B.n824 VSUBS 0.012056f
C1074 B.n825 VSUBS 0.012056f
C1075 B.n826 VSUBS 0.012056f
C1076 B.n827 VSUBS 0.012056f
C1077 B.n828 VSUBS 0.012056f
C1078 B.n829 VSUBS 0.012056f
C1079 B.n830 VSUBS 0.012056f
C1080 B.n831 VSUBS 0.012056f
C1081 B.n832 VSUBS 0.012056f
C1082 B.n833 VSUBS 0.012056f
C1083 B.n834 VSUBS 0.012056f
C1084 B.n835 VSUBS 0.012056f
C1085 B.n836 VSUBS 0.012056f
C1086 B.n837 VSUBS 0.012056f
C1087 B.n838 VSUBS 0.012056f
C1088 B.n839 VSUBS 0.012056f
C1089 B.n840 VSUBS 0.012056f
C1090 B.n841 VSUBS 0.012056f
C1091 B.n842 VSUBS 0.012056f
C1092 B.n843 VSUBS 0.012056f
C1093 B.n844 VSUBS 0.012056f
C1094 B.n845 VSUBS 0.012056f
C1095 B.n846 VSUBS 0.012056f
C1096 B.n847 VSUBS 0.012056f
C1097 B.n848 VSUBS 0.012056f
C1098 B.n849 VSUBS 0.012056f
C1099 B.n850 VSUBS 0.012056f
C1100 B.n851 VSUBS 0.012056f
C1101 B.n852 VSUBS 0.012056f
C1102 B.n853 VSUBS 0.012056f
C1103 B.n854 VSUBS 0.012056f
C1104 B.n855 VSUBS 0.012056f
C1105 B.n856 VSUBS 0.012056f
C1106 B.n857 VSUBS 0.012056f
C1107 B.n858 VSUBS 0.012056f
C1108 B.n859 VSUBS 0.027299f
C1109 VDD2.n0 VSUBS 0.039492f
C1110 VDD2.n1 VSUBS 0.036219f
C1111 VDD2.n2 VSUBS 0.019463f
C1112 VDD2.n3 VSUBS 0.046002f
C1113 VDD2.n4 VSUBS 0.020607f
C1114 VDD2.n5 VSUBS 0.036219f
C1115 VDD2.n6 VSUBS 0.019463f
C1116 VDD2.n7 VSUBS 0.034502f
C1117 VDD2.n8 VSUBS 0.029221f
C1118 VDD2.t9 VSUBS 0.099297f
C1119 VDD2.n9 VSUBS 0.153319f
C1120 VDD2.n10 VSUBS 0.716218f
C1121 VDD2.n11 VSUBS 0.019463f
C1122 VDD2.n12 VSUBS 0.020607f
C1123 VDD2.n13 VSUBS 0.046002f
C1124 VDD2.n14 VSUBS 0.046002f
C1125 VDD2.n15 VSUBS 0.020607f
C1126 VDD2.n16 VSUBS 0.019463f
C1127 VDD2.n17 VSUBS 0.036219f
C1128 VDD2.n18 VSUBS 0.036219f
C1129 VDD2.n19 VSUBS 0.019463f
C1130 VDD2.n20 VSUBS 0.020607f
C1131 VDD2.n21 VSUBS 0.046002f
C1132 VDD2.n22 VSUBS 0.110328f
C1133 VDD2.n23 VSUBS 0.020607f
C1134 VDD2.n24 VSUBS 0.019463f
C1135 VDD2.n25 VSUBS 0.085203f
C1136 VDD2.n26 VSUBS 0.111593f
C1137 VDD2.t0 VSUBS 0.15198f
C1138 VDD2.t1 VSUBS 0.15198f
C1139 VDD2.n27 VSUBS 0.972723f
C1140 VDD2.n28 VSUBS 1.50961f
C1141 VDD2.t3 VSUBS 0.15198f
C1142 VDD2.t4 VSUBS 0.15198f
C1143 VDD2.n29 VSUBS 1.00518f
C1144 VDD2.n30 VSUBS 4.70948f
C1145 VDD2.n31 VSUBS 0.039492f
C1146 VDD2.n32 VSUBS 0.036219f
C1147 VDD2.n33 VSUBS 0.019463f
C1148 VDD2.n34 VSUBS 0.046002f
C1149 VDD2.n35 VSUBS 0.020607f
C1150 VDD2.n36 VSUBS 0.036219f
C1151 VDD2.n37 VSUBS 0.019463f
C1152 VDD2.n38 VSUBS 0.034502f
C1153 VDD2.n39 VSUBS 0.029221f
C1154 VDD2.t6 VSUBS 0.099297f
C1155 VDD2.n40 VSUBS 0.153319f
C1156 VDD2.n41 VSUBS 0.716218f
C1157 VDD2.n42 VSUBS 0.019463f
C1158 VDD2.n43 VSUBS 0.020607f
C1159 VDD2.n44 VSUBS 0.046002f
C1160 VDD2.n45 VSUBS 0.046002f
C1161 VDD2.n46 VSUBS 0.020607f
C1162 VDD2.n47 VSUBS 0.019463f
C1163 VDD2.n48 VSUBS 0.036219f
C1164 VDD2.n49 VSUBS 0.036219f
C1165 VDD2.n50 VSUBS 0.019463f
C1166 VDD2.n51 VSUBS 0.020607f
C1167 VDD2.n52 VSUBS 0.046002f
C1168 VDD2.n53 VSUBS 0.110328f
C1169 VDD2.n54 VSUBS 0.020607f
C1170 VDD2.n55 VSUBS 0.019463f
C1171 VDD2.n56 VSUBS 0.085203f
C1172 VDD2.n57 VSUBS 0.080479f
C1173 VDD2.n58 VSUBS 4.05361f
C1174 VDD2.t7 VSUBS 0.15198f
C1175 VDD2.t8 VSUBS 0.15198f
C1176 VDD2.n59 VSUBS 0.972728f
C1177 VDD2.n60 VSUBS 1.07789f
C1178 VDD2.t2 VSUBS 0.15198f
C1179 VDD2.t5 VSUBS 0.15198f
C1180 VDD2.n61 VSUBS 1.00513f
C1181 VTAIL.t13 VSUBS 0.150759f
C1182 VTAIL.t14 VSUBS 0.150759f
C1183 VTAIL.n0 VSUBS 0.851127f
C1184 VTAIL.n1 VSUBS 1.18858f
C1185 VTAIL.n2 VSUBS 0.039175f
C1186 VTAIL.n3 VSUBS 0.035928f
C1187 VTAIL.n4 VSUBS 0.019306f
C1188 VTAIL.n5 VSUBS 0.045633f
C1189 VTAIL.n6 VSUBS 0.020442f
C1190 VTAIL.n7 VSUBS 0.035928f
C1191 VTAIL.n8 VSUBS 0.019306f
C1192 VTAIL.n9 VSUBS 0.034225f
C1193 VTAIL.n10 VSUBS 0.028986f
C1194 VTAIL.t7 VSUBS 0.0985f
C1195 VTAIL.n11 VSUBS 0.152088f
C1196 VTAIL.n12 VSUBS 0.710464f
C1197 VTAIL.n13 VSUBS 0.019306f
C1198 VTAIL.n14 VSUBS 0.020442f
C1199 VTAIL.n15 VSUBS 0.045633f
C1200 VTAIL.n16 VSUBS 0.045633f
C1201 VTAIL.n17 VSUBS 0.020442f
C1202 VTAIL.n18 VSUBS 0.019306f
C1203 VTAIL.n19 VSUBS 0.035928f
C1204 VTAIL.n20 VSUBS 0.035928f
C1205 VTAIL.n21 VSUBS 0.019306f
C1206 VTAIL.n22 VSUBS 0.020442f
C1207 VTAIL.n23 VSUBS 0.045633f
C1208 VTAIL.n24 VSUBS 0.109442f
C1209 VTAIL.n25 VSUBS 0.020442f
C1210 VTAIL.n26 VSUBS 0.019306f
C1211 VTAIL.n27 VSUBS 0.084519f
C1212 VTAIL.n28 VSUBS 0.055037f
C1213 VTAIL.n29 VSUBS 0.687705f
C1214 VTAIL.t4 VSUBS 0.150759f
C1215 VTAIL.t5 VSUBS 0.150759f
C1216 VTAIL.n30 VSUBS 0.851127f
C1217 VTAIL.n31 VSUBS 1.42835f
C1218 VTAIL.t3 VSUBS 0.150759f
C1219 VTAIL.t0 VSUBS 0.150759f
C1220 VTAIL.n32 VSUBS 0.851127f
C1221 VTAIL.n33 VSUBS 2.84753f
C1222 VTAIL.t9 VSUBS 0.150759f
C1223 VTAIL.t12 VSUBS 0.150759f
C1224 VTAIL.n34 VSUBS 0.851133f
C1225 VTAIL.n35 VSUBS 2.84752f
C1226 VTAIL.t10 VSUBS 0.150759f
C1227 VTAIL.t16 VSUBS 0.150759f
C1228 VTAIL.n36 VSUBS 0.851133f
C1229 VTAIL.n37 VSUBS 1.42834f
C1230 VTAIL.n38 VSUBS 0.039175f
C1231 VTAIL.n39 VSUBS 0.035928f
C1232 VTAIL.n40 VSUBS 0.019306f
C1233 VTAIL.n41 VSUBS 0.045633f
C1234 VTAIL.n42 VSUBS 0.020442f
C1235 VTAIL.n43 VSUBS 0.035928f
C1236 VTAIL.n44 VSUBS 0.019306f
C1237 VTAIL.n45 VSUBS 0.034225f
C1238 VTAIL.n46 VSUBS 0.028986f
C1239 VTAIL.t18 VSUBS 0.0985f
C1240 VTAIL.n47 VSUBS 0.152088f
C1241 VTAIL.n48 VSUBS 0.710464f
C1242 VTAIL.n49 VSUBS 0.019306f
C1243 VTAIL.n50 VSUBS 0.020442f
C1244 VTAIL.n51 VSUBS 0.045633f
C1245 VTAIL.n52 VSUBS 0.045633f
C1246 VTAIL.n53 VSUBS 0.020442f
C1247 VTAIL.n54 VSUBS 0.019306f
C1248 VTAIL.n55 VSUBS 0.035928f
C1249 VTAIL.n56 VSUBS 0.035928f
C1250 VTAIL.n57 VSUBS 0.019306f
C1251 VTAIL.n58 VSUBS 0.020442f
C1252 VTAIL.n59 VSUBS 0.045633f
C1253 VTAIL.n60 VSUBS 0.109442f
C1254 VTAIL.n61 VSUBS 0.020442f
C1255 VTAIL.n62 VSUBS 0.019306f
C1256 VTAIL.n63 VSUBS 0.084519f
C1257 VTAIL.n64 VSUBS 0.055037f
C1258 VTAIL.n65 VSUBS 0.687705f
C1259 VTAIL.t8 VSUBS 0.150759f
C1260 VTAIL.t6 VSUBS 0.150759f
C1261 VTAIL.n66 VSUBS 0.851133f
C1262 VTAIL.n67 VSUBS 1.28214f
C1263 VTAIL.t19 VSUBS 0.150759f
C1264 VTAIL.t2 VSUBS 0.150759f
C1265 VTAIL.n68 VSUBS 0.851133f
C1266 VTAIL.n69 VSUBS 1.42834f
C1267 VTAIL.n70 VSUBS 0.039175f
C1268 VTAIL.n71 VSUBS 0.035928f
C1269 VTAIL.n72 VSUBS 0.019306f
C1270 VTAIL.n73 VSUBS 0.045633f
C1271 VTAIL.n74 VSUBS 0.020442f
C1272 VTAIL.n75 VSUBS 0.035928f
C1273 VTAIL.n76 VSUBS 0.019306f
C1274 VTAIL.n77 VSUBS 0.034225f
C1275 VTAIL.n78 VSUBS 0.028986f
C1276 VTAIL.t1 VSUBS 0.0985f
C1277 VTAIL.n79 VSUBS 0.152088f
C1278 VTAIL.n80 VSUBS 0.710464f
C1279 VTAIL.n81 VSUBS 0.019306f
C1280 VTAIL.n82 VSUBS 0.020442f
C1281 VTAIL.n83 VSUBS 0.045633f
C1282 VTAIL.n84 VSUBS 0.045633f
C1283 VTAIL.n85 VSUBS 0.020442f
C1284 VTAIL.n86 VSUBS 0.019306f
C1285 VTAIL.n87 VSUBS 0.035928f
C1286 VTAIL.n88 VSUBS 0.035928f
C1287 VTAIL.n89 VSUBS 0.019306f
C1288 VTAIL.n90 VSUBS 0.020442f
C1289 VTAIL.n91 VSUBS 0.045633f
C1290 VTAIL.n92 VSUBS 0.109442f
C1291 VTAIL.n93 VSUBS 0.020442f
C1292 VTAIL.n94 VSUBS 0.019306f
C1293 VTAIL.n95 VSUBS 0.084519f
C1294 VTAIL.n96 VSUBS 0.055037f
C1295 VTAIL.n97 VSUBS 1.85189f
C1296 VTAIL.n98 VSUBS 0.039175f
C1297 VTAIL.n99 VSUBS 0.035928f
C1298 VTAIL.n100 VSUBS 0.019306f
C1299 VTAIL.n101 VSUBS 0.045633f
C1300 VTAIL.n102 VSUBS 0.020442f
C1301 VTAIL.n103 VSUBS 0.035928f
C1302 VTAIL.n104 VSUBS 0.019306f
C1303 VTAIL.n105 VSUBS 0.034225f
C1304 VTAIL.n106 VSUBS 0.028986f
C1305 VTAIL.t11 VSUBS 0.0985f
C1306 VTAIL.n107 VSUBS 0.152088f
C1307 VTAIL.n108 VSUBS 0.710464f
C1308 VTAIL.n109 VSUBS 0.019306f
C1309 VTAIL.n110 VSUBS 0.020442f
C1310 VTAIL.n111 VSUBS 0.045633f
C1311 VTAIL.n112 VSUBS 0.045633f
C1312 VTAIL.n113 VSUBS 0.020442f
C1313 VTAIL.n114 VSUBS 0.019306f
C1314 VTAIL.n115 VSUBS 0.035928f
C1315 VTAIL.n116 VSUBS 0.035928f
C1316 VTAIL.n117 VSUBS 0.019306f
C1317 VTAIL.n118 VSUBS 0.020442f
C1318 VTAIL.n119 VSUBS 0.045633f
C1319 VTAIL.n120 VSUBS 0.109442f
C1320 VTAIL.n121 VSUBS 0.020442f
C1321 VTAIL.n122 VSUBS 0.019306f
C1322 VTAIL.n123 VSUBS 0.084519f
C1323 VTAIL.n124 VSUBS 0.055037f
C1324 VTAIL.n125 VSUBS 1.85189f
C1325 VTAIL.t15 VSUBS 0.150759f
C1326 VTAIL.t17 VSUBS 0.150759f
C1327 VTAIL.n126 VSUBS 0.851127f
C1328 VTAIL.n127 VSUBS 1.12071f
C1329 VN.t5 VSUBS 1.67192f
C1330 VN.n0 VSUBS 0.741573f
C1331 VN.n1 VSUBS 0.032487f
C1332 VN.n2 VSUBS 0.063415f
C1333 VN.n3 VSUBS 0.032487f
C1334 VN.n4 VSUBS 0.059352f
C1335 VN.n5 VSUBS 0.032487f
C1336 VN.n6 VSUBS 0.064221f
C1337 VN.n7 VSUBS 0.032487f
C1338 VN.n8 VSUBS 0.060548f
C1339 VN.n9 VSUBS 0.032487f
C1340 VN.t8 VSUBS 1.67192f
C1341 VN.n10 VSUBS 0.064872f
C1342 VN.n11 VSUBS 0.032487f
C1343 VN.n12 VSUBS 0.060548f
C1344 VN.t0 VSUBS 2.08723f
C1345 VN.n13 VSUBS 0.713624f
C1346 VN.t9 VSUBS 1.67192f
C1347 VN.n14 VSUBS 0.727461f
C1348 VN.n15 VSUBS 0.031851f
C1349 VN.n16 VSUBS 0.41275f
C1350 VN.n17 VSUBS 0.032487f
C1351 VN.n18 VSUBS 0.032487f
C1352 VN.n19 VSUBS 0.060548f
C1353 VN.n20 VSUBS 0.064221f
C1354 VN.n21 VSUBS 0.026305f
C1355 VN.n22 VSUBS 0.032487f
C1356 VN.n23 VSUBS 0.032487f
C1357 VN.n24 VSUBS 0.032487f
C1358 VN.n25 VSUBS 0.060548f
C1359 VN.n26 VSUBS 0.060548f
C1360 VN.n27 VSUBS 0.655183f
C1361 VN.n28 VSUBS 0.032487f
C1362 VN.n29 VSUBS 0.032487f
C1363 VN.n30 VSUBS 0.032487f
C1364 VN.n31 VSUBS 0.060548f
C1365 VN.n32 VSUBS 0.064872f
C1366 VN.n33 VSUBS 0.026305f
C1367 VN.n34 VSUBS 0.032487f
C1368 VN.n35 VSUBS 0.032487f
C1369 VN.n36 VSUBS 0.032487f
C1370 VN.n37 VSUBS 0.060548f
C1371 VN.n38 VSUBS 0.060548f
C1372 VN.t6 VSUBS 1.67192f
C1373 VN.n39 VSUBS 0.624528f
C1374 VN.n40 VSUBS 0.031851f
C1375 VN.n41 VSUBS 0.032487f
C1376 VN.n42 VSUBS 0.032487f
C1377 VN.n43 VSUBS 0.032487f
C1378 VN.n44 VSUBS 0.060548f
C1379 VN.n45 VSUBS 0.065343f
C1380 VN.n46 VSUBS 0.02664f
C1381 VN.n47 VSUBS 0.032487f
C1382 VN.n48 VSUBS 0.032487f
C1383 VN.n49 VSUBS 0.032487f
C1384 VN.n50 VSUBS 0.060548f
C1385 VN.n51 VSUBS 0.060548f
C1386 VN.n52 VSUBS 0.033046f
C1387 VN.n53 VSUBS 0.052433f
C1388 VN.n54 VSUBS 0.098649f
C1389 VN.t3 VSUBS 1.67192f
C1390 VN.n55 VSUBS 0.741573f
C1391 VN.n56 VSUBS 0.032487f
C1392 VN.n57 VSUBS 0.063415f
C1393 VN.n58 VSUBS 0.032487f
C1394 VN.n59 VSUBS 0.059352f
C1395 VN.n60 VSUBS 0.032487f
C1396 VN.t2 VSUBS 1.67192f
C1397 VN.n61 VSUBS 0.624528f
C1398 VN.n62 VSUBS 0.064221f
C1399 VN.n63 VSUBS 0.032487f
C1400 VN.n64 VSUBS 0.060548f
C1401 VN.n65 VSUBS 0.032487f
C1402 VN.t1 VSUBS 1.67192f
C1403 VN.n66 VSUBS 0.064872f
C1404 VN.n67 VSUBS 0.032487f
C1405 VN.n68 VSUBS 0.060548f
C1406 VN.t4 VSUBS 2.08723f
C1407 VN.n69 VSUBS 0.713624f
C1408 VN.t7 VSUBS 1.67192f
C1409 VN.n70 VSUBS 0.727461f
C1410 VN.n71 VSUBS 0.031851f
C1411 VN.n72 VSUBS 0.41275f
C1412 VN.n73 VSUBS 0.032487f
C1413 VN.n74 VSUBS 0.032487f
C1414 VN.n75 VSUBS 0.060548f
C1415 VN.n76 VSUBS 0.064221f
C1416 VN.n77 VSUBS 0.026305f
C1417 VN.n78 VSUBS 0.032487f
C1418 VN.n79 VSUBS 0.032487f
C1419 VN.n80 VSUBS 0.032487f
C1420 VN.n81 VSUBS 0.060548f
C1421 VN.n82 VSUBS 0.060548f
C1422 VN.n83 VSUBS 0.655183f
C1423 VN.n84 VSUBS 0.032487f
C1424 VN.n85 VSUBS 0.032487f
C1425 VN.n86 VSUBS 0.032487f
C1426 VN.n87 VSUBS 0.060548f
C1427 VN.n88 VSUBS 0.064872f
C1428 VN.n89 VSUBS 0.026305f
C1429 VN.n90 VSUBS 0.032487f
C1430 VN.n91 VSUBS 0.032487f
C1431 VN.n92 VSUBS 0.032487f
C1432 VN.n93 VSUBS 0.060548f
C1433 VN.n94 VSUBS 0.060548f
C1434 VN.n95 VSUBS 0.031851f
C1435 VN.n96 VSUBS 0.032487f
C1436 VN.n97 VSUBS 0.032487f
C1437 VN.n98 VSUBS 0.032487f
C1438 VN.n99 VSUBS 0.060548f
C1439 VN.n100 VSUBS 0.065343f
C1440 VN.n101 VSUBS 0.02664f
C1441 VN.n102 VSUBS 0.032487f
C1442 VN.n103 VSUBS 0.032487f
C1443 VN.n104 VSUBS 0.032487f
C1444 VN.n105 VSUBS 0.060548f
C1445 VN.n106 VSUBS 0.060548f
C1446 VN.n107 VSUBS 0.033046f
C1447 VN.n108 VSUBS 0.052433f
C1448 VN.n109 VSUBS 2.09132f
.ends

