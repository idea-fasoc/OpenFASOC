* NGSPICE file created from diff_pair_sample_0247.ext - technology: sky130A

.subckt diff_pair_sample_0247 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t3 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=2.33805 ps=14.5 w=14.17 l=3.67
X1 VTAIL.t3 VP.t0 VDD1.t7 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=2.33805 ps=14.5 w=14.17 l=3.67
X2 VTAIL.t14 VN.t1 VDD2.t2 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=5.5263 pd=29.12 as=2.33805 ps=14.5 w=14.17 l=3.67
X3 VTAIL.t13 VN.t2 VDD2.t1 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=2.33805 ps=14.5 w=14.17 l=3.67
X4 VTAIL.t4 VP.t1 VDD1.t6 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=5.5263 pd=29.12 as=2.33805 ps=14.5 w=14.17 l=3.67
X5 VDD2.t0 VN.t3 VTAIL.t12 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=5.5263 ps=29.12 w=14.17 l=3.67
X6 VTAIL.t5 VP.t2 VDD1.t5 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=2.33805 ps=14.5 w=14.17 l=3.67
X7 B.t11 B.t9 B.t10 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=5.5263 pd=29.12 as=0 ps=0 w=14.17 l=3.67
X8 VDD1.t4 VP.t3 VTAIL.t0 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=2.33805 ps=14.5 w=14.17 l=3.67
X9 B.t8 B.t6 B.t7 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=5.5263 pd=29.12 as=0 ps=0 w=14.17 l=3.67
X10 VDD1.t3 VP.t4 VTAIL.t1 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=5.5263 ps=29.12 w=14.17 l=3.67
X11 VDD2.t7 VN.t4 VTAIL.t11 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=5.5263 ps=29.12 w=14.17 l=3.67
X12 VTAIL.t2 VP.t5 VDD1.t2 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=5.5263 pd=29.12 as=2.33805 ps=14.5 w=14.17 l=3.67
X13 B.t5 B.t3 B.t4 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=5.5263 pd=29.12 as=0 ps=0 w=14.17 l=3.67
X14 VDD1.t1 VP.t6 VTAIL.t6 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=2.33805 ps=14.5 w=14.17 l=3.67
X15 VTAIL.t10 VN.t5 VDD2.t6 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=5.5263 pd=29.12 as=2.33805 ps=14.5 w=14.17 l=3.67
X16 VDD2.t5 VN.t6 VTAIL.t9 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=2.33805 ps=14.5 w=14.17 l=3.67
X17 VDD2.t4 VN.t7 VTAIL.t8 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=2.33805 ps=14.5 w=14.17 l=3.67
X18 B.t2 B.t0 B.t1 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=5.5263 pd=29.12 as=0 ps=0 w=14.17 l=3.67
X19 VDD1.t0 VP.t7 VTAIL.t7 w_n4970_n3802# sky130_fd_pr__pfet_01v8 ad=2.33805 pd=14.5 as=5.5263 ps=29.12 w=14.17 l=3.67
R0 VN.n65 VN.n34 161.3
R1 VN.n64 VN.n63 161.3
R2 VN.n62 VN.n35 161.3
R3 VN.n61 VN.n60 161.3
R4 VN.n59 VN.n36 161.3
R5 VN.n58 VN.n57 161.3
R6 VN.n56 VN.n37 161.3
R7 VN.n55 VN.n54 161.3
R8 VN.n53 VN.n38 161.3
R9 VN.n52 VN.n51 161.3
R10 VN.n50 VN.n39 161.3
R11 VN.n49 VN.n48 161.3
R12 VN.n47 VN.n40 161.3
R13 VN.n46 VN.n45 161.3
R14 VN.n44 VN.n41 161.3
R15 VN.n31 VN.n0 161.3
R16 VN.n30 VN.n29 161.3
R17 VN.n28 VN.n1 161.3
R18 VN.n27 VN.n26 161.3
R19 VN.n25 VN.n2 161.3
R20 VN.n24 VN.n23 161.3
R21 VN.n22 VN.n3 161.3
R22 VN.n21 VN.n20 161.3
R23 VN.n19 VN.n4 161.3
R24 VN.n18 VN.n17 161.3
R25 VN.n16 VN.n5 161.3
R26 VN.n15 VN.n14 161.3
R27 VN.n13 VN.n6 161.3
R28 VN.n12 VN.n11 161.3
R29 VN.n10 VN.n7 161.3
R30 VN.n9 VN.t5 125.162
R31 VN.n43 VN.t4 125.162
R32 VN.n32 VN.t3 93.0515
R33 VN.n20 VN.t2 93.0515
R34 VN.n8 VN.t7 93.0515
R35 VN.n66 VN.t1 93.0515
R36 VN.n54 VN.t6 93.0515
R37 VN.n42 VN.t0 93.0515
R38 VN VN.n67 57.8148
R39 VN.n33 VN.n32 57.7148
R40 VN.n67 VN.n66 57.7148
R41 VN.n9 VN.n8 50.4779
R42 VN.n43 VN.n42 50.4779
R43 VN.n14 VN.n13 40.4934
R44 VN.n14 VN.n5 40.4934
R45 VN.n26 VN.n25 40.4934
R46 VN.n26 VN.n1 40.4934
R47 VN.n48 VN.n47 40.4934
R48 VN.n48 VN.n39 40.4934
R49 VN.n60 VN.n59 40.4934
R50 VN.n60 VN.n35 40.4934
R51 VN.n8 VN.n7 24.4675
R52 VN.n12 VN.n7 24.4675
R53 VN.n13 VN.n12 24.4675
R54 VN.n18 VN.n5 24.4675
R55 VN.n19 VN.n18 24.4675
R56 VN.n20 VN.n19 24.4675
R57 VN.n20 VN.n3 24.4675
R58 VN.n24 VN.n3 24.4675
R59 VN.n25 VN.n24 24.4675
R60 VN.n30 VN.n1 24.4675
R61 VN.n31 VN.n30 24.4675
R62 VN.n32 VN.n31 24.4675
R63 VN.n47 VN.n46 24.4675
R64 VN.n46 VN.n41 24.4675
R65 VN.n42 VN.n41 24.4675
R66 VN.n59 VN.n58 24.4675
R67 VN.n58 VN.n37 24.4675
R68 VN.n54 VN.n37 24.4675
R69 VN.n54 VN.n53 24.4675
R70 VN.n53 VN.n52 24.4675
R71 VN.n52 VN.n39 24.4675
R72 VN.n66 VN.n65 24.4675
R73 VN.n65 VN.n64 24.4675
R74 VN.n64 VN.n35 24.4675
R75 VN.n44 VN.n43 2.5265
R76 VN.n10 VN.n9 2.5265
R77 VN.n67 VN.n34 0.417535
R78 VN.n33 VN.n0 0.417535
R79 VN VN.n33 0.394291
R80 VN.n63 VN.n34 0.189894
R81 VN.n63 VN.n62 0.189894
R82 VN.n62 VN.n61 0.189894
R83 VN.n61 VN.n36 0.189894
R84 VN.n57 VN.n36 0.189894
R85 VN.n57 VN.n56 0.189894
R86 VN.n56 VN.n55 0.189894
R87 VN.n55 VN.n38 0.189894
R88 VN.n51 VN.n38 0.189894
R89 VN.n51 VN.n50 0.189894
R90 VN.n50 VN.n49 0.189894
R91 VN.n49 VN.n40 0.189894
R92 VN.n45 VN.n40 0.189894
R93 VN.n45 VN.n44 0.189894
R94 VN.n11 VN.n10 0.189894
R95 VN.n11 VN.n6 0.189894
R96 VN.n15 VN.n6 0.189894
R97 VN.n16 VN.n15 0.189894
R98 VN.n17 VN.n16 0.189894
R99 VN.n17 VN.n4 0.189894
R100 VN.n21 VN.n4 0.189894
R101 VN.n22 VN.n21 0.189894
R102 VN.n23 VN.n22 0.189894
R103 VN.n23 VN.n2 0.189894
R104 VN.n27 VN.n2 0.189894
R105 VN.n28 VN.n27 0.189894
R106 VN.n29 VN.n28 0.189894
R107 VN.n29 VN.n0 0.189894
R108 VDD2.n2 VDD2.n1 71.1684
R109 VDD2.n2 VDD2.n0 71.1684
R110 VDD2 VDD2.n5 71.1656
R111 VDD2.n4 VDD2.n3 69.4996
R112 VDD2.n4 VDD2.n2 51.4481
R113 VDD2.n5 VDD2.t3 2.29443
R114 VDD2.n5 VDD2.t7 2.29443
R115 VDD2.n3 VDD2.t2 2.29443
R116 VDD2.n3 VDD2.t5 2.29443
R117 VDD2.n1 VDD2.t1 2.29443
R118 VDD2.n1 VDD2.t0 2.29443
R119 VDD2.n0 VDD2.t6 2.29443
R120 VDD2.n0 VDD2.t4 2.29443
R121 VDD2 VDD2.n4 1.78283
R122 VTAIL.n626 VTAIL.n554 756.745
R123 VTAIL.n74 VTAIL.n2 756.745
R124 VTAIL.n152 VTAIL.n80 756.745
R125 VTAIL.n232 VTAIL.n160 756.745
R126 VTAIL.n548 VTAIL.n476 756.745
R127 VTAIL.n468 VTAIL.n396 756.745
R128 VTAIL.n390 VTAIL.n318 756.745
R129 VTAIL.n310 VTAIL.n238 756.745
R130 VTAIL.n578 VTAIL.n577 585
R131 VTAIL.n583 VTAIL.n582 585
R132 VTAIL.n585 VTAIL.n584 585
R133 VTAIL.n574 VTAIL.n573 585
R134 VTAIL.n591 VTAIL.n590 585
R135 VTAIL.n593 VTAIL.n592 585
R136 VTAIL.n570 VTAIL.n569 585
R137 VTAIL.n600 VTAIL.n599 585
R138 VTAIL.n601 VTAIL.n568 585
R139 VTAIL.n603 VTAIL.n602 585
R140 VTAIL.n566 VTAIL.n565 585
R141 VTAIL.n609 VTAIL.n608 585
R142 VTAIL.n611 VTAIL.n610 585
R143 VTAIL.n562 VTAIL.n561 585
R144 VTAIL.n617 VTAIL.n616 585
R145 VTAIL.n619 VTAIL.n618 585
R146 VTAIL.n558 VTAIL.n557 585
R147 VTAIL.n625 VTAIL.n624 585
R148 VTAIL.n627 VTAIL.n626 585
R149 VTAIL.n26 VTAIL.n25 585
R150 VTAIL.n31 VTAIL.n30 585
R151 VTAIL.n33 VTAIL.n32 585
R152 VTAIL.n22 VTAIL.n21 585
R153 VTAIL.n39 VTAIL.n38 585
R154 VTAIL.n41 VTAIL.n40 585
R155 VTAIL.n18 VTAIL.n17 585
R156 VTAIL.n48 VTAIL.n47 585
R157 VTAIL.n49 VTAIL.n16 585
R158 VTAIL.n51 VTAIL.n50 585
R159 VTAIL.n14 VTAIL.n13 585
R160 VTAIL.n57 VTAIL.n56 585
R161 VTAIL.n59 VTAIL.n58 585
R162 VTAIL.n10 VTAIL.n9 585
R163 VTAIL.n65 VTAIL.n64 585
R164 VTAIL.n67 VTAIL.n66 585
R165 VTAIL.n6 VTAIL.n5 585
R166 VTAIL.n73 VTAIL.n72 585
R167 VTAIL.n75 VTAIL.n74 585
R168 VTAIL.n104 VTAIL.n103 585
R169 VTAIL.n109 VTAIL.n108 585
R170 VTAIL.n111 VTAIL.n110 585
R171 VTAIL.n100 VTAIL.n99 585
R172 VTAIL.n117 VTAIL.n116 585
R173 VTAIL.n119 VTAIL.n118 585
R174 VTAIL.n96 VTAIL.n95 585
R175 VTAIL.n126 VTAIL.n125 585
R176 VTAIL.n127 VTAIL.n94 585
R177 VTAIL.n129 VTAIL.n128 585
R178 VTAIL.n92 VTAIL.n91 585
R179 VTAIL.n135 VTAIL.n134 585
R180 VTAIL.n137 VTAIL.n136 585
R181 VTAIL.n88 VTAIL.n87 585
R182 VTAIL.n143 VTAIL.n142 585
R183 VTAIL.n145 VTAIL.n144 585
R184 VTAIL.n84 VTAIL.n83 585
R185 VTAIL.n151 VTAIL.n150 585
R186 VTAIL.n153 VTAIL.n152 585
R187 VTAIL.n184 VTAIL.n183 585
R188 VTAIL.n189 VTAIL.n188 585
R189 VTAIL.n191 VTAIL.n190 585
R190 VTAIL.n180 VTAIL.n179 585
R191 VTAIL.n197 VTAIL.n196 585
R192 VTAIL.n199 VTAIL.n198 585
R193 VTAIL.n176 VTAIL.n175 585
R194 VTAIL.n206 VTAIL.n205 585
R195 VTAIL.n207 VTAIL.n174 585
R196 VTAIL.n209 VTAIL.n208 585
R197 VTAIL.n172 VTAIL.n171 585
R198 VTAIL.n215 VTAIL.n214 585
R199 VTAIL.n217 VTAIL.n216 585
R200 VTAIL.n168 VTAIL.n167 585
R201 VTAIL.n223 VTAIL.n222 585
R202 VTAIL.n225 VTAIL.n224 585
R203 VTAIL.n164 VTAIL.n163 585
R204 VTAIL.n231 VTAIL.n230 585
R205 VTAIL.n233 VTAIL.n232 585
R206 VTAIL.n549 VTAIL.n548 585
R207 VTAIL.n547 VTAIL.n546 585
R208 VTAIL.n480 VTAIL.n479 585
R209 VTAIL.n541 VTAIL.n540 585
R210 VTAIL.n539 VTAIL.n538 585
R211 VTAIL.n484 VTAIL.n483 585
R212 VTAIL.n533 VTAIL.n532 585
R213 VTAIL.n531 VTAIL.n530 585
R214 VTAIL.n488 VTAIL.n487 585
R215 VTAIL.n525 VTAIL.n524 585
R216 VTAIL.n523 VTAIL.n490 585
R217 VTAIL.n522 VTAIL.n521 585
R218 VTAIL.n493 VTAIL.n491 585
R219 VTAIL.n516 VTAIL.n515 585
R220 VTAIL.n514 VTAIL.n513 585
R221 VTAIL.n497 VTAIL.n496 585
R222 VTAIL.n508 VTAIL.n507 585
R223 VTAIL.n506 VTAIL.n505 585
R224 VTAIL.n501 VTAIL.n500 585
R225 VTAIL.n469 VTAIL.n468 585
R226 VTAIL.n467 VTAIL.n466 585
R227 VTAIL.n400 VTAIL.n399 585
R228 VTAIL.n461 VTAIL.n460 585
R229 VTAIL.n459 VTAIL.n458 585
R230 VTAIL.n404 VTAIL.n403 585
R231 VTAIL.n453 VTAIL.n452 585
R232 VTAIL.n451 VTAIL.n450 585
R233 VTAIL.n408 VTAIL.n407 585
R234 VTAIL.n445 VTAIL.n444 585
R235 VTAIL.n443 VTAIL.n410 585
R236 VTAIL.n442 VTAIL.n441 585
R237 VTAIL.n413 VTAIL.n411 585
R238 VTAIL.n436 VTAIL.n435 585
R239 VTAIL.n434 VTAIL.n433 585
R240 VTAIL.n417 VTAIL.n416 585
R241 VTAIL.n428 VTAIL.n427 585
R242 VTAIL.n426 VTAIL.n425 585
R243 VTAIL.n421 VTAIL.n420 585
R244 VTAIL.n391 VTAIL.n390 585
R245 VTAIL.n389 VTAIL.n388 585
R246 VTAIL.n322 VTAIL.n321 585
R247 VTAIL.n383 VTAIL.n382 585
R248 VTAIL.n381 VTAIL.n380 585
R249 VTAIL.n326 VTAIL.n325 585
R250 VTAIL.n375 VTAIL.n374 585
R251 VTAIL.n373 VTAIL.n372 585
R252 VTAIL.n330 VTAIL.n329 585
R253 VTAIL.n367 VTAIL.n366 585
R254 VTAIL.n365 VTAIL.n332 585
R255 VTAIL.n364 VTAIL.n363 585
R256 VTAIL.n335 VTAIL.n333 585
R257 VTAIL.n358 VTAIL.n357 585
R258 VTAIL.n356 VTAIL.n355 585
R259 VTAIL.n339 VTAIL.n338 585
R260 VTAIL.n350 VTAIL.n349 585
R261 VTAIL.n348 VTAIL.n347 585
R262 VTAIL.n343 VTAIL.n342 585
R263 VTAIL.n311 VTAIL.n310 585
R264 VTAIL.n309 VTAIL.n308 585
R265 VTAIL.n242 VTAIL.n241 585
R266 VTAIL.n303 VTAIL.n302 585
R267 VTAIL.n301 VTAIL.n300 585
R268 VTAIL.n246 VTAIL.n245 585
R269 VTAIL.n295 VTAIL.n294 585
R270 VTAIL.n293 VTAIL.n292 585
R271 VTAIL.n250 VTAIL.n249 585
R272 VTAIL.n287 VTAIL.n286 585
R273 VTAIL.n285 VTAIL.n252 585
R274 VTAIL.n284 VTAIL.n283 585
R275 VTAIL.n255 VTAIL.n253 585
R276 VTAIL.n278 VTAIL.n277 585
R277 VTAIL.n276 VTAIL.n275 585
R278 VTAIL.n259 VTAIL.n258 585
R279 VTAIL.n270 VTAIL.n269 585
R280 VTAIL.n268 VTAIL.n267 585
R281 VTAIL.n263 VTAIL.n262 585
R282 VTAIL.n579 VTAIL.t12 329.036
R283 VTAIL.n27 VTAIL.t10 329.036
R284 VTAIL.n105 VTAIL.t7 329.036
R285 VTAIL.n185 VTAIL.t2 329.036
R286 VTAIL.n422 VTAIL.t4 329.036
R287 VTAIL.n344 VTAIL.t11 329.036
R288 VTAIL.n264 VTAIL.t14 329.036
R289 VTAIL.n502 VTAIL.t1 329.036
R290 VTAIL.n583 VTAIL.n577 171.744
R291 VTAIL.n584 VTAIL.n583 171.744
R292 VTAIL.n584 VTAIL.n573 171.744
R293 VTAIL.n591 VTAIL.n573 171.744
R294 VTAIL.n592 VTAIL.n591 171.744
R295 VTAIL.n592 VTAIL.n569 171.744
R296 VTAIL.n600 VTAIL.n569 171.744
R297 VTAIL.n601 VTAIL.n600 171.744
R298 VTAIL.n602 VTAIL.n601 171.744
R299 VTAIL.n602 VTAIL.n565 171.744
R300 VTAIL.n609 VTAIL.n565 171.744
R301 VTAIL.n610 VTAIL.n609 171.744
R302 VTAIL.n610 VTAIL.n561 171.744
R303 VTAIL.n617 VTAIL.n561 171.744
R304 VTAIL.n618 VTAIL.n617 171.744
R305 VTAIL.n618 VTAIL.n557 171.744
R306 VTAIL.n625 VTAIL.n557 171.744
R307 VTAIL.n626 VTAIL.n625 171.744
R308 VTAIL.n31 VTAIL.n25 171.744
R309 VTAIL.n32 VTAIL.n31 171.744
R310 VTAIL.n32 VTAIL.n21 171.744
R311 VTAIL.n39 VTAIL.n21 171.744
R312 VTAIL.n40 VTAIL.n39 171.744
R313 VTAIL.n40 VTAIL.n17 171.744
R314 VTAIL.n48 VTAIL.n17 171.744
R315 VTAIL.n49 VTAIL.n48 171.744
R316 VTAIL.n50 VTAIL.n49 171.744
R317 VTAIL.n50 VTAIL.n13 171.744
R318 VTAIL.n57 VTAIL.n13 171.744
R319 VTAIL.n58 VTAIL.n57 171.744
R320 VTAIL.n58 VTAIL.n9 171.744
R321 VTAIL.n65 VTAIL.n9 171.744
R322 VTAIL.n66 VTAIL.n65 171.744
R323 VTAIL.n66 VTAIL.n5 171.744
R324 VTAIL.n73 VTAIL.n5 171.744
R325 VTAIL.n74 VTAIL.n73 171.744
R326 VTAIL.n109 VTAIL.n103 171.744
R327 VTAIL.n110 VTAIL.n109 171.744
R328 VTAIL.n110 VTAIL.n99 171.744
R329 VTAIL.n117 VTAIL.n99 171.744
R330 VTAIL.n118 VTAIL.n117 171.744
R331 VTAIL.n118 VTAIL.n95 171.744
R332 VTAIL.n126 VTAIL.n95 171.744
R333 VTAIL.n127 VTAIL.n126 171.744
R334 VTAIL.n128 VTAIL.n127 171.744
R335 VTAIL.n128 VTAIL.n91 171.744
R336 VTAIL.n135 VTAIL.n91 171.744
R337 VTAIL.n136 VTAIL.n135 171.744
R338 VTAIL.n136 VTAIL.n87 171.744
R339 VTAIL.n143 VTAIL.n87 171.744
R340 VTAIL.n144 VTAIL.n143 171.744
R341 VTAIL.n144 VTAIL.n83 171.744
R342 VTAIL.n151 VTAIL.n83 171.744
R343 VTAIL.n152 VTAIL.n151 171.744
R344 VTAIL.n189 VTAIL.n183 171.744
R345 VTAIL.n190 VTAIL.n189 171.744
R346 VTAIL.n190 VTAIL.n179 171.744
R347 VTAIL.n197 VTAIL.n179 171.744
R348 VTAIL.n198 VTAIL.n197 171.744
R349 VTAIL.n198 VTAIL.n175 171.744
R350 VTAIL.n206 VTAIL.n175 171.744
R351 VTAIL.n207 VTAIL.n206 171.744
R352 VTAIL.n208 VTAIL.n207 171.744
R353 VTAIL.n208 VTAIL.n171 171.744
R354 VTAIL.n215 VTAIL.n171 171.744
R355 VTAIL.n216 VTAIL.n215 171.744
R356 VTAIL.n216 VTAIL.n167 171.744
R357 VTAIL.n223 VTAIL.n167 171.744
R358 VTAIL.n224 VTAIL.n223 171.744
R359 VTAIL.n224 VTAIL.n163 171.744
R360 VTAIL.n231 VTAIL.n163 171.744
R361 VTAIL.n232 VTAIL.n231 171.744
R362 VTAIL.n548 VTAIL.n547 171.744
R363 VTAIL.n547 VTAIL.n479 171.744
R364 VTAIL.n540 VTAIL.n479 171.744
R365 VTAIL.n540 VTAIL.n539 171.744
R366 VTAIL.n539 VTAIL.n483 171.744
R367 VTAIL.n532 VTAIL.n483 171.744
R368 VTAIL.n532 VTAIL.n531 171.744
R369 VTAIL.n531 VTAIL.n487 171.744
R370 VTAIL.n524 VTAIL.n487 171.744
R371 VTAIL.n524 VTAIL.n523 171.744
R372 VTAIL.n523 VTAIL.n522 171.744
R373 VTAIL.n522 VTAIL.n491 171.744
R374 VTAIL.n515 VTAIL.n491 171.744
R375 VTAIL.n515 VTAIL.n514 171.744
R376 VTAIL.n514 VTAIL.n496 171.744
R377 VTAIL.n507 VTAIL.n496 171.744
R378 VTAIL.n507 VTAIL.n506 171.744
R379 VTAIL.n506 VTAIL.n500 171.744
R380 VTAIL.n468 VTAIL.n467 171.744
R381 VTAIL.n467 VTAIL.n399 171.744
R382 VTAIL.n460 VTAIL.n399 171.744
R383 VTAIL.n460 VTAIL.n459 171.744
R384 VTAIL.n459 VTAIL.n403 171.744
R385 VTAIL.n452 VTAIL.n403 171.744
R386 VTAIL.n452 VTAIL.n451 171.744
R387 VTAIL.n451 VTAIL.n407 171.744
R388 VTAIL.n444 VTAIL.n407 171.744
R389 VTAIL.n444 VTAIL.n443 171.744
R390 VTAIL.n443 VTAIL.n442 171.744
R391 VTAIL.n442 VTAIL.n411 171.744
R392 VTAIL.n435 VTAIL.n411 171.744
R393 VTAIL.n435 VTAIL.n434 171.744
R394 VTAIL.n434 VTAIL.n416 171.744
R395 VTAIL.n427 VTAIL.n416 171.744
R396 VTAIL.n427 VTAIL.n426 171.744
R397 VTAIL.n426 VTAIL.n420 171.744
R398 VTAIL.n390 VTAIL.n389 171.744
R399 VTAIL.n389 VTAIL.n321 171.744
R400 VTAIL.n382 VTAIL.n321 171.744
R401 VTAIL.n382 VTAIL.n381 171.744
R402 VTAIL.n381 VTAIL.n325 171.744
R403 VTAIL.n374 VTAIL.n325 171.744
R404 VTAIL.n374 VTAIL.n373 171.744
R405 VTAIL.n373 VTAIL.n329 171.744
R406 VTAIL.n366 VTAIL.n329 171.744
R407 VTAIL.n366 VTAIL.n365 171.744
R408 VTAIL.n365 VTAIL.n364 171.744
R409 VTAIL.n364 VTAIL.n333 171.744
R410 VTAIL.n357 VTAIL.n333 171.744
R411 VTAIL.n357 VTAIL.n356 171.744
R412 VTAIL.n356 VTAIL.n338 171.744
R413 VTAIL.n349 VTAIL.n338 171.744
R414 VTAIL.n349 VTAIL.n348 171.744
R415 VTAIL.n348 VTAIL.n342 171.744
R416 VTAIL.n310 VTAIL.n309 171.744
R417 VTAIL.n309 VTAIL.n241 171.744
R418 VTAIL.n302 VTAIL.n241 171.744
R419 VTAIL.n302 VTAIL.n301 171.744
R420 VTAIL.n301 VTAIL.n245 171.744
R421 VTAIL.n294 VTAIL.n245 171.744
R422 VTAIL.n294 VTAIL.n293 171.744
R423 VTAIL.n293 VTAIL.n249 171.744
R424 VTAIL.n286 VTAIL.n249 171.744
R425 VTAIL.n286 VTAIL.n285 171.744
R426 VTAIL.n285 VTAIL.n284 171.744
R427 VTAIL.n284 VTAIL.n253 171.744
R428 VTAIL.n277 VTAIL.n253 171.744
R429 VTAIL.n277 VTAIL.n276 171.744
R430 VTAIL.n276 VTAIL.n258 171.744
R431 VTAIL.n269 VTAIL.n258 171.744
R432 VTAIL.n269 VTAIL.n268 171.744
R433 VTAIL.n268 VTAIL.n262 171.744
R434 VTAIL.t12 VTAIL.n577 85.8723
R435 VTAIL.t10 VTAIL.n25 85.8723
R436 VTAIL.t7 VTAIL.n103 85.8723
R437 VTAIL.t2 VTAIL.n183 85.8723
R438 VTAIL.t1 VTAIL.n500 85.8723
R439 VTAIL.t4 VTAIL.n420 85.8723
R440 VTAIL.t11 VTAIL.n342 85.8723
R441 VTAIL.t14 VTAIL.n262 85.8723
R442 VTAIL.n475 VTAIL.n474 52.8208
R443 VTAIL.n317 VTAIL.n316 52.8208
R444 VTAIL.n1 VTAIL.n0 52.8208
R445 VTAIL.n159 VTAIL.n158 52.8208
R446 VTAIL.n631 VTAIL.n630 30.052
R447 VTAIL.n79 VTAIL.n78 30.052
R448 VTAIL.n157 VTAIL.n156 30.052
R449 VTAIL.n237 VTAIL.n236 30.052
R450 VTAIL.n553 VTAIL.n552 30.052
R451 VTAIL.n473 VTAIL.n472 30.052
R452 VTAIL.n395 VTAIL.n394 30.052
R453 VTAIL.n315 VTAIL.n314 30.052
R454 VTAIL.n631 VTAIL.n553 28.0307
R455 VTAIL.n315 VTAIL.n237 28.0307
R456 VTAIL.n603 VTAIL.n568 13.1884
R457 VTAIL.n51 VTAIL.n16 13.1884
R458 VTAIL.n129 VTAIL.n94 13.1884
R459 VTAIL.n209 VTAIL.n174 13.1884
R460 VTAIL.n525 VTAIL.n490 13.1884
R461 VTAIL.n445 VTAIL.n410 13.1884
R462 VTAIL.n367 VTAIL.n332 13.1884
R463 VTAIL.n287 VTAIL.n252 13.1884
R464 VTAIL.n599 VTAIL.n598 12.8005
R465 VTAIL.n604 VTAIL.n566 12.8005
R466 VTAIL.n47 VTAIL.n46 12.8005
R467 VTAIL.n52 VTAIL.n14 12.8005
R468 VTAIL.n125 VTAIL.n124 12.8005
R469 VTAIL.n130 VTAIL.n92 12.8005
R470 VTAIL.n205 VTAIL.n204 12.8005
R471 VTAIL.n210 VTAIL.n172 12.8005
R472 VTAIL.n526 VTAIL.n488 12.8005
R473 VTAIL.n521 VTAIL.n492 12.8005
R474 VTAIL.n446 VTAIL.n408 12.8005
R475 VTAIL.n441 VTAIL.n412 12.8005
R476 VTAIL.n368 VTAIL.n330 12.8005
R477 VTAIL.n363 VTAIL.n334 12.8005
R478 VTAIL.n288 VTAIL.n250 12.8005
R479 VTAIL.n283 VTAIL.n254 12.8005
R480 VTAIL.n597 VTAIL.n570 12.0247
R481 VTAIL.n608 VTAIL.n607 12.0247
R482 VTAIL.n45 VTAIL.n18 12.0247
R483 VTAIL.n56 VTAIL.n55 12.0247
R484 VTAIL.n123 VTAIL.n96 12.0247
R485 VTAIL.n134 VTAIL.n133 12.0247
R486 VTAIL.n203 VTAIL.n176 12.0247
R487 VTAIL.n214 VTAIL.n213 12.0247
R488 VTAIL.n530 VTAIL.n529 12.0247
R489 VTAIL.n520 VTAIL.n493 12.0247
R490 VTAIL.n450 VTAIL.n449 12.0247
R491 VTAIL.n440 VTAIL.n413 12.0247
R492 VTAIL.n372 VTAIL.n371 12.0247
R493 VTAIL.n362 VTAIL.n335 12.0247
R494 VTAIL.n292 VTAIL.n291 12.0247
R495 VTAIL.n282 VTAIL.n255 12.0247
R496 VTAIL.n594 VTAIL.n593 11.249
R497 VTAIL.n611 VTAIL.n564 11.249
R498 VTAIL.n42 VTAIL.n41 11.249
R499 VTAIL.n59 VTAIL.n12 11.249
R500 VTAIL.n120 VTAIL.n119 11.249
R501 VTAIL.n137 VTAIL.n90 11.249
R502 VTAIL.n200 VTAIL.n199 11.249
R503 VTAIL.n217 VTAIL.n170 11.249
R504 VTAIL.n533 VTAIL.n486 11.249
R505 VTAIL.n517 VTAIL.n516 11.249
R506 VTAIL.n453 VTAIL.n406 11.249
R507 VTAIL.n437 VTAIL.n436 11.249
R508 VTAIL.n375 VTAIL.n328 11.249
R509 VTAIL.n359 VTAIL.n358 11.249
R510 VTAIL.n295 VTAIL.n248 11.249
R511 VTAIL.n279 VTAIL.n278 11.249
R512 VTAIL.n579 VTAIL.n578 10.7239
R513 VTAIL.n27 VTAIL.n26 10.7239
R514 VTAIL.n105 VTAIL.n104 10.7239
R515 VTAIL.n185 VTAIL.n184 10.7239
R516 VTAIL.n502 VTAIL.n501 10.7239
R517 VTAIL.n422 VTAIL.n421 10.7239
R518 VTAIL.n344 VTAIL.n343 10.7239
R519 VTAIL.n264 VTAIL.n263 10.7239
R520 VTAIL.n590 VTAIL.n572 10.4732
R521 VTAIL.n612 VTAIL.n562 10.4732
R522 VTAIL.n38 VTAIL.n20 10.4732
R523 VTAIL.n60 VTAIL.n10 10.4732
R524 VTAIL.n116 VTAIL.n98 10.4732
R525 VTAIL.n138 VTAIL.n88 10.4732
R526 VTAIL.n196 VTAIL.n178 10.4732
R527 VTAIL.n218 VTAIL.n168 10.4732
R528 VTAIL.n534 VTAIL.n484 10.4732
R529 VTAIL.n513 VTAIL.n495 10.4732
R530 VTAIL.n454 VTAIL.n404 10.4732
R531 VTAIL.n433 VTAIL.n415 10.4732
R532 VTAIL.n376 VTAIL.n326 10.4732
R533 VTAIL.n355 VTAIL.n337 10.4732
R534 VTAIL.n296 VTAIL.n246 10.4732
R535 VTAIL.n275 VTAIL.n257 10.4732
R536 VTAIL.n589 VTAIL.n574 9.69747
R537 VTAIL.n616 VTAIL.n615 9.69747
R538 VTAIL.n37 VTAIL.n22 9.69747
R539 VTAIL.n64 VTAIL.n63 9.69747
R540 VTAIL.n115 VTAIL.n100 9.69747
R541 VTAIL.n142 VTAIL.n141 9.69747
R542 VTAIL.n195 VTAIL.n180 9.69747
R543 VTAIL.n222 VTAIL.n221 9.69747
R544 VTAIL.n538 VTAIL.n537 9.69747
R545 VTAIL.n512 VTAIL.n497 9.69747
R546 VTAIL.n458 VTAIL.n457 9.69747
R547 VTAIL.n432 VTAIL.n417 9.69747
R548 VTAIL.n380 VTAIL.n379 9.69747
R549 VTAIL.n354 VTAIL.n339 9.69747
R550 VTAIL.n300 VTAIL.n299 9.69747
R551 VTAIL.n274 VTAIL.n259 9.69747
R552 VTAIL.n630 VTAIL.n629 9.45567
R553 VTAIL.n78 VTAIL.n77 9.45567
R554 VTAIL.n156 VTAIL.n155 9.45567
R555 VTAIL.n236 VTAIL.n235 9.45567
R556 VTAIL.n552 VTAIL.n551 9.45567
R557 VTAIL.n472 VTAIL.n471 9.45567
R558 VTAIL.n394 VTAIL.n393 9.45567
R559 VTAIL.n314 VTAIL.n313 9.45567
R560 VTAIL.n556 VTAIL.n555 9.3005
R561 VTAIL.n629 VTAIL.n628 9.3005
R562 VTAIL.n621 VTAIL.n620 9.3005
R563 VTAIL.n560 VTAIL.n559 9.3005
R564 VTAIL.n615 VTAIL.n614 9.3005
R565 VTAIL.n613 VTAIL.n612 9.3005
R566 VTAIL.n564 VTAIL.n563 9.3005
R567 VTAIL.n607 VTAIL.n606 9.3005
R568 VTAIL.n605 VTAIL.n604 9.3005
R569 VTAIL.n581 VTAIL.n580 9.3005
R570 VTAIL.n576 VTAIL.n575 9.3005
R571 VTAIL.n587 VTAIL.n586 9.3005
R572 VTAIL.n589 VTAIL.n588 9.3005
R573 VTAIL.n572 VTAIL.n571 9.3005
R574 VTAIL.n595 VTAIL.n594 9.3005
R575 VTAIL.n597 VTAIL.n596 9.3005
R576 VTAIL.n598 VTAIL.n567 9.3005
R577 VTAIL.n623 VTAIL.n622 9.3005
R578 VTAIL.n4 VTAIL.n3 9.3005
R579 VTAIL.n77 VTAIL.n76 9.3005
R580 VTAIL.n69 VTAIL.n68 9.3005
R581 VTAIL.n8 VTAIL.n7 9.3005
R582 VTAIL.n63 VTAIL.n62 9.3005
R583 VTAIL.n61 VTAIL.n60 9.3005
R584 VTAIL.n12 VTAIL.n11 9.3005
R585 VTAIL.n55 VTAIL.n54 9.3005
R586 VTAIL.n53 VTAIL.n52 9.3005
R587 VTAIL.n29 VTAIL.n28 9.3005
R588 VTAIL.n24 VTAIL.n23 9.3005
R589 VTAIL.n35 VTAIL.n34 9.3005
R590 VTAIL.n37 VTAIL.n36 9.3005
R591 VTAIL.n20 VTAIL.n19 9.3005
R592 VTAIL.n43 VTAIL.n42 9.3005
R593 VTAIL.n45 VTAIL.n44 9.3005
R594 VTAIL.n46 VTAIL.n15 9.3005
R595 VTAIL.n71 VTAIL.n70 9.3005
R596 VTAIL.n82 VTAIL.n81 9.3005
R597 VTAIL.n155 VTAIL.n154 9.3005
R598 VTAIL.n147 VTAIL.n146 9.3005
R599 VTAIL.n86 VTAIL.n85 9.3005
R600 VTAIL.n141 VTAIL.n140 9.3005
R601 VTAIL.n139 VTAIL.n138 9.3005
R602 VTAIL.n90 VTAIL.n89 9.3005
R603 VTAIL.n133 VTAIL.n132 9.3005
R604 VTAIL.n131 VTAIL.n130 9.3005
R605 VTAIL.n107 VTAIL.n106 9.3005
R606 VTAIL.n102 VTAIL.n101 9.3005
R607 VTAIL.n113 VTAIL.n112 9.3005
R608 VTAIL.n115 VTAIL.n114 9.3005
R609 VTAIL.n98 VTAIL.n97 9.3005
R610 VTAIL.n121 VTAIL.n120 9.3005
R611 VTAIL.n123 VTAIL.n122 9.3005
R612 VTAIL.n124 VTAIL.n93 9.3005
R613 VTAIL.n149 VTAIL.n148 9.3005
R614 VTAIL.n162 VTAIL.n161 9.3005
R615 VTAIL.n235 VTAIL.n234 9.3005
R616 VTAIL.n227 VTAIL.n226 9.3005
R617 VTAIL.n166 VTAIL.n165 9.3005
R618 VTAIL.n221 VTAIL.n220 9.3005
R619 VTAIL.n219 VTAIL.n218 9.3005
R620 VTAIL.n170 VTAIL.n169 9.3005
R621 VTAIL.n213 VTAIL.n212 9.3005
R622 VTAIL.n211 VTAIL.n210 9.3005
R623 VTAIL.n187 VTAIL.n186 9.3005
R624 VTAIL.n182 VTAIL.n181 9.3005
R625 VTAIL.n193 VTAIL.n192 9.3005
R626 VTAIL.n195 VTAIL.n194 9.3005
R627 VTAIL.n178 VTAIL.n177 9.3005
R628 VTAIL.n201 VTAIL.n200 9.3005
R629 VTAIL.n203 VTAIL.n202 9.3005
R630 VTAIL.n204 VTAIL.n173 9.3005
R631 VTAIL.n229 VTAIL.n228 9.3005
R632 VTAIL.n478 VTAIL.n477 9.3005
R633 VTAIL.n545 VTAIL.n544 9.3005
R634 VTAIL.n543 VTAIL.n542 9.3005
R635 VTAIL.n482 VTAIL.n481 9.3005
R636 VTAIL.n537 VTAIL.n536 9.3005
R637 VTAIL.n535 VTAIL.n534 9.3005
R638 VTAIL.n486 VTAIL.n485 9.3005
R639 VTAIL.n529 VTAIL.n528 9.3005
R640 VTAIL.n527 VTAIL.n526 9.3005
R641 VTAIL.n492 VTAIL.n489 9.3005
R642 VTAIL.n520 VTAIL.n519 9.3005
R643 VTAIL.n518 VTAIL.n517 9.3005
R644 VTAIL.n495 VTAIL.n494 9.3005
R645 VTAIL.n512 VTAIL.n511 9.3005
R646 VTAIL.n510 VTAIL.n509 9.3005
R647 VTAIL.n499 VTAIL.n498 9.3005
R648 VTAIL.n504 VTAIL.n503 9.3005
R649 VTAIL.n551 VTAIL.n550 9.3005
R650 VTAIL.n424 VTAIL.n423 9.3005
R651 VTAIL.n419 VTAIL.n418 9.3005
R652 VTAIL.n430 VTAIL.n429 9.3005
R653 VTAIL.n432 VTAIL.n431 9.3005
R654 VTAIL.n415 VTAIL.n414 9.3005
R655 VTAIL.n438 VTAIL.n437 9.3005
R656 VTAIL.n440 VTAIL.n439 9.3005
R657 VTAIL.n412 VTAIL.n409 9.3005
R658 VTAIL.n471 VTAIL.n470 9.3005
R659 VTAIL.n398 VTAIL.n397 9.3005
R660 VTAIL.n465 VTAIL.n464 9.3005
R661 VTAIL.n463 VTAIL.n462 9.3005
R662 VTAIL.n402 VTAIL.n401 9.3005
R663 VTAIL.n457 VTAIL.n456 9.3005
R664 VTAIL.n455 VTAIL.n454 9.3005
R665 VTAIL.n406 VTAIL.n405 9.3005
R666 VTAIL.n449 VTAIL.n448 9.3005
R667 VTAIL.n447 VTAIL.n446 9.3005
R668 VTAIL.n346 VTAIL.n345 9.3005
R669 VTAIL.n341 VTAIL.n340 9.3005
R670 VTAIL.n352 VTAIL.n351 9.3005
R671 VTAIL.n354 VTAIL.n353 9.3005
R672 VTAIL.n337 VTAIL.n336 9.3005
R673 VTAIL.n360 VTAIL.n359 9.3005
R674 VTAIL.n362 VTAIL.n361 9.3005
R675 VTAIL.n334 VTAIL.n331 9.3005
R676 VTAIL.n393 VTAIL.n392 9.3005
R677 VTAIL.n320 VTAIL.n319 9.3005
R678 VTAIL.n387 VTAIL.n386 9.3005
R679 VTAIL.n385 VTAIL.n384 9.3005
R680 VTAIL.n324 VTAIL.n323 9.3005
R681 VTAIL.n379 VTAIL.n378 9.3005
R682 VTAIL.n377 VTAIL.n376 9.3005
R683 VTAIL.n328 VTAIL.n327 9.3005
R684 VTAIL.n371 VTAIL.n370 9.3005
R685 VTAIL.n369 VTAIL.n368 9.3005
R686 VTAIL.n266 VTAIL.n265 9.3005
R687 VTAIL.n261 VTAIL.n260 9.3005
R688 VTAIL.n272 VTAIL.n271 9.3005
R689 VTAIL.n274 VTAIL.n273 9.3005
R690 VTAIL.n257 VTAIL.n256 9.3005
R691 VTAIL.n280 VTAIL.n279 9.3005
R692 VTAIL.n282 VTAIL.n281 9.3005
R693 VTAIL.n254 VTAIL.n251 9.3005
R694 VTAIL.n313 VTAIL.n312 9.3005
R695 VTAIL.n240 VTAIL.n239 9.3005
R696 VTAIL.n307 VTAIL.n306 9.3005
R697 VTAIL.n305 VTAIL.n304 9.3005
R698 VTAIL.n244 VTAIL.n243 9.3005
R699 VTAIL.n299 VTAIL.n298 9.3005
R700 VTAIL.n297 VTAIL.n296 9.3005
R701 VTAIL.n248 VTAIL.n247 9.3005
R702 VTAIL.n291 VTAIL.n290 9.3005
R703 VTAIL.n289 VTAIL.n288 9.3005
R704 VTAIL.n586 VTAIL.n585 8.92171
R705 VTAIL.n619 VTAIL.n560 8.92171
R706 VTAIL.n34 VTAIL.n33 8.92171
R707 VTAIL.n67 VTAIL.n8 8.92171
R708 VTAIL.n112 VTAIL.n111 8.92171
R709 VTAIL.n145 VTAIL.n86 8.92171
R710 VTAIL.n192 VTAIL.n191 8.92171
R711 VTAIL.n225 VTAIL.n166 8.92171
R712 VTAIL.n541 VTAIL.n482 8.92171
R713 VTAIL.n509 VTAIL.n508 8.92171
R714 VTAIL.n461 VTAIL.n402 8.92171
R715 VTAIL.n429 VTAIL.n428 8.92171
R716 VTAIL.n383 VTAIL.n324 8.92171
R717 VTAIL.n351 VTAIL.n350 8.92171
R718 VTAIL.n303 VTAIL.n244 8.92171
R719 VTAIL.n271 VTAIL.n270 8.92171
R720 VTAIL.n582 VTAIL.n576 8.14595
R721 VTAIL.n620 VTAIL.n558 8.14595
R722 VTAIL.n630 VTAIL.n554 8.14595
R723 VTAIL.n30 VTAIL.n24 8.14595
R724 VTAIL.n68 VTAIL.n6 8.14595
R725 VTAIL.n78 VTAIL.n2 8.14595
R726 VTAIL.n108 VTAIL.n102 8.14595
R727 VTAIL.n146 VTAIL.n84 8.14595
R728 VTAIL.n156 VTAIL.n80 8.14595
R729 VTAIL.n188 VTAIL.n182 8.14595
R730 VTAIL.n226 VTAIL.n164 8.14595
R731 VTAIL.n236 VTAIL.n160 8.14595
R732 VTAIL.n552 VTAIL.n476 8.14595
R733 VTAIL.n542 VTAIL.n480 8.14595
R734 VTAIL.n505 VTAIL.n499 8.14595
R735 VTAIL.n472 VTAIL.n396 8.14595
R736 VTAIL.n462 VTAIL.n400 8.14595
R737 VTAIL.n425 VTAIL.n419 8.14595
R738 VTAIL.n394 VTAIL.n318 8.14595
R739 VTAIL.n384 VTAIL.n322 8.14595
R740 VTAIL.n347 VTAIL.n341 8.14595
R741 VTAIL.n314 VTAIL.n238 8.14595
R742 VTAIL.n304 VTAIL.n242 8.14595
R743 VTAIL.n267 VTAIL.n261 8.14595
R744 VTAIL.n581 VTAIL.n578 7.3702
R745 VTAIL.n624 VTAIL.n623 7.3702
R746 VTAIL.n628 VTAIL.n627 7.3702
R747 VTAIL.n29 VTAIL.n26 7.3702
R748 VTAIL.n72 VTAIL.n71 7.3702
R749 VTAIL.n76 VTAIL.n75 7.3702
R750 VTAIL.n107 VTAIL.n104 7.3702
R751 VTAIL.n150 VTAIL.n149 7.3702
R752 VTAIL.n154 VTAIL.n153 7.3702
R753 VTAIL.n187 VTAIL.n184 7.3702
R754 VTAIL.n230 VTAIL.n229 7.3702
R755 VTAIL.n234 VTAIL.n233 7.3702
R756 VTAIL.n550 VTAIL.n549 7.3702
R757 VTAIL.n546 VTAIL.n545 7.3702
R758 VTAIL.n504 VTAIL.n501 7.3702
R759 VTAIL.n470 VTAIL.n469 7.3702
R760 VTAIL.n466 VTAIL.n465 7.3702
R761 VTAIL.n424 VTAIL.n421 7.3702
R762 VTAIL.n392 VTAIL.n391 7.3702
R763 VTAIL.n388 VTAIL.n387 7.3702
R764 VTAIL.n346 VTAIL.n343 7.3702
R765 VTAIL.n312 VTAIL.n311 7.3702
R766 VTAIL.n308 VTAIL.n307 7.3702
R767 VTAIL.n266 VTAIL.n263 7.3702
R768 VTAIL.n624 VTAIL.n556 6.59444
R769 VTAIL.n627 VTAIL.n556 6.59444
R770 VTAIL.n72 VTAIL.n4 6.59444
R771 VTAIL.n75 VTAIL.n4 6.59444
R772 VTAIL.n150 VTAIL.n82 6.59444
R773 VTAIL.n153 VTAIL.n82 6.59444
R774 VTAIL.n230 VTAIL.n162 6.59444
R775 VTAIL.n233 VTAIL.n162 6.59444
R776 VTAIL.n549 VTAIL.n478 6.59444
R777 VTAIL.n546 VTAIL.n478 6.59444
R778 VTAIL.n469 VTAIL.n398 6.59444
R779 VTAIL.n466 VTAIL.n398 6.59444
R780 VTAIL.n391 VTAIL.n320 6.59444
R781 VTAIL.n388 VTAIL.n320 6.59444
R782 VTAIL.n311 VTAIL.n240 6.59444
R783 VTAIL.n308 VTAIL.n240 6.59444
R784 VTAIL.n582 VTAIL.n581 5.81868
R785 VTAIL.n623 VTAIL.n558 5.81868
R786 VTAIL.n628 VTAIL.n554 5.81868
R787 VTAIL.n30 VTAIL.n29 5.81868
R788 VTAIL.n71 VTAIL.n6 5.81868
R789 VTAIL.n76 VTAIL.n2 5.81868
R790 VTAIL.n108 VTAIL.n107 5.81868
R791 VTAIL.n149 VTAIL.n84 5.81868
R792 VTAIL.n154 VTAIL.n80 5.81868
R793 VTAIL.n188 VTAIL.n187 5.81868
R794 VTAIL.n229 VTAIL.n164 5.81868
R795 VTAIL.n234 VTAIL.n160 5.81868
R796 VTAIL.n550 VTAIL.n476 5.81868
R797 VTAIL.n545 VTAIL.n480 5.81868
R798 VTAIL.n505 VTAIL.n504 5.81868
R799 VTAIL.n470 VTAIL.n396 5.81868
R800 VTAIL.n465 VTAIL.n400 5.81868
R801 VTAIL.n425 VTAIL.n424 5.81868
R802 VTAIL.n392 VTAIL.n318 5.81868
R803 VTAIL.n387 VTAIL.n322 5.81868
R804 VTAIL.n347 VTAIL.n346 5.81868
R805 VTAIL.n312 VTAIL.n238 5.81868
R806 VTAIL.n307 VTAIL.n242 5.81868
R807 VTAIL.n267 VTAIL.n266 5.81868
R808 VTAIL.n585 VTAIL.n576 5.04292
R809 VTAIL.n620 VTAIL.n619 5.04292
R810 VTAIL.n33 VTAIL.n24 5.04292
R811 VTAIL.n68 VTAIL.n67 5.04292
R812 VTAIL.n111 VTAIL.n102 5.04292
R813 VTAIL.n146 VTAIL.n145 5.04292
R814 VTAIL.n191 VTAIL.n182 5.04292
R815 VTAIL.n226 VTAIL.n225 5.04292
R816 VTAIL.n542 VTAIL.n541 5.04292
R817 VTAIL.n508 VTAIL.n499 5.04292
R818 VTAIL.n462 VTAIL.n461 5.04292
R819 VTAIL.n428 VTAIL.n419 5.04292
R820 VTAIL.n384 VTAIL.n383 5.04292
R821 VTAIL.n350 VTAIL.n341 5.04292
R822 VTAIL.n304 VTAIL.n303 5.04292
R823 VTAIL.n270 VTAIL.n261 5.04292
R824 VTAIL.n586 VTAIL.n574 4.26717
R825 VTAIL.n616 VTAIL.n560 4.26717
R826 VTAIL.n34 VTAIL.n22 4.26717
R827 VTAIL.n64 VTAIL.n8 4.26717
R828 VTAIL.n112 VTAIL.n100 4.26717
R829 VTAIL.n142 VTAIL.n86 4.26717
R830 VTAIL.n192 VTAIL.n180 4.26717
R831 VTAIL.n222 VTAIL.n166 4.26717
R832 VTAIL.n538 VTAIL.n482 4.26717
R833 VTAIL.n509 VTAIL.n497 4.26717
R834 VTAIL.n458 VTAIL.n402 4.26717
R835 VTAIL.n429 VTAIL.n417 4.26717
R836 VTAIL.n380 VTAIL.n324 4.26717
R837 VTAIL.n351 VTAIL.n339 4.26717
R838 VTAIL.n300 VTAIL.n244 4.26717
R839 VTAIL.n271 VTAIL.n259 4.26717
R840 VTAIL.n590 VTAIL.n589 3.49141
R841 VTAIL.n615 VTAIL.n562 3.49141
R842 VTAIL.n38 VTAIL.n37 3.49141
R843 VTAIL.n63 VTAIL.n10 3.49141
R844 VTAIL.n116 VTAIL.n115 3.49141
R845 VTAIL.n141 VTAIL.n88 3.49141
R846 VTAIL.n196 VTAIL.n195 3.49141
R847 VTAIL.n221 VTAIL.n168 3.49141
R848 VTAIL.n537 VTAIL.n484 3.49141
R849 VTAIL.n513 VTAIL.n512 3.49141
R850 VTAIL.n457 VTAIL.n404 3.49141
R851 VTAIL.n433 VTAIL.n432 3.49141
R852 VTAIL.n379 VTAIL.n326 3.49141
R853 VTAIL.n355 VTAIL.n354 3.49141
R854 VTAIL.n299 VTAIL.n246 3.49141
R855 VTAIL.n275 VTAIL.n274 3.49141
R856 VTAIL.n317 VTAIL.n315 3.44878
R857 VTAIL.n395 VTAIL.n317 3.44878
R858 VTAIL.n475 VTAIL.n473 3.44878
R859 VTAIL.n553 VTAIL.n475 3.44878
R860 VTAIL.n237 VTAIL.n159 3.44878
R861 VTAIL.n159 VTAIL.n157 3.44878
R862 VTAIL.n79 VTAIL.n1 3.44878
R863 VTAIL VTAIL.n631 3.39059
R864 VTAIL.n593 VTAIL.n572 2.71565
R865 VTAIL.n612 VTAIL.n611 2.71565
R866 VTAIL.n41 VTAIL.n20 2.71565
R867 VTAIL.n60 VTAIL.n59 2.71565
R868 VTAIL.n119 VTAIL.n98 2.71565
R869 VTAIL.n138 VTAIL.n137 2.71565
R870 VTAIL.n199 VTAIL.n178 2.71565
R871 VTAIL.n218 VTAIL.n217 2.71565
R872 VTAIL.n534 VTAIL.n533 2.71565
R873 VTAIL.n516 VTAIL.n495 2.71565
R874 VTAIL.n454 VTAIL.n453 2.71565
R875 VTAIL.n436 VTAIL.n415 2.71565
R876 VTAIL.n376 VTAIL.n375 2.71565
R877 VTAIL.n358 VTAIL.n337 2.71565
R878 VTAIL.n296 VTAIL.n295 2.71565
R879 VTAIL.n278 VTAIL.n257 2.71565
R880 VTAIL.n503 VTAIL.n502 2.41282
R881 VTAIL.n423 VTAIL.n422 2.41282
R882 VTAIL.n345 VTAIL.n344 2.41282
R883 VTAIL.n265 VTAIL.n264 2.41282
R884 VTAIL.n580 VTAIL.n579 2.41282
R885 VTAIL.n28 VTAIL.n27 2.41282
R886 VTAIL.n106 VTAIL.n105 2.41282
R887 VTAIL.n186 VTAIL.n185 2.41282
R888 VTAIL.n0 VTAIL.t8 2.29443
R889 VTAIL.n0 VTAIL.t13 2.29443
R890 VTAIL.n158 VTAIL.t0 2.29443
R891 VTAIL.n158 VTAIL.t5 2.29443
R892 VTAIL.n474 VTAIL.t6 2.29443
R893 VTAIL.n474 VTAIL.t3 2.29443
R894 VTAIL.n316 VTAIL.t9 2.29443
R895 VTAIL.n316 VTAIL.t15 2.29443
R896 VTAIL.n594 VTAIL.n570 1.93989
R897 VTAIL.n608 VTAIL.n564 1.93989
R898 VTAIL.n42 VTAIL.n18 1.93989
R899 VTAIL.n56 VTAIL.n12 1.93989
R900 VTAIL.n120 VTAIL.n96 1.93989
R901 VTAIL.n134 VTAIL.n90 1.93989
R902 VTAIL.n200 VTAIL.n176 1.93989
R903 VTAIL.n214 VTAIL.n170 1.93989
R904 VTAIL.n530 VTAIL.n486 1.93989
R905 VTAIL.n517 VTAIL.n493 1.93989
R906 VTAIL.n450 VTAIL.n406 1.93989
R907 VTAIL.n437 VTAIL.n413 1.93989
R908 VTAIL.n372 VTAIL.n328 1.93989
R909 VTAIL.n359 VTAIL.n335 1.93989
R910 VTAIL.n292 VTAIL.n248 1.93989
R911 VTAIL.n279 VTAIL.n255 1.93989
R912 VTAIL.n599 VTAIL.n597 1.16414
R913 VTAIL.n607 VTAIL.n566 1.16414
R914 VTAIL.n47 VTAIL.n45 1.16414
R915 VTAIL.n55 VTAIL.n14 1.16414
R916 VTAIL.n125 VTAIL.n123 1.16414
R917 VTAIL.n133 VTAIL.n92 1.16414
R918 VTAIL.n205 VTAIL.n203 1.16414
R919 VTAIL.n213 VTAIL.n172 1.16414
R920 VTAIL.n529 VTAIL.n488 1.16414
R921 VTAIL.n521 VTAIL.n520 1.16414
R922 VTAIL.n449 VTAIL.n408 1.16414
R923 VTAIL.n441 VTAIL.n440 1.16414
R924 VTAIL.n371 VTAIL.n330 1.16414
R925 VTAIL.n363 VTAIL.n362 1.16414
R926 VTAIL.n291 VTAIL.n250 1.16414
R927 VTAIL.n283 VTAIL.n282 1.16414
R928 VTAIL.n473 VTAIL.n395 0.470328
R929 VTAIL.n157 VTAIL.n79 0.470328
R930 VTAIL.n598 VTAIL.n568 0.388379
R931 VTAIL.n604 VTAIL.n603 0.388379
R932 VTAIL.n46 VTAIL.n16 0.388379
R933 VTAIL.n52 VTAIL.n51 0.388379
R934 VTAIL.n124 VTAIL.n94 0.388379
R935 VTAIL.n130 VTAIL.n129 0.388379
R936 VTAIL.n204 VTAIL.n174 0.388379
R937 VTAIL.n210 VTAIL.n209 0.388379
R938 VTAIL.n526 VTAIL.n525 0.388379
R939 VTAIL.n492 VTAIL.n490 0.388379
R940 VTAIL.n446 VTAIL.n445 0.388379
R941 VTAIL.n412 VTAIL.n410 0.388379
R942 VTAIL.n368 VTAIL.n367 0.388379
R943 VTAIL.n334 VTAIL.n332 0.388379
R944 VTAIL.n288 VTAIL.n287 0.388379
R945 VTAIL.n254 VTAIL.n252 0.388379
R946 VTAIL.n580 VTAIL.n575 0.155672
R947 VTAIL.n587 VTAIL.n575 0.155672
R948 VTAIL.n588 VTAIL.n587 0.155672
R949 VTAIL.n588 VTAIL.n571 0.155672
R950 VTAIL.n595 VTAIL.n571 0.155672
R951 VTAIL.n596 VTAIL.n595 0.155672
R952 VTAIL.n596 VTAIL.n567 0.155672
R953 VTAIL.n605 VTAIL.n567 0.155672
R954 VTAIL.n606 VTAIL.n605 0.155672
R955 VTAIL.n606 VTAIL.n563 0.155672
R956 VTAIL.n613 VTAIL.n563 0.155672
R957 VTAIL.n614 VTAIL.n613 0.155672
R958 VTAIL.n614 VTAIL.n559 0.155672
R959 VTAIL.n621 VTAIL.n559 0.155672
R960 VTAIL.n622 VTAIL.n621 0.155672
R961 VTAIL.n622 VTAIL.n555 0.155672
R962 VTAIL.n629 VTAIL.n555 0.155672
R963 VTAIL.n28 VTAIL.n23 0.155672
R964 VTAIL.n35 VTAIL.n23 0.155672
R965 VTAIL.n36 VTAIL.n35 0.155672
R966 VTAIL.n36 VTAIL.n19 0.155672
R967 VTAIL.n43 VTAIL.n19 0.155672
R968 VTAIL.n44 VTAIL.n43 0.155672
R969 VTAIL.n44 VTAIL.n15 0.155672
R970 VTAIL.n53 VTAIL.n15 0.155672
R971 VTAIL.n54 VTAIL.n53 0.155672
R972 VTAIL.n54 VTAIL.n11 0.155672
R973 VTAIL.n61 VTAIL.n11 0.155672
R974 VTAIL.n62 VTAIL.n61 0.155672
R975 VTAIL.n62 VTAIL.n7 0.155672
R976 VTAIL.n69 VTAIL.n7 0.155672
R977 VTAIL.n70 VTAIL.n69 0.155672
R978 VTAIL.n70 VTAIL.n3 0.155672
R979 VTAIL.n77 VTAIL.n3 0.155672
R980 VTAIL.n106 VTAIL.n101 0.155672
R981 VTAIL.n113 VTAIL.n101 0.155672
R982 VTAIL.n114 VTAIL.n113 0.155672
R983 VTAIL.n114 VTAIL.n97 0.155672
R984 VTAIL.n121 VTAIL.n97 0.155672
R985 VTAIL.n122 VTAIL.n121 0.155672
R986 VTAIL.n122 VTAIL.n93 0.155672
R987 VTAIL.n131 VTAIL.n93 0.155672
R988 VTAIL.n132 VTAIL.n131 0.155672
R989 VTAIL.n132 VTAIL.n89 0.155672
R990 VTAIL.n139 VTAIL.n89 0.155672
R991 VTAIL.n140 VTAIL.n139 0.155672
R992 VTAIL.n140 VTAIL.n85 0.155672
R993 VTAIL.n147 VTAIL.n85 0.155672
R994 VTAIL.n148 VTAIL.n147 0.155672
R995 VTAIL.n148 VTAIL.n81 0.155672
R996 VTAIL.n155 VTAIL.n81 0.155672
R997 VTAIL.n186 VTAIL.n181 0.155672
R998 VTAIL.n193 VTAIL.n181 0.155672
R999 VTAIL.n194 VTAIL.n193 0.155672
R1000 VTAIL.n194 VTAIL.n177 0.155672
R1001 VTAIL.n201 VTAIL.n177 0.155672
R1002 VTAIL.n202 VTAIL.n201 0.155672
R1003 VTAIL.n202 VTAIL.n173 0.155672
R1004 VTAIL.n211 VTAIL.n173 0.155672
R1005 VTAIL.n212 VTAIL.n211 0.155672
R1006 VTAIL.n212 VTAIL.n169 0.155672
R1007 VTAIL.n219 VTAIL.n169 0.155672
R1008 VTAIL.n220 VTAIL.n219 0.155672
R1009 VTAIL.n220 VTAIL.n165 0.155672
R1010 VTAIL.n227 VTAIL.n165 0.155672
R1011 VTAIL.n228 VTAIL.n227 0.155672
R1012 VTAIL.n228 VTAIL.n161 0.155672
R1013 VTAIL.n235 VTAIL.n161 0.155672
R1014 VTAIL.n551 VTAIL.n477 0.155672
R1015 VTAIL.n544 VTAIL.n477 0.155672
R1016 VTAIL.n544 VTAIL.n543 0.155672
R1017 VTAIL.n543 VTAIL.n481 0.155672
R1018 VTAIL.n536 VTAIL.n481 0.155672
R1019 VTAIL.n536 VTAIL.n535 0.155672
R1020 VTAIL.n535 VTAIL.n485 0.155672
R1021 VTAIL.n528 VTAIL.n485 0.155672
R1022 VTAIL.n528 VTAIL.n527 0.155672
R1023 VTAIL.n527 VTAIL.n489 0.155672
R1024 VTAIL.n519 VTAIL.n489 0.155672
R1025 VTAIL.n519 VTAIL.n518 0.155672
R1026 VTAIL.n518 VTAIL.n494 0.155672
R1027 VTAIL.n511 VTAIL.n494 0.155672
R1028 VTAIL.n511 VTAIL.n510 0.155672
R1029 VTAIL.n510 VTAIL.n498 0.155672
R1030 VTAIL.n503 VTAIL.n498 0.155672
R1031 VTAIL.n471 VTAIL.n397 0.155672
R1032 VTAIL.n464 VTAIL.n397 0.155672
R1033 VTAIL.n464 VTAIL.n463 0.155672
R1034 VTAIL.n463 VTAIL.n401 0.155672
R1035 VTAIL.n456 VTAIL.n401 0.155672
R1036 VTAIL.n456 VTAIL.n455 0.155672
R1037 VTAIL.n455 VTAIL.n405 0.155672
R1038 VTAIL.n448 VTAIL.n405 0.155672
R1039 VTAIL.n448 VTAIL.n447 0.155672
R1040 VTAIL.n447 VTAIL.n409 0.155672
R1041 VTAIL.n439 VTAIL.n409 0.155672
R1042 VTAIL.n439 VTAIL.n438 0.155672
R1043 VTAIL.n438 VTAIL.n414 0.155672
R1044 VTAIL.n431 VTAIL.n414 0.155672
R1045 VTAIL.n431 VTAIL.n430 0.155672
R1046 VTAIL.n430 VTAIL.n418 0.155672
R1047 VTAIL.n423 VTAIL.n418 0.155672
R1048 VTAIL.n393 VTAIL.n319 0.155672
R1049 VTAIL.n386 VTAIL.n319 0.155672
R1050 VTAIL.n386 VTAIL.n385 0.155672
R1051 VTAIL.n385 VTAIL.n323 0.155672
R1052 VTAIL.n378 VTAIL.n323 0.155672
R1053 VTAIL.n378 VTAIL.n377 0.155672
R1054 VTAIL.n377 VTAIL.n327 0.155672
R1055 VTAIL.n370 VTAIL.n327 0.155672
R1056 VTAIL.n370 VTAIL.n369 0.155672
R1057 VTAIL.n369 VTAIL.n331 0.155672
R1058 VTAIL.n361 VTAIL.n331 0.155672
R1059 VTAIL.n361 VTAIL.n360 0.155672
R1060 VTAIL.n360 VTAIL.n336 0.155672
R1061 VTAIL.n353 VTAIL.n336 0.155672
R1062 VTAIL.n353 VTAIL.n352 0.155672
R1063 VTAIL.n352 VTAIL.n340 0.155672
R1064 VTAIL.n345 VTAIL.n340 0.155672
R1065 VTAIL.n313 VTAIL.n239 0.155672
R1066 VTAIL.n306 VTAIL.n239 0.155672
R1067 VTAIL.n306 VTAIL.n305 0.155672
R1068 VTAIL.n305 VTAIL.n243 0.155672
R1069 VTAIL.n298 VTAIL.n243 0.155672
R1070 VTAIL.n298 VTAIL.n297 0.155672
R1071 VTAIL.n297 VTAIL.n247 0.155672
R1072 VTAIL.n290 VTAIL.n247 0.155672
R1073 VTAIL.n290 VTAIL.n289 0.155672
R1074 VTAIL.n289 VTAIL.n251 0.155672
R1075 VTAIL.n281 VTAIL.n251 0.155672
R1076 VTAIL.n281 VTAIL.n280 0.155672
R1077 VTAIL.n280 VTAIL.n256 0.155672
R1078 VTAIL.n273 VTAIL.n256 0.155672
R1079 VTAIL.n273 VTAIL.n272 0.155672
R1080 VTAIL.n272 VTAIL.n260 0.155672
R1081 VTAIL.n265 VTAIL.n260 0.155672
R1082 VTAIL VTAIL.n1 0.0586897
R1083 VP.n22 VP.n19 161.3
R1084 VP.n24 VP.n23 161.3
R1085 VP.n25 VP.n18 161.3
R1086 VP.n27 VP.n26 161.3
R1087 VP.n28 VP.n17 161.3
R1088 VP.n30 VP.n29 161.3
R1089 VP.n31 VP.n16 161.3
R1090 VP.n33 VP.n32 161.3
R1091 VP.n34 VP.n15 161.3
R1092 VP.n36 VP.n35 161.3
R1093 VP.n37 VP.n14 161.3
R1094 VP.n39 VP.n38 161.3
R1095 VP.n40 VP.n13 161.3
R1096 VP.n42 VP.n41 161.3
R1097 VP.n43 VP.n12 161.3
R1098 VP.n81 VP.n0 161.3
R1099 VP.n80 VP.n79 161.3
R1100 VP.n78 VP.n1 161.3
R1101 VP.n77 VP.n76 161.3
R1102 VP.n75 VP.n2 161.3
R1103 VP.n74 VP.n73 161.3
R1104 VP.n72 VP.n3 161.3
R1105 VP.n71 VP.n70 161.3
R1106 VP.n69 VP.n4 161.3
R1107 VP.n68 VP.n67 161.3
R1108 VP.n66 VP.n5 161.3
R1109 VP.n65 VP.n64 161.3
R1110 VP.n63 VP.n6 161.3
R1111 VP.n62 VP.n61 161.3
R1112 VP.n60 VP.n7 161.3
R1113 VP.n59 VP.n58 161.3
R1114 VP.n57 VP.n8 161.3
R1115 VP.n56 VP.n55 161.3
R1116 VP.n54 VP.n9 161.3
R1117 VP.n53 VP.n52 161.3
R1118 VP.n51 VP.n10 161.3
R1119 VP.n50 VP.n49 161.3
R1120 VP.n48 VP.n11 161.3
R1121 VP.n21 VP.t1 125.16
R1122 VP.n82 VP.t7 93.0515
R1123 VP.n70 VP.t2 93.0515
R1124 VP.n58 VP.t3 93.0515
R1125 VP.n46 VP.t5 93.0515
R1126 VP.n20 VP.t6 93.0515
R1127 VP.n32 VP.t0 93.0515
R1128 VP.n44 VP.t4 93.0515
R1129 VP.n47 VP.n45 57.7767
R1130 VP.n47 VP.n46 57.7148
R1131 VP.n83 VP.n82 57.7148
R1132 VP.n45 VP.n44 57.7148
R1133 VP.n21 VP.n20 50.4779
R1134 VP.n52 VP.n51 40.4934
R1135 VP.n52 VP.n9 40.4934
R1136 VP.n64 VP.n63 40.4934
R1137 VP.n64 VP.n5 40.4934
R1138 VP.n76 VP.n75 40.4934
R1139 VP.n76 VP.n1 40.4934
R1140 VP.n38 VP.n13 40.4934
R1141 VP.n38 VP.n37 40.4934
R1142 VP.n26 VP.n17 40.4934
R1143 VP.n26 VP.n25 40.4934
R1144 VP.n46 VP.n11 24.4675
R1145 VP.n50 VP.n11 24.4675
R1146 VP.n51 VP.n50 24.4675
R1147 VP.n56 VP.n9 24.4675
R1148 VP.n57 VP.n56 24.4675
R1149 VP.n58 VP.n57 24.4675
R1150 VP.n58 VP.n7 24.4675
R1151 VP.n62 VP.n7 24.4675
R1152 VP.n63 VP.n62 24.4675
R1153 VP.n68 VP.n5 24.4675
R1154 VP.n69 VP.n68 24.4675
R1155 VP.n70 VP.n69 24.4675
R1156 VP.n70 VP.n3 24.4675
R1157 VP.n74 VP.n3 24.4675
R1158 VP.n75 VP.n74 24.4675
R1159 VP.n80 VP.n1 24.4675
R1160 VP.n81 VP.n80 24.4675
R1161 VP.n82 VP.n81 24.4675
R1162 VP.n42 VP.n13 24.4675
R1163 VP.n43 VP.n42 24.4675
R1164 VP.n44 VP.n43 24.4675
R1165 VP.n30 VP.n17 24.4675
R1166 VP.n31 VP.n30 24.4675
R1167 VP.n32 VP.n31 24.4675
R1168 VP.n32 VP.n15 24.4675
R1169 VP.n36 VP.n15 24.4675
R1170 VP.n37 VP.n36 24.4675
R1171 VP.n20 VP.n19 24.4675
R1172 VP.n24 VP.n19 24.4675
R1173 VP.n25 VP.n24 24.4675
R1174 VP.n22 VP.n21 2.52647
R1175 VP.n45 VP.n12 0.417535
R1176 VP.n48 VP.n47 0.417535
R1177 VP.n83 VP.n0 0.417535
R1178 VP VP.n83 0.394291
R1179 VP.n23 VP.n22 0.189894
R1180 VP.n23 VP.n18 0.189894
R1181 VP.n27 VP.n18 0.189894
R1182 VP.n28 VP.n27 0.189894
R1183 VP.n29 VP.n28 0.189894
R1184 VP.n29 VP.n16 0.189894
R1185 VP.n33 VP.n16 0.189894
R1186 VP.n34 VP.n33 0.189894
R1187 VP.n35 VP.n34 0.189894
R1188 VP.n35 VP.n14 0.189894
R1189 VP.n39 VP.n14 0.189894
R1190 VP.n40 VP.n39 0.189894
R1191 VP.n41 VP.n40 0.189894
R1192 VP.n41 VP.n12 0.189894
R1193 VP.n49 VP.n48 0.189894
R1194 VP.n49 VP.n10 0.189894
R1195 VP.n53 VP.n10 0.189894
R1196 VP.n54 VP.n53 0.189894
R1197 VP.n55 VP.n54 0.189894
R1198 VP.n55 VP.n8 0.189894
R1199 VP.n59 VP.n8 0.189894
R1200 VP.n60 VP.n59 0.189894
R1201 VP.n61 VP.n60 0.189894
R1202 VP.n61 VP.n6 0.189894
R1203 VP.n65 VP.n6 0.189894
R1204 VP.n66 VP.n65 0.189894
R1205 VP.n67 VP.n66 0.189894
R1206 VP.n67 VP.n4 0.189894
R1207 VP.n71 VP.n4 0.189894
R1208 VP.n72 VP.n71 0.189894
R1209 VP.n73 VP.n72 0.189894
R1210 VP.n73 VP.n2 0.189894
R1211 VP.n77 VP.n2 0.189894
R1212 VP.n78 VP.n77 0.189894
R1213 VP.n79 VP.n78 0.189894
R1214 VP.n79 VP.n0 0.189894
R1215 VDD1 VDD1.n0 71.282
R1216 VDD1.n3 VDD1.n2 71.1684
R1217 VDD1.n3 VDD1.n1 71.1684
R1218 VDD1.n5 VDD1.n4 69.4996
R1219 VDD1.n5 VDD1.n3 52.0311
R1220 VDD1.n4 VDD1.t7 2.29443
R1221 VDD1.n4 VDD1.t3 2.29443
R1222 VDD1.n0 VDD1.t6 2.29443
R1223 VDD1.n0 VDD1.t1 2.29443
R1224 VDD1.n2 VDD1.t5 2.29443
R1225 VDD1.n2 VDD1.t0 2.29443
R1226 VDD1.n1 VDD1.t2 2.29443
R1227 VDD1.n1 VDD1.t4 2.29443
R1228 VDD1 VDD1.n5 1.66645
R1229 B.n714 B.n93 585
R1230 B.n716 B.n715 585
R1231 B.n717 B.n92 585
R1232 B.n719 B.n718 585
R1233 B.n720 B.n91 585
R1234 B.n722 B.n721 585
R1235 B.n723 B.n90 585
R1236 B.n725 B.n724 585
R1237 B.n726 B.n89 585
R1238 B.n728 B.n727 585
R1239 B.n729 B.n88 585
R1240 B.n731 B.n730 585
R1241 B.n732 B.n87 585
R1242 B.n734 B.n733 585
R1243 B.n735 B.n86 585
R1244 B.n737 B.n736 585
R1245 B.n738 B.n85 585
R1246 B.n740 B.n739 585
R1247 B.n741 B.n84 585
R1248 B.n743 B.n742 585
R1249 B.n744 B.n83 585
R1250 B.n746 B.n745 585
R1251 B.n747 B.n82 585
R1252 B.n749 B.n748 585
R1253 B.n750 B.n81 585
R1254 B.n752 B.n751 585
R1255 B.n753 B.n80 585
R1256 B.n755 B.n754 585
R1257 B.n756 B.n79 585
R1258 B.n758 B.n757 585
R1259 B.n759 B.n78 585
R1260 B.n761 B.n760 585
R1261 B.n762 B.n77 585
R1262 B.n764 B.n763 585
R1263 B.n765 B.n76 585
R1264 B.n767 B.n766 585
R1265 B.n768 B.n75 585
R1266 B.n770 B.n769 585
R1267 B.n771 B.n74 585
R1268 B.n773 B.n772 585
R1269 B.n774 B.n73 585
R1270 B.n776 B.n775 585
R1271 B.n777 B.n72 585
R1272 B.n779 B.n778 585
R1273 B.n780 B.n71 585
R1274 B.n782 B.n781 585
R1275 B.n783 B.n67 585
R1276 B.n785 B.n784 585
R1277 B.n786 B.n66 585
R1278 B.n788 B.n787 585
R1279 B.n789 B.n65 585
R1280 B.n791 B.n790 585
R1281 B.n792 B.n64 585
R1282 B.n794 B.n793 585
R1283 B.n795 B.n63 585
R1284 B.n797 B.n796 585
R1285 B.n798 B.n62 585
R1286 B.n800 B.n799 585
R1287 B.n802 B.n59 585
R1288 B.n804 B.n803 585
R1289 B.n805 B.n58 585
R1290 B.n807 B.n806 585
R1291 B.n808 B.n57 585
R1292 B.n810 B.n809 585
R1293 B.n811 B.n56 585
R1294 B.n813 B.n812 585
R1295 B.n814 B.n55 585
R1296 B.n816 B.n815 585
R1297 B.n817 B.n54 585
R1298 B.n819 B.n818 585
R1299 B.n820 B.n53 585
R1300 B.n822 B.n821 585
R1301 B.n823 B.n52 585
R1302 B.n825 B.n824 585
R1303 B.n826 B.n51 585
R1304 B.n828 B.n827 585
R1305 B.n829 B.n50 585
R1306 B.n831 B.n830 585
R1307 B.n832 B.n49 585
R1308 B.n834 B.n833 585
R1309 B.n835 B.n48 585
R1310 B.n837 B.n836 585
R1311 B.n838 B.n47 585
R1312 B.n840 B.n839 585
R1313 B.n841 B.n46 585
R1314 B.n843 B.n842 585
R1315 B.n844 B.n45 585
R1316 B.n846 B.n845 585
R1317 B.n847 B.n44 585
R1318 B.n849 B.n848 585
R1319 B.n850 B.n43 585
R1320 B.n852 B.n851 585
R1321 B.n853 B.n42 585
R1322 B.n855 B.n854 585
R1323 B.n856 B.n41 585
R1324 B.n858 B.n857 585
R1325 B.n859 B.n40 585
R1326 B.n861 B.n860 585
R1327 B.n862 B.n39 585
R1328 B.n864 B.n863 585
R1329 B.n865 B.n38 585
R1330 B.n867 B.n866 585
R1331 B.n868 B.n37 585
R1332 B.n870 B.n869 585
R1333 B.n871 B.n36 585
R1334 B.n873 B.n872 585
R1335 B.n713 B.n712 585
R1336 B.n711 B.n94 585
R1337 B.n710 B.n709 585
R1338 B.n708 B.n95 585
R1339 B.n707 B.n706 585
R1340 B.n705 B.n96 585
R1341 B.n704 B.n703 585
R1342 B.n702 B.n97 585
R1343 B.n701 B.n700 585
R1344 B.n699 B.n98 585
R1345 B.n698 B.n697 585
R1346 B.n696 B.n99 585
R1347 B.n695 B.n694 585
R1348 B.n693 B.n100 585
R1349 B.n692 B.n691 585
R1350 B.n690 B.n101 585
R1351 B.n689 B.n688 585
R1352 B.n687 B.n102 585
R1353 B.n686 B.n685 585
R1354 B.n684 B.n103 585
R1355 B.n683 B.n682 585
R1356 B.n681 B.n104 585
R1357 B.n680 B.n679 585
R1358 B.n678 B.n105 585
R1359 B.n677 B.n676 585
R1360 B.n675 B.n106 585
R1361 B.n674 B.n673 585
R1362 B.n672 B.n107 585
R1363 B.n671 B.n670 585
R1364 B.n669 B.n108 585
R1365 B.n668 B.n667 585
R1366 B.n666 B.n109 585
R1367 B.n665 B.n664 585
R1368 B.n663 B.n110 585
R1369 B.n662 B.n661 585
R1370 B.n660 B.n111 585
R1371 B.n659 B.n658 585
R1372 B.n657 B.n112 585
R1373 B.n656 B.n655 585
R1374 B.n654 B.n113 585
R1375 B.n653 B.n652 585
R1376 B.n651 B.n114 585
R1377 B.n650 B.n649 585
R1378 B.n648 B.n115 585
R1379 B.n647 B.n646 585
R1380 B.n645 B.n116 585
R1381 B.n644 B.n643 585
R1382 B.n642 B.n117 585
R1383 B.n641 B.n640 585
R1384 B.n639 B.n118 585
R1385 B.n638 B.n637 585
R1386 B.n636 B.n119 585
R1387 B.n635 B.n634 585
R1388 B.n633 B.n120 585
R1389 B.n632 B.n631 585
R1390 B.n630 B.n121 585
R1391 B.n629 B.n628 585
R1392 B.n627 B.n122 585
R1393 B.n626 B.n625 585
R1394 B.n624 B.n123 585
R1395 B.n623 B.n622 585
R1396 B.n621 B.n124 585
R1397 B.n620 B.n619 585
R1398 B.n618 B.n125 585
R1399 B.n617 B.n616 585
R1400 B.n615 B.n126 585
R1401 B.n614 B.n613 585
R1402 B.n612 B.n127 585
R1403 B.n611 B.n610 585
R1404 B.n609 B.n128 585
R1405 B.n608 B.n607 585
R1406 B.n606 B.n129 585
R1407 B.n605 B.n604 585
R1408 B.n603 B.n130 585
R1409 B.n602 B.n601 585
R1410 B.n600 B.n131 585
R1411 B.n599 B.n598 585
R1412 B.n597 B.n132 585
R1413 B.n596 B.n595 585
R1414 B.n594 B.n133 585
R1415 B.n593 B.n592 585
R1416 B.n591 B.n134 585
R1417 B.n590 B.n589 585
R1418 B.n588 B.n135 585
R1419 B.n587 B.n586 585
R1420 B.n585 B.n136 585
R1421 B.n584 B.n583 585
R1422 B.n582 B.n137 585
R1423 B.n581 B.n580 585
R1424 B.n579 B.n138 585
R1425 B.n578 B.n577 585
R1426 B.n576 B.n139 585
R1427 B.n575 B.n574 585
R1428 B.n573 B.n140 585
R1429 B.n572 B.n571 585
R1430 B.n570 B.n141 585
R1431 B.n569 B.n568 585
R1432 B.n567 B.n142 585
R1433 B.n566 B.n565 585
R1434 B.n564 B.n143 585
R1435 B.n563 B.n562 585
R1436 B.n561 B.n144 585
R1437 B.n560 B.n559 585
R1438 B.n558 B.n145 585
R1439 B.n557 B.n556 585
R1440 B.n555 B.n146 585
R1441 B.n554 B.n553 585
R1442 B.n552 B.n147 585
R1443 B.n551 B.n550 585
R1444 B.n549 B.n148 585
R1445 B.n548 B.n547 585
R1446 B.n546 B.n149 585
R1447 B.n545 B.n544 585
R1448 B.n543 B.n150 585
R1449 B.n542 B.n541 585
R1450 B.n540 B.n151 585
R1451 B.n539 B.n538 585
R1452 B.n537 B.n152 585
R1453 B.n536 B.n535 585
R1454 B.n534 B.n153 585
R1455 B.n533 B.n532 585
R1456 B.n531 B.n154 585
R1457 B.n530 B.n529 585
R1458 B.n528 B.n155 585
R1459 B.n527 B.n526 585
R1460 B.n525 B.n156 585
R1461 B.n524 B.n523 585
R1462 B.n522 B.n157 585
R1463 B.n521 B.n520 585
R1464 B.n519 B.n158 585
R1465 B.n518 B.n517 585
R1466 B.n516 B.n159 585
R1467 B.n515 B.n514 585
R1468 B.n513 B.n160 585
R1469 B.n512 B.n511 585
R1470 B.n351 B.n218 585
R1471 B.n353 B.n352 585
R1472 B.n354 B.n217 585
R1473 B.n356 B.n355 585
R1474 B.n357 B.n216 585
R1475 B.n359 B.n358 585
R1476 B.n360 B.n215 585
R1477 B.n362 B.n361 585
R1478 B.n363 B.n214 585
R1479 B.n365 B.n364 585
R1480 B.n366 B.n213 585
R1481 B.n368 B.n367 585
R1482 B.n369 B.n212 585
R1483 B.n371 B.n370 585
R1484 B.n372 B.n211 585
R1485 B.n374 B.n373 585
R1486 B.n375 B.n210 585
R1487 B.n377 B.n376 585
R1488 B.n378 B.n209 585
R1489 B.n380 B.n379 585
R1490 B.n381 B.n208 585
R1491 B.n383 B.n382 585
R1492 B.n384 B.n207 585
R1493 B.n386 B.n385 585
R1494 B.n387 B.n206 585
R1495 B.n389 B.n388 585
R1496 B.n390 B.n205 585
R1497 B.n392 B.n391 585
R1498 B.n393 B.n204 585
R1499 B.n395 B.n394 585
R1500 B.n396 B.n203 585
R1501 B.n398 B.n397 585
R1502 B.n399 B.n202 585
R1503 B.n401 B.n400 585
R1504 B.n402 B.n201 585
R1505 B.n404 B.n403 585
R1506 B.n405 B.n200 585
R1507 B.n407 B.n406 585
R1508 B.n408 B.n199 585
R1509 B.n410 B.n409 585
R1510 B.n411 B.n198 585
R1511 B.n413 B.n412 585
R1512 B.n414 B.n197 585
R1513 B.n416 B.n415 585
R1514 B.n417 B.n196 585
R1515 B.n419 B.n418 585
R1516 B.n420 B.n195 585
R1517 B.n422 B.n421 585
R1518 B.n424 B.n192 585
R1519 B.n426 B.n425 585
R1520 B.n427 B.n191 585
R1521 B.n429 B.n428 585
R1522 B.n430 B.n190 585
R1523 B.n432 B.n431 585
R1524 B.n433 B.n189 585
R1525 B.n435 B.n434 585
R1526 B.n436 B.n188 585
R1527 B.n438 B.n437 585
R1528 B.n440 B.n439 585
R1529 B.n441 B.n184 585
R1530 B.n443 B.n442 585
R1531 B.n444 B.n183 585
R1532 B.n446 B.n445 585
R1533 B.n447 B.n182 585
R1534 B.n449 B.n448 585
R1535 B.n450 B.n181 585
R1536 B.n452 B.n451 585
R1537 B.n453 B.n180 585
R1538 B.n455 B.n454 585
R1539 B.n456 B.n179 585
R1540 B.n458 B.n457 585
R1541 B.n459 B.n178 585
R1542 B.n461 B.n460 585
R1543 B.n462 B.n177 585
R1544 B.n464 B.n463 585
R1545 B.n465 B.n176 585
R1546 B.n467 B.n466 585
R1547 B.n468 B.n175 585
R1548 B.n470 B.n469 585
R1549 B.n471 B.n174 585
R1550 B.n473 B.n472 585
R1551 B.n474 B.n173 585
R1552 B.n476 B.n475 585
R1553 B.n477 B.n172 585
R1554 B.n479 B.n478 585
R1555 B.n480 B.n171 585
R1556 B.n482 B.n481 585
R1557 B.n483 B.n170 585
R1558 B.n485 B.n484 585
R1559 B.n486 B.n169 585
R1560 B.n488 B.n487 585
R1561 B.n489 B.n168 585
R1562 B.n491 B.n490 585
R1563 B.n492 B.n167 585
R1564 B.n494 B.n493 585
R1565 B.n495 B.n166 585
R1566 B.n497 B.n496 585
R1567 B.n498 B.n165 585
R1568 B.n500 B.n499 585
R1569 B.n501 B.n164 585
R1570 B.n503 B.n502 585
R1571 B.n504 B.n163 585
R1572 B.n506 B.n505 585
R1573 B.n507 B.n162 585
R1574 B.n509 B.n508 585
R1575 B.n510 B.n161 585
R1576 B.n350 B.n349 585
R1577 B.n348 B.n219 585
R1578 B.n347 B.n346 585
R1579 B.n345 B.n220 585
R1580 B.n344 B.n343 585
R1581 B.n342 B.n221 585
R1582 B.n341 B.n340 585
R1583 B.n339 B.n222 585
R1584 B.n338 B.n337 585
R1585 B.n336 B.n223 585
R1586 B.n335 B.n334 585
R1587 B.n333 B.n224 585
R1588 B.n332 B.n331 585
R1589 B.n330 B.n225 585
R1590 B.n329 B.n328 585
R1591 B.n327 B.n226 585
R1592 B.n326 B.n325 585
R1593 B.n324 B.n227 585
R1594 B.n323 B.n322 585
R1595 B.n321 B.n228 585
R1596 B.n320 B.n319 585
R1597 B.n318 B.n229 585
R1598 B.n317 B.n316 585
R1599 B.n315 B.n230 585
R1600 B.n314 B.n313 585
R1601 B.n312 B.n231 585
R1602 B.n311 B.n310 585
R1603 B.n309 B.n232 585
R1604 B.n308 B.n307 585
R1605 B.n306 B.n233 585
R1606 B.n305 B.n304 585
R1607 B.n303 B.n234 585
R1608 B.n302 B.n301 585
R1609 B.n300 B.n235 585
R1610 B.n299 B.n298 585
R1611 B.n297 B.n236 585
R1612 B.n296 B.n295 585
R1613 B.n294 B.n237 585
R1614 B.n293 B.n292 585
R1615 B.n291 B.n238 585
R1616 B.n290 B.n289 585
R1617 B.n288 B.n239 585
R1618 B.n287 B.n286 585
R1619 B.n285 B.n240 585
R1620 B.n284 B.n283 585
R1621 B.n282 B.n241 585
R1622 B.n281 B.n280 585
R1623 B.n279 B.n242 585
R1624 B.n278 B.n277 585
R1625 B.n276 B.n243 585
R1626 B.n275 B.n274 585
R1627 B.n273 B.n244 585
R1628 B.n272 B.n271 585
R1629 B.n270 B.n245 585
R1630 B.n269 B.n268 585
R1631 B.n267 B.n246 585
R1632 B.n266 B.n265 585
R1633 B.n264 B.n247 585
R1634 B.n263 B.n262 585
R1635 B.n261 B.n248 585
R1636 B.n260 B.n259 585
R1637 B.n258 B.n249 585
R1638 B.n257 B.n256 585
R1639 B.n255 B.n250 585
R1640 B.n254 B.n253 585
R1641 B.n252 B.n251 585
R1642 B.n2 B.n0 585
R1643 B.n973 B.n1 585
R1644 B.n972 B.n971 585
R1645 B.n970 B.n3 585
R1646 B.n969 B.n968 585
R1647 B.n967 B.n4 585
R1648 B.n966 B.n965 585
R1649 B.n964 B.n5 585
R1650 B.n963 B.n962 585
R1651 B.n961 B.n6 585
R1652 B.n960 B.n959 585
R1653 B.n958 B.n7 585
R1654 B.n957 B.n956 585
R1655 B.n955 B.n8 585
R1656 B.n954 B.n953 585
R1657 B.n952 B.n9 585
R1658 B.n951 B.n950 585
R1659 B.n949 B.n10 585
R1660 B.n948 B.n947 585
R1661 B.n946 B.n11 585
R1662 B.n945 B.n944 585
R1663 B.n943 B.n12 585
R1664 B.n942 B.n941 585
R1665 B.n940 B.n13 585
R1666 B.n939 B.n938 585
R1667 B.n937 B.n14 585
R1668 B.n936 B.n935 585
R1669 B.n934 B.n15 585
R1670 B.n933 B.n932 585
R1671 B.n931 B.n16 585
R1672 B.n930 B.n929 585
R1673 B.n928 B.n17 585
R1674 B.n927 B.n926 585
R1675 B.n925 B.n18 585
R1676 B.n924 B.n923 585
R1677 B.n922 B.n19 585
R1678 B.n921 B.n920 585
R1679 B.n919 B.n20 585
R1680 B.n918 B.n917 585
R1681 B.n916 B.n21 585
R1682 B.n915 B.n914 585
R1683 B.n913 B.n22 585
R1684 B.n912 B.n911 585
R1685 B.n910 B.n23 585
R1686 B.n909 B.n908 585
R1687 B.n907 B.n24 585
R1688 B.n906 B.n905 585
R1689 B.n904 B.n25 585
R1690 B.n903 B.n902 585
R1691 B.n901 B.n26 585
R1692 B.n900 B.n899 585
R1693 B.n898 B.n27 585
R1694 B.n897 B.n896 585
R1695 B.n895 B.n28 585
R1696 B.n894 B.n893 585
R1697 B.n892 B.n29 585
R1698 B.n891 B.n890 585
R1699 B.n889 B.n30 585
R1700 B.n888 B.n887 585
R1701 B.n886 B.n31 585
R1702 B.n885 B.n884 585
R1703 B.n883 B.n32 585
R1704 B.n882 B.n881 585
R1705 B.n880 B.n33 585
R1706 B.n879 B.n878 585
R1707 B.n877 B.n34 585
R1708 B.n876 B.n875 585
R1709 B.n874 B.n35 585
R1710 B.n975 B.n974 585
R1711 B.n185 B.t5 492.37
R1712 B.n68 B.t7 492.37
R1713 B.n193 B.t2 492.37
R1714 B.n60 B.t10 492.37
R1715 B.n349 B.n218 454.062
R1716 B.n872 B.n35 454.062
R1717 B.n511 B.n510 454.062
R1718 B.n714 B.n713 454.062
R1719 B.n186 B.t4 414.793
R1720 B.n69 B.t8 414.793
R1721 B.n194 B.t1 414.793
R1722 B.n61 B.t11 414.793
R1723 B.n185 B.t3 302.291
R1724 B.n193 B.t0 302.291
R1725 B.n60 B.t9 302.291
R1726 B.n68 B.t6 302.291
R1727 B.n349 B.n348 163.367
R1728 B.n348 B.n347 163.367
R1729 B.n347 B.n220 163.367
R1730 B.n343 B.n220 163.367
R1731 B.n343 B.n342 163.367
R1732 B.n342 B.n341 163.367
R1733 B.n341 B.n222 163.367
R1734 B.n337 B.n222 163.367
R1735 B.n337 B.n336 163.367
R1736 B.n336 B.n335 163.367
R1737 B.n335 B.n224 163.367
R1738 B.n331 B.n224 163.367
R1739 B.n331 B.n330 163.367
R1740 B.n330 B.n329 163.367
R1741 B.n329 B.n226 163.367
R1742 B.n325 B.n226 163.367
R1743 B.n325 B.n324 163.367
R1744 B.n324 B.n323 163.367
R1745 B.n323 B.n228 163.367
R1746 B.n319 B.n228 163.367
R1747 B.n319 B.n318 163.367
R1748 B.n318 B.n317 163.367
R1749 B.n317 B.n230 163.367
R1750 B.n313 B.n230 163.367
R1751 B.n313 B.n312 163.367
R1752 B.n312 B.n311 163.367
R1753 B.n311 B.n232 163.367
R1754 B.n307 B.n232 163.367
R1755 B.n307 B.n306 163.367
R1756 B.n306 B.n305 163.367
R1757 B.n305 B.n234 163.367
R1758 B.n301 B.n234 163.367
R1759 B.n301 B.n300 163.367
R1760 B.n300 B.n299 163.367
R1761 B.n299 B.n236 163.367
R1762 B.n295 B.n236 163.367
R1763 B.n295 B.n294 163.367
R1764 B.n294 B.n293 163.367
R1765 B.n293 B.n238 163.367
R1766 B.n289 B.n238 163.367
R1767 B.n289 B.n288 163.367
R1768 B.n288 B.n287 163.367
R1769 B.n287 B.n240 163.367
R1770 B.n283 B.n240 163.367
R1771 B.n283 B.n282 163.367
R1772 B.n282 B.n281 163.367
R1773 B.n281 B.n242 163.367
R1774 B.n277 B.n242 163.367
R1775 B.n277 B.n276 163.367
R1776 B.n276 B.n275 163.367
R1777 B.n275 B.n244 163.367
R1778 B.n271 B.n244 163.367
R1779 B.n271 B.n270 163.367
R1780 B.n270 B.n269 163.367
R1781 B.n269 B.n246 163.367
R1782 B.n265 B.n246 163.367
R1783 B.n265 B.n264 163.367
R1784 B.n264 B.n263 163.367
R1785 B.n263 B.n248 163.367
R1786 B.n259 B.n248 163.367
R1787 B.n259 B.n258 163.367
R1788 B.n258 B.n257 163.367
R1789 B.n257 B.n250 163.367
R1790 B.n253 B.n250 163.367
R1791 B.n253 B.n252 163.367
R1792 B.n252 B.n2 163.367
R1793 B.n974 B.n2 163.367
R1794 B.n974 B.n973 163.367
R1795 B.n973 B.n972 163.367
R1796 B.n972 B.n3 163.367
R1797 B.n968 B.n3 163.367
R1798 B.n968 B.n967 163.367
R1799 B.n967 B.n966 163.367
R1800 B.n966 B.n5 163.367
R1801 B.n962 B.n5 163.367
R1802 B.n962 B.n961 163.367
R1803 B.n961 B.n960 163.367
R1804 B.n960 B.n7 163.367
R1805 B.n956 B.n7 163.367
R1806 B.n956 B.n955 163.367
R1807 B.n955 B.n954 163.367
R1808 B.n954 B.n9 163.367
R1809 B.n950 B.n9 163.367
R1810 B.n950 B.n949 163.367
R1811 B.n949 B.n948 163.367
R1812 B.n948 B.n11 163.367
R1813 B.n944 B.n11 163.367
R1814 B.n944 B.n943 163.367
R1815 B.n943 B.n942 163.367
R1816 B.n942 B.n13 163.367
R1817 B.n938 B.n13 163.367
R1818 B.n938 B.n937 163.367
R1819 B.n937 B.n936 163.367
R1820 B.n936 B.n15 163.367
R1821 B.n932 B.n15 163.367
R1822 B.n932 B.n931 163.367
R1823 B.n931 B.n930 163.367
R1824 B.n930 B.n17 163.367
R1825 B.n926 B.n17 163.367
R1826 B.n926 B.n925 163.367
R1827 B.n925 B.n924 163.367
R1828 B.n924 B.n19 163.367
R1829 B.n920 B.n19 163.367
R1830 B.n920 B.n919 163.367
R1831 B.n919 B.n918 163.367
R1832 B.n918 B.n21 163.367
R1833 B.n914 B.n21 163.367
R1834 B.n914 B.n913 163.367
R1835 B.n913 B.n912 163.367
R1836 B.n912 B.n23 163.367
R1837 B.n908 B.n23 163.367
R1838 B.n908 B.n907 163.367
R1839 B.n907 B.n906 163.367
R1840 B.n906 B.n25 163.367
R1841 B.n902 B.n25 163.367
R1842 B.n902 B.n901 163.367
R1843 B.n901 B.n900 163.367
R1844 B.n900 B.n27 163.367
R1845 B.n896 B.n27 163.367
R1846 B.n896 B.n895 163.367
R1847 B.n895 B.n894 163.367
R1848 B.n894 B.n29 163.367
R1849 B.n890 B.n29 163.367
R1850 B.n890 B.n889 163.367
R1851 B.n889 B.n888 163.367
R1852 B.n888 B.n31 163.367
R1853 B.n884 B.n31 163.367
R1854 B.n884 B.n883 163.367
R1855 B.n883 B.n882 163.367
R1856 B.n882 B.n33 163.367
R1857 B.n878 B.n33 163.367
R1858 B.n878 B.n877 163.367
R1859 B.n877 B.n876 163.367
R1860 B.n876 B.n35 163.367
R1861 B.n353 B.n218 163.367
R1862 B.n354 B.n353 163.367
R1863 B.n355 B.n354 163.367
R1864 B.n355 B.n216 163.367
R1865 B.n359 B.n216 163.367
R1866 B.n360 B.n359 163.367
R1867 B.n361 B.n360 163.367
R1868 B.n361 B.n214 163.367
R1869 B.n365 B.n214 163.367
R1870 B.n366 B.n365 163.367
R1871 B.n367 B.n366 163.367
R1872 B.n367 B.n212 163.367
R1873 B.n371 B.n212 163.367
R1874 B.n372 B.n371 163.367
R1875 B.n373 B.n372 163.367
R1876 B.n373 B.n210 163.367
R1877 B.n377 B.n210 163.367
R1878 B.n378 B.n377 163.367
R1879 B.n379 B.n378 163.367
R1880 B.n379 B.n208 163.367
R1881 B.n383 B.n208 163.367
R1882 B.n384 B.n383 163.367
R1883 B.n385 B.n384 163.367
R1884 B.n385 B.n206 163.367
R1885 B.n389 B.n206 163.367
R1886 B.n390 B.n389 163.367
R1887 B.n391 B.n390 163.367
R1888 B.n391 B.n204 163.367
R1889 B.n395 B.n204 163.367
R1890 B.n396 B.n395 163.367
R1891 B.n397 B.n396 163.367
R1892 B.n397 B.n202 163.367
R1893 B.n401 B.n202 163.367
R1894 B.n402 B.n401 163.367
R1895 B.n403 B.n402 163.367
R1896 B.n403 B.n200 163.367
R1897 B.n407 B.n200 163.367
R1898 B.n408 B.n407 163.367
R1899 B.n409 B.n408 163.367
R1900 B.n409 B.n198 163.367
R1901 B.n413 B.n198 163.367
R1902 B.n414 B.n413 163.367
R1903 B.n415 B.n414 163.367
R1904 B.n415 B.n196 163.367
R1905 B.n419 B.n196 163.367
R1906 B.n420 B.n419 163.367
R1907 B.n421 B.n420 163.367
R1908 B.n421 B.n192 163.367
R1909 B.n426 B.n192 163.367
R1910 B.n427 B.n426 163.367
R1911 B.n428 B.n427 163.367
R1912 B.n428 B.n190 163.367
R1913 B.n432 B.n190 163.367
R1914 B.n433 B.n432 163.367
R1915 B.n434 B.n433 163.367
R1916 B.n434 B.n188 163.367
R1917 B.n438 B.n188 163.367
R1918 B.n439 B.n438 163.367
R1919 B.n439 B.n184 163.367
R1920 B.n443 B.n184 163.367
R1921 B.n444 B.n443 163.367
R1922 B.n445 B.n444 163.367
R1923 B.n445 B.n182 163.367
R1924 B.n449 B.n182 163.367
R1925 B.n450 B.n449 163.367
R1926 B.n451 B.n450 163.367
R1927 B.n451 B.n180 163.367
R1928 B.n455 B.n180 163.367
R1929 B.n456 B.n455 163.367
R1930 B.n457 B.n456 163.367
R1931 B.n457 B.n178 163.367
R1932 B.n461 B.n178 163.367
R1933 B.n462 B.n461 163.367
R1934 B.n463 B.n462 163.367
R1935 B.n463 B.n176 163.367
R1936 B.n467 B.n176 163.367
R1937 B.n468 B.n467 163.367
R1938 B.n469 B.n468 163.367
R1939 B.n469 B.n174 163.367
R1940 B.n473 B.n174 163.367
R1941 B.n474 B.n473 163.367
R1942 B.n475 B.n474 163.367
R1943 B.n475 B.n172 163.367
R1944 B.n479 B.n172 163.367
R1945 B.n480 B.n479 163.367
R1946 B.n481 B.n480 163.367
R1947 B.n481 B.n170 163.367
R1948 B.n485 B.n170 163.367
R1949 B.n486 B.n485 163.367
R1950 B.n487 B.n486 163.367
R1951 B.n487 B.n168 163.367
R1952 B.n491 B.n168 163.367
R1953 B.n492 B.n491 163.367
R1954 B.n493 B.n492 163.367
R1955 B.n493 B.n166 163.367
R1956 B.n497 B.n166 163.367
R1957 B.n498 B.n497 163.367
R1958 B.n499 B.n498 163.367
R1959 B.n499 B.n164 163.367
R1960 B.n503 B.n164 163.367
R1961 B.n504 B.n503 163.367
R1962 B.n505 B.n504 163.367
R1963 B.n505 B.n162 163.367
R1964 B.n509 B.n162 163.367
R1965 B.n510 B.n509 163.367
R1966 B.n511 B.n160 163.367
R1967 B.n515 B.n160 163.367
R1968 B.n516 B.n515 163.367
R1969 B.n517 B.n516 163.367
R1970 B.n517 B.n158 163.367
R1971 B.n521 B.n158 163.367
R1972 B.n522 B.n521 163.367
R1973 B.n523 B.n522 163.367
R1974 B.n523 B.n156 163.367
R1975 B.n527 B.n156 163.367
R1976 B.n528 B.n527 163.367
R1977 B.n529 B.n528 163.367
R1978 B.n529 B.n154 163.367
R1979 B.n533 B.n154 163.367
R1980 B.n534 B.n533 163.367
R1981 B.n535 B.n534 163.367
R1982 B.n535 B.n152 163.367
R1983 B.n539 B.n152 163.367
R1984 B.n540 B.n539 163.367
R1985 B.n541 B.n540 163.367
R1986 B.n541 B.n150 163.367
R1987 B.n545 B.n150 163.367
R1988 B.n546 B.n545 163.367
R1989 B.n547 B.n546 163.367
R1990 B.n547 B.n148 163.367
R1991 B.n551 B.n148 163.367
R1992 B.n552 B.n551 163.367
R1993 B.n553 B.n552 163.367
R1994 B.n553 B.n146 163.367
R1995 B.n557 B.n146 163.367
R1996 B.n558 B.n557 163.367
R1997 B.n559 B.n558 163.367
R1998 B.n559 B.n144 163.367
R1999 B.n563 B.n144 163.367
R2000 B.n564 B.n563 163.367
R2001 B.n565 B.n564 163.367
R2002 B.n565 B.n142 163.367
R2003 B.n569 B.n142 163.367
R2004 B.n570 B.n569 163.367
R2005 B.n571 B.n570 163.367
R2006 B.n571 B.n140 163.367
R2007 B.n575 B.n140 163.367
R2008 B.n576 B.n575 163.367
R2009 B.n577 B.n576 163.367
R2010 B.n577 B.n138 163.367
R2011 B.n581 B.n138 163.367
R2012 B.n582 B.n581 163.367
R2013 B.n583 B.n582 163.367
R2014 B.n583 B.n136 163.367
R2015 B.n587 B.n136 163.367
R2016 B.n588 B.n587 163.367
R2017 B.n589 B.n588 163.367
R2018 B.n589 B.n134 163.367
R2019 B.n593 B.n134 163.367
R2020 B.n594 B.n593 163.367
R2021 B.n595 B.n594 163.367
R2022 B.n595 B.n132 163.367
R2023 B.n599 B.n132 163.367
R2024 B.n600 B.n599 163.367
R2025 B.n601 B.n600 163.367
R2026 B.n601 B.n130 163.367
R2027 B.n605 B.n130 163.367
R2028 B.n606 B.n605 163.367
R2029 B.n607 B.n606 163.367
R2030 B.n607 B.n128 163.367
R2031 B.n611 B.n128 163.367
R2032 B.n612 B.n611 163.367
R2033 B.n613 B.n612 163.367
R2034 B.n613 B.n126 163.367
R2035 B.n617 B.n126 163.367
R2036 B.n618 B.n617 163.367
R2037 B.n619 B.n618 163.367
R2038 B.n619 B.n124 163.367
R2039 B.n623 B.n124 163.367
R2040 B.n624 B.n623 163.367
R2041 B.n625 B.n624 163.367
R2042 B.n625 B.n122 163.367
R2043 B.n629 B.n122 163.367
R2044 B.n630 B.n629 163.367
R2045 B.n631 B.n630 163.367
R2046 B.n631 B.n120 163.367
R2047 B.n635 B.n120 163.367
R2048 B.n636 B.n635 163.367
R2049 B.n637 B.n636 163.367
R2050 B.n637 B.n118 163.367
R2051 B.n641 B.n118 163.367
R2052 B.n642 B.n641 163.367
R2053 B.n643 B.n642 163.367
R2054 B.n643 B.n116 163.367
R2055 B.n647 B.n116 163.367
R2056 B.n648 B.n647 163.367
R2057 B.n649 B.n648 163.367
R2058 B.n649 B.n114 163.367
R2059 B.n653 B.n114 163.367
R2060 B.n654 B.n653 163.367
R2061 B.n655 B.n654 163.367
R2062 B.n655 B.n112 163.367
R2063 B.n659 B.n112 163.367
R2064 B.n660 B.n659 163.367
R2065 B.n661 B.n660 163.367
R2066 B.n661 B.n110 163.367
R2067 B.n665 B.n110 163.367
R2068 B.n666 B.n665 163.367
R2069 B.n667 B.n666 163.367
R2070 B.n667 B.n108 163.367
R2071 B.n671 B.n108 163.367
R2072 B.n672 B.n671 163.367
R2073 B.n673 B.n672 163.367
R2074 B.n673 B.n106 163.367
R2075 B.n677 B.n106 163.367
R2076 B.n678 B.n677 163.367
R2077 B.n679 B.n678 163.367
R2078 B.n679 B.n104 163.367
R2079 B.n683 B.n104 163.367
R2080 B.n684 B.n683 163.367
R2081 B.n685 B.n684 163.367
R2082 B.n685 B.n102 163.367
R2083 B.n689 B.n102 163.367
R2084 B.n690 B.n689 163.367
R2085 B.n691 B.n690 163.367
R2086 B.n691 B.n100 163.367
R2087 B.n695 B.n100 163.367
R2088 B.n696 B.n695 163.367
R2089 B.n697 B.n696 163.367
R2090 B.n697 B.n98 163.367
R2091 B.n701 B.n98 163.367
R2092 B.n702 B.n701 163.367
R2093 B.n703 B.n702 163.367
R2094 B.n703 B.n96 163.367
R2095 B.n707 B.n96 163.367
R2096 B.n708 B.n707 163.367
R2097 B.n709 B.n708 163.367
R2098 B.n709 B.n94 163.367
R2099 B.n713 B.n94 163.367
R2100 B.n872 B.n871 163.367
R2101 B.n871 B.n870 163.367
R2102 B.n870 B.n37 163.367
R2103 B.n866 B.n37 163.367
R2104 B.n866 B.n865 163.367
R2105 B.n865 B.n864 163.367
R2106 B.n864 B.n39 163.367
R2107 B.n860 B.n39 163.367
R2108 B.n860 B.n859 163.367
R2109 B.n859 B.n858 163.367
R2110 B.n858 B.n41 163.367
R2111 B.n854 B.n41 163.367
R2112 B.n854 B.n853 163.367
R2113 B.n853 B.n852 163.367
R2114 B.n852 B.n43 163.367
R2115 B.n848 B.n43 163.367
R2116 B.n848 B.n847 163.367
R2117 B.n847 B.n846 163.367
R2118 B.n846 B.n45 163.367
R2119 B.n842 B.n45 163.367
R2120 B.n842 B.n841 163.367
R2121 B.n841 B.n840 163.367
R2122 B.n840 B.n47 163.367
R2123 B.n836 B.n47 163.367
R2124 B.n836 B.n835 163.367
R2125 B.n835 B.n834 163.367
R2126 B.n834 B.n49 163.367
R2127 B.n830 B.n49 163.367
R2128 B.n830 B.n829 163.367
R2129 B.n829 B.n828 163.367
R2130 B.n828 B.n51 163.367
R2131 B.n824 B.n51 163.367
R2132 B.n824 B.n823 163.367
R2133 B.n823 B.n822 163.367
R2134 B.n822 B.n53 163.367
R2135 B.n818 B.n53 163.367
R2136 B.n818 B.n817 163.367
R2137 B.n817 B.n816 163.367
R2138 B.n816 B.n55 163.367
R2139 B.n812 B.n55 163.367
R2140 B.n812 B.n811 163.367
R2141 B.n811 B.n810 163.367
R2142 B.n810 B.n57 163.367
R2143 B.n806 B.n57 163.367
R2144 B.n806 B.n805 163.367
R2145 B.n805 B.n804 163.367
R2146 B.n804 B.n59 163.367
R2147 B.n799 B.n59 163.367
R2148 B.n799 B.n798 163.367
R2149 B.n798 B.n797 163.367
R2150 B.n797 B.n63 163.367
R2151 B.n793 B.n63 163.367
R2152 B.n793 B.n792 163.367
R2153 B.n792 B.n791 163.367
R2154 B.n791 B.n65 163.367
R2155 B.n787 B.n65 163.367
R2156 B.n787 B.n786 163.367
R2157 B.n786 B.n785 163.367
R2158 B.n785 B.n67 163.367
R2159 B.n781 B.n67 163.367
R2160 B.n781 B.n780 163.367
R2161 B.n780 B.n779 163.367
R2162 B.n779 B.n72 163.367
R2163 B.n775 B.n72 163.367
R2164 B.n775 B.n774 163.367
R2165 B.n774 B.n773 163.367
R2166 B.n773 B.n74 163.367
R2167 B.n769 B.n74 163.367
R2168 B.n769 B.n768 163.367
R2169 B.n768 B.n767 163.367
R2170 B.n767 B.n76 163.367
R2171 B.n763 B.n76 163.367
R2172 B.n763 B.n762 163.367
R2173 B.n762 B.n761 163.367
R2174 B.n761 B.n78 163.367
R2175 B.n757 B.n78 163.367
R2176 B.n757 B.n756 163.367
R2177 B.n756 B.n755 163.367
R2178 B.n755 B.n80 163.367
R2179 B.n751 B.n80 163.367
R2180 B.n751 B.n750 163.367
R2181 B.n750 B.n749 163.367
R2182 B.n749 B.n82 163.367
R2183 B.n745 B.n82 163.367
R2184 B.n745 B.n744 163.367
R2185 B.n744 B.n743 163.367
R2186 B.n743 B.n84 163.367
R2187 B.n739 B.n84 163.367
R2188 B.n739 B.n738 163.367
R2189 B.n738 B.n737 163.367
R2190 B.n737 B.n86 163.367
R2191 B.n733 B.n86 163.367
R2192 B.n733 B.n732 163.367
R2193 B.n732 B.n731 163.367
R2194 B.n731 B.n88 163.367
R2195 B.n727 B.n88 163.367
R2196 B.n727 B.n726 163.367
R2197 B.n726 B.n725 163.367
R2198 B.n725 B.n90 163.367
R2199 B.n721 B.n90 163.367
R2200 B.n721 B.n720 163.367
R2201 B.n720 B.n719 163.367
R2202 B.n719 B.n92 163.367
R2203 B.n715 B.n92 163.367
R2204 B.n715 B.n714 163.367
R2205 B.n186 B.n185 77.5763
R2206 B.n194 B.n193 77.5763
R2207 B.n61 B.n60 77.5763
R2208 B.n69 B.n68 77.5763
R2209 B.n187 B.n186 59.5399
R2210 B.n423 B.n194 59.5399
R2211 B.n801 B.n61 59.5399
R2212 B.n70 B.n69 59.5399
R2213 B.n712 B.n93 29.5029
R2214 B.n874 B.n873 29.5029
R2215 B.n512 B.n161 29.5029
R2216 B.n351 B.n350 29.5029
R2217 B B.n975 18.0485
R2218 B.n873 B.n36 10.6151
R2219 B.n869 B.n36 10.6151
R2220 B.n869 B.n868 10.6151
R2221 B.n868 B.n867 10.6151
R2222 B.n867 B.n38 10.6151
R2223 B.n863 B.n38 10.6151
R2224 B.n863 B.n862 10.6151
R2225 B.n862 B.n861 10.6151
R2226 B.n861 B.n40 10.6151
R2227 B.n857 B.n40 10.6151
R2228 B.n857 B.n856 10.6151
R2229 B.n856 B.n855 10.6151
R2230 B.n855 B.n42 10.6151
R2231 B.n851 B.n42 10.6151
R2232 B.n851 B.n850 10.6151
R2233 B.n850 B.n849 10.6151
R2234 B.n849 B.n44 10.6151
R2235 B.n845 B.n44 10.6151
R2236 B.n845 B.n844 10.6151
R2237 B.n844 B.n843 10.6151
R2238 B.n843 B.n46 10.6151
R2239 B.n839 B.n46 10.6151
R2240 B.n839 B.n838 10.6151
R2241 B.n838 B.n837 10.6151
R2242 B.n837 B.n48 10.6151
R2243 B.n833 B.n48 10.6151
R2244 B.n833 B.n832 10.6151
R2245 B.n832 B.n831 10.6151
R2246 B.n831 B.n50 10.6151
R2247 B.n827 B.n50 10.6151
R2248 B.n827 B.n826 10.6151
R2249 B.n826 B.n825 10.6151
R2250 B.n825 B.n52 10.6151
R2251 B.n821 B.n52 10.6151
R2252 B.n821 B.n820 10.6151
R2253 B.n820 B.n819 10.6151
R2254 B.n819 B.n54 10.6151
R2255 B.n815 B.n54 10.6151
R2256 B.n815 B.n814 10.6151
R2257 B.n814 B.n813 10.6151
R2258 B.n813 B.n56 10.6151
R2259 B.n809 B.n56 10.6151
R2260 B.n809 B.n808 10.6151
R2261 B.n808 B.n807 10.6151
R2262 B.n807 B.n58 10.6151
R2263 B.n803 B.n58 10.6151
R2264 B.n803 B.n802 10.6151
R2265 B.n800 B.n62 10.6151
R2266 B.n796 B.n62 10.6151
R2267 B.n796 B.n795 10.6151
R2268 B.n795 B.n794 10.6151
R2269 B.n794 B.n64 10.6151
R2270 B.n790 B.n64 10.6151
R2271 B.n790 B.n789 10.6151
R2272 B.n789 B.n788 10.6151
R2273 B.n788 B.n66 10.6151
R2274 B.n784 B.n783 10.6151
R2275 B.n783 B.n782 10.6151
R2276 B.n782 B.n71 10.6151
R2277 B.n778 B.n71 10.6151
R2278 B.n778 B.n777 10.6151
R2279 B.n777 B.n776 10.6151
R2280 B.n776 B.n73 10.6151
R2281 B.n772 B.n73 10.6151
R2282 B.n772 B.n771 10.6151
R2283 B.n771 B.n770 10.6151
R2284 B.n770 B.n75 10.6151
R2285 B.n766 B.n75 10.6151
R2286 B.n766 B.n765 10.6151
R2287 B.n765 B.n764 10.6151
R2288 B.n764 B.n77 10.6151
R2289 B.n760 B.n77 10.6151
R2290 B.n760 B.n759 10.6151
R2291 B.n759 B.n758 10.6151
R2292 B.n758 B.n79 10.6151
R2293 B.n754 B.n79 10.6151
R2294 B.n754 B.n753 10.6151
R2295 B.n753 B.n752 10.6151
R2296 B.n752 B.n81 10.6151
R2297 B.n748 B.n81 10.6151
R2298 B.n748 B.n747 10.6151
R2299 B.n747 B.n746 10.6151
R2300 B.n746 B.n83 10.6151
R2301 B.n742 B.n83 10.6151
R2302 B.n742 B.n741 10.6151
R2303 B.n741 B.n740 10.6151
R2304 B.n740 B.n85 10.6151
R2305 B.n736 B.n85 10.6151
R2306 B.n736 B.n735 10.6151
R2307 B.n735 B.n734 10.6151
R2308 B.n734 B.n87 10.6151
R2309 B.n730 B.n87 10.6151
R2310 B.n730 B.n729 10.6151
R2311 B.n729 B.n728 10.6151
R2312 B.n728 B.n89 10.6151
R2313 B.n724 B.n89 10.6151
R2314 B.n724 B.n723 10.6151
R2315 B.n723 B.n722 10.6151
R2316 B.n722 B.n91 10.6151
R2317 B.n718 B.n91 10.6151
R2318 B.n718 B.n717 10.6151
R2319 B.n717 B.n716 10.6151
R2320 B.n716 B.n93 10.6151
R2321 B.n513 B.n512 10.6151
R2322 B.n514 B.n513 10.6151
R2323 B.n514 B.n159 10.6151
R2324 B.n518 B.n159 10.6151
R2325 B.n519 B.n518 10.6151
R2326 B.n520 B.n519 10.6151
R2327 B.n520 B.n157 10.6151
R2328 B.n524 B.n157 10.6151
R2329 B.n525 B.n524 10.6151
R2330 B.n526 B.n525 10.6151
R2331 B.n526 B.n155 10.6151
R2332 B.n530 B.n155 10.6151
R2333 B.n531 B.n530 10.6151
R2334 B.n532 B.n531 10.6151
R2335 B.n532 B.n153 10.6151
R2336 B.n536 B.n153 10.6151
R2337 B.n537 B.n536 10.6151
R2338 B.n538 B.n537 10.6151
R2339 B.n538 B.n151 10.6151
R2340 B.n542 B.n151 10.6151
R2341 B.n543 B.n542 10.6151
R2342 B.n544 B.n543 10.6151
R2343 B.n544 B.n149 10.6151
R2344 B.n548 B.n149 10.6151
R2345 B.n549 B.n548 10.6151
R2346 B.n550 B.n549 10.6151
R2347 B.n550 B.n147 10.6151
R2348 B.n554 B.n147 10.6151
R2349 B.n555 B.n554 10.6151
R2350 B.n556 B.n555 10.6151
R2351 B.n556 B.n145 10.6151
R2352 B.n560 B.n145 10.6151
R2353 B.n561 B.n560 10.6151
R2354 B.n562 B.n561 10.6151
R2355 B.n562 B.n143 10.6151
R2356 B.n566 B.n143 10.6151
R2357 B.n567 B.n566 10.6151
R2358 B.n568 B.n567 10.6151
R2359 B.n568 B.n141 10.6151
R2360 B.n572 B.n141 10.6151
R2361 B.n573 B.n572 10.6151
R2362 B.n574 B.n573 10.6151
R2363 B.n574 B.n139 10.6151
R2364 B.n578 B.n139 10.6151
R2365 B.n579 B.n578 10.6151
R2366 B.n580 B.n579 10.6151
R2367 B.n580 B.n137 10.6151
R2368 B.n584 B.n137 10.6151
R2369 B.n585 B.n584 10.6151
R2370 B.n586 B.n585 10.6151
R2371 B.n586 B.n135 10.6151
R2372 B.n590 B.n135 10.6151
R2373 B.n591 B.n590 10.6151
R2374 B.n592 B.n591 10.6151
R2375 B.n592 B.n133 10.6151
R2376 B.n596 B.n133 10.6151
R2377 B.n597 B.n596 10.6151
R2378 B.n598 B.n597 10.6151
R2379 B.n598 B.n131 10.6151
R2380 B.n602 B.n131 10.6151
R2381 B.n603 B.n602 10.6151
R2382 B.n604 B.n603 10.6151
R2383 B.n604 B.n129 10.6151
R2384 B.n608 B.n129 10.6151
R2385 B.n609 B.n608 10.6151
R2386 B.n610 B.n609 10.6151
R2387 B.n610 B.n127 10.6151
R2388 B.n614 B.n127 10.6151
R2389 B.n615 B.n614 10.6151
R2390 B.n616 B.n615 10.6151
R2391 B.n616 B.n125 10.6151
R2392 B.n620 B.n125 10.6151
R2393 B.n621 B.n620 10.6151
R2394 B.n622 B.n621 10.6151
R2395 B.n622 B.n123 10.6151
R2396 B.n626 B.n123 10.6151
R2397 B.n627 B.n626 10.6151
R2398 B.n628 B.n627 10.6151
R2399 B.n628 B.n121 10.6151
R2400 B.n632 B.n121 10.6151
R2401 B.n633 B.n632 10.6151
R2402 B.n634 B.n633 10.6151
R2403 B.n634 B.n119 10.6151
R2404 B.n638 B.n119 10.6151
R2405 B.n639 B.n638 10.6151
R2406 B.n640 B.n639 10.6151
R2407 B.n640 B.n117 10.6151
R2408 B.n644 B.n117 10.6151
R2409 B.n645 B.n644 10.6151
R2410 B.n646 B.n645 10.6151
R2411 B.n646 B.n115 10.6151
R2412 B.n650 B.n115 10.6151
R2413 B.n651 B.n650 10.6151
R2414 B.n652 B.n651 10.6151
R2415 B.n652 B.n113 10.6151
R2416 B.n656 B.n113 10.6151
R2417 B.n657 B.n656 10.6151
R2418 B.n658 B.n657 10.6151
R2419 B.n658 B.n111 10.6151
R2420 B.n662 B.n111 10.6151
R2421 B.n663 B.n662 10.6151
R2422 B.n664 B.n663 10.6151
R2423 B.n664 B.n109 10.6151
R2424 B.n668 B.n109 10.6151
R2425 B.n669 B.n668 10.6151
R2426 B.n670 B.n669 10.6151
R2427 B.n670 B.n107 10.6151
R2428 B.n674 B.n107 10.6151
R2429 B.n675 B.n674 10.6151
R2430 B.n676 B.n675 10.6151
R2431 B.n676 B.n105 10.6151
R2432 B.n680 B.n105 10.6151
R2433 B.n681 B.n680 10.6151
R2434 B.n682 B.n681 10.6151
R2435 B.n682 B.n103 10.6151
R2436 B.n686 B.n103 10.6151
R2437 B.n687 B.n686 10.6151
R2438 B.n688 B.n687 10.6151
R2439 B.n688 B.n101 10.6151
R2440 B.n692 B.n101 10.6151
R2441 B.n693 B.n692 10.6151
R2442 B.n694 B.n693 10.6151
R2443 B.n694 B.n99 10.6151
R2444 B.n698 B.n99 10.6151
R2445 B.n699 B.n698 10.6151
R2446 B.n700 B.n699 10.6151
R2447 B.n700 B.n97 10.6151
R2448 B.n704 B.n97 10.6151
R2449 B.n705 B.n704 10.6151
R2450 B.n706 B.n705 10.6151
R2451 B.n706 B.n95 10.6151
R2452 B.n710 B.n95 10.6151
R2453 B.n711 B.n710 10.6151
R2454 B.n712 B.n711 10.6151
R2455 B.n352 B.n351 10.6151
R2456 B.n352 B.n217 10.6151
R2457 B.n356 B.n217 10.6151
R2458 B.n357 B.n356 10.6151
R2459 B.n358 B.n357 10.6151
R2460 B.n358 B.n215 10.6151
R2461 B.n362 B.n215 10.6151
R2462 B.n363 B.n362 10.6151
R2463 B.n364 B.n363 10.6151
R2464 B.n364 B.n213 10.6151
R2465 B.n368 B.n213 10.6151
R2466 B.n369 B.n368 10.6151
R2467 B.n370 B.n369 10.6151
R2468 B.n370 B.n211 10.6151
R2469 B.n374 B.n211 10.6151
R2470 B.n375 B.n374 10.6151
R2471 B.n376 B.n375 10.6151
R2472 B.n376 B.n209 10.6151
R2473 B.n380 B.n209 10.6151
R2474 B.n381 B.n380 10.6151
R2475 B.n382 B.n381 10.6151
R2476 B.n382 B.n207 10.6151
R2477 B.n386 B.n207 10.6151
R2478 B.n387 B.n386 10.6151
R2479 B.n388 B.n387 10.6151
R2480 B.n388 B.n205 10.6151
R2481 B.n392 B.n205 10.6151
R2482 B.n393 B.n392 10.6151
R2483 B.n394 B.n393 10.6151
R2484 B.n394 B.n203 10.6151
R2485 B.n398 B.n203 10.6151
R2486 B.n399 B.n398 10.6151
R2487 B.n400 B.n399 10.6151
R2488 B.n400 B.n201 10.6151
R2489 B.n404 B.n201 10.6151
R2490 B.n405 B.n404 10.6151
R2491 B.n406 B.n405 10.6151
R2492 B.n406 B.n199 10.6151
R2493 B.n410 B.n199 10.6151
R2494 B.n411 B.n410 10.6151
R2495 B.n412 B.n411 10.6151
R2496 B.n412 B.n197 10.6151
R2497 B.n416 B.n197 10.6151
R2498 B.n417 B.n416 10.6151
R2499 B.n418 B.n417 10.6151
R2500 B.n418 B.n195 10.6151
R2501 B.n422 B.n195 10.6151
R2502 B.n425 B.n424 10.6151
R2503 B.n425 B.n191 10.6151
R2504 B.n429 B.n191 10.6151
R2505 B.n430 B.n429 10.6151
R2506 B.n431 B.n430 10.6151
R2507 B.n431 B.n189 10.6151
R2508 B.n435 B.n189 10.6151
R2509 B.n436 B.n435 10.6151
R2510 B.n437 B.n436 10.6151
R2511 B.n441 B.n440 10.6151
R2512 B.n442 B.n441 10.6151
R2513 B.n442 B.n183 10.6151
R2514 B.n446 B.n183 10.6151
R2515 B.n447 B.n446 10.6151
R2516 B.n448 B.n447 10.6151
R2517 B.n448 B.n181 10.6151
R2518 B.n452 B.n181 10.6151
R2519 B.n453 B.n452 10.6151
R2520 B.n454 B.n453 10.6151
R2521 B.n454 B.n179 10.6151
R2522 B.n458 B.n179 10.6151
R2523 B.n459 B.n458 10.6151
R2524 B.n460 B.n459 10.6151
R2525 B.n460 B.n177 10.6151
R2526 B.n464 B.n177 10.6151
R2527 B.n465 B.n464 10.6151
R2528 B.n466 B.n465 10.6151
R2529 B.n466 B.n175 10.6151
R2530 B.n470 B.n175 10.6151
R2531 B.n471 B.n470 10.6151
R2532 B.n472 B.n471 10.6151
R2533 B.n472 B.n173 10.6151
R2534 B.n476 B.n173 10.6151
R2535 B.n477 B.n476 10.6151
R2536 B.n478 B.n477 10.6151
R2537 B.n478 B.n171 10.6151
R2538 B.n482 B.n171 10.6151
R2539 B.n483 B.n482 10.6151
R2540 B.n484 B.n483 10.6151
R2541 B.n484 B.n169 10.6151
R2542 B.n488 B.n169 10.6151
R2543 B.n489 B.n488 10.6151
R2544 B.n490 B.n489 10.6151
R2545 B.n490 B.n167 10.6151
R2546 B.n494 B.n167 10.6151
R2547 B.n495 B.n494 10.6151
R2548 B.n496 B.n495 10.6151
R2549 B.n496 B.n165 10.6151
R2550 B.n500 B.n165 10.6151
R2551 B.n501 B.n500 10.6151
R2552 B.n502 B.n501 10.6151
R2553 B.n502 B.n163 10.6151
R2554 B.n506 B.n163 10.6151
R2555 B.n507 B.n506 10.6151
R2556 B.n508 B.n507 10.6151
R2557 B.n508 B.n161 10.6151
R2558 B.n350 B.n219 10.6151
R2559 B.n346 B.n219 10.6151
R2560 B.n346 B.n345 10.6151
R2561 B.n345 B.n344 10.6151
R2562 B.n344 B.n221 10.6151
R2563 B.n340 B.n221 10.6151
R2564 B.n340 B.n339 10.6151
R2565 B.n339 B.n338 10.6151
R2566 B.n338 B.n223 10.6151
R2567 B.n334 B.n223 10.6151
R2568 B.n334 B.n333 10.6151
R2569 B.n333 B.n332 10.6151
R2570 B.n332 B.n225 10.6151
R2571 B.n328 B.n225 10.6151
R2572 B.n328 B.n327 10.6151
R2573 B.n327 B.n326 10.6151
R2574 B.n326 B.n227 10.6151
R2575 B.n322 B.n227 10.6151
R2576 B.n322 B.n321 10.6151
R2577 B.n321 B.n320 10.6151
R2578 B.n320 B.n229 10.6151
R2579 B.n316 B.n229 10.6151
R2580 B.n316 B.n315 10.6151
R2581 B.n315 B.n314 10.6151
R2582 B.n314 B.n231 10.6151
R2583 B.n310 B.n231 10.6151
R2584 B.n310 B.n309 10.6151
R2585 B.n309 B.n308 10.6151
R2586 B.n308 B.n233 10.6151
R2587 B.n304 B.n233 10.6151
R2588 B.n304 B.n303 10.6151
R2589 B.n303 B.n302 10.6151
R2590 B.n302 B.n235 10.6151
R2591 B.n298 B.n235 10.6151
R2592 B.n298 B.n297 10.6151
R2593 B.n297 B.n296 10.6151
R2594 B.n296 B.n237 10.6151
R2595 B.n292 B.n237 10.6151
R2596 B.n292 B.n291 10.6151
R2597 B.n291 B.n290 10.6151
R2598 B.n290 B.n239 10.6151
R2599 B.n286 B.n239 10.6151
R2600 B.n286 B.n285 10.6151
R2601 B.n285 B.n284 10.6151
R2602 B.n284 B.n241 10.6151
R2603 B.n280 B.n241 10.6151
R2604 B.n280 B.n279 10.6151
R2605 B.n279 B.n278 10.6151
R2606 B.n278 B.n243 10.6151
R2607 B.n274 B.n243 10.6151
R2608 B.n274 B.n273 10.6151
R2609 B.n273 B.n272 10.6151
R2610 B.n272 B.n245 10.6151
R2611 B.n268 B.n245 10.6151
R2612 B.n268 B.n267 10.6151
R2613 B.n267 B.n266 10.6151
R2614 B.n266 B.n247 10.6151
R2615 B.n262 B.n247 10.6151
R2616 B.n262 B.n261 10.6151
R2617 B.n261 B.n260 10.6151
R2618 B.n260 B.n249 10.6151
R2619 B.n256 B.n249 10.6151
R2620 B.n256 B.n255 10.6151
R2621 B.n255 B.n254 10.6151
R2622 B.n254 B.n251 10.6151
R2623 B.n251 B.n0 10.6151
R2624 B.n971 B.n1 10.6151
R2625 B.n971 B.n970 10.6151
R2626 B.n970 B.n969 10.6151
R2627 B.n969 B.n4 10.6151
R2628 B.n965 B.n4 10.6151
R2629 B.n965 B.n964 10.6151
R2630 B.n964 B.n963 10.6151
R2631 B.n963 B.n6 10.6151
R2632 B.n959 B.n6 10.6151
R2633 B.n959 B.n958 10.6151
R2634 B.n958 B.n957 10.6151
R2635 B.n957 B.n8 10.6151
R2636 B.n953 B.n8 10.6151
R2637 B.n953 B.n952 10.6151
R2638 B.n952 B.n951 10.6151
R2639 B.n951 B.n10 10.6151
R2640 B.n947 B.n10 10.6151
R2641 B.n947 B.n946 10.6151
R2642 B.n946 B.n945 10.6151
R2643 B.n945 B.n12 10.6151
R2644 B.n941 B.n12 10.6151
R2645 B.n941 B.n940 10.6151
R2646 B.n940 B.n939 10.6151
R2647 B.n939 B.n14 10.6151
R2648 B.n935 B.n14 10.6151
R2649 B.n935 B.n934 10.6151
R2650 B.n934 B.n933 10.6151
R2651 B.n933 B.n16 10.6151
R2652 B.n929 B.n16 10.6151
R2653 B.n929 B.n928 10.6151
R2654 B.n928 B.n927 10.6151
R2655 B.n927 B.n18 10.6151
R2656 B.n923 B.n18 10.6151
R2657 B.n923 B.n922 10.6151
R2658 B.n922 B.n921 10.6151
R2659 B.n921 B.n20 10.6151
R2660 B.n917 B.n20 10.6151
R2661 B.n917 B.n916 10.6151
R2662 B.n916 B.n915 10.6151
R2663 B.n915 B.n22 10.6151
R2664 B.n911 B.n22 10.6151
R2665 B.n911 B.n910 10.6151
R2666 B.n910 B.n909 10.6151
R2667 B.n909 B.n24 10.6151
R2668 B.n905 B.n24 10.6151
R2669 B.n905 B.n904 10.6151
R2670 B.n904 B.n903 10.6151
R2671 B.n903 B.n26 10.6151
R2672 B.n899 B.n26 10.6151
R2673 B.n899 B.n898 10.6151
R2674 B.n898 B.n897 10.6151
R2675 B.n897 B.n28 10.6151
R2676 B.n893 B.n28 10.6151
R2677 B.n893 B.n892 10.6151
R2678 B.n892 B.n891 10.6151
R2679 B.n891 B.n30 10.6151
R2680 B.n887 B.n30 10.6151
R2681 B.n887 B.n886 10.6151
R2682 B.n886 B.n885 10.6151
R2683 B.n885 B.n32 10.6151
R2684 B.n881 B.n32 10.6151
R2685 B.n881 B.n880 10.6151
R2686 B.n880 B.n879 10.6151
R2687 B.n879 B.n34 10.6151
R2688 B.n875 B.n34 10.6151
R2689 B.n875 B.n874 10.6151
R2690 B.n802 B.n801 9.36635
R2691 B.n784 B.n70 9.36635
R2692 B.n423 B.n422 9.36635
R2693 B.n440 B.n187 9.36635
R2694 B.n975 B.n0 2.81026
R2695 B.n975 B.n1 2.81026
R2696 B.n801 B.n800 1.24928
R2697 B.n70 B.n66 1.24928
R2698 B.n424 B.n423 1.24928
R2699 B.n437 B.n187 1.24928
C0 VDD1 VDD2 2.32923f
C1 B VTAIL 6.17292f
C2 VTAIL w_n4970_n3802# 4.77086f
C3 VDD1 VN 0.153204f
C4 B VP 2.59233f
C5 VP w_n4970_n3802# 11.1208f
C6 VDD2 VN 10.803599f
C7 VDD1 VTAIL 9.1378f
C8 VDD2 VTAIL 9.199389f
C9 B w_n4970_n3802# 12.3615f
C10 VDD1 VP 11.2815f
C11 VN VTAIL 11.4489f
C12 VDD2 VP 0.633072f
C13 VP VN 9.37811f
C14 VDD1 B 2.03462f
C15 VDD1 w_n4970_n3802# 2.34918f
C16 VDD2 B 2.16431f
C17 VDD2 w_n4970_n3802# 2.50877f
C18 VP VTAIL 11.463f
C19 B VN 1.49975f
C20 VN w_n4970_n3802# 10.4725f
C21 VDD2 VSUBS 2.519171f
C22 VDD1 VSUBS 3.34203f
C23 VTAIL VSUBS 1.626927f
C24 VN VSUBS 8.254451f
C25 VP VSUBS 4.77802f
C26 B VSUBS 6.380239f
C27 w_n4970_n3802# VSUBS 0.23194p
C28 B.n0 VSUBS 0.005141f
C29 B.n1 VSUBS 0.005141f
C30 B.n2 VSUBS 0.00813f
C31 B.n3 VSUBS 0.00813f
C32 B.n4 VSUBS 0.00813f
C33 B.n5 VSUBS 0.00813f
C34 B.n6 VSUBS 0.00813f
C35 B.n7 VSUBS 0.00813f
C36 B.n8 VSUBS 0.00813f
C37 B.n9 VSUBS 0.00813f
C38 B.n10 VSUBS 0.00813f
C39 B.n11 VSUBS 0.00813f
C40 B.n12 VSUBS 0.00813f
C41 B.n13 VSUBS 0.00813f
C42 B.n14 VSUBS 0.00813f
C43 B.n15 VSUBS 0.00813f
C44 B.n16 VSUBS 0.00813f
C45 B.n17 VSUBS 0.00813f
C46 B.n18 VSUBS 0.00813f
C47 B.n19 VSUBS 0.00813f
C48 B.n20 VSUBS 0.00813f
C49 B.n21 VSUBS 0.00813f
C50 B.n22 VSUBS 0.00813f
C51 B.n23 VSUBS 0.00813f
C52 B.n24 VSUBS 0.00813f
C53 B.n25 VSUBS 0.00813f
C54 B.n26 VSUBS 0.00813f
C55 B.n27 VSUBS 0.00813f
C56 B.n28 VSUBS 0.00813f
C57 B.n29 VSUBS 0.00813f
C58 B.n30 VSUBS 0.00813f
C59 B.n31 VSUBS 0.00813f
C60 B.n32 VSUBS 0.00813f
C61 B.n33 VSUBS 0.00813f
C62 B.n34 VSUBS 0.00813f
C63 B.n35 VSUBS 0.017178f
C64 B.n36 VSUBS 0.00813f
C65 B.n37 VSUBS 0.00813f
C66 B.n38 VSUBS 0.00813f
C67 B.n39 VSUBS 0.00813f
C68 B.n40 VSUBS 0.00813f
C69 B.n41 VSUBS 0.00813f
C70 B.n42 VSUBS 0.00813f
C71 B.n43 VSUBS 0.00813f
C72 B.n44 VSUBS 0.00813f
C73 B.n45 VSUBS 0.00813f
C74 B.n46 VSUBS 0.00813f
C75 B.n47 VSUBS 0.00813f
C76 B.n48 VSUBS 0.00813f
C77 B.n49 VSUBS 0.00813f
C78 B.n50 VSUBS 0.00813f
C79 B.n51 VSUBS 0.00813f
C80 B.n52 VSUBS 0.00813f
C81 B.n53 VSUBS 0.00813f
C82 B.n54 VSUBS 0.00813f
C83 B.n55 VSUBS 0.00813f
C84 B.n56 VSUBS 0.00813f
C85 B.n57 VSUBS 0.00813f
C86 B.n58 VSUBS 0.00813f
C87 B.n59 VSUBS 0.00813f
C88 B.t11 VSUBS 0.302418f
C89 B.t10 VSUBS 0.352804f
C90 B.t9 VSUBS 2.78538f
C91 B.n60 VSUBS 0.561639f
C92 B.n61 VSUBS 0.331393f
C93 B.n62 VSUBS 0.00813f
C94 B.n63 VSUBS 0.00813f
C95 B.n64 VSUBS 0.00813f
C96 B.n65 VSUBS 0.00813f
C97 B.n66 VSUBS 0.004543f
C98 B.n67 VSUBS 0.00813f
C99 B.t8 VSUBS 0.302422f
C100 B.t7 VSUBS 0.352807f
C101 B.t6 VSUBS 2.78538f
C102 B.n68 VSUBS 0.561635f
C103 B.n69 VSUBS 0.331389f
C104 B.n70 VSUBS 0.018835f
C105 B.n71 VSUBS 0.00813f
C106 B.n72 VSUBS 0.00813f
C107 B.n73 VSUBS 0.00813f
C108 B.n74 VSUBS 0.00813f
C109 B.n75 VSUBS 0.00813f
C110 B.n76 VSUBS 0.00813f
C111 B.n77 VSUBS 0.00813f
C112 B.n78 VSUBS 0.00813f
C113 B.n79 VSUBS 0.00813f
C114 B.n80 VSUBS 0.00813f
C115 B.n81 VSUBS 0.00813f
C116 B.n82 VSUBS 0.00813f
C117 B.n83 VSUBS 0.00813f
C118 B.n84 VSUBS 0.00813f
C119 B.n85 VSUBS 0.00813f
C120 B.n86 VSUBS 0.00813f
C121 B.n87 VSUBS 0.00813f
C122 B.n88 VSUBS 0.00813f
C123 B.n89 VSUBS 0.00813f
C124 B.n90 VSUBS 0.00813f
C125 B.n91 VSUBS 0.00813f
C126 B.n92 VSUBS 0.00813f
C127 B.n93 VSUBS 0.017385f
C128 B.n94 VSUBS 0.00813f
C129 B.n95 VSUBS 0.00813f
C130 B.n96 VSUBS 0.00813f
C131 B.n97 VSUBS 0.00813f
C132 B.n98 VSUBS 0.00813f
C133 B.n99 VSUBS 0.00813f
C134 B.n100 VSUBS 0.00813f
C135 B.n101 VSUBS 0.00813f
C136 B.n102 VSUBS 0.00813f
C137 B.n103 VSUBS 0.00813f
C138 B.n104 VSUBS 0.00813f
C139 B.n105 VSUBS 0.00813f
C140 B.n106 VSUBS 0.00813f
C141 B.n107 VSUBS 0.00813f
C142 B.n108 VSUBS 0.00813f
C143 B.n109 VSUBS 0.00813f
C144 B.n110 VSUBS 0.00813f
C145 B.n111 VSUBS 0.00813f
C146 B.n112 VSUBS 0.00813f
C147 B.n113 VSUBS 0.00813f
C148 B.n114 VSUBS 0.00813f
C149 B.n115 VSUBS 0.00813f
C150 B.n116 VSUBS 0.00813f
C151 B.n117 VSUBS 0.00813f
C152 B.n118 VSUBS 0.00813f
C153 B.n119 VSUBS 0.00813f
C154 B.n120 VSUBS 0.00813f
C155 B.n121 VSUBS 0.00813f
C156 B.n122 VSUBS 0.00813f
C157 B.n123 VSUBS 0.00813f
C158 B.n124 VSUBS 0.00813f
C159 B.n125 VSUBS 0.00813f
C160 B.n126 VSUBS 0.00813f
C161 B.n127 VSUBS 0.00813f
C162 B.n128 VSUBS 0.00813f
C163 B.n129 VSUBS 0.00813f
C164 B.n130 VSUBS 0.00813f
C165 B.n131 VSUBS 0.00813f
C166 B.n132 VSUBS 0.00813f
C167 B.n133 VSUBS 0.00813f
C168 B.n134 VSUBS 0.00813f
C169 B.n135 VSUBS 0.00813f
C170 B.n136 VSUBS 0.00813f
C171 B.n137 VSUBS 0.00813f
C172 B.n138 VSUBS 0.00813f
C173 B.n139 VSUBS 0.00813f
C174 B.n140 VSUBS 0.00813f
C175 B.n141 VSUBS 0.00813f
C176 B.n142 VSUBS 0.00813f
C177 B.n143 VSUBS 0.00813f
C178 B.n144 VSUBS 0.00813f
C179 B.n145 VSUBS 0.00813f
C180 B.n146 VSUBS 0.00813f
C181 B.n147 VSUBS 0.00813f
C182 B.n148 VSUBS 0.00813f
C183 B.n149 VSUBS 0.00813f
C184 B.n150 VSUBS 0.00813f
C185 B.n151 VSUBS 0.00813f
C186 B.n152 VSUBS 0.00813f
C187 B.n153 VSUBS 0.00813f
C188 B.n154 VSUBS 0.00813f
C189 B.n155 VSUBS 0.00813f
C190 B.n156 VSUBS 0.00813f
C191 B.n157 VSUBS 0.00813f
C192 B.n158 VSUBS 0.00813f
C193 B.n159 VSUBS 0.00813f
C194 B.n160 VSUBS 0.00813f
C195 B.n161 VSUBS 0.018449f
C196 B.n162 VSUBS 0.00813f
C197 B.n163 VSUBS 0.00813f
C198 B.n164 VSUBS 0.00813f
C199 B.n165 VSUBS 0.00813f
C200 B.n166 VSUBS 0.00813f
C201 B.n167 VSUBS 0.00813f
C202 B.n168 VSUBS 0.00813f
C203 B.n169 VSUBS 0.00813f
C204 B.n170 VSUBS 0.00813f
C205 B.n171 VSUBS 0.00813f
C206 B.n172 VSUBS 0.00813f
C207 B.n173 VSUBS 0.00813f
C208 B.n174 VSUBS 0.00813f
C209 B.n175 VSUBS 0.00813f
C210 B.n176 VSUBS 0.00813f
C211 B.n177 VSUBS 0.00813f
C212 B.n178 VSUBS 0.00813f
C213 B.n179 VSUBS 0.00813f
C214 B.n180 VSUBS 0.00813f
C215 B.n181 VSUBS 0.00813f
C216 B.n182 VSUBS 0.00813f
C217 B.n183 VSUBS 0.00813f
C218 B.n184 VSUBS 0.00813f
C219 B.t4 VSUBS 0.302422f
C220 B.t5 VSUBS 0.352807f
C221 B.t3 VSUBS 2.78538f
C222 B.n185 VSUBS 0.561635f
C223 B.n186 VSUBS 0.331389f
C224 B.n187 VSUBS 0.018835f
C225 B.n188 VSUBS 0.00813f
C226 B.n189 VSUBS 0.00813f
C227 B.n190 VSUBS 0.00813f
C228 B.n191 VSUBS 0.00813f
C229 B.n192 VSUBS 0.00813f
C230 B.t1 VSUBS 0.302418f
C231 B.t2 VSUBS 0.352804f
C232 B.t0 VSUBS 2.78538f
C233 B.n193 VSUBS 0.561639f
C234 B.n194 VSUBS 0.331393f
C235 B.n195 VSUBS 0.00813f
C236 B.n196 VSUBS 0.00813f
C237 B.n197 VSUBS 0.00813f
C238 B.n198 VSUBS 0.00813f
C239 B.n199 VSUBS 0.00813f
C240 B.n200 VSUBS 0.00813f
C241 B.n201 VSUBS 0.00813f
C242 B.n202 VSUBS 0.00813f
C243 B.n203 VSUBS 0.00813f
C244 B.n204 VSUBS 0.00813f
C245 B.n205 VSUBS 0.00813f
C246 B.n206 VSUBS 0.00813f
C247 B.n207 VSUBS 0.00813f
C248 B.n208 VSUBS 0.00813f
C249 B.n209 VSUBS 0.00813f
C250 B.n210 VSUBS 0.00813f
C251 B.n211 VSUBS 0.00813f
C252 B.n212 VSUBS 0.00813f
C253 B.n213 VSUBS 0.00813f
C254 B.n214 VSUBS 0.00813f
C255 B.n215 VSUBS 0.00813f
C256 B.n216 VSUBS 0.00813f
C257 B.n217 VSUBS 0.00813f
C258 B.n218 VSUBS 0.018449f
C259 B.n219 VSUBS 0.00813f
C260 B.n220 VSUBS 0.00813f
C261 B.n221 VSUBS 0.00813f
C262 B.n222 VSUBS 0.00813f
C263 B.n223 VSUBS 0.00813f
C264 B.n224 VSUBS 0.00813f
C265 B.n225 VSUBS 0.00813f
C266 B.n226 VSUBS 0.00813f
C267 B.n227 VSUBS 0.00813f
C268 B.n228 VSUBS 0.00813f
C269 B.n229 VSUBS 0.00813f
C270 B.n230 VSUBS 0.00813f
C271 B.n231 VSUBS 0.00813f
C272 B.n232 VSUBS 0.00813f
C273 B.n233 VSUBS 0.00813f
C274 B.n234 VSUBS 0.00813f
C275 B.n235 VSUBS 0.00813f
C276 B.n236 VSUBS 0.00813f
C277 B.n237 VSUBS 0.00813f
C278 B.n238 VSUBS 0.00813f
C279 B.n239 VSUBS 0.00813f
C280 B.n240 VSUBS 0.00813f
C281 B.n241 VSUBS 0.00813f
C282 B.n242 VSUBS 0.00813f
C283 B.n243 VSUBS 0.00813f
C284 B.n244 VSUBS 0.00813f
C285 B.n245 VSUBS 0.00813f
C286 B.n246 VSUBS 0.00813f
C287 B.n247 VSUBS 0.00813f
C288 B.n248 VSUBS 0.00813f
C289 B.n249 VSUBS 0.00813f
C290 B.n250 VSUBS 0.00813f
C291 B.n251 VSUBS 0.00813f
C292 B.n252 VSUBS 0.00813f
C293 B.n253 VSUBS 0.00813f
C294 B.n254 VSUBS 0.00813f
C295 B.n255 VSUBS 0.00813f
C296 B.n256 VSUBS 0.00813f
C297 B.n257 VSUBS 0.00813f
C298 B.n258 VSUBS 0.00813f
C299 B.n259 VSUBS 0.00813f
C300 B.n260 VSUBS 0.00813f
C301 B.n261 VSUBS 0.00813f
C302 B.n262 VSUBS 0.00813f
C303 B.n263 VSUBS 0.00813f
C304 B.n264 VSUBS 0.00813f
C305 B.n265 VSUBS 0.00813f
C306 B.n266 VSUBS 0.00813f
C307 B.n267 VSUBS 0.00813f
C308 B.n268 VSUBS 0.00813f
C309 B.n269 VSUBS 0.00813f
C310 B.n270 VSUBS 0.00813f
C311 B.n271 VSUBS 0.00813f
C312 B.n272 VSUBS 0.00813f
C313 B.n273 VSUBS 0.00813f
C314 B.n274 VSUBS 0.00813f
C315 B.n275 VSUBS 0.00813f
C316 B.n276 VSUBS 0.00813f
C317 B.n277 VSUBS 0.00813f
C318 B.n278 VSUBS 0.00813f
C319 B.n279 VSUBS 0.00813f
C320 B.n280 VSUBS 0.00813f
C321 B.n281 VSUBS 0.00813f
C322 B.n282 VSUBS 0.00813f
C323 B.n283 VSUBS 0.00813f
C324 B.n284 VSUBS 0.00813f
C325 B.n285 VSUBS 0.00813f
C326 B.n286 VSUBS 0.00813f
C327 B.n287 VSUBS 0.00813f
C328 B.n288 VSUBS 0.00813f
C329 B.n289 VSUBS 0.00813f
C330 B.n290 VSUBS 0.00813f
C331 B.n291 VSUBS 0.00813f
C332 B.n292 VSUBS 0.00813f
C333 B.n293 VSUBS 0.00813f
C334 B.n294 VSUBS 0.00813f
C335 B.n295 VSUBS 0.00813f
C336 B.n296 VSUBS 0.00813f
C337 B.n297 VSUBS 0.00813f
C338 B.n298 VSUBS 0.00813f
C339 B.n299 VSUBS 0.00813f
C340 B.n300 VSUBS 0.00813f
C341 B.n301 VSUBS 0.00813f
C342 B.n302 VSUBS 0.00813f
C343 B.n303 VSUBS 0.00813f
C344 B.n304 VSUBS 0.00813f
C345 B.n305 VSUBS 0.00813f
C346 B.n306 VSUBS 0.00813f
C347 B.n307 VSUBS 0.00813f
C348 B.n308 VSUBS 0.00813f
C349 B.n309 VSUBS 0.00813f
C350 B.n310 VSUBS 0.00813f
C351 B.n311 VSUBS 0.00813f
C352 B.n312 VSUBS 0.00813f
C353 B.n313 VSUBS 0.00813f
C354 B.n314 VSUBS 0.00813f
C355 B.n315 VSUBS 0.00813f
C356 B.n316 VSUBS 0.00813f
C357 B.n317 VSUBS 0.00813f
C358 B.n318 VSUBS 0.00813f
C359 B.n319 VSUBS 0.00813f
C360 B.n320 VSUBS 0.00813f
C361 B.n321 VSUBS 0.00813f
C362 B.n322 VSUBS 0.00813f
C363 B.n323 VSUBS 0.00813f
C364 B.n324 VSUBS 0.00813f
C365 B.n325 VSUBS 0.00813f
C366 B.n326 VSUBS 0.00813f
C367 B.n327 VSUBS 0.00813f
C368 B.n328 VSUBS 0.00813f
C369 B.n329 VSUBS 0.00813f
C370 B.n330 VSUBS 0.00813f
C371 B.n331 VSUBS 0.00813f
C372 B.n332 VSUBS 0.00813f
C373 B.n333 VSUBS 0.00813f
C374 B.n334 VSUBS 0.00813f
C375 B.n335 VSUBS 0.00813f
C376 B.n336 VSUBS 0.00813f
C377 B.n337 VSUBS 0.00813f
C378 B.n338 VSUBS 0.00813f
C379 B.n339 VSUBS 0.00813f
C380 B.n340 VSUBS 0.00813f
C381 B.n341 VSUBS 0.00813f
C382 B.n342 VSUBS 0.00813f
C383 B.n343 VSUBS 0.00813f
C384 B.n344 VSUBS 0.00813f
C385 B.n345 VSUBS 0.00813f
C386 B.n346 VSUBS 0.00813f
C387 B.n347 VSUBS 0.00813f
C388 B.n348 VSUBS 0.00813f
C389 B.n349 VSUBS 0.017178f
C390 B.n350 VSUBS 0.017178f
C391 B.n351 VSUBS 0.018449f
C392 B.n352 VSUBS 0.00813f
C393 B.n353 VSUBS 0.00813f
C394 B.n354 VSUBS 0.00813f
C395 B.n355 VSUBS 0.00813f
C396 B.n356 VSUBS 0.00813f
C397 B.n357 VSUBS 0.00813f
C398 B.n358 VSUBS 0.00813f
C399 B.n359 VSUBS 0.00813f
C400 B.n360 VSUBS 0.00813f
C401 B.n361 VSUBS 0.00813f
C402 B.n362 VSUBS 0.00813f
C403 B.n363 VSUBS 0.00813f
C404 B.n364 VSUBS 0.00813f
C405 B.n365 VSUBS 0.00813f
C406 B.n366 VSUBS 0.00813f
C407 B.n367 VSUBS 0.00813f
C408 B.n368 VSUBS 0.00813f
C409 B.n369 VSUBS 0.00813f
C410 B.n370 VSUBS 0.00813f
C411 B.n371 VSUBS 0.00813f
C412 B.n372 VSUBS 0.00813f
C413 B.n373 VSUBS 0.00813f
C414 B.n374 VSUBS 0.00813f
C415 B.n375 VSUBS 0.00813f
C416 B.n376 VSUBS 0.00813f
C417 B.n377 VSUBS 0.00813f
C418 B.n378 VSUBS 0.00813f
C419 B.n379 VSUBS 0.00813f
C420 B.n380 VSUBS 0.00813f
C421 B.n381 VSUBS 0.00813f
C422 B.n382 VSUBS 0.00813f
C423 B.n383 VSUBS 0.00813f
C424 B.n384 VSUBS 0.00813f
C425 B.n385 VSUBS 0.00813f
C426 B.n386 VSUBS 0.00813f
C427 B.n387 VSUBS 0.00813f
C428 B.n388 VSUBS 0.00813f
C429 B.n389 VSUBS 0.00813f
C430 B.n390 VSUBS 0.00813f
C431 B.n391 VSUBS 0.00813f
C432 B.n392 VSUBS 0.00813f
C433 B.n393 VSUBS 0.00813f
C434 B.n394 VSUBS 0.00813f
C435 B.n395 VSUBS 0.00813f
C436 B.n396 VSUBS 0.00813f
C437 B.n397 VSUBS 0.00813f
C438 B.n398 VSUBS 0.00813f
C439 B.n399 VSUBS 0.00813f
C440 B.n400 VSUBS 0.00813f
C441 B.n401 VSUBS 0.00813f
C442 B.n402 VSUBS 0.00813f
C443 B.n403 VSUBS 0.00813f
C444 B.n404 VSUBS 0.00813f
C445 B.n405 VSUBS 0.00813f
C446 B.n406 VSUBS 0.00813f
C447 B.n407 VSUBS 0.00813f
C448 B.n408 VSUBS 0.00813f
C449 B.n409 VSUBS 0.00813f
C450 B.n410 VSUBS 0.00813f
C451 B.n411 VSUBS 0.00813f
C452 B.n412 VSUBS 0.00813f
C453 B.n413 VSUBS 0.00813f
C454 B.n414 VSUBS 0.00813f
C455 B.n415 VSUBS 0.00813f
C456 B.n416 VSUBS 0.00813f
C457 B.n417 VSUBS 0.00813f
C458 B.n418 VSUBS 0.00813f
C459 B.n419 VSUBS 0.00813f
C460 B.n420 VSUBS 0.00813f
C461 B.n421 VSUBS 0.00813f
C462 B.n422 VSUBS 0.007651f
C463 B.n423 VSUBS 0.018835f
C464 B.n424 VSUBS 0.004543f
C465 B.n425 VSUBS 0.00813f
C466 B.n426 VSUBS 0.00813f
C467 B.n427 VSUBS 0.00813f
C468 B.n428 VSUBS 0.00813f
C469 B.n429 VSUBS 0.00813f
C470 B.n430 VSUBS 0.00813f
C471 B.n431 VSUBS 0.00813f
C472 B.n432 VSUBS 0.00813f
C473 B.n433 VSUBS 0.00813f
C474 B.n434 VSUBS 0.00813f
C475 B.n435 VSUBS 0.00813f
C476 B.n436 VSUBS 0.00813f
C477 B.n437 VSUBS 0.004543f
C478 B.n438 VSUBS 0.00813f
C479 B.n439 VSUBS 0.00813f
C480 B.n440 VSUBS 0.007651f
C481 B.n441 VSUBS 0.00813f
C482 B.n442 VSUBS 0.00813f
C483 B.n443 VSUBS 0.00813f
C484 B.n444 VSUBS 0.00813f
C485 B.n445 VSUBS 0.00813f
C486 B.n446 VSUBS 0.00813f
C487 B.n447 VSUBS 0.00813f
C488 B.n448 VSUBS 0.00813f
C489 B.n449 VSUBS 0.00813f
C490 B.n450 VSUBS 0.00813f
C491 B.n451 VSUBS 0.00813f
C492 B.n452 VSUBS 0.00813f
C493 B.n453 VSUBS 0.00813f
C494 B.n454 VSUBS 0.00813f
C495 B.n455 VSUBS 0.00813f
C496 B.n456 VSUBS 0.00813f
C497 B.n457 VSUBS 0.00813f
C498 B.n458 VSUBS 0.00813f
C499 B.n459 VSUBS 0.00813f
C500 B.n460 VSUBS 0.00813f
C501 B.n461 VSUBS 0.00813f
C502 B.n462 VSUBS 0.00813f
C503 B.n463 VSUBS 0.00813f
C504 B.n464 VSUBS 0.00813f
C505 B.n465 VSUBS 0.00813f
C506 B.n466 VSUBS 0.00813f
C507 B.n467 VSUBS 0.00813f
C508 B.n468 VSUBS 0.00813f
C509 B.n469 VSUBS 0.00813f
C510 B.n470 VSUBS 0.00813f
C511 B.n471 VSUBS 0.00813f
C512 B.n472 VSUBS 0.00813f
C513 B.n473 VSUBS 0.00813f
C514 B.n474 VSUBS 0.00813f
C515 B.n475 VSUBS 0.00813f
C516 B.n476 VSUBS 0.00813f
C517 B.n477 VSUBS 0.00813f
C518 B.n478 VSUBS 0.00813f
C519 B.n479 VSUBS 0.00813f
C520 B.n480 VSUBS 0.00813f
C521 B.n481 VSUBS 0.00813f
C522 B.n482 VSUBS 0.00813f
C523 B.n483 VSUBS 0.00813f
C524 B.n484 VSUBS 0.00813f
C525 B.n485 VSUBS 0.00813f
C526 B.n486 VSUBS 0.00813f
C527 B.n487 VSUBS 0.00813f
C528 B.n488 VSUBS 0.00813f
C529 B.n489 VSUBS 0.00813f
C530 B.n490 VSUBS 0.00813f
C531 B.n491 VSUBS 0.00813f
C532 B.n492 VSUBS 0.00813f
C533 B.n493 VSUBS 0.00813f
C534 B.n494 VSUBS 0.00813f
C535 B.n495 VSUBS 0.00813f
C536 B.n496 VSUBS 0.00813f
C537 B.n497 VSUBS 0.00813f
C538 B.n498 VSUBS 0.00813f
C539 B.n499 VSUBS 0.00813f
C540 B.n500 VSUBS 0.00813f
C541 B.n501 VSUBS 0.00813f
C542 B.n502 VSUBS 0.00813f
C543 B.n503 VSUBS 0.00813f
C544 B.n504 VSUBS 0.00813f
C545 B.n505 VSUBS 0.00813f
C546 B.n506 VSUBS 0.00813f
C547 B.n507 VSUBS 0.00813f
C548 B.n508 VSUBS 0.00813f
C549 B.n509 VSUBS 0.00813f
C550 B.n510 VSUBS 0.018449f
C551 B.n511 VSUBS 0.017178f
C552 B.n512 VSUBS 0.017178f
C553 B.n513 VSUBS 0.00813f
C554 B.n514 VSUBS 0.00813f
C555 B.n515 VSUBS 0.00813f
C556 B.n516 VSUBS 0.00813f
C557 B.n517 VSUBS 0.00813f
C558 B.n518 VSUBS 0.00813f
C559 B.n519 VSUBS 0.00813f
C560 B.n520 VSUBS 0.00813f
C561 B.n521 VSUBS 0.00813f
C562 B.n522 VSUBS 0.00813f
C563 B.n523 VSUBS 0.00813f
C564 B.n524 VSUBS 0.00813f
C565 B.n525 VSUBS 0.00813f
C566 B.n526 VSUBS 0.00813f
C567 B.n527 VSUBS 0.00813f
C568 B.n528 VSUBS 0.00813f
C569 B.n529 VSUBS 0.00813f
C570 B.n530 VSUBS 0.00813f
C571 B.n531 VSUBS 0.00813f
C572 B.n532 VSUBS 0.00813f
C573 B.n533 VSUBS 0.00813f
C574 B.n534 VSUBS 0.00813f
C575 B.n535 VSUBS 0.00813f
C576 B.n536 VSUBS 0.00813f
C577 B.n537 VSUBS 0.00813f
C578 B.n538 VSUBS 0.00813f
C579 B.n539 VSUBS 0.00813f
C580 B.n540 VSUBS 0.00813f
C581 B.n541 VSUBS 0.00813f
C582 B.n542 VSUBS 0.00813f
C583 B.n543 VSUBS 0.00813f
C584 B.n544 VSUBS 0.00813f
C585 B.n545 VSUBS 0.00813f
C586 B.n546 VSUBS 0.00813f
C587 B.n547 VSUBS 0.00813f
C588 B.n548 VSUBS 0.00813f
C589 B.n549 VSUBS 0.00813f
C590 B.n550 VSUBS 0.00813f
C591 B.n551 VSUBS 0.00813f
C592 B.n552 VSUBS 0.00813f
C593 B.n553 VSUBS 0.00813f
C594 B.n554 VSUBS 0.00813f
C595 B.n555 VSUBS 0.00813f
C596 B.n556 VSUBS 0.00813f
C597 B.n557 VSUBS 0.00813f
C598 B.n558 VSUBS 0.00813f
C599 B.n559 VSUBS 0.00813f
C600 B.n560 VSUBS 0.00813f
C601 B.n561 VSUBS 0.00813f
C602 B.n562 VSUBS 0.00813f
C603 B.n563 VSUBS 0.00813f
C604 B.n564 VSUBS 0.00813f
C605 B.n565 VSUBS 0.00813f
C606 B.n566 VSUBS 0.00813f
C607 B.n567 VSUBS 0.00813f
C608 B.n568 VSUBS 0.00813f
C609 B.n569 VSUBS 0.00813f
C610 B.n570 VSUBS 0.00813f
C611 B.n571 VSUBS 0.00813f
C612 B.n572 VSUBS 0.00813f
C613 B.n573 VSUBS 0.00813f
C614 B.n574 VSUBS 0.00813f
C615 B.n575 VSUBS 0.00813f
C616 B.n576 VSUBS 0.00813f
C617 B.n577 VSUBS 0.00813f
C618 B.n578 VSUBS 0.00813f
C619 B.n579 VSUBS 0.00813f
C620 B.n580 VSUBS 0.00813f
C621 B.n581 VSUBS 0.00813f
C622 B.n582 VSUBS 0.00813f
C623 B.n583 VSUBS 0.00813f
C624 B.n584 VSUBS 0.00813f
C625 B.n585 VSUBS 0.00813f
C626 B.n586 VSUBS 0.00813f
C627 B.n587 VSUBS 0.00813f
C628 B.n588 VSUBS 0.00813f
C629 B.n589 VSUBS 0.00813f
C630 B.n590 VSUBS 0.00813f
C631 B.n591 VSUBS 0.00813f
C632 B.n592 VSUBS 0.00813f
C633 B.n593 VSUBS 0.00813f
C634 B.n594 VSUBS 0.00813f
C635 B.n595 VSUBS 0.00813f
C636 B.n596 VSUBS 0.00813f
C637 B.n597 VSUBS 0.00813f
C638 B.n598 VSUBS 0.00813f
C639 B.n599 VSUBS 0.00813f
C640 B.n600 VSUBS 0.00813f
C641 B.n601 VSUBS 0.00813f
C642 B.n602 VSUBS 0.00813f
C643 B.n603 VSUBS 0.00813f
C644 B.n604 VSUBS 0.00813f
C645 B.n605 VSUBS 0.00813f
C646 B.n606 VSUBS 0.00813f
C647 B.n607 VSUBS 0.00813f
C648 B.n608 VSUBS 0.00813f
C649 B.n609 VSUBS 0.00813f
C650 B.n610 VSUBS 0.00813f
C651 B.n611 VSUBS 0.00813f
C652 B.n612 VSUBS 0.00813f
C653 B.n613 VSUBS 0.00813f
C654 B.n614 VSUBS 0.00813f
C655 B.n615 VSUBS 0.00813f
C656 B.n616 VSUBS 0.00813f
C657 B.n617 VSUBS 0.00813f
C658 B.n618 VSUBS 0.00813f
C659 B.n619 VSUBS 0.00813f
C660 B.n620 VSUBS 0.00813f
C661 B.n621 VSUBS 0.00813f
C662 B.n622 VSUBS 0.00813f
C663 B.n623 VSUBS 0.00813f
C664 B.n624 VSUBS 0.00813f
C665 B.n625 VSUBS 0.00813f
C666 B.n626 VSUBS 0.00813f
C667 B.n627 VSUBS 0.00813f
C668 B.n628 VSUBS 0.00813f
C669 B.n629 VSUBS 0.00813f
C670 B.n630 VSUBS 0.00813f
C671 B.n631 VSUBS 0.00813f
C672 B.n632 VSUBS 0.00813f
C673 B.n633 VSUBS 0.00813f
C674 B.n634 VSUBS 0.00813f
C675 B.n635 VSUBS 0.00813f
C676 B.n636 VSUBS 0.00813f
C677 B.n637 VSUBS 0.00813f
C678 B.n638 VSUBS 0.00813f
C679 B.n639 VSUBS 0.00813f
C680 B.n640 VSUBS 0.00813f
C681 B.n641 VSUBS 0.00813f
C682 B.n642 VSUBS 0.00813f
C683 B.n643 VSUBS 0.00813f
C684 B.n644 VSUBS 0.00813f
C685 B.n645 VSUBS 0.00813f
C686 B.n646 VSUBS 0.00813f
C687 B.n647 VSUBS 0.00813f
C688 B.n648 VSUBS 0.00813f
C689 B.n649 VSUBS 0.00813f
C690 B.n650 VSUBS 0.00813f
C691 B.n651 VSUBS 0.00813f
C692 B.n652 VSUBS 0.00813f
C693 B.n653 VSUBS 0.00813f
C694 B.n654 VSUBS 0.00813f
C695 B.n655 VSUBS 0.00813f
C696 B.n656 VSUBS 0.00813f
C697 B.n657 VSUBS 0.00813f
C698 B.n658 VSUBS 0.00813f
C699 B.n659 VSUBS 0.00813f
C700 B.n660 VSUBS 0.00813f
C701 B.n661 VSUBS 0.00813f
C702 B.n662 VSUBS 0.00813f
C703 B.n663 VSUBS 0.00813f
C704 B.n664 VSUBS 0.00813f
C705 B.n665 VSUBS 0.00813f
C706 B.n666 VSUBS 0.00813f
C707 B.n667 VSUBS 0.00813f
C708 B.n668 VSUBS 0.00813f
C709 B.n669 VSUBS 0.00813f
C710 B.n670 VSUBS 0.00813f
C711 B.n671 VSUBS 0.00813f
C712 B.n672 VSUBS 0.00813f
C713 B.n673 VSUBS 0.00813f
C714 B.n674 VSUBS 0.00813f
C715 B.n675 VSUBS 0.00813f
C716 B.n676 VSUBS 0.00813f
C717 B.n677 VSUBS 0.00813f
C718 B.n678 VSUBS 0.00813f
C719 B.n679 VSUBS 0.00813f
C720 B.n680 VSUBS 0.00813f
C721 B.n681 VSUBS 0.00813f
C722 B.n682 VSUBS 0.00813f
C723 B.n683 VSUBS 0.00813f
C724 B.n684 VSUBS 0.00813f
C725 B.n685 VSUBS 0.00813f
C726 B.n686 VSUBS 0.00813f
C727 B.n687 VSUBS 0.00813f
C728 B.n688 VSUBS 0.00813f
C729 B.n689 VSUBS 0.00813f
C730 B.n690 VSUBS 0.00813f
C731 B.n691 VSUBS 0.00813f
C732 B.n692 VSUBS 0.00813f
C733 B.n693 VSUBS 0.00813f
C734 B.n694 VSUBS 0.00813f
C735 B.n695 VSUBS 0.00813f
C736 B.n696 VSUBS 0.00813f
C737 B.n697 VSUBS 0.00813f
C738 B.n698 VSUBS 0.00813f
C739 B.n699 VSUBS 0.00813f
C740 B.n700 VSUBS 0.00813f
C741 B.n701 VSUBS 0.00813f
C742 B.n702 VSUBS 0.00813f
C743 B.n703 VSUBS 0.00813f
C744 B.n704 VSUBS 0.00813f
C745 B.n705 VSUBS 0.00813f
C746 B.n706 VSUBS 0.00813f
C747 B.n707 VSUBS 0.00813f
C748 B.n708 VSUBS 0.00813f
C749 B.n709 VSUBS 0.00813f
C750 B.n710 VSUBS 0.00813f
C751 B.n711 VSUBS 0.00813f
C752 B.n712 VSUBS 0.018241f
C753 B.n713 VSUBS 0.017178f
C754 B.n714 VSUBS 0.018449f
C755 B.n715 VSUBS 0.00813f
C756 B.n716 VSUBS 0.00813f
C757 B.n717 VSUBS 0.00813f
C758 B.n718 VSUBS 0.00813f
C759 B.n719 VSUBS 0.00813f
C760 B.n720 VSUBS 0.00813f
C761 B.n721 VSUBS 0.00813f
C762 B.n722 VSUBS 0.00813f
C763 B.n723 VSUBS 0.00813f
C764 B.n724 VSUBS 0.00813f
C765 B.n725 VSUBS 0.00813f
C766 B.n726 VSUBS 0.00813f
C767 B.n727 VSUBS 0.00813f
C768 B.n728 VSUBS 0.00813f
C769 B.n729 VSUBS 0.00813f
C770 B.n730 VSUBS 0.00813f
C771 B.n731 VSUBS 0.00813f
C772 B.n732 VSUBS 0.00813f
C773 B.n733 VSUBS 0.00813f
C774 B.n734 VSUBS 0.00813f
C775 B.n735 VSUBS 0.00813f
C776 B.n736 VSUBS 0.00813f
C777 B.n737 VSUBS 0.00813f
C778 B.n738 VSUBS 0.00813f
C779 B.n739 VSUBS 0.00813f
C780 B.n740 VSUBS 0.00813f
C781 B.n741 VSUBS 0.00813f
C782 B.n742 VSUBS 0.00813f
C783 B.n743 VSUBS 0.00813f
C784 B.n744 VSUBS 0.00813f
C785 B.n745 VSUBS 0.00813f
C786 B.n746 VSUBS 0.00813f
C787 B.n747 VSUBS 0.00813f
C788 B.n748 VSUBS 0.00813f
C789 B.n749 VSUBS 0.00813f
C790 B.n750 VSUBS 0.00813f
C791 B.n751 VSUBS 0.00813f
C792 B.n752 VSUBS 0.00813f
C793 B.n753 VSUBS 0.00813f
C794 B.n754 VSUBS 0.00813f
C795 B.n755 VSUBS 0.00813f
C796 B.n756 VSUBS 0.00813f
C797 B.n757 VSUBS 0.00813f
C798 B.n758 VSUBS 0.00813f
C799 B.n759 VSUBS 0.00813f
C800 B.n760 VSUBS 0.00813f
C801 B.n761 VSUBS 0.00813f
C802 B.n762 VSUBS 0.00813f
C803 B.n763 VSUBS 0.00813f
C804 B.n764 VSUBS 0.00813f
C805 B.n765 VSUBS 0.00813f
C806 B.n766 VSUBS 0.00813f
C807 B.n767 VSUBS 0.00813f
C808 B.n768 VSUBS 0.00813f
C809 B.n769 VSUBS 0.00813f
C810 B.n770 VSUBS 0.00813f
C811 B.n771 VSUBS 0.00813f
C812 B.n772 VSUBS 0.00813f
C813 B.n773 VSUBS 0.00813f
C814 B.n774 VSUBS 0.00813f
C815 B.n775 VSUBS 0.00813f
C816 B.n776 VSUBS 0.00813f
C817 B.n777 VSUBS 0.00813f
C818 B.n778 VSUBS 0.00813f
C819 B.n779 VSUBS 0.00813f
C820 B.n780 VSUBS 0.00813f
C821 B.n781 VSUBS 0.00813f
C822 B.n782 VSUBS 0.00813f
C823 B.n783 VSUBS 0.00813f
C824 B.n784 VSUBS 0.007651f
C825 B.n785 VSUBS 0.00813f
C826 B.n786 VSUBS 0.00813f
C827 B.n787 VSUBS 0.00813f
C828 B.n788 VSUBS 0.00813f
C829 B.n789 VSUBS 0.00813f
C830 B.n790 VSUBS 0.00813f
C831 B.n791 VSUBS 0.00813f
C832 B.n792 VSUBS 0.00813f
C833 B.n793 VSUBS 0.00813f
C834 B.n794 VSUBS 0.00813f
C835 B.n795 VSUBS 0.00813f
C836 B.n796 VSUBS 0.00813f
C837 B.n797 VSUBS 0.00813f
C838 B.n798 VSUBS 0.00813f
C839 B.n799 VSUBS 0.00813f
C840 B.n800 VSUBS 0.004543f
C841 B.n801 VSUBS 0.018835f
C842 B.n802 VSUBS 0.007651f
C843 B.n803 VSUBS 0.00813f
C844 B.n804 VSUBS 0.00813f
C845 B.n805 VSUBS 0.00813f
C846 B.n806 VSUBS 0.00813f
C847 B.n807 VSUBS 0.00813f
C848 B.n808 VSUBS 0.00813f
C849 B.n809 VSUBS 0.00813f
C850 B.n810 VSUBS 0.00813f
C851 B.n811 VSUBS 0.00813f
C852 B.n812 VSUBS 0.00813f
C853 B.n813 VSUBS 0.00813f
C854 B.n814 VSUBS 0.00813f
C855 B.n815 VSUBS 0.00813f
C856 B.n816 VSUBS 0.00813f
C857 B.n817 VSUBS 0.00813f
C858 B.n818 VSUBS 0.00813f
C859 B.n819 VSUBS 0.00813f
C860 B.n820 VSUBS 0.00813f
C861 B.n821 VSUBS 0.00813f
C862 B.n822 VSUBS 0.00813f
C863 B.n823 VSUBS 0.00813f
C864 B.n824 VSUBS 0.00813f
C865 B.n825 VSUBS 0.00813f
C866 B.n826 VSUBS 0.00813f
C867 B.n827 VSUBS 0.00813f
C868 B.n828 VSUBS 0.00813f
C869 B.n829 VSUBS 0.00813f
C870 B.n830 VSUBS 0.00813f
C871 B.n831 VSUBS 0.00813f
C872 B.n832 VSUBS 0.00813f
C873 B.n833 VSUBS 0.00813f
C874 B.n834 VSUBS 0.00813f
C875 B.n835 VSUBS 0.00813f
C876 B.n836 VSUBS 0.00813f
C877 B.n837 VSUBS 0.00813f
C878 B.n838 VSUBS 0.00813f
C879 B.n839 VSUBS 0.00813f
C880 B.n840 VSUBS 0.00813f
C881 B.n841 VSUBS 0.00813f
C882 B.n842 VSUBS 0.00813f
C883 B.n843 VSUBS 0.00813f
C884 B.n844 VSUBS 0.00813f
C885 B.n845 VSUBS 0.00813f
C886 B.n846 VSUBS 0.00813f
C887 B.n847 VSUBS 0.00813f
C888 B.n848 VSUBS 0.00813f
C889 B.n849 VSUBS 0.00813f
C890 B.n850 VSUBS 0.00813f
C891 B.n851 VSUBS 0.00813f
C892 B.n852 VSUBS 0.00813f
C893 B.n853 VSUBS 0.00813f
C894 B.n854 VSUBS 0.00813f
C895 B.n855 VSUBS 0.00813f
C896 B.n856 VSUBS 0.00813f
C897 B.n857 VSUBS 0.00813f
C898 B.n858 VSUBS 0.00813f
C899 B.n859 VSUBS 0.00813f
C900 B.n860 VSUBS 0.00813f
C901 B.n861 VSUBS 0.00813f
C902 B.n862 VSUBS 0.00813f
C903 B.n863 VSUBS 0.00813f
C904 B.n864 VSUBS 0.00813f
C905 B.n865 VSUBS 0.00813f
C906 B.n866 VSUBS 0.00813f
C907 B.n867 VSUBS 0.00813f
C908 B.n868 VSUBS 0.00813f
C909 B.n869 VSUBS 0.00813f
C910 B.n870 VSUBS 0.00813f
C911 B.n871 VSUBS 0.00813f
C912 B.n872 VSUBS 0.018449f
C913 B.n873 VSUBS 0.018449f
C914 B.n874 VSUBS 0.017178f
C915 B.n875 VSUBS 0.00813f
C916 B.n876 VSUBS 0.00813f
C917 B.n877 VSUBS 0.00813f
C918 B.n878 VSUBS 0.00813f
C919 B.n879 VSUBS 0.00813f
C920 B.n880 VSUBS 0.00813f
C921 B.n881 VSUBS 0.00813f
C922 B.n882 VSUBS 0.00813f
C923 B.n883 VSUBS 0.00813f
C924 B.n884 VSUBS 0.00813f
C925 B.n885 VSUBS 0.00813f
C926 B.n886 VSUBS 0.00813f
C927 B.n887 VSUBS 0.00813f
C928 B.n888 VSUBS 0.00813f
C929 B.n889 VSUBS 0.00813f
C930 B.n890 VSUBS 0.00813f
C931 B.n891 VSUBS 0.00813f
C932 B.n892 VSUBS 0.00813f
C933 B.n893 VSUBS 0.00813f
C934 B.n894 VSUBS 0.00813f
C935 B.n895 VSUBS 0.00813f
C936 B.n896 VSUBS 0.00813f
C937 B.n897 VSUBS 0.00813f
C938 B.n898 VSUBS 0.00813f
C939 B.n899 VSUBS 0.00813f
C940 B.n900 VSUBS 0.00813f
C941 B.n901 VSUBS 0.00813f
C942 B.n902 VSUBS 0.00813f
C943 B.n903 VSUBS 0.00813f
C944 B.n904 VSUBS 0.00813f
C945 B.n905 VSUBS 0.00813f
C946 B.n906 VSUBS 0.00813f
C947 B.n907 VSUBS 0.00813f
C948 B.n908 VSUBS 0.00813f
C949 B.n909 VSUBS 0.00813f
C950 B.n910 VSUBS 0.00813f
C951 B.n911 VSUBS 0.00813f
C952 B.n912 VSUBS 0.00813f
C953 B.n913 VSUBS 0.00813f
C954 B.n914 VSUBS 0.00813f
C955 B.n915 VSUBS 0.00813f
C956 B.n916 VSUBS 0.00813f
C957 B.n917 VSUBS 0.00813f
C958 B.n918 VSUBS 0.00813f
C959 B.n919 VSUBS 0.00813f
C960 B.n920 VSUBS 0.00813f
C961 B.n921 VSUBS 0.00813f
C962 B.n922 VSUBS 0.00813f
C963 B.n923 VSUBS 0.00813f
C964 B.n924 VSUBS 0.00813f
C965 B.n925 VSUBS 0.00813f
C966 B.n926 VSUBS 0.00813f
C967 B.n927 VSUBS 0.00813f
C968 B.n928 VSUBS 0.00813f
C969 B.n929 VSUBS 0.00813f
C970 B.n930 VSUBS 0.00813f
C971 B.n931 VSUBS 0.00813f
C972 B.n932 VSUBS 0.00813f
C973 B.n933 VSUBS 0.00813f
C974 B.n934 VSUBS 0.00813f
C975 B.n935 VSUBS 0.00813f
C976 B.n936 VSUBS 0.00813f
C977 B.n937 VSUBS 0.00813f
C978 B.n938 VSUBS 0.00813f
C979 B.n939 VSUBS 0.00813f
C980 B.n940 VSUBS 0.00813f
C981 B.n941 VSUBS 0.00813f
C982 B.n942 VSUBS 0.00813f
C983 B.n943 VSUBS 0.00813f
C984 B.n944 VSUBS 0.00813f
C985 B.n945 VSUBS 0.00813f
C986 B.n946 VSUBS 0.00813f
C987 B.n947 VSUBS 0.00813f
C988 B.n948 VSUBS 0.00813f
C989 B.n949 VSUBS 0.00813f
C990 B.n950 VSUBS 0.00813f
C991 B.n951 VSUBS 0.00813f
C992 B.n952 VSUBS 0.00813f
C993 B.n953 VSUBS 0.00813f
C994 B.n954 VSUBS 0.00813f
C995 B.n955 VSUBS 0.00813f
C996 B.n956 VSUBS 0.00813f
C997 B.n957 VSUBS 0.00813f
C998 B.n958 VSUBS 0.00813f
C999 B.n959 VSUBS 0.00813f
C1000 B.n960 VSUBS 0.00813f
C1001 B.n961 VSUBS 0.00813f
C1002 B.n962 VSUBS 0.00813f
C1003 B.n963 VSUBS 0.00813f
C1004 B.n964 VSUBS 0.00813f
C1005 B.n965 VSUBS 0.00813f
C1006 B.n966 VSUBS 0.00813f
C1007 B.n967 VSUBS 0.00813f
C1008 B.n968 VSUBS 0.00813f
C1009 B.n969 VSUBS 0.00813f
C1010 B.n970 VSUBS 0.00813f
C1011 B.n971 VSUBS 0.00813f
C1012 B.n972 VSUBS 0.00813f
C1013 B.n973 VSUBS 0.00813f
C1014 B.n974 VSUBS 0.00813f
C1015 B.n975 VSUBS 0.018408f
C1016 VDD1.t6 VSUBS 0.362069f
C1017 VDD1.t1 VSUBS 0.362069f
C1018 VDD1.n0 VSUBS 2.91896f
C1019 VDD1.t2 VSUBS 0.362069f
C1020 VDD1.t4 VSUBS 0.362069f
C1021 VDD1.n1 VSUBS 2.91682f
C1022 VDD1.t5 VSUBS 0.362069f
C1023 VDD1.t0 VSUBS 0.362069f
C1024 VDD1.n2 VSUBS 2.91682f
C1025 VDD1.n3 VSUBS 6.01494f
C1026 VDD1.t7 VSUBS 0.362069f
C1027 VDD1.t3 VSUBS 0.362069f
C1028 VDD1.n4 VSUBS 2.88905f
C1029 VDD1.n5 VSUBS 4.92112f
C1030 VP.n0 VSUBS 0.047132f
C1031 VP.t7 VSUBS 3.56587f
C1032 VP.n1 VSUBS 0.0498f
C1033 VP.n2 VSUBS 0.025057f
C1034 VP.n3 VSUBS 0.0467f
C1035 VP.n4 VSUBS 0.025057f
C1036 VP.t2 VSUBS 3.56587f
C1037 VP.n5 VSUBS 0.0498f
C1038 VP.n6 VSUBS 0.025057f
C1039 VP.n7 VSUBS 0.0467f
C1040 VP.n8 VSUBS 0.025057f
C1041 VP.t3 VSUBS 3.56587f
C1042 VP.n9 VSUBS 0.0498f
C1043 VP.n10 VSUBS 0.025057f
C1044 VP.n11 VSUBS 0.0467f
C1045 VP.n12 VSUBS 0.047132f
C1046 VP.t4 VSUBS 3.56587f
C1047 VP.n13 VSUBS 0.0498f
C1048 VP.n14 VSUBS 0.025057f
C1049 VP.n15 VSUBS 0.0467f
C1050 VP.n16 VSUBS 0.025057f
C1051 VP.t0 VSUBS 3.56587f
C1052 VP.n17 VSUBS 0.0498f
C1053 VP.n18 VSUBS 0.025057f
C1054 VP.n19 VSUBS 0.0467f
C1055 VP.t1 VSUBS 3.93433f
C1056 VP.t6 VSUBS 3.56587f
C1057 VP.n20 VSUBS 1.34259f
C1058 VP.n21 VSUBS 1.28053f
C1059 VP.n22 VSUBS 0.31931f
C1060 VP.n23 VSUBS 0.025057f
C1061 VP.n24 VSUBS 0.0467f
C1062 VP.n25 VSUBS 0.0498f
C1063 VP.n26 VSUBS 0.020256f
C1064 VP.n27 VSUBS 0.025057f
C1065 VP.n28 VSUBS 0.025057f
C1066 VP.n29 VSUBS 0.025057f
C1067 VP.n30 VSUBS 0.0467f
C1068 VP.n31 VSUBS 0.0467f
C1069 VP.n32 VSUBS 1.26396f
C1070 VP.n33 VSUBS 0.025057f
C1071 VP.n34 VSUBS 0.025057f
C1072 VP.n35 VSUBS 0.025057f
C1073 VP.n36 VSUBS 0.0467f
C1074 VP.n37 VSUBS 0.0498f
C1075 VP.n38 VSUBS 0.020256f
C1076 VP.n39 VSUBS 0.025057f
C1077 VP.n40 VSUBS 0.025057f
C1078 VP.n41 VSUBS 0.025057f
C1079 VP.n42 VSUBS 0.0467f
C1080 VP.n43 VSUBS 0.0467f
C1081 VP.n44 VSUBS 1.35134f
C1082 VP.n45 VSUBS 1.76634f
C1083 VP.t5 VSUBS 3.56587f
C1084 VP.n46 VSUBS 1.35134f
C1085 VP.n47 VSUBS 1.78193f
C1086 VP.n48 VSUBS 0.047132f
C1087 VP.n49 VSUBS 0.025057f
C1088 VP.n50 VSUBS 0.0467f
C1089 VP.n51 VSUBS 0.0498f
C1090 VP.n52 VSUBS 0.020256f
C1091 VP.n53 VSUBS 0.025057f
C1092 VP.n54 VSUBS 0.025057f
C1093 VP.n55 VSUBS 0.025057f
C1094 VP.n56 VSUBS 0.0467f
C1095 VP.n57 VSUBS 0.0467f
C1096 VP.n58 VSUBS 1.26396f
C1097 VP.n59 VSUBS 0.025057f
C1098 VP.n60 VSUBS 0.025057f
C1099 VP.n61 VSUBS 0.025057f
C1100 VP.n62 VSUBS 0.0467f
C1101 VP.n63 VSUBS 0.0498f
C1102 VP.n64 VSUBS 0.020256f
C1103 VP.n65 VSUBS 0.025057f
C1104 VP.n66 VSUBS 0.025057f
C1105 VP.n67 VSUBS 0.025057f
C1106 VP.n68 VSUBS 0.0467f
C1107 VP.n69 VSUBS 0.0467f
C1108 VP.n70 VSUBS 1.26396f
C1109 VP.n71 VSUBS 0.025057f
C1110 VP.n72 VSUBS 0.025057f
C1111 VP.n73 VSUBS 0.025057f
C1112 VP.n74 VSUBS 0.0467f
C1113 VP.n75 VSUBS 0.0498f
C1114 VP.n76 VSUBS 0.020256f
C1115 VP.n77 VSUBS 0.025057f
C1116 VP.n78 VSUBS 0.025057f
C1117 VP.n79 VSUBS 0.025057f
C1118 VP.n80 VSUBS 0.0467f
C1119 VP.n81 VSUBS 0.0467f
C1120 VP.n82 VSUBS 1.35134f
C1121 VP.n83 VSUBS 0.070522f
C1122 VTAIL.t8 VSUBS 0.28282f
C1123 VTAIL.t13 VSUBS 0.28282f
C1124 VTAIL.n0 VSUBS 2.10075f
C1125 VTAIL.n1 VSUBS 0.905636f
C1126 VTAIL.n2 VSUBS 0.027754f
C1127 VTAIL.n3 VSUBS 0.025257f
C1128 VTAIL.n4 VSUBS 0.013572f
C1129 VTAIL.n5 VSUBS 0.03208f
C1130 VTAIL.n6 VSUBS 0.01437f
C1131 VTAIL.n7 VSUBS 0.025257f
C1132 VTAIL.n8 VSUBS 0.013572f
C1133 VTAIL.n9 VSUBS 0.03208f
C1134 VTAIL.n10 VSUBS 0.01437f
C1135 VTAIL.n11 VSUBS 0.025257f
C1136 VTAIL.n12 VSUBS 0.013572f
C1137 VTAIL.n13 VSUBS 0.03208f
C1138 VTAIL.n14 VSUBS 0.01437f
C1139 VTAIL.n15 VSUBS 0.025257f
C1140 VTAIL.n16 VSUBS 0.013971f
C1141 VTAIL.n17 VSUBS 0.03208f
C1142 VTAIL.n18 VSUBS 0.01437f
C1143 VTAIL.n19 VSUBS 0.025257f
C1144 VTAIL.n20 VSUBS 0.013572f
C1145 VTAIL.n21 VSUBS 0.03208f
C1146 VTAIL.n22 VSUBS 0.01437f
C1147 VTAIL.n23 VSUBS 0.025257f
C1148 VTAIL.n24 VSUBS 0.013572f
C1149 VTAIL.n25 VSUBS 0.02406f
C1150 VTAIL.n26 VSUBS 0.024132f
C1151 VTAIL.t10 VSUBS 0.06931f
C1152 VTAIL.n27 VSUBS 0.223695f
C1153 VTAIL.n28 VSUBS 1.48113f
C1154 VTAIL.n29 VSUBS 0.013572f
C1155 VTAIL.n30 VSUBS 0.01437f
C1156 VTAIL.n31 VSUBS 0.03208f
C1157 VTAIL.n32 VSUBS 0.03208f
C1158 VTAIL.n33 VSUBS 0.01437f
C1159 VTAIL.n34 VSUBS 0.013572f
C1160 VTAIL.n35 VSUBS 0.025257f
C1161 VTAIL.n36 VSUBS 0.025257f
C1162 VTAIL.n37 VSUBS 0.013572f
C1163 VTAIL.n38 VSUBS 0.01437f
C1164 VTAIL.n39 VSUBS 0.03208f
C1165 VTAIL.n40 VSUBS 0.03208f
C1166 VTAIL.n41 VSUBS 0.01437f
C1167 VTAIL.n42 VSUBS 0.013572f
C1168 VTAIL.n43 VSUBS 0.025257f
C1169 VTAIL.n44 VSUBS 0.025257f
C1170 VTAIL.n45 VSUBS 0.013572f
C1171 VTAIL.n46 VSUBS 0.013572f
C1172 VTAIL.n47 VSUBS 0.01437f
C1173 VTAIL.n48 VSUBS 0.03208f
C1174 VTAIL.n49 VSUBS 0.03208f
C1175 VTAIL.n50 VSUBS 0.03208f
C1176 VTAIL.n51 VSUBS 0.013971f
C1177 VTAIL.n52 VSUBS 0.013572f
C1178 VTAIL.n53 VSUBS 0.025257f
C1179 VTAIL.n54 VSUBS 0.025257f
C1180 VTAIL.n55 VSUBS 0.013572f
C1181 VTAIL.n56 VSUBS 0.01437f
C1182 VTAIL.n57 VSUBS 0.03208f
C1183 VTAIL.n58 VSUBS 0.03208f
C1184 VTAIL.n59 VSUBS 0.01437f
C1185 VTAIL.n60 VSUBS 0.013572f
C1186 VTAIL.n61 VSUBS 0.025257f
C1187 VTAIL.n62 VSUBS 0.025257f
C1188 VTAIL.n63 VSUBS 0.013572f
C1189 VTAIL.n64 VSUBS 0.01437f
C1190 VTAIL.n65 VSUBS 0.03208f
C1191 VTAIL.n66 VSUBS 0.03208f
C1192 VTAIL.n67 VSUBS 0.01437f
C1193 VTAIL.n68 VSUBS 0.013572f
C1194 VTAIL.n69 VSUBS 0.025257f
C1195 VTAIL.n70 VSUBS 0.025257f
C1196 VTAIL.n71 VSUBS 0.013572f
C1197 VTAIL.n72 VSUBS 0.01437f
C1198 VTAIL.n73 VSUBS 0.03208f
C1199 VTAIL.n74 VSUBS 0.077666f
C1200 VTAIL.n75 VSUBS 0.01437f
C1201 VTAIL.n76 VSUBS 0.013572f
C1202 VTAIL.n77 VSUBS 0.054586f
C1203 VTAIL.n78 VSUBS 0.038937f
C1204 VTAIL.n79 VSUBS 0.338306f
C1205 VTAIL.n80 VSUBS 0.027754f
C1206 VTAIL.n81 VSUBS 0.025257f
C1207 VTAIL.n82 VSUBS 0.013572f
C1208 VTAIL.n83 VSUBS 0.03208f
C1209 VTAIL.n84 VSUBS 0.01437f
C1210 VTAIL.n85 VSUBS 0.025257f
C1211 VTAIL.n86 VSUBS 0.013572f
C1212 VTAIL.n87 VSUBS 0.03208f
C1213 VTAIL.n88 VSUBS 0.01437f
C1214 VTAIL.n89 VSUBS 0.025257f
C1215 VTAIL.n90 VSUBS 0.013572f
C1216 VTAIL.n91 VSUBS 0.03208f
C1217 VTAIL.n92 VSUBS 0.01437f
C1218 VTAIL.n93 VSUBS 0.025257f
C1219 VTAIL.n94 VSUBS 0.013971f
C1220 VTAIL.n95 VSUBS 0.03208f
C1221 VTAIL.n96 VSUBS 0.01437f
C1222 VTAIL.n97 VSUBS 0.025257f
C1223 VTAIL.n98 VSUBS 0.013572f
C1224 VTAIL.n99 VSUBS 0.03208f
C1225 VTAIL.n100 VSUBS 0.01437f
C1226 VTAIL.n101 VSUBS 0.025257f
C1227 VTAIL.n102 VSUBS 0.013572f
C1228 VTAIL.n103 VSUBS 0.02406f
C1229 VTAIL.n104 VSUBS 0.024132f
C1230 VTAIL.t7 VSUBS 0.06931f
C1231 VTAIL.n105 VSUBS 0.223695f
C1232 VTAIL.n106 VSUBS 1.48113f
C1233 VTAIL.n107 VSUBS 0.013572f
C1234 VTAIL.n108 VSUBS 0.01437f
C1235 VTAIL.n109 VSUBS 0.03208f
C1236 VTAIL.n110 VSUBS 0.03208f
C1237 VTAIL.n111 VSUBS 0.01437f
C1238 VTAIL.n112 VSUBS 0.013572f
C1239 VTAIL.n113 VSUBS 0.025257f
C1240 VTAIL.n114 VSUBS 0.025257f
C1241 VTAIL.n115 VSUBS 0.013572f
C1242 VTAIL.n116 VSUBS 0.01437f
C1243 VTAIL.n117 VSUBS 0.03208f
C1244 VTAIL.n118 VSUBS 0.03208f
C1245 VTAIL.n119 VSUBS 0.01437f
C1246 VTAIL.n120 VSUBS 0.013572f
C1247 VTAIL.n121 VSUBS 0.025257f
C1248 VTAIL.n122 VSUBS 0.025257f
C1249 VTAIL.n123 VSUBS 0.013572f
C1250 VTAIL.n124 VSUBS 0.013572f
C1251 VTAIL.n125 VSUBS 0.01437f
C1252 VTAIL.n126 VSUBS 0.03208f
C1253 VTAIL.n127 VSUBS 0.03208f
C1254 VTAIL.n128 VSUBS 0.03208f
C1255 VTAIL.n129 VSUBS 0.013971f
C1256 VTAIL.n130 VSUBS 0.013572f
C1257 VTAIL.n131 VSUBS 0.025257f
C1258 VTAIL.n132 VSUBS 0.025257f
C1259 VTAIL.n133 VSUBS 0.013572f
C1260 VTAIL.n134 VSUBS 0.01437f
C1261 VTAIL.n135 VSUBS 0.03208f
C1262 VTAIL.n136 VSUBS 0.03208f
C1263 VTAIL.n137 VSUBS 0.01437f
C1264 VTAIL.n138 VSUBS 0.013572f
C1265 VTAIL.n139 VSUBS 0.025257f
C1266 VTAIL.n140 VSUBS 0.025257f
C1267 VTAIL.n141 VSUBS 0.013572f
C1268 VTAIL.n142 VSUBS 0.01437f
C1269 VTAIL.n143 VSUBS 0.03208f
C1270 VTAIL.n144 VSUBS 0.03208f
C1271 VTAIL.n145 VSUBS 0.01437f
C1272 VTAIL.n146 VSUBS 0.013572f
C1273 VTAIL.n147 VSUBS 0.025257f
C1274 VTAIL.n148 VSUBS 0.025257f
C1275 VTAIL.n149 VSUBS 0.013572f
C1276 VTAIL.n150 VSUBS 0.01437f
C1277 VTAIL.n151 VSUBS 0.03208f
C1278 VTAIL.n152 VSUBS 0.077666f
C1279 VTAIL.n153 VSUBS 0.01437f
C1280 VTAIL.n154 VSUBS 0.013572f
C1281 VTAIL.n155 VSUBS 0.054586f
C1282 VTAIL.n156 VSUBS 0.038937f
C1283 VTAIL.n157 VSUBS 0.338306f
C1284 VTAIL.t0 VSUBS 0.28282f
C1285 VTAIL.t5 VSUBS 0.28282f
C1286 VTAIL.n158 VSUBS 2.10075f
C1287 VTAIL.n159 VSUBS 1.18154f
C1288 VTAIL.n160 VSUBS 0.027754f
C1289 VTAIL.n161 VSUBS 0.025257f
C1290 VTAIL.n162 VSUBS 0.013572f
C1291 VTAIL.n163 VSUBS 0.03208f
C1292 VTAIL.n164 VSUBS 0.01437f
C1293 VTAIL.n165 VSUBS 0.025257f
C1294 VTAIL.n166 VSUBS 0.013572f
C1295 VTAIL.n167 VSUBS 0.03208f
C1296 VTAIL.n168 VSUBS 0.01437f
C1297 VTAIL.n169 VSUBS 0.025257f
C1298 VTAIL.n170 VSUBS 0.013572f
C1299 VTAIL.n171 VSUBS 0.03208f
C1300 VTAIL.n172 VSUBS 0.01437f
C1301 VTAIL.n173 VSUBS 0.025257f
C1302 VTAIL.n174 VSUBS 0.013971f
C1303 VTAIL.n175 VSUBS 0.03208f
C1304 VTAIL.n176 VSUBS 0.01437f
C1305 VTAIL.n177 VSUBS 0.025257f
C1306 VTAIL.n178 VSUBS 0.013572f
C1307 VTAIL.n179 VSUBS 0.03208f
C1308 VTAIL.n180 VSUBS 0.01437f
C1309 VTAIL.n181 VSUBS 0.025257f
C1310 VTAIL.n182 VSUBS 0.013572f
C1311 VTAIL.n183 VSUBS 0.02406f
C1312 VTAIL.n184 VSUBS 0.024132f
C1313 VTAIL.t2 VSUBS 0.06931f
C1314 VTAIL.n185 VSUBS 0.223695f
C1315 VTAIL.n186 VSUBS 1.48113f
C1316 VTAIL.n187 VSUBS 0.013572f
C1317 VTAIL.n188 VSUBS 0.01437f
C1318 VTAIL.n189 VSUBS 0.03208f
C1319 VTAIL.n190 VSUBS 0.03208f
C1320 VTAIL.n191 VSUBS 0.01437f
C1321 VTAIL.n192 VSUBS 0.013572f
C1322 VTAIL.n193 VSUBS 0.025257f
C1323 VTAIL.n194 VSUBS 0.025257f
C1324 VTAIL.n195 VSUBS 0.013572f
C1325 VTAIL.n196 VSUBS 0.01437f
C1326 VTAIL.n197 VSUBS 0.03208f
C1327 VTAIL.n198 VSUBS 0.03208f
C1328 VTAIL.n199 VSUBS 0.01437f
C1329 VTAIL.n200 VSUBS 0.013572f
C1330 VTAIL.n201 VSUBS 0.025257f
C1331 VTAIL.n202 VSUBS 0.025257f
C1332 VTAIL.n203 VSUBS 0.013572f
C1333 VTAIL.n204 VSUBS 0.013572f
C1334 VTAIL.n205 VSUBS 0.01437f
C1335 VTAIL.n206 VSUBS 0.03208f
C1336 VTAIL.n207 VSUBS 0.03208f
C1337 VTAIL.n208 VSUBS 0.03208f
C1338 VTAIL.n209 VSUBS 0.013971f
C1339 VTAIL.n210 VSUBS 0.013572f
C1340 VTAIL.n211 VSUBS 0.025257f
C1341 VTAIL.n212 VSUBS 0.025257f
C1342 VTAIL.n213 VSUBS 0.013572f
C1343 VTAIL.n214 VSUBS 0.01437f
C1344 VTAIL.n215 VSUBS 0.03208f
C1345 VTAIL.n216 VSUBS 0.03208f
C1346 VTAIL.n217 VSUBS 0.01437f
C1347 VTAIL.n218 VSUBS 0.013572f
C1348 VTAIL.n219 VSUBS 0.025257f
C1349 VTAIL.n220 VSUBS 0.025257f
C1350 VTAIL.n221 VSUBS 0.013572f
C1351 VTAIL.n222 VSUBS 0.01437f
C1352 VTAIL.n223 VSUBS 0.03208f
C1353 VTAIL.n224 VSUBS 0.03208f
C1354 VTAIL.n225 VSUBS 0.01437f
C1355 VTAIL.n226 VSUBS 0.013572f
C1356 VTAIL.n227 VSUBS 0.025257f
C1357 VTAIL.n228 VSUBS 0.025257f
C1358 VTAIL.n229 VSUBS 0.013572f
C1359 VTAIL.n230 VSUBS 0.01437f
C1360 VTAIL.n231 VSUBS 0.03208f
C1361 VTAIL.n232 VSUBS 0.077666f
C1362 VTAIL.n233 VSUBS 0.01437f
C1363 VTAIL.n234 VSUBS 0.013572f
C1364 VTAIL.n235 VSUBS 0.054586f
C1365 VTAIL.n236 VSUBS 0.038937f
C1366 VTAIL.n237 VSUBS 1.91795f
C1367 VTAIL.n238 VSUBS 0.027754f
C1368 VTAIL.n239 VSUBS 0.025257f
C1369 VTAIL.n240 VSUBS 0.013572f
C1370 VTAIL.n241 VSUBS 0.03208f
C1371 VTAIL.n242 VSUBS 0.01437f
C1372 VTAIL.n243 VSUBS 0.025257f
C1373 VTAIL.n244 VSUBS 0.013572f
C1374 VTAIL.n245 VSUBS 0.03208f
C1375 VTAIL.n246 VSUBS 0.01437f
C1376 VTAIL.n247 VSUBS 0.025257f
C1377 VTAIL.n248 VSUBS 0.013572f
C1378 VTAIL.n249 VSUBS 0.03208f
C1379 VTAIL.n250 VSUBS 0.01437f
C1380 VTAIL.n251 VSUBS 0.025257f
C1381 VTAIL.n252 VSUBS 0.013971f
C1382 VTAIL.n253 VSUBS 0.03208f
C1383 VTAIL.n254 VSUBS 0.013572f
C1384 VTAIL.n255 VSUBS 0.01437f
C1385 VTAIL.n256 VSUBS 0.025257f
C1386 VTAIL.n257 VSUBS 0.013572f
C1387 VTAIL.n258 VSUBS 0.03208f
C1388 VTAIL.n259 VSUBS 0.01437f
C1389 VTAIL.n260 VSUBS 0.025257f
C1390 VTAIL.n261 VSUBS 0.013572f
C1391 VTAIL.n262 VSUBS 0.02406f
C1392 VTAIL.n263 VSUBS 0.024132f
C1393 VTAIL.t14 VSUBS 0.06931f
C1394 VTAIL.n264 VSUBS 0.223695f
C1395 VTAIL.n265 VSUBS 1.48113f
C1396 VTAIL.n266 VSUBS 0.013572f
C1397 VTAIL.n267 VSUBS 0.01437f
C1398 VTAIL.n268 VSUBS 0.03208f
C1399 VTAIL.n269 VSUBS 0.03208f
C1400 VTAIL.n270 VSUBS 0.01437f
C1401 VTAIL.n271 VSUBS 0.013572f
C1402 VTAIL.n272 VSUBS 0.025257f
C1403 VTAIL.n273 VSUBS 0.025257f
C1404 VTAIL.n274 VSUBS 0.013572f
C1405 VTAIL.n275 VSUBS 0.01437f
C1406 VTAIL.n276 VSUBS 0.03208f
C1407 VTAIL.n277 VSUBS 0.03208f
C1408 VTAIL.n278 VSUBS 0.01437f
C1409 VTAIL.n279 VSUBS 0.013572f
C1410 VTAIL.n280 VSUBS 0.025257f
C1411 VTAIL.n281 VSUBS 0.025257f
C1412 VTAIL.n282 VSUBS 0.013572f
C1413 VTAIL.n283 VSUBS 0.01437f
C1414 VTAIL.n284 VSUBS 0.03208f
C1415 VTAIL.n285 VSUBS 0.03208f
C1416 VTAIL.n286 VSUBS 0.03208f
C1417 VTAIL.n287 VSUBS 0.013971f
C1418 VTAIL.n288 VSUBS 0.013572f
C1419 VTAIL.n289 VSUBS 0.025257f
C1420 VTAIL.n290 VSUBS 0.025257f
C1421 VTAIL.n291 VSUBS 0.013572f
C1422 VTAIL.n292 VSUBS 0.01437f
C1423 VTAIL.n293 VSUBS 0.03208f
C1424 VTAIL.n294 VSUBS 0.03208f
C1425 VTAIL.n295 VSUBS 0.01437f
C1426 VTAIL.n296 VSUBS 0.013572f
C1427 VTAIL.n297 VSUBS 0.025257f
C1428 VTAIL.n298 VSUBS 0.025257f
C1429 VTAIL.n299 VSUBS 0.013572f
C1430 VTAIL.n300 VSUBS 0.01437f
C1431 VTAIL.n301 VSUBS 0.03208f
C1432 VTAIL.n302 VSUBS 0.03208f
C1433 VTAIL.n303 VSUBS 0.01437f
C1434 VTAIL.n304 VSUBS 0.013572f
C1435 VTAIL.n305 VSUBS 0.025257f
C1436 VTAIL.n306 VSUBS 0.025257f
C1437 VTAIL.n307 VSUBS 0.013572f
C1438 VTAIL.n308 VSUBS 0.01437f
C1439 VTAIL.n309 VSUBS 0.03208f
C1440 VTAIL.n310 VSUBS 0.077666f
C1441 VTAIL.n311 VSUBS 0.01437f
C1442 VTAIL.n312 VSUBS 0.013572f
C1443 VTAIL.n313 VSUBS 0.054586f
C1444 VTAIL.n314 VSUBS 0.038937f
C1445 VTAIL.n315 VSUBS 1.91795f
C1446 VTAIL.t9 VSUBS 0.28282f
C1447 VTAIL.t15 VSUBS 0.28282f
C1448 VTAIL.n316 VSUBS 2.10076f
C1449 VTAIL.n317 VSUBS 1.18153f
C1450 VTAIL.n318 VSUBS 0.027754f
C1451 VTAIL.n319 VSUBS 0.025257f
C1452 VTAIL.n320 VSUBS 0.013572f
C1453 VTAIL.n321 VSUBS 0.03208f
C1454 VTAIL.n322 VSUBS 0.01437f
C1455 VTAIL.n323 VSUBS 0.025257f
C1456 VTAIL.n324 VSUBS 0.013572f
C1457 VTAIL.n325 VSUBS 0.03208f
C1458 VTAIL.n326 VSUBS 0.01437f
C1459 VTAIL.n327 VSUBS 0.025257f
C1460 VTAIL.n328 VSUBS 0.013572f
C1461 VTAIL.n329 VSUBS 0.03208f
C1462 VTAIL.n330 VSUBS 0.01437f
C1463 VTAIL.n331 VSUBS 0.025257f
C1464 VTAIL.n332 VSUBS 0.013971f
C1465 VTAIL.n333 VSUBS 0.03208f
C1466 VTAIL.n334 VSUBS 0.013572f
C1467 VTAIL.n335 VSUBS 0.01437f
C1468 VTAIL.n336 VSUBS 0.025257f
C1469 VTAIL.n337 VSUBS 0.013572f
C1470 VTAIL.n338 VSUBS 0.03208f
C1471 VTAIL.n339 VSUBS 0.01437f
C1472 VTAIL.n340 VSUBS 0.025257f
C1473 VTAIL.n341 VSUBS 0.013572f
C1474 VTAIL.n342 VSUBS 0.02406f
C1475 VTAIL.n343 VSUBS 0.024132f
C1476 VTAIL.t11 VSUBS 0.06931f
C1477 VTAIL.n344 VSUBS 0.223695f
C1478 VTAIL.n345 VSUBS 1.48113f
C1479 VTAIL.n346 VSUBS 0.013572f
C1480 VTAIL.n347 VSUBS 0.01437f
C1481 VTAIL.n348 VSUBS 0.03208f
C1482 VTAIL.n349 VSUBS 0.03208f
C1483 VTAIL.n350 VSUBS 0.01437f
C1484 VTAIL.n351 VSUBS 0.013572f
C1485 VTAIL.n352 VSUBS 0.025257f
C1486 VTAIL.n353 VSUBS 0.025257f
C1487 VTAIL.n354 VSUBS 0.013572f
C1488 VTAIL.n355 VSUBS 0.01437f
C1489 VTAIL.n356 VSUBS 0.03208f
C1490 VTAIL.n357 VSUBS 0.03208f
C1491 VTAIL.n358 VSUBS 0.01437f
C1492 VTAIL.n359 VSUBS 0.013572f
C1493 VTAIL.n360 VSUBS 0.025257f
C1494 VTAIL.n361 VSUBS 0.025257f
C1495 VTAIL.n362 VSUBS 0.013572f
C1496 VTAIL.n363 VSUBS 0.01437f
C1497 VTAIL.n364 VSUBS 0.03208f
C1498 VTAIL.n365 VSUBS 0.03208f
C1499 VTAIL.n366 VSUBS 0.03208f
C1500 VTAIL.n367 VSUBS 0.013971f
C1501 VTAIL.n368 VSUBS 0.013572f
C1502 VTAIL.n369 VSUBS 0.025257f
C1503 VTAIL.n370 VSUBS 0.025257f
C1504 VTAIL.n371 VSUBS 0.013572f
C1505 VTAIL.n372 VSUBS 0.01437f
C1506 VTAIL.n373 VSUBS 0.03208f
C1507 VTAIL.n374 VSUBS 0.03208f
C1508 VTAIL.n375 VSUBS 0.01437f
C1509 VTAIL.n376 VSUBS 0.013572f
C1510 VTAIL.n377 VSUBS 0.025257f
C1511 VTAIL.n378 VSUBS 0.025257f
C1512 VTAIL.n379 VSUBS 0.013572f
C1513 VTAIL.n380 VSUBS 0.01437f
C1514 VTAIL.n381 VSUBS 0.03208f
C1515 VTAIL.n382 VSUBS 0.03208f
C1516 VTAIL.n383 VSUBS 0.01437f
C1517 VTAIL.n384 VSUBS 0.013572f
C1518 VTAIL.n385 VSUBS 0.025257f
C1519 VTAIL.n386 VSUBS 0.025257f
C1520 VTAIL.n387 VSUBS 0.013572f
C1521 VTAIL.n388 VSUBS 0.01437f
C1522 VTAIL.n389 VSUBS 0.03208f
C1523 VTAIL.n390 VSUBS 0.077666f
C1524 VTAIL.n391 VSUBS 0.01437f
C1525 VTAIL.n392 VSUBS 0.013572f
C1526 VTAIL.n393 VSUBS 0.054586f
C1527 VTAIL.n394 VSUBS 0.038937f
C1528 VTAIL.n395 VSUBS 0.338306f
C1529 VTAIL.n396 VSUBS 0.027754f
C1530 VTAIL.n397 VSUBS 0.025257f
C1531 VTAIL.n398 VSUBS 0.013572f
C1532 VTAIL.n399 VSUBS 0.03208f
C1533 VTAIL.n400 VSUBS 0.01437f
C1534 VTAIL.n401 VSUBS 0.025257f
C1535 VTAIL.n402 VSUBS 0.013572f
C1536 VTAIL.n403 VSUBS 0.03208f
C1537 VTAIL.n404 VSUBS 0.01437f
C1538 VTAIL.n405 VSUBS 0.025257f
C1539 VTAIL.n406 VSUBS 0.013572f
C1540 VTAIL.n407 VSUBS 0.03208f
C1541 VTAIL.n408 VSUBS 0.01437f
C1542 VTAIL.n409 VSUBS 0.025257f
C1543 VTAIL.n410 VSUBS 0.013971f
C1544 VTAIL.n411 VSUBS 0.03208f
C1545 VTAIL.n412 VSUBS 0.013572f
C1546 VTAIL.n413 VSUBS 0.01437f
C1547 VTAIL.n414 VSUBS 0.025257f
C1548 VTAIL.n415 VSUBS 0.013572f
C1549 VTAIL.n416 VSUBS 0.03208f
C1550 VTAIL.n417 VSUBS 0.01437f
C1551 VTAIL.n418 VSUBS 0.025257f
C1552 VTAIL.n419 VSUBS 0.013572f
C1553 VTAIL.n420 VSUBS 0.02406f
C1554 VTAIL.n421 VSUBS 0.024132f
C1555 VTAIL.t4 VSUBS 0.06931f
C1556 VTAIL.n422 VSUBS 0.223695f
C1557 VTAIL.n423 VSUBS 1.48113f
C1558 VTAIL.n424 VSUBS 0.013572f
C1559 VTAIL.n425 VSUBS 0.01437f
C1560 VTAIL.n426 VSUBS 0.03208f
C1561 VTAIL.n427 VSUBS 0.03208f
C1562 VTAIL.n428 VSUBS 0.01437f
C1563 VTAIL.n429 VSUBS 0.013572f
C1564 VTAIL.n430 VSUBS 0.025257f
C1565 VTAIL.n431 VSUBS 0.025257f
C1566 VTAIL.n432 VSUBS 0.013572f
C1567 VTAIL.n433 VSUBS 0.01437f
C1568 VTAIL.n434 VSUBS 0.03208f
C1569 VTAIL.n435 VSUBS 0.03208f
C1570 VTAIL.n436 VSUBS 0.01437f
C1571 VTAIL.n437 VSUBS 0.013572f
C1572 VTAIL.n438 VSUBS 0.025257f
C1573 VTAIL.n439 VSUBS 0.025257f
C1574 VTAIL.n440 VSUBS 0.013572f
C1575 VTAIL.n441 VSUBS 0.01437f
C1576 VTAIL.n442 VSUBS 0.03208f
C1577 VTAIL.n443 VSUBS 0.03208f
C1578 VTAIL.n444 VSUBS 0.03208f
C1579 VTAIL.n445 VSUBS 0.013971f
C1580 VTAIL.n446 VSUBS 0.013572f
C1581 VTAIL.n447 VSUBS 0.025257f
C1582 VTAIL.n448 VSUBS 0.025257f
C1583 VTAIL.n449 VSUBS 0.013572f
C1584 VTAIL.n450 VSUBS 0.01437f
C1585 VTAIL.n451 VSUBS 0.03208f
C1586 VTAIL.n452 VSUBS 0.03208f
C1587 VTAIL.n453 VSUBS 0.01437f
C1588 VTAIL.n454 VSUBS 0.013572f
C1589 VTAIL.n455 VSUBS 0.025257f
C1590 VTAIL.n456 VSUBS 0.025257f
C1591 VTAIL.n457 VSUBS 0.013572f
C1592 VTAIL.n458 VSUBS 0.01437f
C1593 VTAIL.n459 VSUBS 0.03208f
C1594 VTAIL.n460 VSUBS 0.03208f
C1595 VTAIL.n461 VSUBS 0.01437f
C1596 VTAIL.n462 VSUBS 0.013572f
C1597 VTAIL.n463 VSUBS 0.025257f
C1598 VTAIL.n464 VSUBS 0.025257f
C1599 VTAIL.n465 VSUBS 0.013572f
C1600 VTAIL.n466 VSUBS 0.01437f
C1601 VTAIL.n467 VSUBS 0.03208f
C1602 VTAIL.n468 VSUBS 0.077666f
C1603 VTAIL.n469 VSUBS 0.01437f
C1604 VTAIL.n470 VSUBS 0.013572f
C1605 VTAIL.n471 VSUBS 0.054586f
C1606 VTAIL.n472 VSUBS 0.038937f
C1607 VTAIL.n473 VSUBS 0.338306f
C1608 VTAIL.t6 VSUBS 0.28282f
C1609 VTAIL.t3 VSUBS 0.28282f
C1610 VTAIL.n474 VSUBS 2.10076f
C1611 VTAIL.n475 VSUBS 1.18153f
C1612 VTAIL.n476 VSUBS 0.027754f
C1613 VTAIL.n477 VSUBS 0.025257f
C1614 VTAIL.n478 VSUBS 0.013572f
C1615 VTAIL.n479 VSUBS 0.03208f
C1616 VTAIL.n480 VSUBS 0.01437f
C1617 VTAIL.n481 VSUBS 0.025257f
C1618 VTAIL.n482 VSUBS 0.013572f
C1619 VTAIL.n483 VSUBS 0.03208f
C1620 VTAIL.n484 VSUBS 0.01437f
C1621 VTAIL.n485 VSUBS 0.025257f
C1622 VTAIL.n486 VSUBS 0.013572f
C1623 VTAIL.n487 VSUBS 0.03208f
C1624 VTAIL.n488 VSUBS 0.01437f
C1625 VTAIL.n489 VSUBS 0.025257f
C1626 VTAIL.n490 VSUBS 0.013971f
C1627 VTAIL.n491 VSUBS 0.03208f
C1628 VTAIL.n492 VSUBS 0.013572f
C1629 VTAIL.n493 VSUBS 0.01437f
C1630 VTAIL.n494 VSUBS 0.025257f
C1631 VTAIL.n495 VSUBS 0.013572f
C1632 VTAIL.n496 VSUBS 0.03208f
C1633 VTAIL.n497 VSUBS 0.01437f
C1634 VTAIL.n498 VSUBS 0.025257f
C1635 VTAIL.n499 VSUBS 0.013572f
C1636 VTAIL.n500 VSUBS 0.02406f
C1637 VTAIL.n501 VSUBS 0.024132f
C1638 VTAIL.t1 VSUBS 0.06931f
C1639 VTAIL.n502 VSUBS 0.223695f
C1640 VTAIL.n503 VSUBS 1.48113f
C1641 VTAIL.n504 VSUBS 0.013572f
C1642 VTAIL.n505 VSUBS 0.01437f
C1643 VTAIL.n506 VSUBS 0.03208f
C1644 VTAIL.n507 VSUBS 0.03208f
C1645 VTAIL.n508 VSUBS 0.01437f
C1646 VTAIL.n509 VSUBS 0.013572f
C1647 VTAIL.n510 VSUBS 0.025257f
C1648 VTAIL.n511 VSUBS 0.025257f
C1649 VTAIL.n512 VSUBS 0.013572f
C1650 VTAIL.n513 VSUBS 0.01437f
C1651 VTAIL.n514 VSUBS 0.03208f
C1652 VTAIL.n515 VSUBS 0.03208f
C1653 VTAIL.n516 VSUBS 0.01437f
C1654 VTAIL.n517 VSUBS 0.013572f
C1655 VTAIL.n518 VSUBS 0.025257f
C1656 VTAIL.n519 VSUBS 0.025257f
C1657 VTAIL.n520 VSUBS 0.013572f
C1658 VTAIL.n521 VSUBS 0.01437f
C1659 VTAIL.n522 VSUBS 0.03208f
C1660 VTAIL.n523 VSUBS 0.03208f
C1661 VTAIL.n524 VSUBS 0.03208f
C1662 VTAIL.n525 VSUBS 0.013971f
C1663 VTAIL.n526 VSUBS 0.013572f
C1664 VTAIL.n527 VSUBS 0.025257f
C1665 VTAIL.n528 VSUBS 0.025257f
C1666 VTAIL.n529 VSUBS 0.013572f
C1667 VTAIL.n530 VSUBS 0.01437f
C1668 VTAIL.n531 VSUBS 0.03208f
C1669 VTAIL.n532 VSUBS 0.03208f
C1670 VTAIL.n533 VSUBS 0.01437f
C1671 VTAIL.n534 VSUBS 0.013572f
C1672 VTAIL.n535 VSUBS 0.025257f
C1673 VTAIL.n536 VSUBS 0.025257f
C1674 VTAIL.n537 VSUBS 0.013572f
C1675 VTAIL.n538 VSUBS 0.01437f
C1676 VTAIL.n539 VSUBS 0.03208f
C1677 VTAIL.n540 VSUBS 0.03208f
C1678 VTAIL.n541 VSUBS 0.01437f
C1679 VTAIL.n542 VSUBS 0.013572f
C1680 VTAIL.n543 VSUBS 0.025257f
C1681 VTAIL.n544 VSUBS 0.025257f
C1682 VTAIL.n545 VSUBS 0.013572f
C1683 VTAIL.n546 VSUBS 0.01437f
C1684 VTAIL.n547 VSUBS 0.03208f
C1685 VTAIL.n548 VSUBS 0.077666f
C1686 VTAIL.n549 VSUBS 0.01437f
C1687 VTAIL.n550 VSUBS 0.013572f
C1688 VTAIL.n551 VSUBS 0.054586f
C1689 VTAIL.n552 VSUBS 0.038937f
C1690 VTAIL.n553 VSUBS 1.91795f
C1691 VTAIL.n554 VSUBS 0.027754f
C1692 VTAIL.n555 VSUBS 0.025257f
C1693 VTAIL.n556 VSUBS 0.013572f
C1694 VTAIL.n557 VSUBS 0.03208f
C1695 VTAIL.n558 VSUBS 0.01437f
C1696 VTAIL.n559 VSUBS 0.025257f
C1697 VTAIL.n560 VSUBS 0.013572f
C1698 VTAIL.n561 VSUBS 0.03208f
C1699 VTAIL.n562 VSUBS 0.01437f
C1700 VTAIL.n563 VSUBS 0.025257f
C1701 VTAIL.n564 VSUBS 0.013572f
C1702 VTAIL.n565 VSUBS 0.03208f
C1703 VTAIL.n566 VSUBS 0.01437f
C1704 VTAIL.n567 VSUBS 0.025257f
C1705 VTAIL.n568 VSUBS 0.013971f
C1706 VTAIL.n569 VSUBS 0.03208f
C1707 VTAIL.n570 VSUBS 0.01437f
C1708 VTAIL.n571 VSUBS 0.025257f
C1709 VTAIL.n572 VSUBS 0.013572f
C1710 VTAIL.n573 VSUBS 0.03208f
C1711 VTAIL.n574 VSUBS 0.01437f
C1712 VTAIL.n575 VSUBS 0.025257f
C1713 VTAIL.n576 VSUBS 0.013572f
C1714 VTAIL.n577 VSUBS 0.02406f
C1715 VTAIL.n578 VSUBS 0.024132f
C1716 VTAIL.t12 VSUBS 0.06931f
C1717 VTAIL.n579 VSUBS 0.223695f
C1718 VTAIL.n580 VSUBS 1.48113f
C1719 VTAIL.n581 VSUBS 0.013572f
C1720 VTAIL.n582 VSUBS 0.01437f
C1721 VTAIL.n583 VSUBS 0.03208f
C1722 VTAIL.n584 VSUBS 0.03208f
C1723 VTAIL.n585 VSUBS 0.01437f
C1724 VTAIL.n586 VSUBS 0.013572f
C1725 VTAIL.n587 VSUBS 0.025257f
C1726 VTAIL.n588 VSUBS 0.025257f
C1727 VTAIL.n589 VSUBS 0.013572f
C1728 VTAIL.n590 VSUBS 0.01437f
C1729 VTAIL.n591 VSUBS 0.03208f
C1730 VTAIL.n592 VSUBS 0.03208f
C1731 VTAIL.n593 VSUBS 0.01437f
C1732 VTAIL.n594 VSUBS 0.013572f
C1733 VTAIL.n595 VSUBS 0.025257f
C1734 VTAIL.n596 VSUBS 0.025257f
C1735 VTAIL.n597 VSUBS 0.013572f
C1736 VTAIL.n598 VSUBS 0.013572f
C1737 VTAIL.n599 VSUBS 0.01437f
C1738 VTAIL.n600 VSUBS 0.03208f
C1739 VTAIL.n601 VSUBS 0.03208f
C1740 VTAIL.n602 VSUBS 0.03208f
C1741 VTAIL.n603 VSUBS 0.013971f
C1742 VTAIL.n604 VSUBS 0.013572f
C1743 VTAIL.n605 VSUBS 0.025257f
C1744 VTAIL.n606 VSUBS 0.025257f
C1745 VTAIL.n607 VSUBS 0.013572f
C1746 VTAIL.n608 VSUBS 0.01437f
C1747 VTAIL.n609 VSUBS 0.03208f
C1748 VTAIL.n610 VSUBS 0.03208f
C1749 VTAIL.n611 VSUBS 0.01437f
C1750 VTAIL.n612 VSUBS 0.013572f
C1751 VTAIL.n613 VSUBS 0.025257f
C1752 VTAIL.n614 VSUBS 0.025257f
C1753 VTAIL.n615 VSUBS 0.013572f
C1754 VTAIL.n616 VSUBS 0.01437f
C1755 VTAIL.n617 VSUBS 0.03208f
C1756 VTAIL.n618 VSUBS 0.03208f
C1757 VTAIL.n619 VSUBS 0.01437f
C1758 VTAIL.n620 VSUBS 0.013572f
C1759 VTAIL.n621 VSUBS 0.025257f
C1760 VTAIL.n622 VSUBS 0.025257f
C1761 VTAIL.n623 VSUBS 0.013572f
C1762 VTAIL.n624 VSUBS 0.01437f
C1763 VTAIL.n625 VSUBS 0.03208f
C1764 VTAIL.n626 VSUBS 0.077666f
C1765 VTAIL.n627 VSUBS 0.01437f
C1766 VTAIL.n628 VSUBS 0.013572f
C1767 VTAIL.n629 VSUBS 0.054586f
C1768 VTAIL.n630 VSUBS 0.038937f
C1769 VTAIL.n631 VSUBS 1.91322f
C1770 VDD2.t6 VSUBS 0.363678f
C1771 VDD2.t4 VSUBS 0.363678f
C1772 VDD2.n0 VSUBS 2.92978f
C1773 VDD2.t1 VSUBS 0.363678f
C1774 VDD2.t0 VSUBS 0.363678f
C1775 VDD2.n1 VSUBS 2.92978f
C1776 VDD2.n2 VSUBS 5.97483f
C1777 VDD2.t2 VSUBS 0.363678f
C1778 VDD2.t5 VSUBS 0.363678f
C1779 VDD2.n3 VSUBS 2.90188f
C1780 VDD2.n4 VSUBS 4.90204f
C1781 VDD2.t3 VSUBS 0.363678f
C1782 VDD2.t7 VSUBS 0.363678f
C1783 VDD2.n5 VSUBS 2.92973f
C1784 VN.n0 VSUBS 0.043197f
C1785 VN.t3 VSUBS 3.26815f
C1786 VN.n1 VSUBS 0.045642f
C1787 VN.n2 VSUBS 0.022965f
C1788 VN.n3 VSUBS 0.042801f
C1789 VN.n4 VSUBS 0.022965f
C1790 VN.t2 VSUBS 3.26815f
C1791 VN.n5 VSUBS 0.045642f
C1792 VN.n6 VSUBS 0.022965f
C1793 VN.n7 VSUBS 0.042801f
C1794 VN.t5 VSUBS 3.60585f
C1795 VN.t7 VSUBS 3.26815f
C1796 VN.n8 VSUBS 1.23049f
C1797 VN.n9 VSUBS 1.17361f
C1798 VN.n10 VSUBS 0.29265f
C1799 VN.n11 VSUBS 0.022965f
C1800 VN.n12 VSUBS 0.042801f
C1801 VN.n13 VSUBS 0.045642f
C1802 VN.n14 VSUBS 0.018565f
C1803 VN.n15 VSUBS 0.022965f
C1804 VN.n16 VSUBS 0.022965f
C1805 VN.n17 VSUBS 0.022965f
C1806 VN.n18 VSUBS 0.042801f
C1807 VN.n19 VSUBS 0.042801f
C1808 VN.n20 VSUBS 1.15843f
C1809 VN.n21 VSUBS 0.022965f
C1810 VN.n22 VSUBS 0.022965f
C1811 VN.n23 VSUBS 0.022965f
C1812 VN.n24 VSUBS 0.042801f
C1813 VN.n25 VSUBS 0.045642f
C1814 VN.n26 VSUBS 0.018565f
C1815 VN.n27 VSUBS 0.022965f
C1816 VN.n28 VSUBS 0.022965f
C1817 VN.n29 VSUBS 0.022965f
C1818 VN.n30 VSUBS 0.042801f
C1819 VN.n31 VSUBS 0.042801f
C1820 VN.n32 VSUBS 1.23852f
C1821 VN.n33 VSUBS 0.064634f
C1822 VN.n34 VSUBS 0.043197f
C1823 VN.t1 VSUBS 3.26815f
C1824 VN.n35 VSUBS 0.045642f
C1825 VN.n36 VSUBS 0.022965f
C1826 VN.n37 VSUBS 0.042801f
C1827 VN.n38 VSUBS 0.022965f
C1828 VN.t6 VSUBS 3.26815f
C1829 VN.n39 VSUBS 0.045642f
C1830 VN.n40 VSUBS 0.022965f
C1831 VN.n41 VSUBS 0.042801f
C1832 VN.t4 VSUBS 3.60585f
C1833 VN.t0 VSUBS 3.26815f
C1834 VN.n42 VSUBS 1.23049f
C1835 VN.n43 VSUBS 1.17361f
C1836 VN.n44 VSUBS 0.29265f
C1837 VN.n45 VSUBS 0.022965f
C1838 VN.n46 VSUBS 0.042801f
C1839 VN.n47 VSUBS 0.045642f
C1840 VN.n48 VSUBS 0.018565f
C1841 VN.n49 VSUBS 0.022965f
C1842 VN.n50 VSUBS 0.022965f
C1843 VN.n51 VSUBS 0.022965f
C1844 VN.n52 VSUBS 0.042801f
C1845 VN.n53 VSUBS 0.042801f
C1846 VN.n54 VSUBS 1.15843f
C1847 VN.n55 VSUBS 0.022965f
C1848 VN.n56 VSUBS 0.022965f
C1849 VN.n57 VSUBS 0.022965f
C1850 VN.n58 VSUBS 0.042801f
C1851 VN.n59 VSUBS 0.045642f
C1852 VN.n60 VSUBS 0.018565f
C1853 VN.n61 VSUBS 0.022965f
C1854 VN.n62 VSUBS 0.022965f
C1855 VN.n63 VSUBS 0.022965f
C1856 VN.n64 VSUBS 0.042801f
C1857 VN.n65 VSUBS 0.042801f
C1858 VN.n66 VSUBS 1.23852f
C1859 VN.n67 VSUBS 1.62427f
.ends

