* NGSPICE file created from diff_pair_sample_1766.ext - technology: sky130A

.subckt diff_pair_sample_1766 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=4.5903 pd=24.32 as=1.94205 ps=12.1 w=11.77 l=3.45
X1 VTAIL.t8 VN.t0 VDD2.t9 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X2 VTAIL.t17 VP.t1 VDD1.t8 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X3 VDD2.t8 VN.t1 VTAIL.t2 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=4.5903 ps=24.32 w=11.77 l=3.45
X4 VDD1.t7 VP.t2 VTAIL.t18 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=4.5903 ps=24.32 w=11.77 l=3.45
X5 VTAIL.t4 VN.t2 VDD2.t7 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X6 VDD2.t6 VN.t3 VTAIL.t6 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X7 VTAIL.t10 VP.t3 VDD1.t6 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X8 VTAIL.t16 VP.t4 VDD1.t5 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X9 VDD2.t5 VN.t4 VTAIL.t3 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=4.5903 pd=24.32 as=1.94205 ps=12.1 w=11.77 l=3.45
X10 B.t11 B.t9 B.t10 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=4.5903 pd=24.32 as=0 ps=0 w=11.77 l=3.45
X11 B.t8 B.t6 B.t7 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=4.5903 pd=24.32 as=0 ps=0 w=11.77 l=3.45
X12 VDD2.t4 VN.t5 VTAIL.t5 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=4.5903 ps=24.32 w=11.77 l=3.45
X13 VDD2.t3 VN.t6 VTAIL.t7 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X14 B.t5 B.t3 B.t4 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=4.5903 pd=24.32 as=0 ps=0 w=11.77 l=3.45
X15 VDD1.t4 VP.t5 VTAIL.t14 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X16 VDD1.t3 VP.t6 VTAIL.t13 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=4.5903 pd=24.32 as=1.94205 ps=12.1 w=11.77 l=3.45
X17 B.t2 B.t0 B.t1 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=4.5903 pd=24.32 as=0 ps=0 w=11.77 l=3.45
X18 VTAIL.t0 VN.t7 VDD2.t2 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X19 VDD1.t2 VP.t7 VTAIL.t11 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X20 VDD2.t1 VN.t8 VTAIL.t9 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=4.5903 pd=24.32 as=1.94205 ps=12.1 w=11.77 l=3.45
X21 VTAIL.t1 VN.t9 VDD2.t0 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X22 VTAIL.t19 VP.t8 VDD1.t1 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=1.94205 ps=12.1 w=11.77 l=3.45
X23 VDD1.t0 VP.t9 VTAIL.t15 w_n5506_n3322# sky130_fd_pr__pfet_01v8 ad=1.94205 pd=12.1 as=4.5903 ps=24.32 w=11.77 l=3.45
R0 VP.n32 VP.n29 161.3
R1 VP.n34 VP.n33 161.3
R2 VP.n35 VP.n28 161.3
R3 VP.n37 VP.n36 161.3
R4 VP.n38 VP.n27 161.3
R5 VP.n40 VP.n39 161.3
R6 VP.n41 VP.n26 161.3
R7 VP.n44 VP.n43 161.3
R8 VP.n45 VP.n25 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n48 VP.n24 161.3
R11 VP.n50 VP.n49 161.3
R12 VP.n51 VP.n23 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n22 161.3
R15 VP.n56 VP.n55 161.3
R16 VP.n58 VP.n57 161.3
R17 VP.n59 VP.n20 161.3
R18 VP.n61 VP.n60 161.3
R19 VP.n62 VP.n19 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n65 VP.n18 161.3
R22 VP.n67 VP.n66 161.3
R23 VP.n117 VP.n116 161.3
R24 VP.n115 VP.n1 161.3
R25 VP.n114 VP.n113 161.3
R26 VP.n112 VP.n2 161.3
R27 VP.n111 VP.n110 161.3
R28 VP.n109 VP.n3 161.3
R29 VP.n108 VP.n107 161.3
R30 VP.n106 VP.n105 161.3
R31 VP.n104 VP.n5 161.3
R32 VP.n103 VP.n102 161.3
R33 VP.n101 VP.n6 161.3
R34 VP.n100 VP.n99 161.3
R35 VP.n98 VP.n7 161.3
R36 VP.n97 VP.n96 161.3
R37 VP.n95 VP.n8 161.3
R38 VP.n94 VP.n93 161.3
R39 VP.n91 VP.n9 161.3
R40 VP.n90 VP.n89 161.3
R41 VP.n88 VP.n10 161.3
R42 VP.n87 VP.n86 161.3
R43 VP.n85 VP.n11 161.3
R44 VP.n84 VP.n83 161.3
R45 VP.n82 VP.n12 161.3
R46 VP.n81 VP.n80 161.3
R47 VP.n78 VP.n13 161.3
R48 VP.n77 VP.n76 161.3
R49 VP.n75 VP.n14 161.3
R50 VP.n74 VP.n73 161.3
R51 VP.n72 VP.n15 161.3
R52 VP.n71 VP.n70 161.3
R53 VP.n31 VP.t6 115.079
R54 VP.n16 VP.t0 82.2199
R55 VP.n79 VP.t8 82.2199
R56 VP.n92 VP.t5 82.2199
R57 VP.n4 VP.t3 82.2199
R58 VP.n0 VP.t9 82.2199
R59 VP.n17 VP.t2 82.2199
R60 VP.n21 VP.t4 82.2199
R61 VP.n42 VP.t7 82.2199
R62 VP.n30 VP.t1 82.2199
R63 VP.n69 VP.n16 74.8979
R64 VP.n118 VP.n0 74.8979
R65 VP.n68 VP.n17 74.8979
R66 VP.n31 VP.n30 73.2461
R67 VP.n69 VP.n68 57.719
R68 VP.n86 VP.n10 54.0911
R69 VP.n99 VP.n6 54.0911
R70 VP.n49 VP.n23 54.0911
R71 VP.n36 VP.n27 54.0911
R72 VP.n77 VP.n14 48.2635
R73 VP.n110 VP.n2 48.2635
R74 VP.n60 VP.n19 48.2635
R75 VP.n73 VP.n14 32.7233
R76 VP.n114 VP.n2 32.7233
R77 VP.n64 VP.n19 32.7233
R78 VP.n90 VP.n10 26.8957
R79 VP.n99 VP.n98 26.8957
R80 VP.n49 VP.n48 26.8957
R81 VP.n40 VP.n27 26.8957
R82 VP.n72 VP.n71 24.4675
R83 VP.n73 VP.n72 24.4675
R84 VP.n78 VP.n77 24.4675
R85 VP.n80 VP.n78 24.4675
R86 VP.n84 VP.n12 24.4675
R87 VP.n85 VP.n84 24.4675
R88 VP.n86 VP.n85 24.4675
R89 VP.n91 VP.n90 24.4675
R90 VP.n93 VP.n91 24.4675
R91 VP.n97 VP.n8 24.4675
R92 VP.n98 VP.n97 24.4675
R93 VP.n103 VP.n6 24.4675
R94 VP.n104 VP.n103 24.4675
R95 VP.n105 VP.n104 24.4675
R96 VP.n109 VP.n108 24.4675
R97 VP.n110 VP.n109 24.4675
R98 VP.n115 VP.n114 24.4675
R99 VP.n116 VP.n115 24.4675
R100 VP.n65 VP.n64 24.4675
R101 VP.n66 VP.n65 24.4675
R102 VP.n53 VP.n23 24.4675
R103 VP.n54 VP.n53 24.4675
R104 VP.n55 VP.n54 24.4675
R105 VP.n59 VP.n58 24.4675
R106 VP.n60 VP.n59 24.4675
R107 VP.n41 VP.n40 24.4675
R108 VP.n43 VP.n41 24.4675
R109 VP.n47 VP.n25 24.4675
R110 VP.n48 VP.n47 24.4675
R111 VP.n34 VP.n29 24.4675
R112 VP.n35 VP.n34 24.4675
R113 VP.n36 VP.n35 24.4675
R114 VP.n80 VP.n79 22.9995
R115 VP.n108 VP.n4 22.9995
R116 VP.n58 VP.n21 22.9995
R117 VP.n71 VP.n16 15.17
R118 VP.n116 VP.n0 15.17
R119 VP.n66 VP.n17 15.17
R120 VP.n93 VP.n92 12.234
R121 VP.n92 VP.n8 12.234
R122 VP.n43 VP.n42 12.234
R123 VP.n42 VP.n25 12.234
R124 VP.n32 VP.n31 4.14768
R125 VP.n79 VP.n12 1.46852
R126 VP.n105 VP.n4 1.46852
R127 VP.n55 VP.n21 1.46852
R128 VP.n30 VP.n29 1.46852
R129 VP.n68 VP.n67 0.354971
R130 VP.n70 VP.n69 0.354971
R131 VP.n118 VP.n117 0.354971
R132 VP VP.n118 0.26696
R133 VP.n33 VP.n32 0.189894
R134 VP.n33 VP.n28 0.189894
R135 VP.n37 VP.n28 0.189894
R136 VP.n38 VP.n37 0.189894
R137 VP.n39 VP.n38 0.189894
R138 VP.n39 VP.n26 0.189894
R139 VP.n44 VP.n26 0.189894
R140 VP.n45 VP.n44 0.189894
R141 VP.n46 VP.n45 0.189894
R142 VP.n46 VP.n24 0.189894
R143 VP.n50 VP.n24 0.189894
R144 VP.n51 VP.n50 0.189894
R145 VP.n52 VP.n51 0.189894
R146 VP.n52 VP.n22 0.189894
R147 VP.n56 VP.n22 0.189894
R148 VP.n57 VP.n56 0.189894
R149 VP.n57 VP.n20 0.189894
R150 VP.n61 VP.n20 0.189894
R151 VP.n62 VP.n61 0.189894
R152 VP.n63 VP.n62 0.189894
R153 VP.n63 VP.n18 0.189894
R154 VP.n67 VP.n18 0.189894
R155 VP.n70 VP.n15 0.189894
R156 VP.n74 VP.n15 0.189894
R157 VP.n75 VP.n74 0.189894
R158 VP.n76 VP.n75 0.189894
R159 VP.n76 VP.n13 0.189894
R160 VP.n81 VP.n13 0.189894
R161 VP.n82 VP.n81 0.189894
R162 VP.n83 VP.n82 0.189894
R163 VP.n83 VP.n11 0.189894
R164 VP.n87 VP.n11 0.189894
R165 VP.n88 VP.n87 0.189894
R166 VP.n89 VP.n88 0.189894
R167 VP.n89 VP.n9 0.189894
R168 VP.n94 VP.n9 0.189894
R169 VP.n95 VP.n94 0.189894
R170 VP.n96 VP.n95 0.189894
R171 VP.n96 VP.n7 0.189894
R172 VP.n100 VP.n7 0.189894
R173 VP.n101 VP.n100 0.189894
R174 VP.n102 VP.n101 0.189894
R175 VP.n102 VP.n5 0.189894
R176 VP.n106 VP.n5 0.189894
R177 VP.n107 VP.n106 0.189894
R178 VP.n107 VP.n3 0.189894
R179 VP.n111 VP.n3 0.189894
R180 VP.n112 VP.n111 0.189894
R181 VP.n113 VP.n112 0.189894
R182 VP.n113 VP.n1 0.189894
R183 VP.n117 VP.n1 0.189894
R184 VTAIL.n11 VTAIL.t5 60.5718
R185 VTAIL.n17 VTAIL.t2 60.5715
R186 VTAIL.n2 VTAIL.t15 60.5715
R187 VTAIL.n16 VTAIL.t18 60.5715
R188 VTAIL.n15 VTAIL.n14 57.8101
R189 VTAIL.n13 VTAIL.n12 57.8101
R190 VTAIL.n10 VTAIL.n9 57.8101
R191 VTAIL.n8 VTAIL.n7 57.8101
R192 VTAIL.n19 VTAIL.n18 57.8098
R193 VTAIL.n1 VTAIL.n0 57.8098
R194 VTAIL.n4 VTAIL.n3 57.8098
R195 VTAIL.n6 VTAIL.n5 57.8098
R196 VTAIL.n8 VTAIL.n6 29.0307
R197 VTAIL.n17 VTAIL.n16 25.7721
R198 VTAIL.n10 VTAIL.n8 3.25912
R199 VTAIL.n11 VTAIL.n10 3.25912
R200 VTAIL.n15 VTAIL.n13 3.25912
R201 VTAIL.n16 VTAIL.n15 3.25912
R202 VTAIL.n6 VTAIL.n4 3.25912
R203 VTAIL.n4 VTAIL.n2 3.25912
R204 VTAIL.n19 VTAIL.n17 3.25912
R205 VTAIL.n18 VTAIL.t7 2.76218
R206 VTAIL.n18 VTAIL.t0 2.76218
R207 VTAIL.n0 VTAIL.t9 2.76218
R208 VTAIL.n0 VTAIL.t8 2.76218
R209 VTAIL.n3 VTAIL.t14 2.76218
R210 VTAIL.n3 VTAIL.t10 2.76218
R211 VTAIL.n5 VTAIL.t12 2.76218
R212 VTAIL.n5 VTAIL.t19 2.76218
R213 VTAIL.n14 VTAIL.t11 2.76218
R214 VTAIL.n14 VTAIL.t16 2.76218
R215 VTAIL.n12 VTAIL.t13 2.76218
R216 VTAIL.n12 VTAIL.t17 2.76218
R217 VTAIL.n9 VTAIL.t6 2.76218
R218 VTAIL.n9 VTAIL.t4 2.76218
R219 VTAIL.n7 VTAIL.t3 2.76218
R220 VTAIL.n7 VTAIL.t1 2.76218
R221 VTAIL VTAIL.n1 2.50266
R222 VTAIL.n13 VTAIL.n11 2.09964
R223 VTAIL.n2 VTAIL.n1 2.09964
R224 VTAIL VTAIL.n19 0.756965
R225 VDD1.n1 VDD1.t3 80.5092
R226 VDD1.n3 VDD1.t9 80.5089
R227 VDD1.n5 VDD1.n4 76.8772
R228 VDD1.n1 VDD1.n0 74.4889
R229 VDD1.n7 VDD1.n6 74.4887
R230 VDD1.n3 VDD1.n2 74.4886
R231 VDD1.n7 VDD1.n5 51.5526
R232 VDD1.n6 VDD1.t5 2.76218
R233 VDD1.n6 VDD1.t7 2.76218
R234 VDD1.n0 VDD1.t8 2.76218
R235 VDD1.n0 VDD1.t2 2.76218
R236 VDD1.n4 VDD1.t6 2.76218
R237 VDD1.n4 VDD1.t0 2.76218
R238 VDD1.n2 VDD1.t1 2.76218
R239 VDD1.n2 VDD1.t4 2.76218
R240 VDD1 VDD1.n7 2.38628
R241 VDD1 VDD1.n1 0.873345
R242 VDD1.n5 VDD1.n3 0.759809
R243 VN.n102 VN.n101 161.3
R244 VN.n100 VN.n53 161.3
R245 VN.n99 VN.n98 161.3
R246 VN.n97 VN.n54 161.3
R247 VN.n96 VN.n95 161.3
R248 VN.n94 VN.n55 161.3
R249 VN.n93 VN.n92 161.3
R250 VN.n91 VN.n90 161.3
R251 VN.n89 VN.n57 161.3
R252 VN.n88 VN.n87 161.3
R253 VN.n86 VN.n58 161.3
R254 VN.n85 VN.n84 161.3
R255 VN.n83 VN.n59 161.3
R256 VN.n82 VN.n81 161.3
R257 VN.n80 VN.n60 161.3
R258 VN.n79 VN.n78 161.3
R259 VN.n77 VN.n61 161.3
R260 VN.n76 VN.n75 161.3
R261 VN.n74 VN.n63 161.3
R262 VN.n73 VN.n72 161.3
R263 VN.n71 VN.n64 161.3
R264 VN.n70 VN.n69 161.3
R265 VN.n68 VN.n65 161.3
R266 VN.n50 VN.n49 161.3
R267 VN.n48 VN.n1 161.3
R268 VN.n47 VN.n46 161.3
R269 VN.n45 VN.n2 161.3
R270 VN.n44 VN.n43 161.3
R271 VN.n42 VN.n3 161.3
R272 VN.n41 VN.n40 161.3
R273 VN.n39 VN.n38 161.3
R274 VN.n37 VN.n5 161.3
R275 VN.n36 VN.n35 161.3
R276 VN.n34 VN.n6 161.3
R277 VN.n33 VN.n32 161.3
R278 VN.n31 VN.n7 161.3
R279 VN.n30 VN.n29 161.3
R280 VN.n28 VN.n8 161.3
R281 VN.n27 VN.n26 161.3
R282 VN.n24 VN.n9 161.3
R283 VN.n23 VN.n22 161.3
R284 VN.n21 VN.n10 161.3
R285 VN.n20 VN.n19 161.3
R286 VN.n18 VN.n11 161.3
R287 VN.n17 VN.n16 161.3
R288 VN.n15 VN.n12 161.3
R289 VN.n14 VN.t8 115.079
R290 VN.n67 VN.t5 115.079
R291 VN.n13 VN.t0 82.2199
R292 VN.n25 VN.t6 82.2199
R293 VN.n4 VN.t7 82.2199
R294 VN.n0 VN.t1 82.2199
R295 VN.n66 VN.t2 82.2199
R296 VN.n62 VN.t3 82.2199
R297 VN.n56 VN.t9 82.2199
R298 VN.n52 VN.t4 82.2199
R299 VN.n51 VN.n0 74.8979
R300 VN.n103 VN.n52 74.8979
R301 VN.n14 VN.n13 73.246
R302 VN.n67 VN.n66 73.246
R303 VN VN.n103 57.8844
R304 VN.n19 VN.n10 54.0911
R305 VN.n32 VN.n6 54.0911
R306 VN.n72 VN.n63 54.0911
R307 VN.n84 VN.n58 54.0911
R308 VN.n43 VN.n2 48.2635
R309 VN.n95 VN.n54 48.2635
R310 VN.n47 VN.n2 32.7233
R311 VN.n99 VN.n54 32.7233
R312 VN.n23 VN.n10 26.8957
R313 VN.n32 VN.n31 26.8957
R314 VN.n76 VN.n63 26.8957
R315 VN.n84 VN.n83 26.8957
R316 VN.n17 VN.n12 24.4675
R317 VN.n18 VN.n17 24.4675
R318 VN.n19 VN.n18 24.4675
R319 VN.n24 VN.n23 24.4675
R320 VN.n26 VN.n24 24.4675
R321 VN.n30 VN.n8 24.4675
R322 VN.n31 VN.n30 24.4675
R323 VN.n36 VN.n6 24.4675
R324 VN.n37 VN.n36 24.4675
R325 VN.n38 VN.n37 24.4675
R326 VN.n42 VN.n41 24.4675
R327 VN.n43 VN.n42 24.4675
R328 VN.n48 VN.n47 24.4675
R329 VN.n49 VN.n48 24.4675
R330 VN.n72 VN.n71 24.4675
R331 VN.n71 VN.n70 24.4675
R332 VN.n70 VN.n65 24.4675
R333 VN.n83 VN.n82 24.4675
R334 VN.n82 VN.n60 24.4675
R335 VN.n78 VN.n77 24.4675
R336 VN.n77 VN.n76 24.4675
R337 VN.n95 VN.n94 24.4675
R338 VN.n94 VN.n93 24.4675
R339 VN.n90 VN.n89 24.4675
R340 VN.n89 VN.n88 24.4675
R341 VN.n88 VN.n58 24.4675
R342 VN.n101 VN.n100 24.4675
R343 VN.n100 VN.n99 24.4675
R344 VN.n41 VN.n4 22.9995
R345 VN.n93 VN.n56 22.9995
R346 VN.n49 VN.n0 15.17
R347 VN.n101 VN.n52 15.17
R348 VN.n26 VN.n25 12.234
R349 VN.n25 VN.n8 12.234
R350 VN.n62 VN.n60 12.234
R351 VN.n78 VN.n62 12.234
R352 VN.n15 VN.n14 4.14771
R353 VN.n68 VN.n67 4.14771
R354 VN.n13 VN.n12 1.46852
R355 VN.n38 VN.n4 1.46852
R356 VN.n66 VN.n65 1.46852
R357 VN.n90 VN.n56 1.46852
R358 VN.n103 VN.n102 0.354971
R359 VN.n51 VN.n50 0.354971
R360 VN VN.n51 0.26696
R361 VN.n102 VN.n53 0.189894
R362 VN.n98 VN.n53 0.189894
R363 VN.n98 VN.n97 0.189894
R364 VN.n97 VN.n96 0.189894
R365 VN.n96 VN.n55 0.189894
R366 VN.n92 VN.n55 0.189894
R367 VN.n92 VN.n91 0.189894
R368 VN.n91 VN.n57 0.189894
R369 VN.n87 VN.n57 0.189894
R370 VN.n87 VN.n86 0.189894
R371 VN.n86 VN.n85 0.189894
R372 VN.n85 VN.n59 0.189894
R373 VN.n81 VN.n59 0.189894
R374 VN.n81 VN.n80 0.189894
R375 VN.n80 VN.n79 0.189894
R376 VN.n79 VN.n61 0.189894
R377 VN.n75 VN.n61 0.189894
R378 VN.n75 VN.n74 0.189894
R379 VN.n74 VN.n73 0.189894
R380 VN.n73 VN.n64 0.189894
R381 VN.n69 VN.n64 0.189894
R382 VN.n69 VN.n68 0.189894
R383 VN.n16 VN.n15 0.189894
R384 VN.n16 VN.n11 0.189894
R385 VN.n20 VN.n11 0.189894
R386 VN.n21 VN.n20 0.189894
R387 VN.n22 VN.n21 0.189894
R388 VN.n22 VN.n9 0.189894
R389 VN.n27 VN.n9 0.189894
R390 VN.n28 VN.n27 0.189894
R391 VN.n29 VN.n28 0.189894
R392 VN.n29 VN.n7 0.189894
R393 VN.n33 VN.n7 0.189894
R394 VN.n34 VN.n33 0.189894
R395 VN.n35 VN.n34 0.189894
R396 VN.n35 VN.n5 0.189894
R397 VN.n39 VN.n5 0.189894
R398 VN.n40 VN.n39 0.189894
R399 VN.n40 VN.n3 0.189894
R400 VN.n44 VN.n3 0.189894
R401 VN.n45 VN.n44 0.189894
R402 VN.n46 VN.n45 0.189894
R403 VN.n46 VN.n1 0.189894
R404 VN.n50 VN.n1 0.189894
R405 VDD2.n1 VDD2.t1 80.5089
R406 VDD2.n4 VDD2.t5 77.2505
R407 VDD2.n3 VDD2.n2 76.8772
R408 VDD2 VDD2.n7 76.8745
R409 VDD2.n6 VDD2.n5 74.4889
R410 VDD2.n1 VDD2.n0 74.4886
R411 VDD2.n4 VDD2.n3 49.3403
R412 VDD2.n6 VDD2.n4 3.25912
R413 VDD2.n7 VDD2.t7 2.76218
R414 VDD2.n7 VDD2.t4 2.76218
R415 VDD2.n5 VDD2.t0 2.76218
R416 VDD2.n5 VDD2.t6 2.76218
R417 VDD2.n2 VDD2.t2 2.76218
R418 VDD2.n2 VDD2.t8 2.76218
R419 VDD2.n0 VDD2.t9 2.76218
R420 VDD2.n0 VDD2.t3 2.76218
R421 VDD2 VDD2.n6 0.873345
R422 VDD2.n3 VDD2.n1 0.759809
R423 B.n728 B.n89 585
R424 B.n730 B.n729 585
R425 B.n731 B.n88 585
R426 B.n733 B.n732 585
R427 B.n734 B.n87 585
R428 B.n736 B.n735 585
R429 B.n737 B.n86 585
R430 B.n739 B.n738 585
R431 B.n740 B.n85 585
R432 B.n742 B.n741 585
R433 B.n743 B.n84 585
R434 B.n745 B.n744 585
R435 B.n746 B.n83 585
R436 B.n748 B.n747 585
R437 B.n749 B.n82 585
R438 B.n751 B.n750 585
R439 B.n752 B.n81 585
R440 B.n754 B.n753 585
R441 B.n755 B.n80 585
R442 B.n757 B.n756 585
R443 B.n758 B.n79 585
R444 B.n760 B.n759 585
R445 B.n761 B.n78 585
R446 B.n763 B.n762 585
R447 B.n764 B.n77 585
R448 B.n766 B.n765 585
R449 B.n767 B.n76 585
R450 B.n769 B.n768 585
R451 B.n770 B.n75 585
R452 B.n772 B.n771 585
R453 B.n773 B.n74 585
R454 B.n775 B.n774 585
R455 B.n776 B.n73 585
R456 B.n778 B.n777 585
R457 B.n779 B.n72 585
R458 B.n781 B.n780 585
R459 B.n782 B.n71 585
R460 B.n784 B.n783 585
R461 B.n785 B.n70 585
R462 B.n787 B.n786 585
R463 B.n788 B.n67 585
R464 B.n791 B.n790 585
R465 B.n792 B.n66 585
R466 B.n794 B.n793 585
R467 B.n795 B.n65 585
R468 B.n797 B.n796 585
R469 B.n798 B.n64 585
R470 B.n800 B.n799 585
R471 B.n801 B.n63 585
R472 B.n803 B.n802 585
R473 B.n805 B.n804 585
R474 B.n806 B.n59 585
R475 B.n808 B.n807 585
R476 B.n809 B.n58 585
R477 B.n811 B.n810 585
R478 B.n812 B.n57 585
R479 B.n814 B.n813 585
R480 B.n815 B.n56 585
R481 B.n817 B.n816 585
R482 B.n818 B.n55 585
R483 B.n820 B.n819 585
R484 B.n821 B.n54 585
R485 B.n823 B.n822 585
R486 B.n824 B.n53 585
R487 B.n826 B.n825 585
R488 B.n827 B.n52 585
R489 B.n829 B.n828 585
R490 B.n830 B.n51 585
R491 B.n832 B.n831 585
R492 B.n833 B.n50 585
R493 B.n835 B.n834 585
R494 B.n836 B.n49 585
R495 B.n838 B.n837 585
R496 B.n839 B.n48 585
R497 B.n841 B.n840 585
R498 B.n842 B.n47 585
R499 B.n844 B.n843 585
R500 B.n845 B.n46 585
R501 B.n847 B.n846 585
R502 B.n848 B.n45 585
R503 B.n850 B.n849 585
R504 B.n851 B.n44 585
R505 B.n853 B.n852 585
R506 B.n854 B.n43 585
R507 B.n856 B.n855 585
R508 B.n857 B.n42 585
R509 B.n859 B.n858 585
R510 B.n860 B.n41 585
R511 B.n862 B.n861 585
R512 B.n863 B.n40 585
R513 B.n865 B.n864 585
R514 B.n727 B.n726 585
R515 B.n725 B.n90 585
R516 B.n724 B.n723 585
R517 B.n722 B.n91 585
R518 B.n721 B.n720 585
R519 B.n719 B.n92 585
R520 B.n718 B.n717 585
R521 B.n716 B.n93 585
R522 B.n715 B.n714 585
R523 B.n713 B.n94 585
R524 B.n712 B.n711 585
R525 B.n710 B.n95 585
R526 B.n709 B.n708 585
R527 B.n707 B.n96 585
R528 B.n706 B.n705 585
R529 B.n704 B.n97 585
R530 B.n703 B.n702 585
R531 B.n701 B.n98 585
R532 B.n700 B.n699 585
R533 B.n698 B.n99 585
R534 B.n697 B.n696 585
R535 B.n695 B.n100 585
R536 B.n694 B.n693 585
R537 B.n692 B.n101 585
R538 B.n691 B.n690 585
R539 B.n689 B.n102 585
R540 B.n688 B.n687 585
R541 B.n686 B.n103 585
R542 B.n685 B.n684 585
R543 B.n683 B.n104 585
R544 B.n682 B.n681 585
R545 B.n680 B.n105 585
R546 B.n679 B.n678 585
R547 B.n677 B.n106 585
R548 B.n676 B.n675 585
R549 B.n674 B.n107 585
R550 B.n673 B.n672 585
R551 B.n671 B.n108 585
R552 B.n670 B.n669 585
R553 B.n668 B.n109 585
R554 B.n667 B.n666 585
R555 B.n665 B.n110 585
R556 B.n664 B.n663 585
R557 B.n662 B.n111 585
R558 B.n661 B.n660 585
R559 B.n659 B.n112 585
R560 B.n658 B.n657 585
R561 B.n656 B.n113 585
R562 B.n655 B.n654 585
R563 B.n653 B.n114 585
R564 B.n652 B.n651 585
R565 B.n650 B.n115 585
R566 B.n649 B.n648 585
R567 B.n647 B.n116 585
R568 B.n646 B.n645 585
R569 B.n644 B.n117 585
R570 B.n643 B.n642 585
R571 B.n641 B.n118 585
R572 B.n640 B.n639 585
R573 B.n638 B.n119 585
R574 B.n637 B.n636 585
R575 B.n635 B.n120 585
R576 B.n634 B.n633 585
R577 B.n632 B.n121 585
R578 B.n631 B.n630 585
R579 B.n629 B.n122 585
R580 B.n628 B.n627 585
R581 B.n626 B.n123 585
R582 B.n625 B.n624 585
R583 B.n623 B.n124 585
R584 B.n622 B.n621 585
R585 B.n620 B.n125 585
R586 B.n619 B.n618 585
R587 B.n617 B.n126 585
R588 B.n616 B.n615 585
R589 B.n614 B.n127 585
R590 B.n613 B.n612 585
R591 B.n611 B.n128 585
R592 B.n610 B.n609 585
R593 B.n608 B.n129 585
R594 B.n607 B.n606 585
R595 B.n605 B.n130 585
R596 B.n604 B.n603 585
R597 B.n602 B.n131 585
R598 B.n601 B.n600 585
R599 B.n599 B.n132 585
R600 B.n598 B.n597 585
R601 B.n596 B.n133 585
R602 B.n595 B.n594 585
R603 B.n593 B.n134 585
R604 B.n592 B.n591 585
R605 B.n590 B.n135 585
R606 B.n589 B.n588 585
R607 B.n587 B.n136 585
R608 B.n586 B.n585 585
R609 B.n584 B.n137 585
R610 B.n583 B.n582 585
R611 B.n581 B.n138 585
R612 B.n580 B.n579 585
R613 B.n578 B.n139 585
R614 B.n577 B.n576 585
R615 B.n575 B.n140 585
R616 B.n574 B.n573 585
R617 B.n572 B.n141 585
R618 B.n571 B.n570 585
R619 B.n569 B.n142 585
R620 B.n568 B.n567 585
R621 B.n566 B.n143 585
R622 B.n565 B.n564 585
R623 B.n563 B.n144 585
R624 B.n562 B.n561 585
R625 B.n560 B.n145 585
R626 B.n559 B.n558 585
R627 B.n557 B.n146 585
R628 B.n556 B.n555 585
R629 B.n554 B.n147 585
R630 B.n553 B.n552 585
R631 B.n551 B.n148 585
R632 B.n550 B.n549 585
R633 B.n548 B.n149 585
R634 B.n547 B.n546 585
R635 B.n545 B.n150 585
R636 B.n544 B.n543 585
R637 B.n542 B.n151 585
R638 B.n541 B.n540 585
R639 B.n539 B.n152 585
R640 B.n538 B.n537 585
R641 B.n536 B.n153 585
R642 B.n535 B.n534 585
R643 B.n533 B.n154 585
R644 B.n532 B.n531 585
R645 B.n530 B.n155 585
R646 B.n529 B.n528 585
R647 B.n527 B.n156 585
R648 B.n526 B.n525 585
R649 B.n524 B.n157 585
R650 B.n523 B.n522 585
R651 B.n521 B.n158 585
R652 B.n520 B.n519 585
R653 B.n518 B.n159 585
R654 B.n517 B.n516 585
R655 B.n515 B.n160 585
R656 B.n514 B.n513 585
R657 B.n512 B.n161 585
R658 B.n511 B.n510 585
R659 B.n509 B.n162 585
R660 B.n508 B.n507 585
R661 B.n506 B.n163 585
R662 B.n505 B.n504 585
R663 B.n503 B.n164 585
R664 B.n502 B.n501 585
R665 B.n364 B.n363 585
R666 B.n365 B.n214 585
R667 B.n367 B.n366 585
R668 B.n368 B.n213 585
R669 B.n370 B.n369 585
R670 B.n371 B.n212 585
R671 B.n373 B.n372 585
R672 B.n374 B.n211 585
R673 B.n376 B.n375 585
R674 B.n377 B.n210 585
R675 B.n379 B.n378 585
R676 B.n380 B.n209 585
R677 B.n382 B.n381 585
R678 B.n383 B.n208 585
R679 B.n385 B.n384 585
R680 B.n386 B.n207 585
R681 B.n388 B.n387 585
R682 B.n389 B.n206 585
R683 B.n391 B.n390 585
R684 B.n392 B.n205 585
R685 B.n394 B.n393 585
R686 B.n395 B.n204 585
R687 B.n397 B.n396 585
R688 B.n398 B.n203 585
R689 B.n400 B.n399 585
R690 B.n401 B.n202 585
R691 B.n403 B.n402 585
R692 B.n404 B.n201 585
R693 B.n406 B.n405 585
R694 B.n407 B.n200 585
R695 B.n409 B.n408 585
R696 B.n410 B.n199 585
R697 B.n412 B.n411 585
R698 B.n413 B.n198 585
R699 B.n415 B.n414 585
R700 B.n416 B.n197 585
R701 B.n418 B.n417 585
R702 B.n419 B.n196 585
R703 B.n421 B.n420 585
R704 B.n422 B.n195 585
R705 B.n424 B.n423 585
R706 B.n426 B.n425 585
R707 B.n427 B.n191 585
R708 B.n429 B.n428 585
R709 B.n430 B.n190 585
R710 B.n432 B.n431 585
R711 B.n433 B.n189 585
R712 B.n435 B.n434 585
R713 B.n436 B.n188 585
R714 B.n438 B.n437 585
R715 B.n440 B.n185 585
R716 B.n442 B.n441 585
R717 B.n443 B.n184 585
R718 B.n445 B.n444 585
R719 B.n446 B.n183 585
R720 B.n448 B.n447 585
R721 B.n449 B.n182 585
R722 B.n451 B.n450 585
R723 B.n452 B.n181 585
R724 B.n454 B.n453 585
R725 B.n455 B.n180 585
R726 B.n457 B.n456 585
R727 B.n458 B.n179 585
R728 B.n460 B.n459 585
R729 B.n461 B.n178 585
R730 B.n463 B.n462 585
R731 B.n464 B.n177 585
R732 B.n466 B.n465 585
R733 B.n467 B.n176 585
R734 B.n469 B.n468 585
R735 B.n470 B.n175 585
R736 B.n472 B.n471 585
R737 B.n473 B.n174 585
R738 B.n475 B.n474 585
R739 B.n476 B.n173 585
R740 B.n478 B.n477 585
R741 B.n479 B.n172 585
R742 B.n481 B.n480 585
R743 B.n482 B.n171 585
R744 B.n484 B.n483 585
R745 B.n485 B.n170 585
R746 B.n487 B.n486 585
R747 B.n488 B.n169 585
R748 B.n490 B.n489 585
R749 B.n491 B.n168 585
R750 B.n493 B.n492 585
R751 B.n494 B.n167 585
R752 B.n496 B.n495 585
R753 B.n497 B.n166 585
R754 B.n499 B.n498 585
R755 B.n500 B.n165 585
R756 B.n362 B.n215 585
R757 B.n361 B.n360 585
R758 B.n359 B.n216 585
R759 B.n358 B.n357 585
R760 B.n356 B.n217 585
R761 B.n355 B.n354 585
R762 B.n353 B.n218 585
R763 B.n352 B.n351 585
R764 B.n350 B.n219 585
R765 B.n349 B.n348 585
R766 B.n347 B.n220 585
R767 B.n346 B.n345 585
R768 B.n344 B.n221 585
R769 B.n343 B.n342 585
R770 B.n341 B.n222 585
R771 B.n340 B.n339 585
R772 B.n338 B.n223 585
R773 B.n337 B.n336 585
R774 B.n335 B.n224 585
R775 B.n334 B.n333 585
R776 B.n332 B.n225 585
R777 B.n331 B.n330 585
R778 B.n329 B.n226 585
R779 B.n328 B.n327 585
R780 B.n326 B.n227 585
R781 B.n325 B.n324 585
R782 B.n323 B.n228 585
R783 B.n322 B.n321 585
R784 B.n320 B.n229 585
R785 B.n319 B.n318 585
R786 B.n317 B.n230 585
R787 B.n316 B.n315 585
R788 B.n314 B.n231 585
R789 B.n313 B.n312 585
R790 B.n311 B.n232 585
R791 B.n310 B.n309 585
R792 B.n308 B.n233 585
R793 B.n307 B.n306 585
R794 B.n305 B.n234 585
R795 B.n304 B.n303 585
R796 B.n302 B.n235 585
R797 B.n301 B.n300 585
R798 B.n299 B.n236 585
R799 B.n298 B.n297 585
R800 B.n296 B.n237 585
R801 B.n295 B.n294 585
R802 B.n293 B.n238 585
R803 B.n292 B.n291 585
R804 B.n290 B.n239 585
R805 B.n289 B.n288 585
R806 B.n287 B.n240 585
R807 B.n286 B.n285 585
R808 B.n284 B.n241 585
R809 B.n283 B.n282 585
R810 B.n281 B.n242 585
R811 B.n280 B.n279 585
R812 B.n278 B.n243 585
R813 B.n277 B.n276 585
R814 B.n275 B.n244 585
R815 B.n274 B.n273 585
R816 B.n272 B.n245 585
R817 B.n271 B.n270 585
R818 B.n269 B.n246 585
R819 B.n268 B.n267 585
R820 B.n266 B.n247 585
R821 B.n265 B.n264 585
R822 B.n263 B.n248 585
R823 B.n262 B.n261 585
R824 B.n260 B.n249 585
R825 B.n259 B.n258 585
R826 B.n257 B.n250 585
R827 B.n256 B.n255 585
R828 B.n254 B.n251 585
R829 B.n253 B.n252 585
R830 B.n2 B.n0 585
R831 B.n977 B.n1 585
R832 B.n976 B.n975 585
R833 B.n974 B.n3 585
R834 B.n973 B.n972 585
R835 B.n971 B.n4 585
R836 B.n970 B.n969 585
R837 B.n968 B.n5 585
R838 B.n967 B.n966 585
R839 B.n965 B.n6 585
R840 B.n964 B.n963 585
R841 B.n962 B.n7 585
R842 B.n961 B.n960 585
R843 B.n959 B.n8 585
R844 B.n958 B.n957 585
R845 B.n956 B.n9 585
R846 B.n955 B.n954 585
R847 B.n953 B.n10 585
R848 B.n952 B.n951 585
R849 B.n950 B.n11 585
R850 B.n949 B.n948 585
R851 B.n947 B.n12 585
R852 B.n946 B.n945 585
R853 B.n944 B.n13 585
R854 B.n943 B.n942 585
R855 B.n941 B.n14 585
R856 B.n940 B.n939 585
R857 B.n938 B.n15 585
R858 B.n937 B.n936 585
R859 B.n935 B.n16 585
R860 B.n934 B.n933 585
R861 B.n932 B.n17 585
R862 B.n931 B.n930 585
R863 B.n929 B.n18 585
R864 B.n928 B.n927 585
R865 B.n926 B.n19 585
R866 B.n925 B.n924 585
R867 B.n923 B.n20 585
R868 B.n922 B.n921 585
R869 B.n920 B.n21 585
R870 B.n919 B.n918 585
R871 B.n917 B.n22 585
R872 B.n916 B.n915 585
R873 B.n914 B.n23 585
R874 B.n913 B.n912 585
R875 B.n911 B.n24 585
R876 B.n910 B.n909 585
R877 B.n908 B.n25 585
R878 B.n907 B.n906 585
R879 B.n905 B.n26 585
R880 B.n904 B.n903 585
R881 B.n902 B.n27 585
R882 B.n901 B.n900 585
R883 B.n899 B.n28 585
R884 B.n898 B.n897 585
R885 B.n896 B.n29 585
R886 B.n895 B.n894 585
R887 B.n893 B.n30 585
R888 B.n892 B.n891 585
R889 B.n890 B.n31 585
R890 B.n889 B.n888 585
R891 B.n887 B.n32 585
R892 B.n886 B.n885 585
R893 B.n884 B.n33 585
R894 B.n883 B.n882 585
R895 B.n881 B.n34 585
R896 B.n880 B.n879 585
R897 B.n878 B.n35 585
R898 B.n877 B.n876 585
R899 B.n875 B.n36 585
R900 B.n874 B.n873 585
R901 B.n872 B.n37 585
R902 B.n871 B.n870 585
R903 B.n869 B.n38 585
R904 B.n868 B.n867 585
R905 B.n866 B.n39 585
R906 B.n979 B.n978 585
R907 B.n364 B.n215 506.916
R908 B.n864 B.n39 506.916
R909 B.n502 B.n165 506.916
R910 B.n726 B.n89 506.916
R911 B.n186 B.t9 291.269
R912 B.n192 B.t3 291.269
R913 B.n60 B.t6 291.269
R914 B.n68 B.t0 291.269
R915 B.n186 B.t11 184.542
R916 B.n68 B.t1 184.542
R917 B.n192 B.t5 184.528
R918 B.n60 B.t7 184.528
R919 B.n360 B.n215 163.367
R920 B.n360 B.n359 163.367
R921 B.n359 B.n358 163.367
R922 B.n358 B.n217 163.367
R923 B.n354 B.n217 163.367
R924 B.n354 B.n353 163.367
R925 B.n353 B.n352 163.367
R926 B.n352 B.n219 163.367
R927 B.n348 B.n219 163.367
R928 B.n348 B.n347 163.367
R929 B.n347 B.n346 163.367
R930 B.n346 B.n221 163.367
R931 B.n342 B.n221 163.367
R932 B.n342 B.n341 163.367
R933 B.n341 B.n340 163.367
R934 B.n340 B.n223 163.367
R935 B.n336 B.n223 163.367
R936 B.n336 B.n335 163.367
R937 B.n335 B.n334 163.367
R938 B.n334 B.n225 163.367
R939 B.n330 B.n225 163.367
R940 B.n330 B.n329 163.367
R941 B.n329 B.n328 163.367
R942 B.n328 B.n227 163.367
R943 B.n324 B.n227 163.367
R944 B.n324 B.n323 163.367
R945 B.n323 B.n322 163.367
R946 B.n322 B.n229 163.367
R947 B.n318 B.n229 163.367
R948 B.n318 B.n317 163.367
R949 B.n317 B.n316 163.367
R950 B.n316 B.n231 163.367
R951 B.n312 B.n231 163.367
R952 B.n312 B.n311 163.367
R953 B.n311 B.n310 163.367
R954 B.n310 B.n233 163.367
R955 B.n306 B.n233 163.367
R956 B.n306 B.n305 163.367
R957 B.n305 B.n304 163.367
R958 B.n304 B.n235 163.367
R959 B.n300 B.n235 163.367
R960 B.n300 B.n299 163.367
R961 B.n299 B.n298 163.367
R962 B.n298 B.n237 163.367
R963 B.n294 B.n237 163.367
R964 B.n294 B.n293 163.367
R965 B.n293 B.n292 163.367
R966 B.n292 B.n239 163.367
R967 B.n288 B.n239 163.367
R968 B.n288 B.n287 163.367
R969 B.n287 B.n286 163.367
R970 B.n286 B.n241 163.367
R971 B.n282 B.n241 163.367
R972 B.n282 B.n281 163.367
R973 B.n281 B.n280 163.367
R974 B.n280 B.n243 163.367
R975 B.n276 B.n243 163.367
R976 B.n276 B.n275 163.367
R977 B.n275 B.n274 163.367
R978 B.n274 B.n245 163.367
R979 B.n270 B.n245 163.367
R980 B.n270 B.n269 163.367
R981 B.n269 B.n268 163.367
R982 B.n268 B.n247 163.367
R983 B.n264 B.n247 163.367
R984 B.n264 B.n263 163.367
R985 B.n263 B.n262 163.367
R986 B.n262 B.n249 163.367
R987 B.n258 B.n249 163.367
R988 B.n258 B.n257 163.367
R989 B.n257 B.n256 163.367
R990 B.n256 B.n251 163.367
R991 B.n252 B.n251 163.367
R992 B.n252 B.n2 163.367
R993 B.n978 B.n2 163.367
R994 B.n978 B.n977 163.367
R995 B.n977 B.n976 163.367
R996 B.n976 B.n3 163.367
R997 B.n972 B.n3 163.367
R998 B.n972 B.n971 163.367
R999 B.n971 B.n970 163.367
R1000 B.n970 B.n5 163.367
R1001 B.n966 B.n5 163.367
R1002 B.n966 B.n965 163.367
R1003 B.n965 B.n964 163.367
R1004 B.n964 B.n7 163.367
R1005 B.n960 B.n7 163.367
R1006 B.n960 B.n959 163.367
R1007 B.n959 B.n958 163.367
R1008 B.n958 B.n9 163.367
R1009 B.n954 B.n9 163.367
R1010 B.n954 B.n953 163.367
R1011 B.n953 B.n952 163.367
R1012 B.n952 B.n11 163.367
R1013 B.n948 B.n11 163.367
R1014 B.n948 B.n947 163.367
R1015 B.n947 B.n946 163.367
R1016 B.n946 B.n13 163.367
R1017 B.n942 B.n13 163.367
R1018 B.n942 B.n941 163.367
R1019 B.n941 B.n940 163.367
R1020 B.n940 B.n15 163.367
R1021 B.n936 B.n15 163.367
R1022 B.n936 B.n935 163.367
R1023 B.n935 B.n934 163.367
R1024 B.n934 B.n17 163.367
R1025 B.n930 B.n17 163.367
R1026 B.n930 B.n929 163.367
R1027 B.n929 B.n928 163.367
R1028 B.n928 B.n19 163.367
R1029 B.n924 B.n19 163.367
R1030 B.n924 B.n923 163.367
R1031 B.n923 B.n922 163.367
R1032 B.n922 B.n21 163.367
R1033 B.n918 B.n21 163.367
R1034 B.n918 B.n917 163.367
R1035 B.n917 B.n916 163.367
R1036 B.n916 B.n23 163.367
R1037 B.n912 B.n23 163.367
R1038 B.n912 B.n911 163.367
R1039 B.n911 B.n910 163.367
R1040 B.n910 B.n25 163.367
R1041 B.n906 B.n25 163.367
R1042 B.n906 B.n905 163.367
R1043 B.n905 B.n904 163.367
R1044 B.n904 B.n27 163.367
R1045 B.n900 B.n27 163.367
R1046 B.n900 B.n899 163.367
R1047 B.n899 B.n898 163.367
R1048 B.n898 B.n29 163.367
R1049 B.n894 B.n29 163.367
R1050 B.n894 B.n893 163.367
R1051 B.n893 B.n892 163.367
R1052 B.n892 B.n31 163.367
R1053 B.n888 B.n31 163.367
R1054 B.n888 B.n887 163.367
R1055 B.n887 B.n886 163.367
R1056 B.n886 B.n33 163.367
R1057 B.n882 B.n33 163.367
R1058 B.n882 B.n881 163.367
R1059 B.n881 B.n880 163.367
R1060 B.n880 B.n35 163.367
R1061 B.n876 B.n35 163.367
R1062 B.n876 B.n875 163.367
R1063 B.n875 B.n874 163.367
R1064 B.n874 B.n37 163.367
R1065 B.n870 B.n37 163.367
R1066 B.n870 B.n869 163.367
R1067 B.n869 B.n868 163.367
R1068 B.n868 B.n39 163.367
R1069 B.n365 B.n364 163.367
R1070 B.n366 B.n365 163.367
R1071 B.n366 B.n213 163.367
R1072 B.n370 B.n213 163.367
R1073 B.n371 B.n370 163.367
R1074 B.n372 B.n371 163.367
R1075 B.n372 B.n211 163.367
R1076 B.n376 B.n211 163.367
R1077 B.n377 B.n376 163.367
R1078 B.n378 B.n377 163.367
R1079 B.n378 B.n209 163.367
R1080 B.n382 B.n209 163.367
R1081 B.n383 B.n382 163.367
R1082 B.n384 B.n383 163.367
R1083 B.n384 B.n207 163.367
R1084 B.n388 B.n207 163.367
R1085 B.n389 B.n388 163.367
R1086 B.n390 B.n389 163.367
R1087 B.n390 B.n205 163.367
R1088 B.n394 B.n205 163.367
R1089 B.n395 B.n394 163.367
R1090 B.n396 B.n395 163.367
R1091 B.n396 B.n203 163.367
R1092 B.n400 B.n203 163.367
R1093 B.n401 B.n400 163.367
R1094 B.n402 B.n401 163.367
R1095 B.n402 B.n201 163.367
R1096 B.n406 B.n201 163.367
R1097 B.n407 B.n406 163.367
R1098 B.n408 B.n407 163.367
R1099 B.n408 B.n199 163.367
R1100 B.n412 B.n199 163.367
R1101 B.n413 B.n412 163.367
R1102 B.n414 B.n413 163.367
R1103 B.n414 B.n197 163.367
R1104 B.n418 B.n197 163.367
R1105 B.n419 B.n418 163.367
R1106 B.n420 B.n419 163.367
R1107 B.n420 B.n195 163.367
R1108 B.n424 B.n195 163.367
R1109 B.n425 B.n424 163.367
R1110 B.n425 B.n191 163.367
R1111 B.n429 B.n191 163.367
R1112 B.n430 B.n429 163.367
R1113 B.n431 B.n430 163.367
R1114 B.n431 B.n189 163.367
R1115 B.n435 B.n189 163.367
R1116 B.n436 B.n435 163.367
R1117 B.n437 B.n436 163.367
R1118 B.n437 B.n185 163.367
R1119 B.n442 B.n185 163.367
R1120 B.n443 B.n442 163.367
R1121 B.n444 B.n443 163.367
R1122 B.n444 B.n183 163.367
R1123 B.n448 B.n183 163.367
R1124 B.n449 B.n448 163.367
R1125 B.n450 B.n449 163.367
R1126 B.n450 B.n181 163.367
R1127 B.n454 B.n181 163.367
R1128 B.n455 B.n454 163.367
R1129 B.n456 B.n455 163.367
R1130 B.n456 B.n179 163.367
R1131 B.n460 B.n179 163.367
R1132 B.n461 B.n460 163.367
R1133 B.n462 B.n461 163.367
R1134 B.n462 B.n177 163.367
R1135 B.n466 B.n177 163.367
R1136 B.n467 B.n466 163.367
R1137 B.n468 B.n467 163.367
R1138 B.n468 B.n175 163.367
R1139 B.n472 B.n175 163.367
R1140 B.n473 B.n472 163.367
R1141 B.n474 B.n473 163.367
R1142 B.n474 B.n173 163.367
R1143 B.n478 B.n173 163.367
R1144 B.n479 B.n478 163.367
R1145 B.n480 B.n479 163.367
R1146 B.n480 B.n171 163.367
R1147 B.n484 B.n171 163.367
R1148 B.n485 B.n484 163.367
R1149 B.n486 B.n485 163.367
R1150 B.n486 B.n169 163.367
R1151 B.n490 B.n169 163.367
R1152 B.n491 B.n490 163.367
R1153 B.n492 B.n491 163.367
R1154 B.n492 B.n167 163.367
R1155 B.n496 B.n167 163.367
R1156 B.n497 B.n496 163.367
R1157 B.n498 B.n497 163.367
R1158 B.n498 B.n165 163.367
R1159 B.n503 B.n502 163.367
R1160 B.n504 B.n503 163.367
R1161 B.n504 B.n163 163.367
R1162 B.n508 B.n163 163.367
R1163 B.n509 B.n508 163.367
R1164 B.n510 B.n509 163.367
R1165 B.n510 B.n161 163.367
R1166 B.n514 B.n161 163.367
R1167 B.n515 B.n514 163.367
R1168 B.n516 B.n515 163.367
R1169 B.n516 B.n159 163.367
R1170 B.n520 B.n159 163.367
R1171 B.n521 B.n520 163.367
R1172 B.n522 B.n521 163.367
R1173 B.n522 B.n157 163.367
R1174 B.n526 B.n157 163.367
R1175 B.n527 B.n526 163.367
R1176 B.n528 B.n527 163.367
R1177 B.n528 B.n155 163.367
R1178 B.n532 B.n155 163.367
R1179 B.n533 B.n532 163.367
R1180 B.n534 B.n533 163.367
R1181 B.n534 B.n153 163.367
R1182 B.n538 B.n153 163.367
R1183 B.n539 B.n538 163.367
R1184 B.n540 B.n539 163.367
R1185 B.n540 B.n151 163.367
R1186 B.n544 B.n151 163.367
R1187 B.n545 B.n544 163.367
R1188 B.n546 B.n545 163.367
R1189 B.n546 B.n149 163.367
R1190 B.n550 B.n149 163.367
R1191 B.n551 B.n550 163.367
R1192 B.n552 B.n551 163.367
R1193 B.n552 B.n147 163.367
R1194 B.n556 B.n147 163.367
R1195 B.n557 B.n556 163.367
R1196 B.n558 B.n557 163.367
R1197 B.n558 B.n145 163.367
R1198 B.n562 B.n145 163.367
R1199 B.n563 B.n562 163.367
R1200 B.n564 B.n563 163.367
R1201 B.n564 B.n143 163.367
R1202 B.n568 B.n143 163.367
R1203 B.n569 B.n568 163.367
R1204 B.n570 B.n569 163.367
R1205 B.n570 B.n141 163.367
R1206 B.n574 B.n141 163.367
R1207 B.n575 B.n574 163.367
R1208 B.n576 B.n575 163.367
R1209 B.n576 B.n139 163.367
R1210 B.n580 B.n139 163.367
R1211 B.n581 B.n580 163.367
R1212 B.n582 B.n581 163.367
R1213 B.n582 B.n137 163.367
R1214 B.n586 B.n137 163.367
R1215 B.n587 B.n586 163.367
R1216 B.n588 B.n587 163.367
R1217 B.n588 B.n135 163.367
R1218 B.n592 B.n135 163.367
R1219 B.n593 B.n592 163.367
R1220 B.n594 B.n593 163.367
R1221 B.n594 B.n133 163.367
R1222 B.n598 B.n133 163.367
R1223 B.n599 B.n598 163.367
R1224 B.n600 B.n599 163.367
R1225 B.n600 B.n131 163.367
R1226 B.n604 B.n131 163.367
R1227 B.n605 B.n604 163.367
R1228 B.n606 B.n605 163.367
R1229 B.n606 B.n129 163.367
R1230 B.n610 B.n129 163.367
R1231 B.n611 B.n610 163.367
R1232 B.n612 B.n611 163.367
R1233 B.n612 B.n127 163.367
R1234 B.n616 B.n127 163.367
R1235 B.n617 B.n616 163.367
R1236 B.n618 B.n617 163.367
R1237 B.n618 B.n125 163.367
R1238 B.n622 B.n125 163.367
R1239 B.n623 B.n622 163.367
R1240 B.n624 B.n623 163.367
R1241 B.n624 B.n123 163.367
R1242 B.n628 B.n123 163.367
R1243 B.n629 B.n628 163.367
R1244 B.n630 B.n629 163.367
R1245 B.n630 B.n121 163.367
R1246 B.n634 B.n121 163.367
R1247 B.n635 B.n634 163.367
R1248 B.n636 B.n635 163.367
R1249 B.n636 B.n119 163.367
R1250 B.n640 B.n119 163.367
R1251 B.n641 B.n640 163.367
R1252 B.n642 B.n641 163.367
R1253 B.n642 B.n117 163.367
R1254 B.n646 B.n117 163.367
R1255 B.n647 B.n646 163.367
R1256 B.n648 B.n647 163.367
R1257 B.n648 B.n115 163.367
R1258 B.n652 B.n115 163.367
R1259 B.n653 B.n652 163.367
R1260 B.n654 B.n653 163.367
R1261 B.n654 B.n113 163.367
R1262 B.n658 B.n113 163.367
R1263 B.n659 B.n658 163.367
R1264 B.n660 B.n659 163.367
R1265 B.n660 B.n111 163.367
R1266 B.n664 B.n111 163.367
R1267 B.n665 B.n664 163.367
R1268 B.n666 B.n665 163.367
R1269 B.n666 B.n109 163.367
R1270 B.n670 B.n109 163.367
R1271 B.n671 B.n670 163.367
R1272 B.n672 B.n671 163.367
R1273 B.n672 B.n107 163.367
R1274 B.n676 B.n107 163.367
R1275 B.n677 B.n676 163.367
R1276 B.n678 B.n677 163.367
R1277 B.n678 B.n105 163.367
R1278 B.n682 B.n105 163.367
R1279 B.n683 B.n682 163.367
R1280 B.n684 B.n683 163.367
R1281 B.n684 B.n103 163.367
R1282 B.n688 B.n103 163.367
R1283 B.n689 B.n688 163.367
R1284 B.n690 B.n689 163.367
R1285 B.n690 B.n101 163.367
R1286 B.n694 B.n101 163.367
R1287 B.n695 B.n694 163.367
R1288 B.n696 B.n695 163.367
R1289 B.n696 B.n99 163.367
R1290 B.n700 B.n99 163.367
R1291 B.n701 B.n700 163.367
R1292 B.n702 B.n701 163.367
R1293 B.n702 B.n97 163.367
R1294 B.n706 B.n97 163.367
R1295 B.n707 B.n706 163.367
R1296 B.n708 B.n707 163.367
R1297 B.n708 B.n95 163.367
R1298 B.n712 B.n95 163.367
R1299 B.n713 B.n712 163.367
R1300 B.n714 B.n713 163.367
R1301 B.n714 B.n93 163.367
R1302 B.n718 B.n93 163.367
R1303 B.n719 B.n718 163.367
R1304 B.n720 B.n719 163.367
R1305 B.n720 B.n91 163.367
R1306 B.n724 B.n91 163.367
R1307 B.n725 B.n724 163.367
R1308 B.n726 B.n725 163.367
R1309 B.n864 B.n863 163.367
R1310 B.n863 B.n862 163.367
R1311 B.n862 B.n41 163.367
R1312 B.n858 B.n41 163.367
R1313 B.n858 B.n857 163.367
R1314 B.n857 B.n856 163.367
R1315 B.n856 B.n43 163.367
R1316 B.n852 B.n43 163.367
R1317 B.n852 B.n851 163.367
R1318 B.n851 B.n850 163.367
R1319 B.n850 B.n45 163.367
R1320 B.n846 B.n45 163.367
R1321 B.n846 B.n845 163.367
R1322 B.n845 B.n844 163.367
R1323 B.n844 B.n47 163.367
R1324 B.n840 B.n47 163.367
R1325 B.n840 B.n839 163.367
R1326 B.n839 B.n838 163.367
R1327 B.n838 B.n49 163.367
R1328 B.n834 B.n49 163.367
R1329 B.n834 B.n833 163.367
R1330 B.n833 B.n832 163.367
R1331 B.n832 B.n51 163.367
R1332 B.n828 B.n51 163.367
R1333 B.n828 B.n827 163.367
R1334 B.n827 B.n826 163.367
R1335 B.n826 B.n53 163.367
R1336 B.n822 B.n53 163.367
R1337 B.n822 B.n821 163.367
R1338 B.n821 B.n820 163.367
R1339 B.n820 B.n55 163.367
R1340 B.n816 B.n55 163.367
R1341 B.n816 B.n815 163.367
R1342 B.n815 B.n814 163.367
R1343 B.n814 B.n57 163.367
R1344 B.n810 B.n57 163.367
R1345 B.n810 B.n809 163.367
R1346 B.n809 B.n808 163.367
R1347 B.n808 B.n59 163.367
R1348 B.n804 B.n59 163.367
R1349 B.n804 B.n803 163.367
R1350 B.n803 B.n63 163.367
R1351 B.n799 B.n63 163.367
R1352 B.n799 B.n798 163.367
R1353 B.n798 B.n797 163.367
R1354 B.n797 B.n65 163.367
R1355 B.n793 B.n65 163.367
R1356 B.n793 B.n792 163.367
R1357 B.n792 B.n791 163.367
R1358 B.n791 B.n67 163.367
R1359 B.n786 B.n67 163.367
R1360 B.n786 B.n785 163.367
R1361 B.n785 B.n784 163.367
R1362 B.n784 B.n71 163.367
R1363 B.n780 B.n71 163.367
R1364 B.n780 B.n779 163.367
R1365 B.n779 B.n778 163.367
R1366 B.n778 B.n73 163.367
R1367 B.n774 B.n73 163.367
R1368 B.n774 B.n773 163.367
R1369 B.n773 B.n772 163.367
R1370 B.n772 B.n75 163.367
R1371 B.n768 B.n75 163.367
R1372 B.n768 B.n767 163.367
R1373 B.n767 B.n766 163.367
R1374 B.n766 B.n77 163.367
R1375 B.n762 B.n77 163.367
R1376 B.n762 B.n761 163.367
R1377 B.n761 B.n760 163.367
R1378 B.n760 B.n79 163.367
R1379 B.n756 B.n79 163.367
R1380 B.n756 B.n755 163.367
R1381 B.n755 B.n754 163.367
R1382 B.n754 B.n81 163.367
R1383 B.n750 B.n81 163.367
R1384 B.n750 B.n749 163.367
R1385 B.n749 B.n748 163.367
R1386 B.n748 B.n83 163.367
R1387 B.n744 B.n83 163.367
R1388 B.n744 B.n743 163.367
R1389 B.n743 B.n742 163.367
R1390 B.n742 B.n85 163.367
R1391 B.n738 B.n85 163.367
R1392 B.n738 B.n737 163.367
R1393 B.n737 B.n736 163.367
R1394 B.n736 B.n87 163.367
R1395 B.n732 B.n87 163.367
R1396 B.n732 B.n731 163.367
R1397 B.n731 B.n730 163.367
R1398 B.n730 B.n89 163.367
R1399 B.n187 B.t10 111.233
R1400 B.n69 B.t2 111.233
R1401 B.n193 B.t4 111.219
R1402 B.n61 B.t8 111.219
R1403 B.n187 B.n186 73.3096
R1404 B.n193 B.n192 73.3096
R1405 B.n61 B.n60 73.3096
R1406 B.n69 B.n68 73.3096
R1407 B.n439 B.n187 59.5399
R1408 B.n194 B.n193 59.5399
R1409 B.n62 B.n61 59.5399
R1410 B.n789 B.n69 59.5399
R1411 B.n866 B.n865 32.9371
R1412 B.n728 B.n727 32.9371
R1413 B.n501 B.n500 32.9371
R1414 B.n363 B.n362 32.9371
R1415 B B.n979 18.0485
R1416 B.n865 B.n40 10.6151
R1417 B.n861 B.n40 10.6151
R1418 B.n861 B.n860 10.6151
R1419 B.n860 B.n859 10.6151
R1420 B.n859 B.n42 10.6151
R1421 B.n855 B.n42 10.6151
R1422 B.n855 B.n854 10.6151
R1423 B.n854 B.n853 10.6151
R1424 B.n853 B.n44 10.6151
R1425 B.n849 B.n44 10.6151
R1426 B.n849 B.n848 10.6151
R1427 B.n848 B.n847 10.6151
R1428 B.n847 B.n46 10.6151
R1429 B.n843 B.n46 10.6151
R1430 B.n843 B.n842 10.6151
R1431 B.n842 B.n841 10.6151
R1432 B.n841 B.n48 10.6151
R1433 B.n837 B.n48 10.6151
R1434 B.n837 B.n836 10.6151
R1435 B.n836 B.n835 10.6151
R1436 B.n835 B.n50 10.6151
R1437 B.n831 B.n50 10.6151
R1438 B.n831 B.n830 10.6151
R1439 B.n830 B.n829 10.6151
R1440 B.n829 B.n52 10.6151
R1441 B.n825 B.n52 10.6151
R1442 B.n825 B.n824 10.6151
R1443 B.n824 B.n823 10.6151
R1444 B.n823 B.n54 10.6151
R1445 B.n819 B.n54 10.6151
R1446 B.n819 B.n818 10.6151
R1447 B.n818 B.n817 10.6151
R1448 B.n817 B.n56 10.6151
R1449 B.n813 B.n56 10.6151
R1450 B.n813 B.n812 10.6151
R1451 B.n812 B.n811 10.6151
R1452 B.n811 B.n58 10.6151
R1453 B.n807 B.n58 10.6151
R1454 B.n807 B.n806 10.6151
R1455 B.n806 B.n805 10.6151
R1456 B.n802 B.n801 10.6151
R1457 B.n801 B.n800 10.6151
R1458 B.n800 B.n64 10.6151
R1459 B.n796 B.n64 10.6151
R1460 B.n796 B.n795 10.6151
R1461 B.n795 B.n794 10.6151
R1462 B.n794 B.n66 10.6151
R1463 B.n790 B.n66 10.6151
R1464 B.n788 B.n787 10.6151
R1465 B.n787 B.n70 10.6151
R1466 B.n783 B.n70 10.6151
R1467 B.n783 B.n782 10.6151
R1468 B.n782 B.n781 10.6151
R1469 B.n781 B.n72 10.6151
R1470 B.n777 B.n72 10.6151
R1471 B.n777 B.n776 10.6151
R1472 B.n776 B.n775 10.6151
R1473 B.n775 B.n74 10.6151
R1474 B.n771 B.n74 10.6151
R1475 B.n771 B.n770 10.6151
R1476 B.n770 B.n769 10.6151
R1477 B.n769 B.n76 10.6151
R1478 B.n765 B.n76 10.6151
R1479 B.n765 B.n764 10.6151
R1480 B.n764 B.n763 10.6151
R1481 B.n763 B.n78 10.6151
R1482 B.n759 B.n78 10.6151
R1483 B.n759 B.n758 10.6151
R1484 B.n758 B.n757 10.6151
R1485 B.n757 B.n80 10.6151
R1486 B.n753 B.n80 10.6151
R1487 B.n753 B.n752 10.6151
R1488 B.n752 B.n751 10.6151
R1489 B.n751 B.n82 10.6151
R1490 B.n747 B.n82 10.6151
R1491 B.n747 B.n746 10.6151
R1492 B.n746 B.n745 10.6151
R1493 B.n745 B.n84 10.6151
R1494 B.n741 B.n84 10.6151
R1495 B.n741 B.n740 10.6151
R1496 B.n740 B.n739 10.6151
R1497 B.n739 B.n86 10.6151
R1498 B.n735 B.n86 10.6151
R1499 B.n735 B.n734 10.6151
R1500 B.n734 B.n733 10.6151
R1501 B.n733 B.n88 10.6151
R1502 B.n729 B.n88 10.6151
R1503 B.n729 B.n728 10.6151
R1504 B.n501 B.n164 10.6151
R1505 B.n505 B.n164 10.6151
R1506 B.n506 B.n505 10.6151
R1507 B.n507 B.n506 10.6151
R1508 B.n507 B.n162 10.6151
R1509 B.n511 B.n162 10.6151
R1510 B.n512 B.n511 10.6151
R1511 B.n513 B.n512 10.6151
R1512 B.n513 B.n160 10.6151
R1513 B.n517 B.n160 10.6151
R1514 B.n518 B.n517 10.6151
R1515 B.n519 B.n518 10.6151
R1516 B.n519 B.n158 10.6151
R1517 B.n523 B.n158 10.6151
R1518 B.n524 B.n523 10.6151
R1519 B.n525 B.n524 10.6151
R1520 B.n525 B.n156 10.6151
R1521 B.n529 B.n156 10.6151
R1522 B.n530 B.n529 10.6151
R1523 B.n531 B.n530 10.6151
R1524 B.n531 B.n154 10.6151
R1525 B.n535 B.n154 10.6151
R1526 B.n536 B.n535 10.6151
R1527 B.n537 B.n536 10.6151
R1528 B.n537 B.n152 10.6151
R1529 B.n541 B.n152 10.6151
R1530 B.n542 B.n541 10.6151
R1531 B.n543 B.n542 10.6151
R1532 B.n543 B.n150 10.6151
R1533 B.n547 B.n150 10.6151
R1534 B.n548 B.n547 10.6151
R1535 B.n549 B.n548 10.6151
R1536 B.n549 B.n148 10.6151
R1537 B.n553 B.n148 10.6151
R1538 B.n554 B.n553 10.6151
R1539 B.n555 B.n554 10.6151
R1540 B.n555 B.n146 10.6151
R1541 B.n559 B.n146 10.6151
R1542 B.n560 B.n559 10.6151
R1543 B.n561 B.n560 10.6151
R1544 B.n561 B.n144 10.6151
R1545 B.n565 B.n144 10.6151
R1546 B.n566 B.n565 10.6151
R1547 B.n567 B.n566 10.6151
R1548 B.n567 B.n142 10.6151
R1549 B.n571 B.n142 10.6151
R1550 B.n572 B.n571 10.6151
R1551 B.n573 B.n572 10.6151
R1552 B.n573 B.n140 10.6151
R1553 B.n577 B.n140 10.6151
R1554 B.n578 B.n577 10.6151
R1555 B.n579 B.n578 10.6151
R1556 B.n579 B.n138 10.6151
R1557 B.n583 B.n138 10.6151
R1558 B.n584 B.n583 10.6151
R1559 B.n585 B.n584 10.6151
R1560 B.n585 B.n136 10.6151
R1561 B.n589 B.n136 10.6151
R1562 B.n590 B.n589 10.6151
R1563 B.n591 B.n590 10.6151
R1564 B.n591 B.n134 10.6151
R1565 B.n595 B.n134 10.6151
R1566 B.n596 B.n595 10.6151
R1567 B.n597 B.n596 10.6151
R1568 B.n597 B.n132 10.6151
R1569 B.n601 B.n132 10.6151
R1570 B.n602 B.n601 10.6151
R1571 B.n603 B.n602 10.6151
R1572 B.n603 B.n130 10.6151
R1573 B.n607 B.n130 10.6151
R1574 B.n608 B.n607 10.6151
R1575 B.n609 B.n608 10.6151
R1576 B.n609 B.n128 10.6151
R1577 B.n613 B.n128 10.6151
R1578 B.n614 B.n613 10.6151
R1579 B.n615 B.n614 10.6151
R1580 B.n615 B.n126 10.6151
R1581 B.n619 B.n126 10.6151
R1582 B.n620 B.n619 10.6151
R1583 B.n621 B.n620 10.6151
R1584 B.n621 B.n124 10.6151
R1585 B.n625 B.n124 10.6151
R1586 B.n626 B.n625 10.6151
R1587 B.n627 B.n626 10.6151
R1588 B.n627 B.n122 10.6151
R1589 B.n631 B.n122 10.6151
R1590 B.n632 B.n631 10.6151
R1591 B.n633 B.n632 10.6151
R1592 B.n633 B.n120 10.6151
R1593 B.n637 B.n120 10.6151
R1594 B.n638 B.n637 10.6151
R1595 B.n639 B.n638 10.6151
R1596 B.n639 B.n118 10.6151
R1597 B.n643 B.n118 10.6151
R1598 B.n644 B.n643 10.6151
R1599 B.n645 B.n644 10.6151
R1600 B.n645 B.n116 10.6151
R1601 B.n649 B.n116 10.6151
R1602 B.n650 B.n649 10.6151
R1603 B.n651 B.n650 10.6151
R1604 B.n651 B.n114 10.6151
R1605 B.n655 B.n114 10.6151
R1606 B.n656 B.n655 10.6151
R1607 B.n657 B.n656 10.6151
R1608 B.n657 B.n112 10.6151
R1609 B.n661 B.n112 10.6151
R1610 B.n662 B.n661 10.6151
R1611 B.n663 B.n662 10.6151
R1612 B.n663 B.n110 10.6151
R1613 B.n667 B.n110 10.6151
R1614 B.n668 B.n667 10.6151
R1615 B.n669 B.n668 10.6151
R1616 B.n669 B.n108 10.6151
R1617 B.n673 B.n108 10.6151
R1618 B.n674 B.n673 10.6151
R1619 B.n675 B.n674 10.6151
R1620 B.n675 B.n106 10.6151
R1621 B.n679 B.n106 10.6151
R1622 B.n680 B.n679 10.6151
R1623 B.n681 B.n680 10.6151
R1624 B.n681 B.n104 10.6151
R1625 B.n685 B.n104 10.6151
R1626 B.n686 B.n685 10.6151
R1627 B.n687 B.n686 10.6151
R1628 B.n687 B.n102 10.6151
R1629 B.n691 B.n102 10.6151
R1630 B.n692 B.n691 10.6151
R1631 B.n693 B.n692 10.6151
R1632 B.n693 B.n100 10.6151
R1633 B.n697 B.n100 10.6151
R1634 B.n698 B.n697 10.6151
R1635 B.n699 B.n698 10.6151
R1636 B.n699 B.n98 10.6151
R1637 B.n703 B.n98 10.6151
R1638 B.n704 B.n703 10.6151
R1639 B.n705 B.n704 10.6151
R1640 B.n705 B.n96 10.6151
R1641 B.n709 B.n96 10.6151
R1642 B.n710 B.n709 10.6151
R1643 B.n711 B.n710 10.6151
R1644 B.n711 B.n94 10.6151
R1645 B.n715 B.n94 10.6151
R1646 B.n716 B.n715 10.6151
R1647 B.n717 B.n716 10.6151
R1648 B.n717 B.n92 10.6151
R1649 B.n721 B.n92 10.6151
R1650 B.n722 B.n721 10.6151
R1651 B.n723 B.n722 10.6151
R1652 B.n723 B.n90 10.6151
R1653 B.n727 B.n90 10.6151
R1654 B.n363 B.n214 10.6151
R1655 B.n367 B.n214 10.6151
R1656 B.n368 B.n367 10.6151
R1657 B.n369 B.n368 10.6151
R1658 B.n369 B.n212 10.6151
R1659 B.n373 B.n212 10.6151
R1660 B.n374 B.n373 10.6151
R1661 B.n375 B.n374 10.6151
R1662 B.n375 B.n210 10.6151
R1663 B.n379 B.n210 10.6151
R1664 B.n380 B.n379 10.6151
R1665 B.n381 B.n380 10.6151
R1666 B.n381 B.n208 10.6151
R1667 B.n385 B.n208 10.6151
R1668 B.n386 B.n385 10.6151
R1669 B.n387 B.n386 10.6151
R1670 B.n387 B.n206 10.6151
R1671 B.n391 B.n206 10.6151
R1672 B.n392 B.n391 10.6151
R1673 B.n393 B.n392 10.6151
R1674 B.n393 B.n204 10.6151
R1675 B.n397 B.n204 10.6151
R1676 B.n398 B.n397 10.6151
R1677 B.n399 B.n398 10.6151
R1678 B.n399 B.n202 10.6151
R1679 B.n403 B.n202 10.6151
R1680 B.n404 B.n403 10.6151
R1681 B.n405 B.n404 10.6151
R1682 B.n405 B.n200 10.6151
R1683 B.n409 B.n200 10.6151
R1684 B.n410 B.n409 10.6151
R1685 B.n411 B.n410 10.6151
R1686 B.n411 B.n198 10.6151
R1687 B.n415 B.n198 10.6151
R1688 B.n416 B.n415 10.6151
R1689 B.n417 B.n416 10.6151
R1690 B.n417 B.n196 10.6151
R1691 B.n421 B.n196 10.6151
R1692 B.n422 B.n421 10.6151
R1693 B.n423 B.n422 10.6151
R1694 B.n427 B.n426 10.6151
R1695 B.n428 B.n427 10.6151
R1696 B.n428 B.n190 10.6151
R1697 B.n432 B.n190 10.6151
R1698 B.n433 B.n432 10.6151
R1699 B.n434 B.n433 10.6151
R1700 B.n434 B.n188 10.6151
R1701 B.n438 B.n188 10.6151
R1702 B.n441 B.n440 10.6151
R1703 B.n441 B.n184 10.6151
R1704 B.n445 B.n184 10.6151
R1705 B.n446 B.n445 10.6151
R1706 B.n447 B.n446 10.6151
R1707 B.n447 B.n182 10.6151
R1708 B.n451 B.n182 10.6151
R1709 B.n452 B.n451 10.6151
R1710 B.n453 B.n452 10.6151
R1711 B.n453 B.n180 10.6151
R1712 B.n457 B.n180 10.6151
R1713 B.n458 B.n457 10.6151
R1714 B.n459 B.n458 10.6151
R1715 B.n459 B.n178 10.6151
R1716 B.n463 B.n178 10.6151
R1717 B.n464 B.n463 10.6151
R1718 B.n465 B.n464 10.6151
R1719 B.n465 B.n176 10.6151
R1720 B.n469 B.n176 10.6151
R1721 B.n470 B.n469 10.6151
R1722 B.n471 B.n470 10.6151
R1723 B.n471 B.n174 10.6151
R1724 B.n475 B.n174 10.6151
R1725 B.n476 B.n475 10.6151
R1726 B.n477 B.n476 10.6151
R1727 B.n477 B.n172 10.6151
R1728 B.n481 B.n172 10.6151
R1729 B.n482 B.n481 10.6151
R1730 B.n483 B.n482 10.6151
R1731 B.n483 B.n170 10.6151
R1732 B.n487 B.n170 10.6151
R1733 B.n488 B.n487 10.6151
R1734 B.n489 B.n488 10.6151
R1735 B.n489 B.n168 10.6151
R1736 B.n493 B.n168 10.6151
R1737 B.n494 B.n493 10.6151
R1738 B.n495 B.n494 10.6151
R1739 B.n495 B.n166 10.6151
R1740 B.n499 B.n166 10.6151
R1741 B.n500 B.n499 10.6151
R1742 B.n362 B.n361 10.6151
R1743 B.n361 B.n216 10.6151
R1744 B.n357 B.n216 10.6151
R1745 B.n357 B.n356 10.6151
R1746 B.n356 B.n355 10.6151
R1747 B.n355 B.n218 10.6151
R1748 B.n351 B.n218 10.6151
R1749 B.n351 B.n350 10.6151
R1750 B.n350 B.n349 10.6151
R1751 B.n349 B.n220 10.6151
R1752 B.n345 B.n220 10.6151
R1753 B.n345 B.n344 10.6151
R1754 B.n344 B.n343 10.6151
R1755 B.n343 B.n222 10.6151
R1756 B.n339 B.n222 10.6151
R1757 B.n339 B.n338 10.6151
R1758 B.n338 B.n337 10.6151
R1759 B.n337 B.n224 10.6151
R1760 B.n333 B.n224 10.6151
R1761 B.n333 B.n332 10.6151
R1762 B.n332 B.n331 10.6151
R1763 B.n331 B.n226 10.6151
R1764 B.n327 B.n226 10.6151
R1765 B.n327 B.n326 10.6151
R1766 B.n326 B.n325 10.6151
R1767 B.n325 B.n228 10.6151
R1768 B.n321 B.n228 10.6151
R1769 B.n321 B.n320 10.6151
R1770 B.n320 B.n319 10.6151
R1771 B.n319 B.n230 10.6151
R1772 B.n315 B.n230 10.6151
R1773 B.n315 B.n314 10.6151
R1774 B.n314 B.n313 10.6151
R1775 B.n313 B.n232 10.6151
R1776 B.n309 B.n232 10.6151
R1777 B.n309 B.n308 10.6151
R1778 B.n308 B.n307 10.6151
R1779 B.n307 B.n234 10.6151
R1780 B.n303 B.n234 10.6151
R1781 B.n303 B.n302 10.6151
R1782 B.n302 B.n301 10.6151
R1783 B.n301 B.n236 10.6151
R1784 B.n297 B.n236 10.6151
R1785 B.n297 B.n296 10.6151
R1786 B.n296 B.n295 10.6151
R1787 B.n295 B.n238 10.6151
R1788 B.n291 B.n238 10.6151
R1789 B.n291 B.n290 10.6151
R1790 B.n290 B.n289 10.6151
R1791 B.n289 B.n240 10.6151
R1792 B.n285 B.n240 10.6151
R1793 B.n285 B.n284 10.6151
R1794 B.n284 B.n283 10.6151
R1795 B.n283 B.n242 10.6151
R1796 B.n279 B.n242 10.6151
R1797 B.n279 B.n278 10.6151
R1798 B.n278 B.n277 10.6151
R1799 B.n277 B.n244 10.6151
R1800 B.n273 B.n244 10.6151
R1801 B.n273 B.n272 10.6151
R1802 B.n272 B.n271 10.6151
R1803 B.n271 B.n246 10.6151
R1804 B.n267 B.n246 10.6151
R1805 B.n267 B.n266 10.6151
R1806 B.n266 B.n265 10.6151
R1807 B.n265 B.n248 10.6151
R1808 B.n261 B.n248 10.6151
R1809 B.n261 B.n260 10.6151
R1810 B.n260 B.n259 10.6151
R1811 B.n259 B.n250 10.6151
R1812 B.n255 B.n250 10.6151
R1813 B.n255 B.n254 10.6151
R1814 B.n254 B.n253 10.6151
R1815 B.n253 B.n0 10.6151
R1816 B.n975 B.n1 10.6151
R1817 B.n975 B.n974 10.6151
R1818 B.n974 B.n973 10.6151
R1819 B.n973 B.n4 10.6151
R1820 B.n969 B.n4 10.6151
R1821 B.n969 B.n968 10.6151
R1822 B.n968 B.n967 10.6151
R1823 B.n967 B.n6 10.6151
R1824 B.n963 B.n6 10.6151
R1825 B.n963 B.n962 10.6151
R1826 B.n962 B.n961 10.6151
R1827 B.n961 B.n8 10.6151
R1828 B.n957 B.n8 10.6151
R1829 B.n957 B.n956 10.6151
R1830 B.n956 B.n955 10.6151
R1831 B.n955 B.n10 10.6151
R1832 B.n951 B.n10 10.6151
R1833 B.n951 B.n950 10.6151
R1834 B.n950 B.n949 10.6151
R1835 B.n949 B.n12 10.6151
R1836 B.n945 B.n12 10.6151
R1837 B.n945 B.n944 10.6151
R1838 B.n944 B.n943 10.6151
R1839 B.n943 B.n14 10.6151
R1840 B.n939 B.n14 10.6151
R1841 B.n939 B.n938 10.6151
R1842 B.n938 B.n937 10.6151
R1843 B.n937 B.n16 10.6151
R1844 B.n933 B.n16 10.6151
R1845 B.n933 B.n932 10.6151
R1846 B.n932 B.n931 10.6151
R1847 B.n931 B.n18 10.6151
R1848 B.n927 B.n18 10.6151
R1849 B.n927 B.n926 10.6151
R1850 B.n926 B.n925 10.6151
R1851 B.n925 B.n20 10.6151
R1852 B.n921 B.n20 10.6151
R1853 B.n921 B.n920 10.6151
R1854 B.n920 B.n919 10.6151
R1855 B.n919 B.n22 10.6151
R1856 B.n915 B.n22 10.6151
R1857 B.n915 B.n914 10.6151
R1858 B.n914 B.n913 10.6151
R1859 B.n913 B.n24 10.6151
R1860 B.n909 B.n24 10.6151
R1861 B.n909 B.n908 10.6151
R1862 B.n908 B.n907 10.6151
R1863 B.n907 B.n26 10.6151
R1864 B.n903 B.n26 10.6151
R1865 B.n903 B.n902 10.6151
R1866 B.n902 B.n901 10.6151
R1867 B.n901 B.n28 10.6151
R1868 B.n897 B.n28 10.6151
R1869 B.n897 B.n896 10.6151
R1870 B.n896 B.n895 10.6151
R1871 B.n895 B.n30 10.6151
R1872 B.n891 B.n30 10.6151
R1873 B.n891 B.n890 10.6151
R1874 B.n890 B.n889 10.6151
R1875 B.n889 B.n32 10.6151
R1876 B.n885 B.n32 10.6151
R1877 B.n885 B.n884 10.6151
R1878 B.n884 B.n883 10.6151
R1879 B.n883 B.n34 10.6151
R1880 B.n879 B.n34 10.6151
R1881 B.n879 B.n878 10.6151
R1882 B.n878 B.n877 10.6151
R1883 B.n877 B.n36 10.6151
R1884 B.n873 B.n36 10.6151
R1885 B.n873 B.n872 10.6151
R1886 B.n872 B.n871 10.6151
R1887 B.n871 B.n38 10.6151
R1888 B.n867 B.n38 10.6151
R1889 B.n867 B.n866 10.6151
R1890 B.n802 B.n62 6.5566
R1891 B.n790 B.n789 6.5566
R1892 B.n426 B.n194 6.5566
R1893 B.n439 B.n438 6.5566
R1894 B.n805 B.n62 4.05904
R1895 B.n789 B.n788 4.05904
R1896 B.n423 B.n194 4.05904
R1897 B.n440 B.n439 4.05904
R1898 B.n979 B.n0 2.81026
R1899 B.n979 B.n1 2.81026
C0 VDD1 B 2.79271f
C1 VDD2 VN 11.008f
C2 VP VN 9.607321f
C3 VDD2 w_n5506_n3322# 3.28293f
C4 VP w_n5506_n3322# 12.7448f
C5 VDD2 VTAIL 10.7349f
C6 VP VTAIL 12.039599f
C7 w_n5506_n3322# VN 12.0254f
C8 VDD2 B 2.94373f
C9 VTAIL VN 12.0254f
C10 VP B 2.71143f
C11 VTAIL w_n5506_n3322# 3.30114f
C12 B VN 1.4969f
C13 B w_n5506_n3322# 11.9113f
C14 B VTAIL 4.00465f
C15 VDD2 VDD1 2.72782f
C16 VP VDD1 11.5408f
C17 VDD1 VN 0.155265f
C18 VDD1 w_n5506_n3322# 3.0952f
C19 VDD1 VTAIL 10.6775f
C20 VP VDD2 0.69198f
C21 VDD2 VSUBS 2.47976f
C22 VDD1 VSUBS 2.305332f
C23 VTAIL VSUBS 1.497694f
C24 VN VSUBS 9.10572f
C25 VP VSUBS 5.319186f
C26 B VSUBS 6.401008f
C27 w_n5506_n3322# VSUBS 0.225239p
C28 B.n0 VSUBS 0.005685f
C29 B.n1 VSUBS 0.005685f
C30 B.n2 VSUBS 0.008991f
C31 B.n3 VSUBS 0.008991f
C32 B.n4 VSUBS 0.008991f
C33 B.n5 VSUBS 0.008991f
C34 B.n6 VSUBS 0.008991f
C35 B.n7 VSUBS 0.008991f
C36 B.n8 VSUBS 0.008991f
C37 B.n9 VSUBS 0.008991f
C38 B.n10 VSUBS 0.008991f
C39 B.n11 VSUBS 0.008991f
C40 B.n12 VSUBS 0.008991f
C41 B.n13 VSUBS 0.008991f
C42 B.n14 VSUBS 0.008991f
C43 B.n15 VSUBS 0.008991f
C44 B.n16 VSUBS 0.008991f
C45 B.n17 VSUBS 0.008991f
C46 B.n18 VSUBS 0.008991f
C47 B.n19 VSUBS 0.008991f
C48 B.n20 VSUBS 0.008991f
C49 B.n21 VSUBS 0.008991f
C50 B.n22 VSUBS 0.008991f
C51 B.n23 VSUBS 0.008991f
C52 B.n24 VSUBS 0.008991f
C53 B.n25 VSUBS 0.008991f
C54 B.n26 VSUBS 0.008991f
C55 B.n27 VSUBS 0.008991f
C56 B.n28 VSUBS 0.008991f
C57 B.n29 VSUBS 0.008991f
C58 B.n30 VSUBS 0.008991f
C59 B.n31 VSUBS 0.008991f
C60 B.n32 VSUBS 0.008991f
C61 B.n33 VSUBS 0.008991f
C62 B.n34 VSUBS 0.008991f
C63 B.n35 VSUBS 0.008991f
C64 B.n36 VSUBS 0.008991f
C65 B.n37 VSUBS 0.008991f
C66 B.n38 VSUBS 0.008991f
C67 B.n39 VSUBS 0.021014f
C68 B.n40 VSUBS 0.008991f
C69 B.n41 VSUBS 0.008991f
C70 B.n42 VSUBS 0.008991f
C71 B.n43 VSUBS 0.008991f
C72 B.n44 VSUBS 0.008991f
C73 B.n45 VSUBS 0.008991f
C74 B.n46 VSUBS 0.008991f
C75 B.n47 VSUBS 0.008991f
C76 B.n48 VSUBS 0.008991f
C77 B.n49 VSUBS 0.008991f
C78 B.n50 VSUBS 0.008991f
C79 B.n51 VSUBS 0.008991f
C80 B.n52 VSUBS 0.008991f
C81 B.n53 VSUBS 0.008991f
C82 B.n54 VSUBS 0.008991f
C83 B.n55 VSUBS 0.008991f
C84 B.n56 VSUBS 0.008991f
C85 B.n57 VSUBS 0.008991f
C86 B.n58 VSUBS 0.008991f
C87 B.n59 VSUBS 0.008991f
C88 B.t8 VSUBS 0.49164f
C89 B.t7 VSUBS 0.524967f
C90 B.t6 VSUBS 2.42139f
C91 B.n60 VSUBS 0.295448f
C92 B.n61 VSUBS 0.09671f
C93 B.n62 VSUBS 0.020831f
C94 B.n63 VSUBS 0.008991f
C95 B.n64 VSUBS 0.008991f
C96 B.n65 VSUBS 0.008991f
C97 B.n66 VSUBS 0.008991f
C98 B.n67 VSUBS 0.008991f
C99 B.t2 VSUBS 0.491631f
C100 B.t1 VSUBS 0.524959f
C101 B.t0 VSUBS 2.42139f
C102 B.n68 VSUBS 0.295456f
C103 B.n69 VSUBS 0.096719f
C104 B.n70 VSUBS 0.008991f
C105 B.n71 VSUBS 0.008991f
C106 B.n72 VSUBS 0.008991f
C107 B.n73 VSUBS 0.008991f
C108 B.n74 VSUBS 0.008991f
C109 B.n75 VSUBS 0.008991f
C110 B.n76 VSUBS 0.008991f
C111 B.n77 VSUBS 0.008991f
C112 B.n78 VSUBS 0.008991f
C113 B.n79 VSUBS 0.008991f
C114 B.n80 VSUBS 0.008991f
C115 B.n81 VSUBS 0.008991f
C116 B.n82 VSUBS 0.008991f
C117 B.n83 VSUBS 0.008991f
C118 B.n84 VSUBS 0.008991f
C119 B.n85 VSUBS 0.008991f
C120 B.n86 VSUBS 0.008991f
C121 B.n87 VSUBS 0.008991f
C122 B.n88 VSUBS 0.008991f
C123 B.n89 VSUBS 0.021297f
C124 B.n90 VSUBS 0.008991f
C125 B.n91 VSUBS 0.008991f
C126 B.n92 VSUBS 0.008991f
C127 B.n93 VSUBS 0.008991f
C128 B.n94 VSUBS 0.008991f
C129 B.n95 VSUBS 0.008991f
C130 B.n96 VSUBS 0.008991f
C131 B.n97 VSUBS 0.008991f
C132 B.n98 VSUBS 0.008991f
C133 B.n99 VSUBS 0.008991f
C134 B.n100 VSUBS 0.008991f
C135 B.n101 VSUBS 0.008991f
C136 B.n102 VSUBS 0.008991f
C137 B.n103 VSUBS 0.008991f
C138 B.n104 VSUBS 0.008991f
C139 B.n105 VSUBS 0.008991f
C140 B.n106 VSUBS 0.008991f
C141 B.n107 VSUBS 0.008991f
C142 B.n108 VSUBS 0.008991f
C143 B.n109 VSUBS 0.008991f
C144 B.n110 VSUBS 0.008991f
C145 B.n111 VSUBS 0.008991f
C146 B.n112 VSUBS 0.008991f
C147 B.n113 VSUBS 0.008991f
C148 B.n114 VSUBS 0.008991f
C149 B.n115 VSUBS 0.008991f
C150 B.n116 VSUBS 0.008991f
C151 B.n117 VSUBS 0.008991f
C152 B.n118 VSUBS 0.008991f
C153 B.n119 VSUBS 0.008991f
C154 B.n120 VSUBS 0.008991f
C155 B.n121 VSUBS 0.008991f
C156 B.n122 VSUBS 0.008991f
C157 B.n123 VSUBS 0.008991f
C158 B.n124 VSUBS 0.008991f
C159 B.n125 VSUBS 0.008991f
C160 B.n126 VSUBS 0.008991f
C161 B.n127 VSUBS 0.008991f
C162 B.n128 VSUBS 0.008991f
C163 B.n129 VSUBS 0.008991f
C164 B.n130 VSUBS 0.008991f
C165 B.n131 VSUBS 0.008991f
C166 B.n132 VSUBS 0.008991f
C167 B.n133 VSUBS 0.008991f
C168 B.n134 VSUBS 0.008991f
C169 B.n135 VSUBS 0.008991f
C170 B.n136 VSUBS 0.008991f
C171 B.n137 VSUBS 0.008991f
C172 B.n138 VSUBS 0.008991f
C173 B.n139 VSUBS 0.008991f
C174 B.n140 VSUBS 0.008991f
C175 B.n141 VSUBS 0.008991f
C176 B.n142 VSUBS 0.008991f
C177 B.n143 VSUBS 0.008991f
C178 B.n144 VSUBS 0.008991f
C179 B.n145 VSUBS 0.008991f
C180 B.n146 VSUBS 0.008991f
C181 B.n147 VSUBS 0.008991f
C182 B.n148 VSUBS 0.008991f
C183 B.n149 VSUBS 0.008991f
C184 B.n150 VSUBS 0.008991f
C185 B.n151 VSUBS 0.008991f
C186 B.n152 VSUBS 0.008991f
C187 B.n153 VSUBS 0.008991f
C188 B.n154 VSUBS 0.008991f
C189 B.n155 VSUBS 0.008991f
C190 B.n156 VSUBS 0.008991f
C191 B.n157 VSUBS 0.008991f
C192 B.n158 VSUBS 0.008991f
C193 B.n159 VSUBS 0.008991f
C194 B.n160 VSUBS 0.008991f
C195 B.n161 VSUBS 0.008991f
C196 B.n162 VSUBS 0.008991f
C197 B.n163 VSUBS 0.008991f
C198 B.n164 VSUBS 0.008991f
C199 B.n165 VSUBS 0.021297f
C200 B.n166 VSUBS 0.008991f
C201 B.n167 VSUBS 0.008991f
C202 B.n168 VSUBS 0.008991f
C203 B.n169 VSUBS 0.008991f
C204 B.n170 VSUBS 0.008991f
C205 B.n171 VSUBS 0.008991f
C206 B.n172 VSUBS 0.008991f
C207 B.n173 VSUBS 0.008991f
C208 B.n174 VSUBS 0.008991f
C209 B.n175 VSUBS 0.008991f
C210 B.n176 VSUBS 0.008991f
C211 B.n177 VSUBS 0.008991f
C212 B.n178 VSUBS 0.008991f
C213 B.n179 VSUBS 0.008991f
C214 B.n180 VSUBS 0.008991f
C215 B.n181 VSUBS 0.008991f
C216 B.n182 VSUBS 0.008991f
C217 B.n183 VSUBS 0.008991f
C218 B.n184 VSUBS 0.008991f
C219 B.n185 VSUBS 0.008991f
C220 B.t10 VSUBS 0.491631f
C221 B.t11 VSUBS 0.524959f
C222 B.t9 VSUBS 2.42139f
C223 B.n186 VSUBS 0.295456f
C224 B.n187 VSUBS 0.096719f
C225 B.n188 VSUBS 0.008991f
C226 B.n189 VSUBS 0.008991f
C227 B.n190 VSUBS 0.008991f
C228 B.n191 VSUBS 0.008991f
C229 B.t4 VSUBS 0.49164f
C230 B.t5 VSUBS 0.524967f
C231 B.t3 VSUBS 2.42139f
C232 B.n192 VSUBS 0.295448f
C233 B.n193 VSUBS 0.09671f
C234 B.n194 VSUBS 0.020831f
C235 B.n195 VSUBS 0.008991f
C236 B.n196 VSUBS 0.008991f
C237 B.n197 VSUBS 0.008991f
C238 B.n198 VSUBS 0.008991f
C239 B.n199 VSUBS 0.008991f
C240 B.n200 VSUBS 0.008991f
C241 B.n201 VSUBS 0.008991f
C242 B.n202 VSUBS 0.008991f
C243 B.n203 VSUBS 0.008991f
C244 B.n204 VSUBS 0.008991f
C245 B.n205 VSUBS 0.008991f
C246 B.n206 VSUBS 0.008991f
C247 B.n207 VSUBS 0.008991f
C248 B.n208 VSUBS 0.008991f
C249 B.n209 VSUBS 0.008991f
C250 B.n210 VSUBS 0.008991f
C251 B.n211 VSUBS 0.008991f
C252 B.n212 VSUBS 0.008991f
C253 B.n213 VSUBS 0.008991f
C254 B.n214 VSUBS 0.008991f
C255 B.n215 VSUBS 0.021014f
C256 B.n216 VSUBS 0.008991f
C257 B.n217 VSUBS 0.008991f
C258 B.n218 VSUBS 0.008991f
C259 B.n219 VSUBS 0.008991f
C260 B.n220 VSUBS 0.008991f
C261 B.n221 VSUBS 0.008991f
C262 B.n222 VSUBS 0.008991f
C263 B.n223 VSUBS 0.008991f
C264 B.n224 VSUBS 0.008991f
C265 B.n225 VSUBS 0.008991f
C266 B.n226 VSUBS 0.008991f
C267 B.n227 VSUBS 0.008991f
C268 B.n228 VSUBS 0.008991f
C269 B.n229 VSUBS 0.008991f
C270 B.n230 VSUBS 0.008991f
C271 B.n231 VSUBS 0.008991f
C272 B.n232 VSUBS 0.008991f
C273 B.n233 VSUBS 0.008991f
C274 B.n234 VSUBS 0.008991f
C275 B.n235 VSUBS 0.008991f
C276 B.n236 VSUBS 0.008991f
C277 B.n237 VSUBS 0.008991f
C278 B.n238 VSUBS 0.008991f
C279 B.n239 VSUBS 0.008991f
C280 B.n240 VSUBS 0.008991f
C281 B.n241 VSUBS 0.008991f
C282 B.n242 VSUBS 0.008991f
C283 B.n243 VSUBS 0.008991f
C284 B.n244 VSUBS 0.008991f
C285 B.n245 VSUBS 0.008991f
C286 B.n246 VSUBS 0.008991f
C287 B.n247 VSUBS 0.008991f
C288 B.n248 VSUBS 0.008991f
C289 B.n249 VSUBS 0.008991f
C290 B.n250 VSUBS 0.008991f
C291 B.n251 VSUBS 0.008991f
C292 B.n252 VSUBS 0.008991f
C293 B.n253 VSUBS 0.008991f
C294 B.n254 VSUBS 0.008991f
C295 B.n255 VSUBS 0.008991f
C296 B.n256 VSUBS 0.008991f
C297 B.n257 VSUBS 0.008991f
C298 B.n258 VSUBS 0.008991f
C299 B.n259 VSUBS 0.008991f
C300 B.n260 VSUBS 0.008991f
C301 B.n261 VSUBS 0.008991f
C302 B.n262 VSUBS 0.008991f
C303 B.n263 VSUBS 0.008991f
C304 B.n264 VSUBS 0.008991f
C305 B.n265 VSUBS 0.008991f
C306 B.n266 VSUBS 0.008991f
C307 B.n267 VSUBS 0.008991f
C308 B.n268 VSUBS 0.008991f
C309 B.n269 VSUBS 0.008991f
C310 B.n270 VSUBS 0.008991f
C311 B.n271 VSUBS 0.008991f
C312 B.n272 VSUBS 0.008991f
C313 B.n273 VSUBS 0.008991f
C314 B.n274 VSUBS 0.008991f
C315 B.n275 VSUBS 0.008991f
C316 B.n276 VSUBS 0.008991f
C317 B.n277 VSUBS 0.008991f
C318 B.n278 VSUBS 0.008991f
C319 B.n279 VSUBS 0.008991f
C320 B.n280 VSUBS 0.008991f
C321 B.n281 VSUBS 0.008991f
C322 B.n282 VSUBS 0.008991f
C323 B.n283 VSUBS 0.008991f
C324 B.n284 VSUBS 0.008991f
C325 B.n285 VSUBS 0.008991f
C326 B.n286 VSUBS 0.008991f
C327 B.n287 VSUBS 0.008991f
C328 B.n288 VSUBS 0.008991f
C329 B.n289 VSUBS 0.008991f
C330 B.n290 VSUBS 0.008991f
C331 B.n291 VSUBS 0.008991f
C332 B.n292 VSUBS 0.008991f
C333 B.n293 VSUBS 0.008991f
C334 B.n294 VSUBS 0.008991f
C335 B.n295 VSUBS 0.008991f
C336 B.n296 VSUBS 0.008991f
C337 B.n297 VSUBS 0.008991f
C338 B.n298 VSUBS 0.008991f
C339 B.n299 VSUBS 0.008991f
C340 B.n300 VSUBS 0.008991f
C341 B.n301 VSUBS 0.008991f
C342 B.n302 VSUBS 0.008991f
C343 B.n303 VSUBS 0.008991f
C344 B.n304 VSUBS 0.008991f
C345 B.n305 VSUBS 0.008991f
C346 B.n306 VSUBS 0.008991f
C347 B.n307 VSUBS 0.008991f
C348 B.n308 VSUBS 0.008991f
C349 B.n309 VSUBS 0.008991f
C350 B.n310 VSUBS 0.008991f
C351 B.n311 VSUBS 0.008991f
C352 B.n312 VSUBS 0.008991f
C353 B.n313 VSUBS 0.008991f
C354 B.n314 VSUBS 0.008991f
C355 B.n315 VSUBS 0.008991f
C356 B.n316 VSUBS 0.008991f
C357 B.n317 VSUBS 0.008991f
C358 B.n318 VSUBS 0.008991f
C359 B.n319 VSUBS 0.008991f
C360 B.n320 VSUBS 0.008991f
C361 B.n321 VSUBS 0.008991f
C362 B.n322 VSUBS 0.008991f
C363 B.n323 VSUBS 0.008991f
C364 B.n324 VSUBS 0.008991f
C365 B.n325 VSUBS 0.008991f
C366 B.n326 VSUBS 0.008991f
C367 B.n327 VSUBS 0.008991f
C368 B.n328 VSUBS 0.008991f
C369 B.n329 VSUBS 0.008991f
C370 B.n330 VSUBS 0.008991f
C371 B.n331 VSUBS 0.008991f
C372 B.n332 VSUBS 0.008991f
C373 B.n333 VSUBS 0.008991f
C374 B.n334 VSUBS 0.008991f
C375 B.n335 VSUBS 0.008991f
C376 B.n336 VSUBS 0.008991f
C377 B.n337 VSUBS 0.008991f
C378 B.n338 VSUBS 0.008991f
C379 B.n339 VSUBS 0.008991f
C380 B.n340 VSUBS 0.008991f
C381 B.n341 VSUBS 0.008991f
C382 B.n342 VSUBS 0.008991f
C383 B.n343 VSUBS 0.008991f
C384 B.n344 VSUBS 0.008991f
C385 B.n345 VSUBS 0.008991f
C386 B.n346 VSUBS 0.008991f
C387 B.n347 VSUBS 0.008991f
C388 B.n348 VSUBS 0.008991f
C389 B.n349 VSUBS 0.008991f
C390 B.n350 VSUBS 0.008991f
C391 B.n351 VSUBS 0.008991f
C392 B.n352 VSUBS 0.008991f
C393 B.n353 VSUBS 0.008991f
C394 B.n354 VSUBS 0.008991f
C395 B.n355 VSUBS 0.008991f
C396 B.n356 VSUBS 0.008991f
C397 B.n357 VSUBS 0.008991f
C398 B.n358 VSUBS 0.008991f
C399 B.n359 VSUBS 0.008991f
C400 B.n360 VSUBS 0.008991f
C401 B.n361 VSUBS 0.008991f
C402 B.n362 VSUBS 0.021014f
C403 B.n363 VSUBS 0.021297f
C404 B.n364 VSUBS 0.021297f
C405 B.n365 VSUBS 0.008991f
C406 B.n366 VSUBS 0.008991f
C407 B.n367 VSUBS 0.008991f
C408 B.n368 VSUBS 0.008991f
C409 B.n369 VSUBS 0.008991f
C410 B.n370 VSUBS 0.008991f
C411 B.n371 VSUBS 0.008991f
C412 B.n372 VSUBS 0.008991f
C413 B.n373 VSUBS 0.008991f
C414 B.n374 VSUBS 0.008991f
C415 B.n375 VSUBS 0.008991f
C416 B.n376 VSUBS 0.008991f
C417 B.n377 VSUBS 0.008991f
C418 B.n378 VSUBS 0.008991f
C419 B.n379 VSUBS 0.008991f
C420 B.n380 VSUBS 0.008991f
C421 B.n381 VSUBS 0.008991f
C422 B.n382 VSUBS 0.008991f
C423 B.n383 VSUBS 0.008991f
C424 B.n384 VSUBS 0.008991f
C425 B.n385 VSUBS 0.008991f
C426 B.n386 VSUBS 0.008991f
C427 B.n387 VSUBS 0.008991f
C428 B.n388 VSUBS 0.008991f
C429 B.n389 VSUBS 0.008991f
C430 B.n390 VSUBS 0.008991f
C431 B.n391 VSUBS 0.008991f
C432 B.n392 VSUBS 0.008991f
C433 B.n393 VSUBS 0.008991f
C434 B.n394 VSUBS 0.008991f
C435 B.n395 VSUBS 0.008991f
C436 B.n396 VSUBS 0.008991f
C437 B.n397 VSUBS 0.008991f
C438 B.n398 VSUBS 0.008991f
C439 B.n399 VSUBS 0.008991f
C440 B.n400 VSUBS 0.008991f
C441 B.n401 VSUBS 0.008991f
C442 B.n402 VSUBS 0.008991f
C443 B.n403 VSUBS 0.008991f
C444 B.n404 VSUBS 0.008991f
C445 B.n405 VSUBS 0.008991f
C446 B.n406 VSUBS 0.008991f
C447 B.n407 VSUBS 0.008991f
C448 B.n408 VSUBS 0.008991f
C449 B.n409 VSUBS 0.008991f
C450 B.n410 VSUBS 0.008991f
C451 B.n411 VSUBS 0.008991f
C452 B.n412 VSUBS 0.008991f
C453 B.n413 VSUBS 0.008991f
C454 B.n414 VSUBS 0.008991f
C455 B.n415 VSUBS 0.008991f
C456 B.n416 VSUBS 0.008991f
C457 B.n417 VSUBS 0.008991f
C458 B.n418 VSUBS 0.008991f
C459 B.n419 VSUBS 0.008991f
C460 B.n420 VSUBS 0.008991f
C461 B.n421 VSUBS 0.008991f
C462 B.n422 VSUBS 0.008991f
C463 B.n423 VSUBS 0.006214f
C464 B.n424 VSUBS 0.008991f
C465 B.n425 VSUBS 0.008991f
C466 B.n426 VSUBS 0.007272f
C467 B.n427 VSUBS 0.008991f
C468 B.n428 VSUBS 0.008991f
C469 B.n429 VSUBS 0.008991f
C470 B.n430 VSUBS 0.008991f
C471 B.n431 VSUBS 0.008991f
C472 B.n432 VSUBS 0.008991f
C473 B.n433 VSUBS 0.008991f
C474 B.n434 VSUBS 0.008991f
C475 B.n435 VSUBS 0.008991f
C476 B.n436 VSUBS 0.008991f
C477 B.n437 VSUBS 0.008991f
C478 B.n438 VSUBS 0.007272f
C479 B.n439 VSUBS 0.020831f
C480 B.n440 VSUBS 0.006214f
C481 B.n441 VSUBS 0.008991f
C482 B.n442 VSUBS 0.008991f
C483 B.n443 VSUBS 0.008991f
C484 B.n444 VSUBS 0.008991f
C485 B.n445 VSUBS 0.008991f
C486 B.n446 VSUBS 0.008991f
C487 B.n447 VSUBS 0.008991f
C488 B.n448 VSUBS 0.008991f
C489 B.n449 VSUBS 0.008991f
C490 B.n450 VSUBS 0.008991f
C491 B.n451 VSUBS 0.008991f
C492 B.n452 VSUBS 0.008991f
C493 B.n453 VSUBS 0.008991f
C494 B.n454 VSUBS 0.008991f
C495 B.n455 VSUBS 0.008991f
C496 B.n456 VSUBS 0.008991f
C497 B.n457 VSUBS 0.008991f
C498 B.n458 VSUBS 0.008991f
C499 B.n459 VSUBS 0.008991f
C500 B.n460 VSUBS 0.008991f
C501 B.n461 VSUBS 0.008991f
C502 B.n462 VSUBS 0.008991f
C503 B.n463 VSUBS 0.008991f
C504 B.n464 VSUBS 0.008991f
C505 B.n465 VSUBS 0.008991f
C506 B.n466 VSUBS 0.008991f
C507 B.n467 VSUBS 0.008991f
C508 B.n468 VSUBS 0.008991f
C509 B.n469 VSUBS 0.008991f
C510 B.n470 VSUBS 0.008991f
C511 B.n471 VSUBS 0.008991f
C512 B.n472 VSUBS 0.008991f
C513 B.n473 VSUBS 0.008991f
C514 B.n474 VSUBS 0.008991f
C515 B.n475 VSUBS 0.008991f
C516 B.n476 VSUBS 0.008991f
C517 B.n477 VSUBS 0.008991f
C518 B.n478 VSUBS 0.008991f
C519 B.n479 VSUBS 0.008991f
C520 B.n480 VSUBS 0.008991f
C521 B.n481 VSUBS 0.008991f
C522 B.n482 VSUBS 0.008991f
C523 B.n483 VSUBS 0.008991f
C524 B.n484 VSUBS 0.008991f
C525 B.n485 VSUBS 0.008991f
C526 B.n486 VSUBS 0.008991f
C527 B.n487 VSUBS 0.008991f
C528 B.n488 VSUBS 0.008991f
C529 B.n489 VSUBS 0.008991f
C530 B.n490 VSUBS 0.008991f
C531 B.n491 VSUBS 0.008991f
C532 B.n492 VSUBS 0.008991f
C533 B.n493 VSUBS 0.008991f
C534 B.n494 VSUBS 0.008991f
C535 B.n495 VSUBS 0.008991f
C536 B.n496 VSUBS 0.008991f
C537 B.n497 VSUBS 0.008991f
C538 B.n498 VSUBS 0.008991f
C539 B.n499 VSUBS 0.008991f
C540 B.n500 VSUBS 0.021297f
C541 B.n501 VSUBS 0.021014f
C542 B.n502 VSUBS 0.021014f
C543 B.n503 VSUBS 0.008991f
C544 B.n504 VSUBS 0.008991f
C545 B.n505 VSUBS 0.008991f
C546 B.n506 VSUBS 0.008991f
C547 B.n507 VSUBS 0.008991f
C548 B.n508 VSUBS 0.008991f
C549 B.n509 VSUBS 0.008991f
C550 B.n510 VSUBS 0.008991f
C551 B.n511 VSUBS 0.008991f
C552 B.n512 VSUBS 0.008991f
C553 B.n513 VSUBS 0.008991f
C554 B.n514 VSUBS 0.008991f
C555 B.n515 VSUBS 0.008991f
C556 B.n516 VSUBS 0.008991f
C557 B.n517 VSUBS 0.008991f
C558 B.n518 VSUBS 0.008991f
C559 B.n519 VSUBS 0.008991f
C560 B.n520 VSUBS 0.008991f
C561 B.n521 VSUBS 0.008991f
C562 B.n522 VSUBS 0.008991f
C563 B.n523 VSUBS 0.008991f
C564 B.n524 VSUBS 0.008991f
C565 B.n525 VSUBS 0.008991f
C566 B.n526 VSUBS 0.008991f
C567 B.n527 VSUBS 0.008991f
C568 B.n528 VSUBS 0.008991f
C569 B.n529 VSUBS 0.008991f
C570 B.n530 VSUBS 0.008991f
C571 B.n531 VSUBS 0.008991f
C572 B.n532 VSUBS 0.008991f
C573 B.n533 VSUBS 0.008991f
C574 B.n534 VSUBS 0.008991f
C575 B.n535 VSUBS 0.008991f
C576 B.n536 VSUBS 0.008991f
C577 B.n537 VSUBS 0.008991f
C578 B.n538 VSUBS 0.008991f
C579 B.n539 VSUBS 0.008991f
C580 B.n540 VSUBS 0.008991f
C581 B.n541 VSUBS 0.008991f
C582 B.n542 VSUBS 0.008991f
C583 B.n543 VSUBS 0.008991f
C584 B.n544 VSUBS 0.008991f
C585 B.n545 VSUBS 0.008991f
C586 B.n546 VSUBS 0.008991f
C587 B.n547 VSUBS 0.008991f
C588 B.n548 VSUBS 0.008991f
C589 B.n549 VSUBS 0.008991f
C590 B.n550 VSUBS 0.008991f
C591 B.n551 VSUBS 0.008991f
C592 B.n552 VSUBS 0.008991f
C593 B.n553 VSUBS 0.008991f
C594 B.n554 VSUBS 0.008991f
C595 B.n555 VSUBS 0.008991f
C596 B.n556 VSUBS 0.008991f
C597 B.n557 VSUBS 0.008991f
C598 B.n558 VSUBS 0.008991f
C599 B.n559 VSUBS 0.008991f
C600 B.n560 VSUBS 0.008991f
C601 B.n561 VSUBS 0.008991f
C602 B.n562 VSUBS 0.008991f
C603 B.n563 VSUBS 0.008991f
C604 B.n564 VSUBS 0.008991f
C605 B.n565 VSUBS 0.008991f
C606 B.n566 VSUBS 0.008991f
C607 B.n567 VSUBS 0.008991f
C608 B.n568 VSUBS 0.008991f
C609 B.n569 VSUBS 0.008991f
C610 B.n570 VSUBS 0.008991f
C611 B.n571 VSUBS 0.008991f
C612 B.n572 VSUBS 0.008991f
C613 B.n573 VSUBS 0.008991f
C614 B.n574 VSUBS 0.008991f
C615 B.n575 VSUBS 0.008991f
C616 B.n576 VSUBS 0.008991f
C617 B.n577 VSUBS 0.008991f
C618 B.n578 VSUBS 0.008991f
C619 B.n579 VSUBS 0.008991f
C620 B.n580 VSUBS 0.008991f
C621 B.n581 VSUBS 0.008991f
C622 B.n582 VSUBS 0.008991f
C623 B.n583 VSUBS 0.008991f
C624 B.n584 VSUBS 0.008991f
C625 B.n585 VSUBS 0.008991f
C626 B.n586 VSUBS 0.008991f
C627 B.n587 VSUBS 0.008991f
C628 B.n588 VSUBS 0.008991f
C629 B.n589 VSUBS 0.008991f
C630 B.n590 VSUBS 0.008991f
C631 B.n591 VSUBS 0.008991f
C632 B.n592 VSUBS 0.008991f
C633 B.n593 VSUBS 0.008991f
C634 B.n594 VSUBS 0.008991f
C635 B.n595 VSUBS 0.008991f
C636 B.n596 VSUBS 0.008991f
C637 B.n597 VSUBS 0.008991f
C638 B.n598 VSUBS 0.008991f
C639 B.n599 VSUBS 0.008991f
C640 B.n600 VSUBS 0.008991f
C641 B.n601 VSUBS 0.008991f
C642 B.n602 VSUBS 0.008991f
C643 B.n603 VSUBS 0.008991f
C644 B.n604 VSUBS 0.008991f
C645 B.n605 VSUBS 0.008991f
C646 B.n606 VSUBS 0.008991f
C647 B.n607 VSUBS 0.008991f
C648 B.n608 VSUBS 0.008991f
C649 B.n609 VSUBS 0.008991f
C650 B.n610 VSUBS 0.008991f
C651 B.n611 VSUBS 0.008991f
C652 B.n612 VSUBS 0.008991f
C653 B.n613 VSUBS 0.008991f
C654 B.n614 VSUBS 0.008991f
C655 B.n615 VSUBS 0.008991f
C656 B.n616 VSUBS 0.008991f
C657 B.n617 VSUBS 0.008991f
C658 B.n618 VSUBS 0.008991f
C659 B.n619 VSUBS 0.008991f
C660 B.n620 VSUBS 0.008991f
C661 B.n621 VSUBS 0.008991f
C662 B.n622 VSUBS 0.008991f
C663 B.n623 VSUBS 0.008991f
C664 B.n624 VSUBS 0.008991f
C665 B.n625 VSUBS 0.008991f
C666 B.n626 VSUBS 0.008991f
C667 B.n627 VSUBS 0.008991f
C668 B.n628 VSUBS 0.008991f
C669 B.n629 VSUBS 0.008991f
C670 B.n630 VSUBS 0.008991f
C671 B.n631 VSUBS 0.008991f
C672 B.n632 VSUBS 0.008991f
C673 B.n633 VSUBS 0.008991f
C674 B.n634 VSUBS 0.008991f
C675 B.n635 VSUBS 0.008991f
C676 B.n636 VSUBS 0.008991f
C677 B.n637 VSUBS 0.008991f
C678 B.n638 VSUBS 0.008991f
C679 B.n639 VSUBS 0.008991f
C680 B.n640 VSUBS 0.008991f
C681 B.n641 VSUBS 0.008991f
C682 B.n642 VSUBS 0.008991f
C683 B.n643 VSUBS 0.008991f
C684 B.n644 VSUBS 0.008991f
C685 B.n645 VSUBS 0.008991f
C686 B.n646 VSUBS 0.008991f
C687 B.n647 VSUBS 0.008991f
C688 B.n648 VSUBS 0.008991f
C689 B.n649 VSUBS 0.008991f
C690 B.n650 VSUBS 0.008991f
C691 B.n651 VSUBS 0.008991f
C692 B.n652 VSUBS 0.008991f
C693 B.n653 VSUBS 0.008991f
C694 B.n654 VSUBS 0.008991f
C695 B.n655 VSUBS 0.008991f
C696 B.n656 VSUBS 0.008991f
C697 B.n657 VSUBS 0.008991f
C698 B.n658 VSUBS 0.008991f
C699 B.n659 VSUBS 0.008991f
C700 B.n660 VSUBS 0.008991f
C701 B.n661 VSUBS 0.008991f
C702 B.n662 VSUBS 0.008991f
C703 B.n663 VSUBS 0.008991f
C704 B.n664 VSUBS 0.008991f
C705 B.n665 VSUBS 0.008991f
C706 B.n666 VSUBS 0.008991f
C707 B.n667 VSUBS 0.008991f
C708 B.n668 VSUBS 0.008991f
C709 B.n669 VSUBS 0.008991f
C710 B.n670 VSUBS 0.008991f
C711 B.n671 VSUBS 0.008991f
C712 B.n672 VSUBS 0.008991f
C713 B.n673 VSUBS 0.008991f
C714 B.n674 VSUBS 0.008991f
C715 B.n675 VSUBS 0.008991f
C716 B.n676 VSUBS 0.008991f
C717 B.n677 VSUBS 0.008991f
C718 B.n678 VSUBS 0.008991f
C719 B.n679 VSUBS 0.008991f
C720 B.n680 VSUBS 0.008991f
C721 B.n681 VSUBS 0.008991f
C722 B.n682 VSUBS 0.008991f
C723 B.n683 VSUBS 0.008991f
C724 B.n684 VSUBS 0.008991f
C725 B.n685 VSUBS 0.008991f
C726 B.n686 VSUBS 0.008991f
C727 B.n687 VSUBS 0.008991f
C728 B.n688 VSUBS 0.008991f
C729 B.n689 VSUBS 0.008991f
C730 B.n690 VSUBS 0.008991f
C731 B.n691 VSUBS 0.008991f
C732 B.n692 VSUBS 0.008991f
C733 B.n693 VSUBS 0.008991f
C734 B.n694 VSUBS 0.008991f
C735 B.n695 VSUBS 0.008991f
C736 B.n696 VSUBS 0.008991f
C737 B.n697 VSUBS 0.008991f
C738 B.n698 VSUBS 0.008991f
C739 B.n699 VSUBS 0.008991f
C740 B.n700 VSUBS 0.008991f
C741 B.n701 VSUBS 0.008991f
C742 B.n702 VSUBS 0.008991f
C743 B.n703 VSUBS 0.008991f
C744 B.n704 VSUBS 0.008991f
C745 B.n705 VSUBS 0.008991f
C746 B.n706 VSUBS 0.008991f
C747 B.n707 VSUBS 0.008991f
C748 B.n708 VSUBS 0.008991f
C749 B.n709 VSUBS 0.008991f
C750 B.n710 VSUBS 0.008991f
C751 B.n711 VSUBS 0.008991f
C752 B.n712 VSUBS 0.008991f
C753 B.n713 VSUBS 0.008991f
C754 B.n714 VSUBS 0.008991f
C755 B.n715 VSUBS 0.008991f
C756 B.n716 VSUBS 0.008991f
C757 B.n717 VSUBS 0.008991f
C758 B.n718 VSUBS 0.008991f
C759 B.n719 VSUBS 0.008991f
C760 B.n720 VSUBS 0.008991f
C761 B.n721 VSUBS 0.008991f
C762 B.n722 VSUBS 0.008991f
C763 B.n723 VSUBS 0.008991f
C764 B.n724 VSUBS 0.008991f
C765 B.n725 VSUBS 0.008991f
C766 B.n726 VSUBS 0.021014f
C767 B.n727 VSUBS 0.022067f
C768 B.n728 VSUBS 0.020243f
C769 B.n729 VSUBS 0.008991f
C770 B.n730 VSUBS 0.008991f
C771 B.n731 VSUBS 0.008991f
C772 B.n732 VSUBS 0.008991f
C773 B.n733 VSUBS 0.008991f
C774 B.n734 VSUBS 0.008991f
C775 B.n735 VSUBS 0.008991f
C776 B.n736 VSUBS 0.008991f
C777 B.n737 VSUBS 0.008991f
C778 B.n738 VSUBS 0.008991f
C779 B.n739 VSUBS 0.008991f
C780 B.n740 VSUBS 0.008991f
C781 B.n741 VSUBS 0.008991f
C782 B.n742 VSUBS 0.008991f
C783 B.n743 VSUBS 0.008991f
C784 B.n744 VSUBS 0.008991f
C785 B.n745 VSUBS 0.008991f
C786 B.n746 VSUBS 0.008991f
C787 B.n747 VSUBS 0.008991f
C788 B.n748 VSUBS 0.008991f
C789 B.n749 VSUBS 0.008991f
C790 B.n750 VSUBS 0.008991f
C791 B.n751 VSUBS 0.008991f
C792 B.n752 VSUBS 0.008991f
C793 B.n753 VSUBS 0.008991f
C794 B.n754 VSUBS 0.008991f
C795 B.n755 VSUBS 0.008991f
C796 B.n756 VSUBS 0.008991f
C797 B.n757 VSUBS 0.008991f
C798 B.n758 VSUBS 0.008991f
C799 B.n759 VSUBS 0.008991f
C800 B.n760 VSUBS 0.008991f
C801 B.n761 VSUBS 0.008991f
C802 B.n762 VSUBS 0.008991f
C803 B.n763 VSUBS 0.008991f
C804 B.n764 VSUBS 0.008991f
C805 B.n765 VSUBS 0.008991f
C806 B.n766 VSUBS 0.008991f
C807 B.n767 VSUBS 0.008991f
C808 B.n768 VSUBS 0.008991f
C809 B.n769 VSUBS 0.008991f
C810 B.n770 VSUBS 0.008991f
C811 B.n771 VSUBS 0.008991f
C812 B.n772 VSUBS 0.008991f
C813 B.n773 VSUBS 0.008991f
C814 B.n774 VSUBS 0.008991f
C815 B.n775 VSUBS 0.008991f
C816 B.n776 VSUBS 0.008991f
C817 B.n777 VSUBS 0.008991f
C818 B.n778 VSUBS 0.008991f
C819 B.n779 VSUBS 0.008991f
C820 B.n780 VSUBS 0.008991f
C821 B.n781 VSUBS 0.008991f
C822 B.n782 VSUBS 0.008991f
C823 B.n783 VSUBS 0.008991f
C824 B.n784 VSUBS 0.008991f
C825 B.n785 VSUBS 0.008991f
C826 B.n786 VSUBS 0.008991f
C827 B.n787 VSUBS 0.008991f
C828 B.n788 VSUBS 0.006214f
C829 B.n789 VSUBS 0.020831f
C830 B.n790 VSUBS 0.007272f
C831 B.n791 VSUBS 0.008991f
C832 B.n792 VSUBS 0.008991f
C833 B.n793 VSUBS 0.008991f
C834 B.n794 VSUBS 0.008991f
C835 B.n795 VSUBS 0.008991f
C836 B.n796 VSUBS 0.008991f
C837 B.n797 VSUBS 0.008991f
C838 B.n798 VSUBS 0.008991f
C839 B.n799 VSUBS 0.008991f
C840 B.n800 VSUBS 0.008991f
C841 B.n801 VSUBS 0.008991f
C842 B.n802 VSUBS 0.007272f
C843 B.n803 VSUBS 0.008991f
C844 B.n804 VSUBS 0.008991f
C845 B.n805 VSUBS 0.006214f
C846 B.n806 VSUBS 0.008991f
C847 B.n807 VSUBS 0.008991f
C848 B.n808 VSUBS 0.008991f
C849 B.n809 VSUBS 0.008991f
C850 B.n810 VSUBS 0.008991f
C851 B.n811 VSUBS 0.008991f
C852 B.n812 VSUBS 0.008991f
C853 B.n813 VSUBS 0.008991f
C854 B.n814 VSUBS 0.008991f
C855 B.n815 VSUBS 0.008991f
C856 B.n816 VSUBS 0.008991f
C857 B.n817 VSUBS 0.008991f
C858 B.n818 VSUBS 0.008991f
C859 B.n819 VSUBS 0.008991f
C860 B.n820 VSUBS 0.008991f
C861 B.n821 VSUBS 0.008991f
C862 B.n822 VSUBS 0.008991f
C863 B.n823 VSUBS 0.008991f
C864 B.n824 VSUBS 0.008991f
C865 B.n825 VSUBS 0.008991f
C866 B.n826 VSUBS 0.008991f
C867 B.n827 VSUBS 0.008991f
C868 B.n828 VSUBS 0.008991f
C869 B.n829 VSUBS 0.008991f
C870 B.n830 VSUBS 0.008991f
C871 B.n831 VSUBS 0.008991f
C872 B.n832 VSUBS 0.008991f
C873 B.n833 VSUBS 0.008991f
C874 B.n834 VSUBS 0.008991f
C875 B.n835 VSUBS 0.008991f
C876 B.n836 VSUBS 0.008991f
C877 B.n837 VSUBS 0.008991f
C878 B.n838 VSUBS 0.008991f
C879 B.n839 VSUBS 0.008991f
C880 B.n840 VSUBS 0.008991f
C881 B.n841 VSUBS 0.008991f
C882 B.n842 VSUBS 0.008991f
C883 B.n843 VSUBS 0.008991f
C884 B.n844 VSUBS 0.008991f
C885 B.n845 VSUBS 0.008991f
C886 B.n846 VSUBS 0.008991f
C887 B.n847 VSUBS 0.008991f
C888 B.n848 VSUBS 0.008991f
C889 B.n849 VSUBS 0.008991f
C890 B.n850 VSUBS 0.008991f
C891 B.n851 VSUBS 0.008991f
C892 B.n852 VSUBS 0.008991f
C893 B.n853 VSUBS 0.008991f
C894 B.n854 VSUBS 0.008991f
C895 B.n855 VSUBS 0.008991f
C896 B.n856 VSUBS 0.008991f
C897 B.n857 VSUBS 0.008991f
C898 B.n858 VSUBS 0.008991f
C899 B.n859 VSUBS 0.008991f
C900 B.n860 VSUBS 0.008991f
C901 B.n861 VSUBS 0.008991f
C902 B.n862 VSUBS 0.008991f
C903 B.n863 VSUBS 0.008991f
C904 B.n864 VSUBS 0.021297f
C905 B.n865 VSUBS 0.021297f
C906 B.n866 VSUBS 0.021014f
C907 B.n867 VSUBS 0.008991f
C908 B.n868 VSUBS 0.008991f
C909 B.n869 VSUBS 0.008991f
C910 B.n870 VSUBS 0.008991f
C911 B.n871 VSUBS 0.008991f
C912 B.n872 VSUBS 0.008991f
C913 B.n873 VSUBS 0.008991f
C914 B.n874 VSUBS 0.008991f
C915 B.n875 VSUBS 0.008991f
C916 B.n876 VSUBS 0.008991f
C917 B.n877 VSUBS 0.008991f
C918 B.n878 VSUBS 0.008991f
C919 B.n879 VSUBS 0.008991f
C920 B.n880 VSUBS 0.008991f
C921 B.n881 VSUBS 0.008991f
C922 B.n882 VSUBS 0.008991f
C923 B.n883 VSUBS 0.008991f
C924 B.n884 VSUBS 0.008991f
C925 B.n885 VSUBS 0.008991f
C926 B.n886 VSUBS 0.008991f
C927 B.n887 VSUBS 0.008991f
C928 B.n888 VSUBS 0.008991f
C929 B.n889 VSUBS 0.008991f
C930 B.n890 VSUBS 0.008991f
C931 B.n891 VSUBS 0.008991f
C932 B.n892 VSUBS 0.008991f
C933 B.n893 VSUBS 0.008991f
C934 B.n894 VSUBS 0.008991f
C935 B.n895 VSUBS 0.008991f
C936 B.n896 VSUBS 0.008991f
C937 B.n897 VSUBS 0.008991f
C938 B.n898 VSUBS 0.008991f
C939 B.n899 VSUBS 0.008991f
C940 B.n900 VSUBS 0.008991f
C941 B.n901 VSUBS 0.008991f
C942 B.n902 VSUBS 0.008991f
C943 B.n903 VSUBS 0.008991f
C944 B.n904 VSUBS 0.008991f
C945 B.n905 VSUBS 0.008991f
C946 B.n906 VSUBS 0.008991f
C947 B.n907 VSUBS 0.008991f
C948 B.n908 VSUBS 0.008991f
C949 B.n909 VSUBS 0.008991f
C950 B.n910 VSUBS 0.008991f
C951 B.n911 VSUBS 0.008991f
C952 B.n912 VSUBS 0.008991f
C953 B.n913 VSUBS 0.008991f
C954 B.n914 VSUBS 0.008991f
C955 B.n915 VSUBS 0.008991f
C956 B.n916 VSUBS 0.008991f
C957 B.n917 VSUBS 0.008991f
C958 B.n918 VSUBS 0.008991f
C959 B.n919 VSUBS 0.008991f
C960 B.n920 VSUBS 0.008991f
C961 B.n921 VSUBS 0.008991f
C962 B.n922 VSUBS 0.008991f
C963 B.n923 VSUBS 0.008991f
C964 B.n924 VSUBS 0.008991f
C965 B.n925 VSUBS 0.008991f
C966 B.n926 VSUBS 0.008991f
C967 B.n927 VSUBS 0.008991f
C968 B.n928 VSUBS 0.008991f
C969 B.n929 VSUBS 0.008991f
C970 B.n930 VSUBS 0.008991f
C971 B.n931 VSUBS 0.008991f
C972 B.n932 VSUBS 0.008991f
C973 B.n933 VSUBS 0.008991f
C974 B.n934 VSUBS 0.008991f
C975 B.n935 VSUBS 0.008991f
C976 B.n936 VSUBS 0.008991f
C977 B.n937 VSUBS 0.008991f
C978 B.n938 VSUBS 0.008991f
C979 B.n939 VSUBS 0.008991f
C980 B.n940 VSUBS 0.008991f
C981 B.n941 VSUBS 0.008991f
C982 B.n942 VSUBS 0.008991f
C983 B.n943 VSUBS 0.008991f
C984 B.n944 VSUBS 0.008991f
C985 B.n945 VSUBS 0.008991f
C986 B.n946 VSUBS 0.008991f
C987 B.n947 VSUBS 0.008991f
C988 B.n948 VSUBS 0.008991f
C989 B.n949 VSUBS 0.008991f
C990 B.n950 VSUBS 0.008991f
C991 B.n951 VSUBS 0.008991f
C992 B.n952 VSUBS 0.008991f
C993 B.n953 VSUBS 0.008991f
C994 B.n954 VSUBS 0.008991f
C995 B.n955 VSUBS 0.008991f
C996 B.n956 VSUBS 0.008991f
C997 B.n957 VSUBS 0.008991f
C998 B.n958 VSUBS 0.008991f
C999 B.n959 VSUBS 0.008991f
C1000 B.n960 VSUBS 0.008991f
C1001 B.n961 VSUBS 0.008991f
C1002 B.n962 VSUBS 0.008991f
C1003 B.n963 VSUBS 0.008991f
C1004 B.n964 VSUBS 0.008991f
C1005 B.n965 VSUBS 0.008991f
C1006 B.n966 VSUBS 0.008991f
C1007 B.n967 VSUBS 0.008991f
C1008 B.n968 VSUBS 0.008991f
C1009 B.n969 VSUBS 0.008991f
C1010 B.n970 VSUBS 0.008991f
C1011 B.n971 VSUBS 0.008991f
C1012 B.n972 VSUBS 0.008991f
C1013 B.n973 VSUBS 0.008991f
C1014 B.n974 VSUBS 0.008991f
C1015 B.n975 VSUBS 0.008991f
C1016 B.n976 VSUBS 0.008991f
C1017 B.n977 VSUBS 0.008991f
C1018 B.n978 VSUBS 0.008991f
C1019 B.n979 VSUBS 0.020359f
C1020 VDD2.t1 VSUBS 2.96231f
C1021 VDD2.t9 VSUBS 0.287361f
C1022 VDD2.t3 VSUBS 0.287361f
C1023 VDD2.n0 VSUBS 2.23529f
C1024 VDD2.n1 VSUBS 1.9497f
C1025 VDD2.t2 VSUBS 0.287361f
C1026 VDD2.t8 VSUBS 0.287361f
C1027 VDD2.n2 VSUBS 2.2711f
C1028 VDD2.n3 VSUBS 4.43765f
C1029 VDD2.t5 VSUBS 2.92135f
C1030 VDD2.n4 VSUBS 4.58784f
C1031 VDD2.t0 VSUBS 0.287361f
C1032 VDD2.t6 VSUBS 0.287361f
C1033 VDD2.n5 VSUBS 2.2353f
C1034 VDD2.n6 VSUBS 0.988901f
C1035 VDD2.t7 VSUBS 0.287361f
C1036 VDD2.t4 VSUBS 0.287361f
C1037 VDD2.n7 VSUBS 2.27104f
C1038 VN.t1 VSUBS 2.7063f
C1039 VN.n0 VSUBS 1.052f
C1040 VN.n1 VSUBS 0.024475f
C1041 VN.n2 VSUBS 0.021874f
C1042 VN.n3 VSUBS 0.024475f
C1043 VN.t7 VSUBS 2.7063f
C1044 VN.n4 VSUBS 0.950912f
C1045 VN.n5 VSUBS 0.024475f
C1046 VN.n6 VSUBS 0.042899f
C1047 VN.n7 VSUBS 0.024475f
C1048 VN.n8 VSUBS 0.034354f
C1049 VN.n9 VSUBS 0.024475f
C1050 VN.n10 VSUBS 0.026729f
C1051 VN.n11 VSUBS 0.024475f
C1052 VN.n12 VSUBS 0.024446f
C1053 VN.t0 VSUBS 2.7063f
C1054 VN.n13 VSUBS 1.026f
C1055 VN.t8 VSUBS 3.0292f
C1056 VN.n14 VSUBS 0.976898f
C1057 VN.n15 VSUBS 0.29202f
C1058 VN.n16 VSUBS 0.024475f
C1059 VN.n17 VSUBS 0.045615f
C1060 VN.n18 VSUBS 0.045615f
C1061 VN.n19 VSUBS 0.042899f
C1062 VN.n20 VSUBS 0.024475f
C1063 VN.n21 VSUBS 0.024475f
C1064 VN.n22 VSUBS 0.024475f
C1065 VN.n23 VSUBS 0.047443f
C1066 VN.n24 VSUBS 0.045615f
C1067 VN.t6 VSUBS 2.7063f
C1068 VN.n25 VSUBS 0.950912f
C1069 VN.n26 VSUBS 0.034354f
C1070 VN.n27 VSUBS 0.024475f
C1071 VN.n28 VSUBS 0.024475f
C1072 VN.n29 VSUBS 0.024475f
C1073 VN.n30 VSUBS 0.045615f
C1074 VN.n31 VSUBS 0.047443f
C1075 VN.n32 VSUBS 0.026729f
C1076 VN.n33 VSUBS 0.024475f
C1077 VN.n34 VSUBS 0.024475f
C1078 VN.n35 VSUBS 0.024475f
C1079 VN.n36 VSUBS 0.045615f
C1080 VN.n37 VSUBS 0.045615f
C1081 VN.n38 VSUBS 0.024446f
C1082 VN.n39 VSUBS 0.024475f
C1083 VN.n40 VSUBS 0.024475f
C1084 VN.n41 VSUBS 0.044263f
C1085 VN.n42 VSUBS 0.045615f
C1086 VN.n43 VSUBS 0.045835f
C1087 VN.n44 VSUBS 0.024475f
C1088 VN.n45 VSUBS 0.024475f
C1089 VN.n46 VSUBS 0.024475f
C1090 VN.n47 VSUBS 0.049363f
C1091 VN.n48 VSUBS 0.045615f
C1092 VN.n49 VSUBS 0.037057f
C1093 VN.n50 VSUBS 0.039502f
C1094 VN.n51 VSUBS 0.060218f
C1095 VN.t4 VSUBS 2.7063f
C1096 VN.n52 VSUBS 1.052f
C1097 VN.n53 VSUBS 0.024475f
C1098 VN.n54 VSUBS 0.021874f
C1099 VN.n55 VSUBS 0.024475f
C1100 VN.t9 VSUBS 2.7063f
C1101 VN.n56 VSUBS 0.950912f
C1102 VN.n57 VSUBS 0.024475f
C1103 VN.n58 VSUBS 0.042899f
C1104 VN.n59 VSUBS 0.024475f
C1105 VN.n60 VSUBS 0.034354f
C1106 VN.n61 VSUBS 0.024475f
C1107 VN.t3 VSUBS 2.7063f
C1108 VN.n62 VSUBS 0.950912f
C1109 VN.n63 VSUBS 0.026729f
C1110 VN.n64 VSUBS 0.024475f
C1111 VN.n65 VSUBS 0.024446f
C1112 VN.t5 VSUBS 3.0292f
C1113 VN.t2 VSUBS 2.7063f
C1114 VN.n66 VSUBS 1.026f
C1115 VN.n67 VSUBS 0.976898f
C1116 VN.n68 VSUBS 0.29202f
C1117 VN.n69 VSUBS 0.024475f
C1118 VN.n70 VSUBS 0.045615f
C1119 VN.n71 VSUBS 0.045615f
C1120 VN.n72 VSUBS 0.042899f
C1121 VN.n73 VSUBS 0.024475f
C1122 VN.n74 VSUBS 0.024475f
C1123 VN.n75 VSUBS 0.024475f
C1124 VN.n76 VSUBS 0.047443f
C1125 VN.n77 VSUBS 0.045615f
C1126 VN.n78 VSUBS 0.034354f
C1127 VN.n79 VSUBS 0.024475f
C1128 VN.n80 VSUBS 0.024475f
C1129 VN.n81 VSUBS 0.024475f
C1130 VN.n82 VSUBS 0.045615f
C1131 VN.n83 VSUBS 0.047443f
C1132 VN.n84 VSUBS 0.026729f
C1133 VN.n85 VSUBS 0.024475f
C1134 VN.n86 VSUBS 0.024475f
C1135 VN.n87 VSUBS 0.024475f
C1136 VN.n88 VSUBS 0.045615f
C1137 VN.n89 VSUBS 0.045615f
C1138 VN.n90 VSUBS 0.024446f
C1139 VN.n91 VSUBS 0.024475f
C1140 VN.n92 VSUBS 0.024475f
C1141 VN.n93 VSUBS 0.044263f
C1142 VN.n94 VSUBS 0.045615f
C1143 VN.n95 VSUBS 0.045835f
C1144 VN.n96 VSUBS 0.024475f
C1145 VN.n97 VSUBS 0.024475f
C1146 VN.n98 VSUBS 0.024475f
C1147 VN.n99 VSUBS 0.049363f
C1148 VN.n100 VSUBS 0.045615f
C1149 VN.n101 VSUBS 0.037057f
C1150 VN.n102 VSUBS 0.039502f
C1151 VN.n103 VSUBS 1.71306f
C1152 VDD1.t3 VSUBS 2.9706f
C1153 VDD1.t8 VSUBS 0.288165f
C1154 VDD1.t2 VSUBS 0.288165f
C1155 VDD1.n0 VSUBS 2.24155f
C1156 VDD1.n1 VSUBS 1.96552f
C1157 VDD1.t9 VSUBS 2.9706f
C1158 VDD1.t1 VSUBS 0.288165f
C1159 VDD1.t4 VSUBS 0.288165f
C1160 VDD1.n2 VSUBS 2.24154f
C1161 VDD1.n3 VSUBS 1.95515f
C1162 VDD1.t6 VSUBS 0.288165f
C1163 VDD1.t0 VSUBS 0.288165f
C1164 VDD1.n4 VSUBS 2.27745f
C1165 VDD1.n5 VSUBS 4.6337f
C1166 VDD1.t5 VSUBS 0.288165f
C1167 VDD1.t7 VSUBS 0.288165f
C1168 VDD1.n6 VSUBS 2.24154f
C1169 VDD1.n7 VSUBS 4.67172f
C1170 VTAIL.t9 VSUBS 0.276978f
C1171 VTAIL.t8 VSUBS 0.276978f
C1172 VTAIL.n0 VSUBS 1.99554f
C1173 VTAIL.n1 VSUBS 1.11677f
C1174 VTAIL.t15 VSUBS 2.63813f
C1175 VTAIL.n2 VSUBS 1.30216f
C1176 VTAIL.t14 VSUBS 0.276978f
C1177 VTAIL.t10 VSUBS 0.276978f
C1178 VTAIL.n3 VSUBS 1.99554f
C1179 VTAIL.n4 VSUBS 1.30062f
C1180 VTAIL.t12 VSUBS 0.276978f
C1181 VTAIL.t19 VSUBS 0.276978f
C1182 VTAIL.n5 VSUBS 1.99554f
C1183 VTAIL.n6 VSUBS 2.99144f
C1184 VTAIL.t3 VSUBS 0.276978f
C1185 VTAIL.t1 VSUBS 0.276978f
C1186 VTAIL.n7 VSUBS 1.99554f
C1187 VTAIL.n8 VSUBS 2.99143f
C1188 VTAIL.t6 VSUBS 0.276978f
C1189 VTAIL.t4 VSUBS 0.276978f
C1190 VTAIL.n9 VSUBS 1.99554f
C1191 VTAIL.n10 VSUBS 1.30061f
C1192 VTAIL.t5 VSUBS 2.63814f
C1193 VTAIL.n11 VSUBS 1.30215f
C1194 VTAIL.t13 VSUBS 0.276978f
C1195 VTAIL.t17 VSUBS 0.276978f
C1196 VTAIL.n12 VSUBS 1.99554f
C1197 VTAIL.n13 VSUBS 1.18935f
C1198 VTAIL.t11 VSUBS 0.276978f
C1199 VTAIL.t16 VSUBS 0.276978f
C1200 VTAIL.n14 VSUBS 1.99554f
C1201 VTAIL.n15 VSUBS 1.30061f
C1202 VTAIL.t18 VSUBS 2.63813f
C1203 VTAIL.n16 VSUBS 2.79156f
C1204 VTAIL.t2 VSUBS 2.63813f
C1205 VTAIL.n17 VSUBS 2.79156f
C1206 VTAIL.t7 VSUBS 0.276978f
C1207 VTAIL.t0 VSUBS 0.276978f
C1208 VTAIL.n18 VSUBS 1.99554f
C1209 VTAIL.n19 VSUBS 1.06052f
C1210 VP.t9 VSUBS 2.94522f
C1211 VP.n0 VSUBS 1.14487f
C1212 VP.n1 VSUBS 0.026635f
C1213 VP.n2 VSUBS 0.023805f
C1214 VP.n3 VSUBS 0.026635f
C1215 VP.t3 VSUBS 2.94522f
C1216 VP.n4 VSUBS 1.03486f
C1217 VP.n5 VSUBS 0.026635f
C1218 VP.n6 VSUBS 0.046686f
C1219 VP.n7 VSUBS 0.026635f
C1220 VP.n8 VSUBS 0.037387f
C1221 VP.n9 VSUBS 0.026635f
C1222 VP.n10 VSUBS 0.029089f
C1223 VP.n11 VSUBS 0.026635f
C1224 VP.n12 VSUBS 0.026604f
C1225 VP.n13 VSUBS 0.026635f
C1226 VP.n14 VSUBS 0.023805f
C1227 VP.n15 VSUBS 0.026635f
C1228 VP.t0 VSUBS 2.94522f
C1229 VP.n16 VSUBS 1.14487f
C1230 VP.t2 VSUBS 2.94522f
C1231 VP.n17 VSUBS 1.14487f
C1232 VP.n18 VSUBS 0.026635f
C1233 VP.n19 VSUBS 0.023805f
C1234 VP.n20 VSUBS 0.026635f
C1235 VP.t4 VSUBS 2.94522f
C1236 VP.n21 VSUBS 1.03486f
C1237 VP.n22 VSUBS 0.026635f
C1238 VP.n23 VSUBS 0.046686f
C1239 VP.n24 VSUBS 0.026635f
C1240 VP.n25 VSUBS 0.037387f
C1241 VP.n26 VSUBS 0.026635f
C1242 VP.n27 VSUBS 0.029089f
C1243 VP.n28 VSUBS 0.026635f
C1244 VP.n29 VSUBS 0.026604f
C1245 VP.t6 VSUBS 3.29663f
C1246 VP.t1 VSUBS 2.94522f
C1247 VP.n30 VSUBS 1.11658f
C1248 VP.n31 VSUBS 1.06314f
C1249 VP.n32 VSUBS 0.317801f
C1250 VP.n33 VSUBS 0.026635f
C1251 VP.n34 VSUBS 0.049642f
C1252 VP.n35 VSUBS 0.049642f
C1253 VP.n36 VSUBS 0.046686f
C1254 VP.n37 VSUBS 0.026635f
C1255 VP.n38 VSUBS 0.026635f
C1256 VP.n39 VSUBS 0.026635f
C1257 VP.n40 VSUBS 0.051632f
C1258 VP.n41 VSUBS 0.049642f
C1259 VP.t7 VSUBS 2.94522f
C1260 VP.n42 VSUBS 1.03486f
C1261 VP.n43 VSUBS 0.037387f
C1262 VP.n44 VSUBS 0.026635f
C1263 VP.n45 VSUBS 0.026635f
C1264 VP.n46 VSUBS 0.026635f
C1265 VP.n47 VSUBS 0.049642f
C1266 VP.n48 VSUBS 0.051632f
C1267 VP.n49 VSUBS 0.029089f
C1268 VP.n50 VSUBS 0.026635f
C1269 VP.n51 VSUBS 0.026635f
C1270 VP.n52 VSUBS 0.026635f
C1271 VP.n53 VSUBS 0.049642f
C1272 VP.n54 VSUBS 0.049642f
C1273 VP.n55 VSUBS 0.026604f
C1274 VP.n56 VSUBS 0.026635f
C1275 VP.n57 VSUBS 0.026635f
C1276 VP.n58 VSUBS 0.048171f
C1277 VP.n59 VSUBS 0.049642f
C1278 VP.n60 VSUBS 0.049881f
C1279 VP.n61 VSUBS 0.026635f
C1280 VP.n62 VSUBS 0.026635f
C1281 VP.n63 VSUBS 0.026635f
C1282 VP.n64 VSUBS 0.053721f
C1283 VP.n65 VSUBS 0.049642f
C1284 VP.n66 VSUBS 0.040328f
C1285 VP.n67 VSUBS 0.042989f
C1286 VP.n68 VSUBS 1.85391f
C1287 VP.n69 VSUBS 1.8705f
C1288 VP.n70 VSUBS 0.042989f
C1289 VP.n71 VSUBS 0.040328f
C1290 VP.n72 VSUBS 0.049642f
C1291 VP.n73 VSUBS 0.053721f
C1292 VP.n74 VSUBS 0.026635f
C1293 VP.n75 VSUBS 0.026635f
C1294 VP.n76 VSUBS 0.026635f
C1295 VP.n77 VSUBS 0.049881f
C1296 VP.n78 VSUBS 0.049642f
C1297 VP.t8 VSUBS 2.94522f
C1298 VP.n79 VSUBS 1.03486f
C1299 VP.n80 VSUBS 0.048171f
C1300 VP.n81 VSUBS 0.026635f
C1301 VP.n82 VSUBS 0.026635f
C1302 VP.n83 VSUBS 0.026635f
C1303 VP.n84 VSUBS 0.049642f
C1304 VP.n85 VSUBS 0.049642f
C1305 VP.n86 VSUBS 0.046686f
C1306 VP.n87 VSUBS 0.026635f
C1307 VP.n88 VSUBS 0.026635f
C1308 VP.n89 VSUBS 0.026635f
C1309 VP.n90 VSUBS 0.051632f
C1310 VP.n91 VSUBS 0.049642f
C1311 VP.t5 VSUBS 2.94522f
C1312 VP.n92 VSUBS 1.03486f
C1313 VP.n93 VSUBS 0.037387f
C1314 VP.n94 VSUBS 0.026635f
C1315 VP.n95 VSUBS 0.026635f
C1316 VP.n96 VSUBS 0.026635f
C1317 VP.n97 VSUBS 0.049642f
C1318 VP.n98 VSUBS 0.051632f
C1319 VP.n99 VSUBS 0.029089f
C1320 VP.n100 VSUBS 0.026635f
C1321 VP.n101 VSUBS 0.026635f
C1322 VP.n102 VSUBS 0.026635f
C1323 VP.n103 VSUBS 0.049642f
C1324 VP.n104 VSUBS 0.049642f
C1325 VP.n105 VSUBS 0.026604f
C1326 VP.n106 VSUBS 0.026635f
C1327 VP.n107 VSUBS 0.026635f
C1328 VP.n108 VSUBS 0.048171f
C1329 VP.n109 VSUBS 0.049642f
C1330 VP.n110 VSUBS 0.049881f
C1331 VP.n111 VSUBS 0.026635f
C1332 VP.n112 VSUBS 0.026635f
C1333 VP.n113 VSUBS 0.026635f
C1334 VP.n114 VSUBS 0.053721f
C1335 VP.n115 VSUBS 0.049642f
C1336 VP.n116 VSUBS 0.040328f
C1337 VP.n117 VSUBS 0.042989f
C1338 VP.n118 VSUBS 0.065535f
.ends

