* NGSPICE file created from diff_pair_sample_0802.ext - technology: sky130A

.subckt diff_pair_sample_0802 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=6.9264 pd=36.3 as=6.9264 ps=36.3 w=17.76 l=2.13
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=6.9264 pd=36.3 as=0 ps=0 w=17.76 l=2.13
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=6.9264 pd=36.3 as=0 ps=0 w=17.76 l=2.13
X3 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.9264 pd=36.3 as=6.9264 ps=36.3 w=17.76 l=2.13
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.9264 pd=36.3 as=0 ps=0 w=17.76 l=2.13
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=6.9264 pd=36.3 as=0 ps=0 w=17.76 l=2.13
X6 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=6.9264 pd=36.3 as=6.9264 ps=36.3 w=17.76 l=2.13
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.9264 pd=36.3 as=6.9264 ps=36.3 w=17.76 l=2.13
R0 VN VN.t1 297.943
R1 VN VN.t0 250.41
R2 VTAIL.n1 VTAIL.t3 42.7728
R3 VTAIL.n3 VTAIL.t2 42.7726
R4 VTAIL.n0 VTAIL.t1 42.7726
R5 VTAIL.n2 VTAIL.t0 42.7726
R6 VTAIL.n1 VTAIL.n0 31.9186
R7 VTAIL.n3 VTAIL.n2 29.7979
R8 VTAIL.n2 VTAIL.n1 1.53067
R9 VTAIL VTAIL.n0 1.05869
R10 VTAIL VTAIL.n3 0.472483
R11 VDD2.n0 VDD2.t1 102.662
R12 VDD2.n0 VDD2.t0 59.4513
R13 VDD2 VDD2.n0 0.588862
R14 B.n575 B.n574 585
R15 B.n575 B.n44 585
R16 B.n578 B.n577 585
R17 B.n579 B.n112 585
R18 B.n581 B.n580 585
R19 B.n583 B.n111 585
R20 B.n586 B.n585 585
R21 B.n587 B.n110 585
R22 B.n589 B.n588 585
R23 B.n591 B.n109 585
R24 B.n594 B.n593 585
R25 B.n595 B.n108 585
R26 B.n597 B.n596 585
R27 B.n599 B.n107 585
R28 B.n602 B.n601 585
R29 B.n603 B.n106 585
R30 B.n605 B.n604 585
R31 B.n607 B.n105 585
R32 B.n610 B.n609 585
R33 B.n611 B.n104 585
R34 B.n613 B.n612 585
R35 B.n615 B.n103 585
R36 B.n618 B.n617 585
R37 B.n619 B.n102 585
R38 B.n621 B.n620 585
R39 B.n623 B.n101 585
R40 B.n626 B.n625 585
R41 B.n627 B.n100 585
R42 B.n629 B.n628 585
R43 B.n631 B.n99 585
R44 B.n634 B.n633 585
R45 B.n635 B.n98 585
R46 B.n637 B.n636 585
R47 B.n639 B.n97 585
R48 B.n642 B.n641 585
R49 B.n643 B.n96 585
R50 B.n645 B.n644 585
R51 B.n647 B.n95 585
R52 B.n650 B.n649 585
R53 B.n651 B.n94 585
R54 B.n653 B.n652 585
R55 B.n655 B.n93 585
R56 B.n658 B.n657 585
R57 B.n659 B.n92 585
R58 B.n661 B.n660 585
R59 B.n663 B.n91 585
R60 B.n666 B.n665 585
R61 B.n667 B.n90 585
R62 B.n669 B.n668 585
R63 B.n671 B.n89 585
R64 B.n674 B.n673 585
R65 B.n675 B.n88 585
R66 B.n677 B.n676 585
R67 B.n679 B.n87 585
R68 B.n682 B.n681 585
R69 B.n683 B.n86 585
R70 B.n685 B.n684 585
R71 B.n687 B.n85 585
R72 B.n690 B.n689 585
R73 B.n691 B.n82 585
R74 B.n694 B.n693 585
R75 B.n696 B.n81 585
R76 B.n699 B.n698 585
R77 B.n700 B.n80 585
R78 B.n702 B.n701 585
R79 B.n704 B.n79 585
R80 B.n707 B.n706 585
R81 B.n708 B.n75 585
R82 B.n710 B.n709 585
R83 B.n712 B.n74 585
R84 B.n715 B.n714 585
R85 B.n716 B.n73 585
R86 B.n718 B.n717 585
R87 B.n720 B.n72 585
R88 B.n723 B.n722 585
R89 B.n724 B.n71 585
R90 B.n726 B.n725 585
R91 B.n728 B.n70 585
R92 B.n731 B.n730 585
R93 B.n732 B.n69 585
R94 B.n734 B.n733 585
R95 B.n736 B.n68 585
R96 B.n739 B.n738 585
R97 B.n740 B.n67 585
R98 B.n742 B.n741 585
R99 B.n744 B.n66 585
R100 B.n747 B.n746 585
R101 B.n748 B.n65 585
R102 B.n750 B.n749 585
R103 B.n752 B.n64 585
R104 B.n755 B.n754 585
R105 B.n756 B.n63 585
R106 B.n758 B.n757 585
R107 B.n760 B.n62 585
R108 B.n763 B.n762 585
R109 B.n764 B.n61 585
R110 B.n766 B.n765 585
R111 B.n768 B.n60 585
R112 B.n771 B.n770 585
R113 B.n772 B.n59 585
R114 B.n774 B.n773 585
R115 B.n776 B.n58 585
R116 B.n779 B.n778 585
R117 B.n780 B.n57 585
R118 B.n782 B.n781 585
R119 B.n784 B.n56 585
R120 B.n787 B.n786 585
R121 B.n788 B.n55 585
R122 B.n790 B.n789 585
R123 B.n792 B.n54 585
R124 B.n795 B.n794 585
R125 B.n796 B.n53 585
R126 B.n798 B.n797 585
R127 B.n800 B.n52 585
R128 B.n803 B.n802 585
R129 B.n804 B.n51 585
R130 B.n806 B.n805 585
R131 B.n808 B.n50 585
R132 B.n811 B.n810 585
R133 B.n812 B.n49 585
R134 B.n814 B.n813 585
R135 B.n816 B.n48 585
R136 B.n819 B.n818 585
R137 B.n820 B.n47 585
R138 B.n822 B.n821 585
R139 B.n824 B.n46 585
R140 B.n827 B.n826 585
R141 B.n828 B.n45 585
R142 B.n573 B.n43 585
R143 B.n831 B.n43 585
R144 B.n572 B.n42 585
R145 B.n832 B.n42 585
R146 B.n571 B.n41 585
R147 B.n833 B.n41 585
R148 B.n570 B.n569 585
R149 B.n569 B.n37 585
R150 B.n568 B.n36 585
R151 B.n839 B.n36 585
R152 B.n567 B.n35 585
R153 B.n840 B.n35 585
R154 B.n566 B.n34 585
R155 B.n841 B.n34 585
R156 B.n565 B.n564 585
R157 B.n564 B.n30 585
R158 B.n563 B.n29 585
R159 B.n847 B.n29 585
R160 B.n562 B.n28 585
R161 B.n848 B.n28 585
R162 B.n561 B.n27 585
R163 B.n849 B.n27 585
R164 B.n560 B.n559 585
R165 B.n559 B.n23 585
R166 B.n558 B.n22 585
R167 B.n855 B.n22 585
R168 B.n557 B.n21 585
R169 B.n856 B.n21 585
R170 B.n556 B.n20 585
R171 B.n857 B.n20 585
R172 B.n555 B.n554 585
R173 B.n554 B.n16 585
R174 B.n553 B.n15 585
R175 B.n863 B.n15 585
R176 B.n552 B.n14 585
R177 B.n864 B.n14 585
R178 B.n551 B.n13 585
R179 B.n865 B.n13 585
R180 B.n550 B.n549 585
R181 B.n549 B.n12 585
R182 B.n548 B.n547 585
R183 B.n548 B.n8 585
R184 B.n546 B.n7 585
R185 B.n872 B.n7 585
R186 B.n545 B.n6 585
R187 B.n873 B.n6 585
R188 B.n544 B.n5 585
R189 B.n874 B.n5 585
R190 B.n543 B.n542 585
R191 B.n542 B.n4 585
R192 B.n541 B.n113 585
R193 B.n541 B.n540 585
R194 B.n531 B.n114 585
R195 B.n115 B.n114 585
R196 B.n533 B.n532 585
R197 B.n534 B.n533 585
R198 B.n530 B.n119 585
R199 B.n123 B.n119 585
R200 B.n529 B.n528 585
R201 B.n528 B.n527 585
R202 B.n121 B.n120 585
R203 B.n122 B.n121 585
R204 B.n520 B.n519 585
R205 B.n521 B.n520 585
R206 B.n518 B.n128 585
R207 B.n128 B.n127 585
R208 B.n517 B.n516 585
R209 B.n516 B.n515 585
R210 B.n130 B.n129 585
R211 B.n131 B.n130 585
R212 B.n508 B.n507 585
R213 B.n509 B.n508 585
R214 B.n506 B.n136 585
R215 B.n136 B.n135 585
R216 B.n505 B.n504 585
R217 B.n504 B.n503 585
R218 B.n138 B.n137 585
R219 B.n139 B.n138 585
R220 B.n496 B.n495 585
R221 B.n497 B.n496 585
R222 B.n494 B.n144 585
R223 B.n144 B.n143 585
R224 B.n493 B.n492 585
R225 B.n492 B.n491 585
R226 B.n146 B.n145 585
R227 B.n147 B.n146 585
R228 B.n484 B.n483 585
R229 B.n485 B.n484 585
R230 B.n482 B.n152 585
R231 B.n152 B.n151 585
R232 B.n481 B.n480 585
R233 B.n480 B.n479 585
R234 B.n476 B.n156 585
R235 B.n475 B.n474 585
R236 B.n472 B.n157 585
R237 B.n472 B.n155 585
R238 B.n471 B.n470 585
R239 B.n469 B.n468 585
R240 B.n467 B.n159 585
R241 B.n465 B.n464 585
R242 B.n463 B.n160 585
R243 B.n462 B.n461 585
R244 B.n459 B.n161 585
R245 B.n457 B.n456 585
R246 B.n455 B.n162 585
R247 B.n454 B.n453 585
R248 B.n451 B.n163 585
R249 B.n449 B.n448 585
R250 B.n447 B.n164 585
R251 B.n446 B.n445 585
R252 B.n443 B.n165 585
R253 B.n441 B.n440 585
R254 B.n439 B.n166 585
R255 B.n438 B.n437 585
R256 B.n435 B.n167 585
R257 B.n433 B.n432 585
R258 B.n431 B.n168 585
R259 B.n430 B.n429 585
R260 B.n427 B.n169 585
R261 B.n425 B.n424 585
R262 B.n423 B.n170 585
R263 B.n422 B.n421 585
R264 B.n419 B.n171 585
R265 B.n417 B.n416 585
R266 B.n415 B.n172 585
R267 B.n414 B.n413 585
R268 B.n411 B.n173 585
R269 B.n409 B.n408 585
R270 B.n407 B.n174 585
R271 B.n406 B.n405 585
R272 B.n403 B.n175 585
R273 B.n401 B.n400 585
R274 B.n399 B.n176 585
R275 B.n398 B.n397 585
R276 B.n395 B.n177 585
R277 B.n393 B.n392 585
R278 B.n391 B.n178 585
R279 B.n390 B.n389 585
R280 B.n387 B.n179 585
R281 B.n385 B.n384 585
R282 B.n383 B.n180 585
R283 B.n382 B.n381 585
R284 B.n379 B.n181 585
R285 B.n377 B.n376 585
R286 B.n375 B.n182 585
R287 B.n374 B.n373 585
R288 B.n371 B.n183 585
R289 B.n369 B.n368 585
R290 B.n367 B.n184 585
R291 B.n366 B.n365 585
R292 B.n363 B.n185 585
R293 B.n361 B.n360 585
R294 B.n358 B.n186 585
R295 B.n357 B.n356 585
R296 B.n354 B.n189 585
R297 B.n352 B.n351 585
R298 B.n350 B.n190 585
R299 B.n349 B.n348 585
R300 B.n346 B.n191 585
R301 B.n344 B.n343 585
R302 B.n342 B.n192 585
R303 B.n340 B.n339 585
R304 B.n337 B.n195 585
R305 B.n335 B.n334 585
R306 B.n333 B.n196 585
R307 B.n332 B.n331 585
R308 B.n329 B.n197 585
R309 B.n327 B.n326 585
R310 B.n325 B.n198 585
R311 B.n324 B.n323 585
R312 B.n321 B.n199 585
R313 B.n319 B.n318 585
R314 B.n317 B.n200 585
R315 B.n316 B.n315 585
R316 B.n313 B.n201 585
R317 B.n311 B.n310 585
R318 B.n309 B.n202 585
R319 B.n308 B.n307 585
R320 B.n305 B.n203 585
R321 B.n303 B.n302 585
R322 B.n301 B.n204 585
R323 B.n300 B.n299 585
R324 B.n297 B.n205 585
R325 B.n295 B.n294 585
R326 B.n293 B.n206 585
R327 B.n292 B.n291 585
R328 B.n289 B.n207 585
R329 B.n287 B.n286 585
R330 B.n285 B.n208 585
R331 B.n284 B.n283 585
R332 B.n281 B.n209 585
R333 B.n279 B.n278 585
R334 B.n277 B.n210 585
R335 B.n276 B.n275 585
R336 B.n273 B.n211 585
R337 B.n271 B.n270 585
R338 B.n269 B.n212 585
R339 B.n268 B.n267 585
R340 B.n265 B.n213 585
R341 B.n263 B.n262 585
R342 B.n261 B.n214 585
R343 B.n260 B.n259 585
R344 B.n257 B.n215 585
R345 B.n255 B.n254 585
R346 B.n253 B.n216 585
R347 B.n252 B.n251 585
R348 B.n249 B.n217 585
R349 B.n247 B.n246 585
R350 B.n245 B.n218 585
R351 B.n244 B.n243 585
R352 B.n241 B.n219 585
R353 B.n239 B.n238 585
R354 B.n237 B.n220 585
R355 B.n236 B.n235 585
R356 B.n233 B.n221 585
R357 B.n231 B.n230 585
R358 B.n229 B.n222 585
R359 B.n228 B.n227 585
R360 B.n225 B.n223 585
R361 B.n154 B.n153 585
R362 B.n478 B.n477 585
R363 B.n479 B.n478 585
R364 B.n150 B.n149 585
R365 B.n151 B.n150 585
R366 B.n487 B.n486 585
R367 B.n486 B.n485 585
R368 B.n488 B.n148 585
R369 B.n148 B.n147 585
R370 B.n490 B.n489 585
R371 B.n491 B.n490 585
R372 B.n142 B.n141 585
R373 B.n143 B.n142 585
R374 B.n499 B.n498 585
R375 B.n498 B.n497 585
R376 B.n500 B.n140 585
R377 B.n140 B.n139 585
R378 B.n502 B.n501 585
R379 B.n503 B.n502 585
R380 B.n134 B.n133 585
R381 B.n135 B.n134 585
R382 B.n511 B.n510 585
R383 B.n510 B.n509 585
R384 B.n512 B.n132 585
R385 B.n132 B.n131 585
R386 B.n514 B.n513 585
R387 B.n515 B.n514 585
R388 B.n126 B.n125 585
R389 B.n127 B.n126 585
R390 B.n523 B.n522 585
R391 B.n522 B.n521 585
R392 B.n524 B.n124 585
R393 B.n124 B.n122 585
R394 B.n526 B.n525 585
R395 B.n527 B.n526 585
R396 B.n118 B.n117 585
R397 B.n123 B.n118 585
R398 B.n536 B.n535 585
R399 B.n535 B.n534 585
R400 B.n537 B.n116 585
R401 B.n116 B.n115 585
R402 B.n539 B.n538 585
R403 B.n540 B.n539 585
R404 B.n3 B.n0 585
R405 B.n4 B.n3 585
R406 B.n871 B.n1 585
R407 B.n872 B.n871 585
R408 B.n870 B.n869 585
R409 B.n870 B.n8 585
R410 B.n868 B.n9 585
R411 B.n12 B.n9 585
R412 B.n867 B.n866 585
R413 B.n866 B.n865 585
R414 B.n11 B.n10 585
R415 B.n864 B.n11 585
R416 B.n862 B.n861 585
R417 B.n863 B.n862 585
R418 B.n860 B.n17 585
R419 B.n17 B.n16 585
R420 B.n859 B.n858 585
R421 B.n858 B.n857 585
R422 B.n19 B.n18 585
R423 B.n856 B.n19 585
R424 B.n854 B.n853 585
R425 B.n855 B.n854 585
R426 B.n852 B.n24 585
R427 B.n24 B.n23 585
R428 B.n851 B.n850 585
R429 B.n850 B.n849 585
R430 B.n26 B.n25 585
R431 B.n848 B.n26 585
R432 B.n846 B.n845 585
R433 B.n847 B.n846 585
R434 B.n844 B.n31 585
R435 B.n31 B.n30 585
R436 B.n843 B.n842 585
R437 B.n842 B.n841 585
R438 B.n33 B.n32 585
R439 B.n840 B.n33 585
R440 B.n838 B.n837 585
R441 B.n839 B.n838 585
R442 B.n836 B.n38 585
R443 B.n38 B.n37 585
R444 B.n835 B.n834 585
R445 B.n834 B.n833 585
R446 B.n40 B.n39 585
R447 B.n832 B.n40 585
R448 B.n830 B.n829 585
R449 B.n831 B.n830 585
R450 B.n875 B.n874 585
R451 B.n873 B.n2 585
R452 B.n830 B.n45 487.695
R453 B.n575 B.n43 487.695
R454 B.n480 B.n154 487.695
R455 B.n478 B.n156 487.695
R456 B.n76 B.t6 408.154
R457 B.n83 B.t13 408.154
R458 B.n193 B.t2 408.154
R459 B.n187 B.t10 408.154
R460 B.n576 B.n44 256.663
R461 B.n582 B.n44 256.663
R462 B.n584 B.n44 256.663
R463 B.n590 B.n44 256.663
R464 B.n592 B.n44 256.663
R465 B.n598 B.n44 256.663
R466 B.n600 B.n44 256.663
R467 B.n606 B.n44 256.663
R468 B.n608 B.n44 256.663
R469 B.n614 B.n44 256.663
R470 B.n616 B.n44 256.663
R471 B.n622 B.n44 256.663
R472 B.n624 B.n44 256.663
R473 B.n630 B.n44 256.663
R474 B.n632 B.n44 256.663
R475 B.n638 B.n44 256.663
R476 B.n640 B.n44 256.663
R477 B.n646 B.n44 256.663
R478 B.n648 B.n44 256.663
R479 B.n654 B.n44 256.663
R480 B.n656 B.n44 256.663
R481 B.n662 B.n44 256.663
R482 B.n664 B.n44 256.663
R483 B.n670 B.n44 256.663
R484 B.n672 B.n44 256.663
R485 B.n678 B.n44 256.663
R486 B.n680 B.n44 256.663
R487 B.n686 B.n44 256.663
R488 B.n688 B.n44 256.663
R489 B.n695 B.n44 256.663
R490 B.n697 B.n44 256.663
R491 B.n703 B.n44 256.663
R492 B.n705 B.n44 256.663
R493 B.n711 B.n44 256.663
R494 B.n713 B.n44 256.663
R495 B.n719 B.n44 256.663
R496 B.n721 B.n44 256.663
R497 B.n727 B.n44 256.663
R498 B.n729 B.n44 256.663
R499 B.n735 B.n44 256.663
R500 B.n737 B.n44 256.663
R501 B.n743 B.n44 256.663
R502 B.n745 B.n44 256.663
R503 B.n751 B.n44 256.663
R504 B.n753 B.n44 256.663
R505 B.n759 B.n44 256.663
R506 B.n761 B.n44 256.663
R507 B.n767 B.n44 256.663
R508 B.n769 B.n44 256.663
R509 B.n775 B.n44 256.663
R510 B.n777 B.n44 256.663
R511 B.n783 B.n44 256.663
R512 B.n785 B.n44 256.663
R513 B.n791 B.n44 256.663
R514 B.n793 B.n44 256.663
R515 B.n799 B.n44 256.663
R516 B.n801 B.n44 256.663
R517 B.n807 B.n44 256.663
R518 B.n809 B.n44 256.663
R519 B.n815 B.n44 256.663
R520 B.n817 B.n44 256.663
R521 B.n823 B.n44 256.663
R522 B.n825 B.n44 256.663
R523 B.n473 B.n155 256.663
R524 B.n158 B.n155 256.663
R525 B.n466 B.n155 256.663
R526 B.n460 B.n155 256.663
R527 B.n458 B.n155 256.663
R528 B.n452 B.n155 256.663
R529 B.n450 B.n155 256.663
R530 B.n444 B.n155 256.663
R531 B.n442 B.n155 256.663
R532 B.n436 B.n155 256.663
R533 B.n434 B.n155 256.663
R534 B.n428 B.n155 256.663
R535 B.n426 B.n155 256.663
R536 B.n420 B.n155 256.663
R537 B.n418 B.n155 256.663
R538 B.n412 B.n155 256.663
R539 B.n410 B.n155 256.663
R540 B.n404 B.n155 256.663
R541 B.n402 B.n155 256.663
R542 B.n396 B.n155 256.663
R543 B.n394 B.n155 256.663
R544 B.n388 B.n155 256.663
R545 B.n386 B.n155 256.663
R546 B.n380 B.n155 256.663
R547 B.n378 B.n155 256.663
R548 B.n372 B.n155 256.663
R549 B.n370 B.n155 256.663
R550 B.n364 B.n155 256.663
R551 B.n362 B.n155 256.663
R552 B.n355 B.n155 256.663
R553 B.n353 B.n155 256.663
R554 B.n347 B.n155 256.663
R555 B.n345 B.n155 256.663
R556 B.n338 B.n155 256.663
R557 B.n336 B.n155 256.663
R558 B.n330 B.n155 256.663
R559 B.n328 B.n155 256.663
R560 B.n322 B.n155 256.663
R561 B.n320 B.n155 256.663
R562 B.n314 B.n155 256.663
R563 B.n312 B.n155 256.663
R564 B.n306 B.n155 256.663
R565 B.n304 B.n155 256.663
R566 B.n298 B.n155 256.663
R567 B.n296 B.n155 256.663
R568 B.n290 B.n155 256.663
R569 B.n288 B.n155 256.663
R570 B.n282 B.n155 256.663
R571 B.n280 B.n155 256.663
R572 B.n274 B.n155 256.663
R573 B.n272 B.n155 256.663
R574 B.n266 B.n155 256.663
R575 B.n264 B.n155 256.663
R576 B.n258 B.n155 256.663
R577 B.n256 B.n155 256.663
R578 B.n250 B.n155 256.663
R579 B.n248 B.n155 256.663
R580 B.n242 B.n155 256.663
R581 B.n240 B.n155 256.663
R582 B.n234 B.n155 256.663
R583 B.n232 B.n155 256.663
R584 B.n226 B.n155 256.663
R585 B.n224 B.n155 256.663
R586 B.n877 B.n876 256.663
R587 B.n826 B.n824 163.367
R588 B.n822 B.n47 163.367
R589 B.n818 B.n816 163.367
R590 B.n814 B.n49 163.367
R591 B.n810 B.n808 163.367
R592 B.n806 B.n51 163.367
R593 B.n802 B.n800 163.367
R594 B.n798 B.n53 163.367
R595 B.n794 B.n792 163.367
R596 B.n790 B.n55 163.367
R597 B.n786 B.n784 163.367
R598 B.n782 B.n57 163.367
R599 B.n778 B.n776 163.367
R600 B.n774 B.n59 163.367
R601 B.n770 B.n768 163.367
R602 B.n766 B.n61 163.367
R603 B.n762 B.n760 163.367
R604 B.n758 B.n63 163.367
R605 B.n754 B.n752 163.367
R606 B.n750 B.n65 163.367
R607 B.n746 B.n744 163.367
R608 B.n742 B.n67 163.367
R609 B.n738 B.n736 163.367
R610 B.n734 B.n69 163.367
R611 B.n730 B.n728 163.367
R612 B.n726 B.n71 163.367
R613 B.n722 B.n720 163.367
R614 B.n718 B.n73 163.367
R615 B.n714 B.n712 163.367
R616 B.n710 B.n75 163.367
R617 B.n706 B.n704 163.367
R618 B.n702 B.n80 163.367
R619 B.n698 B.n696 163.367
R620 B.n694 B.n82 163.367
R621 B.n689 B.n687 163.367
R622 B.n685 B.n86 163.367
R623 B.n681 B.n679 163.367
R624 B.n677 B.n88 163.367
R625 B.n673 B.n671 163.367
R626 B.n669 B.n90 163.367
R627 B.n665 B.n663 163.367
R628 B.n661 B.n92 163.367
R629 B.n657 B.n655 163.367
R630 B.n653 B.n94 163.367
R631 B.n649 B.n647 163.367
R632 B.n645 B.n96 163.367
R633 B.n641 B.n639 163.367
R634 B.n637 B.n98 163.367
R635 B.n633 B.n631 163.367
R636 B.n629 B.n100 163.367
R637 B.n625 B.n623 163.367
R638 B.n621 B.n102 163.367
R639 B.n617 B.n615 163.367
R640 B.n613 B.n104 163.367
R641 B.n609 B.n607 163.367
R642 B.n605 B.n106 163.367
R643 B.n601 B.n599 163.367
R644 B.n597 B.n108 163.367
R645 B.n593 B.n591 163.367
R646 B.n589 B.n110 163.367
R647 B.n585 B.n583 163.367
R648 B.n581 B.n112 163.367
R649 B.n577 B.n575 163.367
R650 B.n480 B.n152 163.367
R651 B.n484 B.n152 163.367
R652 B.n484 B.n146 163.367
R653 B.n492 B.n146 163.367
R654 B.n492 B.n144 163.367
R655 B.n496 B.n144 163.367
R656 B.n496 B.n138 163.367
R657 B.n504 B.n138 163.367
R658 B.n504 B.n136 163.367
R659 B.n508 B.n136 163.367
R660 B.n508 B.n130 163.367
R661 B.n516 B.n130 163.367
R662 B.n516 B.n128 163.367
R663 B.n520 B.n128 163.367
R664 B.n520 B.n121 163.367
R665 B.n528 B.n121 163.367
R666 B.n528 B.n119 163.367
R667 B.n533 B.n119 163.367
R668 B.n533 B.n114 163.367
R669 B.n541 B.n114 163.367
R670 B.n542 B.n541 163.367
R671 B.n542 B.n5 163.367
R672 B.n6 B.n5 163.367
R673 B.n7 B.n6 163.367
R674 B.n548 B.n7 163.367
R675 B.n549 B.n548 163.367
R676 B.n549 B.n13 163.367
R677 B.n14 B.n13 163.367
R678 B.n15 B.n14 163.367
R679 B.n554 B.n15 163.367
R680 B.n554 B.n20 163.367
R681 B.n21 B.n20 163.367
R682 B.n22 B.n21 163.367
R683 B.n559 B.n22 163.367
R684 B.n559 B.n27 163.367
R685 B.n28 B.n27 163.367
R686 B.n29 B.n28 163.367
R687 B.n564 B.n29 163.367
R688 B.n564 B.n34 163.367
R689 B.n35 B.n34 163.367
R690 B.n36 B.n35 163.367
R691 B.n569 B.n36 163.367
R692 B.n569 B.n41 163.367
R693 B.n42 B.n41 163.367
R694 B.n43 B.n42 163.367
R695 B.n474 B.n472 163.367
R696 B.n472 B.n471 163.367
R697 B.n468 B.n467 163.367
R698 B.n465 B.n160 163.367
R699 B.n461 B.n459 163.367
R700 B.n457 B.n162 163.367
R701 B.n453 B.n451 163.367
R702 B.n449 B.n164 163.367
R703 B.n445 B.n443 163.367
R704 B.n441 B.n166 163.367
R705 B.n437 B.n435 163.367
R706 B.n433 B.n168 163.367
R707 B.n429 B.n427 163.367
R708 B.n425 B.n170 163.367
R709 B.n421 B.n419 163.367
R710 B.n417 B.n172 163.367
R711 B.n413 B.n411 163.367
R712 B.n409 B.n174 163.367
R713 B.n405 B.n403 163.367
R714 B.n401 B.n176 163.367
R715 B.n397 B.n395 163.367
R716 B.n393 B.n178 163.367
R717 B.n389 B.n387 163.367
R718 B.n385 B.n180 163.367
R719 B.n381 B.n379 163.367
R720 B.n377 B.n182 163.367
R721 B.n373 B.n371 163.367
R722 B.n369 B.n184 163.367
R723 B.n365 B.n363 163.367
R724 B.n361 B.n186 163.367
R725 B.n356 B.n354 163.367
R726 B.n352 B.n190 163.367
R727 B.n348 B.n346 163.367
R728 B.n344 B.n192 163.367
R729 B.n339 B.n337 163.367
R730 B.n335 B.n196 163.367
R731 B.n331 B.n329 163.367
R732 B.n327 B.n198 163.367
R733 B.n323 B.n321 163.367
R734 B.n319 B.n200 163.367
R735 B.n315 B.n313 163.367
R736 B.n311 B.n202 163.367
R737 B.n307 B.n305 163.367
R738 B.n303 B.n204 163.367
R739 B.n299 B.n297 163.367
R740 B.n295 B.n206 163.367
R741 B.n291 B.n289 163.367
R742 B.n287 B.n208 163.367
R743 B.n283 B.n281 163.367
R744 B.n279 B.n210 163.367
R745 B.n275 B.n273 163.367
R746 B.n271 B.n212 163.367
R747 B.n267 B.n265 163.367
R748 B.n263 B.n214 163.367
R749 B.n259 B.n257 163.367
R750 B.n255 B.n216 163.367
R751 B.n251 B.n249 163.367
R752 B.n247 B.n218 163.367
R753 B.n243 B.n241 163.367
R754 B.n239 B.n220 163.367
R755 B.n235 B.n233 163.367
R756 B.n231 B.n222 163.367
R757 B.n227 B.n225 163.367
R758 B.n478 B.n150 163.367
R759 B.n486 B.n150 163.367
R760 B.n486 B.n148 163.367
R761 B.n490 B.n148 163.367
R762 B.n490 B.n142 163.367
R763 B.n498 B.n142 163.367
R764 B.n498 B.n140 163.367
R765 B.n502 B.n140 163.367
R766 B.n502 B.n134 163.367
R767 B.n510 B.n134 163.367
R768 B.n510 B.n132 163.367
R769 B.n514 B.n132 163.367
R770 B.n514 B.n126 163.367
R771 B.n522 B.n126 163.367
R772 B.n522 B.n124 163.367
R773 B.n526 B.n124 163.367
R774 B.n526 B.n118 163.367
R775 B.n535 B.n118 163.367
R776 B.n535 B.n116 163.367
R777 B.n539 B.n116 163.367
R778 B.n539 B.n3 163.367
R779 B.n875 B.n3 163.367
R780 B.n871 B.n2 163.367
R781 B.n871 B.n870 163.367
R782 B.n870 B.n9 163.367
R783 B.n866 B.n9 163.367
R784 B.n866 B.n11 163.367
R785 B.n862 B.n11 163.367
R786 B.n862 B.n17 163.367
R787 B.n858 B.n17 163.367
R788 B.n858 B.n19 163.367
R789 B.n854 B.n19 163.367
R790 B.n854 B.n24 163.367
R791 B.n850 B.n24 163.367
R792 B.n850 B.n26 163.367
R793 B.n846 B.n26 163.367
R794 B.n846 B.n31 163.367
R795 B.n842 B.n31 163.367
R796 B.n842 B.n33 163.367
R797 B.n838 B.n33 163.367
R798 B.n838 B.n38 163.367
R799 B.n834 B.n38 163.367
R800 B.n834 B.n40 163.367
R801 B.n830 B.n40 163.367
R802 B.n83 B.t14 116.523
R803 B.n193 B.t5 116.523
R804 B.n76 B.t8 116.501
R805 B.n187 B.t12 116.501
R806 B.n825 B.n45 71.676
R807 B.n824 B.n823 71.676
R808 B.n817 B.n47 71.676
R809 B.n816 B.n815 71.676
R810 B.n809 B.n49 71.676
R811 B.n808 B.n807 71.676
R812 B.n801 B.n51 71.676
R813 B.n800 B.n799 71.676
R814 B.n793 B.n53 71.676
R815 B.n792 B.n791 71.676
R816 B.n785 B.n55 71.676
R817 B.n784 B.n783 71.676
R818 B.n777 B.n57 71.676
R819 B.n776 B.n775 71.676
R820 B.n769 B.n59 71.676
R821 B.n768 B.n767 71.676
R822 B.n761 B.n61 71.676
R823 B.n760 B.n759 71.676
R824 B.n753 B.n63 71.676
R825 B.n752 B.n751 71.676
R826 B.n745 B.n65 71.676
R827 B.n744 B.n743 71.676
R828 B.n737 B.n67 71.676
R829 B.n736 B.n735 71.676
R830 B.n729 B.n69 71.676
R831 B.n728 B.n727 71.676
R832 B.n721 B.n71 71.676
R833 B.n720 B.n719 71.676
R834 B.n713 B.n73 71.676
R835 B.n712 B.n711 71.676
R836 B.n705 B.n75 71.676
R837 B.n704 B.n703 71.676
R838 B.n697 B.n80 71.676
R839 B.n696 B.n695 71.676
R840 B.n688 B.n82 71.676
R841 B.n687 B.n686 71.676
R842 B.n680 B.n86 71.676
R843 B.n679 B.n678 71.676
R844 B.n672 B.n88 71.676
R845 B.n671 B.n670 71.676
R846 B.n664 B.n90 71.676
R847 B.n663 B.n662 71.676
R848 B.n656 B.n92 71.676
R849 B.n655 B.n654 71.676
R850 B.n648 B.n94 71.676
R851 B.n647 B.n646 71.676
R852 B.n640 B.n96 71.676
R853 B.n639 B.n638 71.676
R854 B.n632 B.n98 71.676
R855 B.n631 B.n630 71.676
R856 B.n624 B.n100 71.676
R857 B.n623 B.n622 71.676
R858 B.n616 B.n102 71.676
R859 B.n615 B.n614 71.676
R860 B.n608 B.n104 71.676
R861 B.n607 B.n606 71.676
R862 B.n600 B.n106 71.676
R863 B.n599 B.n598 71.676
R864 B.n592 B.n108 71.676
R865 B.n591 B.n590 71.676
R866 B.n584 B.n110 71.676
R867 B.n583 B.n582 71.676
R868 B.n576 B.n112 71.676
R869 B.n577 B.n576 71.676
R870 B.n582 B.n581 71.676
R871 B.n585 B.n584 71.676
R872 B.n590 B.n589 71.676
R873 B.n593 B.n592 71.676
R874 B.n598 B.n597 71.676
R875 B.n601 B.n600 71.676
R876 B.n606 B.n605 71.676
R877 B.n609 B.n608 71.676
R878 B.n614 B.n613 71.676
R879 B.n617 B.n616 71.676
R880 B.n622 B.n621 71.676
R881 B.n625 B.n624 71.676
R882 B.n630 B.n629 71.676
R883 B.n633 B.n632 71.676
R884 B.n638 B.n637 71.676
R885 B.n641 B.n640 71.676
R886 B.n646 B.n645 71.676
R887 B.n649 B.n648 71.676
R888 B.n654 B.n653 71.676
R889 B.n657 B.n656 71.676
R890 B.n662 B.n661 71.676
R891 B.n665 B.n664 71.676
R892 B.n670 B.n669 71.676
R893 B.n673 B.n672 71.676
R894 B.n678 B.n677 71.676
R895 B.n681 B.n680 71.676
R896 B.n686 B.n685 71.676
R897 B.n689 B.n688 71.676
R898 B.n695 B.n694 71.676
R899 B.n698 B.n697 71.676
R900 B.n703 B.n702 71.676
R901 B.n706 B.n705 71.676
R902 B.n711 B.n710 71.676
R903 B.n714 B.n713 71.676
R904 B.n719 B.n718 71.676
R905 B.n722 B.n721 71.676
R906 B.n727 B.n726 71.676
R907 B.n730 B.n729 71.676
R908 B.n735 B.n734 71.676
R909 B.n738 B.n737 71.676
R910 B.n743 B.n742 71.676
R911 B.n746 B.n745 71.676
R912 B.n751 B.n750 71.676
R913 B.n754 B.n753 71.676
R914 B.n759 B.n758 71.676
R915 B.n762 B.n761 71.676
R916 B.n767 B.n766 71.676
R917 B.n770 B.n769 71.676
R918 B.n775 B.n774 71.676
R919 B.n778 B.n777 71.676
R920 B.n783 B.n782 71.676
R921 B.n786 B.n785 71.676
R922 B.n791 B.n790 71.676
R923 B.n794 B.n793 71.676
R924 B.n799 B.n798 71.676
R925 B.n802 B.n801 71.676
R926 B.n807 B.n806 71.676
R927 B.n810 B.n809 71.676
R928 B.n815 B.n814 71.676
R929 B.n818 B.n817 71.676
R930 B.n823 B.n822 71.676
R931 B.n826 B.n825 71.676
R932 B.n473 B.n156 71.676
R933 B.n471 B.n158 71.676
R934 B.n467 B.n466 71.676
R935 B.n460 B.n160 71.676
R936 B.n459 B.n458 71.676
R937 B.n452 B.n162 71.676
R938 B.n451 B.n450 71.676
R939 B.n444 B.n164 71.676
R940 B.n443 B.n442 71.676
R941 B.n436 B.n166 71.676
R942 B.n435 B.n434 71.676
R943 B.n428 B.n168 71.676
R944 B.n427 B.n426 71.676
R945 B.n420 B.n170 71.676
R946 B.n419 B.n418 71.676
R947 B.n412 B.n172 71.676
R948 B.n411 B.n410 71.676
R949 B.n404 B.n174 71.676
R950 B.n403 B.n402 71.676
R951 B.n396 B.n176 71.676
R952 B.n395 B.n394 71.676
R953 B.n388 B.n178 71.676
R954 B.n387 B.n386 71.676
R955 B.n380 B.n180 71.676
R956 B.n379 B.n378 71.676
R957 B.n372 B.n182 71.676
R958 B.n371 B.n370 71.676
R959 B.n364 B.n184 71.676
R960 B.n363 B.n362 71.676
R961 B.n355 B.n186 71.676
R962 B.n354 B.n353 71.676
R963 B.n347 B.n190 71.676
R964 B.n346 B.n345 71.676
R965 B.n338 B.n192 71.676
R966 B.n337 B.n336 71.676
R967 B.n330 B.n196 71.676
R968 B.n329 B.n328 71.676
R969 B.n322 B.n198 71.676
R970 B.n321 B.n320 71.676
R971 B.n314 B.n200 71.676
R972 B.n313 B.n312 71.676
R973 B.n306 B.n202 71.676
R974 B.n305 B.n304 71.676
R975 B.n298 B.n204 71.676
R976 B.n297 B.n296 71.676
R977 B.n290 B.n206 71.676
R978 B.n289 B.n288 71.676
R979 B.n282 B.n208 71.676
R980 B.n281 B.n280 71.676
R981 B.n274 B.n210 71.676
R982 B.n273 B.n272 71.676
R983 B.n266 B.n212 71.676
R984 B.n265 B.n264 71.676
R985 B.n258 B.n214 71.676
R986 B.n257 B.n256 71.676
R987 B.n250 B.n216 71.676
R988 B.n249 B.n248 71.676
R989 B.n242 B.n218 71.676
R990 B.n241 B.n240 71.676
R991 B.n234 B.n220 71.676
R992 B.n233 B.n232 71.676
R993 B.n226 B.n222 71.676
R994 B.n225 B.n224 71.676
R995 B.n474 B.n473 71.676
R996 B.n468 B.n158 71.676
R997 B.n466 B.n465 71.676
R998 B.n461 B.n460 71.676
R999 B.n458 B.n457 71.676
R1000 B.n453 B.n452 71.676
R1001 B.n450 B.n449 71.676
R1002 B.n445 B.n444 71.676
R1003 B.n442 B.n441 71.676
R1004 B.n437 B.n436 71.676
R1005 B.n434 B.n433 71.676
R1006 B.n429 B.n428 71.676
R1007 B.n426 B.n425 71.676
R1008 B.n421 B.n420 71.676
R1009 B.n418 B.n417 71.676
R1010 B.n413 B.n412 71.676
R1011 B.n410 B.n409 71.676
R1012 B.n405 B.n404 71.676
R1013 B.n402 B.n401 71.676
R1014 B.n397 B.n396 71.676
R1015 B.n394 B.n393 71.676
R1016 B.n389 B.n388 71.676
R1017 B.n386 B.n385 71.676
R1018 B.n381 B.n380 71.676
R1019 B.n378 B.n377 71.676
R1020 B.n373 B.n372 71.676
R1021 B.n370 B.n369 71.676
R1022 B.n365 B.n364 71.676
R1023 B.n362 B.n361 71.676
R1024 B.n356 B.n355 71.676
R1025 B.n353 B.n352 71.676
R1026 B.n348 B.n347 71.676
R1027 B.n345 B.n344 71.676
R1028 B.n339 B.n338 71.676
R1029 B.n336 B.n335 71.676
R1030 B.n331 B.n330 71.676
R1031 B.n328 B.n327 71.676
R1032 B.n323 B.n322 71.676
R1033 B.n320 B.n319 71.676
R1034 B.n315 B.n314 71.676
R1035 B.n312 B.n311 71.676
R1036 B.n307 B.n306 71.676
R1037 B.n304 B.n303 71.676
R1038 B.n299 B.n298 71.676
R1039 B.n296 B.n295 71.676
R1040 B.n291 B.n290 71.676
R1041 B.n288 B.n287 71.676
R1042 B.n283 B.n282 71.676
R1043 B.n280 B.n279 71.676
R1044 B.n275 B.n274 71.676
R1045 B.n272 B.n271 71.676
R1046 B.n267 B.n266 71.676
R1047 B.n264 B.n263 71.676
R1048 B.n259 B.n258 71.676
R1049 B.n256 B.n255 71.676
R1050 B.n251 B.n250 71.676
R1051 B.n248 B.n247 71.676
R1052 B.n243 B.n242 71.676
R1053 B.n240 B.n239 71.676
R1054 B.n235 B.n234 71.676
R1055 B.n232 B.n231 71.676
R1056 B.n227 B.n226 71.676
R1057 B.n224 B.n154 71.676
R1058 B.n876 B.n875 71.676
R1059 B.n876 B.n2 71.676
R1060 B.n84 B.t15 68.8148
R1061 B.n194 B.t4 68.8148
R1062 B.n77 B.t9 68.791
R1063 B.n188 B.t11 68.791
R1064 B.n479 B.n155 61.6024
R1065 B.n831 B.n44 61.6024
R1066 B.n78 B.n77 59.5399
R1067 B.n692 B.n84 59.5399
R1068 B.n341 B.n194 59.5399
R1069 B.n359 B.n188 59.5399
R1070 B.n77 B.n76 47.7096
R1071 B.n84 B.n83 47.7096
R1072 B.n194 B.n193 47.7096
R1073 B.n188 B.n187 47.7096
R1074 B.n479 B.n151 32.4728
R1075 B.n485 B.n151 32.4728
R1076 B.n485 B.n147 32.4728
R1077 B.n491 B.n147 32.4728
R1078 B.n491 B.n143 32.4728
R1079 B.n497 B.n143 32.4728
R1080 B.n503 B.n139 32.4728
R1081 B.n503 B.n135 32.4728
R1082 B.n509 B.n135 32.4728
R1083 B.n509 B.n131 32.4728
R1084 B.n515 B.n131 32.4728
R1085 B.n515 B.n127 32.4728
R1086 B.n521 B.n127 32.4728
R1087 B.n521 B.n122 32.4728
R1088 B.n527 B.n122 32.4728
R1089 B.n527 B.n123 32.4728
R1090 B.n534 B.n115 32.4728
R1091 B.n540 B.n115 32.4728
R1092 B.n540 B.n4 32.4728
R1093 B.n874 B.n4 32.4728
R1094 B.n874 B.n873 32.4728
R1095 B.n873 B.n872 32.4728
R1096 B.n872 B.n8 32.4728
R1097 B.n12 B.n8 32.4728
R1098 B.n865 B.n12 32.4728
R1099 B.n864 B.n863 32.4728
R1100 B.n863 B.n16 32.4728
R1101 B.n857 B.n16 32.4728
R1102 B.n857 B.n856 32.4728
R1103 B.n856 B.n855 32.4728
R1104 B.n855 B.n23 32.4728
R1105 B.n849 B.n23 32.4728
R1106 B.n849 B.n848 32.4728
R1107 B.n848 B.n847 32.4728
R1108 B.n847 B.n30 32.4728
R1109 B.n841 B.n840 32.4728
R1110 B.n840 B.n839 32.4728
R1111 B.n839 B.n37 32.4728
R1112 B.n833 B.n37 32.4728
R1113 B.n833 B.n832 32.4728
R1114 B.n832 B.n831 32.4728
R1115 B.n477 B.n476 31.6883
R1116 B.n481 B.n153 31.6883
R1117 B.n574 B.n573 31.6883
R1118 B.n829 B.n828 31.6883
R1119 B.n497 B.t3 27.2199
R1120 B.n841 B.t7 27.2199
R1121 B.n534 B.t1 23.3997
R1122 B.n865 B.t0 23.3997
R1123 B B.n877 18.0485
R1124 B.n477 B.n149 10.6151
R1125 B.n487 B.n149 10.6151
R1126 B.n488 B.n487 10.6151
R1127 B.n489 B.n488 10.6151
R1128 B.n489 B.n141 10.6151
R1129 B.n499 B.n141 10.6151
R1130 B.n500 B.n499 10.6151
R1131 B.n501 B.n500 10.6151
R1132 B.n501 B.n133 10.6151
R1133 B.n511 B.n133 10.6151
R1134 B.n512 B.n511 10.6151
R1135 B.n513 B.n512 10.6151
R1136 B.n513 B.n125 10.6151
R1137 B.n523 B.n125 10.6151
R1138 B.n524 B.n523 10.6151
R1139 B.n525 B.n524 10.6151
R1140 B.n525 B.n117 10.6151
R1141 B.n536 B.n117 10.6151
R1142 B.n537 B.n536 10.6151
R1143 B.n538 B.n537 10.6151
R1144 B.n538 B.n0 10.6151
R1145 B.n476 B.n475 10.6151
R1146 B.n475 B.n157 10.6151
R1147 B.n470 B.n157 10.6151
R1148 B.n470 B.n469 10.6151
R1149 B.n469 B.n159 10.6151
R1150 B.n464 B.n159 10.6151
R1151 B.n464 B.n463 10.6151
R1152 B.n463 B.n462 10.6151
R1153 B.n462 B.n161 10.6151
R1154 B.n456 B.n161 10.6151
R1155 B.n456 B.n455 10.6151
R1156 B.n455 B.n454 10.6151
R1157 B.n454 B.n163 10.6151
R1158 B.n448 B.n163 10.6151
R1159 B.n448 B.n447 10.6151
R1160 B.n447 B.n446 10.6151
R1161 B.n446 B.n165 10.6151
R1162 B.n440 B.n165 10.6151
R1163 B.n440 B.n439 10.6151
R1164 B.n439 B.n438 10.6151
R1165 B.n438 B.n167 10.6151
R1166 B.n432 B.n167 10.6151
R1167 B.n432 B.n431 10.6151
R1168 B.n431 B.n430 10.6151
R1169 B.n430 B.n169 10.6151
R1170 B.n424 B.n169 10.6151
R1171 B.n424 B.n423 10.6151
R1172 B.n423 B.n422 10.6151
R1173 B.n422 B.n171 10.6151
R1174 B.n416 B.n171 10.6151
R1175 B.n416 B.n415 10.6151
R1176 B.n415 B.n414 10.6151
R1177 B.n414 B.n173 10.6151
R1178 B.n408 B.n173 10.6151
R1179 B.n408 B.n407 10.6151
R1180 B.n407 B.n406 10.6151
R1181 B.n406 B.n175 10.6151
R1182 B.n400 B.n175 10.6151
R1183 B.n400 B.n399 10.6151
R1184 B.n399 B.n398 10.6151
R1185 B.n398 B.n177 10.6151
R1186 B.n392 B.n177 10.6151
R1187 B.n392 B.n391 10.6151
R1188 B.n391 B.n390 10.6151
R1189 B.n390 B.n179 10.6151
R1190 B.n384 B.n179 10.6151
R1191 B.n384 B.n383 10.6151
R1192 B.n383 B.n382 10.6151
R1193 B.n382 B.n181 10.6151
R1194 B.n376 B.n181 10.6151
R1195 B.n376 B.n375 10.6151
R1196 B.n375 B.n374 10.6151
R1197 B.n374 B.n183 10.6151
R1198 B.n368 B.n183 10.6151
R1199 B.n368 B.n367 10.6151
R1200 B.n367 B.n366 10.6151
R1201 B.n366 B.n185 10.6151
R1202 B.n360 B.n185 10.6151
R1203 B.n358 B.n357 10.6151
R1204 B.n357 B.n189 10.6151
R1205 B.n351 B.n189 10.6151
R1206 B.n351 B.n350 10.6151
R1207 B.n350 B.n349 10.6151
R1208 B.n349 B.n191 10.6151
R1209 B.n343 B.n191 10.6151
R1210 B.n343 B.n342 10.6151
R1211 B.n340 B.n195 10.6151
R1212 B.n334 B.n195 10.6151
R1213 B.n334 B.n333 10.6151
R1214 B.n333 B.n332 10.6151
R1215 B.n332 B.n197 10.6151
R1216 B.n326 B.n197 10.6151
R1217 B.n326 B.n325 10.6151
R1218 B.n325 B.n324 10.6151
R1219 B.n324 B.n199 10.6151
R1220 B.n318 B.n199 10.6151
R1221 B.n318 B.n317 10.6151
R1222 B.n317 B.n316 10.6151
R1223 B.n316 B.n201 10.6151
R1224 B.n310 B.n201 10.6151
R1225 B.n310 B.n309 10.6151
R1226 B.n309 B.n308 10.6151
R1227 B.n308 B.n203 10.6151
R1228 B.n302 B.n203 10.6151
R1229 B.n302 B.n301 10.6151
R1230 B.n301 B.n300 10.6151
R1231 B.n300 B.n205 10.6151
R1232 B.n294 B.n205 10.6151
R1233 B.n294 B.n293 10.6151
R1234 B.n293 B.n292 10.6151
R1235 B.n292 B.n207 10.6151
R1236 B.n286 B.n207 10.6151
R1237 B.n286 B.n285 10.6151
R1238 B.n285 B.n284 10.6151
R1239 B.n284 B.n209 10.6151
R1240 B.n278 B.n209 10.6151
R1241 B.n278 B.n277 10.6151
R1242 B.n277 B.n276 10.6151
R1243 B.n276 B.n211 10.6151
R1244 B.n270 B.n211 10.6151
R1245 B.n270 B.n269 10.6151
R1246 B.n269 B.n268 10.6151
R1247 B.n268 B.n213 10.6151
R1248 B.n262 B.n213 10.6151
R1249 B.n262 B.n261 10.6151
R1250 B.n261 B.n260 10.6151
R1251 B.n260 B.n215 10.6151
R1252 B.n254 B.n215 10.6151
R1253 B.n254 B.n253 10.6151
R1254 B.n253 B.n252 10.6151
R1255 B.n252 B.n217 10.6151
R1256 B.n246 B.n217 10.6151
R1257 B.n246 B.n245 10.6151
R1258 B.n245 B.n244 10.6151
R1259 B.n244 B.n219 10.6151
R1260 B.n238 B.n219 10.6151
R1261 B.n238 B.n237 10.6151
R1262 B.n237 B.n236 10.6151
R1263 B.n236 B.n221 10.6151
R1264 B.n230 B.n221 10.6151
R1265 B.n230 B.n229 10.6151
R1266 B.n229 B.n228 10.6151
R1267 B.n228 B.n223 10.6151
R1268 B.n223 B.n153 10.6151
R1269 B.n482 B.n481 10.6151
R1270 B.n483 B.n482 10.6151
R1271 B.n483 B.n145 10.6151
R1272 B.n493 B.n145 10.6151
R1273 B.n494 B.n493 10.6151
R1274 B.n495 B.n494 10.6151
R1275 B.n495 B.n137 10.6151
R1276 B.n505 B.n137 10.6151
R1277 B.n506 B.n505 10.6151
R1278 B.n507 B.n506 10.6151
R1279 B.n507 B.n129 10.6151
R1280 B.n517 B.n129 10.6151
R1281 B.n518 B.n517 10.6151
R1282 B.n519 B.n518 10.6151
R1283 B.n519 B.n120 10.6151
R1284 B.n529 B.n120 10.6151
R1285 B.n530 B.n529 10.6151
R1286 B.n532 B.n530 10.6151
R1287 B.n532 B.n531 10.6151
R1288 B.n531 B.n113 10.6151
R1289 B.n543 B.n113 10.6151
R1290 B.n544 B.n543 10.6151
R1291 B.n545 B.n544 10.6151
R1292 B.n546 B.n545 10.6151
R1293 B.n547 B.n546 10.6151
R1294 B.n550 B.n547 10.6151
R1295 B.n551 B.n550 10.6151
R1296 B.n552 B.n551 10.6151
R1297 B.n553 B.n552 10.6151
R1298 B.n555 B.n553 10.6151
R1299 B.n556 B.n555 10.6151
R1300 B.n557 B.n556 10.6151
R1301 B.n558 B.n557 10.6151
R1302 B.n560 B.n558 10.6151
R1303 B.n561 B.n560 10.6151
R1304 B.n562 B.n561 10.6151
R1305 B.n563 B.n562 10.6151
R1306 B.n565 B.n563 10.6151
R1307 B.n566 B.n565 10.6151
R1308 B.n567 B.n566 10.6151
R1309 B.n568 B.n567 10.6151
R1310 B.n570 B.n568 10.6151
R1311 B.n571 B.n570 10.6151
R1312 B.n572 B.n571 10.6151
R1313 B.n573 B.n572 10.6151
R1314 B.n869 B.n1 10.6151
R1315 B.n869 B.n868 10.6151
R1316 B.n868 B.n867 10.6151
R1317 B.n867 B.n10 10.6151
R1318 B.n861 B.n10 10.6151
R1319 B.n861 B.n860 10.6151
R1320 B.n860 B.n859 10.6151
R1321 B.n859 B.n18 10.6151
R1322 B.n853 B.n18 10.6151
R1323 B.n853 B.n852 10.6151
R1324 B.n852 B.n851 10.6151
R1325 B.n851 B.n25 10.6151
R1326 B.n845 B.n25 10.6151
R1327 B.n845 B.n844 10.6151
R1328 B.n844 B.n843 10.6151
R1329 B.n843 B.n32 10.6151
R1330 B.n837 B.n32 10.6151
R1331 B.n837 B.n836 10.6151
R1332 B.n836 B.n835 10.6151
R1333 B.n835 B.n39 10.6151
R1334 B.n829 B.n39 10.6151
R1335 B.n828 B.n827 10.6151
R1336 B.n827 B.n46 10.6151
R1337 B.n821 B.n46 10.6151
R1338 B.n821 B.n820 10.6151
R1339 B.n820 B.n819 10.6151
R1340 B.n819 B.n48 10.6151
R1341 B.n813 B.n48 10.6151
R1342 B.n813 B.n812 10.6151
R1343 B.n812 B.n811 10.6151
R1344 B.n811 B.n50 10.6151
R1345 B.n805 B.n50 10.6151
R1346 B.n805 B.n804 10.6151
R1347 B.n804 B.n803 10.6151
R1348 B.n803 B.n52 10.6151
R1349 B.n797 B.n52 10.6151
R1350 B.n797 B.n796 10.6151
R1351 B.n796 B.n795 10.6151
R1352 B.n795 B.n54 10.6151
R1353 B.n789 B.n54 10.6151
R1354 B.n789 B.n788 10.6151
R1355 B.n788 B.n787 10.6151
R1356 B.n787 B.n56 10.6151
R1357 B.n781 B.n56 10.6151
R1358 B.n781 B.n780 10.6151
R1359 B.n780 B.n779 10.6151
R1360 B.n779 B.n58 10.6151
R1361 B.n773 B.n58 10.6151
R1362 B.n773 B.n772 10.6151
R1363 B.n772 B.n771 10.6151
R1364 B.n771 B.n60 10.6151
R1365 B.n765 B.n60 10.6151
R1366 B.n765 B.n764 10.6151
R1367 B.n764 B.n763 10.6151
R1368 B.n763 B.n62 10.6151
R1369 B.n757 B.n62 10.6151
R1370 B.n757 B.n756 10.6151
R1371 B.n756 B.n755 10.6151
R1372 B.n755 B.n64 10.6151
R1373 B.n749 B.n64 10.6151
R1374 B.n749 B.n748 10.6151
R1375 B.n748 B.n747 10.6151
R1376 B.n747 B.n66 10.6151
R1377 B.n741 B.n66 10.6151
R1378 B.n741 B.n740 10.6151
R1379 B.n740 B.n739 10.6151
R1380 B.n739 B.n68 10.6151
R1381 B.n733 B.n68 10.6151
R1382 B.n733 B.n732 10.6151
R1383 B.n732 B.n731 10.6151
R1384 B.n731 B.n70 10.6151
R1385 B.n725 B.n70 10.6151
R1386 B.n725 B.n724 10.6151
R1387 B.n724 B.n723 10.6151
R1388 B.n723 B.n72 10.6151
R1389 B.n717 B.n72 10.6151
R1390 B.n717 B.n716 10.6151
R1391 B.n716 B.n715 10.6151
R1392 B.n715 B.n74 10.6151
R1393 B.n709 B.n708 10.6151
R1394 B.n708 B.n707 10.6151
R1395 B.n707 B.n79 10.6151
R1396 B.n701 B.n79 10.6151
R1397 B.n701 B.n700 10.6151
R1398 B.n700 B.n699 10.6151
R1399 B.n699 B.n81 10.6151
R1400 B.n693 B.n81 10.6151
R1401 B.n691 B.n690 10.6151
R1402 B.n690 B.n85 10.6151
R1403 B.n684 B.n85 10.6151
R1404 B.n684 B.n683 10.6151
R1405 B.n683 B.n682 10.6151
R1406 B.n682 B.n87 10.6151
R1407 B.n676 B.n87 10.6151
R1408 B.n676 B.n675 10.6151
R1409 B.n675 B.n674 10.6151
R1410 B.n674 B.n89 10.6151
R1411 B.n668 B.n89 10.6151
R1412 B.n668 B.n667 10.6151
R1413 B.n667 B.n666 10.6151
R1414 B.n666 B.n91 10.6151
R1415 B.n660 B.n91 10.6151
R1416 B.n660 B.n659 10.6151
R1417 B.n659 B.n658 10.6151
R1418 B.n658 B.n93 10.6151
R1419 B.n652 B.n93 10.6151
R1420 B.n652 B.n651 10.6151
R1421 B.n651 B.n650 10.6151
R1422 B.n650 B.n95 10.6151
R1423 B.n644 B.n95 10.6151
R1424 B.n644 B.n643 10.6151
R1425 B.n643 B.n642 10.6151
R1426 B.n642 B.n97 10.6151
R1427 B.n636 B.n97 10.6151
R1428 B.n636 B.n635 10.6151
R1429 B.n635 B.n634 10.6151
R1430 B.n634 B.n99 10.6151
R1431 B.n628 B.n99 10.6151
R1432 B.n628 B.n627 10.6151
R1433 B.n627 B.n626 10.6151
R1434 B.n626 B.n101 10.6151
R1435 B.n620 B.n101 10.6151
R1436 B.n620 B.n619 10.6151
R1437 B.n619 B.n618 10.6151
R1438 B.n618 B.n103 10.6151
R1439 B.n612 B.n103 10.6151
R1440 B.n612 B.n611 10.6151
R1441 B.n611 B.n610 10.6151
R1442 B.n610 B.n105 10.6151
R1443 B.n604 B.n105 10.6151
R1444 B.n604 B.n603 10.6151
R1445 B.n603 B.n602 10.6151
R1446 B.n602 B.n107 10.6151
R1447 B.n596 B.n107 10.6151
R1448 B.n596 B.n595 10.6151
R1449 B.n595 B.n594 10.6151
R1450 B.n594 B.n109 10.6151
R1451 B.n588 B.n109 10.6151
R1452 B.n588 B.n587 10.6151
R1453 B.n587 B.n586 10.6151
R1454 B.n586 B.n111 10.6151
R1455 B.n580 B.n111 10.6151
R1456 B.n580 B.n579 10.6151
R1457 B.n579 B.n578 10.6151
R1458 B.n578 B.n574 10.6151
R1459 B.n123 B.t1 9.07365
R1460 B.t0 B.n864 9.07365
R1461 B.n877 B.n0 8.11757
R1462 B.n877 B.n1 8.11757
R1463 B.n359 B.n358 6.5566
R1464 B.n342 B.n341 6.5566
R1465 B.n709 B.n78 6.5566
R1466 B.n693 B.n692 6.5566
R1467 B.t3 B.n139 5.25338
R1468 B.t7 B.n30 5.25338
R1469 B.n360 B.n359 4.05904
R1470 B.n341 B.n340 4.05904
R1471 B.n78 B.n74 4.05904
R1472 B.n692 B.n691 4.05904
R1473 VP.n0 VP.t1 297.846
R1474 VP.n0 VP.t0 250.073
R1475 VP VP.n0 0.336784
R1476 VDD1 VDD1.t1 103.718
R1477 VDD1 VDD1.t0 60.0397
C0 VTAIL VDD2 6.64856f
C1 VTAIL VDD1 6.60329f
C2 VDD2 VP 0.31355f
C3 VDD1 VP 4.02401f
C4 VDD2 VN 3.86201f
C5 VN VDD1 0.147572f
C6 VDD2 VDD1 0.619414f
C7 VTAIL VP 3.24363f
C8 VTAIL VN 3.22919f
C9 VN VP 6.3086f
C10 VDD2 B 5.300968f
C11 VDD1 B 8.73683f
C12 VTAIL B 9.435796f
C13 VN B 11.71732f
C14 VP B 6.215725f
C15 VDD1.t0 B 3.25735f
C16 VDD1.t1 B 3.99015f
C17 VP.t1 B 4.2525f
C18 VP.t0 B 3.77778f
C19 VP.n0 B 5.40371f
C20 VDD2.t1 B 3.94318f
C21 VDD2.t0 B 3.24657f
C22 VDD2.n0 B 3.20393f
C23 VTAIL.t1 B 3.09778f
C24 VTAIL.n0 B 1.83921f
C25 VTAIL.t3 B 3.09779f
C26 VTAIL.n1 B 1.86889f
C27 VTAIL.t0 B 3.09778f
C28 VTAIL.n2 B 1.73554f
C29 VTAIL.t2 B 3.09778f
C30 VTAIL.n3 B 1.66901f
C31 VN.t0 B 3.73837f
C32 VN.t1 B 4.20887f
.ends

