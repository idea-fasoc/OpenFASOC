* NGSPICE file created from diff_pair_sample_1015.ext - technology: sky130A

.subckt diff_pair_sample_1015 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t3 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=1.7199 pd=9.6 as=0.72765 ps=4.74 w=4.41 l=1.41
X1 VTAIL.t14 VN.t1 VDD2.t5 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=0.72765 ps=4.74 w=4.41 l=1.41
X2 VTAIL.t6 VP.t0 VDD1.t7 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=1.7199 pd=9.6 as=0.72765 ps=4.74 w=4.41 l=1.41
X3 VTAIL.t5 VP.t1 VDD1.t6 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=1.7199 pd=9.6 as=0.72765 ps=4.74 w=4.41 l=1.41
X4 VDD2.t0 VN.t2 VTAIL.t13 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=1.7199 ps=9.6 w=4.41 l=1.41
X5 VDD1.t5 VP.t2 VTAIL.t1 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=0.72765 ps=4.74 w=4.41 l=1.41
X6 VDD2.t4 VN.t3 VTAIL.t12 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=1.7199 ps=9.6 w=4.41 l=1.41
X7 VTAIL.t2 VP.t3 VDD1.t4 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=0.72765 ps=4.74 w=4.41 l=1.41
X8 VTAIL.t11 VN.t4 VDD2.t6 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=1.7199 pd=9.6 as=0.72765 ps=4.74 w=4.41 l=1.41
X9 B.t11 B.t9 B.t10 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=1.7199 pd=9.6 as=0 ps=0 w=4.41 l=1.41
X10 VDD2.t7 VN.t5 VTAIL.t10 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=0.72765 ps=4.74 w=4.41 l=1.41
X11 VDD1.t3 VP.t4 VTAIL.t4 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=1.7199 ps=9.6 w=4.41 l=1.41
X12 B.t8 B.t6 B.t7 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=1.7199 pd=9.6 as=0 ps=0 w=4.41 l=1.41
X13 VTAIL.t7 VP.t5 VDD1.t2 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=0.72765 ps=4.74 w=4.41 l=1.41
X14 B.t5 B.t3 B.t4 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=1.7199 pd=9.6 as=0 ps=0 w=4.41 l=1.41
X15 VDD2.t1 VN.t6 VTAIL.t9 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=0.72765 ps=4.74 w=4.41 l=1.41
X16 VDD1.t1 VP.t6 VTAIL.t3 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=0.72765 ps=4.74 w=4.41 l=1.41
X17 VTAIL.t8 VN.t7 VDD2.t2 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=0.72765 ps=4.74 w=4.41 l=1.41
X18 B.t2 B.t0 B.t1 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=1.7199 pd=9.6 as=0 ps=0 w=4.41 l=1.41
X19 VDD1.t0 VP.t7 VTAIL.t0 w_n2710_n1850# sky130_fd_pr__pfet_01v8 ad=0.72765 pd=4.74 as=1.7199 ps=9.6 w=4.41 l=1.41
R0 VN.n18 VN.n17 180.385
R1 VN.n37 VN.n36 180.385
R2 VN.n35 VN.n19 161.3
R3 VN.n34 VN.n33 161.3
R4 VN.n32 VN.n20 161.3
R5 VN.n31 VN.n30 161.3
R6 VN.n28 VN.n21 161.3
R7 VN.n27 VN.n26 161.3
R8 VN.n25 VN.n22 161.3
R9 VN.n16 VN.n0 161.3
R10 VN.n15 VN.n14 161.3
R11 VN.n13 VN.n1 161.3
R12 VN.n12 VN.n11 161.3
R13 VN.n9 VN.n2 161.3
R14 VN.n8 VN.n7 161.3
R15 VN.n6 VN.n3 161.3
R16 VN.n5 VN.t4 106.62
R17 VN.n24 VN.t3 106.62
R18 VN.n4 VN.t5 75.3771
R19 VN.n10 VN.t1 75.3771
R20 VN.n17 VN.t2 75.3771
R21 VN.n23 VN.t7 75.3771
R22 VN.n29 VN.t6 75.3771
R23 VN.n36 VN.t0 75.3771
R24 VN.n15 VN.n1 56.5193
R25 VN.n34 VN.n20 56.5193
R26 VN.n5 VN.n4 47.8106
R27 VN.n24 VN.n23 47.8106
R28 VN.n8 VN.n3 40.4934
R29 VN.n9 VN.n8 40.4934
R30 VN.n27 VN.n22 40.4934
R31 VN.n28 VN.n27 40.4934
R32 VN VN.n37 39.7903
R33 VN.n11 VN.n1 24.4675
R34 VN.n16 VN.n15 24.4675
R35 VN.n30 VN.n20 24.4675
R36 VN.n35 VN.n34 24.4675
R37 VN.n25 VN.n24 18.2406
R38 VN.n6 VN.n5 18.2406
R39 VN.n4 VN.n3 18.1061
R40 VN.n10 VN.n9 18.1061
R41 VN.n23 VN.n22 18.1061
R42 VN.n29 VN.n28 18.1061
R43 VN.n11 VN.n10 6.36192
R44 VN.n30 VN.n29 6.36192
R45 VN.n17 VN.n16 5.38324
R46 VN.n36 VN.n35 5.38324
R47 VN.n37 VN.n19 0.189894
R48 VN.n33 VN.n19 0.189894
R49 VN.n33 VN.n32 0.189894
R50 VN.n32 VN.n31 0.189894
R51 VN.n31 VN.n21 0.189894
R52 VN.n26 VN.n21 0.189894
R53 VN.n26 VN.n25 0.189894
R54 VN.n7 VN.n6 0.189894
R55 VN.n7 VN.n2 0.189894
R56 VN.n12 VN.n2 0.189894
R57 VN.n13 VN.n12 0.189894
R58 VN.n14 VN.n13 0.189894
R59 VN.n14 VN.n0 0.189894
R60 VN.n18 VN.n0 0.189894
R61 VN VN.n18 0.0516364
R62 VDD2.n2 VDD2.n1 113.153
R63 VDD2.n2 VDD2.n0 113.153
R64 VDD2 VDD2.n5 113.151
R65 VDD2.n4 VDD2.n3 112.46
R66 VDD2.n4 VDD2.n2 34.267
R67 VDD2.n5 VDD2.t2 7.37125
R68 VDD2.n5 VDD2.t4 7.37125
R69 VDD2.n3 VDD2.t3 7.37125
R70 VDD2.n3 VDD2.t1 7.37125
R71 VDD2.n1 VDD2.t5 7.37125
R72 VDD2.n1 VDD2.t0 7.37125
R73 VDD2.n0 VDD2.t6 7.37125
R74 VDD2.n0 VDD2.t7 7.37125
R75 VDD2 VDD2.n4 0.80869
R76 VTAIL.n11 VTAIL.t5 103.151
R77 VTAIL.n10 VTAIL.t12 103.151
R78 VTAIL.n7 VTAIL.t15 103.151
R79 VTAIL.n15 VTAIL.t13 103.151
R80 VTAIL.n2 VTAIL.t11 103.151
R81 VTAIL.n3 VTAIL.t4 103.151
R82 VTAIL.n6 VTAIL.t6 103.151
R83 VTAIL.n14 VTAIL.t0 103.151
R84 VTAIL.n13 VTAIL.n12 95.7806
R85 VTAIL.n9 VTAIL.n8 95.7806
R86 VTAIL.n1 VTAIL.n0 95.7803
R87 VTAIL.n5 VTAIL.n4 95.7803
R88 VTAIL.n15 VTAIL.n14 17.6686
R89 VTAIL.n7 VTAIL.n6 17.6686
R90 VTAIL.n0 VTAIL.t10 7.37125
R91 VTAIL.n0 VTAIL.t14 7.37125
R92 VTAIL.n4 VTAIL.t1 7.37125
R93 VTAIL.n4 VTAIL.t7 7.37125
R94 VTAIL.n12 VTAIL.t3 7.37125
R95 VTAIL.n12 VTAIL.t2 7.37125
R96 VTAIL.n8 VTAIL.t9 7.37125
R97 VTAIL.n8 VTAIL.t8 7.37125
R98 VTAIL.n9 VTAIL.n7 1.5005
R99 VTAIL.n10 VTAIL.n9 1.5005
R100 VTAIL.n13 VTAIL.n11 1.5005
R101 VTAIL.n14 VTAIL.n13 1.5005
R102 VTAIL.n6 VTAIL.n5 1.5005
R103 VTAIL.n5 VTAIL.n3 1.5005
R104 VTAIL.n2 VTAIL.n1 1.5005
R105 VTAIL VTAIL.n15 1.44231
R106 VTAIL.n11 VTAIL.n10 0.470328
R107 VTAIL.n3 VTAIL.n2 0.470328
R108 VTAIL VTAIL.n1 0.0586897
R109 VP.n26 VP.n25 180.385
R110 VP.n46 VP.n45 180.385
R111 VP.n24 VP.n23 180.385
R112 VP.n12 VP.n9 161.3
R113 VP.n14 VP.n13 161.3
R114 VP.n15 VP.n8 161.3
R115 VP.n18 VP.n17 161.3
R116 VP.n19 VP.n7 161.3
R117 VP.n21 VP.n20 161.3
R118 VP.n22 VP.n6 161.3
R119 VP.n44 VP.n0 161.3
R120 VP.n43 VP.n42 161.3
R121 VP.n41 VP.n1 161.3
R122 VP.n40 VP.n39 161.3
R123 VP.n37 VP.n2 161.3
R124 VP.n36 VP.n35 161.3
R125 VP.n34 VP.n3 161.3
R126 VP.n33 VP.n32 161.3
R127 VP.n30 VP.n4 161.3
R128 VP.n29 VP.n28 161.3
R129 VP.n27 VP.n5 161.3
R130 VP.n11 VP.t1 106.62
R131 VP.n25 VP.t0 75.3771
R132 VP.n31 VP.t2 75.3771
R133 VP.n38 VP.t5 75.3771
R134 VP.n45 VP.t4 75.3771
R135 VP.n23 VP.t7 75.3771
R136 VP.n16 VP.t3 75.3771
R137 VP.n10 VP.t6 75.3771
R138 VP.n30 VP.n29 56.5193
R139 VP.n43 VP.n1 56.5193
R140 VP.n21 VP.n7 56.5193
R141 VP.n11 VP.n10 47.8106
R142 VP.n36 VP.n3 40.4934
R143 VP.n37 VP.n36 40.4934
R144 VP.n15 VP.n14 40.4934
R145 VP.n14 VP.n9 40.4934
R146 VP.n26 VP.n24 39.4096
R147 VP.n29 VP.n5 24.4675
R148 VP.n32 VP.n30 24.4675
R149 VP.n39 VP.n1 24.4675
R150 VP.n44 VP.n43 24.4675
R151 VP.n22 VP.n21 24.4675
R152 VP.n17 VP.n7 24.4675
R153 VP.n12 VP.n11 18.2406
R154 VP.n31 VP.n3 18.1061
R155 VP.n38 VP.n37 18.1061
R156 VP.n16 VP.n15 18.1061
R157 VP.n10 VP.n9 18.1061
R158 VP.n32 VP.n31 6.36192
R159 VP.n39 VP.n38 6.36192
R160 VP.n17 VP.n16 6.36192
R161 VP.n25 VP.n5 5.38324
R162 VP.n45 VP.n44 5.38324
R163 VP.n23 VP.n22 5.38324
R164 VP.n13 VP.n12 0.189894
R165 VP.n13 VP.n8 0.189894
R166 VP.n18 VP.n8 0.189894
R167 VP.n19 VP.n18 0.189894
R168 VP.n20 VP.n19 0.189894
R169 VP.n20 VP.n6 0.189894
R170 VP.n24 VP.n6 0.189894
R171 VP.n27 VP.n26 0.189894
R172 VP.n28 VP.n27 0.189894
R173 VP.n28 VP.n4 0.189894
R174 VP.n33 VP.n4 0.189894
R175 VP.n34 VP.n33 0.189894
R176 VP.n35 VP.n34 0.189894
R177 VP.n35 VP.n2 0.189894
R178 VP.n40 VP.n2 0.189894
R179 VP.n41 VP.n40 0.189894
R180 VP.n42 VP.n41 0.189894
R181 VP.n42 VP.n0 0.189894
R182 VP.n46 VP.n0 0.189894
R183 VP VP.n46 0.0516364
R184 VDD1 VDD1.n0 113.267
R185 VDD1.n3 VDD1.n2 113.153
R186 VDD1.n3 VDD1.n1 113.153
R187 VDD1.n5 VDD1.n4 112.46
R188 VDD1.n5 VDD1.n3 34.85
R189 VDD1.n4 VDD1.t4 7.37125
R190 VDD1.n4 VDD1.t0 7.37125
R191 VDD1.n0 VDD1.t6 7.37125
R192 VDD1.n0 VDD1.t1 7.37125
R193 VDD1.n2 VDD1.t2 7.37125
R194 VDD1.n2 VDD1.t3 7.37125
R195 VDD1.n1 VDD1.t7 7.37125
R196 VDD1.n1 VDD1.t5 7.37125
R197 VDD1 VDD1.n5 0.69231
R198 B.n246 B.n81 585
R199 B.n245 B.n244 585
R200 B.n243 B.n82 585
R201 B.n242 B.n241 585
R202 B.n240 B.n83 585
R203 B.n239 B.n238 585
R204 B.n237 B.n84 585
R205 B.n236 B.n235 585
R206 B.n234 B.n85 585
R207 B.n233 B.n232 585
R208 B.n231 B.n86 585
R209 B.n230 B.n229 585
R210 B.n228 B.n87 585
R211 B.n227 B.n226 585
R212 B.n225 B.n88 585
R213 B.n224 B.n223 585
R214 B.n222 B.n89 585
R215 B.n221 B.n220 585
R216 B.n219 B.n90 585
R217 B.n218 B.n217 585
R218 B.n213 B.n91 585
R219 B.n212 B.n211 585
R220 B.n210 B.n92 585
R221 B.n209 B.n208 585
R222 B.n207 B.n93 585
R223 B.n206 B.n205 585
R224 B.n204 B.n94 585
R225 B.n203 B.n202 585
R226 B.n201 B.n95 585
R227 B.n199 B.n198 585
R228 B.n197 B.n98 585
R229 B.n196 B.n195 585
R230 B.n194 B.n99 585
R231 B.n193 B.n192 585
R232 B.n191 B.n100 585
R233 B.n190 B.n189 585
R234 B.n188 B.n101 585
R235 B.n187 B.n186 585
R236 B.n185 B.n102 585
R237 B.n184 B.n183 585
R238 B.n182 B.n103 585
R239 B.n181 B.n180 585
R240 B.n179 B.n104 585
R241 B.n178 B.n177 585
R242 B.n176 B.n105 585
R243 B.n175 B.n174 585
R244 B.n173 B.n106 585
R245 B.n172 B.n171 585
R246 B.n248 B.n247 585
R247 B.n249 B.n80 585
R248 B.n251 B.n250 585
R249 B.n252 B.n79 585
R250 B.n254 B.n253 585
R251 B.n255 B.n78 585
R252 B.n257 B.n256 585
R253 B.n258 B.n77 585
R254 B.n260 B.n259 585
R255 B.n261 B.n76 585
R256 B.n263 B.n262 585
R257 B.n264 B.n75 585
R258 B.n266 B.n265 585
R259 B.n267 B.n74 585
R260 B.n269 B.n268 585
R261 B.n270 B.n73 585
R262 B.n272 B.n271 585
R263 B.n273 B.n72 585
R264 B.n275 B.n274 585
R265 B.n276 B.n71 585
R266 B.n278 B.n277 585
R267 B.n279 B.n70 585
R268 B.n281 B.n280 585
R269 B.n282 B.n69 585
R270 B.n284 B.n283 585
R271 B.n285 B.n68 585
R272 B.n287 B.n286 585
R273 B.n288 B.n67 585
R274 B.n290 B.n289 585
R275 B.n291 B.n66 585
R276 B.n293 B.n292 585
R277 B.n294 B.n65 585
R278 B.n296 B.n295 585
R279 B.n297 B.n64 585
R280 B.n299 B.n298 585
R281 B.n300 B.n63 585
R282 B.n302 B.n301 585
R283 B.n303 B.n62 585
R284 B.n305 B.n304 585
R285 B.n306 B.n61 585
R286 B.n308 B.n307 585
R287 B.n309 B.n60 585
R288 B.n311 B.n310 585
R289 B.n312 B.n59 585
R290 B.n314 B.n313 585
R291 B.n315 B.n58 585
R292 B.n317 B.n316 585
R293 B.n318 B.n57 585
R294 B.n320 B.n319 585
R295 B.n321 B.n56 585
R296 B.n323 B.n322 585
R297 B.n324 B.n55 585
R298 B.n326 B.n325 585
R299 B.n327 B.n54 585
R300 B.n329 B.n328 585
R301 B.n330 B.n53 585
R302 B.n332 B.n331 585
R303 B.n333 B.n52 585
R304 B.n335 B.n334 585
R305 B.n336 B.n51 585
R306 B.n338 B.n337 585
R307 B.n339 B.n50 585
R308 B.n341 B.n340 585
R309 B.n342 B.n49 585
R310 B.n344 B.n343 585
R311 B.n345 B.n48 585
R312 B.n347 B.n346 585
R313 B.n348 B.n47 585
R314 B.n422 B.n421 585
R315 B.n420 B.n19 585
R316 B.n419 B.n418 585
R317 B.n417 B.n20 585
R318 B.n416 B.n415 585
R319 B.n414 B.n21 585
R320 B.n413 B.n412 585
R321 B.n411 B.n22 585
R322 B.n410 B.n409 585
R323 B.n408 B.n23 585
R324 B.n407 B.n406 585
R325 B.n405 B.n24 585
R326 B.n404 B.n403 585
R327 B.n402 B.n25 585
R328 B.n401 B.n400 585
R329 B.n399 B.n26 585
R330 B.n398 B.n397 585
R331 B.n396 B.n27 585
R332 B.n395 B.n394 585
R333 B.n393 B.n392 585
R334 B.n391 B.n31 585
R335 B.n390 B.n389 585
R336 B.n388 B.n32 585
R337 B.n387 B.n386 585
R338 B.n385 B.n33 585
R339 B.n384 B.n383 585
R340 B.n382 B.n34 585
R341 B.n381 B.n380 585
R342 B.n379 B.n35 585
R343 B.n377 B.n376 585
R344 B.n375 B.n38 585
R345 B.n374 B.n373 585
R346 B.n372 B.n39 585
R347 B.n371 B.n370 585
R348 B.n369 B.n40 585
R349 B.n368 B.n367 585
R350 B.n366 B.n41 585
R351 B.n365 B.n364 585
R352 B.n363 B.n42 585
R353 B.n362 B.n361 585
R354 B.n360 B.n43 585
R355 B.n359 B.n358 585
R356 B.n357 B.n44 585
R357 B.n356 B.n355 585
R358 B.n354 B.n45 585
R359 B.n353 B.n352 585
R360 B.n351 B.n46 585
R361 B.n350 B.n349 585
R362 B.n423 B.n18 585
R363 B.n425 B.n424 585
R364 B.n426 B.n17 585
R365 B.n428 B.n427 585
R366 B.n429 B.n16 585
R367 B.n431 B.n430 585
R368 B.n432 B.n15 585
R369 B.n434 B.n433 585
R370 B.n435 B.n14 585
R371 B.n437 B.n436 585
R372 B.n438 B.n13 585
R373 B.n440 B.n439 585
R374 B.n441 B.n12 585
R375 B.n443 B.n442 585
R376 B.n444 B.n11 585
R377 B.n446 B.n445 585
R378 B.n447 B.n10 585
R379 B.n449 B.n448 585
R380 B.n450 B.n9 585
R381 B.n452 B.n451 585
R382 B.n453 B.n8 585
R383 B.n455 B.n454 585
R384 B.n456 B.n7 585
R385 B.n458 B.n457 585
R386 B.n459 B.n6 585
R387 B.n461 B.n460 585
R388 B.n462 B.n5 585
R389 B.n464 B.n463 585
R390 B.n465 B.n4 585
R391 B.n467 B.n466 585
R392 B.n468 B.n3 585
R393 B.n470 B.n469 585
R394 B.n471 B.n0 585
R395 B.n2 B.n1 585
R396 B.n124 B.n123 585
R397 B.n125 B.n122 585
R398 B.n127 B.n126 585
R399 B.n128 B.n121 585
R400 B.n130 B.n129 585
R401 B.n131 B.n120 585
R402 B.n133 B.n132 585
R403 B.n134 B.n119 585
R404 B.n136 B.n135 585
R405 B.n137 B.n118 585
R406 B.n139 B.n138 585
R407 B.n140 B.n117 585
R408 B.n142 B.n141 585
R409 B.n143 B.n116 585
R410 B.n145 B.n144 585
R411 B.n146 B.n115 585
R412 B.n148 B.n147 585
R413 B.n149 B.n114 585
R414 B.n151 B.n150 585
R415 B.n152 B.n113 585
R416 B.n154 B.n153 585
R417 B.n155 B.n112 585
R418 B.n157 B.n156 585
R419 B.n158 B.n111 585
R420 B.n160 B.n159 585
R421 B.n161 B.n110 585
R422 B.n163 B.n162 585
R423 B.n164 B.n109 585
R424 B.n166 B.n165 585
R425 B.n167 B.n108 585
R426 B.n169 B.n168 585
R427 B.n170 B.n107 585
R428 B.n172 B.n107 545.355
R429 B.n248 B.n81 545.355
R430 B.n350 B.n47 545.355
R431 B.n423 B.n422 545.355
R432 B.n96 B.t0 280.466
R433 B.n214 B.t6 280.466
R434 B.n36 B.t3 280.466
R435 B.n28 B.t9 280.466
R436 B.n473 B.n472 256.663
R437 B.n472 B.n471 235.042
R438 B.n472 B.n2 235.042
R439 B.n173 B.n172 163.367
R440 B.n174 B.n173 163.367
R441 B.n174 B.n105 163.367
R442 B.n178 B.n105 163.367
R443 B.n179 B.n178 163.367
R444 B.n180 B.n179 163.367
R445 B.n180 B.n103 163.367
R446 B.n184 B.n103 163.367
R447 B.n185 B.n184 163.367
R448 B.n186 B.n185 163.367
R449 B.n186 B.n101 163.367
R450 B.n190 B.n101 163.367
R451 B.n191 B.n190 163.367
R452 B.n192 B.n191 163.367
R453 B.n192 B.n99 163.367
R454 B.n196 B.n99 163.367
R455 B.n197 B.n196 163.367
R456 B.n198 B.n197 163.367
R457 B.n198 B.n95 163.367
R458 B.n203 B.n95 163.367
R459 B.n204 B.n203 163.367
R460 B.n205 B.n204 163.367
R461 B.n205 B.n93 163.367
R462 B.n209 B.n93 163.367
R463 B.n210 B.n209 163.367
R464 B.n211 B.n210 163.367
R465 B.n211 B.n91 163.367
R466 B.n218 B.n91 163.367
R467 B.n219 B.n218 163.367
R468 B.n220 B.n219 163.367
R469 B.n220 B.n89 163.367
R470 B.n224 B.n89 163.367
R471 B.n225 B.n224 163.367
R472 B.n226 B.n225 163.367
R473 B.n226 B.n87 163.367
R474 B.n230 B.n87 163.367
R475 B.n231 B.n230 163.367
R476 B.n232 B.n231 163.367
R477 B.n232 B.n85 163.367
R478 B.n236 B.n85 163.367
R479 B.n237 B.n236 163.367
R480 B.n238 B.n237 163.367
R481 B.n238 B.n83 163.367
R482 B.n242 B.n83 163.367
R483 B.n243 B.n242 163.367
R484 B.n244 B.n243 163.367
R485 B.n244 B.n81 163.367
R486 B.n346 B.n47 163.367
R487 B.n346 B.n345 163.367
R488 B.n345 B.n344 163.367
R489 B.n344 B.n49 163.367
R490 B.n340 B.n49 163.367
R491 B.n340 B.n339 163.367
R492 B.n339 B.n338 163.367
R493 B.n338 B.n51 163.367
R494 B.n334 B.n51 163.367
R495 B.n334 B.n333 163.367
R496 B.n333 B.n332 163.367
R497 B.n332 B.n53 163.367
R498 B.n328 B.n53 163.367
R499 B.n328 B.n327 163.367
R500 B.n327 B.n326 163.367
R501 B.n326 B.n55 163.367
R502 B.n322 B.n55 163.367
R503 B.n322 B.n321 163.367
R504 B.n321 B.n320 163.367
R505 B.n320 B.n57 163.367
R506 B.n316 B.n57 163.367
R507 B.n316 B.n315 163.367
R508 B.n315 B.n314 163.367
R509 B.n314 B.n59 163.367
R510 B.n310 B.n59 163.367
R511 B.n310 B.n309 163.367
R512 B.n309 B.n308 163.367
R513 B.n308 B.n61 163.367
R514 B.n304 B.n61 163.367
R515 B.n304 B.n303 163.367
R516 B.n303 B.n302 163.367
R517 B.n302 B.n63 163.367
R518 B.n298 B.n63 163.367
R519 B.n298 B.n297 163.367
R520 B.n297 B.n296 163.367
R521 B.n296 B.n65 163.367
R522 B.n292 B.n65 163.367
R523 B.n292 B.n291 163.367
R524 B.n291 B.n290 163.367
R525 B.n290 B.n67 163.367
R526 B.n286 B.n67 163.367
R527 B.n286 B.n285 163.367
R528 B.n285 B.n284 163.367
R529 B.n284 B.n69 163.367
R530 B.n280 B.n69 163.367
R531 B.n280 B.n279 163.367
R532 B.n279 B.n278 163.367
R533 B.n278 B.n71 163.367
R534 B.n274 B.n71 163.367
R535 B.n274 B.n273 163.367
R536 B.n273 B.n272 163.367
R537 B.n272 B.n73 163.367
R538 B.n268 B.n73 163.367
R539 B.n268 B.n267 163.367
R540 B.n267 B.n266 163.367
R541 B.n266 B.n75 163.367
R542 B.n262 B.n75 163.367
R543 B.n262 B.n261 163.367
R544 B.n261 B.n260 163.367
R545 B.n260 B.n77 163.367
R546 B.n256 B.n77 163.367
R547 B.n256 B.n255 163.367
R548 B.n255 B.n254 163.367
R549 B.n254 B.n79 163.367
R550 B.n250 B.n79 163.367
R551 B.n250 B.n249 163.367
R552 B.n249 B.n248 163.367
R553 B.n422 B.n19 163.367
R554 B.n418 B.n19 163.367
R555 B.n418 B.n417 163.367
R556 B.n417 B.n416 163.367
R557 B.n416 B.n21 163.367
R558 B.n412 B.n21 163.367
R559 B.n412 B.n411 163.367
R560 B.n411 B.n410 163.367
R561 B.n410 B.n23 163.367
R562 B.n406 B.n23 163.367
R563 B.n406 B.n405 163.367
R564 B.n405 B.n404 163.367
R565 B.n404 B.n25 163.367
R566 B.n400 B.n25 163.367
R567 B.n400 B.n399 163.367
R568 B.n399 B.n398 163.367
R569 B.n398 B.n27 163.367
R570 B.n394 B.n27 163.367
R571 B.n394 B.n393 163.367
R572 B.n393 B.n31 163.367
R573 B.n389 B.n31 163.367
R574 B.n389 B.n388 163.367
R575 B.n388 B.n387 163.367
R576 B.n387 B.n33 163.367
R577 B.n383 B.n33 163.367
R578 B.n383 B.n382 163.367
R579 B.n382 B.n381 163.367
R580 B.n381 B.n35 163.367
R581 B.n376 B.n35 163.367
R582 B.n376 B.n375 163.367
R583 B.n375 B.n374 163.367
R584 B.n374 B.n39 163.367
R585 B.n370 B.n39 163.367
R586 B.n370 B.n369 163.367
R587 B.n369 B.n368 163.367
R588 B.n368 B.n41 163.367
R589 B.n364 B.n41 163.367
R590 B.n364 B.n363 163.367
R591 B.n363 B.n362 163.367
R592 B.n362 B.n43 163.367
R593 B.n358 B.n43 163.367
R594 B.n358 B.n357 163.367
R595 B.n357 B.n356 163.367
R596 B.n356 B.n45 163.367
R597 B.n352 B.n45 163.367
R598 B.n352 B.n351 163.367
R599 B.n351 B.n350 163.367
R600 B.n424 B.n423 163.367
R601 B.n424 B.n17 163.367
R602 B.n428 B.n17 163.367
R603 B.n429 B.n428 163.367
R604 B.n430 B.n429 163.367
R605 B.n430 B.n15 163.367
R606 B.n434 B.n15 163.367
R607 B.n435 B.n434 163.367
R608 B.n436 B.n435 163.367
R609 B.n436 B.n13 163.367
R610 B.n440 B.n13 163.367
R611 B.n441 B.n440 163.367
R612 B.n442 B.n441 163.367
R613 B.n442 B.n11 163.367
R614 B.n446 B.n11 163.367
R615 B.n447 B.n446 163.367
R616 B.n448 B.n447 163.367
R617 B.n448 B.n9 163.367
R618 B.n452 B.n9 163.367
R619 B.n453 B.n452 163.367
R620 B.n454 B.n453 163.367
R621 B.n454 B.n7 163.367
R622 B.n458 B.n7 163.367
R623 B.n459 B.n458 163.367
R624 B.n460 B.n459 163.367
R625 B.n460 B.n5 163.367
R626 B.n464 B.n5 163.367
R627 B.n465 B.n464 163.367
R628 B.n466 B.n465 163.367
R629 B.n466 B.n3 163.367
R630 B.n470 B.n3 163.367
R631 B.n471 B.n470 163.367
R632 B.n124 B.n2 163.367
R633 B.n125 B.n124 163.367
R634 B.n126 B.n125 163.367
R635 B.n126 B.n121 163.367
R636 B.n130 B.n121 163.367
R637 B.n131 B.n130 163.367
R638 B.n132 B.n131 163.367
R639 B.n132 B.n119 163.367
R640 B.n136 B.n119 163.367
R641 B.n137 B.n136 163.367
R642 B.n138 B.n137 163.367
R643 B.n138 B.n117 163.367
R644 B.n142 B.n117 163.367
R645 B.n143 B.n142 163.367
R646 B.n144 B.n143 163.367
R647 B.n144 B.n115 163.367
R648 B.n148 B.n115 163.367
R649 B.n149 B.n148 163.367
R650 B.n150 B.n149 163.367
R651 B.n150 B.n113 163.367
R652 B.n154 B.n113 163.367
R653 B.n155 B.n154 163.367
R654 B.n156 B.n155 163.367
R655 B.n156 B.n111 163.367
R656 B.n160 B.n111 163.367
R657 B.n161 B.n160 163.367
R658 B.n162 B.n161 163.367
R659 B.n162 B.n109 163.367
R660 B.n166 B.n109 163.367
R661 B.n167 B.n166 163.367
R662 B.n168 B.n167 163.367
R663 B.n168 B.n107 163.367
R664 B.n214 B.t7 158.641
R665 B.n36 B.t5 158.641
R666 B.n96 B.t1 158.637
R667 B.n28 B.t11 158.637
R668 B.n215 B.t8 124.894
R669 B.n37 B.t4 124.894
R670 B.n97 B.t2 124.891
R671 B.n29 B.t10 124.891
R672 B.n200 B.n97 59.5399
R673 B.n216 B.n215 59.5399
R674 B.n378 B.n37 59.5399
R675 B.n30 B.n29 59.5399
R676 B.n247 B.n246 35.4346
R677 B.n421 B.n18 35.4346
R678 B.n349 B.n348 35.4346
R679 B.n171 B.n170 35.4346
R680 B.n97 B.n96 33.746
R681 B.n215 B.n214 33.746
R682 B.n37 B.n36 33.746
R683 B.n29 B.n28 33.746
R684 B B.n473 18.0485
R685 B.n425 B.n18 10.6151
R686 B.n426 B.n425 10.6151
R687 B.n427 B.n426 10.6151
R688 B.n427 B.n16 10.6151
R689 B.n431 B.n16 10.6151
R690 B.n432 B.n431 10.6151
R691 B.n433 B.n432 10.6151
R692 B.n433 B.n14 10.6151
R693 B.n437 B.n14 10.6151
R694 B.n438 B.n437 10.6151
R695 B.n439 B.n438 10.6151
R696 B.n439 B.n12 10.6151
R697 B.n443 B.n12 10.6151
R698 B.n444 B.n443 10.6151
R699 B.n445 B.n444 10.6151
R700 B.n445 B.n10 10.6151
R701 B.n449 B.n10 10.6151
R702 B.n450 B.n449 10.6151
R703 B.n451 B.n450 10.6151
R704 B.n451 B.n8 10.6151
R705 B.n455 B.n8 10.6151
R706 B.n456 B.n455 10.6151
R707 B.n457 B.n456 10.6151
R708 B.n457 B.n6 10.6151
R709 B.n461 B.n6 10.6151
R710 B.n462 B.n461 10.6151
R711 B.n463 B.n462 10.6151
R712 B.n463 B.n4 10.6151
R713 B.n467 B.n4 10.6151
R714 B.n468 B.n467 10.6151
R715 B.n469 B.n468 10.6151
R716 B.n469 B.n0 10.6151
R717 B.n421 B.n420 10.6151
R718 B.n420 B.n419 10.6151
R719 B.n419 B.n20 10.6151
R720 B.n415 B.n20 10.6151
R721 B.n415 B.n414 10.6151
R722 B.n414 B.n413 10.6151
R723 B.n413 B.n22 10.6151
R724 B.n409 B.n22 10.6151
R725 B.n409 B.n408 10.6151
R726 B.n408 B.n407 10.6151
R727 B.n407 B.n24 10.6151
R728 B.n403 B.n24 10.6151
R729 B.n403 B.n402 10.6151
R730 B.n402 B.n401 10.6151
R731 B.n401 B.n26 10.6151
R732 B.n397 B.n26 10.6151
R733 B.n397 B.n396 10.6151
R734 B.n396 B.n395 10.6151
R735 B.n392 B.n391 10.6151
R736 B.n391 B.n390 10.6151
R737 B.n390 B.n32 10.6151
R738 B.n386 B.n32 10.6151
R739 B.n386 B.n385 10.6151
R740 B.n385 B.n384 10.6151
R741 B.n384 B.n34 10.6151
R742 B.n380 B.n34 10.6151
R743 B.n380 B.n379 10.6151
R744 B.n377 B.n38 10.6151
R745 B.n373 B.n38 10.6151
R746 B.n373 B.n372 10.6151
R747 B.n372 B.n371 10.6151
R748 B.n371 B.n40 10.6151
R749 B.n367 B.n40 10.6151
R750 B.n367 B.n366 10.6151
R751 B.n366 B.n365 10.6151
R752 B.n365 B.n42 10.6151
R753 B.n361 B.n42 10.6151
R754 B.n361 B.n360 10.6151
R755 B.n360 B.n359 10.6151
R756 B.n359 B.n44 10.6151
R757 B.n355 B.n44 10.6151
R758 B.n355 B.n354 10.6151
R759 B.n354 B.n353 10.6151
R760 B.n353 B.n46 10.6151
R761 B.n349 B.n46 10.6151
R762 B.n348 B.n347 10.6151
R763 B.n347 B.n48 10.6151
R764 B.n343 B.n48 10.6151
R765 B.n343 B.n342 10.6151
R766 B.n342 B.n341 10.6151
R767 B.n341 B.n50 10.6151
R768 B.n337 B.n50 10.6151
R769 B.n337 B.n336 10.6151
R770 B.n336 B.n335 10.6151
R771 B.n335 B.n52 10.6151
R772 B.n331 B.n52 10.6151
R773 B.n331 B.n330 10.6151
R774 B.n330 B.n329 10.6151
R775 B.n329 B.n54 10.6151
R776 B.n325 B.n54 10.6151
R777 B.n325 B.n324 10.6151
R778 B.n324 B.n323 10.6151
R779 B.n323 B.n56 10.6151
R780 B.n319 B.n56 10.6151
R781 B.n319 B.n318 10.6151
R782 B.n318 B.n317 10.6151
R783 B.n317 B.n58 10.6151
R784 B.n313 B.n58 10.6151
R785 B.n313 B.n312 10.6151
R786 B.n312 B.n311 10.6151
R787 B.n311 B.n60 10.6151
R788 B.n307 B.n60 10.6151
R789 B.n307 B.n306 10.6151
R790 B.n306 B.n305 10.6151
R791 B.n305 B.n62 10.6151
R792 B.n301 B.n62 10.6151
R793 B.n301 B.n300 10.6151
R794 B.n300 B.n299 10.6151
R795 B.n299 B.n64 10.6151
R796 B.n295 B.n64 10.6151
R797 B.n295 B.n294 10.6151
R798 B.n294 B.n293 10.6151
R799 B.n293 B.n66 10.6151
R800 B.n289 B.n66 10.6151
R801 B.n289 B.n288 10.6151
R802 B.n288 B.n287 10.6151
R803 B.n287 B.n68 10.6151
R804 B.n283 B.n68 10.6151
R805 B.n283 B.n282 10.6151
R806 B.n282 B.n281 10.6151
R807 B.n281 B.n70 10.6151
R808 B.n277 B.n70 10.6151
R809 B.n277 B.n276 10.6151
R810 B.n276 B.n275 10.6151
R811 B.n275 B.n72 10.6151
R812 B.n271 B.n72 10.6151
R813 B.n271 B.n270 10.6151
R814 B.n270 B.n269 10.6151
R815 B.n269 B.n74 10.6151
R816 B.n265 B.n74 10.6151
R817 B.n265 B.n264 10.6151
R818 B.n264 B.n263 10.6151
R819 B.n263 B.n76 10.6151
R820 B.n259 B.n76 10.6151
R821 B.n259 B.n258 10.6151
R822 B.n258 B.n257 10.6151
R823 B.n257 B.n78 10.6151
R824 B.n253 B.n78 10.6151
R825 B.n253 B.n252 10.6151
R826 B.n252 B.n251 10.6151
R827 B.n251 B.n80 10.6151
R828 B.n247 B.n80 10.6151
R829 B.n123 B.n1 10.6151
R830 B.n123 B.n122 10.6151
R831 B.n127 B.n122 10.6151
R832 B.n128 B.n127 10.6151
R833 B.n129 B.n128 10.6151
R834 B.n129 B.n120 10.6151
R835 B.n133 B.n120 10.6151
R836 B.n134 B.n133 10.6151
R837 B.n135 B.n134 10.6151
R838 B.n135 B.n118 10.6151
R839 B.n139 B.n118 10.6151
R840 B.n140 B.n139 10.6151
R841 B.n141 B.n140 10.6151
R842 B.n141 B.n116 10.6151
R843 B.n145 B.n116 10.6151
R844 B.n146 B.n145 10.6151
R845 B.n147 B.n146 10.6151
R846 B.n147 B.n114 10.6151
R847 B.n151 B.n114 10.6151
R848 B.n152 B.n151 10.6151
R849 B.n153 B.n152 10.6151
R850 B.n153 B.n112 10.6151
R851 B.n157 B.n112 10.6151
R852 B.n158 B.n157 10.6151
R853 B.n159 B.n158 10.6151
R854 B.n159 B.n110 10.6151
R855 B.n163 B.n110 10.6151
R856 B.n164 B.n163 10.6151
R857 B.n165 B.n164 10.6151
R858 B.n165 B.n108 10.6151
R859 B.n169 B.n108 10.6151
R860 B.n170 B.n169 10.6151
R861 B.n171 B.n106 10.6151
R862 B.n175 B.n106 10.6151
R863 B.n176 B.n175 10.6151
R864 B.n177 B.n176 10.6151
R865 B.n177 B.n104 10.6151
R866 B.n181 B.n104 10.6151
R867 B.n182 B.n181 10.6151
R868 B.n183 B.n182 10.6151
R869 B.n183 B.n102 10.6151
R870 B.n187 B.n102 10.6151
R871 B.n188 B.n187 10.6151
R872 B.n189 B.n188 10.6151
R873 B.n189 B.n100 10.6151
R874 B.n193 B.n100 10.6151
R875 B.n194 B.n193 10.6151
R876 B.n195 B.n194 10.6151
R877 B.n195 B.n98 10.6151
R878 B.n199 B.n98 10.6151
R879 B.n202 B.n201 10.6151
R880 B.n202 B.n94 10.6151
R881 B.n206 B.n94 10.6151
R882 B.n207 B.n206 10.6151
R883 B.n208 B.n207 10.6151
R884 B.n208 B.n92 10.6151
R885 B.n212 B.n92 10.6151
R886 B.n213 B.n212 10.6151
R887 B.n217 B.n213 10.6151
R888 B.n221 B.n90 10.6151
R889 B.n222 B.n221 10.6151
R890 B.n223 B.n222 10.6151
R891 B.n223 B.n88 10.6151
R892 B.n227 B.n88 10.6151
R893 B.n228 B.n227 10.6151
R894 B.n229 B.n228 10.6151
R895 B.n229 B.n86 10.6151
R896 B.n233 B.n86 10.6151
R897 B.n234 B.n233 10.6151
R898 B.n235 B.n234 10.6151
R899 B.n235 B.n84 10.6151
R900 B.n239 B.n84 10.6151
R901 B.n240 B.n239 10.6151
R902 B.n241 B.n240 10.6151
R903 B.n241 B.n82 10.6151
R904 B.n245 B.n82 10.6151
R905 B.n246 B.n245 10.6151
R906 B.n395 B.n30 9.36635
R907 B.n378 B.n377 9.36635
R908 B.n200 B.n199 9.36635
R909 B.n216 B.n90 9.36635
R910 B.n473 B.n0 8.11757
R911 B.n473 B.n1 8.11757
R912 B.n392 B.n30 1.24928
R913 B.n379 B.n378 1.24928
R914 B.n201 B.n200 1.24928
R915 B.n217 B.n216 1.24928
C0 B VDD2 1.14109f
C1 VN VDD2 2.98503f
C2 VTAIL VP 3.44441f
C3 VTAIL w_n2710_n1850# 2.33598f
C4 B VP 1.45134f
C5 B w_n2710_n1850# 6.17044f
C6 VDD1 VDD2 1.18364f
C7 VN VP 4.81123f
C8 VN w_n2710_n1850# 5.05338f
C9 VDD1 VP 3.22765f
C10 VDD1 w_n2710_n1850# 1.35752f
C11 VTAIL B 2.06689f
C12 VTAIL VN 3.43031f
C13 VN B 0.873928f
C14 VDD1 VTAIL 4.94557f
C15 VDD2 VP 0.397596f
C16 w_n2710_n1850# VDD2 1.42194f
C17 VDD1 B 1.08234f
C18 VDD1 VN 0.153715f
C19 w_n2710_n1850# VP 5.40134f
C20 VTAIL VDD2 4.99201f
C21 VDD2 VSUBS 1.175641f
C22 VDD1 VSUBS 1.605918f
C23 VTAIL VSUBS 0.533388f
C24 VN VSUBS 4.8892f
C25 VP VSUBS 1.89803f
C26 B VSUBS 2.875876f
C27 w_n2710_n1850# VSUBS 62.991196f
C28 B.n0 VSUBS 0.008225f
C29 B.n1 VSUBS 0.008225f
C30 B.n2 VSUBS 0.012164f
C31 B.n3 VSUBS 0.009322f
C32 B.n4 VSUBS 0.009322f
C33 B.n5 VSUBS 0.009322f
C34 B.n6 VSUBS 0.009322f
C35 B.n7 VSUBS 0.009322f
C36 B.n8 VSUBS 0.009322f
C37 B.n9 VSUBS 0.009322f
C38 B.n10 VSUBS 0.009322f
C39 B.n11 VSUBS 0.009322f
C40 B.n12 VSUBS 0.009322f
C41 B.n13 VSUBS 0.009322f
C42 B.n14 VSUBS 0.009322f
C43 B.n15 VSUBS 0.009322f
C44 B.n16 VSUBS 0.009322f
C45 B.n17 VSUBS 0.009322f
C46 B.n18 VSUBS 0.022448f
C47 B.n19 VSUBS 0.009322f
C48 B.n20 VSUBS 0.009322f
C49 B.n21 VSUBS 0.009322f
C50 B.n22 VSUBS 0.009322f
C51 B.n23 VSUBS 0.009322f
C52 B.n24 VSUBS 0.009322f
C53 B.n25 VSUBS 0.009322f
C54 B.n26 VSUBS 0.009322f
C55 B.n27 VSUBS 0.009322f
C56 B.t10 VSUBS 0.158124f
C57 B.t11 VSUBS 0.173644f
C58 B.t9 VSUBS 0.385212f
C59 B.n28 VSUBS 0.114508f
C60 B.n29 VSUBS 0.086253f
C61 B.n30 VSUBS 0.021597f
C62 B.n31 VSUBS 0.009322f
C63 B.n32 VSUBS 0.009322f
C64 B.n33 VSUBS 0.009322f
C65 B.n34 VSUBS 0.009322f
C66 B.n35 VSUBS 0.009322f
C67 B.t4 VSUBS 0.158124f
C68 B.t5 VSUBS 0.173643f
C69 B.t3 VSUBS 0.385212f
C70 B.n36 VSUBS 0.114509f
C71 B.n37 VSUBS 0.086253f
C72 B.n38 VSUBS 0.009322f
C73 B.n39 VSUBS 0.009322f
C74 B.n40 VSUBS 0.009322f
C75 B.n41 VSUBS 0.009322f
C76 B.n42 VSUBS 0.009322f
C77 B.n43 VSUBS 0.009322f
C78 B.n44 VSUBS 0.009322f
C79 B.n45 VSUBS 0.009322f
C80 B.n46 VSUBS 0.009322f
C81 B.n47 VSUBS 0.022448f
C82 B.n48 VSUBS 0.009322f
C83 B.n49 VSUBS 0.009322f
C84 B.n50 VSUBS 0.009322f
C85 B.n51 VSUBS 0.009322f
C86 B.n52 VSUBS 0.009322f
C87 B.n53 VSUBS 0.009322f
C88 B.n54 VSUBS 0.009322f
C89 B.n55 VSUBS 0.009322f
C90 B.n56 VSUBS 0.009322f
C91 B.n57 VSUBS 0.009322f
C92 B.n58 VSUBS 0.009322f
C93 B.n59 VSUBS 0.009322f
C94 B.n60 VSUBS 0.009322f
C95 B.n61 VSUBS 0.009322f
C96 B.n62 VSUBS 0.009322f
C97 B.n63 VSUBS 0.009322f
C98 B.n64 VSUBS 0.009322f
C99 B.n65 VSUBS 0.009322f
C100 B.n66 VSUBS 0.009322f
C101 B.n67 VSUBS 0.009322f
C102 B.n68 VSUBS 0.009322f
C103 B.n69 VSUBS 0.009322f
C104 B.n70 VSUBS 0.009322f
C105 B.n71 VSUBS 0.009322f
C106 B.n72 VSUBS 0.009322f
C107 B.n73 VSUBS 0.009322f
C108 B.n74 VSUBS 0.009322f
C109 B.n75 VSUBS 0.009322f
C110 B.n76 VSUBS 0.009322f
C111 B.n77 VSUBS 0.009322f
C112 B.n78 VSUBS 0.009322f
C113 B.n79 VSUBS 0.009322f
C114 B.n80 VSUBS 0.009322f
C115 B.n81 VSUBS 0.023612f
C116 B.n82 VSUBS 0.009322f
C117 B.n83 VSUBS 0.009322f
C118 B.n84 VSUBS 0.009322f
C119 B.n85 VSUBS 0.009322f
C120 B.n86 VSUBS 0.009322f
C121 B.n87 VSUBS 0.009322f
C122 B.n88 VSUBS 0.009322f
C123 B.n89 VSUBS 0.009322f
C124 B.n90 VSUBS 0.008773f
C125 B.n91 VSUBS 0.009322f
C126 B.n92 VSUBS 0.009322f
C127 B.n93 VSUBS 0.009322f
C128 B.n94 VSUBS 0.009322f
C129 B.n95 VSUBS 0.009322f
C130 B.t2 VSUBS 0.158124f
C131 B.t1 VSUBS 0.173644f
C132 B.t0 VSUBS 0.385212f
C133 B.n96 VSUBS 0.114508f
C134 B.n97 VSUBS 0.086253f
C135 B.n98 VSUBS 0.009322f
C136 B.n99 VSUBS 0.009322f
C137 B.n100 VSUBS 0.009322f
C138 B.n101 VSUBS 0.009322f
C139 B.n102 VSUBS 0.009322f
C140 B.n103 VSUBS 0.009322f
C141 B.n104 VSUBS 0.009322f
C142 B.n105 VSUBS 0.009322f
C143 B.n106 VSUBS 0.009322f
C144 B.n107 VSUBS 0.022448f
C145 B.n108 VSUBS 0.009322f
C146 B.n109 VSUBS 0.009322f
C147 B.n110 VSUBS 0.009322f
C148 B.n111 VSUBS 0.009322f
C149 B.n112 VSUBS 0.009322f
C150 B.n113 VSUBS 0.009322f
C151 B.n114 VSUBS 0.009322f
C152 B.n115 VSUBS 0.009322f
C153 B.n116 VSUBS 0.009322f
C154 B.n117 VSUBS 0.009322f
C155 B.n118 VSUBS 0.009322f
C156 B.n119 VSUBS 0.009322f
C157 B.n120 VSUBS 0.009322f
C158 B.n121 VSUBS 0.009322f
C159 B.n122 VSUBS 0.009322f
C160 B.n123 VSUBS 0.009322f
C161 B.n124 VSUBS 0.009322f
C162 B.n125 VSUBS 0.009322f
C163 B.n126 VSUBS 0.009322f
C164 B.n127 VSUBS 0.009322f
C165 B.n128 VSUBS 0.009322f
C166 B.n129 VSUBS 0.009322f
C167 B.n130 VSUBS 0.009322f
C168 B.n131 VSUBS 0.009322f
C169 B.n132 VSUBS 0.009322f
C170 B.n133 VSUBS 0.009322f
C171 B.n134 VSUBS 0.009322f
C172 B.n135 VSUBS 0.009322f
C173 B.n136 VSUBS 0.009322f
C174 B.n137 VSUBS 0.009322f
C175 B.n138 VSUBS 0.009322f
C176 B.n139 VSUBS 0.009322f
C177 B.n140 VSUBS 0.009322f
C178 B.n141 VSUBS 0.009322f
C179 B.n142 VSUBS 0.009322f
C180 B.n143 VSUBS 0.009322f
C181 B.n144 VSUBS 0.009322f
C182 B.n145 VSUBS 0.009322f
C183 B.n146 VSUBS 0.009322f
C184 B.n147 VSUBS 0.009322f
C185 B.n148 VSUBS 0.009322f
C186 B.n149 VSUBS 0.009322f
C187 B.n150 VSUBS 0.009322f
C188 B.n151 VSUBS 0.009322f
C189 B.n152 VSUBS 0.009322f
C190 B.n153 VSUBS 0.009322f
C191 B.n154 VSUBS 0.009322f
C192 B.n155 VSUBS 0.009322f
C193 B.n156 VSUBS 0.009322f
C194 B.n157 VSUBS 0.009322f
C195 B.n158 VSUBS 0.009322f
C196 B.n159 VSUBS 0.009322f
C197 B.n160 VSUBS 0.009322f
C198 B.n161 VSUBS 0.009322f
C199 B.n162 VSUBS 0.009322f
C200 B.n163 VSUBS 0.009322f
C201 B.n164 VSUBS 0.009322f
C202 B.n165 VSUBS 0.009322f
C203 B.n166 VSUBS 0.009322f
C204 B.n167 VSUBS 0.009322f
C205 B.n168 VSUBS 0.009322f
C206 B.n169 VSUBS 0.009322f
C207 B.n170 VSUBS 0.022448f
C208 B.n171 VSUBS 0.023612f
C209 B.n172 VSUBS 0.023612f
C210 B.n173 VSUBS 0.009322f
C211 B.n174 VSUBS 0.009322f
C212 B.n175 VSUBS 0.009322f
C213 B.n176 VSUBS 0.009322f
C214 B.n177 VSUBS 0.009322f
C215 B.n178 VSUBS 0.009322f
C216 B.n179 VSUBS 0.009322f
C217 B.n180 VSUBS 0.009322f
C218 B.n181 VSUBS 0.009322f
C219 B.n182 VSUBS 0.009322f
C220 B.n183 VSUBS 0.009322f
C221 B.n184 VSUBS 0.009322f
C222 B.n185 VSUBS 0.009322f
C223 B.n186 VSUBS 0.009322f
C224 B.n187 VSUBS 0.009322f
C225 B.n188 VSUBS 0.009322f
C226 B.n189 VSUBS 0.009322f
C227 B.n190 VSUBS 0.009322f
C228 B.n191 VSUBS 0.009322f
C229 B.n192 VSUBS 0.009322f
C230 B.n193 VSUBS 0.009322f
C231 B.n194 VSUBS 0.009322f
C232 B.n195 VSUBS 0.009322f
C233 B.n196 VSUBS 0.009322f
C234 B.n197 VSUBS 0.009322f
C235 B.n198 VSUBS 0.009322f
C236 B.n199 VSUBS 0.008773f
C237 B.n200 VSUBS 0.021597f
C238 B.n201 VSUBS 0.005209f
C239 B.n202 VSUBS 0.009322f
C240 B.n203 VSUBS 0.009322f
C241 B.n204 VSUBS 0.009322f
C242 B.n205 VSUBS 0.009322f
C243 B.n206 VSUBS 0.009322f
C244 B.n207 VSUBS 0.009322f
C245 B.n208 VSUBS 0.009322f
C246 B.n209 VSUBS 0.009322f
C247 B.n210 VSUBS 0.009322f
C248 B.n211 VSUBS 0.009322f
C249 B.n212 VSUBS 0.009322f
C250 B.n213 VSUBS 0.009322f
C251 B.t8 VSUBS 0.158124f
C252 B.t7 VSUBS 0.173643f
C253 B.t6 VSUBS 0.385212f
C254 B.n214 VSUBS 0.114509f
C255 B.n215 VSUBS 0.086253f
C256 B.n216 VSUBS 0.021597f
C257 B.n217 VSUBS 0.005209f
C258 B.n218 VSUBS 0.009322f
C259 B.n219 VSUBS 0.009322f
C260 B.n220 VSUBS 0.009322f
C261 B.n221 VSUBS 0.009322f
C262 B.n222 VSUBS 0.009322f
C263 B.n223 VSUBS 0.009322f
C264 B.n224 VSUBS 0.009322f
C265 B.n225 VSUBS 0.009322f
C266 B.n226 VSUBS 0.009322f
C267 B.n227 VSUBS 0.009322f
C268 B.n228 VSUBS 0.009322f
C269 B.n229 VSUBS 0.009322f
C270 B.n230 VSUBS 0.009322f
C271 B.n231 VSUBS 0.009322f
C272 B.n232 VSUBS 0.009322f
C273 B.n233 VSUBS 0.009322f
C274 B.n234 VSUBS 0.009322f
C275 B.n235 VSUBS 0.009322f
C276 B.n236 VSUBS 0.009322f
C277 B.n237 VSUBS 0.009322f
C278 B.n238 VSUBS 0.009322f
C279 B.n239 VSUBS 0.009322f
C280 B.n240 VSUBS 0.009322f
C281 B.n241 VSUBS 0.009322f
C282 B.n242 VSUBS 0.009322f
C283 B.n243 VSUBS 0.009322f
C284 B.n244 VSUBS 0.009322f
C285 B.n245 VSUBS 0.009322f
C286 B.n246 VSUBS 0.022597f
C287 B.n247 VSUBS 0.023463f
C288 B.n248 VSUBS 0.022448f
C289 B.n249 VSUBS 0.009322f
C290 B.n250 VSUBS 0.009322f
C291 B.n251 VSUBS 0.009322f
C292 B.n252 VSUBS 0.009322f
C293 B.n253 VSUBS 0.009322f
C294 B.n254 VSUBS 0.009322f
C295 B.n255 VSUBS 0.009322f
C296 B.n256 VSUBS 0.009322f
C297 B.n257 VSUBS 0.009322f
C298 B.n258 VSUBS 0.009322f
C299 B.n259 VSUBS 0.009322f
C300 B.n260 VSUBS 0.009322f
C301 B.n261 VSUBS 0.009322f
C302 B.n262 VSUBS 0.009322f
C303 B.n263 VSUBS 0.009322f
C304 B.n264 VSUBS 0.009322f
C305 B.n265 VSUBS 0.009322f
C306 B.n266 VSUBS 0.009322f
C307 B.n267 VSUBS 0.009322f
C308 B.n268 VSUBS 0.009322f
C309 B.n269 VSUBS 0.009322f
C310 B.n270 VSUBS 0.009322f
C311 B.n271 VSUBS 0.009322f
C312 B.n272 VSUBS 0.009322f
C313 B.n273 VSUBS 0.009322f
C314 B.n274 VSUBS 0.009322f
C315 B.n275 VSUBS 0.009322f
C316 B.n276 VSUBS 0.009322f
C317 B.n277 VSUBS 0.009322f
C318 B.n278 VSUBS 0.009322f
C319 B.n279 VSUBS 0.009322f
C320 B.n280 VSUBS 0.009322f
C321 B.n281 VSUBS 0.009322f
C322 B.n282 VSUBS 0.009322f
C323 B.n283 VSUBS 0.009322f
C324 B.n284 VSUBS 0.009322f
C325 B.n285 VSUBS 0.009322f
C326 B.n286 VSUBS 0.009322f
C327 B.n287 VSUBS 0.009322f
C328 B.n288 VSUBS 0.009322f
C329 B.n289 VSUBS 0.009322f
C330 B.n290 VSUBS 0.009322f
C331 B.n291 VSUBS 0.009322f
C332 B.n292 VSUBS 0.009322f
C333 B.n293 VSUBS 0.009322f
C334 B.n294 VSUBS 0.009322f
C335 B.n295 VSUBS 0.009322f
C336 B.n296 VSUBS 0.009322f
C337 B.n297 VSUBS 0.009322f
C338 B.n298 VSUBS 0.009322f
C339 B.n299 VSUBS 0.009322f
C340 B.n300 VSUBS 0.009322f
C341 B.n301 VSUBS 0.009322f
C342 B.n302 VSUBS 0.009322f
C343 B.n303 VSUBS 0.009322f
C344 B.n304 VSUBS 0.009322f
C345 B.n305 VSUBS 0.009322f
C346 B.n306 VSUBS 0.009322f
C347 B.n307 VSUBS 0.009322f
C348 B.n308 VSUBS 0.009322f
C349 B.n309 VSUBS 0.009322f
C350 B.n310 VSUBS 0.009322f
C351 B.n311 VSUBS 0.009322f
C352 B.n312 VSUBS 0.009322f
C353 B.n313 VSUBS 0.009322f
C354 B.n314 VSUBS 0.009322f
C355 B.n315 VSUBS 0.009322f
C356 B.n316 VSUBS 0.009322f
C357 B.n317 VSUBS 0.009322f
C358 B.n318 VSUBS 0.009322f
C359 B.n319 VSUBS 0.009322f
C360 B.n320 VSUBS 0.009322f
C361 B.n321 VSUBS 0.009322f
C362 B.n322 VSUBS 0.009322f
C363 B.n323 VSUBS 0.009322f
C364 B.n324 VSUBS 0.009322f
C365 B.n325 VSUBS 0.009322f
C366 B.n326 VSUBS 0.009322f
C367 B.n327 VSUBS 0.009322f
C368 B.n328 VSUBS 0.009322f
C369 B.n329 VSUBS 0.009322f
C370 B.n330 VSUBS 0.009322f
C371 B.n331 VSUBS 0.009322f
C372 B.n332 VSUBS 0.009322f
C373 B.n333 VSUBS 0.009322f
C374 B.n334 VSUBS 0.009322f
C375 B.n335 VSUBS 0.009322f
C376 B.n336 VSUBS 0.009322f
C377 B.n337 VSUBS 0.009322f
C378 B.n338 VSUBS 0.009322f
C379 B.n339 VSUBS 0.009322f
C380 B.n340 VSUBS 0.009322f
C381 B.n341 VSUBS 0.009322f
C382 B.n342 VSUBS 0.009322f
C383 B.n343 VSUBS 0.009322f
C384 B.n344 VSUBS 0.009322f
C385 B.n345 VSUBS 0.009322f
C386 B.n346 VSUBS 0.009322f
C387 B.n347 VSUBS 0.009322f
C388 B.n348 VSUBS 0.022448f
C389 B.n349 VSUBS 0.023612f
C390 B.n350 VSUBS 0.023612f
C391 B.n351 VSUBS 0.009322f
C392 B.n352 VSUBS 0.009322f
C393 B.n353 VSUBS 0.009322f
C394 B.n354 VSUBS 0.009322f
C395 B.n355 VSUBS 0.009322f
C396 B.n356 VSUBS 0.009322f
C397 B.n357 VSUBS 0.009322f
C398 B.n358 VSUBS 0.009322f
C399 B.n359 VSUBS 0.009322f
C400 B.n360 VSUBS 0.009322f
C401 B.n361 VSUBS 0.009322f
C402 B.n362 VSUBS 0.009322f
C403 B.n363 VSUBS 0.009322f
C404 B.n364 VSUBS 0.009322f
C405 B.n365 VSUBS 0.009322f
C406 B.n366 VSUBS 0.009322f
C407 B.n367 VSUBS 0.009322f
C408 B.n368 VSUBS 0.009322f
C409 B.n369 VSUBS 0.009322f
C410 B.n370 VSUBS 0.009322f
C411 B.n371 VSUBS 0.009322f
C412 B.n372 VSUBS 0.009322f
C413 B.n373 VSUBS 0.009322f
C414 B.n374 VSUBS 0.009322f
C415 B.n375 VSUBS 0.009322f
C416 B.n376 VSUBS 0.009322f
C417 B.n377 VSUBS 0.008773f
C418 B.n378 VSUBS 0.021597f
C419 B.n379 VSUBS 0.005209f
C420 B.n380 VSUBS 0.009322f
C421 B.n381 VSUBS 0.009322f
C422 B.n382 VSUBS 0.009322f
C423 B.n383 VSUBS 0.009322f
C424 B.n384 VSUBS 0.009322f
C425 B.n385 VSUBS 0.009322f
C426 B.n386 VSUBS 0.009322f
C427 B.n387 VSUBS 0.009322f
C428 B.n388 VSUBS 0.009322f
C429 B.n389 VSUBS 0.009322f
C430 B.n390 VSUBS 0.009322f
C431 B.n391 VSUBS 0.009322f
C432 B.n392 VSUBS 0.005209f
C433 B.n393 VSUBS 0.009322f
C434 B.n394 VSUBS 0.009322f
C435 B.n395 VSUBS 0.008773f
C436 B.n396 VSUBS 0.009322f
C437 B.n397 VSUBS 0.009322f
C438 B.n398 VSUBS 0.009322f
C439 B.n399 VSUBS 0.009322f
C440 B.n400 VSUBS 0.009322f
C441 B.n401 VSUBS 0.009322f
C442 B.n402 VSUBS 0.009322f
C443 B.n403 VSUBS 0.009322f
C444 B.n404 VSUBS 0.009322f
C445 B.n405 VSUBS 0.009322f
C446 B.n406 VSUBS 0.009322f
C447 B.n407 VSUBS 0.009322f
C448 B.n408 VSUBS 0.009322f
C449 B.n409 VSUBS 0.009322f
C450 B.n410 VSUBS 0.009322f
C451 B.n411 VSUBS 0.009322f
C452 B.n412 VSUBS 0.009322f
C453 B.n413 VSUBS 0.009322f
C454 B.n414 VSUBS 0.009322f
C455 B.n415 VSUBS 0.009322f
C456 B.n416 VSUBS 0.009322f
C457 B.n417 VSUBS 0.009322f
C458 B.n418 VSUBS 0.009322f
C459 B.n419 VSUBS 0.009322f
C460 B.n420 VSUBS 0.009322f
C461 B.n421 VSUBS 0.023612f
C462 B.n422 VSUBS 0.023612f
C463 B.n423 VSUBS 0.022448f
C464 B.n424 VSUBS 0.009322f
C465 B.n425 VSUBS 0.009322f
C466 B.n426 VSUBS 0.009322f
C467 B.n427 VSUBS 0.009322f
C468 B.n428 VSUBS 0.009322f
C469 B.n429 VSUBS 0.009322f
C470 B.n430 VSUBS 0.009322f
C471 B.n431 VSUBS 0.009322f
C472 B.n432 VSUBS 0.009322f
C473 B.n433 VSUBS 0.009322f
C474 B.n434 VSUBS 0.009322f
C475 B.n435 VSUBS 0.009322f
C476 B.n436 VSUBS 0.009322f
C477 B.n437 VSUBS 0.009322f
C478 B.n438 VSUBS 0.009322f
C479 B.n439 VSUBS 0.009322f
C480 B.n440 VSUBS 0.009322f
C481 B.n441 VSUBS 0.009322f
C482 B.n442 VSUBS 0.009322f
C483 B.n443 VSUBS 0.009322f
C484 B.n444 VSUBS 0.009322f
C485 B.n445 VSUBS 0.009322f
C486 B.n446 VSUBS 0.009322f
C487 B.n447 VSUBS 0.009322f
C488 B.n448 VSUBS 0.009322f
C489 B.n449 VSUBS 0.009322f
C490 B.n450 VSUBS 0.009322f
C491 B.n451 VSUBS 0.009322f
C492 B.n452 VSUBS 0.009322f
C493 B.n453 VSUBS 0.009322f
C494 B.n454 VSUBS 0.009322f
C495 B.n455 VSUBS 0.009322f
C496 B.n456 VSUBS 0.009322f
C497 B.n457 VSUBS 0.009322f
C498 B.n458 VSUBS 0.009322f
C499 B.n459 VSUBS 0.009322f
C500 B.n460 VSUBS 0.009322f
C501 B.n461 VSUBS 0.009322f
C502 B.n462 VSUBS 0.009322f
C503 B.n463 VSUBS 0.009322f
C504 B.n464 VSUBS 0.009322f
C505 B.n465 VSUBS 0.009322f
C506 B.n466 VSUBS 0.009322f
C507 B.n467 VSUBS 0.009322f
C508 B.n468 VSUBS 0.009322f
C509 B.n469 VSUBS 0.009322f
C510 B.n470 VSUBS 0.009322f
C511 B.n471 VSUBS 0.012164f
C512 B.n472 VSUBS 0.012958f
C513 B.n473 VSUBS 0.025768f
C514 VDD1.t6 VSUBS 0.086828f
C515 VDD1.t1 VSUBS 0.086828f
C516 VDD1.n0 VSUBS 0.529191f
C517 VDD1.t7 VSUBS 0.086828f
C518 VDD1.t5 VSUBS 0.086828f
C519 VDD1.n1 VSUBS 0.528581f
C520 VDD1.t2 VSUBS 0.086828f
C521 VDD1.t3 VSUBS 0.086828f
C522 VDD1.n2 VSUBS 0.528581f
C523 VDD1.n3 VSUBS 2.49509f
C524 VDD1.t4 VSUBS 0.086828f
C525 VDD1.t0 VSUBS 0.086828f
C526 VDD1.n4 VSUBS 0.525195f
C527 VDD1.n5 VSUBS 2.12259f
C528 VP.n0 VSUBS 0.052657f
C529 VP.t4 VSUBS 0.848247f
C530 VP.n1 VSUBS 0.075403f
C531 VP.n2 VSUBS 0.052657f
C532 VP.t5 VSUBS 0.848247f
C533 VP.n3 VSUBS 0.092058f
C534 VP.n4 VSUBS 0.052657f
C535 VP.n5 VSUBS 0.060347f
C536 VP.n6 VSUBS 0.052657f
C537 VP.t7 VSUBS 0.848247f
C538 VP.n7 VSUBS 0.075403f
C539 VP.n8 VSUBS 0.052657f
C540 VP.t3 VSUBS 0.848247f
C541 VP.n9 VSUBS 0.092058f
C542 VP.t1 VSUBS 1.00798f
C543 VP.t6 VSUBS 0.848247f
C544 VP.n10 VSUBS 0.459394f
C545 VP.n11 VSUBS 0.460717f
C546 VP.n12 VSUBS 0.325409f
C547 VP.n13 VSUBS 0.052657f
C548 VP.n14 VSUBS 0.042568f
C549 VP.n15 VSUBS 0.092058f
C550 VP.n16 VSUBS 0.354321f
C551 VP.n17 VSUBS 0.062285f
C552 VP.n18 VSUBS 0.052657f
C553 VP.n19 VSUBS 0.052657f
C554 VP.n20 VSUBS 0.052657f
C555 VP.n21 VSUBS 0.078337f
C556 VP.n22 VSUBS 0.060347f
C557 VP.n23 VSUBS 0.44381f
C558 VP.n24 VSUBS 1.96061f
C559 VP.t0 VSUBS 0.848247f
C560 VP.n25 VSUBS 0.44381f
C561 VP.n26 VSUBS 2.00864f
C562 VP.n27 VSUBS 0.052657f
C563 VP.n28 VSUBS 0.052657f
C564 VP.n29 VSUBS 0.078337f
C565 VP.n30 VSUBS 0.075403f
C566 VP.t2 VSUBS 0.848247f
C567 VP.n31 VSUBS 0.354321f
C568 VP.n32 VSUBS 0.062285f
C569 VP.n33 VSUBS 0.052657f
C570 VP.n34 VSUBS 0.052657f
C571 VP.n35 VSUBS 0.052657f
C572 VP.n36 VSUBS 0.042568f
C573 VP.n37 VSUBS 0.092058f
C574 VP.n38 VSUBS 0.354321f
C575 VP.n39 VSUBS 0.062285f
C576 VP.n40 VSUBS 0.052657f
C577 VP.n41 VSUBS 0.052657f
C578 VP.n42 VSUBS 0.052657f
C579 VP.n43 VSUBS 0.078337f
C580 VP.n44 VSUBS 0.060347f
C581 VP.n45 VSUBS 0.44381f
C582 VP.n46 VSUBS 0.051395f
C583 VTAIL.t10 VSUBS 0.101829f
C584 VTAIL.t14 VSUBS 0.101829f
C585 VTAIL.n0 VSUBS 0.542488f
C586 VTAIL.n1 VSUBS 0.607775f
C587 VTAIL.t11 VSUBS 0.768871f
C588 VTAIL.n2 VSUBS 0.697864f
C589 VTAIL.t4 VSUBS 0.768871f
C590 VTAIL.n3 VSUBS 0.697864f
C591 VTAIL.t1 VSUBS 0.101829f
C592 VTAIL.t7 VSUBS 0.101829f
C593 VTAIL.n4 VSUBS 0.542488f
C594 VTAIL.n5 VSUBS 0.743526f
C595 VTAIL.t6 VSUBS 0.768871f
C596 VTAIL.n6 VSUBS 1.54972f
C597 VTAIL.t15 VSUBS 0.768874f
C598 VTAIL.n7 VSUBS 1.54972f
C599 VTAIL.t9 VSUBS 0.101829f
C600 VTAIL.t8 VSUBS 0.101829f
C601 VTAIL.n8 VSUBS 0.542491f
C602 VTAIL.n9 VSUBS 0.743523f
C603 VTAIL.t12 VSUBS 0.768874f
C604 VTAIL.n10 VSUBS 0.697861f
C605 VTAIL.t5 VSUBS 0.768874f
C606 VTAIL.n11 VSUBS 0.697861f
C607 VTAIL.t3 VSUBS 0.101829f
C608 VTAIL.t2 VSUBS 0.101829f
C609 VTAIL.n12 VSUBS 0.542491f
C610 VTAIL.n13 VSUBS 0.743523f
C611 VTAIL.t0 VSUBS 0.768871f
C612 VTAIL.n14 VSUBS 1.54972f
C613 VTAIL.t13 VSUBS 0.768871f
C614 VTAIL.n15 VSUBS 1.54424f
C615 VDD2.t6 VSUBS 0.086741f
C616 VDD2.t7 VSUBS 0.086741f
C617 VDD2.n0 VSUBS 0.528054f
C618 VDD2.t5 VSUBS 0.086741f
C619 VDD2.t0 VSUBS 0.086741f
C620 VDD2.n1 VSUBS 0.528054f
C621 VDD2.n2 VSUBS 2.43979f
C622 VDD2.t3 VSUBS 0.086741f
C623 VDD2.t1 VSUBS 0.086741f
C624 VDD2.n3 VSUBS 0.524674f
C625 VDD2.n4 VSUBS 2.09069f
C626 VDD2.t2 VSUBS 0.086741f
C627 VDD2.t4 VSUBS 0.086741f
C628 VDD2.n5 VSUBS 0.528034f
C629 VN.n0 VSUBS 0.050866f
C630 VN.t2 VSUBS 0.819391f
C631 VN.n1 VSUBS 0.072838f
C632 VN.n2 VSUBS 0.050866f
C633 VN.t1 VSUBS 0.819391f
C634 VN.n3 VSUBS 0.088926f
C635 VN.t4 VSUBS 0.973692f
C636 VN.t5 VSUBS 0.819391f
C637 VN.n4 VSUBS 0.443766f
C638 VN.n5 VSUBS 0.445045f
C639 VN.n6 VSUBS 0.314339f
C640 VN.n7 VSUBS 0.050866f
C641 VN.n8 VSUBS 0.04112f
C642 VN.n9 VSUBS 0.088926f
C643 VN.n10 VSUBS 0.342267f
C644 VN.n11 VSUBS 0.060166f
C645 VN.n12 VSUBS 0.050866f
C646 VN.n13 VSUBS 0.050866f
C647 VN.n14 VSUBS 0.050866f
C648 VN.n15 VSUBS 0.075672f
C649 VN.n16 VSUBS 0.058294f
C650 VN.n17 VSUBS 0.428713f
C651 VN.n18 VSUBS 0.049647f
C652 VN.n19 VSUBS 0.050866f
C653 VN.t0 VSUBS 0.819391f
C654 VN.n20 VSUBS 0.072838f
C655 VN.n21 VSUBS 0.050866f
C656 VN.t6 VSUBS 0.819391f
C657 VN.n22 VSUBS 0.088926f
C658 VN.t3 VSUBS 0.973692f
C659 VN.t7 VSUBS 0.819391f
C660 VN.n23 VSUBS 0.443766f
C661 VN.n24 VSUBS 0.445045f
C662 VN.n25 VSUBS 0.314339f
C663 VN.n26 VSUBS 0.050866f
C664 VN.n27 VSUBS 0.04112f
C665 VN.n28 VSUBS 0.088926f
C666 VN.n29 VSUBS 0.342267f
C667 VN.n30 VSUBS 0.060166f
C668 VN.n31 VSUBS 0.050866f
C669 VN.n32 VSUBS 0.050866f
C670 VN.n33 VSUBS 0.050866f
C671 VN.n34 VSUBS 0.075672f
C672 VN.n35 VSUBS 0.058294f
C673 VN.n36 VSUBS 0.428713f
C674 VN.n37 VSUBS 1.92744f
.ends

