* NGSPICE file created from diff_pair_sample_0127.ext - technology: sky130A

.subckt diff_pair_sample_0127 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t11 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=5.0895 ps=26.88 w=13.05 l=3.48
X1 VTAIL.t3 VP.t0 VDD1.t9 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
X2 VTAIL.t8 VP.t1 VDD1.t8 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
X3 VDD2.t8 VN.t1 VTAIL.t13 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
X4 VDD2.t7 VN.t2 VTAIL.t10 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
X5 B.t11 B.t9 B.t10 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=5.0895 pd=26.88 as=0 ps=0 w=13.05 l=3.48
X6 VDD1.t7 VP.t2 VTAIL.t9 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
X7 VDD1.t6 VP.t3 VTAIL.t1 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=5.0895 ps=26.88 w=13.05 l=3.48
X8 VDD2.t6 VN.t3 VTAIL.t17 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=5.0895 ps=26.88 w=13.05 l=3.48
X9 VTAIL.t16 VN.t4 VDD2.t5 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
X10 VDD2.t4 VN.t5 VTAIL.t15 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=5.0895 pd=26.88 as=2.15325 ps=13.38 w=13.05 l=3.48
X11 B.t8 B.t6 B.t7 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=5.0895 pd=26.88 as=0 ps=0 w=13.05 l=3.48
X12 VDD1.t5 VP.t4 VTAIL.t4 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=5.0895 pd=26.88 as=2.15325 ps=13.38 w=13.05 l=3.48
X13 VDD1.t4 VP.t5 VTAIL.t6 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=5.0895 ps=26.88 w=13.05 l=3.48
X14 B.t5 B.t3 B.t4 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=5.0895 pd=26.88 as=0 ps=0 w=13.05 l=3.48
X15 VTAIL.t2 VP.t6 VDD1.t3 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
X16 B.t2 B.t0 B.t1 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=5.0895 pd=26.88 as=0 ps=0 w=13.05 l=3.48
X17 VDD2.t3 VN.t6 VTAIL.t12 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=5.0895 pd=26.88 as=2.15325 ps=13.38 w=13.05 l=3.48
X18 VTAIL.t18 VN.t7 VDD2.t2 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
X19 VDD1.t2 VP.t7 VTAIL.t0 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=5.0895 pd=26.88 as=2.15325 ps=13.38 w=13.05 l=3.48
X20 VTAIL.t7 VP.t8 VDD1.t1 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
X21 VDD1.t0 VP.t9 VTAIL.t5 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
X22 VTAIL.t14 VN.t8 VDD2.t1 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
X23 VTAIL.t19 VN.t9 VDD2.t0 w_n5542_n3578# sky130_fd_pr__pfet_01v8 ad=2.15325 pd=13.38 as=2.15325 ps=13.38 w=13.05 l=3.48
R0 VN.n100 VN.n99 161.3
R1 VN.n98 VN.n52 161.3
R2 VN.n97 VN.n96 161.3
R3 VN.n95 VN.n53 161.3
R4 VN.n94 VN.n93 161.3
R5 VN.n92 VN.n54 161.3
R6 VN.n91 VN.n90 161.3
R7 VN.n89 VN.n55 161.3
R8 VN.n88 VN.n87 161.3
R9 VN.n86 VN.n56 161.3
R10 VN.n85 VN.n84 161.3
R11 VN.n83 VN.n58 161.3
R12 VN.n82 VN.n81 161.3
R13 VN.n80 VN.n59 161.3
R14 VN.n79 VN.n78 161.3
R15 VN.n77 VN.n60 161.3
R16 VN.n76 VN.n75 161.3
R17 VN.n74 VN.n61 161.3
R18 VN.n73 VN.n72 161.3
R19 VN.n71 VN.n62 161.3
R20 VN.n70 VN.n69 161.3
R21 VN.n68 VN.n63 161.3
R22 VN.n67 VN.n66 161.3
R23 VN.n49 VN.n48 161.3
R24 VN.n47 VN.n1 161.3
R25 VN.n46 VN.n45 161.3
R26 VN.n44 VN.n2 161.3
R27 VN.n43 VN.n42 161.3
R28 VN.n41 VN.n3 161.3
R29 VN.n40 VN.n39 161.3
R30 VN.n38 VN.n4 161.3
R31 VN.n37 VN.n36 161.3
R32 VN.n34 VN.n5 161.3
R33 VN.n33 VN.n32 161.3
R34 VN.n31 VN.n6 161.3
R35 VN.n30 VN.n29 161.3
R36 VN.n28 VN.n7 161.3
R37 VN.n27 VN.n26 161.3
R38 VN.n25 VN.n8 161.3
R39 VN.n24 VN.n23 161.3
R40 VN.n22 VN.n9 161.3
R41 VN.n21 VN.n20 161.3
R42 VN.n19 VN.n10 161.3
R43 VN.n18 VN.n17 161.3
R44 VN.n16 VN.n11 161.3
R45 VN.n15 VN.n14 161.3
R46 VN.n65 VN.t3 123.005
R47 VN.n13 VN.t6 123.005
R48 VN.n8 VN.t2 90.3755
R49 VN.n12 VN.t8 90.3755
R50 VN.n35 VN.t7 90.3755
R51 VN.n0 VN.t0 90.3755
R52 VN.n60 VN.t1 90.3755
R53 VN.n64 VN.t4 90.3755
R54 VN.n57 VN.t9 90.3755
R55 VN.n51 VN.t5 90.3755
R56 VN.n50 VN.n0 84.1953
R57 VN.n101 VN.n51 84.1953
R58 VN.n13 VN.n12 59.3004
R59 VN.n65 VN.n64 59.3004
R60 VN VN.n101 58.8806
R61 VN.n42 VN.n2 56.5193
R62 VN.n93 VN.n53 56.5193
R63 VN.n21 VN.n10 49.7204
R64 VN.n29 VN.n6 49.7204
R65 VN.n73 VN.n62 49.7204
R66 VN.n81 VN.n58 49.7204
R67 VN.n17 VN.n10 31.2664
R68 VN.n33 VN.n6 31.2664
R69 VN.n69 VN.n62 31.2664
R70 VN.n85 VN.n58 31.2664
R71 VN.n16 VN.n15 24.4675
R72 VN.n17 VN.n16 24.4675
R73 VN.n22 VN.n21 24.4675
R74 VN.n23 VN.n22 24.4675
R75 VN.n23 VN.n8 24.4675
R76 VN.n27 VN.n8 24.4675
R77 VN.n28 VN.n27 24.4675
R78 VN.n29 VN.n28 24.4675
R79 VN.n34 VN.n33 24.4675
R80 VN.n36 VN.n34 24.4675
R81 VN.n40 VN.n4 24.4675
R82 VN.n41 VN.n40 24.4675
R83 VN.n42 VN.n41 24.4675
R84 VN.n46 VN.n2 24.4675
R85 VN.n47 VN.n46 24.4675
R86 VN.n48 VN.n47 24.4675
R87 VN.n69 VN.n68 24.4675
R88 VN.n68 VN.n67 24.4675
R89 VN.n81 VN.n80 24.4675
R90 VN.n80 VN.n79 24.4675
R91 VN.n79 VN.n60 24.4675
R92 VN.n75 VN.n60 24.4675
R93 VN.n75 VN.n74 24.4675
R94 VN.n74 VN.n73 24.4675
R95 VN.n93 VN.n92 24.4675
R96 VN.n92 VN.n91 24.4675
R97 VN.n91 VN.n55 24.4675
R98 VN.n87 VN.n86 24.4675
R99 VN.n86 VN.n85 24.4675
R100 VN.n99 VN.n98 24.4675
R101 VN.n98 VN.n97 24.4675
R102 VN.n97 VN.n53 24.4675
R103 VN.n15 VN.n12 15.17
R104 VN.n36 VN.n35 15.17
R105 VN.n67 VN.n64 15.17
R106 VN.n87 VN.n57 15.17
R107 VN.n35 VN.n4 9.29796
R108 VN.n57 VN.n55 9.29796
R109 VN.n48 VN.n0 5.87258
R110 VN.n99 VN.n51 5.87258
R111 VN.n66 VN.n65 3.29162
R112 VN.n14 VN.n13 3.29162
R113 VN.n101 VN.n100 0.354971
R114 VN.n50 VN.n49 0.354971
R115 VN VN.n50 0.26696
R116 VN.n100 VN.n52 0.189894
R117 VN.n96 VN.n52 0.189894
R118 VN.n96 VN.n95 0.189894
R119 VN.n95 VN.n94 0.189894
R120 VN.n94 VN.n54 0.189894
R121 VN.n90 VN.n54 0.189894
R122 VN.n90 VN.n89 0.189894
R123 VN.n89 VN.n88 0.189894
R124 VN.n88 VN.n56 0.189894
R125 VN.n84 VN.n56 0.189894
R126 VN.n84 VN.n83 0.189894
R127 VN.n83 VN.n82 0.189894
R128 VN.n82 VN.n59 0.189894
R129 VN.n78 VN.n59 0.189894
R130 VN.n78 VN.n77 0.189894
R131 VN.n77 VN.n76 0.189894
R132 VN.n76 VN.n61 0.189894
R133 VN.n72 VN.n61 0.189894
R134 VN.n72 VN.n71 0.189894
R135 VN.n71 VN.n70 0.189894
R136 VN.n70 VN.n63 0.189894
R137 VN.n66 VN.n63 0.189894
R138 VN.n14 VN.n11 0.189894
R139 VN.n18 VN.n11 0.189894
R140 VN.n19 VN.n18 0.189894
R141 VN.n20 VN.n19 0.189894
R142 VN.n20 VN.n9 0.189894
R143 VN.n24 VN.n9 0.189894
R144 VN.n25 VN.n24 0.189894
R145 VN.n26 VN.n25 0.189894
R146 VN.n26 VN.n7 0.189894
R147 VN.n30 VN.n7 0.189894
R148 VN.n31 VN.n30 0.189894
R149 VN.n32 VN.n31 0.189894
R150 VN.n32 VN.n5 0.189894
R151 VN.n37 VN.n5 0.189894
R152 VN.n38 VN.n37 0.189894
R153 VN.n39 VN.n38 0.189894
R154 VN.n39 VN.n3 0.189894
R155 VN.n43 VN.n3 0.189894
R156 VN.n44 VN.n43 0.189894
R157 VN.n45 VN.n44 0.189894
R158 VN.n45 VN.n1 0.189894
R159 VN.n49 VN.n1 0.189894
R160 VTAIL.n11 VTAIL.t17 62.1945
R161 VTAIL.n17 VTAIL.t11 62.1934
R162 VTAIL.n2 VTAIL.t6 62.1934
R163 VTAIL.n16 VTAIL.t1 62.1934
R164 VTAIL.n15 VTAIL.n14 59.7037
R165 VTAIL.n13 VTAIL.n12 59.7037
R166 VTAIL.n10 VTAIL.n9 59.7037
R167 VTAIL.n8 VTAIL.n7 59.7037
R168 VTAIL.n19 VTAIL.n18 59.7025
R169 VTAIL.n1 VTAIL.n0 59.7025
R170 VTAIL.n4 VTAIL.n3 59.7025
R171 VTAIL.n6 VTAIL.n5 59.7025
R172 VTAIL.n8 VTAIL.n6 30.1858
R173 VTAIL.n17 VTAIL.n16 26.9014
R174 VTAIL.n10 VTAIL.n8 3.28498
R175 VTAIL.n11 VTAIL.n10 3.28498
R176 VTAIL.n15 VTAIL.n13 3.28498
R177 VTAIL.n16 VTAIL.n15 3.28498
R178 VTAIL.n6 VTAIL.n4 3.28498
R179 VTAIL.n4 VTAIL.n2 3.28498
R180 VTAIL.n19 VTAIL.n17 3.28498
R181 VTAIL VTAIL.n1 2.52205
R182 VTAIL.n18 VTAIL.t10 2.4913
R183 VTAIL.n18 VTAIL.t18 2.4913
R184 VTAIL.n0 VTAIL.t12 2.4913
R185 VTAIL.n0 VTAIL.t14 2.4913
R186 VTAIL.n3 VTAIL.t9 2.4913
R187 VTAIL.n3 VTAIL.t8 2.4913
R188 VTAIL.n5 VTAIL.t0 2.4913
R189 VTAIL.n5 VTAIL.t7 2.4913
R190 VTAIL.n14 VTAIL.t5 2.4913
R191 VTAIL.n14 VTAIL.t2 2.4913
R192 VTAIL.n12 VTAIL.t4 2.4913
R193 VTAIL.n12 VTAIL.t3 2.4913
R194 VTAIL.n9 VTAIL.t13 2.4913
R195 VTAIL.n9 VTAIL.t16 2.4913
R196 VTAIL.n7 VTAIL.t15 2.4913
R197 VTAIL.n7 VTAIL.t19 2.4913
R198 VTAIL.n13 VTAIL.n11 2.11257
R199 VTAIL.n2 VTAIL.n1 2.11257
R200 VTAIL VTAIL.n19 0.763431
R201 VDD2.n1 VDD2.t3 82.1566
R202 VDD2.n4 VDD2.t4 78.8733
R203 VDD2.n3 VDD2.n2 78.7893
R204 VDD2 VDD2.n7 78.7865
R205 VDD2.n6 VDD2.n5 76.3825
R206 VDD2.n1 VDD2.n0 76.3813
R207 VDD2.n4 VDD2.n3 50.5666
R208 VDD2.n6 VDD2.n4 3.28498
R209 VDD2.n7 VDD2.t5 2.4913
R210 VDD2.n7 VDD2.t6 2.4913
R211 VDD2.n5 VDD2.t0 2.4913
R212 VDD2.n5 VDD2.t8 2.4913
R213 VDD2.n2 VDD2.t2 2.4913
R214 VDD2.n2 VDD2.t9 2.4913
R215 VDD2.n0 VDD2.t1 2.4913
R216 VDD2.n0 VDD2.t7 2.4913
R217 VDD2 VDD2.n6 0.87981
R218 VDD2.n3 VDD2.n1 0.766275
R219 VP.n32 VP.n31 161.3
R220 VP.n33 VP.n28 161.3
R221 VP.n35 VP.n34 161.3
R222 VP.n36 VP.n27 161.3
R223 VP.n38 VP.n37 161.3
R224 VP.n39 VP.n26 161.3
R225 VP.n41 VP.n40 161.3
R226 VP.n42 VP.n25 161.3
R227 VP.n44 VP.n43 161.3
R228 VP.n45 VP.n24 161.3
R229 VP.n47 VP.n46 161.3
R230 VP.n48 VP.n23 161.3
R231 VP.n50 VP.n49 161.3
R232 VP.n51 VP.n22 161.3
R233 VP.n54 VP.n53 161.3
R234 VP.n55 VP.n21 161.3
R235 VP.n57 VP.n56 161.3
R236 VP.n58 VP.n20 161.3
R237 VP.n60 VP.n59 161.3
R238 VP.n61 VP.n19 161.3
R239 VP.n63 VP.n62 161.3
R240 VP.n64 VP.n18 161.3
R241 VP.n66 VP.n65 161.3
R242 VP.n117 VP.n116 161.3
R243 VP.n115 VP.n1 161.3
R244 VP.n114 VP.n113 161.3
R245 VP.n112 VP.n2 161.3
R246 VP.n111 VP.n110 161.3
R247 VP.n109 VP.n3 161.3
R248 VP.n108 VP.n107 161.3
R249 VP.n106 VP.n4 161.3
R250 VP.n105 VP.n104 161.3
R251 VP.n102 VP.n5 161.3
R252 VP.n101 VP.n100 161.3
R253 VP.n99 VP.n6 161.3
R254 VP.n98 VP.n97 161.3
R255 VP.n96 VP.n7 161.3
R256 VP.n95 VP.n94 161.3
R257 VP.n93 VP.n8 161.3
R258 VP.n92 VP.n91 161.3
R259 VP.n90 VP.n9 161.3
R260 VP.n89 VP.n88 161.3
R261 VP.n87 VP.n10 161.3
R262 VP.n86 VP.n85 161.3
R263 VP.n84 VP.n11 161.3
R264 VP.n83 VP.n82 161.3
R265 VP.n81 VP.n80 161.3
R266 VP.n79 VP.n13 161.3
R267 VP.n78 VP.n77 161.3
R268 VP.n76 VP.n14 161.3
R269 VP.n75 VP.n74 161.3
R270 VP.n73 VP.n15 161.3
R271 VP.n72 VP.n71 161.3
R272 VP.n70 VP.n16 161.3
R273 VP.n30 VP.t4 123.004
R274 VP.n8 VP.t2 90.3755
R275 VP.n68 VP.t7 90.3755
R276 VP.n12 VP.t8 90.3755
R277 VP.n103 VP.t1 90.3755
R278 VP.n0 VP.t5 90.3755
R279 VP.n25 VP.t9 90.3755
R280 VP.n17 VP.t3 90.3755
R281 VP.n52 VP.t6 90.3755
R282 VP.n29 VP.t0 90.3755
R283 VP.n69 VP.n68 84.1953
R284 VP.n118 VP.n0 84.1953
R285 VP.n67 VP.n17 84.1953
R286 VP.n30 VP.n29 59.3004
R287 VP.n69 VP.n67 58.7152
R288 VP.n74 VP.n14 56.5193
R289 VP.n110 VP.n2 56.5193
R290 VP.n59 VP.n19 56.5193
R291 VP.n89 VP.n10 49.7204
R292 VP.n97 VP.n6 49.7204
R293 VP.n46 VP.n23 49.7204
R294 VP.n38 VP.n27 49.7204
R295 VP.n85 VP.n10 31.2664
R296 VP.n101 VP.n6 31.2664
R297 VP.n50 VP.n23 31.2664
R298 VP.n34 VP.n27 31.2664
R299 VP.n72 VP.n16 24.4675
R300 VP.n73 VP.n72 24.4675
R301 VP.n74 VP.n73 24.4675
R302 VP.n78 VP.n14 24.4675
R303 VP.n79 VP.n78 24.4675
R304 VP.n80 VP.n79 24.4675
R305 VP.n84 VP.n83 24.4675
R306 VP.n85 VP.n84 24.4675
R307 VP.n90 VP.n89 24.4675
R308 VP.n91 VP.n90 24.4675
R309 VP.n91 VP.n8 24.4675
R310 VP.n95 VP.n8 24.4675
R311 VP.n96 VP.n95 24.4675
R312 VP.n97 VP.n96 24.4675
R313 VP.n102 VP.n101 24.4675
R314 VP.n104 VP.n102 24.4675
R315 VP.n108 VP.n4 24.4675
R316 VP.n109 VP.n108 24.4675
R317 VP.n110 VP.n109 24.4675
R318 VP.n114 VP.n2 24.4675
R319 VP.n115 VP.n114 24.4675
R320 VP.n116 VP.n115 24.4675
R321 VP.n63 VP.n19 24.4675
R322 VP.n64 VP.n63 24.4675
R323 VP.n65 VP.n64 24.4675
R324 VP.n51 VP.n50 24.4675
R325 VP.n53 VP.n51 24.4675
R326 VP.n57 VP.n21 24.4675
R327 VP.n58 VP.n57 24.4675
R328 VP.n59 VP.n58 24.4675
R329 VP.n39 VP.n38 24.4675
R330 VP.n40 VP.n39 24.4675
R331 VP.n40 VP.n25 24.4675
R332 VP.n44 VP.n25 24.4675
R333 VP.n45 VP.n44 24.4675
R334 VP.n46 VP.n45 24.4675
R335 VP.n33 VP.n32 24.4675
R336 VP.n34 VP.n33 24.4675
R337 VP.n83 VP.n12 15.17
R338 VP.n104 VP.n103 15.17
R339 VP.n53 VP.n52 15.17
R340 VP.n32 VP.n29 15.17
R341 VP.n80 VP.n12 9.29796
R342 VP.n103 VP.n4 9.29796
R343 VP.n52 VP.n21 9.29796
R344 VP.n68 VP.n16 5.87258
R345 VP.n116 VP.n0 5.87258
R346 VP.n65 VP.n17 5.87258
R347 VP.n31 VP.n30 3.29161
R348 VP.n67 VP.n66 0.354971
R349 VP.n70 VP.n69 0.354971
R350 VP.n118 VP.n117 0.354971
R351 VP VP.n118 0.26696
R352 VP.n31 VP.n28 0.189894
R353 VP.n35 VP.n28 0.189894
R354 VP.n36 VP.n35 0.189894
R355 VP.n37 VP.n36 0.189894
R356 VP.n37 VP.n26 0.189894
R357 VP.n41 VP.n26 0.189894
R358 VP.n42 VP.n41 0.189894
R359 VP.n43 VP.n42 0.189894
R360 VP.n43 VP.n24 0.189894
R361 VP.n47 VP.n24 0.189894
R362 VP.n48 VP.n47 0.189894
R363 VP.n49 VP.n48 0.189894
R364 VP.n49 VP.n22 0.189894
R365 VP.n54 VP.n22 0.189894
R366 VP.n55 VP.n54 0.189894
R367 VP.n56 VP.n55 0.189894
R368 VP.n56 VP.n20 0.189894
R369 VP.n60 VP.n20 0.189894
R370 VP.n61 VP.n60 0.189894
R371 VP.n62 VP.n61 0.189894
R372 VP.n62 VP.n18 0.189894
R373 VP.n66 VP.n18 0.189894
R374 VP.n71 VP.n70 0.189894
R375 VP.n71 VP.n15 0.189894
R376 VP.n75 VP.n15 0.189894
R377 VP.n76 VP.n75 0.189894
R378 VP.n77 VP.n76 0.189894
R379 VP.n77 VP.n13 0.189894
R380 VP.n81 VP.n13 0.189894
R381 VP.n82 VP.n81 0.189894
R382 VP.n82 VP.n11 0.189894
R383 VP.n86 VP.n11 0.189894
R384 VP.n87 VP.n86 0.189894
R385 VP.n88 VP.n87 0.189894
R386 VP.n88 VP.n9 0.189894
R387 VP.n92 VP.n9 0.189894
R388 VP.n93 VP.n92 0.189894
R389 VP.n94 VP.n93 0.189894
R390 VP.n94 VP.n7 0.189894
R391 VP.n98 VP.n7 0.189894
R392 VP.n99 VP.n98 0.189894
R393 VP.n100 VP.n99 0.189894
R394 VP.n100 VP.n5 0.189894
R395 VP.n105 VP.n5 0.189894
R396 VP.n106 VP.n105 0.189894
R397 VP.n107 VP.n106 0.189894
R398 VP.n107 VP.n3 0.189894
R399 VP.n111 VP.n3 0.189894
R400 VP.n112 VP.n111 0.189894
R401 VP.n113 VP.n112 0.189894
R402 VP.n113 VP.n1 0.189894
R403 VP.n117 VP.n1 0.189894
R404 VDD1.n1 VDD1.t5 82.1578
R405 VDD1.n3 VDD1.t2 82.1566
R406 VDD1.n5 VDD1.n4 78.7893
R407 VDD1.n1 VDD1.n0 76.3825
R408 VDD1.n7 VDD1.n6 76.3814
R409 VDD1.n3 VDD1.n2 76.3813
R410 VDD1.n7 VDD1.n5 52.7918
R411 VDD1.n6 VDD1.t3 2.4913
R412 VDD1.n6 VDD1.t6 2.4913
R413 VDD1.n0 VDD1.t9 2.4913
R414 VDD1.n0 VDD1.t0 2.4913
R415 VDD1.n4 VDD1.t8 2.4913
R416 VDD1.n4 VDD1.t4 2.4913
R417 VDD1.n2 VDD1.t1 2.4913
R418 VDD1.n2 VDD1.t7 2.4913
R419 VDD1 VDD1.n7 2.40567
R420 VDD1 VDD1.n1 0.87981
R421 VDD1.n5 VDD1.n3 0.766275
R422 B.n521 B.n520 585
R423 B.n519 B.n170 585
R424 B.n518 B.n517 585
R425 B.n516 B.n171 585
R426 B.n515 B.n514 585
R427 B.n513 B.n172 585
R428 B.n512 B.n511 585
R429 B.n510 B.n173 585
R430 B.n509 B.n508 585
R431 B.n507 B.n174 585
R432 B.n506 B.n505 585
R433 B.n504 B.n175 585
R434 B.n503 B.n502 585
R435 B.n501 B.n176 585
R436 B.n500 B.n499 585
R437 B.n498 B.n177 585
R438 B.n497 B.n496 585
R439 B.n495 B.n178 585
R440 B.n494 B.n493 585
R441 B.n492 B.n179 585
R442 B.n491 B.n490 585
R443 B.n489 B.n180 585
R444 B.n488 B.n487 585
R445 B.n486 B.n181 585
R446 B.n485 B.n484 585
R447 B.n483 B.n182 585
R448 B.n482 B.n481 585
R449 B.n480 B.n183 585
R450 B.n479 B.n478 585
R451 B.n477 B.n184 585
R452 B.n476 B.n475 585
R453 B.n474 B.n185 585
R454 B.n473 B.n472 585
R455 B.n471 B.n186 585
R456 B.n470 B.n469 585
R457 B.n468 B.n187 585
R458 B.n467 B.n466 585
R459 B.n465 B.n188 585
R460 B.n464 B.n463 585
R461 B.n462 B.n189 585
R462 B.n461 B.n460 585
R463 B.n459 B.n190 585
R464 B.n458 B.n457 585
R465 B.n456 B.n191 585
R466 B.n455 B.n454 585
R467 B.n453 B.n452 585
R468 B.n451 B.n195 585
R469 B.n450 B.n449 585
R470 B.n448 B.n196 585
R471 B.n447 B.n446 585
R472 B.n445 B.n197 585
R473 B.n444 B.n443 585
R474 B.n442 B.n198 585
R475 B.n441 B.n440 585
R476 B.n438 B.n199 585
R477 B.n437 B.n436 585
R478 B.n435 B.n202 585
R479 B.n434 B.n433 585
R480 B.n432 B.n203 585
R481 B.n431 B.n430 585
R482 B.n429 B.n204 585
R483 B.n428 B.n427 585
R484 B.n426 B.n205 585
R485 B.n425 B.n424 585
R486 B.n423 B.n206 585
R487 B.n422 B.n421 585
R488 B.n420 B.n207 585
R489 B.n419 B.n418 585
R490 B.n417 B.n208 585
R491 B.n416 B.n415 585
R492 B.n414 B.n209 585
R493 B.n413 B.n412 585
R494 B.n411 B.n210 585
R495 B.n410 B.n409 585
R496 B.n408 B.n211 585
R497 B.n407 B.n406 585
R498 B.n405 B.n212 585
R499 B.n404 B.n403 585
R500 B.n402 B.n213 585
R501 B.n401 B.n400 585
R502 B.n399 B.n214 585
R503 B.n398 B.n397 585
R504 B.n396 B.n215 585
R505 B.n395 B.n394 585
R506 B.n393 B.n216 585
R507 B.n392 B.n391 585
R508 B.n390 B.n217 585
R509 B.n389 B.n388 585
R510 B.n387 B.n218 585
R511 B.n386 B.n385 585
R512 B.n384 B.n219 585
R513 B.n383 B.n382 585
R514 B.n381 B.n220 585
R515 B.n380 B.n379 585
R516 B.n378 B.n221 585
R517 B.n377 B.n376 585
R518 B.n375 B.n222 585
R519 B.n374 B.n373 585
R520 B.n372 B.n223 585
R521 B.n522 B.n169 585
R522 B.n524 B.n523 585
R523 B.n525 B.n168 585
R524 B.n527 B.n526 585
R525 B.n528 B.n167 585
R526 B.n530 B.n529 585
R527 B.n531 B.n166 585
R528 B.n533 B.n532 585
R529 B.n534 B.n165 585
R530 B.n536 B.n535 585
R531 B.n537 B.n164 585
R532 B.n539 B.n538 585
R533 B.n540 B.n163 585
R534 B.n542 B.n541 585
R535 B.n543 B.n162 585
R536 B.n545 B.n544 585
R537 B.n546 B.n161 585
R538 B.n548 B.n547 585
R539 B.n549 B.n160 585
R540 B.n551 B.n550 585
R541 B.n552 B.n159 585
R542 B.n554 B.n553 585
R543 B.n555 B.n158 585
R544 B.n557 B.n556 585
R545 B.n558 B.n157 585
R546 B.n560 B.n559 585
R547 B.n561 B.n156 585
R548 B.n563 B.n562 585
R549 B.n564 B.n155 585
R550 B.n566 B.n565 585
R551 B.n567 B.n154 585
R552 B.n569 B.n568 585
R553 B.n570 B.n153 585
R554 B.n572 B.n571 585
R555 B.n573 B.n152 585
R556 B.n575 B.n574 585
R557 B.n576 B.n151 585
R558 B.n578 B.n577 585
R559 B.n579 B.n150 585
R560 B.n581 B.n580 585
R561 B.n582 B.n149 585
R562 B.n584 B.n583 585
R563 B.n585 B.n148 585
R564 B.n587 B.n586 585
R565 B.n588 B.n147 585
R566 B.n590 B.n589 585
R567 B.n591 B.n146 585
R568 B.n593 B.n592 585
R569 B.n594 B.n145 585
R570 B.n596 B.n595 585
R571 B.n597 B.n144 585
R572 B.n599 B.n598 585
R573 B.n600 B.n143 585
R574 B.n602 B.n601 585
R575 B.n603 B.n142 585
R576 B.n605 B.n604 585
R577 B.n606 B.n141 585
R578 B.n608 B.n607 585
R579 B.n609 B.n140 585
R580 B.n611 B.n610 585
R581 B.n612 B.n139 585
R582 B.n614 B.n613 585
R583 B.n615 B.n138 585
R584 B.n617 B.n616 585
R585 B.n618 B.n137 585
R586 B.n620 B.n619 585
R587 B.n621 B.n136 585
R588 B.n623 B.n622 585
R589 B.n624 B.n135 585
R590 B.n626 B.n625 585
R591 B.n627 B.n134 585
R592 B.n629 B.n628 585
R593 B.n630 B.n133 585
R594 B.n632 B.n631 585
R595 B.n633 B.n132 585
R596 B.n635 B.n634 585
R597 B.n636 B.n131 585
R598 B.n638 B.n637 585
R599 B.n639 B.n130 585
R600 B.n641 B.n640 585
R601 B.n642 B.n129 585
R602 B.n644 B.n643 585
R603 B.n645 B.n128 585
R604 B.n647 B.n646 585
R605 B.n648 B.n127 585
R606 B.n650 B.n649 585
R607 B.n651 B.n126 585
R608 B.n653 B.n652 585
R609 B.n654 B.n125 585
R610 B.n656 B.n655 585
R611 B.n657 B.n124 585
R612 B.n659 B.n658 585
R613 B.n660 B.n123 585
R614 B.n662 B.n661 585
R615 B.n663 B.n122 585
R616 B.n665 B.n664 585
R617 B.n666 B.n121 585
R618 B.n668 B.n667 585
R619 B.n669 B.n120 585
R620 B.n671 B.n670 585
R621 B.n672 B.n119 585
R622 B.n674 B.n673 585
R623 B.n675 B.n118 585
R624 B.n677 B.n676 585
R625 B.n678 B.n117 585
R626 B.n680 B.n679 585
R627 B.n681 B.n116 585
R628 B.n683 B.n682 585
R629 B.n684 B.n115 585
R630 B.n686 B.n685 585
R631 B.n687 B.n114 585
R632 B.n689 B.n688 585
R633 B.n690 B.n113 585
R634 B.n692 B.n691 585
R635 B.n693 B.n112 585
R636 B.n695 B.n694 585
R637 B.n696 B.n111 585
R638 B.n698 B.n697 585
R639 B.n699 B.n110 585
R640 B.n701 B.n700 585
R641 B.n702 B.n109 585
R642 B.n704 B.n703 585
R643 B.n705 B.n108 585
R644 B.n707 B.n706 585
R645 B.n708 B.n107 585
R646 B.n710 B.n709 585
R647 B.n711 B.n106 585
R648 B.n713 B.n712 585
R649 B.n714 B.n105 585
R650 B.n716 B.n715 585
R651 B.n717 B.n104 585
R652 B.n719 B.n718 585
R653 B.n720 B.n103 585
R654 B.n722 B.n721 585
R655 B.n723 B.n102 585
R656 B.n725 B.n724 585
R657 B.n726 B.n101 585
R658 B.n728 B.n727 585
R659 B.n729 B.n100 585
R660 B.n731 B.n730 585
R661 B.n732 B.n99 585
R662 B.n734 B.n733 585
R663 B.n735 B.n98 585
R664 B.n737 B.n736 585
R665 B.n738 B.n97 585
R666 B.n740 B.n739 585
R667 B.n741 B.n96 585
R668 B.n743 B.n742 585
R669 B.n744 B.n95 585
R670 B.n746 B.n745 585
R671 B.n747 B.n94 585
R672 B.n749 B.n748 585
R673 B.n899 B.n898 585
R674 B.n897 B.n40 585
R675 B.n896 B.n895 585
R676 B.n894 B.n41 585
R677 B.n893 B.n892 585
R678 B.n891 B.n42 585
R679 B.n890 B.n889 585
R680 B.n888 B.n43 585
R681 B.n887 B.n886 585
R682 B.n885 B.n44 585
R683 B.n884 B.n883 585
R684 B.n882 B.n45 585
R685 B.n881 B.n880 585
R686 B.n879 B.n46 585
R687 B.n878 B.n877 585
R688 B.n876 B.n47 585
R689 B.n875 B.n874 585
R690 B.n873 B.n48 585
R691 B.n872 B.n871 585
R692 B.n870 B.n49 585
R693 B.n869 B.n868 585
R694 B.n867 B.n50 585
R695 B.n866 B.n865 585
R696 B.n864 B.n51 585
R697 B.n863 B.n862 585
R698 B.n861 B.n52 585
R699 B.n860 B.n859 585
R700 B.n858 B.n53 585
R701 B.n857 B.n856 585
R702 B.n855 B.n54 585
R703 B.n854 B.n853 585
R704 B.n852 B.n55 585
R705 B.n851 B.n850 585
R706 B.n849 B.n56 585
R707 B.n848 B.n847 585
R708 B.n846 B.n57 585
R709 B.n845 B.n844 585
R710 B.n843 B.n58 585
R711 B.n842 B.n841 585
R712 B.n840 B.n59 585
R713 B.n839 B.n838 585
R714 B.n837 B.n60 585
R715 B.n836 B.n835 585
R716 B.n834 B.n61 585
R717 B.n833 B.n832 585
R718 B.n831 B.n830 585
R719 B.n829 B.n65 585
R720 B.n828 B.n827 585
R721 B.n826 B.n66 585
R722 B.n825 B.n824 585
R723 B.n823 B.n67 585
R724 B.n822 B.n821 585
R725 B.n820 B.n68 585
R726 B.n819 B.n818 585
R727 B.n816 B.n69 585
R728 B.n815 B.n814 585
R729 B.n813 B.n72 585
R730 B.n812 B.n811 585
R731 B.n810 B.n73 585
R732 B.n809 B.n808 585
R733 B.n807 B.n74 585
R734 B.n806 B.n805 585
R735 B.n804 B.n75 585
R736 B.n803 B.n802 585
R737 B.n801 B.n76 585
R738 B.n800 B.n799 585
R739 B.n798 B.n77 585
R740 B.n797 B.n796 585
R741 B.n795 B.n78 585
R742 B.n794 B.n793 585
R743 B.n792 B.n79 585
R744 B.n791 B.n790 585
R745 B.n789 B.n80 585
R746 B.n788 B.n787 585
R747 B.n786 B.n81 585
R748 B.n785 B.n784 585
R749 B.n783 B.n82 585
R750 B.n782 B.n781 585
R751 B.n780 B.n83 585
R752 B.n779 B.n778 585
R753 B.n777 B.n84 585
R754 B.n776 B.n775 585
R755 B.n774 B.n85 585
R756 B.n773 B.n772 585
R757 B.n771 B.n86 585
R758 B.n770 B.n769 585
R759 B.n768 B.n87 585
R760 B.n767 B.n766 585
R761 B.n765 B.n88 585
R762 B.n764 B.n763 585
R763 B.n762 B.n89 585
R764 B.n761 B.n760 585
R765 B.n759 B.n90 585
R766 B.n758 B.n757 585
R767 B.n756 B.n91 585
R768 B.n755 B.n754 585
R769 B.n753 B.n92 585
R770 B.n752 B.n751 585
R771 B.n750 B.n93 585
R772 B.n900 B.n39 585
R773 B.n902 B.n901 585
R774 B.n903 B.n38 585
R775 B.n905 B.n904 585
R776 B.n906 B.n37 585
R777 B.n908 B.n907 585
R778 B.n909 B.n36 585
R779 B.n911 B.n910 585
R780 B.n912 B.n35 585
R781 B.n914 B.n913 585
R782 B.n915 B.n34 585
R783 B.n917 B.n916 585
R784 B.n918 B.n33 585
R785 B.n920 B.n919 585
R786 B.n921 B.n32 585
R787 B.n923 B.n922 585
R788 B.n924 B.n31 585
R789 B.n926 B.n925 585
R790 B.n927 B.n30 585
R791 B.n929 B.n928 585
R792 B.n930 B.n29 585
R793 B.n932 B.n931 585
R794 B.n933 B.n28 585
R795 B.n935 B.n934 585
R796 B.n936 B.n27 585
R797 B.n938 B.n937 585
R798 B.n939 B.n26 585
R799 B.n941 B.n940 585
R800 B.n942 B.n25 585
R801 B.n944 B.n943 585
R802 B.n945 B.n24 585
R803 B.n947 B.n946 585
R804 B.n948 B.n23 585
R805 B.n950 B.n949 585
R806 B.n951 B.n22 585
R807 B.n953 B.n952 585
R808 B.n954 B.n21 585
R809 B.n956 B.n955 585
R810 B.n957 B.n20 585
R811 B.n959 B.n958 585
R812 B.n960 B.n19 585
R813 B.n962 B.n961 585
R814 B.n963 B.n18 585
R815 B.n965 B.n964 585
R816 B.n966 B.n17 585
R817 B.n968 B.n967 585
R818 B.n969 B.n16 585
R819 B.n971 B.n970 585
R820 B.n972 B.n15 585
R821 B.n974 B.n973 585
R822 B.n975 B.n14 585
R823 B.n977 B.n976 585
R824 B.n978 B.n13 585
R825 B.n980 B.n979 585
R826 B.n981 B.n12 585
R827 B.n983 B.n982 585
R828 B.n984 B.n11 585
R829 B.n986 B.n985 585
R830 B.n987 B.n10 585
R831 B.n989 B.n988 585
R832 B.n990 B.n9 585
R833 B.n992 B.n991 585
R834 B.n993 B.n8 585
R835 B.n995 B.n994 585
R836 B.n996 B.n7 585
R837 B.n998 B.n997 585
R838 B.n999 B.n6 585
R839 B.n1001 B.n1000 585
R840 B.n1002 B.n5 585
R841 B.n1004 B.n1003 585
R842 B.n1005 B.n4 585
R843 B.n1007 B.n1006 585
R844 B.n1008 B.n3 585
R845 B.n1010 B.n1009 585
R846 B.n1011 B.n0 585
R847 B.n2 B.n1 585
R848 B.n261 B.n260 585
R849 B.n263 B.n262 585
R850 B.n264 B.n259 585
R851 B.n266 B.n265 585
R852 B.n267 B.n258 585
R853 B.n269 B.n268 585
R854 B.n270 B.n257 585
R855 B.n272 B.n271 585
R856 B.n273 B.n256 585
R857 B.n275 B.n274 585
R858 B.n276 B.n255 585
R859 B.n278 B.n277 585
R860 B.n279 B.n254 585
R861 B.n281 B.n280 585
R862 B.n282 B.n253 585
R863 B.n284 B.n283 585
R864 B.n285 B.n252 585
R865 B.n287 B.n286 585
R866 B.n288 B.n251 585
R867 B.n290 B.n289 585
R868 B.n291 B.n250 585
R869 B.n293 B.n292 585
R870 B.n294 B.n249 585
R871 B.n296 B.n295 585
R872 B.n297 B.n248 585
R873 B.n299 B.n298 585
R874 B.n300 B.n247 585
R875 B.n302 B.n301 585
R876 B.n303 B.n246 585
R877 B.n305 B.n304 585
R878 B.n306 B.n245 585
R879 B.n308 B.n307 585
R880 B.n309 B.n244 585
R881 B.n311 B.n310 585
R882 B.n312 B.n243 585
R883 B.n314 B.n313 585
R884 B.n315 B.n242 585
R885 B.n317 B.n316 585
R886 B.n318 B.n241 585
R887 B.n320 B.n319 585
R888 B.n321 B.n240 585
R889 B.n323 B.n322 585
R890 B.n324 B.n239 585
R891 B.n326 B.n325 585
R892 B.n327 B.n238 585
R893 B.n329 B.n328 585
R894 B.n330 B.n237 585
R895 B.n332 B.n331 585
R896 B.n333 B.n236 585
R897 B.n335 B.n334 585
R898 B.n336 B.n235 585
R899 B.n338 B.n337 585
R900 B.n339 B.n234 585
R901 B.n341 B.n340 585
R902 B.n342 B.n233 585
R903 B.n344 B.n343 585
R904 B.n345 B.n232 585
R905 B.n347 B.n346 585
R906 B.n348 B.n231 585
R907 B.n350 B.n349 585
R908 B.n351 B.n230 585
R909 B.n353 B.n352 585
R910 B.n354 B.n229 585
R911 B.n356 B.n355 585
R912 B.n357 B.n228 585
R913 B.n359 B.n358 585
R914 B.n360 B.n227 585
R915 B.n362 B.n361 585
R916 B.n363 B.n226 585
R917 B.n365 B.n364 585
R918 B.n366 B.n225 585
R919 B.n368 B.n367 585
R920 B.n369 B.n224 585
R921 B.n371 B.n370 585
R922 B.n370 B.n223 473.281
R923 B.n520 B.n169 473.281
R924 B.n748 B.n93 473.281
R925 B.n898 B.n39 473.281
R926 B.n200 B.t3 299.45
R927 B.n192 B.t6 299.45
R928 B.n70 B.t9 299.45
R929 B.n62 B.t0 299.45
R930 B.n1013 B.n1012 256.663
R931 B.n1012 B.n1011 235.042
R932 B.n1012 B.n2 235.042
R933 B.n192 B.t7 183.297
R934 B.n70 B.t11 183.297
R935 B.n200 B.t4 183.28
R936 B.n62 B.t2 183.28
R937 B.n374 B.n223 163.367
R938 B.n375 B.n374 163.367
R939 B.n376 B.n375 163.367
R940 B.n376 B.n221 163.367
R941 B.n380 B.n221 163.367
R942 B.n381 B.n380 163.367
R943 B.n382 B.n381 163.367
R944 B.n382 B.n219 163.367
R945 B.n386 B.n219 163.367
R946 B.n387 B.n386 163.367
R947 B.n388 B.n387 163.367
R948 B.n388 B.n217 163.367
R949 B.n392 B.n217 163.367
R950 B.n393 B.n392 163.367
R951 B.n394 B.n393 163.367
R952 B.n394 B.n215 163.367
R953 B.n398 B.n215 163.367
R954 B.n399 B.n398 163.367
R955 B.n400 B.n399 163.367
R956 B.n400 B.n213 163.367
R957 B.n404 B.n213 163.367
R958 B.n405 B.n404 163.367
R959 B.n406 B.n405 163.367
R960 B.n406 B.n211 163.367
R961 B.n410 B.n211 163.367
R962 B.n411 B.n410 163.367
R963 B.n412 B.n411 163.367
R964 B.n412 B.n209 163.367
R965 B.n416 B.n209 163.367
R966 B.n417 B.n416 163.367
R967 B.n418 B.n417 163.367
R968 B.n418 B.n207 163.367
R969 B.n422 B.n207 163.367
R970 B.n423 B.n422 163.367
R971 B.n424 B.n423 163.367
R972 B.n424 B.n205 163.367
R973 B.n428 B.n205 163.367
R974 B.n429 B.n428 163.367
R975 B.n430 B.n429 163.367
R976 B.n430 B.n203 163.367
R977 B.n434 B.n203 163.367
R978 B.n435 B.n434 163.367
R979 B.n436 B.n435 163.367
R980 B.n436 B.n199 163.367
R981 B.n441 B.n199 163.367
R982 B.n442 B.n441 163.367
R983 B.n443 B.n442 163.367
R984 B.n443 B.n197 163.367
R985 B.n447 B.n197 163.367
R986 B.n448 B.n447 163.367
R987 B.n449 B.n448 163.367
R988 B.n449 B.n195 163.367
R989 B.n453 B.n195 163.367
R990 B.n454 B.n453 163.367
R991 B.n454 B.n191 163.367
R992 B.n458 B.n191 163.367
R993 B.n459 B.n458 163.367
R994 B.n460 B.n459 163.367
R995 B.n460 B.n189 163.367
R996 B.n464 B.n189 163.367
R997 B.n465 B.n464 163.367
R998 B.n466 B.n465 163.367
R999 B.n466 B.n187 163.367
R1000 B.n470 B.n187 163.367
R1001 B.n471 B.n470 163.367
R1002 B.n472 B.n471 163.367
R1003 B.n472 B.n185 163.367
R1004 B.n476 B.n185 163.367
R1005 B.n477 B.n476 163.367
R1006 B.n478 B.n477 163.367
R1007 B.n478 B.n183 163.367
R1008 B.n482 B.n183 163.367
R1009 B.n483 B.n482 163.367
R1010 B.n484 B.n483 163.367
R1011 B.n484 B.n181 163.367
R1012 B.n488 B.n181 163.367
R1013 B.n489 B.n488 163.367
R1014 B.n490 B.n489 163.367
R1015 B.n490 B.n179 163.367
R1016 B.n494 B.n179 163.367
R1017 B.n495 B.n494 163.367
R1018 B.n496 B.n495 163.367
R1019 B.n496 B.n177 163.367
R1020 B.n500 B.n177 163.367
R1021 B.n501 B.n500 163.367
R1022 B.n502 B.n501 163.367
R1023 B.n502 B.n175 163.367
R1024 B.n506 B.n175 163.367
R1025 B.n507 B.n506 163.367
R1026 B.n508 B.n507 163.367
R1027 B.n508 B.n173 163.367
R1028 B.n512 B.n173 163.367
R1029 B.n513 B.n512 163.367
R1030 B.n514 B.n513 163.367
R1031 B.n514 B.n171 163.367
R1032 B.n518 B.n171 163.367
R1033 B.n519 B.n518 163.367
R1034 B.n520 B.n519 163.367
R1035 B.n748 B.n747 163.367
R1036 B.n747 B.n746 163.367
R1037 B.n746 B.n95 163.367
R1038 B.n742 B.n95 163.367
R1039 B.n742 B.n741 163.367
R1040 B.n741 B.n740 163.367
R1041 B.n740 B.n97 163.367
R1042 B.n736 B.n97 163.367
R1043 B.n736 B.n735 163.367
R1044 B.n735 B.n734 163.367
R1045 B.n734 B.n99 163.367
R1046 B.n730 B.n99 163.367
R1047 B.n730 B.n729 163.367
R1048 B.n729 B.n728 163.367
R1049 B.n728 B.n101 163.367
R1050 B.n724 B.n101 163.367
R1051 B.n724 B.n723 163.367
R1052 B.n723 B.n722 163.367
R1053 B.n722 B.n103 163.367
R1054 B.n718 B.n103 163.367
R1055 B.n718 B.n717 163.367
R1056 B.n717 B.n716 163.367
R1057 B.n716 B.n105 163.367
R1058 B.n712 B.n105 163.367
R1059 B.n712 B.n711 163.367
R1060 B.n711 B.n710 163.367
R1061 B.n710 B.n107 163.367
R1062 B.n706 B.n107 163.367
R1063 B.n706 B.n705 163.367
R1064 B.n705 B.n704 163.367
R1065 B.n704 B.n109 163.367
R1066 B.n700 B.n109 163.367
R1067 B.n700 B.n699 163.367
R1068 B.n699 B.n698 163.367
R1069 B.n698 B.n111 163.367
R1070 B.n694 B.n111 163.367
R1071 B.n694 B.n693 163.367
R1072 B.n693 B.n692 163.367
R1073 B.n692 B.n113 163.367
R1074 B.n688 B.n113 163.367
R1075 B.n688 B.n687 163.367
R1076 B.n687 B.n686 163.367
R1077 B.n686 B.n115 163.367
R1078 B.n682 B.n115 163.367
R1079 B.n682 B.n681 163.367
R1080 B.n681 B.n680 163.367
R1081 B.n680 B.n117 163.367
R1082 B.n676 B.n117 163.367
R1083 B.n676 B.n675 163.367
R1084 B.n675 B.n674 163.367
R1085 B.n674 B.n119 163.367
R1086 B.n670 B.n119 163.367
R1087 B.n670 B.n669 163.367
R1088 B.n669 B.n668 163.367
R1089 B.n668 B.n121 163.367
R1090 B.n664 B.n121 163.367
R1091 B.n664 B.n663 163.367
R1092 B.n663 B.n662 163.367
R1093 B.n662 B.n123 163.367
R1094 B.n658 B.n123 163.367
R1095 B.n658 B.n657 163.367
R1096 B.n657 B.n656 163.367
R1097 B.n656 B.n125 163.367
R1098 B.n652 B.n125 163.367
R1099 B.n652 B.n651 163.367
R1100 B.n651 B.n650 163.367
R1101 B.n650 B.n127 163.367
R1102 B.n646 B.n127 163.367
R1103 B.n646 B.n645 163.367
R1104 B.n645 B.n644 163.367
R1105 B.n644 B.n129 163.367
R1106 B.n640 B.n129 163.367
R1107 B.n640 B.n639 163.367
R1108 B.n639 B.n638 163.367
R1109 B.n638 B.n131 163.367
R1110 B.n634 B.n131 163.367
R1111 B.n634 B.n633 163.367
R1112 B.n633 B.n632 163.367
R1113 B.n632 B.n133 163.367
R1114 B.n628 B.n133 163.367
R1115 B.n628 B.n627 163.367
R1116 B.n627 B.n626 163.367
R1117 B.n626 B.n135 163.367
R1118 B.n622 B.n135 163.367
R1119 B.n622 B.n621 163.367
R1120 B.n621 B.n620 163.367
R1121 B.n620 B.n137 163.367
R1122 B.n616 B.n137 163.367
R1123 B.n616 B.n615 163.367
R1124 B.n615 B.n614 163.367
R1125 B.n614 B.n139 163.367
R1126 B.n610 B.n139 163.367
R1127 B.n610 B.n609 163.367
R1128 B.n609 B.n608 163.367
R1129 B.n608 B.n141 163.367
R1130 B.n604 B.n141 163.367
R1131 B.n604 B.n603 163.367
R1132 B.n603 B.n602 163.367
R1133 B.n602 B.n143 163.367
R1134 B.n598 B.n143 163.367
R1135 B.n598 B.n597 163.367
R1136 B.n597 B.n596 163.367
R1137 B.n596 B.n145 163.367
R1138 B.n592 B.n145 163.367
R1139 B.n592 B.n591 163.367
R1140 B.n591 B.n590 163.367
R1141 B.n590 B.n147 163.367
R1142 B.n586 B.n147 163.367
R1143 B.n586 B.n585 163.367
R1144 B.n585 B.n584 163.367
R1145 B.n584 B.n149 163.367
R1146 B.n580 B.n149 163.367
R1147 B.n580 B.n579 163.367
R1148 B.n579 B.n578 163.367
R1149 B.n578 B.n151 163.367
R1150 B.n574 B.n151 163.367
R1151 B.n574 B.n573 163.367
R1152 B.n573 B.n572 163.367
R1153 B.n572 B.n153 163.367
R1154 B.n568 B.n153 163.367
R1155 B.n568 B.n567 163.367
R1156 B.n567 B.n566 163.367
R1157 B.n566 B.n155 163.367
R1158 B.n562 B.n155 163.367
R1159 B.n562 B.n561 163.367
R1160 B.n561 B.n560 163.367
R1161 B.n560 B.n157 163.367
R1162 B.n556 B.n157 163.367
R1163 B.n556 B.n555 163.367
R1164 B.n555 B.n554 163.367
R1165 B.n554 B.n159 163.367
R1166 B.n550 B.n159 163.367
R1167 B.n550 B.n549 163.367
R1168 B.n549 B.n548 163.367
R1169 B.n548 B.n161 163.367
R1170 B.n544 B.n161 163.367
R1171 B.n544 B.n543 163.367
R1172 B.n543 B.n542 163.367
R1173 B.n542 B.n163 163.367
R1174 B.n538 B.n163 163.367
R1175 B.n538 B.n537 163.367
R1176 B.n537 B.n536 163.367
R1177 B.n536 B.n165 163.367
R1178 B.n532 B.n165 163.367
R1179 B.n532 B.n531 163.367
R1180 B.n531 B.n530 163.367
R1181 B.n530 B.n167 163.367
R1182 B.n526 B.n167 163.367
R1183 B.n526 B.n525 163.367
R1184 B.n525 B.n524 163.367
R1185 B.n524 B.n169 163.367
R1186 B.n898 B.n897 163.367
R1187 B.n897 B.n896 163.367
R1188 B.n896 B.n41 163.367
R1189 B.n892 B.n41 163.367
R1190 B.n892 B.n891 163.367
R1191 B.n891 B.n890 163.367
R1192 B.n890 B.n43 163.367
R1193 B.n886 B.n43 163.367
R1194 B.n886 B.n885 163.367
R1195 B.n885 B.n884 163.367
R1196 B.n884 B.n45 163.367
R1197 B.n880 B.n45 163.367
R1198 B.n880 B.n879 163.367
R1199 B.n879 B.n878 163.367
R1200 B.n878 B.n47 163.367
R1201 B.n874 B.n47 163.367
R1202 B.n874 B.n873 163.367
R1203 B.n873 B.n872 163.367
R1204 B.n872 B.n49 163.367
R1205 B.n868 B.n49 163.367
R1206 B.n868 B.n867 163.367
R1207 B.n867 B.n866 163.367
R1208 B.n866 B.n51 163.367
R1209 B.n862 B.n51 163.367
R1210 B.n862 B.n861 163.367
R1211 B.n861 B.n860 163.367
R1212 B.n860 B.n53 163.367
R1213 B.n856 B.n53 163.367
R1214 B.n856 B.n855 163.367
R1215 B.n855 B.n854 163.367
R1216 B.n854 B.n55 163.367
R1217 B.n850 B.n55 163.367
R1218 B.n850 B.n849 163.367
R1219 B.n849 B.n848 163.367
R1220 B.n848 B.n57 163.367
R1221 B.n844 B.n57 163.367
R1222 B.n844 B.n843 163.367
R1223 B.n843 B.n842 163.367
R1224 B.n842 B.n59 163.367
R1225 B.n838 B.n59 163.367
R1226 B.n838 B.n837 163.367
R1227 B.n837 B.n836 163.367
R1228 B.n836 B.n61 163.367
R1229 B.n832 B.n61 163.367
R1230 B.n832 B.n831 163.367
R1231 B.n831 B.n65 163.367
R1232 B.n827 B.n65 163.367
R1233 B.n827 B.n826 163.367
R1234 B.n826 B.n825 163.367
R1235 B.n825 B.n67 163.367
R1236 B.n821 B.n67 163.367
R1237 B.n821 B.n820 163.367
R1238 B.n820 B.n819 163.367
R1239 B.n819 B.n69 163.367
R1240 B.n814 B.n69 163.367
R1241 B.n814 B.n813 163.367
R1242 B.n813 B.n812 163.367
R1243 B.n812 B.n73 163.367
R1244 B.n808 B.n73 163.367
R1245 B.n808 B.n807 163.367
R1246 B.n807 B.n806 163.367
R1247 B.n806 B.n75 163.367
R1248 B.n802 B.n75 163.367
R1249 B.n802 B.n801 163.367
R1250 B.n801 B.n800 163.367
R1251 B.n800 B.n77 163.367
R1252 B.n796 B.n77 163.367
R1253 B.n796 B.n795 163.367
R1254 B.n795 B.n794 163.367
R1255 B.n794 B.n79 163.367
R1256 B.n790 B.n79 163.367
R1257 B.n790 B.n789 163.367
R1258 B.n789 B.n788 163.367
R1259 B.n788 B.n81 163.367
R1260 B.n784 B.n81 163.367
R1261 B.n784 B.n783 163.367
R1262 B.n783 B.n782 163.367
R1263 B.n782 B.n83 163.367
R1264 B.n778 B.n83 163.367
R1265 B.n778 B.n777 163.367
R1266 B.n777 B.n776 163.367
R1267 B.n776 B.n85 163.367
R1268 B.n772 B.n85 163.367
R1269 B.n772 B.n771 163.367
R1270 B.n771 B.n770 163.367
R1271 B.n770 B.n87 163.367
R1272 B.n766 B.n87 163.367
R1273 B.n766 B.n765 163.367
R1274 B.n765 B.n764 163.367
R1275 B.n764 B.n89 163.367
R1276 B.n760 B.n89 163.367
R1277 B.n760 B.n759 163.367
R1278 B.n759 B.n758 163.367
R1279 B.n758 B.n91 163.367
R1280 B.n754 B.n91 163.367
R1281 B.n754 B.n753 163.367
R1282 B.n753 B.n752 163.367
R1283 B.n752 B.n93 163.367
R1284 B.n902 B.n39 163.367
R1285 B.n903 B.n902 163.367
R1286 B.n904 B.n903 163.367
R1287 B.n904 B.n37 163.367
R1288 B.n908 B.n37 163.367
R1289 B.n909 B.n908 163.367
R1290 B.n910 B.n909 163.367
R1291 B.n910 B.n35 163.367
R1292 B.n914 B.n35 163.367
R1293 B.n915 B.n914 163.367
R1294 B.n916 B.n915 163.367
R1295 B.n916 B.n33 163.367
R1296 B.n920 B.n33 163.367
R1297 B.n921 B.n920 163.367
R1298 B.n922 B.n921 163.367
R1299 B.n922 B.n31 163.367
R1300 B.n926 B.n31 163.367
R1301 B.n927 B.n926 163.367
R1302 B.n928 B.n927 163.367
R1303 B.n928 B.n29 163.367
R1304 B.n932 B.n29 163.367
R1305 B.n933 B.n932 163.367
R1306 B.n934 B.n933 163.367
R1307 B.n934 B.n27 163.367
R1308 B.n938 B.n27 163.367
R1309 B.n939 B.n938 163.367
R1310 B.n940 B.n939 163.367
R1311 B.n940 B.n25 163.367
R1312 B.n944 B.n25 163.367
R1313 B.n945 B.n944 163.367
R1314 B.n946 B.n945 163.367
R1315 B.n946 B.n23 163.367
R1316 B.n950 B.n23 163.367
R1317 B.n951 B.n950 163.367
R1318 B.n952 B.n951 163.367
R1319 B.n952 B.n21 163.367
R1320 B.n956 B.n21 163.367
R1321 B.n957 B.n956 163.367
R1322 B.n958 B.n957 163.367
R1323 B.n958 B.n19 163.367
R1324 B.n962 B.n19 163.367
R1325 B.n963 B.n962 163.367
R1326 B.n964 B.n963 163.367
R1327 B.n964 B.n17 163.367
R1328 B.n968 B.n17 163.367
R1329 B.n969 B.n968 163.367
R1330 B.n970 B.n969 163.367
R1331 B.n970 B.n15 163.367
R1332 B.n974 B.n15 163.367
R1333 B.n975 B.n974 163.367
R1334 B.n976 B.n975 163.367
R1335 B.n976 B.n13 163.367
R1336 B.n980 B.n13 163.367
R1337 B.n981 B.n980 163.367
R1338 B.n982 B.n981 163.367
R1339 B.n982 B.n11 163.367
R1340 B.n986 B.n11 163.367
R1341 B.n987 B.n986 163.367
R1342 B.n988 B.n987 163.367
R1343 B.n988 B.n9 163.367
R1344 B.n992 B.n9 163.367
R1345 B.n993 B.n992 163.367
R1346 B.n994 B.n993 163.367
R1347 B.n994 B.n7 163.367
R1348 B.n998 B.n7 163.367
R1349 B.n999 B.n998 163.367
R1350 B.n1000 B.n999 163.367
R1351 B.n1000 B.n5 163.367
R1352 B.n1004 B.n5 163.367
R1353 B.n1005 B.n1004 163.367
R1354 B.n1006 B.n1005 163.367
R1355 B.n1006 B.n3 163.367
R1356 B.n1010 B.n3 163.367
R1357 B.n1011 B.n1010 163.367
R1358 B.n261 B.n2 163.367
R1359 B.n262 B.n261 163.367
R1360 B.n262 B.n259 163.367
R1361 B.n266 B.n259 163.367
R1362 B.n267 B.n266 163.367
R1363 B.n268 B.n267 163.367
R1364 B.n268 B.n257 163.367
R1365 B.n272 B.n257 163.367
R1366 B.n273 B.n272 163.367
R1367 B.n274 B.n273 163.367
R1368 B.n274 B.n255 163.367
R1369 B.n278 B.n255 163.367
R1370 B.n279 B.n278 163.367
R1371 B.n280 B.n279 163.367
R1372 B.n280 B.n253 163.367
R1373 B.n284 B.n253 163.367
R1374 B.n285 B.n284 163.367
R1375 B.n286 B.n285 163.367
R1376 B.n286 B.n251 163.367
R1377 B.n290 B.n251 163.367
R1378 B.n291 B.n290 163.367
R1379 B.n292 B.n291 163.367
R1380 B.n292 B.n249 163.367
R1381 B.n296 B.n249 163.367
R1382 B.n297 B.n296 163.367
R1383 B.n298 B.n297 163.367
R1384 B.n298 B.n247 163.367
R1385 B.n302 B.n247 163.367
R1386 B.n303 B.n302 163.367
R1387 B.n304 B.n303 163.367
R1388 B.n304 B.n245 163.367
R1389 B.n308 B.n245 163.367
R1390 B.n309 B.n308 163.367
R1391 B.n310 B.n309 163.367
R1392 B.n310 B.n243 163.367
R1393 B.n314 B.n243 163.367
R1394 B.n315 B.n314 163.367
R1395 B.n316 B.n315 163.367
R1396 B.n316 B.n241 163.367
R1397 B.n320 B.n241 163.367
R1398 B.n321 B.n320 163.367
R1399 B.n322 B.n321 163.367
R1400 B.n322 B.n239 163.367
R1401 B.n326 B.n239 163.367
R1402 B.n327 B.n326 163.367
R1403 B.n328 B.n327 163.367
R1404 B.n328 B.n237 163.367
R1405 B.n332 B.n237 163.367
R1406 B.n333 B.n332 163.367
R1407 B.n334 B.n333 163.367
R1408 B.n334 B.n235 163.367
R1409 B.n338 B.n235 163.367
R1410 B.n339 B.n338 163.367
R1411 B.n340 B.n339 163.367
R1412 B.n340 B.n233 163.367
R1413 B.n344 B.n233 163.367
R1414 B.n345 B.n344 163.367
R1415 B.n346 B.n345 163.367
R1416 B.n346 B.n231 163.367
R1417 B.n350 B.n231 163.367
R1418 B.n351 B.n350 163.367
R1419 B.n352 B.n351 163.367
R1420 B.n352 B.n229 163.367
R1421 B.n356 B.n229 163.367
R1422 B.n357 B.n356 163.367
R1423 B.n358 B.n357 163.367
R1424 B.n358 B.n227 163.367
R1425 B.n362 B.n227 163.367
R1426 B.n363 B.n362 163.367
R1427 B.n364 B.n363 163.367
R1428 B.n364 B.n225 163.367
R1429 B.n368 B.n225 163.367
R1430 B.n369 B.n368 163.367
R1431 B.n370 B.n369 163.367
R1432 B.n193 B.t8 109.406
R1433 B.n71 B.t10 109.406
R1434 B.n201 B.t5 109.389
R1435 B.n63 B.t1 109.389
R1436 B.n201 B.n200 73.8914
R1437 B.n193 B.n192 73.8914
R1438 B.n71 B.n70 73.8914
R1439 B.n63 B.n62 73.8914
R1440 B.n439 B.n201 59.5399
R1441 B.n194 B.n193 59.5399
R1442 B.n817 B.n71 59.5399
R1443 B.n64 B.n63 59.5399
R1444 B.n900 B.n899 30.7517
R1445 B.n750 B.n749 30.7517
R1446 B.n522 B.n521 30.7517
R1447 B.n372 B.n371 30.7517
R1448 B B.n1013 18.0485
R1449 B.n901 B.n900 10.6151
R1450 B.n901 B.n38 10.6151
R1451 B.n905 B.n38 10.6151
R1452 B.n906 B.n905 10.6151
R1453 B.n907 B.n906 10.6151
R1454 B.n907 B.n36 10.6151
R1455 B.n911 B.n36 10.6151
R1456 B.n912 B.n911 10.6151
R1457 B.n913 B.n912 10.6151
R1458 B.n913 B.n34 10.6151
R1459 B.n917 B.n34 10.6151
R1460 B.n918 B.n917 10.6151
R1461 B.n919 B.n918 10.6151
R1462 B.n919 B.n32 10.6151
R1463 B.n923 B.n32 10.6151
R1464 B.n924 B.n923 10.6151
R1465 B.n925 B.n924 10.6151
R1466 B.n925 B.n30 10.6151
R1467 B.n929 B.n30 10.6151
R1468 B.n930 B.n929 10.6151
R1469 B.n931 B.n930 10.6151
R1470 B.n931 B.n28 10.6151
R1471 B.n935 B.n28 10.6151
R1472 B.n936 B.n935 10.6151
R1473 B.n937 B.n936 10.6151
R1474 B.n937 B.n26 10.6151
R1475 B.n941 B.n26 10.6151
R1476 B.n942 B.n941 10.6151
R1477 B.n943 B.n942 10.6151
R1478 B.n943 B.n24 10.6151
R1479 B.n947 B.n24 10.6151
R1480 B.n948 B.n947 10.6151
R1481 B.n949 B.n948 10.6151
R1482 B.n949 B.n22 10.6151
R1483 B.n953 B.n22 10.6151
R1484 B.n954 B.n953 10.6151
R1485 B.n955 B.n954 10.6151
R1486 B.n955 B.n20 10.6151
R1487 B.n959 B.n20 10.6151
R1488 B.n960 B.n959 10.6151
R1489 B.n961 B.n960 10.6151
R1490 B.n961 B.n18 10.6151
R1491 B.n965 B.n18 10.6151
R1492 B.n966 B.n965 10.6151
R1493 B.n967 B.n966 10.6151
R1494 B.n967 B.n16 10.6151
R1495 B.n971 B.n16 10.6151
R1496 B.n972 B.n971 10.6151
R1497 B.n973 B.n972 10.6151
R1498 B.n973 B.n14 10.6151
R1499 B.n977 B.n14 10.6151
R1500 B.n978 B.n977 10.6151
R1501 B.n979 B.n978 10.6151
R1502 B.n979 B.n12 10.6151
R1503 B.n983 B.n12 10.6151
R1504 B.n984 B.n983 10.6151
R1505 B.n985 B.n984 10.6151
R1506 B.n985 B.n10 10.6151
R1507 B.n989 B.n10 10.6151
R1508 B.n990 B.n989 10.6151
R1509 B.n991 B.n990 10.6151
R1510 B.n991 B.n8 10.6151
R1511 B.n995 B.n8 10.6151
R1512 B.n996 B.n995 10.6151
R1513 B.n997 B.n996 10.6151
R1514 B.n997 B.n6 10.6151
R1515 B.n1001 B.n6 10.6151
R1516 B.n1002 B.n1001 10.6151
R1517 B.n1003 B.n1002 10.6151
R1518 B.n1003 B.n4 10.6151
R1519 B.n1007 B.n4 10.6151
R1520 B.n1008 B.n1007 10.6151
R1521 B.n1009 B.n1008 10.6151
R1522 B.n1009 B.n0 10.6151
R1523 B.n899 B.n40 10.6151
R1524 B.n895 B.n40 10.6151
R1525 B.n895 B.n894 10.6151
R1526 B.n894 B.n893 10.6151
R1527 B.n893 B.n42 10.6151
R1528 B.n889 B.n42 10.6151
R1529 B.n889 B.n888 10.6151
R1530 B.n888 B.n887 10.6151
R1531 B.n887 B.n44 10.6151
R1532 B.n883 B.n44 10.6151
R1533 B.n883 B.n882 10.6151
R1534 B.n882 B.n881 10.6151
R1535 B.n881 B.n46 10.6151
R1536 B.n877 B.n46 10.6151
R1537 B.n877 B.n876 10.6151
R1538 B.n876 B.n875 10.6151
R1539 B.n875 B.n48 10.6151
R1540 B.n871 B.n48 10.6151
R1541 B.n871 B.n870 10.6151
R1542 B.n870 B.n869 10.6151
R1543 B.n869 B.n50 10.6151
R1544 B.n865 B.n50 10.6151
R1545 B.n865 B.n864 10.6151
R1546 B.n864 B.n863 10.6151
R1547 B.n863 B.n52 10.6151
R1548 B.n859 B.n52 10.6151
R1549 B.n859 B.n858 10.6151
R1550 B.n858 B.n857 10.6151
R1551 B.n857 B.n54 10.6151
R1552 B.n853 B.n54 10.6151
R1553 B.n853 B.n852 10.6151
R1554 B.n852 B.n851 10.6151
R1555 B.n851 B.n56 10.6151
R1556 B.n847 B.n56 10.6151
R1557 B.n847 B.n846 10.6151
R1558 B.n846 B.n845 10.6151
R1559 B.n845 B.n58 10.6151
R1560 B.n841 B.n58 10.6151
R1561 B.n841 B.n840 10.6151
R1562 B.n840 B.n839 10.6151
R1563 B.n839 B.n60 10.6151
R1564 B.n835 B.n60 10.6151
R1565 B.n835 B.n834 10.6151
R1566 B.n834 B.n833 10.6151
R1567 B.n830 B.n829 10.6151
R1568 B.n829 B.n828 10.6151
R1569 B.n828 B.n66 10.6151
R1570 B.n824 B.n66 10.6151
R1571 B.n824 B.n823 10.6151
R1572 B.n823 B.n822 10.6151
R1573 B.n822 B.n68 10.6151
R1574 B.n818 B.n68 10.6151
R1575 B.n816 B.n815 10.6151
R1576 B.n815 B.n72 10.6151
R1577 B.n811 B.n72 10.6151
R1578 B.n811 B.n810 10.6151
R1579 B.n810 B.n809 10.6151
R1580 B.n809 B.n74 10.6151
R1581 B.n805 B.n74 10.6151
R1582 B.n805 B.n804 10.6151
R1583 B.n804 B.n803 10.6151
R1584 B.n803 B.n76 10.6151
R1585 B.n799 B.n76 10.6151
R1586 B.n799 B.n798 10.6151
R1587 B.n798 B.n797 10.6151
R1588 B.n797 B.n78 10.6151
R1589 B.n793 B.n78 10.6151
R1590 B.n793 B.n792 10.6151
R1591 B.n792 B.n791 10.6151
R1592 B.n791 B.n80 10.6151
R1593 B.n787 B.n80 10.6151
R1594 B.n787 B.n786 10.6151
R1595 B.n786 B.n785 10.6151
R1596 B.n785 B.n82 10.6151
R1597 B.n781 B.n82 10.6151
R1598 B.n781 B.n780 10.6151
R1599 B.n780 B.n779 10.6151
R1600 B.n779 B.n84 10.6151
R1601 B.n775 B.n84 10.6151
R1602 B.n775 B.n774 10.6151
R1603 B.n774 B.n773 10.6151
R1604 B.n773 B.n86 10.6151
R1605 B.n769 B.n86 10.6151
R1606 B.n769 B.n768 10.6151
R1607 B.n768 B.n767 10.6151
R1608 B.n767 B.n88 10.6151
R1609 B.n763 B.n88 10.6151
R1610 B.n763 B.n762 10.6151
R1611 B.n762 B.n761 10.6151
R1612 B.n761 B.n90 10.6151
R1613 B.n757 B.n90 10.6151
R1614 B.n757 B.n756 10.6151
R1615 B.n756 B.n755 10.6151
R1616 B.n755 B.n92 10.6151
R1617 B.n751 B.n92 10.6151
R1618 B.n751 B.n750 10.6151
R1619 B.n749 B.n94 10.6151
R1620 B.n745 B.n94 10.6151
R1621 B.n745 B.n744 10.6151
R1622 B.n744 B.n743 10.6151
R1623 B.n743 B.n96 10.6151
R1624 B.n739 B.n96 10.6151
R1625 B.n739 B.n738 10.6151
R1626 B.n738 B.n737 10.6151
R1627 B.n737 B.n98 10.6151
R1628 B.n733 B.n98 10.6151
R1629 B.n733 B.n732 10.6151
R1630 B.n732 B.n731 10.6151
R1631 B.n731 B.n100 10.6151
R1632 B.n727 B.n100 10.6151
R1633 B.n727 B.n726 10.6151
R1634 B.n726 B.n725 10.6151
R1635 B.n725 B.n102 10.6151
R1636 B.n721 B.n102 10.6151
R1637 B.n721 B.n720 10.6151
R1638 B.n720 B.n719 10.6151
R1639 B.n719 B.n104 10.6151
R1640 B.n715 B.n104 10.6151
R1641 B.n715 B.n714 10.6151
R1642 B.n714 B.n713 10.6151
R1643 B.n713 B.n106 10.6151
R1644 B.n709 B.n106 10.6151
R1645 B.n709 B.n708 10.6151
R1646 B.n708 B.n707 10.6151
R1647 B.n707 B.n108 10.6151
R1648 B.n703 B.n108 10.6151
R1649 B.n703 B.n702 10.6151
R1650 B.n702 B.n701 10.6151
R1651 B.n701 B.n110 10.6151
R1652 B.n697 B.n110 10.6151
R1653 B.n697 B.n696 10.6151
R1654 B.n696 B.n695 10.6151
R1655 B.n695 B.n112 10.6151
R1656 B.n691 B.n112 10.6151
R1657 B.n691 B.n690 10.6151
R1658 B.n690 B.n689 10.6151
R1659 B.n689 B.n114 10.6151
R1660 B.n685 B.n114 10.6151
R1661 B.n685 B.n684 10.6151
R1662 B.n684 B.n683 10.6151
R1663 B.n683 B.n116 10.6151
R1664 B.n679 B.n116 10.6151
R1665 B.n679 B.n678 10.6151
R1666 B.n678 B.n677 10.6151
R1667 B.n677 B.n118 10.6151
R1668 B.n673 B.n118 10.6151
R1669 B.n673 B.n672 10.6151
R1670 B.n672 B.n671 10.6151
R1671 B.n671 B.n120 10.6151
R1672 B.n667 B.n120 10.6151
R1673 B.n667 B.n666 10.6151
R1674 B.n666 B.n665 10.6151
R1675 B.n665 B.n122 10.6151
R1676 B.n661 B.n122 10.6151
R1677 B.n661 B.n660 10.6151
R1678 B.n660 B.n659 10.6151
R1679 B.n659 B.n124 10.6151
R1680 B.n655 B.n124 10.6151
R1681 B.n655 B.n654 10.6151
R1682 B.n654 B.n653 10.6151
R1683 B.n653 B.n126 10.6151
R1684 B.n649 B.n126 10.6151
R1685 B.n649 B.n648 10.6151
R1686 B.n648 B.n647 10.6151
R1687 B.n647 B.n128 10.6151
R1688 B.n643 B.n128 10.6151
R1689 B.n643 B.n642 10.6151
R1690 B.n642 B.n641 10.6151
R1691 B.n641 B.n130 10.6151
R1692 B.n637 B.n130 10.6151
R1693 B.n637 B.n636 10.6151
R1694 B.n636 B.n635 10.6151
R1695 B.n635 B.n132 10.6151
R1696 B.n631 B.n132 10.6151
R1697 B.n631 B.n630 10.6151
R1698 B.n630 B.n629 10.6151
R1699 B.n629 B.n134 10.6151
R1700 B.n625 B.n134 10.6151
R1701 B.n625 B.n624 10.6151
R1702 B.n624 B.n623 10.6151
R1703 B.n623 B.n136 10.6151
R1704 B.n619 B.n136 10.6151
R1705 B.n619 B.n618 10.6151
R1706 B.n618 B.n617 10.6151
R1707 B.n617 B.n138 10.6151
R1708 B.n613 B.n138 10.6151
R1709 B.n613 B.n612 10.6151
R1710 B.n612 B.n611 10.6151
R1711 B.n611 B.n140 10.6151
R1712 B.n607 B.n140 10.6151
R1713 B.n607 B.n606 10.6151
R1714 B.n606 B.n605 10.6151
R1715 B.n605 B.n142 10.6151
R1716 B.n601 B.n142 10.6151
R1717 B.n601 B.n600 10.6151
R1718 B.n600 B.n599 10.6151
R1719 B.n599 B.n144 10.6151
R1720 B.n595 B.n144 10.6151
R1721 B.n595 B.n594 10.6151
R1722 B.n594 B.n593 10.6151
R1723 B.n593 B.n146 10.6151
R1724 B.n589 B.n146 10.6151
R1725 B.n589 B.n588 10.6151
R1726 B.n588 B.n587 10.6151
R1727 B.n587 B.n148 10.6151
R1728 B.n583 B.n148 10.6151
R1729 B.n583 B.n582 10.6151
R1730 B.n582 B.n581 10.6151
R1731 B.n581 B.n150 10.6151
R1732 B.n577 B.n150 10.6151
R1733 B.n577 B.n576 10.6151
R1734 B.n576 B.n575 10.6151
R1735 B.n575 B.n152 10.6151
R1736 B.n571 B.n152 10.6151
R1737 B.n571 B.n570 10.6151
R1738 B.n570 B.n569 10.6151
R1739 B.n569 B.n154 10.6151
R1740 B.n565 B.n154 10.6151
R1741 B.n565 B.n564 10.6151
R1742 B.n564 B.n563 10.6151
R1743 B.n563 B.n156 10.6151
R1744 B.n559 B.n156 10.6151
R1745 B.n559 B.n558 10.6151
R1746 B.n558 B.n557 10.6151
R1747 B.n557 B.n158 10.6151
R1748 B.n553 B.n158 10.6151
R1749 B.n553 B.n552 10.6151
R1750 B.n552 B.n551 10.6151
R1751 B.n551 B.n160 10.6151
R1752 B.n547 B.n160 10.6151
R1753 B.n547 B.n546 10.6151
R1754 B.n546 B.n545 10.6151
R1755 B.n545 B.n162 10.6151
R1756 B.n541 B.n162 10.6151
R1757 B.n541 B.n540 10.6151
R1758 B.n540 B.n539 10.6151
R1759 B.n539 B.n164 10.6151
R1760 B.n535 B.n164 10.6151
R1761 B.n535 B.n534 10.6151
R1762 B.n534 B.n533 10.6151
R1763 B.n533 B.n166 10.6151
R1764 B.n529 B.n166 10.6151
R1765 B.n529 B.n528 10.6151
R1766 B.n528 B.n527 10.6151
R1767 B.n527 B.n168 10.6151
R1768 B.n523 B.n168 10.6151
R1769 B.n523 B.n522 10.6151
R1770 B.n260 B.n1 10.6151
R1771 B.n263 B.n260 10.6151
R1772 B.n264 B.n263 10.6151
R1773 B.n265 B.n264 10.6151
R1774 B.n265 B.n258 10.6151
R1775 B.n269 B.n258 10.6151
R1776 B.n270 B.n269 10.6151
R1777 B.n271 B.n270 10.6151
R1778 B.n271 B.n256 10.6151
R1779 B.n275 B.n256 10.6151
R1780 B.n276 B.n275 10.6151
R1781 B.n277 B.n276 10.6151
R1782 B.n277 B.n254 10.6151
R1783 B.n281 B.n254 10.6151
R1784 B.n282 B.n281 10.6151
R1785 B.n283 B.n282 10.6151
R1786 B.n283 B.n252 10.6151
R1787 B.n287 B.n252 10.6151
R1788 B.n288 B.n287 10.6151
R1789 B.n289 B.n288 10.6151
R1790 B.n289 B.n250 10.6151
R1791 B.n293 B.n250 10.6151
R1792 B.n294 B.n293 10.6151
R1793 B.n295 B.n294 10.6151
R1794 B.n295 B.n248 10.6151
R1795 B.n299 B.n248 10.6151
R1796 B.n300 B.n299 10.6151
R1797 B.n301 B.n300 10.6151
R1798 B.n301 B.n246 10.6151
R1799 B.n305 B.n246 10.6151
R1800 B.n306 B.n305 10.6151
R1801 B.n307 B.n306 10.6151
R1802 B.n307 B.n244 10.6151
R1803 B.n311 B.n244 10.6151
R1804 B.n312 B.n311 10.6151
R1805 B.n313 B.n312 10.6151
R1806 B.n313 B.n242 10.6151
R1807 B.n317 B.n242 10.6151
R1808 B.n318 B.n317 10.6151
R1809 B.n319 B.n318 10.6151
R1810 B.n319 B.n240 10.6151
R1811 B.n323 B.n240 10.6151
R1812 B.n324 B.n323 10.6151
R1813 B.n325 B.n324 10.6151
R1814 B.n325 B.n238 10.6151
R1815 B.n329 B.n238 10.6151
R1816 B.n330 B.n329 10.6151
R1817 B.n331 B.n330 10.6151
R1818 B.n331 B.n236 10.6151
R1819 B.n335 B.n236 10.6151
R1820 B.n336 B.n335 10.6151
R1821 B.n337 B.n336 10.6151
R1822 B.n337 B.n234 10.6151
R1823 B.n341 B.n234 10.6151
R1824 B.n342 B.n341 10.6151
R1825 B.n343 B.n342 10.6151
R1826 B.n343 B.n232 10.6151
R1827 B.n347 B.n232 10.6151
R1828 B.n348 B.n347 10.6151
R1829 B.n349 B.n348 10.6151
R1830 B.n349 B.n230 10.6151
R1831 B.n353 B.n230 10.6151
R1832 B.n354 B.n353 10.6151
R1833 B.n355 B.n354 10.6151
R1834 B.n355 B.n228 10.6151
R1835 B.n359 B.n228 10.6151
R1836 B.n360 B.n359 10.6151
R1837 B.n361 B.n360 10.6151
R1838 B.n361 B.n226 10.6151
R1839 B.n365 B.n226 10.6151
R1840 B.n366 B.n365 10.6151
R1841 B.n367 B.n366 10.6151
R1842 B.n367 B.n224 10.6151
R1843 B.n371 B.n224 10.6151
R1844 B.n373 B.n372 10.6151
R1845 B.n373 B.n222 10.6151
R1846 B.n377 B.n222 10.6151
R1847 B.n378 B.n377 10.6151
R1848 B.n379 B.n378 10.6151
R1849 B.n379 B.n220 10.6151
R1850 B.n383 B.n220 10.6151
R1851 B.n384 B.n383 10.6151
R1852 B.n385 B.n384 10.6151
R1853 B.n385 B.n218 10.6151
R1854 B.n389 B.n218 10.6151
R1855 B.n390 B.n389 10.6151
R1856 B.n391 B.n390 10.6151
R1857 B.n391 B.n216 10.6151
R1858 B.n395 B.n216 10.6151
R1859 B.n396 B.n395 10.6151
R1860 B.n397 B.n396 10.6151
R1861 B.n397 B.n214 10.6151
R1862 B.n401 B.n214 10.6151
R1863 B.n402 B.n401 10.6151
R1864 B.n403 B.n402 10.6151
R1865 B.n403 B.n212 10.6151
R1866 B.n407 B.n212 10.6151
R1867 B.n408 B.n407 10.6151
R1868 B.n409 B.n408 10.6151
R1869 B.n409 B.n210 10.6151
R1870 B.n413 B.n210 10.6151
R1871 B.n414 B.n413 10.6151
R1872 B.n415 B.n414 10.6151
R1873 B.n415 B.n208 10.6151
R1874 B.n419 B.n208 10.6151
R1875 B.n420 B.n419 10.6151
R1876 B.n421 B.n420 10.6151
R1877 B.n421 B.n206 10.6151
R1878 B.n425 B.n206 10.6151
R1879 B.n426 B.n425 10.6151
R1880 B.n427 B.n426 10.6151
R1881 B.n427 B.n204 10.6151
R1882 B.n431 B.n204 10.6151
R1883 B.n432 B.n431 10.6151
R1884 B.n433 B.n432 10.6151
R1885 B.n433 B.n202 10.6151
R1886 B.n437 B.n202 10.6151
R1887 B.n438 B.n437 10.6151
R1888 B.n440 B.n198 10.6151
R1889 B.n444 B.n198 10.6151
R1890 B.n445 B.n444 10.6151
R1891 B.n446 B.n445 10.6151
R1892 B.n446 B.n196 10.6151
R1893 B.n450 B.n196 10.6151
R1894 B.n451 B.n450 10.6151
R1895 B.n452 B.n451 10.6151
R1896 B.n456 B.n455 10.6151
R1897 B.n457 B.n456 10.6151
R1898 B.n457 B.n190 10.6151
R1899 B.n461 B.n190 10.6151
R1900 B.n462 B.n461 10.6151
R1901 B.n463 B.n462 10.6151
R1902 B.n463 B.n188 10.6151
R1903 B.n467 B.n188 10.6151
R1904 B.n468 B.n467 10.6151
R1905 B.n469 B.n468 10.6151
R1906 B.n469 B.n186 10.6151
R1907 B.n473 B.n186 10.6151
R1908 B.n474 B.n473 10.6151
R1909 B.n475 B.n474 10.6151
R1910 B.n475 B.n184 10.6151
R1911 B.n479 B.n184 10.6151
R1912 B.n480 B.n479 10.6151
R1913 B.n481 B.n480 10.6151
R1914 B.n481 B.n182 10.6151
R1915 B.n485 B.n182 10.6151
R1916 B.n486 B.n485 10.6151
R1917 B.n487 B.n486 10.6151
R1918 B.n487 B.n180 10.6151
R1919 B.n491 B.n180 10.6151
R1920 B.n492 B.n491 10.6151
R1921 B.n493 B.n492 10.6151
R1922 B.n493 B.n178 10.6151
R1923 B.n497 B.n178 10.6151
R1924 B.n498 B.n497 10.6151
R1925 B.n499 B.n498 10.6151
R1926 B.n499 B.n176 10.6151
R1927 B.n503 B.n176 10.6151
R1928 B.n504 B.n503 10.6151
R1929 B.n505 B.n504 10.6151
R1930 B.n505 B.n174 10.6151
R1931 B.n509 B.n174 10.6151
R1932 B.n510 B.n509 10.6151
R1933 B.n511 B.n510 10.6151
R1934 B.n511 B.n172 10.6151
R1935 B.n515 B.n172 10.6151
R1936 B.n516 B.n515 10.6151
R1937 B.n517 B.n516 10.6151
R1938 B.n517 B.n170 10.6151
R1939 B.n521 B.n170 10.6151
R1940 B.n1013 B.n0 8.11757
R1941 B.n1013 B.n1 8.11757
R1942 B.n830 B.n64 6.5566
R1943 B.n818 B.n817 6.5566
R1944 B.n440 B.n439 6.5566
R1945 B.n452 B.n194 6.5566
R1946 B.n833 B.n64 4.05904
R1947 B.n817 B.n816 4.05904
R1948 B.n439 B.n438 4.05904
R1949 B.n455 B.n194 4.05904
C0 w_n5542_n3578# VDD1 3.19559f
C1 B VN 1.51956f
C2 B VDD1 2.9072f
C3 VTAIL VN 13.130799f
C4 VDD1 VTAIL 11.211901f
C5 VP VN 9.894401f
C6 VDD1 VP 12.6973f
C7 VDD2 VN 12.1608f
C8 VDD1 VDD2 2.74804f
C9 w_n5542_n3578# B 12.3206f
C10 w_n5542_n3578# VTAIL 3.48222f
C11 B VTAIL 4.31689f
C12 w_n5542_n3578# VP 12.8725f
C13 B VP 2.74229f
C14 VP VTAIL 13.1451f
C15 w_n5542_n3578# VDD2 3.38488f
C16 B VDD2 3.05939f
C17 VDD2 VTAIL 11.2693f
C18 VP VDD2 0.69597f
C19 VDD1 VN 0.155414f
C20 w_n5542_n3578# VN 12.1483f
C21 VDD2 VSUBS 2.49327f
C22 VDD1 VSUBS 2.348135f
C23 VTAIL VSUBS 1.546175f
C24 VN VSUBS 9.18068f
C25 VP VSUBS 5.396679f
C26 B VSUBS 6.546034f
C27 w_n5542_n3578# VSUBS 0.243737p
C28 B.n0 VSUBS 0.007624f
C29 B.n1 VSUBS 0.007624f
C30 B.n2 VSUBS 0.011275f
C31 B.n3 VSUBS 0.00864f
C32 B.n4 VSUBS 0.00864f
C33 B.n5 VSUBS 0.00864f
C34 B.n6 VSUBS 0.00864f
C35 B.n7 VSUBS 0.00864f
C36 B.n8 VSUBS 0.00864f
C37 B.n9 VSUBS 0.00864f
C38 B.n10 VSUBS 0.00864f
C39 B.n11 VSUBS 0.00864f
C40 B.n12 VSUBS 0.00864f
C41 B.n13 VSUBS 0.00864f
C42 B.n14 VSUBS 0.00864f
C43 B.n15 VSUBS 0.00864f
C44 B.n16 VSUBS 0.00864f
C45 B.n17 VSUBS 0.00864f
C46 B.n18 VSUBS 0.00864f
C47 B.n19 VSUBS 0.00864f
C48 B.n20 VSUBS 0.00864f
C49 B.n21 VSUBS 0.00864f
C50 B.n22 VSUBS 0.00864f
C51 B.n23 VSUBS 0.00864f
C52 B.n24 VSUBS 0.00864f
C53 B.n25 VSUBS 0.00864f
C54 B.n26 VSUBS 0.00864f
C55 B.n27 VSUBS 0.00864f
C56 B.n28 VSUBS 0.00864f
C57 B.n29 VSUBS 0.00864f
C58 B.n30 VSUBS 0.00864f
C59 B.n31 VSUBS 0.00864f
C60 B.n32 VSUBS 0.00864f
C61 B.n33 VSUBS 0.00864f
C62 B.n34 VSUBS 0.00864f
C63 B.n35 VSUBS 0.00864f
C64 B.n36 VSUBS 0.00864f
C65 B.n37 VSUBS 0.00864f
C66 B.n38 VSUBS 0.00864f
C67 B.n39 VSUBS 0.019057f
C68 B.n40 VSUBS 0.00864f
C69 B.n41 VSUBS 0.00864f
C70 B.n42 VSUBS 0.00864f
C71 B.n43 VSUBS 0.00864f
C72 B.n44 VSUBS 0.00864f
C73 B.n45 VSUBS 0.00864f
C74 B.n46 VSUBS 0.00864f
C75 B.n47 VSUBS 0.00864f
C76 B.n48 VSUBS 0.00864f
C77 B.n49 VSUBS 0.00864f
C78 B.n50 VSUBS 0.00864f
C79 B.n51 VSUBS 0.00864f
C80 B.n52 VSUBS 0.00864f
C81 B.n53 VSUBS 0.00864f
C82 B.n54 VSUBS 0.00864f
C83 B.n55 VSUBS 0.00864f
C84 B.n56 VSUBS 0.00864f
C85 B.n57 VSUBS 0.00864f
C86 B.n58 VSUBS 0.00864f
C87 B.n59 VSUBS 0.00864f
C88 B.n60 VSUBS 0.00864f
C89 B.n61 VSUBS 0.00864f
C90 B.t1 VSUBS 0.529464f
C91 B.t2 VSUBS 0.562072f
C92 B.t0 VSUBS 2.58886f
C93 B.n62 VSUBS 0.319946f
C94 B.n63 VSUBS 0.093205f
C95 B.n64 VSUBS 0.020018f
C96 B.n65 VSUBS 0.00864f
C97 B.n66 VSUBS 0.00864f
C98 B.n67 VSUBS 0.00864f
C99 B.n68 VSUBS 0.00864f
C100 B.n69 VSUBS 0.00864f
C101 B.t10 VSUBS 0.529452f
C102 B.t11 VSUBS 0.562062f
C103 B.t9 VSUBS 2.58886f
C104 B.n70 VSUBS 0.319956f
C105 B.n71 VSUBS 0.093217f
C106 B.n72 VSUBS 0.00864f
C107 B.n73 VSUBS 0.00864f
C108 B.n74 VSUBS 0.00864f
C109 B.n75 VSUBS 0.00864f
C110 B.n76 VSUBS 0.00864f
C111 B.n77 VSUBS 0.00864f
C112 B.n78 VSUBS 0.00864f
C113 B.n79 VSUBS 0.00864f
C114 B.n80 VSUBS 0.00864f
C115 B.n81 VSUBS 0.00864f
C116 B.n82 VSUBS 0.00864f
C117 B.n83 VSUBS 0.00864f
C118 B.n84 VSUBS 0.00864f
C119 B.n85 VSUBS 0.00864f
C120 B.n86 VSUBS 0.00864f
C121 B.n87 VSUBS 0.00864f
C122 B.n88 VSUBS 0.00864f
C123 B.n89 VSUBS 0.00864f
C124 B.n90 VSUBS 0.00864f
C125 B.n91 VSUBS 0.00864f
C126 B.n92 VSUBS 0.00864f
C127 B.n93 VSUBS 0.019824f
C128 B.n94 VSUBS 0.00864f
C129 B.n95 VSUBS 0.00864f
C130 B.n96 VSUBS 0.00864f
C131 B.n97 VSUBS 0.00864f
C132 B.n98 VSUBS 0.00864f
C133 B.n99 VSUBS 0.00864f
C134 B.n100 VSUBS 0.00864f
C135 B.n101 VSUBS 0.00864f
C136 B.n102 VSUBS 0.00864f
C137 B.n103 VSUBS 0.00864f
C138 B.n104 VSUBS 0.00864f
C139 B.n105 VSUBS 0.00864f
C140 B.n106 VSUBS 0.00864f
C141 B.n107 VSUBS 0.00864f
C142 B.n108 VSUBS 0.00864f
C143 B.n109 VSUBS 0.00864f
C144 B.n110 VSUBS 0.00864f
C145 B.n111 VSUBS 0.00864f
C146 B.n112 VSUBS 0.00864f
C147 B.n113 VSUBS 0.00864f
C148 B.n114 VSUBS 0.00864f
C149 B.n115 VSUBS 0.00864f
C150 B.n116 VSUBS 0.00864f
C151 B.n117 VSUBS 0.00864f
C152 B.n118 VSUBS 0.00864f
C153 B.n119 VSUBS 0.00864f
C154 B.n120 VSUBS 0.00864f
C155 B.n121 VSUBS 0.00864f
C156 B.n122 VSUBS 0.00864f
C157 B.n123 VSUBS 0.00864f
C158 B.n124 VSUBS 0.00864f
C159 B.n125 VSUBS 0.00864f
C160 B.n126 VSUBS 0.00864f
C161 B.n127 VSUBS 0.00864f
C162 B.n128 VSUBS 0.00864f
C163 B.n129 VSUBS 0.00864f
C164 B.n130 VSUBS 0.00864f
C165 B.n131 VSUBS 0.00864f
C166 B.n132 VSUBS 0.00864f
C167 B.n133 VSUBS 0.00864f
C168 B.n134 VSUBS 0.00864f
C169 B.n135 VSUBS 0.00864f
C170 B.n136 VSUBS 0.00864f
C171 B.n137 VSUBS 0.00864f
C172 B.n138 VSUBS 0.00864f
C173 B.n139 VSUBS 0.00864f
C174 B.n140 VSUBS 0.00864f
C175 B.n141 VSUBS 0.00864f
C176 B.n142 VSUBS 0.00864f
C177 B.n143 VSUBS 0.00864f
C178 B.n144 VSUBS 0.00864f
C179 B.n145 VSUBS 0.00864f
C180 B.n146 VSUBS 0.00864f
C181 B.n147 VSUBS 0.00864f
C182 B.n148 VSUBS 0.00864f
C183 B.n149 VSUBS 0.00864f
C184 B.n150 VSUBS 0.00864f
C185 B.n151 VSUBS 0.00864f
C186 B.n152 VSUBS 0.00864f
C187 B.n153 VSUBS 0.00864f
C188 B.n154 VSUBS 0.00864f
C189 B.n155 VSUBS 0.00864f
C190 B.n156 VSUBS 0.00864f
C191 B.n157 VSUBS 0.00864f
C192 B.n158 VSUBS 0.00864f
C193 B.n159 VSUBS 0.00864f
C194 B.n160 VSUBS 0.00864f
C195 B.n161 VSUBS 0.00864f
C196 B.n162 VSUBS 0.00864f
C197 B.n163 VSUBS 0.00864f
C198 B.n164 VSUBS 0.00864f
C199 B.n165 VSUBS 0.00864f
C200 B.n166 VSUBS 0.00864f
C201 B.n167 VSUBS 0.00864f
C202 B.n168 VSUBS 0.00864f
C203 B.n169 VSUBS 0.019057f
C204 B.n170 VSUBS 0.00864f
C205 B.n171 VSUBS 0.00864f
C206 B.n172 VSUBS 0.00864f
C207 B.n173 VSUBS 0.00864f
C208 B.n174 VSUBS 0.00864f
C209 B.n175 VSUBS 0.00864f
C210 B.n176 VSUBS 0.00864f
C211 B.n177 VSUBS 0.00864f
C212 B.n178 VSUBS 0.00864f
C213 B.n179 VSUBS 0.00864f
C214 B.n180 VSUBS 0.00864f
C215 B.n181 VSUBS 0.00864f
C216 B.n182 VSUBS 0.00864f
C217 B.n183 VSUBS 0.00864f
C218 B.n184 VSUBS 0.00864f
C219 B.n185 VSUBS 0.00864f
C220 B.n186 VSUBS 0.00864f
C221 B.n187 VSUBS 0.00864f
C222 B.n188 VSUBS 0.00864f
C223 B.n189 VSUBS 0.00864f
C224 B.n190 VSUBS 0.00864f
C225 B.n191 VSUBS 0.00864f
C226 B.t8 VSUBS 0.529452f
C227 B.t7 VSUBS 0.562062f
C228 B.t6 VSUBS 2.58886f
C229 B.n192 VSUBS 0.319956f
C230 B.n193 VSUBS 0.093217f
C231 B.n194 VSUBS 0.020018f
C232 B.n195 VSUBS 0.00864f
C233 B.n196 VSUBS 0.00864f
C234 B.n197 VSUBS 0.00864f
C235 B.n198 VSUBS 0.00864f
C236 B.n199 VSUBS 0.00864f
C237 B.t5 VSUBS 0.529464f
C238 B.t4 VSUBS 0.562072f
C239 B.t3 VSUBS 2.58886f
C240 B.n200 VSUBS 0.319946f
C241 B.n201 VSUBS 0.093205f
C242 B.n202 VSUBS 0.00864f
C243 B.n203 VSUBS 0.00864f
C244 B.n204 VSUBS 0.00864f
C245 B.n205 VSUBS 0.00864f
C246 B.n206 VSUBS 0.00864f
C247 B.n207 VSUBS 0.00864f
C248 B.n208 VSUBS 0.00864f
C249 B.n209 VSUBS 0.00864f
C250 B.n210 VSUBS 0.00864f
C251 B.n211 VSUBS 0.00864f
C252 B.n212 VSUBS 0.00864f
C253 B.n213 VSUBS 0.00864f
C254 B.n214 VSUBS 0.00864f
C255 B.n215 VSUBS 0.00864f
C256 B.n216 VSUBS 0.00864f
C257 B.n217 VSUBS 0.00864f
C258 B.n218 VSUBS 0.00864f
C259 B.n219 VSUBS 0.00864f
C260 B.n220 VSUBS 0.00864f
C261 B.n221 VSUBS 0.00864f
C262 B.n222 VSUBS 0.00864f
C263 B.n223 VSUBS 0.019824f
C264 B.n224 VSUBS 0.00864f
C265 B.n225 VSUBS 0.00864f
C266 B.n226 VSUBS 0.00864f
C267 B.n227 VSUBS 0.00864f
C268 B.n228 VSUBS 0.00864f
C269 B.n229 VSUBS 0.00864f
C270 B.n230 VSUBS 0.00864f
C271 B.n231 VSUBS 0.00864f
C272 B.n232 VSUBS 0.00864f
C273 B.n233 VSUBS 0.00864f
C274 B.n234 VSUBS 0.00864f
C275 B.n235 VSUBS 0.00864f
C276 B.n236 VSUBS 0.00864f
C277 B.n237 VSUBS 0.00864f
C278 B.n238 VSUBS 0.00864f
C279 B.n239 VSUBS 0.00864f
C280 B.n240 VSUBS 0.00864f
C281 B.n241 VSUBS 0.00864f
C282 B.n242 VSUBS 0.00864f
C283 B.n243 VSUBS 0.00864f
C284 B.n244 VSUBS 0.00864f
C285 B.n245 VSUBS 0.00864f
C286 B.n246 VSUBS 0.00864f
C287 B.n247 VSUBS 0.00864f
C288 B.n248 VSUBS 0.00864f
C289 B.n249 VSUBS 0.00864f
C290 B.n250 VSUBS 0.00864f
C291 B.n251 VSUBS 0.00864f
C292 B.n252 VSUBS 0.00864f
C293 B.n253 VSUBS 0.00864f
C294 B.n254 VSUBS 0.00864f
C295 B.n255 VSUBS 0.00864f
C296 B.n256 VSUBS 0.00864f
C297 B.n257 VSUBS 0.00864f
C298 B.n258 VSUBS 0.00864f
C299 B.n259 VSUBS 0.00864f
C300 B.n260 VSUBS 0.00864f
C301 B.n261 VSUBS 0.00864f
C302 B.n262 VSUBS 0.00864f
C303 B.n263 VSUBS 0.00864f
C304 B.n264 VSUBS 0.00864f
C305 B.n265 VSUBS 0.00864f
C306 B.n266 VSUBS 0.00864f
C307 B.n267 VSUBS 0.00864f
C308 B.n268 VSUBS 0.00864f
C309 B.n269 VSUBS 0.00864f
C310 B.n270 VSUBS 0.00864f
C311 B.n271 VSUBS 0.00864f
C312 B.n272 VSUBS 0.00864f
C313 B.n273 VSUBS 0.00864f
C314 B.n274 VSUBS 0.00864f
C315 B.n275 VSUBS 0.00864f
C316 B.n276 VSUBS 0.00864f
C317 B.n277 VSUBS 0.00864f
C318 B.n278 VSUBS 0.00864f
C319 B.n279 VSUBS 0.00864f
C320 B.n280 VSUBS 0.00864f
C321 B.n281 VSUBS 0.00864f
C322 B.n282 VSUBS 0.00864f
C323 B.n283 VSUBS 0.00864f
C324 B.n284 VSUBS 0.00864f
C325 B.n285 VSUBS 0.00864f
C326 B.n286 VSUBS 0.00864f
C327 B.n287 VSUBS 0.00864f
C328 B.n288 VSUBS 0.00864f
C329 B.n289 VSUBS 0.00864f
C330 B.n290 VSUBS 0.00864f
C331 B.n291 VSUBS 0.00864f
C332 B.n292 VSUBS 0.00864f
C333 B.n293 VSUBS 0.00864f
C334 B.n294 VSUBS 0.00864f
C335 B.n295 VSUBS 0.00864f
C336 B.n296 VSUBS 0.00864f
C337 B.n297 VSUBS 0.00864f
C338 B.n298 VSUBS 0.00864f
C339 B.n299 VSUBS 0.00864f
C340 B.n300 VSUBS 0.00864f
C341 B.n301 VSUBS 0.00864f
C342 B.n302 VSUBS 0.00864f
C343 B.n303 VSUBS 0.00864f
C344 B.n304 VSUBS 0.00864f
C345 B.n305 VSUBS 0.00864f
C346 B.n306 VSUBS 0.00864f
C347 B.n307 VSUBS 0.00864f
C348 B.n308 VSUBS 0.00864f
C349 B.n309 VSUBS 0.00864f
C350 B.n310 VSUBS 0.00864f
C351 B.n311 VSUBS 0.00864f
C352 B.n312 VSUBS 0.00864f
C353 B.n313 VSUBS 0.00864f
C354 B.n314 VSUBS 0.00864f
C355 B.n315 VSUBS 0.00864f
C356 B.n316 VSUBS 0.00864f
C357 B.n317 VSUBS 0.00864f
C358 B.n318 VSUBS 0.00864f
C359 B.n319 VSUBS 0.00864f
C360 B.n320 VSUBS 0.00864f
C361 B.n321 VSUBS 0.00864f
C362 B.n322 VSUBS 0.00864f
C363 B.n323 VSUBS 0.00864f
C364 B.n324 VSUBS 0.00864f
C365 B.n325 VSUBS 0.00864f
C366 B.n326 VSUBS 0.00864f
C367 B.n327 VSUBS 0.00864f
C368 B.n328 VSUBS 0.00864f
C369 B.n329 VSUBS 0.00864f
C370 B.n330 VSUBS 0.00864f
C371 B.n331 VSUBS 0.00864f
C372 B.n332 VSUBS 0.00864f
C373 B.n333 VSUBS 0.00864f
C374 B.n334 VSUBS 0.00864f
C375 B.n335 VSUBS 0.00864f
C376 B.n336 VSUBS 0.00864f
C377 B.n337 VSUBS 0.00864f
C378 B.n338 VSUBS 0.00864f
C379 B.n339 VSUBS 0.00864f
C380 B.n340 VSUBS 0.00864f
C381 B.n341 VSUBS 0.00864f
C382 B.n342 VSUBS 0.00864f
C383 B.n343 VSUBS 0.00864f
C384 B.n344 VSUBS 0.00864f
C385 B.n345 VSUBS 0.00864f
C386 B.n346 VSUBS 0.00864f
C387 B.n347 VSUBS 0.00864f
C388 B.n348 VSUBS 0.00864f
C389 B.n349 VSUBS 0.00864f
C390 B.n350 VSUBS 0.00864f
C391 B.n351 VSUBS 0.00864f
C392 B.n352 VSUBS 0.00864f
C393 B.n353 VSUBS 0.00864f
C394 B.n354 VSUBS 0.00864f
C395 B.n355 VSUBS 0.00864f
C396 B.n356 VSUBS 0.00864f
C397 B.n357 VSUBS 0.00864f
C398 B.n358 VSUBS 0.00864f
C399 B.n359 VSUBS 0.00864f
C400 B.n360 VSUBS 0.00864f
C401 B.n361 VSUBS 0.00864f
C402 B.n362 VSUBS 0.00864f
C403 B.n363 VSUBS 0.00864f
C404 B.n364 VSUBS 0.00864f
C405 B.n365 VSUBS 0.00864f
C406 B.n366 VSUBS 0.00864f
C407 B.n367 VSUBS 0.00864f
C408 B.n368 VSUBS 0.00864f
C409 B.n369 VSUBS 0.00864f
C410 B.n370 VSUBS 0.019057f
C411 B.n371 VSUBS 0.019057f
C412 B.n372 VSUBS 0.019824f
C413 B.n373 VSUBS 0.00864f
C414 B.n374 VSUBS 0.00864f
C415 B.n375 VSUBS 0.00864f
C416 B.n376 VSUBS 0.00864f
C417 B.n377 VSUBS 0.00864f
C418 B.n378 VSUBS 0.00864f
C419 B.n379 VSUBS 0.00864f
C420 B.n380 VSUBS 0.00864f
C421 B.n381 VSUBS 0.00864f
C422 B.n382 VSUBS 0.00864f
C423 B.n383 VSUBS 0.00864f
C424 B.n384 VSUBS 0.00864f
C425 B.n385 VSUBS 0.00864f
C426 B.n386 VSUBS 0.00864f
C427 B.n387 VSUBS 0.00864f
C428 B.n388 VSUBS 0.00864f
C429 B.n389 VSUBS 0.00864f
C430 B.n390 VSUBS 0.00864f
C431 B.n391 VSUBS 0.00864f
C432 B.n392 VSUBS 0.00864f
C433 B.n393 VSUBS 0.00864f
C434 B.n394 VSUBS 0.00864f
C435 B.n395 VSUBS 0.00864f
C436 B.n396 VSUBS 0.00864f
C437 B.n397 VSUBS 0.00864f
C438 B.n398 VSUBS 0.00864f
C439 B.n399 VSUBS 0.00864f
C440 B.n400 VSUBS 0.00864f
C441 B.n401 VSUBS 0.00864f
C442 B.n402 VSUBS 0.00864f
C443 B.n403 VSUBS 0.00864f
C444 B.n404 VSUBS 0.00864f
C445 B.n405 VSUBS 0.00864f
C446 B.n406 VSUBS 0.00864f
C447 B.n407 VSUBS 0.00864f
C448 B.n408 VSUBS 0.00864f
C449 B.n409 VSUBS 0.00864f
C450 B.n410 VSUBS 0.00864f
C451 B.n411 VSUBS 0.00864f
C452 B.n412 VSUBS 0.00864f
C453 B.n413 VSUBS 0.00864f
C454 B.n414 VSUBS 0.00864f
C455 B.n415 VSUBS 0.00864f
C456 B.n416 VSUBS 0.00864f
C457 B.n417 VSUBS 0.00864f
C458 B.n418 VSUBS 0.00864f
C459 B.n419 VSUBS 0.00864f
C460 B.n420 VSUBS 0.00864f
C461 B.n421 VSUBS 0.00864f
C462 B.n422 VSUBS 0.00864f
C463 B.n423 VSUBS 0.00864f
C464 B.n424 VSUBS 0.00864f
C465 B.n425 VSUBS 0.00864f
C466 B.n426 VSUBS 0.00864f
C467 B.n427 VSUBS 0.00864f
C468 B.n428 VSUBS 0.00864f
C469 B.n429 VSUBS 0.00864f
C470 B.n430 VSUBS 0.00864f
C471 B.n431 VSUBS 0.00864f
C472 B.n432 VSUBS 0.00864f
C473 B.n433 VSUBS 0.00864f
C474 B.n434 VSUBS 0.00864f
C475 B.n435 VSUBS 0.00864f
C476 B.n436 VSUBS 0.00864f
C477 B.n437 VSUBS 0.00864f
C478 B.n438 VSUBS 0.005972f
C479 B.n439 VSUBS 0.020018f
C480 B.n440 VSUBS 0.006988f
C481 B.n441 VSUBS 0.00864f
C482 B.n442 VSUBS 0.00864f
C483 B.n443 VSUBS 0.00864f
C484 B.n444 VSUBS 0.00864f
C485 B.n445 VSUBS 0.00864f
C486 B.n446 VSUBS 0.00864f
C487 B.n447 VSUBS 0.00864f
C488 B.n448 VSUBS 0.00864f
C489 B.n449 VSUBS 0.00864f
C490 B.n450 VSUBS 0.00864f
C491 B.n451 VSUBS 0.00864f
C492 B.n452 VSUBS 0.006988f
C493 B.n453 VSUBS 0.00864f
C494 B.n454 VSUBS 0.00864f
C495 B.n455 VSUBS 0.005972f
C496 B.n456 VSUBS 0.00864f
C497 B.n457 VSUBS 0.00864f
C498 B.n458 VSUBS 0.00864f
C499 B.n459 VSUBS 0.00864f
C500 B.n460 VSUBS 0.00864f
C501 B.n461 VSUBS 0.00864f
C502 B.n462 VSUBS 0.00864f
C503 B.n463 VSUBS 0.00864f
C504 B.n464 VSUBS 0.00864f
C505 B.n465 VSUBS 0.00864f
C506 B.n466 VSUBS 0.00864f
C507 B.n467 VSUBS 0.00864f
C508 B.n468 VSUBS 0.00864f
C509 B.n469 VSUBS 0.00864f
C510 B.n470 VSUBS 0.00864f
C511 B.n471 VSUBS 0.00864f
C512 B.n472 VSUBS 0.00864f
C513 B.n473 VSUBS 0.00864f
C514 B.n474 VSUBS 0.00864f
C515 B.n475 VSUBS 0.00864f
C516 B.n476 VSUBS 0.00864f
C517 B.n477 VSUBS 0.00864f
C518 B.n478 VSUBS 0.00864f
C519 B.n479 VSUBS 0.00864f
C520 B.n480 VSUBS 0.00864f
C521 B.n481 VSUBS 0.00864f
C522 B.n482 VSUBS 0.00864f
C523 B.n483 VSUBS 0.00864f
C524 B.n484 VSUBS 0.00864f
C525 B.n485 VSUBS 0.00864f
C526 B.n486 VSUBS 0.00864f
C527 B.n487 VSUBS 0.00864f
C528 B.n488 VSUBS 0.00864f
C529 B.n489 VSUBS 0.00864f
C530 B.n490 VSUBS 0.00864f
C531 B.n491 VSUBS 0.00864f
C532 B.n492 VSUBS 0.00864f
C533 B.n493 VSUBS 0.00864f
C534 B.n494 VSUBS 0.00864f
C535 B.n495 VSUBS 0.00864f
C536 B.n496 VSUBS 0.00864f
C537 B.n497 VSUBS 0.00864f
C538 B.n498 VSUBS 0.00864f
C539 B.n499 VSUBS 0.00864f
C540 B.n500 VSUBS 0.00864f
C541 B.n501 VSUBS 0.00864f
C542 B.n502 VSUBS 0.00864f
C543 B.n503 VSUBS 0.00864f
C544 B.n504 VSUBS 0.00864f
C545 B.n505 VSUBS 0.00864f
C546 B.n506 VSUBS 0.00864f
C547 B.n507 VSUBS 0.00864f
C548 B.n508 VSUBS 0.00864f
C549 B.n509 VSUBS 0.00864f
C550 B.n510 VSUBS 0.00864f
C551 B.n511 VSUBS 0.00864f
C552 B.n512 VSUBS 0.00864f
C553 B.n513 VSUBS 0.00864f
C554 B.n514 VSUBS 0.00864f
C555 B.n515 VSUBS 0.00864f
C556 B.n516 VSUBS 0.00864f
C557 B.n517 VSUBS 0.00864f
C558 B.n518 VSUBS 0.00864f
C559 B.n519 VSUBS 0.00864f
C560 B.n520 VSUBS 0.019824f
C561 B.n521 VSUBS 0.01874f
C562 B.n522 VSUBS 0.020141f
C563 B.n523 VSUBS 0.00864f
C564 B.n524 VSUBS 0.00864f
C565 B.n525 VSUBS 0.00864f
C566 B.n526 VSUBS 0.00864f
C567 B.n527 VSUBS 0.00864f
C568 B.n528 VSUBS 0.00864f
C569 B.n529 VSUBS 0.00864f
C570 B.n530 VSUBS 0.00864f
C571 B.n531 VSUBS 0.00864f
C572 B.n532 VSUBS 0.00864f
C573 B.n533 VSUBS 0.00864f
C574 B.n534 VSUBS 0.00864f
C575 B.n535 VSUBS 0.00864f
C576 B.n536 VSUBS 0.00864f
C577 B.n537 VSUBS 0.00864f
C578 B.n538 VSUBS 0.00864f
C579 B.n539 VSUBS 0.00864f
C580 B.n540 VSUBS 0.00864f
C581 B.n541 VSUBS 0.00864f
C582 B.n542 VSUBS 0.00864f
C583 B.n543 VSUBS 0.00864f
C584 B.n544 VSUBS 0.00864f
C585 B.n545 VSUBS 0.00864f
C586 B.n546 VSUBS 0.00864f
C587 B.n547 VSUBS 0.00864f
C588 B.n548 VSUBS 0.00864f
C589 B.n549 VSUBS 0.00864f
C590 B.n550 VSUBS 0.00864f
C591 B.n551 VSUBS 0.00864f
C592 B.n552 VSUBS 0.00864f
C593 B.n553 VSUBS 0.00864f
C594 B.n554 VSUBS 0.00864f
C595 B.n555 VSUBS 0.00864f
C596 B.n556 VSUBS 0.00864f
C597 B.n557 VSUBS 0.00864f
C598 B.n558 VSUBS 0.00864f
C599 B.n559 VSUBS 0.00864f
C600 B.n560 VSUBS 0.00864f
C601 B.n561 VSUBS 0.00864f
C602 B.n562 VSUBS 0.00864f
C603 B.n563 VSUBS 0.00864f
C604 B.n564 VSUBS 0.00864f
C605 B.n565 VSUBS 0.00864f
C606 B.n566 VSUBS 0.00864f
C607 B.n567 VSUBS 0.00864f
C608 B.n568 VSUBS 0.00864f
C609 B.n569 VSUBS 0.00864f
C610 B.n570 VSUBS 0.00864f
C611 B.n571 VSUBS 0.00864f
C612 B.n572 VSUBS 0.00864f
C613 B.n573 VSUBS 0.00864f
C614 B.n574 VSUBS 0.00864f
C615 B.n575 VSUBS 0.00864f
C616 B.n576 VSUBS 0.00864f
C617 B.n577 VSUBS 0.00864f
C618 B.n578 VSUBS 0.00864f
C619 B.n579 VSUBS 0.00864f
C620 B.n580 VSUBS 0.00864f
C621 B.n581 VSUBS 0.00864f
C622 B.n582 VSUBS 0.00864f
C623 B.n583 VSUBS 0.00864f
C624 B.n584 VSUBS 0.00864f
C625 B.n585 VSUBS 0.00864f
C626 B.n586 VSUBS 0.00864f
C627 B.n587 VSUBS 0.00864f
C628 B.n588 VSUBS 0.00864f
C629 B.n589 VSUBS 0.00864f
C630 B.n590 VSUBS 0.00864f
C631 B.n591 VSUBS 0.00864f
C632 B.n592 VSUBS 0.00864f
C633 B.n593 VSUBS 0.00864f
C634 B.n594 VSUBS 0.00864f
C635 B.n595 VSUBS 0.00864f
C636 B.n596 VSUBS 0.00864f
C637 B.n597 VSUBS 0.00864f
C638 B.n598 VSUBS 0.00864f
C639 B.n599 VSUBS 0.00864f
C640 B.n600 VSUBS 0.00864f
C641 B.n601 VSUBS 0.00864f
C642 B.n602 VSUBS 0.00864f
C643 B.n603 VSUBS 0.00864f
C644 B.n604 VSUBS 0.00864f
C645 B.n605 VSUBS 0.00864f
C646 B.n606 VSUBS 0.00864f
C647 B.n607 VSUBS 0.00864f
C648 B.n608 VSUBS 0.00864f
C649 B.n609 VSUBS 0.00864f
C650 B.n610 VSUBS 0.00864f
C651 B.n611 VSUBS 0.00864f
C652 B.n612 VSUBS 0.00864f
C653 B.n613 VSUBS 0.00864f
C654 B.n614 VSUBS 0.00864f
C655 B.n615 VSUBS 0.00864f
C656 B.n616 VSUBS 0.00864f
C657 B.n617 VSUBS 0.00864f
C658 B.n618 VSUBS 0.00864f
C659 B.n619 VSUBS 0.00864f
C660 B.n620 VSUBS 0.00864f
C661 B.n621 VSUBS 0.00864f
C662 B.n622 VSUBS 0.00864f
C663 B.n623 VSUBS 0.00864f
C664 B.n624 VSUBS 0.00864f
C665 B.n625 VSUBS 0.00864f
C666 B.n626 VSUBS 0.00864f
C667 B.n627 VSUBS 0.00864f
C668 B.n628 VSUBS 0.00864f
C669 B.n629 VSUBS 0.00864f
C670 B.n630 VSUBS 0.00864f
C671 B.n631 VSUBS 0.00864f
C672 B.n632 VSUBS 0.00864f
C673 B.n633 VSUBS 0.00864f
C674 B.n634 VSUBS 0.00864f
C675 B.n635 VSUBS 0.00864f
C676 B.n636 VSUBS 0.00864f
C677 B.n637 VSUBS 0.00864f
C678 B.n638 VSUBS 0.00864f
C679 B.n639 VSUBS 0.00864f
C680 B.n640 VSUBS 0.00864f
C681 B.n641 VSUBS 0.00864f
C682 B.n642 VSUBS 0.00864f
C683 B.n643 VSUBS 0.00864f
C684 B.n644 VSUBS 0.00864f
C685 B.n645 VSUBS 0.00864f
C686 B.n646 VSUBS 0.00864f
C687 B.n647 VSUBS 0.00864f
C688 B.n648 VSUBS 0.00864f
C689 B.n649 VSUBS 0.00864f
C690 B.n650 VSUBS 0.00864f
C691 B.n651 VSUBS 0.00864f
C692 B.n652 VSUBS 0.00864f
C693 B.n653 VSUBS 0.00864f
C694 B.n654 VSUBS 0.00864f
C695 B.n655 VSUBS 0.00864f
C696 B.n656 VSUBS 0.00864f
C697 B.n657 VSUBS 0.00864f
C698 B.n658 VSUBS 0.00864f
C699 B.n659 VSUBS 0.00864f
C700 B.n660 VSUBS 0.00864f
C701 B.n661 VSUBS 0.00864f
C702 B.n662 VSUBS 0.00864f
C703 B.n663 VSUBS 0.00864f
C704 B.n664 VSUBS 0.00864f
C705 B.n665 VSUBS 0.00864f
C706 B.n666 VSUBS 0.00864f
C707 B.n667 VSUBS 0.00864f
C708 B.n668 VSUBS 0.00864f
C709 B.n669 VSUBS 0.00864f
C710 B.n670 VSUBS 0.00864f
C711 B.n671 VSUBS 0.00864f
C712 B.n672 VSUBS 0.00864f
C713 B.n673 VSUBS 0.00864f
C714 B.n674 VSUBS 0.00864f
C715 B.n675 VSUBS 0.00864f
C716 B.n676 VSUBS 0.00864f
C717 B.n677 VSUBS 0.00864f
C718 B.n678 VSUBS 0.00864f
C719 B.n679 VSUBS 0.00864f
C720 B.n680 VSUBS 0.00864f
C721 B.n681 VSUBS 0.00864f
C722 B.n682 VSUBS 0.00864f
C723 B.n683 VSUBS 0.00864f
C724 B.n684 VSUBS 0.00864f
C725 B.n685 VSUBS 0.00864f
C726 B.n686 VSUBS 0.00864f
C727 B.n687 VSUBS 0.00864f
C728 B.n688 VSUBS 0.00864f
C729 B.n689 VSUBS 0.00864f
C730 B.n690 VSUBS 0.00864f
C731 B.n691 VSUBS 0.00864f
C732 B.n692 VSUBS 0.00864f
C733 B.n693 VSUBS 0.00864f
C734 B.n694 VSUBS 0.00864f
C735 B.n695 VSUBS 0.00864f
C736 B.n696 VSUBS 0.00864f
C737 B.n697 VSUBS 0.00864f
C738 B.n698 VSUBS 0.00864f
C739 B.n699 VSUBS 0.00864f
C740 B.n700 VSUBS 0.00864f
C741 B.n701 VSUBS 0.00864f
C742 B.n702 VSUBS 0.00864f
C743 B.n703 VSUBS 0.00864f
C744 B.n704 VSUBS 0.00864f
C745 B.n705 VSUBS 0.00864f
C746 B.n706 VSUBS 0.00864f
C747 B.n707 VSUBS 0.00864f
C748 B.n708 VSUBS 0.00864f
C749 B.n709 VSUBS 0.00864f
C750 B.n710 VSUBS 0.00864f
C751 B.n711 VSUBS 0.00864f
C752 B.n712 VSUBS 0.00864f
C753 B.n713 VSUBS 0.00864f
C754 B.n714 VSUBS 0.00864f
C755 B.n715 VSUBS 0.00864f
C756 B.n716 VSUBS 0.00864f
C757 B.n717 VSUBS 0.00864f
C758 B.n718 VSUBS 0.00864f
C759 B.n719 VSUBS 0.00864f
C760 B.n720 VSUBS 0.00864f
C761 B.n721 VSUBS 0.00864f
C762 B.n722 VSUBS 0.00864f
C763 B.n723 VSUBS 0.00864f
C764 B.n724 VSUBS 0.00864f
C765 B.n725 VSUBS 0.00864f
C766 B.n726 VSUBS 0.00864f
C767 B.n727 VSUBS 0.00864f
C768 B.n728 VSUBS 0.00864f
C769 B.n729 VSUBS 0.00864f
C770 B.n730 VSUBS 0.00864f
C771 B.n731 VSUBS 0.00864f
C772 B.n732 VSUBS 0.00864f
C773 B.n733 VSUBS 0.00864f
C774 B.n734 VSUBS 0.00864f
C775 B.n735 VSUBS 0.00864f
C776 B.n736 VSUBS 0.00864f
C777 B.n737 VSUBS 0.00864f
C778 B.n738 VSUBS 0.00864f
C779 B.n739 VSUBS 0.00864f
C780 B.n740 VSUBS 0.00864f
C781 B.n741 VSUBS 0.00864f
C782 B.n742 VSUBS 0.00864f
C783 B.n743 VSUBS 0.00864f
C784 B.n744 VSUBS 0.00864f
C785 B.n745 VSUBS 0.00864f
C786 B.n746 VSUBS 0.00864f
C787 B.n747 VSUBS 0.00864f
C788 B.n748 VSUBS 0.019057f
C789 B.n749 VSUBS 0.019057f
C790 B.n750 VSUBS 0.019824f
C791 B.n751 VSUBS 0.00864f
C792 B.n752 VSUBS 0.00864f
C793 B.n753 VSUBS 0.00864f
C794 B.n754 VSUBS 0.00864f
C795 B.n755 VSUBS 0.00864f
C796 B.n756 VSUBS 0.00864f
C797 B.n757 VSUBS 0.00864f
C798 B.n758 VSUBS 0.00864f
C799 B.n759 VSUBS 0.00864f
C800 B.n760 VSUBS 0.00864f
C801 B.n761 VSUBS 0.00864f
C802 B.n762 VSUBS 0.00864f
C803 B.n763 VSUBS 0.00864f
C804 B.n764 VSUBS 0.00864f
C805 B.n765 VSUBS 0.00864f
C806 B.n766 VSUBS 0.00864f
C807 B.n767 VSUBS 0.00864f
C808 B.n768 VSUBS 0.00864f
C809 B.n769 VSUBS 0.00864f
C810 B.n770 VSUBS 0.00864f
C811 B.n771 VSUBS 0.00864f
C812 B.n772 VSUBS 0.00864f
C813 B.n773 VSUBS 0.00864f
C814 B.n774 VSUBS 0.00864f
C815 B.n775 VSUBS 0.00864f
C816 B.n776 VSUBS 0.00864f
C817 B.n777 VSUBS 0.00864f
C818 B.n778 VSUBS 0.00864f
C819 B.n779 VSUBS 0.00864f
C820 B.n780 VSUBS 0.00864f
C821 B.n781 VSUBS 0.00864f
C822 B.n782 VSUBS 0.00864f
C823 B.n783 VSUBS 0.00864f
C824 B.n784 VSUBS 0.00864f
C825 B.n785 VSUBS 0.00864f
C826 B.n786 VSUBS 0.00864f
C827 B.n787 VSUBS 0.00864f
C828 B.n788 VSUBS 0.00864f
C829 B.n789 VSUBS 0.00864f
C830 B.n790 VSUBS 0.00864f
C831 B.n791 VSUBS 0.00864f
C832 B.n792 VSUBS 0.00864f
C833 B.n793 VSUBS 0.00864f
C834 B.n794 VSUBS 0.00864f
C835 B.n795 VSUBS 0.00864f
C836 B.n796 VSUBS 0.00864f
C837 B.n797 VSUBS 0.00864f
C838 B.n798 VSUBS 0.00864f
C839 B.n799 VSUBS 0.00864f
C840 B.n800 VSUBS 0.00864f
C841 B.n801 VSUBS 0.00864f
C842 B.n802 VSUBS 0.00864f
C843 B.n803 VSUBS 0.00864f
C844 B.n804 VSUBS 0.00864f
C845 B.n805 VSUBS 0.00864f
C846 B.n806 VSUBS 0.00864f
C847 B.n807 VSUBS 0.00864f
C848 B.n808 VSUBS 0.00864f
C849 B.n809 VSUBS 0.00864f
C850 B.n810 VSUBS 0.00864f
C851 B.n811 VSUBS 0.00864f
C852 B.n812 VSUBS 0.00864f
C853 B.n813 VSUBS 0.00864f
C854 B.n814 VSUBS 0.00864f
C855 B.n815 VSUBS 0.00864f
C856 B.n816 VSUBS 0.005972f
C857 B.n817 VSUBS 0.020018f
C858 B.n818 VSUBS 0.006988f
C859 B.n819 VSUBS 0.00864f
C860 B.n820 VSUBS 0.00864f
C861 B.n821 VSUBS 0.00864f
C862 B.n822 VSUBS 0.00864f
C863 B.n823 VSUBS 0.00864f
C864 B.n824 VSUBS 0.00864f
C865 B.n825 VSUBS 0.00864f
C866 B.n826 VSUBS 0.00864f
C867 B.n827 VSUBS 0.00864f
C868 B.n828 VSUBS 0.00864f
C869 B.n829 VSUBS 0.00864f
C870 B.n830 VSUBS 0.006988f
C871 B.n831 VSUBS 0.00864f
C872 B.n832 VSUBS 0.00864f
C873 B.n833 VSUBS 0.005972f
C874 B.n834 VSUBS 0.00864f
C875 B.n835 VSUBS 0.00864f
C876 B.n836 VSUBS 0.00864f
C877 B.n837 VSUBS 0.00864f
C878 B.n838 VSUBS 0.00864f
C879 B.n839 VSUBS 0.00864f
C880 B.n840 VSUBS 0.00864f
C881 B.n841 VSUBS 0.00864f
C882 B.n842 VSUBS 0.00864f
C883 B.n843 VSUBS 0.00864f
C884 B.n844 VSUBS 0.00864f
C885 B.n845 VSUBS 0.00864f
C886 B.n846 VSUBS 0.00864f
C887 B.n847 VSUBS 0.00864f
C888 B.n848 VSUBS 0.00864f
C889 B.n849 VSUBS 0.00864f
C890 B.n850 VSUBS 0.00864f
C891 B.n851 VSUBS 0.00864f
C892 B.n852 VSUBS 0.00864f
C893 B.n853 VSUBS 0.00864f
C894 B.n854 VSUBS 0.00864f
C895 B.n855 VSUBS 0.00864f
C896 B.n856 VSUBS 0.00864f
C897 B.n857 VSUBS 0.00864f
C898 B.n858 VSUBS 0.00864f
C899 B.n859 VSUBS 0.00864f
C900 B.n860 VSUBS 0.00864f
C901 B.n861 VSUBS 0.00864f
C902 B.n862 VSUBS 0.00864f
C903 B.n863 VSUBS 0.00864f
C904 B.n864 VSUBS 0.00864f
C905 B.n865 VSUBS 0.00864f
C906 B.n866 VSUBS 0.00864f
C907 B.n867 VSUBS 0.00864f
C908 B.n868 VSUBS 0.00864f
C909 B.n869 VSUBS 0.00864f
C910 B.n870 VSUBS 0.00864f
C911 B.n871 VSUBS 0.00864f
C912 B.n872 VSUBS 0.00864f
C913 B.n873 VSUBS 0.00864f
C914 B.n874 VSUBS 0.00864f
C915 B.n875 VSUBS 0.00864f
C916 B.n876 VSUBS 0.00864f
C917 B.n877 VSUBS 0.00864f
C918 B.n878 VSUBS 0.00864f
C919 B.n879 VSUBS 0.00864f
C920 B.n880 VSUBS 0.00864f
C921 B.n881 VSUBS 0.00864f
C922 B.n882 VSUBS 0.00864f
C923 B.n883 VSUBS 0.00864f
C924 B.n884 VSUBS 0.00864f
C925 B.n885 VSUBS 0.00864f
C926 B.n886 VSUBS 0.00864f
C927 B.n887 VSUBS 0.00864f
C928 B.n888 VSUBS 0.00864f
C929 B.n889 VSUBS 0.00864f
C930 B.n890 VSUBS 0.00864f
C931 B.n891 VSUBS 0.00864f
C932 B.n892 VSUBS 0.00864f
C933 B.n893 VSUBS 0.00864f
C934 B.n894 VSUBS 0.00864f
C935 B.n895 VSUBS 0.00864f
C936 B.n896 VSUBS 0.00864f
C937 B.n897 VSUBS 0.00864f
C938 B.n898 VSUBS 0.019824f
C939 B.n899 VSUBS 0.019824f
C940 B.n900 VSUBS 0.019057f
C941 B.n901 VSUBS 0.00864f
C942 B.n902 VSUBS 0.00864f
C943 B.n903 VSUBS 0.00864f
C944 B.n904 VSUBS 0.00864f
C945 B.n905 VSUBS 0.00864f
C946 B.n906 VSUBS 0.00864f
C947 B.n907 VSUBS 0.00864f
C948 B.n908 VSUBS 0.00864f
C949 B.n909 VSUBS 0.00864f
C950 B.n910 VSUBS 0.00864f
C951 B.n911 VSUBS 0.00864f
C952 B.n912 VSUBS 0.00864f
C953 B.n913 VSUBS 0.00864f
C954 B.n914 VSUBS 0.00864f
C955 B.n915 VSUBS 0.00864f
C956 B.n916 VSUBS 0.00864f
C957 B.n917 VSUBS 0.00864f
C958 B.n918 VSUBS 0.00864f
C959 B.n919 VSUBS 0.00864f
C960 B.n920 VSUBS 0.00864f
C961 B.n921 VSUBS 0.00864f
C962 B.n922 VSUBS 0.00864f
C963 B.n923 VSUBS 0.00864f
C964 B.n924 VSUBS 0.00864f
C965 B.n925 VSUBS 0.00864f
C966 B.n926 VSUBS 0.00864f
C967 B.n927 VSUBS 0.00864f
C968 B.n928 VSUBS 0.00864f
C969 B.n929 VSUBS 0.00864f
C970 B.n930 VSUBS 0.00864f
C971 B.n931 VSUBS 0.00864f
C972 B.n932 VSUBS 0.00864f
C973 B.n933 VSUBS 0.00864f
C974 B.n934 VSUBS 0.00864f
C975 B.n935 VSUBS 0.00864f
C976 B.n936 VSUBS 0.00864f
C977 B.n937 VSUBS 0.00864f
C978 B.n938 VSUBS 0.00864f
C979 B.n939 VSUBS 0.00864f
C980 B.n940 VSUBS 0.00864f
C981 B.n941 VSUBS 0.00864f
C982 B.n942 VSUBS 0.00864f
C983 B.n943 VSUBS 0.00864f
C984 B.n944 VSUBS 0.00864f
C985 B.n945 VSUBS 0.00864f
C986 B.n946 VSUBS 0.00864f
C987 B.n947 VSUBS 0.00864f
C988 B.n948 VSUBS 0.00864f
C989 B.n949 VSUBS 0.00864f
C990 B.n950 VSUBS 0.00864f
C991 B.n951 VSUBS 0.00864f
C992 B.n952 VSUBS 0.00864f
C993 B.n953 VSUBS 0.00864f
C994 B.n954 VSUBS 0.00864f
C995 B.n955 VSUBS 0.00864f
C996 B.n956 VSUBS 0.00864f
C997 B.n957 VSUBS 0.00864f
C998 B.n958 VSUBS 0.00864f
C999 B.n959 VSUBS 0.00864f
C1000 B.n960 VSUBS 0.00864f
C1001 B.n961 VSUBS 0.00864f
C1002 B.n962 VSUBS 0.00864f
C1003 B.n963 VSUBS 0.00864f
C1004 B.n964 VSUBS 0.00864f
C1005 B.n965 VSUBS 0.00864f
C1006 B.n966 VSUBS 0.00864f
C1007 B.n967 VSUBS 0.00864f
C1008 B.n968 VSUBS 0.00864f
C1009 B.n969 VSUBS 0.00864f
C1010 B.n970 VSUBS 0.00864f
C1011 B.n971 VSUBS 0.00864f
C1012 B.n972 VSUBS 0.00864f
C1013 B.n973 VSUBS 0.00864f
C1014 B.n974 VSUBS 0.00864f
C1015 B.n975 VSUBS 0.00864f
C1016 B.n976 VSUBS 0.00864f
C1017 B.n977 VSUBS 0.00864f
C1018 B.n978 VSUBS 0.00864f
C1019 B.n979 VSUBS 0.00864f
C1020 B.n980 VSUBS 0.00864f
C1021 B.n981 VSUBS 0.00864f
C1022 B.n982 VSUBS 0.00864f
C1023 B.n983 VSUBS 0.00864f
C1024 B.n984 VSUBS 0.00864f
C1025 B.n985 VSUBS 0.00864f
C1026 B.n986 VSUBS 0.00864f
C1027 B.n987 VSUBS 0.00864f
C1028 B.n988 VSUBS 0.00864f
C1029 B.n989 VSUBS 0.00864f
C1030 B.n990 VSUBS 0.00864f
C1031 B.n991 VSUBS 0.00864f
C1032 B.n992 VSUBS 0.00864f
C1033 B.n993 VSUBS 0.00864f
C1034 B.n994 VSUBS 0.00864f
C1035 B.n995 VSUBS 0.00864f
C1036 B.n996 VSUBS 0.00864f
C1037 B.n997 VSUBS 0.00864f
C1038 B.n998 VSUBS 0.00864f
C1039 B.n999 VSUBS 0.00864f
C1040 B.n1000 VSUBS 0.00864f
C1041 B.n1001 VSUBS 0.00864f
C1042 B.n1002 VSUBS 0.00864f
C1043 B.n1003 VSUBS 0.00864f
C1044 B.n1004 VSUBS 0.00864f
C1045 B.n1005 VSUBS 0.00864f
C1046 B.n1006 VSUBS 0.00864f
C1047 B.n1007 VSUBS 0.00864f
C1048 B.n1008 VSUBS 0.00864f
C1049 B.n1009 VSUBS 0.00864f
C1050 B.n1010 VSUBS 0.00864f
C1051 B.n1011 VSUBS 0.011275f
C1052 B.n1012 VSUBS 0.012011f
C1053 B.n1013 VSUBS 0.023885f
C1054 VDD1.t5 VSUBS 3.3118f
C1055 VDD1.t9 VSUBS 0.313921f
C1056 VDD1.t0 VSUBS 0.313921f
C1057 VDD1.n0 VSUBS 2.51285f
C1058 VDD1.n1 VSUBS 1.90327f
C1059 VDD1.t2 VSUBS 3.31178f
C1060 VDD1.t1 VSUBS 0.313921f
C1061 VDD1.t7 VSUBS 0.313921f
C1062 VDD1.n2 VSUBS 2.51283f
C1063 VDD1.n3 VSUBS 1.89309f
C1064 VDD1.t8 VSUBS 0.313921f
C1065 VDD1.t4 VSUBS 0.313921f
C1066 VDD1.n4 VSUBS 2.54714f
C1067 VDD1.n5 VSUBS 4.65503f
C1068 VDD1.t3 VSUBS 0.313921f
C1069 VDD1.t6 VSUBS 0.313921f
C1070 VDD1.n6 VSUBS 2.51283f
C1071 VDD1.n7 VSUBS 4.70584f
C1072 VP.t5 VSUBS 3.17128f
C1073 VP.n0 VSUBS 1.20057f
C1074 VP.n1 VSUBS 0.025571f
C1075 VP.n2 VSUBS 0.039825f
C1076 VP.n3 VSUBS 0.025571f
C1077 VP.n4 VSUBS 0.033069f
C1078 VP.n5 VSUBS 0.025571f
C1079 VP.n6 VSUBS 0.023799f
C1080 VP.n7 VSUBS 0.025571f
C1081 VP.t2 VSUBS 3.17128f
C1082 VP.n8 VSUBS 1.13246f
C1083 VP.n9 VSUBS 0.025571f
C1084 VP.n10 VSUBS 0.023799f
C1085 VP.n11 VSUBS 0.025571f
C1086 VP.t8 VSUBS 3.17128f
C1087 VP.n12 VSUBS 1.10833f
C1088 VP.n13 VSUBS 0.025571f
C1089 VP.n14 VSUBS 0.034837f
C1090 VP.n15 VSUBS 0.025571f
C1091 VP.n16 VSUBS 0.029775f
C1092 VP.t3 VSUBS 3.17128f
C1093 VP.n17 VSUBS 1.20057f
C1094 VP.n18 VSUBS 0.025571f
C1095 VP.n19 VSUBS 0.039825f
C1096 VP.n20 VSUBS 0.025571f
C1097 VP.n21 VSUBS 0.033069f
C1098 VP.n22 VSUBS 0.025571f
C1099 VP.n23 VSUBS 0.023799f
C1100 VP.n24 VSUBS 0.025571f
C1101 VP.t9 VSUBS 3.17128f
C1102 VP.n25 VSUBS 1.13246f
C1103 VP.n26 VSUBS 0.025571f
C1104 VP.n27 VSUBS 0.023799f
C1105 VP.n28 VSUBS 0.025571f
C1106 VP.t0 VSUBS 3.17128f
C1107 VP.n29 VSUBS 1.19875f
C1108 VP.t4 VSUBS 3.51542f
C1109 VP.n30 VSUBS 1.14303f
C1110 VP.n31 VSUBS 0.316863f
C1111 VP.n32 VSUBS 0.038716f
C1112 VP.n33 VSUBS 0.047657f
C1113 VP.n34 VSUBS 0.051341f
C1114 VP.n35 VSUBS 0.025571f
C1115 VP.n36 VSUBS 0.025571f
C1116 VP.n37 VSUBS 0.025571f
C1117 VP.n38 VSUBS 0.047179f
C1118 VP.n39 VSUBS 0.047657f
C1119 VP.n40 VSUBS 0.047657f
C1120 VP.n41 VSUBS 0.025571f
C1121 VP.n42 VSUBS 0.025571f
C1122 VP.n43 VSUBS 0.025571f
C1123 VP.n44 VSUBS 0.047657f
C1124 VP.n45 VSUBS 0.047657f
C1125 VP.n46 VSUBS 0.047179f
C1126 VP.n47 VSUBS 0.025571f
C1127 VP.n48 VSUBS 0.025571f
C1128 VP.n49 VSUBS 0.025571f
C1129 VP.n50 VSUBS 0.051341f
C1130 VP.n51 VSUBS 0.047657f
C1131 VP.t6 VSUBS 3.17128f
C1132 VP.n52 VSUBS 1.10833f
C1133 VP.n53 VSUBS 0.038716f
C1134 VP.n54 VSUBS 0.025571f
C1135 VP.n55 VSUBS 0.025571f
C1136 VP.n56 VSUBS 0.025571f
C1137 VP.n57 VSUBS 0.047657f
C1138 VP.n58 VSUBS 0.047657f
C1139 VP.n59 VSUBS 0.034837f
C1140 VP.n60 VSUBS 0.025571f
C1141 VP.n61 VSUBS 0.025571f
C1142 VP.n62 VSUBS 0.025571f
C1143 VP.n63 VSUBS 0.047657f
C1144 VP.n64 VSUBS 0.047657f
C1145 VP.n65 VSUBS 0.029775f
C1146 VP.n66 VSUBS 0.04127f
C1147 VP.n67 VSUBS 1.82725f
C1148 VP.t7 VSUBS 3.17128f
C1149 VP.n68 VSUBS 1.20057f
C1150 VP.n69 VSUBS 1.8429f
C1151 VP.n70 VSUBS 0.04127f
C1152 VP.n71 VSUBS 0.025571f
C1153 VP.n72 VSUBS 0.047657f
C1154 VP.n73 VSUBS 0.047657f
C1155 VP.n74 VSUBS 0.039825f
C1156 VP.n75 VSUBS 0.025571f
C1157 VP.n76 VSUBS 0.025571f
C1158 VP.n77 VSUBS 0.025571f
C1159 VP.n78 VSUBS 0.047657f
C1160 VP.n79 VSUBS 0.047657f
C1161 VP.n80 VSUBS 0.033069f
C1162 VP.n81 VSUBS 0.025571f
C1163 VP.n82 VSUBS 0.025571f
C1164 VP.n83 VSUBS 0.038716f
C1165 VP.n84 VSUBS 0.047657f
C1166 VP.n85 VSUBS 0.051341f
C1167 VP.n86 VSUBS 0.025571f
C1168 VP.n87 VSUBS 0.025571f
C1169 VP.n88 VSUBS 0.025571f
C1170 VP.n89 VSUBS 0.047179f
C1171 VP.n90 VSUBS 0.047657f
C1172 VP.n91 VSUBS 0.047657f
C1173 VP.n92 VSUBS 0.025571f
C1174 VP.n93 VSUBS 0.025571f
C1175 VP.n94 VSUBS 0.025571f
C1176 VP.n95 VSUBS 0.047657f
C1177 VP.n96 VSUBS 0.047657f
C1178 VP.n97 VSUBS 0.047179f
C1179 VP.n98 VSUBS 0.025571f
C1180 VP.n99 VSUBS 0.025571f
C1181 VP.n100 VSUBS 0.025571f
C1182 VP.n101 VSUBS 0.051341f
C1183 VP.n102 VSUBS 0.047657f
C1184 VP.t1 VSUBS 3.17128f
C1185 VP.n103 VSUBS 1.10833f
C1186 VP.n104 VSUBS 0.038716f
C1187 VP.n105 VSUBS 0.025571f
C1188 VP.n106 VSUBS 0.025571f
C1189 VP.n107 VSUBS 0.025571f
C1190 VP.n108 VSUBS 0.047657f
C1191 VP.n109 VSUBS 0.047657f
C1192 VP.n110 VSUBS 0.034837f
C1193 VP.n111 VSUBS 0.025571f
C1194 VP.n112 VSUBS 0.025571f
C1195 VP.n113 VSUBS 0.025571f
C1196 VP.n114 VSUBS 0.047657f
C1197 VP.n115 VSUBS 0.047657f
C1198 VP.n116 VSUBS 0.029775f
C1199 VP.n117 VSUBS 0.04127f
C1200 VP.n118 VSUBS 0.071862f
C1201 VDD2.t3 VSUBS 3.32321f
C1202 VDD2.t1 VSUBS 0.315004f
C1203 VDD2.t7 VSUBS 0.315004f
C1204 VDD2.n0 VSUBS 2.5215f
C1205 VDD2.n1 VSUBS 1.89962f
C1206 VDD2.t2 VSUBS 0.315004f
C1207 VDD2.t9 VSUBS 0.315004f
C1208 VDD2.n2 VSUBS 2.55593f
C1209 VDD2.n3 VSUBS 4.48781f
C1210 VDD2.t4 VSUBS 3.28381f
C1211 VDD2.n4 VSUBS 4.6526f
C1212 VDD2.t0 VSUBS 0.315004f
C1213 VDD2.t8 VSUBS 0.315004f
C1214 VDD2.n5 VSUBS 2.52152f
C1215 VDD2.n6 VSUBS 0.963344f
C1216 VDD2.t5 VSUBS 0.315004f
C1217 VDD2.t6 VSUBS 0.315004f
C1218 VDD2.n7 VSUBS 2.55587f
C1219 VTAIL.t12 VSUBS 0.302111f
C1220 VTAIL.t14 VSUBS 0.302111f
C1221 VTAIL.n0 VSUBS 2.27155f
C1222 VTAIL.n1 VSUBS 1.07521f
C1223 VTAIL.t6 VSUBS 2.98361f
C1224 VTAIL.n2 VSUBS 1.25911f
C1225 VTAIL.t9 VSUBS 0.302111f
C1226 VTAIL.t8 VSUBS 0.302111f
C1227 VTAIL.n3 VSUBS 2.27155f
C1228 VTAIL.n4 VSUBS 1.2579f
C1229 VTAIL.t0 VSUBS 0.302111f
C1230 VTAIL.t7 VSUBS 0.302111f
C1231 VTAIL.n5 VSUBS 2.27155f
C1232 VTAIL.n6 VSUBS 3.02786f
C1233 VTAIL.t15 VSUBS 0.302111f
C1234 VTAIL.t19 VSUBS 0.302111f
C1235 VTAIL.n7 VSUBS 2.27157f
C1236 VTAIL.n8 VSUBS 3.02784f
C1237 VTAIL.t13 VSUBS 0.302111f
C1238 VTAIL.t16 VSUBS 0.302111f
C1239 VTAIL.n9 VSUBS 2.27157f
C1240 VTAIL.n10 VSUBS 1.25788f
C1241 VTAIL.t17 VSUBS 2.98364f
C1242 VTAIL.n11 VSUBS 1.25908f
C1243 VTAIL.t4 VSUBS 0.302111f
C1244 VTAIL.t3 VSUBS 0.302111f
C1245 VTAIL.n12 VSUBS 2.27157f
C1246 VTAIL.n13 VSUBS 1.14721f
C1247 VTAIL.t5 VSUBS 0.302111f
C1248 VTAIL.t2 VSUBS 0.302111f
C1249 VTAIL.n14 VSUBS 2.27157f
C1250 VTAIL.n15 VSUBS 1.25788f
C1251 VTAIL.t1 VSUBS 2.98361f
C1252 VTAIL.n16 VSUBS 2.82969f
C1253 VTAIL.t11 VSUBS 2.98361f
C1254 VTAIL.n17 VSUBS 2.82969f
C1255 VTAIL.t10 VSUBS 0.302111f
C1256 VTAIL.t18 VSUBS 0.302111f
C1257 VTAIL.n18 VSUBS 2.27155f
C1258 VTAIL.n19 VSUBS 1.01987f
C1259 VN.t0 VSUBS 2.92196f
C1260 VN.n0 VSUBS 1.10618f
C1261 VN.n1 VSUBS 0.02356f
C1262 VN.n2 VSUBS 0.036694f
C1263 VN.n3 VSUBS 0.02356f
C1264 VN.n4 VSUBS 0.03047f
C1265 VN.n5 VSUBS 0.02356f
C1266 VN.n6 VSUBS 0.021928f
C1267 VN.n7 VSUBS 0.02356f
C1268 VN.t2 VSUBS 2.92196f
C1269 VN.n8 VSUBS 1.04343f
C1270 VN.n9 VSUBS 0.02356f
C1271 VN.n10 VSUBS 0.021928f
C1272 VN.n11 VSUBS 0.02356f
C1273 VN.t8 VSUBS 2.92196f
C1274 VN.n12 VSUBS 1.10451f
C1275 VN.t6 VSUBS 3.23904f
C1276 VN.n13 VSUBS 1.05317f
C1277 VN.n14 VSUBS 0.291951f
C1278 VN.n15 VSUBS 0.035673f
C1279 VN.n16 VSUBS 0.04391f
C1280 VN.n17 VSUBS 0.047305f
C1281 VN.n18 VSUBS 0.02356f
C1282 VN.n19 VSUBS 0.02356f
C1283 VN.n20 VSUBS 0.02356f
C1284 VN.n21 VSUBS 0.04347f
C1285 VN.n22 VSUBS 0.04391f
C1286 VN.n23 VSUBS 0.04391f
C1287 VN.n24 VSUBS 0.02356f
C1288 VN.n25 VSUBS 0.02356f
C1289 VN.n26 VSUBS 0.02356f
C1290 VN.n27 VSUBS 0.04391f
C1291 VN.n28 VSUBS 0.04391f
C1292 VN.n29 VSUBS 0.04347f
C1293 VN.n30 VSUBS 0.02356f
C1294 VN.n31 VSUBS 0.02356f
C1295 VN.n32 VSUBS 0.02356f
C1296 VN.n33 VSUBS 0.047305f
C1297 VN.n34 VSUBS 0.04391f
C1298 VN.t7 VSUBS 2.92196f
C1299 VN.n35 VSUBS 1.02119f
C1300 VN.n36 VSUBS 0.035673f
C1301 VN.n37 VSUBS 0.02356f
C1302 VN.n38 VSUBS 0.02356f
C1303 VN.n39 VSUBS 0.02356f
C1304 VN.n40 VSUBS 0.04391f
C1305 VN.n41 VSUBS 0.04391f
C1306 VN.n42 VSUBS 0.032098f
C1307 VN.n43 VSUBS 0.02356f
C1308 VN.n44 VSUBS 0.02356f
C1309 VN.n45 VSUBS 0.02356f
C1310 VN.n46 VSUBS 0.04391f
C1311 VN.n47 VSUBS 0.04391f
C1312 VN.n48 VSUBS 0.027434f
C1313 VN.n49 VSUBS 0.038026f
C1314 VN.n50 VSUBS 0.066212f
C1315 VN.t5 VSUBS 2.92196f
C1316 VN.n51 VSUBS 1.10618f
C1317 VN.n52 VSUBS 0.02356f
C1318 VN.n53 VSUBS 0.036694f
C1319 VN.n54 VSUBS 0.02356f
C1320 VN.n55 VSUBS 0.03047f
C1321 VN.n56 VSUBS 0.02356f
C1322 VN.t9 VSUBS 2.92196f
C1323 VN.n57 VSUBS 1.02119f
C1324 VN.n58 VSUBS 0.021928f
C1325 VN.n59 VSUBS 0.02356f
C1326 VN.t1 VSUBS 2.92196f
C1327 VN.n60 VSUBS 1.04343f
C1328 VN.n61 VSUBS 0.02356f
C1329 VN.n62 VSUBS 0.021928f
C1330 VN.n63 VSUBS 0.02356f
C1331 VN.t4 VSUBS 2.92196f
C1332 VN.n64 VSUBS 1.10451f
C1333 VN.t3 VSUBS 3.23904f
C1334 VN.n65 VSUBS 1.05317f
C1335 VN.n66 VSUBS 0.291951f
C1336 VN.n67 VSUBS 0.035673f
C1337 VN.n68 VSUBS 0.04391f
C1338 VN.n69 VSUBS 0.047305f
C1339 VN.n70 VSUBS 0.02356f
C1340 VN.n71 VSUBS 0.02356f
C1341 VN.n72 VSUBS 0.02356f
C1342 VN.n73 VSUBS 0.04347f
C1343 VN.n74 VSUBS 0.04391f
C1344 VN.n75 VSUBS 0.04391f
C1345 VN.n76 VSUBS 0.02356f
C1346 VN.n77 VSUBS 0.02356f
C1347 VN.n78 VSUBS 0.02356f
C1348 VN.n79 VSUBS 0.04391f
C1349 VN.n80 VSUBS 0.04391f
C1350 VN.n81 VSUBS 0.04347f
C1351 VN.n82 VSUBS 0.02356f
C1352 VN.n83 VSUBS 0.02356f
C1353 VN.n84 VSUBS 0.02356f
C1354 VN.n85 VSUBS 0.047305f
C1355 VN.n86 VSUBS 0.04391f
C1356 VN.n87 VSUBS 0.035673f
C1357 VN.n88 VSUBS 0.02356f
C1358 VN.n89 VSUBS 0.02356f
C1359 VN.n90 VSUBS 0.02356f
C1360 VN.n91 VSUBS 0.04391f
C1361 VN.n92 VSUBS 0.04391f
C1362 VN.n93 VSUBS 0.032098f
C1363 VN.n94 VSUBS 0.02356f
C1364 VN.n95 VSUBS 0.02356f
C1365 VN.n96 VSUBS 0.02356f
C1366 VN.n97 VSUBS 0.04391f
C1367 VN.n98 VSUBS 0.04391f
C1368 VN.n99 VSUBS 0.027434f
C1369 VN.n100 VSUBS 0.038026f
C1370 VN.n101 VSUBS 1.69274f
.ends

