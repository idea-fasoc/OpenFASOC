* NGSPICE file created from diff_pair_sample_0183.ext - technology: sky130A

.subckt diff_pair_sample_0183 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t19 B.t4 sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=3.37
X1 VTAIL.t3 VP.t0 VDD1.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X2 VDD1.t8 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=3.37
X3 VTAIL.t9 VP.t2 VDD1.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X4 VDD2.t8 VN.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=3.37
X5 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=3.37
X6 VTAIL.t5 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X7 VTAIL.t13 VN.t2 VDD2.t7 B.t9 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X8 VDD1.t5 VP.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X9 VTAIL.t11 VN.t3 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X10 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=3.37
X11 VTAIL.t12 VN.t4 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X12 VTAIL.t17 VN.t5 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X13 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=3.37
X14 VDD2.t3 VN.t6 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=3.37
X15 VTAIL.t0 VP.t5 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X16 VDD2.t2 VN.t7 VTAIL.t10 B.t2 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=3.37
X17 VDD2.t1 VN.t8 VTAIL.t16 B.t6 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X18 VDD1.t3 VP.t6 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=3.37
X19 VDD2.t0 VN.t9 VTAIL.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X20 VDD1.t2 VP.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=1.98 ps=12.33 w=12 l=3.37
X21 VDD1.t1 VP.t8 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.98 pd=12.33 as=4.68 ps=24.78 w=12 l=3.37
X22 VDD1.t0 VP.t9 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=1.98 ps=12.33 w=12 l=3.37
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.68 pd=24.78 as=0 ps=0 w=12 l=3.37
R0 VN.n98 VN.n97 161.3
R1 VN.n96 VN.n51 161.3
R2 VN.n95 VN.n94 161.3
R3 VN.n93 VN.n52 161.3
R4 VN.n92 VN.n91 161.3
R5 VN.n90 VN.n53 161.3
R6 VN.n89 VN.n88 161.3
R7 VN.n87 VN.n54 161.3
R8 VN.n86 VN.n85 161.3
R9 VN.n84 VN.n55 161.3
R10 VN.n83 VN.n82 161.3
R11 VN.n81 VN.n57 161.3
R12 VN.n80 VN.n79 161.3
R13 VN.n78 VN.n58 161.3
R14 VN.n77 VN.n76 161.3
R15 VN.n75 VN.n74 161.3
R16 VN.n73 VN.n60 161.3
R17 VN.n72 VN.n71 161.3
R18 VN.n70 VN.n61 161.3
R19 VN.n69 VN.n68 161.3
R20 VN.n67 VN.n62 161.3
R21 VN.n66 VN.n65 161.3
R22 VN.n48 VN.n47 161.3
R23 VN.n46 VN.n1 161.3
R24 VN.n45 VN.n44 161.3
R25 VN.n43 VN.n2 161.3
R26 VN.n42 VN.n41 161.3
R27 VN.n40 VN.n3 161.3
R28 VN.n39 VN.n38 161.3
R29 VN.n37 VN.n4 161.3
R30 VN.n36 VN.n35 161.3
R31 VN.n33 VN.n5 161.3
R32 VN.n32 VN.n31 161.3
R33 VN.n30 VN.n6 161.3
R34 VN.n29 VN.n28 161.3
R35 VN.n27 VN.n7 161.3
R36 VN.n26 VN.n25 161.3
R37 VN.n24 VN.n23 161.3
R38 VN.n22 VN.n9 161.3
R39 VN.n21 VN.n20 161.3
R40 VN.n19 VN.n10 161.3
R41 VN.n18 VN.n17 161.3
R42 VN.n16 VN.n11 161.3
R43 VN.n15 VN.n14 161.3
R44 VN.n64 VN.t6 118.828
R45 VN.n13 VN.t0 118.828
R46 VN.n12 VN.t4 85.8165
R47 VN.n8 VN.t8 85.8165
R48 VN.n34 VN.t2 85.8165
R49 VN.n0 VN.t7 85.8165
R50 VN.n63 VN.t5 85.8165
R51 VN.n59 VN.t9 85.8165
R52 VN.n56 VN.t3 85.8165
R53 VN.n50 VN.t1 85.8165
R54 VN.n49 VN.n0 82.868
R55 VN.n99 VN.n50 82.868
R56 VN VN.n99 57.483
R57 VN.n41 VN.n2 56.5617
R58 VN.n91 VN.n52 56.5617
R59 VN.n13 VN.n12 52.6179
R60 VN.n64 VN.n63 52.6179
R61 VN.n17 VN.n10 50.2647
R62 VN.n32 VN.n6 50.2647
R63 VN.n68 VN.n61 50.2647
R64 VN.n83 VN.n57 50.2647
R65 VN.n21 VN.n10 30.8893
R66 VN.n28 VN.n6 30.8893
R67 VN.n72 VN.n61 30.8893
R68 VN.n79 VN.n57 30.8893
R69 VN.n16 VN.n15 24.5923
R70 VN.n17 VN.n16 24.5923
R71 VN.n22 VN.n21 24.5923
R72 VN.n23 VN.n22 24.5923
R73 VN.n27 VN.n26 24.5923
R74 VN.n28 VN.n27 24.5923
R75 VN.n33 VN.n32 24.5923
R76 VN.n35 VN.n33 24.5923
R77 VN.n39 VN.n4 24.5923
R78 VN.n40 VN.n39 24.5923
R79 VN.n41 VN.n40 24.5923
R80 VN.n45 VN.n2 24.5923
R81 VN.n46 VN.n45 24.5923
R82 VN.n47 VN.n46 24.5923
R83 VN.n68 VN.n67 24.5923
R84 VN.n67 VN.n66 24.5923
R85 VN.n79 VN.n78 24.5923
R86 VN.n78 VN.n77 24.5923
R87 VN.n74 VN.n73 24.5923
R88 VN.n73 VN.n72 24.5923
R89 VN.n91 VN.n90 24.5923
R90 VN.n90 VN.n89 24.5923
R91 VN.n89 VN.n54 24.5923
R92 VN.n85 VN.n84 24.5923
R93 VN.n84 VN.n83 24.5923
R94 VN.n97 VN.n96 24.5923
R95 VN.n96 VN.n95 24.5923
R96 VN.n95 VN.n52 24.5923
R97 VN.n15 VN.n12 22.1332
R98 VN.n35 VN.n34 22.1332
R99 VN.n66 VN.n63 22.1332
R100 VN.n85 VN.n56 22.1332
R101 VN.n23 VN.n8 12.2964
R102 VN.n26 VN.n8 12.2964
R103 VN.n77 VN.n59 12.2964
R104 VN.n74 VN.n59 12.2964
R105 VN.n47 VN.n0 7.37805
R106 VN.n97 VN.n50 7.37805
R107 VN.n65 VN.n64 3.23081
R108 VN.n14 VN.n13 3.23081
R109 VN.n34 VN.n4 2.45968
R110 VN.n56 VN.n54 2.45968
R111 VN.n99 VN.n98 0.354861
R112 VN.n49 VN.n48 0.354861
R113 VN VN.n49 0.267071
R114 VN.n98 VN.n51 0.189894
R115 VN.n94 VN.n51 0.189894
R116 VN.n94 VN.n93 0.189894
R117 VN.n93 VN.n92 0.189894
R118 VN.n92 VN.n53 0.189894
R119 VN.n88 VN.n53 0.189894
R120 VN.n88 VN.n87 0.189894
R121 VN.n87 VN.n86 0.189894
R122 VN.n86 VN.n55 0.189894
R123 VN.n82 VN.n55 0.189894
R124 VN.n82 VN.n81 0.189894
R125 VN.n81 VN.n80 0.189894
R126 VN.n80 VN.n58 0.189894
R127 VN.n76 VN.n58 0.189894
R128 VN.n76 VN.n75 0.189894
R129 VN.n75 VN.n60 0.189894
R130 VN.n71 VN.n60 0.189894
R131 VN.n71 VN.n70 0.189894
R132 VN.n70 VN.n69 0.189894
R133 VN.n69 VN.n62 0.189894
R134 VN.n65 VN.n62 0.189894
R135 VN.n14 VN.n11 0.189894
R136 VN.n18 VN.n11 0.189894
R137 VN.n19 VN.n18 0.189894
R138 VN.n20 VN.n19 0.189894
R139 VN.n20 VN.n9 0.189894
R140 VN.n24 VN.n9 0.189894
R141 VN.n25 VN.n24 0.189894
R142 VN.n25 VN.n7 0.189894
R143 VN.n29 VN.n7 0.189894
R144 VN.n30 VN.n29 0.189894
R145 VN.n31 VN.n30 0.189894
R146 VN.n31 VN.n5 0.189894
R147 VN.n36 VN.n5 0.189894
R148 VN.n37 VN.n36 0.189894
R149 VN.n38 VN.n37 0.189894
R150 VN.n38 VN.n3 0.189894
R151 VN.n42 VN.n3 0.189894
R152 VN.n43 VN.n42 0.189894
R153 VN.n44 VN.n43 0.189894
R154 VN.n44 VN.n1 0.189894
R155 VN.n48 VN.n1 0.189894
R156 VTAIL.n272 VTAIL.n212 289.615
R157 VTAIL.n62 VTAIL.n2 289.615
R158 VTAIL.n206 VTAIL.n146 289.615
R159 VTAIL.n136 VTAIL.n76 289.615
R160 VTAIL.n232 VTAIL.n231 185
R161 VTAIL.n237 VTAIL.n236 185
R162 VTAIL.n239 VTAIL.n238 185
R163 VTAIL.n228 VTAIL.n227 185
R164 VTAIL.n245 VTAIL.n244 185
R165 VTAIL.n247 VTAIL.n246 185
R166 VTAIL.n224 VTAIL.n223 185
R167 VTAIL.n254 VTAIL.n253 185
R168 VTAIL.n255 VTAIL.n222 185
R169 VTAIL.n257 VTAIL.n256 185
R170 VTAIL.n220 VTAIL.n219 185
R171 VTAIL.n263 VTAIL.n262 185
R172 VTAIL.n265 VTAIL.n264 185
R173 VTAIL.n216 VTAIL.n215 185
R174 VTAIL.n271 VTAIL.n270 185
R175 VTAIL.n273 VTAIL.n272 185
R176 VTAIL.n22 VTAIL.n21 185
R177 VTAIL.n27 VTAIL.n26 185
R178 VTAIL.n29 VTAIL.n28 185
R179 VTAIL.n18 VTAIL.n17 185
R180 VTAIL.n35 VTAIL.n34 185
R181 VTAIL.n37 VTAIL.n36 185
R182 VTAIL.n14 VTAIL.n13 185
R183 VTAIL.n44 VTAIL.n43 185
R184 VTAIL.n45 VTAIL.n12 185
R185 VTAIL.n47 VTAIL.n46 185
R186 VTAIL.n10 VTAIL.n9 185
R187 VTAIL.n53 VTAIL.n52 185
R188 VTAIL.n55 VTAIL.n54 185
R189 VTAIL.n6 VTAIL.n5 185
R190 VTAIL.n61 VTAIL.n60 185
R191 VTAIL.n63 VTAIL.n62 185
R192 VTAIL.n207 VTAIL.n206 185
R193 VTAIL.n205 VTAIL.n204 185
R194 VTAIL.n150 VTAIL.n149 185
R195 VTAIL.n199 VTAIL.n198 185
R196 VTAIL.n197 VTAIL.n196 185
R197 VTAIL.n154 VTAIL.n153 185
R198 VTAIL.n191 VTAIL.n190 185
R199 VTAIL.n189 VTAIL.n156 185
R200 VTAIL.n188 VTAIL.n187 185
R201 VTAIL.n159 VTAIL.n157 185
R202 VTAIL.n182 VTAIL.n181 185
R203 VTAIL.n180 VTAIL.n179 185
R204 VTAIL.n163 VTAIL.n162 185
R205 VTAIL.n174 VTAIL.n173 185
R206 VTAIL.n172 VTAIL.n171 185
R207 VTAIL.n167 VTAIL.n166 185
R208 VTAIL.n137 VTAIL.n136 185
R209 VTAIL.n135 VTAIL.n134 185
R210 VTAIL.n80 VTAIL.n79 185
R211 VTAIL.n129 VTAIL.n128 185
R212 VTAIL.n127 VTAIL.n126 185
R213 VTAIL.n84 VTAIL.n83 185
R214 VTAIL.n121 VTAIL.n120 185
R215 VTAIL.n119 VTAIL.n86 185
R216 VTAIL.n118 VTAIL.n117 185
R217 VTAIL.n89 VTAIL.n87 185
R218 VTAIL.n112 VTAIL.n111 185
R219 VTAIL.n110 VTAIL.n109 185
R220 VTAIL.n93 VTAIL.n92 185
R221 VTAIL.n104 VTAIL.n103 185
R222 VTAIL.n102 VTAIL.n101 185
R223 VTAIL.n97 VTAIL.n96 185
R224 VTAIL.n233 VTAIL.t10 149.524
R225 VTAIL.n23 VTAIL.t8 149.524
R226 VTAIL.n168 VTAIL.t2 149.524
R227 VTAIL.n98 VTAIL.t18 149.524
R228 VTAIL.n237 VTAIL.n231 104.615
R229 VTAIL.n238 VTAIL.n237 104.615
R230 VTAIL.n238 VTAIL.n227 104.615
R231 VTAIL.n245 VTAIL.n227 104.615
R232 VTAIL.n246 VTAIL.n245 104.615
R233 VTAIL.n246 VTAIL.n223 104.615
R234 VTAIL.n254 VTAIL.n223 104.615
R235 VTAIL.n255 VTAIL.n254 104.615
R236 VTAIL.n256 VTAIL.n255 104.615
R237 VTAIL.n256 VTAIL.n219 104.615
R238 VTAIL.n263 VTAIL.n219 104.615
R239 VTAIL.n264 VTAIL.n263 104.615
R240 VTAIL.n264 VTAIL.n215 104.615
R241 VTAIL.n271 VTAIL.n215 104.615
R242 VTAIL.n272 VTAIL.n271 104.615
R243 VTAIL.n27 VTAIL.n21 104.615
R244 VTAIL.n28 VTAIL.n27 104.615
R245 VTAIL.n28 VTAIL.n17 104.615
R246 VTAIL.n35 VTAIL.n17 104.615
R247 VTAIL.n36 VTAIL.n35 104.615
R248 VTAIL.n36 VTAIL.n13 104.615
R249 VTAIL.n44 VTAIL.n13 104.615
R250 VTAIL.n45 VTAIL.n44 104.615
R251 VTAIL.n46 VTAIL.n45 104.615
R252 VTAIL.n46 VTAIL.n9 104.615
R253 VTAIL.n53 VTAIL.n9 104.615
R254 VTAIL.n54 VTAIL.n53 104.615
R255 VTAIL.n54 VTAIL.n5 104.615
R256 VTAIL.n61 VTAIL.n5 104.615
R257 VTAIL.n62 VTAIL.n61 104.615
R258 VTAIL.n206 VTAIL.n205 104.615
R259 VTAIL.n205 VTAIL.n149 104.615
R260 VTAIL.n198 VTAIL.n149 104.615
R261 VTAIL.n198 VTAIL.n197 104.615
R262 VTAIL.n197 VTAIL.n153 104.615
R263 VTAIL.n190 VTAIL.n153 104.615
R264 VTAIL.n190 VTAIL.n189 104.615
R265 VTAIL.n189 VTAIL.n188 104.615
R266 VTAIL.n188 VTAIL.n157 104.615
R267 VTAIL.n181 VTAIL.n157 104.615
R268 VTAIL.n181 VTAIL.n180 104.615
R269 VTAIL.n180 VTAIL.n162 104.615
R270 VTAIL.n173 VTAIL.n162 104.615
R271 VTAIL.n173 VTAIL.n172 104.615
R272 VTAIL.n172 VTAIL.n166 104.615
R273 VTAIL.n136 VTAIL.n135 104.615
R274 VTAIL.n135 VTAIL.n79 104.615
R275 VTAIL.n128 VTAIL.n79 104.615
R276 VTAIL.n128 VTAIL.n127 104.615
R277 VTAIL.n127 VTAIL.n83 104.615
R278 VTAIL.n120 VTAIL.n83 104.615
R279 VTAIL.n120 VTAIL.n119 104.615
R280 VTAIL.n119 VTAIL.n118 104.615
R281 VTAIL.n118 VTAIL.n87 104.615
R282 VTAIL.n111 VTAIL.n87 104.615
R283 VTAIL.n111 VTAIL.n110 104.615
R284 VTAIL.n110 VTAIL.n92 104.615
R285 VTAIL.n103 VTAIL.n92 104.615
R286 VTAIL.n103 VTAIL.n102 104.615
R287 VTAIL.n102 VTAIL.n96 104.615
R288 VTAIL.t10 VTAIL.n231 52.3082
R289 VTAIL.t8 VTAIL.n21 52.3082
R290 VTAIL.t2 VTAIL.n166 52.3082
R291 VTAIL.t18 VTAIL.n96 52.3082
R292 VTAIL.n145 VTAIL.n144 42.8739
R293 VTAIL.n143 VTAIL.n142 42.8739
R294 VTAIL.n75 VTAIL.n74 42.8739
R295 VTAIL.n73 VTAIL.n72 42.8739
R296 VTAIL.n279 VTAIL.n278 42.8737
R297 VTAIL.n1 VTAIL.n0 42.8737
R298 VTAIL.n69 VTAIL.n68 42.8737
R299 VTAIL.n71 VTAIL.n70 42.8737
R300 VTAIL.n277 VTAIL.n276 29.8581
R301 VTAIL.n67 VTAIL.n66 29.8581
R302 VTAIL.n211 VTAIL.n210 29.8581
R303 VTAIL.n141 VTAIL.n140 29.8581
R304 VTAIL.n73 VTAIL.n71 29.091
R305 VTAIL.n277 VTAIL.n211 25.9014
R306 VTAIL.n257 VTAIL.n222 13.1884
R307 VTAIL.n47 VTAIL.n12 13.1884
R308 VTAIL.n191 VTAIL.n156 13.1884
R309 VTAIL.n121 VTAIL.n86 13.1884
R310 VTAIL.n253 VTAIL.n252 12.8005
R311 VTAIL.n258 VTAIL.n220 12.8005
R312 VTAIL.n43 VTAIL.n42 12.8005
R313 VTAIL.n48 VTAIL.n10 12.8005
R314 VTAIL.n192 VTAIL.n154 12.8005
R315 VTAIL.n187 VTAIL.n158 12.8005
R316 VTAIL.n122 VTAIL.n84 12.8005
R317 VTAIL.n117 VTAIL.n88 12.8005
R318 VTAIL.n251 VTAIL.n224 12.0247
R319 VTAIL.n262 VTAIL.n261 12.0247
R320 VTAIL.n41 VTAIL.n14 12.0247
R321 VTAIL.n52 VTAIL.n51 12.0247
R322 VTAIL.n196 VTAIL.n195 12.0247
R323 VTAIL.n186 VTAIL.n159 12.0247
R324 VTAIL.n126 VTAIL.n125 12.0247
R325 VTAIL.n116 VTAIL.n89 12.0247
R326 VTAIL.n248 VTAIL.n247 11.249
R327 VTAIL.n265 VTAIL.n218 11.249
R328 VTAIL.n38 VTAIL.n37 11.249
R329 VTAIL.n55 VTAIL.n8 11.249
R330 VTAIL.n199 VTAIL.n152 11.249
R331 VTAIL.n183 VTAIL.n182 11.249
R332 VTAIL.n129 VTAIL.n82 11.249
R333 VTAIL.n113 VTAIL.n112 11.249
R334 VTAIL.n244 VTAIL.n226 10.4732
R335 VTAIL.n266 VTAIL.n216 10.4732
R336 VTAIL.n34 VTAIL.n16 10.4732
R337 VTAIL.n56 VTAIL.n6 10.4732
R338 VTAIL.n200 VTAIL.n150 10.4732
R339 VTAIL.n179 VTAIL.n161 10.4732
R340 VTAIL.n130 VTAIL.n80 10.4732
R341 VTAIL.n109 VTAIL.n91 10.4732
R342 VTAIL.n233 VTAIL.n232 10.2747
R343 VTAIL.n23 VTAIL.n22 10.2747
R344 VTAIL.n168 VTAIL.n167 10.2747
R345 VTAIL.n98 VTAIL.n97 10.2747
R346 VTAIL.n243 VTAIL.n228 9.69747
R347 VTAIL.n270 VTAIL.n269 9.69747
R348 VTAIL.n33 VTAIL.n18 9.69747
R349 VTAIL.n60 VTAIL.n59 9.69747
R350 VTAIL.n204 VTAIL.n203 9.69747
R351 VTAIL.n178 VTAIL.n163 9.69747
R352 VTAIL.n134 VTAIL.n133 9.69747
R353 VTAIL.n108 VTAIL.n93 9.69747
R354 VTAIL.n276 VTAIL.n275 9.45567
R355 VTAIL.n66 VTAIL.n65 9.45567
R356 VTAIL.n210 VTAIL.n209 9.45567
R357 VTAIL.n140 VTAIL.n139 9.45567
R358 VTAIL.n275 VTAIL.n274 9.3005
R359 VTAIL.n214 VTAIL.n213 9.3005
R360 VTAIL.n269 VTAIL.n268 9.3005
R361 VTAIL.n267 VTAIL.n266 9.3005
R362 VTAIL.n218 VTAIL.n217 9.3005
R363 VTAIL.n261 VTAIL.n260 9.3005
R364 VTAIL.n259 VTAIL.n258 9.3005
R365 VTAIL.n235 VTAIL.n234 9.3005
R366 VTAIL.n230 VTAIL.n229 9.3005
R367 VTAIL.n241 VTAIL.n240 9.3005
R368 VTAIL.n243 VTAIL.n242 9.3005
R369 VTAIL.n226 VTAIL.n225 9.3005
R370 VTAIL.n249 VTAIL.n248 9.3005
R371 VTAIL.n251 VTAIL.n250 9.3005
R372 VTAIL.n252 VTAIL.n221 9.3005
R373 VTAIL.n65 VTAIL.n64 9.3005
R374 VTAIL.n4 VTAIL.n3 9.3005
R375 VTAIL.n59 VTAIL.n58 9.3005
R376 VTAIL.n57 VTAIL.n56 9.3005
R377 VTAIL.n8 VTAIL.n7 9.3005
R378 VTAIL.n51 VTAIL.n50 9.3005
R379 VTAIL.n49 VTAIL.n48 9.3005
R380 VTAIL.n25 VTAIL.n24 9.3005
R381 VTAIL.n20 VTAIL.n19 9.3005
R382 VTAIL.n31 VTAIL.n30 9.3005
R383 VTAIL.n33 VTAIL.n32 9.3005
R384 VTAIL.n16 VTAIL.n15 9.3005
R385 VTAIL.n39 VTAIL.n38 9.3005
R386 VTAIL.n41 VTAIL.n40 9.3005
R387 VTAIL.n42 VTAIL.n11 9.3005
R388 VTAIL.n170 VTAIL.n169 9.3005
R389 VTAIL.n165 VTAIL.n164 9.3005
R390 VTAIL.n176 VTAIL.n175 9.3005
R391 VTAIL.n178 VTAIL.n177 9.3005
R392 VTAIL.n161 VTAIL.n160 9.3005
R393 VTAIL.n184 VTAIL.n183 9.3005
R394 VTAIL.n186 VTAIL.n185 9.3005
R395 VTAIL.n158 VTAIL.n155 9.3005
R396 VTAIL.n209 VTAIL.n208 9.3005
R397 VTAIL.n148 VTAIL.n147 9.3005
R398 VTAIL.n203 VTAIL.n202 9.3005
R399 VTAIL.n201 VTAIL.n200 9.3005
R400 VTAIL.n152 VTAIL.n151 9.3005
R401 VTAIL.n195 VTAIL.n194 9.3005
R402 VTAIL.n193 VTAIL.n192 9.3005
R403 VTAIL.n100 VTAIL.n99 9.3005
R404 VTAIL.n95 VTAIL.n94 9.3005
R405 VTAIL.n106 VTAIL.n105 9.3005
R406 VTAIL.n108 VTAIL.n107 9.3005
R407 VTAIL.n91 VTAIL.n90 9.3005
R408 VTAIL.n114 VTAIL.n113 9.3005
R409 VTAIL.n116 VTAIL.n115 9.3005
R410 VTAIL.n88 VTAIL.n85 9.3005
R411 VTAIL.n139 VTAIL.n138 9.3005
R412 VTAIL.n78 VTAIL.n77 9.3005
R413 VTAIL.n133 VTAIL.n132 9.3005
R414 VTAIL.n131 VTAIL.n130 9.3005
R415 VTAIL.n82 VTAIL.n81 9.3005
R416 VTAIL.n125 VTAIL.n124 9.3005
R417 VTAIL.n123 VTAIL.n122 9.3005
R418 VTAIL.n240 VTAIL.n239 8.92171
R419 VTAIL.n273 VTAIL.n214 8.92171
R420 VTAIL.n30 VTAIL.n29 8.92171
R421 VTAIL.n63 VTAIL.n4 8.92171
R422 VTAIL.n207 VTAIL.n148 8.92171
R423 VTAIL.n175 VTAIL.n174 8.92171
R424 VTAIL.n137 VTAIL.n78 8.92171
R425 VTAIL.n105 VTAIL.n104 8.92171
R426 VTAIL.n236 VTAIL.n230 8.14595
R427 VTAIL.n274 VTAIL.n212 8.14595
R428 VTAIL.n26 VTAIL.n20 8.14595
R429 VTAIL.n64 VTAIL.n2 8.14595
R430 VTAIL.n208 VTAIL.n146 8.14595
R431 VTAIL.n171 VTAIL.n165 8.14595
R432 VTAIL.n138 VTAIL.n76 8.14595
R433 VTAIL.n101 VTAIL.n95 8.14595
R434 VTAIL.n235 VTAIL.n232 7.3702
R435 VTAIL.n25 VTAIL.n22 7.3702
R436 VTAIL.n170 VTAIL.n167 7.3702
R437 VTAIL.n100 VTAIL.n97 7.3702
R438 VTAIL.n236 VTAIL.n235 5.81868
R439 VTAIL.n276 VTAIL.n212 5.81868
R440 VTAIL.n26 VTAIL.n25 5.81868
R441 VTAIL.n66 VTAIL.n2 5.81868
R442 VTAIL.n210 VTAIL.n146 5.81868
R443 VTAIL.n171 VTAIL.n170 5.81868
R444 VTAIL.n140 VTAIL.n76 5.81868
R445 VTAIL.n101 VTAIL.n100 5.81868
R446 VTAIL.n239 VTAIL.n230 5.04292
R447 VTAIL.n274 VTAIL.n273 5.04292
R448 VTAIL.n29 VTAIL.n20 5.04292
R449 VTAIL.n64 VTAIL.n63 5.04292
R450 VTAIL.n208 VTAIL.n207 5.04292
R451 VTAIL.n174 VTAIL.n165 5.04292
R452 VTAIL.n138 VTAIL.n137 5.04292
R453 VTAIL.n104 VTAIL.n95 5.04292
R454 VTAIL.n240 VTAIL.n228 4.26717
R455 VTAIL.n270 VTAIL.n214 4.26717
R456 VTAIL.n30 VTAIL.n18 4.26717
R457 VTAIL.n60 VTAIL.n4 4.26717
R458 VTAIL.n204 VTAIL.n148 4.26717
R459 VTAIL.n175 VTAIL.n163 4.26717
R460 VTAIL.n134 VTAIL.n78 4.26717
R461 VTAIL.n105 VTAIL.n93 4.26717
R462 VTAIL.n244 VTAIL.n243 3.49141
R463 VTAIL.n269 VTAIL.n216 3.49141
R464 VTAIL.n34 VTAIL.n33 3.49141
R465 VTAIL.n59 VTAIL.n6 3.49141
R466 VTAIL.n203 VTAIL.n150 3.49141
R467 VTAIL.n179 VTAIL.n178 3.49141
R468 VTAIL.n133 VTAIL.n80 3.49141
R469 VTAIL.n109 VTAIL.n108 3.49141
R470 VTAIL.n75 VTAIL.n73 3.19016
R471 VTAIL.n141 VTAIL.n75 3.19016
R472 VTAIL.n145 VTAIL.n143 3.19016
R473 VTAIL.n211 VTAIL.n145 3.19016
R474 VTAIL.n71 VTAIL.n69 3.19016
R475 VTAIL.n69 VTAIL.n67 3.19016
R476 VTAIL.n279 VTAIL.n277 3.19016
R477 VTAIL.n234 VTAIL.n233 2.84303
R478 VTAIL.n24 VTAIL.n23 2.84303
R479 VTAIL.n169 VTAIL.n168 2.84303
R480 VTAIL.n99 VTAIL.n98 2.84303
R481 VTAIL.n247 VTAIL.n226 2.71565
R482 VTAIL.n266 VTAIL.n265 2.71565
R483 VTAIL.n37 VTAIL.n16 2.71565
R484 VTAIL.n56 VTAIL.n55 2.71565
R485 VTAIL.n200 VTAIL.n199 2.71565
R486 VTAIL.n182 VTAIL.n161 2.71565
R487 VTAIL.n130 VTAIL.n129 2.71565
R488 VTAIL.n112 VTAIL.n91 2.71565
R489 VTAIL VTAIL.n1 2.45093
R490 VTAIL.n143 VTAIL.n141 2.06516
R491 VTAIL.n67 VTAIL.n1 2.06516
R492 VTAIL.n248 VTAIL.n224 1.93989
R493 VTAIL.n262 VTAIL.n218 1.93989
R494 VTAIL.n38 VTAIL.n14 1.93989
R495 VTAIL.n52 VTAIL.n8 1.93989
R496 VTAIL.n196 VTAIL.n152 1.93989
R497 VTAIL.n183 VTAIL.n159 1.93989
R498 VTAIL.n126 VTAIL.n82 1.93989
R499 VTAIL.n113 VTAIL.n89 1.93989
R500 VTAIL.n278 VTAIL.t16 1.6505
R501 VTAIL.n278 VTAIL.t13 1.6505
R502 VTAIL.n0 VTAIL.t19 1.6505
R503 VTAIL.n0 VTAIL.t12 1.6505
R504 VTAIL.n68 VTAIL.t7 1.6505
R505 VTAIL.n68 VTAIL.t5 1.6505
R506 VTAIL.n70 VTAIL.t1 1.6505
R507 VTAIL.n70 VTAIL.t3 1.6505
R508 VTAIL.n144 VTAIL.t6 1.6505
R509 VTAIL.n144 VTAIL.t9 1.6505
R510 VTAIL.n142 VTAIL.t4 1.6505
R511 VTAIL.n142 VTAIL.t0 1.6505
R512 VTAIL.n74 VTAIL.t15 1.6505
R513 VTAIL.n74 VTAIL.t17 1.6505
R514 VTAIL.n72 VTAIL.t14 1.6505
R515 VTAIL.n72 VTAIL.t11 1.6505
R516 VTAIL.n253 VTAIL.n251 1.16414
R517 VTAIL.n261 VTAIL.n220 1.16414
R518 VTAIL.n43 VTAIL.n41 1.16414
R519 VTAIL.n51 VTAIL.n10 1.16414
R520 VTAIL.n195 VTAIL.n154 1.16414
R521 VTAIL.n187 VTAIL.n186 1.16414
R522 VTAIL.n125 VTAIL.n84 1.16414
R523 VTAIL.n117 VTAIL.n116 1.16414
R524 VTAIL VTAIL.n279 0.739724
R525 VTAIL.n252 VTAIL.n222 0.388379
R526 VTAIL.n258 VTAIL.n257 0.388379
R527 VTAIL.n42 VTAIL.n12 0.388379
R528 VTAIL.n48 VTAIL.n47 0.388379
R529 VTAIL.n192 VTAIL.n191 0.388379
R530 VTAIL.n158 VTAIL.n156 0.388379
R531 VTAIL.n122 VTAIL.n121 0.388379
R532 VTAIL.n88 VTAIL.n86 0.388379
R533 VTAIL.n234 VTAIL.n229 0.155672
R534 VTAIL.n241 VTAIL.n229 0.155672
R535 VTAIL.n242 VTAIL.n241 0.155672
R536 VTAIL.n242 VTAIL.n225 0.155672
R537 VTAIL.n249 VTAIL.n225 0.155672
R538 VTAIL.n250 VTAIL.n249 0.155672
R539 VTAIL.n250 VTAIL.n221 0.155672
R540 VTAIL.n259 VTAIL.n221 0.155672
R541 VTAIL.n260 VTAIL.n259 0.155672
R542 VTAIL.n260 VTAIL.n217 0.155672
R543 VTAIL.n267 VTAIL.n217 0.155672
R544 VTAIL.n268 VTAIL.n267 0.155672
R545 VTAIL.n268 VTAIL.n213 0.155672
R546 VTAIL.n275 VTAIL.n213 0.155672
R547 VTAIL.n24 VTAIL.n19 0.155672
R548 VTAIL.n31 VTAIL.n19 0.155672
R549 VTAIL.n32 VTAIL.n31 0.155672
R550 VTAIL.n32 VTAIL.n15 0.155672
R551 VTAIL.n39 VTAIL.n15 0.155672
R552 VTAIL.n40 VTAIL.n39 0.155672
R553 VTAIL.n40 VTAIL.n11 0.155672
R554 VTAIL.n49 VTAIL.n11 0.155672
R555 VTAIL.n50 VTAIL.n49 0.155672
R556 VTAIL.n50 VTAIL.n7 0.155672
R557 VTAIL.n57 VTAIL.n7 0.155672
R558 VTAIL.n58 VTAIL.n57 0.155672
R559 VTAIL.n58 VTAIL.n3 0.155672
R560 VTAIL.n65 VTAIL.n3 0.155672
R561 VTAIL.n209 VTAIL.n147 0.155672
R562 VTAIL.n202 VTAIL.n147 0.155672
R563 VTAIL.n202 VTAIL.n201 0.155672
R564 VTAIL.n201 VTAIL.n151 0.155672
R565 VTAIL.n194 VTAIL.n151 0.155672
R566 VTAIL.n194 VTAIL.n193 0.155672
R567 VTAIL.n193 VTAIL.n155 0.155672
R568 VTAIL.n185 VTAIL.n155 0.155672
R569 VTAIL.n185 VTAIL.n184 0.155672
R570 VTAIL.n184 VTAIL.n160 0.155672
R571 VTAIL.n177 VTAIL.n160 0.155672
R572 VTAIL.n177 VTAIL.n176 0.155672
R573 VTAIL.n176 VTAIL.n164 0.155672
R574 VTAIL.n169 VTAIL.n164 0.155672
R575 VTAIL.n139 VTAIL.n77 0.155672
R576 VTAIL.n132 VTAIL.n77 0.155672
R577 VTAIL.n132 VTAIL.n131 0.155672
R578 VTAIL.n131 VTAIL.n81 0.155672
R579 VTAIL.n124 VTAIL.n81 0.155672
R580 VTAIL.n124 VTAIL.n123 0.155672
R581 VTAIL.n123 VTAIL.n85 0.155672
R582 VTAIL.n115 VTAIL.n85 0.155672
R583 VTAIL.n115 VTAIL.n114 0.155672
R584 VTAIL.n114 VTAIL.n90 0.155672
R585 VTAIL.n107 VTAIL.n90 0.155672
R586 VTAIL.n107 VTAIL.n106 0.155672
R587 VTAIL.n106 VTAIL.n94 0.155672
R588 VTAIL.n99 VTAIL.n94 0.155672
R589 VDD2.n129 VDD2.n69 289.615
R590 VDD2.n60 VDD2.n0 289.615
R591 VDD2.n130 VDD2.n129 185
R592 VDD2.n128 VDD2.n127 185
R593 VDD2.n73 VDD2.n72 185
R594 VDD2.n122 VDD2.n121 185
R595 VDD2.n120 VDD2.n119 185
R596 VDD2.n77 VDD2.n76 185
R597 VDD2.n114 VDD2.n113 185
R598 VDD2.n112 VDD2.n79 185
R599 VDD2.n111 VDD2.n110 185
R600 VDD2.n82 VDD2.n80 185
R601 VDD2.n105 VDD2.n104 185
R602 VDD2.n103 VDD2.n102 185
R603 VDD2.n86 VDD2.n85 185
R604 VDD2.n97 VDD2.n96 185
R605 VDD2.n95 VDD2.n94 185
R606 VDD2.n90 VDD2.n89 185
R607 VDD2.n20 VDD2.n19 185
R608 VDD2.n25 VDD2.n24 185
R609 VDD2.n27 VDD2.n26 185
R610 VDD2.n16 VDD2.n15 185
R611 VDD2.n33 VDD2.n32 185
R612 VDD2.n35 VDD2.n34 185
R613 VDD2.n12 VDD2.n11 185
R614 VDD2.n42 VDD2.n41 185
R615 VDD2.n43 VDD2.n10 185
R616 VDD2.n45 VDD2.n44 185
R617 VDD2.n8 VDD2.n7 185
R618 VDD2.n51 VDD2.n50 185
R619 VDD2.n53 VDD2.n52 185
R620 VDD2.n4 VDD2.n3 185
R621 VDD2.n59 VDD2.n58 185
R622 VDD2.n61 VDD2.n60 185
R623 VDD2.n91 VDD2.t8 149.524
R624 VDD2.n21 VDD2.t9 149.524
R625 VDD2.n129 VDD2.n128 104.615
R626 VDD2.n128 VDD2.n72 104.615
R627 VDD2.n121 VDD2.n72 104.615
R628 VDD2.n121 VDD2.n120 104.615
R629 VDD2.n120 VDD2.n76 104.615
R630 VDD2.n113 VDD2.n76 104.615
R631 VDD2.n113 VDD2.n112 104.615
R632 VDD2.n112 VDD2.n111 104.615
R633 VDD2.n111 VDD2.n80 104.615
R634 VDD2.n104 VDD2.n80 104.615
R635 VDD2.n104 VDD2.n103 104.615
R636 VDD2.n103 VDD2.n85 104.615
R637 VDD2.n96 VDD2.n85 104.615
R638 VDD2.n96 VDD2.n95 104.615
R639 VDD2.n95 VDD2.n89 104.615
R640 VDD2.n25 VDD2.n19 104.615
R641 VDD2.n26 VDD2.n25 104.615
R642 VDD2.n26 VDD2.n15 104.615
R643 VDD2.n33 VDD2.n15 104.615
R644 VDD2.n34 VDD2.n33 104.615
R645 VDD2.n34 VDD2.n11 104.615
R646 VDD2.n42 VDD2.n11 104.615
R647 VDD2.n43 VDD2.n42 104.615
R648 VDD2.n44 VDD2.n43 104.615
R649 VDD2.n44 VDD2.n7 104.615
R650 VDD2.n51 VDD2.n7 104.615
R651 VDD2.n52 VDD2.n51 104.615
R652 VDD2.n52 VDD2.n3 104.615
R653 VDD2.n59 VDD2.n3 104.615
R654 VDD2.n60 VDD2.n59 104.615
R655 VDD2.n68 VDD2.n67 61.8894
R656 VDD2 VDD2.n137 61.8866
R657 VDD2.n136 VDD2.n135 59.5527
R658 VDD2.n66 VDD2.n65 59.5525
R659 VDD2.t8 VDD2.n89 52.3082
R660 VDD2.t9 VDD2.n19 52.3082
R661 VDD2.n66 VDD2.n64 49.7265
R662 VDD2.n134 VDD2.n68 49.211
R663 VDD2.n134 VDD2.n133 46.5369
R664 VDD2.n114 VDD2.n79 13.1884
R665 VDD2.n45 VDD2.n10 13.1884
R666 VDD2.n115 VDD2.n77 12.8005
R667 VDD2.n110 VDD2.n81 12.8005
R668 VDD2.n41 VDD2.n40 12.8005
R669 VDD2.n46 VDD2.n8 12.8005
R670 VDD2.n119 VDD2.n118 12.0247
R671 VDD2.n109 VDD2.n82 12.0247
R672 VDD2.n39 VDD2.n12 12.0247
R673 VDD2.n50 VDD2.n49 12.0247
R674 VDD2.n122 VDD2.n75 11.249
R675 VDD2.n106 VDD2.n105 11.249
R676 VDD2.n36 VDD2.n35 11.249
R677 VDD2.n53 VDD2.n6 11.249
R678 VDD2.n123 VDD2.n73 10.4732
R679 VDD2.n102 VDD2.n84 10.4732
R680 VDD2.n32 VDD2.n14 10.4732
R681 VDD2.n54 VDD2.n4 10.4732
R682 VDD2.n91 VDD2.n90 10.2747
R683 VDD2.n21 VDD2.n20 10.2747
R684 VDD2.n127 VDD2.n126 9.69747
R685 VDD2.n101 VDD2.n86 9.69747
R686 VDD2.n31 VDD2.n16 9.69747
R687 VDD2.n58 VDD2.n57 9.69747
R688 VDD2.n133 VDD2.n132 9.45567
R689 VDD2.n64 VDD2.n63 9.45567
R690 VDD2.n93 VDD2.n92 9.3005
R691 VDD2.n88 VDD2.n87 9.3005
R692 VDD2.n99 VDD2.n98 9.3005
R693 VDD2.n101 VDD2.n100 9.3005
R694 VDD2.n84 VDD2.n83 9.3005
R695 VDD2.n107 VDD2.n106 9.3005
R696 VDD2.n109 VDD2.n108 9.3005
R697 VDD2.n81 VDD2.n78 9.3005
R698 VDD2.n132 VDD2.n131 9.3005
R699 VDD2.n71 VDD2.n70 9.3005
R700 VDD2.n126 VDD2.n125 9.3005
R701 VDD2.n124 VDD2.n123 9.3005
R702 VDD2.n75 VDD2.n74 9.3005
R703 VDD2.n118 VDD2.n117 9.3005
R704 VDD2.n116 VDD2.n115 9.3005
R705 VDD2.n63 VDD2.n62 9.3005
R706 VDD2.n2 VDD2.n1 9.3005
R707 VDD2.n57 VDD2.n56 9.3005
R708 VDD2.n55 VDD2.n54 9.3005
R709 VDD2.n6 VDD2.n5 9.3005
R710 VDD2.n49 VDD2.n48 9.3005
R711 VDD2.n47 VDD2.n46 9.3005
R712 VDD2.n23 VDD2.n22 9.3005
R713 VDD2.n18 VDD2.n17 9.3005
R714 VDD2.n29 VDD2.n28 9.3005
R715 VDD2.n31 VDD2.n30 9.3005
R716 VDD2.n14 VDD2.n13 9.3005
R717 VDD2.n37 VDD2.n36 9.3005
R718 VDD2.n39 VDD2.n38 9.3005
R719 VDD2.n40 VDD2.n9 9.3005
R720 VDD2.n130 VDD2.n71 8.92171
R721 VDD2.n98 VDD2.n97 8.92171
R722 VDD2.n28 VDD2.n27 8.92171
R723 VDD2.n61 VDD2.n2 8.92171
R724 VDD2.n131 VDD2.n69 8.14595
R725 VDD2.n94 VDD2.n88 8.14595
R726 VDD2.n24 VDD2.n18 8.14595
R727 VDD2.n62 VDD2.n0 8.14595
R728 VDD2.n93 VDD2.n90 7.3702
R729 VDD2.n23 VDD2.n20 7.3702
R730 VDD2.n133 VDD2.n69 5.81868
R731 VDD2.n94 VDD2.n93 5.81868
R732 VDD2.n24 VDD2.n23 5.81868
R733 VDD2.n64 VDD2.n0 5.81868
R734 VDD2.n131 VDD2.n130 5.04292
R735 VDD2.n97 VDD2.n88 5.04292
R736 VDD2.n27 VDD2.n18 5.04292
R737 VDD2.n62 VDD2.n61 5.04292
R738 VDD2.n127 VDD2.n71 4.26717
R739 VDD2.n98 VDD2.n86 4.26717
R740 VDD2.n28 VDD2.n16 4.26717
R741 VDD2.n58 VDD2.n2 4.26717
R742 VDD2.n126 VDD2.n73 3.49141
R743 VDD2.n102 VDD2.n101 3.49141
R744 VDD2.n32 VDD2.n31 3.49141
R745 VDD2.n57 VDD2.n4 3.49141
R746 VDD2.n136 VDD2.n134 3.19016
R747 VDD2.n92 VDD2.n91 2.84303
R748 VDD2.n22 VDD2.n21 2.84303
R749 VDD2.n123 VDD2.n122 2.71565
R750 VDD2.n105 VDD2.n84 2.71565
R751 VDD2.n35 VDD2.n14 2.71565
R752 VDD2.n54 VDD2.n53 2.71565
R753 VDD2.n119 VDD2.n75 1.93989
R754 VDD2.n106 VDD2.n82 1.93989
R755 VDD2.n36 VDD2.n12 1.93989
R756 VDD2.n50 VDD2.n6 1.93989
R757 VDD2.n137 VDD2.t4 1.6505
R758 VDD2.n137 VDD2.t3 1.6505
R759 VDD2.n135 VDD2.t6 1.6505
R760 VDD2.n135 VDD2.t0 1.6505
R761 VDD2.n67 VDD2.t7 1.6505
R762 VDD2.n67 VDD2.t2 1.6505
R763 VDD2.n65 VDD2.t5 1.6505
R764 VDD2.n65 VDD2.t1 1.6505
R765 VDD2.n118 VDD2.n77 1.16414
R766 VDD2.n110 VDD2.n109 1.16414
R767 VDD2.n41 VDD2.n39 1.16414
R768 VDD2.n49 VDD2.n8 1.16414
R769 VDD2 VDD2.n136 0.856103
R770 VDD2.n68 VDD2.n66 0.742568
R771 VDD2.n115 VDD2.n114 0.388379
R772 VDD2.n81 VDD2.n79 0.388379
R773 VDD2.n40 VDD2.n10 0.388379
R774 VDD2.n46 VDD2.n45 0.388379
R775 VDD2.n132 VDD2.n70 0.155672
R776 VDD2.n125 VDD2.n70 0.155672
R777 VDD2.n125 VDD2.n124 0.155672
R778 VDD2.n124 VDD2.n74 0.155672
R779 VDD2.n117 VDD2.n74 0.155672
R780 VDD2.n117 VDD2.n116 0.155672
R781 VDD2.n116 VDD2.n78 0.155672
R782 VDD2.n108 VDD2.n78 0.155672
R783 VDD2.n108 VDD2.n107 0.155672
R784 VDD2.n107 VDD2.n83 0.155672
R785 VDD2.n100 VDD2.n83 0.155672
R786 VDD2.n100 VDD2.n99 0.155672
R787 VDD2.n99 VDD2.n87 0.155672
R788 VDD2.n92 VDD2.n87 0.155672
R789 VDD2.n22 VDD2.n17 0.155672
R790 VDD2.n29 VDD2.n17 0.155672
R791 VDD2.n30 VDD2.n29 0.155672
R792 VDD2.n30 VDD2.n13 0.155672
R793 VDD2.n37 VDD2.n13 0.155672
R794 VDD2.n38 VDD2.n37 0.155672
R795 VDD2.n38 VDD2.n9 0.155672
R796 VDD2.n47 VDD2.n9 0.155672
R797 VDD2.n48 VDD2.n47 0.155672
R798 VDD2.n48 VDD2.n5 0.155672
R799 VDD2.n55 VDD2.n5 0.155672
R800 VDD2.n56 VDD2.n55 0.155672
R801 VDD2.n56 VDD2.n1 0.155672
R802 VDD2.n63 VDD2.n1 0.155672
R803 B.n1066 B.n1065 585
R804 B.n1067 B.n1066 585
R805 B.n369 B.n180 585
R806 B.n368 B.n367 585
R807 B.n366 B.n365 585
R808 B.n364 B.n363 585
R809 B.n362 B.n361 585
R810 B.n360 B.n359 585
R811 B.n358 B.n357 585
R812 B.n356 B.n355 585
R813 B.n354 B.n353 585
R814 B.n352 B.n351 585
R815 B.n350 B.n349 585
R816 B.n348 B.n347 585
R817 B.n346 B.n345 585
R818 B.n344 B.n343 585
R819 B.n342 B.n341 585
R820 B.n340 B.n339 585
R821 B.n338 B.n337 585
R822 B.n336 B.n335 585
R823 B.n334 B.n333 585
R824 B.n332 B.n331 585
R825 B.n330 B.n329 585
R826 B.n328 B.n327 585
R827 B.n326 B.n325 585
R828 B.n324 B.n323 585
R829 B.n322 B.n321 585
R830 B.n320 B.n319 585
R831 B.n318 B.n317 585
R832 B.n316 B.n315 585
R833 B.n314 B.n313 585
R834 B.n312 B.n311 585
R835 B.n310 B.n309 585
R836 B.n308 B.n307 585
R837 B.n306 B.n305 585
R838 B.n304 B.n303 585
R839 B.n302 B.n301 585
R840 B.n300 B.n299 585
R841 B.n298 B.n297 585
R842 B.n296 B.n295 585
R843 B.n294 B.n293 585
R844 B.n292 B.n291 585
R845 B.n290 B.n289 585
R846 B.n287 B.n286 585
R847 B.n285 B.n284 585
R848 B.n283 B.n282 585
R849 B.n281 B.n280 585
R850 B.n279 B.n278 585
R851 B.n277 B.n276 585
R852 B.n275 B.n274 585
R853 B.n273 B.n272 585
R854 B.n271 B.n270 585
R855 B.n269 B.n268 585
R856 B.n267 B.n266 585
R857 B.n265 B.n264 585
R858 B.n263 B.n262 585
R859 B.n261 B.n260 585
R860 B.n259 B.n258 585
R861 B.n257 B.n256 585
R862 B.n255 B.n254 585
R863 B.n253 B.n252 585
R864 B.n251 B.n250 585
R865 B.n249 B.n248 585
R866 B.n247 B.n246 585
R867 B.n245 B.n244 585
R868 B.n243 B.n242 585
R869 B.n241 B.n240 585
R870 B.n239 B.n238 585
R871 B.n237 B.n236 585
R872 B.n235 B.n234 585
R873 B.n233 B.n232 585
R874 B.n231 B.n230 585
R875 B.n229 B.n228 585
R876 B.n227 B.n226 585
R877 B.n225 B.n224 585
R878 B.n223 B.n222 585
R879 B.n221 B.n220 585
R880 B.n219 B.n218 585
R881 B.n217 B.n216 585
R882 B.n215 B.n214 585
R883 B.n213 B.n212 585
R884 B.n211 B.n210 585
R885 B.n209 B.n208 585
R886 B.n207 B.n206 585
R887 B.n205 B.n204 585
R888 B.n203 B.n202 585
R889 B.n201 B.n200 585
R890 B.n199 B.n198 585
R891 B.n197 B.n196 585
R892 B.n195 B.n194 585
R893 B.n193 B.n192 585
R894 B.n191 B.n190 585
R895 B.n189 B.n188 585
R896 B.n187 B.n186 585
R897 B.n1064 B.n133 585
R898 B.n1068 B.n133 585
R899 B.n1063 B.n132 585
R900 B.n1069 B.n132 585
R901 B.n1062 B.n1061 585
R902 B.n1061 B.n128 585
R903 B.n1060 B.n127 585
R904 B.n1075 B.n127 585
R905 B.n1059 B.n126 585
R906 B.n1076 B.n126 585
R907 B.n1058 B.n125 585
R908 B.n1077 B.n125 585
R909 B.n1057 B.n1056 585
R910 B.n1056 B.n121 585
R911 B.n1055 B.n120 585
R912 B.n1083 B.n120 585
R913 B.n1054 B.n119 585
R914 B.n1084 B.n119 585
R915 B.n1053 B.n118 585
R916 B.n1085 B.n118 585
R917 B.n1052 B.n1051 585
R918 B.n1051 B.n114 585
R919 B.n1050 B.n113 585
R920 B.n1091 B.n113 585
R921 B.n1049 B.n112 585
R922 B.n1092 B.n112 585
R923 B.n1048 B.n111 585
R924 B.n1093 B.n111 585
R925 B.n1047 B.n1046 585
R926 B.n1046 B.n107 585
R927 B.n1045 B.n106 585
R928 B.n1099 B.n106 585
R929 B.n1044 B.n105 585
R930 B.n1100 B.n105 585
R931 B.n1043 B.n104 585
R932 B.n1101 B.n104 585
R933 B.n1042 B.n1041 585
R934 B.n1041 B.n100 585
R935 B.n1040 B.n99 585
R936 B.n1107 B.n99 585
R937 B.n1039 B.n98 585
R938 B.n1108 B.n98 585
R939 B.n1038 B.n97 585
R940 B.n1109 B.n97 585
R941 B.n1037 B.n1036 585
R942 B.n1036 B.n96 585
R943 B.n1035 B.n92 585
R944 B.n1115 B.n92 585
R945 B.n1034 B.n91 585
R946 B.n1116 B.n91 585
R947 B.n1033 B.n90 585
R948 B.n1117 B.n90 585
R949 B.n1032 B.n1031 585
R950 B.n1031 B.n86 585
R951 B.n1030 B.n85 585
R952 B.n1123 B.n85 585
R953 B.n1029 B.n84 585
R954 B.n1124 B.n84 585
R955 B.n1028 B.n83 585
R956 B.n1125 B.n83 585
R957 B.n1027 B.n1026 585
R958 B.n1026 B.n79 585
R959 B.n1025 B.n78 585
R960 B.n1131 B.n78 585
R961 B.n1024 B.n77 585
R962 B.n1132 B.n77 585
R963 B.n1023 B.n76 585
R964 B.n1133 B.n76 585
R965 B.n1022 B.n1021 585
R966 B.n1021 B.n72 585
R967 B.n1020 B.n71 585
R968 B.n1139 B.n71 585
R969 B.n1019 B.n70 585
R970 B.n1140 B.n70 585
R971 B.n1018 B.n69 585
R972 B.n1141 B.n69 585
R973 B.n1017 B.n1016 585
R974 B.n1016 B.n65 585
R975 B.n1015 B.n64 585
R976 B.n1147 B.n64 585
R977 B.n1014 B.n63 585
R978 B.n1148 B.n63 585
R979 B.n1013 B.n62 585
R980 B.n1149 B.n62 585
R981 B.n1012 B.n1011 585
R982 B.n1011 B.n58 585
R983 B.n1010 B.n57 585
R984 B.n1155 B.n57 585
R985 B.n1009 B.n56 585
R986 B.n1156 B.n56 585
R987 B.n1008 B.n55 585
R988 B.n1157 B.n55 585
R989 B.n1007 B.n1006 585
R990 B.n1006 B.n51 585
R991 B.n1005 B.n50 585
R992 B.n1163 B.n50 585
R993 B.n1004 B.n49 585
R994 B.n1164 B.n49 585
R995 B.n1003 B.n48 585
R996 B.n1165 B.n48 585
R997 B.n1002 B.n1001 585
R998 B.n1001 B.n44 585
R999 B.n1000 B.n43 585
R1000 B.n1171 B.n43 585
R1001 B.n999 B.n42 585
R1002 B.n1172 B.n42 585
R1003 B.n998 B.n41 585
R1004 B.n1173 B.n41 585
R1005 B.n997 B.n996 585
R1006 B.n996 B.n37 585
R1007 B.n995 B.n36 585
R1008 B.n1179 B.n36 585
R1009 B.n994 B.n35 585
R1010 B.n1180 B.n35 585
R1011 B.n993 B.n34 585
R1012 B.n1181 B.n34 585
R1013 B.n992 B.n991 585
R1014 B.n991 B.n30 585
R1015 B.n990 B.n29 585
R1016 B.n1187 B.n29 585
R1017 B.n989 B.n28 585
R1018 B.n1188 B.n28 585
R1019 B.n988 B.n27 585
R1020 B.n1189 B.n27 585
R1021 B.n987 B.n986 585
R1022 B.n986 B.n23 585
R1023 B.n985 B.n22 585
R1024 B.n1195 B.n22 585
R1025 B.n984 B.n21 585
R1026 B.n1196 B.n21 585
R1027 B.n983 B.n20 585
R1028 B.n1197 B.n20 585
R1029 B.n982 B.n981 585
R1030 B.n981 B.n19 585
R1031 B.n980 B.n15 585
R1032 B.n1203 B.n15 585
R1033 B.n979 B.n14 585
R1034 B.n1204 B.n14 585
R1035 B.n978 B.n13 585
R1036 B.n1205 B.n13 585
R1037 B.n977 B.n976 585
R1038 B.n976 B.n12 585
R1039 B.n975 B.n974 585
R1040 B.n975 B.n8 585
R1041 B.n973 B.n7 585
R1042 B.n1212 B.n7 585
R1043 B.n972 B.n6 585
R1044 B.n1213 B.n6 585
R1045 B.n971 B.n5 585
R1046 B.n1214 B.n5 585
R1047 B.n970 B.n969 585
R1048 B.n969 B.n4 585
R1049 B.n968 B.n370 585
R1050 B.n968 B.n967 585
R1051 B.n958 B.n371 585
R1052 B.n372 B.n371 585
R1053 B.n960 B.n959 585
R1054 B.n961 B.n960 585
R1055 B.n957 B.n377 585
R1056 B.n377 B.n376 585
R1057 B.n956 B.n955 585
R1058 B.n955 B.n954 585
R1059 B.n379 B.n378 585
R1060 B.n947 B.n379 585
R1061 B.n946 B.n945 585
R1062 B.n948 B.n946 585
R1063 B.n944 B.n384 585
R1064 B.n384 B.n383 585
R1065 B.n943 B.n942 585
R1066 B.n942 B.n941 585
R1067 B.n386 B.n385 585
R1068 B.n387 B.n386 585
R1069 B.n934 B.n933 585
R1070 B.n935 B.n934 585
R1071 B.n932 B.n392 585
R1072 B.n392 B.n391 585
R1073 B.n931 B.n930 585
R1074 B.n930 B.n929 585
R1075 B.n394 B.n393 585
R1076 B.n395 B.n394 585
R1077 B.n922 B.n921 585
R1078 B.n923 B.n922 585
R1079 B.n920 B.n400 585
R1080 B.n400 B.n399 585
R1081 B.n919 B.n918 585
R1082 B.n918 B.n917 585
R1083 B.n402 B.n401 585
R1084 B.n403 B.n402 585
R1085 B.n910 B.n909 585
R1086 B.n911 B.n910 585
R1087 B.n908 B.n408 585
R1088 B.n408 B.n407 585
R1089 B.n907 B.n906 585
R1090 B.n906 B.n905 585
R1091 B.n410 B.n409 585
R1092 B.n411 B.n410 585
R1093 B.n898 B.n897 585
R1094 B.n899 B.n898 585
R1095 B.n896 B.n416 585
R1096 B.n416 B.n415 585
R1097 B.n895 B.n894 585
R1098 B.n894 B.n893 585
R1099 B.n418 B.n417 585
R1100 B.n419 B.n418 585
R1101 B.n886 B.n885 585
R1102 B.n887 B.n886 585
R1103 B.n884 B.n423 585
R1104 B.n427 B.n423 585
R1105 B.n883 B.n882 585
R1106 B.n882 B.n881 585
R1107 B.n425 B.n424 585
R1108 B.n426 B.n425 585
R1109 B.n874 B.n873 585
R1110 B.n875 B.n874 585
R1111 B.n872 B.n432 585
R1112 B.n432 B.n431 585
R1113 B.n871 B.n870 585
R1114 B.n870 B.n869 585
R1115 B.n434 B.n433 585
R1116 B.n435 B.n434 585
R1117 B.n862 B.n861 585
R1118 B.n863 B.n862 585
R1119 B.n860 B.n440 585
R1120 B.n440 B.n439 585
R1121 B.n859 B.n858 585
R1122 B.n858 B.n857 585
R1123 B.n442 B.n441 585
R1124 B.n443 B.n442 585
R1125 B.n850 B.n849 585
R1126 B.n851 B.n850 585
R1127 B.n848 B.n448 585
R1128 B.n448 B.n447 585
R1129 B.n847 B.n846 585
R1130 B.n846 B.n845 585
R1131 B.n450 B.n449 585
R1132 B.n451 B.n450 585
R1133 B.n838 B.n837 585
R1134 B.n839 B.n838 585
R1135 B.n836 B.n456 585
R1136 B.n456 B.n455 585
R1137 B.n835 B.n834 585
R1138 B.n834 B.n833 585
R1139 B.n458 B.n457 585
R1140 B.n459 B.n458 585
R1141 B.n826 B.n825 585
R1142 B.n827 B.n826 585
R1143 B.n824 B.n464 585
R1144 B.n464 B.n463 585
R1145 B.n823 B.n822 585
R1146 B.n822 B.n821 585
R1147 B.n466 B.n465 585
R1148 B.n814 B.n466 585
R1149 B.n813 B.n812 585
R1150 B.n815 B.n813 585
R1151 B.n811 B.n471 585
R1152 B.n471 B.n470 585
R1153 B.n810 B.n809 585
R1154 B.n809 B.n808 585
R1155 B.n473 B.n472 585
R1156 B.n474 B.n473 585
R1157 B.n801 B.n800 585
R1158 B.n802 B.n801 585
R1159 B.n799 B.n479 585
R1160 B.n479 B.n478 585
R1161 B.n798 B.n797 585
R1162 B.n797 B.n796 585
R1163 B.n481 B.n480 585
R1164 B.n482 B.n481 585
R1165 B.n789 B.n788 585
R1166 B.n790 B.n789 585
R1167 B.n787 B.n487 585
R1168 B.n487 B.n486 585
R1169 B.n786 B.n785 585
R1170 B.n785 B.n784 585
R1171 B.n489 B.n488 585
R1172 B.n490 B.n489 585
R1173 B.n777 B.n776 585
R1174 B.n778 B.n777 585
R1175 B.n775 B.n494 585
R1176 B.n498 B.n494 585
R1177 B.n774 B.n773 585
R1178 B.n773 B.n772 585
R1179 B.n496 B.n495 585
R1180 B.n497 B.n496 585
R1181 B.n765 B.n764 585
R1182 B.n766 B.n765 585
R1183 B.n763 B.n503 585
R1184 B.n503 B.n502 585
R1185 B.n762 B.n761 585
R1186 B.n761 B.n760 585
R1187 B.n505 B.n504 585
R1188 B.n506 B.n505 585
R1189 B.n753 B.n752 585
R1190 B.n754 B.n753 585
R1191 B.n751 B.n511 585
R1192 B.n511 B.n510 585
R1193 B.n745 B.n744 585
R1194 B.n743 B.n559 585
R1195 B.n742 B.n558 585
R1196 B.n747 B.n558 585
R1197 B.n741 B.n740 585
R1198 B.n739 B.n738 585
R1199 B.n737 B.n736 585
R1200 B.n735 B.n734 585
R1201 B.n733 B.n732 585
R1202 B.n731 B.n730 585
R1203 B.n729 B.n728 585
R1204 B.n727 B.n726 585
R1205 B.n725 B.n724 585
R1206 B.n723 B.n722 585
R1207 B.n721 B.n720 585
R1208 B.n719 B.n718 585
R1209 B.n717 B.n716 585
R1210 B.n715 B.n714 585
R1211 B.n713 B.n712 585
R1212 B.n711 B.n710 585
R1213 B.n709 B.n708 585
R1214 B.n707 B.n706 585
R1215 B.n705 B.n704 585
R1216 B.n703 B.n702 585
R1217 B.n701 B.n700 585
R1218 B.n699 B.n698 585
R1219 B.n697 B.n696 585
R1220 B.n695 B.n694 585
R1221 B.n693 B.n692 585
R1222 B.n691 B.n690 585
R1223 B.n689 B.n688 585
R1224 B.n687 B.n686 585
R1225 B.n685 B.n684 585
R1226 B.n683 B.n682 585
R1227 B.n681 B.n680 585
R1228 B.n679 B.n678 585
R1229 B.n677 B.n676 585
R1230 B.n675 B.n674 585
R1231 B.n673 B.n672 585
R1232 B.n671 B.n670 585
R1233 B.n669 B.n668 585
R1234 B.n667 B.n666 585
R1235 B.n665 B.n664 585
R1236 B.n662 B.n661 585
R1237 B.n660 B.n659 585
R1238 B.n658 B.n657 585
R1239 B.n656 B.n655 585
R1240 B.n654 B.n653 585
R1241 B.n652 B.n651 585
R1242 B.n650 B.n649 585
R1243 B.n648 B.n647 585
R1244 B.n646 B.n645 585
R1245 B.n644 B.n643 585
R1246 B.n642 B.n641 585
R1247 B.n640 B.n639 585
R1248 B.n638 B.n637 585
R1249 B.n636 B.n635 585
R1250 B.n634 B.n633 585
R1251 B.n632 B.n631 585
R1252 B.n630 B.n629 585
R1253 B.n628 B.n627 585
R1254 B.n626 B.n625 585
R1255 B.n624 B.n623 585
R1256 B.n622 B.n621 585
R1257 B.n620 B.n619 585
R1258 B.n618 B.n617 585
R1259 B.n616 B.n615 585
R1260 B.n614 B.n613 585
R1261 B.n612 B.n611 585
R1262 B.n610 B.n609 585
R1263 B.n608 B.n607 585
R1264 B.n606 B.n605 585
R1265 B.n604 B.n603 585
R1266 B.n602 B.n601 585
R1267 B.n600 B.n599 585
R1268 B.n598 B.n597 585
R1269 B.n596 B.n595 585
R1270 B.n594 B.n593 585
R1271 B.n592 B.n591 585
R1272 B.n590 B.n589 585
R1273 B.n588 B.n587 585
R1274 B.n586 B.n585 585
R1275 B.n584 B.n583 585
R1276 B.n582 B.n581 585
R1277 B.n580 B.n579 585
R1278 B.n578 B.n577 585
R1279 B.n576 B.n575 585
R1280 B.n574 B.n573 585
R1281 B.n572 B.n571 585
R1282 B.n570 B.n569 585
R1283 B.n568 B.n567 585
R1284 B.n566 B.n565 585
R1285 B.n513 B.n512 585
R1286 B.n750 B.n749 585
R1287 B.n509 B.n508 585
R1288 B.n510 B.n509 585
R1289 B.n756 B.n755 585
R1290 B.n755 B.n754 585
R1291 B.n757 B.n507 585
R1292 B.n507 B.n506 585
R1293 B.n759 B.n758 585
R1294 B.n760 B.n759 585
R1295 B.n501 B.n500 585
R1296 B.n502 B.n501 585
R1297 B.n768 B.n767 585
R1298 B.n767 B.n766 585
R1299 B.n769 B.n499 585
R1300 B.n499 B.n497 585
R1301 B.n771 B.n770 585
R1302 B.n772 B.n771 585
R1303 B.n493 B.n492 585
R1304 B.n498 B.n493 585
R1305 B.n780 B.n779 585
R1306 B.n779 B.n778 585
R1307 B.n781 B.n491 585
R1308 B.n491 B.n490 585
R1309 B.n783 B.n782 585
R1310 B.n784 B.n783 585
R1311 B.n485 B.n484 585
R1312 B.n486 B.n485 585
R1313 B.n792 B.n791 585
R1314 B.n791 B.n790 585
R1315 B.n793 B.n483 585
R1316 B.n483 B.n482 585
R1317 B.n795 B.n794 585
R1318 B.n796 B.n795 585
R1319 B.n477 B.n476 585
R1320 B.n478 B.n477 585
R1321 B.n804 B.n803 585
R1322 B.n803 B.n802 585
R1323 B.n805 B.n475 585
R1324 B.n475 B.n474 585
R1325 B.n807 B.n806 585
R1326 B.n808 B.n807 585
R1327 B.n469 B.n468 585
R1328 B.n470 B.n469 585
R1329 B.n817 B.n816 585
R1330 B.n816 B.n815 585
R1331 B.n818 B.n467 585
R1332 B.n814 B.n467 585
R1333 B.n820 B.n819 585
R1334 B.n821 B.n820 585
R1335 B.n462 B.n461 585
R1336 B.n463 B.n462 585
R1337 B.n829 B.n828 585
R1338 B.n828 B.n827 585
R1339 B.n830 B.n460 585
R1340 B.n460 B.n459 585
R1341 B.n832 B.n831 585
R1342 B.n833 B.n832 585
R1343 B.n454 B.n453 585
R1344 B.n455 B.n454 585
R1345 B.n841 B.n840 585
R1346 B.n840 B.n839 585
R1347 B.n842 B.n452 585
R1348 B.n452 B.n451 585
R1349 B.n844 B.n843 585
R1350 B.n845 B.n844 585
R1351 B.n446 B.n445 585
R1352 B.n447 B.n446 585
R1353 B.n853 B.n852 585
R1354 B.n852 B.n851 585
R1355 B.n854 B.n444 585
R1356 B.n444 B.n443 585
R1357 B.n856 B.n855 585
R1358 B.n857 B.n856 585
R1359 B.n438 B.n437 585
R1360 B.n439 B.n438 585
R1361 B.n865 B.n864 585
R1362 B.n864 B.n863 585
R1363 B.n866 B.n436 585
R1364 B.n436 B.n435 585
R1365 B.n868 B.n867 585
R1366 B.n869 B.n868 585
R1367 B.n430 B.n429 585
R1368 B.n431 B.n430 585
R1369 B.n877 B.n876 585
R1370 B.n876 B.n875 585
R1371 B.n878 B.n428 585
R1372 B.n428 B.n426 585
R1373 B.n880 B.n879 585
R1374 B.n881 B.n880 585
R1375 B.n422 B.n421 585
R1376 B.n427 B.n422 585
R1377 B.n889 B.n888 585
R1378 B.n888 B.n887 585
R1379 B.n890 B.n420 585
R1380 B.n420 B.n419 585
R1381 B.n892 B.n891 585
R1382 B.n893 B.n892 585
R1383 B.n414 B.n413 585
R1384 B.n415 B.n414 585
R1385 B.n901 B.n900 585
R1386 B.n900 B.n899 585
R1387 B.n902 B.n412 585
R1388 B.n412 B.n411 585
R1389 B.n904 B.n903 585
R1390 B.n905 B.n904 585
R1391 B.n406 B.n405 585
R1392 B.n407 B.n406 585
R1393 B.n913 B.n912 585
R1394 B.n912 B.n911 585
R1395 B.n914 B.n404 585
R1396 B.n404 B.n403 585
R1397 B.n916 B.n915 585
R1398 B.n917 B.n916 585
R1399 B.n398 B.n397 585
R1400 B.n399 B.n398 585
R1401 B.n925 B.n924 585
R1402 B.n924 B.n923 585
R1403 B.n926 B.n396 585
R1404 B.n396 B.n395 585
R1405 B.n928 B.n927 585
R1406 B.n929 B.n928 585
R1407 B.n390 B.n389 585
R1408 B.n391 B.n390 585
R1409 B.n937 B.n936 585
R1410 B.n936 B.n935 585
R1411 B.n938 B.n388 585
R1412 B.n388 B.n387 585
R1413 B.n940 B.n939 585
R1414 B.n941 B.n940 585
R1415 B.n382 B.n381 585
R1416 B.n383 B.n382 585
R1417 B.n950 B.n949 585
R1418 B.n949 B.n948 585
R1419 B.n951 B.n380 585
R1420 B.n947 B.n380 585
R1421 B.n953 B.n952 585
R1422 B.n954 B.n953 585
R1423 B.n375 B.n374 585
R1424 B.n376 B.n375 585
R1425 B.n963 B.n962 585
R1426 B.n962 B.n961 585
R1427 B.n964 B.n373 585
R1428 B.n373 B.n372 585
R1429 B.n966 B.n965 585
R1430 B.n967 B.n966 585
R1431 B.n3 B.n0 585
R1432 B.n4 B.n3 585
R1433 B.n1211 B.n1 585
R1434 B.n1212 B.n1211 585
R1435 B.n1210 B.n1209 585
R1436 B.n1210 B.n8 585
R1437 B.n1208 B.n9 585
R1438 B.n12 B.n9 585
R1439 B.n1207 B.n1206 585
R1440 B.n1206 B.n1205 585
R1441 B.n11 B.n10 585
R1442 B.n1204 B.n11 585
R1443 B.n1202 B.n1201 585
R1444 B.n1203 B.n1202 585
R1445 B.n1200 B.n16 585
R1446 B.n19 B.n16 585
R1447 B.n1199 B.n1198 585
R1448 B.n1198 B.n1197 585
R1449 B.n18 B.n17 585
R1450 B.n1196 B.n18 585
R1451 B.n1194 B.n1193 585
R1452 B.n1195 B.n1194 585
R1453 B.n1192 B.n24 585
R1454 B.n24 B.n23 585
R1455 B.n1191 B.n1190 585
R1456 B.n1190 B.n1189 585
R1457 B.n26 B.n25 585
R1458 B.n1188 B.n26 585
R1459 B.n1186 B.n1185 585
R1460 B.n1187 B.n1186 585
R1461 B.n1184 B.n31 585
R1462 B.n31 B.n30 585
R1463 B.n1183 B.n1182 585
R1464 B.n1182 B.n1181 585
R1465 B.n33 B.n32 585
R1466 B.n1180 B.n33 585
R1467 B.n1178 B.n1177 585
R1468 B.n1179 B.n1178 585
R1469 B.n1176 B.n38 585
R1470 B.n38 B.n37 585
R1471 B.n1175 B.n1174 585
R1472 B.n1174 B.n1173 585
R1473 B.n40 B.n39 585
R1474 B.n1172 B.n40 585
R1475 B.n1170 B.n1169 585
R1476 B.n1171 B.n1170 585
R1477 B.n1168 B.n45 585
R1478 B.n45 B.n44 585
R1479 B.n1167 B.n1166 585
R1480 B.n1166 B.n1165 585
R1481 B.n47 B.n46 585
R1482 B.n1164 B.n47 585
R1483 B.n1162 B.n1161 585
R1484 B.n1163 B.n1162 585
R1485 B.n1160 B.n52 585
R1486 B.n52 B.n51 585
R1487 B.n1159 B.n1158 585
R1488 B.n1158 B.n1157 585
R1489 B.n54 B.n53 585
R1490 B.n1156 B.n54 585
R1491 B.n1154 B.n1153 585
R1492 B.n1155 B.n1154 585
R1493 B.n1152 B.n59 585
R1494 B.n59 B.n58 585
R1495 B.n1151 B.n1150 585
R1496 B.n1150 B.n1149 585
R1497 B.n61 B.n60 585
R1498 B.n1148 B.n61 585
R1499 B.n1146 B.n1145 585
R1500 B.n1147 B.n1146 585
R1501 B.n1144 B.n66 585
R1502 B.n66 B.n65 585
R1503 B.n1143 B.n1142 585
R1504 B.n1142 B.n1141 585
R1505 B.n68 B.n67 585
R1506 B.n1140 B.n68 585
R1507 B.n1138 B.n1137 585
R1508 B.n1139 B.n1138 585
R1509 B.n1136 B.n73 585
R1510 B.n73 B.n72 585
R1511 B.n1135 B.n1134 585
R1512 B.n1134 B.n1133 585
R1513 B.n75 B.n74 585
R1514 B.n1132 B.n75 585
R1515 B.n1130 B.n1129 585
R1516 B.n1131 B.n1130 585
R1517 B.n1128 B.n80 585
R1518 B.n80 B.n79 585
R1519 B.n1127 B.n1126 585
R1520 B.n1126 B.n1125 585
R1521 B.n82 B.n81 585
R1522 B.n1124 B.n82 585
R1523 B.n1122 B.n1121 585
R1524 B.n1123 B.n1122 585
R1525 B.n1120 B.n87 585
R1526 B.n87 B.n86 585
R1527 B.n1119 B.n1118 585
R1528 B.n1118 B.n1117 585
R1529 B.n89 B.n88 585
R1530 B.n1116 B.n89 585
R1531 B.n1114 B.n1113 585
R1532 B.n1115 B.n1114 585
R1533 B.n1112 B.n93 585
R1534 B.n96 B.n93 585
R1535 B.n1111 B.n1110 585
R1536 B.n1110 B.n1109 585
R1537 B.n95 B.n94 585
R1538 B.n1108 B.n95 585
R1539 B.n1106 B.n1105 585
R1540 B.n1107 B.n1106 585
R1541 B.n1104 B.n101 585
R1542 B.n101 B.n100 585
R1543 B.n1103 B.n1102 585
R1544 B.n1102 B.n1101 585
R1545 B.n103 B.n102 585
R1546 B.n1100 B.n103 585
R1547 B.n1098 B.n1097 585
R1548 B.n1099 B.n1098 585
R1549 B.n1096 B.n108 585
R1550 B.n108 B.n107 585
R1551 B.n1095 B.n1094 585
R1552 B.n1094 B.n1093 585
R1553 B.n110 B.n109 585
R1554 B.n1092 B.n110 585
R1555 B.n1090 B.n1089 585
R1556 B.n1091 B.n1090 585
R1557 B.n1088 B.n115 585
R1558 B.n115 B.n114 585
R1559 B.n1087 B.n1086 585
R1560 B.n1086 B.n1085 585
R1561 B.n117 B.n116 585
R1562 B.n1084 B.n117 585
R1563 B.n1082 B.n1081 585
R1564 B.n1083 B.n1082 585
R1565 B.n1080 B.n122 585
R1566 B.n122 B.n121 585
R1567 B.n1079 B.n1078 585
R1568 B.n1078 B.n1077 585
R1569 B.n124 B.n123 585
R1570 B.n1076 B.n124 585
R1571 B.n1074 B.n1073 585
R1572 B.n1075 B.n1074 585
R1573 B.n1072 B.n129 585
R1574 B.n129 B.n128 585
R1575 B.n1071 B.n1070 585
R1576 B.n1070 B.n1069 585
R1577 B.n131 B.n130 585
R1578 B.n1068 B.n131 585
R1579 B.n1215 B.n1214 585
R1580 B.n1213 B.n2 585
R1581 B.n186 B.n131 468.476
R1582 B.n1066 B.n133 468.476
R1583 B.n749 B.n511 468.476
R1584 B.n745 B.n509 468.476
R1585 B.n181 B.t22 353.765
R1586 B.n562 B.t13 353.765
R1587 B.n183 B.t16 353.765
R1588 B.n560 B.t20 353.765
R1589 B.n183 B.t14 294.789
R1590 B.n181 B.t21 294.789
R1591 B.n562 B.t10 294.789
R1592 B.n560 B.t18 294.789
R1593 B.n182 B.t23 282.009
R1594 B.n563 B.t12 282.009
R1595 B.n184 B.t17 282.009
R1596 B.n561 B.t19 282.009
R1597 B.n1067 B.n179 256.663
R1598 B.n1067 B.n178 256.663
R1599 B.n1067 B.n177 256.663
R1600 B.n1067 B.n176 256.663
R1601 B.n1067 B.n175 256.663
R1602 B.n1067 B.n174 256.663
R1603 B.n1067 B.n173 256.663
R1604 B.n1067 B.n172 256.663
R1605 B.n1067 B.n171 256.663
R1606 B.n1067 B.n170 256.663
R1607 B.n1067 B.n169 256.663
R1608 B.n1067 B.n168 256.663
R1609 B.n1067 B.n167 256.663
R1610 B.n1067 B.n166 256.663
R1611 B.n1067 B.n165 256.663
R1612 B.n1067 B.n164 256.663
R1613 B.n1067 B.n163 256.663
R1614 B.n1067 B.n162 256.663
R1615 B.n1067 B.n161 256.663
R1616 B.n1067 B.n160 256.663
R1617 B.n1067 B.n159 256.663
R1618 B.n1067 B.n158 256.663
R1619 B.n1067 B.n157 256.663
R1620 B.n1067 B.n156 256.663
R1621 B.n1067 B.n155 256.663
R1622 B.n1067 B.n154 256.663
R1623 B.n1067 B.n153 256.663
R1624 B.n1067 B.n152 256.663
R1625 B.n1067 B.n151 256.663
R1626 B.n1067 B.n150 256.663
R1627 B.n1067 B.n149 256.663
R1628 B.n1067 B.n148 256.663
R1629 B.n1067 B.n147 256.663
R1630 B.n1067 B.n146 256.663
R1631 B.n1067 B.n145 256.663
R1632 B.n1067 B.n144 256.663
R1633 B.n1067 B.n143 256.663
R1634 B.n1067 B.n142 256.663
R1635 B.n1067 B.n141 256.663
R1636 B.n1067 B.n140 256.663
R1637 B.n1067 B.n139 256.663
R1638 B.n1067 B.n138 256.663
R1639 B.n1067 B.n137 256.663
R1640 B.n1067 B.n136 256.663
R1641 B.n1067 B.n135 256.663
R1642 B.n1067 B.n134 256.663
R1643 B.n747 B.n746 256.663
R1644 B.n747 B.n514 256.663
R1645 B.n747 B.n515 256.663
R1646 B.n747 B.n516 256.663
R1647 B.n747 B.n517 256.663
R1648 B.n747 B.n518 256.663
R1649 B.n747 B.n519 256.663
R1650 B.n747 B.n520 256.663
R1651 B.n747 B.n521 256.663
R1652 B.n747 B.n522 256.663
R1653 B.n747 B.n523 256.663
R1654 B.n747 B.n524 256.663
R1655 B.n747 B.n525 256.663
R1656 B.n747 B.n526 256.663
R1657 B.n747 B.n527 256.663
R1658 B.n747 B.n528 256.663
R1659 B.n747 B.n529 256.663
R1660 B.n747 B.n530 256.663
R1661 B.n747 B.n531 256.663
R1662 B.n747 B.n532 256.663
R1663 B.n747 B.n533 256.663
R1664 B.n747 B.n534 256.663
R1665 B.n747 B.n535 256.663
R1666 B.n747 B.n536 256.663
R1667 B.n747 B.n537 256.663
R1668 B.n747 B.n538 256.663
R1669 B.n747 B.n539 256.663
R1670 B.n747 B.n540 256.663
R1671 B.n747 B.n541 256.663
R1672 B.n747 B.n542 256.663
R1673 B.n747 B.n543 256.663
R1674 B.n747 B.n544 256.663
R1675 B.n747 B.n545 256.663
R1676 B.n747 B.n546 256.663
R1677 B.n747 B.n547 256.663
R1678 B.n747 B.n548 256.663
R1679 B.n747 B.n549 256.663
R1680 B.n747 B.n550 256.663
R1681 B.n747 B.n551 256.663
R1682 B.n747 B.n552 256.663
R1683 B.n747 B.n553 256.663
R1684 B.n747 B.n554 256.663
R1685 B.n747 B.n555 256.663
R1686 B.n747 B.n556 256.663
R1687 B.n747 B.n557 256.663
R1688 B.n748 B.n747 256.663
R1689 B.n1217 B.n1216 256.663
R1690 B.n190 B.n189 163.367
R1691 B.n194 B.n193 163.367
R1692 B.n198 B.n197 163.367
R1693 B.n202 B.n201 163.367
R1694 B.n206 B.n205 163.367
R1695 B.n210 B.n209 163.367
R1696 B.n214 B.n213 163.367
R1697 B.n218 B.n217 163.367
R1698 B.n222 B.n221 163.367
R1699 B.n226 B.n225 163.367
R1700 B.n230 B.n229 163.367
R1701 B.n234 B.n233 163.367
R1702 B.n238 B.n237 163.367
R1703 B.n242 B.n241 163.367
R1704 B.n246 B.n245 163.367
R1705 B.n250 B.n249 163.367
R1706 B.n254 B.n253 163.367
R1707 B.n258 B.n257 163.367
R1708 B.n262 B.n261 163.367
R1709 B.n266 B.n265 163.367
R1710 B.n270 B.n269 163.367
R1711 B.n274 B.n273 163.367
R1712 B.n278 B.n277 163.367
R1713 B.n282 B.n281 163.367
R1714 B.n286 B.n285 163.367
R1715 B.n291 B.n290 163.367
R1716 B.n295 B.n294 163.367
R1717 B.n299 B.n298 163.367
R1718 B.n303 B.n302 163.367
R1719 B.n307 B.n306 163.367
R1720 B.n311 B.n310 163.367
R1721 B.n315 B.n314 163.367
R1722 B.n319 B.n318 163.367
R1723 B.n323 B.n322 163.367
R1724 B.n327 B.n326 163.367
R1725 B.n331 B.n330 163.367
R1726 B.n335 B.n334 163.367
R1727 B.n339 B.n338 163.367
R1728 B.n343 B.n342 163.367
R1729 B.n347 B.n346 163.367
R1730 B.n351 B.n350 163.367
R1731 B.n355 B.n354 163.367
R1732 B.n359 B.n358 163.367
R1733 B.n363 B.n362 163.367
R1734 B.n367 B.n366 163.367
R1735 B.n1066 B.n180 163.367
R1736 B.n753 B.n511 163.367
R1737 B.n753 B.n505 163.367
R1738 B.n761 B.n505 163.367
R1739 B.n761 B.n503 163.367
R1740 B.n765 B.n503 163.367
R1741 B.n765 B.n496 163.367
R1742 B.n773 B.n496 163.367
R1743 B.n773 B.n494 163.367
R1744 B.n777 B.n494 163.367
R1745 B.n777 B.n489 163.367
R1746 B.n785 B.n489 163.367
R1747 B.n785 B.n487 163.367
R1748 B.n789 B.n487 163.367
R1749 B.n789 B.n481 163.367
R1750 B.n797 B.n481 163.367
R1751 B.n797 B.n479 163.367
R1752 B.n801 B.n479 163.367
R1753 B.n801 B.n473 163.367
R1754 B.n809 B.n473 163.367
R1755 B.n809 B.n471 163.367
R1756 B.n813 B.n471 163.367
R1757 B.n813 B.n466 163.367
R1758 B.n822 B.n466 163.367
R1759 B.n822 B.n464 163.367
R1760 B.n826 B.n464 163.367
R1761 B.n826 B.n458 163.367
R1762 B.n834 B.n458 163.367
R1763 B.n834 B.n456 163.367
R1764 B.n838 B.n456 163.367
R1765 B.n838 B.n450 163.367
R1766 B.n846 B.n450 163.367
R1767 B.n846 B.n448 163.367
R1768 B.n850 B.n448 163.367
R1769 B.n850 B.n442 163.367
R1770 B.n858 B.n442 163.367
R1771 B.n858 B.n440 163.367
R1772 B.n862 B.n440 163.367
R1773 B.n862 B.n434 163.367
R1774 B.n870 B.n434 163.367
R1775 B.n870 B.n432 163.367
R1776 B.n874 B.n432 163.367
R1777 B.n874 B.n425 163.367
R1778 B.n882 B.n425 163.367
R1779 B.n882 B.n423 163.367
R1780 B.n886 B.n423 163.367
R1781 B.n886 B.n418 163.367
R1782 B.n894 B.n418 163.367
R1783 B.n894 B.n416 163.367
R1784 B.n898 B.n416 163.367
R1785 B.n898 B.n410 163.367
R1786 B.n906 B.n410 163.367
R1787 B.n906 B.n408 163.367
R1788 B.n910 B.n408 163.367
R1789 B.n910 B.n402 163.367
R1790 B.n918 B.n402 163.367
R1791 B.n918 B.n400 163.367
R1792 B.n922 B.n400 163.367
R1793 B.n922 B.n394 163.367
R1794 B.n930 B.n394 163.367
R1795 B.n930 B.n392 163.367
R1796 B.n934 B.n392 163.367
R1797 B.n934 B.n386 163.367
R1798 B.n942 B.n386 163.367
R1799 B.n942 B.n384 163.367
R1800 B.n946 B.n384 163.367
R1801 B.n946 B.n379 163.367
R1802 B.n955 B.n379 163.367
R1803 B.n955 B.n377 163.367
R1804 B.n960 B.n377 163.367
R1805 B.n960 B.n371 163.367
R1806 B.n968 B.n371 163.367
R1807 B.n969 B.n968 163.367
R1808 B.n969 B.n5 163.367
R1809 B.n6 B.n5 163.367
R1810 B.n7 B.n6 163.367
R1811 B.n975 B.n7 163.367
R1812 B.n976 B.n975 163.367
R1813 B.n976 B.n13 163.367
R1814 B.n14 B.n13 163.367
R1815 B.n15 B.n14 163.367
R1816 B.n981 B.n15 163.367
R1817 B.n981 B.n20 163.367
R1818 B.n21 B.n20 163.367
R1819 B.n22 B.n21 163.367
R1820 B.n986 B.n22 163.367
R1821 B.n986 B.n27 163.367
R1822 B.n28 B.n27 163.367
R1823 B.n29 B.n28 163.367
R1824 B.n991 B.n29 163.367
R1825 B.n991 B.n34 163.367
R1826 B.n35 B.n34 163.367
R1827 B.n36 B.n35 163.367
R1828 B.n996 B.n36 163.367
R1829 B.n996 B.n41 163.367
R1830 B.n42 B.n41 163.367
R1831 B.n43 B.n42 163.367
R1832 B.n1001 B.n43 163.367
R1833 B.n1001 B.n48 163.367
R1834 B.n49 B.n48 163.367
R1835 B.n50 B.n49 163.367
R1836 B.n1006 B.n50 163.367
R1837 B.n1006 B.n55 163.367
R1838 B.n56 B.n55 163.367
R1839 B.n57 B.n56 163.367
R1840 B.n1011 B.n57 163.367
R1841 B.n1011 B.n62 163.367
R1842 B.n63 B.n62 163.367
R1843 B.n64 B.n63 163.367
R1844 B.n1016 B.n64 163.367
R1845 B.n1016 B.n69 163.367
R1846 B.n70 B.n69 163.367
R1847 B.n71 B.n70 163.367
R1848 B.n1021 B.n71 163.367
R1849 B.n1021 B.n76 163.367
R1850 B.n77 B.n76 163.367
R1851 B.n78 B.n77 163.367
R1852 B.n1026 B.n78 163.367
R1853 B.n1026 B.n83 163.367
R1854 B.n84 B.n83 163.367
R1855 B.n85 B.n84 163.367
R1856 B.n1031 B.n85 163.367
R1857 B.n1031 B.n90 163.367
R1858 B.n91 B.n90 163.367
R1859 B.n92 B.n91 163.367
R1860 B.n1036 B.n92 163.367
R1861 B.n1036 B.n97 163.367
R1862 B.n98 B.n97 163.367
R1863 B.n99 B.n98 163.367
R1864 B.n1041 B.n99 163.367
R1865 B.n1041 B.n104 163.367
R1866 B.n105 B.n104 163.367
R1867 B.n106 B.n105 163.367
R1868 B.n1046 B.n106 163.367
R1869 B.n1046 B.n111 163.367
R1870 B.n112 B.n111 163.367
R1871 B.n113 B.n112 163.367
R1872 B.n1051 B.n113 163.367
R1873 B.n1051 B.n118 163.367
R1874 B.n119 B.n118 163.367
R1875 B.n120 B.n119 163.367
R1876 B.n1056 B.n120 163.367
R1877 B.n1056 B.n125 163.367
R1878 B.n126 B.n125 163.367
R1879 B.n127 B.n126 163.367
R1880 B.n1061 B.n127 163.367
R1881 B.n1061 B.n132 163.367
R1882 B.n133 B.n132 163.367
R1883 B.n559 B.n558 163.367
R1884 B.n740 B.n558 163.367
R1885 B.n738 B.n737 163.367
R1886 B.n734 B.n733 163.367
R1887 B.n730 B.n729 163.367
R1888 B.n726 B.n725 163.367
R1889 B.n722 B.n721 163.367
R1890 B.n718 B.n717 163.367
R1891 B.n714 B.n713 163.367
R1892 B.n710 B.n709 163.367
R1893 B.n706 B.n705 163.367
R1894 B.n702 B.n701 163.367
R1895 B.n698 B.n697 163.367
R1896 B.n694 B.n693 163.367
R1897 B.n690 B.n689 163.367
R1898 B.n686 B.n685 163.367
R1899 B.n682 B.n681 163.367
R1900 B.n678 B.n677 163.367
R1901 B.n674 B.n673 163.367
R1902 B.n670 B.n669 163.367
R1903 B.n666 B.n665 163.367
R1904 B.n661 B.n660 163.367
R1905 B.n657 B.n656 163.367
R1906 B.n653 B.n652 163.367
R1907 B.n649 B.n648 163.367
R1908 B.n645 B.n644 163.367
R1909 B.n641 B.n640 163.367
R1910 B.n637 B.n636 163.367
R1911 B.n633 B.n632 163.367
R1912 B.n629 B.n628 163.367
R1913 B.n625 B.n624 163.367
R1914 B.n621 B.n620 163.367
R1915 B.n617 B.n616 163.367
R1916 B.n613 B.n612 163.367
R1917 B.n609 B.n608 163.367
R1918 B.n605 B.n604 163.367
R1919 B.n601 B.n600 163.367
R1920 B.n597 B.n596 163.367
R1921 B.n593 B.n592 163.367
R1922 B.n589 B.n588 163.367
R1923 B.n585 B.n584 163.367
R1924 B.n581 B.n580 163.367
R1925 B.n577 B.n576 163.367
R1926 B.n573 B.n572 163.367
R1927 B.n569 B.n568 163.367
R1928 B.n565 B.n513 163.367
R1929 B.n755 B.n509 163.367
R1930 B.n755 B.n507 163.367
R1931 B.n759 B.n507 163.367
R1932 B.n759 B.n501 163.367
R1933 B.n767 B.n501 163.367
R1934 B.n767 B.n499 163.367
R1935 B.n771 B.n499 163.367
R1936 B.n771 B.n493 163.367
R1937 B.n779 B.n493 163.367
R1938 B.n779 B.n491 163.367
R1939 B.n783 B.n491 163.367
R1940 B.n783 B.n485 163.367
R1941 B.n791 B.n485 163.367
R1942 B.n791 B.n483 163.367
R1943 B.n795 B.n483 163.367
R1944 B.n795 B.n477 163.367
R1945 B.n803 B.n477 163.367
R1946 B.n803 B.n475 163.367
R1947 B.n807 B.n475 163.367
R1948 B.n807 B.n469 163.367
R1949 B.n816 B.n469 163.367
R1950 B.n816 B.n467 163.367
R1951 B.n820 B.n467 163.367
R1952 B.n820 B.n462 163.367
R1953 B.n828 B.n462 163.367
R1954 B.n828 B.n460 163.367
R1955 B.n832 B.n460 163.367
R1956 B.n832 B.n454 163.367
R1957 B.n840 B.n454 163.367
R1958 B.n840 B.n452 163.367
R1959 B.n844 B.n452 163.367
R1960 B.n844 B.n446 163.367
R1961 B.n852 B.n446 163.367
R1962 B.n852 B.n444 163.367
R1963 B.n856 B.n444 163.367
R1964 B.n856 B.n438 163.367
R1965 B.n864 B.n438 163.367
R1966 B.n864 B.n436 163.367
R1967 B.n868 B.n436 163.367
R1968 B.n868 B.n430 163.367
R1969 B.n876 B.n430 163.367
R1970 B.n876 B.n428 163.367
R1971 B.n880 B.n428 163.367
R1972 B.n880 B.n422 163.367
R1973 B.n888 B.n422 163.367
R1974 B.n888 B.n420 163.367
R1975 B.n892 B.n420 163.367
R1976 B.n892 B.n414 163.367
R1977 B.n900 B.n414 163.367
R1978 B.n900 B.n412 163.367
R1979 B.n904 B.n412 163.367
R1980 B.n904 B.n406 163.367
R1981 B.n912 B.n406 163.367
R1982 B.n912 B.n404 163.367
R1983 B.n916 B.n404 163.367
R1984 B.n916 B.n398 163.367
R1985 B.n924 B.n398 163.367
R1986 B.n924 B.n396 163.367
R1987 B.n928 B.n396 163.367
R1988 B.n928 B.n390 163.367
R1989 B.n936 B.n390 163.367
R1990 B.n936 B.n388 163.367
R1991 B.n940 B.n388 163.367
R1992 B.n940 B.n382 163.367
R1993 B.n949 B.n382 163.367
R1994 B.n949 B.n380 163.367
R1995 B.n953 B.n380 163.367
R1996 B.n953 B.n375 163.367
R1997 B.n962 B.n375 163.367
R1998 B.n962 B.n373 163.367
R1999 B.n966 B.n373 163.367
R2000 B.n966 B.n3 163.367
R2001 B.n1215 B.n3 163.367
R2002 B.n1211 B.n2 163.367
R2003 B.n1211 B.n1210 163.367
R2004 B.n1210 B.n9 163.367
R2005 B.n1206 B.n9 163.367
R2006 B.n1206 B.n11 163.367
R2007 B.n1202 B.n11 163.367
R2008 B.n1202 B.n16 163.367
R2009 B.n1198 B.n16 163.367
R2010 B.n1198 B.n18 163.367
R2011 B.n1194 B.n18 163.367
R2012 B.n1194 B.n24 163.367
R2013 B.n1190 B.n24 163.367
R2014 B.n1190 B.n26 163.367
R2015 B.n1186 B.n26 163.367
R2016 B.n1186 B.n31 163.367
R2017 B.n1182 B.n31 163.367
R2018 B.n1182 B.n33 163.367
R2019 B.n1178 B.n33 163.367
R2020 B.n1178 B.n38 163.367
R2021 B.n1174 B.n38 163.367
R2022 B.n1174 B.n40 163.367
R2023 B.n1170 B.n40 163.367
R2024 B.n1170 B.n45 163.367
R2025 B.n1166 B.n45 163.367
R2026 B.n1166 B.n47 163.367
R2027 B.n1162 B.n47 163.367
R2028 B.n1162 B.n52 163.367
R2029 B.n1158 B.n52 163.367
R2030 B.n1158 B.n54 163.367
R2031 B.n1154 B.n54 163.367
R2032 B.n1154 B.n59 163.367
R2033 B.n1150 B.n59 163.367
R2034 B.n1150 B.n61 163.367
R2035 B.n1146 B.n61 163.367
R2036 B.n1146 B.n66 163.367
R2037 B.n1142 B.n66 163.367
R2038 B.n1142 B.n68 163.367
R2039 B.n1138 B.n68 163.367
R2040 B.n1138 B.n73 163.367
R2041 B.n1134 B.n73 163.367
R2042 B.n1134 B.n75 163.367
R2043 B.n1130 B.n75 163.367
R2044 B.n1130 B.n80 163.367
R2045 B.n1126 B.n80 163.367
R2046 B.n1126 B.n82 163.367
R2047 B.n1122 B.n82 163.367
R2048 B.n1122 B.n87 163.367
R2049 B.n1118 B.n87 163.367
R2050 B.n1118 B.n89 163.367
R2051 B.n1114 B.n89 163.367
R2052 B.n1114 B.n93 163.367
R2053 B.n1110 B.n93 163.367
R2054 B.n1110 B.n95 163.367
R2055 B.n1106 B.n95 163.367
R2056 B.n1106 B.n101 163.367
R2057 B.n1102 B.n101 163.367
R2058 B.n1102 B.n103 163.367
R2059 B.n1098 B.n103 163.367
R2060 B.n1098 B.n108 163.367
R2061 B.n1094 B.n108 163.367
R2062 B.n1094 B.n110 163.367
R2063 B.n1090 B.n110 163.367
R2064 B.n1090 B.n115 163.367
R2065 B.n1086 B.n115 163.367
R2066 B.n1086 B.n117 163.367
R2067 B.n1082 B.n117 163.367
R2068 B.n1082 B.n122 163.367
R2069 B.n1078 B.n122 163.367
R2070 B.n1078 B.n124 163.367
R2071 B.n1074 B.n124 163.367
R2072 B.n1074 B.n129 163.367
R2073 B.n1070 B.n129 163.367
R2074 B.n1070 B.n131 163.367
R2075 B.n747 B.n510 74.5012
R2076 B.n1068 B.n1067 74.5012
R2077 B.n184 B.n183 71.7581
R2078 B.n182 B.n181 71.7581
R2079 B.n563 B.n562 71.7581
R2080 B.n561 B.n560 71.7581
R2081 B.n186 B.n134 71.676
R2082 B.n190 B.n135 71.676
R2083 B.n194 B.n136 71.676
R2084 B.n198 B.n137 71.676
R2085 B.n202 B.n138 71.676
R2086 B.n206 B.n139 71.676
R2087 B.n210 B.n140 71.676
R2088 B.n214 B.n141 71.676
R2089 B.n218 B.n142 71.676
R2090 B.n222 B.n143 71.676
R2091 B.n226 B.n144 71.676
R2092 B.n230 B.n145 71.676
R2093 B.n234 B.n146 71.676
R2094 B.n238 B.n147 71.676
R2095 B.n242 B.n148 71.676
R2096 B.n246 B.n149 71.676
R2097 B.n250 B.n150 71.676
R2098 B.n254 B.n151 71.676
R2099 B.n258 B.n152 71.676
R2100 B.n262 B.n153 71.676
R2101 B.n266 B.n154 71.676
R2102 B.n270 B.n155 71.676
R2103 B.n274 B.n156 71.676
R2104 B.n278 B.n157 71.676
R2105 B.n282 B.n158 71.676
R2106 B.n286 B.n159 71.676
R2107 B.n291 B.n160 71.676
R2108 B.n295 B.n161 71.676
R2109 B.n299 B.n162 71.676
R2110 B.n303 B.n163 71.676
R2111 B.n307 B.n164 71.676
R2112 B.n311 B.n165 71.676
R2113 B.n315 B.n166 71.676
R2114 B.n319 B.n167 71.676
R2115 B.n323 B.n168 71.676
R2116 B.n327 B.n169 71.676
R2117 B.n331 B.n170 71.676
R2118 B.n335 B.n171 71.676
R2119 B.n339 B.n172 71.676
R2120 B.n343 B.n173 71.676
R2121 B.n347 B.n174 71.676
R2122 B.n351 B.n175 71.676
R2123 B.n355 B.n176 71.676
R2124 B.n359 B.n177 71.676
R2125 B.n363 B.n178 71.676
R2126 B.n367 B.n179 71.676
R2127 B.n180 B.n179 71.676
R2128 B.n366 B.n178 71.676
R2129 B.n362 B.n177 71.676
R2130 B.n358 B.n176 71.676
R2131 B.n354 B.n175 71.676
R2132 B.n350 B.n174 71.676
R2133 B.n346 B.n173 71.676
R2134 B.n342 B.n172 71.676
R2135 B.n338 B.n171 71.676
R2136 B.n334 B.n170 71.676
R2137 B.n330 B.n169 71.676
R2138 B.n326 B.n168 71.676
R2139 B.n322 B.n167 71.676
R2140 B.n318 B.n166 71.676
R2141 B.n314 B.n165 71.676
R2142 B.n310 B.n164 71.676
R2143 B.n306 B.n163 71.676
R2144 B.n302 B.n162 71.676
R2145 B.n298 B.n161 71.676
R2146 B.n294 B.n160 71.676
R2147 B.n290 B.n159 71.676
R2148 B.n285 B.n158 71.676
R2149 B.n281 B.n157 71.676
R2150 B.n277 B.n156 71.676
R2151 B.n273 B.n155 71.676
R2152 B.n269 B.n154 71.676
R2153 B.n265 B.n153 71.676
R2154 B.n261 B.n152 71.676
R2155 B.n257 B.n151 71.676
R2156 B.n253 B.n150 71.676
R2157 B.n249 B.n149 71.676
R2158 B.n245 B.n148 71.676
R2159 B.n241 B.n147 71.676
R2160 B.n237 B.n146 71.676
R2161 B.n233 B.n145 71.676
R2162 B.n229 B.n144 71.676
R2163 B.n225 B.n143 71.676
R2164 B.n221 B.n142 71.676
R2165 B.n217 B.n141 71.676
R2166 B.n213 B.n140 71.676
R2167 B.n209 B.n139 71.676
R2168 B.n205 B.n138 71.676
R2169 B.n201 B.n137 71.676
R2170 B.n197 B.n136 71.676
R2171 B.n193 B.n135 71.676
R2172 B.n189 B.n134 71.676
R2173 B.n746 B.n745 71.676
R2174 B.n740 B.n514 71.676
R2175 B.n737 B.n515 71.676
R2176 B.n733 B.n516 71.676
R2177 B.n729 B.n517 71.676
R2178 B.n725 B.n518 71.676
R2179 B.n721 B.n519 71.676
R2180 B.n717 B.n520 71.676
R2181 B.n713 B.n521 71.676
R2182 B.n709 B.n522 71.676
R2183 B.n705 B.n523 71.676
R2184 B.n701 B.n524 71.676
R2185 B.n697 B.n525 71.676
R2186 B.n693 B.n526 71.676
R2187 B.n689 B.n527 71.676
R2188 B.n685 B.n528 71.676
R2189 B.n681 B.n529 71.676
R2190 B.n677 B.n530 71.676
R2191 B.n673 B.n531 71.676
R2192 B.n669 B.n532 71.676
R2193 B.n665 B.n533 71.676
R2194 B.n660 B.n534 71.676
R2195 B.n656 B.n535 71.676
R2196 B.n652 B.n536 71.676
R2197 B.n648 B.n537 71.676
R2198 B.n644 B.n538 71.676
R2199 B.n640 B.n539 71.676
R2200 B.n636 B.n540 71.676
R2201 B.n632 B.n541 71.676
R2202 B.n628 B.n542 71.676
R2203 B.n624 B.n543 71.676
R2204 B.n620 B.n544 71.676
R2205 B.n616 B.n545 71.676
R2206 B.n612 B.n546 71.676
R2207 B.n608 B.n547 71.676
R2208 B.n604 B.n548 71.676
R2209 B.n600 B.n549 71.676
R2210 B.n596 B.n550 71.676
R2211 B.n592 B.n551 71.676
R2212 B.n588 B.n552 71.676
R2213 B.n584 B.n553 71.676
R2214 B.n580 B.n554 71.676
R2215 B.n576 B.n555 71.676
R2216 B.n572 B.n556 71.676
R2217 B.n568 B.n557 71.676
R2218 B.n748 B.n513 71.676
R2219 B.n746 B.n559 71.676
R2220 B.n738 B.n514 71.676
R2221 B.n734 B.n515 71.676
R2222 B.n730 B.n516 71.676
R2223 B.n726 B.n517 71.676
R2224 B.n722 B.n518 71.676
R2225 B.n718 B.n519 71.676
R2226 B.n714 B.n520 71.676
R2227 B.n710 B.n521 71.676
R2228 B.n706 B.n522 71.676
R2229 B.n702 B.n523 71.676
R2230 B.n698 B.n524 71.676
R2231 B.n694 B.n525 71.676
R2232 B.n690 B.n526 71.676
R2233 B.n686 B.n527 71.676
R2234 B.n682 B.n528 71.676
R2235 B.n678 B.n529 71.676
R2236 B.n674 B.n530 71.676
R2237 B.n670 B.n531 71.676
R2238 B.n666 B.n532 71.676
R2239 B.n661 B.n533 71.676
R2240 B.n657 B.n534 71.676
R2241 B.n653 B.n535 71.676
R2242 B.n649 B.n536 71.676
R2243 B.n645 B.n537 71.676
R2244 B.n641 B.n538 71.676
R2245 B.n637 B.n539 71.676
R2246 B.n633 B.n540 71.676
R2247 B.n629 B.n541 71.676
R2248 B.n625 B.n542 71.676
R2249 B.n621 B.n543 71.676
R2250 B.n617 B.n544 71.676
R2251 B.n613 B.n545 71.676
R2252 B.n609 B.n546 71.676
R2253 B.n605 B.n547 71.676
R2254 B.n601 B.n548 71.676
R2255 B.n597 B.n549 71.676
R2256 B.n593 B.n550 71.676
R2257 B.n589 B.n551 71.676
R2258 B.n585 B.n552 71.676
R2259 B.n581 B.n553 71.676
R2260 B.n577 B.n554 71.676
R2261 B.n573 B.n555 71.676
R2262 B.n569 B.n556 71.676
R2263 B.n565 B.n557 71.676
R2264 B.n749 B.n748 71.676
R2265 B.n1216 B.n1215 71.676
R2266 B.n1216 B.n2 71.676
R2267 B.n185 B.n184 59.5399
R2268 B.n288 B.n182 59.5399
R2269 B.n564 B.n563 59.5399
R2270 B.n663 B.n561 59.5399
R2271 B.n754 B.n510 43.3001
R2272 B.n754 B.n506 43.3001
R2273 B.n760 B.n506 43.3001
R2274 B.n760 B.n502 43.3001
R2275 B.n766 B.n502 43.3001
R2276 B.n766 B.n497 43.3001
R2277 B.n772 B.n497 43.3001
R2278 B.n772 B.n498 43.3001
R2279 B.n778 B.n490 43.3001
R2280 B.n784 B.n490 43.3001
R2281 B.n784 B.n486 43.3001
R2282 B.n790 B.n486 43.3001
R2283 B.n790 B.n482 43.3001
R2284 B.n796 B.n482 43.3001
R2285 B.n796 B.n478 43.3001
R2286 B.n802 B.n478 43.3001
R2287 B.n802 B.n474 43.3001
R2288 B.n808 B.n474 43.3001
R2289 B.n808 B.n470 43.3001
R2290 B.n815 B.n470 43.3001
R2291 B.n815 B.n814 43.3001
R2292 B.n821 B.n463 43.3001
R2293 B.n827 B.n463 43.3001
R2294 B.n827 B.n459 43.3001
R2295 B.n833 B.n459 43.3001
R2296 B.n833 B.n455 43.3001
R2297 B.n839 B.n455 43.3001
R2298 B.n839 B.n451 43.3001
R2299 B.n845 B.n451 43.3001
R2300 B.n845 B.n447 43.3001
R2301 B.n851 B.n447 43.3001
R2302 B.n857 B.n443 43.3001
R2303 B.n857 B.n439 43.3001
R2304 B.n863 B.n439 43.3001
R2305 B.n863 B.n435 43.3001
R2306 B.n869 B.n435 43.3001
R2307 B.n869 B.n431 43.3001
R2308 B.n875 B.n431 43.3001
R2309 B.n875 B.n426 43.3001
R2310 B.n881 B.n426 43.3001
R2311 B.n881 B.n427 43.3001
R2312 B.n887 B.n419 43.3001
R2313 B.n893 B.n419 43.3001
R2314 B.n893 B.n415 43.3001
R2315 B.n899 B.n415 43.3001
R2316 B.n899 B.n411 43.3001
R2317 B.n905 B.n411 43.3001
R2318 B.n905 B.n407 43.3001
R2319 B.n911 B.n407 43.3001
R2320 B.n911 B.n403 43.3001
R2321 B.n917 B.n403 43.3001
R2322 B.n923 B.n399 43.3001
R2323 B.n923 B.n395 43.3001
R2324 B.n929 B.n395 43.3001
R2325 B.n929 B.n391 43.3001
R2326 B.n935 B.n391 43.3001
R2327 B.n935 B.n387 43.3001
R2328 B.n941 B.n387 43.3001
R2329 B.n941 B.n383 43.3001
R2330 B.n948 B.n383 43.3001
R2331 B.n948 B.n947 43.3001
R2332 B.n954 B.n376 43.3001
R2333 B.n961 B.n376 43.3001
R2334 B.n961 B.n372 43.3001
R2335 B.n967 B.n372 43.3001
R2336 B.n967 B.n4 43.3001
R2337 B.n1214 B.n4 43.3001
R2338 B.n1214 B.n1213 43.3001
R2339 B.n1213 B.n1212 43.3001
R2340 B.n1212 B.n8 43.3001
R2341 B.n12 B.n8 43.3001
R2342 B.n1205 B.n12 43.3001
R2343 B.n1205 B.n1204 43.3001
R2344 B.n1204 B.n1203 43.3001
R2345 B.n1197 B.n19 43.3001
R2346 B.n1197 B.n1196 43.3001
R2347 B.n1196 B.n1195 43.3001
R2348 B.n1195 B.n23 43.3001
R2349 B.n1189 B.n23 43.3001
R2350 B.n1189 B.n1188 43.3001
R2351 B.n1188 B.n1187 43.3001
R2352 B.n1187 B.n30 43.3001
R2353 B.n1181 B.n30 43.3001
R2354 B.n1181 B.n1180 43.3001
R2355 B.n1179 B.n37 43.3001
R2356 B.n1173 B.n37 43.3001
R2357 B.n1173 B.n1172 43.3001
R2358 B.n1172 B.n1171 43.3001
R2359 B.n1171 B.n44 43.3001
R2360 B.n1165 B.n44 43.3001
R2361 B.n1165 B.n1164 43.3001
R2362 B.n1164 B.n1163 43.3001
R2363 B.n1163 B.n51 43.3001
R2364 B.n1157 B.n51 43.3001
R2365 B.n1156 B.n1155 43.3001
R2366 B.n1155 B.n58 43.3001
R2367 B.n1149 B.n58 43.3001
R2368 B.n1149 B.n1148 43.3001
R2369 B.n1148 B.n1147 43.3001
R2370 B.n1147 B.n65 43.3001
R2371 B.n1141 B.n65 43.3001
R2372 B.n1141 B.n1140 43.3001
R2373 B.n1140 B.n1139 43.3001
R2374 B.n1139 B.n72 43.3001
R2375 B.n1133 B.n1132 43.3001
R2376 B.n1132 B.n1131 43.3001
R2377 B.n1131 B.n79 43.3001
R2378 B.n1125 B.n79 43.3001
R2379 B.n1125 B.n1124 43.3001
R2380 B.n1124 B.n1123 43.3001
R2381 B.n1123 B.n86 43.3001
R2382 B.n1117 B.n86 43.3001
R2383 B.n1117 B.n1116 43.3001
R2384 B.n1116 B.n1115 43.3001
R2385 B.n1109 B.n96 43.3001
R2386 B.n1109 B.n1108 43.3001
R2387 B.n1108 B.n1107 43.3001
R2388 B.n1107 B.n100 43.3001
R2389 B.n1101 B.n100 43.3001
R2390 B.n1101 B.n1100 43.3001
R2391 B.n1100 B.n1099 43.3001
R2392 B.n1099 B.n107 43.3001
R2393 B.n1093 B.n107 43.3001
R2394 B.n1093 B.n1092 43.3001
R2395 B.n1092 B.n1091 43.3001
R2396 B.n1091 B.n114 43.3001
R2397 B.n1085 B.n114 43.3001
R2398 B.n1084 B.n1083 43.3001
R2399 B.n1083 B.n121 43.3001
R2400 B.n1077 B.n121 43.3001
R2401 B.n1077 B.n1076 43.3001
R2402 B.n1076 B.n1075 43.3001
R2403 B.n1075 B.n128 43.3001
R2404 B.n1069 B.n128 43.3001
R2405 B.n1069 B.n1068 43.3001
R2406 B.n814 B.t1 40.1163
R2407 B.n96 B.t2 40.1163
R2408 B.n498 B.t11 36.2957
R2409 B.t15 B.n1084 36.2957
R2410 B.n851 B.t3 35.0222
R2411 B.n1133 B.t9 35.0222
R2412 B.n744 B.n508 30.4395
R2413 B.n751 B.n750 30.4395
R2414 B.n1065 B.n1064 30.4395
R2415 B.n187 B.n130 30.4395
R2416 B.n427 B.t7 29.9281
R2417 B.t6 B.n1156 29.9281
R2418 B.n917 B.t5 24.8341
R2419 B.t0 B.n1179 24.8341
R2420 B.n954 B.t8 23.5606
R2421 B.n1203 B.t4 23.5606
R2422 B.n947 B.t8 19.74
R2423 B.n19 B.t4 19.74
R2424 B.t5 B.n399 18.4665
R2425 B.n1180 B.t0 18.4665
R2426 B B.n1217 18.0485
R2427 B.n887 B.t7 13.3724
R2428 B.n1157 B.t6 13.3724
R2429 B.n756 B.n508 10.6151
R2430 B.n757 B.n756 10.6151
R2431 B.n758 B.n757 10.6151
R2432 B.n758 B.n500 10.6151
R2433 B.n768 B.n500 10.6151
R2434 B.n769 B.n768 10.6151
R2435 B.n770 B.n769 10.6151
R2436 B.n770 B.n492 10.6151
R2437 B.n780 B.n492 10.6151
R2438 B.n781 B.n780 10.6151
R2439 B.n782 B.n781 10.6151
R2440 B.n782 B.n484 10.6151
R2441 B.n792 B.n484 10.6151
R2442 B.n793 B.n792 10.6151
R2443 B.n794 B.n793 10.6151
R2444 B.n794 B.n476 10.6151
R2445 B.n804 B.n476 10.6151
R2446 B.n805 B.n804 10.6151
R2447 B.n806 B.n805 10.6151
R2448 B.n806 B.n468 10.6151
R2449 B.n817 B.n468 10.6151
R2450 B.n818 B.n817 10.6151
R2451 B.n819 B.n818 10.6151
R2452 B.n819 B.n461 10.6151
R2453 B.n829 B.n461 10.6151
R2454 B.n830 B.n829 10.6151
R2455 B.n831 B.n830 10.6151
R2456 B.n831 B.n453 10.6151
R2457 B.n841 B.n453 10.6151
R2458 B.n842 B.n841 10.6151
R2459 B.n843 B.n842 10.6151
R2460 B.n843 B.n445 10.6151
R2461 B.n853 B.n445 10.6151
R2462 B.n854 B.n853 10.6151
R2463 B.n855 B.n854 10.6151
R2464 B.n855 B.n437 10.6151
R2465 B.n865 B.n437 10.6151
R2466 B.n866 B.n865 10.6151
R2467 B.n867 B.n866 10.6151
R2468 B.n867 B.n429 10.6151
R2469 B.n877 B.n429 10.6151
R2470 B.n878 B.n877 10.6151
R2471 B.n879 B.n878 10.6151
R2472 B.n879 B.n421 10.6151
R2473 B.n889 B.n421 10.6151
R2474 B.n890 B.n889 10.6151
R2475 B.n891 B.n890 10.6151
R2476 B.n891 B.n413 10.6151
R2477 B.n901 B.n413 10.6151
R2478 B.n902 B.n901 10.6151
R2479 B.n903 B.n902 10.6151
R2480 B.n903 B.n405 10.6151
R2481 B.n913 B.n405 10.6151
R2482 B.n914 B.n913 10.6151
R2483 B.n915 B.n914 10.6151
R2484 B.n915 B.n397 10.6151
R2485 B.n925 B.n397 10.6151
R2486 B.n926 B.n925 10.6151
R2487 B.n927 B.n926 10.6151
R2488 B.n927 B.n389 10.6151
R2489 B.n937 B.n389 10.6151
R2490 B.n938 B.n937 10.6151
R2491 B.n939 B.n938 10.6151
R2492 B.n939 B.n381 10.6151
R2493 B.n950 B.n381 10.6151
R2494 B.n951 B.n950 10.6151
R2495 B.n952 B.n951 10.6151
R2496 B.n952 B.n374 10.6151
R2497 B.n963 B.n374 10.6151
R2498 B.n964 B.n963 10.6151
R2499 B.n965 B.n964 10.6151
R2500 B.n965 B.n0 10.6151
R2501 B.n744 B.n743 10.6151
R2502 B.n743 B.n742 10.6151
R2503 B.n742 B.n741 10.6151
R2504 B.n741 B.n739 10.6151
R2505 B.n739 B.n736 10.6151
R2506 B.n736 B.n735 10.6151
R2507 B.n735 B.n732 10.6151
R2508 B.n732 B.n731 10.6151
R2509 B.n731 B.n728 10.6151
R2510 B.n728 B.n727 10.6151
R2511 B.n727 B.n724 10.6151
R2512 B.n724 B.n723 10.6151
R2513 B.n723 B.n720 10.6151
R2514 B.n720 B.n719 10.6151
R2515 B.n719 B.n716 10.6151
R2516 B.n716 B.n715 10.6151
R2517 B.n715 B.n712 10.6151
R2518 B.n712 B.n711 10.6151
R2519 B.n711 B.n708 10.6151
R2520 B.n708 B.n707 10.6151
R2521 B.n707 B.n704 10.6151
R2522 B.n704 B.n703 10.6151
R2523 B.n703 B.n700 10.6151
R2524 B.n700 B.n699 10.6151
R2525 B.n699 B.n696 10.6151
R2526 B.n696 B.n695 10.6151
R2527 B.n695 B.n692 10.6151
R2528 B.n692 B.n691 10.6151
R2529 B.n691 B.n688 10.6151
R2530 B.n688 B.n687 10.6151
R2531 B.n687 B.n684 10.6151
R2532 B.n684 B.n683 10.6151
R2533 B.n683 B.n680 10.6151
R2534 B.n680 B.n679 10.6151
R2535 B.n679 B.n676 10.6151
R2536 B.n676 B.n675 10.6151
R2537 B.n675 B.n672 10.6151
R2538 B.n672 B.n671 10.6151
R2539 B.n671 B.n668 10.6151
R2540 B.n668 B.n667 10.6151
R2541 B.n667 B.n664 10.6151
R2542 B.n662 B.n659 10.6151
R2543 B.n659 B.n658 10.6151
R2544 B.n658 B.n655 10.6151
R2545 B.n655 B.n654 10.6151
R2546 B.n654 B.n651 10.6151
R2547 B.n651 B.n650 10.6151
R2548 B.n650 B.n647 10.6151
R2549 B.n647 B.n646 10.6151
R2550 B.n643 B.n642 10.6151
R2551 B.n642 B.n639 10.6151
R2552 B.n639 B.n638 10.6151
R2553 B.n638 B.n635 10.6151
R2554 B.n635 B.n634 10.6151
R2555 B.n634 B.n631 10.6151
R2556 B.n631 B.n630 10.6151
R2557 B.n630 B.n627 10.6151
R2558 B.n627 B.n626 10.6151
R2559 B.n626 B.n623 10.6151
R2560 B.n623 B.n622 10.6151
R2561 B.n622 B.n619 10.6151
R2562 B.n619 B.n618 10.6151
R2563 B.n618 B.n615 10.6151
R2564 B.n615 B.n614 10.6151
R2565 B.n614 B.n611 10.6151
R2566 B.n611 B.n610 10.6151
R2567 B.n610 B.n607 10.6151
R2568 B.n607 B.n606 10.6151
R2569 B.n606 B.n603 10.6151
R2570 B.n603 B.n602 10.6151
R2571 B.n602 B.n599 10.6151
R2572 B.n599 B.n598 10.6151
R2573 B.n598 B.n595 10.6151
R2574 B.n595 B.n594 10.6151
R2575 B.n594 B.n591 10.6151
R2576 B.n591 B.n590 10.6151
R2577 B.n590 B.n587 10.6151
R2578 B.n587 B.n586 10.6151
R2579 B.n586 B.n583 10.6151
R2580 B.n583 B.n582 10.6151
R2581 B.n582 B.n579 10.6151
R2582 B.n579 B.n578 10.6151
R2583 B.n578 B.n575 10.6151
R2584 B.n575 B.n574 10.6151
R2585 B.n574 B.n571 10.6151
R2586 B.n571 B.n570 10.6151
R2587 B.n570 B.n567 10.6151
R2588 B.n567 B.n566 10.6151
R2589 B.n566 B.n512 10.6151
R2590 B.n750 B.n512 10.6151
R2591 B.n752 B.n751 10.6151
R2592 B.n752 B.n504 10.6151
R2593 B.n762 B.n504 10.6151
R2594 B.n763 B.n762 10.6151
R2595 B.n764 B.n763 10.6151
R2596 B.n764 B.n495 10.6151
R2597 B.n774 B.n495 10.6151
R2598 B.n775 B.n774 10.6151
R2599 B.n776 B.n775 10.6151
R2600 B.n776 B.n488 10.6151
R2601 B.n786 B.n488 10.6151
R2602 B.n787 B.n786 10.6151
R2603 B.n788 B.n787 10.6151
R2604 B.n788 B.n480 10.6151
R2605 B.n798 B.n480 10.6151
R2606 B.n799 B.n798 10.6151
R2607 B.n800 B.n799 10.6151
R2608 B.n800 B.n472 10.6151
R2609 B.n810 B.n472 10.6151
R2610 B.n811 B.n810 10.6151
R2611 B.n812 B.n811 10.6151
R2612 B.n812 B.n465 10.6151
R2613 B.n823 B.n465 10.6151
R2614 B.n824 B.n823 10.6151
R2615 B.n825 B.n824 10.6151
R2616 B.n825 B.n457 10.6151
R2617 B.n835 B.n457 10.6151
R2618 B.n836 B.n835 10.6151
R2619 B.n837 B.n836 10.6151
R2620 B.n837 B.n449 10.6151
R2621 B.n847 B.n449 10.6151
R2622 B.n848 B.n847 10.6151
R2623 B.n849 B.n848 10.6151
R2624 B.n849 B.n441 10.6151
R2625 B.n859 B.n441 10.6151
R2626 B.n860 B.n859 10.6151
R2627 B.n861 B.n860 10.6151
R2628 B.n861 B.n433 10.6151
R2629 B.n871 B.n433 10.6151
R2630 B.n872 B.n871 10.6151
R2631 B.n873 B.n872 10.6151
R2632 B.n873 B.n424 10.6151
R2633 B.n883 B.n424 10.6151
R2634 B.n884 B.n883 10.6151
R2635 B.n885 B.n884 10.6151
R2636 B.n885 B.n417 10.6151
R2637 B.n895 B.n417 10.6151
R2638 B.n896 B.n895 10.6151
R2639 B.n897 B.n896 10.6151
R2640 B.n897 B.n409 10.6151
R2641 B.n907 B.n409 10.6151
R2642 B.n908 B.n907 10.6151
R2643 B.n909 B.n908 10.6151
R2644 B.n909 B.n401 10.6151
R2645 B.n919 B.n401 10.6151
R2646 B.n920 B.n919 10.6151
R2647 B.n921 B.n920 10.6151
R2648 B.n921 B.n393 10.6151
R2649 B.n931 B.n393 10.6151
R2650 B.n932 B.n931 10.6151
R2651 B.n933 B.n932 10.6151
R2652 B.n933 B.n385 10.6151
R2653 B.n943 B.n385 10.6151
R2654 B.n944 B.n943 10.6151
R2655 B.n945 B.n944 10.6151
R2656 B.n945 B.n378 10.6151
R2657 B.n956 B.n378 10.6151
R2658 B.n957 B.n956 10.6151
R2659 B.n959 B.n957 10.6151
R2660 B.n959 B.n958 10.6151
R2661 B.n958 B.n370 10.6151
R2662 B.n970 B.n370 10.6151
R2663 B.n971 B.n970 10.6151
R2664 B.n972 B.n971 10.6151
R2665 B.n973 B.n972 10.6151
R2666 B.n974 B.n973 10.6151
R2667 B.n977 B.n974 10.6151
R2668 B.n978 B.n977 10.6151
R2669 B.n979 B.n978 10.6151
R2670 B.n980 B.n979 10.6151
R2671 B.n982 B.n980 10.6151
R2672 B.n983 B.n982 10.6151
R2673 B.n984 B.n983 10.6151
R2674 B.n985 B.n984 10.6151
R2675 B.n987 B.n985 10.6151
R2676 B.n988 B.n987 10.6151
R2677 B.n989 B.n988 10.6151
R2678 B.n990 B.n989 10.6151
R2679 B.n992 B.n990 10.6151
R2680 B.n993 B.n992 10.6151
R2681 B.n994 B.n993 10.6151
R2682 B.n995 B.n994 10.6151
R2683 B.n997 B.n995 10.6151
R2684 B.n998 B.n997 10.6151
R2685 B.n999 B.n998 10.6151
R2686 B.n1000 B.n999 10.6151
R2687 B.n1002 B.n1000 10.6151
R2688 B.n1003 B.n1002 10.6151
R2689 B.n1004 B.n1003 10.6151
R2690 B.n1005 B.n1004 10.6151
R2691 B.n1007 B.n1005 10.6151
R2692 B.n1008 B.n1007 10.6151
R2693 B.n1009 B.n1008 10.6151
R2694 B.n1010 B.n1009 10.6151
R2695 B.n1012 B.n1010 10.6151
R2696 B.n1013 B.n1012 10.6151
R2697 B.n1014 B.n1013 10.6151
R2698 B.n1015 B.n1014 10.6151
R2699 B.n1017 B.n1015 10.6151
R2700 B.n1018 B.n1017 10.6151
R2701 B.n1019 B.n1018 10.6151
R2702 B.n1020 B.n1019 10.6151
R2703 B.n1022 B.n1020 10.6151
R2704 B.n1023 B.n1022 10.6151
R2705 B.n1024 B.n1023 10.6151
R2706 B.n1025 B.n1024 10.6151
R2707 B.n1027 B.n1025 10.6151
R2708 B.n1028 B.n1027 10.6151
R2709 B.n1029 B.n1028 10.6151
R2710 B.n1030 B.n1029 10.6151
R2711 B.n1032 B.n1030 10.6151
R2712 B.n1033 B.n1032 10.6151
R2713 B.n1034 B.n1033 10.6151
R2714 B.n1035 B.n1034 10.6151
R2715 B.n1037 B.n1035 10.6151
R2716 B.n1038 B.n1037 10.6151
R2717 B.n1039 B.n1038 10.6151
R2718 B.n1040 B.n1039 10.6151
R2719 B.n1042 B.n1040 10.6151
R2720 B.n1043 B.n1042 10.6151
R2721 B.n1044 B.n1043 10.6151
R2722 B.n1045 B.n1044 10.6151
R2723 B.n1047 B.n1045 10.6151
R2724 B.n1048 B.n1047 10.6151
R2725 B.n1049 B.n1048 10.6151
R2726 B.n1050 B.n1049 10.6151
R2727 B.n1052 B.n1050 10.6151
R2728 B.n1053 B.n1052 10.6151
R2729 B.n1054 B.n1053 10.6151
R2730 B.n1055 B.n1054 10.6151
R2731 B.n1057 B.n1055 10.6151
R2732 B.n1058 B.n1057 10.6151
R2733 B.n1059 B.n1058 10.6151
R2734 B.n1060 B.n1059 10.6151
R2735 B.n1062 B.n1060 10.6151
R2736 B.n1063 B.n1062 10.6151
R2737 B.n1064 B.n1063 10.6151
R2738 B.n1209 B.n1 10.6151
R2739 B.n1209 B.n1208 10.6151
R2740 B.n1208 B.n1207 10.6151
R2741 B.n1207 B.n10 10.6151
R2742 B.n1201 B.n10 10.6151
R2743 B.n1201 B.n1200 10.6151
R2744 B.n1200 B.n1199 10.6151
R2745 B.n1199 B.n17 10.6151
R2746 B.n1193 B.n17 10.6151
R2747 B.n1193 B.n1192 10.6151
R2748 B.n1192 B.n1191 10.6151
R2749 B.n1191 B.n25 10.6151
R2750 B.n1185 B.n25 10.6151
R2751 B.n1185 B.n1184 10.6151
R2752 B.n1184 B.n1183 10.6151
R2753 B.n1183 B.n32 10.6151
R2754 B.n1177 B.n32 10.6151
R2755 B.n1177 B.n1176 10.6151
R2756 B.n1176 B.n1175 10.6151
R2757 B.n1175 B.n39 10.6151
R2758 B.n1169 B.n39 10.6151
R2759 B.n1169 B.n1168 10.6151
R2760 B.n1168 B.n1167 10.6151
R2761 B.n1167 B.n46 10.6151
R2762 B.n1161 B.n46 10.6151
R2763 B.n1161 B.n1160 10.6151
R2764 B.n1160 B.n1159 10.6151
R2765 B.n1159 B.n53 10.6151
R2766 B.n1153 B.n53 10.6151
R2767 B.n1153 B.n1152 10.6151
R2768 B.n1152 B.n1151 10.6151
R2769 B.n1151 B.n60 10.6151
R2770 B.n1145 B.n60 10.6151
R2771 B.n1145 B.n1144 10.6151
R2772 B.n1144 B.n1143 10.6151
R2773 B.n1143 B.n67 10.6151
R2774 B.n1137 B.n67 10.6151
R2775 B.n1137 B.n1136 10.6151
R2776 B.n1136 B.n1135 10.6151
R2777 B.n1135 B.n74 10.6151
R2778 B.n1129 B.n74 10.6151
R2779 B.n1129 B.n1128 10.6151
R2780 B.n1128 B.n1127 10.6151
R2781 B.n1127 B.n81 10.6151
R2782 B.n1121 B.n81 10.6151
R2783 B.n1121 B.n1120 10.6151
R2784 B.n1120 B.n1119 10.6151
R2785 B.n1119 B.n88 10.6151
R2786 B.n1113 B.n88 10.6151
R2787 B.n1113 B.n1112 10.6151
R2788 B.n1112 B.n1111 10.6151
R2789 B.n1111 B.n94 10.6151
R2790 B.n1105 B.n94 10.6151
R2791 B.n1105 B.n1104 10.6151
R2792 B.n1104 B.n1103 10.6151
R2793 B.n1103 B.n102 10.6151
R2794 B.n1097 B.n102 10.6151
R2795 B.n1097 B.n1096 10.6151
R2796 B.n1096 B.n1095 10.6151
R2797 B.n1095 B.n109 10.6151
R2798 B.n1089 B.n109 10.6151
R2799 B.n1089 B.n1088 10.6151
R2800 B.n1088 B.n1087 10.6151
R2801 B.n1087 B.n116 10.6151
R2802 B.n1081 B.n116 10.6151
R2803 B.n1081 B.n1080 10.6151
R2804 B.n1080 B.n1079 10.6151
R2805 B.n1079 B.n123 10.6151
R2806 B.n1073 B.n123 10.6151
R2807 B.n1073 B.n1072 10.6151
R2808 B.n1072 B.n1071 10.6151
R2809 B.n1071 B.n130 10.6151
R2810 B.n188 B.n187 10.6151
R2811 B.n191 B.n188 10.6151
R2812 B.n192 B.n191 10.6151
R2813 B.n195 B.n192 10.6151
R2814 B.n196 B.n195 10.6151
R2815 B.n199 B.n196 10.6151
R2816 B.n200 B.n199 10.6151
R2817 B.n203 B.n200 10.6151
R2818 B.n204 B.n203 10.6151
R2819 B.n207 B.n204 10.6151
R2820 B.n208 B.n207 10.6151
R2821 B.n211 B.n208 10.6151
R2822 B.n212 B.n211 10.6151
R2823 B.n215 B.n212 10.6151
R2824 B.n216 B.n215 10.6151
R2825 B.n219 B.n216 10.6151
R2826 B.n220 B.n219 10.6151
R2827 B.n223 B.n220 10.6151
R2828 B.n224 B.n223 10.6151
R2829 B.n227 B.n224 10.6151
R2830 B.n228 B.n227 10.6151
R2831 B.n231 B.n228 10.6151
R2832 B.n232 B.n231 10.6151
R2833 B.n235 B.n232 10.6151
R2834 B.n236 B.n235 10.6151
R2835 B.n239 B.n236 10.6151
R2836 B.n240 B.n239 10.6151
R2837 B.n243 B.n240 10.6151
R2838 B.n244 B.n243 10.6151
R2839 B.n247 B.n244 10.6151
R2840 B.n248 B.n247 10.6151
R2841 B.n251 B.n248 10.6151
R2842 B.n252 B.n251 10.6151
R2843 B.n255 B.n252 10.6151
R2844 B.n256 B.n255 10.6151
R2845 B.n259 B.n256 10.6151
R2846 B.n260 B.n259 10.6151
R2847 B.n263 B.n260 10.6151
R2848 B.n264 B.n263 10.6151
R2849 B.n267 B.n264 10.6151
R2850 B.n268 B.n267 10.6151
R2851 B.n272 B.n271 10.6151
R2852 B.n275 B.n272 10.6151
R2853 B.n276 B.n275 10.6151
R2854 B.n279 B.n276 10.6151
R2855 B.n280 B.n279 10.6151
R2856 B.n283 B.n280 10.6151
R2857 B.n284 B.n283 10.6151
R2858 B.n287 B.n284 10.6151
R2859 B.n292 B.n289 10.6151
R2860 B.n293 B.n292 10.6151
R2861 B.n296 B.n293 10.6151
R2862 B.n297 B.n296 10.6151
R2863 B.n300 B.n297 10.6151
R2864 B.n301 B.n300 10.6151
R2865 B.n304 B.n301 10.6151
R2866 B.n305 B.n304 10.6151
R2867 B.n308 B.n305 10.6151
R2868 B.n309 B.n308 10.6151
R2869 B.n312 B.n309 10.6151
R2870 B.n313 B.n312 10.6151
R2871 B.n316 B.n313 10.6151
R2872 B.n317 B.n316 10.6151
R2873 B.n320 B.n317 10.6151
R2874 B.n321 B.n320 10.6151
R2875 B.n324 B.n321 10.6151
R2876 B.n325 B.n324 10.6151
R2877 B.n328 B.n325 10.6151
R2878 B.n329 B.n328 10.6151
R2879 B.n332 B.n329 10.6151
R2880 B.n333 B.n332 10.6151
R2881 B.n336 B.n333 10.6151
R2882 B.n337 B.n336 10.6151
R2883 B.n340 B.n337 10.6151
R2884 B.n341 B.n340 10.6151
R2885 B.n344 B.n341 10.6151
R2886 B.n345 B.n344 10.6151
R2887 B.n348 B.n345 10.6151
R2888 B.n349 B.n348 10.6151
R2889 B.n352 B.n349 10.6151
R2890 B.n353 B.n352 10.6151
R2891 B.n356 B.n353 10.6151
R2892 B.n357 B.n356 10.6151
R2893 B.n360 B.n357 10.6151
R2894 B.n361 B.n360 10.6151
R2895 B.n364 B.n361 10.6151
R2896 B.n365 B.n364 10.6151
R2897 B.n368 B.n365 10.6151
R2898 B.n369 B.n368 10.6151
R2899 B.n1065 B.n369 10.6151
R2900 B.t3 B.n443 8.27836
R2901 B.t9 B.n72 8.27836
R2902 B.n1217 B.n0 8.11757
R2903 B.n1217 B.n1 8.11757
R2904 B.n778 B.t11 7.00484
R2905 B.n1085 B.t15 7.00484
R2906 B.n663 B.n662 6.5566
R2907 B.n646 B.n564 6.5566
R2908 B.n271 B.n185 6.5566
R2909 B.n288 B.n287 6.5566
R2910 B.n664 B.n663 4.05904
R2911 B.n643 B.n564 4.05904
R2912 B.n268 B.n185 4.05904
R2913 B.n289 B.n288 4.05904
R2914 B.n821 B.t1 3.18429
R2915 B.n1115 B.t2 3.18429
R2916 VP.n32 VP.n31 161.3
R2917 VP.n33 VP.n28 161.3
R2918 VP.n35 VP.n34 161.3
R2919 VP.n36 VP.n27 161.3
R2920 VP.n38 VP.n37 161.3
R2921 VP.n39 VP.n26 161.3
R2922 VP.n41 VP.n40 161.3
R2923 VP.n43 VP.n42 161.3
R2924 VP.n44 VP.n24 161.3
R2925 VP.n46 VP.n45 161.3
R2926 VP.n47 VP.n23 161.3
R2927 VP.n49 VP.n48 161.3
R2928 VP.n50 VP.n22 161.3
R2929 VP.n53 VP.n52 161.3
R2930 VP.n54 VP.n21 161.3
R2931 VP.n56 VP.n55 161.3
R2932 VP.n57 VP.n20 161.3
R2933 VP.n59 VP.n58 161.3
R2934 VP.n60 VP.n19 161.3
R2935 VP.n62 VP.n61 161.3
R2936 VP.n63 VP.n18 161.3
R2937 VP.n65 VP.n64 161.3
R2938 VP.n115 VP.n114 161.3
R2939 VP.n113 VP.n1 161.3
R2940 VP.n112 VP.n111 161.3
R2941 VP.n110 VP.n2 161.3
R2942 VP.n109 VP.n108 161.3
R2943 VP.n107 VP.n3 161.3
R2944 VP.n106 VP.n105 161.3
R2945 VP.n104 VP.n4 161.3
R2946 VP.n103 VP.n102 161.3
R2947 VP.n100 VP.n5 161.3
R2948 VP.n99 VP.n98 161.3
R2949 VP.n97 VP.n6 161.3
R2950 VP.n96 VP.n95 161.3
R2951 VP.n94 VP.n7 161.3
R2952 VP.n93 VP.n92 161.3
R2953 VP.n91 VP.n90 161.3
R2954 VP.n89 VP.n9 161.3
R2955 VP.n88 VP.n87 161.3
R2956 VP.n86 VP.n10 161.3
R2957 VP.n85 VP.n84 161.3
R2958 VP.n83 VP.n11 161.3
R2959 VP.n82 VP.n81 161.3
R2960 VP.n80 VP.n79 161.3
R2961 VP.n78 VP.n13 161.3
R2962 VP.n77 VP.n76 161.3
R2963 VP.n75 VP.n14 161.3
R2964 VP.n74 VP.n73 161.3
R2965 VP.n72 VP.n15 161.3
R2966 VP.n71 VP.n70 161.3
R2967 VP.n69 VP.n16 161.3
R2968 VP.n30 VP.t9 118.828
R2969 VP.n67 VP.t6 85.8165
R2970 VP.n12 VP.t0 85.8165
R2971 VP.n8 VP.t7 85.8165
R2972 VP.n101 VP.t3 85.8165
R2973 VP.n0 VP.t8 85.8165
R2974 VP.n17 VP.t1 85.8165
R2975 VP.n51 VP.t2 85.8165
R2976 VP.n25 VP.t4 85.8165
R2977 VP.n29 VP.t5 85.8165
R2978 VP.n68 VP.n67 82.868
R2979 VP.n116 VP.n0 82.868
R2980 VP.n66 VP.n17 82.868
R2981 VP.n68 VP.n66 57.3177
R2982 VP.n73 VP.n14 56.5617
R2983 VP.n108 VP.n2 56.5617
R2984 VP.n58 VP.n19 56.5617
R2985 VP.n30 VP.n29 52.6179
R2986 VP.n84 VP.n10 50.2647
R2987 VP.n99 VP.n6 50.2647
R2988 VP.n49 VP.n23 50.2647
R2989 VP.n34 VP.n27 50.2647
R2990 VP.n88 VP.n10 30.8893
R2991 VP.n95 VP.n6 30.8893
R2992 VP.n45 VP.n23 30.8893
R2993 VP.n38 VP.n27 30.8893
R2994 VP.n71 VP.n16 24.5923
R2995 VP.n72 VP.n71 24.5923
R2996 VP.n73 VP.n72 24.5923
R2997 VP.n77 VP.n14 24.5923
R2998 VP.n78 VP.n77 24.5923
R2999 VP.n79 VP.n78 24.5923
R3000 VP.n83 VP.n82 24.5923
R3001 VP.n84 VP.n83 24.5923
R3002 VP.n89 VP.n88 24.5923
R3003 VP.n90 VP.n89 24.5923
R3004 VP.n94 VP.n93 24.5923
R3005 VP.n95 VP.n94 24.5923
R3006 VP.n100 VP.n99 24.5923
R3007 VP.n102 VP.n100 24.5923
R3008 VP.n106 VP.n4 24.5923
R3009 VP.n107 VP.n106 24.5923
R3010 VP.n108 VP.n107 24.5923
R3011 VP.n112 VP.n2 24.5923
R3012 VP.n113 VP.n112 24.5923
R3013 VP.n114 VP.n113 24.5923
R3014 VP.n62 VP.n19 24.5923
R3015 VP.n63 VP.n62 24.5923
R3016 VP.n64 VP.n63 24.5923
R3017 VP.n50 VP.n49 24.5923
R3018 VP.n52 VP.n50 24.5923
R3019 VP.n56 VP.n21 24.5923
R3020 VP.n57 VP.n56 24.5923
R3021 VP.n58 VP.n57 24.5923
R3022 VP.n39 VP.n38 24.5923
R3023 VP.n40 VP.n39 24.5923
R3024 VP.n44 VP.n43 24.5923
R3025 VP.n45 VP.n44 24.5923
R3026 VP.n33 VP.n32 24.5923
R3027 VP.n34 VP.n33 24.5923
R3028 VP.n82 VP.n12 22.1332
R3029 VP.n102 VP.n101 22.1332
R3030 VP.n52 VP.n51 22.1332
R3031 VP.n32 VP.n29 22.1332
R3032 VP.n90 VP.n8 12.2964
R3033 VP.n93 VP.n8 12.2964
R3034 VP.n40 VP.n25 12.2964
R3035 VP.n43 VP.n25 12.2964
R3036 VP.n67 VP.n16 7.37805
R3037 VP.n114 VP.n0 7.37805
R3038 VP.n64 VP.n17 7.37805
R3039 VP.n31 VP.n30 3.2308
R3040 VP.n79 VP.n12 2.45968
R3041 VP.n101 VP.n4 2.45968
R3042 VP.n51 VP.n21 2.45968
R3043 VP.n66 VP.n65 0.354861
R3044 VP.n69 VP.n68 0.354861
R3045 VP.n116 VP.n115 0.354861
R3046 VP VP.n116 0.267071
R3047 VP.n31 VP.n28 0.189894
R3048 VP.n35 VP.n28 0.189894
R3049 VP.n36 VP.n35 0.189894
R3050 VP.n37 VP.n36 0.189894
R3051 VP.n37 VP.n26 0.189894
R3052 VP.n41 VP.n26 0.189894
R3053 VP.n42 VP.n41 0.189894
R3054 VP.n42 VP.n24 0.189894
R3055 VP.n46 VP.n24 0.189894
R3056 VP.n47 VP.n46 0.189894
R3057 VP.n48 VP.n47 0.189894
R3058 VP.n48 VP.n22 0.189894
R3059 VP.n53 VP.n22 0.189894
R3060 VP.n54 VP.n53 0.189894
R3061 VP.n55 VP.n54 0.189894
R3062 VP.n55 VP.n20 0.189894
R3063 VP.n59 VP.n20 0.189894
R3064 VP.n60 VP.n59 0.189894
R3065 VP.n61 VP.n60 0.189894
R3066 VP.n61 VP.n18 0.189894
R3067 VP.n65 VP.n18 0.189894
R3068 VP.n70 VP.n69 0.189894
R3069 VP.n70 VP.n15 0.189894
R3070 VP.n74 VP.n15 0.189894
R3071 VP.n75 VP.n74 0.189894
R3072 VP.n76 VP.n75 0.189894
R3073 VP.n76 VP.n13 0.189894
R3074 VP.n80 VP.n13 0.189894
R3075 VP.n81 VP.n80 0.189894
R3076 VP.n81 VP.n11 0.189894
R3077 VP.n85 VP.n11 0.189894
R3078 VP.n86 VP.n85 0.189894
R3079 VP.n87 VP.n86 0.189894
R3080 VP.n87 VP.n9 0.189894
R3081 VP.n91 VP.n9 0.189894
R3082 VP.n92 VP.n91 0.189894
R3083 VP.n92 VP.n7 0.189894
R3084 VP.n96 VP.n7 0.189894
R3085 VP.n97 VP.n96 0.189894
R3086 VP.n98 VP.n97 0.189894
R3087 VP.n98 VP.n5 0.189894
R3088 VP.n103 VP.n5 0.189894
R3089 VP.n104 VP.n103 0.189894
R3090 VP.n105 VP.n104 0.189894
R3091 VP.n105 VP.n3 0.189894
R3092 VP.n109 VP.n3 0.189894
R3093 VP.n110 VP.n109 0.189894
R3094 VP.n111 VP.n110 0.189894
R3095 VP.n111 VP.n1 0.189894
R3096 VP.n115 VP.n1 0.189894
R3097 VDD1.n60 VDD1.n0 289.615
R3098 VDD1.n127 VDD1.n67 289.615
R3099 VDD1.n61 VDD1.n60 185
R3100 VDD1.n59 VDD1.n58 185
R3101 VDD1.n4 VDD1.n3 185
R3102 VDD1.n53 VDD1.n52 185
R3103 VDD1.n51 VDD1.n50 185
R3104 VDD1.n8 VDD1.n7 185
R3105 VDD1.n45 VDD1.n44 185
R3106 VDD1.n43 VDD1.n10 185
R3107 VDD1.n42 VDD1.n41 185
R3108 VDD1.n13 VDD1.n11 185
R3109 VDD1.n36 VDD1.n35 185
R3110 VDD1.n34 VDD1.n33 185
R3111 VDD1.n17 VDD1.n16 185
R3112 VDD1.n28 VDD1.n27 185
R3113 VDD1.n26 VDD1.n25 185
R3114 VDD1.n21 VDD1.n20 185
R3115 VDD1.n87 VDD1.n86 185
R3116 VDD1.n92 VDD1.n91 185
R3117 VDD1.n94 VDD1.n93 185
R3118 VDD1.n83 VDD1.n82 185
R3119 VDD1.n100 VDD1.n99 185
R3120 VDD1.n102 VDD1.n101 185
R3121 VDD1.n79 VDD1.n78 185
R3122 VDD1.n109 VDD1.n108 185
R3123 VDD1.n110 VDD1.n77 185
R3124 VDD1.n112 VDD1.n111 185
R3125 VDD1.n75 VDD1.n74 185
R3126 VDD1.n118 VDD1.n117 185
R3127 VDD1.n120 VDD1.n119 185
R3128 VDD1.n71 VDD1.n70 185
R3129 VDD1.n126 VDD1.n125 185
R3130 VDD1.n128 VDD1.n127 185
R3131 VDD1.n22 VDD1.t0 149.524
R3132 VDD1.n88 VDD1.t3 149.524
R3133 VDD1.n60 VDD1.n59 104.615
R3134 VDD1.n59 VDD1.n3 104.615
R3135 VDD1.n52 VDD1.n3 104.615
R3136 VDD1.n52 VDD1.n51 104.615
R3137 VDD1.n51 VDD1.n7 104.615
R3138 VDD1.n44 VDD1.n7 104.615
R3139 VDD1.n44 VDD1.n43 104.615
R3140 VDD1.n43 VDD1.n42 104.615
R3141 VDD1.n42 VDD1.n11 104.615
R3142 VDD1.n35 VDD1.n11 104.615
R3143 VDD1.n35 VDD1.n34 104.615
R3144 VDD1.n34 VDD1.n16 104.615
R3145 VDD1.n27 VDD1.n16 104.615
R3146 VDD1.n27 VDD1.n26 104.615
R3147 VDD1.n26 VDD1.n20 104.615
R3148 VDD1.n92 VDD1.n86 104.615
R3149 VDD1.n93 VDD1.n92 104.615
R3150 VDD1.n93 VDD1.n82 104.615
R3151 VDD1.n100 VDD1.n82 104.615
R3152 VDD1.n101 VDD1.n100 104.615
R3153 VDD1.n101 VDD1.n78 104.615
R3154 VDD1.n109 VDD1.n78 104.615
R3155 VDD1.n110 VDD1.n109 104.615
R3156 VDD1.n111 VDD1.n110 104.615
R3157 VDD1.n111 VDD1.n74 104.615
R3158 VDD1.n118 VDD1.n74 104.615
R3159 VDD1.n119 VDD1.n118 104.615
R3160 VDD1.n119 VDD1.n70 104.615
R3161 VDD1.n126 VDD1.n70 104.615
R3162 VDD1.n127 VDD1.n126 104.615
R3163 VDD1.n135 VDD1.n134 61.8894
R3164 VDD1.n66 VDD1.n65 59.5527
R3165 VDD1.n137 VDD1.n136 59.5525
R3166 VDD1.n133 VDD1.n132 59.5525
R3167 VDD1.t0 VDD1.n20 52.3082
R3168 VDD1.t3 VDD1.n86 52.3082
R3169 VDD1.n137 VDD1.n135 51.3888
R3170 VDD1.n66 VDD1.n64 49.7265
R3171 VDD1.n133 VDD1.n131 49.7265
R3172 VDD1.n45 VDD1.n10 13.1884
R3173 VDD1.n112 VDD1.n77 13.1884
R3174 VDD1.n46 VDD1.n8 12.8005
R3175 VDD1.n41 VDD1.n12 12.8005
R3176 VDD1.n108 VDD1.n107 12.8005
R3177 VDD1.n113 VDD1.n75 12.8005
R3178 VDD1.n50 VDD1.n49 12.0247
R3179 VDD1.n40 VDD1.n13 12.0247
R3180 VDD1.n106 VDD1.n79 12.0247
R3181 VDD1.n117 VDD1.n116 12.0247
R3182 VDD1.n53 VDD1.n6 11.249
R3183 VDD1.n37 VDD1.n36 11.249
R3184 VDD1.n103 VDD1.n102 11.249
R3185 VDD1.n120 VDD1.n73 11.249
R3186 VDD1.n54 VDD1.n4 10.4732
R3187 VDD1.n33 VDD1.n15 10.4732
R3188 VDD1.n99 VDD1.n81 10.4732
R3189 VDD1.n121 VDD1.n71 10.4732
R3190 VDD1.n22 VDD1.n21 10.2747
R3191 VDD1.n88 VDD1.n87 10.2747
R3192 VDD1.n58 VDD1.n57 9.69747
R3193 VDD1.n32 VDD1.n17 9.69747
R3194 VDD1.n98 VDD1.n83 9.69747
R3195 VDD1.n125 VDD1.n124 9.69747
R3196 VDD1.n64 VDD1.n63 9.45567
R3197 VDD1.n131 VDD1.n130 9.45567
R3198 VDD1.n24 VDD1.n23 9.3005
R3199 VDD1.n19 VDD1.n18 9.3005
R3200 VDD1.n30 VDD1.n29 9.3005
R3201 VDD1.n32 VDD1.n31 9.3005
R3202 VDD1.n15 VDD1.n14 9.3005
R3203 VDD1.n38 VDD1.n37 9.3005
R3204 VDD1.n40 VDD1.n39 9.3005
R3205 VDD1.n12 VDD1.n9 9.3005
R3206 VDD1.n63 VDD1.n62 9.3005
R3207 VDD1.n2 VDD1.n1 9.3005
R3208 VDD1.n57 VDD1.n56 9.3005
R3209 VDD1.n55 VDD1.n54 9.3005
R3210 VDD1.n6 VDD1.n5 9.3005
R3211 VDD1.n49 VDD1.n48 9.3005
R3212 VDD1.n47 VDD1.n46 9.3005
R3213 VDD1.n130 VDD1.n129 9.3005
R3214 VDD1.n69 VDD1.n68 9.3005
R3215 VDD1.n124 VDD1.n123 9.3005
R3216 VDD1.n122 VDD1.n121 9.3005
R3217 VDD1.n73 VDD1.n72 9.3005
R3218 VDD1.n116 VDD1.n115 9.3005
R3219 VDD1.n114 VDD1.n113 9.3005
R3220 VDD1.n90 VDD1.n89 9.3005
R3221 VDD1.n85 VDD1.n84 9.3005
R3222 VDD1.n96 VDD1.n95 9.3005
R3223 VDD1.n98 VDD1.n97 9.3005
R3224 VDD1.n81 VDD1.n80 9.3005
R3225 VDD1.n104 VDD1.n103 9.3005
R3226 VDD1.n106 VDD1.n105 9.3005
R3227 VDD1.n107 VDD1.n76 9.3005
R3228 VDD1.n61 VDD1.n2 8.92171
R3229 VDD1.n29 VDD1.n28 8.92171
R3230 VDD1.n95 VDD1.n94 8.92171
R3231 VDD1.n128 VDD1.n69 8.92171
R3232 VDD1.n62 VDD1.n0 8.14595
R3233 VDD1.n25 VDD1.n19 8.14595
R3234 VDD1.n91 VDD1.n85 8.14595
R3235 VDD1.n129 VDD1.n67 8.14595
R3236 VDD1.n24 VDD1.n21 7.3702
R3237 VDD1.n90 VDD1.n87 7.3702
R3238 VDD1.n64 VDD1.n0 5.81868
R3239 VDD1.n25 VDD1.n24 5.81868
R3240 VDD1.n91 VDD1.n90 5.81868
R3241 VDD1.n131 VDD1.n67 5.81868
R3242 VDD1.n62 VDD1.n61 5.04292
R3243 VDD1.n28 VDD1.n19 5.04292
R3244 VDD1.n94 VDD1.n85 5.04292
R3245 VDD1.n129 VDD1.n128 5.04292
R3246 VDD1.n58 VDD1.n2 4.26717
R3247 VDD1.n29 VDD1.n17 4.26717
R3248 VDD1.n95 VDD1.n83 4.26717
R3249 VDD1.n125 VDD1.n69 4.26717
R3250 VDD1.n57 VDD1.n4 3.49141
R3251 VDD1.n33 VDD1.n32 3.49141
R3252 VDD1.n99 VDD1.n98 3.49141
R3253 VDD1.n124 VDD1.n71 3.49141
R3254 VDD1.n23 VDD1.n22 2.84303
R3255 VDD1.n89 VDD1.n88 2.84303
R3256 VDD1.n54 VDD1.n53 2.71565
R3257 VDD1.n36 VDD1.n15 2.71565
R3258 VDD1.n102 VDD1.n81 2.71565
R3259 VDD1.n121 VDD1.n120 2.71565
R3260 VDD1 VDD1.n137 2.33455
R3261 VDD1.n50 VDD1.n6 1.93989
R3262 VDD1.n37 VDD1.n13 1.93989
R3263 VDD1.n103 VDD1.n79 1.93989
R3264 VDD1.n117 VDD1.n73 1.93989
R3265 VDD1.n136 VDD1.t7 1.6505
R3266 VDD1.n136 VDD1.t8 1.6505
R3267 VDD1.n65 VDD1.t4 1.6505
R3268 VDD1.n65 VDD1.t5 1.6505
R3269 VDD1.n134 VDD1.t6 1.6505
R3270 VDD1.n134 VDD1.t1 1.6505
R3271 VDD1.n132 VDD1.t9 1.6505
R3272 VDD1.n132 VDD1.t2 1.6505
R3273 VDD1.n49 VDD1.n8 1.16414
R3274 VDD1.n41 VDD1.n40 1.16414
R3275 VDD1.n108 VDD1.n106 1.16414
R3276 VDD1.n116 VDD1.n75 1.16414
R3277 VDD1 VDD1.n66 0.856103
R3278 VDD1.n135 VDD1.n133 0.742568
R3279 VDD1.n46 VDD1.n45 0.388379
R3280 VDD1.n12 VDD1.n10 0.388379
R3281 VDD1.n107 VDD1.n77 0.388379
R3282 VDD1.n113 VDD1.n112 0.388379
R3283 VDD1.n63 VDD1.n1 0.155672
R3284 VDD1.n56 VDD1.n1 0.155672
R3285 VDD1.n56 VDD1.n55 0.155672
R3286 VDD1.n55 VDD1.n5 0.155672
R3287 VDD1.n48 VDD1.n5 0.155672
R3288 VDD1.n48 VDD1.n47 0.155672
R3289 VDD1.n47 VDD1.n9 0.155672
R3290 VDD1.n39 VDD1.n9 0.155672
R3291 VDD1.n39 VDD1.n38 0.155672
R3292 VDD1.n38 VDD1.n14 0.155672
R3293 VDD1.n31 VDD1.n14 0.155672
R3294 VDD1.n31 VDD1.n30 0.155672
R3295 VDD1.n30 VDD1.n18 0.155672
R3296 VDD1.n23 VDD1.n18 0.155672
R3297 VDD1.n89 VDD1.n84 0.155672
R3298 VDD1.n96 VDD1.n84 0.155672
R3299 VDD1.n97 VDD1.n96 0.155672
R3300 VDD1.n97 VDD1.n80 0.155672
R3301 VDD1.n104 VDD1.n80 0.155672
R3302 VDD1.n105 VDD1.n104 0.155672
R3303 VDD1.n105 VDD1.n76 0.155672
R3304 VDD1.n114 VDD1.n76 0.155672
R3305 VDD1.n115 VDD1.n114 0.155672
R3306 VDD1.n115 VDD1.n72 0.155672
R3307 VDD1.n122 VDD1.n72 0.155672
R3308 VDD1.n123 VDD1.n122 0.155672
R3309 VDD1.n123 VDD1.n68 0.155672
R3310 VDD1.n130 VDD1.n68 0.155672
C0 VTAIL VP 12.157f
C1 VN VDD1 0.155502f
C2 VN VDD2 11.17f
C3 VTAIL VDD1 10.7207f
C4 VP VDD1 11.6928f
C5 VTAIL VDD2 10.7775f
C6 VP VDD2 0.682204f
C7 VDD1 VDD2 2.67631f
C8 VN VTAIL 12.1427f
C9 VN VP 9.53026f
C10 VDD2 B 8.116954f
C11 VDD1 B 8.080063f
C12 VTAIL B 8.79783f
C13 VN B 21.80971f
C14 VP B 20.387285f
C15 VDD1.n0 B 0.033119f
C16 VDD1.n1 B 0.025003f
C17 VDD1.n2 B 0.013435f
C18 VDD1.n3 B 0.031756f
C19 VDD1.n4 B 0.014226f
C20 VDD1.n5 B 0.025003f
C21 VDD1.n6 B 0.013435f
C22 VDD1.n7 B 0.031756f
C23 VDD1.n8 B 0.014226f
C24 VDD1.n9 B 0.025003f
C25 VDD1.n10 B 0.013831f
C26 VDD1.n11 B 0.031756f
C27 VDD1.n12 B 0.013435f
C28 VDD1.n13 B 0.014226f
C29 VDD1.n14 B 0.025003f
C30 VDD1.n15 B 0.013435f
C31 VDD1.n16 B 0.031756f
C32 VDD1.n17 B 0.014226f
C33 VDD1.n18 B 0.025003f
C34 VDD1.n19 B 0.013435f
C35 VDD1.n20 B 0.023817f
C36 VDD1.n21 B 0.022449f
C37 VDD1.t0 B 0.053634f
C38 VDD1.n22 B 0.180267f
C39 VDD1.n23 B 1.26135f
C40 VDD1.n24 B 0.013435f
C41 VDD1.n25 B 0.014226f
C42 VDD1.n26 B 0.031756f
C43 VDD1.n27 B 0.031756f
C44 VDD1.n28 B 0.014226f
C45 VDD1.n29 B 0.013435f
C46 VDD1.n30 B 0.025003f
C47 VDD1.n31 B 0.025003f
C48 VDD1.n32 B 0.013435f
C49 VDD1.n33 B 0.014226f
C50 VDD1.n34 B 0.031756f
C51 VDD1.n35 B 0.031756f
C52 VDD1.n36 B 0.014226f
C53 VDD1.n37 B 0.013435f
C54 VDD1.n38 B 0.025003f
C55 VDD1.n39 B 0.025003f
C56 VDD1.n40 B 0.013435f
C57 VDD1.n41 B 0.014226f
C58 VDD1.n42 B 0.031756f
C59 VDD1.n43 B 0.031756f
C60 VDD1.n44 B 0.031756f
C61 VDD1.n45 B 0.013831f
C62 VDD1.n46 B 0.013435f
C63 VDD1.n47 B 0.025003f
C64 VDD1.n48 B 0.025003f
C65 VDD1.n49 B 0.013435f
C66 VDD1.n50 B 0.014226f
C67 VDD1.n51 B 0.031756f
C68 VDD1.n52 B 0.031756f
C69 VDD1.n53 B 0.014226f
C70 VDD1.n54 B 0.013435f
C71 VDD1.n55 B 0.025003f
C72 VDD1.n56 B 0.025003f
C73 VDD1.n57 B 0.013435f
C74 VDD1.n58 B 0.014226f
C75 VDD1.n59 B 0.031756f
C76 VDD1.n60 B 0.065167f
C77 VDD1.n61 B 0.014226f
C78 VDD1.n62 B 0.013435f
C79 VDD1.n63 B 0.053694f
C80 VDD1.n64 B 0.072686f
C81 VDD1.t4 B 0.237095f
C82 VDD1.t5 B 0.237095f
C83 VDD1.n65 B 2.10979f
C84 VDD1.n66 B 0.819084f
C85 VDD1.n67 B 0.033119f
C86 VDD1.n68 B 0.025003f
C87 VDD1.n69 B 0.013435f
C88 VDD1.n70 B 0.031756f
C89 VDD1.n71 B 0.014226f
C90 VDD1.n72 B 0.025003f
C91 VDD1.n73 B 0.013435f
C92 VDD1.n74 B 0.031756f
C93 VDD1.n75 B 0.014226f
C94 VDD1.n76 B 0.025003f
C95 VDD1.n77 B 0.013831f
C96 VDD1.n78 B 0.031756f
C97 VDD1.n79 B 0.014226f
C98 VDD1.n80 B 0.025003f
C99 VDD1.n81 B 0.013435f
C100 VDD1.n82 B 0.031756f
C101 VDD1.n83 B 0.014226f
C102 VDD1.n84 B 0.025003f
C103 VDD1.n85 B 0.013435f
C104 VDD1.n86 B 0.023817f
C105 VDD1.n87 B 0.022449f
C106 VDD1.t3 B 0.053634f
C107 VDD1.n88 B 0.180267f
C108 VDD1.n89 B 1.26135f
C109 VDD1.n90 B 0.013435f
C110 VDD1.n91 B 0.014226f
C111 VDD1.n92 B 0.031756f
C112 VDD1.n93 B 0.031756f
C113 VDD1.n94 B 0.014226f
C114 VDD1.n95 B 0.013435f
C115 VDD1.n96 B 0.025003f
C116 VDD1.n97 B 0.025003f
C117 VDD1.n98 B 0.013435f
C118 VDD1.n99 B 0.014226f
C119 VDD1.n100 B 0.031756f
C120 VDD1.n101 B 0.031756f
C121 VDD1.n102 B 0.014226f
C122 VDD1.n103 B 0.013435f
C123 VDD1.n104 B 0.025003f
C124 VDD1.n105 B 0.025003f
C125 VDD1.n106 B 0.013435f
C126 VDD1.n107 B 0.013435f
C127 VDD1.n108 B 0.014226f
C128 VDD1.n109 B 0.031756f
C129 VDD1.n110 B 0.031756f
C130 VDD1.n111 B 0.031756f
C131 VDD1.n112 B 0.013831f
C132 VDD1.n113 B 0.013435f
C133 VDD1.n114 B 0.025003f
C134 VDD1.n115 B 0.025003f
C135 VDD1.n116 B 0.013435f
C136 VDD1.n117 B 0.014226f
C137 VDD1.n118 B 0.031756f
C138 VDD1.n119 B 0.031756f
C139 VDD1.n120 B 0.014226f
C140 VDD1.n121 B 0.013435f
C141 VDD1.n122 B 0.025003f
C142 VDD1.n123 B 0.025003f
C143 VDD1.n124 B 0.013435f
C144 VDD1.n125 B 0.014226f
C145 VDD1.n126 B 0.031756f
C146 VDD1.n127 B 0.065167f
C147 VDD1.n128 B 0.014226f
C148 VDD1.n129 B 0.013435f
C149 VDD1.n130 B 0.053694f
C150 VDD1.n131 B 0.072686f
C151 VDD1.t9 B 0.237095f
C152 VDD1.t2 B 0.237095f
C153 VDD1.n132 B 2.10978f
C154 VDD1.n133 B 0.810727f
C155 VDD1.t6 B 0.237095f
C156 VDD1.t1 B 0.237095f
C157 VDD1.n134 B 2.13491f
C158 VDD1.n135 B 3.45556f
C159 VDD1.t7 B 0.237095f
C160 VDD1.t8 B 0.237095f
C161 VDD1.n136 B 2.10978f
C162 VDD1.n137 B 3.49677f
C163 VP.t8 B 2.03318f
C164 VP.n0 B 0.779557f
C165 VP.n1 B 0.018453f
C166 VP.n2 B 0.024271f
C167 VP.n3 B 0.018453f
C168 VP.n4 B 0.019015f
C169 VP.n5 B 0.018453f
C170 VP.n6 B 0.017398f
C171 VP.n7 B 0.018453f
C172 VP.t7 B 2.03318f
C173 VP.n8 B 0.713982f
C174 VP.n9 B 0.018453f
C175 VP.n10 B 0.017398f
C176 VP.n11 B 0.018453f
C177 VP.t0 B 2.03318f
C178 VP.n12 B 0.713982f
C179 VP.n13 B 0.018453f
C180 VP.n14 B 0.029376f
C181 VP.n15 B 0.018453f
C182 VP.n16 B 0.022394f
C183 VP.t1 B 2.03318f
C184 VP.n17 B 0.779557f
C185 VP.n18 B 0.018453f
C186 VP.n19 B 0.024271f
C187 VP.n20 B 0.018453f
C188 VP.n21 B 0.019015f
C189 VP.n22 B 0.018453f
C190 VP.n23 B 0.017398f
C191 VP.n24 B 0.018453f
C192 VP.t4 B 2.03318f
C193 VP.n25 B 0.713982f
C194 VP.n26 B 0.018453f
C195 VP.n27 B 0.017398f
C196 VP.n28 B 0.018453f
C197 VP.t5 B 2.03318f
C198 VP.n29 B 0.783734f
C199 VP.t9 B 2.26858f
C200 VP.n30 B 0.741771f
C201 VP.n31 B 0.22569f
C202 VP.n32 B 0.032529f
C203 VP.n33 B 0.034219f
C204 VP.n34 B 0.033701f
C205 VP.n35 B 0.018453f
C206 VP.n36 B 0.018453f
C207 VP.n37 B 0.018453f
C208 VP.n38 B 0.036767f
C209 VP.n39 B 0.034219f
C210 VP.n40 B 0.025772f
C211 VP.n41 B 0.018453f
C212 VP.n42 B 0.018453f
C213 VP.n43 B 0.025772f
C214 VP.n44 B 0.034219f
C215 VP.n45 B 0.036767f
C216 VP.n46 B 0.018453f
C217 VP.n47 B 0.018453f
C218 VP.n48 B 0.018453f
C219 VP.n49 B 0.033701f
C220 VP.n50 B 0.034219f
C221 VP.t2 B 2.03318f
C222 VP.n51 B 0.713982f
C223 VP.n52 B 0.032529f
C224 VP.n53 B 0.018453f
C225 VP.n54 B 0.018453f
C226 VP.n55 B 0.018453f
C227 VP.n56 B 0.034219f
C228 VP.n57 B 0.034219f
C229 VP.n58 B 0.029376f
C230 VP.n59 B 0.018453f
C231 VP.n60 B 0.018453f
C232 VP.n61 B 0.018453f
C233 VP.n62 B 0.034219f
C234 VP.n63 B 0.034219f
C235 VP.n64 B 0.022394f
C236 VP.n65 B 0.029777f
C237 VP.n66 B 1.27422f
C238 VP.t6 B 2.03318f
C239 VP.n67 B 0.779557f
C240 VP.n68 B 1.28583f
C241 VP.n69 B 0.029777f
C242 VP.n70 B 0.018453f
C243 VP.n71 B 0.034219f
C244 VP.n72 B 0.034219f
C245 VP.n73 B 0.024271f
C246 VP.n74 B 0.018453f
C247 VP.n75 B 0.018453f
C248 VP.n76 B 0.018453f
C249 VP.n77 B 0.034219f
C250 VP.n78 B 0.034219f
C251 VP.n79 B 0.019015f
C252 VP.n80 B 0.018453f
C253 VP.n81 B 0.018453f
C254 VP.n82 B 0.032529f
C255 VP.n83 B 0.034219f
C256 VP.n84 B 0.033701f
C257 VP.n85 B 0.018453f
C258 VP.n86 B 0.018453f
C259 VP.n87 B 0.018453f
C260 VP.n88 B 0.036767f
C261 VP.n89 B 0.034219f
C262 VP.n90 B 0.025772f
C263 VP.n91 B 0.018453f
C264 VP.n92 B 0.018453f
C265 VP.n93 B 0.025772f
C266 VP.n94 B 0.034219f
C267 VP.n95 B 0.036767f
C268 VP.n96 B 0.018453f
C269 VP.n97 B 0.018453f
C270 VP.n98 B 0.018453f
C271 VP.n99 B 0.033701f
C272 VP.n100 B 0.034219f
C273 VP.t3 B 2.03318f
C274 VP.n101 B 0.713982f
C275 VP.n102 B 0.032529f
C276 VP.n103 B 0.018453f
C277 VP.n104 B 0.018453f
C278 VP.n105 B 0.018453f
C279 VP.n106 B 0.034219f
C280 VP.n107 B 0.034219f
C281 VP.n108 B 0.029376f
C282 VP.n109 B 0.018453f
C283 VP.n110 B 0.018453f
C284 VP.n111 B 0.018453f
C285 VP.n112 B 0.034219f
C286 VP.n113 B 0.034219f
C287 VP.n114 B 0.022394f
C288 VP.n115 B 0.029777f
C289 VP.n116 B 0.049939f
C290 VDD2.n0 B 0.032712f
C291 VDD2.n1 B 0.024695f
C292 VDD2.n2 B 0.01327f
C293 VDD2.n3 B 0.031366f
C294 VDD2.n4 B 0.014051f
C295 VDD2.n5 B 0.024695f
C296 VDD2.n6 B 0.01327f
C297 VDD2.n7 B 0.031366f
C298 VDD2.n8 B 0.014051f
C299 VDD2.n9 B 0.024695f
C300 VDD2.n10 B 0.01366f
C301 VDD2.n11 B 0.031366f
C302 VDD2.n12 B 0.014051f
C303 VDD2.n13 B 0.024695f
C304 VDD2.n14 B 0.01327f
C305 VDD2.n15 B 0.031366f
C306 VDD2.n16 B 0.014051f
C307 VDD2.n17 B 0.024695f
C308 VDD2.n18 B 0.01327f
C309 VDD2.n19 B 0.023524f
C310 VDD2.n20 B 0.022173f
C311 VDD2.t9 B 0.052975f
C312 VDD2.n21 B 0.178049f
C313 VDD2.n22 B 1.24583f
C314 VDD2.n23 B 0.01327f
C315 VDD2.n24 B 0.014051f
C316 VDD2.n25 B 0.031366f
C317 VDD2.n26 B 0.031366f
C318 VDD2.n27 B 0.014051f
C319 VDD2.n28 B 0.01327f
C320 VDD2.n29 B 0.024695f
C321 VDD2.n30 B 0.024695f
C322 VDD2.n31 B 0.01327f
C323 VDD2.n32 B 0.014051f
C324 VDD2.n33 B 0.031366f
C325 VDD2.n34 B 0.031366f
C326 VDD2.n35 B 0.014051f
C327 VDD2.n36 B 0.01327f
C328 VDD2.n37 B 0.024695f
C329 VDD2.n38 B 0.024695f
C330 VDD2.n39 B 0.01327f
C331 VDD2.n40 B 0.01327f
C332 VDD2.n41 B 0.014051f
C333 VDD2.n42 B 0.031366f
C334 VDD2.n43 B 0.031366f
C335 VDD2.n44 B 0.031366f
C336 VDD2.n45 B 0.01366f
C337 VDD2.n46 B 0.01327f
C338 VDD2.n47 B 0.024695f
C339 VDD2.n48 B 0.024695f
C340 VDD2.n49 B 0.01327f
C341 VDD2.n50 B 0.014051f
C342 VDD2.n51 B 0.031366f
C343 VDD2.n52 B 0.031366f
C344 VDD2.n53 B 0.014051f
C345 VDD2.n54 B 0.01327f
C346 VDD2.n55 B 0.024695f
C347 VDD2.n56 B 0.024695f
C348 VDD2.n57 B 0.01327f
C349 VDD2.n58 B 0.014051f
C350 VDD2.n59 B 0.031366f
C351 VDD2.n60 B 0.064366f
C352 VDD2.n61 B 0.014051f
C353 VDD2.n62 B 0.01327f
C354 VDD2.n63 B 0.053033f
C355 VDD2.n64 B 0.071792f
C356 VDD2.t5 B 0.234178f
C357 VDD2.t1 B 0.234178f
C358 VDD2.n65 B 2.08383f
C359 VDD2.n66 B 0.800753f
C360 VDD2.t7 B 0.234178f
C361 VDD2.t2 B 0.234178f
C362 VDD2.n67 B 2.10864f
C363 VDD2.n68 B 3.26869f
C364 VDD2.n69 B 0.032712f
C365 VDD2.n70 B 0.024695f
C366 VDD2.n71 B 0.01327f
C367 VDD2.n72 B 0.031366f
C368 VDD2.n73 B 0.014051f
C369 VDD2.n74 B 0.024695f
C370 VDD2.n75 B 0.01327f
C371 VDD2.n76 B 0.031366f
C372 VDD2.n77 B 0.014051f
C373 VDD2.n78 B 0.024695f
C374 VDD2.n79 B 0.01366f
C375 VDD2.n80 B 0.031366f
C376 VDD2.n81 B 0.01327f
C377 VDD2.n82 B 0.014051f
C378 VDD2.n83 B 0.024695f
C379 VDD2.n84 B 0.01327f
C380 VDD2.n85 B 0.031366f
C381 VDD2.n86 B 0.014051f
C382 VDD2.n87 B 0.024695f
C383 VDD2.n88 B 0.01327f
C384 VDD2.n89 B 0.023524f
C385 VDD2.n90 B 0.022173f
C386 VDD2.t8 B 0.052975f
C387 VDD2.n91 B 0.178049f
C388 VDD2.n92 B 1.24583f
C389 VDD2.n93 B 0.01327f
C390 VDD2.n94 B 0.014051f
C391 VDD2.n95 B 0.031366f
C392 VDD2.n96 B 0.031366f
C393 VDD2.n97 B 0.014051f
C394 VDD2.n98 B 0.01327f
C395 VDD2.n99 B 0.024695f
C396 VDD2.n100 B 0.024695f
C397 VDD2.n101 B 0.01327f
C398 VDD2.n102 B 0.014051f
C399 VDD2.n103 B 0.031366f
C400 VDD2.n104 B 0.031366f
C401 VDD2.n105 B 0.014051f
C402 VDD2.n106 B 0.01327f
C403 VDD2.n107 B 0.024695f
C404 VDD2.n108 B 0.024695f
C405 VDD2.n109 B 0.01327f
C406 VDD2.n110 B 0.014051f
C407 VDD2.n111 B 0.031366f
C408 VDD2.n112 B 0.031366f
C409 VDD2.n113 B 0.031366f
C410 VDD2.n114 B 0.01366f
C411 VDD2.n115 B 0.01327f
C412 VDD2.n116 B 0.024695f
C413 VDD2.n117 B 0.024695f
C414 VDD2.n118 B 0.01327f
C415 VDD2.n119 B 0.014051f
C416 VDD2.n120 B 0.031366f
C417 VDD2.n121 B 0.031366f
C418 VDD2.n122 B 0.014051f
C419 VDD2.n123 B 0.01327f
C420 VDD2.n124 B 0.024695f
C421 VDD2.n125 B 0.024695f
C422 VDD2.n126 B 0.01327f
C423 VDD2.n127 B 0.014051f
C424 VDD2.n128 B 0.031366f
C425 VDD2.n129 B 0.064366f
C426 VDD2.n130 B 0.014051f
C427 VDD2.n131 B 0.01327f
C428 VDD2.n132 B 0.053033f
C429 VDD2.n133 B 0.05261f
C430 VDD2.n134 B 3.14921f
C431 VDD2.t6 B 0.234178f
C432 VDD2.t0 B 0.234178f
C433 VDD2.n135 B 2.08383f
C434 VDD2.n136 B 0.529142f
C435 VDD2.t4 B 0.234178f
C436 VDD2.t3 B 0.234178f
C437 VDD2.n137 B 2.10859f
C438 VTAIL.t19 B 0.242287f
C439 VTAIL.t12 B 0.242287f
C440 VTAIL.n0 B 2.07445f
C441 VTAIL.n1 B 0.632952f
C442 VTAIL.n2 B 0.033845f
C443 VTAIL.n3 B 0.02555f
C444 VTAIL.n4 B 0.01373f
C445 VTAIL.n5 B 0.032452f
C446 VTAIL.n6 B 0.014537f
C447 VTAIL.n7 B 0.02555f
C448 VTAIL.n8 B 0.01373f
C449 VTAIL.n9 B 0.032452f
C450 VTAIL.n10 B 0.014537f
C451 VTAIL.n11 B 0.02555f
C452 VTAIL.n12 B 0.014133f
C453 VTAIL.n13 B 0.032452f
C454 VTAIL.n14 B 0.014537f
C455 VTAIL.n15 B 0.02555f
C456 VTAIL.n16 B 0.01373f
C457 VTAIL.n17 B 0.032452f
C458 VTAIL.n18 B 0.014537f
C459 VTAIL.n19 B 0.02555f
C460 VTAIL.n20 B 0.01373f
C461 VTAIL.n21 B 0.024339f
C462 VTAIL.n22 B 0.022941f
C463 VTAIL.t8 B 0.054809f
C464 VTAIL.n23 B 0.184214f
C465 VTAIL.n24 B 1.28897f
C466 VTAIL.n25 B 0.01373f
C467 VTAIL.n26 B 0.014537f
C468 VTAIL.n27 B 0.032452f
C469 VTAIL.n28 B 0.032452f
C470 VTAIL.n29 B 0.014537f
C471 VTAIL.n30 B 0.01373f
C472 VTAIL.n31 B 0.02555f
C473 VTAIL.n32 B 0.02555f
C474 VTAIL.n33 B 0.01373f
C475 VTAIL.n34 B 0.014537f
C476 VTAIL.n35 B 0.032452f
C477 VTAIL.n36 B 0.032452f
C478 VTAIL.n37 B 0.014537f
C479 VTAIL.n38 B 0.01373f
C480 VTAIL.n39 B 0.02555f
C481 VTAIL.n40 B 0.02555f
C482 VTAIL.n41 B 0.01373f
C483 VTAIL.n42 B 0.01373f
C484 VTAIL.n43 B 0.014537f
C485 VTAIL.n44 B 0.032452f
C486 VTAIL.n45 B 0.032452f
C487 VTAIL.n46 B 0.032452f
C488 VTAIL.n47 B 0.014133f
C489 VTAIL.n48 B 0.01373f
C490 VTAIL.n49 B 0.02555f
C491 VTAIL.n50 B 0.02555f
C492 VTAIL.n51 B 0.01373f
C493 VTAIL.n52 B 0.014537f
C494 VTAIL.n53 B 0.032452f
C495 VTAIL.n54 B 0.032452f
C496 VTAIL.n55 B 0.014537f
C497 VTAIL.n56 B 0.01373f
C498 VTAIL.n57 B 0.02555f
C499 VTAIL.n58 B 0.02555f
C500 VTAIL.n59 B 0.01373f
C501 VTAIL.n60 B 0.014537f
C502 VTAIL.n61 B 0.032452f
C503 VTAIL.n62 B 0.066594f
C504 VTAIL.n63 B 0.014537f
C505 VTAIL.n64 B 0.01373f
C506 VTAIL.n65 B 0.05487f
C507 VTAIL.n66 B 0.036753f
C508 VTAIL.n67 B 0.452042f
C509 VTAIL.t7 B 0.242287f
C510 VTAIL.t5 B 0.242287f
C511 VTAIL.n68 B 2.07445f
C512 VTAIL.n69 B 0.786431f
C513 VTAIL.t1 B 0.242287f
C514 VTAIL.t3 B 0.242287f
C515 VTAIL.n70 B 2.07445f
C516 VTAIL.n71 B 2.24778f
C517 VTAIL.t14 B 0.242287f
C518 VTAIL.t11 B 0.242287f
C519 VTAIL.n72 B 2.07446f
C520 VTAIL.n73 B 2.24776f
C521 VTAIL.t15 B 0.242287f
C522 VTAIL.t17 B 0.242287f
C523 VTAIL.n74 B 2.07446f
C524 VTAIL.n75 B 0.786418f
C525 VTAIL.n76 B 0.033845f
C526 VTAIL.n77 B 0.02555f
C527 VTAIL.n78 B 0.01373f
C528 VTAIL.n79 B 0.032452f
C529 VTAIL.n80 B 0.014537f
C530 VTAIL.n81 B 0.02555f
C531 VTAIL.n82 B 0.01373f
C532 VTAIL.n83 B 0.032452f
C533 VTAIL.n84 B 0.014537f
C534 VTAIL.n85 B 0.02555f
C535 VTAIL.n86 B 0.014133f
C536 VTAIL.n87 B 0.032452f
C537 VTAIL.n88 B 0.01373f
C538 VTAIL.n89 B 0.014537f
C539 VTAIL.n90 B 0.02555f
C540 VTAIL.n91 B 0.01373f
C541 VTAIL.n92 B 0.032452f
C542 VTAIL.n93 B 0.014537f
C543 VTAIL.n94 B 0.02555f
C544 VTAIL.n95 B 0.01373f
C545 VTAIL.n96 B 0.024339f
C546 VTAIL.n97 B 0.022941f
C547 VTAIL.t18 B 0.054809f
C548 VTAIL.n98 B 0.184214f
C549 VTAIL.n99 B 1.28897f
C550 VTAIL.n100 B 0.01373f
C551 VTAIL.n101 B 0.014537f
C552 VTAIL.n102 B 0.032452f
C553 VTAIL.n103 B 0.032452f
C554 VTAIL.n104 B 0.014537f
C555 VTAIL.n105 B 0.01373f
C556 VTAIL.n106 B 0.02555f
C557 VTAIL.n107 B 0.02555f
C558 VTAIL.n108 B 0.01373f
C559 VTAIL.n109 B 0.014537f
C560 VTAIL.n110 B 0.032452f
C561 VTAIL.n111 B 0.032452f
C562 VTAIL.n112 B 0.014537f
C563 VTAIL.n113 B 0.01373f
C564 VTAIL.n114 B 0.02555f
C565 VTAIL.n115 B 0.02555f
C566 VTAIL.n116 B 0.01373f
C567 VTAIL.n117 B 0.014537f
C568 VTAIL.n118 B 0.032452f
C569 VTAIL.n119 B 0.032452f
C570 VTAIL.n120 B 0.032452f
C571 VTAIL.n121 B 0.014133f
C572 VTAIL.n122 B 0.01373f
C573 VTAIL.n123 B 0.02555f
C574 VTAIL.n124 B 0.02555f
C575 VTAIL.n125 B 0.01373f
C576 VTAIL.n126 B 0.014537f
C577 VTAIL.n127 B 0.032452f
C578 VTAIL.n128 B 0.032452f
C579 VTAIL.n129 B 0.014537f
C580 VTAIL.n130 B 0.01373f
C581 VTAIL.n131 B 0.02555f
C582 VTAIL.n132 B 0.02555f
C583 VTAIL.n133 B 0.01373f
C584 VTAIL.n134 B 0.014537f
C585 VTAIL.n135 B 0.032452f
C586 VTAIL.n136 B 0.066594f
C587 VTAIL.n137 B 0.014537f
C588 VTAIL.n138 B 0.01373f
C589 VTAIL.n139 B 0.05487f
C590 VTAIL.n140 B 0.036753f
C591 VTAIL.n141 B 0.452042f
C592 VTAIL.t4 B 0.242287f
C593 VTAIL.t0 B 0.242287f
C594 VTAIL.n142 B 2.07446f
C595 VTAIL.n143 B 0.693798f
C596 VTAIL.t6 B 0.242287f
C597 VTAIL.t9 B 0.242287f
C598 VTAIL.n144 B 2.07446f
C599 VTAIL.n145 B 0.786418f
C600 VTAIL.n146 B 0.033845f
C601 VTAIL.n147 B 0.02555f
C602 VTAIL.n148 B 0.01373f
C603 VTAIL.n149 B 0.032452f
C604 VTAIL.n150 B 0.014537f
C605 VTAIL.n151 B 0.02555f
C606 VTAIL.n152 B 0.01373f
C607 VTAIL.n153 B 0.032452f
C608 VTAIL.n154 B 0.014537f
C609 VTAIL.n155 B 0.02555f
C610 VTAIL.n156 B 0.014133f
C611 VTAIL.n157 B 0.032452f
C612 VTAIL.n158 B 0.01373f
C613 VTAIL.n159 B 0.014537f
C614 VTAIL.n160 B 0.02555f
C615 VTAIL.n161 B 0.01373f
C616 VTAIL.n162 B 0.032452f
C617 VTAIL.n163 B 0.014537f
C618 VTAIL.n164 B 0.02555f
C619 VTAIL.n165 B 0.01373f
C620 VTAIL.n166 B 0.024339f
C621 VTAIL.n167 B 0.022941f
C622 VTAIL.t2 B 0.054809f
C623 VTAIL.n168 B 0.184214f
C624 VTAIL.n169 B 1.28897f
C625 VTAIL.n170 B 0.01373f
C626 VTAIL.n171 B 0.014537f
C627 VTAIL.n172 B 0.032452f
C628 VTAIL.n173 B 0.032452f
C629 VTAIL.n174 B 0.014537f
C630 VTAIL.n175 B 0.01373f
C631 VTAIL.n176 B 0.02555f
C632 VTAIL.n177 B 0.02555f
C633 VTAIL.n178 B 0.01373f
C634 VTAIL.n179 B 0.014537f
C635 VTAIL.n180 B 0.032452f
C636 VTAIL.n181 B 0.032452f
C637 VTAIL.n182 B 0.014537f
C638 VTAIL.n183 B 0.01373f
C639 VTAIL.n184 B 0.02555f
C640 VTAIL.n185 B 0.02555f
C641 VTAIL.n186 B 0.01373f
C642 VTAIL.n187 B 0.014537f
C643 VTAIL.n188 B 0.032452f
C644 VTAIL.n189 B 0.032452f
C645 VTAIL.n190 B 0.032452f
C646 VTAIL.n191 B 0.014133f
C647 VTAIL.n192 B 0.01373f
C648 VTAIL.n193 B 0.02555f
C649 VTAIL.n194 B 0.02555f
C650 VTAIL.n195 B 0.01373f
C651 VTAIL.n196 B 0.014537f
C652 VTAIL.n197 B 0.032452f
C653 VTAIL.n198 B 0.032452f
C654 VTAIL.n199 B 0.014537f
C655 VTAIL.n200 B 0.01373f
C656 VTAIL.n201 B 0.02555f
C657 VTAIL.n202 B 0.02555f
C658 VTAIL.n203 B 0.01373f
C659 VTAIL.n204 B 0.014537f
C660 VTAIL.n205 B 0.032452f
C661 VTAIL.n206 B 0.066594f
C662 VTAIL.n207 B 0.014537f
C663 VTAIL.n208 B 0.01373f
C664 VTAIL.n209 B 0.05487f
C665 VTAIL.n210 B 0.036753f
C666 VTAIL.n211 B 1.74341f
C667 VTAIL.n212 B 0.033845f
C668 VTAIL.n213 B 0.02555f
C669 VTAIL.n214 B 0.01373f
C670 VTAIL.n215 B 0.032452f
C671 VTAIL.n216 B 0.014537f
C672 VTAIL.n217 B 0.02555f
C673 VTAIL.n218 B 0.01373f
C674 VTAIL.n219 B 0.032452f
C675 VTAIL.n220 B 0.014537f
C676 VTAIL.n221 B 0.02555f
C677 VTAIL.n222 B 0.014133f
C678 VTAIL.n223 B 0.032452f
C679 VTAIL.n224 B 0.014537f
C680 VTAIL.n225 B 0.02555f
C681 VTAIL.n226 B 0.01373f
C682 VTAIL.n227 B 0.032452f
C683 VTAIL.n228 B 0.014537f
C684 VTAIL.n229 B 0.02555f
C685 VTAIL.n230 B 0.01373f
C686 VTAIL.n231 B 0.024339f
C687 VTAIL.n232 B 0.022941f
C688 VTAIL.t10 B 0.054809f
C689 VTAIL.n233 B 0.184214f
C690 VTAIL.n234 B 1.28897f
C691 VTAIL.n235 B 0.01373f
C692 VTAIL.n236 B 0.014537f
C693 VTAIL.n237 B 0.032452f
C694 VTAIL.n238 B 0.032452f
C695 VTAIL.n239 B 0.014537f
C696 VTAIL.n240 B 0.01373f
C697 VTAIL.n241 B 0.02555f
C698 VTAIL.n242 B 0.02555f
C699 VTAIL.n243 B 0.01373f
C700 VTAIL.n244 B 0.014537f
C701 VTAIL.n245 B 0.032452f
C702 VTAIL.n246 B 0.032452f
C703 VTAIL.n247 B 0.014537f
C704 VTAIL.n248 B 0.01373f
C705 VTAIL.n249 B 0.02555f
C706 VTAIL.n250 B 0.02555f
C707 VTAIL.n251 B 0.01373f
C708 VTAIL.n252 B 0.01373f
C709 VTAIL.n253 B 0.014537f
C710 VTAIL.n254 B 0.032452f
C711 VTAIL.n255 B 0.032452f
C712 VTAIL.n256 B 0.032452f
C713 VTAIL.n257 B 0.014133f
C714 VTAIL.n258 B 0.01373f
C715 VTAIL.n259 B 0.02555f
C716 VTAIL.n260 B 0.02555f
C717 VTAIL.n261 B 0.01373f
C718 VTAIL.n262 B 0.014537f
C719 VTAIL.n263 B 0.032452f
C720 VTAIL.n264 B 0.032452f
C721 VTAIL.n265 B 0.014537f
C722 VTAIL.n266 B 0.01373f
C723 VTAIL.n267 B 0.02555f
C724 VTAIL.n268 B 0.02555f
C725 VTAIL.n269 B 0.01373f
C726 VTAIL.n270 B 0.014537f
C727 VTAIL.n271 B 0.032452f
C728 VTAIL.n272 B 0.066594f
C729 VTAIL.n273 B 0.014537f
C730 VTAIL.n274 B 0.01373f
C731 VTAIL.n275 B 0.05487f
C732 VTAIL.n276 B 0.036753f
C733 VTAIL.n277 B 1.74341f
C734 VTAIL.t16 B 0.242287f
C735 VTAIL.t13 B 0.242287f
C736 VTAIL.n278 B 2.07445f
C737 VTAIL.n279 B 0.58469f
C738 VN.t7 B 1.9951f
C739 VN.n0 B 0.764959f
C740 VN.n1 B 0.018107f
C741 VN.n2 B 0.023817f
C742 VN.n3 B 0.018107f
C743 VN.n4 B 0.018659f
C744 VN.n5 B 0.018107f
C745 VN.n6 B 0.017072f
C746 VN.n7 B 0.018107f
C747 VN.t8 B 1.9951f
C748 VN.n8 B 0.700612f
C749 VN.n9 B 0.018107f
C750 VN.n10 B 0.017072f
C751 VN.n11 B 0.018107f
C752 VN.t4 B 1.9951f
C753 VN.n12 B 0.769057f
C754 VN.t0 B 2.2261f
C755 VN.n13 B 0.727879f
C756 VN.n14 B 0.221463f
C757 VN.n15 B 0.03192f
C758 VN.n16 B 0.033578f
C759 VN.n17 B 0.03307f
C760 VN.n18 B 0.018107f
C761 VN.n19 B 0.018107f
C762 VN.n20 B 0.018107f
C763 VN.n21 B 0.036079f
C764 VN.n22 B 0.033578f
C765 VN.n23 B 0.02529f
C766 VN.n24 B 0.018107f
C767 VN.n25 B 0.018107f
C768 VN.n26 B 0.02529f
C769 VN.n27 B 0.033578f
C770 VN.n28 B 0.036079f
C771 VN.n29 B 0.018107f
C772 VN.n30 B 0.018107f
C773 VN.n31 B 0.018107f
C774 VN.n32 B 0.03307f
C775 VN.n33 B 0.033578f
C776 VN.t2 B 1.9951f
C777 VN.n34 B 0.700612f
C778 VN.n35 B 0.03192f
C779 VN.n36 B 0.018107f
C780 VN.n37 B 0.018107f
C781 VN.n38 B 0.018107f
C782 VN.n39 B 0.033578f
C783 VN.n40 B 0.033578f
C784 VN.n41 B 0.028826f
C785 VN.n42 B 0.018107f
C786 VN.n43 B 0.018107f
C787 VN.n44 B 0.018107f
C788 VN.n45 B 0.033578f
C789 VN.n46 B 0.033578f
C790 VN.n47 B 0.021974f
C791 VN.n48 B 0.02922f
C792 VN.n49 B 0.049004f
C793 VN.t1 B 1.9951f
C794 VN.n50 B 0.764959f
C795 VN.n51 B 0.018107f
C796 VN.n52 B 0.023817f
C797 VN.n53 B 0.018107f
C798 VN.n54 B 0.018659f
C799 VN.n55 B 0.018107f
C800 VN.t3 B 1.9951f
C801 VN.n56 B 0.700612f
C802 VN.n57 B 0.017072f
C803 VN.n58 B 0.018107f
C804 VN.t9 B 1.9951f
C805 VN.n59 B 0.700612f
C806 VN.n60 B 0.018107f
C807 VN.n61 B 0.017072f
C808 VN.n62 B 0.018107f
C809 VN.t5 B 1.9951f
C810 VN.n63 B 0.769057f
C811 VN.t6 B 2.2261f
C812 VN.n64 B 0.727879f
C813 VN.n65 B 0.221463f
C814 VN.n66 B 0.03192f
C815 VN.n67 B 0.033578f
C816 VN.n68 B 0.03307f
C817 VN.n69 B 0.018107f
C818 VN.n70 B 0.018107f
C819 VN.n71 B 0.018107f
C820 VN.n72 B 0.036079f
C821 VN.n73 B 0.033578f
C822 VN.n74 B 0.02529f
C823 VN.n75 B 0.018107f
C824 VN.n76 B 0.018107f
C825 VN.n77 B 0.02529f
C826 VN.n78 B 0.033578f
C827 VN.n79 B 0.036079f
C828 VN.n80 B 0.018107f
C829 VN.n81 B 0.018107f
C830 VN.n82 B 0.018107f
C831 VN.n83 B 0.03307f
C832 VN.n84 B 0.033578f
C833 VN.n85 B 0.03192f
C834 VN.n86 B 0.018107f
C835 VN.n87 B 0.018107f
C836 VN.n88 B 0.018107f
C837 VN.n89 B 0.033578f
C838 VN.n90 B 0.033578f
C839 VN.n91 B 0.028826f
C840 VN.n92 B 0.018107f
C841 VN.n93 B 0.018107f
C842 VN.n94 B 0.018107f
C843 VN.n95 B 0.033578f
C844 VN.n96 B 0.033578f
C845 VN.n97 B 0.021974f
C846 VN.n98 B 0.02922f
C847 VN.n99 B 1.25745f
.ends

