* NGSPICE file created from diff_pair_sample_1188.ext - technology: sky130A

.subckt diff_pair_sample_1188 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t8 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X1 VDD2.t6 VN.t1 VTAIL.t9 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X2 VTAIL.t11 VN.t2 VDD2.t5 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X3 B.t11 B.t9 B.t10 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=6.8445 pd=35.88 as=0 ps=0 w=17.55 l=1.09
X4 VTAIL.t15 VN.t3 VDD2.t4 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=6.8445 pd=35.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X5 VDD1.t7 VP.t0 VTAIL.t5 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X6 VTAIL.t7 VP.t1 VDD1.t6 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=6.8445 pd=35.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X7 VTAIL.t14 VN.t4 VDD2.t3 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=6.8445 pd=35.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X8 VDD2.t2 VN.t5 VTAIL.t13 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=6.8445 ps=35.88 w=17.55 l=1.09
X9 VTAIL.t1 VP.t2 VDD1.t5 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X10 B.t8 B.t6 B.t7 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=6.8445 pd=35.88 as=0 ps=0 w=17.55 l=1.09
X11 VDD1.t4 VP.t3 VTAIL.t6 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X12 VDD1.t3 VP.t4 VTAIL.t0 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=6.8445 ps=35.88 w=17.55 l=1.09
X13 B.t5 B.t3 B.t4 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=6.8445 pd=35.88 as=0 ps=0 w=17.55 l=1.09
X14 VTAIL.t10 VN.t6 VDD2.t1 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X15 VDD2.t0 VN.t7 VTAIL.t12 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=6.8445 ps=35.88 w=17.55 l=1.09
X16 VDD1.t2 VP.t5 VTAIL.t4 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=6.8445 ps=35.88 w=17.55 l=1.09
X17 VTAIL.t3 VP.t6 VDD1.t1 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=2.89575 pd=17.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X18 VTAIL.t2 VP.t7 VDD1.t0 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=6.8445 pd=35.88 as=2.89575 ps=17.88 w=17.55 l=1.09
X19 B.t2 B.t0 B.t1 w_n2390_n4478# sky130_fd_pr__pfet_01v8 ad=6.8445 pd=35.88 as=0 ps=0 w=17.55 l=1.09
R0 VN.n3 VN.t4 446.76
R1 VN.n16 VN.t5 446.76
R2 VN.n11 VN.t7 424.293
R3 VN.n24 VN.t3 424.293
R4 VN.n4 VN.t0 388.033
R5 VN.n1 VN.t2 388.033
R6 VN.n17 VN.t6 388.033
R7 VN.n14 VN.t1 388.033
R8 VN.n23 VN.n13 161.3
R9 VN.n22 VN.n21 161.3
R10 VN.n20 VN.n19 161.3
R11 VN.n18 VN.n15 161.3
R12 VN.n10 VN.n0 161.3
R13 VN.n9 VN.n8 161.3
R14 VN.n7 VN.n6 161.3
R15 VN.n5 VN.n2 161.3
R16 VN.n25 VN.n24 80.6037
R17 VN.n12 VN.n11 80.6037
R18 VN.n6 VN.n5 56.5193
R19 VN.n19 VN.n18 56.5193
R20 VN VN.n25 48.4688
R21 VN.n11 VN.n10 48.4452
R22 VN.n24 VN.n23 48.4452
R23 VN.n4 VN.n3 34.0975
R24 VN.n17 VN.n16 34.0975
R25 VN.n16 VN.n15 28.4044
R26 VN.n3 VN.n2 28.4044
R27 VN.n10 VN.n9 24.4675
R28 VN.n23 VN.n22 24.4675
R29 VN.n5 VN.n4 22.5101
R30 VN.n6 VN.n1 22.5101
R31 VN.n18 VN.n17 22.5101
R32 VN.n19 VN.n14 22.5101
R33 VN.n9 VN.n1 1.95786
R34 VN.n22 VN.n14 1.95786
R35 VN.n25 VN.n13 0.285035
R36 VN.n12 VN.n0 0.285035
R37 VN.n21 VN.n13 0.189894
R38 VN.n21 VN.n20 0.189894
R39 VN.n20 VN.n15 0.189894
R40 VN.n7 VN.n2 0.189894
R41 VN.n8 VN.n7 0.189894
R42 VN.n8 VN.n0 0.189894
R43 VN VN.n12 0.146778
R44 VTAIL.n786 VTAIL.n694 756.745
R45 VTAIL.n94 VTAIL.n2 756.745
R46 VTAIL.n192 VTAIL.n100 756.745
R47 VTAIL.n292 VTAIL.n200 756.745
R48 VTAIL.n688 VTAIL.n596 756.745
R49 VTAIL.n588 VTAIL.n496 756.745
R50 VTAIL.n490 VTAIL.n398 756.745
R51 VTAIL.n390 VTAIL.n298 756.745
R52 VTAIL.n727 VTAIL.n726 585
R53 VTAIL.n729 VTAIL.n728 585
R54 VTAIL.n722 VTAIL.n721 585
R55 VTAIL.n735 VTAIL.n734 585
R56 VTAIL.n737 VTAIL.n736 585
R57 VTAIL.n718 VTAIL.n717 585
R58 VTAIL.n743 VTAIL.n742 585
R59 VTAIL.n745 VTAIL.n744 585
R60 VTAIL.n714 VTAIL.n713 585
R61 VTAIL.n751 VTAIL.n750 585
R62 VTAIL.n753 VTAIL.n752 585
R63 VTAIL.n710 VTAIL.n709 585
R64 VTAIL.n759 VTAIL.n758 585
R65 VTAIL.n761 VTAIL.n760 585
R66 VTAIL.n706 VTAIL.n705 585
R67 VTAIL.n768 VTAIL.n767 585
R68 VTAIL.n769 VTAIL.n704 585
R69 VTAIL.n771 VTAIL.n770 585
R70 VTAIL.n702 VTAIL.n701 585
R71 VTAIL.n777 VTAIL.n776 585
R72 VTAIL.n779 VTAIL.n778 585
R73 VTAIL.n698 VTAIL.n697 585
R74 VTAIL.n785 VTAIL.n784 585
R75 VTAIL.n787 VTAIL.n786 585
R76 VTAIL.n35 VTAIL.n34 585
R77 VTAIL.n37 VTAIL.n36 585
R78 VTAIL.n30 VTAIL.n29 585
R79 VTAIL.n43 VTAIL.n42 585
R80 VTAIL.n45 VTAIL.n44 585
R81 VTAIL.n26 VTAIL.n25 585
R82 VTAIL.n51 VTAIL.n50 585
R83 VTAIL.n53 VTAIL.n52 585
R84 VTAIL.n22 VTAIL.n21 585
R85 VTAIL.n59 VTAIL.n58 585
R86 VTAIL.n61 VTAIL.n60 585
R87 VTAIL.n18 VTAIL.n17 585
R88 VTAIL.n67 VTAIL.n66 585
R89 VTAIL.n69 VTAIL.n68 585
R90 VTAIL.n14 VTAIL.n13 585
R91 VTAIL.n76 VTAIL.n75 585
R92 VTAIL.n77 VTAIL.n12 585
R93 VTAIL.n79 VTAIL.n78 585
R94 VTAIL.n10 VTAIL.n9 585
R95 VTAIL.n85 VTAIL.n84 585
R96 VTAIL.n87 VTAIL.n86 585
R97 VTAIL.n6 VTAIL.n5 585
R98 VTAIL.n93 VTAIL.n92 585
R99 VTAIL.n95 VTAIL.n94 585
R100 VTAIL.n133 VTAIL.n132 585
R101 VTAIL.n135 VTAIL.n134 585
R102 VTAIL.n128 VTAIL.n127 585
R103 VTAIL.n141 VTAIL.n140 585
R104 VTAIL.n143 VTAIL.n142 585
R105 VTAIL.n124 VTAIL.n123 585
R106 VTAIL.n149 VTAIL.n148 585
R107 VTAIL.n151 VTAIL.n150 585
R108 VTAIL.n120 VTAIL.n119 585
R109 VTAIL.n157 VTAIL.n156 585
R110 VTAIL.n159 VTAIL.n158 585
R111 VTAIL.n116 VTAIL.n115 585
R112 VTAIL.n165 VTAIL.n164 585
R113 VTAIL.n167 VTAIL.n166 585
R114 VTAIL.n112 VTAIL.n111 585
R115 VTAIL.n174 VTAIL.n173 585
R116 VTAIL.n175 VTAIL.n110 585
R117 VTAIL.n177 VTAIL.n176 585
R118 VTAIL.n108 VTAIL.n107 585
R119 VTAIL.n183 VTAIL.n182 585
R120 VTAIL.n185 VTAIL.n184 585
R121 VTAIL.n104 VTAIL.n103 585
R122 VTAIL.n191 VTAIL.n190 585
R123 VTAIL.n193 VTAIL.n192 585
R124 VTAIL.n233 VTAIL.n232 585
R125 VTAIL.n235 VTAIL.n234 585
R126 VTAIL.n228 VTAIL.n227 585
R127 VTAIL.n241 VTAIL.n240 585
R128 VTAIL.n243 VTAIL.n242 585
R129 VTAIL.n224 VTAIL.n223 585
R130 VTAIL.n249 VTAIL.n248 585
R131 VTAIL.n251 VTAIL.n250 585
R132 VTAIL.n220 VTAIL.n219 585
R133 VTAIL.n257 VTAIL.n256 585
R134 VTAIL.n259 VTAIL.n258 585
R135 VTAIL.n216 VTAIL.n215 585
R136 VTAIL.n265 VTAIL.n264 585
R137 VTAIL.n267 VTAIL.n266 585
R138 VTAIL.n212 VTAIL.n211 585
R139 VTAIL.n274 VTAIL.n273 585
R140 VTAIL.n275 VTAIL.n210 585
R141 VTAIL.n277 VTAIL.n276 585
R142 VTAIL.n208 VTAIL.n207 585
R143 VTAIL.n283 VTAIL.n282 585
R144 VTAIL.n285 VTAIL.n284 585
R145 VTAIL.n204 VTAIL.n203 585
R146 VTAIL.n291 VTAIL.n290 585
R147 VTAIL.n293 VTAIL.n292 585
R148 VTAIL.n689 VTAIL.n688 585
R149 VTAIL.n687 VTAIL.n686 585
R150 VTAIL.n600 VTAIL.n599 585
R151 VTAIL.n681 VTAIL.n680 585
R152 VTAIL.n679 VTAIL.n678 585
R153 VTAIL.n604 VTAIL.n603 585
R154 VTAIL.n608 VTAIL.n606 585
R155 VTAIL.n673 VTAIL.n672 585
R156 VTAIL.n671 VTAIL.n670 585
R157 VTAIL.n610 VTAIL.n609 585
R158 VTAIL.n665 VTAIL.n664 585
R159 VTAIL.n663 VTAIL.n662 585
R160 VTAIL.n614 VTAIL.n613 585
R161 VTAIL.n657 VTAIL.n656 585
R162 VTAIL.n655 VTAIL.n654 585
R163 VTAIL.n618 VTAIL.n617 585
R164 VTAIL.n649 VTAIL.n648 585
R165 VTAIL.n647 VTAIL.n646 585
R166 VTAIL.n622 VTAIL.n621 585
R167 VTAIL.n641 VTAIL.n640 585
R168 VTAIL.n639 VTAIL.n638 585
R169 VTAIL.n626 VTAIL.n625 585
R170 VTAIL.n633 VTAIL.n632 585
R171 VTAIL.n631 VTAIL.n630 585
R172 VTAIL.n589 VTAIL.n588 585
R173 VTAIL.n587 VTAIL.n586 585
R174 VTAIL.n500 VTAIL.n499 585
R175 VTAIL.n581 VTAIL.n580 585
R176 VTAIL.n579 VTAIL.n578 585
R177 VTAIL.n504 VTAIL.n503 585
R178 VTAIL.n508 VTAIL.n506 585
R179 VTAIL.n573 VTAIL.n572 585
R180 VTAIL.n571 VTAIL.n570 585
R181 VTAIL.n510 VTAIL.n509 585
R182 VTAIL.n565 VTAIL.n564 585
R183 VTAIL.n563 VTAIL.n562 585
R184 VTAIL.n514 VTAIL.n513 585
R185 VTAIL.n557 VTAIL.n556 585
R186 VTAIL.n555 VTAIL.n554 585
R187 VTAIL.n518 VTAIL.n517 585
R188 VTAIL.n549 VTAIL.n548 585
R189 VTAIL.n547 VTAIL.n546 585
R190 VTAIL.n522 VTAIL.n521 585
R191 VTAIL.n541 VTAIL.n540 585
R192 VTAIL.n539 VTAIL.n538 585
R193 VTAIL.n526 VTAIL.n525 585
R194 VTAIL.n533 VTAIL.n532 585
R195 VTAIL.n531 VTAIL.n530 585
R196 VTAIL.n491 VTAIL.n490 585
R197 VTAIL.n489 VTAIL.n488 585
R198 VTAIL.n402 VTAIL.n401 585
R199 VTAIL.n483 VTAIL.n482 585
R200 VTAIL.n481 VTAIL.n480 585
R201 VTAIL.n406 VTAIL.n405 585
R202 VTAIL.n410 VTAIL.n408 585
R203 VTAIL.n475 VTAIL.n474 585
R204 VTAIL.n473 VTAIL.n472 585
R205 VTAIL.n412 VTAIL.n411 585
R206 VTAIL.n467 VTAIL.n466 585
R207 VTAIL.n465 VTAIL.n464 585
R208 VTAIL.n416 VTAIL.n415 585
R209 VTAIL.n459 VTAIL.n458 585
R210 VTAIL.n457 VTAIL.n456 585
R211 VTAIL.n420 VTAIL.n419 585
R212 VTAIL.n451 VTAIL.n450 585
R213 VTAIL.n449 VTAIL.n448 585
R214 VTAIL.n424 VTAIL.n423 585
R215 VTAIL.n443 VTAIL.n442 585
R216 VTAIL.n441 VTAIL.n440 585
R217 VTAIL.n428 VTAIL.n427 585
R218 VTAIL.n435 VTAIL.n434 585
R219 VTAIL.n433 VTAIL.n432 585
R220 VTAIL.n391 VTAIL.n390 585
R221 VTAIL.n389 VTAIL.n388 585
R222 VTAIL.n302 VTAIL.n301 585
R223 VTAIL.n383 VTAIL.n382 585
R224 VTAIL.n381 VTAIL.n380 585
R225 VTAIL.n306 VTAIL.n305 585
R226 VTAIL.n310 VTAIL.n308 585
R227 VTAIL.n375 VTAIL.n374 585
R228 VTAIL.n373 VTAIL.n372 585
R229 VTAIL.n312 VTAIL.n311 585
R230 VTAIL.n367 VTAIL.n366 585
R231 VTAIL.n365 VTAIL.n364 585
R232 VTAIL.n316 VTAIL.n315 585
R233 VTAIL.n359 VTAIL.n358 585
R234 VTAIL.n357 VTAIL.n356 585
R235 VTAIL.n320 VTAIL.n319 585
R236 VTAIL.n351 VTAIL.n350 585
R237 VTAIL.n349 VTAIL.n348 585
R238 VTAIL.n324 VTAIL.n323 585
R239 VTAIL.n343 VTAIL.n342 585
R240 VTAIL.n341 VTAIL.n340 585
R241 VTAIL.n328 VTAIL.n327 585
R242 VTAIL.n335 VTAIL.n334 585
R243 VTAIL.n333 VTAIL.n332 585
R244 VTAIL.n725 VTAIL.t12 327.466
R245 VTAIL.n33 VTAIL.t14 327.466
R246 VTAIL.n131 VTAIL.t4 327.466
R247 VTAIL.n231 VTAIL.t7 327.466
R248 VTAIL.n629 VTAIL.t0 327.466
R249 VTAIL.n529 VTAIL.t2 327.466
R250 VTAIL.n431 VTAIL.t13 327.466
R251 VTAIL.n331 VTAIL.t15 327.466
R252 VTAIL.n728 VTAIL.n727 171.744
R253 VTAIL.n728 VTAIL.n721 171.744
R254 VTAIL.n735 VTAIL.n721 171.744
R255 VTAIL.n736 VTAIL.n735 171.744
R256 VTAIL.n736 VTAIL.n717 171.744
R257 VTAIL.n743 VTAIL.n717 171.744
R258 VTAIL.n744 VTAIL.n743 171.744
R259 VTAIL.n744 VTAIL.n713 171.744
R260 VTAIL.n751 VTAIL.n713 171.744
R261 VTAIL.n752 VTAIL.n751 171.744
R262 VTAIL.n752 VTAIL.n709 171.744
R263 VTAIL.n759 VTAIL.n709 171.744
R264 VTAIL.n760 VTAIL.n759 171.744
R265 VTAIL.n760 VTAIL.n705 171.744
R266 VTAIL.n768 VTAIL.n705 171.744
R267 VTAIL.n769 VTAIL.n768 171.744
R268 VTAIL.n770 VTAIL.n769 171.744
R269 VTAIL.n770 VTAIL.n701 171.744
R270 VTAIL.n777 VTAIL.n701 171.744
R271 VTAIL.n778 VTAIL.n777 171.744
R272 VTAIL.n778 VTAIL.n697 171.744
R273 VTAIL.n785 VTAIL.n697 171.744
R274 VTAIL.n786 VTAIL.n785 171.744
R275 VTAIL.n36 VTAIL.n35 171.744
R276 VTAIL.n36 VTAIL.n29 171.744
R277 VTAIL.n43 VTAIL.n29 171.744
R278 VTAIL.n44 VTAIL.n43 171.744
R279 VTAIL.n44 VTAIL.n25 171.744
R280 VTAIL.n51 VTAIL.n25 171.744
R281 VTAIL.n52 VTAIL.n51 171.744
R282 VTAIL.n52 VTAIL.n21 171.744
R283 VTAIL.n59 VTAIL.n21 171.744
R284 VTAIL.n60 VTAIL.n59 171.744
R285 VTAIL.n60 VTAIL.n17 171.744
R286 VTAIL.n67 VTAIL.n17 171.744
R287 VTAIL.n68 VTAIL.n67 171.744
R288 VTAIL.n68 VTAIL.n13 171.744
R289 VTAIL.n76 VTAIL.n13 171.744
R290 VTAIL.n77 VTAIL.n76 171.744
R291 VTAIL.n78 VTAIL.n77 171.744
R292 VTAIL.n78 VTAIL.n9 171.744
R293 VTAIL.n85 VTAIL.n9 171.744
R294 VTAIL.n86 VTAIL.n85 171.744
R295 VTAIL.n86 VTAIL.n5 171.744
R296 VTAIL.n93 VTAIL.n5 171.744
R297 VTAIL.n94 VTAIL.n93 171.744
R298 VTAIL.n134 VTAIL.n133 171.744
R299 VTAIL.n134 VTAIL.n127 171.744
R300 VTAIL.n141 VTAIL.n127 171.744
R301 VTAIL.n142 VTAIL.n141 171.744
R302 VTAIL.n142 VTAIL.n123 171.744
R303 VTAIL.n149 VTAIL.n123 171.744
R304 VTAIL.n150 VTAIL.n149 171.744
R305 VTAIL.n150 VTAIL.n119 171.744
R306 VTAIL.n157 VTAIL.n119 171.744
R307 VTAIL.n158 VTAIL.n157 171.744
R308 VTAIL.n158 VTAIL.n115 171.744
R309 VTAIL.n165 VTAIL.n115 171.744
R310 VTAIL.n166 VTAIL.n165 171.744
R311 VTAIL.n166 VTAIL.n111 171.744
R312 VTAIL.n174 VTAIL.n111 171.744
R313 VTAIL.n175 VTAIL.n174 171.744
R314 VTAIL.n176 VTAIL.n175 171.744
R315 VTAIL.n176 VTAIL.n107 171.744
R316 VTAIL.n183 VTAIL.n107 171.744
R317 VTAIL.n184 VTAIL.n183 171.744
R318 VTAIL.n184 VTAIL.n103 171.744
R319 VTAIL.n191 VTAIL.n103 171.744
R320 VTAIL.n192 VTAIL.n191 171.744
R321 VTAIL.n234 VTAIL.n233 171.744
R322 VTAIL.n234 VTAIL.n227 171.744
R323 VTAIL.n241 VTAIL.n227 171.744
R324 VTAIL.n242 VTAIL.n241 171.744
R325 VTAIL.n242 VTAIL.n223 171.744
R326 VTAIL.n249 VTAIL.n223 171.744
R327 VTAIL.n250 VTAIL.n249 171.744
R328 VTAIL.n250 VTAIL.n219 171.744
R329 VTAIL.n257 VTAIL.n219 171.744
R330 VTAIL.n258 VTAIL.n257 171.744
R331 VTAIL.n258 VTAIL.n215 171.744
R332 VTAIL.n265 VTAIL.n215 171.744
R333 VTAIL.n266 VTAIL.n265 171.744
R334 VTAIL.n266 VTAIL.n211 171.744
R335 VTAIL.n274 VTAIL.n211 171.744
R336 VTAIL.n275 VTAIL.n274 171.744
R337 VTAIL.n276 VTAIL.n275 171.744
R338 VTAIL.n276 VTAIL.n207 171.744
R339 VTAIL.n283 VTAIL.n207 171.744
R340 VTAIL.n284 VTAIL.n283 171.744
R341 VTAIL.n284 VTAIL.n203 171.744
R342 VTAIL.n291 VTAIL.n203 171.744
R343 VTAIL.n292 VTAIL.n291 171.744
R344 VTAIL.n688 VTAIL.n687 171.744
R345 VTAIL.n687 VTAIL.n599 171.744
R346 VTAIL.n680 VTAIL.n599 171.744
R347 VTAIL.n680 VTAIL.n679 171.744
R348 VTAIL.n679 VTAIL.n603 171.744
R349 VTAIL.n608 VTAIL.n603 171.744
R350 VTAIL.n672 VTAIL.n608 171.744
R351 VTAIL.n672 VTAIL.n671 171.744
R352 VTAIL.n671 VTAIL.n609 171.744
R353 VTAIL.n664 VTAIL.n609 171.744
R354 VTAIL.n664 VTAIL.n663 171.744
R355 VTAIL.n663 VTAIL.n613 171.744
R356 VTAIL.n656 VTAIL.n613 171.744
R357 VTAIL.n656 VTAIL.n655 171.744
R358 VTAIL.n655 VTAIL.n617 171.744
R359 VTAIL.n648 VTAIL.n617 171.744
R360 VTAIL.n648 VTAIL.n647 171.744
R361 VTAIL.n647 VTAIL.n621 171.744
R362 VTAIL.n640 VTAIL.n621 171.744
R363 VTAIL.n640 VTAIL.n639 171.744
R364 VTAIL.n639 VTAIL.n625 171.744
R365 VTAIL.n632 VTAIL.n625 171.744
R366 VTAIL.n632 VTAIL.n631 171.744
R367 VTAIL.n588 VTAIL.n587 171.744
R368 VTAIL.n587 VTAIL.n499 171.744
R369 VTAIL.n580 VTAIL.n499 171.744
R370 VTAIL.n580 VTAIL.n579 171.744
R371 VTAIL.n579 VTAIL.n503 171.744
R372 VTAIL.n508 VTAIL.n503 171.744
R373 VTAIL.n572 VTAIL.n508 171.744
R374 VTAIL.n572 VTAIL.n571 171.744
R375 VTAIL.n571 VTAIL.n509 171.744
R376 VTAIL.n564 VTAIL.n509 171.744
R377 VTAIL.n564 VTAIL.n563 171.744
R378 VTAIL.n563 VTAIL.n513 171.744
R379 VTAIL.n556 VTAIL.n513 171.744
R380 VTAIL.n556 VTAIL.n555 171.744
R381 VTAIL.n555 VTAIL.n517 171.744
R382 VTAIL.n548 VTAIL.n517 171.744
R383 VTAIL.n548 VTAIL.n547 171.744
R384 VTAIL.n547 VTAIL.n521 171.744
R385 VTAIL.n540 VTAIL.n521 171.744
R386 VTAIL.n540 VTAIL.n539 171.744
R387 VTAIL.n539 VTAIL.n525 171.744
R388 VTAIL.n532 VTAIL.n525 171.744
R389 VTAIL.n532 VTAIL.n531 171.744
R390 VTAIL.n490 VTAIL.n489 171.744
R391 VTAIL.n489 VTAIL.n401 171.744
R392 VTAIL.n482 VTAIL.n401 171.744
R393 VTAIL.n482 VTAIL.n481 171.744
R394 VTAIL.n481 VTAIL.n405 171.744
R395 VTAIL.n410 VTAIL.n405 171.744
R396 VTAIL.n474 VTAIL.n410 171.744
R397 VTAIL.n474 VTAIL.n473 171.744
R398 VTAIL.n473 VTAIL.n411 171.744
R399 VTAIL.n466 VTAIL.n411 171.744
R400 VTAIL.n466 VTAIL.n465 171.744
R401 VTAIL.n465 VTAIL.n415 171.744
R402 VTAIL.n458 VTAIL.n415 171.744
R403 VTAIL.n458 VTAIL.n457 171.744
R404 VTAIL.n457 VTAIL.n419 171.744
R405 VTAIL.n450 VTAIL.n419 171.744
R406 VTAIL.n450 VTAIL.n449 171.744
R407 VTAIL.n449 VTAIL.n423 171.744
R408 VTAIL.n442 VTAIL.n423 171.744
R409 VTAIL.n442 VTAIL.n441 171.744
R410 VTAIL.n441 VTAIL.n427 171.744
R411 VTAIL.n434 VTAIL.n427 171.744
R412 VTAIL.n434 VTAIL.n433 171.744
R413 VTAIL.n390 VTAIL.n389 171.744
R414 VTAIL.n389 VTAIL.n301 171.744
R415 VTAIL.n382 VTAIL.n301 171.744
R416 VTAIL.n382 VTAIL.n381 171.744
R417 VTAIL.n381 VTAIL.n305 171.744
R418 VTAIL.n310 VTAIL.n305 171.744
R419 VTAIL.n374 VTAIL.n310 171.744
R420 VTAIL.n374 VTAIL.n373 171.744
R421 VTAIL.n373 VTAIL.n311 171.744
R422 VTAIL.n366 VTAIL.n311 171.744
R423 VTAIL.n366 VTAIL.n365 171.744
R424 VTAIL.n365 VTAIL.n315 171.744
R425 VTAIL.n358 VTAIL.n315 171.744
R426 VTAIL.n358 VTAIL.n357 171.744
R427 VTAIL.n357 VTAIL.n319 171.744
R428 VTAIL.n350 VTAIL.n319 171.744
R429 VTAIL.n350 VTAIL.n349 171.744
R430 VTAIL.n349 VTAIL.n323 171.744
R431 VTAIL.n342 VTAIL.n323 171.744
R432 VTAIL.n342 VTAIL.n341 171.744
R433 VTAIL.n341 VTAIL.n327 171.744
R434 VTAIL.n334 VTAIL.n327 171.744
R435 VTAIL.n334 VTAIL.n333 171.744
R436 VTAIL.n727 VTAIL.t12 85.8723
R437 VTAIL.n35 VTAIL.t14 85.8723
R438 VTAIL.n133 VTAIL.t4 85.8723
R439 VTAIL.n233 VTAIL.t7 85.8723
R440 VTAIL.n631 VTAIL.t0 85.8723
R441 VTAIL.n531 VTAIL.t2 85.8723
R442 VTAIL.n433 VTAIL.t13 85.8723
R443 VTAIL.n333 VTAIL.t15 85.8723
R444 VTAIL.n595 VTAIL.n594 52.9253
R445 VTAIL.n397 VTAIL.n396 52.9253
R446 VTAIL.n1 VTAIL.n0 52.9251
R447 VTAIL.n199 VTAIL.n198 52.9251
R448 VTAIL.n791 VTAIL.n790 32.7672
R449 VTAIL.n99 VTAIL.n98 32.7672
R450 VTAIL.n197 VTAIL.n196 32.7672
R451 VTAIL.n297 VTAIL.n296 32.7672
R452 VTAIL.n693 VTAIL.n692 32.7672
R453 VTAIL.n593 VTAIL.n592 32.7672
R454 VTAIL.n495 VTAIL.n494 32.7672
R455 VTAIL.n395 VTAIL.n394 32.7672
R456 VTAIL.n791 VTAIL.n693 28.7203
R457 VTAIL.n395 VTAIL.n297 28.7203
R458 VTAIL.n726 VTAIL.n725 16.3895
R459 VTAIL.n34 VTAIL.n33 16.3895
R460 VTAIL.n132 VTAIL.n131 16.3895
R461 VTAIL.n232 VTAIL.n231 16.3895
R462 VTAIL.n630 VTAIL.n629 16.3895
R463 VTAIL.n530 VTAIL.n529 16.3895
R464 VTAIL.n432 VTAIL.n431 16.3895
R465 VTAIL.n332 VTAIL.n331 16.3895
R466 VTAIL.n771 VTAIL.n702 13.1884
R467 VTAIL.n79 VTAIL.n10 13.1884
R468 VTAIL.n177 VTAIL.n108 13.1884
R469 VTAIL.n277 VTAIL.n208 13.1884
R470 VTAIL.n606 VTAIL.n604 13.1884
R471 VTAIL.n506 VTAIL.n504 13.1884
R472 VTAIL.n408 VTAIL.n406 13.1884
R473 VTAIL.n308 VTAIL.n306 13.1884
R474 VTAIL.n729 VTAIL.n724 12.8005
R475 VTAIL.n772 VTAIL.n704 12.8005
R476 VTAIL.n776 VTAIL.n775 12.8005
R477 VTAIL.n37 VTAIL.n32 12.8005
R478 VTAIL.n80 VTAIL.n12 12.8005
R479 VTAIL.n84 VTAIL.n83 12.8005
R480 VTAIL.n135 VTAIL.n130 12.8005
R481 VTAIL.n178 VTAIL.n110 12.8005
R482 VTAIL.n182 VTAIL.n181 12.8005
R483 VTAIL.n235 VTAIL.n230 12.8005
R484 VTAIL.n278 VTAIL.n210 12.8005
R485 VTAIL.n282 VTAIL.n281 12.8005
R486 VTAIL.n678 VTAIL.n677 12.8005
R487 VTAIL.n674 VTAIL.n673 12.8005
R488 VTAIL.n633 VTAIL.n628 12.8005
R489 VTAIL.n578 VTAIL.n577 12.8005
R490 VTAIL.n574 VTAIL.n573 12.8005
R491 VTAIL.n533 VTAIL.n528 12.8005
R492 VTAIL.n480 VTAIL.n479 12.8005
R493 VTAIL.n476 VTAIL.n475 12.8005
R494 VTAIL.n435 VTAIL.n430 12.8005
R495 VTAIL.n380 VTAIL.n379 12.8005
R496 VTAIL.n376 VTAIL.n375 12.8005
R497 VTAIL.n335 VTAIL.n330 12.8005
R498 VTAIL.n730 VTAIL.n722 12.0247
R499 VTAIL.n767 VTAIL.n766 12.0247
R500 VTAIL.n779 VTAIL.n700 12.0247
R501 VTAIL.n38 VTAIL.n30 12.0247
R502 VTAIL.n75 VTAIL.n74 12.0247
R503 VTAIL.n87 VTAIL.n8 12.0247
R504 VTAIL.n136 VTAIL.n128 12.0247
R505 VTAIL.n173 VTAIL.n172 12.0247
R506 VTAIL.n185 VTAIL.n106 12.0247
R507 VTAIL.n236 VTAIL.n228 12.0247
R508 VTAIL.n273 VTAIL.n272 12.0247
R509 VTAIL.n285 VTAIL.n206 12.0247
R510 VTAIL.n681 VTAIL.n602 12.0247
R511 VTAIL.n670 VTAIL.n607 12.0247
R512 VTAIL.n634 VTAIL.n626 12.0247
R513 VTAIL.n581 VTAIL.n502 12.0247
R514 VTAIL.n570 VTAIL.n507 12.0247
R515 VTAIL.n534 VTAIL.n526 12.0247
R516 VTAIL.n483 VTAIL.n404 12.0247
R517 VTAIL.n472 VTAIL.n409 12.0247
R518 VTAIL.n436 VTAIL.n428 12.0247
R519 VTAIL.n383 VTAIL.n304 12.0247
R520 VTAIL.n372 VTAIL.n309 12.0247
R521 VTAIL.n336 VTAIL.n328 12.0247
R522 VTAIL.n734 VTAIL.n733 11.249
R523 VTAIL.n765 VTAIL.n706 11.249
R524 VTAIL.n780 VTAIL.n698 11.249
R525 VTAIL.n42 VTAIL.n41 11.249
R526 VTAIL.n73 VTAIL.n14 11.249
R527 VTAIL.n88 VTAIL.n6 11.249
R528 VTAIL.n140 VTAIL.n139 11.249
R529 VTAIL.n171 VTAIL.n112 11.249
R530 VTAIL.n186 VTAIL.n104 11.249
R531 VTAIL.n240 VTAIL.n239 11.249
R532 VTAIL.n271 VTAIL.n212 11.249
R533 VTAIL.n286 VTAIL.n204 11.249
R534 VTAIL.n682 VTAIL.n600 11.249
R535 VTAIL.n669 VTAIL.n610 11.249
R536 VTAIL.n638 VTAIL.n637 11.249
R537 VTAIL.n582 VTAIL.n500 11.249
R538 VTAIL.n569 VTAIL.n510 11.249
R539 VTAIL.n538 VTAIL.n537 11.249
R540 VTAIL.n484 VTAIL.n402 11.249
R541 VTAIL.n471 VTAIL.n412 11.249
R542 VTAIL.n440 VTAIL.n439 11.249
R543 VTAIL.n384 VTAIL.n302 11.249
R544 VTAIL.n371 VTAIL.n312 11.249
R545 VTAIL.n340 VTAIL.n339 11.249
R546 VTAIL.n737 VTAIL.n720 10.4732
R547 VTAIL.n762 VTAIL.n761 10.4732
R548 VTAIL.n784 VTAIL.n783 10.4732
R549 VTAIL.n45 VTAIL.n28 10.4732
R550 VTAIL.n70 VTAIL.n69 10.4732
R551 VTAIL.n92 VTAIL.n91 10.4732
R552 VTAIL.n143 VTAIL.n126 10.4732
R553 VTAIL.n168 VTAIL.n167 10.4732
R554 VTAIL.n190 VTAIL.n189 10.4732
R555 VTAIL.n243 VTAIL.n226 10.4732
R556 VTAIL.n268 VTAIL.n267 10.4732
R557 VTAIL.n290 VTAIL.n289 10.4732
R558 VTAIL.n686 VTAIL.n685 10.4732
R559 VTAIL.n666 VTAIL.n665 10.4732
R560 VTAIL.n641 VTAIL.n624 10.4732
R561 VTAIL.n586 VTAIL.n585 10.4732
R562 VTAIL.n566 VTAIL.n565 10.4732
R563 VTAIL.n541 VTAIL.n524 10.4732
R564 VTAIL.n488 VTAIL.n487 10.4732
R565 VTAIL.n468 VTAIL.n467 10.4732
R566 VTAIL.n443 VTAIL.n426 10.4732
R567 VTAIL.n388 VTAIL.n387 10.4732
R568 VTAIL.n368 VTAIL.n367 10.4732
R569 VTAIL.n343 VTAIL.n326 10.4732
R570 VTAIL.n738 VTAIL.n718 9.69747
R571 VTAIL.n758 VTAIL.n708 9.69747
R572 VTAIL.n787 VTAIL.n696 9.69747
R573 VTAIL.n46 VTAIL.n26 9.69747
R574 VTAIL.n66 VTAIL.n16 9.69747
R575 VTAIL.n95 VTAIL.n4 9.69747
R576 VTAIL.n144 VTAIL.n124 9.69747
R577 VTAIL.n164 VTAIL.n114 9.69747
R578 VTAIL.n193 VTAIL.n102 9.69747
R579 VTAIL.n244 VTAIL.n224 9.69747
R580 VTAIL.n264 VTAIL.n214 9.69747
R581 VTAIL.n293 VTAIL.n202 9.69747
R582 VTAIL.n689 VTAIL.n598 9.69747
R583 VTAIL.n662 VTAIL.n612 9.69747
R584 VTAIL.n642 VTAIL.n622 9.69747
R585 VTAIL.n589 VTAIL.n498 9.69747
R586 VTAIL.n562 VTAIL.n512 9.69747
R587 VTAIL.n542 VTAIL.n522 9.69747
R588 VTAIL.n491 VTAIL.n400 9.69747
R589 VTAIL.n464 VTAIL.n414 9.69747
R590 VTAIL.n444 VTAIL.n424 9.69747
R591 VTAIL.n391 VTAIL.n300 9.69747
R592 VTAIL.n364 VTAIL.n314 9.69747
R593 VTAIL.n344 VTAIL.n324 9.69747
R594 VTAIL.n790 VTAIL.n789 9.45567
R595 VTAIL.n98 VTAIL.n97 9.45567
R596 VTAIL.n196 VTAIL.n195 9.45567
R597 VTAIL.n296 VTAIL.n295 9.45567
R598 VTAIL.n692 VTAIL.n691 9.45567
R599 VTAIL.n592 VTAIL.n591 9.45567
R600 VTAIL.n494 VTAIL.n493 9.45567
R601 VTAIL.n394 VTAIL.n393 9.45567
R602 VTAIL.n789 VTAIL.n788 9.3005
R603 VTAIL.n696 VTAIL.n695 9.3005
R604 VTAIL.n783 VTAIL.n782 9.3005
R605 VTAIL.n781 VTAIL.n780 9.3005
R606 VTAIL.n700 VTAIL.n699 9.3005
R607 VTAIL.n775 VTAIL.n774 9.3005
R608 VTAIL.n747 VTAIL.n746 9.3005
R609 VTAIL.n716 VTAIL.n715 9.3005
R610 VTAIL.n741 VTAIL.n740 9.3005
R611 VTAIL.n739 VTAIL.n738 9.3005
R612 VTAIL.n720 VTAIL.n719 9.3005
R613 VTAIL.n733 VTAIL.n732 9.3005
R614 VTAIL.n731 VTAIL.n730 9.3005
R615 VTAIL.n724 VTAIL.n723 9.3005
R616 VTAIL.n749 VTAIL.n748 9.3005
R617 VTAIL.n712 VTAIL.n711 9.3005
R618 VTAIL.n755 VTAIL.n754 9.3005
R619 VTAIL.n757 VTAIL.n756 9.3005
R620 VTAIL.n708 VTAIL.n707 9.3005
R621 VTAIL.n763 VTAIL.n762 9.3005
R622 VTAIL.n765 VTAIL.n764 9.3005
R623 VTAIL.n766 VTAIL.n703 9.3005
R624 VTAIL.n773 VTAIL.n772 9.3005
R625 VTAIL.n97 VTAIL.n96 9.3005
R626 VTAIL.n4 VTAIL.n3 9.3005
R627 VTAIL.n91 VTAIL.n90 9.3005
R628 VTAIL.n89 VTAIL.n88 9.3005
R629 VTAIL.n8 VTAIL.n7 9.3005
R630 VTAIL.n83 VTAIL.n82 9.3005
R631 VTAIL.n55 VTAIL.n54 9.3005
R632 VTAIL.n24 VTAIL.n23 9.3005
R633 VTAIL.n49 VTAIL.n48 9.3005
R634 VTAIL.n47 VTAIL.n46 9.3005
R635 VTAIL.n28 VTAIL.n27 9.3005
R636 VTAIL.n41 VTAIL.n40 9.3005
R637 VTAIL.n39 VTAIL.n38 9.3005
R638 VTAIL.n32 VTAIL.n31 9.3005
R639 VTAIL.n57 VTAIL.n56 9.3005
R640 VTAIL.n20 VTAIL.n19 9.3005
R641 VTAIL.n63 VTAIL.n62 9.3005
R642 VTAIL.n65 VTAIL.n64 9.3005
R643 VTAIL.n16 VTAIL.n15 9.3005
R644 VTAIL.n71 VTAIL.n70 9.3005
R645 VTAIL.n73 VTAIL.n72 9.3005
R646 VTAIL.n74 VTAIL.n11 9.3005
R647 VTAIL.n81 VTAIL.n80 9.3005
R648 VTAIL.n195 VTAIL.n194 9.3005
R649 VTAIL.n102 VTAIL.n101 9.3005
R650 VTAIL.n189 VTAIL.n188 9.3005
R651 VTAIL.n187 VTAIL.n186 9.3005
R652 VTAIL.n106 VTAIL.n105 9.3005
R653 VTAIL.n181 VTAIL.n180 9.3005
R654 VTAIL.n153 VTAIL.n152 9.3005
R655 VTAIL.n122 VTAIL.n121 9.3005
R656 VTAIL.n147 VTAIL.n146 9.3005
R657 VTAIL.n145 VTAIL.n144 9.3005
R658 VTAIL.n126 VTAIL.n125 9.3005
R659 VTAIL.n139 VTAIL.n138 9.3005
R660 VTAIL.n137 VTAIL.n136 9.3005
R661 VTAIL.n130 VTAIL.n129 9.3005
R662 VTAIL.n155 VTAIL.n154 9.3005
R663 VTAIL.n118 VTAIL.n117 9.3005
R664 VTAIL.n161 VTAIL.n160 9.3005
R665 VTAIL.n163 VTAIL.n162 9.3005
R666 VTAIL.n114 VTAIL.n113 9.3005
R667 VTAIL.n169 VTAIL.n168 9.3005
R668 VTAIL.n171 VTAIL.n170 9.3005
R669 VTAIL.n172 VTAIL.n109 9.3005
R670 VTAIL.n179 VTAIL.n178 9.3005
R671 VTAIL.n295 VTAIL.n294 9.3005
R672 VTAIL.n202 VTAIL.n201 9.3005
R673 VTAIL.n289 VTAIL.n288 9.3005
R674 VTAIL.n287 VTAIL.n286 9.3005
R675 VTAIL.n206 VTAIL.n205 9.3005
R676 VTAIL.n281 VTAIL.n280 9.3005
R677 VTAIL.n253 VTAIL.n252 9.3005
R678 VTAIL.n222 VTAIL.n221 9.3005
R679 VTAIL.n247 VTAIL.n246 9.3005
R680 VTAIL.n245 VTAIL.n244 9.3005
R681 VTAIL.n226 VTAIL.n225 9.3005
R682 VTAIL.n239 VTAIL.n238 9.3005
R683 VTAIL.n237 VTAIL.n236 9.3005
R684 VTAIL.n230 VTAIL.n229 9.3005
R685 VTAIL.n255 VTAIL.n254 9.3005
R686 VTAIL.n218 VTAIL.n217 9.3005
R687 VTAIL.n261 VTAIL.n260 9.3005
R688 VTAIL.n263 VTAIL.n262 9.3005
R689 VTAIL.n214 VTAIL.n213 9.3005
R690 VTAIL.n269 VTAIL.n268 9.3005
R691 VTAIL.n271 VTAIL.n270 9.3005
R692 VTAIL.n272 VTAIL.n209 9.3005
R693 VTAIL.n279 VTAIL.n278 9.3005
R694 VTAIL.n616 VTAIL.n615 9.3005
R695 VTAIL.n659 VTAIL.n658 9.3005
R696 VTAIL.n661 VTAIL.n660 9.3005
R697 VTAIL.n612 VTAIL.n611 9.3005
R698 VTAIL.n667 VTAIL.n666 9.3005
R699 VTAIL.n669 VTAIL.n668 9.3005
R700 VTAIL.n607 VTAIL.n605 9.3005
R701 VTAIL.n675 VTAIL.n674 9.3005
R702 VTAIL.n691 VTAIL.n690 9.3005
R703 VTAIL.n598 VTAIL.n597 9.3005
R704 VTAIL.n685 VTAIL.n684 9.3005
R705 VTAIL.n683 VTAIL.n682 9.3005
R706 VTAIL.n602 VTAIL.n601 9.3005
R707 VTAIL.n677 VTAIL.n676 9.3005
R708 VTAIL.n653 VTAIL.n652 9.3005
R709 VTAIL.n651 VTAIL.n650 9.3005
R710 VTAIL.n620 VTAIL.n619 9.3005
R711 VTAIL.n645 VTAIL.n644 9.3005
R712 VTAIL.n643 VTAIL.n642 9.3005
R713 VTAIL.n624 VTAIL.n623 9.3005
R714 VTAIL.n637 VTAIL.n636 9.3005
R715 VTAIL.n635 VTAIL.n634 9.3005
R716 VTAIL.n628 VTAIL.n627 9.3005
R717 VTAIL.n516 VTAIL.n515 9.3005
R718 VTAIL.n559 VTAIL.n558 9.3005
R719 VTAIL.n561 VTAIL.n560 9.3005
R720 VTAIL.n512 VTAIL.n511 9.3005
R721 VTAIL.n567 VTAIL.n566 9.3005
R722 VTAIL.n569 VTAIL.n568 9.3005
R723 VTAIL.n507 VTAIL.n505 9.3005
R724 VTAIL.n575 VTAIL.n574 9.3005
R725 VTAIL.n591 VTAIL.n590 9.3005
R726 VTAIL.n498 VTAIL.n497 9.3005
R727 VTAIL.n585 VTAIL.n584 9.3005
R728 VTAIL.n583 VTAIL.n582 9.3005
R729 VTAIL.n502 VTAIL.n501 9.3005
R730 VTAIL.n577 VTAIL.n576 9.3005
R731 VTAIL.n553 VTAIL.n552 9.3005
R732 VTAIL.n551 VTAIL.n550 9.3005
R733 VTAIL.n520 VTAIL.n519 9.3005
R734 VTAIL.n545 VTAIL.n544 9.3005
R735 VTAIL.n543 VTAIL.n542 9.3005
R736 VTAIL.n524 VTAIL.n523 9.3005
R737 VTAIL.n537 VTAIL.n536 9.3005
R738 VTAIL.n535 VTAIL.n534 9.3005
R739 VTAIL.n528 VTAIL.n527 9.3005
R740 VTAIL.n418 VTAIL.n417 9.3005
R741 VTAIL.n461 VTAIL.n460 9.3005
R742 VTAIL.n463 VTAIL.n462 9.3005
R743 VTAIL.n414 VTAIL.n413 9.3005
R744 VTAIL.n469 VTAIL.n468 9.3005
R745 VTAIL.n471 VTAIL.n470 9.3005
R746 VTAIL.n409 VTAIL.n407 9.3005
R747 VTAIL.n477 VTAIL.n476 9.3005
R748 VTAIL.n493 VTAIL.n492 9.3005
R749 VTAIL.n400 VTAIL.n399 9.3005
R750 VTAIL.n487 VTAIL.n486 9.3005
R751 VTAIL.n485 VTAIL.n484 9.3005
R752 VTAIL.n404 VTAIL.n403 9.3005
R753 VTAIL.n479 VTAIL.n478 9.3005
R754 VTAIL.n455 VTAIL.n454 9.3005
R755 VTAIL.n453 VTAIL.n452 9.3005
R756 VTAIL.n422 VTAIL.n421 9.3005
R757 VTAIL.n447 VTAIL.n446 9.3005
R758 VTAIL.n445 VTAIL.n444 9.3005
R759 VTAIL.n426 VTAIL.n425 9.3005
R760 VTAIL.n439 VTAIL.n438 9.3005
R761 VTAIL.n437 VTAIL.n436 9.3005
R762 VTAIL.n430 VTAIL.n429 9.3005
R763 VTAIL.n318 VTAIL.n317 9.3005
R764 VTAIL.n361 VTAIL.n360 9.3005
R765 VTAIL.n363 VTAIL.n362 9.3005
R766 VTAIL.n314 VTAIL.n313 9.3005
R767 VTAIL.n369 VTAIL.n368 9.3005
R768 VTAIL.n371 VTAIL.n370 9.3005
R769 VTAIL.n309 VTAIL.n307 9.3005
R770 VTAIL.n377 VTAIL.n376 9.3005
R771 VTAIL.n393 VTAIL.n392 9.3005
R772 VTAIL.n300 VTAIL.n299 9.3005
R773 VTAIL.n387 VTAIL.n386 9.3005
R774 VTAIL.n385 VTAIL.n384 9.3005
R775 VTAIL.n304 VTAIL.n303 9.3005
R776 VTAIL.n379 VTAIL.n378 9.3005
R777 VTAIL.n355 VTAIL.n354 9.3005
R778 VTAIL.n353 VTAIL.n352 9.3005
R779 VTAIL.n322 VTAIL.n321 9.3005
R780 VTAIL.n347 VTAIL.n346 9.3005
R781 VTAIL.n345 VTAIL.n344 9.3005
R782 VTAIL.n326 VTAIL.n325 9.3005
R783 VTAIL.n339 VTAIL.n338 9.3005
R784 VTAIL.n337 VTAIL.n336 9.3005
R785 VTAIL.n330 VTAIL.n329 9.3005
R786 VTAIL.n742 VTAIL.n741 8.92171
R787 VTAIL.n757 VTAIL.n710 8.92171
R788 VTAIL.n788 VTAIL.n694 8.92171
R789 VTAIL.n50 VTAIL.n49 8.92171
R790 VTAIL.n65 VTAIL.n18 8.92171
R791 VTAIL.n96 VTAIL.n2 8.92171
R792 VTAIL.n148 VTAIL.n147 8.92171
R793 VTAIL.n163 VTAIL.n116 8.92171
R794 VTAIL.n194 VTAIL.n100 8.92171
R795 VTAIL.n248 VTAIL.n247 8.92171
R796 VTAIL.n263 VTAIL.n216 8.92171
R797 VTAIL.n294 VTAIL.n200 8.92171
R798 VTAIL.n690 VTAIL.n596 8.92171
R799 VTAIL.n661 VTAIL.n614 8.92171
R800 VTAIL.n646 VTAIL.n645 8.92171
R801 VTAIL.n590 VTAIL.n496 8.92171
R802 VTAIL.n561 VTAIL.n514 8.92171
R803 VTAIL.n546 VTAIL.n545 8.92171
R804 VTAIL.n492 VTAIL.n398 8.92171
R805 VTAIL.n463 VTAIL.n416 8.92171
R806 VTAIL.n448 VTAIL.n447 8.92171
R807 VTAIL.n392 VTAIL.n298 8.92171
R808 VTAIL.n363 VTAIL.n316 8.92171
R809 VTAIL.n348 VTAIL.n347 8.92171
R810 VTAIL.n745 VTAIL.n716 8.14595
R811 VTAIL.n754 VTAIL.n753 8.14595
R812 VTAIL.n53 VTAIL.n24 8.14595
R813 VTAIL.n62 VTAIL.n61 8.14595
R814 VTAIL.n151 VTAIL.n122 8.14595
R815 VTAIL.n160 VTAIL.n159 8.14595
R816 VTAIL.n251 VTAIL.n222 8.14595
R817 VTAIL.n260 VTAIL.n259 8.14595
R818 VTAIL.n658 VTAIL.n657 8.14595
R819 VTAIL.n649 VTAIL.n620 8.14595
R820 VTAIL.n558 VTAIL.n557 8.14595
R821 VTAIL.n549 VTAIL.n520 8.14595
R822 VTAIL.n460 VTAIL.n459 8.14595
R823 VTAIL.n451 VTAIL.n422 8.14595
R824 VTAIL.n360 VTAIL.n359 8.14595
R825 VTAIL.n351 VTAIL.n322 8.14595
R826 VTAIL.n746 VTAIL.n714 7.3702
R827 VTAIL.n750 VTAIL.n712 7.3702
R828 VTAIL.n54 VTAIL.n22 7.3702
R829 VTAIL.n58 VTAIL.n20 7.3702
R830 VTAIL.n152 VTAIL.n120 7.3702
R831 VTAIL.n156 VTAIL.n118 7.3702
R832 VTAIL.n252 VTAIL.n220 7.3702
R833 VTAIL.n256 VTAIL.n218 7.3702
R834 VTAIL.n654 VTAIL.n616 7.3702
R835 VTAIL.n650 VTAIL.n618 7.3702
R836 VTAIL.n554 VTAIL.n516 7.3702
R837 VTAIL.n550 VTAIL.n518 7.3702
R838 VTAIL.n456 VTAIL.n418 7.3702
R839 VTAIL.n452 VTAIL.n420 7.3702
R840 VTAIL.n356 VTAIL.n318 7.3702
R841 VTAIL.n352 VTAIL.n320 7.3702
R842 VTAIL.n749 VTAIL.n714 6.59444
R843 VTAIL.n750 VTAIL.n749 6.59444
R844 VTAIL.n57 VTAIL.n22 6.59444
R845 VTAIL.n58 VTAIL.n57 6.59444
R846 VTAIL.n155 VTAIL.n120 6.59444
R847 VTAIL.n156 VTAIL.n155 6.59444
R848 VTAIL.n255 VTAIL.n220 6.59444
R849 VTAIL.n256 VTAIL.n255 6.59444
R850 VTAIL.n654 VTAIL.n653 6.59444
R851 VTAIL.n653 VTAIL.n618 6.59444
R852 VTAIL.n554 VTAIL.n553 6.59444
R853 VTAIL.n553 VTAIL.n518 6.59444
R854 VTAIL.n456 VTAIL.n455 6.59444
R855 VTAIL.n455 VTAIL.n420 6.59444
R856 VTAIL.n356 VTAIL.n355 6.59444
R857 VTAIL.n355 VTAIL.n320 6.59444
R858 VTAIL.n746 VTAIL.n745 5.81868
R859 VTAIL.n753 VTAIL.n712 5.81868
R860 VTAIL.n54 VTAIL.n53 5.81868
R861 VTAIL.n61 VTAIL.n20 5.81868
R862 VTAIL.n152 VTAIL.n151 5.81868
R863 VTAIL.n159 VTAIL.n118 5.81868
R864 VTAIL.n252 VTAIL.n251 5.81868
R865 VTAIL.n259 VTAIL.n218 5.81868
R866 VTAIL.n657 VTAIL.n616 5.81868
R867 VTAIL.n650 VTAIL.n649 5.81868
R868 VTAIL.n557 VTAIL.n516 5.81868
R869 VTAIL.n550 VTAIL.n549 5.81868
R870 VTAIL.n459 VTAIL.n418 5.81868
R871 VTAIL.n452 VTAIL.n451 5.81868
R872 VTAIL.n359 VTAIL.n318 5.81868
R873 VTAIL.n352 VTAIL.n351 5.81868
R874 VTAIL.n742 VTAIL.n716 5.04292
R875 VTAIL.n754 VTAIL.n710 5.04292
R876 VTAIL.n790 VTAIL.n694 5.04292
R877 VTAIL.n50 VTAIL.n24 5.04292
R878 VTAIL.n62 VTAIL.n18 5.04292
R879 VTAIL.n98 VTAIL.n2 5.04292
R880 VTAIL.n148 VTAIL.n122 5.04292
R881 VTAIL.n160 VTAIL.n116 5.04292
R882 VTAIL.n196 VTAIL.n100 5.04292
R883 VTAIL.n248 VTAIL.n222 5.04292
R884 VTAIL.n260 VTAIL.n216 5.04292
R885 VTAIL.n296 VTAIL.n200 5.04292
R886 VTAIL.n692 VTAIL.n596 5.04292
R887 VTAIL.n658 VTAIL.n614 5.04292
R888 VTAIL.n646 VTAIL.n620 5.04292
R889 VTAIL.n592 VTAIL.n496 5.04292
R890 VTAIL.n558 VTAIL.n514 5.04292
R891 VTAIL.n546 VTAIL.n520 5.04292
R892 VTAIL.n494 VTAIL.n398 5.04292
R893 VTAIL.n460 VTAIL.n416 5.04292
R894 VTAIL.n448 VTAIL.n422 5.04292
R895 VTAIL.n394 VTAIL.n298 5.04292
R896 VTAIL.n360 VTAIL.n316 5.04292
R897 VTAIL.n348 VTAIL.n322 5.04292
R898 VTAIL.n741 VTAIL.n718 4.26717
R899 VTAIL.n758 VTAIL.n757 4.26717
R900 VTAIL.n788 VTAIL.n787 4.26717
R901 VTAIL.n49 VTAIL.n26 4.26717
R902 VTAIL.n66 VTAIL.n65 4.26717
R903 VTAIL.n96 VTAIL.n95 4.26717
R904 VTAIL.n147 VTAIL.n124 4.26717
R905 VTAIL.n164 VTAIL.n163 4.26717
R906 VTAIL.n194 VTAIL.n193 4.26717
R907 VTAIL.n247 VTAIL.n224 4.26717
R908 VTAIL.n264 VTAIL.n263 4.26717
R909 VTAIL.n294 VTAIL.n293 4.26717
R910 VTAIL.n690 VTAIL.n689 4.26717
R911 VTAIL.n662 VTAIL.n661 4.26717
R912 VTAIL.n645 VTAIL.n622 4.26717
R913 VTAIL.n590 VTAIL.n589 4.26717
R914 VTAIL.n562 VTAIL.n561 4.26717
R915 VTAIL.n545 VTAIL.n522 4.26717
R916 VTAIL.n492 VTAIL.n491 4.26717
R917 VTAIL.n464 VTAIL.n463 4.26717
R918 VTAIL.n447 VTAIL.n424 4.26717
R919 VTAIL.n392 VTAIL.n391 4.26717
R920 VTAIL.n364 VTAIL.n363 4.26717
R921 VTAIL.n347 VTAIL.n324 4.26717
R922 VTAIL.n725 VTAIL.n723 3.70982
R923 VTAIL.n33 VTAIL.n31 3.70982
R924 VTAIL.n131 VTAIL.n129 3.70982
R925 VTAIL.n231 VTAIL.n229 3.70982
R926 VTAIL.n629 VTAIL.n627 3.70982
R927 VTAIL.n529 VTAIL.n527 3.70982
R928 VTAIL.n431 VTAIL.n429 3.70982
R929 VTAIL.n331 VTAIL.n329 3.70982
R930 VTAIL.n738 VTAIL.n737 3.49141
R931 VTAIL.n761 VTAIL.n708 3.49141
R932 VTAIL.n784 VTAIL.n696 3.49141
R933 VTAIL.n46 VTAIL.n45 3.49141
R934 VTAIL.n69 VTAIL.n16 3.49141
R935 VTAIL.n92 VTAIL.n4 3.49141
R936 VTAIL.n144 VTAIL.n143 3.49141
R937 VTAIL.n167 VTAIL.n114 3.49141
R938 VTAIL.n190 VTAIL.n102 3.49141
R939 VTAIL.n244 VTAIL.n243 3.49141
R940 VTAIL.n267 VTAIL.n214 3.49141
R941 VTAIL.n290 VTAIL.n202 3.49141
R942 VTAIL.n686 VTAIL.n598 3.49141
R943 VTAIL.n665 VTAIL.n612 3.49141
R944 VTAIL.n642 VTAIL.n641 3.49141
R945 VTAIL.n586 VTAIL.n498 3.49141
R946 VTAIL.n565 VTAIL.n512 3.49141
R947 VTAIL.n542 VTAIL.n541 3.49141
R948 VTAIL.n488 VTAIL.n400 3.49141
R949 VTAIL.n467 VTAIL.n414 3.49141
R950 VTAIL.n444 VTAIL.n443 3.49141
R951 VTAIL.n388 VTAIL.n300 3.49141
R952 VTAIL.n367 VTAIL.n314 3.49141
R953 VTAIL.n344 VTAIL.n343 3.49141
R954 VTAIL.n734 VTAIL.n720 2.71565
R955 VTAIL.n762 VTAIL.n706 2.71565
R956 VTAIL.n783 VTAIL.n698 2.71565
R957 VTAIL.n42 VTAIL.n28 2.71565
R958 VTAIL.n70 VTAIL.n14 2.71565
R959 VTAIL.n91 VTAIL.n6 2.71565
R960 VTAIL.n140 VTAIL.n126 2.71565
R961 VTAIL.n168 VTAIL.n112 2.71565
R962 VTAIL.n189 VTAIL.n104 2.71565
R963 VTAIL.n240 VTAIL.n226 2.71565
R964 VTAIL.n268 VTAIL.n212 2.71565
R965 VTAIL.n289 VTAIL.n204 2.71565
R966 VTAIL.n685 VTAIL.n600 2.71565
R967 VTAIL.n666 VTAIL.n610 2.71565
R968 VTAIL.n638 VTAIL.n624 2.71565
R969 VTAIL.n585 VTAIL.n500 2.71565
R970 VTAIL.n566 VTAIL.n510 2.71565
R971 VTAIL.n538 VTAIL.n524 2.71565
R972 VTAIL.n487 VTAIL.n402 2.71565
R973 VTAIL.n468 VTAIL.n412 2.71565
R974 VTAIL.n440 VTAIL.n426 2.71565
R975 VTAIL.n387 VTAIL.n302 2.71565
R976 VTAIL.n368 VTAIL.n312 2.71565
R977 VTAIL.n340 VTAIL.n326 2.71565
R978 VTAIL.n733 VTAIL.n722 1.93989
R979 VTAIL.n767 VTAIL.n765 1.93989
R980 VTAIL.n780 VTAIL.n779 1.93989
R981 VTAIL.n41 VTAIL.n30 1.93989
R982 VTAIL.n75 VTAIL.n73 1.93989
R983 VTAIL.n88 VTAIL.n87 1.93989
R984 VTAIL.n139 VTAIL.n128 1.93989
R985 VTAIL.n173 VTAIL.n171 1.93989
R986 VTAIL.n186 VTAIL.n185 1.93989
R987 VTAIL.n239 VTAIL.n228 1.93989
R988 VTAIL.n273 VTAIL.n271 1.93989
R989 VTAIL.n286 VTAIL.n285 1.93989
R990 VTAIL.n682 VTAIL.n681 1.93989
R991 VTAIL.n670 VTAIL.n669 1.93989
R992 VTAIL.n637 VTAIL.n626 1.93989
R993 VTAIL.n582 VTAIL.n581 1.93989
R994 VTAIL.n570 VTAIL.n569 1.93989
R995 VTAIL.n537 VTAIL.n526 1.93989
R996 VTAIL.n484 VTAIL.n483 1.93989
R997 VTAIL.n472 VTAIL.n471 1.93989
R998 VTAIL.n439 VTAIL.n428 1.93989
R999 VTAIL.n384 VTAIL.n383 1.93989
R1000 VTAIL.n372 VTAIL.n371 1.93989
R1001 VTAIL.n339 VTAIL.n328 1.93989
R1002 VTAIL.n0 VTAIL.t8 1.85264
R1003 VTAIL.n0 VTAIL.t11 1.85264
R1004 VTAIL.n198 VTAIL.t6 1.85264
R1005 VTAIL.n198 VTAIL.t3 1.85264
R1006 VTAIL.n594 VTAIL.t5 1.85264
R1007 VTAIL.n594 VTAIL.t1 1.85264
R1008 VTAIL.n396 VTAIL.t9 1.85264
R1009 VTAIL.n396 VTAIL.t10 1.85264
R1010 VTAIL.n397 VTAIL.n395 1.22464
R1011 VTAIL.n495 VTAIL.n397 1.22464
R1012 VTAIL.n595 VTAIL.n593 1.22464
R1013 VTAIL.n693 VTAIL.n595 1.22464
R1014 VTAIL.n297 VTAIL.n199 1.22464
R1015 VTAIL.n199 VTAIL.n197 1.22464
R1016 VTAIL.n99 VTAIL.n1 1.22464
R1017 VTAIL VTAIL.n791 1.16645
R1018 VTAIL.n730 VTAIL.n729 1.16414
R1019 VTAIL.n766 VTAIL.n704 1.16414
R1020 VTAIL.n776 VTAIL.n700 1.16414
R1021 VTAIL.n38 VTAIL.n37 1.16414
R1022 VTAIL.n74 VTAIL.n12 1.16414
R1023 VTAIL.n84 VTAIL.n8 1.16414
R1024 VTAIL.n136 VTAIL.n135 1.16414
R1025 VTAIL.n172 VTAIL.n110 1.16414
R1026 VTAIL.n182 VTAIL.n106 1.16414
R1027 VTAIL.n236 VTAIL.n235 1.16414
R1028 VTAIL.n272 VTAIL.n210 1.16414
R1029 VTAIL.n282 VTAIL.n206 1.16414
R1030 VTAIL.n678 VTAIL.n602 1.16414
R1031 VTAIL.n673 VTAIL.n607 1.16414
R1032 VTAIL.n634 VTAIL.n633 1.16414
R1033 VTAIL.n578 VTAIL.n502 1.16414
R1034 VTAIL.n573 VTAIL.n507 1.16414
R1035 VTAIL.n534 VTAIL.n533 1.16414
R1036 VTAIL.n480 VTAIL.n404 1.16414
R1037 VTAIL.n475 VTAIL.n409 1.16414
R1038 VTAIL.n436 VTAIL.n435 1.16414
R1039 VTAIL.n380 VTAIL.n304 1.16414
R1040 VTAIL.n375 VTAIL.n309 1.16414
R1041 VTAIL.n336 VTAIL.n335 1.16414
R1042 VTAIL.n593 VTAIL.n495 0.470328
R1043 VTAIL.n197 VTAIL.n99 0.470328
R1044 VTAIL.n726 VTAIL.n724 0.388379
R1045 VTAIL.n772 VTAIL.n771 0.388379
R1046 VTAIL.n775 VTAIL.n702 0.388379
R1047 VTAIL.n34 VTAIL.n32 0.388379
R1048 VTAIL.n80 VTAIL.n79 0.388379
R1049 VTAIL.n83 VTAIL.n10 0.388379
R1050 VTAIL.n132 VTAIL.n130 0.388379
R1051 VTAIL.n178 VTAIL.n177 0.388379
R1052 VTAIL.n181 VTAIL.n108 0.388379
R1053 VTAIL.n232 VTAIL.n230 0.388379
R1054 VTAIL.n278 VTAIL.n277 0.388379
R1055 VTAIL.n281 VTAIL.n208 0.388379
R1056 VTAIL.n677 VTAIL.n604 0.388379
R1057 VTAIL.n674 VTAIL.n606 0.388379
R1058 VTAIL.n630 VTAIL.n628 0.388379
R1059 VTAIL.n577 VTAIL.n504 0.388379
R1060 VTAIL.n574 VTAIL.n506 0.388379
R1061 VTAIL.n530 VTAIL.n528 0.388379
R1062 VTAIL.n479 VTAIL.n406 0.388379
R1063 VTAIL.n476 VTAIL.n408 0.388379
R1064 VTAIL.n432 VTAIL.n430 0.388379
R1065 VTAIL.n379 VTAIL.n306 0.388379
R1066 VTAIL.n376 VTAIL.n308 0.388379
R1067 VTAIL.n332 VTAIL.n330 0.388379
R1068 VTAIL.n731 VTAIL.n723 0.155672
R1069 VTAIL.n732 VTAIL.n731 0.155672
R1070 VTAIL.n732 VTAIL.n719 0.155672
R1071 VTAIL.n739 VTAIL.n719 0.155672
R1072 VTAIL.n740 VTAIL.n739 0.155672
R1073 VTAIL.n740 VTAIL.n715 0.155672
R1074 VTAIL.n747 VTAIL.n715 0.155672
R1075 VTAIL.n748 VTAIL.n747 0.155672
R1076 VTAIL.n748 VTAIL.n711 0.155672
R1077 VTAIL.n755 VTAIL.n711 0.155672
R1078 VTAIL.n756 VTAIL.n755 0.155672
R1079 VTAIL.n756 VTAIL.n707 0.155672
R1080 VTAIL.n763 VTAIL.n707 0.155672
R1081 VTAIL.n764 VTAIL.n763 0.155672
R1082 VTAIL.n764 VTAIL.n703 0.155672
R1083 VTAIL.n773 VTAIL.n703 0.155672
R1084 VTAIL.n774 VTAIL.n773 0.155672
R1085 VTAIL.n774 VTAIL.n699 0.155672
R1086 VTAIL.n781 VTAIL.n699 0.155672
R1087 VTAIL.n782 VTAIL.n781 0.155672
R1088 VTAIL.n782 VTAIL.n695 0.155672
R1089 VTAIL.n789 VTAIL.n695 0.155672
R1090 VTAIL.n39 VTAIL.n31 0.155672
R1091 VTAIL.n40 VTAIL.n39 0.155672
R1092 VTAIL.n40 VTAIL.n27 0.155672
R1093 VTAIL.n47 VTAIL.n27 0.155672
R1094 VTAIL.n48 VTAIL.n47 0.155672
R1095 VTAIL.n48 VTAIL.n23 0.155672
R1096 VTAIL.n55 VTAIL.n23 0.155672
R1097 VTAIL.n56 VTAIL.n55 0.155672
R1098 VTAIL.n56 VTAIL.n19 0.155672
R1099 VTAIL.n63 VTAIL.n19 0.155672
R1100 VTAIL.n64 VTAIL.n63 0.155672
R1101 VTAIL.n64 VTAIL.n15 0.155672
R1102 VTAIL.n71 VTAIL.n15 0.155672
R1103 VTAIL.n72 VTAIL.n71 0.155672
R1104 VTAIL.n72 VTAIL.n11 0.155672
R1105 VTAIL.n81 VTAIL.n11 0.155672
R1106 VTAIL.n82 VTAIL.n81 0.155672
R1107 VTAIL.n82 VTAIL.n7 0.155672
R1108 VTAIL.n89 VTAIL.n7 0.155672
R1109 VTAIL.n90 VTAIL.n89 0.155672
R1110 VTAIL.n90 VTAIL.n3 0.155672
R1111 VTAIL.n97 VTAIL.n3 0.155672
R1112 VTAIL.n137 VTAIL.n129 0.155672
R1113 VTAIL.n138 VTAIL.n137 0.155672
R1114 VTAIL.n138 VTAIL.n125 0.155672
R1115 VTAIL.n145 VTAIL.n125 0.155672
R1116 VTAIL.n146 VTAIL.n145 0.155672
R1117 VTAIL.n146 VTAIL.n121 0.155672
R1118 VTAIL.n153 VTAIL.n121 0.155672
R1119 VTAIL.n154 VTAIL.n153 0.155672
R1120 VTAIL.n154 VTAIL.n117 0.155672
R1121 VTAIL.n161 VTAIL.n117 0.155672
R1122 VTAIL.n162 VTAIL.n161 0.155672
R1123 VTAIL.n162 VTAIL.n113 0.155672
R1124 VTAIL.n169 VTAIL.n113 0.155672
R1125 VTAIL.n170 VTAIL.n169 0.155672
R1126 VTAIL.n170 VTAIL.n109 0.155672
R1127 VTAIL.n179 VTAIL.n109 0.155672
R1128 VTAIL.n180 VTAIL.n179 0.155672
R1129 VTAIL.n180 VTAIL.n105 0.155672
R1130 VTAIL.n187 VTAIL.n105 0.155672
R1131 VTAIL.n188 VTAIL.n187 0.155672
R1132 VTAIL.n188 VTAIL.n101 0.155672
R1133 VTAIL.n195 VTAIL.n101 0.155672
R1134 VTAIL.n237 VTAIL.n229 0.155672
R1135 VTAIL.n238 VTAIL.n237 0.155672
R1136 VTAIL.n238 VTAIL.n225 0.155672
R1137 VTAIL.n245 VTAIL.n225 0.155672
R1138 VTAIL.n246 VTAIL.n245 0.155672
R1139 VTAIL.n246 VTAIL.n221 0.155672
R1140 VTAIL.n253 VTAIL.n221 0.155672
R1141 VTAIL.n254 VTAIL.n253 0.155672
R1142 VTAIL.n254 VTAIL.n217 0.155672
R1143 VTAIL.n261 VTAIL.n217 0.155672
R1144 VTAIL.n262 VTAIL.n261 0.155672
R1145 VTAIL.n262 VTAIL.n213 0.155672
R1146 VTAIL.n269 VTAIL.n213 0.155672
R1147 VTAIL.n270 VTAIL.n269 0.155672
R1148 VTAIL.n270 VTAIL.n209 0.155672
R1149 VTAIL.n279 VTAIL.n209 0.155672
R1150 VTAIL.n280 VTAIL.n279 0.155672
R1151 VTAIL.n280 VTAIL.n205 0.155672
R1152 VTAIL.n287 VTAIL.n205 0.155672
R1153 VTAIL.n288 VTAIL.n287 0.155672
R1154 VTAIL.n288 VTAIL.n201 0.155672
R1155 VTAIL.n295 VTAIL.n201 0.155672
R1156 VTAIL.n691 VTAIL.n597 0.155672
R1157 VTAIL.n684 VTAIL.n597 0.155672
R1158 VTAIL.n684 VTAIL.n683 0.155672
R1159 VTAIL.n683 VTAIL.n601 0.155672
R1160 VTAIL.n676 VTAIL.n601 0.155672
R1161 VTAIL.n676 VTAIL.n675 0.155672
R1162 VTAIL.n675 VTAIL.n605 0.155672
R1163 VTAIL.n668 VTAIL.n605 0.155672
R1164 VTAIL.n668 VTAIL.n667 0.155672
R1165 VTAIL.n667 VTAIL.n611 0.155672
R1166 VTAIL.n660 VTAIL.n611 0.155672
R1167 VTAIL.n660 VTAIL.n659 0.155672
R1168 VTAIL.n659 VTAIL.n615 0.155672
R1169 VTAIL.n652 VTAIL.n615 0.155672
R1170 VTAIL.n652 VTAIL.n651 0.155672
R1171 VTAIL.n651 VTAIL.n619 0.155672
R1172 VTAIL.n644 VTAIL.n619 0.155672
R1173 VTAIL.n644 VTAIL.n643 0.155672
R1174 VTAIL.n643 VTAIL.n623 0.155672
R1175 VTAIL.n636 VTAIL.n623 0.155672
R1176 VTAIL.n636 VTAIL.n635 0.155672
R1177 VTAIL.n635 VTAIL.n627 0.155672
R1178 VTAIL.n591 VTAIL.n497 0.155672
R1179 VTAIL.n584 VTAIL.n497 0.155672
R1180 VTAIL.n584 VTAIL.n583 0.155672
R1181 VTAIL.n583 VTAIL.n501 0.155672
R1182 VTAIL.n576 VTAIL.n501 0.155672
R1183 VTAIL.n576 VTAIL.n575 0.155672
R1184 VTAIL.n575 VTAIL.n505 0.155672
R1185 VTAIL.n568 VTAIL.n505 0.155672
R1186 VTAIL.n568 VTAIL.n567 0.155672
R1187 VTAIL.n567 VTAIL.n511 0.155672
R1188 VTAIL.n560 VTAIL.n511 0.155672
R1189 VTAIL.n560 VTAIL.n559 0.155672
R1190 VTAIL.n559 VTAIL.n515 0.155672
R1191 VTAIL.n552 VTAIL.n515 0.155672
R1192 VTAIL.n552 VTAIL.n551 0.155672
R1193 VTAIL.n551 VTAIL.n519 0.155672
R1194 VTAIL.n544 VTAIL.n519 0.155672
R1195 VTAIL.n544 VTAIL.n543 0.155672
R1196 VTAIL.n543 VTAIL.n523 0.155672
R1197 VTAIL.n536 VTAIL.n523 0.155672
R1198 VTAIL.n536 VTAIL.n535 0.155672
R1199 VTAIL.n535 VTAIL.n527 0.155672
R1200 VTAIL.n493 VTAIL.n399 0.155672
R1201 VTAIL.n486 VTAIL.n399 0.155672
R1202 VTAIL.n486 VTAIL.n485 0.155672
R1203 VTAIL.n485 VTAIL.n403 0.155672
R1204 VTAIL.n478 VTAIL.n403 0.155672
R1205 VTAIL.n478 VTAIL.n477 0.155672
R1206 VTAIL.n477 VTAIL.n407 0.155672
R1207 VTAIL.n470 VTAIL.n407 0.155672
R1208 VTAIL.n470 VTAIL.n469 0.155672
R1209 VTAIL.n469 VTAIL.n413 0.155672
R1210 VTAIL.n462 VTAIL.n413 0.155672
R1211 VTAIL.n462 VTAIL.n461 0.155672
R1212 VTAIL.n461 VTAIL.n417 0.155672
R1213 VTAIL.n454 VTAIL.n417 0.155672
R1214 VTAIL.n454 VTAIL.n453 0.155672
R1215 VTAIL.n453 VTAIL.n421 0.155672
R1216 VTAIL.n446 VTAIL.n421 0.155672
R1217 VTAIL.n446 VTAIL.n445 0.155672
R1218 VTAIL.n445 VTAIL.n425 0.155672
R1219 VTAIL.n438 VTAIL.n425 0.155672
R1220 VTAIL.n438 VTAIL.n437 0.155672
R1221 VTAIL.n437 VTAIL.n429 0.155672
R1222 VTAIL.n393 VTAIL.n299 0.155672
R1223 VTAIL.n386 VTAIL.n299 0.155672
R1224 VTAIL.n386 VTAIL.n385 0.155672
R1225 VTAIL.n385 VTAIL.n303 0.155672
R1226 VTAIL.n378 VTAIL.n303 0.155672
R1227 VTAIL.n378 VTAIL.n377 0.155672
R1228 VTAIL.n377 VTAIL.n307 0.155672
R1229 VTAIL.n370 VTAIL.n307 0.155672
R1230 VTAIL.n370 VTAIL.n369 0.155672
R1231 VTAIL.n369 VTAIL.n313 0.155672
R1232 VTAIL.n362 VTAIL.n313 0.155672
R1233 VTAIL.n362 VTAIL.n361 0.155672
R1234 VTAIL.n361 VTAIL.n317 0.155672
R1235 VTAIL.n354 VTAIL.n317 0.155672
R1236 VTAIL.n354 VTAIL.n353 0.155672
R1237 VTAIL.n353 VTAIL.n321 0.155672
R1238 VTAIL.n346 VTAIL.n321 0.155672
R1239 VTAIL.n346 VTAIL.n345 0.155672
R1240 VTAIL.n345 VTAIL.n325 0.155672
R1241 VTAIL.n338 VTAIL.n325 0.155672
R1242 VTAIL.n338 VTAIL.n337 0.155672
R1243 VTAIL.n337 VTAIL.n329 0.155672
R1244 VTAIL VTAIL.n1 0.0586897
R1245 VDD2.n2 VDD2.n1 70.1606
R1246 VDD2.n2 VDD2.n0 70.1606
R1247 VDD2 VDD2.n5 70.1577
R1248 VDD2.n4 VDD2.n3 69.6041
R1249 VDD2.n4 VDD2.n2 44.3532
R1250 VDD2.n5 VDD2.t1 1.85264
R1251 VDD2.n5 VDD2.t2 1.85264
R1252 VDD2.n3 VDD2.t4 1.85264
R1253 VDD2.n3 VDD2.t6 1.85264
R1254 VDD2.n1 VDD2.t5 1.85264
R1255 VDD2.n1 VDD2.t0 1.85264
R1256 VDD2.n0 VDD2.t3 1.85264
R1257 VDD2.n0 VDD2.t7 1.85264
R1258 VDD2 VDD2.n4 0.670759
R1259 B.n142 B.t0 591.534
R1260 B.n150 B.t9 591.534
R1261 B.n46 B.t6 591.534
R1262 B.n52 B.t3 591.534
R1263 B.n514 B.n83 585
R1264 B.n516 B.n515 585
R1265 B.n517 B.n82 585
R1266 B.n519 B.n518 585
R1267 B.n520 B.n81 585
R1268 B.n522 B.n521 585
R1269 B.n523 B.n80 585
R1270 B.n525 B.n524 585
R1271 B.n526 B.n79 585
R1272 B.n528 B.n527 585
R1273 B.n529 B.n78 585
R1274 B.n531 B.n530 585
R1275 B.n532 B.n77 585
R1276 B.n534 B.n533 585
R1277 B.n535 B.n76 585
R1278 B.n537 B.n536 585
R1279 B.n538 B.n75 585
R1280 B.n540 B.n539 585
R1281 B.n541 B.n74 585
R1282 B.n543 B.n542 585
R1283 B.n544 B.n73 585
R1284 B.n546 B.n545 585
R1285 B.n547 B.n72 585
R1286 B.n549 B.n548 585
R1287 B.n550 B.n71 585
R1288 B.n552 B.n551 585
R1289 B.n553 B.n70 585
R1290 B.n555 B.n554 585
R1291 B.n556 B.n69 585
R1292 B.n558 B.n557 585
R1293 B.n559 B.n68 585
R1294 B.n561 B.n560 585
R1295 B.n562 B.n67 585
R1296 B.n564 B.n563 585
R1297 B.n565 B.n66 585
R1298 B.n567 B.n566 585
R1299 B.n568 B.n65 585
R1300 B.n570 B.n569 585
R1301 B.n571 B.n64 585
R1302 B.n573 B.n572 585
R1303 B.n574 B.n63 585
R1304 B.n576 B.n575 585
R1305 B.n577 B.n62 585
R1306 B.n579 B.n578 585
R1307 B.n580 B.n61 585
R1308 B.n582 B.n581 585
R1309 B.n583 B.n60 585
R1310 B.n585 B.n584 585
R1311 B.n586 B.n59 585
R1312 B.n588 B.n587 585
R1313 B.n589 B.n58 585
R1314 B.n591 B.n590 585
R1315 B.n592 B.n57 585
R1316 B.n594 B.n593 585
R1317 B.n595 B.n56 585
R1318 B.n597 B.n596 585
R1319 B.n598 B.n55 585
R1320 B.n600 B.n599 585
R1321 B.n602 B.n601 585
R1322 B.n603 B.n51 585
R1323 B.n605 B.n604 585
R1324 B.n606 B.n50 585
R1325 B.n608 B.n607 585
R1326 B.n609 B.n49 585
R1327 B.n611 B.n610 585
R1328 B.n612 B.n48 585
R1329 B.n614 B.n613 585
R1330 B.n616 B.n45 585
R1331 B.n618 B.n617 585
R1332 B.n619 B.n44 585
R1333 B.n621 B.n620 585
R1334 B.n622 B.n43 585
R1335 B.n624 B.n623 585
R1336 B.n625 B.n42 585
R1337 B.n627 B.n626 585
R1338 B.n628 B.n41 585
R1339 B.n630 B.n629 585
R1340 B.n631 B.n40 585
R1341 B.n633 B.n632 585
R1342 B.n634 B.n39 585
R1343 B.n636 B.n635 585
R1344 B.n637 B.n38 585
R1345 B.n639 B.n638 585
R1346 B.n640 B.n37 585
R1347 B.n642 B.n641 585
R1348 B.n643 B.n36 585
R1349 B.n645 B.n644 585
R1350 B.n646 B.n35 585
R1351 B.n648 B.n647 585
R1352 B.n649 B.n34 585
R1353 B.n651 B.n650 585
R1354 B.n652 B.n33 585
R1355 B.n654 B.n653 585
R1356 B.n655 B.n32 585
R1357 B.n657 B.n656 585
R1358 B.n658 B.n31 585
R1359 B.n660 B.n659 585
R1360 B.n661 B.n30 585
R1361 B.n663 B.n662 585
R1362 B.n664 B.n29 585
R1363 B.n666 B.n665 585
R1364 B.n667 B.n28 585
R1365 B.n669 B.n668 585
R1366 B.n670 B.n27 585
R1367 B.n672 B.n671 585
R1368 B.n673 B.n26 585
R1369 B.n675 B.n674 585
R1370 B.n676 B.n25 585
R1371 B.n678 B.n677 585
R1372 B.n679 B.n24 585
R1373 B.n681 B.n680 585
R1374 B.n682 B.n23 585
R1375 B.n684 B.n683 585
R1376 B.n685 B.n22 585
R1377 B.n687 B.n686 585
R1378 B.n688 B.n21 585
R1379 B.n690 B.n689 585
R1380 B.n691 B.n20 585
R1381 B.n693 B.n692 585
R1382 B.n694 B.n19 585
R1383 B.n696 B.n695 585
R1384 B.n697 B.n18 585
R1385 B.n699 B.n698 585
R1386 B.n700 B.n17 585
R1387 B.n702 B.n701 585
R1388 B.n513 B.n512 585
R1389 B.n511 B.n84 585
R1390 B.n510 B.n509 585
R1391 B.n508 B.n85 585
R1392 B.n507 B.n506 585
R1393 B.n505 B.n86 585
R1394 B.n504 B.n503 585
R1395 B.n502 B.n87 585
R1396 B.n501 B.n500 585
R1397 B.n499 B.n88 585
R1398 B.n498 B.n497 585
R1399 B.n496 B.n89 585
R1400 B.n495 B.n494 585
R1401 B.n493 B.n90 585
R1402 B.n492 B.n491 585
R1403 B.n490 B.n91 585
R1404 B.n489 B.n488 585
R1405 B.n487 B.n92 585
R1406 B.n486 B.n485 585
R1407 B.n484 B.n93 585
R1408 B.n483 B.n482 585
R1409 B.n481 B.n94 585
R1410 B.n480 B.n479 585
R1411 B.n478 B.n95 585
R1412 B.n477 B.n476 585
R1413 B.n475 B.n96 585
R1414 B.n474 B.n473 585
R1415 B.n472 B.n97 585
R1416 B.n471 B.n470 585
R1417 B.n469 B.n98 585
R1418 B.n468 B.n467 585
R1419 B.n466 B.n99 585
R1420 B.n465 B.n464 585
R1421 B.n463 B.n100 585
R1422 B.n462 B.n461 585
R1423 B.n460 B.n101 585
R1424 B.n459 B.n458 585
R1425 B.n457 B.n102 585
R1426 B.n456 B.n455 585
R1427 B.n454 B.n103 585
R1428 B.n453 B.n452 585
R1429 B.n451 B.n104 585
R1430 B.n450 B.n449 585
R1431 B.n448 B.n105 585
R1432 B.n447 B.n446 585
R1433 B.n445 B.n106 585
R1434 B.n444 B.n443 585
R1435 B.n442 B.n107 585
R1436 B.n441 B.n440 585
R1437 B.n439 B.n108 585
R1438 B.n438 B.n437 585
R1439 B.n436 B.n109 585
R1440 B.n435 B.n434 585
R1441 B.n433 B.n110 585
R1442 B.n432 B.n431 585
R1443 B.n430 B.n111 585
R1444 B.n429 B.n428 585
R1445 B.n427 B.n112 585
R1446 B.n426 B.n425 585
R1447 B.n237 B.n236 585
R1448 B.n238 B.n179 585
R1449 B.n240 B.n239 585
R1450 B.n241 B.n178 585
R1451 B.n243 B.n242 585
R1452 B.n244 B.n177 585
R1453 B.n246 B.n245 585
R1454 B.n247 B.n176 585
R1455 B.n249 B.n248 585
R1456 B.n250 B.n175 585
R1457 B.n252 B.n251 585
R1458 B.n253 B.n174 585
R1459 B.n255 B.n254 585
R1460 B.n256 B.n173 585
R1461 B.n258 B.n257 585
R1462 B.n259 B.n172 585
R1463 B.n261 B.n260 585
R1464 B.n262 B.n171 585
R1465 B.n264 B.n263 585
R1466 B.n265 B.n170 585
R1467 B.n267 B.n266 585
R1468 B.n268 B.n169 585
R1469 B.n270 B.n269 585
R1470 B.n271 B.n168 585
R1471 B.n273 B.n272 585
R1472 B.n274 B.n167 585
R1473 B.n276 B.n275 585
R1474 B.n277 B.n166 585
R1475 B.n279 B.n278 585
R1476 B.n280 B.n165 585
R1477 B.n282 B.n281 585
R1478 B.n283 B.n164 585
R1479 B.n285 B.n284 585
R1480 B.n286 B.n163 585
R1481 B.n288 B.n287 585
R1482 B.n289 B.n162 585
R1483 B.n291 B.n290 585
R1484 B.n292 B.n161 585
R1485 B.n294 B.n293 585
R1486 B.n295 B.n160 585
R1487 B.n297 B.n296 585
R1488 B.n298 B.n159 585
R1489 B.n300 B.n299 585
R1490 B.n301 B.n158 585
R1491 B.n303 B.n302 585
R1492 B.n304 B.n157 585
R1493 B.n306 B.n305 585
R1494 B.n307 B.n156 585
R1495 B.n309 B.n308 585
R1496 B.n310 B.n155 585
R1497 B.n312 B.n311 585
R1498 B.n313 B.n154 585
R1499 B.n315 B.n314 585
R1500 B.n316 B.n153 585
R1501 B.n318 B.n317 585
R1502 B.n319 B.n152 585
R1503 B.n321 B.n320 585
R1504 B.n322 B.n149 585
R1505 B.n325 B.n324 585
R1506 B.n326 B.n148 585
R1507 B.n328 B.n327 585
R1508 B.n329 B.n147 585
R1509 B.n331 B.n330 585
R1510 B.n332 B.n146 585
R1511 B.n334 B.n333 585
R1512 B.n335 B.n145 585
R1513 B.n337 B.n336 585
R1514 B.n339 B.n338 585
R1515 B.n340 B.n141 585
R1516 B.n342 B.n341 585
R1517 B.n343 B.n140 585
R1518 B.n345 B.n344 585
R1519 B.n346 B.n139 585
R1520 B.n348 B.n347 585
R1521 B.n349 B.n138 585
R1522 B.n351 B.n350 585
R1523 B.n352 B.n137 585
R1524 B.n354 B.n353 585
R1525 B.n355 B.n136 585
R1526 B.n357 B.n356 585
R1527 B.n358 B.n135 585
R1528 B.n360 B.n359 585
R1529 B.n361 B.n134 585
R1530 B.n363 B.n362 585
R1531 B.n364 B.n133 585
R1532 B.n366 B.n365 585
R1533 B.n367 B.n132 585
R1534 B.n369 B.n368 585
R1535 B.n370 B.n131 585
R1536 B.n372 B.n371 585
R1537 B.n373 B.n130 585
R1538 B.n375 B.n374 585
R1539 B.n376 B.n129 585
R1540 B.n378 B.n377 585
R1541 B.n379 B.n128 585
R1542 B.n381 B.n380 585
R1543 B.n382 B.n127 585
R1544 B.n384 B.n383 585
R1545 B.n385 B.n126 585
R1546 B.n387 B.n386 585
R1547 B.n388 B.n125 585
R1548 B.n390 B.n389 585
R1549 B.n391 B.n124 585
R1550 B.n393 B.n392 585
R1551 B.n394 B.n123 585
R1552 B.n396 B.n395 585
R1553 B.n397 B.n122 585
R1554 B.n399 B.n398 585
R1555 B.n400 B.n121 585
R1556 B.n402 B.n401 585
R1557 B.n403 B.n120 585
R1558 B.n405 B.n404 585
R1559 B.n406 B.n119 585
R1560 B.n408 B.n407 585
R1561 B.n409 B.n118 585
R1562 B.n411 B.n410 585
R1563 B.n412 B.n117 585
R1564 B.n414 B.n413 585
R1565 B.n415 B.n116 585
R1566 B.n417 B.n416 585
R1567 B.n418 B.n115 585
R1568 B.n420 B.n419 585
R1569 B.n421 B.n114 585
R1570 B.n423 B.n422 585
R1571 B.n424 B.n113 585
R1572 B.n235 B.n180 585
R1573 B.n234 B.n233 585
R1574 B.n232 B.n181 585
R1575 B.n231 B.n230 585
R1576 B.n229 B.n182 585
R1577 B.n228 B.n227 585
R1578 B.n226 B.n183 585
R1579 B.n225 B.n224 585
R1580 B.n223 B.n184 585
R1581 B.n222 B.n221 585
R1582 B.n220 B.n185 585
R1583 B.n219 B.n218 585
R1584 B.n217 B.n186 585
R1585 B.n216 B.n215 585
R1586 B.n214 B.n187 585
R1587 B.n213 B.n212 585
R1588 B.n211 B.n188 585
R1589 B.n210 B.n209 585
R1590 B.n208 B.n189 585
R1591 B.n207 B.n206 585
R1592 B.n205 B.n190 585
R1593 B.n204 B.n203 585
R1594 B.n202 B.n191 585
R1595 B.n201 B.n200 585
R1596 B.n199 B.n192 585
R1597 B.n198 B.n197 585
R1598 B.n196 B.n193 585
R1599 B.n195 B.n194 585
R1600 B.n2 B.n0 585
R1601 B.n745 B.n1 585
R1602 B.n744 B.n743 585
R1603 B.n742 B.n3 585
R1604 B.n741 B.n740 585
R1605 B.n739 B.n4 585
R1606 B.n738 B.n737 585
R1607 B.n736 B.n5 585
R1608 B.n735 B.n734 585
R1609 B.n733 B.n6 585
R1610 B.n732 B.n731 585
R1611 B.n730 B.n7 585
R1612 B.n729 B.n728 585
R1613 B.n727 B.n8 585
R1614 B.n726 B.n725 585
R1615 B.n724 B.n9 585
R1616 B.n723 B.n722 585
R1617 B.n721 B.n10 585
R1618 B.n720 B.n719 585
R1619 B.n718 B.n11 585
R1620 B.n717 B.n716 585
R1621 B.n715 B.n12 585
R1622 B.n714 B.n713 585
R1623 B.n712 B.n13 585
R1624 B.n711 B.n710 585
R1625 B.n709 B.n14 585
R1626 B.n708 B.n707 585
R1627 B.n706 B.n15 585
R1628 B.n705 B.n704 585
R1629 B.n703 B.n16 585
R1630 B.n747 B.n746 585
R1631 B.n236 B.n235 535.745
R1632 B.n703 B.n702 535.745
R1633 B.n426 B.n113 535.745
R1634 B.n512 B.n83 535.745
R1635 B.n142 B.t2 503.187
R1636 B.n52 B.t4 503.187
R1637 B.n150 B.t11 503.185
R1638 B.n46 B.t7 503.185
R1639 B.n143 B.t1 475.647
R1640 B.n53 B.t5 475.647
R1641 B.n151 B.t10 475.647
R1642 B.n47 B.t8 475.647
R1643 B.n235 B.n234 163.367
R1644 B.n234 B.n181 163.367
R1645 B.n230 B.n181 163.367
R1646 B.n230 B.n229 163.367
R1647 B.n229 B.n228 163.367
R1648 B.n228 B.n183 163.367
R1649 B.n224 B.n183 163.367
R1650 B.n224 B.n223 163.367
R1651 B.n223 B.n222 163.367
R1652 B.n222 B.n185 163.367
R1653 B.n218 B.n185 163.367
R1654 B.n218 B.n217 163.367
R1655 B.n217 B.n216 163.367
R1656 B.n216 B.n187 163.367
R1657 B.n212 B.n187 163.367
R1658 B.n212 B.n211 163.367
R1659 B.n211 B.n210 163.367
R1660 B.n210 B.n189 163.367
R1661 B.n206 B.n189 163.367
R1662 B.n206 B.n205 163.367
R1663 B.n205 B.n204 163.367
R1664 B.n204 B.n191 163.367
R1665 B.n200 B.n191 163.367
R1666 B.n200 B.n199 163.367
R1667 B.n199 B.n198 163.367
R1668 B.n198 B.n193 163.367
R1669 B.n194 B.n193 163.367
R1670 B.n194 B.n2 163.367
R1671 B.n746 B.n2 163.367
R1672 B.n746 B.n745 163.367
R1673 B.n745 B.n744 163.367
R1674 B.n744 B.n3 163.367
R1675 B.n740 B.n3 163.367
R1676 B.n740 B.n739 163.367
R1677 B.n739 B.n738 163.367
R1678 B.n738 B.n5 163.367
R1679 B.n734 B.n5 163.367
R1680 B.n734 B.n733 163.367
R1681 B.n733 B.n732 163.367
R1682 B.n732 B.n7 163.367
R1683 B.n728 B.n7 163.367
R1684 B.n728 B.n727 163.367
R1685 B.n727 B.n726 163.367
R1686 B.n726 B.n9 163.367
R1687 B.n722 B.n9 163.367
R1688 B.n722 B.n721 163.367
R1689 B.n721 B.n720 163.367
R1690 B.n720 B.n11 163.367
R1691 B.n716 B.n11 163.367
R1692 B.n716 B.n715 163.367
R1693 B.n715 B.n714 163.367
R1694 B.n714 B.n13 163.367
R1695 B.n710 B.n13 163.367
R1696 B.n710 B.n709 163.367
R1697 B.n709 B.n708 163.367
R1698 B.n708 B.n15 163.367
R1699 B.n704 B.n15 163.367
R1700 B.n704 B.n703 163.367
R1701 B.n236 B.n179 163.367
R1702 B.n240 B.n179 163.367
R1703 B.n241 B.n240 163.367
R1704 B.n242 B.n241 163.367
R1705 B.n242 B.n177 163.367
R1706 B.n246 B.n177 163.367
R1707 B.n247 B.n246 163.367
R1708 B.n248 B.n247 163.367
R1709 B.n248 B.n175 163.367
R1710 B.n252 B.n175 163.367
R1711 B.n253 B.n252 163.367
R1712 B.n254 B.n253 163.367
R1713 B.n254 B.n173 163.367
R1714 B.n258 B.n173 163.367
R1715 B.n259 B.n258 163.367
R1716 B.n260 B.n259 163.367
R1717 B.n260 B.n171 163.367
R1718 B.n264 B.n171 163.367
R1719 B.n265 B.n264 163.367
R1720 B.n266 B.n265 163.367
R1721 B.n266 B.n169 163.367
R1722 B.n270 B.n169 163.367
R1723 B.n271 B.n270 163.367
R1724 B.n272 B.n271 163.367
R1725 B.n272 B.n167 163.367
R1726 B.n276 B.n167 163.367
R1727 B.n277 B.n276 163.367
R1728 B.n278 B.n277 163.367
R1729 B.n278 B.n165 163.367
R1730 B.n282 B.n165 163.367
R1731 B.n283 B.n282 163.367
R1732 B.n284 B.n283 163.367
R1733 B.n284 B.n163 163.367
R1734 B.n288 B.n163 163.367
R1735 B.n289 B.n288 163.367
R1736 B.n290 B.n289 163.367
R1737 B.n290 B.n161 163.367
R1738 B.n294 B.n161 163.367
R1739 B.n295 B.n294 163.367
R1740 B.n296 B.n295 163.367
R1741 B.n296 B.n159 163.367
R1742 B.n300 B.n159 163.367
R1743 B.n301 B.n300 163.367
R1744 B.n302 B.n301 163.367
R1745 B.n302 B.n157 163.367
R1746 B.n306 B.n157 163.367
R1747 B.n307 B.n306 163.367
R1748 B.n308 B.n307 163.367
R1749 B.n308 B.n155 163.367
R1750 B.n312 B.n155 163.367
R1751 B.n313 B.n312 163.367
R1752 B.n314 B.n313 163.367
R1753 B.n314 B.n153 163.367
R1754 B.n318 B.n153 163.367
R1755 B.n319 B.n318 163.367
R1756 B.n320 B.n319 163.367
R1757 B.n320 B.n149 163.367
R1758 B.n325 B.n149 163.367
R1759 B.n326 B.n325 163.367
R1760 B.n327 B.n326 163.367
R1761 B.n327 B.n147 163.367
R1762 B.n331 B.n147 163.367
R1763 B.n332 B.n331 163.367
R1764 B.n333 B.n332 163.367
R1765 B.n333 B.n145 163.367
R1766 B.n337 B.n145 163.367
R1767 B.n338 B.n337 163.367
R1768 B.n338 B.n141 163.367
R1769 B.n342 B.n141 163.367
R1770 B.n343 B.n342 163.367
R1771 B.n344 B.n343 163.367
R1772 B.n344 B.n139 163.367
R1773 B.n348 B.n139 163.367
R1774 B.n349 B.n348 163.367
R1775 B.n350 B.n349 163.367
R1776 B.n350 B.n137 163.367
R1777 B.n354 B.n137 163.367
R1778 B.n355 B.n354 163.367
R1779 B.n356 B.n355 163.367
R1780 B.n356 B.n135 163.367
R1781 B.n360 B.n135 163.367
R1782 B.n361 B.n360 163.367
R1783 B.n362 B.n361 163.367
R1784 B.n362 B.n133 163.367
R1785 B.n366 B.n133 163.367
R1786 B.n367 B.n366 163.367
R1787 B.n368 B.n367 163.367
R1788 B.n368 B.n131 163.367
R1789 B.n372 B.n131 163.367
R1790 B.n373 B.n372 163.367
R1791 B.n374 B.n373 163.367
R1792 B.n374 B.n129 163.367
R1793 B.n378 B.n129 163.367
R1794 B.n379 B.n378 163.367
R1795 B.n380 B.n379 163.367
R1796 B.n380 B.n127 163.367
R1797 B.n384 B.n127 163.367
R1798 B.n385 B.n384 163.367
R1799 B.n386 B.n385 163.367
R1800 B.n386 B.n125 163.367
R1801 B.n390 B.n125 163.367
R1802 B.n391 B.n390 163.367
R1803 B.n392 B.n391 163.367
R1804 B.n392 B.n123 163.367
R1805 B.n396 B.n123 163.367
R1806 B.n397 B.n396 163.367
R1807 B.n398 B.n397 163.367
R1808 B.n398 B.n121 163.367
R1809 B.n402 B.n121 163.367
R1810 B.n403 B.n402 163.367
R1811 B.n404 B.n403 163.367
R1812 B.n404 B.n119 163.367
R1813 B.n408 B.n119 163.367
R1814 B.n409 B.n408 163.367
R1815 B.n410 B.n409 163.367
R1816 B.n410 B.n117 163.367
R1817 B.n414 B.n117 163.367
R1818 B.n415 B.n414 163.367
R1819 B.n416 B.n415 163.367
R1820 B.n416 B.n115 163.367
R1821 B.n420 B.n115 163.367
R1822 B.n421 B.n420 163.367
R1823 B.n422 B.n421 163.367
R1824 B.n422 B.n113 163.367
R1825 B.n427 B.n426 163.367
R1826 B.n428 B.n427 163.367
R1827 B.n428 B.n111 163.367
R1828 B.n432 B.n111 163.367
R1829 B.n433 B.n432 163.367
R1830 B.n434 B.n433 163.367
R1831 B.n434 B.n109 163.367
R1832 B.n438 B.n109 163.367
R1833 B.n439 B.n438 163.367
R1834 B.n440 B.n439 163.367
R1835 B.n440 B.n107 163.367
R1836 B.n444 B.n107 163.367
R1837 B.n445 B.n444 163.367
R1838 B.n446 B.n445 163.367
R1839 B.n446 B.n105 163.367
R1840 B.n450 B.n105 163.367
R1841 B.n451 B.n450 163.367
R1842 B.n452 B.n451 163.367
R1843 B.n452 B.n103 163.367
R1844 B.n456 B.n103 163.367
R1845 B.n457 B.n456 163.367
R1846 B.n458 B.n457 163.367
R1847 B.n458 B.n101 163.367
R1848 B.n462 B.n101 163.367
R1849 B.n463 B.n462 163.367
R1850 B.n464 B.n463 163.367
R1851 B.n464 B.n99 163.367
R1852 B.n468 B.n99 163.367
R1853 B.n469 B.n468 163.367
R1854 B.n470 B.n469 163.367
R1855 B.n470 B.n97 163.367
R1856 B.n474 B.n97 163.367
R1857 B.n475 B.n474 163.367
R1858 B.n476 B.n475 163.367
R1859 B.n476 B.n95 163.367
R1860 B.n480 B.n95 163.367
R1861 B.n481 B.n480 163.367
R1862 B.n482 B.n481 163.367
R1863 B.n482 B.n93 163.367
R1864 B.n486 B.n93 163.367
R1865 B.n487 B.n486 163.367
R1866 B.n488 B.n487 163.367
R1867 B.n488 B.n91 163.367
R1868 B.n492 B.n91 163.367
R1869 B.n493 B.n492 163.367
R1870 B.n494 B.n493 163.367
R1871 B.n494 B.n89 163.367
R1872 B.n498 B.n89 163.367
R1873 B.n499 B.n498 163.367
R1874 B.n500 B.n499 163.367
R1875 B.n500 B.n87 163.367
R1876 B.n504 B.n87 163.367
R1877 B.n505 B.n504 163.367
R1878 B.n506 B.n505 163.367
R1879 B.n506 B.n85 163.367
R1880 B.n510 B.n85 163.367
R1881 B.n511 B.n510 163.367
R1882 B.n512 B.n511 163.367
R1883 B.n702 B.n17 163.367
R1884 B.n698 B.n17 163.367
R1885 B.n698 B.n697 163.367
R1886 B.n697 B.n696 163.367
R1887 B.n696 B.n19 163.367
R1888 B.n692 B.n19 163.367
R1889 B.n692 B.n691 163.367
R1890 B.n691 B.n690 163.367
R1891 B.n690 B.n21 163.367
R1892 B.n686 B.n21 163.367
R1893 B.n686 B.n685 163.367
R1894 B.n685 B.n684 163.367
R1895 B.n684 B.n23 163.367
R1896 B.n680 B.n23 163.367
R1897 B.n680 B.n679 163.367
R1898 B.n679 B.n678 163.367
R1899 B.n678 B.n25 163.367
R1900 B.n674 B.n25 163.367
R1901 B.n674 B.n673 163.367
R1902 B.n673 B.n672 163.367
R1903 B.n672 B.n27 163.367
R1904 B.n668 B.n27 163.367
R1905 B.n668 B.n667 163.367
R1906 B.n667 B.n666 163.367
R1907 B.n666 B.n29 163.367
R1908 B.n662 B.n29 163.367
R1909 B.n662 B.n661 163.367
R1910 B.n661 B.n660 163.367
R1911 B.n660 B.n31 163.367
R1912 B.n656 B.n31 163.367
R1913 B.n656 B.n655 163.367
R1914 B.n655 B.n654 163.367
R1915 B.n654 B.n33 163.367
R1916 B.n650 B.n33 163.367
R1917 B.n650 B.n649 163.367
R1918 B.n649 B.n648 163.367
R1919 B.n648 B.n35 163.367
R1920 B.n644 B.n35 163.367
R1921 B.n644 B.n643 163.367
R1922 B.n643 B.n642 163.367
R1923 B.n642 B.n37 163.367
R1924 B.n638 B.n37 163.367
R1925 B.n638 B.n637 163.367
R1926 B.n637 B.n636 163.367
R1927 B.n636 B.n39 163.367
R1928 B.n632 B.n39 163.367
R1929 B.n632 B.n631 163.367
R1930 B.n631 B.n630 163.367
R1931 B.n630 B.n41 163.367
R1932 B.n626 B.n41 163.367
R1933 B.n626 B.n625 163.367
R1934 B.n625 B.n624 163.367
R1935 B.n624 B.n43 163.367
R1936 B.n620 B.n43 163.367
R1937 B.n620 B.n619 163.367
R1938 B.n619 B.n618 163.367
R1939 B.n618 B.n45 163.367
R1940 B.n613 B.n45 163.367
R1941 B.n613 B.n612 163.367
R1942 B.n612 B.n611 163.367
R1943 B.n611 B.n49 163.367
R1944 B.n607 B.n49 163.367
R1945 B.n607 B.n606 163.367
R1946 B.n606 B.n605 163.367
R1947 B.n605 B.n51 163.367
R1948 B.n601 B.n51 163.367
R1949 B.n601 B.n600 163.367
R1950 B.n600 B.n55 163.367
R1951 B.n596 B.n55 163.367
R1952 B.n596 B.n595 163.367
R1953 B.n595 B.n594 163.367
R1954 B.n594 B.n57 163.367
R1955 B.n590 B.n57 163.367
R1956 B.n590 B.n589 163.367
R1957 B.n589 B.n588 163.367
R1958 B.n588 B.n59 163.367
R1959 B.n584 B.n59 163.367
R1960 B.n584 B.n583 163.367
R1961 B.n583 B.n582 163.367
R1962 B.n582 B.n61 163.367
R1963 B.n578 B.n61 163.367
R1964 B.n578 B.n577 163.367
R1965 B.n577 B.n576 163.367
R1966 B.n576 B.n63 163.367
R1967 B.n572 B.n63 163.367
R1968 B.n572 B.n571 163.367
R1969 B.n571 B.n570 163.367
R1970 B.n570 B.n65 163.367
R1971 B.n566 B.n65 163.367
R1972 B.n566 B.n565 163.367
R1973 B.n565 B.n564 163.367
R1974 B.n564 B.n67 163.367
R1975 B.n560 B.n67 163.367
R1976 B.n560 B.n559 163.367
R1977 B.n559 B.n558 163.367
R1978 B.n558 B.n69 163.367
R1979 B.n554 B.n69 163.367
R1980 B.n554 B.n553 163.367
R1981 B.n553 B.n552 163.367
R1982 B.n552 B.n71 163.367
R1983 B.n548 B.n71 163.367
R1984 B.n548 B.n547 163.367
R1985 B.n547 B.n546 163.367
R1986 B.n546 B.n73 163.367
R1987 B.n542 B.n73 163.367
R1988 B.n542 B.n541 163.367
R1989 B.n541 B.n540 163.367
R1990 B.n540 B.n75 163.367
R1991 B.n536 B.n75 163.367
R1992 B.n536 B.n535 163.367
R1993 B.n535 B.n534 163.367
R1994 B.n534 B.n77 163.367
R1995 B.n530 B.n77 163.367
R1996 B.n530 B.n529 163.367
R1997 B.n529 B.n528 163.367
R1998 B.n528 B.n79 163.367
R1999 B.n524 B.n79 163.367
R2000 B.n524 B.n523 163.367
R2001 B.n523 B.n522 163.367
R2002 B.n522 B.n81 163.367
R2003 B.n518 B.n81 163.367
R2004 B.n518 B.n517 163.367
R2005 B.n517 B.n516 163.367
R2006 B.n516 B.n83 163.367
R2007 B.n144 B.n143 59.5399
R2008 B.n323 B.n151 59.5399
R2009 B.n615 B.n47 59.5399
R2010 B.n54 B.n53 59.5399
R2011 B.n701 B.n16 34.8103
R2012 B.n514 B.n513 34.8103
R2013 B.n425 B.n424 34.8103
R2014 B.n237 B.n180 34.8103
R2015 B.n143 B.n142 27.5399
R2016 B.n151 B.n150 27.5399
R2017 B.n47 B.n46 27.5399
R2018 B.n53 B.n52 27.5399
R2019 B B.n747 18.0485
R2020 B.n701 B.n700 10.6151
R2021 B.n700 B.n699 10.6151
R2022 B.n699 B.n18 10.6151
R2023 B.n695 B.n18 10.6151
R2024 B.n695 B.n694 10.6151
R2025 B.n694 B.n693 10.6151
R2026 B.n693 B.n20 10.6151
R2027 B.n689 B.n20 10.6151
R2028 B.n689 B.n688 10.6151
R2029 B.n688 B.n687 10.6151
R2030 B.n687 B.n22 10.6151
R2031 B.n683 B.n22 10.6151
R2032 B.n683 B.n682 10.6151
R2033 B.n682 B.n681 10.6151
R2034 B.n681 B.n24 10.6151
R2035 B.n677 B.n24 10.6151
R2036 B.n677 B.n676 10.6151
R2037 B.n676 B.n675 10.6151
R2038 B.n675 B.n26 10.6151
R2039 B.n671 B.n26 10.6151
R2040 B.n671 B.n670 10.6151
R2041 B.n670 B.n669 10.6151
R2042 B.n669 B.n28 10.6151
R2043 B.n665 B.n28 10.6151
R2044 B.n665 B.n664 10.6151
R2045 B.n664 B.n663 10.6151
R2046 B.n663 B.n30 10.6151
R2047 B.n659 B.n30 10.6151
R2048 B.n659 B.n658 10.6151
R2049 B.n658 B.n657 10.6151
R2050 B.n657 B.n32 10.6151
R2051 B.n653 B.n32 10.6151
R2052 B.n653 B.n652 10.6151
R2053 B.n652 B.n651 10.6151
R2054 B.n651 B.n34 10.6151
R2055 B.n647 B.n34 10.6151
R2056 B.n647 B.n646 10.6151
R2057 B.n646 B.n645 10.6151
R2058 B.n645 B.n36 10.6151
R2059 B.n641 B.n36 10.6151
R2060 B.n641 B.n640 10.6151
R2061 B.n640 B.n639 10.6151
R2062 B.n639 B.n38 10.6151
R2063 B.n635 B.n38 10.6151
R2064 B.n635 B.n634 10.6151
R2065 B.n634 B.n633 10.6151
R2066 B.n633 B.n40 10.6151
R2067 B.n629 B.n40 10.6151
R2068 B.n629 B.n628 10.6151
R2069 B.n628 B.n627 10.6151
R2070 B.n627 B.n42 10.6151
R2071 B.n623 B.n42 10.6151
R2072 B.n623 B.n622 10.6151
R2073 B.n622 B.n621 10.6151
R2074 B.n621 B.n44 10.6151
R2075 B.n617 B.n44 10.6151
R2076 B.n617 B.n616 10.6151
R2077 B.n614 B.n48 10.6151
R2078 B.n610 B.n48 10.6151
R2079 B.n610 B.n609 10.6151
R2080 B.n609 B.n608 10.6151
R2081 B.n608 B.n50 10.6151
R2082 B.n604 B.n50 10.6151
R2083 B.n604 B.n603 10.6151
R2084 B.n603 B.n602 10.6151
R2085 B.n599 B.n598 10.6151
R2086 B.n598 B.n597 10.6151
R2087 B.n597 B.n56 10.6151
R2088 B.n593 B.n56 10.6151
R2089 B.n593 B.n592 10.6151
R2090 B.n592 B.n591 10.6151
R2091 B.n591 B.n58 10.6151
R2092 B.n587 B.n58 10.6151
R2093 B.n587 B.n586 10.6151
R2094 B.n586 B.n585 10.6151
R2095 B.n585 B.n60 10.6151
R2096 B.n581 B.n60 10.6151
R2097 B.n581 B.n580 10.6151
R2098 B.n580 B.n579 10.6151
R2099 B.n579 B.n62 10.6151
R2100 B.n575 B.n62 10.6151
R2101 B.n575 B.n574 10.6151
R2102 B.n574 B.n573 10.6151
R2103 B.n573 B.n64 10.6151
R2104 B.n569 B.n64 10.6151
R2105 B.n569 B.n568 10.6151
R2106 B.n568 B.n567 10.6151
R2107 B.n567 B.n66 10.6151
R2108 B.n563 B.n66 10.6151
R2109 B.n563 B.n562 10.6151
R2110 B.n562 B.n561 10.6151
R2111 B.n561 B.n68 10.6151
R2112 B.n557 B.n68 10.6151
R2113 B.n557 B.n556 10.6151
R2114 B.n556 B.n555 10.6151
R2115 B.n555 B.n70 10.6151
R2116 B.n551 B.n70 10.6151
R2117 B.n551 B.n550 10.6151
R2118 B.n550 B.n549 10.6151
R2119 B.n549 B.n72 10.6151
R2120 B.n545 B.n72 10.6151
R2121 B.n545 B.n544 10.6151
R2122 B.n544 B.n543 10.6151
R2123 B.n543 B.n74 10.6151
R2124 B.n539 B.n74 10.6151
R2125 B.n539 B.n538 10.6151
R2126 B.n538 B.n537 10.6151
R2127 B.n537 B.n76 10.6151
R2128 B.n533 B.n76 10.6151
R2129 B.n533 B.n532 10.6151
R2130 B.n532 B.n531 10.6151
R2131 B.n531 B.n78 10.6151
R2132 B.n527 B.n78 10.6151
R2133 B.n527 B.n526 10.6151
R2134 B.n526 B.n525 10.6151
R2135 B.n525 B.n80 10.6151
R2136 B.n521 B.n80 10.6151
R2137 B.n521 B.n520 10.6151
R2138 B.n520 B.n519 10.6151
R2139 B.n519 B.n82 10.6151
R2140 B.n515 B.n82 10.6151
R2141 B.n515 B.n514 10.6151
R2142 B.n425 B.n112 10.6151
R2143 B.n429 B.n112 10.6151
R2144 B.n430 B.n429 10.6151
R2145 B.n431 B.n430 10.6151
R2146 B.n431 B.n110 10.6151
R2147 B.n435 B.n110 10.6151
R2148 B.n436 B.n435 10.6151
R2149 B.n437 B.n436 10.6151
R2150 B.n437 B.n108 10.6151
R2151 B.n441 B.n108 10.6151
R2152 B.n442 B.n441 10.6151
R2153 B.n443 B.n442 10.6151
R2154 B.n443 B.n106 10.6151
R2155 B.n447 B.n106 10.6151
R2156 B.n448 B.n447 10.6151
R2157 B.n449 B.n448 10.6151
R2158 B.n449 B.n104 10.6151
R2159 B.n453 B.n104 10.6151
R2160 B.n454 B.n453 10.6151
R2161 B.n455 B.n454 10.6151
R2162 B.n455 B.n102 10.6151
R2163 B.n459 B.n102 10.6151
R2164 B.n460 B.n459 10.6151
R2165 B.n461 B.n460 10.6151
R2166 B.n461 B.n100 10.6151
R2167 B.n465 B.n100 10.6151
R2168 B.n466 B.n465 10.6151
R2169 B.n467 B.n466 10.6151
R2170 B.n467 B.n98 10.6151
R2171 B.n471 B.n98 10.6151
R2172 B.n472 B.n471 10.6151
R2173 B.n473 B.n472 10.6151
R2174 B.n473 B.n96 10.6151
R2175 B.n477 B.n96 10.6151
R2176 B.n478 B.n477 10.6151
R2177 B.n479 B.n478 10.6151
R2178 B.n479 B.n94 10.6151
R2179 B.n483 B.n94 10.6151
R2180 B.n484 B.n483 10.6151
R2181 B.n485 B.n484 10.6151
R2182 B.n485 B.n92 10.6151
R2183 B.n489 B.n92 10.6151
R2184 B.n490 B.n489 10.6151
R2185 B.n491 B.n490 10.6151
R2186 B.n491 B.n90 10.6151
R2187 B.n495 B.n90 10.6151
R2188 B.n496 B.n495 10.6151
R2189 B.n497 B.n496 10.6151
R2190 B.n497 B.n88 10.6151
R2191 B.n501 B.n88 10.6151
R2192 B.n502 B.n501 10.6151
R2193 B.n503 B.n502 10.6151
R2194 B.n503 B.n86 10.6151
R2195 B.n507 B.n86 10.6151
R2196 B.n508 B.n507 10.6151
R2197 B.n509 B.n508 10.6151
R2198 B.n509 B.n84 10.6151
R2199 B.n513 B.n84 10.6151
R2200 B.n238 B.n237 10.6151
R2201 B.n239 B.n238 10.6151
R2202 B.n239 B.n178 10.6151
R2203 B.n243 B.n178 10.6151
R2204 B.n244 B.n243 10.6151
R2205 B.n245 B.n244 10.6151
R2206 B.n245 B.n176 10.6151
R2207 B.n249 B.n176 10.6151
R2208 B.n250 B.n249 10.6151
R2209 B.n251 B.n250 10.6151
R2210 B.n251 B.n174 10.6151
R2211 B.n255 B.n174 10.6151
R2212 B.n256 B.n255 10.6151
R2213 B.n257 B.n256 10.6151
R2214 B.n257 B.n172 10.6151
R2215 B.n261 B.n172 10.6151
R2216 B.n262 B.n261 10.6151
R2217 B.n263 B.n262 10.6151
R2218 B.n263 B.n170 10.6151
R2219 B.n267 B.n170 10.6151
R2220 B.n268 B.n267 10.6151
R2221 B.n269 B.n268 10.6151
R2222 B.n269 B.n168 10.6151
R2223 B.n273 B.n168 10.6151
R2224 B.n274 B.n273 10.6151
R2225 B.n275 B.n274 10.6151
R2226 B.n275 B.n166 10.6151
R2227 B.n279 B.n166 10.6151
R2228 B.n280 B.n279 10.6151
R2229 B.n281 B.n280 10.6151
R2230 B.n281 B.n164 10.6151
R2231 B.n285 B.n164 10.6151
R2232 B.n286 B.n285 10.6151
R2233 B.n287 B.n286 10.6151
R2234 B.n287 B.n162 10.6151
R2235 B.n291 B.n162 10.6151
R2236 B.n292 B.n291 10.6151
R2237 B.n293 B.n292 10.6151
R2238 B.n293 B.n160 10.6151
R2239 B.n297 B.n160 10.6151
R2240 B.n298 B.n297 10.6151
R2241 B.n299 B.n298 10.6151
R2242 B.n299 B.n158 10.6151
R2243 B.n303 B.n158 10.6151
R2244 B.n304 B.n303 10.6151
R2245 B.n305 B.n304 10.6151
R2246 B.n305 B.n156 10.6151
R2247 B.n309 B.n156 10.6151
R2248 B.n310 B.n309 10.6151
R2249 B.n311 B.n310 10.6151
R2250 B.n311 B.n154 10.6151
R2251 B.n315 B.n154 10.6151
R2252 B.n316 B.n315 10.6151
R2253 B.n317 B.n316 10.6151
R2254 B.n317 B.n152 10.6151
R2255 B.n321 B.n152 10.6151
R2256 B.n322 B.n321 10.6151
R2257 B.n324 B.n148 10.6151
R2258 B.n328 B.n148 10.6151
R2259 B.n329 B.n328 10.6151
R2260 B.n330 B.n329 10.6151
R2261 B.n330 B.n146 10.6151
R2262 B.n334 B.n146 10.6151
R2263 B.n335 B.n334 10.6151
R2264 B.n336 B.n335 10.6151
R2265 B.n340 B.n339 10.6151
R2266 B.n341 B.n340 10.6151
R2267 B.n341 B.n140 10.6151
R2268 B.n345 B.n140 10.6151
R2269 B.n346 B.n345 10.6151
R2270 B.n347 B.n346 10.6151
R2271 B.n347 B.n138 10.6151
R2272 B.n351 B.n138 10.6151
R2273 B.n352 B.n351 10.6151
R2274 B.n353 B.n352 10.6151
R2275 B.n353 B.n136 10.6151
R2276 B.n357 B.n136 10.6151
R2277 B.n358 B.n357 10.6151
R2278 B.n359 B.n358 10.6151
R2279 B.n359 B.n134 10.6151
R2280 B.n363 B.n134 10.6151
R2281 B.n364 B.n363 10.6151
R2282 B.n365 B.n364 10.6151
R2283 B.n365 B.n132 10.6151
R2284 B.n369 B.n132 10.6151
R2285 B.n370 B.n369 10.6151
R2286 B.n371 B.n370 10.6151
R2287 B.n371 B.n130 10.6151
R2288 B.n375 B.n130 10.6151
R2289 B.n376 B.n375 10.6151
R2290 B.n377 B.n376 10.6151
R2291 B.n377 B.n128 10.6151
R2292 B.n381 B.n128 10.6151
R2293 B.n382 B.n381 10.6151
R2294 B.n383 B.n382 10.6151
R2295 B.n383 B.n126 10.6151
R2296 B.n387 B.n126 10.6151
R2297 B.n388 B.n387 10.6151
R2298 B.n389 B.n388 10.6151
R2299 B.n389 B.n124 10.6151
R2300 B.n393 B.n124 10.6151
R2301 B.n394 B.n393 10.6151
R2302 B.n395 B.n394 10.6151
R2303 B.n395 B.n122 10.6151
R2304 B.n399 B.n122 10.6151
R2305 B.n400 B.n399 10.6151
R2306 B.n401 B.n400 10.6151
R2307 B.n401 B.n120 10.6151
R2308 B.n405 B.n120 10.6151
R2309 B.n406 B.n405 10.6151
R2310 B.n407 B.n406 10.6151
R2311 B.n407 B.n118 10.6151
R2312 B.n411 B.n118 10.6151
R2313 B.n412 B.n411 10.6151
R2314 B.n413 B.n412 10.6151
R2315 B.n413 B.n116 10.6151
R2316 B.n417 B.n116 10.6151
R2317 B.n418 B.n417 10.6151
R2318 B.n419 B.n418 10.6151
R2319 B.n419 B.n114 10.6151
R2320 B.n423 B.n114 10.6151
R2321 B.n424 B.n423 10.6151
R2322 B.n233 B.n180 10.6151
R2323 B.n233 B.n232 10.6151
R2324 B.n232 B.n231 10.6151
R2325 B.n231 B.n182 10.6151
R2326 B.n227 B.n182 10.6151
R2327 B.n227 B.n226 10.6151
R2328 B.n226 B.n225 10.6151
R2329 B.n225 B.n184 10.6151
R2330 B.n221 B.n184 10.6151
R2331 B.n221 B.n220 10.6151
R2332 B.n220 B.n219 10.6151
R2333 B.n219 B.n186 10.6151
R2334 B.n215 B.n186 10.6151
R2335 B.n215 B.n214 10.6151
R2336 B.n214 B.n213 10.6151
R2337 B.n213 B.n188 10.6151
R2338 B.n209 B.n188 10.6151
R2339 B.n209 B.n208 10.6151
R2340 B.n208 B.n207 10.6151
R2341 B.n207 B.n190 10.6151
R2342 B.n203 B.n190 10.6151
R2343 B.n203 B.n202 10.6151
R2344 B.n202 B.n201 10.6151
R2345 B.n201 B.n192 10.6151
R2346 B.n197 B.n192 10.6151
R2347 B.n197 B.n196 10.6151
R2348 B.n196 B.n195 10.6151
R2349 B.n195 B.n0 10.6151
R2350 B.n743 B.n1 10.6151
R2351 B.n743 B.n742 10.6151
R2352 B.n742 B.n741 10.6151
R2353 B.n741 B.n4 10.6151
R2354 B.n737 B.n4 10.6151
R2355 B.n737 B.n736 10.6151
R2356 B.n736 B.n735 10.6151
R2357 B.n735 B.n6 10.6151
R2358 B.n731 B.n6 10.6151
R2359 B.n731 B.n730 10.6151
R2360 B.n730 B.n729 10.6151
R2361 B.n729 B.n8 10.6151
R2362 B.n725 B.n8 10.6151
R2363 B.n725 B.n724 10.6151
R2364 B.n724 B.n723 10.6151
R2365 B.n723 B.n10 10.6151
R2366 B.n719 B.n10 10.6151
R2367 B.n719 B.n718 10.6151
R2368 B.n718 B.n717 10.6151
R2369 B.n717 B.n12 10.6151
R2370 B.n713 B.n12 10.6151
R2371 B.n713 B.n712 10.6151
R2372 B.n712 B.n711 10.6151
R2373 B.n711 B.n14 10.6151
R2374 B.n707 B.n14 10.6151
R2375 B.n707 B.n706 10.6151
R2376 B.n706 B.n705 10.6151
R2377 B.n705 B.n16 10.6151
R2378 B.n615 B.n614 6.5566
R2379 B.n602 B.n54 6.5566
R2380 B.n324 B.n323 6.5566
R2381 B.n336 B.n144 6.5566
R2382 B.n616 B.n615 4.05904
R2383 B.n599 B.n54 4.05904
R2384 B.n323 B.n322 4.05904
R2385 B.n339 B.n144 4.05904
R2386 B.n747 B.n0 2.81026
R2387 B.n747 B.n1 2.81026
R2388 VP.n7 VP.t7 446.76
R2389 VP.n17 VP.t1 424.293
R2390 VP.n29 VP.t5 424.293
R2391 VP.n15 VP.t4 424.293
R2392 VP.n22 VP.t3 388.033
R2393 VP.n1 VP.t6 388.033
R2394 VP.n5 VP.t2 388.033
R2395 VP.n8 VP.t0 388.033
R2396 VP.n9 VP.n6 161.3
R2397 VP.n11 VP.n10 161.3
R2398 VP.n13 VP.n12 161.3
R2399 VP.n14 VP.n4 161.3
R2400 VP.n28 VP.n0 161.3
R2401 VP.n27 VP.n26 161.3
R2402 VP.n25 VP.n24 161.3
R2403 VP.n23 VP.n2 161.3
R2404 VP.n21 VP.n20 161.3
R2405 VP.n19 VP.n3 161.3
R2406 VP.n16 VP.n15 80.6037
R2407 VP.n30 VP.n29 80.6037
R2408 VP.n18 VP.n17 80.6037
R2409 VP.n24 VP.n23 56.5193
R2410 VP.n10 VP.n9 56.5193
R2411 VP.n17 VP.n3 48.4452
R2412 VP.n29 VP.n28 48.4452
R2413 VP.n15 VP.n14 48.4452
R2414 VP.n18 VP.n16 48.1832
R2415 VP.n8 VP.n7 34.0975
R2416 VP.n7 VP.n6 28.4044
R2417 VP.n21 VP.n3 24.4675
R2418 VP.n28 VP.n27 24.4675
R2419 VP.n14 VP.n13 24.4675
R2420 VP.n23 VP.n22 22.5101
R2421 VP.n24 VP.n1 22.5101
R2422 VP.n10 VP.n5 22.5101
R2423 VP.n9 VP.n8 22.5101
R2424 VP.n22 VP.n21 1.95786
R2425 VP.n27 VP.n1 1.95786
R2426 VP.n13 VP.n5 1.95786
R2427 VP.n16 VP.n4 0.285035
R2428 VP.n19 VP.n18 0.285035
R2429 VP.n30 VP.n0 0.285035
R2430 VP.n11 VP.n6 0.189894
R2431 VP.n12 VP.n11 0.189894
R2432 VP.n12 VP.n4 0.189894
R2433 VP.n20 VP.n19 0.189894
R2434 VP.n20 VP.n2 0.189894
R2435 VP.n25 VP.n2 0.189894
R2436 VP.n26 VP.n25 0.189894
R2437 VP.n26 VP.n0 0.189894
R2438 VP VP.n30 0.146778
R2439 VDD1 VDD1.n0 70.2743
R2440 VDD1.n3 VDD1.n2 70.1606
R2441 VDD1.n3 VDD1.n1 70.1606
R2442 VDD1.n5 VDD1.n4 69.6039
R2443 VDD1.n5 VDD1.n3 44.9362
R2444 VDD1.n4 VDD1.t5 1.85264
R2445 VDD1.n4 VDD1.t3 1.85264
R2446 VDD1.n0 VDD1.t0 1.85264
R2447 VDD1.n0 VDD1.t7 1.85264
R2448 VDD1.n2 VDD1.t1 1.85264
R2449 VDD1.n2 VDD1.t2 1.85264
R2450 VDD1.n1 VDD1.t6 1.85264
R2451 VDD1.n1 VDD1.t4 1.85264
R2452 VDD1 VDD1.n5 0.554379
C0 VDD2 B 1.38746f
C1 w_n2390_n4478# VN 4.54303f
C2 VP w_n2390_n4478# 4.84885f
C3 w_n2390_n4478# VTAIL 5.50256f
C4 VDD1 w_n2390_n4478# 1.59695f
C5 B w_n2390_n4478# 9.360139f
C6 VP VN 6.84406f
C7 VDD2 w_n2390_n4478# 1.64812f
C8 VN VTAIL 9.37532f
C9 VP VTAIL 9.38943f
C10 VDD1 VN 0.149053f
C11 B VN 0.938219f
C12 VDD1 VP 9.889481f
C13 B VP 1.44283f
C14 VDD2 VN 9.68012f
C15 VDD2 VP 0.359046f
C16 VDD1 VTAIL 12.415701f
C17 B VTAIL 5.72409f
C18 VDD1 B 1.33873f
C19 VDD2 VTAIL 12.46f
C20 VDD1 VDD2 1.02147f
C21 VDD2 VSUBS 1.555074f
C22 VDD1 VSUBS 1.928169f
C23 VTAIL VSUBS 1.289083f
C24 VN VSUBS 5.37256f
C25 VP VSUBS 2.264868f
C26 B VSUBS 3.789273f
C27 w_n2390_n4478# VSUBS 0.130924p
C28 VDD1.t0 VSUBS 0.358715f
C29 VDD1.t7 VSUBS 0.358715f
C30 VDD1.n0 VSUBS 2.97915f
C31 VDD1.t6 VSUBS 0.358715f
C32 VDD1.t4 VSUBS 0.358715f
C33 VDD1.n1 VSUBS 2.97799f
C34 VDD1.t1 VSUBS 0.358715f
C35 VDD1.t2 VSUBS 0.358715f
C36 VDD1.n2 VSUBS 2.97799f
C37 VDD1.n3 VSUBS 3.47836f
C38 VDD1.t5 VSUBS 0.358715f
C39 VDD1.t3 VSUBS 0.358715f
C40 VDD1.n4 VSUBS 2.9727f
C41 VDD1.n5 VSUBS 3.27387f
C42 VP.n0 VSUBS 0.057263f
C43 VP.t6 VSUBS 2.25691f
C44 VP.n1 VSUBS 0.806355f
C45 VP.n2 VSUBS 0.042914f
C46 VP.t3 VSUBS 2.25691f
C47 VP.n3 VSUBS 0.049965f
C48 VP.n4 VSUBS 0.057263f
C49 VP.t4 VSUBS 2.32857f
C50 VP.t2 VSUBS 2.25691f
C51 VP.n5 VSUBS 0.806355f
C52 VP.n6 VSUBS 0.221767f
C53 VP.t0 VSUBS 2.25691f
C54 VP.t7 VSUBS 2.37323f
C55 VP.n7 VSUBS 0.86337f
C56 VP.n8 VSUBS 0.87216f
C57 VP.n9 VSUBS 0.059487f
C58 VP.n10 VSUBS 0.059487f
C59 VP.n11 VSUBS 0.042914f
C60 VP.n12 VSUBS 0.042914f
C61 VP.n13 VSUBS 0.043653f
C62 VP.n14 VSUBS 0.049965f
C63 VP.n15 VSUBS 0.87816f
C64 VP.n16 VSUBS 2.22088f
C65 VP.t1 VSUBS 2.32857f
C66 VP.n17 VSUBS 0.87816f
C67 VP.n18 VSUBS 2.25289f
C68 VP.n19 VSUBS 0.057263f
C69 VP.n20 VSUBS 0.042914f
C70 VP.n21 VSUBS 0.043653f
C71 VP.n22 VSUBS 0.806355f
C72 VP.n23 VSUBS 0.059487f
C73 VP.n24 VSUBS 0.059487f
C74 VP.n25 VSUBS 0.042914f
C75 VP.n26 VSUBS 0.042914f
C76 VP.n27 VSUBS 0.043653f
C77 VP.n28 VSUBS 0.049965f
C78 VP.t5 VSUBS 2.32857f
C79 VP.n29 VSUBS 0.87816f
C80 VP.n30 VSUBS 0.04019f
C81 B.n0 VSUBS 0.004608f
C82 B.n1 VSUBS 0.004608f
C83 B.n2 VSUBS 0.007286f
C84 B.n3 VSUBS 0.007286f
C85 B.n4 VSUBS 0.007286f
C86 B.n5 VSUBS 0.007286f
C87 B.n6 VSUBS 0.007286f
C88 B.n7 VSUBS 0.007286f
C89 B.n8 VSUBS 0.007286f
C90 B.n9 VSUBS 0.007286f
C91 B.n10 VSUBS 0.007286f
C92 B.n11 VSUBS 0.007286f
C93 B.n12 VSUBS 0.007286f
C94 B.n13 VSUBS 0.007286f
C95 B.n14 VSUBS 0.007286f
C96 B.n15 VSUBS 0.007286f
C97 B.n16 VSUBS 0.017561f
C98 B.n17 VSUBS 0.007286f
C99 B.n18 VSUBS 0.007286f
C100 B.n19 VSUBS 0.007286f
C101 B.n20 VSUBS 0.007286f
C102 B.n21 VSUBS 0.007286f
C103 B.n22 VSUBS 0.007286f
C104 B.n23 VSUBS 0.007286f
C105 B.n24 VSUBS 0.007286f
C106 B.n25 VSUBS 0.007286f
C107 B.n26 VSUBS 0.007286f
C108 B.n27 VSUBS 0.007286f
C109 B.n28 VSUBS 0.007286f
C110 B.n29 VSUBS 0.007286f
C111 B.n30 VSUBS 0.007286f
C112 B.n31 VSUBS 0.007286f
C113 B.n32 VSUBS 0.007286f
C114 B.n33 VSUBS 0.007286f
C115 B.n34 VSUBS 0.007286f
C116 B.n35 VSUBS 0.007286f
C117 B.n36 VSUBS 0.007286f
C118 B.n37 VSUBS 0.007286f
C119 B.n38 VSUBS 0.007286f
C120 B.n39 VSUBS 0.007286f
C121 B.n40 VSUBS 0.007286f
C122 B.n41 VSUBS 0.007286f
C123 B.n42 VSUBS 0.007286f
C124 B.n43 VSUBS 0.007286f
C125 B.n44 VSUBS 0.007286f
C126 B.n45 VSUBS 0.007286f
C127 B.t8 VSUBS 0.354194f
C128 B.t7 VSUBS 0.371684f
C129 B.t6 VSUBS 0.827982f
C130 B.n46 VSUBS 0.491948f
C131 B.n47 VSUBS 0.329969f
C132 B.n48 VSUBS 0.007286f
C133 B.n49 VSUBS 0.007286f
C134 B.n50 VSUBS 0.007286f
C135 B.n51 VSUBS 0.007286f
C136 B.t5 VSUBS 0.354197f
C137 B.t4 VSUBS 0.371688f
C138 B.t3 VSUBS 0.827982f
C139 B.n52 VSUBS 0.491945f
C140 B.n53 VSUBS 0.329965f
C141 B.n54 VSUBS 0.016882f
C142 B.n55 VSUBS 0.007286f
C143 B.n56 VSUBS 0.007286f
C144 B.n57 VSUBS 0.007286f
C145 B.n58 VSUBS 0.007286f
C146 B.n59 VSUBS 0.007286f
C147 B.n60 VSUBS 0.007286f
C148 B.n61 VSUBS 0.007286f
C149 B.n62 VSUBS 0.007286f
C150 B.n63 VSUBS 0.007286f
C151 B.n64 VSUBS 0.007286f
C152 B.n65 VSUBS 0.007286f
C153 B.n66 VSUBS 0.007286f
C154 B.n67 VSUBS 0.007286f
C155 B.n68 VSUBS 0.007286f
C156 B.n69 VSUBS 0.007286f
C157 B.n70 VSUBS 0.007286f
C158 B.n71 VSUBS 0.007286f
C159 B.n72 VSUBS 0.007286f
C160 B.n73 VSUBS 0.007286f
C161 B.n74 VSUBS 0.007286f
C162 B.n75 VSUBS 0.007286f
C163 B.n76 VSUBS 0.007286f
C164 B.n77 VSUBS 0.007286f
C165 B.n78 VSUBS 0.007286f
C166 B.n79 VSUBS 0.007286f
C167 B.n80 VSUBS 0.007286f
C168 B.n81 VSUBS 0.007286f
C169 B.n82 VSUBS 0.007286f
C170 B.n83 VSUBS 0.018014f
C171 B.n84 VSUBS 0.007286f
C172 B.n85 VSUBS 0.007286f
C173 B.n86 VSUBS 0.007286f
C174 B.n87 VSUBS 0.007286f
C175 B.n88 VSUBS 0.007286f
C176 B.n89 VSUBS 0.007286f
C177 B.n90 VSUBS 0.007286f
C178 B.n91 VSUBS 0.007286f
C179 B.n92 VSUBS 0.007286f
C180 B.n93 VSUBS 0.007286f
C181 B.n94 VSUBS 0.007286f
C182 B.n95 VSUBS 0.007286f
C183 B.n96 VSUBS 0.007286f
C184 B.n97 VSUBS 0.007286f
C185 B.n98 VSUBS 0.007286f
C186 B.n99 VSUBS 0.007286f
C187 B.n100 VSUBS 0.007286f
C188 B.n101 VSUBS 0.007286f
C189 B.n102 VSUBS 0.007286f
C190 B.n103 VSUBS 0.007286f
C191 B.n104 VSUBS 0.007286f
C192 B.n105 VSUBS 0.007286f
C193 B.n106 VSUBS 0.007286f
C194 B.n107 VSUBS 0.007286f
C195 B.n108 VSUBS 0.007286f
C196 B.n109 VSUBS 0.007286f
C197 B.n110 VSUBS 0.007286f
C198 B.n111 VSUBS 0.007286f
C199 B.n112 VSUBS 0.007286f
C200 B.n113 VSUBS 0.018014f
C201 B.n114 VSUBS 0.007286f
C202 B.n115 VSUBS 0.007286f
C203 B.n116 VSUBS 0.007286f
C204 B.n117 VSUBS 0.007286f
C205 B.n118 VSUBS 0.007286f
C206 B.n119 VSUBS 0.007286f
C207 B.n120 VSUBS 0.007286f
C208 B.n121 VSUBS 0.007286f
C209 B.n122 VSUBS 0.007286f
C210 B.n123 VSUBS 0.007286f
C211 B.n124 VSUBS 0.007286f
C212 B.n125 VSUBS 0.007286f
C213 B.n126 VSUBS 0.007286f
C214 B.n127 VSUBS 0.007286f
C215 B.n128 VSUBS 0.007286f
C216 B.n129 VSUBS 0.007286f
C217 B.n130 VSUBS 0.007286f
C218 B.n131 VSUBS 0.007286f
C219 B.n132 VSUBS 0.007286f
C220 B.n133 VSUBS 0.007286f
C221 B.n134 VSUBS 0.007286f
C222 B.n135 VSUBS 0.007286f
C223 B.n136 VSUBS 0.007286f
C224 B.n137 VSUBS 0.007286f
C225 B.n138 VSUBS 0.007286f
C226 B.n139 VSUBS 0.007286f
C227 B.n140 VSUBS 0.007286f
C228 B.n141 VSUBS 0.007286f
C229 B.t1 VSUBS 0.354197f
C230 B.t2 VSUBS 0.371688f
C231 B.t0 VSUBS 0.827982f
C232 B.n142 VSUBS 0.491945f
C233 B.n143 VSUBS 0.329965f
C234 B.n144 VSUBS 0.016882f
C235 B.n145 VSUBS 0.007286f
C236 B.n146 VSUBS 0.007286f
C237 B.n147 VSUBS 0.007286f
C238 B.n148 VSUBS 0.007286f
C239 B.n149 VSUBS 0.007286f
C240 B.t10 VSUBS 0.354194f
C241 B.t11 VSUBS 0.371684f
C242 B.t9 VSUBS 0.827982f
C243 B.n150 VSUBS 0.491948f
C244 B.n151 VSUBS 0.329969f
C245 B.n152 VSUBS 0.007286f
C246 B.n153 VSUBS 0.007286f
C247 B.n154 VSUBS 0.007286f
C248 B.n155 VSUBS 0.007286f
C249 B.n156 VSUBS 0.007286f
C250 B.n157 VSUBS 0.007286f
C251 B.n158 VSUBS 0.007286f
C252 B.n159 VSUBS 0.007286f
C253 B.n160 VSUBS 0.007286f
C254 B.n161 VSUBS 0.007286f
C255 B.n162 VSUBS 0.007286f
C256 B.n163 VSUBS 0.007286f
C257 B.n164 VSUBS 0.007286f
C258 B.n165 VSUBS 0.007286f
C259 B.n166 VSUBS 0.007286f
C260 B.n167 VSUBS 0.007286f
C261 B.n168 VSUBS 0.007286f
C262 B.n169 VSUBS 0.007286f
C263 B.n170 VSUBS 0.007286f
C264 B.n171 VSUBS 0.007286f
C265 B.n172 VSUBS 0.007286f
C266 B.n173 VSUBS 0.007286f
C267 B.n174 VSUBS 0.007286f
C268 B.n175 VSUBS 0.007286f
C269 B.n176 VSUBS 0.007286f
C270 B.n177 VSUBS 0.007286f
C271 B.n178 VSUBS 0.007286f
C272 B.n179 VSUBS 0.007286f
C273 B.n180 VSUBS 0.017561f
C274 B.n181 VSUBS 0.007286f
C275 B.n182 VSUBS 0.007286f
C276 B.n183 VSUBS 0.007286f
C277 B.n184 VSUBS 0.007286f
C278 B.n185 VSUBS 0.007286f
C279 B.n186 VSUBS 0.007286f
C280 B.n187 VSUBS 0.007286f
C281 B.n188 VSUBS 0.007286f
C282 B.n189 VSUBS 0.007286f
C283 B.n190 VSUBS 0.007286f
C284 B.n191 VSUBS 0.007286f
C285 B.n192 VSUBS 0.007286f
C286 B.n193 VSUBS 0.007286f
C287 B.n194 VSUBS 0.007286f
C288 B.n195 VSUBS 0.007286f
C289 B.n196 VSUBS 0.007286f
C290 B.n197 VSUBS 0.007286f
C291 B.n198 VSUBS 0.007286f
C292 B.n199 VSUBS 0.007286f
C293 B.n200 VSUBS 0.007286f
C294 B.n201 VSUBS 0.007286f
C295 B.n202 VSUBS 0.007286f
C296 B.n203 VSUBS 0.007286f
C297 B.n204 VSUBS 0.007286f
C298 B.n205 VSUBS 0.007286f
C299 B.n206 VSUBS 0.007286f
C300 B.n207 VSUBS 0.007286f
C301 B.n208 VSUBS 0.007286f
C302 B.n209 VSUBS 0.007286f
C303 B.n210 VSUBS 0.007286f
C304 B.n211 VSUBS 0.007286f
C305 B.n212 VSUBS 0.007286f
C306 B.n213 VSUBS 0.007286f
C307 B.n214 VSUBS 0.007286f
C308 B.n215 VSUBS 0.007286f
C309 B.n216 VSUBS 0.007286f
C310 B.n217 VSUBS 0.007286f
C311 B.n218 VSUBS 0.007286f
C312 B.n219 VSUBS 0.007286f
C313 B.n220 VSUBS 0.007286f
C314 B.n221 VSUBS 0.007286f
C315 B.n222 VSUBS 0.007286f
C316 B.n223 VSUBS 0.007286f
C317 B.n224 VSUBS 0.007286f
C318 B.n225 VSUBS 0.007286f
C319 B.n226 VSUBS 0.007286f
C320 B.n227 VSUBS 0.007286f
C321 B.n228 VSUBS 0.007286f
C322 B.n229 VSUBS 0.007286f
C323 B.n230 VSUBS 0.007286f
C324 B.n231 VSUBS 0.007286f
C325 B.n232 VSUBS 0.007286f
C326 B.n233 VSUBS 0.007286f
C327 B.n234 VSUBS 0.007286f
C328 B.n235 VSUBS 0.017561f
C329 B.n236 VSUBS 0.018014f
C330 B.n237 VSUBS 0.018014f
C331 B.n238 VSUBS 0.007286f
C332 B.n239 VSUBS 0.007286f
C333 B.n240 VSUBS 0.007286f
C334 B.n241 VSUBS 0.007286f
C335 B.n242 VSUBS 0.007286f
C336 B.n243 VSUBS 0.007286f
C337 B.n244 VSUBS 0.007286f
C338 B.n245 VSUBS 0.007286f
C339 B.n246 VSUBS 0.007286f
C340 B.n247 VSUBS 0.007286f
C341 B.n248 VSUBS 0.007286f
C342 B.n249 VSUBS 0.007286f
C343 B.n250 VSUBS 0.007286f
C344 B.n251 VSUBS 0.007286f
C345 B.n252 VSUBS 0.007286f
C346 B.n253 VSUBS 0.007286f
C347 B.n254 VSUBS 0.007286f
C348 B.n255 VSUBS 0.007286f
C349 B.n256 VSUBS 0.007286f
C350 B.n257 VSUBS 0.007286f
C351 B.n258 VSUBS 0.007286f
C352 B.n259 VSUBS 0.007286f
C353 B.n260 VSUBS 0.007286f
C354 B.n261 VSUBS 0.007286f
C355 B.n262 VSUBS 0.007286f
C356 B.n263 VSUBS 0.007286f
C357 B.n264 VSUBS 0.007286f
C358 B.n265 VSUBS 0.007286f
C359 B.n266 VSUBS 0.007286f
C360 B.n267 VSUBS 0.007286f
C361 B.n268 VSUBS 0.007286f
C362 B.n269 VSUBS 0.007286f
C363 B.n270 VSUBS 0.007286f
C364 B.n271 VSUBS 0.007286f
C365 B.n272 VSUBS 0.007286f
C366 B.n273 VSUBS 0.007286f
C367 B.n274 VSUBS 0.007286f
C368 B.n275 VSUBS 0.007286f
C369 B.n276 VSUBS 0.007286f
C370 B.n277 VSUBS 0.007286f
C371 B.n278 VSUBS 0.007286f
C372 B.n279 VSUBS 0.007286f
C373 B.n280 VSUBS 0.007286f
C374 B.n281 VSUBS 0.007286f
C375 B.n282 VSUBS 0.007286f
C376 B.n283 VSUBS 0.007286f
C377 B.n284 VSUBS 0.007286f
C378 B.n285 VSUBS 0.007286f
C379 B.n286 VSUBS 0.007286f
C380 B.n287 VSUBS 0.007286f
C381 B.n288 VSUBS 0.007286f
C382 B.n289 VSUBS 0.007286f
C383 B.n290 VSUBS 0.007286f
C384 B.n291 VSUBS 0.007286f
C385 B.n292 VSUBS 0.007286f
C386 B.n293 VSUBS 0.007286f
C387 B.n294 VSUBS 0.007286f
C388 B.n295 VSUBS 0.007286f
C389 B.n296 VSUBS 0.007286f
C390 B.n297 VSUBS 0.007286f
C391 B.n298 VSUBS 0.007286f
C392 B.n299 VSUBS 0.007286f
C393 B.n300 VSUBS 0.007286f
C394 B.n301 VSUBS 0.007286f
C395 B.n302 VSUBS 0.007286f
C396 B.n303 VSUBS 0.007286f
C397 B.n304 VSUBS 0.007286f
C398 B.n305 VSUBS 0.007286f
C399 B.n306 VSUBS 0.007286f
C400 B.n307 VSUBS 0.007286f
C401 B.n308 VSUBS 0.007286f
C402 B.n309 VSUBS 0.007286f
C403 B.n310 VSUBS 0.007286f
C404 B.n311 VSUBS 0.007286f
C405 B.n312 VSUBS 0.007286f
C406 B.n313 VSUBS 0.007286f
C407 B.n314 VSUBS 0.007286f
C408 B.n315 VSUBS 0.007286f
C409 B.n316 VSUBS 0.007286f
C410 B.n317 VSUBS 0.007286f
C411 B.n318 VSUBS 0.007286f
C412 B.n319 VSUBS 0.007286f
C413 B.n320 VSUBS 0.007286f
C414 B.n321 VSUBS 0.007286f
C415 B.n322 VSUBS 0.005036f
C416 B.n323 VSUBS 0.016882f
C417 B.n324 VSUBS 0.005893f
C418 B.n325 VSUBS 0.007286f
C419 B.n326 VSUBS 0.007286f
C420 B.n327 VSUBS 0.007286f
C421 B.n328 VSUBS 0.007286f
C422 B.n329 VSUBS 0.007286f
C423 B.n330 VSUBS 0.007286f
C424 B.n331 VSUBS 0.007286f
C425 B.n332 VSUBS 0.007286f
C426 B.n333 VSUBS 0.007286f
C427 B.n334 VSUBS 0.007286f
C428 B.n335 VSUBS 0.007286f
C429 B.n336 VSUBS 0.005893f
C430 B.n337 VSUBS 0.007286f
C431 B.n338 VSUBS 0.007286f
C432 B.n339 VSUBS 0.005036f
C433 B.n340 VSUBS 0.007286f
C434 B.n341 VSUBS 0.007286f
C435 B.n342 VSUBS 0.007286f
C436 B.n343 VSUBS 0.007286f
C437 B.n344 VSUBS 0.007286f
C438 B.n345 VSUBS 0.007286f
C439 B.n346 VSUBS 0.007286f
C440 B.n347 VSUBS 0.007286f
C441 B.n348 VSUBS 0.007286f
C442 B.n349 VSUBS 0.007286f
C443 B.n350 VSUBS 0.007286f
C444 B.n351 VSUBS 0.007286f
C445 B.n352 VSUBS 0.007286f
C446 B.n353 VSUBS 0.007286f
C447 B.n354 VSUBS 0.007286f
C448 B.n355 VSUBS 0.007286f
C449 B.n356 VSUBS 0.007286f
C450 B.n357 VSUBS 0.007286f
C451 B.n358 VSUBS 0.007286f
C452 B.n359 VSUBS 0.007286f
C453 B.n360 VSUBS 0.007286f
C454 B.n361 VSUBS 0.007286f
C455 B.n362 VSUBS 0.007286f
C456 B.n363 VSUBS 0.007286f
C457 B.n364 VSUBS 0.007286f
C458 B.n365 VSUBS 0.007286f
C459 B.n366 VSUBS 0.007286f
C460 B.n367 VSUBS 0.007286f
C461 B.n368 VSUBS 0.007286f
C462 B.n369 VSUBS 0.007286f
C463 B.n370 VSUBS 0.007286f
C464 B.n371 VSUBS 0.007286f
C465 B.n372 VSUBS 0.007286f
C466 B.n373 VSUBS 0.007286f
C467 B.n374 VSUBS 0.007286f
C468 B.n375 VSUBS 0.007286f
C469 B.n376 VSUBS 0.007286f
C470 B.n377 VSUBS 0.007286f
C471 B.n378 VSUBS 0.007286f
C472 B.n379 VSUBS 0.007286f
C473 B.n380 VSUBS 0.007286f
C474 B.n381 VSUBS 0.007286f
C475 B.n382 VSUBS 0.007286f
C476 B.n383 VSUBS 0.007286f
C477 B.n384 VSUBS 0.007286f
C478 B.n385 VSUBS 0.007286f
C479 B.n386 VSUBS 0.007286f
C480 B.n387 VSUBS 0.007286f
C481 B.n388 VSUBS 0.007286f
C482 B.n389 VSUBS 0.007286f
C483 B.n390 VSUBS 0.007286f
C484 B.n391 VSUBS 0.007286f
C485 B.n392 VSUBS 0.007286f
C486 B.n393 VSUBS 0.007286f
C487 B.n394 VSUBS 0.007286f
C488 B.n395 VSUBS 0.007286f
C489 B.n396 VSUBS 0.007286f
C490 B.n397 VSUBS 0.007286f
C491 B.n398 VSUBS 0.007286f
C492 B.n399 VSUBS 0.007286f
C493 B.n400 VSUBS 0.007286f
C494 B.n401 VSUBS 0.007286f
C495 B.n402 VSUBS 0.007286f
C496 B.n403 VSUBS 0.007286f
C497 B.n404 VSUBS 0.007286f
C498 B.n405 VSUBS 0.007286f
C499 B.n406 VSUBS 0.007286f
C500 B.n407 VSUBS 0.007286f
C501 B.n408 VSUBS 0.007286f
C502 B.n409 VSUBS 0.007286f
C503 B.n410 VSUBS 0.007286f
C504 B.n411 VSUBS 0.007286f
C505 B.n412 VSUBS 0.007286f
C506 B.n413 VSUBS 0.007286f
C507 B.n414 VSUBS 0.007286f
C508 B.n415 VSUBS 0.007286f
C509 B.n416 VSUBS 0.007286f
C510 B.n417 VSUBS 0.007286f
C511 B.n418 VSUBS 0.007286f
C512 B.n419 VSUBS 0.007286f
C513 B.n420 VSUBS 0.007286f
C514 B.n421 VSUBS 0.007286f
C515 B.n422 VSUBS 0.007286f
C516 B.n423 VSUBS 0.007286f
C517 B.n424 VSUBS 0.018014f
C518 B.n425 VSUBS 0.017561f
C519 B.n426 VSUBS 0.017561f
C520 B.n427 VSUBS 0.007286f
C521 B.n428 VSUBS 0.007286f
C522 B.n429 VSUBS 0.007286f
C523 B.n430 VSUBS 0.007286f
C524 B.n431 VSUBS 0.007286f
C525 B.n432 VSUBS 0.007286f
C526 B.n433 VSUBS 0.007286f
C527 B.n434 VSUBS 0.007286f
C528 B.n435 VSUBS 0.007286f
C529 B.n436 VSUBS 0.007286f
C530 B.n437 VSUBS 0.007286f
C531 B.n438 VSUBS 0.007286f
C532 B.n439 VSUBS 0.007286f
C533 B.n440 VSUBS 0.007286f
C534 B.n441 VSUBS 0.007286f
C535 B.n442 VSUBS 0.007286f
C536 B.n443 VSUBS 0.007286f
C537 B.n444 VSUBS 0.007286f
C538 B.n445 VSUBS 0.007286f
C539 B.n446 VSUBS 0.007286f
C540 B.n447 VSUBS 0.007286f
C541 B.n448 VSUBS 0.007286f
C542 B.n449 VSUBS 0.007286f
C543 B.n450 VSUBS 0.007286f
C544 B.n451 VSUBS 0.007286f
C545 B.n452 VSUBS 0.007286f
C546 B.n453 VSUBS 0.007286f
C547 B.n454 VSUBS 0.007286f
C548 B.n455 VSUBS 0.007286f
C549 B.n456 VSUBS 0.007286f
C550 B.n457 VSUBS 0.007286f
C551 B.n458 VSUBS 0.007286f
C552 B.n459 VSUBS 0.007286f
C553 B.n460 VSUBS 0.007286f
C554 B.n461 VSUBS 0.007286f
C555 B.n462 VSUBS 0.007286f
C556 B.n463 VSUBS 0.007286f
C557 B.n464 VSUBS 0.007286f
C558 B.n465 VSUBS 0.007286f
C559 B.n466 VSUBS 0.007286f
C560 B.n467 VSUBS 0.007286f
C561 B.n468 VSUBS 0.007286f
C562 B.n469 VSUBS 0.007286f
C563 B.n470 VSUBS 0.007286f
C564 B.n471 VSUBS 0.007286f
C565 B.n472 VSUBS 0.007286f
C566 B.n473 VSUBS 0.007286f
C567 B.n474 VSUBS 0.007286f
C568 B.n475 VSUBS 0.007286f
C569 B.n476 VSUBS 0.007286f
C570 B.n477 VSUBS 0.007286f
C571 B.n478 VSUBS 0.007286f
C572 B.n479 VSUBS 0.007286f
C573 B.n480 VSUBS 0.007286f
C574 B.n481 VSUBS 0.007286f
C575 B.n482 VSUBS 0.007286f
C576 B.n483 VSUBS 0.007286f
C577 B.n484 VSUBS 0.007286f
C578 B.n485 VSUBS 0.007286f
C579 B.n486 VSUBS 0.007286f
C580 B.n487 VSUBS 0.007286f
C581 B.n488 VSUBS 0.007286f
C582 B.n489 VSUBS 0.007286f
C583 B.n490 VSUBS 0.007286f
C584 B.n491 VSUBS 0.007286f
C585 B.n492 VSUBS 0.007286f
C586 B.n493 VSUBS 0.007286f
C587 B.n494 VSUBS 0.007286f
C588 B.n495 VSUBS 0.007286f
C589 B.n496 VSUBS 0.007286f
C590 B.n497 VSUBS 0.007286f
C591 B.n498 VSUBS 0.007286f
C592 B.n499 VSUBS 0.007286f
C593 B.n500 VSUBS 0.007286f
C594 B.n501 VSUBS 0.007286f
C595 B.n502 VSUBS 0.007286f
C596 B.n503 VSUBS 0.007286f
C597 B.n504 VSUBS 0.007286f
C598 B.n505 VSUBS 0.007286f
C599 B.n506 VSUBS 0.007286f
C600 B.n507 VSUBS 0.007286f
C601 B.n508 VSUBS 0.007286f
C602 B.n509 VSUBS 0.007286f
C603 B.n510 VSUBS 0.007286f
C604 B.n511 VSUBS 0.007286f
C605 B.n512 VSUBS 0.017561f
C606 B.n513 VSUBS 0.018369f
C607 B.n514 VSUBS 0.017206f
C608 B.n515 VSUBS 0.007286f
C609 B.n516 VSUBS 0.007286f
C610 B.n517 VSUBS 0.007286f
C611 B.n518 VSUBS 0.007286f
C612 B.n519 VSUBS 0.007286f
C613 B.n520 VSUBS 0.007286f
C614 B.n521 VSUBS 0.007286f
C615 B.n522 VSUBS 0.007286f
C616 B.n523 VSUBS 0.007286f
C617 B.n524 VSUBS 0.007286f
C618 B.n525 VSUBS 0.007286f
C619 B.n526 VSUBS 0.007286f
C620 B.n527 VSUBS 0.007286f
C621 B.n528 VSUBS 0.007286f
C622 B.n529 VSUBS 0.007286f
C623 B.n530 VSUBS 0.007286f
C624 B.n531 VSUBS 0.007286f
C625 B.n532 VSUBS 0.007286f
C626 B.n533 VSUBS 0.007286f
C627 B.n534 VSUBS 0.007286f
C628 B.n535 VSUBS 0.007286f
C629 B.n536 VSUBS 0.007286f
C630 B.n537 VSUBS 0.007286f
C631 B.n538 VSUBS 0.007286f
C632 B.n539 VSUBS 0.007286f
C633 B.n540 VSUBS 0.007286f
C634 B.n541 VSUBS 0.007286f
C635 B.n542 VSUBS 0.007286f
C636 B.n543 VSUBS 0.007286f
C637 B.n544 VSUBS 0.007286f
C638 B.n545 VSUBS 0.007286f
C639 B.n546 VSUBS 0.007286f
C640 B.n547 VSUBS 0.007286f
C641 B.n548 VSUBS 0.007286f
C642 B.n549 VSUBS 0.007286f
C643 B.n550 VSUBS 0.007286f
C644 B.n551 VSUBS 0.007286f
C645 B.n552 VSUBS 0.007286f
C646 B.n553 VSUBS 0.007286f
C647 B.n554 VSUBS 0.007286f
C648 B.n555 VSUBS 0.007286f
C649 B.n556 VSUBS 0.007286f
C650 B.n557 VSUBS 0.007286f
C651 B.n558 VSUBS 0.007286f
C652 B.n559 VSUBS 0.007286f
C653 B.n560 VSUBS 0.007286f
C654 B.n561 VSUBS 0.007286f
C655 B.n562 VSUBS 0.007286f
C656 B.n563 VSUBS 0.007286f
C657 B.n564 VSUBS 0.007286f
C658 B.n565 VSUBS 0.007286f
C659 B.n566 VSUBS 0.007286f
C660 B.n567 VSUBS 0.007286f
C661 B.n568 VSUBS 0.007286f
C662 B.n569 VSUBS 0.007286f
C663 B.n570 VSUBS 0.007286f
C664 B.n571 VSUBS 0.007286f
C665 B.n572 VSUBS 0.007286f
C666 B.n573 VSUBS 0.007286f
C667 B.n574 VSUBS 0.007286f
C668 B.n575 VSUBS 0.007286f
C669 B.n576 VSUBS 0.007286f
C670 B.n577 VSUBS 0.007286f
C671 B.n578 VSUBS 0.007286f
C672 B.n579 VSUBS 0.007286f
C673 B.n580 VSUBS 0.007286f
C674 B.n581 VSUBS 0.007286f
C675 B.n582 VSUBS 0.007286f
C676 B.n583 VSUBS 0.007286f
C677 B.n584 VSUBS 0.007286f
C678 B.n585 VSUBS 0.007286f
C679 B.n586 VSUBS 0.007286f
C680 B.n587 VSUBS 0.007286f
C681 B.n588 VSUBS 0.007286f
C682 B.n589 VSUBS 0.007286f
C683 B.n590 VSUBS 0.007286f
C684 B.n591 VSUBS 0.007286f
C685 B.n592 VSUBS 0.007286f
C686 B.n593 VSUBS 0.007286f
C687 B.n594 VSUBS 0.007286f
C688 B.n595 VSUBS 0.007286f
C689 B.n596 VSUBS 0.007286f
C690 B.n597 VSUBS 0.007286f
C691 B.n598 VSUBS 0.007286f
C692 B.n599 VSUBS 0.005036f
C693 B.n600 VSUBS 0.007286f
C694 B.n601 VSUBS 0.007286f
C695 B.n602 VSUBS 0.005893f
C696 B.n603 VSUBS 0.007286f
C697 B.n604 VSUBS 0.007286f
C698 B.n605 VSUBS 0.007286f
C699 B.n606 VSUBS 0.007286f
C700 B.n607 VSUBS 0.007286f
C701 B.n608 VSUBS 0.007286f
C702 B.n609 VSUBS 0.007286f
C703 B.n610 VSUBS 0.007286f
C704 B.n611 VSUBS 0.007286f
C705 B.n612 VSUBS 0.007286f
C706 B.n613 VSUBS 0.007286f
C707 B.n614 VSUBS 0.005893f
C708 B.n615 VSUBS 0.016882f
C709 B.n616 VSUBS 0.005036f
C710 B.n617 VSUBS 0.007286f
C711 B.n618 VSUBS 0.007286f
C712 B.n619 VSUBS 0.007286f
C713 B.n620 VSUBS 0.007286f
C714 B.n621 VSUBS 0.007286f
C715 B.n622 VSUBS 0.007286f
C716 B.n623 VSUBS 0.007286f
C717 B.n624 VSUBS 0.007286f
C718 B.n625 VSUBS 0.007286f
C719 B.n626 VSUBS 0.007286f
C720 B.n627 VSUBS 0.007286f
C721 B.n628 VSUBS 0.007286f
C722 B.n629 VSUBS 0.007286f
C723 B.n630 VSUBS 0.007286f
C724 B.n631 VSUBS 0.007286f
C725 B.n632 VSUBS 0.007286f
C726 B.n633 VSUBS 0.007286f
C727 B.n634 VSUBS 0.007286f
C728 B.n635 VSUBS 0.007286f
C729 B.n636 VSUBS 0.007286f
C730 B.n637 VSUBS 0.007286f
C731 B.n638 VSUBS 0.007286f
C732 B.n639 VSUBS 0.007286f
C733 B.n640 VSUBS 0.007286f
C734 B.n641 VSUBS 0.007286f
C735 B.n642 VSUBS 0.007286f
C736 B.n643 VSUBS 0.007286f
C737 B.n644 VSUBS 0.007286f
C738 B.n645 VSUBS 0.007286f
C739 B.n646 VSUBS 0.007286f
C740 B.n647 VSUBS 0.007286f
C741 B.n648 VSUBS 0.007286f
C742 B.n649 VSUBS 0.007286f
C743 B.n650 VSUBS 0.007286f
C744 B.n651 VSUBS 0.007286f
C745 B.n652 VSUBS 0.007286f
C746 B.n653 VSUBS 0.007286f
C747 B.n654 VSUBS 0.007286f
C748 B.n655 VSUBS 0.007286f
C749 B.n656 VSUBS 0.007286f
C750 B.n657 VSUBS 0.007286f
C751 B.n658 VSUBS 0.007286f
C752 B.n659 VSUBS 0.007286f
C753 B.n660 VSUBS 0.007286f
C754 B.n661 VSUBS 0.007286f
C755 B.n662 VSUBS 0.007286f
C756 B.n663 VSUBS 0.007286f
C757 B.n664 VSUBS 0.007286f
C758 B.n665 VSUBS 0.007286f
C759 B.n666 VSUBS 0.007286f
C760 B.n667 VSUBS 0.007286f
C761 B.n668 VSUBS 0.007286f
C762 B.n669 VSUBS 0.007286f
C763 B.n670 VSUBS 0.007286f
C764 B.n671 VSUBS 0.007286f
C765 B.n672 VSUBS 0.007286f
C766 B.n673 VSUBS 0.007286f
C767 B.n674 VSUBS 0.007286f
C768 B.n675 VSUBS 0.007286f
C769 B.n676 VSUBS 0.007286f
C770 B.n677 VSUBS 0.007286f
C771 B.n678 VSUBS 0.007286f
C772 B.n679 VSUBS 0.007286f
C773 B.n680 VSUBS 0.007286f
C774 B.n681 VSUBS 0.007286f
C775 B.n682 VSUBS 0.007286f
C776 B.n683 VSUBS 0.007286f
C777 B.n684 VSUBS 0.007286f
C778 B.n685 VSUBS 0.007286f
C779 B.n686 VSUBS 0.007286f
C780 B.n687 VSUBS 0.007286f
C781 B.n688 VSUBS 0.007286f
C782 B.n689 VSUBS 0.007286f
C783 B.n690 VSUBS 0.007286f
C784 B.n691 VSUBS 0.007286f
C785 B.n692 VSUBS 0.007286f
C786 B.n693 VSUBS 0.007286f
C787 B.n694 VSUBS 0.007286f
C788 B.n695 VSUBS 0.007286f
C789 B.n696 VSUBS 0.007286f
C790 B.n697 VSUBS 0.007286f
C791 B.n698 VSUBS 0.007286f
C792 B.n699 VSUBS 0.007286f
C793 B.n700 VSUBS 0.007286f
C794 B.n701 VSUBS 0.018014f
C795 B.n702 VSUBS 0.018014f
C796 B.n703 VSUBS 0.017561f
C797 B.n704 VSUBS 0.007286f
C798 B.n705 VSUBS 0.007286f
C799 B.n706 VSUBS 0.007286f
C800 B.n707 VSUBS 0.007286f
C801 B.n708 VSUBS 0.007286f
C802 B.n709 VSUBS 0.007286f
C803 B.n710 VSUBS 0.007286f
C804 B.n711 VSUBS 0.007286f
C805 B.n712 VSUBS 0.007286f
C806 B.n713 VSUBS 0.007286f
C807 B.n714 VSUBS 0.007286f
C808 B.n715 VSUBS 0.007286f
C809 B.n716 VSUBS 0.007286f
C810 B.n717 VSUBS 0.007286f
C811 B.n718 VSUBS 0.007286f
C812 B.n719 VSUBS 0.007286f
C813 B.n720 VSUBS 0.007286f
C814 B.n721 VSUBS 0.007286f
C815 B.n722 VSUBS 0.007286f
C816 B.n723 VSUBS 0.007286f
C817 B.n724 VSUBS 0.007286f
C818 B.n725 VSUBS 0.007286f
C819 B.n726 VSUBS 0.007286f
C820 B.n727 VSUBS 0.007286f
C821 B.n728 VSUBS 0.007286f
C822 B.n729 VSUBS 0.007286f
C823 B.n730 VSUBS 0.007286f
C824 B.n731 VSUBS 0.007286f
C825 B.n732 VSUBS 0.007286f
C826 B.n733 VSUBS 0.007286f
C827 B.n734 VSUBS 0.007286f
C828 B.n735 VSUBS 0.007286f
C829 B.n736 VSUBS 0.007286f
C830 B.n737 VSUBS 0.007286f
C831 B.n738 VSUBS 0.007286f
C832 B.n739 VSUBS 0.007286f
C833 B.n740 VSUBS 0.007286f
C834 B.n741 VSUBS 0.007286f
C835 B.n742 VSUBS 0.007286f
C836 B.n743 VSUBS 0.007286f
C837 B.n744 VSUBS 0.007286f
C838 B.n745 VSUBS 0.007286f
C839 B.n746 VSUBS 0.007286f
C840 B.n747 VSUBS 0.016499f
C841 VDD2.t3 VSUBS 0.358643f
C842 VDD2.t7 VSUBS 0.358643f
C843 VDD2.n0 VSUBS 2.97739f
C844 VDD2.t5 VSUBS 0.358643f
C845 VDD2.t0 VSUBS 0.358643f
C846 VDD2.n1 VSUBS 2.97739f
C847 VDD2.n2 VSUBS 3.4231f
C848 VDD2.t4 VSUBS 0.358643f
C849 VDD2.t6 VSUBS 0.358643f
C850 VDD2.n3 VSUBS 2.97211f
C851 VDD2.n4 VSUBS 3.24194f
C852 VDD2.t1 VSUBS 0.358643f
C853 VDD2.t2 VSUBS 0.358643f
C854 VDD2.n5 VSUBS 2.97735f
C855 VTAIL.t8 VSUBS 0.324604f
C856 VTAIL.t11 VSUBS 0.324604f
C857 VTAIL.n0 VSUBS 2.54702f
C858 VTAIL.n1 VSUBS 0.666087f
C859 VTAIL.n2 VSUBS 0.025521f
C860 VTAIL.n3 VSUBS 0.023406f
C861 VTAIL.n4 VSUBS 0.012577f
C862 VTAIL.n5 VSUBS 0.029728f
C863 VTAIL.n6 VSUBS 0.013317f
C864 VTAIL.n7 VSUBS 0.023406f
C865 VTAIL.n8 VSUBS 0.012577f
C866 VTAIL.n9 VSUBS 0.029728f
C867 VTAIL.n10 VSUBS 0.012947f
C868 VTAIL.n11 VSUBS 0.023406f
C869 VTAIL.n12 VSUBS 0.013317f
C870 VTAIL.n13 VSUBS 0.029728f
C871 VTAIL.n14 VSUBS 0.013317f
C872 VTAIL.n15 VSUBS 0.023406f
C873 VTAIL.n16 VSUBS 0.012577f
C874 VTAIL.n17 VSUBS 0.029728f
C875 VTAIL.n18 VSUBS 0.013317f
C876 VTAIL.n19 VSUBS 0.023406f
C877 VTAIL.n20 VSUBS 0.012577f
C878 VTAIL.n21 VSUBS 0.029728f
C879 VTAIL.n22 VSUBS 0.013317f
C880 VTAIL.n23 VSUBS 0.023406f
C881 VTAIL.n24 VSUBS 0.012577f
C882 VTAIL.n25 VSUBS 0.029728f
C883 VTAIL.n26 VSUBS 0.013317f
C884 VTAIL.n27 VSUBS 0.023406f
C885 VTAIL.n28 VSUBS 0.012577f
C886 VTAIL.n29 VSUBS 0.029728f
C887 VTAIL.n30 VSUBS 0.013317f
C888 VTAIL.n31 VSUBS 1.76546f
C889 VTAIL.n32 VSUBS 0.012577f
C890 VTAIL.t14 VSUBS 0.06379f
C891 VTAIL.n33 VSUBS 0.182595f
C892 VTAIL.n34 VSUBS 0.018912f
C893 VTAIL.n35 VSUBS 0.022296f
C894 VTAIL.n36 VSUBS 0.029728f
C895 VTAIL.n37 VSUBS 0.013317f
C896 VTAIL.n38 VSUBS 0.012577f
C897 VTAIL.n39 VSUBS 0.023406f
C898 VTAIL.n40 VSUBS 0.023406f
C899 VTAIL.n41 VSUBS 0.012577f
C900 VTAIL.n42 VSUBS 0.013317f
C901 VTAIL.n43 VSUBS 0.029728f
C902 VTAIL.n44 VSUBS 0.029728f
C903 VTAIL.n45 VSUBS 0.013317f
C904 VTAIL.n46 VSUBS 0.012577f
C905 VTAIL.n47 VSUBS 0.023406f
C906 VTAIL.n48 VSUBS 0.023406f
C907 VTAIL.n49 VSUBS 0.012577f
C908 VTAIL.n50 VSUBS 0.013317f
C909 VTAIL.n51 VSUBS 0.029728f
C910 VTAIL.n52 VSUBS 0.029728f
C911 VTAIL.n53 VSUBS 0.013317f
C912 VTAIL.n54 VSUBS 0.012577f
C913 VTAIL.n55 VSUBS 0.023406f
C914 VTAIL.n56 VSUBS 0.023406f
C915 VTAIL.n57 VSUBS 0.012577f
C916 VTAIL.n58 VSUBS 0.013317f
C917 VTAIL.n59 VSUBS 0.029728f
C918 VTAIL.n60 VSUBS 0.029728f
C919 VTAIL.n61 VSUBS 0.013317f
C920 VTAIL.n62 VSUBS 0.012577f
C921 VTAIL.n63 VSUBS 0.023406f
C922 VTAIL.n64 VSUBS 0.023406f
C923 VTAIL.n65 VSUBS 0.012577f
C924 VTAIL.n66 VSUBS 0.013317f
C925 VTAIL.n67 VSUBS 0.029728f
C926 VTAIL.n68 VSUBS 0.029728f
C927 VTAIL.n69 VSUBS 0.013317f
C928 VTAIL.n70 VSUBS 0.012577f
C929 VTAIL.n71 VSUBS 0.023406f
C930 VTAIL.n72 VSUBS 0.023406f
C931 VTAIL.n73 VSUBS 0.012577f
C932 VTAIL.n74 VSUBS 0.012577f
C933 VTAIL.n75 VSUBS 0.013317f
C934 VTAIL.n76 VSUBS 0.029728f
C935 VTAIL.n77 VSUBS 0.029728f
C936 VTAIL.n78 VSUBS 0.029728f
C937 VTAIL.n79 VSUBS 0.012947f
C938 VTAIL.n80 VSUBS 0.012577f
C939 VTAIL.n81 VSUBS 0.023406f
C940 VTAIL.n82 VSUBS 0.023406f
C941 VTAIL.n83 VSUBS 0.012577f
C942 VTAIL.n84 VSUBS 0.013317f
C943 VTAIL.n85 VSUBS 0.029728f
C944 VTAIL.n86 VSUBS 0.029728f
C945 VTAIL.n87 VSUBS 0.013317f
C946 VTAIL.n88 VSUBS 0.012577f
C947 VTAIL.n89 VSUBS 0.023406f
C948 VTAIL.n90 VSUBS 0.023406f
C949 VTAIL.n91 VSUBS 0.012577f
C950 VTAIL.n92 VSUBS 0.013317f
C951 VTAIL.n93 VSUBS 0.029728f
C952 VTAIL.n94 VSUBS 0.071297f
C953 VTAIL.n95 VSUBS 0.013317f
C954 VTAIL.n96 VSUBS 0.012577f
C955 VTAIL.n97 VSUBS 0.055061f
C956 VTAIL.n98 VSUBS 0.035854f
C957 VTAIL.n99 VSUBS 0.148288f
C958 VTAIL.n100 VSUBS 0.025521f
C959 VTAIL.n101 VSUBS 0.023406f
C960 VTAIL.n102 VSUBS 0.012577f
C961 VTAIL.n103 VSUBS 0.029728f
C962 VTAIL.n104 VSUBS 0.013317f
C963 VTAIL.n105 VSUBS 0.023406f
C964 VTAIL.n106 VSUBS 0.012577f
C965 VTAIL.n107 VSUBS 0.029728f
C966 VTAIL.n108 VSUBS 0.012947f
C967 VTAIL.n109 VSUBS 0.023406f
C968 VTAIL.n110 VSUBS 0.013317f
C969 VTAIL.n111 VSUBS 0.029728f
C970 VTAIL.n112 VSUBS 0.013317f
C971 VTAIL.n113 VSUBS 0.023406f
C972 VTAIL.n114 VSUBS 0.012577f
C973 VTAIL.n115 VSUBS 0.029728f
C974 VTAIL.n116 VSUBS 0.013317f
C975 VTAIL.n117 VSUBS 0.023406f
C976 VTAIL.n118 VSUBS 0.012577f
C977 VTAIL.n119 VSUBS 0.029728f
C978 VTAIL.n120 VSUBS 0.013317f
C979 VTAIL.n121 VSUBS 0.023406f
C980 VTAIL.n122 VSUBS 0.012577f
C981 VTAIL.n123 VSUBS 0.029728f
C982 VTAIL.n124 VSUBS 0.013317f
C983 VTAIL.n125 VSUBS 0.023406f
C984 VTAIL.n126 VSUBS 0.012577f
C985 VTAIL.n127 VSUBS 0.029728f
C986 VTAIL.n128 VSUBS 0.013317f
C987 VTAIL.n129 VSUBS 1.76546f
C988 VTAIL.n130 VSUBS 0.012577f
C989 VTAIL.t4 VSUBS 0.06379f
C990 VTAIL.n131 VSUBS 0.182595f
C991 VTAIL.n132 VSUBS 0.018912f
C992 VTAIL.n133 VSUBS 0.022296f
C993 VTAIL.n134 VSUBS 0.029728f
C994 VTAIL.n135 VSUBS 0.013317f
C995 VTAIL.n136 VSUBS 0.012577f
C996 VTAIL.n137 VSUBS 0.023406f
C997 VTAIL.n138 VSUBS 0.023406f
C998 VTAIL.n139 VSUBS 0.012577f
C999 VTAIL.n140 VSUBS 0.013317f
C1000 VTAIL.n141 VSUBS 0.029728f
C1001 VTAIL.n142 VSUBS 0.029728f
C1002 VTAIL.n143 VSUBS 0.013317f
C1003 VTAIL.n144 VSUBS 0.012577f
C1004 VTAIL.n145 VSUBS 0.023406f
C1005 VTAIL.n146 VSUBS 0.023406f
C1006 VTAIL.n147 VSUBS 0.012577f
C1007 VTAIL.n148 VSUBS 0.013317f
C1008 VTAIL.n149 VSUBS 0.029728f
C1009 VTAIL.n150 VSUBS 0.029728f
C1010 VTAIL.n151 VSUBS 0.013317f
C1011 VTAIL.n152 VSUBS 0.012577f
C1012 VTAIL.n153 VSUBS 0.023406f
C1013 VTAIL.n154 VSUBS 0.023406f
C1014 VTAIL.n155 VSUBS 0.012577f
C1015 VTAIL.n156 VSUBS 0.013317f
C1016 VTAIL.n157 VSUBS 0.029728f
C1017 VTAIL.n158 VSUBS 0.029728f
C1018 VTAIL.n159 VSUBS 0.013317f
C1019 VTAIL.n160 VSUBS 0.012577f
C1020 VTAIL.n161 VSUBS 0.023406f
C1021 VTAIL.n162 VSUBS 0.023406f
C1022 VTAIL.n163 VSUBS 0.012577f
C1023 VTAIL.n164 VSUBS 0.013317f
C1024 VTAIL.n165 VSUBS 0.029728f
C1025 VTAIL.n166 VSUBS 0.029728f
C1026 VTAIL.n167 VSUBS 0.013317f
C1027 VTAIL.n168 VSUBS 0.012577f
C1028 VTAIL.n169 VSUBS 0.023406f
C1029 VTAIL.n170 VSUBS 0.023406f
C1030 VTAIL.n171 VSUBS 0.012577f
C1031 VTAIL.n172 VSUBS 0.012577f
C1032 VTAIL.n173 VSUBS 0.013317f
C1033 VTAIL.n174 VSUBS 0.029728f
C1034 VTAIL.n175 VSUBS 0.029728f
C1035 VTAIL.n176 VSUBS 0.029728f
C1036 VTAIL.n177 VSUBS 0.012947f
C1037 VTAIL.n178 VSUBS 0.012577f
C1038 VTAIL.n179 VSUBS 0.023406f
C1039 VTAIL.n180 VSUBS 0.023406f
C1040 VTAIL.n181 VSUBS 0.012577f
C1041 VTAIL.n182 VSUBS 0.013317f
C1042 VTAIL.n183 VSUBS 0.029728f
C1043 VTAIL.n184 VSUBS 0.029728f
C1044 VTAIL.n185 VSUBS 0.013317f
C1045 VTAIL.n186 VSUBS 0.012577f
C1046 VTAIL.n187 VSUBS 0.023406f
C1047 VTAIL.n188 VSUBS 0.023406f
C1048 VTAIL.n189 VSUBS 0.012577f
C1049 VTAIL.n190 VSUBS 0.013317f
C1050 VTAIL.n191 VSUBS 0.029728f
C1051 VTAIL.n192 VSUBS 0.071297f
C1052 VTAIL.n193 VSUBS 0.013317f
C1053 VTAIL.n194 VSUBS 0.012577f
C1054 VTAIL.n195 VSUBS 0.055061f
C1055 VTAIL.n196 VSUBS 0.035854f
C1056 VTAIL.n197 VSUBS 0.148288f
C1057 VTAIL.t6 VSUBS 0.324604f
C1058 VTAIL.t3 VSUBS 0.324604f
C1059 VTAIL.n198 VSUBS 2.54702f
C1060 VTAIL.n199 VSUBS 0.754022f
C1061 VTAIL.n200 VSUBS 0.025521f
C1062 VTAIL.n201 VSUBS 0.023406f
C1063 VTAIL.n202 VSUBS 0.012577f
C1064 VTAIL.n203 VSUBS 0.029728f
C1065 VTAIL.n204 VSUBS 0.013317f
C1066 VTAIL.n205 VSUBS 0.023406f
C1067 VTAIL.n206 VSUBS 0.012577f
C1068 VTAIL.n207 VSUBS 0.029728f
C1069 VTAIL.n208 VSUBS 0.012947f
C1070 VTAIL.n209 VSUBS 0.023406f
C1071 VTAIL.n210 VSUBS 0.013317f
C1072 VTAIL.n211 VSUBS 0.029728f
C1073 VTAIL.n212 VSUBS 0.013317f
C1074 VTAIL.n213 VSUBS 0.023406f
C1075 VTAIL.n214 VSUBS 0.012577f
C1076 VTAIL.n215 VSUBS 0.029728f
C1077 VTAIL.n216 VSUBS 0.013317f
C1078 VTAIL.n217 VSUBS 0.023406f
C1079 VTAIL.n218 VSUBS 0.012577f
C1080 VTAIL.n219 VSUBS 0.029728f
C1081 VTAIL.n220 VSUBS 0.013317f
C1082 VTAIL.n221 VSUBS 0.023406f
C1083 VTAIL.n222 VSUBS 0.012577f
C1084 VTAIL.n223 VSUBS 0.029728f
C1085 VTAIL.n224 VSUBS 0.013317f
C1086 VTAIL.n225 VSUBS 0.023406f
C1087 VTAIL.n226 VSUBS 0.012577f
C1088 VTAIL.n227 VSUBS 0.029728f
C1089 VTAIL.n228 VSUBS 0.013317f
C1090 VTAIL.n229 VSUBS 1.76546f
C1091 VTAIL.n230 VSUBS 0.012577f
C1092 VTAIL.t7 VSUBS 0.06379f
C1093 VTAIL.n231 VSUBS 0.182595f
C1094 VTAIL.n232 VSUBS 0.018912f
C1095 VTAIL.n233 VSUBS 0.022296f
C1096 VTAIL.n234 VSUBS 0.029728f
C1097 VTAIL.n235 VSUBS 0.013317f
C1098 VTAIL.n236 VSUBS 0.012577f
C1099 VTAIL.n237 VSUBS 0.023406f
C1100 VTAIL.n238 VSUBS 0.023406f
C1101 VTAIL.n239 VSUBS 0.012577f
C1102 VTAIL.n240 VSUBS 0.013317f
C1103 VTAIL.n241 VSUBS 0.029728f
C1104 VTAIL.n242 VSUBS 0.029728f
C1105 VTAIL.n243 VSUBS 0.013317f
C1106 VTAIL.n244 VSUBS 0.012577f
C1107 VTAIL.n245 VSUBS 0.023406f
C1108 VTAIL.n246 VSUBS 0.023406f
C1109 VTAIL.n247 VSUBS 0.012577f
C1110 VTAIL.n248 VSUBS 0.013317f
C1111 VTAIL.n249 VSUBS 0.029728f
C1112 VTAIL.n250 VSUBS 0.029728f
C1113 VTAIL.n251 VSUBS 0.013317f
C1114 VTAIL.n252 VSUBS 0.012577f
C1115 VTAIL.n253 VSUBS 0.023406f
C1116 VTAIL.n254 VSUBS 0.023406f
C1117 VTAIL.n255 VSUBS 0.012577f
C1118 VTAIL.n256 VSUBS 0.013317f
C1119 VTAIL.n257 VSUBS 0.029728f
C1120 VTAIL.n258 VSUBS 0.029728f
C1121 VTAIL.n259 VSUBS 0.013317f
C1122 VTAIL.n260 VSUBS 0.012577f
C1123 VTAIL.n261 VSUBS 0.023406f
C1124 VTAIL.n262 VSUBS 0.023406f
C1125 VTAIL.n263 VSUBS 0.012577f
C1126 VTAIL.n264 VSUBS 0.013317f
C1127 VTAIL.n265 VSUBS 0.029728f
C1128 VTAIL.n266 VSUBS 0.029728f
C1129 VTAIL.n267 VSUBS 0.013317f
C1130 VTAIL.n268 VSUBS 0.012577f
C1131 VTAIL.n269 VSUBS 0.023406f
C1132 VTAIL.n270 VSUBS 0.023406f
C1133 VTAIL.n271 VSUBS 0.012577f
C1134 VTAIL.n272 VSUBS 0.012577f
C1135 VTAIL.n273 VSUBS 0.013317f
C1136 VTAIL.n274 VSUBS 0.029728f
C1137 VTAIL.n275 VSUBS 0.029728f
C1138 VTAIL.n276 VSUBS 0.029728f
C1139 VTAIL.n277 VSUBS 0.012947f
C1140 VTAIL.n278 VSUBS 0.012577f
C1141 VTAIL.n279 VSUBS 0.023406f
C1142 VTAIL.n280 VSUBS 0.023406f
C1143 VTAIL.n281 VSUBS 0.012577f
C1144 VTAIL.n282 VSUBS 0.013317f
C1145 VTAIL.n283 VSUBS 0.029728f
C1146 VTAIL.n284 VSUBS 0.029728f
C1147 VTAIL.n285 VSUBS 0.013317f
C1148 VTAIL.n286 VSUBS 0.012577f
C1149 VTAIL.n287 VSUBS 0.023406f
C1150 VTAIL.n288 VSUBS 0.023406f
C1151 VTAIL.n289 VSUBS 0.012577f
C1152 VTAIL.n290 VSUBS 0.013317f
C1153 VTAIL.n291 VSUBS 0.029728f
C1154 VTAIL.n292 VSUBS 0.071297f
C1155 VTAIL.n293 VSUBS 0.013317f
C1156 VTAIL.n294 VSUBS 0.012577f
C1157 VTAIL.n295 VSUBS 0.055061f
C1158 VTAIL.n296 VSUBS 0.035854f
C1159 VTAIL.n297 VSUBS 1.66415f
C1160 VTAIL.n298 VSUBS 0.025521f
C1161 VTAIL.n299 VSUBS 0.023406f
C1162 VTAIL.n300 VSUBS 0.012577f
C1163 VTAIL.n301 VSUBS 0.029728f
C1164 VTAIL.n302 VSUBS 0.013317f
C1165 VTAIL.n303 VSUBS 0.023406f
C1166 VTAIL.n304 VSUBS 0.012577f
C1167 VTAIL.n305 VSUBS 0.029728f
C1168 VTAIL.n306 VSUBS 0.012947f
C1169 VTAIL.n307 VSUBS 0.023406f
C1170 VTAIL.n308 VSUBS 0.012947f
C1171 VTAIL.n309 VSUBS 0.012577f
C1172 VTAIL.n310 VSUBS 0.029728f
C1173 VTAIL.n311 VSUBS 0.029728f
C1174 VTAIL.n312 VSUBS 0.013317f
C1175 VTAIL.n313 VSUBS 0.023406f
C1176 VTAIL.n314 VSUBS 0.012577f
C1177 VTAIL.n315 VSUBS 0.029728f
C1178 VTAIL.n316 VSUBS 0.013317f
C1179 VTAIL.n317 VSUBS 0.023406f
C1180 VTAIL.n318 VSUBS 0.012577f
C1181 VTAIL.n319 VSUBS 0.029728f
C1182 VTAIL.n320 VSUBS 0.013317f
C1183 VTAIL.n321 VSUBS 0.023406f
C1184 VTAIL.n322 VSUBS 0.012577f
C1185 VTAIL.n323 VSUBS 0.029728f
C1186 VTAIL.n324 VSUBS 0.013317f
C1187 VTAIL.n325 VSUBS 0.023406f
C1188 VTAIL.n326 VSUBS 0.012577f
C1189 VTAIL.n327 VSUBS 0.029728f
C1190 VTAIL.n328 VSUBS 0.013317f
C1191 VTAIL.n329 VSUBS 1.76546f
C1192 VTAIL.n330 VSUBS 0.012577f
C1193 VTAIL.t15 VSUBS 0.06379f
C1194 VTAIL.n331 VSUBS 0.182595f
C1195 VTAIL.n332 VSUBS 0.018912f
C1196 VTAIL.n333 VSUBS 0.022296f
C1197 VTAIL.n334 VSUBS 0.029728f
C1198 VTAIL.n335 VSUBS 0.013317f
C1199 VTAIL.n336 VSUBS 0.012577f
C1200 VTAIL.n337 VSUBS 0.023406f
C1201 VTAIL.n338 VSUBS 0.023406f
C1202 VTAIL.n339 VSUBS 0.012577f
C1203 VTAIL.n340 VSUBS 0.013317f
C1204 VTAIL.n341 VSUBS 0.029728f
C1205 VTAIL.n342 VSUBS 0.029728f
C1206 VTAIL.n343 VSUBS 0.013317f
C1207 VTAIL.n344 VSUBS 0.012577f
C1208 VTAIL.n345 VSUBS 0.023406f
C1209 VTAIL.n346 VSUBS 0.023406f
C1210 VTAIL.n347 VSUBS 0.012577f
C1211 VTAIL.n348 VSUBS 0.013317f
C1212 VTAIL.n349 VSUBS 0.029728f
C1213 VTAIL.n350 VSUBS 0.029728f
C1214 VTAIL.n351 VSUBS 0.013317f
C1215 VTAIL.n352 VSUBS 0.012577f
C1216 VTAIL.n353 VSUBS 0.023406f
C1217 VTAIL.n354 VSUBS 0.023406f
C1218 VTAIL.n355 VSUBS 0.012577f
C1219 VTAIL.n356 VSUBS 0.013317f
C1220 VTAIL.n357 VSUBS 0.029728f
C1221 VTAIL.n358 VSUBS 0.029728f
C1222 VTAIL.n359 VSUBS 0.013317f
C1223 VTAIL.n360 VSUBS 0.012577f
C1224 VTAIL.n361 VSUBS 0.023406f
C1225 VTAIL.n362 VSUBS 0.023406f
C1226 VTAIL.n363 VSUBS 0.012577f
C1227 VTAIL.n364 VSUBS 0.013317f
C1228 VTAIL.n365 VSUBS 0.029728f
C1229 VTAIL.n366 VSUBS 0.029728f
C1230 VTAIL.n367 VSUBS 0.013317f
C1231 VTAIL.n368 VSUBS 0.012577f
C1232 VTAIL.n369 VSUBS 0.023406f
C1233 VTAIL.n370 VSUBS 0.023406f
C1234 VTAIL.n371 VSUBS 0.012577f
C1235 VTAIL.n372 VSUBS 0.013317f
C1236 VTAIL.n373 VSUBS 0.029728f
C1237 VTAIL.n374 VSUBS 0.029728f
C1238 VTAIL.n375 VSUBS 0.013317f
C1239 VTAIL.n376 VSUBS 0.012577f
C1240 VTAIL.n377 VSUBS 0.023406f
C1241 VTAIL.n378 VSUBS 0.023406f
C1242 VTAIL.n379 VSUBS 0.012577f
C1243 VTAIL.n380 VSUBS 0.013317f
C1244 VTAIL.n381 VSUBS 0.029728f
C1245 VTAIL.n382 VSUBS 0.029728f
C1246 VTAIL.n383 VSUBS 0.013317f
C1247 VTAIL.n384 VSUBS 0.012577f
C1248 VTAIL.n385 VSUBS 0.023406f
C1249 VTAIL.n386 VSUBS 0.023406f
C1250 VTAIL.n387 VSUBS 0.012577f
C1251 VTAIL.n388 VSUBS 0.013317f
C1252 VTAIL.n389 VSUBS 0.029728f
C1253 VTAIL.n390 VSUBS 0.071297f
C1254 VTAIL.n391 VSUBS 0.013317f
C1255 VTAIL.n392 VSUBS 0.012577f
C1256 VTAIL.n393 VSUBS 0.055061f
C1257 VTAIL.n394 VSUBS 0.035854f
C1258 VTAIL.n395 VSUBS 1.66415f
C1259 VTAIL.t9 VSUBS 0.324604f
C1260 VTAIL.t10 VSUBS 0.324604f
C1261 VTAIL.n396 VSUBS 2.54704f
C1262 VTAIL.n397 VSUBS 0.754006f
C1263 VTAIL.n398 VSUBS 0.025521f
C1264 VTAIL.n399 VSUBS 0.023406f
C1265 VTAIL.n400 VSUBS 0.012577f
C1266 VTAIL.n401 VSUBS 0.029728f
C1267 VTAIL.n402 VSUBS 0.013317f
C1268 VTAIL.n403 VSUBS 0.023406f
C1269 VTAIL.n404 VSUBS 0.012577f
C1270 VTAIL.n405 VSUBS 0.029728f
C1271 VTAIL.n406 VSUBS 0.012947f
C1272 VTAIL.n407 VSUBS 0.023406f
C1273 VTAIL.n408 VSUBS 0.012947f
C1274 VTAIL.n409 VSUBS 0.012577f
C1275 VTAIL.n410 VSUBS 0.029728f
C1276 VTAIL.n411 VSUBS 0.029728f
C1277 VTAIL.n412 VSUBS 0.013317f
C1278 VTAIL.n413 VSUBS 0.023406f
C1279 VTAIL.n414 VSUBS 0.012577f
C1280 VTAIL.n415 VSUBS 0.029728f
C1281 VTAIL.n416 VSUBS 0.013317f
C1282 VTAIL.n417 VSUBS 0.023406f
C1283 VTAIL.n418 VSUBS 0.012577f
C1284 VTAIL.n419 VSUBS 0.029728f
C1285 VTAIL.n420 VSUBS 0.013317f
C1286 VTAIL.n421 VSUBS 0.023406f
C1287 VTAIL.n422 VSUBS 0.012577f
C1288 VTAIL.n423 VSUBS 0.029728f
C1289 VTAIL.n424 VSUBS 0.013317f
C1290 VTAIL.n425 VSUBS 0.023406f
C1291 VTAIL.n426 VSUBS 0.012577f
C1292 VTAIL.n427 VSUBS 0.029728f
C1293 VTAIL.n428 VSUBS 0.013317f
C1294 VTAIL.n429 VSUBS 1.76546f
C1295 VTAIL.n430 VSUBS 0.012577f
C1296 VTAIL.t13 VSUBS 0.06379f
C1297 VTAIL.n431 VSUBS 0.182595f
C1298 VTAIL.n432 VSUBS 0.018912f
C1299 VTAIL.n433 VSUBS 0.022296f
C1300 VTAIL.n434 VSUBS 0.029728f
C1301 VTAIL.n435 VSUBS 0.013317f
C1302 VTAIL.n436 VSUBS 0.012577f
C1303 VTAIL.n437 VSUBS 0.023406f
C1304 VTAIL.n438 VSUBS 0.023406f
C1305 VTAIL.n439 VSUBS 0.012577f
C1306 VTAIL.n440 VSUBS 0.013317f
C1307 VTAIL.n441 VSUBS 0.029728f
C1308 VTAIL.n442 VSUBS 0.029728f
C1309 VTAIL.n443 VSUBS 0.013317f
C1310 VTAIL.n444 VSUBS 0.012577f
C1311 VTAIL.n445 VSUBS 0.023406f
C1312 VTAIL.n446 VSUBS 0.023406f
C1313 VTAIL.n447 VSUBS 0.012577f
C1314 VTAIL.n448 VSUBS 0.013317f
C1315 VTAIL.n449 VSUBS 0.029728f
C1316 VTAIL.n450 VSUBS 0.029728f
C1317 VTAIL.n451 VSUBS 0.013317f
C1318 VTAIL.n452 VSUBS 0.012577f
C1319 VTAIL.n453 VSUBS 0.023406f
C1320 VTAIL.n454 VSUBS 0.023406f
C1321 VTAIL.n455 VSUBS 0.012577f
C1322 VTAIL.n456 VSUBS 0.013317f
C1323 VTAIL.n457 VSUBS 0.029728f
C1324 VTAIL.n458 VSUBS 0.029728f
C1325 VTAIL.n459 VSUBS 0.013317f
C1326 VTAIL.n460 VSUBS 0.012577f
C1327 VTAIL.n461 VSUBS 0.023406f
C1328 VTAIL.n462 VSUBS 0.023406f
C1329 VTAIL.n463 VSUBS 0.012577f
C1330 VTAIL.n464 VSUBS 0.013317f
C1331 VTAIL.n465 VSUBS 0.029728f
C1332 VTAIL.n466 VSUBS 0.029728f
C1333 VTAIL.n467 VSUBS 0.013317f
C1334 VTAIL.n468 VSUBS 0.012577f
C1335 VTAIL.n469 VSUBS 0.023406f
C1336 VTAIL.n470 VSUBS 0.023406f
C1337 VTAIL.n471 VSUBS 0.012577f
C1338 VTAIL.n472 VSUBS 0.013317f
C1339 VTAIL.n473 VSUBS 0.029728f
C1340 VTAIL.n474 VSUBS 0.029728f
C1341 VTAIL.n475 VSUBS 0.013317f
C1342 VTAIL.n476 VSUBS 0.012577f
C1343 VTAIL.n477 VSUBS 0.023406f
C1344 VTAIL.n478 VSUBS 0.023406f
C1345 VTAIL.n479 VSUBS 0.012577f
C1346 VTAIL.n480 VSUBS 0.013317f
C1347 VTAIL.n481 VSUBS 0.029728f
C1348 VTAIL.n482 VSUBS 0.029728f
C1349 VTAIL.n483 VSUBS 0.013317f
C1350 VTAIL.n484 VSUBS 0.012577f
C1351 VTAIL.n485 VSUBS 0.023406f
C1352 VTAIL.n486 VSUBS 0.023406f
C1353 VTAIL.n487 VSUBS 0.012577f
C1354 VTAIL.n488 VSUBS 0.013317f
C1355 VTAIL.n489 VSUBS 0.029728f
C1356 VTAIL.n490 VSUBS 0.071297f
C1357 VTAIL.n491 VSUBS 0.013317f
C1358 VTAIL.n492 VSUBS 0.012577f
C1359 VTAIL.n493 VSUBS 0.055061f
C1360 VTAIL.n494 VSUBS 0.035854f
C1361 VTAIL.n495 VSUBS 0.148288f
C1362 VTAIL.n496 VSUBS 0.025521f
C1363 VTAIL.n497 VSUBS 0.023406f
C1364 VTAIL.n498 VSUBS 0.012577f
C1365 VTAIL.n499 VSUBS 0.029728f
C1366 VTAIL.n500 VSUBS 0.013317f
C1367 VTAIL.n501 VSUBS 0.023406f
C1368 VTAIL.n502 VSUBS 0.012577f
C1369 VTAIL.n503 VSUBS 0.029728f
C1370 VTAIL.n504 VSUBS 0.012947f
C1371 VTAIL.n505 VSUBS 0.023406f
C1372 VTAIL.n506 VSUBS 0.012947f
C1373 VTAIL.n507 VSUBS 0.012577f
C1374 VTAIL.n508 VSUBS 0.029728f
C1375 VTAIL.n509 VSUBS 0.029728f
C1376 VTAIL.n510 VSUBS 0.013317f
C1377 VTAIL.n511 VSUBS 0.023406f
C1378 VTAIL.n512 VSUBS 0.012577f
C1379 VTAIL.n513 VSUBS 0.029728f
C1380 VTAIL.n514 VSUBS 0.013317f
C1381 VTAIL.n515 VSUBS 0.023406f
C1382 VTAIL.n516 VSUBS 0.012577f
C1383 VTAIL.n517 VSUBS 0.029728f
C1384 VTAIL.n518 VSUBS 0.013317f
C1385 VTAIL.n519 VSUBS 0.023406f
C1386 VTAIL.n520 VSUBS 0.012577f
C1387 VTAIL.n521 VSUBS 0.029728f
C1388 VTAIL.n522 VSUBS 0.013317f
C1389 VTAIL.n523 VSUBS 0.023406f
C1390 VTAIL.n524 VSUBS 0.012577f
C1391 VTAIL.n525 VSUBS 0.029728f
C1392 VTAIL.n526 VSUBS 0.013317f
C1393 VTAIL.n527 VSUBS 1.76546f
C1394 VTAIL.n528 VSUBS 0.012577f
C1395 VTAIL.t2 VSUBS 0.06379f
C1396 VTAIL.n529 VSUBS 0.182595f
C1397 VTAIL.n530 VSUBS 0.018912f
C1398 VTAIL.n531 VSUBS 0.022296f
C1399 VTAIL.n532 VSUBS 0.029728f
C1400 VTAIL.n533 VSUBS 0.013317f
C1401 VTAIL.n534 VSUBS 0.012577f
C1402 VTAIL.n535 VSUBS 0.023406f
C1403 VTAIL.n536 VSUBS 0.023406f
C1404 VTAIL.n537 VSUBS 0.012577f
C1405 VTAIL.n538 VSUBS 0.013317f
C1406 VTAIL.n539 VSUBS 0.029728f
C1407 VTAIL.n540 VSUBS 0.029728f
C1408 VTAIL.n541 VSUBS 0.013317f
C1409 VTAIL.n542 VSUBS 0.012577f
C1410 VTAIL.n543 VSUBS 0.023406f
C1411 VTAIL.n544 VSUBS 0.023406f
C1412 VTAIL.n545 VSUBS 0.012577f
C1413 VTAIL.n546 VSUBS 0.013317f
C1414 VTAIL.n547 VSUBS 0.029728f
C1415 VTAIL.n548 VSUBS 0.029728f
C1416 VTAIL.n549 VSUBS 0.013317f
C1417 VTAIL.n550 VSUBS 0.012577f
C1418 VTAIL.n551 VSUBS 0.023406f
C1419 VTAIL.n552 VSUBS 0.023406f
C1420 VTAIL.n553 VSUBS 0.012577f
C1421 VTAIL.n554 VSUBS 0.013317f
C1422 VTAIL.n555 VSUBS 0.029728f
C1423 VTAIL.n556 VSUBS 0.029728f
C1424 VTAIL.n557 VSUBS 0.013317f
C1425 VTAIL.n558 VSUBS 0.012577f
C1426 VTAIL.n559 VSUBS 0.023406f
C1427 VTAIL.n560 VSUBS 0.023406f
C1428 VTAIL.n561 VSUBS 0.012577f
C1429 VTAIL.n562 VSUBS 0.013317f
C1430 VTAIL.n563 VSUBS 0.029728f
C1431 VTAIL.n564 VSUBS 0.029728f
C1432 VTAIL.n565 VSUBS 0.013317f
C1433 VTAIL.n566 VSUBS 0.012577f
C1434 VTAIL.n567 VSUBS 0.023406f
C1435 VTAIL.n568 VSUBS 0.023406f
C1436 VTAIL.n569 VSUBS 0.012577f
C1437 VTAIL.n570 VSUBS 0.013317f
C1438 VTAIL.n571 VSUBS 0.029728f
C1439 VTAIL.n572 VSUBS 0.029728f
C1440 VTAIL.n573 VSUBS 0.013317f
C1441 VTAIL.n574 VSUBS 0.012577f
C1442 VTAIL.n575 VSUBS 0.023406f
C1443 VTAIL.n576 VSUBS 0.023406f
C1444 VTAIL.n577 VSUBS 0.012577f
C1445 VTAIL.n578 VSUBS 0.013317f
C1446 VTAIL.n579 VSUBS 0.029728f
C1447 VTAIL.n580 VSUBS 0.029728f
C1448 VTAIL.n581 VSUBS 0.013317f
C1449 VTAIL.n582 VSUBS 0.012577f
C1450 VTAIL.n583 VSUBS 0.023406f
C1451 VTAIL.n584 VSUBS 0.023406f
C1452 VTAIL.n585 VSUBS 0.012577f
C1453 VTAIL.n586 VSUBS 0.013317f
C1454 VTAIL.n587 VSUBS 0.029728f
C1455 VTAIL.n588 VSUBS 0.071297f
C1456 VTAIL.n589 VSUBS 0.013317f
C1457 VTAIL.n590 VSUBS 0.012577f
C1458 VTAIL.n591 VSUBS 0.055061f
C1459 VTAIL.n592 VSUBS 0.035854f
C1460 VTAIL.n593 VSUBS 0.148288f
C1461 VTAIL.t5 VSUBS 0.324604f
C1462 VTAIL.t1 VSUBS 0.324604f
C1463 VTAIL.n594 VSUBS 2.54704f
C1464 VTAIL.n595 VSUBS 0.754006f
C1465 VTAIL.n596 VSUBS 0.025521f
C1466 VTAIL.n597 VSUBS 0.023406f
C1467 VTAIL.n598 VSUBS 0.012577f
C1468 VTAIL.n599 VSUBS 0.029728f
C1469 VTAIL.n600 VSUBS 0.013317f
C1470 VTAIL.n601 VSUBS 0.023406f
C1471 VTAIL.n602 VSUBS 0.012577f
C1472 VTAIL.n603 VSUBS 0.029728f
C1473 VTAIL.n604 VSUBS 0.012947f
C1474 VTAIL.n605 VSUBS 0.023406f
C1475 VTAIL.n606 VSUBS 0.012947f
C1476 VTAIL.n607 VSUBS 0.012577f
C1477 VTAIL.n608 VSUBS 0.029728f
C1478 VTAIL.n609 VSUBS 0.029728f
C1479 VTAIL.n610 VSUBS 0.013317f
C1480 VTAIL.n611 VSUBS 0.023406f
C1481 VTAIL.n612 VSUBS 0.012577f
C1482 VTAIL.n613 VSUBS 0.029728f
C1483 VTAIL.n614 VSUBS 0.013317f
C1484 VTAIL.n615 VSUBS 0.023406f
C1485 VTAIL.n616 VSUBS 0.012577f
C1486 VTAIL.n617 VSUBS 0.029728f
C1487 VTAIL.n618 VSUBS 0.013317f
C1488 VTAIL.n619 VSUBS 0.023406f
C1489 VTAIL.n620 VSUBS 0.012577f
C1490 VTAIL.n621 VSUBS 0.029728f
C1491 VTAIL.n622 VSUBS 0.013317f
C1492 VTAIL.n623 VSUBS 0.023406f
C1493 VTAIL.n624 VSUBS 0.012577f
C1494 VTAIL.n625 VSUBS 0.029728f
C1495 VTAIL.n626 VSUBS 0.013317f
C1496 VTAIL.n627 VSUBS 1.76546f
C1497 VTAIL.n628 VSUBS 0.012577f
C1498 VTAIL.t0 VSUBS 0.06379f
C1499 VTAIL.n629 VSUBS 0.182595f
C1500 VTAIL.n630 VSUBS 0.018912f
C1501 VTAIL.n631 VSUBS 0.022296f
C1502 VTAIL.n632 VSUBS 0.029728f
C1503 VTAIL.n633 VSUBS 0.013317f
C1504 VTAIL.n634 VSUBS 0.012577f
C1505 VTAIL.n635 VSUBS 0.023406f
C1506 VTAIL.n636 VSUBS 0.023406f
C1507 VTAIL.n637 VSUBS 0.012577f
C1508 VTAIL.n638 VSUBS 0.013317f
C1509 VTAIL.n639 VSUBS 0.029728f
C1510 VTAIL.n640 VSUBS 0.029728f
C1511 VTAIL.n641 VSUBS 0.013317f
C1512 VTAIL.n642 VSUBS 0.012577f
C1513 VTAIL.n643 VSUBS 0.023406f
C1514 VTAIL.n644 VSUBS 0.023406f
C1515 VTAIL.n645 VSUBS 0.012577f
C1516 VTAIL.n646 VSUBS 0.013317f
C1517 VTAIL.n647 VSUBS 0.029728f
C1518 VTAIL.n648 VSUBS 0.029728f
C1519 VTAIL.n649 VSUBS 0.013317f
C1520 VTAIL.n650 VSUBS 0.012577f
C1521 VTAIL.n651 VSUBS 0.023406f
C1522 VTAIL.n652 VSUBS 0.023406f
C1523 VTAIL.n653 VSUBS 0.012577f
C1524 VTAIL.n654 VSUBS 0.013317f
C1525 VTAIL.n655 VSUBS 0.029728f
C1526 VTAIL.n656 VSUBS 0.029728f
C1527 VTAIL.n657 VSUBS 0.013317f
C1528 VTAIL.n658 VSUBS 0.012577f
C1529 VTAIL.n659 VSUBS 0.023406f
C1530 VTAIL.n660 VSUBS 0.023406f
C1531 VTAIL.n661 VSUBS 0.012577f
C1532 VTAIL.n662 VSUBS 0.013317f
C1533 VTAIL.n663 VSUBS 0.029728f
C1534 VTAIL.n664 VSUBS 0.029728f
C1535 VTAIL.n665 VSUBS 0.013317f
C1536 VTAIL.n666 VSUBS 0.012577f
C1537 VTAIL.n667 VSUBS 0.023406f
C1538 VTAIL.n668 VSUBS 0.023406f
C1539 VTAIL.n669 VSUBS 0.012577f
C1540 VTAIL.n670 VSUBS 0.013317f
C1541 VTAIL.n671 VSUBS 0.029728f
C1542 VTAIL.n672 VSUBS 0.029728f
C1543 VTAIL.n673 VSUBS 0.013317f
C1544 VTAIL.n674 VSUBS 0.012577f
C1545 VTAIL.n675 VSUBS 0.023406f
C1546 VTAIL.n676 VSUBS 0.023406f
C1547 VTAIL.n677 VSUBS 0.012577f
C1548 VTAIL.n678 VSUBS 0.013317f
C1549 VTAIL.n679 VSUBS 0.029728f
C1550 VTAIL.n680 VSUBS 0.029728f
C1551 VTAIL.n681 VSUBS 0.013317f
C1552 VTAIL.n682 VSUBS 0.012577f
C1553 VTAIL.n683 VSUBS 0.023406f
C1554 VTAIL.n684 VSUBS 0.023406f
C1555 VTAIL.n685 VSUBS 0.012577f
C1556 VTAIL.n686 VSUBS 0.013317f
C1557 VTAIL.n687 VSUBS 0.029728f
C1558 VTAIL.n688 VSUBS 0.071297f
C1559 VTAIL.n689 VSUBS 0.013317f
C1560 VTAIL.n690 VSUBS 0.012577f
C1561 VTAIL.n691 VSUBS 0.055061f
C1562 VTAIL.n692 VSUBS 0.035854f
C1563 VTAIL.n693 VSUBS 1.66415f
C1564 VTAIL.n694 VSUBS 0.025521f
C1565 VTAIL.n695 VSUBS 0.023406f
C1566 VTAIL.n696 VSUBS 0.012577f
C1567 VTAIL.n697 VSUBS 0.029728f
C1568 VTAIL.n698 VSUBS 0.013317f
C1569 VTAIL.n699 VSUBS 0.023406f
C1570 VTAIL.n700 VSUBS 0.012577f
C1571 VTAIL.n701 VSUBS 0.029728f
C1572 VTAIL.n702 VSUBS 0.012947f
C1573 VTAIL.n703 VSUBS 0.023406f
C1574 VTAIL.n704 VSUBS 0.013317f
C1575 VTAIL.n705 VSUBS 0.029728f
C1576 VTAIL.n706 VSUBS 0.013317f
C1577 VTAIL.n707 VSUBS 0.023406f
C1578 VTAIL.n708 VSUBS 0.012577f
C1579 VTAIL.n709 VSUBS 0.029728f
C1580 VTAIL.n710 VSUBS 0.013317f
C1581 VTAIL.n711 VSUBS 0.023406f
C1582 VTAIL.n712 VSUBS 0.012577f
C1583 VTAIL.n713 VSUBS 0.029728f
C1584 VTAIL.n714 VSUBS 0.013317f
C1585 VTAIL.n715 VSUBS 0.023406f
C1586 VTAIL.n716 VSUBS 0.012577f
C1587 VTAIL.n717 VSUBS 0.029728f
C1588 VTAIL.n718 VSUBS 0.013317f
C1589 VTAIL.n719 VSUBS 0.023406f
C1590 VTAIL.n720 VSUBS 0.012577f
C1591 VTAIL.n721 VSUBS 0.029728f
C1592 VTAIL.n722 VSUBS 0.013317f
C1593 VTAIL.n723 VSUBS 1.76546f
C1594 VTAIL.n724 VSUBS 0.012577f
C1595 VTAIL.t12 VSUBS 0.06379f
C1596 VTAIL.n725 VSUBS 0.182595f
C1597 VTAIL.n726 VSUBS 0.018912f
C1598 VTAIL.n727 VSUBS 0.022296f
C1599 VTAIL.n728 VSUBS 0.029728f
C1600 VTAIL.n729 VSUBS 0.013317f
C1601 VTAIL.n730 VSUBS 0.012577f
C1602 VTAIL.n731 VSUBS 0.023406f
C1603 VTAIL.n732 VSUBS 0.023406f
C1604 VTAIL.n733 VSUBS 0.012577f
C1605 VTAIL.n734 VSUBS 0.013317f
C1606 VTAIL.n735 VSUBS 0.029728f
C1607 VTAIL.n736 VSUBS 0.029728f
C1608 VTAIL.n737 VSUBS 0.013317f
C1609 VTAIL.n738 VSUBS 0.012577f
C1610 VTAIL.n739 VSUBS 0.023406f
C1611 VTAIL.n740 VSUBS 0.023406f
C1612 VTAIL.n741 VSUBS 0.012577f
C1613 VTAIL.n742 VSUBS 0.013317f
C1614 VTAIL.n743 VSUBS 0.029728f
C1615 VTAIL.n744 VSUBS 0.029728f
C1616 VTAIL.n745 VSUBS 0.013317f
C1617 VTAIL.n746 VSUBS 0.012577f
C1618 VTAIL.n747 VSUBS 0.023406f
C1619 VTAIL.n748 VSUBS 0.023406f
C1620 VTAIL.n749 VSUBS 0.012577f
C1621 VTAIL.n750 VSUBS 0.013317f
C1622 VTAIL.n751 VSUBS 0.029728f
C1623 VTAIL.n752 VSUBS 0.029728f
C1624 VTAIL.n753 VSUBS 0.013317f
C1625 VTAIL.n754 VSUBS 0.012577f
C1626 VTAIL.n755 VSUBS 0.023406f
C1627 VTAIL.n756 VSUBS 0.023406f
C1628 VTAIL.n757 VSUBS 0.012577f
C1629 VTAIL.n758 VSUBS 0.013317f
C1630 VTAIL.n759 VSUBS 0.029728f
C1631 VTAIL.n760 VSUBS 0.029728f
C1632 VTAIL.n761 VSUBS 0.013317f
C1633 VTAIL.n762 VSUBS 0.012577f
C1634 VTAIL.n763 VSUBS 0.023406f
C1635 VTAIL.n764 VSUBS 0.023406f
C1636 VTAIL.n765 VSUBS 0.012577f
C1637 VTAIL.n766 VSUBS 0.012577f
C1638 VTAIL.n767 VSUBS 0.013317f
C1639 VTAIL.n768 VSUBS 0.029728f
C1640 VTAIL.n769 VSUBS 0.029728f
C1641 VTAIL.n770 VSUBS 0.029728f
C1642 VTAIL.n771 VSUBS 0.012947f
C1643 VTAIL.n772 VSUBS 0.012577f
C1644 VTAIL.n773 VSUBS 0.023406f
C1645 VTAIL.n774 VSUBS 0.023406f
C1646 VTAIL.n775 VSUBS 0.012577f
C1647 VTAIL.n776 VSUBS 0.013317f
C1648 VTAIL.n777 VSUBS 0.029728f
C1649 VTAIL.n778 VSUBS 0.029728f
C1650 VTAIL.n779 VSUBS 0.013317f
C1651 VTAIL.n780 VSUBS 0.012577f
C1652 VTAIL.n781 VSUBS 0.023406f
C1653 VTAIL.n782 VSUBS 0.023406f
C1654 VTAIL.n783 VSUBS 0.012577f
C1655 VTAIL.n784 VSUBS 0.013317f
C1656 VTAIL.n785 VSUBS 0.029728f
C1657 VTAIL.n786 VSUBS 0.071297f
C1658 VTAIL.n787 VSUBS 0.013317f
C1659 VTAIL.n788 VSUBS 0.012577f
C1660 VTAIL.n789 VSUBS 0.055061f
C1661 VTAIL.n790 VSUBS 0.035854f
C1662 VTAIL.n791 VSUBS 1.65976f
C1663 VN.n0 VSUBS 0.056227f
C1664 VN.t2 VSUBS 2.21606f
C1665 VN.n1 VSUBS 0.791761f
C1666 VN.n2 VSUBS 0.217753f
C1667 VN.t0 VSUBS 2.21606f
C1668 VN.t4 VSUBS 2.33028f
C1669 VN.n3 VSUBS 0.847745f
C1670 VN.n4 VSUBS 0.856375f
C1671 VN.n5 VSUBS 0.058411f
C1672 VN.n6 VSUBS 0.058411f
C1673 VN.n7 VSUBS 0.042137f
C1674 VN.n8 VSUBS 0.042137f
C1675 VN.n9 VSUBS 0.042863f
C1676 VN.n10 VSUBS 0.04906f
C1677 VN.t7 VSUBS 2.28643f
C1678 VN.n11 VSUBS 0.862267f
C1679 VN.n12 VSUBS 0.039463f
C1680 VN.n13 VSUBS 0.056227f
C1681 VN.t1 VSUBS 2.21606f
C1682 VN.n14 VSUBS 0.791761f
C1683 VN.n15 VSUBS 0.217753f
C1684 VN.t6 VSUBS 2.21606f
C1685 VN.t5 VSUBS 2.33028f
C1686 VN.n16 VSUBS 0.847745f
C1687 VN.n17 VSUBS 0.856375f
C1688 VN.n18 VSUBS 0.058411f
C1689 VN.n19 VSUBS 0.058411f
C1690 VN.n20 VSUBS 0.042137f
C1691 VN.n21 VSUBS 0.042137f
C1692 VN.n22 VSUBS 0.042863f
C1693 VN.n23 VSUBS 0.04906f
C1694 VN.t3 VSUBS 2.28643f
C1695 VN.n24 VSUBS 0.862267f
C1696 VN.n25 VSUBS 2.20379f
.ends

