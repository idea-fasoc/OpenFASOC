* NGSPICE file created from diff_pair_sample_0992.ext - technology: sky130A

.subckt diff_pair_sample_0992 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t2 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=1.6797 pd=10.51 as=3.9702 ps=21.14 w=10.18 l=3.99
X1 VDD2.t3 VN.t0 VTAIL.t0 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=1.6797 pd=10.51 as=3.9702 ps=21.14 w=10.18 l=3.99
X2 B.t11 B.t9 B.t10 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=3.9702 pd=21.14 as=0 ps=0 w=10.18 l=3.99
X3 VDD2.t2 VN.t1 VTAIL.t1 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=1.6797 pd=10.51 as=3.9702 ps=21.14 w=10.18 l=3.99
X4 VTAIL.t6 VN.t2 VDD2.t1 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=3.9702 pd=21.14 as=1.6797 ps=10.51 w=10.18 l=3.99
X5 VDD1.t2 VP.t1 VTAIL.t3 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=1.6797 pd=10.51 as=3.9702 ps=21.14 w=10.18 l=3.99
X6 VTAIL.t7 VN.t3 VDD2.t0 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=3.9702 pd=21.14 as=1.6797 ps=10.51 w=10.18 l=3.99
X7 B.t8 B.t6 B.t7 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=3.9702 pd=21.14 as=0 ps=0 w=10.18 l=3.99
X8 VTAIL.t5 VP.t2 VDD1.t1 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=3.9702 pd=21.14 as=1.6797 ps=10.51 w=10.18 l=3.99
X9 B.t5 B.t3 B.t4 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=3.9702 pd=21.14 as=0 ps=0 w=10.18 l=3.99
X10 B.t2 B.t0 B.t1 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=3.9702 pd=21.14 as=0 ps=0 w=10.18 l=3.99
X11 VTAIL.t4 VP.t3 VDD1.t0 w_n3562_n3004# sky130_fd_pr__pfet_01v8 ad=3.9702 pd=21.14 as=1.6797 ps=10.51 w=10.18 l=3.99
R0 VP.n18 VP.n0 161.3
R1 VP.n17 VP.n16 161.3
R2 VP.n15 VP.n1 161.3
R3 VP.n14 VP.n13 161.3
R4 VP.n12 VP.n2 161.3
R5 VP.n11 VP.n10 161.3
R6 VP.n9 VP.n3 161.3
R7 VP.n8 VP.n7 161.3
R8 VP.n4 VP.t2 95.3548
R9 VP.n4 VP.t1 93.9101
R10 VP.n6 VP.n5 62.2146
R11 VP.n20 VP.n19 62.2146
R12 VP.n6 VP.t3 61.4887
R13 VP.n19 VP.t0 61.4887
R14 VP.n13 VP.n12 56.5617
R15 VP.n5 VP.n4 51.0472
R16 VP.n7 VP.n3 24.5923
R17 VP.n11 VP.n3 24.5923
R18 VP.n12 VP.n11 24.5923
R19 VP.n13 VP.n1 24.5923
R20 VP.n17 VP.n1 24.5923
R21 VP.n18 VP.n17 24.5923
R22 VP.n7 VP.n6 20.1658
R23 VP.n19 VP.n18 20.1658
R24 VP.n8 VP.n5 0.417304
R25 VP.n20 VP.n0 0.417304
R26 VP VP.n20 0.394524
R27 VP.n9 VP.n8 0.189894
R28 VP.n10 VP.n9 0.189894
R29 VP.n10 VP.n2 0.189894
R30 VP.n14 VP.n2 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n16 VP.n15 0.189894
R33 VP.n16 VP.n0 0.189894
R34 VTAIL.n426 VTAIL.n378 756.745
R35 VTAIL.n48 VTAIL.n0 756.745
R36 VTAIL.n102 VTAIL.n54 756.745
R37 VTAIL.n156 VTAIL.n108 756.745
R38 VTAIL.n372 VTAIL.n324 756.745
R39 VTAIL.n318 VTAIL.n270 756.745
R40 VTAIL.n264 VTAIL.n216 756.745
R41 VTAIL.n210 VTAIL.n162 756.745
R42 VTAIL.n394 VTAIL.n393 585
R43 VTAIL.n399 VTAIL.n398 585
R44 VTAIL.n401 VTAIL.n400 585
R45 VTAIL.n390 VTAIL.n389 585
R46 VTAIL.n407 VTAIL.n406 585
R47 VTAIL.n409 VTAIL.n408 585
R48 VTAIL.n386 VTAIL.n385 585
R49 VTAIL.n416 VTAIL.n415 585
R50 VTAIL.n417 VTAIL.n384 585
R51 VTAIL.n419 VTAIL.n418 585
R52 VTAIL.n382 VTAIL.n381 585
R53 VTAIL.n425 VTAIL.n424 585
R54 VTAIL.n427 VTAIL.n426 585
R55 VTAIL.n16 VTAIL.n15 585
R56 VTAIL.n21 VTAIL.n20 585
R57 VTAIL.n23 VTAIL.n22 585
R58 VTAIL.n12 VTAIL.n11 585
R59 VTAIL.n29 VTAIL.n28 585
R60 VTAIL.n31 VTAIL.n30 585
R61 VTAIL.n8 VTAIL.n7 585
R62 VTAIL.n38 VTAIL.n37 585
R63 VTAIL.n39 VTAIL.n6 585
R64 VTAIL.n41 VTAIL.n40 585
R65 VTAIL.n4 VTAIL.n3 585
R66 VTAIL.n47 VTAIL.n46 585
R67 VTAIL.n49 VTAIL.n48 585
R68 VTAIL.n70 VTAIL.n69 585
R69 VTAIL.n75 VTAIL.n74 585
R70 VTAIL.n77 VTAIL.n76 585
R71 VTAIL.n66 VTAIL.n65 585
R72 VTAIL.n83 VTAIL.n82 585
R73 VTAIL.n85 VTAIL.n84 585
R74 VTAIL.n62 VTAIL.n61 585
R75 VTAIL.n92 VTAIL.n91 585
R76 VTAIL.n93 VTAIL.n60 585
R77 VTAIL.n95 VTAIL.n94 585
R78 VTAIL.n58 VTAIL.n57 585
R79 VTAIL.n101 VTAIL.n100 585
R80 VTAIL.n103 VTAIL.n102 585
R81 VTAIL.n124 VTAIL.n123 585
R82 VTAIL.n129 VTAIL.n128 585
R83 VTAIL.n131 VTAIL.n130 585
R84 VTAIL.n120 VTAIL.n119 585
R85 VTAIL.n137 VTAIL.n136 585
R86 VTAIL.n139 VTAIL.n138 585
R87 VTAIL.n116 VTAIL.n115 585
R88 VTAIL.n146 VTAIL.n145 585
R89 VTAIL.n147 VTAIL.n114 585
R90 VTAIL.n149 VTAIL.n148 585
R91 VTAIL.n112 VTAIL.n111 585
R92 VTAIL.n155 VTAIL.n154 585
R93 VTAIL.n157 VTAIL.n156 585
R94 VTAIL.n373 VTAIL.n372 585
R95 VTAIL.n371 VTAIL.n370 585
R96 VTAIL.n328 VTAIL.n327 585
R97 VTAIL.n365 VTAIL.n364 585
R98 VTAIL.n363 VTAIL.n330 585
R99 VTAIL.n362 VTAIL.n361 585
R100 VTAIL.n333 VTAIL.n331 585
R101 VTAIL.n356 VTAIL.n355 585
R102 VTAIL.n354 VTAIL.n353 585
R103 VTAIL.n337 VTAIL.n336 585
R104 VTAIL.n348 VTAIL.n347 585
R105 VTAIL.n346 VTAIL.n345 585
R106 VTAIL.n341 VTAIL.n340 585
R107 VTAIL.n319 VTAIL.n318 585
R108 VTAIL.n317 VTAIL.n316 585
R109 VTAIL.n274 VTAIL.n273 585
R110 VTAIL.n311 VTAIL.n310 585
R111 VTAIL.n309 VTAIL.n276 585
R112 VTAIL.n308 VTAIL.n307 585
R113 VTAIL.n279 VTAIL.n277 585
R114 VTAIL.n302 VTAIL.n301 585
R115 VTAIL.n300 VTAIL.n299 585
R116 VTAIL.n283 VTAIL.n282 585
R117 VTAIL.n294 VTAIL.n293 585
R118 VTAIL.n292 VTAIL.n291 585
R119 VTAIL.n287 VTAIL.n286 585
R120 VTAIL.n265 VTAIL.n264 585
R121 VTAIL.n263 VTAIL.n262 585
R122 VTAIL.n220 VTAIL.n219 585
R123 VTAIL.n257 VTAIL.n256 585
R124 VTAIL.n255 VTAIL.n222 585
R125 VTAIL.n254 VTAIL.n253 585
R126 VTAIL.n225 VTAIL.n223 585
R127 VTAIL.n248 VTAIL.n247 585
R128 VTAIL.n246 VTAIL.n245 585
R129 VTAIL.n229 VTAIL.n228 585
R130 VTAIL.n240 VTAIL.n239 585
R131 VTAIL.n238 VTAIL.n237 585
R132 VTAIL.n233 VTAIL.n232 585
R133 VTAIL.n211 VTAIL.n210 585
R134 VTAIL.n209 VTAIL.n208 585
R135 VTAIL.n166 VTAIL.n165 585
R136 VTAIL.n203 VTAIL.n202 585
R137 VTAIL.n201 VTAIL.n168 585
R138 VTAIL.n200 VTAIL.n199 585
R139 VTAIL.n171 VTAIL.n169 585
R140 VTAIL.n194 VTAIL.n193 585
R141 VTAIL.n192 VTAIL.n191 585
R142 VTAIL.n175 VTAIL.n174 585
R143 VTAIL.n186 VTAIL.n185 585
R144 VTAIL.n184 VTAIL.n183 585
R145 VTAIL.n179 VTAIL.n178 585
R146 VTAIL.n395 VTAIL.t0 329.038
R147 VTAIL.n17 VTAIL.t6 329.038
R148 VTAIL.n71 VTAIL.t2 329.038
R149 VTAIL.n125 VTAIL.t4 329.038
R150 VTAIL.n342 VTAIL.t3 329.038
R151 VTAIL.n288 VTAIL.t5 329.038
R152 VTAIL.n234 VTAIL.t1 329.038
R153 VTAIL.n180 VTAIL.t7 329.038
R154 VTAIL.n399 VTAIL.n393 171.744
R155 VTAIL.n400 VTAIL.n399 171.744
R156 VTAIL.n400 VTAIL.n389 171.744
R157 VTAIL.n407 VTAIL.n389 171.744
R158 VTAIL.n408 VTAIL.n407 171.744
R159 VTAIL.n408 VTAIL.n385 171.744
R160 VTAIL.n416 VTAIL.n385 171.744
R161 VTAIL.n417 VTAIL.n416 171.744
R162 VTAIL.n418 VTAIL.n417 171.744
R163 VTAIL.n418 VTAIL.n381 171.744
R164 VTAIL.n425 VTAIL.n381 171.744
R165 VTAIL.n426 VTAIL.n425 171.744
R166 VTAIL.n21 VTAIL.n15 171.744
R167 VTAIL.n22 VTAIL.n21 171.744
R168 VTAIL.n22 VTAIL.n11 171.744
R169 VTAIL.n29 VTAIL.n11 171.744
R170 VTAIL.n30 VTAIL.n29 171.744
R171 VTAIL.n30 VTAIL.n7 171.744
R172 VTAIL.n38 VTAIL.n7 171.744
R173 VTAIL.n39 VTAIL.n38 171.744
R174 VTAIL.n40 VTAIL.n39 171.744
R175 VTAIL.n40 VTAIL.n3 171.744
R176 VTAIL.n47 VTAIL.n3 171.744
R177 VTAIL.n48 VTAIL.n47 171.744
R178 VTAIL.n75 VTAIL.n69 171.744
R179 VTAIL.n76 VTAIL.n75 171.744
R180 VTAIL.n76 VTAIL.n65 171.744
R181 VTAIL.n83 VTAIL.n65 171.744
R182 VTAIL.n84 VTAIL.n83 171.744
R183 VTAIL.n84 VTAIL.n61 171.744
R184 VTAIL.n92 VTAIL.n61 171.744
R185 VTAIL.n93 VTAIL.n92 171.744
R186 VTAIL.n94 VTAIL.n93 171.744
R187 VTAIL.n94 VTAIL.n57 171.744
R188 VTAIL.n101 VTAIL.n57 171.744
R189 VTAIL.n102 VTAIL.n101 171.744
R190 VTAIL.n129 VTAIL.n123 171.744
R191 VTAIL.n130 VTAIL.n129 171.744
R192 VTAIL.n130 VTAIL.n119 171.744
R193 VTAIL.n137 VTAIL.n119 171.744
R194 VTAIL.n138 VTAIL.n137 171.744
R195 VTAIL.n138 VTAIL.n115 171.744
R196 VTAIL.n146 VTAIL.n115 171.744
R197 VTAIL.n147 VTAIL.n146 171.744
R198 VTAIL.n148 VTAIL.n147 171.744
R199 VTAIL.n148 VTAIL.n111 171.744
R200 VTAIL.n155 VTAIL.n111 171.744
R201 VTAIL.n156 VTAIL.n155 171.744
R202 VTAIL.n372 VTAIL.n371 171.744
R203 VTAIL.n371 VTAIL.n327 171.744
R204 VTAIL.n364 VTAIL.n327 171.744
R205 VTAIL.n364 VTAIL.n363 171.744
R206 VTAIL.n363 VTAIL.n362 171.744
R207 VTAIL.n362 VTAIL.n331 171.744
R208 VTAIL.n355 VTAIL.n331 171.744
R209 VTAIL.n355 VTAIL.n354 171.744
R210 VTAIL.n354 VTAIL.n336 171.744
R211 VTAIL.n347 VTAIL.n336 171.744
R212 VTAIL.n347 VTAIL.n346 171.744
R213 VTAIL.n346 VTAIL.n340 171.744
R214 VTAIL.n318 VTAIL.n317 171.744
R215 VTAIL.n317 VTAIL.n273 171.744
R216 VTAIL.n310 VTAIL.n273 171.744
R217 VTAIL.n310 VTAIL.n309 171.744
R218 VTAIL.n309 VTAIL.n308 171.744
R219 VTAIL.n308 VTAIL.n277 171.744
R220 VTAIL.n301 VTAIL.n277 171.744
R221 VTAIL.n301 VTAIL.n300 171.744
R222 VTAIL.n300 VTAIL.n282 171.744
R223 VTAIL.n293 VTAIL.n282 171.744
R224 VTAIL.n293 VTAIL.n292 171.744
R225 VTAIL.n292 VTAIL.n286 171.744
R226 VTAIL.n264 VTAIL.n263 171.744
R227 VTAIL.n263 VTAIL.n219 171.744
R228 VTAIL.n256 VTAIL.n219 171.744
R229 VTAIL.n256 VTAIL.n255 171.744
R230 VTAIL.n255 VTAIL.n254 171.744
R231 VTAIL.n254 VTAIL.n223 171.744
R232 VTAIL.n247 VTAIL.n223 171.744
R233 VTAIL.n247 VTAIL.n246 171.744
R234 VTAIL.n246 VTAIL.n228 171.744
R235 VTAIL.n239 VTAIL.n228 171.744
R236 VTAIL.n239 VTAIL.n238 171.744
R237 VTAIL.n238 VTAIL.n232 171.744
R238 VTAIL.n210 VTAIL.n209 171.744
R239 VTAIL.n209 VTAIL.n165 171.744
R240 VTAIL.n202 VTAIL.n165 171.744
R241 VTAIL.n202 VTAIL.n201 171.744
R242 VTAIL.n201 VTAIL.n200 171.744
R243 VTAIL.n200 VTAIL.n169 171.744
R244 VTAIL.n193 VTAIL.n169 171.744
R245 VTAIL.n193 VTAIL.n192 171.744
R246 VTAIL.n192 VTAIL.n174 171.744
R247 VTAIL.n185 VTAIL.n174 171.744
R248 VTAIL.n185 VTAIL.n184 171.744
R249 VTAIL.n184 VTAIL.n178 171.744
R250 VTAIL.t0 VTAIL.n393 85.8723
R251 VTAIL.t6 VTAIL.n15 85.8723
R252 VTAIL.t2 VTAIL.n69 85.8723
R253 VTAIL.t4 VTAIL.n123 85.8723
R254 VTAIL.t3 VTAIL.n340 85.8723
R255 VTAIL.t5 VTAIL.n286 85.8723
R256 VTAIL.t1 VTAIL.n232 85.8723
R257 VTAIL.t7 VTAIL.n178 85.8723
R258 VTAIL.n431 VTAIL.n430 36.452
R259 VTAIL.n53 VTAIL.n52 36.452
R260 VTAIL.n107 VTAIL.n106 36.452
R261 VTAIL.n161 VTAIL.n160 36.452
R262 VTAIL.n377 VTAIL.n376 36.452
R263 VTAIL.n323 VTAIL.n322 36.452
R264 VTAIL.n269 VTAIL.n268 36.452
R265 VTAIL.n215 VTAIL.n214 36.452
R266 VTAIL.n431 VTAIL.n377 24.8669
R267 VTAIL.n215 VTAIL.n161 24.8669
R268 VTAIL.n419 VTAIL.n384 13.1884
R269 VTAIL.n41 VTAIL.n6 13.1884
R270 VTAIL.n95 VTAIL.n60 13.1884
R271 VTAIL.n149 VTAIL.n114 13.1884
R272 VTAIL.n365 VTAIL.n330 13.1884
R273 VTAIL.n311 VTAIL.n276 13.1884
R274 VTAIL.n257 VTAIL.n222 13.1884
R275 VTAIL.n203 VTAIL.n168 13.1884
R276 VTAIL.n415 VTAIL.n414 12.8005
R277 VTAIL.n420 VTAIL.n382 12.8005
R278 VTAIL.n37 VTAIL.n36 12.8005
R279 VTAIL.n42 VTAIL.n4 12.8005
R280 VTAIL.n91 VTAIL.n90 12.8005
R281 VTAIL.n96 VTAIL.n58 12.8005
R282 VTAIL.n145 VTAIL.n144 12.8005
R283 VTAIL.n150 VTAIL.n112 12.8005
R284 VTAIL.n366 VTAIL.n328 12.8005
R285 VTAIL.n361 VTAIL.n332 12.8005
R286 VTAIL.n312 VTAIL.n274 12.8005
R287 VTAIL.n307 VTAIL.n278 12.8005
R288 VTAIL.n258 VTAIL.n220 12.8005
R289 VTAIL.n253 VTAIL.n224 12.8005
R290 VTAIL.n204 VTAIL.n166 12.8005
R291 VTAIL.n199 VTAIL.n170 12.8005
R292 VTAIL.n413 VTAIL.n386 12.0247
R293 VTAIL.n424 VTAIL.n423 12.0247
R294 VTAIL.n35 VTAIL.n8 12.0247
R295 VTAIL.n46 VTAIL.n45 12.0247
R296 VTAIL.n89 VTAIL.n62 12.0247
R297 VTAIL.n100 VTAIL.n99 12.0247
R298 VTAIL.n143 VTAIL.n116 12.0247
R299 VTAIL.n154 VTAIL.n153 12.0247
R300 VTAIL.n370 VTAIL.n369 12.0247
R301 VTAIL.n360 VTAIL.n333 12.0247
R302 VTAIL.n316 VTAIL.n315 12.0247
R303 VTAIL.n306 VTAIL.n279 12.0247
R304 VTAIL.n262 VTAIL.n261 12.0247
R305 VTAIL.n252 VTAIL.n225 12.0247
R306 VTAIL.n208 VTAIL.n207 12.0247
R307 VTAIL.n198 VTAIL.n171 12.0247
R308 VTAIL.n410 VTAIL.n409 11.249
R309 VTAIL.n427 VTAIL.n380 11.249
R310 VTAIL.n32 VTAIL.n31 11.249
R311 VTAIL.n49 VTAIL.n2 11.249
R312 VTAIL.n86 VTAIL.n85 11.249
R313 VTAIL.n103 VTAIL.n56 11.249
R314 VTAIL.n140 VTAIL.n139 11.249
R315 VTAIL.n157 VTAIL.n110 11.249
R316 VTAIL.n373 VTAIL.n326 11.249
R317 VTAIL.n357 VTAIL.n356 11.249
R318 VTAIL.n319 VTAIL.n272 11.249
R319 VTAIL.n303 VTAIL.n302 11.249
R320 VTAIL.n265 VTAIL.n218 11.249
R321 VTAIL.n249 VTAIL.n248 11.249
R322 VTAIL.n211 VTAIL.n164 11.249
R323 VTAIL.n195 VTAIL.n194 11.249
R324 VTAIL.n395 VTAIL.n394 10.7239
R325 VTAIL.n17 VTAIL.n16 10.7239
R326 VTAIL.n71 VTAIL.n70 10.7239
R327 VTAIL.n125 VTAIL.n124 10.7239
R328 VTAIL.n342 VTAIL.n341 10.7239
R329 VTAIL.n288 VTAIL.n287 10.7239
R330 VTAIL.n234 VTAIL.n233 10.7239
R331 VTAIL.n180 VTAIL.n179 10.7239
R332 VTAIL.n406 VTAIL.n388 10.4732
R333 VTAIL.n428 VTAIL.n378 10.4732
R334 VTAIL.n28 VTAIL.n10 10.4732
R335 VTAIL.n50 VTAIL.n0 10.4732
R336 VTAIL.n82 VTAIL.n64 10.4732
R337 VTAIL.n104 VTAIL.n54 10.4732
R338 VTAIL.n136 VTAIL.n118 10.4732
R339 VTAIL.n158 VTAIL.n108 10.4732
R340 VTAIL.n374 VTAIL.n324 10.4732
R341 VTAIL.n353 VTAIL.n335 10.4732
R342 VTAIL.n320 VTAIL.n270 10.4732
R343 VTAIL.n299 VTAIL.n281 10.4732
R344 VTAIL.n266 VTAIL.n216 10.4732
R345 VTAIL.n245 VTAIL.n227 10.4732
R346 VTAIL.n212 VTAIL.n162 10.4732
R347 VTAIL.n191 VTAIL.n173 10.4732
R348 VTAIL.n405 VTAIL.n390 9.69747
R349 VTAIL.n27 VTAIL.n12 9.69747
R350 VTAIL.n81 VTAIL.n66 9.69747
R351 VTAIL.n135 VTAIL.n120 9.69747
R352 VTAIL.n352 VTAIL.n337 9.69747
R353 VTAIL.n298 VTAIL.n283 9.69747
R354 VTAIL.n244 VTAIL.n229 9.69747
R355 VTAIL.n190 VTAIL.n175 9.69747
R356 VTAIL.n430 VTAIL.n429 9.45567
R357 VTAIL.n52 VTAIL.n51 9.45567
R358 VTAIL.n106 VTAIL.n105 9.45567
R359 VTAIL.n160 VTAIL.n159 9.45567
R360 VTAIL.n376 VTAIL.n375 9.45567
R361 VTAIL.n322 VTAIL.n321 9.45567
R362 VTAIL.n268 VTAIL.n267 9.45567
R363 VTAIL.n214 VTAIL.n213 9.45567
R364 VTAIL.n429 VTAIL.n428 9.3005
R365 VTAIL.n380 VTAIL.n379 9.3005
R366 VTAIL.n423 VTAIL.n422 9.3005
R367 VTAIL.n421 VTAIL.n420 9.3005
R368 VTAIL.n397 VTAIL.n396 9.3005
R369 VTAIL.n392 VTAIL.n391 9.3005
R370 VTAIL.n403 VTAIL.n402 9.3005
R371 VTAIL.n405 VTAIL.n404 9.3005
R372 VTAIL.n388 VTAIL.n387 9.3005
R373 VTAIL.n411 VTAIL.n410 9.3005
R374 VTAIL.n413 VTAIL.n412 9.3005
R375 VTAIL.n414 VTAIL.n383 9.3005
R376 VTAIL.n51 VTAIL.n50 9.3005
R377 VTAIL.n2 VTAIL.n1 9.3005
R378 VTAIL.n45 VTAIL.n44 9.3005
R379 VTAIL.n43 VTAIL.n42 9.3005
R380 VTAIL.n19 VTAIL.n18 9.3005
R381 VTAIL.n14 VTAIL.n13 9.3005
R382 VTAIL.n25 VTAIL.n24 9.3005
R383 VTAIL.n27 VTAIL.n26 9.3005
R384 VTAIL.n10 VTAIL.n9 9.3005
R385 VTAIL.n33 VTAIL.n32 9.3005
R386 VTAIL.n35 VTAIL.n34 9.3005
R387 VTAIL.n36 VTAIL.n5 9.3005
R388 VTAIL.n105 VTAIL.n104 9.3005
R389 VTAIL.n56 VTAIL.n55 9.3005
R390 VTAIL.n99 VTAIL.n98 9.3005
R391 VTAIL.n97 VTAIL.n96 9.3005
R392 VTAIL.n73 VTAIL.n72 9.3005
R393 VTAIL.n68 VTAIL.n67 9.3005
R394 VTAIL.n79 VTAIL.n78 9.3005
R395 VTAIL.n81 VTAIL.n80 9.3005
R396 VTAIL.n64 VTAIL.n63 9.3005
R397 VTAIL.n87 VTAIL.n86 9.3005
R398 VTAIL.n89 VTAIL.n88 9.3005
R399 VTAIL.n90 VTAIL.n59 9.3005
R400 VTAIL.n159 VTAIL.n158 9.3005
R401 VTAIL.n110 VTAIL.n109 9.3005
R402 VTAIL.n153 VTAIL.n152 9.3005
R403 VTAIL.n151 VTAIL.n150 9.3005
R404 VTAIL.n127 VTAIL.n126 9.3005
R405 VTAIL.n122 VTAIL.n121 9.3005
R406 VTAIL.n133 VTAIL.n132 9.3005
R407 VTAIL.n135 VTAIL.n134 9.3005
R408 VTAIL.n118 VTAIL.n117 9.3005
R409 VTAIL.n141 VTAIL.n140 9.3005
R410 VTAIL.n143 VTAIL.n142 9.3005
R411 VTAIL.n144 VTAIL.n113 9.3005
R412 VTAIL.n344 VTAIL.n343 9.3005
R413 VTAIL.n339 VTAIL.n338 9.3005
R414 VTAIL.n350 VTAIL.n349 9.3005
R415 VTAIL.n352 VTAIL.n351 9.3005
R416 VTAIL.n335 VTAIL.n334 9.3005
R417 VTAIL.n358 VTAIL.n357 9.3005
R418 VTAIL.n360 VTAIL.n359 9.3005
R419 VTAIL.n332 VTAIL.n329 9.3005
R420 VTAIL.n375 VTAIL.n374 9.3005
R421 VTAIL.n326 VTAIL.n325 9.3005
R422 VTAIL.n369 VTAIL.n368 9.3005
R423 VTAIL.n367 VTAIL.n366 9.3005
R424 VTAIL.n290 VTAIL.n289 9.3005
R425 VTAIL.n285 VTAIL.n284 9.3005
R426 VTAIL.n296 VTAIL.n295 9.3005
R427 VTAIL.n298 VTAIL.n297 9.3005
R428 VTAIL.n281 VTAIL.n280 9.3005
R429 VTAIL.n304 VTAIL.n303 9.3005
R430 VTAIL.n306 VTAIL.n305 9.3005
R431 VTAIL.n278 VTAIL.n275 9.3005
R432 VTAIL.n321 VTAIL.n320 9.3005
R433 VTAIL.n272 VTAIL.n271 9.3005
R434 VTAIL.n315 VTAIL.n314 9.3005
R435 VTAIL.n313 VTAIL.n312 9.3005
R436 VTAIL.n236 VTAIL.n235 9.3005
R437 VTAIL.n231 VTAIL.n230 9.3005
R438 VTAIL.n242 VTAIL.n241 9.3005
R439 VTAIL.n244 VTAIL.n243 9.3005
R440 VTAIL.n227 VTAIL.n226 9.3005
R441 VTAIL.n250 VTAIL.n249 9.3005
R442 VTAIL.n252 VTAIL.n251 9.3005
R443 VTAIL.n224 VTAIL.n221 9.3005
R444 VTAIL.n267 VTAIL.n266 9.3005
R445 VTAIL.n218 VTAIL.n217 9.3005
R446 VTAIL.n261 VTAIL.n260 9.3005
R447 VTAIL.n259 VTAIL.n258 9.3005
R448 VTAIL.n182 VTAIL.n181 9.3005
R449 VTAIL.n177 VTAIL.n176 9.3005
R450 VTAIL.n188 VTAIL.n187 9.3005
R451 VTAIL.n190 VTAIL.n189 9.3005
R452 VTAIL.n173 VTAIL.n172 9.3005
R453 VTAIL.n196 VTAIL.n195 9.3005
R454 VTAIL.n198 VTAIL.n197 9.3005
R455 VTAIL.n170 VTAIL.n167 9.3005
R456 VTAIL.n213 VTAIL.n212 9.3005
R457 VTAIL.n164 VTAIL.n163 9.3005
R458 VTAIL.n207 VTAIL.n206 9.3005
R459 VTAIL.n205 VTAIL.n204 9.3005
R460 VTAIL.n402 VTAIL.n401 8.92171
R461 VTAIL.n24 VTAIL.n23 8.92171
R462 VTAIL.n78 VTAIL.n77 8.92171
R463 VTAIL.n132 VTAIL.n131 8.92171
R464 VTAIL.n349 VTAIL.n348 8.92171
R465 VTAIL.n295 VTAIL.n294 8.92171
R466 VTAIL.n241 VTAIL.n240 8.92171
R467 VTAIL.n187 VTAIL.n186 8.92171
R468 VTAIL.n398 VTAIL.n392 8.14595
R469 VTAIL.n20 VTAIL.n14 8.14595
R470 VTAIL.n74 VTAIL.n68 8.14595
R471 VTAIL.n128 VTAIL.n122 8.14595
R472 VTAIL.n345 VTAIL.n339 8.14595
R473 VTAIL.n291 VTAIL.n285 8.14595
R474 VTAIL.n237 VTAIL.n231 8.14595
R475 VTAIL.n183 VTAIL.n177 8.14595
R476 VTAIL.n397 VTAIL.n394 7.3702
R477 VTAIL.n19 VTAIL.n16 7.3702
R478 VTAIL.n73 VTAIL.n70 7.3702
R479 VTAIL.n127 VTAIL.n124 7.3702
R480 VTAIL.n344 VTAIL.n341 7.3702
R481 VTAIL.n290 VTAIL.n287 7.3702
R482 VTAIL.n236 VTAIL.n233 7.3702
R483 VTAIL.n182 VTAIL.n179 7.3702
R484 VTAIL.n398 VTAIL.n397 5.81868
R485 VTAIL.n20 VTAIL.n19 5.81868
R486 VTAIL.n74 VTAIL.n73 5.81868
R487 VTAIL.n128 VTAIL.n127 5.81868
R488 VTAIL.n345 VTAIL.n344 5.81868
R489 VTAIL.n291 VTAIL.n290 5.81868
R490 VTAIL.n237 VTAIL.n236 5.81868
R491 VTAIL.n183 VTAIL.n182 5.81868
R492 VTAIL.n401 VTAIL.n392 5.04292
R493 VTAIL.n23 VTAIL.n14 5.04292
R494 VTAIL.n77 VTAIL.n68 5.04292
R495 VTAIL.n131 VTAIL.n122 5.04292
R496 VTAIL.n348 VTAIL.n339 5.04292
R497 VTAIL.n294 VTAIL.n285 5.04292
R498 VTAIL.n240 VTAIL.n231 5.04292
R499 VTAIL.n186 VTAIL.n177 5.04292
R500 VTAIL.n402 VTAIL.n390 4.26717
R501 VTAIL.n24 VTAIL.n12 4.26717
R502 VTAIL.n78 VTAIL.n66 4.26717
R503 VTAIL.n132 VTAIL.n120 4.26717
R504 VTAIL.n349 VTAIL.n337 4.26717
R505 VTAIL.n295 VTAIL.n283 4.26717
R506 VTAIL.n241 VTAIL.n229 4.26717
R507 VTAIL.n187 VTAIL.n175 4.26717
R508 VTAIL.n269 VTAIL.n215 3.72464
R509 VTAIL.n377 VTAIL.n323 3.72464
R510 VTAIL.n161 VTAIL.n107 3.72464
R511 VTAIL.n406 VTAIL.n405 3.49141
R512 VTAIL.n430 VTAIL.n378 3.49141
R513 VTAIL.n28 VTAIL.n27 3.49141
R514 VTAIL.n52 VTAIL.n0 3.49141
R515 VTAIL.n82 VTAIL.n81 3.49141
R516 VTAIL.n106 VTAIL.n54 3.49141
R517 VTAIL.n136 VTAIL.n135 3.49141
R518 VTAIL.n160 VTAIL.n108 3.49141
R519 VTAIL.n376 VTAIL.n324 3.49141
R520 VTAIL.n353 VTAIL.n352 3.49141
R521 VTAIL.n322 VTAIL.n270 3.49141
R522 VTAIL.n299 VTAIL.n298 3.49141
R523 VTAIL.n268 VTAIL.n216 3.49141
R524 VTAIL.n245 VTAIL.n244 3.49141
R525 VTAIL.n214 VTAIL.n162 3.49141
R526 VTAIL.n191 VTAIL.n190 3.49141
R527 VTAIL.n409 VTAIL.n388 2.71565
R528 VTAIL.n428 VTAIL.n427 2.71565
R529 VTAIL.n31 VTAIL.n10 2.71565
R530 VTAIL.n50 VTAIL.n49 2.71565
R531 VTAIL.n85 VTAIL.n64 2.71565
R532 VTAIL.n104 VTAIL.n103 2.71565
R533 VTAIL.n139 VTAIL.n118 2.71565
R534 VTAIL.n158 VTAIL.n157 2.71565
R535 VTAIL.n374 VTAIL.n373 2.71565
R536 VTAIL.n356 VTAIL.n335 2.71565
R537 VTAIL.n320 VTAIL.n319 2.71565
R538 VTAIL.n302 VTAIL.n281 2.71565
R539 VTAIL.n266 VTAIL.n265 2.71565
R540 VTAIL.n248 VTAIL.n227 2.71565
R541 VTAIL.n212 VTAIL.n211 2.71565
R542 VTAIL.n194 VTAIL.n173 2.71565
R543 VTAIL.n396 VTAIL.n395 2.41283
R544 VTAIL.n18 VTAIL.n17 2.41283
R545 VTAIL.n72 VTAIL.n71 2.41283
R546 VTAIL.n126 VTAIL.n125 2.41283
R547 VTAIL.n343 VTAIL.n342 2.41283
R548 VTAIL.n289 VTAIL.n288 2.41283
R549 VTAIL.n235 VTAIL.n234 2.41283
R550 VTAIL.n181 VTAIL.n180 2.41283
R551 VTAIL.n410 VTAIL.n386 1.93989
R552 VTAIL.n424 VTAIL.n380 1.93989
R553 VTAIL.n32 VTAIL.n8 1.93989
R554 VTAIL.n46 VTAIL.n2 1.93989
R555 VTAIL.n86 VTAIL.n62 1.93989
R556 VTAIL.n100 VTAIL.n56 1.93989
R557 VTAIL.n140 VTAIL.n116 1.93989
R558 VTAIL.n154 VTAIL.n110 1.93989
R559 VTAIL.n370 VTAIL.n326 1.93989
R560 VTAIL.n357 VTAIL.n333 1.93989
R561 VTAIL.n316 VTAIL.n272 1.93989
R562 VTAIL.n303 VTAIL.n279 1.93989
R563 VTAIL.n262 VTAIL.n218 1.93989
R564 VTAIL.n249 VTAIL.n225 1.93989
R565 VTAIL.n208 VTAIL.n164 1.93989
R566 VTAIL.n195 VTAIL.n171 1.93989
R567 VTAIL VTAIL.n53 1.92076
R568 VTAIL VTAIL.n431 1.80438
R569 VTAIL.n415 VTAIL.n413 1.16414
R570 VTAIL.n423 VTAIL.n382 1.16414
R571 VTAIL.n37 VTAIL.n35 1.16414
R572 VTAIL.n45 VTAIL.n4 1.16414
R573 VTAIL.n91 VTAIL.n89 1.16414
R574 VTAIL.n99 VTAIL.n58 1.16414
R575 VTAIL.n145 VTAIL.n143 1.16414
R576 VTAIL.n153 VTAIL.n112 1.16414
R577 VTAIL.n369 VTAIL.n328 1.16414
R578 VTAIL.n361 VTAIL.n360 1.16414
R579 VTAIL.n315 VTAIL.n274 1.16414
R580 VTAIL.n307 VTAIL.n306 1.16414
R581 VTAIL.n261 VTAIL.n220 1.16414
R582 VTAIL.n253 VTAIL.n252 1.16414
R583 VTAIL.n207 VTAIL.n166 1.16414
R584 VTAIL.n199 VTAIL.n198 1.16414
R585 VTAIL.n323 VTAIL.n269 0.470328
R586 VTAIL.n107 VTAIL.n53 0.470328
R587 VTAIL.n414 VTAIL.n384 0.388379
R588 VTAIL.n420 VTAIL.n419 0.388379
R589 VTAIL.n36 VTAIL.n6 0.388379
R590 VTAIL.n42 VTAIL.n41 0.388379
R591 VTAIL.n90 VTAIL.n60 0.388379
R592 VTAIL.n96 VTAIL.n95 0.388379
R593 VTAIL.n144 VTAIL.n114 0.388379
R594 VTAIL.n150 VTAIL.n149 0.388379
R595 VTAIL.n366 VTAIL.n365 0.388379
R596 VTAIL.n332 VTAIL.n330 0.388379
R597 VTAIL.n312 VTAIL.n311 0.388379
R598 VTAIL.n278 VTAIL.n276 0.388379
R599 VTAIL.n258 VTAIL.n257 0.388379
R600 VTAIL.n224 VTAIL.n222 0.388379
R601 VTAIL.n204 VTAIL.n203 0.388379
R602 VTAIL.n170 VTAIL.n168 0.388379
R603 VTAIL.n396 VTAIL.n391 0.155672
R604 VTAIL.n403 VTAIL.n391 0.155672
R605 VTAIL.n404 VTAIL.n403 0.155672
R606 VTAIL.n404 VTAIL.n387 0.155672
R607 VTAIL.n411 VTAIL.n387 0.155672
R608 VTAIL.n412 VTAIL.n411 0.155672
R609 VTAIL.n412 VTAIL.n383 0.155672
R610 VTAIL.n421 VTAIL.n383 0.155672
R611 VTAIL.n422 VTAIL.n421 0.155672
R612 VTAIL.n422 VTAIL.n379 0.155672
R613 VTAIL.n429 VTAIL.n379 0.155672
R614 VTAIL.n18 VTAIL.n13 0.155672
R615 VTAIL.n25 VTAIL.n13 0.155672
R616 VTAIL.n26 VTAIL.n25 0.155672
R617 VTAIL.n26 VTAIL.n9 0.155672
R618 VTAIL.n33 VTAIL.n9 0.155672
R619 VTAIL.n34 VTAIL.n33 0.155672
R620 VTAIL.n34 VTAIL.n5 0.155672
R621 VTAIL.n43 VTAIL.n5 0.155672
R622 VTAIL.n44 VTAIL.n43 0.155672
R623 VTAIL.n44 VTAIL.n1 0.155672
R624 VTAIL.n51 VTAIL.n1 0.155672
R625 VTAIL.n72 VTAIL.n67 0.155672
R626 VTAIL.n79 VTAIL.n67 0.155672
R627 VTAIL.n80 VTAIL.n79 0.155672
R628 VTAIL.n80 VTAIL.n63 0.155672
R629 VTAIL.n87 VTAIL.n63 0.155672
R630 VTAIL.n88 VTAIL.n87 0.155672
R631 VTAIL.n88 VTAIL.n59 0.155672
R632 VTAIL.n97 VTAIL.n59 0.155672
R633 VTAIL.n98 VTAIL.n97 0.155672
R634 VTAIL.n98 VTAIL.n55 0.155672
R635 VTAIL.n105 VTAIL.n55 0.155672
R636 VTAIL.n126 VTAIL.n121 0.155672
R637 VTAIL.n133 VTAIL.n121 0.155672
R638 VTAIL.n134 VTAIL.n133 0.155672
R639 VTAIL.n134 VTAIL.n117 0.155672
R640 VTAIL.n141 VTAIL.n117 0.155672
R641 VTAIL.n142 VTAIL.n141 0.155672
R642 VTAIL.n142 VTAIL.n113 0.155672
R643 VTAIL.n151 VTAIL.n113 0.155672
R644 VTAIL.n152 VTAIL.n151 0.155672
R645 VTAIL.n152 VTAIL.n109 0.155672
R646 VTAIL.n159 VTAIL.n109 0.155672
R647 VTAIL.n375 VTAIL.n325 0.155672
R648 VTAIL.n368 VTAIL.n325 0.155672
R649 VTAIL.n368 VTAIL.n367 0.155672
R650 VTAIL.n367 VTAIL.n329 0.155672
R651 VTAIL.n359 VTAIL.n329 0.155672
R652 VTAIL.n359 VTAIL.n358 0.155672
R653 VTAIL.n358 VTAIL.n334 0.155672
R654 VTAIL.n351 VTAIL.n334 0.155672
R655 VTAIL.n351 VTAIL.n350 0.155672
R656 VTAIL.n350 VTAIL.n338 0.155672
R657 VTAIL.n343 VTAIL.n338 0.155672
R658 VTAIL.n321 VTAIL.n271 0.155672
R659 VTAIL.n314 VTAIL.n271 0.155672
R660 VTAIL.n314 VTAIL.n313 0.155672
R661 VTAIL.n313 VTAIL.n275 0.155672
R662 VTAIL.n305 VTAIL.n275 0.155672
R663 VTAIL.n305 VTAIL.n304 0.155672
R664 VTAIL.n304 VTAIL.n280 0.155672
R665 VTAIL.n297 VTAIL.n280 0.155672
R666 VTAIL.n297 VTAIL.n296 0.155672
R667 VTAIL.n296 VTAIL.n284 0.155672
R668 VTAIL.n289 VTAIL.n284 0.155672
R669 VTAIL.n267 VTAIL.n217 0.155672
R670 VTAIL.n260 VTAIL.n217 0.155672
R671 VTAIL.n260 VTAIL.n259 0.155672
R672 VTAIL.n259 VTAIL.n221 0.155672
R673 VTAIL.n251 VTAIL.n221 0.155672
R674 VTAIL.n251 VTAIL.n250 0.155672
R675 VTAIL.n250 VTAIL.n226 0.155672
R676 VTAIL.n243 VTAIL.n226 0.155672
R677 VTAIL.n243 VTAIL.n242 0.155672
R678 VTAIL.n242 VTAIL.n230 0.155672
R679 VTAIL.n235 VTAIL.n230 0.155672
R680 VTAIL.n213 VTAIL.n163 0.155672
R681 VTAIL.n206 VTAIL.n163 0.155672
R682 VTAIL.n206 VTAIL.n205 0.155672
R683 VTAIL.n205 VTAIL.n167 0.155672
R684 VTAIL.n197 VTAIL.n167 0.155672
R685 VTAIL.n197 VTAIL.n196 0.155672
R686 VTAIL.n196 VTAIL.n172 0.155672
R687 VTAIL.n189 VTAIL.n172 0.155672
R688 VTAIL.n189 VTAIL.n188 0.155672
R689 VTAIL.n188 VTAIL.n176 0.155672
R690 VTAIL.n181 VTAIL.n176 0.155672
R691 VDD1 VDD1.n1 125.573
R692 VDD1 VDD1.n0 81.4436
R693 VDD1.n0 VDD1.t1 3.19353
R694 VDD1.n0 VDD1.t2 3.19353
R695 VDD1.n1 VDD1.t0 3.19353
R696 VDD1.n1 VDD1.t3 3.19353
R697 VN.n0 VN.t2 95.3552
R698 VN.n1 VN.t1 95.3552
R699 VN.n0 VN.t0 93.9101
R700 VN.n1 VN.t3 93.9101
R701 VN VN.n1 51.085
R702 VN VN.n0 1.72517
R703 VDD2.n2 VDD2.n0 125.049
R704 VDD2.n2 VDD2.n1 81.3855
R705 VDD2.n1 VDD2.t0 3.19353
R706 VDD2.n1 VDD2.t2 3.19353
R707 VDD2.n0 VDD2.t1 3.19353
R708 VDD2.n0 VDD2.t3 3.19353
R709 VDD2 VDD2.n2 0.0586897
R710 B.n517 B.n70 585
R711 B.n519 B.n518 585
R712 B.n520 B.n69 585
R713 B.n522 B.n521 585
R714 B.n523 B.n68 585
R715 B.n525 B.n524 585
R716 B.n526 B.n67 585
R717 B.n528 B.n527 585
R718 B.n529 B.n66 585
R719 B.n531 B.n530 585
R720 B.n532 B.n65 585
R721 B.n534 B.n533 585
R722 B.n535 B.n64 585
R723 B.n537 B.n536 585
R724 B.n538 B.n63 585
R725 B.n540 B.n539 585
R726 B.n541 B.n62 585
R727 B.n543 B.n542 585
R728 B.n544 B.n61 585
R729 B.n546 B.n545 585
R730 B.n547 B.n60 585
R731 B.n549 B.n548 585
R732 B.n550 B.n59 585
R733 B.n552 B.n551 585
R734 B.n553 B.n58 585
R735 B.n555 B.n554 585
R736 B.n556 B.n57 585
R737 B.n558 B.n557 585
R738 B.n559 B.n56 585
R739 B.n561 B.n560 585
R740 B.n562 B.n55 585
R741 B.n564 B.n563 585
R742 B.n565 B.n54 585
R743 B.n567 B.n566 585
R744 B.n568 B.n53 585
R745 B.n570 B.n569 585
R746 B.n572 B.n571 585
R747 B.n573 B.n49 585
R748 B.n575 B.n574 585
R749 B.n576 B.n48 585
R750 B.n578 B.n577 585
R751 B.n579 B.n47 585
R752 B.n581 B.n580 585
R753 B.n582 B.n46 585
R754 B.n584 B.n583 585
R755 B.n585 B.n43 585
R756 B.n588 B.n587 585
R757 B.n589 B.n42 585
R758 B.n591 B.n590 585
R759 B.n592 B.n41 585
R760 B.n594 B.n593 585
R761 B.n595 B.n40 585
R762 B.n597 B.n596 585
R763 B.n598 B.n39 585
R764 B.n600 B.n599 585
R765 B.n601 B.n38 585
R766 B.n603 B.n602 585
R767 B.n604 B.n37 585
R768 B.n606 B.n605 585
R769 B.n607 B.n36 585
R770 B.n609 B.n608 585
R771 B.n610 B.n35 585
R772 B.n612 B.n611 585
R773 B.n613 B.n34 585
R774 B.n615 B.n614 585
R775 B.n616 B.n33 585
R776 B.n618 B.n617 585
R777 B.n619 B.n32 585
R778 B.n621 B.n620 585
R779 B.n622 B.n31 585
R780 B.n624 B.n623 585
R781 B.n625 B.n30 585
R782 B.n627 B.n626 585
R783 B.n628 B.n29 585
R784 B.n630 B.n629 585
R785 B.n631 B.n28 585
R786 B.n633 B.n632 585
R787 B.n634 B.n27 585
R788 B.n636 B.n635 585
R789 B.n637 B.n26 585
R790 B.n639 B.n638 585
R791 B.n640 B.n25 585
R792 B.n516 B.n515 585
R793 B.n514 B.n71 585
R794 B.n513 B.n512 585
R795 B.n511 B.n72 585
R796 B.n510 B.n509 585
R797 B.n508 B.n73 585
R798 B.n507 B.n506 585
R799 B.n505 B.n74 585
R800 B.n504 B.n503 585
R801 B.n502 B.n75 585
R802 B.n501 B.n500 585
R803 B.n499 B.n76 585
R804 B.n498 B.n497 585
R805 B.n496 B.n77 585
R806 B.n495 B.n494 585
R807 B.n493 B.n78 585
R808 B.n492 B.n491 585
R809 B.n490 B.n79 585
R810 B.n489 B.n488 585
R811 B.n487 B.n80 585
R812 B.n486 B.n485 585
R813 B.n484 B.n81 585
R814 B.n483 B.n482 585
R815 B.n481 B.n82 585
R816 B.n480 B.n479 585
R817 B.n478 B.n83 585
R818 B.n477 B.n476 585
R819 B.n475 B.n84 585
R820 B.n474 B.n473 585
R821 B.n472 B.n85 585
R822 B.n471 B.n470 585
R823 B.n469 B.n86 585
R824 B.n468 B.n467 585
R825 B.n466 B.n87 585
R826 B.n465 B.n464 585
R827 B.n463 B.n88 585
R828 B.n462 B.n461 585
R829 B.n460 B.n89 585
R830 B.n459 B.n458 585
R831 B.n457 B.n90 585
R832 B.n456 B.n455 585
R833 B.n454 B.n91 585
R834 B.n453 B.n452 585
R835 B.n451 B.n92 585
R836 B.n450 B.n449 585
R837 B.n448 B.n93 585
R838 B.n447 B.n446 585
R839 B.n445 B.n94 585
R840 B.n444 B.n443 585
R841 B.n442 B.n95 585
R842 B.n441 B.n440 585
R843 B.n439 B.n96 585
R844 B.n438 B.n437 585
R845 B.n436 B.n97 585
R846 B.n435 B.n434 585
R847 B.n433 B.n98 585
R848 B.n432 B.n431 585
R849 B.n430 B.n99 585
R850 B.n429 B.n428 585
R851 B.n427 B.n100 585
R852 B.n426 B.n425 585
R853 B.n424 B.n101 585
R854 B.n423 B.n422 585
R855 B.n421 B.n102 585
R856 B.n420 B.n419 585
R857 B.n418 B.n103 585
R858 B.n417 B.n416 585
R859 B.n415 B.n104 585
R860 B.n414 B.n413 585
R861 B.n412 B.n105 585
R862 B.n411 B.n410 585
R863 B.n409 B.n106 585
R864 B.n408 B.n407 585
R865 B.n406 B.n107 585
R866 B.n405 B.n404 585
R867 B.n403 B.n108 585
R868 B.n402 B.n401 585
R869 B.n400 B.n109 585
R870 B.n399 B.n398 585
R871 B.n397 B.n110 585
R872 B.n396 B.n395 585
R873 B.n394 B.n111 585
R874 B.n393 B.n392 585
R875 B.n391 B.n112 585
R876 B.n390 B.n389 585
R877 B.n388 B.n113 585
R878 B.n387 B.n386 585
R879 B.n385 B.n114 585
R880 B.n384 B.n383 585
R881 B.n382 B.n115 585
R882 B.n381 B.n380 585
R883 B.n379 B.n116 585
R884 B.n378 B.n377 585
R885 B.n253 B.n162 585
R886 B.n255 B.n254 585
R887 B.n256 B.n161 585
R888 B.n258 B.n257 585
R889 B.n259 B.n160 585
R890 B.n261 B.n260 585
R891 B.n262 B.n159 585
R892 B.n264 B.n263 585
R893 B.n265 B.n158 585
R894 B.n267 B.n266 585
R895 B.n268 B.n157 585
R896 B.n270 B.n269 585
R897 B.n271 B.n156 585
R898 B.n273 B.n272 585
R899 B.n274 B.n155 585
R900 B.n276 B.n275 585
R901 B.n277 B.n154 585
R902 B.n279 B.n278 585
R903 B.n280 B.n153 585
R904 B.n282 B.n281 585
R905 B.n283 B.n152 585
R906 B.n285 B.n284 585
R907 B.n286 B.n151 585
R908 B.n288 B.n287 585
R909 B.n289 B.n150 585
R910 B.n291 B.n290 585
R911 B.n292 B.n149 585
R912 B.n294 B.n293 585
R913 B.n295 B.n148 585
R914 B.n297 B.n296 585
R915 B.n298 B.n147 585
R916 B.n300 B.n299 585
R917 B.n301 B.n146 585
R918 B.n303 B.n302 585
R919 B.n304 B.n145 585
R920 B.n306 B.n305 585
R921 B.n308 B.n307 585
R922 B.n309 B.n141 585
R923 B.n311 B.n310 585
R924 B.n312 B.n140 585
R925 B.n314 B.n313 585
R926 B.n315 B.n139 585
R927 B.n317 B.n316 585
R928 B.n318 B.n138 585
R929 B.n320 B.n319 585
R930 B.n321 B.n135 585
R931 B.n324 B.n323 585
R932 B.n325 B.n134 585
R933 B.n327 B.n326 585
R934 B.n328 B.n133 585
R935 B.n330 B.n329 585
R936 B.n331 B.n132 585
R937 B.n333 B.n332 585
R938 B.n334 B.n131 585
R939 B.n336 B.n335 585
R940 B.n337 B.n130 585
R941 B.n339 B.n338 585
R942 B.n340 B.n129 585
R943 B.n342 B.n341 585
R944 B.n343 B.n128 585
R945 B.n345 B.n344 585
R946 B.n346 B.n127 585
R947 B.n348 B.n347 585
R948 B.n349 B.n126 585
R949 B.n351 B.n350 585
R950 B.n352 B.n125 585
R951 B.n354 B.n353 585
R952 B.n355 B.n124 585
R953 B.n357 B.n356 585
R954 B.n358 B.n123 585
R955 B.n360 B.n359 585
R956 B.n361 B.n122 585
R957 B.n363 B.n362 585
R958 B.n364 B.n121 585
R959 B.n366 B.n365 585
R960 B.n367 B.n120 585
R961 B.n369 B.n368 585
R962 B.n370 B.n119 585
R963 B.n372 B.n371 585
R964 B.n373 B.n118 585
R965 B.n375 B.n374 585
R966 B.n376 B.n117 585
R967 B.n252 B.n251 585
R968 B.n250 B.n163 585
R969 B.n249 B.n248 585
R970 B.n247 B.n164 585
R971 B.n246 B.n245 585
R972 B.n244 B.n165 585
R973 B.n243 B.n242 585
R974 B.n241 B.n166 585
R975 B.n240 B.n239 585
R976 B.n238 B.n167 585
R977 B.n237 B.n236 585
R978 B.n235 B.n168 585
R979 B.n234 B.n233 585
R980 B.n232 B.n169 585
R981 B.n231 B.n230 585
R982 B.n229 B.n170 585
R983 B.n228 B.n227 585
R984 B.n226 B.n171 585
R985 B.n225 B.n224 585
R986 B.n223 B.n172 585
R987 B.n222 B.n221 585
R988 B.n220 B.n173 585
R989 B.n219 B.n218 585
R990 B.n217 B.n174 585
R991 B.n216 B.n215 585
R992 B.n214 B.n175 585
R993 B.n213 B.n212 585
R994 B.n211 B.n176 585
R995 B.n210 B.n209 585
R996 B.n208 B.n177 585
R997 B.n207 B.n206 585
R998 B.n205 B.n178 585
R999 B.n204 B.n203 585
R1000 B.n202 B.n179 585
R1001 B.n201 B.n200 585
R1002 B.n199 B.n180 585
R1003 B.n198 B.n197 585
R1004 B.n196 B.n181 585
R1005 B.n195 B.n194 585
R1006 B.n193 B.n182 585
R1007 B.n192 B.n191 585
R1008 B.n190 B.n183 585
R1009 B.n189 B.n188 585
R1010 B.n187 B.n184 585
R1011 B.n186 B.n185 585
R1012 B.n2 B.n0 585
R1013 B.n709 B.n1 585
R1014 B.n708 B.n707 585
R1015 B.n706 B.n3 585
R1016 B.n705 B.n704 585
R1017 B.n703 B.n4 585
R1018 B.n702 B.n701 585
R1019 B.n700 B.n5 585
R1020 B.n699 B.n698 585
R1021 B.n697 B.n6 585
R1022 B.n696 B.n695 585
R1023 B.n694 B.n7 585
R1024 B.n693 B.n692 585
R1025 B.n691 B.n8 585
R1026 B.n690 B.n689 585
R1027 B.n688 B.n9 585
R1028 B.n687 B.n686 585
R1029 B.n685 B.n10 585
R1030 B.n684 B.n683 585
R1031 B.n682 B.n11 585
R1032 B.n681 B.n680 585
R1033 B.n679 B.n12 585
R1034 B.n678 B.n677 585
R1035 B.n676 B.n13 585
R1036 B.n675 B.n674 585
R1037 B.n673 B.n14 585
R1038 B.n672 B.n671 585
R1039 B.n670 B.n15 585
R1040 B.n669 B.n668 585
R1041 B.n667 B.n16 585
R1042 B.n666 B.n665 585
R1043 B.n664 B.n17 585
R1044 B.n663 B.n662 585
R1045 B.n661 B.n18 585
R1046 B.n660 B.n659 585
R1047 B.n658 B.n19 585
R1048 B.n657 B.n656 585
R1049 B.n655 B.n20 585
R1050 B.n654 B.n653 585
R1051 B.n652 B.n21 585
R1052 B.n651 B.n650 585
R1053 B.n649 B.n22 585
R1054 B.n648 B.n647 585
R1055 B.n646 B.n23 585
R1056 B.n645 B.n644 585
R1057 B.n643 B.n24 585
R1058 B.n642 B.n641 585
R1059 B.n711 B.n710 585
R1060 B.n253 B.n252 545.355
R1061 B.n642 B.n25 545.355
R1062 B.n378 B.n117 545.355
R1063 B.n517 B.n516 545.355
R1064 B.n136 B.t11 426.849
R1065 B.n50 B.t4 426.849
R1066 B.n142 B.t2 426.849
R1067 B.n44 B.t7 426.849
R1068 B.n137 B.t10 343.067
R1069 B.n51 B.t5 343.067
R1070 B.n143 B.t1 343.067
R1071 B.n45 B.t8 343.067
R1072 B.n136 B.t9 270.973
R1073 B.n142 B.t0 270.973
R1074 B.n44 B.t6 270.973
R1075 B.n50 B.t3 270.973
R1076 B.n252 B.n163 163.367
R1077 B.n248 B.n163 163.367
R1078 B.n248 B.n247 163.367
R1079 B.n247 B.n246 163.367
R1080 B.n246 B.n165 163.367
R1081 B.n242 B.n165 163.367
R1082 B.n242 B.n241 163.367
R1083 B.n241 B.n240 163.367
R1084 B.n240 B.n167 163.367
R1085 B.n236 B.n167 163.367
R1086 B.n236 B.n235 163.367
R1087 B.n235 B.n234 163.367
R1088 B.n234 B.n169 163.367
R1089 B.n230 B.n169 163.367
R1090 B.n230 B.n229 163.367
R1091 B.n229 B.n228 163.367
R1092 B.n228 B.n171 163.367
R1093 B.n224 B.n171 163.367
R1094 B.n224 B.n223 163.367
R1095 B.n223 B.n222 163.367
R1096 B.n222 B.n173 163.367
R1097 B.n218 B.n173 163.367
R1098 B.n218 B.n217 163.367
R1099 B.n217 B.n216 163.367
R1100 B.n216 B.n175 163.367
R1101 B.n212 B.n175 163.367
R1102 B.n212 B.n211 163.367
R1103 B.n211 B.n210 163.367
R1104 B.n210 B.n177 163.367
R1105 B.n206 B.n177 163.367
R1106 B.n206 B.n205 163.367
R1107 B.n205 B.n204 163.367
R1108 B.n204 B.n179 163.367
R1109 B.n200 B.n179 163.367
R1110 B.n200 B.n199 163.367
R1111 B.n199 B.n198 163.367
R1112 B.n198 B.n181 163.367
R1113 B.n194 B.n181 163.367
R1114 B.n194 B.n193 163.367
R1115 B.n193 B.n192 163.367
R1116 B.n192 B.n183 163.367
R1117 B.n188 B.n183 163.367
R1118 B.n188 B.n187 163.367
R1119 B.n187 B.n186 163.367
R1120 B.n186 B.n2 163.367
R1121 B.n710 B.n2 163.367
R1122 B.n710 B.n709 163.367
R1123 B.n709 B.n708 163.367
R1124 B.n708 B.n3 163.367
R1125 B.n704 B.n3 163.367
R1126 B.n704 B.n703 163.367
R1127 B.n703 B.n702 163.367
R1128 B.n702 B.n5 163.367
R1129 B.n698 B.n5 163.367
R1130 B.n698 B.n697 163.367
R1131 B.n697 B.n696 163.367
R1132 B.n696 B.n7 163.367
R1133 B.n692 B.n7 163.367
R1134 B.n692 B.n691 163.367
R1135 B.n691 B.n690 163.367
R1136 B.n690 B.n9 163.367
R1137 B.n686 B.n9 163.367
R1138 B.n686 B.n685 163.367
R1139 B.n685 B.n684 163.367
R1140 B.n684 B.n11 163.367
R1141 B.n680 B.n11 163.367
R1142 B.n680 B.n679 163.367
R1143 B.n679 B.n678 163.367
R1144 B.n678 B.n13 163.367
R1145 B.n674 B.n13 163.367
R1146 B.n674 B.n673 163.367
R1147 B.n673 B.n672 163.367
R1148 B.n672 B.n15 163.367
R1149 B.n668 B.n15 163.367
R1150 B.n668 B.n667 163.367
R1151 B.n667 B.n666 163.367
R1152 B.n666 B.n17 163.367
R1153 B.n662 B.n17 163.367
R1154 B.n662 B.n661 163.367
R1155 B.n661 B.n660 163.367
R1156 B.n660 B.n19 163.367
R1157 B.n656 B.n19 163.367
R1158 B.n656 B.n655 163.367
R1159 B.n655 B.n654 163.367
R1160 B.n654 B.n21 163.367
R1161 B.n650 B.n21 163.367
R1162 B.n650 B.n649 163.367
R1163 B.n649 B.n648 163.367
R1164 B.n648 B.n23 163.367
R1165 B.n644 B.n23 163.367
R1166 B.n644 B.n643 163.367
R1167 B.n643 B.n642 163.367
R1168 B.n254 B.n253 163.367
R1169 B.n254 B.n161 163.367
R1170 B.n258 B.n161 163.367
R1171 B.n259 B.n258 163.367
R1172 B.n260 B.n259 163.367
R1173 B.n260 B.n159 163.367
R1174 B.n264 B.n159 163.367
R1175 B.n265 B.n264 163.367
R1176 B.n266 B.n265 163.367
R1177 B.n266 B.n157 163.367
R1178 B.n270 B.n157 163.367
R1179 B.n271 B.n270 163.367
R1180 B.n272 B.n271 163.367
R1181 B.n272 B.n155 163.367
R1182 B.n276 B.n155 163.367
R1183 B.n277 B.n276 163.367
R1184 B.n278 B.n277 163.367
R1185 B.n278 B.n153 163.367
R1186 B.n282 B.n153 163.367
R1187 B.n283 B.n282 163.367
R1188 B.n284 B.n283 163.367
R1189 B.n284 B.n151 163.367
R1190 B.n288 B.n151 163.367
R1191 B.n289 B.n288 163.367
R1192 B.n290 B.n289 163.367
R1193 B.n290 B.n149 163.367
R1194 B.n294 B.n149 163.367
R1195 B.n295 B.n294 163.367
R1196 B.n296 B.n295 163.367
R1197 B.n296 B.n147 163.367
R1198 B.n300 B.n147 163.367
R1199 B.n301 B.n300 163.367
R1200 B.n302 B.n301 163.367
R1201 B.n302 B.n145 163.367
R1202 B.n306 B.n145 163.367
R1203 B.n307 B.n306 163.367
R1204 B.n307 B.n141 163.367
R1205 B.n311 B.n141 163.367
R1206 B.n312 B.n311 163.367
R1207 B.n313 B.n312 163.367
R1208 B.n313 B.n139 163.367
R1209 B.n317 B.n139 163.367
R1210 B.n318 B.n317 163.367
R1211 B.n319 B.n318 163.367
R1212 B.n319 B.n135 163.367
R1213 B.n324 B.n135 163.367
R1214 B.n325 B.n324 163.367
R1215 B.n326 B.n325 163.367
R1216 B.n326 B.n133 163.367
R1217 B.n330 B.n133 163.367
R1218 B.n331 B.n330 163.367
R1219 B.n332 B.n331 163.367
R1220 B.n332 B.n131 163.367
R1221 B.n336 B.n131 163.367
R1222 B.n337 B.n336 163.367
R1223 B.n338 B.n337 163.367
R1224 B.n338 B.n129 163.367
R1225 B.n342 B.n129 163.367
R1226 B.n343 B.n342 163.367
R1227 B.n344 B.n343 163.367
R1228 B.n344 B.n127 163.367
R1229 B.n348 B.n127 163.367
R1230 B.n349 B.n348 163.367
R1231 B.n350 B.n349 163.367
R1232 B.n350 B.n125 163.367
R1233 B.n354 B.n125 163.367
R1234 B.n355 B.n354 163.367
R1235 B.n356 B.n355 163.367
R1236 B.n356 B.n123 163.367
R1237 B.n360 B.n123 163.367
R1238 B.n361 B.n360 163.367
R1239 B.n362 B.n361 163.367
R1240 B.n362 B.n121 163.367
R1241 B.n366 B.n121 163.367
R1242 B.n367 B.n366 163.367
R1243 B.n368 B.n367 163.367
R1244 B.n368 B.n119 163.367
R1245 B.n372 B.n119 163.367
R1246 B.n373 B.n372 163.367
R1247 B.n374 B.n373 163.367
R1248 B.n374 B.n117 163.367
R1249 B.n379 B.n378 163.367
R1250 B.n380 B.n379 163.367
R1251 B.n380 B.n115 163.367
R1252 B.n384 B.n115 163.367
R1253 B.n385 B.n384 163.367
R1254 B.n386 B.n385 163.367
R1255 B.n386 B.n113 163.367
R1256 B.n390 B.n113 163.367
R1257 B.n391 B.n390 163.367
R1258 B.n392 B.n391 163.367
R1259 B.n392 B.n111 163.367
R1260 B.n396 B.n111 163.367
R1261 B.n397 B.n396 163.367
R1262 B.n398 B.n397 163.367
R1263 B.n398 B.n109 163.367
R1264 B.n402 B.n109 163.367
R1265 B.n403 B.n402 163.367
R1266 B.n404 B.n403 163.367
R1267 B.n404 B.n107 163.367
R1268 B.n408 B.n107 163.367
R1269 B.n409 B.n408 163.367
R1270 B.n410 B.n409 163.367
R1271 B.n410 B.n105 163.367
R1272 B.n414 B.n105 163.367
R1273 B.n415 B.n414 163.367
R1274 B.n416 B.n415 163.367
R1275 B.n416 B.n103 163.367
R1276 B.n420 B.n103 163.367
R1277 B.n421 B.n420 163.367
R1278 B.n422 B.n421 163.367
R1279 B.n422 B.n101 163.367
R1280 B.n426 B.n101 163.367
R1281 B.n427 B.n426 163.367
R1282 B.n428 B.n427 163.367
R1283 B.n428 B.n99 163.367
R1284 B.n432 B.n99 163.367
R1285 B.n433 B.n432 163.367
R1286 B.n434 B.n433 163.367
R1287 B.n434 B.n97 163.367
R1288 B.n438 B.n97 163.367
R1289 B.n439 B.n438 163.367
R1290 B.n440 B.n439 163.367
R1291 B.n440 B.n95 163.367
R1292 B.n444 B.n95 163.367
R1293 B.n445 B.n444 163.367
R1294 B.n446 B.n445 163.367
R1295 B.n446 B.n93 163.367
R1296 B.n450 B.n93 163.367
R1297 B.n451 B.n450 163.367
R1298 B.n452 B.n451 163.367
R1299 B.n452 B.n91 163.367
R1300 B.n456 B.n91 163.367
R1301 B.n457 B.n456 163.367
R1302 B.n458 B.n457 163.367
R1303 B.n458 B.n89 163.367
R1304 B.n462 B.n89 163.367
R1305 B.n463 B.n462 163.367
R1306 B.n464 B.n463 163.367
R1307 B.n464 B.n87 163.367
R1308 B.n468 B.n87 163.367
R1309 B.n469 B.n468 163.367
R1310 B.n470 B.n469 163.367
R1311 B.n470 B.n85 163.367
R1312 B.n474 B.n85 163.367
R1313 B.n475 B.n474 163.367
R1314 B.n476 B.n475 163.367
R1315 B.n476 B.n83 163.367
R1316 B.n480 B.n83 163.367
R1317 B.n481 B.n480 163.367
R1318 B.n482 B.n481 163.367
R1319 B.n482 B.n81 163.367
R1320 B.n486 B.n81 163.367
R1321 B.n487 B.n486 163.367
R1322 B.n488 B.n487 163.367
R1323 B.n488 B.n79 163.367
R1324 B.n492 B.n79 163.367
R1325 B.n493 B.n492 163.367
R1326 B.n494 B.n493 163.367
R1327 B.n494 B.n77 163.367
R1328 B.n498 B.n77 163.367
R1329 B.n499 B.n498 163.367
R1330 B.n500 B.n499 163.367
R1331 B.n500 B.n75 163.367
R1332 B.n504 B.n75 163.367
R1333 B.n505 B.n504 163.367
R1334 B.n506 B.n505 163.367
R1335 B.n506 B.n73 163.367
R1336 B.n510 B.n73 163.367
R1337 B.n511 B.n510 163.367
R1338 B.n512 B.n511 163.367
R1339 B.n512 B.n71 163.367
R1340 B.n516 B.n71 163.367
R1341 B.n638 B.n25 163.367
R1342 B.n638 B.n637 163.367
R1343 B.n637 B.n636 163.367
R1344 B.n636 B.n27 163.367
R1345 B.n632 B.n27 163.367
R1346 B.n632 B.n631 163.367
R1347 B.n631 B.n630 163.367
R1348 B.n630 B.n29 163.367
R1349 B.n626 B.n29 163.367
R1350 B.n626 B.n625 163.367
R1351 B.n625 B.n624 163.367
R1352 B.n624 B.n31 163.367
R1353 B.n620 B.n31 163.367
R1354 B.n620 B.n619 163.367
R1355 B.n619 B.n618 163.367
R1356 B.n618 B.n33 163.367
R1357 B.n614 B.n33 163.367
R1358 B.n614 B.n613 163.367
R1359 B.n613 B.n612 163.367
R1360 B.n612 B.n35 163.367
R1361 B.n608 B.n35 163.367
R1362 B.n608 B.n607 163.367
R1363 B.n607 B.n606 163.367
R1364 B.n606 B.n37 163.367
R1365 B.n602 B.n37 163.367
R1366 B.n602 B.n601 163.367
R1367 B.n601 B.n600 163.367
R1368 B.n600 B.n39 163.367
R1369 B.n596 B.n39 163.367
R1370 B.n596 B.n595 163.367
R1371 B.n595 B.n594 163.367
R1372 B.n594 B.n41 163.367
R1373 B.n590 B.n41 163.367
R1374 B.n590 B.n589 163.367
R1375 B.n589 B.n588 163.367
R1376 B.n588 B.n43 163.367
R1377 B.n583 B.n43 163.367
R1378 B.n583 B.n582 163.367
R1379 B.n582 B.n581 163.367
R1380 B.n581 B.n47 163.367
R1381 B.n577 B.n47 163.367
R1382 B.n577 B.n576 163.367
R1383 B.n576 B.n575 163.367
R1384 B.n575 B.n49 163.367
R1385 B.n571 B.n49 163.367
R1386 B.n571 B.n570 163.367
R1387 B.n570 B.n53 163.367
R1388 B.n566 B.n53 163.367
R1389 B.n566 B.n565 163.367
R1390 B.n565 B.n564 163.367
R1391 B.n564 B.n55 163.367
R1392 B.n560 B.n55 163.367
R1393 B.n560 B.n559 163.367
R1394 B.n559 B.n558 163.367
R1395 B.n558 B.n57 163.367
R1396 B.n554 B.n57 163.367
R1397 B.n554 B.n553 163.367
R1398 B.n553 B.n552 163.367
R1399 B.n552 B.n59 163.367
R1400 B.n548 B.n59 163.367
R1401 B.n548 B.n547 163.367
R1402 B.n547 B.n546 163.367
R1403 B.n546 B.n61 163.367
R1404 B.n542 B.n61 163.367
R1405 B.n542 B.n541 163.367
R1406 B.n541 B.n540 163.367
R1407 B.n540 B.n63 163.367
R1408 B.n536 B.n63 163.367
R1409 B.n536 B.n535 163.367
R1410 B.n535 B.n534 163.367
R1411 B.n534 B.n65 163.367
R1412 B.n530 B.n65 163.367
R1413 B.n530 B.n529 163.367
R1414 B.n529 B.n528 163.367
R1415 B.n528 B.n67 163.367
R1416 B.n524 B.n67 163.367
R1417 B.n524 B.n523 163.367
R1418 B.n523 B.n522 163.367
R1419 B.n522 B.n69 163.367
R1420 B.n518 B.n69 163.367
R1421 B.n518 B.n517 163.367
R1422 B.n137 B.n136 83.7823
R1423 B.n143 B.n142 83.7823
R1424 B.n45 B.n44 83.7823
R1425 B.n51 B.n50 83.7823
R1426 B.n322 B.n137 59.5399
R1427 B.n144 B.n143 59.5399
R1428 B.n586 B.n45 59.5399
R1429 B.n52 B.n51 59.5399
R1430 B.n515 B.n70 35.4346
R1431 B.n641 B.n640 35.4346
R1432 B.n377 B.n376 35.4346
R1433 B.n251 B.n162 35.4346
R1434 B B.n711 18.0485
R1435 B.n640 B.n639 10.6151
R1436 B.n639 B.n26 10.6151
R1437 B.n635 B.n26 10.6151
R1438 B.n635 B.n634 10.6151
R1439 B.n634 B.n633 10.6151
R1440 B.n633 B.n28 10.6151
R1441 B.n629 B.n28 10.6151
R1442 B.n629 B.n628 10.6151
R1443 B.n628 B.n627 10.6151
R1444 B.n627 B.n30 10.6151
R1445 B.n623 B.n30 10.6151
R1446 B.n623 B.n622 10.6151
R1447 B.n622 B.n621 10.6151
R1448 B.n621 B.n32 10.6151
R1449 B.n617 B.n32 10.6151
R1450 B.n617 B.n616 10.6151
R1451 B.n616 B.n615 10.6151
R1452 B.n615 B.n34 10.6151
R1453 B.n611 B.n34 10.6151
R1454 B.n611 B.n610 10.6151
R1455 B.n610 B.n609 10.6151
R1456 B.n609 B.n36 10.6151
R1457 B.n605 B.n36 10.6151
R1458 B.n605 B.n604 10.6151
R1459 B.n604 B.n603 10.6151
R1460 B.n603 B.n38 10.6151
R1461 B.n599 B.n38 10.6151
R1462 B.n599 B.n598 10.6151
R1463 B.n598 B.n597 10.6151
R1464 B.n597 B.n40 10.6151
R1465 B.n593 B.n40 10.6151
R1466 B.n593 B.n592 10.6151
R1467 B.n592 B.n591 10.6151
R1468 B.n591 B.n42 10.6151
R1469 B.n587 B.n42 10.6151
R1470 B.n585 B.n584 10.6151
R1471 B.n584 B.n46 10.6151
R1472 B.n580 B.n46 10.6151
R1473 B.n580 B.n579 10.6151
R1474 B.n579 B.n578 10.6151
R1475 B.n578 B.n48 10.6151
R1476 B.n574 B.n48 10.6151
R1477 B.n574 B.n573 10.6151
R1478 B.n573 B.n572 10.6151
R1479 B.n569 B.n568 10.6151
R1480 B.n568 B.n567 10.6151
R1481 B.n567 B.n54 10.6151
R1482 B.n563 B.n54 10.6151
R1483 B.n563 B.n562 10.6151
R1484 B.n562 B.n561 10.6151
R1485 B.n561 B.n56 10.6151
R1486 B.n557 B.n56 10.6151
R1487 B.n557 B.n556 10.6151
R1488 B.n556 B.n555 10.6151
R1489 B.n555 B.n58 10.6151
R1490 B.n551 B.n58 10.6151
R1491 B.n551 B.n550 10.6151
R1492 B.n550 B.n549 10.6151
R1493 B.n549 B.n60 10.6151
R1494 B.n545 B.n60 10.6151
R1495 B.n545 B.n544 10.6151
R1496 B.n544 B.n543 10.6151
R1497 B.n543 B.n62 10.6151
R1498 B.n539 B.n62 10.6151
R1499 B.n539 B.n538 10.6151
R1500 B.n538 B.n537 10.6151
R1501 B.n537 B.n64 10.6151
R1502 B.n533 B.n64 10.6151
R1503 B.n533 B.n532 10.6151
R1504 B.n532 B.n531 10.6151
R1505 B.n531 B.n66 10.6151
R1506 B.n527 B.n66 10.6151
R1507 B.n527 B.n526 10.6151
R1508 B.n526 B.n525 10.6151
R1509 B.n525 B.n68 10.6151
R1510 B.n521 B.n68 10.6151
R1511 B.n521 B.n520 10.6151
R1512 B.n520 B.n519 10.6151
R1513 B.n519 B.n70 10.6151
R1514 B.n377 B.n116 10.6151
R1515 B.n381 B.n116 10.6151
R1516 B.n382 B.n381 10.6151
R1517 B.n383 B.n382 10.6151
R1518 B.n383 B.n114 10.6151
R1519 B.n387 B.n114 10.6151
R1520 B.n388 B.n387 10.6151
R1521 B.n389 B.n388 10.6151
R1522 B.n389 B.n112 10.6151
R1523 B.n393 B.n112 10.6151
R1524 B.n394 B.n393 10.6151
R1525 B.n395 B.n394 10.6151
R1526 B.n395 B.n110 10.6151
R1527 B.n399 B.n110 10.6151
R1528 B.n400 B.n399 10.6151
R1529 B.n401 B.n400 10.6151
R1530 B.n401 B.n108 10.6151
R1531 B.n405 B.n108 10.6151
R1532 B.n406 B.n405 10.6151
R1533 B.n407 B.n406 10.6151
R1534 B.n407 B.n106 10.6151
R1535 B.n411 B.n106 10.6151
R1536 B.n412 B.n411 10.6151
R1537 B.n413 B.n412 10.6151
R1538 B.n413 B.n104 10.6151
R1539 B.n417 B.n104 10.6151
R1540 B.n418 B.n417 10.6151
R1541 B.n419 B.n418 10.6151
R1542 B.n419 B.n102 10.6151
R1543 B.n423 B.n102 10.6151
R1544 B.n424 B.n423 10.6151
R1545 B.n425 B.n424 10.6151
R1546 B.n425 B.n100 10.6151
R1547 B.n429 B.n100 10.6151
R1548 B.n430 B.n429 10.6151
R1549 B.n431 B.n430 10.6151
R1550 B.n431 B.n98 10.6151
R1551 B.n435 B.n98 10.6151
R1552 B.n436 B.n435 10.6151
R1553 B.n437 B.n436 10.6151
R1554 B.n437 B.n96 10.6151
R1555 B.n441 B.n96 10.6151
R1556 B.n442 B.n441 10.6151
R1557 B.n443 B.n442 10.6151
R1558 B.n443 B.n94 10.6151
R1559 B.n447 B.n94 10.6151
R1560 B.n448 B.n447 10.6151
R1561 B.n449 B.n448 10.6151
R1562 B.n449 B.n92 10.6151
R1563 B.n453 B.n92 10.6151
R1564 B.n454 B.n453 10.6151
R1565 B.n455 B.n454 10.6151
R1566 B.n455 B.n90 10.6151
R1567 B.n459 B.n90 10.6151
R1568 B.n460 B.n459 10.6151
R1569 B.n461 B.n460 10.6151
R1570 B.n461 B.n88 10.6151
R1571 B.n465 B.n88 10.6151
R1572 B.n466 B.n465 10.6151
R1573 B.n467 B.n466 10.6151
R1574 B.n467 B.n86 10.6151
R1575 B.n471 B.n86 10.6151
R1576 B.n472 B.n471 10.6151
R1577 B.n473 B.n472 10.6151
R1578 B.n473 B.n84 10.6151
R1579 B.n477 B.n84 10.6151
R1580 B.n478 B.n477 10.6151
R1581 B.n479 B.n478 10.6151
R1582 B.n479 B.n82 10.6151
R1583 B.n483 B.n82 10.6151
R1584 B.n484 B.n483 10.6151
R1585 B.n485 B.n484 10.6151
R1586 B.n485 B.n80 10.6151
R1587 B.n489 B.n80 10.6151
R1588 B.n490 B.n489 10.6151
R1589 B.n491 B.n490 10.6151
R1590 B.n491 B.n78 10.6151
R1591 B.n495 B.n78 10.6151
R1592 B.n496 B.n495 10.6151
R1593 B.n497 B.n496 10.6151
R1594 B.n497 B.n76 10.6151
R1595 B.n501 B.n76 10.6151
R1596 B.n502 B.n501 10.6151
R1597 B.n503 B.n502 10.6151
R1598 B.n503 B.n74 10.6151
R1599 B.n507 B.n74 10.6151
R1600 B.n508 B.n507 10.6151
R1601 B.n509 B.n508 10.6151
R1602 B.n509 B.n72 10.6151
R1603 B.n513 B.n72 10.6151
R1604 B.n514 B.n513 10.6151
R1605 B.n515 B.n514 10.6151
R1606 B.n255 B.n162 10.6151
R1607 B.n256 B.n255 10.6151
R1608 B.n257 B.n256 10.6151
R1609 B.n257 B.n160 10.6151
R1610 B.n261 B.n160 10.6151
R1611 B.n262 B.n261 10.6151
R1612 B.n263 B.n262 10.6151
R1613 B.n263 B.n158 10.6151
R1614 B.n267 B.n158 10.6151
R1615 B.n268 B.n267 10.6151
R1616 B.n269 B.n268 10.6151
R1617 B.n269 B.n156 10.6151
R1618 B.n273 B.n156 10.6151
R1619 B.n274 B.n273 10.6151
R1620 B.n275 B.n274 10.6151
R1621 B.n275 B.n154 10.6151
R1622 B.n279 B.n154 10.6151
R1623 B.n280 B.n279 10.6151
R1624 B.n281 B.n280 10.6151
R1625 B.n281 B.n152 10.6151
R1626 B.n285 B.n152 10.6151
R1627 B.n286 B.n285 10.6151
R1628 B.n287 B.n286 10.6151
R1629 B.n287 B.n150 10.6151
R1630 B.n291 B.n150 10.6151
R1631 B.n292 B.n291 10.6151
R1632 B.n293 B.n292 10.6151
R1633 B.n293 B.n148 10.6151
R1634 B.n297 B.n148 10.6151
R1635 B.n298 B.n297 10.6151
R1636 B.n299 B.n298 10.6151
R1637 B.n299 B.n146 10.6151
R1638 B.n303 B.n146 10.6151
R1639 B.n304 B.n303 10.6151
R1640 B.n305 B.n304 10.6151
R1641 B.n309 B.n308 10.6151
R1642 B.n310 B.n309 10.6151
R1643 B.n310 B.n140 10.6151
R1644 B.n314 B.n140 10.6151
R1645 B.n315 B.n314 10.6151
R1646 B.n316 B.n315 10.6151
R1647 B.n316 B.n138 10.6151
R1648 B.n320 B.n138 10.6151
R1649 B.n321 B.n320 10.6151
R1650 B.n323 B.n134 10.6151
R1651 B.n327 B.n134 10.6151
R1652 B.n328 B.n327 10.6151
R1653 B.n329 B.n328 10.6151
R1654 B.n329 B.n132 10.6151
R1655 B.n333 B.n132 10.6151
R1656 B.n334 B.n333 10.6151
R1657 B.n335 B.n334 10.6151
R1658 B.n335 B.n130 10.6151
R1659 B.n339 B.n130 10.6151
R1660 B.n340 B.n339 10.6151
R1661 B.n341 B.n340 10.6151
R1662 B.n341 B.n128 10.6151
R1663 B.n345 B.n128 10.6151
R1664 B.n346 B.n345 10.6151
R1665 B.n347 B.n346 10.6151
R1666 B.n347 B.n126 10.6151
R1667 B.n351 B.n126 10.6151
R1668 B.n352 B.n351 10.6151
R1669 B.n353 B.n352 10.6151
R1670 B.n353 B.n124 10.6151
R1671 B.n357 B.n124 10.6151
R1672 B.n358 B.n357 10.6151
R1673 B.n359 B.n358 10.6151
R1674 B.n359 B.n122 10.6151
R1675 B.n363 B.n122 10.6151
R1676 B.n364 B.n363 10.6151
R1677 B.n365 B.n364 10.6151
R1678 B.n365 B.n120 10.6151
R1679 B.n369 B.n120 10.6151
R1680 B.n370 B.n369 10.6151
R1681 B.n371 B.n370 10.6151
R1682 B.n371 B.n118 10.6151
R1683 B.n375 B.n118 10.6151
R1684 B.n376 B.n375 10.6151
R1685 B.n251 B.n250 10.6151
R1686 B.n250 B.n249 10.6151
R1687 B.n249 B.n164 10.6151
R1688 B.n245 B.n164 10.6151
R1689 B.n245 B.n244 10.6151
R1690 B.n244 B.n243 10.6151
R1691 B.n243 B.n166 10.6151
R1692 B.n239 B.n166 10.6151
R1693 B.n239 B.n238 10.6151
R1694 B.n238 B.n237 10.6151
R1695 B.n237 B.n168 10.6151
R1696 B.n233 B.n168 10.6151
R1697 B.n233 B.n232 10.6151
R1698 B.n232 B.n231 10.6151
R1699 B.n231 B.n170 10.6151
R1700 B.n227 B.n170 10.6151
R1701 B.n227 B.n226 10.6151
R1702 B.n226 B.n225 10.6151
R1703 B.n225 B.n172 10.6151
R1704 B.n221 B.n172 10.6151
R1705 B.n221 B.n220 10.6151
R1706 B.n220 B.n219 10.6151
R1707 B.n219 B.n174 10.6151
R1708 B.n215 B.n174 10.6151
R1709 B.n215 B.n214 10.6151
R1710 B.n214 B.n213 10.6151
R1711 B.n213 B.n176 10.6151
R1712 B.n209 B.n176 10.6151
R1713 B.n209 B.n208 10.6151
R1714 B.n208 B.n207 10.6151
R1715 B.n207 B.n178 10.6151
R1716 B.n203 B.n178 10.6151
R1717 B.n203 B.n202 10.6151
R1718 B.n202 B.n201 10.6151
R1719 B.n201 B.n180 10.6151
R1720 B.n197 B.n180 10.6151
R1721 B.n197 B.n196 10.6151
R1722 B.n196 B.n195 10.6151
R1723 B.n195 B.n182 10.6151
R1724 B.n191 B.n182 10.6151
R1725 B.n191 B.n190 10.6151
R1726 B.n190 B.n189 10.6151
R1727 B.n189 B.n184 10.6151
R1728 B.n185 B.n184 10.6151
R1729 B.n185 B.n0 10.6151
R1730 B.n707 B.n1 10.6151
R1731 B.n707 B.n706 10.6151
R1732 B.n706 B.n705 10.6151
R1733 B.n705 B.n4 10.6151
R1734 B.n701 B.n4 10.6151
R1735 B.n701 B.n700 10.6151
R1736 B.n700 B.n699 10.6151
R1737 B.n699 B.n6 10.6151
R1738 B.n695 B.n6 10.6151
R1739 B.n695 B.n694 10.6151
R1740 B.n694 B.n693 10.6151
R1741 B.n693 B.n8 10.6151
R1742 B.n689 B.n8 10.6151
R1743 B.n689 B.n688 10.6151
R1744 B.n688 B.n687 10.6151
R1745 B.n687 B.n10 10.6151
R1746 B.n683 B.n10 10.6151
R1747 B.n683 B.n682 10.6151
R1748 B.n682 B.n681 10.6151
R1749 B.n681 B.n12 10.6151
R1750 B.n677 B.n12 10.6151
R1751 B.n677 B.n676 10.6151
R1752 B.n676 B.n675 10.6151
R1753 B.n675 B.n14 10.6151
R1754 B.n671 B.n14 10.6151
R1755 B.n671 B.n670 10.6151
R1756 B.n670 B.n669 10.6151
R1757 B.n669 B.n16 10.6151
R1758 B.n665 B.n16 10.6151
R1759 B.n665 B.n664 10.6151
R1760 B.n664 B.n663 10.6151
R1761 B.n663 B.n18 10.6151
R1762 B.n659 B.n18 10.6151
R1763 B.n659 B.n658 10.6151
R1764 B.n658 B.n657 10.6151
R1765 B.n657 B.n20 10.6151
R1766 B.n653 B.n20 10.6151
R1767 B.n653 B.n652 10.6151
R1768 B.n652 B.n651 10.6151
R1769 B.n651 B.n22 10.6151
R1770 B.n647 B.n22 10.6151
R1771 B.n647 B.n646 10.6151
R1772 B.n646 B.n645 10.6151
R1773 B.n645 B.n24 10.6151
R1774 B.n641 B.n24 10.6151
R1775 B.n587 B.n586 9.36635
R1776 B.n569 B.n52 9.36635
R1777 B.n305 B.n144 9.36635
R1778 B.n323 B.n322 9.36635
R1779 B.n711 B.n0 2.81026
R1780 B.n711 B.n1 2.81026
R1781 B.n586 B.n585 1.24928
R1782 B.n572 B.n52 1.24928
R1783 B.n308 B.n144 1.24928
R1784 B.n322 B.n321 1.24928
C0 w_n3562_n3004# VP 6.71281f
C1 VP VDD1 4.67339f
C2 w_n3562_n3004# VN 6.25139f
C3 VN VDD1 0.150749f
C4 VP VDD2 0.483246f
C5 VN VDD2 4.34198f
C6 B VP 2.12806f
C7 B VN 1.35588f
C8 VP VTAIL 4.56469f
C9 VN VTAIL 4.55058f
C10 w_n3562_n3004# VDD1 1.66554f
C11 w_n3562_n3004# VDD2 1.75228f
C12 VDD2 VDD1 1.36932f
C13 B w_n3562_n3004# 10.445f
C14 B VDD1 1.45929f
C15 B VDD2 1.53443f
C16 VN VP 6.85311f
C17 w_n3562_n3004# VTAIL 3.62501f
C18 VDD1 VTAIL 5.44815f
C19 VDD2 VTAIL 5.51168f
C20 B VTAIL 4.86006f
C21 VDD2 VSUBS 1.124157f
C22 VDD1 VSUBS 6.335889f
C23 VTAIL VSUBS 1.329561f
C24 VN VSUBS 6.24546f
C25 VP VSUBS 2.979949f
C26 B VSUBS 5.318808f
C27 w_n3562_n3004# VSUBS 0.132122p
C28 B.n0 VSUBS 0.00463f
C29 B.n1 VSUBS 0.00463f
C30 B.n2 VSUBS 0.007322f
C31 B.n3 VSUBS 0.007322f
C32 B.n4 VSUBS 0.007322f
C33 B.n5 VSUBS 0.007322f
C34 B.n6 VSUBS 0.007322f
C35 B.n7 VSUBS 0.007322f
C36 B.n8 VSUBS 0.007322f
C37 B.n9 VSUBS 0.007322f
C38 B.n10 VSUBS 0.007322f
C39 B.n11 VSUBS 0.007322f
C40 B.n12 VSUBS 0.007322f
C41 B.n13 VSUBS 0.007322f
C42 B.n14 VSUBS 0.007322f
C43 B.n15 VSUBS 0.007322f
C44 B.n16 VSUBS 0.007322f
C45 B.n17 VSUBS 0.007322f
C46 B.n18 VSUBS 0.007322f
C47 B.n19 VSUBS 0.007322f
C48 B.n20 VSUBS 0.007322f
C49 B.n21 VSUBS 0.007322f
C50 B.n22 VSUBS 0.007322f
C51 B.n23 VSUBS 0.007322f
C52 B.n24 VSUBS 0.007322f
C53 B.n25 VSUBS 0.018586f
C54 B.n26 VSUBS 0.007322f
C55 B.n27 VSUBS 0.007322f
C56 B.n28 VSUBS 0.007322f
C57 B.n29 VSUBS 0.007322f
C58 B.n30 VSUBS 0.007322f
C59 B.n31 VSUBS 0.007322f
C60 B.n32 VSUBS 0.007322f
C61 B.n33 VSUBS 0.007322f
C62 B.n34 VSUBS 0.007322f
C63 B.n35 VSUBS 0.007322f
C64 B.n36 VSUBS 0.007322f
C65 B.n37 VSUBS 0.007322f
C66 B.n38 VSUBS 0.007322f
C67 B.n39 VSUBS 0.007322f
C68 B.n40 VSUBS 0.007322f
C69 B.n41 VSUBS 0.007322f
C70 B.n42 VSUBS 0.007322f
C71 B.n43 VSUBS 0.007322f
C72 B.t8 VSUBS 0.179509f
C73 B.t7 VSUBS 0.224929f
C74 B.t6 VSUBS 2.00302f
C75 B.n44 VSUBS 0.359657f
C76 B.n45 VSUBS 0.241847f
C77 B.n46 VSUBS 0.007322f
C78 B.n47 VSUBS 0.007322f
C79 B.n48 VSUBS 0.007322f
C80 B.n49 VSUBS 0.007322f
C81 B.t5 VSUBS 0.179512f
C82 B.t4 VSUBS 0.224931f
C83 B.t3 VSUBS 2.00302f
C84 B.n50 VSUBS 0.359654f
C85 B.n51 VSUBS 0.241844f
C86 B.n52 VSUBS 0.016965f
C87 B.n53 VSUBS 0.007322f
C88 B.n54 VSUBS 0.007322f
C89 B.n55 VSUBS 0.007322f
C90 B.n56 VSUBS 0.007322f
C91 B.n57 VSUBS 0.007322f
C92 B.n58 VSUBS 0.007322f
C93 B.n59 VSUBS 0.007322f
C94 B.n60 VSUBS 0.007322f
C95 B.n61 VSUBS 0.007322f
C96 B.n62 VSUBS 0.007322f
C97 B.n63 VSUBS 0.007322f
C98 B.n64 VSUBS 0.007322f
C99 B.n65 VSUBS 0.007322f
C100 B.n66 VSUBS 0.007322f
C101 B.n67 VSUBS 0.007322f
C102 B.n68 VSUBS 0.007322f
C103 B.n69 VSUBS 0.007322f
C104 B.n70 VSUBS 0.017789f
C105 B.n71 VSUBS 0.007322f
C106 B.n72 VSUBS 0.007322f
C107 B.n73 VSUBS 0.007322f
C108 B.n74 VSUBS 0.007322f
C109 B.n75 VSUBS 0.007322f
C110 B.n76 VSUBS 0.007322f
C111 B.n77 VSUBS 0.007322f
C112 B.n78 VSUBS 0.007322f
C113 B.n79 VSUBS 0.007322f
C114 B.n80 VSUBS 0.007322f
C115 B.n81 VSUBS 0.007322f
C116 B.n82 VSUBS 0.007322f
C117 B.n83 VSUBS 0.007322f
C118 B.n84 VSUBS 0.007322f
C119 B.n85 VSUBS 0.007322f
C120 B.n86 VSUBS 0.007322f
C121 B.n87 VSUBS 0.007322f
C122 B.n88 VSUBS 0.007322f
C123 B.n89 VSUBS 0.007322f
C124 B.n90 VSUBS 0.007322f
C125 B.n91 VSUBS 0.007322f
C126 B.n92 VSUBS 0.007322f
C127 B.n93 VSUBS 0.007322f
C128 B.n94 VSUBS 0.007322f
C129 B.n95 VSUBS 0.007322f
C130 B.n96 VSUBS 0.007322f
C131 B.n97 VSUBS 0.007322f
C132 B.n98 VSUBS 0.007322f
C133 B.n99 VSUBS 0.007322f
C134 B.n100 VSUBS 0.007322f
C135 B.n101 VSUBS 0.007322f
C136 B.n102 VSUBS 0.007322f
C137 B.n103 VSUBS 0.007322f
C138 B.n104 VSUBS 0.007322f
C139 B.n105 VSUBS 0.007322f
C140 B.n106 VSUBS 0.007322f
C141 B.n107 VSUBS 0.007322f
C142 B.n108 VSUBS 0.007322f
C143 B.n109 VSUBS 0.007322f
C144 B.n110 VSUBS 0.007322f
C145 B.n111 VSUBS 0.007322f
C146 B.n112 VSUBS 0.007322f
C147 B.n113 VSUBS 0.007322f
C148 B.n114 VSUBS 0.007322f
C149 B.n115 VSUBS 0.007322f
C150 B.n116 VSUBS 0.007322f
C151 B.n117 VSUBS 0.018586f
C152 B.n118 VSUBS 0.007322f
C153 B.n119 VSUBS 0.007322f
C154 B.n120 VSUBS 0.007322f
C155 B.n121 VSUBS 0.007322f
C156 B.n122 VSUBS 0.007322f
C157 B.n123 VSUBS 0.007322f
C158 B.n124 VSUBS 0.007322f
C159 B.n125 VSUBS 0.007322f
C160 B.n126 VSUBS 0.007322f
C161 B.n127 VSUBS 0.007322f
C162 B.n128 VSUBS 0.007322f
C163 B.n129 VSUBS 0.007322f
C164 B.n130 VSUBS 0.007322f
C165 B.n131 VSUBS 0.007322f
C166 B.n132 VSUBS 0.007322f
C167 B.n133 VSUBS 0.007322f
C168 B.n134 VSUBS 0.007322f
C169 B.n135 VSUBS 0.007322f
C170 B.t10 VSUBS 0.179512f
C171 B.t11 VSUBS 0.224931f
C172 B.t9 VSUBS 2.00302f
C173 B.n136 VSUBS 0.359654f
C174 B.n137 VSUBS 0.241844f
C175 B.n138 VSUBS 0.007322f
C176 B.n139 VSUBS 0.007322f
C177 B.n140 VSUBS 0.007322f
C178 B.n141 VSUBS 0.007322f
C179 B.t1 VSUBS 0.179509f
C180 B.t2 VSUBS 0.224929f
C181 B.t0 VSUBS 2.00302f
C182 B.n142 VSUBS 0.359657f
C183 B.n143 VSUBS 0.241847f
C184 B.n144 VSUBS 0.016965f
C185 B.n145 VSUBS 0.007322f
C186 B.n146 VSUBS 0.007322f
C187 B.n147 VSUBS 0.007322f
C188 B.n148 VSUBS 0.007322f
C189 B.n149 VSUBS 0.007322f
C190 B.n150 VSUBS 0.007322f
C191 B.n151 VSUBS 0.007322f
C192 B.n152 VSUBS 0.007322f
C193 B.n153 VSUBS 0.007322f
C194 B.n154 VSUBS 0.007322f
C195 B.n155 VSUBS 0.007322f
C196 B.n156 VSUBS 0.007322f
C197 B.n157 VSUBS 0.007322f
C198 B.n158 VSUBS 0.007322f
C199 B.n159 VSUBS 0.007322f
C200 B.n160 VSUBS 0.007322f
C201 B.n161 VSUBS 0.007322f
C202 B.n162 VSUBS 0.018586f
C203 B.n163 VSUBS 0.007322f
C204 B.n164 VSUBS 0.007322f
C205 B.n165 VSUBS 0.007322f
C206 B.n166 VSUBS 0.007322f
C207 B.n167 VSUBS 0.007322f
C208 B.n168 VSUBS 0.007322f
C209 B.n169 VSUBS 0.007322f
C210 B.n170 VSUBS 0.007322f
C211 B.n171 VSUBS 0.007322f
C212 B.n172 VSUBS 0.007322f
C213 B.n173 VSUBS 0.007322f
C214 B.n174 VSUBS 0.007322f
C215 B.n175 VSUBS 0.007322f
C216 B.n176 VSUBS 0.007322f
C217 B.n177 VSUBS 0.007322f
C218 B.n178 VSUBS 0.007322f
C219 B.n179 VSUBS 0.007322f
C220 B.n180 VSUBS 0.007322f
C221 B.n181 VSUBS 0.007322f
C222 B.n182 VSUBS 0.007322f
C223 B.n183 VSUBS 0.007322f
C224 B.n184 VSUBS 0.007322f
C225 B.n185 VSUBS 0.007322f
C226 B.n186 VSUBS 0.007322f
C227 B.n187 VSUBS 0.007322f
C228 B.n188 VSUBS 0.007322f
C229 B.n189 VSUBS 0.007322f
C230 B.n190 VSUBS 0.007322f
C231 B.n191 VSUBS 0.007322f
C232 B.n192 VSUBS 0.007322f
C233 B.n193 VSUBS 0.007322f
C234 B.n194 VSUBS 0.007322f
C235 B.n195 VSUBS 0.007322f
C236 B.n196 VSUBS 0.007322f
C237 B.n197 VSUBS 0.007322f
C238 B.n198 VSUBS 0.007322f
C239 B.n199 VSUBS 0.007322f
C240 B.n200 VSUBS 0.007322f
C241 B.n201 VSUBS 0.007322f
C242 B.n202 VSUBS 0.007322f
C243 B.n203 VSUBS 0.007322f
C244 B.n204 VSUBS 0.007322f
C245 B.n205 VSUBS 0.007322f
C246 B.n206 VSUBS 0.007322f
C247 B.n207 VSUBS 0.007322f
C248 B.n208 VSUBS 0.007322f
C249 B.n209 VSUBS 0.007322f
C250 B.n210 VSUBS 0.007322f
C251 B.n211 VSUBS 0.007322f
C252 B.n212 VSUBS 0.007322f
C253 B.n213 VSUBS 0.007322f
C254 B.n214 VSUBS 0.007322f
C255 B.n215 VSUBS 0.007322f
C256 B.n216 VSUBS 0.007322f
C257 B.n217 VSUBS 0.007322f
C258 B.n218 VSUBS 0.007322f
C259 B.n219 VSUBS 0.007322f
C260 B.n220 VSUBS 0.007322f
C261 B.n221 VSUBS 0.007322f
C262 B.n222 VSUBS 0.007322f
C263 B.n223 VSUBS 0.007322f
C264 B.n224 VSUBS 0.007322f
C265 B.n225 VSUBS 0.007322f
C266 B.n226 VSUBS 0.007322f
C267 B.n227 VSUBS 0.007322f
C268 B.n228 VSUBS 0.007322f
C269 B.n229 VSUBS 0.007322f
C270 B.n230 VSUBS 0.007322f
C271 B.n231 VSUBS 0.007322f
C272 B.n232 VSUBS 0.007322f
C273 B.n233 VSUBS 0.007322f
C274 B.n234 VSUBS 0.007322f
C275 B.n235 VSUBS 0.007322f
C276 B.n236 VSUBS 0.007322f
C277 B.n237 VSUBS 0.007322f
C278 B.n238 VSUBS 0.007322f
C279 B.n239 VSUBS 0.007322f
C280 B.n240 VSUBS 0.007322f
C281 B.n241 VSUBS 0.007322f
C282 B.n242 VSUBS 0.007322f
C283 B.n243 VSUBS 0.007322f
C284 B.n244 VSUBS 0.007322f
C285 B.n245 VSUBS 0.007322f
C286 B.n246 VSUBS 0.007322f
C287 B.n247 VSUBS 0.007322f
C288 B.n248 VSUBS 0.007322f
C289 B.n249 VSUBS 0.007322f
C290 B.n250 VSUBS 0.007322f
C291 B.n251 VSUBS 0.017594f
C292 B.n252 VSUBS 0.017594f
C293 B.n253 VSUBS 0.018586f
C294 B.n254 VSUBS 0.007322f
C295 B.n255 VSUBS 0.007322f
C296 B.n256 VSUBS 0.007322f
C297 B.n257 VSUBS 0.007322f
C298 B.n258 VSUBS 0.007322f
C299 B.n259 VSUBS 0.007322f
C300 B.n260 VSUBS 0.007322f
C301 B.n261 VSUBS 0.007322f
C302 B.n262 VSUBS 0.007322f
C303 B.n263 VSUBS 0.007322f
C304 B.n264 VSUBS 0.007322f
C305 B.n265 VSUBS 0.007322f
C306 B.n266 VSUBS 0.007322f
C307 B.n267 VSUBS 0.007322f
C308 B.n268 VSUBS 0.007322f
C309 B.n269 VSUBS 0.007322f
C310 B.n270 VSUBS 0.007322f
C311 B.n271 VSUBS 0.007322f
C312 B.n272 VSUBS 0.007322f
C313 B.n273 VSUBS 0.007322f
C314 B.n274 VSUBS 0.007322f
C315 B.n275 VSUBS 0.007322f
C316 B.n276 VSUBS 0.007322f
C317 B.n277 VSUBS 0.007322f
C318 B.n278 VSUBS 0.007322f
C319 B.n279 VSUBS 0.007322f
C320 B.n280 VSUBS 0.007322f
C321 B.n281 VSUBS 0.007322f
C322 B.n282 VSUBS 0.007322f
C323 B.n283 VSUBS 0.007322f
C324 B.n284 VSUBS 0.007322f
C325 B.n285 VSUBS 0.007322f
C326 B.n286 VSUBS 0.007322f
C327 B.n287 VSUBS 0.007322f
C328 B.n288 VSUBS 0.007322f
C329 B.n289 VSUBS 0.007322f
C330 B.n290 VSUBS 0.007322f
C331 B.n291 VSUBS 0.007322f
C332 B.n292 VSUBS 0.007322f
C333 B.n293 VSUBS 0.007322f
C334 B.n294 VSUBS 0.007322f
C335 B.n295 VSUBS 0.007322f
C336 B.n296 VSUBS 0.007322f
C337 B.n297 VSUBS 0.007322f
C338 B.n298 VSUBS 0.007322f
C339 B.n299 VSUBS 0.007322f
C340 B.n300 VSUBS 0.007322f
C341 B.n301 VSUBS 0.007322f
C342 B.n302 VSUBS 0.007322f
C343 B.n303 VSUBS 0.007322f
C344 B.n304 VSUBS 0.007322f
C345 B.n305 VSUBS 0.006891f
C346 B.n306 VSUBS 0.007322f
C347 B.n307 VSUBS 0.007322f
C348 B.n308 VSUBS 0.004092f
C349 B.n309 VSUBS 0.007322f
C350 B.n310 VSUBS 0.007322f
C351 B.n311 VSUBS 0.007322f
C352 B.n312 VSUBS 0.007322f
C353 B.n313 VSUBS 0.007322f
C354 B.n314 VSUBS 0.007322f
C355 B.n315 VSUBS 0.007322f
C356 B.n316 VSUBS 0.007322f
C357 B.n317 VSUBS 0.007322f
C358 B.n318 VSUBS 0.007322f
C359 B.n319 VSUBS 0.007322f
C360 B.n320 VSUBS 0.007322f
C361 B.n321 VSUBS 0.004092f
C362 B.n322 VSUBS 0.016965f
C363 B.n323 VSUBS 0.006891f
C364 B.n324 VSUBS 0.007322f
C365 B.n325 VSUBS 0.007322f
C366 B.n326 VSUBS 0.007322f
C367 B.n327 VSUBS 0.007322f
C368 B.n328 VSUBS 0.007322f
C369 B.n329 VSUBS 0.007322f
C370 B.n330 VSUBS 0.007322f
C371 B.n331 VSUBS 0.007322f
C372 B.n332 VSUBS 0.007322f
C373 B.n333 VSUBS 0.007322f
C374 B.n334 VSUBS 0.007322f
C375 B.n335 VSUBS 0.007322f
C376 B.n336 VSUBS 0.007322f
C377 B.n337 VSUBS 0.007322f
C378 B.n338 VSUBS 0.007322f
C379 B.n339 VSUBS 0.007322f
C380 B.n340 VSUBS 0.007322f
C381 B.n341 VSUBS 0.007322f
C382 B.n342 VSUBS 0.007322f
C383 B.n343 VSUBS 0.007322f
C384 B.n344 VSUBS 0.007322f
C385 B.n345 VSUBS 0.007322f
C386 B.n346 VSUBS 0.007322f
C387 B.n347 VSUBS 0.007322f
C388 B.n348 VSUBS 0.007322f
C389 B.n349 VSUBS 0.007322f
C390 B.n350 VSUBS 0.007322f
C391 B.n351 VSUBS 0.007322f
C392 B.n352 VSUBS 0.007322f
C393 B.n353 VSUBS 0.007322f
C394 B.n354 VSUBS 0.007322f
C395 B.n355 VSUBS 0.007322f
C396 B.n356 VSUBS 0.007322f
C397 B.n357 VSUBS 0.007322f
C398 B.n358 VSUBS 0.007322f
C399 B.n359 VSUBS 0.007322f
C400 B.n360 VSUBS 0.007322f
C401 B.n361 VSUBS 0.007322f
C402 B.n362 VSUBS 0.007322f
C403 B.n363 VSUBS 0.007322f
C404 B.n364 VSUBS 0.007322f
C405 B.n365 VSUBS 0.007322f
C406 B.n366 VSUBS 0.007322f
C407 B.n367 VSUBS 0.007322f
C408 B.n368 VSUBS 0.007322f
C409 B.n369 VSUBS 0.007322f
C410 B.n370 VSUBS 0.007322f
C411 B.n371 VSUBS 0.007322f
C412 B.n372 VSUBS 0.007322f
C413 B.n373 VSUBS 0.007322f
C414 B.n374 VSUBS 0.007322f
C415 B.n375 VSUBS 0.007322f
C416 B.n376 VSUBS 0.018586f
C417 B.n377 VSUBS 0.017594f
C418 B.n378 VSUBS 0.017594f
C419 B.n379 VSUBS 0.007322f
C420 B.n380 VSUBS 0.007322f
C421 B.n381 VSUBS 0.007322f
C422 B.n382 VSUBS 0.007322f
C423 B.n383 VSUBS 0.007322f
C424 B.n384 VSUBS 0.007322f
C425 B.n385 VSUBS 0.007322f
C426 B.n386 VSUBS 0.007322f
C427 B.n387 VSUBS 0.007322f
C428 B.n388 VSUBS 0.007322f
C429 B.n389 VSUBS 0.007322f
C430 B.n390 VSUBS 0.007322f
C431 B.n391 VSUBS 0.007322f
C432 B.n392 VSUBS 0.007322f
C433 B.n393 VSUBS 0.007322f
C434 B.n394 VSUBS 0.007322f
C435 B.n395 VSUBS 0.007322f
C436 B.n396 VSUBS 0.007322f
C437 B.n397 VSUBS 0.007322f
C438 B.n398 VSUBS 0.007322f
C439 B.n399 VSUBS 0.007322f
C440 B.n400 VSUBS 0.007322f
C441 B.n401 VSUBS 0.007322f
C442 B.n402 VSUBS 0.007322f
C443 B.n403 VSUBS 0.007322f
C444 B.n404 VSUBS 0.007322f
C445 B.n405 VSUBS 0.007322f
C446 B.n406 VSUBS 0.007322f
C447 B.n407 VSUBS 0.007322f
C448 B.n408 VSUBS 0.007322f
C449 B.n409 VSUBS 0.007322f
C450 B.n410 VSUBS 0.007322f
C451 B.n411 VSUBS 0.007322f
C452 B.n412 VSUBS 0.007322f
C453 B.n413 VSUBS 0.007322f
C454 B.n414 VSUBS 0.007322f
C455 B.n415 VSUBS 0.007322f
C456 B.n416 VSUBS 0.007322f
C457 B.n417 VSUBS 0.007322f
C458 B.n418 VSUBS 0.007322f
C459 B.n419 VSUBS 0.007322f
C460 B.n420 VSUBS 0.007322f
C461 B.n421 VSUBS 0.007322f
C462 B.n422 VSUBS 0.007322f
C463 B.n423 VSUBS 0.007322f
C464 B.n424 VSUBS 0.007322f
C465 B.n425 VSUBS 0.007322f
C466 B.n426 VSUBS 0.007322f
C467 B.n427 VSUBS 0.007322f
C468 B.n428 VSUBS 0.007322f
C469 B.n429 VSUBS 0.007322f
C470 B.n430 VSUBS 0.007322f
C471 B.n431 VSUBS 0.007322f
C472 B.n432 VSUBS 0.007322f
C473 B.n433 VSUBS 0.007322f
C474 B.n434 VSUBS 0.007322f
C475 B.n435 VSUBS 0.007322f
C476 B.n436 VSUBS 0.007322f
C477 B.n437 VSUBS 0.007322f
C478 B.n438 VSUBS 0.007322f
C479 B.n439 VSUBS 0.007322f
C480 B.n440 VSUBS 0.007322f
C481 B.n441 VSUBS 0.007322f
C482 B.n442 VSUBS 0.007322f
C483 B.n443 VSUBS 0.007322f
C484 B.n444 VSUBS 0.007322f
C485 B.n445 VSUBS 0.007322f
C486 B.n446 VSUBS 0.007322f
C487 B.n447 VSUBS 0.007322f
C488 B.n448 VSUBS 0.007322f
C489 B.n449 VSUBS 0.007322f
C490 B.n450 VSUBS 0.007322f
C491 B.n451 VSUBS 0.007322f
C492 B.n452 VSUBS 0.007322f
C493 B.n453 VSUBS 0.007322f
C494 B.n454 VSUBS 0.007322f
C495 B.n455 VSUBS 0.007322f
C496 B.n456 VSUBS 0.007322f
C497 B.n457 VSUBS 0.007322f
C498 B.n458 VSUBS 0.007322f
C499 B.n459 VSUBS 0.007322f
C500 B.n460 VSUBS 0.007322f
C501 B.n461 VSUBS 0.007322f
C502 B.n462 VSUBS 0.007322f
C503 B.n463 VSUBS 0.007322f
C504 B.n464 VSUBS 0.007322f
C505 B.n465 VSUBS 0.007322f
C506 B.n466 VSUBS 0.007322f
C507 B.n467 VSUBS 0.007322f
C508 B.n468 VSUBS 0.007322f
C509 B.n469 VSUBS 0.007322f
C510 B.n470 VSUBS 0.007322f
C511 B.n471 VSUBS 0.007322f
C512 B.n472 VSUBS 0.007322f
C513 B.n473 VSUBS 0.007322f
C514 B.n474 VSUBS 0.007322f
C515 B.n475 VSUBS 0.007322f
C516 B.n476 VSUBS 0.007322f
C517 B.n477 VSUBS 0.007322f
C518 B.n478 VSUBS 0.007322f
C519 B.n479 VSUBS 0.007322f
C520 B.n480 VSUBS 0.007322f
C521 B.n481 VSUBS 0.007322f
C522 B.n482 VSUBS 0.007322f
C523 B.n483 VSUBS 0.007322f
C524 B.n484 VSUBS 0.007322f
C525 B.n485 VSUBS 0.007322f
C526 B.n486 VSUBS 0.007322f
C527 B.n487 VSUBS 0.007322f
C528 B.n488 VSUBS 0.007322f
C529 B.n489 VSUBS 0.007322f
C530 B.n490 VSUBS 0.007322f
C531 B.n491 VSUBS 0.007322f
C532 B.n492 VSUBS 0.007322f
C533 B.n493 VSUBS 0.007322f
C534 B.n494 VSUBS 0.007322f
C535 B.n495 VSUBS 0.007322f
C536 B.n496 VSUBS 0.007322f
C537 B.n497 VSUBS 0.007322f
C538 B.n498 VSUBS 0.007322f
C539 B.n499 VSUBS 0.007322f
C540 B.n500 VSUBS 0.007322f
C541 B.n501 VSUBS 0.007322f
C542 B.n502 VSUBS 0.007322f
C543 B.n503 VSUBS 0.007322f
C544 B.n504 VSUBS 0.007322f
C545 B.n505 VSUBS 0.007322f
C546 B.n506 VSUBS 0.007322f
C547 B.n507 VSUBS 0.007322f
C548 B.n508 VSUBS 0.007322f
C549 B.n509 VSUBS 0.007322f
C550 B.n510 VSUBS 0.007322f
C551 B.n511 VSUBS 0.007322f
C552 B.n512 VSUBS 0.007322f
C553 B.n513 VSUBS 0.007322f
C554 B.n514 VSUBS 0.007322f
C555 B.n515 VSUBS 0.018392f
C556 B.n516 VSUBS 0.017594f
C557 B.n517 VSUBS 0.018586f
C558 B.n518 VSUBS 0.007322f
C559 B.n519 VSUBS 0.007322f
C560 B.n520 VSUBS 0.007322f
C561 B.n521 VSUBS 0.007322f
C562 B.n522 VSUBS 0.007322f
C563 B.n523 VSUBS 0.007322f
C564 B.n524 VSUBS 0.007322f
C565 B.n525 VSUBS 0.007322f
C566 B.n526 VSUBS 0.007322f
C567 B.n527 VSUBS 0.007322f
C568 B.n528 VSUBS 0.007322f
C569 B.n529 VSUBS 0.007322f
C570 B.n530 VSUBS 0.007322f
C571 B.n531 VSUBS 0.007322f
C572 B.n532 VSUBS 0.007322f
C573 B.n533 VSUBS 0.007322f
C574 B.n534 VSUBS 0.007322f
C575 B.n535 VSUBS 0.007322f
C576 B.n536 VSUBS 0.007322f
C577 B.n537 VSUBS 0.007322f
C578 B.n538 VSUBS 0.007322f
C579 B.n539 VSUBS 0.007322f
C580 B.n540 VSUBS 0.007322f
C581 B.n541 VSUBS 0.007322f
C582 B.n542 VSUBS 0.007322f
C583 B.n543 VSUBS 0.007322f
C584 B.n544 VSUBS 0.007322f
C585 B.n545 VSUBS 0.007322f
C586 B.n546 VSUBS 0.007322f
C587 B.n547 VSUBS 0.007322f
C588 B.n548 VSUBS 0.007322f
C589 B.n549 VSUBS 0.007322f
C590 B.n550 VSUBS 0.007322f
C591 B.n551 VSUBS 0.007322f
C592 B.n552 VSUBS 0.007322f
C593 B.n553 VSUBS 0.007322f
C594 B.n554 VSUBS 0.007322f
C595 B.n555 VSUBS 0.007322f
C596 B.n556 VSUBS 0.007322f
C597 B.n557 VSUBS 0.007322f
C598 B.n558 VSUBS 0.007322f
C599 B.n559 VSUBS 0.007322f
C600 B.n560 VSUBS 0.007322f
C601 B.n561 VSUBS 0.007322f
C602 B.n562 VSUBS 0.007322f
C603 B.n563 VSUBS 0.007322f
C604 B.n564 VSUBS 0.007322f
C605 B.n565 VSUBS 0.007322f
C606 B.n566 VSUBS 0.007322f
C607 B.n567 VSUBS 0.007322f
C608 B.n568 VSUBS 0.007322f
C609 B.n569 VSUBS 0.006891f
C610 B.n570 VSUBS 0.007322f
C611 B.n571 VSUBS 0.007322f
C612 B.n572 VSUBS 0.004092f
C613 B.n573 VSUBS 0.007322f
C614 B.n574 VSUBS 0.007322f
C615 B.n575 VSUBS 0.007322f
C616 B.n576 VSUBS 0.007322f
C617 B.n577 VSUBS 0.007322f
C618 B.n578 VSUBS 0.007322f
C619 B.n579 VSUBS 0.007322f
C620 B.n580 VSUBS 0.007322f
C621 B.n581 VSUBS 0.007322f
C622 B.n582 VSUBS 0.007322f
C623 B.n583 VSUBS 0.007322f
C624 B.n584 VSUBS 0.007322f
C625 B.n585 VSUBS 0.004092f
C626 B.n586 VSUBS 0.016965f
C627 B.n587 VSUBS 0.006891f
C628 B.n588 VSUBS 0.007322f
C629 B.n589 VSUBS 0.007322f
C630 B.n590 VSUBS 0.007322f
C631 B.n591 VSUBS 0.007322f
C632 B.n592 VSUBS 0.007322f
C633 B.n593 VSUBS 0.007322f
C634 B.n594 VSUBS 0.007322f
C635 B.n595 VSUBS 0.007322f
C636 B.n596 VSUBS 0.007322f
C637 B.n597 VSUBS 0.007322f
C638 B.n598 VSUBS 0.007322f
C639 B.n599 VSUBS 0.007322f
C640 B.n600 VSUBS 0.007322f
C641 B.n601 VSUBS 0.007322f
C642 B.n602 VSUBS 0.007322f
C643 B.n603 VSUBS 0.007322f
C644 B.n604 VSUBS 0.007322f
C645 B.n605 VSUBS 0.007322f
C646 B.n606 VSUBS 0.007322f
C647 B.n607 VSUBS 0.007322f
C648 B.n608 VSUBS 0.007322f
C649 B.n609 VSUBS 0.007322f
C650 B.n610 VSUBS 0.007322f
C651 B.n611 VSUBS 0.007322f
C652 B.n612 VSUBS 0.007322f
C653 B.n613 VSUBS 0.007322f
C654 B.n614 VSUBS 0.007322f
C655 B.n615 VSUBS 0.007322f
C656 B.n616 VSUBS 0.007322f
C657 B.n617 VSUBS 0.007322f
C658 B.n618 VSUBS 0.007322f
C659 B.n619 VSUBS 0.007322f
C660 B.n620 VSUBS 0.007322f
C661 B.n621 VSUBS 0.007322f
C662 B.n622 VSUBS 0.007322f
C663 B.n623 VSUBS 0.007322f
C664 B.n624 VSUBS 0.007322f
C665 B.n625 VSUBS 0.007322f
C666 B.n626 VSUBS 0.007322f
C667 B.n627 VSUBS 0.007322f
C668 B.n628 VSUBS 0.007322f
C669 B.n629 VSUBS 0.007322f
C670 B.n630 VSUBS 0.007322f
C671 B.n631 VSUBS 0.007322f
C672 B.n632 VSUBS 0.007322f
C673 B.n633 VSUBS 0.007322f
C674 B.n634 VSUBS 0.007322f
C675 B.n635 VSUBS 0.007322f
C676 B.n636 VSUBS 0.007322f
C677 B.n637 VSUBS 0.007322f
C678 B.n638 VSUBS 0.007322f
C679 B.n639 VSUBS 0.007322f
C680 B.n640 VSUBS 0.018586f
C681 B.n641 VSUBS 0.017594f
C682 B.n642 VSUBS 0.017594f
C683 B.n643 VSUBS 0.007322f
C684 B.n644 VSUBS 0.007322f
C685 B.n645 VSUBS 0.007322f
C686 B.n646 VSUBS 0.007322f
C687 B.n647 VSUBS 0.007322f
C688 B.n648 VSUBS 0.007322f
C689 B.n649 VSUBS 0.007322f
C690 B.n650 VSUBS 0.007322f
C691 B.n651 VSUBS 0.007322f
C692 B.n652 VSUBS 0.007322f
C693 B.n653 VSUBS 0.007322f
C694 B.n654 VSUBS 0.007322f
C695 B.n655 VSUBS 0.007322f
C696 B.n656 VSUBS 0.007322f
C697 B.n657 VSUBS 0.007322f
C698 B.n658 VSUBS 0.007322f
C699 B.n659 VSUBS 0.007322f
C700 B.n660 VSUBS 0.007322f
C701 B.n661 VSUBS 0.007322f
C702 B.n662 VSUBS 0.007322f
C703 B.n663 VSUBS 0.007322f
C704 B.n664 VSUBS 0.007322f
C705 B.n665 VSUBS 0.007322f
C706 B.n666 VSUBS 0.007322f
C707 B.n667 VSUBS 0.007322f
C708 B.n668 VSUBS 0.007322f
C709 B.n669 VSUBS 0.007322f
C710 B.n670 VSUBS 0.007322f
C711 B.n671 VSUBS 0.007322f
C712 B.n672 VSUBS 0.007322f
C713 B.n673 VSUBS 0.007322f
C714 B.n674 VSUBS 0.007322f
C715 B.n675 VSUBS 0.007322f
C716 B.n676 VSUBS 0.007322f
C717 B.n677 VSUBS 0.007322f
C718 B.n678 VSUBS 0.007322f
C719 B.n679 VSUBS 0.007322f
C720 B.n680 VSUBS 0.007322f
C721 B.n681 VSUBS 0.007322f
C722 B.n682 VSUBS 0.007322f
C723 B.n683 VSUBS 0.007322f
C724 B.n684 VSUBS 0.007322f
C725 B.n685 VSUBS 0.007322f
C726 B.n686 VSUBS 0.007322f
C727 B.n687 VSUBS 0.007322f
C728 B.n688 VSUBS 0.007322f
C729 B.n689 VSUBS 0.007322f
C730 B.n690 VSUBS 0.007322f
C731 B.n691 VSUBS 0.007322f
C732 B.n692 VSUBS 0.007322f
C733 B.n693 VSUBS 0.007322f
C734 B.n694 VSUBS 0.007322f
C735 B.n695 VSUBS 0.007322f
C736 B.n696 VSUBS 0.007322f
C737 B.n697 VSUBS 0.007322f
C738 B.n698 VSUBS 0.007322f
C739 B.n699 VSUBS 0.007322f
C740 B.n700 VSUBS 0.007322f
C741 B.n701 VSUBS 0.007322f
C742 B.n702 VSUBS 0.007322f
C743 B.n703 VSUBS 0.007322f
C744 B.n704 VSUBS 0.007322f
C745 B.n705 VSUBS 0.007322f
C746 B.n706 VSUBS 0.007322f
C747 B.n707 VSUBS 0.007322f
C748 B.n708 VSUBS 0.007322f
C749 B.n709 VSUBS 0.007322f
C750 B.n710 VSUBS 0.007322f
C751 B.n711 VSUBS 0.01658f
C752 VDD2.t1 VSUBS 0.221097f
C753 VDD2.t3 VSUBS 0.221097f
C754 VDD2.n0 VSUBS 2.36628f
C755 VDD2.t0 VSUBS 0.221097f
C756 VDD2.t2 VSUBS 0.221097f
C757 VDD2.n1 VSUBS 1.68798f
C758 VDD2.n2 VSUBS 4.52563f
C759 VN.t2 VSUBS 3.54773f
C760 VN.t0 VSUBS 3.52866f
C761 VN.n0 VSUBS 2.08642f
C762 VN.t1 VSUBS 3.54773f
C763 VN.t3 VSUBS 3.52866f
C764 VN.n1 VSUBS 3.90004f
C765 VDD1.t1 VSUBS 0.225529f
C766 VDD1.t2 VSUBS 0.225529f
C767 VDD1.n0 VSUBS 1.72242f
C768 VDD1.t0 VSUBS 0.225529f
C769 VDD1.t3 VSUBS 0.225529f
C770 VDD1.n1 VSUBS 2.43856f
C771 VTAIL.n0 VSUBS 0.029168f
C772 VTAIL.n1 VSUBS 0.025653f
C773 VTAIL.n2 VSUBS 0.013785f
C774 VTAIL.n3 VSUBS 0.032583f
C775 VTAIL.n4 VSUBS 0.014596f
C776 VTAIL.n5 VSUBS 0.025653f
C777 VTAIL.n6 VSUBS 0.01419f
C778 VTAIL.n7 VSUBS 0.032583f
C779 VTAIL.n8 VSUBS 0.014596f
C780 VTAIL.n9 VSUBS 0.025653f
C781 VTAIL.n10 VSUBS 0.013785f
C782 VTAIL.n11 VSUBS 0.032583f
C783 VTAIL.n12 VSUBS 0.014596f
C784 VTAIL.n13 VSUBS 0.025653f
C785 VTAIL.n14 VSUBS 0.013785f
C786 VTAIL.n15 VSUBS 0.024437f
C787 VTAIL.n16 VSUBS 0.02451f
C788 VTAIL.t6 VSUBS 0.070084f
C789 VTAIL.n17 VSUBS 0.18095f
C790 VTAIL.n18 VSUBS 1.0558f
C791 VTAIL.n19 VSUBS 0.013785f
C792 VTAIL.n20 VSUBS 0.014596f
C793 VTAIL.n21 VSUBS 0.032583f
C794 VTAIL.n22 VSUBS 0.032583f
C795 VTAIL.n23 VSUBS 0.014596f
C796 VTAIL.n24 VSUBS 0.013785f
C797 VTAIL.n25 VSUBS 0.025653f
C798 VTAIL.n26 VSUBS 0.025653f
C799 VTAIL.n27 VSUBS 0.013785f
C800 VTAIL.n28 VSUBS 0.014596f
C801 VTAIL.n29 VSUBS 0.032583f
C802 VTAIL.n30 VSUBS 0.032583f
C803 VTAIL.n31 VSUBS 0.014596f
C804 VTAIL.n32 VSUBS 0.013785f
C805 VTAIL.n33 VSUBS 0.025653f
C806 VTAIL.n34 VSUBS 0.025653f
C807 VTAIL.n35 VSUBS 0.013785f
C808 VTAIL.n36 VSUBS 0.013785f
C809 VTAIL.n37 VSUBS 0.014596f
C810 VTAIL.n38 VSUBS 0.032583f
C811 VTAIL.n39 VSUBS 0.032583f
C812 VTAIL.n40 VSUBS 0.032583f
C813 VTAIL.n41 VSUBS 0.01419f
C814 VTAIL.n42 VSUBS 0.013785f
C815 VTAIL.n43 VSUBS 0.025653f
C816 VTAIL.n44 VSUBS 0.025653f
C817 VTAIL.n45 VSUBS 0.013785f
C818 VTAIL.n46 VSUBS 0.014596f
C819 VTAIL.n47 VSUBS 0.032583f
C820 VTAIL.n48 VSUBS 0.082218f
C821 VTAIL.n49 VSUBS 0.014596f
C822 VTAIL.n50 VSUBS 0.013785f
C823 VTAIL.n51 VSUBS 0.067006f
C824 VTAIL.n52 VSUBS 0.041719f
C825 VTAIL.n53 VSUBS 0.223841f
C826 VTAIL.n54 VSUBS 0.029168f
C827 VTAIL.n55 VSUBS 0.025653f
C828 VTAIL.n56 VSUBS 0.013785f
C829 VTAIL.n57 VSUBS 0.032583f
C830 VTAIL.n58 VSUBS 0.014596f
C831 VTAIL.n59 VSUBS 0.025653f
C832 VTAIL.n60 VSUBS 0.01419f
C833 VTAIL.n61 VSUBS 0.032583f
C834 VTAIL.n62 VSUBS 0.014596f
C835 VTAIL.n63 VSUBS 0.025653f
C836 VTAIL.n64 VSUBS 0.013785f
C837 VTAIL.n65 VSUBS 0.032583f
C838 VTAIL.n66 VSUBS 0.014596f
C839 VTAIL.n67 VSUBS 0.025653f
C840 VTAIL.n68 VSUBS 0.013785f
C841 VTAIL.n69 VSUBS 0.024437f
C842 VTAIL.n70 VSUBS 0.02451f
C843 VTAIL.t2 VSUBS 0.070084f
C844 VTAIL.n71 VSUBS 0.18095f
C845 VTAIL.n72 VSUBS 1.0558f
C846 VTAIL.n73 VSUBS 0.013785f
C847 VTAIL.n74 VSUBS 0.014596f
C848 VTAIL.n75 VSUBS 0.032583f
C849 VTAIL.n76 VSUBS 0.032583f
C850 VTAIL.n77 VSUBS 0.014596f
C851 VTAIL.n78 VSUBS 0.013785f
C852 VTAIL.n79 VSUBS 0.025653f
C853 VTAIL.n80 VSUBS 0.025653f
C854 VTAIL.n81 VSUBS 0.013785f
C855 VTAIL.n82 VSUBS 0.014596f
C856 VTAIL.n83 VSUBS 0.032583f
C857 VTAIL.n84 VSUBS 0.032583f
C858 VTAIL.n85 VSUBS 0.014596f
C859 VTAIL.n86 VSUBS 0.013785f
C860 VTAIL.n87 VSUBS 0.025653f
C861 VTAIL.n88 VSUBS 0.025653f
C862 VTAIL.n89 VSUBS 0.013785f
C863 VTAIL.n90 VSUBS 0.013785f
C864 VTAIL.n91 VSUBS 0.014596f
C865 VTAIL.n92 VSUBS 0.032583f
C866 VTAIL.n93 VSUBS 0.032583f
C867 VTAIL.n94 VSUBS 0.032583f
C868 VTAIL.n95 VSUBS 0.01419f
C869 VTAIL.n96 VSUBS 0.013785f
C870 VTAIL.n97 VSUBS 0.025653f
C871 VTAIL.n98 VSUBS 0.025653f
C872 VTAIL.n99 VSUBS 0.013785f
C873 VTAIL.n100 VSUBS 0.014596f
C874 VTAIL.n101 VSUBS 0.032583f
C875 VTAIL.n102 VSUBS 0.082218f
C876 VTAIL.n103 VSUBS 0.014596f
C877 VTAIL.n104 VSUBS 0.013785f
C878 VTAIL.n105 VSUBS 0.067006f
C879 VTAIL.n106 VSUBS 0.041719f
C880 VTAIL.n107 VSUBS 0.372951f
C881 VTAIL.n108 VSUBS 0.029168f
C882 VTAIL.n109 VSUBS 0.025653f
C883 VTAIL.n110 VSUBS 0.013785f
C884 VTAIL.n111 VSUBS 0.032583f
C885 VTAIL.n112 VSUBS 0.014596f
C886 VTAIL.n113 VSUBS 0.025653f
C887 VTAIL.n114 VSUBS 0.01419f
C888 VTAIL.n115 VSUBS 0.032583f
C889 VTAIL.n116 VSUBS 0.014596f
C890 VTAIL.n117 VSUBS 0.025653f
C891 VTAIL.n118 VSUBS 0.013785f
C892 VTAIL.n119 VSUBS 0.032583f
C893 VTAIL.n120 VSUBS 0.014596f
C894 VTAIL.n121 VSUBS 0.025653f
C895 VTAIL.n122 VSUBS 0.013785f
C896 VTAIL.n123 VSUBS 0.024437f
C897 VTAIL.n124 VSUBS 0.02451f
C898 VTAIL.t4 VSUBS 0.070084f
C899 VTAIL.n125 VSUBS 0.18095f
C900 VTAIL.n126 VSUBS 1.0558f
C901 VTAIL.n127 VSUBS 0.013785f
C902 VTAIL.n128 VSUBS 0.014596f
C903 VTAIL.n129 VSUBS 0.032583f
C904 VTAIL.n130 VSUBS 0.032583f
C905 VTAIL.n131 VSUBS 0.014596f
C906 VTAIL.n132 VSUBS 0.013785f
C907 VTAIL.n133 VSUBS 0.025653f
C908 VTAIL.n134 VSUBS 0.025653f
C909 VTAIL.n135 VSUBS 0.013785f
C910 VTAIL.n136 VSUBS 0.014596f
C911 VTAIL.n137 VSUBS 0.032583f
C912 VTAIL.n138 VSUBS 0.032583f
C913 VTAIL.n139 VSUBS 0.014596f
C914 VTAIL.n140 VSUBS 0.013785f
C915 VTAIL.n141 VSUBS 0.025653f
C916 VTAIL.n142 VSUBS 0.025653f
C917 VTAIL.n143 VSUBS 0.013785f
C918 VTAIL.n144 VSUBS 0.013785f
C919 VTAIL.n145 VSUBS 0.014596f
C920 VTAIL.n146 VSUBS 0.032583f
C921 VTAIL.n147 VSUBS 0.032583f
C922 VTAIL.n148 VSUBS 0.032583f
C923 VTAIL.n149 VSUBS 0.01419f
C924 VTAIL.n150 VSUBS 0.013785f
C925 VTAIL.n151 VSUBS 0.025653f
C926 VTAIL.n152 VSUBS 0.025653f
C927 VTAIL.n153 VSUBS 0.013785f
C928 VTAIL.n154 VSUBS 0.014596f
C929 VTAIL.n155 VSUBS 0.032583f
C930 VTAIL.n156 VSUBS 0.082218f
C931 VTAIL.n157 VSUBS 0.014596f
C932 VTAIL.n158 VSUBS 0.013785f
C933 VTAIL.n159 VSUBS 0.067006f
C934 VTAIL.n160 VSUBS 0.041719f
C935 VTAIL.n161 VSUBS 1.71585f
C936 VTAIL.n162 VSUBS 0.029168f
C937 VTAIL.n163 VSUBS 0.025653f
C938 VTAIL.n164 VSUBS 0.013785f
C939 VTAIL.n165 VSUBS 0.032583f
C940 VTAIL.n166 VSUBS 0.014596f
C941 VTAIL.n167 VSUBS 0.025653f
C942 VTAIL.n168 VSUBS 0.01419f
C943 VTAIL.n169 VSUBS 0.032583f
C944 VTAIL.n170 VSUBS 0.013785f
C945 VTAIL.n171 VSUBS 0.014596f
C946 VTAIL.n172 VSUBS 0.025653f
C947 VTAIL.n173 VSUBS 0.013785f
C948 VTAIL.n174 VSUBS 0.032583f
C949 VTAIL.n175 VSUBS 0.014596f
C950 VTAIL.n176 VSUBS 0.025653f
C951 VTAIL.n177 VSUBS 0.013785f
C952 VTAIL.n178 VSUBS 0.024437f
C953 VTAIL.n179 VSUBS 0.02451f
C954 VTAIL.t7 VSUBS 0.070084f
C955 VTAIL.n180 VSUBS 0.18095f
C956 VTAIL.n181 VSUBS 1.0558f
C957 VTAIL.n182 VSUBS 0.013785f
C958 VTAIL.n183 VSUBS 0.014596f
C959 VTAIL.n184 VSUBS 0.032583f
C960 VTAIL.n185 VSUBS 0.032583f
C961 VTAIL.n186 VSUBS 0.014596f
C962 VTAIL.n187 VSUBS 0.013785f
C963 VTAIL.n188 VSUBS 0.025653f
C964 VTAIL.n189 VSUBS 0.025653f
C965 VTAIL.n190 VSUBS 0.013785f
C966 VTAIL.n191 VSUBS 0.014596f
C967 VTAIL.n192 VSUBS 0.032583f
C968 VTAIL.n193 VSUBS 0.032583f
C969 VTAIL.n194 VSUBS 0.014596f
C970 VTAIL.n195 VSUBS 0.013785f
C971 VTAIL.n196 VSUBS 0.025653f
C972 VTAIL.n197 VSUBS 0.025653f
C973 VTAIL.n198 VSUBS 0.013785f
C974 VTAIL.n199 VSUBS 0.014596f
C975 VTAIL.n200 VSUBS 0.032583f
C976 VTAIL.n201 VSUBS 0.032583f
C977 VTAIL.n202 VSUBS 0.032583f
C978 VTAIL.n203 VSUBS 0.01419f
C979 VTAIL.n204 VSUBS 0.013785f
C980 VTAIL.n205 VSUBS 0.025653f
C981 VTAIL.n206 VSUBS 0.025653f
C982 VTAIL.n207 VSUBS 0.013785f
C983 VTAIL.n208 VSUBS 0.014596f
C984 VTAIL.n209 VSUBS 0.032583f
C985 VTAIL.n210 VSUBS 0.082218f
C986 VTAIL.n211 VSUBS 0.014596f
C987 VTAIL.n212 VSUBS 0.013785f
C988 VTAIL.n213 VSUBS 0.067006f
C989 VTAIL.n214 VSUBS 0.041719f
C990 VTAIL.n215 VSUBS 1.71585f
C991 VTAIL.n216 VSUBS 0.029168f
C992 VTAIL.n217 VSUBS 0.025653f
C993 VTAIL.n218 VSUBS 0.013785f
C994 VTAIL.n219 VSUBS 0.032583f
C995 VTAIL.n220 VSUBS 0.014596f
C996 VTAIL.n221 VSUBS 0.025653f
C997 VTAIL.n222 VSUBS 0.01419f
C998 VTAIL.n223 VSUBS 0.032583f
C999 VTAIL.n224 VSUBS 0.013785f
C1000 VTAIL.n225 VSUBS 0.014596f
C1001 VTAIL.n226 VSUBS 0.025653f
C1002 VTAIL.n227 VSUBS 0.013785f
C1003 VTAIL.n228 VSUBS 0.032583f
C1004 VTAIL.n229 VSUBS 0.014596f
C1005 VTAIL.n230 VSUBS 0.025653f
C1006 VTAIL.n231 VSUBS 0.013785f
C1007 VTAIL.n232 VSUBS 0.024437f
C1008 VTAIL.n233 VSUBS 0.02451f
C1009 VTAIL.t1 VSUBS 0.070084f
C1010 VTAIL.n234 VSUBS 0.18095f
C1011 VTAIL.n235 VSUBS 1.0558f
C1012 VTAIL.n236 VSUBS 0.013785f
C1013 VTAIL.n237 VSUBS 0.014596f
C1014 VTAIL.n238 VSUBS 0.032583f
C1015 VTAIL.n239 VSUBS 0.032583f
C1016 VTAIL.n240 VSUBS 0.014596f
C1017 VTAIL.n241 VSUBS 0.013785f
C1018 VTAIL.n242 VSUBS 0.025653f
C1019 VTAIL.n243 VSUBS 0.025653f
C1020 VTAIL.n244 VSUBS 0.013785f
C1021 VTAIL.n245 VSUBS 0.014596f
C1022 VTAIL.n246 VSUBS 0.032583f
C1023 VTAIL.n247 VSUBS 0.032583f
C1024 VTAIL.n248 VSUBS 0.014596f
C1025 VTAIL.n249 VSUBS 0.013785f
C1026 VTAIL.n250 VSUBS 0.025653f
C1027 VTAIL.n251 VSUBS 0.025653f
C1028 VTAIL.n252 VSUBS 0.013785f
C1029 VTAIL.n253 VSUBS 0.014596f
C1030 VTAIL.n254 VSUBS 0.032583f
C1031 VTAIL.n255 VSUBS 0.032583f
C1032 VTAIL.n256 VSUBS 0.032583f
C1033 VTAIL.n257 VSUBS 0.01419f
C1034 VTAIL.n258 VSUBS 0.013785f
C1035 VTAIL.n259 VSUBS 0.025653f
C1036 VTAIL.n260 VSUBS 0.025653f
C1037 VTAIL.n261 VSUBS 0.013785f
C1038 VTAIL.n262 VSUBS 0.014596f
C1039 VTAIL.n263 VSUBS 0.032583f
C1040 VTAIL.n264 VSUBS 0.082218f
C1041 VTAIL.n265 VSUBS 0.014596f
C1042 VTAIL.n266 VSUBS 0.013785f
C1043 VTAIL.n267 VSUBS 0.067006f
C1044 VTAIL.n268 VSUBS 0.041719f
C1045 VTAIL.n269 VSUBS 0.372951f
C1046 VTAIL.n270 VSUBS 0.029168f
C1047 VTAIL.n271 VSUBS 0.025653f
C1048 VTAIL.n272 VSUBS 0.013785f
C1049 VTAIL.n273 VSUBS 0.032583f
C1050 VTAIL.n274 VSUBS 0.014596f
C1051 VTAIL.n275 VSUBS 0.025653f
C1052 VTAIL.n276 VSUBS 0.01419f
C1053 VTAIL.n277 VSUBS 0.032583f
C1054 VTAIL.n278 VSUBS 0.013785f
C1055 VTAIL.n279 VSUBS 0.014596f
C1056 VTAIL.n280 VSUBS 0.025653f
C1057 VTAIL.n281 VSUBS 0.013785f
C1058 VTAIL.n282 VSUBS 0.032583f
C1059 VTAIL.n283 VSUBS 0.014596f
C1060 VTAIL.n284 VSUBS 0.025653f
C1061 VTAIL.n285 VSUBS 0.013785f
C1062 VTAIL.n286 VSUBS 0.024437f
C1063 VTAIL.n287 VSUBS 0.02451f
C1064 VTAIL.t5 VSUBS 0.070084f
C1065 VTAIL.n288 VSUBS 0.18095f
C1066 VTAIL.n289 VSUBS 1.0558f
C1067 VTAIL.n290 VSUBS 0.013785f
C1068 VTAIL.n291 VSUBS 0.014596f
C1069 VTAIL.n292 VSUBS 0.032583f
C1070 VTAIL.n293 VSUBS 0.032583f
C1071 VTAIL.n294 VSUBS 0.014596f
C1072 VTAIL.n295 VSUBS 0.013785f
C1073 VTAIL.n296 VSUBS 0.025653f
C1074 VTAIL.n297 VSUBS 0.025653f
C1075 VTAIL.n298 VSUBS 0.013785f
C1076 VTAIL.n299 VSUBS 0.014596f
C1077 VTAIL.n300 VSUBS 0.032583f
C1078 VTAIL.n301 VSUBS 0.032583f
C1079 VTAIL.n302 VSUBS 0.014596f
C1080 VTAIL.n303 VSUBS 0.013785f
C1081 VTAIL.n304 VSUBS 0.025653f
C1082 VTAIL.n305 VSUBS 0.025653f
C1083 VTAIL.n306 VSUBS 0.013785f
C1084 VTAIL.n307 VSUBS 0.014596f
C1085 VTAIL.n308 VSUBS 0.032583f
C1086 VTAIL.n309 VSUBS 0.032583f
C1087 VTAIL.n310 VSUBS 0.032583f
C1088 VTAIL.n311 VSUBS 0.01419f
C1089 VTAIL.n312 VSUBS 0.013785f
C1090 VTAIL.n313 VSUBS 0.025653f
C1091 VTAIL.n314 VSUBS 0.025653f
C1092 VTAIL.n315 VSUBS 0.013785f
C1093 VTAIL.n316 VSUBS 0.014596f
C1094 VTAIL.n317 VSUBS 0.032583f
C1095 VTAIL.n318 VSUBS 0.082218f
C1096 VTAIL.n319 VSUBS 0.014596f
C1097 VTAIL.n320 VSUBS 0.013785f
C1098 VTAIL.n321 VSUBS 0.067006f
C1099 VTAIL.n322 VSUBS 0.041719f
C1100 VTAIL.n323 VSUBS 0.372951f
C1101 VTAIL.n324 VSUBS 0.029168f
C1102 VTAIL.n325 VSUBS 0.025653f
C1103 VTAIL.n326 VSUBS 0.013785f
C1104 VTAIL.n327 VSUBS 0.032583f
C1105 VTAIL.n328 VSUBS 0.014596f
C1106 VTAIL.n329 VSUBS 0.025653f
C1107 VTAIL.n330 VSUBS 0.01419f
C1108 VTAIL.n331 VSUBS 0.032583f
C1109 VTAIL.n332 VSUBS 0.013785f
C1110 VTAIL.n333 VSUBS 0.014596f
C1111 VTAIL.n334 VSUBS 0.025653f
C1112 VTAIL.n335 VSUBS 0.013785f
C1113 VTAIL.n336 VSUBS 0.032583f
C1114 VTAIL.n337 VSUBS 0.014596f
C1115 VTAIL.n338 VSUBS 0.025653f
C1116 VTAIL.n339 VSUBS 0.013785f
C1117 VTAIL.n340 VSUBS 0.024437f
C1118 VTAIL.n341 VSUBS 0.02451f
C1119 VTAIL.t3 VSUBS 0.070084f
C1120 VTAIL.n342 VSUBS 0.18095f
C1121 VTAIL.n343 VSUBS 1.0558f
C1122 VTAIL.n344 VSUBS 0.013785f
C1123 VTAIL.n345 VSUBS 0.014596f
C1124 VTAIL.n346 VSUBS 0.032583f
C1125 VTAIL.n347 VSUBS 0.032583f
C1126 VTAIL.n348 VSUBS 0.014596f
C1127 VTAIL.n349 VSUBS 0.013785f
C1128 VTAIL.n350 VSUBS 0.025653f
C1129 VTAIL.n351 VSUBS 0.025653f
C1130 VTAIL.n352 VSUBS 0.013785f
C1131 VTAIL.n353 VSUBS 0.014596f
C1132 VTAIL.n354 VSUBS 0.032583f
C1133 VTAIL.n355 VSUBS 0.032583f
C1134 VTAIL.n356 VSUBS 0.014596f
C1135 VTAIL.n357 VSUBS 0.013785f
C1136 VTAIL.n358 VSUBS 0.025653f
C1137 VTAIL.n359 VSUBS 0.025653f
C1138 VTAIL.n360 VSUBS 0.013785f
C1139 VTAIL.n361 VSUBS 0.014596f
C1140 VTAIL.n362 VSUBS 0.032583f
C1141 VTAIL.n363 VSUBS 0.032583f
C1142 VTAIL.n364 VSUBS 0.032583f
C1143 VTAIL.n365 VSUBS 0.01419f
C1144 VTAIL.n366 VSUBS 0.013785f
C1145 VTAIL.n367 VSUBS 0.025653f
C1146 VTAIL.n368 VSUBS 0.025653f
C1147 VTAIL.n369 VSUBS 0.013785f
C1148 VTAIL.n370 VSUBS 0.014596f
C1149 VTAIL.n371 VSUBS 0.032583f
C1150 VTAIL.n372 VSUBS 0.082218f
C1151 VTAIL.n373 VSUBS 0.014596f
C1152 VTAIL.n374 VSUBS 0.013785f
C1153 VTAIL.n375 VSUBS 0.067006f
C1154 VTAIL.n376 VSUBS 0.041719f
C1155 VTAIL.n377 VSUBS 1.71585f
C1156 VTAIL.n378 VSUBS 0.029168f
C1157 VTAIL.n379 VSUBS 0.025653f
C1158 VTAIL.n380 VSUBS 0.013785f
C1159 VTAIL.n381 VSUBS 0.032583f
C1160 VTAIL.n382 VSUBS 0.014596f
C1161 VTAIL.n383 VSUBS 0.025653f
C1162 VTAIL.n384 VSUBS 0.01419f
C1163 VTAIL.n385 VSUBS 0.032583f
C1164 VTAIL.n386 VSUBS 0.014596f
C1165 VTAIL.n387 VSUBS 0.025653f
C1166 VTAIL.n388 VSUBS 0.013785f
C1167 VTAIL.n389 VSUBS 0.032583f
C1168 VTAIL.n390 VSUBS 0.014596f
C1169 VTAIL.n391 VSUBS 0.025653f
C1170 VTAIL.n392 VSUBS 0.013785f
C1171 VTAIL.n393 VSUBS 0.024437f
C1172 VTAIL.n394 VSUBS 0.02451f
C1173 VTAIL.t0 VSUBS 0.070084f
C1174 VTAIL.n395 VSUBS 0.18095f
C1175 VTAIL.n396 VSUBS 1.0558f
C1176 VTAIL.n397 VSUBS 0.013785f
C1177 VTAIL.n398 VSUBS 0.014596f
C1178 VTAIL.n399 VSUBS 0.032583f
C1179 VTAIL.n400 VSUBS 0.032583f
C1180 VTAIL.n401 VSUBS 0.014596f
C1181 VTAIL.n402 VSUBS 0.013785f
C1182 VTAIL.n403 VSUBS 0.025653f
C1183 VTAIL.n404 VSUBS 0.025653f
C1184 VTAIL.n405 VSUBS 0.013785f
C1185 VTAIL.n406 VSUBS 0.014596f
C1186 VTAIL.n407 VSUBS 0.032583f
C1187 VTAIL.n408 VSUBS 0.032583f
C1188 VTAIL.n409 VSUBS 0.014596f
C1189 VTAIL.n410 VSUBS 0.013785f
C1190 VTAIL.n411 VSUBS 0.025653f
C1191 VTAIL.n412 VSUBS 0.025653f
C1192 VTAIL.n413 VSUBS 0.013785f
C1193 VTAIL.n414 VSUBS 0.013785f
C1194 VTAIL.n415 VSUBS 0.014596f
C1195 VTAIL.n416 VSUBS 0.032583f
C1196 VTAIL.n417 VSUBS 0.032583f
C1197 VTAIL.n418 VSUBS 0.032583f
C1198 VTAIL.n419 VSUBS 0.01419f
C1199 VTAIL.n420 VSUBS 0.013785f
C1200 VTAIL.n421 VSUBS 0.025653f
C1201 VTAIL.n422 VSUBS 0.025653f
C1202 VTAIL.n423 VSUBS 0.013785f
C1203 VTAIL.n424 VSUBS 0.014596f
C1204 VTAIL.n425 VSUBS 0.032583f
C1205 VTAIL.n426 VSUBS 0.082218f
C1206 VTAIL.n427 VSUBS 0.014596f
C1207 VTAIL.n428 VSUBS 0.013785f
C1208 VTAIL.n429 VSUBS 0.067006f
C1209 VTAIL.n430 VSUBS 0.041719f
C1210 VTAIL.n431 VSUBS 1.55712f
C1211 VP.n0 VSUBS 0.059593f
C1212 VP.t0 VSUBS 3.48925f
C1213 VP.n1 VSUBS 0.058767f
C1214 VP.n2 VSUBS 0.031691f
C1215 VP.n3 VSUBS 0.058767f
C1216 VP.t1 VSUBS 3.99881f
C1217 VP.t2 VSUBS 4.02041f
C1218 VP.n4 VSUBS 4.41153f
C1219 VP.n5 VSUBS 1.91187f
C1220 VP.t3 VSUBS 3.48925f
C1221 VP.n6 VSUBS 1.3696f
C1222 VP.n7 VSUBS 0.053545f
C1223 VP.n8 VSUBS 0.059593f
C1224 VP.n9 VSUBS 0.031691f
C1225 VP.n10 VSUBS 0.031691f
C1226 VP.n11 VSUBS 0.058767f
C1227 VP.n12 VSUBS 0.046067f
C1228 VP.n13 VSUBS 0.046067f
C1229 VP.n14 VSUBS 0.031691f
C1230 VP.n15 VSUBS 0.031691f
C1231 VP.n16 VSUBS 0.031691f
C1232 VP.n17 VSUBS 0.058767f
C1233 VP.n18 VSUBS 0.053545f
C1234 VP.n19 VSUBS 1.3696f
C1235 VP.n20 VSUBS 0.101432f
.ends

