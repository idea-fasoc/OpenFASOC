* NGSPICE file created from diff_pair_sample_0309.ext - technology: sky130A

.subckt diff_pair_sample_0309 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=7.4997 pd=39.24 as=0 ps=0 w=19.23 l=0.35
X1 VDD1.t7 VP.t0 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=7.4997 ps=39.24 w=19.23 l=0.35
X2 VDD1.t6 VP.t1 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=3.17295 ps=19.56 w=19.23 l=0.35
X3 VTAIL.t1 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=7.4997 pd=39.24 as=3.17295 ps=19.56 w=19.23 l=0.35
X4 VDD1.t5 VP.t2 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=7.4997 ps=39.24 w=19.23 l=0.35
X5 VTAIL.t8 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4997 pd=39.24 as=3.17295 ps=19.56 w=19.23 l=0.35
X6 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=7.4997 pd=39.24 as=0 ps=0 w=19.23 l=0.35
X7 VDD2.t6 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=7.4997 ps=39.24 w=19.23 l=0.35
X8 VTAIL.t2 VN.t2 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=3.17295 ps=19.56 w=19.23 l=0.35
X9 VDD2.t4 VN.t3 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=7.4997 ps=39.24 w=19.23 l=0.35
X10 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.4997 pd=39.24 as=0 ps=0 w=19.23 l=0.35
X11 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.4997 pd=39.24 as=0 ps=0 w=19.23 l=0.35
X12 VTAIL.t6 VN.t4 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=7.4997 pd=39.24 as=3.17295 ps=19.56 w=19.23 l=0.35
X13 VDD2.t2 VN.t5 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=3.17295 ps=19.56 w=19.23 l=0.35
X14 VDD2.t1 VN.t6 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=3.17295 ps=19.56 w=19.23 l=0.35
X15 VTAIL.t14 VP.t4 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=3.17295 ps=19.56 w=19.23 l=0.35
X16 VTAIL.t10 VP.t5 VDD1.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=3.17295 ps=19.56 w=19.23 l=0.35
X17 VTAIL.t5 VN.t7 VDD2.t0 B.t6 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=3.17295 ps=19.56 w=19.23 l=0.35
X18 VDD1.t1 VP.t6 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=3.17295 pd=19.56 as=3.17295 ps=19.56 w=19.23 l=0.35
X19 VTAIL.t12 VP.t7 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=7.4997 pd=39.24 as=3.17295 ps=19.56 w=19.23 l=0.35
R0 B.n181 B.t19 1535.69
R1 B.n175 B.t15 1535.69
R2 B.n70 B.t12 1535.69
R3 B.n77 B.t8 1535.69
R4 B.n564 B.n563 585
R5 B.n564 B.n36 585
R6 B.n567 B.n566 585
R7 B.n568 B.n108 585
R8 B.n570 B.n569 585
R9 B.n572 B.n107 585
R10 B.n575 B.n574 585
R11 B.n576 B.n106 585
R12 B.n578 B.n577 585
R13 B.n580 B.n105 585
R14 B.n583 B.n582 585
R15 B.n584 B.n104 585
R16 B.n586 B.n585 585
R17 B.n588 B.n103 585
R18 B.n591 B.n590 585
R19 B.n592 B.n102 585
R20 B.n594 B.n593 585
R21 B.n596 B.n101 585
R22 B.n599 B.n598 585
R23 B.n600 B.n100 585
R24 B.n602 B.n601 585
R25 B.n604 B.n99 585
R26 B.n607 B.n606 585
R27 B.n608 B.n98 585
R28 B.n610 B.n609 585
R29 B.n612 B.n97 585
R30 B.n615 B.n614 585
R31 B.n616 B.n96 585
R32 B.n618 B.n617 585
R33 B.n620 B.n95 585
R34 B.n623 B.n622 585
R35 B.n624 B.n94 585
R36 B.n626 B.n625 585
R37 B.n628 B.n93 585
R38 B.n631 B.n630 585
R39 B.n632 B.n92 585
R40 B.n634 B.n633 585
R41 B.n636 B.n91 585
R42 B.n639 B.n638 585
R43 B.n640 B.n90 585
R44 B.n642 B.n641 585
R45 B.n644 B.n89 585
R46 B.n647 B.n646 585
R47 B.n648 B.n88 585
R48 B.n650 B.n649 585
R49 B.n652 B.n87 585
R50 B.n655 B.n654 585
R51 B.n656 B.n86 585
R52 B.n658 B.n657 585
R53 B.n660 B.n85 585
R54 B.n663 B.n662 585
R55 B.n664 B.n84 585
R56 B.n666 B.n665 585
R57 B.n668 B.n83 585
R58 B.n671 B.n670 585
R59 B.n672 B.n82 585
R60 B.n674 B.n673 585
R61 B.n676 B.n81 585
R62 B.n679 B.n678 585
R63 B.n680 B.n80 585
R64 B.n682 B.n681 585
R65 B.n684 B.n79 585
R66 B.n687 B.n686 585
R67 B.n688 B.n76 585
R68 B.n691 B.n690 585
R69 B.n693 B.n75 585
R70 B.n696 B.n695 585
R71 B.n697 B.n74 585
R72 B.n699 B.n698 585
R73 B.n701 B.n73 585
R74 B.n704 B.n703 585
R75 B.n705 B.n69 585
R76 B.n707 B.n706 585
R77 B.n709 B.n68 585
R78 B.n712 B.n711 585
R79 B.n713 B.n67 585
R80 B.n715 B.n714 585
R81 B.n717 B.n66 585
R82 B.n720 B.n719 585
R83 B.n721 B.n65 585
R84 B.n723 B.n722 585
R85 B.n725 B.n64 585
R86 B.n728 B.n727 585
R87 B.n729 B.n63 585
R88 B.n731 B.n730 585
R89 B.n733 B.n62 585
R90 B.n736 B.n735 585
R91 B.n737 B.n61 585
R92 B.n739 B.n738 585
R93 B.n741 B.n60 585
R94 B.n744 B.n743 585
R95 B.n745 B.n59 585
R96 B.n747 B.n746 585
R97 B.n749 B.n58 585
R98 B.n752 B.n751 585
R99 B.n753 B.n57 585
R100 B.n755 B.n754 585
R101 B.n757 B.n56 585
R102 B.n760 B.n759 585
R103 B.n761 B.n55 585
R104 B.n763 B.n762 585
R105 B.n765 B.n54 585
R106 B.n768 B.n767 585
R107 B.n769 B.n53 585
R108 B.n771 B.n770 585
R109 B.n773 B.n52 585
R110 B.n776 B.n775 585
R111 B.n777 B.n51 585
R112 B.n779 B.n778 585
R113 B.n781 B.n50 585
R114 B.n784 B.n783 585
R115 B.n785 B.n49 585
R116 B.n787 B.n786 585
R117 B.n789 B.n48 585
R118 B.n792 B.n791 585
R119 B.n793 B.n47 585
R120 B.n795 B.n794 585
R121 B.n797 B.n46 585
R122 B.n800 B.n799 585
R123 B.n801 B.n45 585
R124 B.n803 B.n802 585
R125 B.n805 B.n44 585
R126 B.n808 B.n807 585
R127 B.n809 B.n43 585
R128 B.n811 B.n810 585
R129 B.n813 B.n42 585
R130 B.n816 B.n815 585
R131 B.n817 B.n41 585
R132 B.n819 B.n818 585
R133 B.n821 B.n40 585
R134 B.n824 B.n823 585
R135 B.n825 B.n39 585
R136 B.n827 B.n826 585
R137 B.n829 B.n38 585
R138 B.n832 B.n831 585
R139 B.n833 B.n37 585
R140 B.n562 B.n35 585
R141 B.n836 B.n35 585
R142 B.n561 B.n34 585
R143 B.n837 B.n34 585
R144 B.n560 B.n33 585
R145 B.n838 B.n33 585
R146 B.n559 B.n558 585
R147 B.n558 B.n29 585
R148 B.n557 B.n28 585
R149 B.n844 B.n28 585
R150 B.n556 B.n27 585
R151 B.n845 B.n27 585
R152 B.n555 B.n26 585
R153 B.n846 B.n26 585
R154 B.n554 B.n553 585
R155 B.n553 B.n22 585
R156 B.n552 B.n21 585
R157 B.n852 B.n21 585
R158 B.n551 B.n20 585
R159 B.n853 B.n20 585
R160 B.n550 B.n19 585
R161 B.n854 B.n19 585
R162 B.n549 B.n548 585
R163 B.n548 B.n18 585
R164 B.n547 B.n14 585
R165 B.n860 B.n14 585
R166 B.n546 B.n13 585
R167 B.n861 B.n13 585
R168 B.n545 B.n12 585
R169 B.n862 B.n12 585
R170 B.n544 B.n543 585
R171 B.n543 B.n11 585
R172 B.n542 B.n7 585
R173 B.n868 B.n7 585
R174 B.n541 B.n6 585
R175 B.n869 B.n6 585
R176 B.n540 B.n5 585
R177 B.n870 B.n5 585
R178 B.n539 B.n538 585
R179 B.n538 B.n4 585
R180 B.n537 B.n109 585
R181 B.n537 B.n536 585
R182 B.n526 B.n110 585
R183 B.n529 B.n110 585
R184 B.n528 B.n527 585
R185 B.n530 B.n528 585
R186 B.n525 B.n114 585
R187 B.n117 B.n114 585
R188 B.n524 B.n523 585
R189 B.n523 B.n522 585
R190 B.n116 B.n115 585
R191 B.n515 B.n116 585
R192 B.n514 B.n513 585
R193 B.n516 B.n514 585
R194 B.n512 B.n121 585
R195 B.n125 B.n121 585
R196 B.n511 B.n510 585
R197 B.n510 B.n509 585
R198 B.n123 B.n122 585
R199 B.n124 B.n123 585
R200 B.n502 B.n501 585
R201 B.n503 B.n502 585
R202 B.n500 B.n130 585
R203 B.n130 B.n129 585
R204 B.n499 B.n498 585
R205 B.n498 B.n497 585
R206 B.n132 B.n131 585
R207 B.n133 B.n132 585
R208 B.n490 B.n489 585
R209 B.n491 B.n490 585
R210 B.n488 B.n138 585
R211 B.n138 B.n137 585
R212 B.n487 B.n486 585
R213 B.n486 B.n485 585
R214 B.n482 B.n142 585
R215 B.n481 B.n480 585
R216 B.n478 B.n143 585
R217 B.n478 B.n141 585
R218 B.n477 B.n476 585
R219 B.n475 B.n474 585
R220 B.n473 B.n145 585
R221 B.n471 B.n470 585
R222 B.n469 B.n146 585
R223 B.n468 B.n467 585
R224 B.n465 B.n147 585
R225 B.n463 B.n462 585
R226 B.n461 B.n148 585
R227 B.n460 B.n459 585
R228 B.n457 B.n149 585
R229 B.n455 B.n454 585
R230 B.n453 B.n150 585
R231 B.n452 B.n451 585
R232 B.n449 B.n151 585
R233 B.n447 B.n446 585
R234 B.n445 B.n152 585
R235 B.n444 B.n443 585
R236 B.n441 B.n153 585
R237 B.n439 B.n438 585
R238 B.n437 B.n154 585
R239 B.n436 B.n435 585
R240 B.n433 B.n155 585
R241 B.n431 B.n430 585
R242 B.n429 B.n156 585
R243 B.n428 B.n427 585
R244 B.n425 B.n157 585
R245 B.n423 B.n422 585
R246 B.n421 B.n158 585
R247 B.n420 B.n419 585
R248 B.n417 B.n159 585
R249 B.n415 B.n414 585
R250 B.n413 B.n160 585
R251 B.n412 B.n411 585
R252 B.n409 B.n161 585
R253 B.n407 B.n406 585
R254 B.n405 B.n162 585
R255 B.n404 B.n403 585
R256 B.n401 B.n163 585
R257 B.n399 B.n398 585
R258 B.n397 B.n164 585
R259 B.n396 B.n395 585
R260 B.n393 B.n165 585
R261 B.n391 B.n390 585
R262 B.n389 B.n166 585
R263 B.n388 B.n387 585
R264 B.n385 B.n167 585
R265 B.n383 B.n382 585
R266 B.n381 B.n168 585
R267 B.n380 B.n379 585
R268 B.n377 B.n169 585
R269 B.n375 B.n374 585
R270 B.n373 B.n170 585
R271 B.n372 B.n371 585
R272 B.n369 B.n171 585
R273 B.n367 B.n366 585
R274 B.n365 B.n172 585
R275 B.n364 B.n363 585
R276 B.n361 B.n173 585
R277 B.n359 B.n358 585
R278 B.n356 B.n174 585
R279 B.n355 B.n354 585
R280 B.n352 B.n177 585
R281 B.n350 B.n349 585
R282 B.n348 B.n178 585
R283 B.n347 B.n346 585
R284 B.n344 B.n179 585
R285 B.n342 B.n341 585
R286 B.n340 B.n180 585
R287 B.n338 B.n337 585
R288 B.n335 B.n183 585
R289 B.n333 B.n332 585
R290 B.n331 B.n184 585
R291 B.n330 B.n329 585
R292 B.n327 B.n185 585
R293 B.n325 B.n324 585
R294 B.n323 B.n186 585
R295 B.n322 B.n321 585
R296 B.n319 B.n187 585
R297 B.n317 B.n316 585
R298 B.n315 B.n188 585
R299 B.n314 B.n313 585
R300 B.n311 B.n189 585
R301 B.n309 B.n308 585
R302 B.n307 B.n190 585
R303 B.n306 B.n305 585
R304 B.n303 B.n191 585
R305 B.n301 B.n300 585
R306 B.n299 B.n192 585
R307 B.n298 B.n297 585
R308 B.n295 B.n193 585
R309 B.n293 B.n292 585
R310 B.n291 B.n194 585
R311 B.n290 B.n289 585
R312 B.n287 B.n195 585
R313 B.n285 B.n284 585
R314 B.n283 B.n196 585
R315 B.n282 B.n281 585
R316 B.n279 B.n197 585
R317 B.n277 B.n276 585
R318 B.n275 B.n198 585
R319 B.n274 B.n273 585
R320 B.n271 B.n199 585
R321 B.n269 B.n268 585
R322 B.n267 B.n200 585
R323 B.n266 B.n265 585
R324 B.n263 B.n201 585
R325 B.n261 B.n260 585
R326 B.n259 B.n202 585
R327 B.n258 B.n257 585
R328 B.n255 B.n203 585
R329 B.n253 B.n252 585
R330 B.n251 B.n204 585
R331 B.n250 B.n249 585
R332 B.n247 B.n205 585
R333 B.n245 B.n244 585
R334 B.n243 B.n206 585
R335 B.n242 B.n241 585
R336 B.n239 B.n207 585
R337 B.n237 B.n236 585
R338 B.n235 B.n208 585
R339 B.n234 B.n233 585
R340 B.n231 B.n209 585
R341 B.n229 B.n228 585
R342 B.n227 B.n210 585
R343 B.n226 B.n225 585
R344 B.n223 B.n211 585
R345 B.n221 B.n220 585
R346 B.n219 B.n212 585
R347 B.n218 B.n217 585
R348 B.n215 B.n213 585
R349 B.n140 B.n139 585
R350 B.n484 B.n483 585
R351 B.n485 B.n484 585
R352 B.n136 B.n135 585
R353 B.n137 B.n136 585
R354 B.n493 B.n492 585
R355 B.n492 B.n491 585
R356 B.n494 B.n134 585
R357 B.n134 B.n133 585
R358 B.n496 B.n495 585
R359 B.n497 B.n496 585
R360 B.n128 B.n127 585
R361 B.n129 B.n128 585
R362 B.n505 B.n504 585
R363 B.n504 B.n503 585
R364 B.n506 B.n126 585
R365 B.n126 B.n124 585
R366 B.n508 B.n507 585
R367 B.n509 B.n508 585
R368 B.n120 B.n119 585
R369 B.n125 B.n120 585
R370 B.n518 B.n517 585
R371 B.n517 B.n516 585
R372 B.n519 B.n118 585
R373 B.n515 B.n118 585
R374 B.n521 B.n520 585
R375 B.n522 B.n521 585
R376 B.n113 B.n112 585
R377 B.n117 B.n113 585
R378 B.n532 B.n531 585
R379 B.n531 B.n530 585
R380 B.n533 B.n111 585
R381 B.n529 B.n111 585
R382 B.n535 B.n534 585
R383 B.n536 B.n535 585
R384 B.n2 B.n0 585
R385 B.n4 B.n2 585
R386 B.n3 B.n1 585
R387 B.n869 B.n3 585
R388 B.n867 B.n866 585
R389 B.n868 B.n867 585
R390 B.n865 B.n8 585
R391 B.n11 B.n8 585
R392 B.n864 B.n863 585
R393 B.n863 B.n862 585
R394 B.n10 B.n9 585
R395 B.n861 B.n10 585
R396 B.n859 B.n858 585
R397 B.n860 B.n859 585
R398 B.n857 B.n15 585
R399 B.n18 B.n15 585
R400 B.n856 B.n855 585
R401 B.n855 B.n854 585
R402 B.n17 B.n16 585
R403 B.n853 B.n17 585
R404 B.n851 B.n850 585
R405 B.n852 B.n851 585
R406 B.n849 B.n23 585
R407 B.n23 B.n22 585
R408 B.n848 B.n847 585
R409 B.n847 B.n846 585
R410 B.n25 B.n24 585
R411 B.n845 B.n25 585
R412 B.n843 B.n842 585
R413 B.n844 B.n843 585
R414 B.n841 B.n30 585
R415 B.n30 B.n29 585
R416 B.n840 B.n839 585
R417 B.n839 B.n838 585
R418 B.n32 B.n31 585
R419 B.n837 B.n32 585
R420 B.n835 B.n834 585
R421 B.n836 B.n835 585
R422 B.n872 B.n871 585
R423 B.n871 B.n870 585
R424 B.n484 B.n142 545.355
R425 B.n835 B.n37 545.355
R426 B.n486 B.n140 545.355
R427 B.n564 B.n35 545.355
R428 B.n565 B.n36 256.663
R429 B.n571 B.n36 256.663
R430 B.n573 B.n36 256.663
R431 B.n579 B.n36 256.663
R432 B.n581 B.n36 256.663
R433 B.n587 B.n36 256.663
R434 B.n589 B.n36 256.663
R435 B.n595 B.n36 256.663
R436 B.n597 B.n36 256.663
R437 B.n603 B.n36 256.663
R438 B.n605 B.n36 256.663
R439 B.n611 B.n36 256.663
R440 B.n613 B.n36 256.663
R441 B.n619 B.n36 256.663
R442 B.n621 B.n36 256.663
R443 B.n627 B.n36 256.663
R444 B.n629 B.n36 256.663
R445 B.n635 B.n36 256.663
R446 B.n637 B.n36 256.663
R447 B.n643 B.n36 256.663
R448 B.n645 B.n36 256.663
R449 B.n651 B.n36 256.663
R450 B.n653 B.n36 256.663
R451 B.n659 B.n36 256.663
R452 B.n661 B.n36 256.663
R453 B.n667 B.n36 256.663
R454 B.n669 B.n36 256.663
R455 B.n675 B.n36 256.663
R456 B.n677 B.n36 256.663
R457 B.n683 B.n36 256.663
R458 B.n685 B.n36 256.663
R459 B.n692 B.n36 256.663
R460 B.n694 B.n36 256.663
R461 B.n700 B.n36 256.663
R462 B.n702 B.n36 256.663
R463 B.n708 B.n36 256.663
R464 B.n710 B.n36 256.663
R465 B.n716 B.n36 256.663
R466 B.n718 B.n36 256.663
R467 B.n724 B.n36 256.663
R468 B.n726 B.n36 256.663
R469 B.n732 B.n36 256.663
R470 B.n734 B.n36 256.663
R471 B.n740 B.n36 256.663
R472 B.n742 B.n36 256.663
R473 B.n748 B.n36 256.663
R474 B.n750 B.n36 256.663
R475 B.n756 B.n36 256.663
R476 B.n758 B.n36 256.663
R477 B.n764 B.n36 256.663
R478 B.n766 B.n36 256.663
R479 B.n772 B.n36 256.663
R480 B.n774 B.n36 256.663
R481 B.n780 B.n36 256.663
R482 B.n782 B.n36 256.663
R483 B.n788 B.n36 256.663
R484 B.n790 B.n36 256.663
R485 B.n796 B.n36 256.663
R486 B.n798 B.n36 256.663
R487 B.n804 B.n36 256.663
R488 B.n806 B.n36 256.663
R489 B.n812 B.n36 256.663
R490 B.n814 B.n36 256.663
R491 B.n820 B.n36 256.663
R492 B.n822 B.n36 256.663
R493 B.n828 B.n36 256.663
R494 B.n830 B.n36 256.663
R495 B.n479 B.n141 256.663
R496 B.n144 B.n141 256.663
R497 B.n472 B.n141 256.663
R498 B.n466 B.n141 256.663
R499 B.n464 B.n141 256.663
R500 B.n458 B.n141 256.663
R501 B.n456 B.n141 256.663
R502 B.n450 B.n141 256.663
R503 B.n448 B.n141 256.663
R504 B.n442 B.n141 256.663
R505 B.n440 B.n141 256.663
R506 B.n434 B.n141 256.663
R507 B.n432 B.n141 256.663
R508 B.n426 B.n141 256.663
R509 B.n424 B.n141 256.663
R510 B.n418 B.n141 256.663
R511 B.n416 B.n141 256.663
R512 B.n410 B.n141 256.663
R513 B.n408 B.n141 256.663
R514 B.n402 B.n141 256.663
R515 B.n400 B.n141 256.663
R516 B.n394 B.n141 256.663
R517 B.n392 B.n141 256.663
R518 B.n386 B.n141 256.663
R519 B.n384 B.n141 256.663
R520 B.n378 B.n141 256.663
R521 B.n376 B.n141 256.663
R522 B.n370 B.n141 256.663
R523 B.n368 B.n141 256.663
R524 B.n362 B.n141 256.663
R525 B.n360 B.n141 256.663
R526 B.n353 B.n141 256.663
R527 B.n351 B.n141 256.663
R528 B.n345 B.n141 256.663
R529 B.n343 B.n141 256.663
R530 B.n336 B.n141 256.663
R531 B.n334 B.n141 256.663
R532 B.n328 B.n141 256.663
R533 B.n326 B.n141 256.663
R534 B.n320 B.n141 256.663
R535 B.n318 B.n141 256.663
R536 B.n312 B.n141 256.663
R537 B.n310 B.n141 256.663
R538 B.n304 B.n141 256.663
R539 B.n302 B.n141 256.663
R540 B.n296 B.n141 256.663
R541 B.n294 B.n141 256.663
R542 B.n288 B.n141 256.663
R543 B.n286 B.n141 256.663
R544 B.n280 B.n141 256.663
R545 B.n278 B.n141 256.663
R546 B.n272 B.n141 256.663
R547 B.n270 B.n141 256.663
R548 B.n264 B.n141 256.663
R549 B.n262 B.n141 256.663
R550 B.n256 B.n141 256.663
R551 B.n254 B.n141 256.663
R552 B.n248 B.n141 256.663
R553 B.n246 B.n141 256.663
R554 B.n240 B.n141 256.663
R555 B.n238 B.n141 256.663
R556 B.n232 B.n141 256.663
R557 B.n230 B.n141 256.663
R558 B.n224 B.n141 256.663
R559 B.n222 B.n141 256.663
R560 B.n216 B.n141 256.663
R561 B.n214 B.n141 256.663
R562 B.n484 B.n136 163.367
R563 B.n492 B.n136 163.367
R564 B.n492 B.n134 163.367
R565 B.n496 B.n134 163.367
R566 B.n496 B.n128 163.367
R567 B.n504 B.n128 163.367
R568 B.n504 B.n126 163.367
R569 B.n508 B.n126 163.367
R570 B.n508 B.n120 163.367
R571 B.n517 B.n120 163.367
R572 B.n517 B.n118 163.367
R573 B.n521 B.n118 163.367
R574 B.n521 B.n113 163.367
R575 B.n531 B.n113 163.367
R576 B.n531 B.n111 163.367
R577 B.n535 B.n111 163.367
R578 B.n535 B.n2 163.367
R579 B.n871 B.n2 163.367
R580 B.n871 B.n3 163.367
R581 B.n867 B.n3 163.367
R582 B.n867 B.n8 163.367
R583 B.n863 B.n8 163.367
R584 B.n863 B.n10 163.367
R585 B.n859 B.n10 163.367
R586 B.n859 B.n15 163.367
R587 B.n855 B.n15 163.367
R588 B.n855 B.n17 163.367
R589 B.n851 B.n17 163.367
R590 B.n851 B.n23 163.367
R591 B.n847 B.n23 163.367
R592 B.n847 B.n25 163.367
R593 B.n843 B.n25 163.367
R594 B.n843 B.n30 163.367
R595 B.n839 B.n30 163.367
R596 B.n839 B.n32 163.367
R597 B.n835 B.n32 163.367
R598 B.n480 B.n478 163.367
R599 B.n478 B.n477 163.367
R600 B.n474 B.n473 163.367
R601 B.n471 B.n146 163.367
R602 B.n467 B.n465 163.367
R603 B.n463 B.n148 163.367
R604 B.n459 B.n457 163.367
R605 B.n455 B.n150 163.367
R606 B.n451 B.n449 163.367
R607 B.n447 B.n152 163.367
R608 B.n443 B.n441 163.367
R609 B.n439 B.n154 163.367
R610 B.n435 B.n433 163.367
R611 B.n431 B.n156 163.367
R612 B.n427 B.n425 163.367
R613 B.n423 B.n158 163.367
R614 B.n419 B.n417 163.367
R615 B.n415 B.n160 163.367
R616 B.n411 B.n409 163.367
R617 B.n407 B.n162 163.367
R618 B.n403 B.n401 163.367
R619 B.n399 B.n164 163.367
R620 B.n395 B.n393 163.367
R621 B.n391 B.n166 163.367
R622 B.n387 B.n385 163.367
R623 B.n383 B.n168 163.367
R624 B.n379 B.n377 163.367
R625 B.n375 B.n170 163.367
R626 B.n371 B.n369 163.367
R627 B.n367 B.n172 163.367
R628 B.n363 B.n361 163.367
R629 B.n359 B.n174 163.367
R630 B.n354 B.n352 163.367
R631 B.n350 B.n178 163.367
R632 B.n346 B.n344 163.367
R633 B.n342 B.n180 163.367
R634 B.n337 B.n335 163.367
R635 B.n333 B.n184 163.367
R636 B.n329 B.n327 163.367
R637 B.n325 B.n186 163.367
R638 B.n321 B.n319 163.367
R639 B.n317 B.n188 163.367
R640 B.n313 B.n311 163.367
R641 B.n309 B.n190 163.367
R642 B.n305 B.n303 163.367
R643 B.n301 B.n192 163.367
R644 B.n297 B.n295 163.367
R645 B.n293 B.n194 163.367
R646 B.n289 B.n287 163.367
R647 B.n285 B.n196 163.367
R648 B.n281 B.n279 163.367
R649 B.n277 B.n198 163.367
R650 B.n273 B.n271 163.367
R651 B.n269 B.n200 163.367
R652 B.n265 B.n263 163.367
R653 B.n261 B.n202 163.367
R654 B.n257 B.n255 163.367
R655 B.n253 B.n204 163.367
R656 B.n249 B.n247 163.367
R657 B.n245 B.n206 163.367
R658 B.n241 B.n239 163.367
R659 B.n237 B.n208 163.367
R660 B.n233 B.n231 163.367
R661 B.n229 B.n210 163.367
R662 B.n225 B.n223 163.367
R663 B.n221 B.n212 163.367
R664 B.n217 B.n215 163.367
R665 B.n486 B.n138 163.367
R666 B.n490 B.n138 163.367
R667 B.n490 B.n132 163.367
R668 B.n498 B.n132 163.367
R669 B.n498 B.n130 163.367
R670 B.n502 B.n130 163.367
R671 B.n502 B.n123 163.367
R672 B.n510 B.n123 163.367
R673 B.n510 B.n121 163.367
R674 B.n514 B.n121 163.367
R675 B.n514 B.n116 163.367
R676 B.n523 B.n116 163.367
R677 B.n523 B.n114 163.367
R678 B.n528 B.n114 163.367
R679 B.n528 B.n110 163.367
R680 B.n537 B.n110 163.367
R681 B.n538 B.n537 163.367
R682 B.n538 B.n5 163.367
R683 B.n6 B.n5 163.367
R684 B.n7 B.n6 163.367
R685 B.n543 B.n7 163.367
R686 B.n543 B.n12 163.367
R687 B.n13 B.n12 163.367
R688 B.n14 B.n13 163.367
R689 B.n548 B.n14 163.367
R690 B.n548 B.n19 163.367
R691 B.n20 B.n19 163.367
R692 B.n21 B.n20 163.367
R693 B.n553 B.n21 163.367
R694 B.n553 B.n26 163.367
R695 B.n27 B.n26 163.367
R696 B.n28 B.n27 163.367
R697 B.n558 B.n28 163.367
R698 B.n558 B.n33 163.367
R699 B.n34 B.n33 163.367
R700 B.n35 B.n34 163.367
R701 B.n831 B.n829 163.367
R702 B.n827 B.n39 163.367
R703 B.n823 B.n821 163.367
R704 B.n819 B.n41 163.367
R705 B.n815 B.n813 163.367
R706 B.n811 B.n43 163.367
R707 B.n807 B.n805 163.367
R708 B.n803 B.n45 163.367
R709 B.n799 B.n797 163.367
R710 B.n795 B.n47 163.367
R711 B.n791 B.n789 163.367
R712 B.n787 B.n49 163.367
R713 B.n783 B.n781 163.367
R714 B.n779 B.n51 163.367
R715 B.n775 B.n773 163.367
R716 B.n771 B.n53 163.367
R717 B.n767 B.n765 163.367
R718 B.n763 B.n55 163.367
R719 B.n759 B.n757 163.367
R720 B.n755 B.n57 163.367
R721 B.n751 B.n749 163.367
R722 B.n747 B.n59 163.367
R723 B.n743 B.n741 163.367
R724 B.n739 B.n61 163.367
R725 B.n735 B.n733 163.367
R726 B.n731 B.n63 163.367
R727 B.n727 B.n725 163.367
R728 B.n723 B.n65 163.367
R729 B.n719 B.n717 163.367
R730 B.n715 B.n67 163.367
R731 B.n711 B.n709 163.367
R732 B.n707 B.n69 163.367
R733 B.n703 B.n701 163.367
R734 B.n699 B.n74 163.367
R735 B.n695 B.n693 163.367
R736 B.n691 B.n76 163.367
R737 B.n686 B.n684 163.367
R738 B.n682 B.n80 163.367
R739 B.n678 B.n676 163.367
R740 B.n674 B.n82 163.367
R741 B.n670 B.n668 163.367
R742 B.n666 B.n84 163.367
R743 B.n662 B.n660 163.367
R744 B.n658 B.n86 163.367
R745 B.n654 B.n652 163.367
R746 B.n650 B.n88 163.367
R747 B.n646 B.n644 163.367
R748 B.n642 B.n90 163.367
R749 B.n638 B.n636 163.367
R750 B.n634 B.n92 163.367
R751 B.n630 B.n628 163.367
R752 B.n626 B.n94 163.367
R753 B.n622 B.n620 163.367
R754 B.n618 B.n96 163.367
R755 B.n614 B.n612 163.367
R756 B.n610 B.n98 163.367
R757 B.n606 B.n604 163.367
R758 B.n602 B.n100 163.367
R759 B.n598 B.n596 163.367
R760 B.n594 B.n102 163.367
R761 B.n590 B.n588 163.367
R762 B.n586 B.n104 163.367
R763 B.n582 B.n580 163.367
R764 B.n578 B.n106 163.367
R765 B.n574 B.n572 163.367
R766 B.n570 B.n108 163.367
R767 B.n566 B.n564 163.367
R768 B.n181 B.t21 84.0528
R769 B.n77 B.t10 84.0528
R770 B.n175 B.t18 84.027
R771 B.n70 B.t13 84.027
R772 B.n479 B.n142 71.676
R773 B.n477 B.n144 71.676
R774 B.n473 B.n472 71.676
R775 B.n466 B.n146 71.676
R776 B.n465 B.n464 71.676
R777 B.n458 B.n148 71.676
R778 B.n457 B.n456 71.676
R779 B.n450 B.n150 71.676
R780 B.n449 B.n448 71.676
R781 B.n442 B.n152 71.676
R782 B.n441 B.n440 71.676
R783 B.n434 B.n154 71.676
R784 B.n433 B.n432 71.676
R785 B.n426 B.n156 71.676
R786 B.n425 B.n424 71.676
R787 B.n418 B.n158 71.676
R788 B.n417 B.n416 71.676
R789 B.n410 B.n160 71.676
R790 B.n409 B.n408 71.676
R791 B.n402 B.n162 71.676
R792 B.n401 B.n400 71.676
R793 B.n394 B.n164 71.676
R794 B.n393 B.n392 71.676
R795 B.n386 B.n166 71.676
R796 B.n385 B.n384 71.676
R797 B.n378 B.n168 71.676
R798 B.n377 B.n376 71.676
R799 B.n370 B.n170 71.676
R800 B.n369 B.n368 71.676
R801 B.n362 B.n172 71.676
R802 B.n361 B.n360 71.676
R803 B.n353 B.n174 71.676
R804 B.n352 B.n351 71.676
R805 B.n345 B.n178 71.676
R806 B.n344 B.n343 71.676
R807 B.n336 B.n180 71.676
R808 B.n335 B.n334 71.676
R809 B.n328 B.n184 71.676
R810 B.n327 B.n326 71.676
R811 B.n320 B.n186 71.676
R812 B.n319 B.n318 71.676
R813 B.n312 B.n188 71.676
R814 B.n311 B.n310 71.676
R815 B.n304 B.n190 71.676
R816 B.n303 B.n302 71.676
R817 B.n296 B.n192 71.676
R818 B.n295 B.n294 71.676
R819 B.n288 B.n194 71.676
R820 B.n287 B.n286 71.676
R821 B.n280 B.n196 71.676
R822 B.n279 B.n278 71.676
R823 B.n272 B.n198 71.676
R824 B.n271 B.n270 71.676
R825 B.n264 B.n200 71.676
R826 B.n263 B.n262 71.676
R827 B.n256 B.n202 71.676
R828 B.n255 B.n254 71.676
R829 B.n248 B.n204 71.676
R830 B.n247 B.n246 71.676
R831 B.n240 B.n206 71.676
R832 B.n239 B.n238 71.676
R833 B.n232 B.n208 71.676
R834 B.n231 B.n230 71.676
R835 B.n224 B.n210 71.676
R836 B.n223 B.n222 71.676
R837 B.n216 B.n212 71.676
R838 B.n215 B.n214 71.676
R839 B.n830 B.n37 71.676
R840 B.n829 B.n828 71.676
R841 B.n822 B.n39 71.676
R842 B.n821 B.n820 71.676
R843 B.n814 B.n41 71.676
R844 B.n813 B.n812 71.676
R845 B.n806 B.n43 71.676
R846 B.n805 B.n804 71.676
R847 B.n798 B.n45 71.676
R848 B.n797 B.n796 71.676
R849 B.n790 B.n47 71.676
R850 B.n789 B.n788 71.676
R851 B.n782 B.n49 71.676
R852 B.n781 B.n780 71.676
R853 B.n774 B.n51 71.676
R854 B.n773 B.n772 71.676
R855 B.n766 B.n53 71.676
R856 B.n765 B.n764 71.676
R857 B.n758 B.n55 71.676
R858 B.n757 B.n756 71.676
R859 B.n750 B.n57 71.676
R860 B.n749 B.n748 71.676
R861 B.n742 B.n59 71.676
R862 B.n741 B.n740 71.676
R863 B.n734 B.n61 71.676
R864 B.n733 B.n732 71.676
R865 B.n726 B.n63 71.676
R866 B.n725 B.n724 71.676
R867 B.n718 B.n65 71.676
R868 B.n717 B.n716 71.676
R869 B.n710 B.n67 71.676
R870 B.n709 B.n708 71.676
R871 B.n702 B.n69 71.676
R872 B.n701 B.n700 71.676
R873 B.n694 B.n74 71.676
R874 B.n693 B.n692 71.676
R875 B.n685 B.n76 71.676
R876 B.n684 B.n683 71.676
R877 B.n677 B.n80 71.676
R878 B.n676 B.n675 71.676
R879 B.n669 B.n82 71.676
R880 B.n668 B.n667 71.676
R881 B.n661 B.n84 71.676
R882 B.n660 B.n659 71.676
R883 B.n653 B.n86 71.676
R884 B.n652 B.n651 71.676
R885 B.n645 B.n88 71.676
R886 B.n644 B.n643 71.676
R887 B.n637 B.n90 71.676
R888 B.n636 B.n635 71.676
R889 B.n629 B.n92 71.676
R890 B.n628 B.n627 71.676
R891 B.n621 B.n94 71.676
R892 B.n620 B.n619 71.676
R893 B.n613 B.n96 71.676
R894 B.n612 B.n611 71.676
R895 B.n605 B.n98 71.676
R896 B.n604 B.n603 71.676
R897 B.n597 B.n100 71.676
R898 B.n596 B.n595 71.676
R899 B.n589 B.n102 71.676
R900 B.n588 B.n587 71.676
R901 B.n581 B.n104 71.676
R902 B.n580 B.n579 71.676
R903 B.n573 B.n106 71.676
R904 B.n572 B.n571 71.676
R905 B.n565 B.n108 71.676
R906 B.n566 B.n565 71.676
R907 B.n571 B.n570 71.676
R908 B.n574 B.n573 71.676
R909 B.n579 B.n578 71.676
R910 B.n582 B.n581 71.676
R911 B.n587 B.n586 71.676
R912 B.n590 B.n589 71.676
R913 B.n595 B.n594 71.676
R914 B.n598 B.n597 71.676
R915 B.n603 B.n602 71.676
R916 B.n606 B.n605 71.676
R917 B.n611 B.n610 71.676
R918 B.n614 B.n613 71.676
R919 B.n619 B.n618 71.676
R920 B.n622 B.n621 71.676
R921 B.n627 B.n626 71.676
R922 B.n630 B.n629 71.676
R923 B.n635 B.n634 71.676
R924 B.n638 B.n637 71.676
R925 B.n643 B.n642 71.676
R926 B.n646 B.n645 71.676
R927 B.n651 B.n650 71.676
R928 B.n654 B.n653 71.676
R929 B.n659 B.n658 71.676
R930 B.n662 B.n661 71.676
R931 B.n667 B.n666 71.676
R932 B.n670 B.n669 71.676
R933 B.n675 B.n674 71.676
R934 B.n678 B.n677 71.676
R935 B.n683 B.n682 71.676
R936 B.n686 B.n685 71.676
R937 B.n692 B.n691 71.676
R938 B.n695 B.n694 71.676
R939 B.n700 B.n699 71.676
R940 B.n703 B.n702 71.676
R941 B.n708 B.n707 71.676
R942 B.n711 B.n710 71.676
R943 B.n716 B.n715 71.676
R944 B.n719 B.n718 71.676
R945 B.n724 B.n723 71.676
R946 B.n727 B.n726 71.676
R947 B.n732 B.n731 71.676
R948 B.n735 B.n734 71.676
R949 B.n740 B.n739 71.676
R950 B.n743 B.n742 71.676
R951 B.n748 B.n747 71.676
R952 B.n751 B.n750 71.676
R953 B.n756 B.n755 71.676
R954 B.n759 B.n758 71.676
R955 B.n764 B.n763 71.676
R956 B.n767 B.n766 71.676
R957 B.n772 B.n771 71.676
R958 B.n775 B.n774 71.676
R959 B.n780 B.n779 71.676
R960 B.n783 B.n782 71.676
R961 B.n788 B.n787 71.676
R962 B.n791 B.n790 71.676
R963 B.n796 B.n795 71.676
R964 B.n799 B.n798 71.676
R965 B.n804 B.n803 71.676
R966 B.n807 B.n806 71.676
R967 B.n812 B.n811 71.676
R968 B.n815 B.n814 71.676
R969 B.n820 B.n819 71.676
R970 B.n823 B.n822 71.676
R971 B.n828 B.n827 71.676
R972 B.n831 B.n830 71.676
R973 B.n480 B.n479 71.676
R974 B.n474 B.n144 71.676
R975 B.n472 B.n471 71.676
R976 B.n467 B.n466 71.676
R977 B.n464 B.n463 71.676
R978 B.n459 B.n458 71.676
R979 B.n456 B.n455 71.676
R980 B.n451 B.n450 71.676
R981 B.n448 B.n447 71.676
R982 B.n443 B.n442 71.676
R983 B.n440 B.n439 71.676
R984 B.n435 B.n434 71.676
R985 B.n432 B.n431 71.676
R986 B.n427 B.n426 71.676
R987 B.n424 B.n423 71.676
R988 B.n419 B.n418 71.676
R989 B.n416 B.n415 71.676
R990 B.n411 B.n410 71.676
R991 B.n408 B.n407 71.676
R992 B.n403 B.n402 71.676
R993 B.n400 B.n399 71.676
R994 B.n395 B.n394 71.676
R995 B.n392 B.n391 71.676
R996 B.n387 B.n386 71.676
R997 B.n384 B.n383 71.676
R998 B.n379 B.n378 71.676
R999 B.n376 B.n375 71.676
R1000 B.n371 B.n370 71.676
R1001 B.n368 B.n367 71.676
R1002 B.n363 B.n362 71.676
R1003 B.n360 B.n359 71.676
R1004 B.n354 B.n353 71.676
R1005 B.n351 B.n350 71.676
R1006 B.n346 B.n345 71.676
R1007 B.n343 B.n342 71.676
R1008 B.n337 B.n336 71.676
R1009 B.n334 B.n333 71.676
R1010 B.n329 B.n328 71.676
R1011 B.n326 B.n325 71.676
R1012 B.n321 B.n320 71.676
R1013 B.n318 B.n317 71.676
R1014 B.n313 B.n312 71.676
R1015 B.n310 B.n309 71.676
R1016 B.n305 B.n304 71.676
R1017 B.n302 B.n301 71.676
R1018 B.n297 B.n296 71.676
R1019 B.n294 B.n293 71.676
R1020 B.n289 B.n288 71.676
R1021 B.n286 B.n285 71.676
R1022 B.n281 B.n280 71.676
R1023 B.n278 B.n277 71.676
R1024 B.n273 B.n272 71.676
R1025 B.n270 B.n269 71.676
R1026 B.n265 B.n264 71.676
R1027 B.n262 B.n261 71.676
R1028 B.n257 B.n256 71.676
R1029 B.n254 B.n253 71.676
R1030 B.n249 B.n248 71.676
R1031 B.n246 B.n245 71.676
R1032 B.n241 B.n240 71.676
R1033 B.n238 B.n237 71.676
R1034 B.n233 B.n232 71.676
R1035 B.n230 B.n229 71.676
R1036 B.n225 B.n224 71.676
R1037 B.n222 B.n221 71.676
R1038 B.n217 B.n216 71.676
R1039 B.n214 B.n140 71.676
R1040 B.n182 B.t20 70.8649
R1041 B.n78 B.t11 70.8649
R1042 B.n176 B.t17 70.8391
R1043 B.n71 B.t14 70.8391
R1044 B.n339 B.n182 59.5399
R1045 B.n357 B.n176 59.5399
R1046 B.n72 B.n71 59.5399
R1047 B.n689 B.n78 59.5399
R1048 B.n485 B.n141 58.8048
R1049 B.n836 B.n36 58.8048
R1050 B.n834 B.n833 35.4346
R1051 B.n487 B.n139 35.4346
R1052 B.n483 B.n482 35.4346
R1053 B.n563 B.n562 35.4346
R1054 B.n485 B.n137 30.5249
R1055 B.n491 B.n137 30.5249
R1056 B.n491 B.n133 30.5249
R1057 B.n497 B.n133 30.5249
R1058 B.n503 B.n129 30.5249
R1059 B.n503 B.n124 30.5249
R1060 B.n509 B.n124 30.5249
R1061 B.n509 B.n125 30.5249
R1062 B.n516 B.n515 30.5249
R1063 B.n522 B.n117 30.5249
R1064 B.n530 B.n529 30.5249
R1065 B.n536 B.n4 30.5249
R1066 B.n870 B.n4 30.5249
R1067 B.n870 B.n869 30.5249
R1068 B.n869 B.n868 30.5249
R1069 B.n862 B.n11 30.5249
R1070 B.n861 B.n860 30.5249
R1071 B.n854 B.n18 30.5249
R1072 B.n853 B.n852 30.5249
R1073 B.n852 B.n22 30.5249
R1074 B.n846 B.n22 30.5249
R1075 B.n846 B.n845 30.5249
R1076 B.n844 B.n29 30.5249
R1077 B.n838 B.n29 30.5249
R1078 B.n838 B.n837 30.5249
R1079 B.n837 B.n836 30.5249
R1080 B.t16 B.n129 24.6893
R1081 B.n845 B.t9 24.6893
R1082 B.n516 B.t7 18.4049
R1083 B.n522 B.t4 18.4049
R1084 B.n530 B.t3 18.4049
R1085 B.n536 B.t0 18.4049
R1086 B.n868 B.t2 18.4049
R1087 B.n862 B.t1 18.4049
R1088 B.n860 B.t6 18.4049
R1089 B.n854 B.t5 18.4049
R1090 B B.n872 18.0485
R1091 B.n182 B.n181 13.1884
R1092 B.n176 B.n175 13.1884
R1093 B.n71 B.n70 13.1884
R1094 B.n78 B.n77 13.1884
R1095 B.n125 B.t7 12.1205
R1096 B.n515 B.t4 12.1205
R1097 B.n117 B.t3 12.1205
R1098 B.n529 B.t0 12.1205
R1099 B.n11 B.t2 12.1205
R1100 B.t1 B.n861 12.1205
R1101 B.n18 B.t6 12.1205
R1102 B.t5 B.n853 12.1205
R1103 B.n833 B.n832 10.6151
R1104 B.n832 B.n38 10.6151
R1105 B.n826 B.n38 10.6151
R1106 B.n826 B.n825 10.6151
R1107 B.n825 B.n824 10.6151
R1108 B.n824 B.n40 10.6151
R1109 B.n818 B.n40 10.6151
R1110 B.n818 B.n817 10.6151
R1111 B.n817 B.n816 10.6151
R1112 B.n816 B.n42 10.6151
R1113 B.n810 B.n42 10.6151
R1114 B.n810 B.n809 10.6151
R1115 B.n809 B.n808 10.6151
R1116 B.n808 B.n44 10.6151
R1117 B.n802 B.n44 10.6151
R1118 B.n802 B.n801 10.6151
R1119 B.n801 B.n800 10.6151
R1120 B.n800 B.n46 10.6151
R1121 B.n794 B.n46 10.6151
R1122 B.n794 B.n793 10.6151
R1123 B.n793 B.n792 10.6151
R1124 B.n792 B.n48 10.6151
R1125 B.n786 B.n48 10.6151
R1126 B.n786 B.n785 10.6151
R1127 B.n785 B.n784 10.6151
R1128 B.n784 B.n50 10.6151
R1129 B.n778 B.n50 10.6151
R1130 B.n778 B.n777 10.6151
R1131 B.n777 B.n776 10.6151
R1132 B.n776 B.n52 10.6151
R1133 B.n770 B.n52 10.6151
R1134 B.n770 B.n769 10.6151
R1135 B.n769 B.n768 10.6151
R1136 B.n768 B.n54 10.6151
R1137 B.n762 B.n54 10.6151
R1138 B.n762 B.n761 10.6151
R1139 B.n761 B.n760 10.6151
R1140 B.n760 B.n56 10.6151
R1141 B.n754 B.n56 10.6151
R1142 B.n754 B.n753 10.6151
R1143 B.n753 B.n752 10.6151
R1144 B.n752 B.n58 10.6151
R1145 B.n746 B.n58 10.6151
R1146 B.n746 B.n745 10.6151
R1147 B.n745 B.n744 10.6151
R1148 B.n744 B.n60 10.6151
R1149 B.n738 B.n60 10.6151
R1150 B.n738 B.n737 10.6151
R1151 B.n737 B.n736 10.6151
R1152 B.n736 B.n62 10.6151
R1153 B.n730 B.n62 10.6151
R1154 B.n730 B.n729 10.6151
R1155 B.n729 B.n728 10.6151
R1156 B.n728 B.n64 10.6151
R1157 B.n722 B.n64 10.6151
R1158 B.n722 B.n721 10.6151
R1159 B.n721 B.n720 10.6151
R1160 B.n720 B.n66 10.6151
R1161 B.n714 B.n66 10.6151
R1162 B.n714 B.n713 10.6151
R1163 B.n713 B.n712 10.6151
R1164 B.n712 B.n68 10.6151
R1165 B.n706 B.n705 10.6151
R1166 B.n705 B.n704 10.6151
R1167 B.n704 B.n73 10.6151
R1168 B.n698 B.n73 10.6151
R1169 B.n698 B.n697 10.6151
R1170 B.n697 B.n696 10.6151
R1171 B.n696 B.n75 10.6151
R1172 B.n690 B.n75 10.6151
R1173 B.n688 B.n687 10.6151
R1174 B.n687 B.n79 10.6151
R1175 B.n681 B.n79 10.6151
R1176 B.n681 B.n680 10.6151
R1177 B.n680 B.n679 10.6151
R1178 B.n679 B.n81 10.6151
R1179 B.n673 B.n81 10.6151
R1180 B.n673 B.n672 10.6151
R1181 B.n672 B.n671 10.6151
R1182 B.n671 B.n83 10.6151
R1183 B.n665 B.n83 10.6151
R1184 B.n665 B.n664 10.6151
R1185 B.n664 B.n663 10.6151
R1186 B.n663 B.n85 10.6151
R1187 B.n657 B.n85 10.6151
R1188 B.n657 B.n656 10.6151
R1189 B.n656 B.n655 10.6151
R1190 B.n655 B.n87 10.6151
R1191 B.n649 B.n87 10.6151
R1192 B.n649 B.n648 10.6151
R1193 B.n648 B.n647 10.6151
R1194 B.n647 B.n89 10.6151
R1195 B.n641 B.n89 10.6151
R1196 B.n641 B.n640 10.6151
R1197 B.n640 B.n639 10.6151
R1198 B.n639 B.n91 10.6151
R1199 B.n633 B.n91 10.6151
R1200 B.n633 B.n632 10.6151
R1201 B.n632 B.n631 10.6151
R1202 B.n631 B.n93 10.6151
R1203 B.n625 B.n93 10.6151
R1204 B.n625 B.n624 10.6151
R1205 B.n624 B.n623 10.6151
R1206 B.n623 B.n95 10.6151
R1207 B.n617 B.n95 10.6151
R1208 B.n617 B.n616 10.6151
R1209 B.n616 B.n615 10.6151
R1210 B.n615 B.n97 10.6151
R1211 B.n609 B.n97 10.6151
R1212 B.n609 B.n608 10.6151
R1213 B.n608 B.n607 10.6151
R1214 B.n607 B.n99 10.6151
R1215 B.n601 B.n99 10.6151
R1216 B.n601 B.n600 10.6151
R1217 B.n600 B.n599 10.6151
R1218 B.n599 B.n101 10.6151
R1219 B.n593 B.n101 10.6151
R1220 B.n593 B.n592 10.6151
R1221 B.n592 B.n591 10.6151
R1222 B.n591 B.n103 10.6151
R1223 B.n585 B.n103 10.6151
R1224 B.n585 B.n584 10.6151
R1225 B.n584 B.n583 10.6151
R1226 B.n583 B.n105 10.6151
R1227 B.n577 B.n105 10.6151
R1228 B.n577 B.n576 10.6151
R1229 B.n576 B.n575 10.6151
R1230 B.n575 B.n107 10.6151
R1231 B.n569 B.n107 10.6151
R1232 B.n569 B.n568 10.6151
R1233 B.n568 B.n567 10.6151
R1234 B.n567 B.n563 10.6151
R1235 B.n488 B.n487 10.6151
R1236 B.n489 B.n488 10.6151
R1237 B.n489 B.n131 10.6151
R1238 B.n499 B.n131 10.6151
R1239 B.n500 B.n499 10.6151
R1240 B.n501 B.n500 10.6151
R1241 B.n501 B.n122 10.6151
R1242 B.n511 B.n122 10.6151
R1243 B.n512 B.n511 10.6151
R1244 B.n513 B.n512 10.6151
R1245 B.n513 B.n115 10.6151
R1246 B.n524 B.n115 10.6151
R1247 B.n525 B.n524 10.6151
R1248 B.n527 B.n525 10.6151
R1249 B.n527 B.n526 10.6151
R1250 B.n526 B.n109 10.6151
R1251 B.n539 B.n109 10.6151
R1252 B.n540 B.n539 10.6151
R1253 B.n541 B.n540 10.6151
R1254 B.n542 B.n541 10.6151
R1255 B.n544 B.n542 10.6151
R1256 B.n545 B.n544 10.6151
R1257 B.n546 B.n545 10.6151
R1258 B.n547 B.n546 10.6151
R1259 B.n549 B.n547 10.6151
R1260 B.n550 B.n549 10.6151
R1261 B.n551 B.n550 10.6151
R1262 B.n552 B.n551 10.6151
R1263 B.n554 B.n552 10.6151
R1264 B.n555 B.n554 10.6151
R1265 B.n556 B.n555 10.6151
R1266 B.n557 B.n556 10.6151
R1267 B.n559 B.n557 10.6151
R1268 B.n560 B.n559 10.6151
R1269 B.n561 B.n560 10.6151
R1270 B.n562 B.n561 10.6151
R1271 B.n482 B.n481 10.6151
R1272 B.n481 B.n143 10.6151
R1273 B.n476 B.n143 10.6151
R1274 B.n476 B.n475 10.6151
R1275 B.n475 B.n145 10.6151
R1276 B.n470 B.n145 10.6151
R1277 B.n470 B.n469 10.6151
R1278 B.n469 B.n468 10.6151
R1279 B.n468 B.n147 10.6151
R1280 B.n462 B.n147 10.6151
R1281 B.n462 B.n461 10.6151
R1282 B.n461 B.n460 10.6151
R1283 B.n460 B.n149 10.6151
R1284 B.n454 B.n149 10.6151
R1285 B.n454 B.n453 10.6151
R1286 B.n453 B.n452 10.6151
R1287 B.n452 B.n151 10.6151
R1288 B.n446 B.n151 10.6151
R1289 B.n446 B.n445 10.6151
R1290 B.n445 B.n444 10.6151
R1291 B.n444 B.n153 10.6151
R1292 B.n438 B.n153 10.6151
R1293 B.n438 B.n437 10.6151
R1294 B.n437 B.n436 10.6151
R1295 B.n436 B.n155 10.6151
R1296 B.n430 B.n155 10.6151
R1297 B.n430 B.n429 10.6151
R1298 B.n429 B.n428 10.6151
R1299 B.n428 B.n157 10.6151
R1300 B.n422 B.n157 10.6151
R1301 B.n422 B.n421 10.6151
R1302 B.n421 B.n420 10.6151
R1303 B.n420 B.n159 10.6151
R1304 B.n414 B.n159 10.6151
R1305 B.n414 B.n413 10.6151
R1306 B.n413 B.n412 10.6151
R1307 B.n412 B.n161 10.6151
R1308 B.n406 B.n161 10.6151
R1309 B.n406 B.n405 10.6151
R1310 B.n405 B.n404 10.6151
R1311 B.n404 B.n163 10.6151
R1312 B.n398 B.n163 10.6151
R1313 B.n398 B.n397 10.6151
R1314 B.n397 B.n396 10.6151
R1315 B.n396 B.n165 10.6151
R1316 B.n390 B.n165 10.6151
R1317 B.n390 B.n389 10.6151
R1318 B.n389 B.n388 10.6151
R1319 B.n388 B.n167 10.6151
R1320 B.n382 B.n167 10.6151
R1321 B.n382 B.n381 10.6151
R1322 B.n381 B.n380 10.6151
R1323 B.n380 B.n169 10.6151
R1324 B.n374 B.n169 10.6151
R1325 B.n374 B.n373 10.6151
R1326 B.n373 B.n372 10.6151
R1327 B.n372 B.n171 10.6151
R1328 B.n366 B.n171 10.6151
R1329 B.n366 B.n365 10.6151
R1330 B.n365 B.n364 10.6151
R1331 B.n364 B.n173 10.6151
R1332 B.n358 B.n173 10.6151
R1333 B.n356 B.n355 10.6151
R1334 B.n355 B.n177 10.6151
R1335 B.n349 B.n177 10.6151
R1336 B.n349 B.n348 10.6151
R1337 B.n348 B.n347 10.6151
R1338 B.n347 B.n179 10.6151
R1339 B.n341 B.n179 10.6151
R1340 B.n341 B.n340 10.6151
R1341 B.n338 B.n183 10.6151
R1342 B.n332 B.n183 10.6151
R1343 B.n332 B.n331 10.6151
R1344 B.n331 B.n330 10.6151
R1345 B.n330 B.n185 10.6151
R1346 B.n324 B.n185 10.6151
R1347 B.n324 B.n323 10.6151
R1348 B.n323 B.n322 10.6151
R1349 B.n322 B.n187 10.6151
R1350 B.n316 B.n187 10.6151
R1351 B.n316 B.n315 10.6151
R1352 B.n315 B.n314 10.6151
R1353 B.n314 B.n189 10.6151
R1354 B.n308 B.n189 10.6151
R1355 B.n308 B.n307 10.6151
R1356 B.n307 B.n306 10.6151
R1357 B.n306 B.n191 10.6151
R1358 B.n300 B.n191 10.6151
R1359 B.n300 B.n299 10.6151
R1360 B.n299 B.n298 10.6151
R1361 B.n298 B.n193 10.6151
R1362 B.n292 B.n193 10.6151
R1363 B.n292 B.n291 10.6151
R1364 B.n291 B.n290 10.6151
R1365 B.n290 B.n195 10.6151
R1366 B.n284 B.n195 10.6151
R1367 B.n284 B.n283 10.6151
R1368 B.n283 B.n282 10.6151
R1369 B.n282 B.n197 10.6151
R1370 B.n276 B.n197 10.6151
R1371 B.n276 B.n275 10.6151
R1372 B.n275 B.n274 10.6151
R1373 B.n274 B.n199 10.6151
R1374 B.n268 B.n199 10.6151
R1375 B.n268 B.n267 10.6151
R1376 B.n267 B.n266 10.6151
R1377 B.n266 B.n201 10.6151
R1378 B.n260 B.n201 10.6151
R1379 B.n260 B.n259 10.6151
R1380 B.n259 B.n258 10.6151
R1381 B.n258 B.n203 10.6151
R1382 B.n252 B.n203 10.6151
R1383 B.n252 B.n251 10.6151
R1384 B.n251 B.n250 10.6151
R1385 B.n250 B.n205 10.6151
R1386 B.n244 B.n205 10.6151
R1387 B.n244 B.n243 10.6151
R1388 B.n243 B.n242 10.6151
R1389 B.n242 B.n207 10.6151
R1390 B.n236 B.n207 10.6151
R1391 B.n236 B.n235 10.6151
R1392 B.n235 B.n234 10.6151
R1393 B.n234 B.n209 10.6151
R1394 B.n228 B.n209 10.6151
R1395 B.n228 B.n227 10.6151
R1396 B.n227 B.n226 10.6151
R1397 B.n226 B.n211 10.6151
R1398 B.n220 B.n211 10.6151
R1399 B.n220 B.n219 10.6151
R1400 B.n219 B.n218 10.6151
R1401 B.n218 B.n213 10.6151
R1402 B.n213 B.n139 10.6151
R1403 B.n483 B.n135 10.6151
R1404 B.n493 B.n135 10.6151
R1405 B.n494 B.n493 10.6151
R1406 B.n495 B.n494 10.6151
R1407 B.n495 B.n127 10.6151
R1408 B.n505 B.n127 10.6151
R1409 B.n506 B.n505 10.6151
R1410 B.n507 B.n506 10.6151
R1411 B.n507 B.n119 10.6151
R1412 B.n518 B.n119 10.6151
R1413 B.n519 B.n518 10.6151
R1414 B.n520 B.n519 10.6151
R1415 B.n520 B.n112 10.6151
R1416 B.n532 B.n112 10.6151
R1417 B.n533 B.n532 10.6151
R1418 B.n534 B.n533 10.6151
R1419 B.n534 B.n0 10.6151
R1420 B.n866 B.n1 10.6151
R1421 B.n866 B.n865 10.6151
R1422 B.n865 B.n864 10.6151
R1423 B.n864 B.n9 10.6151
R1424 B.n858 B.n9 10.6151
R1425 B.n858 B.n857 10.6151
R1426 B.n857 B.n856 10.6151
R1427 B.n856 B.n16 10.6151
R1428 B.n850 B.n16 10.6151
R1429 B.n850 B.n849 10.6151
R1430 B.n849 B.n848 10.6151
R1431 B.n848 B.n24 10.6151
R1432 B.n842 B.n24 10.6151
R1433 B.n842 B.n841 10.6151
R1434 B.n841 B.n840 10.6151
R1435 B.n840 B.n31 10.6151
R1436 B.n834 B.n31 10.6151
R1437 B.n706 B.n72 6.5566
R1438 B.n690 B.n689 6.5566
R1439 B.n357 B.n356 6.5566
R1440 B.n340 B.n339 6.5566
R1441 B.n497 B.t16 5.83604
R1442 B.t9 B.n844 5.83604
R1443 B.n72 B.n68 4.05904
R1444 B.n689 B.n688 4.05904
R1445 B.n358 B.n357 4.05904
R1446 B.n339 B.n338 4.05904
R1447 B.n872 B.n0 2.81026
R1448 B.n872 B.n1 2.81026
R1449 VP.n3 VP.t7 1466.45
R1450 VP.n12 VP.t2 1450.92
R1451 VP.n1 VP.t3 1450.92
R1452 VP.n6 VP.t0 1450.92
R1453 VP.n10 VP.t1 1437.05
R1454 VP.n11 VP.t4 1437.05
R1455 VP.n5 VP.t5 1437.05
R1456 VP.n4 VP.t6 1437.05
R1457 VP.n13 VP.n12 161.3
R1458 VP.n5 VP.n2 161.3
R1459 VP.n7 VP.n6 161.3
R1460 VP.n11 VP.n0 161.3
R1461 VP.n10 VP.n9 161.3
R1462 VP.n8 VP.n1 161.3
R1463 VP.n3 VP.n2 73.1314
R1464 VP.n11 VP.n10 48.2005
R1465 VP.n5 VP.n4 48.2005
R1466 VP.n8 VP.n7 45.9172
R1467 VP.n10 VP.n1 34.3247
R1468 VP.n12 VP.n11 34.3247
R1469 VP.n6 VP.n5 34.3247
R1470 VP.n4 VP.n3 15.5045
R1471 VP.n7 VP.n2 0.189894
R1472 VP.n9 VP.n8 0.189894
R1473 VP.n9 VP.n0 0.189894
R1474 VP.n13 VP.n0 0.189894
R1475 VP VP.n13 0.0516364
R1476 VTAIL.n11 VTAIL.t12 43.2165
R1477 VTAIL.n10 VTAIL.t0 43.2165
R1478 VTAIL.n7 VTAIL.t6 43.2165
R1479 VTAIL.n14 VTAIL.t9 43.2163
R1480 VTAIL.n15 VTAIL.t4 43.2163
R1481 VTAIL.n2 VTAIL.t1 43.2163
R1482 VTAIL.n3 VTAIL.t13 43.2163
R1483 VTAIL.n6 VTAIL.t8 43.2163
R1484 VTAIL.n13 VTAIL.n12 42.1869
R1485 VTAIL.n9 VTAIL.n8 42.1869
R1486 VTAIL.n1 VTAIL.n0 42.1868
R1487 VTAIL.n5 VTAIL.n4 42.1868
R1488 VTAIL.n15 VTAIL.n14 29.5307
R1489 VTAIL.n7 VTAIL.n6 29.5307
R1490 VTAIL.n0 VTAIL.t3 1.03014
R1491 VTAIL.n0 VTAIL.t5 1.03014
R1492 VTAIL.n4 VTAIL.t7 1.03014
R1493 VTAIL.n4 VTAIL.t14 1.03014
R1494 VTAIL.n12 VTAIL.t11 1.03014
R1495 VTAIL.n12 VTAIL.t10 1.03014
R1496 VTAIL.n8 VTAIL.t15 1.03014
R1497 VTAIL.n8 VTAIL.t2 1.03014
R1498 VTAIL.n9 VTAIL.n7 0.586707
R1499 VTAIL.n10 VTAIL.n9 0.586707
R1500 VTAIL.n13 VTAIL.n11 0.586707
R1501 VTAIL.n14 VTAIL.n13 0.586707
R1502 VTAIL.n6 VTAIL.n5 0.586707
R1503 VTAIL.n5 VTAIL.n3 0.586707
R1504 VTAIL.n2 VTAIL.n1 0.586707
R1505 VTAIL VTAIL.n15 0.528517
R1506 VTAIL.n11 VTAIL.n10 0.470328
R1507 VTAIL.n3 VTAIL.n2 0.470328
R1508 VTAIL VTAIL.n1 0.0586897
R1509 VDD1 VDD1.n0 59.217
R1510 VDD1.n3 VDD1.n2 59.1034
R1511 VDD1.n3 VDD1.n1 59.1034
R1512 VDD1.n5 VDD1.n4 58.8655
R1513 VDD1.n5 VDD1.n3 43.5138
R1514 VDD1.n4 VDD1.t2 1.03014
R1515 VDD1.n4 VDD1.t7 1.03014
R1516 VDD1.n0 VDD1.t0 1.03014
R1517 VDD1.n0 VDD1.t1 1.03014
R1518 VDD1.n2 VDD1.t3 1.03014
R1519 VDD1.n2 VDD1.t5 1.03014
R1520 VDD1.n1 VDD1.t4 1.03014
R1521 VDD1.n1 VDD1.t6 1.03014
R1522 VDD1 VDD1.n5 0.235414
R1523 VN.n1 VN.t0 1466.45
R1524 VN.n7 VN.t1 1466.45
R1525 VN.n4 VN.t3 1450.92
R1526 VN.n10 VN.t4 1450.92
R1527 VN.n2 VN.t5 1437.05
R1528 VN.n3 VN.t7 1437.05
R1529 VN.n8 VN.t2 1437.05
R1530 VN.n9 VN.t6 1437.05
R1531 VN.n5 VN.n4 161.3
R1532 VN.n11 VN.n10 161.3
R1533 VN.n9 VN.n6 161.3
R1534 VN.n3 VN.n0 161.3
R1535 VN.n7 VN.n6 73.1314
R1536 VN.n1 VN.n0 73.1314
R1537 VN.n3 VN.n2 48.2005
R1538 VN.n9 VN.n8 48.2005
R1539 VN VN.n11 46.2979
R1540 VN.n4 VN.n3 34.3247
R1541 VN.n10 VN.n9 34.3247
R1542 VN.n8 VN.n7 15.5045
R1543 VN.n2 VN.n1 15.5045
R1544 VN.n11 VN.n6 0.189894
R1545 VN.n5 VN.n0 0.189894
R1546 VN VN.n5 0.0516364
R1547 VDD2.n2 VDD2.n1 59.1034
R1548 VDD2.n2 VDD2.n0 59.1034
R1549 VDD2 VDD2.n5 59.1004
R1550 VDD2.n4 VDD2.n3 58.8657
R1551 VDD2.n4 VDD2.n2 42.9308
R1552 VDD2.n5 VDD2.t5 1.03014
R1553 VDD2.n5 VDD2.t6 1.03014
R1554 VDD2.n3 VDD2.t3 1.03014
R1555 VDD2.n3 VDD2.t1 1.03014
R1556 VDD2.n1 VDD2.t0 1.03014
R1557 VDD2.n1 VDD2.t4 1.03014
R1558 VDD2.n0 VDD2.t7 1.03014
R1559 VDD2.n0 VDD2.t2 1.03014
R1560 VDD2 VDD2.n4 0.351793
C0 VP VDD2 0.279925f
C1 VN VDD1 0.147339f
C2 VN VTAIL 4.9958f
C3 VP VDD1 5.8285f
C4 VP VTAIL 5.0099f
C5 VDD2 VDD1 0.653877f
C6 VP VN 6.249f
C7 VDD2 VTAIL 23.461302f
C8 VTAIL VDD1 23.421999f
C9 VDD2 VN 5.69617f
C10 VDD2 B 3.751082f
C11 VDD1 B 3.947458f
C12 VTAIL B 12.482347f
C13 VN B 8.42509f
C14 VP B 5.749989f
C15 VDD2.t7 B 0.4952f
C16 VDD2.t2 B 0.4952f
C17 VDD2.n0 B 4.520471f
C18 VDD2.t0 B 0.4952f
C19 VDD2.t4 B 0.4952f
C20 VDD2.n1 B 4.520471f
C21 VDD2.n2 B 3.16468f
C22 VDD2.t3 B 0.4952f
C23 VDD2.t1 B 0.4952f
C24 VDD2.n3 B 4.51894f
C25 VDD2.n4 B 3.55811f
C26 VDD2.t5 B 0.4952f
C27 VDD2.t6 B 0.4952f
C28 VDD2.n5 B 4.52042f
C29 VN.n0 B 0.173155f
C30 VN.t0 B 1.02912f
C31 VN.n1 B 0.384921f
C32 VN.t5 B 1.02137f
C33 VN.n2 B 0.396905f
C34 VN.t7 B 1.02137f
C35 VN.n3 B 0.396905f
C36 VN.t3 B 1.025f
C37 VN.n4 B 0.388647f
C38 VN.n5 B 0.041503f
C39 VN.n6 B 0.173155f
C40 VN.t4 B 1.025f
C41 VN.t2 B 1.02137f
C42 VN.t1 B 1.02912f
C43 VN.n7 B 0.384921f
C44 VN.n8 B 0.396905f
C45 VN.t6 B 1.02137f
C46 VN.n9 B 0.396905f
C47 VN.n10 B 0.388647f
C48 VN.n11 B 2.58899f
C49 VDD1.t0 B 0.493167f
C50 VDD1.t1 B 0.493167f
C51 VDD1.n0 B 4.50268f
C52 VDD1.t4 B 0.493167f
C53 VDD1.t6 B 0.493167f
C54 VDD1.n1 B 4.50192f
C55 VDD1.t3 B 0.493167f
C56 VDD1.t5 B 0.493167f
C57 VDD1.n2 B 4.50192f
C58 VDD1.n3 B 3.2207f
C59 VDD1.t2 B 0.493167f
C60 VDD1.t7 B 0.493167f
C61 VDD1.n4 B 4.50038f
C62 VDD1.n5 B 3.5822f
C63 VTAIL.t3 B 0.343896f
C64 VTAIL.t5 B 0.343896f
C65 VTAIL.n0 B 3.06419f
C66 VTAIL.n1 B 0.281853f
C67 VTAIL.t1 B 3.91492f
C68 VTAIL.n2 B 0.39904f
C69 VTAIL.t13 B 3.91492f
C70 VTAIL.n3 B 0.39904f
C71 VTAIL.t7 B 0.343896f
C72 VTAIL.t14 B 0.343896f
C73 VTAIL.n4 B 3.06419f
C74 VTAIL.n5 B 0.320357f
C75 VTAIL.t8 B 3.91492f
C76 VTAIL.n6 B 1.92378f
C77 VTAIL.t6 B 3.91492f
C78 VTAIL.n7 B 1.92378f
C79 VTAIL.t15 B 0.343896f
C80 VTAIL.t2 B 0.343896f
C81 VTAIL.n8 B 3.06418f
C82 VTAIL.n9 B 0.320364f
C83 VTAIL.t0 B 3.91492f
C84 VTAIL.n10 B 0.399035f
C85 VTAIL.t12 B 3.91492f
C86 VTAIL.n11 B 0.399035f
C87 VTAIL.t11 B 0.343896f
C88 VTAIL.t10 B 0.343896f
C89 VTAIL.n12 B 3.06418f
C90 VTAIL.n13 B 0.320364f
C91 VTAIL.t9 B 3.91492f
C92 VTAIL.n14 B 1.92378f
C93 VTAIL.t4 B 3.91492f
C94 VTAIL.n15 B 1.91954f
C95 VP.n0 B 0.054113f
C96 VP.t3 B 1.03568f
C97 VP.n1 B 0.392696f
C98 VP.n2 B 0.174959f
C99 VP.t5 B 1.03201f
C100 VP.t6 B 1.03201f
C101 VP.t7 B 1.03984f
C102 VP.n3 B 0.388931f
C103 VP.n4 B 0.40104f
C104 VP.n5 B 0.40104f
C105 VP.t0 B 1.03568f
C106 VP.n6 B 0.392696f
C107 VP.n7 B 2.58062f
C108 VP.n8 B 2.62298f
C109 VP.n9 B 0.054113f
C110 VP.t1 B 1.03201f
C111 VP.n10 B 0.40104f
C112 VP.t4 B 1.03201f
C113 VP.n11 B 0.40104f
C114 VP.t2 B 1.03568f
C115 VP.n12 B 0.392696f
C116 VP.n13 B 0.041936f
.ends

