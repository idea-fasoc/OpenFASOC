* NGSPICE file created from opamp_sample_0015.ext - technology: sky130A

.subckt opamp_sample_0015 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 VOUT.t107 a_n16612_8244.t12 VDD.t197 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X1 a_n7261_9606.t7 a_n7183_9410.t22 VDD.t97 VDD.t96 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.64
X2 VN.t6 GND.t172 GND.t174 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X3 GND.t171 GND.t169 VP.t6 GND.t170 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X4 GND.t185 CS_BIAS.t20 VOUT.t23 GND.t176 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X5 VDD.t196 a_n16612_8244.t13 VOUT.t106 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X6 VDD.t195 a_n16612_8244.t14 VOUT.t105 VDD.t149 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X7 VOUT.t42 CS_BIAS.t21 GND.t227 GND.t18 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X8 a_n16612_8244.t3 VN.t7 a_n7864_n440.t19 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=1.8759 ps=10.4 w=4.81 l=7.38
X9 VDD.t194 a_n16612_8244.t15 VOUT.t104 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0.35805 ps=2.5 w=2.17 l=3.65
X10 a_n7261_9606.t17 a_n7183_9410.t12 a_n7183_9410.t9 VDD.t0 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.64
X11 VDD.t193 a_n16612_8244.t16 VOUT.t103 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X12 VOUT.t102 a_n16612_8244.t17 VDD.t192 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X13 a_n7864_n440.t18 VN.t8 a_n16612_8244.t3 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X14 GND.t229 CS_BIAS.t18 CS_BIAS.t19 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X15 a_n5588_7572.t8 a_n7183_9410.t23 VDD.t99 VDD.t98 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X16 VOUT.t26 CS_BIAS.t22 GND.t188 GND.t18 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X17 VOUT.t19 CS_BIAS.t23 GND.t181 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X18 VDD.t83 VDD.t81 VDD.t82 VDD.t54 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.64
X19 VDD.t80 VDD.t78 VDD.t79 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X20 VDD.t191 a_n16612_8244.t18 VOUT.t101 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X21 a_n7864_n440.t9 VP.t7 a_n7183_9410.t2 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X22 GND.t168 GND.t166 GND.t167 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X23 GND.t165 GND.t163 GND.t164 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X24 VOUT.t100 a_n16612_8244.t19 VDD.t190 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X25 VDD.t189 a_n16612_8244.t20 VOUT.t99 VDD.t147 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0.35805 ps=2.5 w=2.17 l=3.65
X26 VOUT.t98 a_n16612_8244.t21 VDD.t188 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X27 GND.t15 CS_BIAS.t16 CS_BIAS.t17 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X28 VDD.t77 VDD.t75 VDD.t76 VDD.t9 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.64
X29 GND.t162 GND.t160 VP.t5 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X30 VOUT.t33 CS_BIAS.t24 GND.t215 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X31 GND.t233 CS_BIAS.t25 VOUT.t109 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X32 a_n7864_n440.t8 VP.t8 a_n7183_9410.t4 GND.t235 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X33 VDD.t74 VDD.t72 VDD.t73 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X34 VDD.t71 VDD.t69 VDD.t70 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X35 GND.t159 GND.t157 GND.t158 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X36 VDD.t115 a_n7183_9410.t24 a_n7261_9606.t6 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.64
X37 GND.t156 GND.t154 VP.t4 GND.t155 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X38 a_n7183_9410.t4 VP.t9 a_n7864_n440.t7 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X39 VDD.t68 VDD.t66 VDD.t67 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X40 a_n5588_7572.t18 a_n7183_9410.t25 a_n16612_8244.t6 VDD.t116 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X41 GND.t153 GND.t151 GND.t152 GND.t43 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X42 GND.t150 GND.t148 GND.t149 GND.t47 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X43 GND.t147 GND.t145 GND.t146 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X44 VDD.t65 VDD.t63 VDD.t64 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X45 VOUT.t97 a_n16612_8244.t22 VDD.t187 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.8463 ps=5.12 w=2.17 l=3.65
X46 VDD.t62 VDD.t60 VDD.t61 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X47 VOUT.t96 a_n16612_8244.t23 VDD.t186 VDD.t156 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X48 VOUT.t28 CS_BIAS.t26 GND.t190 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X49 VDD.t185 a_n16612_8244.t24 VOUT.t95 VDD.t149 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X50 VDD.t184 a_n16612_8244.t25 VOUT.t94 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X51 VDD.t59 VDD.t57 VDD.t58 VDD.t41 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.64
X52 VDD.t183 a_n16612_8244.t26 VOUT.t93 VDD.t124 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X53 VOUT.t114 a_n5588_7572.t0 sky130_fd_pr__cap_mim_m3_1 l=18.26 w=14.66
X54 GND.t144 GND.t142 GND.t143 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X55 VDD.t201 a_n7183_9410.t26 a_n7261_9606.t5 VDD.t200 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.64
X56 GND.t141 GND.t139 VP.t3 GND.t140 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X57 a_n7864_n440.t24 DIFFPAIR_BIAS.t10 GND.t204 GND.t203 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=1.0803 ps=6.32 w=2.77 l=2.19
X58 VOUT.t14 CS_BIAS.t27 GND.t175 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X59 a_n7261_9606.t4 a_n7183_9410.t27 VDD.t203 VDD.t202 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X60 GND.t138 GND.t136 GND.t137 GND.t104 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0 ps=0 w=4.81 l=7.38
X61 DIFFPAIR_BIAS.t9 DIFFPAIR_BIAS.t8 GND.t206 GND.t205 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=1.0803 ps=6.32 w=2.77 l=2.19
X62 VDD.t181 a_n16612_8244.t27 VOUT.t92 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X63 a_n16612_8244.t0 a_n7183_9410.t28 a_n5588_7572.t17 VDD.t0 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.64
X64 a_n7183_9410.t9 a_n7183_9410.t8 a_n7261_9606.t16 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X65 GND.t135 GND.t133 GND.t134 GND.t43 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X66 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.t6 GND.t208 GND.t207 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=1.0803 ps=6.32 w=2.77 l=2.19
X67 GND.t223 CS_BIAS.t28 VOUT.t39 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X68 VOUT.t91 a_n16612_8244.t28 VDD.t182 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.8463 ps=5.12 w=2.17 l=3.65
X69 VOUT.t90 a_n16612_8244.t29 VDD.t180 VDD.t156 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X70 a_n8273_9606# a_n8273_9606# a_n8273_9606# VDD.t101 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=4.29 ps=23.56 w=5.5 l=3.64
X71 VDD.t56 VDD.t53 VDD.t55 VDD.t54 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.64
X72 VDD.t52 VDD.t50 VDD.t51 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X73 VDD.t179 a_n16612_8244.t30 VOUT.t89 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X74 a_n7183_9410.t5 VP.t10 a_n7864_n440.t6 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=1.8759 ps=10.4 w=4.81 l=7.38
X75 VDD.t178 a_n16612_8244.t31 VOUT.t88 VDD.t147 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0.35805 ps=2.5 w=2.17 l=3.65
X76 VOUT.t0 CS_BIAS.t29 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X77 VDD.t177 a_n16612_8244.t32 VOUT.t87 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X78 a_n7261_9606.t3 a_n7183_9410.t29 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X79 a_n7864_n440.t5 VP.t11 a_n7183_9410.t5 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X80 a_n16612_8244.t1 a_n7183_9410.t30 a_n5588_7572.t16 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X81 GND.t132 GND.t130 GND.t131 GND.t47 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X82 VOUT.t86 a_n16612_8244.t33 VDD.t126 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X83 GND.t7 CS_BIAS.t30 VOUT.t3 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X84 a_n7261_9606.t15 a_n7183_9410.t15 a_n7183_9410.t16 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X85 VOUT.t11 CS_BIAS.t31 GND.t32 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X86 VDD.t176 a_n16612_8244.t34 VOUT.t85 VDD.t124 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X87 a_n7864_n440.t17 VN.t9 a_n16612_8244.t2 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X88 GND.t234 CS_BIAS.t32 VOUT.t110 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X89 GND.t218 CS_BIAS.t33 VOUT.t35 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X90 VOUT.t37 CS_BIAS.t34 GND.t220 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X91 VDD.t175 a_n16612_8244.t35 VOUT.t84 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X92 VDD.t106 a_n7183_9410.t31 a_n5588_7572.t7 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X93 GND.t129 GND.t126 GND.t128 GND.t127 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=0 ps=0 w=2.77 l=2.19
X94 VOUT.t8 CS_BIAS.t35 GND.t26 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X95 VOUT.t5 CS_BIAS.t36 GND.t20 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X96 CS_BIAS.t15 CS_BIAS.t14 GND.t224 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X97 GND.t182 CS_BIAS.t37 VOUT.t20 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X98 GND.t221 CS_BIAS.t12 CS_BIAS.t13 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X99 a_n7864_n440.t16 VN.t10 a_n16612_8244.t10 GND.t235 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X100 VDD.t112 a_n7183_9410.t32 a_n5588_7572.t6 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.64
X101 GND.t116 GND.t114 GND.t115 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X102 GND.t125 GND.t123 GND.t124 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X103 a_n16612_8244.t10 VN.t11 a_n7864_n440.t15 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X104 a_n16612_8244.t7 VN.t12 a_n7864_n440.t14 GND.t24 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0.79365 ps=5.14 w=4.81 l=7.38
X105 VN.t5 GND.t120 GND.t122 GND.t121 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X106 GND.t193 CS_BIAS.t38 VOUT.t31 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X107 VDD.t174 a_n16612_8244.t36 VOUT.t83 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0.35805 ps=2.5 w=2.17 l=3.65
X108 a_n5588_7572.t15 a_n7183_9410.t33 a_n16612_8244.t9 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X109 VOUT.t82 a_n16612_8244.t37 VDD.t173 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X110 VOUT.t81 a_n16612_8244.t38 VDD.t172 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X111 VOUT.t115 a_n5588_7572.t0 sky130_fd_pr__cap_mim_m3_1 l=18.26 w=14.66
X112 VDD.t171 a_n16612_8244.t39 VOUT.t80 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0.35805 ps=2.5 w=2.17 l=3.65
X113 GND.t119 GND.t117 VN.t4 GND.t118 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X114 GND.t216 CS_BIAS.t39 VOUT.t34 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X115 VP.t2 GND.t111 GND.t113 GND.t112 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X116 a_n7864_n440.t23 DIFFPAIR_BIAS.t11 GND.t202 GND.t201 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=1.0803 ps=6.32 w=2.77 l=2.19
X117 CS_BIAS.t11 CS_BIAS.t10 GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X118 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 GND.t210 GND.t209 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=1.0803 ps=6.32 w=2.77 l=2.19
X119 GND.t110 GND.t107 GND.t109 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X120 a_n7183_9410.t2 VP.t12 a_n7864_n440.t4 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=1.8759 ps=10.4 w=4.81 l=7.38
X121 VOUT.t79 a_n16612_8244.t40 VDD.t170 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X122 a_n16612_8244.t9 a_n7183_9410.t34 a_n5588_7572.t14 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.64
X123 VDD.t49 VDD.t47 VDD.t48 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X124 GND.t217 CS_BIAS.t8 CS_BIAS.t9 GND.t176 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X125 GND.t106 GND.t103 GND.t105 GND.t104 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0 ps=0 w=4.81 l=7.38
X126 GND.t49 GND.t46 GND.t48 GND.t47 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X127 a_n7183_9410.t1 VP.t13 a_n7864_n440.t3 GND.t12 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0.79365 ps=5.14 w=4.81 l=7.38
X128 GND.t102 GND.t100 GND.t101 GND.t43 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X129 VOUT.t29 CS_BIAS.t40 GND.t191 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X130 VDD.t46 VDD.t44 VDD.t45 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X131 VOUT.t78 a_n16612_8244.t41 VDD.t169 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.8463 ps=5.12 w=2.17 l=3.65
X132 a_n16612_8244.t8 a_n7183_9410.t35 a_n5588_7572.t13 VDD.t108 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X133 VOUT.t116 a_n5588_7572.t0 sky130_fd_pr__cap_mim_m3_1 l=18.26 w=14.66
X134 VOUT.t77 a_n16612_8244.t42 VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X135 VOUT.t1 CS_BIAS.t41 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X136 VOUT.t76 a_n16612_8244.t43 VDD.t168 VDD.t156 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X137 a_n7183_9410.t16 a_n7183_9410.t21 a_n7261_9606.t14 VDD.t116 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X138 VDD.t160 a_n16612_8244.t44 VOUT.t75 VDD.t124 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X139 VDD.t167 a_n16612_8244.t45 VOUT.t74 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X140 VOUT.t73 a_n16612_8244.t46 VDD.t162 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X141 GND.t99 GND.t97 GND.t98 GND.t75 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0 ps=0 w=4.81 l=7.38
X142 GND.t96 GND.t94 GND.t95 GND.t43 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X143 GND.t93 GND.t91 GND.t92 GND.t47 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X144 CS_BIAS.t7 CS_BIAS.t6 GND.t228 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X145 VDD.t199 a_n7183_9410.t36 a_n7261_9606.t2 VDD.t198 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X146 VOUT.t72 a_n16612_8244.t47 VDD.t166 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.8463 ps=5.12 w=2.17 l=3.65
X147 a_n16612_8244.t11 a_n7183_9410.t37 a_n5588_7572.t12 VDD.t107 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.64
X148 VOUT.t117 a_n5588_7572.t0 sky130_fd_pr__cap_mim_m3_1 l=18.26 w=14.66
X149 VOUT.t111 CS_BIAS.t42 GND.t237 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X150 GND.t239 CS_BIAS.t43 VOUT.t113 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X151 VDD.t161 a_n16612_8244.t48 VOUT.t71 VDD.t149 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X152 GND.t90 GND.t88 VN.t3 GND.t89 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X153 VOUT.t25 CS_BIAS.t44 GND.t187 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X154 VOUT.t70 a_n16612_8244.t49 VDD.t165 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.8463 ps=5.12 w=2.17 l=3.65
X155 a_n7261_9606.t13 a_n7183_9410.t13 a_n7183_9410.t11 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X156 a_n7864_n440.t22 DIFFPAIR_BIAS.t12 GND.t200 GND.t199 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=1.0803 ps=6.32 w=2.77 l=2.19
X157 VDD.t164 a_n16612_8244.t50 VOUT.t69 VDD.t147 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0.35805 ps=2.5 w=2.17 l=3.65
X158 a_n7864_n440.t21 DIFFPAIR_BIAS.t13 GND.t198 GND.t197 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=1.0803 ps=6.32 w=2.77 l=2.19
X159 VDD.t43 VDD.t40 VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.64
X160 a_n5588_7572.t11 a_n7183_9410.t38 a_n16612_8244.t1 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X161 VOUT.t68 a_n16612_8244.t51 VDD.t163 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X162 GND.t222 CS_BIAS.t45 VOUT.t38 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X163 a_n7261_9606.t1 a_n7183_9410.t39 VDD.t85 VDD.t84 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.64
X164 VOUT.t22 CS_BIAS.t46 GND.t184 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X165 VOUT.t67 a_n16612_8244.t52 VDD.t159 VDD.t158 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.8463 ps=5.12 w=2.17 l=3.65
X166 VOUT.t66 a_n16612_8244.t53 VDD.t157 VDD.t156 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X167 VDD.t39 VDD.t37 VDD.t38 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X168 VOUT.t118 a_n5588_7572.t0 sky130_fd_pr__cap_mim_m3_1 l=18.26 w=14.66
X169 GND.t232 CS_BIAS.t47 VOUT.t108 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X170 a_n7183_9410.t3 VP.t14 a_n7864_n440.t2 GND.t24 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0.79365 ps=5.14 w=4.81 l=7.38
X171 VDD.t155 a_n16612_8244.t54 VOUT.t65 VDD.t154 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X172 GND.t225 CS_BIAS.t48 VOUT.t40 GND.t176 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X173 GND.t5 CS_BIAS.t49 VOUT.t2 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X174 GND.t180 CS_BIAS.t50 VOUT.t18 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X175 a_n5588_7572.t5 a_n7183_9410.t40 VDD.t92 VDD.t91 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.64
X176 VOUT.t27 CS_BIAS.t51 GND.t189 GND.t18 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X177 VOUT.t30 CS_BIAS.t52 GND.t192 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X178 VOUT.t64 a_n16612_8244.t55 VDD.t153 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X179 VOUT.t63 a_n16612_8244.t56 VDD.t152 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X180 a_n7183_9410.t11 a_n7183_9410.t10 a_n7261_9606.t12 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X181 VOUT.t62 a_n16612_8244.t57 VDD.t151 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X182 VOUT.t36 CS_BIAS.t53 GND.t219 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X183 VOUT.t16 CS_BIAS.t54 GND.t178 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X184 VDD.t36 VDD.t34 VDD.t35 VDD.t5 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.64
X185 GND.t33 CS_BIAS.t55 VOUT.t12 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X186 VOUT.t119 a_n5588_7572.t0 sky130_fd_pr__cap_mim_m3_1 l=18.26 w=14.66
X187 a_n5588_7572.t4 a_n7183_9410.t41 VDD.t94 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X188 a_n16612_8244.t2 VN.t13 a_n7864_n440.t13 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=1.8759 ps=10.4 w=4.81 l=7.38
X189 VDD.t150 a_n16612_8244.t58 VOUT.t61 VDD.t149 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X190 VOUT.t120 a_n5588_7572.t0 sky130_fd_pr__cap_mim_m3_1 l=18.26 w=14.66
X191 a_n16612_8244.t4 VN.t14 a_n7864_n440.t12 GND.t12 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0.79365 ps=5.14 w=4.81 l=7.38
X192 GND.t87 GND.t85 VN.t2 GND.t86 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X193 a_n16612_8244.t5 VN.t15 a_n7864_n440.t11 GND.t13 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X194 VOUT.t10 CS_BIAS.t56 GND.t29 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X195 GND.t84 GND.t82 GND.t83 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X196 a_n7261_9606.t11 a_n7183_9410.t19 a_n7183_9410.t20 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.64
X197 VDD.t148 a_n16612_8244.t59 VOUT.t60 VDD.t147 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0.35805 ps=2.5 w=2.17 l=3.65
X198 VDD.t103 a_n7183_9410.t42 a_n5588_7572.t3 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.64
X199 GND.t179 CS_BIAS.t57 VOUT.t17 GND.t176 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X200 GND.t177 CS_BIAS.t58 VOUT.t15 GND.t176 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X201 a_n7864_n440.t10 VN.t16 a_n16612_8244.t5 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X202 VOUT.t43 CS_BIAS.t59 GND.t230 GND.t18 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X203 GND.t45 GND.t42 GND.t44 GND.t43 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X204 a_n7261_9606.t10 a_n7183_9410.t17 a_n7183_9410.t18 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.64
X205 a_7389_9606# a_7389_9606# a_7389_9606# VDD.t117 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=4.29 ps=23.56 w=5.5 l=3.64
X206 VDD.t146 a_n16612_8244.t60 VOUT.t59 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X207 VDD.t145 a_n16612_8244.t61 VOUT.t58 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0.35805 ps=2.5 w=2.17 l=3.65
X208 VDD.t33 VDD.t31 VDD.t32 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X209 GND.t81 GND.t78 GND.t80 GND.t79 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=0 ps=0 w=2.77 l=2.19
X210 GND.t77 GND.t74 GND.t76 GND.t75 sky130_fd_pr__nfet_01v8 ad=1.8759 pd=10.4 as=0 ps=0 w=4.81 l=7.38
X211 VDD.t30 VDD.t27 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X212 GND.t73 GND.t71 VN.t1 GND.t72 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X213 VOUT.t121 a_n5588_7572.t0 sky130_fd_pr__cap_mim_m3_1 l=18.26 w=14.66
X214 VOUT.t57 a_n16612_8244.t62 VDD.t143 VDD.t142 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X215 VDD.t26 VDD.t23 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X216 GND.t70 GND.t68 GND.t69 GND.t47 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X217 VOUT.t7 CS_BIAS.t60 GND.t22 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X218 CS_BIAS.t5 CS_BIAS.t4 GND.t236 GND.t18 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X219 GND.t67 GND.t65 GND.t66 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X220 VOUT.t56 a_n16612_8244.t63 VDD.t141 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X221 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t212 GND.t211 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=1.0803 ps=6.32 w=2.77 l=2.19
X222 VDD.t139 a_n16612_8244.t64 VOUT.t55 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X223 VDD.t138 a_n16612_8244.t65 VOUT.t54 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X224 a_n16612_8244.t6 a_n7183_9410.t43 a_n5588_7572.t10 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=2.145 ps=11.78 w=5.5 l=3.64
X225 VP.t1 GND.t62 GND.t64 GND.t63 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X226 VOUT.t53 a_n16612_8244.t66 VDD.t136 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X227 VOUT.t52 a_n16612_8244.t67 VDD.t134 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X228 a_n7261_9606.t9 a_n7183_9410.t14 a_n7183_9410.t7 VDD.t107 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.64
X229 VDD.t133 a_n16612_8244.t68 VOUT.t51 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X230 VDD.t22 VDD.t20 VDD.t21 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X231 VDD.t19 VDD.t16 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X232 VOUT.t41 CS_BIAS.t61 GND.t226 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X233 VDD.t15 VDD.t12 VDD.t14 VDD.t13 sky130_fd_pr__pfet_01v8 ad=0.8463 pd=5.12 as=0 ps=0 w=2.17 l=3.65
X234 VOUT.t50 a_n16612_8244.t69 VDD.t132 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.8463 ps=5.12 w=2.17 l=3.65
X235 GND.t61 GND.t59 GND.t60 GND.t47 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X236 VOUT.t49 a_n16612_8244.t70 VDD.t131 VDD.t127 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X237 VOUT.t4 CS_BIAS.t62 GND.t19 GND.t18 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X238 CS_BIAS.t3 CS_BIAS.t2 GND.t31 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X239 VDD.t130 a_n16612_8244.t71 VOUT.t48 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X240 VDD.t11 VDD.t8 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.64
X241 VOUT.t13 CS_BIAS.t63 GND.t34 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X242 a_n5588_7572.t9 a_n7183_9410.t44 a_n16612_8244.t8 VDD.t90 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X243 GND.t58 GND.t56 GND.t57 GND.t43 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X244 a_n7183_9410.t7 a_n7183_9410.t6 a_n7261_9606.t8 VDD.t3 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X245 VDD.t125 a_n16612_8244.t72 VOUT.t47 VDD.t124 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X246 VOUT.t46 a_n16612_8244.t73 VDD.t123 VDD.t122 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X247 VDD.t121 a_n16612_8244.t74 VOUT.t45 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.35805 ps=2.5 w=2.17 l=3.65
X248 VN.t0 GND.t53 GND.t55 GND.t54 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X249 GND.t52 GND.t50 GND.t51 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X250 GND.t238 CS_BIAS.t64 VOUT.t112 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X251 VDD.t110 a_n7183_9410.t45 a_n7261_9606.t0 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X252 VDD.t7 VDD.t4 VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0 ps=0 w=5.5 l=3.64
X253 VOUT.t21 CS_BIAS.t65 GND.t183 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X254 VOUT.t9 CS_BIAS.t66 GND.t28 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.7917 ps=4.84 w=2.03 l=4.49
X255 a_n5588_7572.t2 a_n7183_9410.t46 VDD.t87 VDD.t86 sky130_fd_pr__pfet_01v8 ad=2.145 pd=11.78 as=0.9075 ps=5.83 w=5.5 l=3.64
X256 GND.t194 CS_BIAS.t67 VOUT.t32 GND.t176 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X257 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t214 GND.t213 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=1.0803 ps=6.32 w=2.77 l=2.19
X258 a_n7864_n440.t1 VP.t15 a_n7183_9410.t0 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X259 a_n7183_9410.t0 VP.t16 a_n7864_n440.t0 GND.t13 sky130_fd_pr__nfet_01v8 ad=0.79365 pd=5.14 as=0.79365 ps=5.14 w=4.81 l=7.38
X260 VOUT.t44 a_n16612_8244.t75 VDD.t119 VDD.t118 sky130_fd_pr__pfet_01v8 ad=0.35805 pd=2.5 as=0.8463 ps=5.12 w=2.17 l=3.65
X261 CS_BIAS.t1 CS_BIAS.t0 GND.t231 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0.33495 ps=2.36 w=2.03 l=4.49
X262 GND.t41 GND.t38 GND.t40 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.7917 pd=4.84 as=0 ps=0 w=2.03 l=4.49
X263 VDD.t89 a_n7183_9410.t47 a_n5588_7572.t1 VDD.t88 sky130_fd_pr__pfet_01v8 ad=0.9075 pd=5.83 as=0.9075 ps=5.83 w=5.5 l=3.64
X264 VP.t0 GND.t35 GND.t37 GND.t36 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X265 VOUT.t24 CS_BIAS.t68 GND.t186 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
X266 a_n7864_n440.t20 DIFFPAIR_BIAS.t14 GND.t196 GND.t195 sky130_fd_pr__nfet_01v8 ad=1.0803 pd=6.32 as=1.0803 ps=6.32 w=2.77 l=2.19
X267 VOUT.t6 CS_BIAS.t69 GND.t21 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.33495 pd=2.36 as=0.33495 ps=2.36 w=2.03 l=4.49
R0 a_n16612_8244.n65 a_n16612_8244.n8 28.5074
R1 a_n16612_8244.n66 a_n16612_8244.n9 28.5074
R2 a_n16612_8244.n52 a_n16612_8244.n9 4.72068
R3 a_n16612_8244.n10 a_n16612_8244.n9 4.72068
R4 a_n16612_8244.n53 a_n16612_8244.n9 4.72068
R5 a_n16612_8244.n63 a_n16612_8244.n11 28.5074
R6 a_n16612_8244.n64 a_n16612_8244.n0 28.5074
R7 a_n16612_8244.n50 a_n16612_8244.n0 4.72068
R8 a_n16612_8244.n12 a_n16612_8244.n0 4.72068
R9 a_n16612_8244.n51 a_n16612_8244.n0 4.72068
R10 a_n16612_8244.n61 a_n16612_8244.n13 28.5074
R11 a_n16612_8244.n62 a_n16612_8244.n0 28.5074
R12 a_n16612_8244.n49 a_n16612_8244.n0 4.72068
R13 a_n16612_8244.n59 a_n16612_8244.n15 28.5074
R14 a_n16612_8244.n60 a_n16612_8244.n16 28.5074
R15 a_n16612_8244.n46 a_n16612_8244.n16 4.72068
R16 a_n16612_8244.n17 a_n16612_8244.n16 4.72068
R17 a_n16612_8244.n47 a_n16612_8244.n16 4.72068
R18 a_n16612_8244.n2 a_n16612_8244.n18 4.72081
R19 a_n16612_8244.n2 a_n16612_8244.n44 4.72081
R20 a_n16612_8244.n2 a_n16612_8244.n3 4.72081
R21 a_n16612_8244.n2 a_n16612_8244.n45 4.72081
R22 a_n16612_8244.n1 a_n16612_8244.n19 4.72081
R23 a_n16612_8244.n1 a_n16612_8244.n42 4.72081
R24 a_n16612_8244.n1 a_n16612_8244.n4 4.72081
R25 a_n16612_8244.n1 a_n16612_8244.n43 4.72081
R26 a_n16612_8244.n1 a_n16612_8244.n20 4.72081
R27 a_n16612_8244.n1 a_n16612_8244.n41 4.72081
R28 a_n16612_8244.n6 a_n16612_8244.n21 4.72081
R29 a_n16612_8244.n6 a_n16612_8244.n38 4.72081
R30 a_n16612_8244.n6 a_n16612_8244.n7 4.72081
R31 a_n16612_8244.n6 a_n16612_8244.n39 4.72081
R32 a_n16612_8244.t0 a_n16612_8244.n37 122.654
R33 a_n16612_8244.n36 a_n16612_8244.t11 120.944
R34 a_n16612_8244.n36 a_n16612_8244.t9 116.743
R35 a_n16612_8244.n23 a_n16612_8244.t7 91.7461
R36 a_n16612_8244.n58 a_n16612_8244.t4 91.746
R37 a_n16612_8244.n8 a_n16612_8244.n28 2.39583
R38 a_n16612_8244.n11 a_n16612_8244.n29 2.39583
R39 a_n16612_8244.n13 a_n16612_8244.n30 2.39583
R40 a_n16612_8244.n15 a_n16612_8244.n31 2.39583
R41 a_n16612_8244.n2 a_n16612_8244.t31 47.5269
R42 a_n16612_8244.n1 a_n16612_8244.t50 47.5269
R43 a_n16612_8244.n1 a_n16612_8244.t20 47.5269
R44 a_n16612_8244.n6 a_n16612_8244.t59 47.5269
R45 a_n16612_8244.n8 a_n16612_8244.t22 47.5267
R46 a_n16612_8244.n11 a_n16612_8244.t41 47.5267
R47 a_n16612_8244.n13 a_n16612_8244.t52 47.5267
R48 a_n16612_8244.n15 a_n16612_8244.t28 47.5267
R49 a_n16612_8244.n35 a_n16612_8244.n102 64.9585
R50 a_n16612_8244.n102 a_n16612_8244.n53 58.1796
R51 a_n16612_8244.n53 a_n16612_8244.n103 62.0943
R52 a_n16612_8244.n103 a_n16612_8244.n10 59.1583
R53 a_n16612_8244.n10 a_n16612_8244.n104 61.1157
R54 a_n16612_8244.n104 a_n16612_8244.n52 60.137
R55 a_n16612_8244.n52 a_n16612_8244.n105 60.137
R56 a_n16612_8244.n105 a_n16612_8244.n66 42.0477
R57 a_n16612_8244.n66 a_n16612_8244.n65 115.168
R58 a_n16612_8244.n65 a_n16612_8244.n106 40.0903
R59 a_n16612_8244.n106 a_n16612_8244.n28 64.2457
R60 a_n16612_8244.n34 a_n16612_8244.n97 64.9585
R61 a_n16612_8244.n97 a_n16612_8244.n51 58.1796
R62 a_n16612_8244.n51 a_n16612_8244.n98 62.0943
R63 a_n16612_8244.n98 a_n16612_8244.n12 59.1583
R64 a_n16612_8244.n12 a_n16612_8244.n99 61.1157
R65 a_n16612_8244.n99 a_n16612_8244.n50 60.137
R66 a_n16612_8244.n50 a_n16612_8244.n100 60.137
R67 a_n16612_8244.n100 a_n16612_8244.n64 42.0477
R68 a_n16612_8244.n64 a_n16612_8244.n63 115.168
R69 a_n16612_8244.n63 a_n16612_8244.n101 40.0903
R70 a_n16612_8244.n101 a_n16612_8244.n29 64.2457
R71 a_n16612_8244.n33 a_n16612_8244.n92 64.9585
R72 a_n16612_8244.n92 a_n16612_8244.n49 58.1796
R73 a_n16612_8244.n49 a_n16612_8244.n93 62.0943
R74 a_n16612_8244.n93 a_n16612_8244.n14 59.1583
R75 a_n16612_8244.n14 a_n16612_8244.n94 61.1157
R76 a_n16612_8244.n94 a_n16612_8244.n48 60.137
R77 a_n16612_8244.n48 a_n16612_8244.n95 60.137
R78 a_n16612_8244.n95 a_n16612_8244.n62 42.0477
R79 a_n16612_8244.n62 a_n16612_8244.n61 115.168
R80 a_n16612_8244.n61 a_n16612_8244.n96 40.0903
R81 a_n16612_8244.n96 a_n16612_8244.n30 64.2457
R82 a_n16612_8244.n32 a_n16612_8244.n87 64.9585
R83 a_n16612_8244.n87 a_n16612_8244.n47 58.1796
R84 a_n16612_8244.n47 a_n16612_8244.n88 62.0943
R85 a_n16612_8244.n88 a_n16612_8244.n17 59.1583
R86 a_n16612_8244.n17 a_n16612_8244.n89 61.1157
R87 a_n16612_8244.n89 a_n16612_8244.n46 60.137
R88 a_n16612_8244.n46 a_n16612_8244.n90 60.137
R89 a_n16612_8244.n90 a_n16612_8244.n60 42.0477
R90 a_n16612_8244.n60 a_n16612_8244.n59 115.168
R91 a_n16612_8244.n36 a_n16612_8244.t1 115.034
R92 a_n16612_8244.n37 a_n16612_8244.t8 115.034
R93 a_n16612_8244.n37 a_n16612_8244.t6 115.034
R94 a_n16612_8244.n58 a_n16612_8244.t2 86.7987
R95 a_n16612_8244.n23 a_n16612_8244.t5 84.3065
R96 a_n16612_8244.n23 a_n16612_8244.t3 84.3065
R97 a_n16612_8244.n58 a_n16612_8244.t10 84.3062
R98 a_n16612_8244.n59 a_n16612_8244.n91 40.0903
R99 a_n16612_8244.n91 a_n16612_8244.n31 64.2457
R100 a_n16612_8244.n82 a_n16612_8244.n24 65.6131
R101 a_n16612_8244.n45 a_n16612_8244.n82 59.1584
R102 a_n16612_8244.n83 a_n16612_8244.n45 61.115
R103 a_n16612_8244.n84 a_n16612_8244.n3 60.1363
R104 a_n16612_8244.n44 a_n16612_8244.n84 61.1158
R105 a_n16612_8244.n85 a_n16612_8244.n44 59.1577
R106 a_n16612_8244.n18 a_n16612_8244.n85 62.0944
R107 a_n16612_8244.n86 a_n16612_8244.n18 58.179
R108 a_n16612_8244.n77 a_n16612_8244.n25 65.6131
R109 a_n16612_8244.n43 a_n16612_8244.n77 59.1584
R110 a_n16612_8244.n78 a_n16612_8244.n43 61.115
R111 a_n16612_8244.n79 a_n16612_8244.n4 60.1363
R112 a_n16612_8244.n42 a_n16612_8244.n79 61.1158
R113 a_n16612_8244.n80 a_n16612_8244.n42 59.1577
R114 a_n16612_8244.n19 a_n16612_8244.n80 62.0944
R115 a_n16612_8244.n81 a_n16612_8244.n19 58.179
R116 a_n16612_8244.n72 a_n16612_8244.n26 65.6131
R117 a_n16612_8244.n41 a_n16612_8244.n72 59.1584
R118 a_n16612_8244.n73 a_n16612_8244.n41 61.115
R119 a_n16612_8244.n74 a_n16612_8244.n5 60.1363
R120 a_n16612_8244.n40 a_n16612_8244.n74 61.1158
R121 a_n16612_8244.n75 a_n16612_8244.n40 59.1577
R122 a_n16612_8244.n20 a_n16612_8244.n75 62.0944
R123 a_n16612_8244.n76 a_n16612_8244.n20 58.179
R124 a_n16612_8244.n67 a_n16612_8244.n27 65.6131
R125 a_n16612_8244.n39 a_n16612_8244.n67 59.1584
R126 a_n16612_8244.n68 a_n16612_8244.n39 61.115
R127 a_n16612_8244.n69 a_n16612_8244.n7 60.1363
R128 a_n16612_8244.n38 a_n16612_8244.n69 61.1158
R129 a_n16612_8244.n70 a_n16612_8244.n38 59.1577
R130 a_n16612_8244.n21 a_n16612_8244.n70 62.0944
R131 a_n16612_8244.n71 a_n16612_8244.n21 58.179
R132 a_n16612_8244.n86 a_n16612_8244.n54 64.9587
R133 a_n16612_8244.n81 a_n16612_8244.n55 64.9587
R134 a_n16612_8244.n76 a_n16612_8244.n56 64.9587
R135 a_n16612_8244.n71 a_n16612_8244.n57 64.9587
R136 a_n16612_8244.n35 a_n16612_8244.t39 46.7928
R137 a_n16612_8244.n102 a_n16612_8244.t46 14.3284
R138 a_n16612_8244.n103 a_n16612_8244.t74 14.3284
R139 a_n16612_8244.n104 a_n16612_8244.t19 14.3284
R140 a_n16612_8244.n105 a_n16612_8244.t45 14.3284
R141 a_n16612_8244.n106 a_n16612_8244.t57 14.3284
R142 a_n16612_8244.n28 a_n16612_8244.t60 43.8466
R143 a_n16612_8244.n34 a_n16612_8244.t61 46.7928
R144 a_n16612_8244.n97 a_n16612_8244.t67 14.3284
R145 a_n16612_8244.n98 a_n16612_8244.t30 14.3284
R146 a_n16612_8244.n99 a_n16612_8244.t38 14.3284
R147 a_n16612_8244.n100 a_n16612_8244.t65 14.3284
R148 a_n16612_8244.n101 a_n16612_8244.t12 14.3284
R149 a_n16612_8244.n29 a_n16612_8244.t18 43.8466
R150 a_n16612_8244.n33 a_n16612_8244.t36 46.7928
R151 a_n16612_8244.n92 a_n16612_8244.t70 14.3284
R152 a_n16612_8244.n93 a_n16612_8244.t27 14.3284
R153 a_n16612_8244.n94 a_n16612_8244.t66 14.3284
R154 a_n16612_8244.n95 a_n16612_8244.t25 14.3284
R155 a_n16612_8244.n96 a_n16612_8244.t63 14.3284
R156 a_n16612_8244.n30 a_n16612_8244.t32 43.8466
R157 a_n16612_8244.n32 a_n16612_8244.t15 46.7928
R158 a_n16612_8244.n87 a_n16612_8244.t42 14.3284
R159 a_n16612_8244.n88 a_n16612_8244.t68 14.3284
R160 a_n16612_8244.n89 a_n16612_8244.t40 14.3284
R161 a_n16612_8244.n90 a_n16612_8244.t64 14.3284
R162 a_n16612_8244.n91 a_n16612_8244.t37 14.3284
R163 a_n16612_8244.n31 a_n16612_8244.t71 43.8466
R164 a_n16612_8244.n24 a_n16612_8244.t23 43.1259
R165 a_n16612_8244.n82 a_n16612_8244.t16 14.3284
R166 a_n16612_8244.n83 a_n16612_8244.t51 14.3284
R167 a_n16612_8244.n84 a_n16612_8244.t26 14.3284
R168 a_n16612_8244.n85 a_n16612_8244.t62 14.3284
R169 a_n16612_8244.n86 a_n16612_8244.t58 14.3284
R170 a_n16612_8244.n54 a_n16612_8244.t47 46.7925
R171 a_n16612_8244.n25 a_n16612_8244.t43 43.1259
R172 a_n16612_8244.n77 a_n16612_8244.t35 14.3284
R173 a_n16612_8244.n78 a_n16612_8244.t73 14.3284
R174 a_n16612_8244.n79 a_n16612_8244.t44 14.3284
R175 a_n16612_8244.n80 a_n16612_8244.t21 14.3284
R176 a_n16612_8244.n81 a_n16612_8244.t14 14.3284
R177 a_n16612_8244.n55 a_n16612_8244.t69 46.7925
R178 a_n16612_8244.n26 a_n16612_8244.t53 43.1259
R179 a_n16612_8244.n72 a_n16612_8244.t13 14.3284
R180 a_n16612_8244.n73 a_n16612_8244.t56 14.3284
R181 a_n16612_8244.n74 a_n16612_8244.t34 14.3284
R182 a_n16612_8244.n75 a_n16612_8244.t17 14.3284
R183 a_n16612_8244.n76 a_n16612_8244.t48 14.3284
R184 a_n16612_8244.n56 a_n16612_8244.t75 46.7925
R185 a_n16612_8244.n27 a_n16612_8244.t29 43.1259
R186 a_n16612_8244.n67 a_n16612_8244.t54 14.3284
R187 a_n16612_8244.n68 a_n16612_8244.t33 14.3284
R188 a_n16612_8244.n69 a_n16612_8244.t72 14.3284
R189 a_n16612_8244.n70 a_n16612_8244.t55 14.3284
R190 a_n16612_8244.n71 a_n16612_8244.t24 14.3284
R191 a_n16612_8244.n57 a_n16612_8244.t49 46.7925
R192 a_n16612_8244.n83 a_n16612_8244.n3 60.1371
R193 a_n16612_8244.n78 a_n16612_8244.n4 60.1371
R194 a_n16612_8244.n73 a_n16612_8244.n5 60.1371
R195 a_n16612_8244.n68 a_n16612_8244.n7 60.1371
R196 a_n16612_8244.n107 a_n16612_8244.n22 11.4887
R197 a_n16612_8244.n23 a_n16612_8244.n58 45.3758
R198 a_n16612_8244.n107 a_n16612_8244.n36 38.8494
R199 a_n16612_8244.n37 a_n16612_8244.n107 23.2907
R200 a_n16612_8244.n22 a_n16612_8244.n23 15.6869
R201 a_n16612_8244.n22 a_n16612_8244.n0 10.7595
R202 a_n16612_8244.n1 a_n16612_8244.n5 9.9172
R203 a_n16612_8244.n1 a_n16612_8244.n40 9.9172
R204 a_n16612_8244.n48 a_n16612_8244.n0 9.91707
R205 a_n16612_8244.n14 a_n16612_8244.n0 9.91707
R206 a_n16612_8244.n6 a_n16612_8244.n27 9.03267
R207 a_n16612_8244.n1 a_n16612_8244.n26 9.03267
R208 a_n16612_8244.n1 a_n16612_8244.n25 9.03267
R209 a_n16612_8244.n2 a_n16612_8244.n24 9.03267
R210 a_n16612_8244.n0 a_n16612_8244.n9 8.92416
R211 a_n16612_8244.n1 a_n16612_8244.n2 8.92416
R212 a_n16612_8244.n22 a_n16612_8244.n1 8.59153
R213 a_n16612_8244.n16 a_n16612_8244.n32 7.76898
R214 a_n16612_8244.n0 a_n16612_8244.n33 7.76898
R215 a_n16612_8244.n0 a_n16612_8244.n34 7.76898
R216 a_n16612_8244.n9 a_n16612_8244.n35 7.76898
R217 a_n16612_8244.n16 a_n16612_8244.n15 7.36253
R218 a_n16612_8244.n0 a_n16612_8244.n13 7.36253
R219 a_n16612_8244.n0 a_n16612_8244.n11 7.36253
R220 a_n16612_8244.n9 a_n16612_8244.n8 7.36253
R221 a_n16612_8244.n0 a_n16612_8244.n16 7.06052
R222 a_n16612_8244.n1 a_n16612_8244.n6 7.06052
R223 a_n16612_8244.n6 a_n16612_8244.n57 6.82204
R224 a_n16612_8244.n1 a_n16612_8244.n56 6.82204
R225 a_n16612_8244.n1 a_n16612_8244.n55 6.82204
R226 a_n16612_8244.n2 a_n16612_8244.n54 6.82204
R227 VDD.n3915 VDD.n167 507.805
R228 VDD.n3839 VDD.n165 507.805
R229 VDD.n3609 VDD.n393 507.805
R230 VDD.n3607 VDD.n395 507.805
R231 VDD.n2166 VDD.n1140 507.805
R232 VDD.n1966 VDD.n1198 507.805
R233 VDD.n1591 VDD.n1444 507.805
R234 VDD.n1587 VDD.n1442 507.805
R235 VDD.n3082 VDD.n705 342.44
R236 VDD.n3429 VDD.n418 342.44
R237 VDD.n3439 VDD.n410 342.44
R238 VDD.n3036 VDD.n2710 342.44
R239 VDD.n2644 VDD.n745 342.44
R240 VDD.n2597 VDD.n2596 342.44
R241 VDD.n1112 VDD.n1030 342.44
R242 VDD.n2191 VDD.n1013 342.44
R243 VDD.n3393 VDD.n3392 342.44
R244 VDD.n3351 VDD.n3350 342.44
R245 VDD.n2899 VDD.n2898 342.44
R246 VDD.n2850 VDD.n701 342.44
R247 VDD.n2698 VDD.n733 342.44
R248 VDD.n2651 VDD.n732 342.44
R249 VDD.n2054 VDD.n1042 342.44
R250 VDD.n2194 VDD.n1017 342.44
R251 VDD.n1447 VDD.t19 249.659
R252 VDD.n1538 VDD.t62 249.659
R253 VDD.n1492 VDD.t39 249.659
R254 VDD.n1573 VDD.t52 249.659
R255 VDD.n2082 VDD.t70 249.659
R256 VDD.n2105 VDD.t48 249.659
R257 VDD.n2128 VDD.t73 249.659
R258 VDD.n1168 VDD.t29 249.659
R259 VDD.n3841 VDD.t32 249.659
R260 VDD.n219 VDD.t79 249.659
R261 VDD.n3879 VDD.t67 249.659
R262 VDD.n179 VDD.t25 249.659
R263 VDD.n3472 VDD.t46 249.659
R264 VDD.n3489 VDD.t15 249.659
R265 VDD.n3507 VDD.t65 249.659
R266 VDD.n3523 VDD.t22 249.659
R267 VDD.n1989 VDD.t4 245.631
R268 VDD.n736 VDD.t53 245.631
R269 VDD.n1045 VDD.t34 245.631
R270 VDD.n747 VDD.t81 245.631
R271 VDD.n2848 VDD.t75 245.631
R272 VDD.n406 VDD.t40 245.631
R273 VDD.n2724 VDD.t8 245.631
R274 VDD.n445 VDD.t57 245.631
R275 VDD.n1447 VDD.t16 223.552
R276 VDD.n1538 VDD.t60 223.552
R277 VDD.n1492 VDD.t37 223.552
R278 VDD.n1573 VDD.t50 223.552
R279 VDD.n2082 VDD.t69 223.552
R280 VDD.n2105 VDD.t47 223.552
R281 VDD.n2128 VDD.t72 223.552
R282 VDD.n1168 VDD.t27 223.552
R283 VDD.n3841 VDD.t31 223.552
R284 VDD.n219 VDD.t78 223.552
R285 VDD.n3879 VDD.t66 223.552
R286 VDD.n179 VDD.t23 223.552
R287 VDD.n3472 VDD.t44 223.552
R288 VDD.n3489 VDD.t12 223.552
R289 VDD.n3507 VDD.t63 223.552
R290 VDD.n3523 VDD.t20 223.552
R291 VDD.n1989 VDD.t7 190.422
R292 VDD.n736 VDD.t55 190.422
R293 VDD.n1045 VDD.t36 190.422
R294 VDD.n747 VDD.t82 190.422
R295 VDD.n2848 VDD.t77 190.422
R296 VDD.n406 VDD.t42 190.422
R297 VDD.n2724 VDD.t11 190.422
R298 VDD.n445 VDD.t58 190.422
R299 VDD.n2165 VDD.t117 187.581
R300 VDD.t101 VDD.n394 187.581
R301 VDD.n3394 VDD.n3393 185
R302 VDD.n3393 VDD.n415 185
R303 VDD.n3395 VDD.n416 185
R304 VDD.n3434 VDD.n416 185
R305 VDD.n3396 VDD.n425 185
R306 VDD.n425 VDD.n413 185
R307 VDD.n3398 VDD.n3397 185
R308 VDD.n3399 VDD.n3398 185
R309 VDD.n426 VDD.n424 185
R310 VDD.n424 VDD.n421 185
R311 VDD.n3330 VDD.n452 185
R312 VDD.n3340 VDD.n452 185
R313 VDD.n3331 VDD.n460 185
R314 VDD.n460 VDD.n450 185
R315 VDD.n3333 VDD.n3332 185
R316 VDD.n3334 VDD.n3333 185
R317 VDD.n3329 VDD.n459 185
R318 VDD.n459 VDD.n456 185
R319 VDD.n3328 VDD.n3327 185
R320 VDD.n3327 VDD.n3326 185
R321 VDD.n462 VDD.n461 185
R322 VDD.n463 VDD.n462 185
R323 VDD.n3319 VDD.n3318 185
R324 VDD.n3320 VDD.n3319 185
R325 VDD.n3317 VDD.n472 185
R326 VDD.n472 VDD.n469 185
R327 VDD.n3316 VDD.n3315 185
R328 VDD.n3315 VDD.n3314 185
R329 VDD.n474 VDD.n473 185
R330 VDD.n475 VDD.n474 185
R331 VDD.n3307 VDD.n3306 185
R332 VDD.n3308 VDD.n3307 185
R333 VDD.n3305 VDD.n484 185
R334 VDD.n484 VDD.n481 185
R335 VDD.n3304 VDD.n3303 185
R336 VDD.n3303 VDD.n3302 185
R337 VDD.n486 VDD.n485 185
R338 VDD.n487 VDD.n486 185
R339 VDD.n3295 VDD.n3294 185
R340 VDD.n3296 VDD.n3295 185
R341 VDD.n3293 VDD.n496 185
R342 VDD.n496 VDD.n493 185
R343 VDD.n3292 VDD.n3291 185
R344 VDD.n3291 VDD.n3290 185
R345 VDD.n498 VDD.n497 185
R346 VDD.n507 VDD.n498 185
R347 VDD.n3283 VDD.n3282 185
R348 VDD.n3284 VDD.n3283 185
R349 VDD.n3281 VDD.n508 185
R350 VDD.n508 VDD.n504 185
R351 VDD.n3280 VDD.n3279 185
R352 VDD.n3279 VDD.n3278 185
R353 VDD.n510 VDD.n509 185
R354 VDD.n511 VDD.n510 185
R355 VDD.n3271 VDD.n3270 185
R356 VDD.n3272 VDD.n3271 185
R357 VDD.n3269 VDD.n520 185
R358 VDD.n520 VDD.n517 185
R359 VDD.n3268 VDD.n3267 185
R360 VDD.n3267 VDD.n3266 185
R361 VDD.n522 VDD.n521 185
R362 VDD.n523 VDD.n522 185
R363 VDD.n3259 VDD.n3258 185
R364 VDD.n3260 VDD.n3259 185
R365 VDD.n3257 VDD.n532 185
R366 VDD.n532 VDD.n529 185
R367 VDD.n3256 VDD.n3255 185
R368 VDD.n3255 VDD.n3254 185
R369 VDD.n534 VDD.n533 185
R370 VDD.n543 VDD.n534 185
R371 VDD.n3247 VDD.n3246 185
R372 VDD.n3248 VDD.n3247 185
R373 VDD.n3245 VDD.n544 185
R374 VDD.n544 VDD.n540 185
R375 VDD.n3244 VDD.n3243 185
R376 VDD.n3243 VDD.n3242 185
R377 VDD.n546 VDD.n545 185
R378 VDD.n547 VDD.n546 185
R379 VDD.n3235 VDD.n3234 185
R380 VDD.n3236 VDD.n3235 185
R381 VDD.n3233 VDD.n556 185
R382 VDD.n556 VDD.n553 185
R383 VDD.n3232 VDD.n3231 185
R384 VDD.n3231 VDD.n3230 185
R385 VDD.n558 VDD.n557 185
R386 VDD.n559 VDD.n558 185
R387 VDD.n3223 VDD.n3222 185
R388 VDD.n3224 VDD.n3223 185
R389 VDD.n3221 VDD.n568 185
R390 VDD.n568 VDD.n565 185
R391 VDD.n3220 VDD.n3219 185
R392 VDD.n3219 VDD.t108 185
R393 VDD.n570 VDD.n569 185
R394 VDD.n571 VDD.n570 185
R395 VDD.n3212 VDD.n3211 185
R396 VDD.n3213 VDD.n3212 185
R397 VDD.n3210 VDD.n580 185
R398 VDD.n580 VDD.n577 185
R399 VDD.n3209 VDD.n3208 185
R400 VDD.n3208 VDD.n3207 185
R401 VDD.n582 VDD.n581 185
R402 VDD.n591 VDD.n582 185
R403 VDD.n3200 VDD.n3199 185
R404 VDD.n3201 VDD.n3200 185
R405 VDD.n3198 VDD.n592 185
R406 VDD.n592 VDD.n588 185
R407 VDD.n3197 VDD.n3196 185
R408 VDD.n3196 VDD.n3195 185
R409 VDD.n594 VDD.n593 185
R410 VDD.n595 VDD.n594 185
R411 VDD.n3188 VDD.n3187 185
R412 VDD.n3189 VDD.n3188 185
R413 VDD.n3186 VDD.n604 185
R414 VDD.n604 VDD.n601 185
R415 VDD.n3185 VDD.n3184 185
R416 VDD.n3184 VDD.n3183 185
R417 VDD.n606 VDD.n605 185
R418 VDD.n607 VDD.n606 185
R419 VDD.n3176 VDD.n3175 185
R420 VDD.n3177 VDD.n3176 185
R421 VDD.n3174 VDD.n616 185
R422 VDD.n616 VDD.n613 185
R423 VDD.n3173 VDD.n3172 185
R424 VDD.n3172 VDD.n3171 185
R425 VDD.n618 VDD.n617 185
R426 VDD.n627 VDD.n618 185
R427 VDD.n3164 VDD.n3163 185
R428 VDD.n3165 VDD.n3164 185
R429 VDD.n3162 VDD.n628 185
R430 VDD.n628 VDD.n624 185
R431 VDD.n3161 VDD.n3160 185
R432 VDD.n3160 VDD.n3159 185
R433 VDD.n630 VDD.n629 185
R434 VDD.n631 VDD.n630 185
R435 VDD.n3152 VDD.n3151 185
R436 VDD.n3153 VDD.n3152 185
R437 VDD.n3150 VDD.n640 185
R438 VDD.n640 VDD.n637 185
R439 VDD.n3149 VDD.n3148 185
R440 VDD.n3148 VDD.n3147 185
R441 VDD.n642 VDD.n641 185
R442 VDD.n643 VDD.n642 185
R443 VDD.n3140 VDD.n3139 185
R444 VDD.n3141 VDD.n3140 185
R445 VDD.n3138 VDD.n652 185
R446 VDD.n652 VDD.n649 185
R447 VDD.n3137 VDD.n3136 185
R448 VDD.n3136 VDD.n3135 185
R449 VDD.n654 VDD.n653 185
R450 VDD.n663 VDD.n654 185
R451 VDD.n3128 VDD.n3127 185
R452 VDD.n3129 VDD.n3128 185
R453 VDD.n3126 VDD.n664 185
R454 VDD.n664 VDD.n660 185
R455 VDD.n3125 VDD.n3124 185
R456 VDD.n3124 VDD.n3123 185
R457 VDD.n666 VDD.n665 185
R458 VDD.n667 VDD.n666 185
R459 VDD.n3116 VDD.n3115 185
R460 VDD.n3117 VDD.n3116 185
R461 VDD.n3114 VDD.n676 185
R462 VDD.n676 VDD.n673 185
R463 VDD.n3113 VDD.n3112 185
R464 VDD.n3112 VDD.n3111 185
R465 VDD.n678 VDD.n677 185
R466 VDD.n679 VDD.n678 185
R467 VDD.n3104 VDD.n3103 185
R468 VDD.n3105 VDD.n3104 185
R469 VDD.n3102 VDD.n687 185
R470 VDD.n3026 VDD.n687 185
R471 VDD.n3101 VDD.n3100 185
R472 VDD.n3100 VDD.n3099 185
R473 VDD.n689 VDD.n688 185
R474 VDD.n690 VDD.n689 185
R475 VDD.n3092 VDD.n3091 185
R476 VDD.n3093 VDD.n3092 185
R477 VDD.n3090 VDD.n699 185
R478 VDD.n699 VDD.n696 185
R479 VDD.n3089 VDD.n3088 185
R480 VDD.n3088 VDD.n3087 185
R481 VDD.n701 VDD.n700 185
R482 VDD.n702 VDD.n701 185
R483 VDD.n2851 VDD.n2850 185
R484 VDD.n2853 VDD.n2852 185
R485 VDD.n2855 VDD.n2854 185
R486 VDD.n2857 VDD.n2856 185
R487 VDD.n2859 VDD.n2858 185
R488 VDD.n2861 VDD.n2860 185
R489 VDD.n2863 VDD.n2862 185
R490 VDD.n2865 VDD.n2864 185
R491 VDD.n2867 VDD.n2866 185
R492 VDD.n2869 VDD.n2868 185
R493 VDD.n2871 VDD.n2870 185
R494 VDD.n2873 VDD.n2872 185
R495 VDD.n2875 VDD.n2874 185
R496 VDD.n2877 VDD.n2876 185
R497 VDD.n2879 VDD.n2878 185
R498 VDD.n2881 VDD.n2880 185
R499 VDD.n2883 VDD.n2882 185
R500 VDD.n2885 VDD.n2884 185
R501 VDD.n2887 VDD.n2886 185
R502 VDD.n2889 VDD.n2888 185
R503 VDD.n2891 VDD.n2890 185
R504 VDD.n2894 VDD.n2893 185
R505 VDD.n2896 VDD.n2895 185
R506 VDD.n2898 VDD.n2897 185
R507 VDD.n3352 VDD.n3351 185
R508 VDD.n3353 VDD.n444 185
R509 VDD.n3355 VDD.n3354 185
R510 VDD.n3357 VDD.n442 185
R511 VDD.n3359 VDD.n3358 185
R512 VDD.n3360 VDD.n441 185
R513 VDD.n3362 VDD.n3361 185
R514 VDD.n3364 VDD.n439 185
R515 VDD.n3366 VDD.n3365 185
R516 VDD.n3367 VDD.n438 185
R517 VDD.n3369 VDD.n3368 185
R518 VDD.n3371 VDD.n437 185
R519 VDD.n3373 VDD.n3372 185
R520 VDD.n3374 VDD.n434 185
R521 VDD.n3376 VDD.n3375 185
R522 VDD.n3378 VDD.n432 185
R523 VDD.n3380 VDD.n3379 185
R524 VDD.n3381 VDD.n431 185
R525 VDD.n3383 VDD.n3382 185
R526 VDD.n3385 VDD.n429 185
R527 VDD.n3387 VDD.n3386 185
R528 VDD.n3388 VDD.n428 185
R529 VDD.n3390 VDD.n3389 185
R530 VDD.n3392 VDD.n427 185
R531 VDD.n3350 VDD.n3348 185
R532 VDD.n3350 VDD.n415 185
R533 VDD.n3347 VDD.n414 185
R534 VDD.n3434 VDD.n414 185
R535 VDD.n3346 VDD.n3345 185
R536 VDD.n3345 VDD.n413 185
R537 VDD.n3344 VDD.n423 185
R538 VDD.n3399 VDD.n423 185
R539 VDD.n3343 VDD.n3342 185
R540 VDD.n3342 VDD.n421 185
R541 VDD.n3341 VDD.n448 185
R542 VDD.n3341 VDD.n3340 185
R543 VDD.n2908 VDD.n449 185
R544 VDD.n450 VDD.n449 185
R545 VDD.n2909 VDD.n458 185
R546 VDD.n3334 VDD.n458 185
R547 VDD.n2911 VDD.n2910 185
R548 VDD.n2910 VDD.n456 185
R549 VDD.n2912 VDD.n465 185
R550 VDD.n3326 VDD.n465 185
R551 VDD.n2914 VDD.n2913 185
R552 VDD.n2913 VDD.n463 185
R553 VDD.n2915 VDD.n471 185
R554 VDD.n3320 VDD.n471 185
R555 VDD.n2917 VDD.n2916 185
R556 VDD.n2916 VDD.n469 185
R557 VDD.n2918 VDD.n477 185
R558 VDD.n3314 VDD.n477 185
R559 VDD.n2920 VDD.n2919 185
R560 VDD.n2919 VDD.n475 185
R561 VDD.n2921 VDD.n483 185
R562 VDD.n3308 VDD.n483 185
R563 VDD.n2923 VDD.n2922 185
R564 VDD.n2922 VDD.n481 185
R565 VDD.n2924 VDD.n489 185
R566 VDD.n3302 VDD.n489 185
R567 VDD.n2926 VDD.n2925 185
R568 VDD.n2925 VDD.n487 185
R569 VDD.n2927 VDD.n495 185
R570 VDD.n3296 VDD.n495 185
R571 VDD.n2929 VDD.n2928 185
R572 VDD.n2928 VDD.n493 185
R573 VDD.n2930 VDD.n500 185
R574 VDD.n3290 VDD.n500 185
R575 VDD.n2932 VDD.n2931 185
R576 VDD.n2931 VDD.n507 185
R577 VDD.n2933 VDD.n506 185
R578 VDD.n3284 VDD.n506 185
R579 VDD.n2935 VDD.n2934 185
R580 VDD.n2934 VDD.n504 185
R581 VDD.n2936 VDD.n513 185
R582 VDD.n3278 VDD.n513 185
R583 VDD.n2938 VDD.n2937 185
R584 VDD.n2937 VDD.n511 185
R585 VDD.n2939 VDD.n519 185
R586 VDD.n3272 VDD.n519 185
R587 VDD.n2941 VDD.n2940 185
R588 VDD.n2940 VDD.n517 185
R589 VDD.n2942 VDD.n525 185
R590 VDD.n3266 VDD.n525 185
R591 VDD.n2944 VDD.n2943 185
R592 VDD.n2943 VDD.n523 185
R593 VDD.n2945 VDD.n531 185
R594 VDD.n3260 VDD.n531 185
R595 VDD.n2947 VDD.n2946 185
R596 VDD.n2946 VDD.n529 185
R597 VDD.n2948 VDD.n536 185
R598 VDD.n3254 VDD.n536 185
R599 VDD.n2950 VDD.n2949 185
R600 VDD.n2949 VDD.n543 185
R601 VDD.n2951 VDD.n542 185
R602 VDD.n3248 VDD.n542 185
R603 VDD.n2953 VDD.n2952 185
R604 VDD.n2952 VDD.n540 185
R605 VDD.n2954 VDD.n549 185
R606 VDD.n3242 VDD.n549 185
R607 VDD.n2956 VDD.n2955 185
R608 VDD.n2955 VDD.n547 185
R609 VDD.n2957 VDD.n555 185
R610 VDD.n3236 VDD.n555 185
R611 VDD.n2959 VDD.n2958 185
R612 VDD.n2958 VDD.n553 185
R613 VDD.n2960 VDD.n561 185
R614 VDD.n3230 VDD.n561 185
R615 VDD.n2962 VDD.n2961 185
R616 VDD.n2961 VDD.n559 185
R617 VDD.n2963 VDD.n567 185
R618 VDD.n3224 VDD.n567 185
R619 VDD.n2965 VDD.n2964 185
R620 VDD.n2964 VDD.n565 185
R621 VDD.n2966 VDD.n572 185
R622 VDD.t108 VDD.n572 185
R623 VDD.n2968 VDD.n2967 185
R624 VDD.n2967 VDD.n571 185
R625 VDD.n2969 VDD.n579 185
R626 VDD.n3213 VDD.n579 185
R627 VDD.n2971 VDD.n2970 185
R628 VDD.n2970 VDD.n577 185
R629 VDD.n2972 VDD.n584 185
R630 VDD.n3207 VDD.n584 185
R631 VDD.n2974 VDD.n2973 185
R632 VDD.n2973 VDD.n591 185
R633 VDD.n2975 VDD.n590 185
R634 VDD.n3201 VDD.n590 185
R635 VDD.n2977 VDD.n2976 185
R636 VDD.n2976 VDD.n588 185
R637 VDD.n2978 VDD.n597 185
R638 VDD.n3195 VDD.n597 185
R639 VDD.n2980 VDD.n2979 185
R640 VDD.n2979 VDD.n595 185
R641 VDD.n2981 VDD.n603 185
R642 VDD.n3189 VDD.n603 185
R643 VDD.n2983 VDD.n2982 185
R644 VDD.n2982 VDD.n601 185
R645 VDD.n2984 VDD.n609 185
R646 VDD.n3183 VDD.n609 185
R647 VDD.n2986 VDD.n2985 185
R648 VDD.n2985 VDD.n607 185
R649 VDD.n2987 VDD.n615 185
R650 VDD.n3177 VDD.n615 185
R651 VDD.n2989 VDD.n2988 185
R652 VDD.n2988 VDD.n613 185
R653 VDD.n2990 VDD.n620 185
R654 VDD.n3171 VDD.n620 185
R655 VDD.n2992 VDD.n2991 185
R656 VDD.n2991 VDD.n627 185
R657 VDD.n2993 VDD.n626 185
R658 VDD.n3165 VDD.n626 185
R659 VDD.n2995 VDD.n2994 185
R660 VDD.n2994 VDD.n624 185
R661 VDD.n2996 VDD.n633 185
R662 VDD.n3159 VDD.n633 185
R663 VDD.n2998 VDD.n2997 185
R664 VDD.n2997 VDD.n631 185
R665 VDD.n2999 VDD.n639 185
R666 VDD.n3153 VDD.n639 185
R667 VDD.n3001 VDD.n3000 185
R668 VDD.n3000 VDD.n637 185
R669 VDD.n3002 VDD.n645 185
R670 VDD.n3147 VDD.n645 185
R671 VDD.n3004 VDD.n3003 185
R672 VDD.n3003 VDD.n643 185
R673 VDD.n3005 VDD.n651 185
R674 VDD.n3141 VDD.n651 185
R675 VDD.n3007 VDD.n3006 185
R676 VDD.n3006 VDD.n649 185
R677 VDD.n3008 VDD.n656 185
R678 VDD.n3135 VDD.n656 185
R679 VDD.n3010 VDD.n3009 185
R680 VDD.n3009 VDD.n663 185
R681 VDD.n3011 VDD.n662 185
R682 VDD.n3129 VDD.n662 185
R683 VDD.n3013 VDD.n3012 185
R684 VDD.n3012 VDD.n660 185
R685 VDD.n3014 VDD.n669 185
R686 VDD.n3123 VDD.n669 185
R687 VDD.n3016 VDD.n3015 185
R688 VDD.n3015 VDD.n667 185
R689 VDD.n3017 VDD.n675 185
R690 VDD.n3117 VDD.n675 185
R691 VDD.n3019 VDD.n3018 185
R692 VDD.n3018 VDD.n673 185
R693 VDD.n3020 VDD.n681 185
R694 VDD.n3111 VDD.n681 185
R695 VDD.n3022 VDD.n3021 185
R696 VDD.n3021 VDD.n679 185
R697 VDD.n3023 VDD.n686 185
R698 VDD.n3105 VDD.n686 185
R699 VDD.n3025 VDD.n3024 185
R700 VDD.n3026 VDD.n3025 185
R701 VDD.n2907 VDD.n692 185
R702 VDD.n3099 VDD.n692 185
R703 VDD.n2906 VDD.n2905 185
R704 VDD.n2905 VDD.n690 185
R705 VDD.n2904 VDD.n698 185
R706 VDD.n3093 VDD.n698 185
R707 VDD.n2903 VDD.n2902 185
R708 VDD.n2902 VDD.n696 185
R709 VDD.n2901 VDD.n704 185
R710 VDD.n3087 VDD.n704 185
R711 VDD.n2900 VDD.n2899 185
R712 VDD.n2899 VDD.n702 185
R713 VDD.n1961 VDD.n1140 185
R714 VDD.n1142 VDD.n1140 185
R715 VDD.n1963 VDD.n1962 185
R716 VDD.n1964 VDD.n1963 185
R717 VDD.n1204 VDD.n1203 185
R718 VDD.n1203 VDD.n1202 185
R719 VDD.n1957 VDD.n1956 185
R720 VDD.n1956 VDD.n1955 185
R721 VDD.n1207 VDD.n1206 185
R722 VDD.t28 VDD.n1207 185
R723 VDD.n1945 VDD.n1944 185
R724 VDD.n1946 VDD.n1945 185
R725 VDD.n1216 VDD.n1215 185
R726 VDD.n1215 VDD.n1214 185
R727 VDD.n1940 VDD.n1939 185
R728 VDD.n1939 VDD.n1938 185
R729 VDD.n1219 VDD.n1218 185
R730 VDD.n1220 VDD.n1219 185
R731 VDD.n1929 VDD.n1928 185
R732 VDD.n1930 VDD.n1929 185
R733 VDD.n1228 VDD.n1227 185
R734 VDD.n1227 VDD.n1226 185
R735 VDD.n1924 VDD.n1923 185
R736 VDD.n1923 VDD.n1922 185
R737 VDD.n1231 VDD.n1230 185
R738 VDD.n1232 VDD.n1231 185
R739 VDD.n1913 VDD.n1912 185
R740 VDD.n1914 VDD.n1913 185
R741 VDD.n1240 VDD.n1239 185
R742 VDD.n1239 VDD.n1238 185
R743 VDD.n1908 VDD.n1907 185
R744 VDD.n1907 VDD.n1906 185
R745 VDD.n1243 VDD.n1242 185
R746 VDD.n1244 VDD.n1243 185
R747 VDD.n1897 VDD.n1896 185
R748 VDD.n1898 VDD.n1897 185
R749 VDD.n1252 VDD.n1251 185
R750 VDD.n1251 VDD.n1250 185
R751 VDD.n1892 VDD.n1891 185
R752 VDD.n1891 VDD.n1890 185
R753 VDD.n1255 VDD.n1254 185
R754 VDD.n1256 VDD.n1255 185
R755 VDD.n1881 VDD.n1880 185
R756 VDD.n1882 VDD.n1881 185
R757 VDD.n1264 VDD.n1263 185
R758 VDD.n1263 VDD.n1262 185
R759 VDD.n1876 VDD.n1875 185
R760 VDD.n1875 VDD.n1874 185
R761 VDD.n1267 VDD.n1266 185
R762 VDD.n1268 VDD.n1267 185
R763 VDD.n1865 VDD.n1864 185
R764 VDD.n1866 VDD.n1865 185
R765 VDD.n1276 VDD.n1275 185
R766 VDD.n1275 VDD.n1274 185
R767 VDD.n1860 VDD.n1859 185
R768 VDD.n1859 VDD.n1858 185
R769 VDD.n1279 VDD.n1278 185
R770 VDD.n1280 VDD.n1279 185
R771 VDD.n1849 VDD.n1848 185
R772 VDD.n1850 VDD.n1849 185
R773 VDD.n1288 VDD.n1287 185
R774 VDD.n1287 VDD.n1286 185
R775 VDD.n1844 VDD.n1843 185
R776 VDD.n1843 VDD.n1842 185
R777 VDD.n1291 VDD.n1290 185
R778 VDD.n1292 VDD.n1291 185
R779 VDD.n1833 VDD.n1832 185
R780 VDD.n1834 VDD.n1833 185
R781 VDD.n1300 VDD.n1299 185
R782 VDD.n1299 VDD.n1298 185
R783 VDD.n1828 VDD.n1827 185
R784 VDD.n1827 VDD.n1826 185
R785 VDD.n1303 VDD.n1302 185
R786 VDD.n1304 VDD.n1303 185
R787 VDD.n1817 VDD.n1816 185
R788 VDD.n1818 VDD.n1817 185
R789 VDD.n1312 VDD.n1311 185
R790 VDD.n1311 VDD.n1310 185
R791 VDD.n1812 VDD.n1811 185
R792 VDD.n1811 VDD.n1810 185
R793 VDD.n1315 VDD.n1314 185
R794 VDD.n1316 VDD.n1315 185
R795 VDD.n1801 VDD.n1800 185
R796 VDD.n1802 VDD.n1801 185
R797 VDD.n1324 VDD.n1323 185
R798 VDD.n1323 VDD.n1322 185
R799 VDD.n1764 VDD.n1763 185
R800 VDD.n1763 VDD.n1762 185
R801 VDD.n1327 VDD.n1326 185
R802 VDD.n1328 VDD.n1327 185
R803 VDD.n1753 VDD.n1752 185
R804 VDD.n1754 VDD.n1753 185
R805 VDD.n1335 VDD.n1334 185
R806 VDD.n1745 VDD.n1334 185
R807 VDD.n1748 VDD.n1747 185
R808 VDD.n1747 VDD.n1746 185
R809 VDD.n1338 VDD.n1337 185
R810 VDD.n1339 VDD.n1338 185
R811 VDD.n1736 VDD.n1735 185
R812 VDD.n1737 VDD.n1736 185
R813 VDD.n1347 VDD.n1346 185
R814 VDD.n1346 VDD.n1345 185
R815 VDD.n1731 VDD.n1730 185
R816 VDD.n1730 VDD.n1729 185
R817 VDD.n1350 VDD.n1349 185
R818 VDD.n1351 VDD.n1350 185
R819 VDD.n1720 VDD.n1719 185
R820 VDD.n1721 VDD.n1720 185
R821 VDD.n1358 VDD.n1357 185
R822 VDD.n1712 VDD.n1357 185
R823 VDD.n1715 VDD.n1714 185
R824 VDD.n1714 VDD.n1713 185
R825 VDD.n1361 VDD.n1360 185
R826 VDD.n1362 VDD.n1361 185
R827 VDD.n1703 VDD.n1702 185
R828 VDD.n1704 VDD.n1703 185
R829 VDD.n1370 VDD.n1369 185
R830 VDD.n1369 VDD.n1368 185
R831 VDD.n1698 VDD.n1697 185
R832 VDD.n1697 VDD.n1696 185
R833 VDD.n1373 VDD.n1372 185
R834 VDD.n1374 VDD.n1373 185
R835 VDD.n1687 VDD.n1686 185
R836 VDD.n1688 VDD.n1687 185
R837 VDD.n1381 VDD.n1380 185
R838 VDD.n1679 VDD.n1380 185
R839 VDD.n1682 VDD.n1681 185
R840 VDD.n1681 VDD.n1680 185
R841 VDD.n1384 VDD.n1383 185
R842 VDD.n1385 VDD.n1384 185
R843 VDD.n1670 VDD.n1669 185
R844 VDD.n1671 VDD.n1670 185
R845 VDD.n1393 VDD.n1392 185
R846 VDD.n1392 VDD.n1391 185
R847 VDD.n1665 VDD.n1664 185
R848 VDD.n1664 VDD.n1663 185
R849 VDD.n1396 VDD.n1395 185
R850 VDD.n1397 VDD.n1396 185
R851 VDD.n1654 VDD.n1653 185
R852 VDD.n1655 VDD.n1654 185
R853 VDD.n1404 VDD.n1403 185
R854 VDD.n1646 VDD.n1403 185
R855 VDD.n1649 VDD.n1648 185
R856 VDD.n1648 VDD.n1647 185
R857 VDD.n1407 VDD.n1406 185
R858 VDD.n1408 VDD.n1407 185
R859 VDD.n1637 VDD.n1636 185
R860 VDD.n1638 VDD.n1637 185
R861 VDD.n1416 VDD.n1415 185
R862 VDD.n1415 VDD.n1414 185
R863 VDD.n1632 VDD.n1631 185
R864 VDD.n1631 VDD.n1630 185
R865 VDD.n1419 VDD.n1418 185
R866 VDD.n1420 VDD.n1419 185
R867 VDD.n1621 VDD.n1620 185
R868 VDD.n1622 VDD.n1621 185
R869 VDD.n1428 VDD.n1427 185
R870 VDD.n1427 VDD.n1426 185
R871 VDD.n1616 VDD.n1615 185
R872 VDD.n1615 VDD.n1614 185
R873 VDD.n1431 VDD.n1430 185
R874 VDD.t17 VDD.n1431 185
R875 VDD.n1605 VDD.n1604 185
R876 VDD.n1606 VDD.n1605 185
R877 VDD.n1439 VDD.n1438 185
R878 VDD.n1438 VDD.n1437 185
R879 VDD.n1600 VDD.n1599 185
R880 VDD.n1599 VDD.n1598 185
R881 VDD.n1442 VDD.n1441 185
R882 VDD.n1443 VDD.n1442 185
R883 VDD.n1587 VDD.n1586 185
R884 VDD.n1585 VDD.n1469 185
R885 VDD.n1471 VDD.n1468 185
R886 VDD.n1589 VDD.n1468 185
R887 VDD.n1581 VDD.n1473 185
R888 VDD.n1580 VDD.n1474 185
R889 VDD.n1579 VDD.n1475 185
R890 VDD.n1571 VDD.n1476 185
R891 VDD.n1575 VDD.n1572 185
R892 VDD.n1570 VDD.n1478 185
R893 VDD.n1569 VDD.n1479 185
R894 VDD.n1482 VDD.n1480 185
R895 VDD.n1565 VDD.n1483 185
R896 VDD.n1564 VDD.n1484 185
R897 VDD.n1563 VDD.n1485 185
R898 VDD.n1488 VDD.n1486 185
R899 VDD.n1559 VDD.n1489 185
R900 VDD.n1558 VDD.n1490 185
R901 VDD.n1557 VDD.n1491 185
R902 VDD.n1554 VDD.n1496 185
R903 VDD.n1553 VDD.n1497 185
R904 VDD.n1552 VDD.n1498 185
R905 VDD.n1500 VDD.n1499 185
R906 VDD.n1548 VDD.n1502 185
R907 VDD.n1547 VDD.n1503 185
R908 VDD.n1546 VDD.n1504 185
R909 VDD.n1506 VDD.n1505 185
R910 VDD.n1542 VDD.n1508 185
R911 VDD.n1541 VDD.n1509 185
R912 VDD.n1537 VDD.n1510 185
R913 VDD.n1512 VDD.n1511 185
R914 VDD.n1533 VDD.n1514 185
R915 VDD.n1532 VDD.n1515 185
R916 VDD.n1531 VDD.n1516 185
R917 VDD.n1518 VDD.n1517 185
R918 VDD.n1527 VDD.n1520 185
R919 VDD.n1526 VDD.n1521 185
R920 VDD.n1525 VDD.n1522 185
R921 VDD.n1523 VDD.n1450 185
R922 VDD.n1592 VDD.n1591 185
R923 VDD.n2081 VDD.n1198 185
R924 VDD.n2086 VDD.n2085 185
R925 VDD.n2088 VDD.n2087 185
R926 VDD.n2090 VDD.n2089 185
R927 VDD.n2092 VDD.n2091 185
R928 VDD.n2094 VDD.n2093 185
R929 VDD.n2096 VDD.n2095 185
R930 VDD.n2098 VDD.n2097 185
R931 VDD.n2100 VDD.n2099 185
R932 VDD.n2102 VDD.n2101 185
R933 VDD.n2104 VDD.n2103 185
R934 VDD.n2109 VDD.n2108 185
R935 VDD.n2111 VDD.n2110 185
R936 VDD.n2113 VDD.n2112 185
R937 VDD.n2115 VDD.n2114 185
R938 VDD.n2117 VDD.n2116 185
R939 VDD.n2119 VDD.n2118 185
R940 VDD.n2121 VDD.n2120 185
R941 VDD.n2123 VDD.n2122 185
R942 VDD.n2125 VDD.n2124 185
R943 VDD.n2127 VDD.n2126 185
R944 VDD.n2132 VDD.n2131 185
R945 VDD.n2134 VDD.n2133 185
R946 VDD.n2136 VDD.n2135 185
R947 VDD.n2138 VDD.n2137 185
R948 VDD.n2140 VDD.n2139 185
R949 VDD.n2142 VDD.n2141 185
R950 VDD.n2144 VDD.n2143 185
R951 VDD.n2146 VDD.n2145 185
R952 VDD.n2149 VDD.n2148 185
R953 VDD.n2147 VDD.n1167 185
R954 VDD.n2154 VDD.n2153 185
R955 VDD.n2156 VDD.n2155 185
R956 VDD.n2158 VDD.n2157 185
R957 VDD.n2160 VDD.n2159 185
R958 VDD.n2161 VDD.n1161 185
R959 VDD.n2163 VDD.n2162 185
R960 VDD.n1141 VDD.n1139 185
R961 VDD.n2167 VDD.n2166 185
R962 VDD.n2166 VDD.n2165 185
R963 VDD.n1967 VDD.n1966 185
R964 VDD.n1966 VDD.n1142 185
R965 VDD.n1965 VDD.n1200 185
R966 VDD.n1965 VDD.n1964 185
R967 VDD.n1210 VDD.n1201 185
R968 VDD.n1202 VDD.n1201 185
R969 VDD.n1954 VDD.n1953 185
R970 VDD.n1955 VDD.n1954 185
R971 VDD.n1209 VDD.n1208 185
R972 VDD.n1208 VDD.t28 185
R973 VDD.n1948 VDD.n1947 185
R974 VDD.n1947 VDD.n1946 185
R975 VDD.n1213 VDD.n1212 185
R976 VDD.n1214 VDD.n1213 185
R977 VDD.n1937 VDD.n1936 185
R978 VDD.n1938 VDD.n1937 185
R979 VDD.n1222 VDD.n1221 185
R980 VDD.n1221 VDD.n1220 185
R981 VDD.n1932 VDD.n1931 185
R982 VDD.n1931 VDD.n1930 185
R983 VDD.n1225 VDD.n1224 185
R984 VDD.n1226 VDD.n1225 185
R985 VDD.n1921 VDD.n1920 185
R986 VDD.n1922 VDD.n1921 185
R987 VDD.n1234 VDD.n1233 185
R988 VDD.n1233 VDD.n1232 185
R989 VDD.n1916 VDD.n1915 185
R990 VDD.n1915 VDD.n1914 185
R991 VDD.n1237 VDD.n1236 185
R992 VDD.n1238 VDD.n1237 185
R993 VDD.n1905 VDD.n1904 185
R994 VDD.n1906 VDD.n1905 185
R995 VDD.n1246 VDD.n1245 185
R996 VDD.n1245 VDD.n1244 185
R997 VDD.n1900 VDD.n1899 185
R998 VDD.n1899 VDD.n1898 185
R999 VDD.n1249 VDD.n1248 185
R1000 VDD.n1250 VDD.n1249 185
R1001 VDD.n1889 VDD.n1888 185
R1002 VDD.n1890 VDD.n1889 185
R1003 VDD.n1258 VDD.n1257 185
R1004 VDD.n1257 VDD.n1256 185
R1005 VDD.n1884 VDD.n1883 185
R1006 VDD.n1883 VDD.n1882 185
R1007 VDD.n1261 VDD.n1260 185
R1008 VDD.n1262 VDD.n1261 185
R1009 VDD.n1873 VDD.n1872 185
R1010 VDD.n1874 VDD.n1873 185
R1011 VDD.n1270 VDD.n1269 185
R1012 VDD.n1269 VDD.n1268 185
R1013 VDD.n1868 VDD.n1867 185
R1014 VDD.n1867 VDD.n1866 185
R1015 VDD.n1273 VDD.n1272 185
R1016 VDD.n1274 VDD.n1273 185
R1017 VDD.n1857 VDD.n1856 185
R1018 VDD.n1858 VDD.n1857 185
R1019 VDD.n1282 VDD.n1281 185
R1020 VDD.n1281 VDD.n1280 185
R1021 VDD.n1852 VDD.n1851 185
R1022 VDD.n1851 VDD.n1850 185
R1023 VDD.n1285 VDD.n1284 185
R1024 VDD.n1286 VDD.n1285 185
R1025 VDD.n1841 VDD.n1840 185
R1026 VDD.n1842 VDD.n1841 185
R1027 VDD.n1294 VDD.n1293 185
R1028 VDD.n1293 VDD.n1292 185
R1029 VDD.n1836 VDD.n1835 185
R1030 VDD.n1835 VDD.n1834 185
R1031 VDD.n1297 VDD.n1296 185
R1032 VDD.n1298 VDD.n1297 185
R1033 VDD.n1825 VDD.n1824 185
R1034 VDD.n1826 VDD.n1825 185
R1035 VDD.n1306 VDD.n1305 185
R1036 VDD.n1305 VDD.n1304 185
R1037 VDD.n1820 VDD.n1819 185
R1038 VDD.n1819 VDD.n1818 185
R1039 VDD.n1309 VDD.n1308 185
R1040 VDD.n1310 VDD.n1309 185
R1041 VDD.n1809 VDD.n1808 185
R1042 VDD.n1810 VDD.n1809 185
R1043 VDD.n1318 VDD.n1317 185
R1044 VDD.n1317 VDD.n1316 185
R1045 VDD.n1804 VDD.n1803 185
R1046 VDD.n1803 VDD.n1802 185
R1047 VDD.n1321 VDD.n1320 185
R1048 VDD.n1322 VDD.n1321 185
R1049 VDD.n1761 VDD.n1760 185
R1050 VDD.n1762 VDD.n1761 185
R1051 VDD.n1330 VDD.n1329 185
R1052 VDD.n1329 VDD.n1328 185
R1053 VDD.n1756 VDD.n1755 185
R1054 VDD.n1755 VDD.n1754 185
R1055 VDD.n1333 VDD.n1332 185
R1056 VDD.n1745 VDD.n1333 185
R1057 VDD.n1744 VDD.n1743 185
R1058 VDD.n1746 VDD.n1744 185
R1059 VDD.n1341 VDD.n1340 185
R1060 VDD.n1340 VDD.n1339 185
R1061 VDD.n1739 VDD.n1738 185
R1062 VDD.n1738 VDD.n1737 185
R1063 VDD.n1344 VDD.n1343 185
R1064 VDD.n1345 VDD.n1344 185
R1065 VDD.n1728 VDD.n1727 185
R1066 VDD.n1729 VDD.n1728 185
R1067 VDD.n1353 VDD.n1352 185
R1068 VDD.n1352 VDD.n1351 185
R1069 VDD.n1723 VDD.n1722 185
R1070 VDD.n1722 VDD.n1721 185
R1071 VDD.n1356 VDD.n1355 185
R1072 VDD.n1712 VDD.n1356 185
R1073 VDD.n1711 VDD.n1710 185
R1074 VDD.n1713 VDD.n1711 185
R1075 VDD.n1364 VDD.n1363 185
R1076 VDD.n1363 VDD.n1362 185
R1077 VDD.n1706 VDD.n1705 185
R1078 VDD.n1705 VDD.n1704 185
R1079 VDD.n1367 VDD.n1366 185
R1080 VDD.n1368 VDD.n1367 185
R1081 VDD.n1695 VDD.n1694 185
R1082 VDD.n1696 VDD.n1695 185
R1083 VDD.n1376 VDD.n1375 185
R1084 VDD.n1375 VDD.n1374 185
R1085 VDD.n1690 VDD.n1689 185
R1086 VDD.n1689 VDD.n1688 185
R1087 VDD.n1379 VDD.n1378 185
R1088 VDD.n1679 VDD.n1379 185
R1089 VDD.n1678 VDD.n1677 185
R1090 VDD.n1680 VDD.n1678 185
R1091 VDD.n1387 VDD.n1386 185
R1092 VDD.n1386 VDD.n1385 185
R1093 VDD.n1673 VDD.n1672 185
R1094 VDD.n1672 VDD.n1671 185
R1095 VDD.n1390 VDD.n1389 185
R1096 VDD.n1391 VDD.n1390 185
R1097 VDD.n1662 VDD.n1661 185
R1098 VDD.n1663 VDD.n1662 185
R1099 VDD.n1399 VDD.n1398 185
R1100 VDD.n1398 VDD.n1397 185
R1101 VDD.n1657 VDD.n1656 185
R1102 VDD.n1656 VDD.n1655 185
R1103 VDD.n1402 VDD.n1401 185
R1104 VDD.n1646 VDD.n1402 185
R1105 VDD.n1645 VDD.n1644 185
R1106 VDD.n1647 VDD.n1645 185
R1107 VDD.n1410 VDD.n1409 185
R1108 VDD.n1409 VDD.n1408 185
R1109 VDD.n1640 VDD.n1639 185
R1110 VDD.n1639 VDD.n1638 185
R1111 VDD.n1413 VDD.n1412 185
R1112 VDD.n1414 VDD.n1413 185
R1113 VDD.n1629 VDD.n1628 185
R1114 VDD.n1630 VDD.n1629 185
R1115 VDD.n1422 VDD.n1421 185
R1116 VDD.n1421 VDD.n1420 185
R1117 VDD.n1624 VDD.n1623 185
R1118 VDD.n1623 VDD.n1622 185
R1119 VDD.n1425 VDD.n1424 185
R1120 VDD.n1426 VDD.n1425 185
R1121 VDD.n1613 VDD.n1612 185
R1122 VDD.n1614 VDD.n1613 185
R1123 VDD.n1433 VDD.n1432 185
R1124 VDD.n1432 VDD.t17 185
R1125 VDD.n1608 VDD.n1607 185
R1126 VDD.n1607 VDD.n1606 185
R1127 VDD.n1436 VDD.n1435 185
R1128 VDD.n1437 VDD.n1436 185
R1129 VDD.n1597 VDD.n1596 185
R1130 VDD.n1598 VDD.n1597 185
R1131 VDD.n1445 VDD.n1444 185
R1132 VDD.n1444 VDD.n1443 185
R1133 VDD.n2646 VDD.n745 185
R1134 VDD.n745 VDD.n708 185
R1135 VDD.n2648 VDD.n2647 185
R1136 VDD.n2649 VDD.n2648 185
R1137 VDD.n746 VDD.n744 185
R1138 VDD.n744 VDD.n741 185
R1139 VDD.n2589 VDD.n2588 185
R1140 VDD.n2590 VDD.n2589 185
R1141 VDD.n2587 VDD.n754 185
R1142 VDD.n754 VDD.n751 185
R1143 VDD.n2586 VDD.n2585 185
R1144 VDD.n2585 VDD.n2584 185
R1145 VDD.n756 VDD.n755 185
R1146 VDD.n2399 VDD.n756 185
R1147 VDD.n2572 VDD.n2571 185
R1148 VDD.n2573 VDD.n2572 185
R1149 VDD.n2570 VDD.n766 185
R1150 VDD.n766 VDD.n763 185
R1151 VDD.n2569 VDD.n2568 185
R1152 VDD.n2568 VDD.n2567 185
R1153 VDD.n768 VDD.n767 185
R1154 VDD.n769 VDD.n768 185
R1155 VDD.n2560 VDD.n2559 185
R1156 VDD.n2561 VDD.n2560 185
R1157 VDD.n2558 VDD.n778 185
R1158 VDD.n778 VDD.n775 185
R1159 VDD.n2557 VDD.n2556 185
R1160 VDD.n2556 VDD.n2555 185
R1161 VDD.n780 VDD.n779 185
R1162 VDD.n781 VDD.n780 185
R1163 VDD.n2548 VDD.n2547 185
R1164 VDD.n2549 VDD.n2548 185
R1165 VDD.n2546 VDD.n790 185
R1166 VDD.n790 VDD.n787 185
R1167 VDD.n2545 VDD.n2544 185
R1168 VDD.n2544 VDD.n2543 185
R1169 VDD.n792 VDD.n791 185
R1170 VDD.n793 VDD.n792 185
R1171 VDD.n2536 VDD.n2535 185
R1172 VDD.n2537 VDD.n2536 185
R1173 VDD.n2534 VDD.n802 185
R1174 VDD.n802 VDD.n799 185
R1175 VDD.n2533 VDD.n2532 185
R1176 VDD.n2532 VDD.n2531 185
R1177 VDD.n804 VDD.n803 185
R1178 VDD.n813 VDD.n804 185
R1179 VDD.n2524 VDD.n2523 185
R1180 VDD.n2525 VDD.n2524 185
R1181 VDD.n2522 VDD.n814 185
R1182 VDD.n814 VDD.n810 185
R1183 VDD.n2521 VDD.n2520 185
R1184 VDD.n2520 VDD.n2519 185
R1185 VDD.n816 VDD.n815 185
R1186 VDD.n817 VDD.n816 185
R1187 VDD.n2512 VDD.n2511 185
R1188 VDD.n2513 VDD.n2512 185
R1189 VDD.n2510 VDD.n826 185
R1190 VDD.n826 VDD.n823 185
R1191 VDD.n2509 VDD.n2508 185
R1192 VDD.n2508 VDD.n2507 185
R1193 VDD.n828 VDD.n827 185
R1194 VDD.n829 VDD.n828 185
R1195 VDD.n2500 VDD.n2499 185
R1196 VDD.n2501 VDD.n2500 185
R1197 VDD.n2498 VDD.n838 185
R1198 VDD.n838 VDD.n835 185
R1199 VDD.n2497 VDD.n2496 185
R1200 VDD.n2496 VDD.n2495 185
R1201 VDD.n840 VDD.n839 185
R1202 VDD.n849 VDD.n840 185
R1203 VDD.n2488 VDD.n2487 185
R1204 VDD.n2489 VDD.n2488 185
R1205 VDD.n2486 VDD.n850 185
R1206 VDD.n850 VDD.n846 185
R1207 VDD.n2485 VDD.n2484 185
R1208 VDD.n2484 VDD.n2483 185
R1209 VDD.n852 VDD.n851 185
R1210 VDD.n853 VDD.n852 185
R1211 VDD.n2476 VDD.n2475 185
R1212 VDD.n2477 VDD.n2476 185
R1213 VDD.n2474 VDD.n862 185
R1214 VDD.n862 VDD.n859 185
R1215 VDD.n2473 VDD.n2472 185
R1216 VDD.n2472 VDD.n2471 185
R1217 VDD.n864 VDD.n863 185
R1218 VDD.n865 VDD.n864 185
R1219 VDD.n2464 VDD.n2463 185
R1220 VDD.n2465 VDD.n2464 185
R1221 VDD.n2462 VDD.n874 185
R1222 VDD.n874 VDD.n871 185
R1223 VDD.n2461 VDD.n2460 185
R1224 VDD.n2460 VDD.t100 185
R1225 VDD.n876 VDD.n875 185
R1226 VDD.n877 VDD.n876 185
R1227 VDD.n2329 VDD.n2328 185
R1228 VDD.n2330 VDD.n2329 185
R1229 VDD.n2327 VDD.n890 185
R1230 VDD.n890 VDD.n887 185
R1231 VDD.n2326 VDD.n2325 185
R1232 VDD.n2325 VDD.n2324 185
R1233 VDD.n892 VDD.n891 185
R1234 VDD.n893 VDD.n892 185
R1235 VDD.n2312 VDD.n2311 185
R1236 VDD.n2313 VDD.n2312 185
R1237 VDD.n2310 VDD.n903 185
R1238 VDD.n903 VDD.n900 185
R1239 VDD.n2309 VDD.n2308 185
R1240 VDD.n2308 VDD.n2307 185
R1241 VDD.n905 VDD.n904 185
R1242 VDD.n906 VDD.n905 185
R1243 VDD.n2300 VDD.n2299 185
R1244 VDD.n2301 VDD.n2300 185
R1245 VDD.n2298 VDD.n915 185
R1246 VDD.n915 VDD.n912 185
R1247 VDD.n2297 VDD.n2296 185
R1248 VDD.n2296 VDD.n2295 185
R1249 VDD.n917 VDD.n916 185
R1250 VDD.n926 VDD.n917 185
R1251 VDD.n2288 VDD.n2287 185
R1252 VDD.n2289 VDD.n2288 185
R1253 VDD.n2286 VDD.n927 185
R1254 VDD.n927 VDD.n923 185
R1255 VDD.n2285 VDD.n2284 185
R1256 VDD.n2284 VDD.n2283 185
R1257 VDD.n929 VDD.n928 185
R1258 VDD.n930 VDD.n929 185
R1259 VDD.n2276 VDD.n2275 185
R1260 VDD.n2277 VDD.n2276 185
R1261 VDD.n2274 VDD.n939 185
R1262 VDD.n939 VDD.n936 185
R1263 VDD.n2273 VDD.n2272 185
R1264 VDD.n2272 VDD.n2271 185
R1265 VDD.n941 VDD.n940 185
R1266 VDD.n942 VDD.n941 185
R1267 VDD.n2264 VDD.n2263 185
R1268 VDD.n2265 VDD.n2264 185
R1269 VDD.n2262 VDD.n951 185
R1270 VDD.n951 VDD.n948 185
R1271 VDD.n2261 VDD.n2260 185
R1272 VDD.n2260 VDD.n2259 185
R1273 VDD.n953 VDD.n952 185
R1274 VDD.n962 VDD.n953 185
R1275 VDD.n2252 VDD.n2251 185
R1276 VDD.n2253 VDD.n2252 185
R1277 VDD.n2250 VDD.n963 185
R1278 VDD.n963 VDD.n959 185
R1279 VDD.n2249 VDD.n2248 185
R1280 VDD.n2248 VDD.n2247 185
R1281 VDD.n965 VDD.n964 185
R1282 VDD.n966 VDD.n965 185
R1283 VDD.n2240 VDD.n2239 185
R1284 VDD.n2241 VDD.n2240 185
R1285 VDD.n2238 VDD.n975 185
R1286 VDD.n975 VDD.n972 185
R1287 VDD.n2237 VDD.n2236 185
R1288 VDD.n2236 VDD.n2235 185
R1289 VDD.n977 VDD.n976 185
R1290 VDD.n978 VDD.n977 185
R1291 VDD.n2228 VDD.n2227 185
R1292 VDD.n2229 VDD.n2228 185
R1293 VDD.n2226 VDD.n987 185
R1294 VDD.n987 VDD.n984 185
R1295 VDD.n2225 VDD.n2224 185
R1296 VDD.n2224 VDD.n2223 185
R1297 VDD.n989 VDD.n988 185
R1298 VDD.n997 VDD.n989 185
R1299 VDD.n2216 VDD.n2215 185
R1300 VDD.n2217 VDD.n2216 185
R1301 VDD.n2214 VDD.n998 185
R1302 VDD.n1004 VDD.n998 185
R1303 VDD.n2213 VDD.n2212 185
R1304 VDD.n2212 VDD.n2211 185
R1305 VDD.n1000 VDD.n999 185
R1306 VDD.n1001 VDD.n1000 185
R1307 VDD.n2204 VDD.n2203 185
R1308 VDD.n2205 VDD.n2204 185
R1309 VDD.n2202 VDD.n1011 185
R1310 VDD.n1011 VDD.n1008 185
R1311 VDD.n2201 VDD.n2200 185
R1312 VDD.n2200 VDD.n2199 185
R1313 VDD.n1013 VDD.n1012 185
R1314 VDD.n1014 VDD.n1013 185
R1315 VDD.n2191 VDD.n2190 185
R1316 VDD.n2189 VDD.n1044 185
R1317 VDD.n2188 VDD.n1043 185
R1318 VDD.n2193 VDD.n1043 185
R1319 VDD.n2187 VDD.n2186 185
R1320 VDD.n2185 VDD.n2184 185
R1321 VDD.n2183 VDD.n2182 185
R1322 VDD.n2181 VDD.n2180 185
R1323 VDD.n2179 VDD.n2178 185
R1324 VDD.n2177 VDD.n2176 185
R1325 VDD.n2175 VDD.n2174 185
R1326 VDD.n2173 VDD.n2172 185
R1327 VDD.n2171 VDD.n2170 185
R1328 VDD.n1136 VDD.n1135 185
R1329 VDD.n1134 VDD.n1133 185
R1330 VDD.n1132 VDD.n1131 185
R1331 VDD.n1130 VDD.n1129 185
R1332 VDD.n1128 VDD.n1127 185
R1333 VDD.n1126 VDD.n1125 185
R1334 VDD.n1124 VDD.n1123 185
R1335 VDD.n1122 VDD.n1121 185
R1336 VDD.n1120 VDD.n1119 185
R1337 VDD.n1118 VDD.n1117 185
R1338 VDD.n1116 VDD.n1115 185
R1339 VDD.n1114 VDD.n1030 185
R1340 VDD.n2193 VDD.n1030 185
R1341 VDD.n2598 VDD.n2597 185
R1342 VDD.n2600 VDD.n2599 185
R1343 VDD.n2602 VDD.n2601 185
R1344 VDD.n2605 VDD.n2604 185
R1345 VDD.n2607 VDD.n2606 185
R1346 VDD.n2609 VDD.n2608 185
R1347 VDD.n2611 VDD.n2610 185
R1348 VDD.n2613 VDD.n2612 185
R1349 VDD.n2615 VDD.n2614 185
R1350 VDD.n2617 VDD.n2616 185
R1351 VDD.n2619 VDD.n2618 185
R1352 VDD.n2621 VDD.n2620 185
R1353 VDD.n2623 VDD.n2622 185
R1354 VDD.n2625 VDD.n2624 185
R1355 VDD.n2627 VDD.n2626 185
R1356 VDD.n2629 VDD.n2628 185
R1357 VDD.n2631 VDD.n2630 185
R1358 VDD.n2633 VDD.n2632 185
R1359 VDD.n2635 VDD.n2634 185
R1360 VDD.n2637 VDD.n2636 185
R1361 VDD.n2639 VDD.n2638 185
R1362 VDD.n2641 VDD.n2640 185
R1363 VDD.n2643 VDD.n2642 185
R1364 VDD.n2645 VDD.n2644 185
R1365 VDD.n2596 VDD.n2595 185
R1366 VDD.n2596 VDD.n708 185
R1367 VDD.n2594 VDD.n742 185
R1368 VDD.n2649 VDD.n742 185
R1369 VDD.n2593 VDD.n2592 185
R1370 VDD.n2592 VDD.n741 185
R1371 VDD.n2591 VDD.n749 185
R1372 VDD.n2591 VDD.n2590 185
R1373 VDD.n883 VDD.n750 185
R1374 VDD.n751 VDD.n750 185
R1375 VDD.n884 VDD.n757 185
R1376 VDD.n2584 VDD.n757 185
R1377 VDD.n2401 VDD.n2400 185
R1378 VDD.n2400 VDD.n2399 185
R1379 VDD.n2402 VDD.n764 185
R1380 VDD.n2573 VDD.n764 185
R1381 VDD.n2404 VDD.n2403 185
R1382 VDD.n2403 VDD.n763 185
R1383 VDD.n2405 VDD.n770 185
R1384 VDD.n2567 VDD.n770 185
R1385 VDD.n2407 VDD.n2406 185
R1386 VDD.n2406 VDD.n769 185
R1387 VDD.n2408 VDD.n776 185
R1388 VDD.n2561 VDD.n776 185
R1389 VDD.n2410 VDD.n2409 185
R1390 VDD.n2409 VDD.n775 185
R1391 VDD.n2411 VDD.n782 185
R1392 VDD.n2555 VDD.n782 185
R1393 VDD.n2413 VDD.n2412 185
R1394 VDD.n2412 VDD.n781 185
R1395 VDD.n2414 VDD.n788 185
R1396 VDD.n2549 VDD.n788 185
R1397 VDD.n2416 VDD.n2415 185
R1398 VDD.n2415 VDD.n787 185
R1399 VDD.n2417 VDD.n794 185
R1400 VDD.n2543 VDD.n794 185
R1401 VDD.n2419 VDD.n2418 185
R1402 VDD.n2418 VDD.n793 185
R1403 VDD.n2420 VDD.n800 185
R1404 VDD.n2537 VDD.n800 185
R1405 VDD.n2422 VDD.n2421 185
R1406 VDD.n2421 VDD.n799 185
R1407 VDD.n2423 VDD.n805 185
R1408 VDD.n2531 VDD.n805 185
R1409 VDD.n2425 VDD.n2424 185
R1410 VDD.n2424 VDD.n813 185
R1411 VDD.n2426 VDD.n811 185
R1412 VDD.n2525 VDD.n811 185
R1413 VDD.n2428 VDD.n2427 185
R1414 VDD.n2427 VDD.n810 185
R1415 VDD.n2429 VDD.n818 185
R1416 VDD.n2519 VDD.n818 185
R1417 VDD.n2431 VDD.n2430 185
R1418 VDD.n2430 VDD.n817 185
R1419 VDD.n2432 VDD.n824 185
R1420 VDD.n2513 VDD.n824 185
R1421 VDD.n2434 VDD.n2433 185
R1422 VDD.n2433 VDD.n823 185
R1423 VDD.n2435 VDD.n830 185
R1424 VDD.n2507 VDD.n830 185
R1425 VDD.n2437 VDD.n2436 185
R1426 VDD.n2436 VDD.n829 185
R1427 VDD.n2438 VDD.n836 185
R1428 VDD.n2501 VDD.n836 185
R1429 VDD.n2440 VDD.n2439 185
R1430 VDD.n2439 VDD.n835 185
R1431 VDD.n2441 VDD.n841 185
R1432 VDD.n2495 VDD.n841 185
R1433 VDD.n2443 VDD.n2442 185
R1434 VDD.n2442 VDD.n849 185
R1435 VDD.n2444 VDD.n847 185
R1436 VDD.n2489 VDD.n847 185
R1437 VDD.n2446 VDD.n2445 185
R1438 VDD.n2445 VDD.n846 185
R1439 VDD.n2447 VDD.n854 185
R1440 VDD.n2483 VDD.n854 185
R1441 VDD.n2449 VDD.n2448 185
R1442 VDD.n2448 VDD.n853 185
R1443 VDD.n2450 VDD.n860 185
R1444 VDD.n2477 VDD.n860 185
R1445 VDD.n2452 VDD.n2451 185
R1446 VDD.n2451 VDD.n859 185
R1447 VDD.n2453 VDD.n866 185
R1448 VDD.n2471 VDD.n866 185
R1449 VDD.n2455 VDD.n2454 185
R1450 VDD.n2454 VDD.n865 185
R1451 VDD.n2456 VDD.n872 185
R1452 VDD.n2465 VDD.n872 185
R1453 VDD.n2457 VDD.n881 185
R1454 VDD.n881 VDD.n871 185
R1455 VDD.n2459 VDD.n2458 185
R1456 VDD.t100 VDD.n2459 185
R1457 VDD.n882 VDD.n880 185
R1458 VDD.n880 VDD.n877 185
R1459 VDD.n1048 VDD.n888 185
R1460 VDD.n2330 VDD.n888 185
R1461 VDD.n1050 VDD.n1049 185
R1462 VDD.n1049 VDD.n887 185
R1463 VDD.n1051 VDD.n894 185
R1464 VDD.n2324 VDD.n894 185
R1465 VDD.n1053 VDD.n1052 185
R1466 VDD.n1052 VDD.n893 185
R1467 VDD.n1054 VDD.n901 185
R1468 VDD.n2313 VDD.n901 185
R1469 VDD.n1056 VDD.n1055 185
R1470 VDD.n1055 VDD.n900 185
R1471 VDD.n1057 VDD.n907 185
R1472 VDD.n2307 VDD.n907 185
R1473 VDD.n1059 VDD.n1058 185
R1474 VDD.n1058 VDD.n906 185
R1475 VDD.n1060 VDD.n913 185
R1476 VDD.n2301 VDD.n913 185
R1477 VDD.n1062 VDD.n1061 185
R1478 VDD.n1061 VDD.n912 185
R1479 VDD.n1063 VDD.n918 185
R1480 VDD.n2295 VDD.n918 185
R1481 VDD.n1065 VDD.n1064 185
R1482 VDD.n1064 VDD.n926 185
R1483 VDD.n1066 VDD.n924 185
R1484 VDD.n2289 VDD.n924 185
R1485 VDD.n1068 VDD.n1067 185
R1486 VDD.n1067 VDD.n923 185
R1487 VDD.n1069 VDD.n931 185
R1488 VDD.n2283 VDD.n931 185
R1489 VDD.n1071 VDD.n1070 185
R1490 VDD.n1070 VDD.n930 185
R1491 VDD.n1072 VDD.n937 185
R1492 VDD.n2277 VDD.n937 185
R1493 VDD.n1074 VDD.n1073 185
R1494 VDD.n1073 VDD.n936 185
R1495 VDD.n1075 VDD.n943 185
R1496 VDD.n2271 VDD.n943 185
R1497 VDD.n1077 VDD.n1076 185
R1498 VDD.n1076 VDD.n942 185
R1499 VDD.n1078 VDD.n949 185
R1500 VDD.n2265 VDD.n949 185
R1501 VDD.n1080 VDD.n1079 185
R1502 VDD.n1079 VDD.n948 185
R1503 VDD.n1081 VDD.n954 185
R1504 VDD.n2259 VDD.n954 185
R1505 VDD.n1083 VDD.n1082 185
R1506 VDD.n1082 VDD.n962 185
R1507 VDD.n1084 VDD.n960 185
R1508 VDD.n2253 VDD.n960 185
R1509 VDD.n1086 VDD.n1085 185
R1510 VDD.n1085 VDD.n959 185
R1511 VDD.n1087 VDD.n967 185
R1512 VDD.n2247 VDD.n967 185
R1513 VDD.n1089 VDD.n1088 185
R1514 VDD.n1088 VDD.n966 185
R1515 VDD.n1090 VDD.n973 185
R1516 VDD.n2241 VDD.n973 185
R1517 VDD.n1092 VDD.n1091 185
R1518 VDD.n1091 VDD.n972 185
R1519 VDD.n1093 VDD.n979 185
R1520 VDD.n2235 VDD.n979 185
R1521 VDD.n1095 VDD.n1094 185
R1522 VDD.n1094 VDD.n978 185
R1523 VDD.n1096 VDD.n985 185
R1524 VDD.n2229 VDD.n985 185
R1525 VDD.n1098 VDD.n1097 185
R1526 VDD.n1097 VDD.n984 185
R1527 VDD.n1099 VDD.n990 185
R1528 VDD.n2223 VDD.n990 185
R1529 VDD.n1101 VDD.n1100 185
R1530 VDD.n1100 VDD.n997 185
R1531 VDD.n1102 VDD.n995 185
R1532 VDD.n2217 VDD.n995 185
R1533 VDD.n1104 VDD.n1103 185
R1534 VDD.n1103 VDD.n1004 185
R1535 VDD.n1105 VDD.n1002 185
R1536 VDD.n2211 VDD.n1002 185
R1537 VDD.n1107 VDD.n1106 185
R1538 VDD.n1106 VDD.n1001 185
R1539 VDD.n1108 VDD.n1009 185
R1540 VDD.n2205 VDD.n1009 185
R1541 VDD.n1110 VDD.n1109 185
R1542 VDD.n1109 VDD.n1008 185
R1543 VDD.n1111 VDD.n1015 185
R1544 VDD.n2199 VDD.n1015 185
R1545 VDD.n1113 VDD.n1112 185
R1546 VDD.n1112 VDD.n1014 185
R1547 VDD.n3915 VDD.n3914 185
R1548 VDD.n3916 VDD.n3915 185
R1549 VDD.n162 VDD.n161 185
R1550 VDD.n3917 VDD.n162 185
R1551 VDD.n3920 VDD.n3919 185
R1552 VDD.n3919 VDD.n3918 185
R1553 VDD.n3921 VDD.n156 185
R1554 VDD.n156 VDD.n155 185
R1555 VDD.n3923 VDD.n3922 185
R1556 VDD.t24 VDD.n3923 185
R1557 VDD.n151 VDD.n150 185
R1558 VDD.n3924 VDD.n151 185
R1559 VDD.n3927 VDD.n3926 185
R1560 VDD.n3926 VDD.n3925 185
R1561 VDD.n3928 VDD.n145 185
R1562 VDD.n145 VDD.n144 185
R1563 VDD.n3930 VDD.n3929 185
R1564 VDD.n3931 VDD.n3930 185
R1565 VDD.n140 VDD.n139 185
R1566 VDD.n3932 VDD.n140 185
R1567 VDD.n3935 VDD.n3934 185
R1568 VDD.n3934 VDD.n3933 185
R1569 VDD.n3936 VDD.n134 185
R1570 VDD.n134 VDD.n133 185
R1571 VDD.n3938 VDD.n3937 185
R1572 VDD.n3939 VDD.n3938 185
R1573 VDD.n129 VDD.n128 185
R1574 VDD.n3940 VDD.n129 185
R1575 VDD.n3943 VDD.n3942 185
R1576 VDD.n3942 VDD.n3941 185
R1577 VDD.n3944 VDD.n123 185
R1578 VDD.n123 VDD.n122 185
R1579 VDD.n3946 VDD.n3945 185
R1580 VDD.n3947 VDD.n3946 185
R1581 VDD.n118 VDD.n117 185
R1582 VDD.n3948 VDD.n118 185
R1583 VDD.n3951 VDD.n3950 185
R1584 VDD.n3950 VDD.n3949 185
R1585 VDD.n3952 VDD.n112 185
R1586 VDD.n112 VDD.n111 185
R1587 VDD.n3954 VDD.n3953 185
R1588 VDD.n3955 VDD.n3954 185
R1589 VDD.n107 VDD.n106 185
R1590 VDD.n3956 VDD.n107 185
R1591 VDD.n3959 VDD.n3958 185
R1592 VDD.n3958 VDD.n3957 185
R1593 VDD.n3960 VDD.n101 185
R1594 VDD.n101 VDD.n100 185
R1595 VDD.n3962 VDD.n3961 185
R1596 VDD.n3963 VDD.n3962 185
R1597 VDD.n96 VDD.n95 185
R1598 VDD.n3964 VDD.n96 185
R1599 VDD.n3967 VDD.n3966 185
R1600 VDD.n3966 VDD.n3965 185
R1601 VDD.n3968 VDD.n90 185
R1602 VDD.n90 VDD.n89 185
R1603 VDD.n3970 VDD.n3969 185
R1604 VDD.n3971 VDD.n3970 185
R1605 VDD.n85 VDD.n84 185
R1606 VDD.n3972 VDD.n85 185
R1607 VDD.n3975 VDD.n3974 185
R1608 VDD.n3974 VDD.n3973 185
R1609 VDD.n3976 VDD.n79 185
R1610 VDD.n79 VDD.n78 185
R1611 VDD.n3978 VDD.n3977 185
R1612 VDD.n3979 VDD.n3978 185
R1613 VDD.n74 VDD.n73 185
R1614 VDD.n3980 VDD.n74 185
R1615 VDD.n3983 VDD.n3982 185
R1616 VDD.n3982 VDD.n3981 185
R1617 VDD.n3984 VDD.n68 185
R1618 VDD.n68 VDD.n67 185
R1619 VDD.n3986 VDD.n3985 185
R1620 VDD.n3987 VDD.n3986 185
R1621 VDD.n63 VDD.n62 185
R1622 VDD.n3988 VDD.n63 185
R1623 VDD.n3991 VDD.n3990 185
R1624 VDD.n3990 VDD.n3989 185
R1625 VDD.n3992 VDD.n58 185
R1626 VDD.n58 VDD.n57 185
R1627 VDD.n3994 VDD.n3993 185
R1628 VDD.n3995 VDD.n3994 185
R1629 VDD.n52 VDD.n50 185
R1630 VDD.n3996 VDD.n52 185
R1631 VDD.n3999 VDD.n3998 185
R1632 VDD.n3998 VDD.n3997 185
R1633 VDD.n51 VDD.n49 185
R1634 VDD.n53 VDD.n51 185
R1635 VDD.n3766 VDD.n3765 185
R1636 VDD.n3767 VDD.n3766 185
R1637 VDD.n277 VDD.n276 185
R1638 VDD.n276 VDD.n275 185
R1639 VDD.n3761 VDD.n3760 185
R1640 VDD.n3760 VDD.n3759 185
R1641 VDD.n280 VDD.n279 185
R1642 VDD.n281 VDD.n280 185
R1643 VDD.n3750 VDD.n3749 185
R1644 VDD.n3751 VDD.n3750 185
R1645 VDD.n289 VDD.n288 185
R1646 VDD.n288 VDD.n287 185
R1647 VDD.n3745 VDD.n3744 185
R1648 VDD.n3744 VDD.n3743 185
R1649 VDD.n292 VDD.n291 185
R1650 VDD.n293 VDD.n292 185
R1651 VDD.n3734 VDD.n3733 185
R1652 VDD.n3735 VDD.n3734 185
R1653 VDD.n301 VDD.n300 185
R1654 VDD.n300 VDD.n299 185
R1655 VDD.n3729 VDD.n3728 185
R1656 VDD.n3728 VDD.n3727 185
R1657 VDD.n304 VDD.n303 185
R1658 VDD.n305 VDD.n304 185
R1659 VDD.n3718 VDD.n3717 185
R1660 VDD.n3719 VDD.n3718 185
R1661 VDD.n313 VDD.n312 185
R1662 VDD.n312 VDD.n311 185
R1663 VDD.n3713 VDD.n3712 185
R1664 VDD.n3712 VDD.n3711 185
R1665 VDD.n316 VDD.n315 185
R1666 VDD.n317 VDD.n316 185
R1667 VDD.n3702 VDD.n3701 185
R1668 VDD.n3703 VDD.n3702 185
R1669 VDD.n325 VDD.n324 185
R1670 VDD.n324 VDD.n323 185
R1671 VDD.n3697 VDD.n3696 185
R1672 VDD.n3696 VDD.n3695 185
R1673 VDD.n328 VDD.n327 185
R1674 VDD.n329 VDD.n328 185
R1675 VDD.n3686 VDD.n3685 185
R1676 VDD.n3687 VDD.n3686 185
R1677 VDD.n337 VDD.n336 185
R1678 VDD.n336 VDD.n335 185
R1679 VDD.n3681 VDD.n3680 185
R1680 VDD.n3680 VDD.n3679 185
R1681 VDD.n340 VDD.n339 185
R1682 VDD.n341 VDD.n340 185
R1683 VDD.n3670 VDD.n3669 185
R1684 VDD.n3671 VDD.n3670 185
R1685 VDD.n349 VDD.n348 185
R1686 VDD.n348 VDD.n347 185
R1687 VDD.n3665 VDD.n3664 185
R1688 VDD.n3664 VDD.n3663 185
R1689 VDD.n352 VDD.n351 185
R1690 VDD.n353 VDD.n352 185
R1691 VDD.n3654 VDD.n3653 185
R1692 VDD.n3655 VDD.n3654 185
R1693 VDD.n361 VDD.n360 185
R1694 VDD.n360 VDD.n359 185
R1695 VDD.n3649 VDD.n3648 185
R1696 VDD.n3648 VDD.n3647 185
R1697 VDD.n364 VDD.n363 185
R1698 VDD.n365 VDD.n364 185
R1699 VDD.n3638 VDD.n3637 185
R1700 VDD.n3639 VDD.n3638 185
R1701 VDD.n373 VDD.n372 185
R1702 VDD.n372 VDD.n371 185
R1703 VDD.n3633 VDD.n3632 185
R1704 VDD.n3632 VDD.n3631 185
R1705 VDD.n376 VDD.n375 185
R1706 VDD.n377 VDD.n376 185
R1707 VDD.n3623 VDD.n3622 185
R1708 VDD.t13 VDD.n3623 185
R1709 VDD.n385 VDD.n384 185
R1710 VDD.n384 VDD.n383 185
R1711 VDD.n3618 VDD.n3617 185
R1712 VDD.n3617 VDD.n3616 185
R1713 VDD.n388 VDD.n387 185
R1714 VDD.n389 VDD.n388 185
R1715 VDD.n3607 VDD.n3606 185
R1716 VDD.n3608 VDD.n3607 185
R1717 VDD.n3603 VDD.n395 185
R1718 VDD.n3602 VDD.n3601 185
R1719 VDD.n3599 VDD.n3462 185
R1720 VDD.n3599 VDD.n394 185
R1721 VDD.n3598 VDD.n3597 185
R1722 VDD.n3596 VDD.n3595 185
R1723 VDD.n3594 VDD.n3467 185
R1724 VDD.n3592 VDD.n3591 185
R1725 VDD.n3590 VDD.n3468 185
R1726 VDD.n3589 VDD.n3588 185
R1727 VDD.n3586 VDD.n3475 185
R1728 VDD.n3584 VDD.n3583 185
R1729 VDD.n3582 VDD.n3476 185
R1730 VDD.n3581 VDD.n3580 185
R1731 VDD.n3578 VDD.n3481 185
R1732 VDD.n3576 VDD.n3575 185
R1733 VDD.n3574 VDD.n3482 185
R1734 VDD.n3573 VDD.n3572 185
R1735 VDD.n3570 VDD.n3487 185
R1736 VDD.n3568 VDD.n3567 185
R1737 VDD.n3566 VDD.n3488 185
R1738 VDD.n3565 VDD.n3564 185
R1739 VDD.n3562 VDD.n3496 185
R1740 VDD.n3560 VDD.n3559 185
R1741 VDD.n3558 VDD.n3497 185
R1742 VDD.n3557 VDD.n3556 185
R1743 VDD.n3554 VDD.n3502 185
R1744 VDD.n3552 VDD.n3551 185
R1745 VDD.n3550 VDD.n3503 185
R1746 VDD.n3548 VDD.n3547 185
R1747 VDD.n3545 VDD.n3510 185
R1748 VDD.n3543 VDD.n3542 185
R1749 VDD.n3541 VDD.n3511 185
R1750 VDD.n3540 VDD.n3539 185
R1751 VDD.n3537 VDD.n3516 185
R1752 VDD.n3535 VDD.n3534 185
R1753 VDD.n3533 VDD.n3517 185
R1754 VDD.n3532 VDD.n3531 185
R1755 VDD.n3529 VDD.n3527 185
R1756 VDD.n3522 VDD.n393 185
R1757 VDD.n3840 VDD.n3839 185
R1758 VDD.n3844 VDD.n235 185
R1759 VDD.n3846 VDD.n3845 185
R1760 VDD.n3848 VDD.n233 185
R1761 VDD.n3850 VDD.n3849 185
R1762 VDD.n3851 VDD.n228 185
R1763 VDD.n3853 VDD.n3852 185
R1764 VDD.n3855 VDD.n226 185
R1765 VDD.n3857 VDD.n3856 185
R1766 VDD.n3858 VDD.n218 185
R1767 VDD.n3860 VDD.n3859 185
R1768 VDD.n3862 VDD.n216 185
R1769 VDD.n3864 VDD.n3863 185
R1770 VDD.n3865 VDD.n211 185
R1771 VDD.n3867 VDD.n3866 185
R1772 VDD.n3869 VDD.n209 185
R1773 VDD.n3871 VDD.n3870 185
R1774 VDD.n3872 VDD.n204 185
R1775 VDD.n3874 VDD.n3873 185
R1776 VDD.n3876 VDD.n202 185
R1777 VDD.n3878 VDD.n3877 185
R1778 VDD.n3882 VDD.n197 185
R1779 VDD.n3884 VDD.n3883 185
R1780 VDD.n3886 VDD.n195 185
R1781 VDD.n3888 VDD.n3887 185
R1782 VDD.n3889 VDD.n190 185
R1783 VDD.n3891 VDD.n3890 185
R1784 VDD.n3893 VDD.n188 185
R1785 VDD.n3895 VDD.n3894 185
R1786 VDD.n3896 VDD.n183 185
R1787 VDD.n3898 VDD.n3897 185
R1788 VDD.n3900 VDD.n181 185
R1789 VDD.n3902 VDD.n3901 185
R1790 VDD.n3903 VDD.n174 185
R1791 VDD.n3905 VDD.n3904 185
R1792 VDD.n3907 VDD.n172 185
R1793 VDD.n3909 VDD.n3908 185
R1794 VDD.n3910 VDD.n170 185
R1795 VDD.n3911 VDD.n167 185
R1796 VDD.n167 VDD.n166 185
R1797 VDD.n3835 VDD.n165 185
R1798 VDD.n3916 VDD.n165 185
R1799 VDD.n3834 VDD.n164 185
R1800 VDD.n3917 VDD.n164 185
R1801 VDD.n3833 VDD.n163 185
R1802 VDD.n3918 VDD.n163 185
R1803 VDD.n241 VDD.n240 185
R1804 VDD.n240 VDD.n155 185
R1805 VDD.n3829 VDD.n154 185
R1806 VDD.t24 VDD.n154 185
R1807 VDD.n3828 VDD.n153 185
R1808 VDD.n3924 VDD.n153 185
R1809 VDD.n3827 VDD.n152 185
R1810 VDD.n3925 VDD.n152 185
R1811 VDD.n244 VDD.n243 185
R1812 VDD.n243 VDD.n144 185
R1813 VDD.n3823 VDD.n143 185
R1814 VDD.n3931 VDD.n143 185
R1815 VDD.n3822 VDD.n142 185
R1816 VDD.n3932 VDD.n142 185
R1817 VDD.n3821 VDD.n141 185
R1818 VDD.n3933 VDD.n141 185
R1819 VDD.n247 VDD.n246 185
R1820 VDD.n246 VDD.n133 185
R1821 VDD.n3817 VDD.n132 185
R1822 VDD.n3939 VDD.n132 185
R1823 VDD.n3816 VDD.n131 185
R1824 VDD.n3940 VDD.n131 185
R1825 VDD.n3815 VDD.n130 185
R1826 VDD.n3941 VDD.n130 185
R1827 VDD.n250 VDD.n249 185
R1828 VDD.n249 VDD.n122 185
R1829 VDD.n3811 VDD.n121 185
R1830 VDD.n3947 VDD.n121 185
R1831 VDD.n3810 VDD.n120 185
R1832 VDD.n3948 VDD.n120 185
R1833 VDD.n3809 VDD.n119 185
R1834 VDD.n3949 VDD.n119 185
R1835 VDD.n253 VDD.n252 185
R1836 VDD.n252 VDD.n111 185
R1837 VDD.n3805 VDD.n110 185
R1838 VDD.n3955 VDD.n110 185
R1839 VDD.n3804 VDD.n109 185
R1840 VDD.n3956 VDD.n109 185
R1841 VDD.n3803 VDD.n108 185
R1842 VDD.n3957 VDD.n108 185
R1843 VDD.n256 VDD.n255 185
R1844 VDD.n255 VDD.n100 185
R1845 VDD.n3799 VDD.n99 185
R1846 VDD.n3963 VDD.n99 185
R1847 VDD.n3798 VDD.n98 185
R1848 VDD.n3964 VDD.n98 185
R1849 VDD.n3797 VDD.n97 185
R1850 VDD.n3965 VDD.n97 185
R1851 VDD.n259 VDD.n258 185
R1852 VDD.n258 VDD.n89 185
R1853 VDD.n3793 VDD.n88 185
R1854 VDD.n3971 VDD.n88 185
R1855 VDD.n3792 VDD.n87 185
R1856 VDD.n3972 VDD.n87 185
R1857 VDD.n3791 VDD.n86 185
R1858 VDD.n3973 VDD.n86 185
R1859 VDD.n262 VDD.n261 185
R1860 VDD.n261 VDD.n78 185
R1861 VDD.n3787 VDD.n77 185
R1862 VDD.n3979 VDD.n77 185
R1863 VDD.n3786 VDD.n76 185
R1864 VDD.n3980 VDD.n76 185
R1865 VDD.n3785 VDD.n75 185
R1866 VDD.n3981 VDD.n75 185
R1867 VDD.n265 VDD.n264 185
R1868 VDD.n264 VDD.n67 185
R1869 VDD.n3781 VDD.n66 185
R1870 VDD.n3987 VDD.n66 185
R1871 VDD.n3780 VDD.n65 185
R1872 VDD.n3988 VDD.n65 185
R1873 VDD.n3779 VDD.n64 185
R1874 VDD.n3989 VDD.n64 185
R1875 VDD.n268 VDD.n267 185
R1876 VDD.n267 VDD.n57 185
R1877 VDD.n3775 VDD.n56 185
R1878 VDD.n3995 VDD.n56 185
R1879 VDD.n3774 VDD.n55 185
R1880 VDD.n3996 VDD.n55 185
R1881 VDD.n3773 VDD.n54 185
R1882 VDD.n3997 VDD.n54 185
R1883 VDD.n274 VDD.n270 185
R1884 VDD.n274 VDD.n53 185
R1885 VDD.n3769 VDD.n3768 185
R1886 VDD.n3768 VDD.n3767 185
R1887 VDD.n273 VDD.n272 185
R1888 VDD.n275 VDD.n273 185
R1889 VDD.n3758 VDD.n3757 185
R1890 VDD.n3759 VDD.n3758 185
R1891 VDD.n283 VDD.n282 185
R1892 VDD.n282 VDD.n281 185
R1893 VDD.n3753 VDD.n3752 185
R1894 VDD.n3752 VDD.n3751 185
R1895 VDD.n286 VDD.n285 185
R1896 VDD.n287 VDD.n286 185
R1897 VDD.n3742 VDD.n3741 185
R1898 VDD.n3743 VDD.n3742 185
R1899 VDD.n295 VDD.n294 185
R1900 VDD.n294 VDD.n293 185
R1901 VDD.n3737 VDD.n3736 185
R1902 VDD.n3736 VDD.n3735 185
R1903 VDD.n298 VDD.n297 185
R1904 VDD.n299 VDD.n298 185
R1905 VDD.n3726 VDD.n3725 185
R1906 VDD.n3727 VDD.n3726 185
R1907 VDD.n307 VDD.n306 185
R1908 VDD.n306 VDD.n305 185
R1909 VDD.n3721 VDD.n3720 185
R1910 VDD.n3720 VDD.n3719 185
R1911 VDD.n310 VDD.n309 185
R1912 VDD.n311 VDD.n310 185
R1913 VDD.n3710 VDD.n3709 185
R1914 VDD.n3711 VDD.n3710 185
R1915 VDD.n319 VDD.n318 185
R1916 VDD.n318 VDD.n317 185
R1917 VDD.n3705 VDD.n3704 185
R1918 VDD.n3704 VDD.n3703 185
R1919 VDD.n322 VDD.n321 185
R1920 VDD.n323 VDD.n322 185
R1921 VDD.n3694 VDD.n3693 185
R1922 VDD.n3695 VDD.n3694 185
R1923 VDD.n331 VDD.n330 185
R1924 VDD.n330 VDD.n329 185
R1925 VDD.n3689 VDD.n3688 185
R1926 VDD.n3688 VDD.n3687 185
R1927 VDD.n334 VDD.n333 185
R1928 VDD.n335 VDD.n334 185
R1929 VDD.n3678 VDD.n3677 185
R1930 VDD.n3679 VDD.n3678 185
R1931 VDD.n343 VDD.n342 185
R1932 VDD.n342 VDD.n341 185
R1933 VDD.n3673 VDD.n3672 185
R1934 VDD.n3672 VDD.n3671 185
R1935 VDD.n346 VDD.n345 185
R1936 VDD.n347 VDD.n346 185
R1937 VDD.n3662 VDD.n3661 185
R1938 VDD.n3663 VDD.n3662 185
R1939 VDD.n355 VDD.n354 185
R1940 VDD.n354 VDD.n353 185
R1941 VDD.n3657 VDD.n3656 185
R1942 VDD.n3656 VDD.n3655 185
R1943 VDD.n358 VDD.n357 185
R1944 VDD.n359 VDD.n358 185
R1945 VDD.n3646 VDD.n3645 185
R1946 VDD.n3647 VDD.n3646 185
R1947 VDD.n367 VDD.n366 185
R1948 VDD.n366 VDD.n365 185
R1949 VDD.n3641 VDD.n3640 185
R1950 VDD.n3640 VDD.n3639 185
R1951 VDD.n370 VDD.n369 185
R1952 VDD.n371 VDD.n370 185
R1953 VDD.n3630 VDD.n3629 185
R1954 VDD.n3631 VDD.n3630 185
R1955 VDD.n379 VDD.n378 185
R1956 VDD.n378 VDD.n377 185
R1957 VDD.n3625 VDD.n3624 185
R1958 VDD.n3624 VDD.t13 185
R1959 VDD.n382 VDD.n381 185
R1960 VDD.n383 VDD.n382 185
R1961 VDD.n3615 VDD.n3614 185
R1962 VDD.n3616 VDD.n3615 185
R1963 VDD.n391 VDD.n390 185
R1964 VDD.n390 VDD.n389 185
R1965 VDD.n3610 VDD.n3609 185
R1966 VDD.n3609 VDD.n3608 185
R1967 VDD.n3083 VDD.n3082 185
R1968 VDD.n707 VDD.n706 185
R1969 VDD.n3079 VDD.n3078 185
R1970 VDD.n3080 VDD.n3079 185
R1971 VDD.n3077 VDD.n2723 185
R1972 VDD.n3076 VDD.n3075 185
R1973 VDD.n3074 VDD.n3073 185
R1974 VDD.n3072 VDD.n3071 185
R1975 VDD.n3070 VDD.n3069 185
R1976 VDD.n3068 VDD.n3067 185
R1977 VDD.n3066 VDD.n3065 185
R1978 VDD.n3064 VDD.n3063 185
R1979 VDD.n3062 VDD.n3061 185
R1980 VDD.n3060 VDD.n3059 185
R1981 VDD.n3058 VDD.n3057 185
R1982 VDD.n3056 VDD.n3055 185
R1983 VDD.n3054 VDD.n3053 185
R1984 VDD.n3052 VDD.n3051 185
R1985 VDD.n3050 VDD.n3049 185
R1986 VDD.n3048 VDD.n3047 185
R1987 VDD.n3046 VDD.n3045 185
R1988 VDD.n3044 VDD.n3043 185
R1989 VDD.n3042 VDD.n3041 185
R1990 VDD.n3040 VDD.n3039 185
R1991 VDD.n3038 VDD.n2710 185
R1992 VDD.n3080 VDD.n2710 185
R1993 VDD.n3439 VDD.n3438 185
R1994 VDD.n3441 VDD.n408 185
R1995 VDD.n3443 VDD.n3442 185
R1996 VDD.n3445 VDD.n405 185
R1997 VDD.n3447 VDD.n3446 185
R1998 VDD.n3449 VDD.n403 185
R1999 VDD.n3451 VDD.n3450 185
R2000 VDD.n3452 VDD.n402 185
R2001 VDD.n3454 VDD.n3453 185
R2002 VDD.n3456 VDD.n401 185
R2003 VDD.n3457 VDD.n398 185
R2004 VDD.n3460 VDD.n3459 185
R2005 VDD.n399 VDD.n397 185
R2006 VDD.n3412 VDD.n3409 185
R2007 VDD.n3414 VDD.n3413 185
R2008 VDD.n3415 VDD.n3408 185
R2009 VDD.n3417 VDD.n3416 185
R2010 VDD.n3419 VDD.n3406 185
R2011 VDD.n3421 VDD.n3420 185
R2012 VDD.n3422 VDD.n3405 185
R2013 VDD.n3424 VDD.n3423 185
R2014 VDD.n3426 VDD.n3404 185
R2015 VDD.n3427 VDD.n3403 185
R2016 VDD.n3430 VDD.n3429 185
R2017 VDD.n3437 VDD.n410 185
R2018 VDD.n415 VDD.n410 185
R2019 VDD.n3436 VDD.n3435 185
R2020 VDD.n3435 VDD.n3434 185
R2021 VDD.n412 VDD.n411 185
R2022 VDD.n413 VDD.n412 185
R2023 VDD.n2727 VDD.n422 185
R2024 VDD.n3399 VDD.n422 185
R2025 VDD.n2729 VDD.n2728 185
R2026 VDD.n2728 VDD.n421 185
R2027 VDD.n2730 VDD.n451 185
R2028 VDD.n3340 VDD.n451 185
R2029 VDD.n2732 VDD.n2731 185
R2030 VDD.n2731 VDD.n450 185
R2031 VDD.n2733 VDD.n457 185
R2032 VDD.n3334 VDD.n457 185
R2033 VDD.n2735 VDD.n2734 185
R2034 VDD.n2734 VDD.n456 185
R2035 VDD.n2736 VDD.n464 185
R2036 VDD.n3326 VDD.n464 185
R2037 VDD.n2738 VDD.n2737 185
R2038 VDD.n2737 VDD.n463 185
R2039 VDD.n2739 VDD.n470 185
R2040 VDD.n3320 VDD.n470 185
R2041 VDD.n2741 VDD.n2740 185
R2042 VDD.n2740 VDD.n469 185
R2043 VDD.n2742 VDD.n476 185
R2044 VDD.n3314 VDD.n476 185
R2045 VDD.n2744 VDD.n2743 185
R2046 VDD.n2743 VDD.n475 185
R2047 VDD.n2745 VDD.n482 185
R2048 VDD.n3308 VDD.n482 185
R2049 VDD.n2747 VDD.n2746 185
R2050 VDD.n2746 VDD.n481 185
R2051 VDD.n2748 VDD.n488 185
R2052 VDD.n3302 VDD.n488 185
R2053 VDD.n2750 VDD.n2749 185
R2054 VDD.n2749 VDD.n487 185
R2055 VDD.n2751 VDD.n494 185
R2056 VDD.n3296 VDD.n494 185
R2057 VDD.n2753 VDD.n2752 185
R2058 VDD.n2752 VDD.n493 185
R2059 VDD.n2754 VDD.n499 185
R2060 VDD.n3290 VDD.n499 185
R2061 VDD.n2756 VDD.n2755 185
R2062 VDD.n2755 VDD.n507 185
R2063 VDD.n2757 VDD.n505 185
R2064 VDD.n3284 VDD.n505 185
R2065 VDD.n2759 VDD.n2758 185
R2066 VDD.n2758 VDD.n504 185
R2067 VDD.n2760 VDD.n512 185
R2068 VDD.n3278 VDD.n512 185
R2069 VDD.n2762 VDD.n2761 185
R2070 VDD.n2761 VDD.n511 185
R2071 VDD.n2763 VDD.n518 185
R2072 VDD.n3272 VDD.n518 185
R2073 VDD.n2765 VDD.n2764 185
R2074 VDD.n2764 VDD.n517 185
R2075 VDD.n2766 VDD.n524 185
R2076 VDD.n3266 VDD.n524 185
R2077 VDD.n2768 VDD.n2767 185
R2078 VDD.n2767 VDD.n523 185
R2079 VDD.n2769 VDD.n530 185
R2080 VDD.n3260 VDD.n530 185
R2081 VDD.n2771 VDD.n2770 185
R2082 VDD.n2770 VDD.n529 185
R2083 VDD.n2772 VDD.n535 185
R2084 VDD.n3254 VDD.n535 185
R2085 VDD.n2774 VDD.n2773 185
R2086 VDD.n2773 VDD.n543 185
R2087 VDD.n2775 VDD.n541 185
R2088 VDD.n3248 VDD.n541 185
R2089 VDD.n2777 VDD.n2776 185
R2090 VDD.n2776 VDD.n540 185
R2091 VDD.n2778 VDD.n548 185
R2092 VDD.n3242 VDD.n548 185
R2093 VDD.n2780 VDD.n2779 185
R2094 VDD.n2779 VDD.n547 185
R2095 VDD.n2781 VDD.n554 185
R2096 VDD.n3236 VDD.n554 185
R2097 VDD.n2783 VDD.n2782 185
R2098 VDD.n2782 VDD.n553 185
R2099 VDD.n2784 VDD.n560 185
R2100 VDD.n3230 VDD.n560 185
R2101 VDD.n2786 VDD.n2785 185
R2102 VDD.n2785 VDD.n559 185
R2103 VDD.n2787 VDD.n566 185
R2104 VDD.n3224 VDD.n566 185
R2105 VDD.n2789 VDD.n2788 185
R2106 VDD.n2788 VDD.n565 185
R2107 VDD.n2790 VDD.n573 185
R2108 VDD.t108 VDD.n573 185
R2109 VDD.n2792 VDD.n2791 185
R2110 VDD.n2791 VDD.n571 185
R2111 VDD.n2793 VDD.n578 185
R2112 VDD.n3213 VDD.n578 185
R2113 VDD.n2795 VDD.n2794 185
R2114 VDD.n2794 VDD.n577 185
R2115 VDD.n2796 VDD.n583 185
R2116 VDD.n3207 VDD.n583 185
R2117 VDD.n2798 VDD.n2797 185
R2118 VDD.n2797 VDD.n591 185
R2119 VDD.n2799 VDD.n589 185
R2120 VDD.n3201 VDD.n589 185
R2121 VDD.n2801 VDD.n2800 185
R2122 VDD.n2800 VDD.n588 185
R2123 VDD.n2802 VDD.n596 185
R2124 VDD.n3195 VDD.n596 185
R2125 VDD.n2804 VDD.n2803 185
R2126 VDD.n2803 VDD.n595 185
R2127 VDD.n2805 VDD.n602 185
R2128 VDD.n3189 VDD.n602 185
R2129 VDD.n2807 VDD.n2806 185
R2130 VDD.n2806 VDD.n601 185
R2131 VDD.n2808 VDD.n608 185
R2132 VDD.n3183 VDD.n608 185
R2133 VDD.n2810 VDD.n2809 185
R2134 VDD.n2809 VDD.n607 185
R2135 VDD.n2811 VDD.n614 185
R2136 VDD.n3177 VDD.n614 185
R2137 VDD.n2813 VDD.n2812 185
R2138 VDD.n2812 VDD.n613 185
R2139 VDD.n2814 VDD.n619 185
R2140 VDD.n3171 VDD.n619 185
R2141 VDD.n2816 VDD.n2815 185
R2142 VDD.n2815 VDD.n627 185
R2143 VDD.n2817 VDD.n625 185
R2144 VDD.n3165 VDD.n625 185
R2145 VDD.n2819 VDD.n2818 185
R2146 VDD.n2818 VDD.n624 185
R2147 VDD.n2820 VDD.n632 185
R2148 VDD.n3159 VDD.n632 185
R2149 VDD.n2822 VDD.n2821 185
R2150 VDD.n2821 VDD.n631 185
R2151 VDD.n2823 VDD.n638 185
R2152 VDD.n3153 VDD.n638 185
R2153 VDD.n2825 VDD.n2824 185
R2154 VDD.n2824 VDD.n637 185
R2155 VDD.n2826 VDD.n644 185
R2156 VDD.n3147 VDD.n644 185
R2157 VDD.n2828 VDD.n2827 185
R2158 VDD.n2827 VDD.n643 185
R2159 VDD.n2829 VDD.n650 185
R2160 VDD.n3141 VDD.n650 185
R2161 VDD.n2831 VDD.n2830 185
R2162 VDD.n2830 VDD.n649 185
R2163 VDD.n2832 VDD.n655 185
R2164 VDD.n3135 VDD.n655 185
R2165 VDD.n2834 VDD.n2833 185
R2166 VDD.n2833 VDD.n663 185
R2167 VDD.n2835 VDD.n661 185
R2168 VDD.n3129 VDD.n661 185
R2169 VDD.n2837 VDD.n2836 185
R2170 VDD.n2836 VDD.n660 185
R2171 VDD.n2838 VDD.n668 185
R2172 VDD.n3123 VDD.n668 185
R2173 VDD.n2840 VDD.n2839 185
R2174 VDD.n2839 VDD.n667 185
R2175 VDD.n2841 VDD.n674 185
R2176 VDD.n3117 VDD.n674 185
R2177 VDD.n2843 VDD.n2842 185
R2178 VDD.n2842 VDD.n673 185
R2179 VDD.n2844 VDD.n680 185
R2180 VDD.n3111 VDD.n680 185
R2181 VDD.n2846 VDD.n2845 185
R2182 VDD.n2845 VDD.n679 185
R2183 VDD.n2847 VDD.n685 185
R2184 VDD.n3105 VDD.n685 185
R2185 VDD.n3028 VDD.n3027 185
R2186 VDD.n3027 VDD.n3026 185
R2187 VDD.n3029 VDD.n691 185
R2188 VDD.n3099 VDD.n691 185
R2189 VDD.n3031 VDD.n3030 185
R2190 VDD.n3030 VDD.n690 185
R2191 VDD.n3032 VDD.n697 185
R2192 VDD.n3093 VDD.n697 185
R2193 VDD.n3034 VDD.n3033 185
R2194 VDD.n3033 VDD.n696 185
R2195 VDD.n3035 VDD.n703 185
R2196 VDD.n3087 VDD.n703 185
R2197 VDD.n3037 VDD.n3036 185
R2198 VDD.n3036 VDD.n702 185
R2199 VDD.n3084 VDD.n705 185
R2200 VDD.n705 VDD.n702 185
R2201 VDD.n3086 VDD.n3085 185
R2202 VDD.n3087 VDD.n3086 185
R2203 VDD.n695 VDD.n694 185
R2204 VDD.n696 VDD.n695 185
R2205 VDD.n3095 VDD.n3094 185
R2206 VDD.n3094 VDD.n3093 185
R2207 VDD.n3096 VDD.n693 185
R2208 VDD.n693 VDD.n690 185
R2209 VDD.n3098 VDD.n3097 185
R2210 VDD.n3099 VDD.n3098 185
R2211 VDD.n684 VDD.n683 185
R2212 VDD.n3026 VDD.n684 185
R2213 VDD.n3107 VDD.n3106 185
R2214 VDD.n3106 VDD.n3105 185
R2215 VDD.n3108 VDD.n682 185
R2216 VDD.n682 VDD.n679 185
R2217 VDD.n3110 VDD.n3109 185
R2218 VDD.n3111 VDD.n3110 185
R2219 VDD.n672 VDD.n671 185
R2220 VDD.n673 VDD.n672 185
R2221 VDD.n3119 VDD.n3118 185
R2222 VDD.n3118 VDD.n3117 185
R2223 VDD.n3120 VDD.n670 185
R2224 VDD.n670 VDD.n667 185
R2225 VDD.n3122 VDD.n3121 185
R2226 VDD.n3123 VDD.n3122 185
R2227 VDD.n659 VDD.n658 185
R2228 VDD.n660 VDD.n659 185
R2229 VDD.n3131 VDD.n3130 185
R2230 VDD.n3130 VDD.n3129 185
R2231 VDD.n3132 VDD.n657 185
R2232 VDD.n663 VDD.n657 185
R2233 VDD.n3134 VDD.n3133 185
R2234 VDD.n3135 VDD.n3134 185
R2235 VDD.n648 VDD.n647 185
R2236 VDD.n649 VDD.n648 185
R2237 VDD.n3143 VDD.n3142 185
R2238 VDD.n3142 VDD.n3141 185
R2239 VDD.n3144 VDD.n646 185
R2240 VDD.n646 VDD.n643 185
R2241 VDD.n3146 VDD.n3145 185
R2242 VDD.n3147 VDD.n3146 185
R2243 VDD.n636 VDD.n635 185
R2244 VDD.n637 VDD.n636 185
R2245 VDD.n3155 VDD.n3154 185
R2246 VDD.n3154 VDD.n3153 185
R2247 VDD.n3156 VDD.n634 185
R2248 VDD.n634 VDD.n631 185
R2249 VDD.n3158 VDD.n3157 185
R2250 VDD.n3159 VDD.n3158 185
R2251 VDD.n623 VDD.n622 185
R2252 VDD.n624 VDD.n623 185
R2253 VDD.n3167 VDD.n3166 185
R2254 VDD.n3166 VDD.n3165 185
R2255 VDD.n3168 VDD.n621 185
R2256 VDD.n627 VDD.n621 185
R2257 VDD.n3170 VDD.n3169 185
R2258 VDD.n3171 VDD.n3170 185
R2259 VDD.n612 VDD.n611 185
R2260 VDD.n613 VDD.n612 185
R2261 VDD.n3179 VDD.n3178 185
R2262 VDD.n3178 VDD.n3177 185
R2263 VDD.n3180 VDD.n610 185
R2264 VDD.n610 VDD.n607 185
R2265 VDD.n3182 VDD.n3181 185
R2266 VDD.n3183 VDD.n3182 185
R2267 VDD.n600 VDD.n599 185
R2268 VDD.n601 VDD.n600 185
R2269 VDD.n3191 VDD.n3190 185
R2270 VDD.n3190 VDD.n3189 185
R2271 VDD.n3192 VDD.n598 185
R2272 VDD.n598 VDD.n595 185
R2273 VDD.n3194 VDD.n3193 185
R2274 VDD.n3195 VDD.n3194 185
R2275 VDD.n587 VDD.n586 185
R2276 VDD.n588 VDD.n587 185
R2277 VDD.n3203 VDD.n3202 185
R2278 VDD.n3202 VDD.n3201 185
R2279 VDD.n3204 VDD.n585 185
R2280 VDD.n591 VDD.n585 185
R2281 VDD.n3206 VDD.n3205 185
R2282 VDD.n3207 VDD.n3206 185
R2283 VDD.n576 VDD.n575 185
R2284 VDD.n577 VDD.n576 185
R2285 VDD.n3215 VDD.n3214 185
R2286 VDD.n3214 VDD.n3213 185
R2287 VDD.n3216 VDD.n574 185
R2288 VDD.n574 VDD.n571 185
R2289 VDD.n3218 VDD.n3217 185
R2290 VDD.t108 VDD.n3218 185
R2291 VDD.n564 VDD.n563 185
R2292 VDD.n565 VDD.n564 185
R2293 VDD.n3226 VDD.n3225 185
R2294 VDD.n3225 VDD.n3224 185
R2295 VDD.n3227 VDD.n562 185
R2296 VDD.n562 VDD.n559 185
R2297 VDD.n3229 VDD.n3228 185
R2298 VDD.n3230 VDD.n3229 185
R2299 VDD.n552 VDD.n551 185
R2300 VDD.n553 VDD.n552 185
R2301 VDD.n3238 VDD.n3237 185
R2302 VDD.n3237 VDD.n3236 185
R2303 VDD.n3239 VDD.n550 185
R2304 VDD.n550 VDD.n547 185
R2305 VDD.n3241 VDD.n3240 185
R2306 VDD.n3242 VDD.n3241 185
R2307 VDD.n539 VDD.n538 185
R2308 VDD.n540 VDD.n539 185
R2309 VDD.n3250 VDD.n3249 185
R2310 VDD.n3249 VDD.n3248 185
R2311 VDD.n3251 VDD.n537 185
R2312 VDD.n543 VDD.n537 185
R2313 VDD.n3253 VDD.n3252 185
R2314 VDD.n3254 VDD.n3253 185
R2315 VDD.n528 VDD.n527 185
R2316 VDD.n529 VDD.n528 185
R2317 VDD.n3262 VDD.n3261 185
R2318 VDD.n3261 VDD.n3260 185
R2319 VDD.n3263 VDD.n526 185
R2320 VDD.n526 VDD.n523 185
R2321 VDD.n3265 VDD.n3264 185
R2322 VDD.n3266 VDD.n3265 185
R2323 VDD.n516 VDD.n515 185
R2324 VDD.n517 VDD.n516 185
R2325 VDD.n3274 VDD.n3273 185
R2326 VDD.n3273 VDD.n3272 185
R2327 VDD.n3275 VDD.n514 185
R2328 VDD.n514 VDD.n511 185
R2329 VDD.n3277 VDD.n3276 185
R2330 VDD.n3278 VDD.n3277 185
R2331 VDD.n503 VDD.n502 185
R2332 VDD.n504 VDD.n503 185
R2333 VDD.n3286 VDD.n3285 185
R2334 VDD.n3285 VDD.n3284 185
R2335 VDD.n3287 VDD.n501 185
R2336 VDD.n507 VDD.n501 185
R2337 VDD.n3289 VDD.n3288 185
R2338 VDD.n3290 VDD.n3289 185
R2339 VDD.n492 VDD.n491 185
R2340 VDD.n493 VDD.n492 185
R2341 VDD.n3298 VDD.n3297 185
R2342 VDD.n3297 VDD.n3296 185
R2343 VDD.n3299 VDD.n490 185
R2344 VDD.n490 VDD.n487 185
R2345 VDD.n3301 VDD.n3300 185
R2346 VDD.n3302 VDD.n3301 185
R2347 VDD.n480 VDD.n479 185
R2348 VDD.n481 VDD.n480 185
R2349 VDD.n3310 VDD.n3309 185
R2350 VDD.n3309 VDD.n3308 185
R2351 VDD.n3311 VDD.n478 185
R2352 VDD.n478 VDD.n475 185
R2353 VDD.n3313 VDD.n3312 185
R2354 VDD.n3314 VDD.n3313 185
R2355 VDD.n468 VDD.n467 185
R2356 VDD.n469 VDD.n468 185
R2357 VDD.n3322 VDD.n3321 185
R2358 VDD.n3321 VDD.n3320 185
R2359 VDD.n3323 VDD.n466 185
R2360 VDD.n466 VDD.n463 185
R2361 VDD.n3325 VDD.n3324 185
R2362 VDD.n3326 VDD.n3325 185
R2363 VDD.n455 VDD.n454 185
R2364 VDD.n456 VDD.n455 185
R2365 VDD.n3336 VDD.n3335 185
R2366 VDD.n3335 VDD.n3334 185
R2367 VDD.n3337 VDD.n453 185
R2368 VDD.n453 VDD.n450 185
R2369 VDD.n3339 VDD.n3338 185
R2370 VDD.n3340 VDD.n3339 185
R2371 VDD.n420 VDD.n419 185
R2372 VDD.n421 VDD.n420 185
R2373 VDD.n3401 VDD.n3400 185
R2374 VDD.n3400 VDD.n3399 185
R2375 VDD.n3402 VDD.n417 185
R2376 VDD.n417 VDD.n413 185
R2377 VDD.n3433 VDD.n3432 185
R2378 VDD.n3434 VDD.n3433 185
R2379 VDD.n3431 VDD.n418 185
R2380 VDD.n418 VDD.n415 185
R2381 VDD.n735 VDD.n733 185
R2382 VDD.n733 VDD.n708 185
R2383 VDD.n2577 VDD.n743 185
R2384 VDD.n2649 VDD.n743 185
R2385 VDD.n2579 VDD.n2578 185
R2386 VDD.n2578 VDD.n741 185
R2387 VDD.n2580 VDD.n753 185
R2388 VDD.n2590 VDD.n753 185
R2389 VDD.n2581 VDD.n760 185
R2390 VDD.n760 VDD.n751 185
R2391 VDD.n2583 VDD.n2582 185
R2392 VDD.n2584 VDD.n2583 185
R2393 VDD.n2576 VDD.n759 185
R2394 VDD.n2399 VDD.n759 185
R2395 VDD.n2575 VDD.n2574 185
R2396 VDD.n2574 VDD.n2573 185
R2397 VDD.n762 VDD.n761 185
R2398 VDD.n763 VDD.n762 185
R2399 VDD.n2566 VDD.n2565 185
R2400 VDD.n2567 VDD.n2566 185
R2401 VDD.n2564 VDD.n772 185
R2402 VDD.n772 VDD.n769 185
R2403 VDD.n2563 VDD.n2562 185
R2404 VDD.n2562 VDD.n2561 185
R2405 VDD.n774 VDD.n773 185
R2406 VDD.n775 VDD.n774 185
R2407 VDD.n2554 VDD.n2553 185
R2408 VDD.n2555 VDD.n2554 185
R2409 VDD.n2552 VDD.n784 185
R2410 VDD.n784 VDD.n781 185
R2411 VDD.n2551 VDD.n2550 185
R2412 VDD.n2550 VDD.n2549 185
R2413 VDD.n786 VDD.n785 185
R2414 VDD.n787 VDD.n786 185
R2415 VDD.n2542 VDD.n2541 185
R2416 VDD.n2543 VDD.n2542 185
R2417 VDD.n2540 VDD.n796 185
R2418 VDD.n796 VDD.n793 185
R2419 VDD.n2539 VDD.n2538 185
R2420 VDD.n2538 VDD.n2537 185
R2421 VDD.n798 VDD.n797 185
R2422 VDD.n799 VDD.n798 185
R2423 VDD.n2530 VDD.n2529 185
R2424 VDD.n2531 VDD.n2530 185
R2425 VDD.n2528 VDD.n807 185
R2426 VDD.n813 VDD.n807 185
R2427 VDD.n2527 VDD.n2526 185
R2428 VDD.n2526 VDD.n2525 185
R2429 VDD.n809 VDD.n808 185
R2430 VDD.n810 VDD.n809 185
R2431 VDD.n2518 VDD.n2517 185
R2432 VDD.n2519 VDD.n2518 185
R2433 VDD.n2516 VDD.n820 185
R2434 VDD.n820 VDD.n817 185
R2435 VDD.n2515 VDD.n2514 185
R2436 VDD.n2514 VDD.n2513 185
R2437 VDD.n822 VDD.n821 185
R2438 VDD.n823 VDD.n822 185
R2439 VDD.n2506 VDD.n2505 185
R2440 VDD.n2507 VDD.n2506 185
R2441 VDD.n2504 VDD.n832 185
R2442 VDD.n832 VDD.n829 185
R2443 VDD.n2503 VDD.n2502 185
R2444 VDD.n2502 VDD.n2501 185
R2445 VDD.n834 VDD.n833 185
R2446 VDD.n835 VDD.n834 185
R2447 VDD.n2494 VDD.n2493 185
R2448 VDD.n2495 VDD.n2494 185
R2449 VDD.n2492 VDD.n843 185
R2450 VDD.n849 VDD.n843 185
R2451 VDD.n2491 VDD.n2490 185
R2452 VDD.n2490 VDD.n2489 185
R2453 VDD.n845 VDD.n844 185
R2454 VDD.n846 VDD.n845 185
R2455 VDD.n2482 VDD.n2481 185
R2456 VDD.n2483 VDD.n2482 185
R2457 VDD.n2480 VDD.n856 185
R2458 VDD.n856 VDD.n853 185
R2459 VDD.n2479 VDD.n2478 185
R2460 VDD.n2478 VDD.n2477 185
R2461 VDD.n858 VDD.n857 185
R2462 VDD.n859 VDD.n858 185
R2463 VDD.n2470 VDD.n2469 185
R2464 VDD.n2471 VDD.n2470 185
R2465 VDD.n2468 VDD.n868 185
R2466 VDD.n868 VDD.n865 185
R2467 VDD.n2467 VDD.n2466 185
R2468 VDD.n2466 VDD.n2465 185
R2469 VDD.n870 VDD.n869 185
R2470 VDD.n871 VDD.n870 185
R2471 VDD.n2317 VDD.n878 185
R2472 VDD.t100 VDD.n878 185
R2473 VDD.n2319 VDD.n2318 185
R2474 VDD.n2318 VDD.n877 185
R2475 VDD.n2320 VDD.n889 185
R2476 VDD.n2330 VDD.n889 185
R2477 VDD.n2321 VDD.n897 185
R2478 VDD.n897 VDD.n887 185
R2479 VDD.n2323 VDD.n2322 185
R2480 VDD.n2324 VDD.n2323 185
R2481 VDD.n2316 VDD.n896 185
R2482 VDD.n896 VDD.n893 185
R2483 VDD.n2315 VDD.n2314 185
R2484 VDD.n2314 VDD.n2313 185
R2485 VDD.n899 VDD.n898 185
R2486 VDD.n900 VDD.n899 185
R2487 VDD.n2306 VDD.n2305 185
R2488 VDD.n2307 VDD.n2306 185
R2489 VDD.n2304 VDD.n909 185
R2490 VDD.n909 VDD.n906 185
R2491 VDD.n2303 VDD.n2302 185
R2492 VDD.n2302 VDD.n2301 185
R2493 VDD.n911 VDD.n910 185
R2494 VDD.n912 VDD.n911 185
R2495 VDD.n2294 VDD.n2293 185
R2496 VDD.n2295 VDD.n2294 185
R2497 VDD.n2292 VDD.n920 185
R2498 VDD.n926 VDD.n920 185
R2499 VDD.n2291 VDD.n2290 185
R2500 VDD.n2290 VDD.n2289 185
R2501 VDD.n922 VDD.n921 185
R2502 VDD.n923 VDD.n922 185
R2503 VDD.n2282 VDD.n2281 185
R2504 VDD.n2283 VDD.n2282 185
R2505 VDD.n2280 VDD.n933 185
R2506 VDD.n933 VDD.n930 185
R2507 VDD.n2279 VDD.n2278 185
R2508 VDD.n2278 VDD.n2277 185
R2509 VDD.n935 VDD.n934 185
R2510 VDD.n936 VDD.n935 185
R2511 VDD.n2270 VDD.n2269 185
R2512 VDD.n2271 VDD.n2270 185
R2513 VDD.n2268 VDD.n945 185
R2514 VDD.n945 VDD.n942 185
R2515 VDD.n2267 VDD.n2266 185
R2516 VDD.n2266 VDD.n2265 185
R2517 VDD.n947 VDD.n946 185
R2518 VDD.n948 VDD.n947 185
R2519 VDD.n2258 VDD.n2257 185
R2520 VDD.n2259 VDD.n2258 185
R2521 VDD.n2256 VDD.n956 185
R2522 VDD.n962 VDD.n956 185
R2523 VDD.n2255 VDD.n2254 185
R2524 VDD.n2254 VDD.n2253 185
R2525 VDD.n958 VDD.n957 185
R2526 VDD.n959 VDD.n958 185
R2527 VDD.n2246 VDD.n2245 185
R2528 VDD.n2247 VDD.n2246 185
R2529 VDD.n2244 VDD.n969 185
R2530 VDD.n969 VDD.n966 185
R2531 VDD.n2243 VDD.n2242 185
R2532 VDD.n2242 VDD.n2241 185
R2533 VDD.n971 VDD.n970 185
R2534 VDD.n972 VDD.n971 185
R2535 VDD.n2234 VDD.n2233 185
R2536 VDD.n2235 VDD.n2234 185
R2537 VDD.n2232 VDD.n981 185
R2538 VDD.n981 VDD.n978 185
R2539 VDD.n2231 VDD.n2230 185
R2540 VDD.n2230 VDD.n2229 185
R2541 VDD.n983 VDD.n982 185
R2542 VDD.n984 VDD.n983 185
R2543 VDD.n2222 VDD.n2221 185
R2544 VDD.n2223 VDD.n2222 185
R2545 VDD.n2220 VDD.n992 185
R2546 VDD.n997 VDD.n992 185
R2547 VDD.n2219 VDD.n2218 185
R2548 VDD.n2218 VDD.n2217 185
R2549 VDD.n994 VDD.n993 185
R2550 VDD.n1004 VDD.n994 185
R2551 VDD.n2210 VDD.n2209 185
R2552 VDD.n2211 VDD.n2210 185
R2553 VDD.n2208 VDD.n1005 185
R2554 VDD.n1005 VDD.n1001 185
R2555 VDD.n2207 VDD.n2206 185
R2556 VDD.n2206 VDD.n2205 185
R2557 VDD.n1007 VDD.n1006 185
R2558 VDD.n1008 VDD.n1007 185
R2559 VDD.n2198 VDD.n2197 185
R2560 VDD.n2199 VDD.n2198 185
R2561 VDD.n2196 VDD.n1017 185
R2562 VDD.n1017 VDD.n1014 185
R2563 VDD.n2653 VDD.n732 185
R2564 VDD.n2699 VDD.n732 185
R2565 VDD.n2655 VDD.n2654 185
R2566 VDD.n2657 VDD.n2656 185
R2567 VDD.n2659 VDD.n2658 185
R2568 VDD.n2661 VDD.n2660 185
R2569 VDD.n2663 VDD.n2662 185
R2570 VDD.n2665 VDD.n2664 185
R2571 VDD.n2667 VDD.n2666 185
R2572 VDD.n2669 VDD.n2668 185
R2573 VDD.n2671 VDD.n2670 185
R2574 VDD.n2673 VDD.n2672 185
R2575 VDD.n2675 VDD.n2674 185
R2576 VDD.n2677 VDD.n2676 185
R2577 VDD.n2679 VDD.n2678 185
R2578 VDD.n2681 VDD.n2680 185
R2579 VDD.n2683 VDD.n2682 185
R2580 VDD.n2685 VDD.n2684 185
R2581 VDD.n2687 VDD.n2686 185
R2582 VDD.n2689 VDD.n2688 185
R2583 VDD.n2691 VDD.n2690 185
R2584 VDD.n2693 VDD.n2692 185
R2585 VDD.n2695 VDD.n2694 185
R2586 VDD.n2696 VDD.n734 185
R2587 VDD.n2698 VDD.n2697 185
R2588 VDD.n2699 VDD.n2698 185
R2589 VDD.n2652 VDD.n2651 185
R2590 VDD.n2651 VDD.n708 185
R2591 VDD.n2650 VDD.n739 185
R2592 VDD.n2650 VDD.n2649 185
R2593 VDD.n2392 VDD.n740 185
R2594 VDD.n741 VDD.n740 185
R2595 VDD.n2393 VDD.n752 185
R2596 VDD.n2590 VDD.n752 185
R2597 VDD.n2395 VDD.n2394 185
R2598 VDD.n2394 VDD.n751 185
R2599 VDD.n2396 VDD.n758 185
R2600 VDD.n2584 VDD.n758 185
R2601 VDD.n2398 VDD.n2397 185
R2602 VDD.n2399 VDD.n2398 185
R2603 VDD.n2391 VDD.n765 185
R2604 VDD.n2573 VDD.n765 185
R2605 VDD.n2390 VDD.n2389 185
R2606 VDD.n2389 VDD.n763 185
R2607 VDD.n2388 VDD.n771 185
R2608 VDD.n2567 VDD.n771 185
R2609 VDD.n2387 VDD.n2386 185
R2610 VDD.n2386 VDD.n769 185
R2611 VDD.n2385 VDD.n777 185
R2612 VDD.n2561 VDD.n777 185
R2613 VDD.n2384 VDD.n2383 185
R2614 VDD.n2383 VDD.n775 185
R2615 VDD.n2382 VDD.n783 185
R2616 VDD.n2555 VDD.n783 185
R2617 VDD.n2381 VDD.n2380 185
R2618 VDD.n2380 VDD.n781 185
R2619 VDD.n2379 VDD.n789 185
R2620 VDD.n2549 VDD.n789 185
R2621 VDD.n2378 VDD.n2377 185
R2622 VDD.n2377 VDD.n787 185
R2623 VDD.n2376 VDD.n795 185
R2624 VDD.n2543 VDD.n795 185
R2625 VDD.n2375 VDD.n2374 185
R2626 VDD.n2374 VDD.n793 185
R2627 VDD.n2373 VDD.n801 185
R2628 VDD.n2537 VDD.n801 185
R2629 VDD.n2372 VDD.n2371 185
R2630 VDD.n2371 VDD.n799 185
R2631 VDD.n2370 VDD.n806 185
R2632 VDD.n2531 VDD.n806 185
R2633 VDD.n2369 VDD.n2368 185
R2634 VDD.n2368 VDD.n813 185
R2635 VDD.n2367 VDD.n812 185
R2636 VDD.n2525 VDD.n812 185
R2637 VDD.n2366 VDD.n2365 185
R2638 VDD.n2365 VDD.n810 185
R2639 VDD.n2364 VDD.n819 185
R2640 VDD.n2519 VDD.n819 185
R2641 VDD.n2363 VDD.n2362 185
R2642 VDD.n2362 VDD.n817 185
R2643 VDD.n2361 VDD.n825 185
R2644 VDD.n2513 VDD.n825 185
R2645 VDD.n2360 VDD.n2359 185
R2646 VDD.n2359 VDD.n823 185
R2647 VDD.n2358 VDD.n831 185
R2648 VDD.n2507 VDD.n831 185
R2649 VDD.n2357 VDD.n2356 185
R2650 VDD.n2356 VDD.n829 185
R2651 VDD.n2355 VDD.n837 185
R2652 VDD.n2501 VDD.n837 185
R2653 VDD.n2354 VDD.n2353 185
R2654 VDD.n2353 VDD.n835 185
R2655 VDD.n2352 VDD.n842 185
R2656 VDD.n2495 VDD.n842 185
R2657 VDD.n2351 VDD.n2350 185
R2658 VDD.n2350 VDD.n849 185
R2659 VDD.n2349 VDD.n848 185
R2660 VDD.n2489 VDD.n848 185
R2661 VDD.n2348 VDD.n2347 185
R2662 VDD.n2347 VDD.n846 185
R2663 VDD.n2346 VDD.n855 185
R2664 VDD.n2483 VDD.n855 185
R2665 VDD.n2345 VDD.n2344 185
R2666 VDD.n2344 VDD.n853 185
R2667 VDD.n2343 VDD.n861 185
R2668 VDD.n2477 VDD.n861 185
R2669 VDD.n2342 VDD.n2341 185
R2670 VDD.n2341 VDD.n859 185
R2671 VDD.n2340 VDD.n867 185
R2672 VDD.n2471 VDD.n867 185
R2673 VDD.n2339 VDD.n2338 185
R2674 VDD.n2338 VDD.n865 185
R2675 VDD.n2337 VDD.n873 185
R2676 VDD.n2465 VDD.n873 185
R2677 VDD.n2336 VDD.n2335 185
R2678 VDD.n2335 VDD.n871 185
R2679 VDD.n2334 VDD.n879 185
R2680 VDD.t100 VDD.n879 185
R2681 VDD.n2333 VDD.n2332 185
R2682 VDD.n2332 VDD.n877 185
R2683 VDD.n2331 VDD.n885 185
R2684 VDD.n2331 VDD.n2330 185
R2685 VDD.n1992 VDD.n886 185
R2686 VDD.n887 VDD.n886 185
R2687 VDD.n1993 VDD.n895 185
R2688 VDD.n2324 VDD.n895 185
R2689 VDD.n1995 VDD.n1994 185
R2690 VDD.n1994 VDD.n893 185
R2691 VDD.n1996 VDD.n902 185
R2692 VDD.n2313 VDD.n902 185
R2693 VDD.n1998 VDD.n1997 185
R2694 VDD.n1997 VDD.n900 185
R2695 VDD.n1999 VDD.n908 185
R2696 VDD.n2307 VDD.n908 185
R2697 VDD.n2001 VDD.n2000 185
R2698 VDD.n2000 VDD.n906 185
R2699 VDD.n2002 VDD.n914 185
R2700 VDD.n2301 VDD.n914 185
R2701 VDD.n2004 VDD.n2003 185
R2702 VDD.n2003 VDD.n912 185
R2703 VDD.n2005 VDD.n919 185
R2704 VDD.n2295 VDD.n919 185
R2705 VDD.n2007 VDD.n2006 185
R2706 VDD.n2006 VDD.n926 185
R2707 VDD.n2008 VDD.n925 185
R2708 VDD.n2289 VDD.n925 185
R2709 VDD.n2010 VDD.n2009 185
R2710 VDD.n2009 VDD.n923 185
R2711 VDD.n2011 VDD.n932 185
R2712 VDD.n2283 VDD.n932 185
R2713 VDD.n2013 VDD.n2012 185
R2714 VDD.n2012 VDD.n930 185
R2715 VDD.n2014 VDD.n938 185
R2716 VDD.n2277 VDD.n938 185
R2717 VDD.n2016 VDD.n2015 185
R2718 VDD.n2015 VDD.n936 185
R2719 VDD.n2017 VDD.n944 185
R2720 VDD.n2271 VDD.n944 185
R2721 VDD.n2019 VDD.n2018 185
R2722 VDD.n2018 VDD.n942 185
R2723 VDD.n2020 VDD.n950 185
R2724 VDD.n2265 VDD.n950 185
R2725 VDD.n2022 VDD.n2021 185
R2726 VDD.n2021 VDD.n948 185
R2727 VDD.n2023 VDD.n955 185
R2728 VDD.n2259 VDD.n955 185
R2729 VDD.n2025 VDD.n2024 185
R2730 VDD.n2024 VDD.n962 185
R2731 VDD.n2026 VDD.n961 185
R2732 VDD.n2253 VDD.n961 185
R2733 VDD.n2028 VDD.n2027 185
R2734 VDD.n2027 VDD.n959 185
R2735 VDD.n2029 VDD.n968 185
R2736 VDD.n2247 VDD.n968 185
R2737 VDD.n2031 VDD.n2030 185
R2738 VDD.n2030 VDD.n966 185
R2739 VDD.n2032 VDD.n974 185
R2740 VDD.n2241 VDD.n974 185
R2741 VDD.n2034 VDD.n2033 185
R2742 VDD.n2033 VDD.n972 185
R2743 VDD.n2035 VDD.n980 185
R2744 VDD.n2235 VDD.n980 185
R2745 VDD.n2037 VDD.n2036 185
R2746 VDD.n2036 VDD.n978 185
R2747 VDD.n2038 VDD.n986 185
R2748 VDD.n2229 VDD.n986 185
R2749 VDD.n2040 VDD.n2039 185
R2750 VDD.n2039 VDD.n984 185
R2751 VDD.n2041 VDD.n991 185
R2752 VDD.n2223 VDD.n991 185
R2753 VDD.n2043 VDD.n2042 185
R2754 VDD.n2042 VDD.n997 185
R2755 VDD.n2044 VDD.n996 185
R2756 VDD.n2217 VDD.n996 185
R2757 VDD.n2046 VDD.n2045 185
R2758 VDD.n2045 VDD.n1004 185
R2759 VDD.n2047 VDD.n1003 185
R2760 VDD.n2211 VDD.n1003 185
R2761 VDD.n2049 VDD.n2048 185
R2762 VDD.n2048 VDD.n1001 185
R2763 VDD.n2050 VDD.n1010 185
R2764 VDD.n2205 VDD.n1010 185
R2765 VDD.n2052 VDD.n2051 185
R2766 VDD.n2051 VDD.n1008 185
R2767 VDD.n2053 VDD.n1016 185
R2768 VDD.n2199 VDD.n1016 185
R2769 VDD.n2055 VDD.n2054 185
R2770 VDD.n2054 VDD.n1014 185
R2771 VDD.n2195 VDD.n2194 185
R2772 VDD.n2194 VDD.n2193 185
R2773 VDD.n1019 VDD.n1018 185
R2774 VDD.n1970 VDD.n1969 185
R2775 VDD.n1972 VDD.n1971 185
R2776 VDD.n1974 VDD.n1973 185
R2777 VDD.n1976 VDD.n1975 185
R2778 VDD.n1978 VDD.n1977 185
R2779 VDD.n1980 VDD.n1979 185
R2780 VDD.n1982 VDD.n1981 185
R2781 VDD.n1984 VDD.n1983 185
R2782 VDD.n1986 VDD.n1985 185
R2783 VDD.n1988 VDD.n1987 185
R2784 VDD.n2078 VDD.n2077 185
R2785 VDD.n2076 VDD.n2075 185
R2786 VDD.n2074 VDD.n2073 185
R2787 VDD.n2072 VDD.n2071 185
R2788 VDD.n2070 VDD.n2069 185
R2789 VDD.n2068 VDD.n2067 185
R2790 VDD.n2066 VDD.n2065 185
R2791 VDD.n2064 VDD.n2063 185
R2792 VDD.n2062 VDD.n2061 185
R2793 VDD.n2060 VDD.n2059 185
R2794 VDD.n2058 VDD.n2057 185
R2795 VDD.n2056 VDD.n1042 185
R2796 VDD.n2193 VDD.n1042 185
R2797 VDD.n40 VDD.t194 179
R2798 VDD.n32 VDD.t174 179
R2799 VDD.n24 VDD.t145 179
R2800 VDD.n17 VDD.t171 179
R2801 VDD.n1790 VDD.t165 179
R2802 VDD.n1782 VDD.t119 179
R2803 VDD.n1774 VDD.t132 179
R2804 VDD.n1767 VDD.t166 179
R2805 VDD.n45 VDD.t182 177.286
R2806 VDD.n37 VDD.t159 177.286
R2807 VDD.n29 VDD.t169 177.286
R2808 VDD.n22 VDD.t187 177.286
R2809 VDD.n1795 VDD.t148 177.286
R2810 VDD.n1787 VDD.t189 177.286
R2811 VDD.n1779 VDD.t164 177.286
R2812 VDD.n1772 VDD.t178 177.286
R2813 VDD.n1448 VDD.t18 172.47
R2814 VDD.n1539 VDD.t61 172.47
R2815 VDD.n1493 VDD.t38 172.47
R2816 VDD.n1574 VDD.t51 172.47
R2817 VDD.n2083 VDD.t71 172.47
R2818 VDD.n2106 VDD.t49 172.47
R2819 VDD.n2129 VDD.t74 172.47
R2820 VDD.n1169 VDD.t30 172.47
R2821 VDD.n3842 VDD.t33 172.47
R2822 VDD.n220 VDD.t80 172.47
R2823 VDD.n3880 VDD.t68 172.47
R2824 VDD.n180 VDD.t26 172.47
R2825 VDD.n3473 VDD.t45 172.47
R2826 VDD.n3490 VDD.t14 172.47
R2827 VDD.n3508 VDD.t64 172.47
R2828 VDD.n3524 VDD.t21 172.47
R2829 VDD.n44 VDD.n43 162.306
R2830 VDD.n42 VDD.n41 162.306
R2831 VDD.n40 VDD.n39 162.306
R2832 VDD.n36 VDD.n35 162.306
R2833 VDD.n34 VDD.n33 162.306
R2834 VDD.n32 VDD.n31 162.306
R2835 VDD.n28 VDD.n27 162.306
R2836 VDD.n26 VDD.n25 162.306
R2837 VDD.n24 VDD.n23 162.306
R2838 VDD.n21 VDD.n20 162.306
R2839 VDD.n19 VDD.n18 162.306
R2840 VDD.n17 VDD.n16 162.306
R2841 VDD.n1790 VDD.n1789 162.306
R2842 VDD.n1792 VDD.n1791 162.306
R2843 VDD.n1794 VDD.n1793 162.306
R2844 VDD.n1782 VDD.n1781 162.306
R2845 VDD.n1784 VDD.n1783 162.306
R2846 VDD.n1786 VDD.n1785 162.306
R2847 VDD.n1774 VDD.n1773 162.306
R2848 VDD.n1776 VDD.n1775 162.306
R2849 VDD.n1778 VDD.n1777 162.306
R2850 VDD.n1767 VDD.n1766 162.306
R2851 VDD.n1769 VDD.n1768 162.306
R2852 VDD.n1771 VDD.n1770 162.306
R2853 VDD.t117 VDD.t91 153.089
R2854 VDD.t114 VDD.t101 153.089
R2855 VDD.n170 VDD.n167 146.341
R2856 VDD.n3908 VDD.n3907 146.341
R2857 VDD.n3905 VDD.n174 146.341
R2858 VDD.n3901 VDD.n3900 146.341
R2859 VDD.n3898 VDD.n183 146.341
R2860 VDD.n3894 VDD.n3893 146.341
R2861 VDD.n3891 VDD.n190 146.341
R2862 VDD.n3887 VDD.n3886 146.341
R2863 VDD.n3884 VDD.n197 146.341
R2864 VDD.n3877 VDD.n3876 146.341
R2865 VDD.n3874 VDD.n204 146.341
R2866 VDD.n3870 VDD.n3869 146.341
R2867 VDD.n3867 VDD.n211 146.341
R2868 VDD.n3863 VDD.n3862 146.341
R2869 VDD.n3860 VDD.n218 146.341
R2870 VDD.n3856 VDD.n3855 146.341
R2871 VDD.n3853 VDD.n228 146.341
R2872 VDD.n3849 VDD.n3848 146.341
R2873 VDD.n3846 VDD.n235 146.341
R2874 VDD.n3609 VDD.n390 146.341
R2875 VDD.n3615 VDD.n390 146.341
R2876 VDD.n3615 VDD.n382 146.341
R2877 VDD.n3624 VDD.n382 146.341
R2878 VDD.n3624 VDD.n378 146.341
R2879 VDD.n3630 VDD.n378 146.341
R2880 VDD.n3630 VDD.n370 146.341
R2881 VDD.n3640 VDD.n370 146.341
R2882 VDD.n3640 VDD.n366 146.341
R2883 VDD.n3646 VDD.n366 146.341
R2884 VDD.n3646 VDD.n358 146.341
R2885 VDD.n3656 VDD.n358 146.341
R2886 VDD.n3656 VDD.n354 146.341
R2887 VDD.n3662 VDD.n354 146.341
R2888 VDD.n3662 VDD.n346 146.341
R2889 VDD.n3672 VDD.n346 146.341
R2890 VDD.n3672 VDD.n342 146.341
R2891 VDD.n3678 VDD.n342 146.341
R2892 VDD.n3678 VDD.n334 146.341
R2893 VDD.n3688 VDD.n334 146.341
R2894 VDD.n3688 VDD.n330 146.341
R2895 VDD.n3694 VDD.n330 146.341
R2896 VDD.n3694 VDD.n322 146.341
R2897 VDD.n3704 VDD.n322 146.341
R2898 VDD.n3704 VDD.n318 146.341
R2899 VDD.n3710 VDD.n318 146.341
R2900 VDD.n3710 VDD.n310 146.341
R2901 VDD.n3720 VDD.n310 146.341
R2902 VDD.n3720 VDD.n306 146.341
R2903 VDD.n3726 VDD.n306 146.341
R2904 VDD.n3726 VDD.n298 146.341
R2905 VDD.n3736 VDD.n298 146.341
R2906 VDD.n3736 VDD.n294 146.341
R2907 VDD.n3742 VDD.n294 146.341
R2908 VDD.n3742 VDD.n286 146.341
R2909 VDD.n3752 VDD.n286 146.341
R2910 VDD.n3752 VDD.n282 146.341
R2911 VDD.n3758 VDD.n282 146.341
R2912 VDD.n3758 VDD.n273 146.341
R2913 VDD.n3768 VDD.n273 146.341
R2914 VDD.n3768 VDD.n274 146.341
R2915 VDD.n274 VDD.n54 146.341
R2916 VDD.n55 VDD.n54 146.341
R2917 VDD.n56 VDD.n55 146.341
R2918 VDD.n267 VDD.n56 146.341
R2919 VDD.n267 VDD.n64 146.341
R2920 VDD.n65 VDD.n64 146.341
R2921 VDD.n66 VDD.n65 146.341
R2922 VDD.n264 VDD.n66 146.341
R2923 VDD.n264 VDD.n75 146.341
R2924 VDD.n76 VDD.n75 146.341
R2925 VDD.n77 VDD.n76 146.341
R2926 VDD.n261 VDD.n77 146.341
R2927 VDD.n261 VDD.n86 146.341
R2928 VDD.n87 VDD.n86 146.341
R2929 VDD.n88 VDD.n87 146.341
R2930 VDD.n258 VDD.n88 146.341
R2931 VDD.n258 VDD.n97 146.341
R2932 VDD.n98 VDD.n97 146.341
R2933 VDD.n99 VDD.n98 146.341
R2934 VDD.n255 VDD.n99 146.341
R2935 VDD.n255 VDD.n108 146.341
R2936 VDD.n109 VDD.n108 146.341
R2937 VDD.n110 VDD.n109 146.341
R2938 VDD.n252 VDD.n110 146.341
R2939 VDD.n252 VDD.n119 146.341
R2940 VDD.n120 VDD.n119 146.341
R2941 VDD.n121 VDD.n120 146.341
R2942 VDD.n249 VDD.n121 146.341
R2943 VDD.n249 VDD.n130 146.341
R2944 VDD.n131 VDD.n130 146.341
R2945 VDD.n132 VDD.n131 146.341
R2946 VDD.n246 VDD.n132 146.341
R2947 VDD.n246 VDD.n141 146.341
R2948 VDD.n142 VDD.n141 146.341
R2949 VDD.n143 VDD.n142 146.341
R2950 VDD.n243 VDD.n143 146.341
R2951 VDD.n243 VDD.n152 146.341
R2952 VDD.n153 VDD.n152 146.341
R2953 VDD.n154 VDD.n153 146.341
R2954 VDD.n240 VDD.n154 146.341
R2955 VDD.n240 VDD.n163 146.341
R2956 VDD.n164 VDD.n163 146.341
R2957 VDD.n165 VDD.n164 146.341
R2958 VDD.n3601 VDD.n3599 146.341
R2959 VDD.n3599 VDD.n3598 146.341
R2960 VDD.n3595 VDD.n3594 146.341
R2961 VDD.n3592 VDD.n3468 146.341
R2962 VDD.n3588 VDD.n3586 146.341
R2963 VDD.n3584 VDD.n3476 146.341
R2964 VDD.n3580 VDD.n3578 146.341
R2965 VDD.n3576 VDD.n3482 146.341
R2966 VDD.n3572 VDD.n3570 146.341
R2967 VDD.n3568 VDD.n3488 146.341
R2968 VDD.n3564 VDD.n3562 146.341
R2969 VDD.n3560 VDD.n3497 146.341
R2970 VDD.n3556 VDD.n3554 146.341
R2971 VDD.n3552 VDD.n3503 146.341
R2972 VDD.n3547 VDD.n3545 146.341
R2973 VDD.n3543 VDD.n3511 146.341
R2974 VDD.n3539 VDD.n3537 146.341
R2975 VDD.n3535 VDD.n3517 146.341
R2976 VDD.n3531 VDD.n3529 146.341
R2977 VDD.n3607 VDD.n388 146.341
R2978 VDD.n3617 VDD.n388 146.341
R2979 VDD.n3617 VDD.n384 146.341
R2980 VDD.n3623 VDD.n384 146.341
R2981 VDD.n3623 VDD.n376 146.341
R2982 VDD.n3632 VDD.n376 146.341
R2983 VDD.n3632 VDD.n372 146.341
R2984 VDD.n3638 VDD.n372 146.341
R2985 VDD.n3638 VDD.n364 146.341
R2986 VDD.n3648 VDD.n364 146.341
R2987 VDD.n3648 VDD.n360 146.341
R2988 VDD.n3654 VDD.n360 146.341
R2989 VDD.n3654 VDD.n352 146.341
R2990 VDD.n3664 VDD.n352 146.341
R2991 VDD.n3664 VDD.n348 146.341
R2992 VDD.n3670 VDD.n348 146.341
R2993 VDD.n3670 VDD.n340 146.341
R2994 VDD.n3680 VDD.n340 146.341
R2995 VDD.n3680 VDD.n336 146.341
R2996 VDD.n3686 VDD.n336 146.341
R2997 VDD.n3686 VDD.n328 146.341
R2998 VDD.n3696 VDD.n328 146.341
R2999 VDD.n3696 VDD.n324 146.341
R3000 VDD.n3702 VDD.n324 146.341
R3001 VDD.n3702 VDD.n316 146.341
R3002 VDD.n3712 VDD.n316 146.341
R3003 VDD.n3712 VDD.n312 146.341
R3004 VDD.n3718 VDD.n312 146.341
R3005 VDD.n3718 VDD.n304 146.341
R3006 VDD.n3728 VDD.n304 146.341
R3007 VDD.n3728 VDD.n300 146.341
R3008 VDD.n3734 VDD.n300 146.341
R3009 VDD.n3734 VDD.n292 146.341
R3010 VDD.n3744 VDD.n292 146.341
R3011 VDD.n3744 VDD.n288 146.341
R3012 VDD.n3750 VDD.n288 146.341
R3013 VDD.n3750 VDD.n280 146.341
R3014 VDD.n3760 VDD.n280 146.341
R3015 VDD.n3760 VDD.n276 146.341
R3016 VDD.n3766 VDD.n276 146.341
R3017 VDD.n3766 VDD.n51 146.341
R3018 VDD.n3998 VDD.n51 146.341
R3019 VDD.n3998 VDD.n52 146.341
R3020 VDD.n3994 VDD.n52 146.341
R3021 VDD.n3994 VDD.n58 146.341
R3022 VDD.n3990 VDD.n58 146.341
R3023 VDD.n3990 VDD.n63 146.341
R3024 VDD.n3986 VDD.n63 146.341
R3025 VDD.n3986 VDD.n68 146.341
R3026 VDD.n3982 VDD.n68 146.341
R3027 VDD.n3982 VDD.n74 146.341
R3028 VDD.n3978 VDD.n74 146.341
R3029 VDD.n3978 VDD.n79 146.341
R3030 VDD.n3974 VDD.n79 146.341
R3031 VDD.n3974 VDD.n85 146.341
R3032 VDD.n3970 VDD.n85 146.341
R3033 VDD.n3970 VDD.n90 146.341
R3034 VDD.n3966 VDD.n90 146.341
R3035 VDD.n3966 VDD.n96 146.341
R3036 VDD.n3962 VDD.n96 146.341
R3037 VDD.n3962 VDD.n101 146.341
R3038 VDD.n3958 VDD.n101 146.341
R3039 VDD.n3958 VDD.n107 146.341
R3040 VDD.n3954 VDD.n107 146.341
R3041 VDD.n3954 VDD.n112 146.341
R3042 VDD.n3950 VDD.n112 146.341
R3043 VDD.n3950 VDD.n118 146.341
R3044 VDD.n3946 VDD.n118 146.341
R3045 VDD.n3946 VDD.n123 146.341
R3046 VDD.n3942 VDD.n123 146.341
R3047 VDD.n3942 VDD.n129 146.341
R3048 VDD.n3938 VDD.n129 146.341
R3049 VDD.n3938 VDD.n134 146.341
R3050 VDD.n3934 VDD.n134 146.341
R3051 VDD.n3934 VDD.n140 146.341
R3052 VDD.n3930 VDD.n140 146.341
R3053 VDD.n3930 VDD.n145 146.341
R3054 VDD.n3926 VDD.n145 146.341
R3055 VDD.n3926 VDD.n151 146.341
R3056 VDD.n3923 VDD.n151 146.341
R3057 VDD.n3923 VDD.n156 146.341
R3058 VDD.n3919 VDD.n156 146.341
R3059 VDD.n3919 VDD.n162 146.341
R3060 VDD.n3915 VDD.n162 146.341
R3061 VDD.n2166 VDD.n1141 146.341
R3062 VDD.n2163 VDD.n1161 146.341
R3063 VDD.n2159 VDD.n2158 146.341
R3064 VDD.n2155 VDD.n2154 146.341
R3065 VDD.n2148 VDD.n2147 146.341
R3066 VDD.n2145 VDD.n2144 146.341
R3067 VDD.n2141 VDD.n2140 146.341
R3068 VDD.n2137 VDD.n2136 146.341
R3069 VDD.n2133 VDD.n2132 146.341
R3070 VDD.n2126 VDD.n2125 146.341
R3071 VDD.n2122 VDD.n2121 146.341
R3072 VDD.n2118 VDD.n2117 146.341
R3073 VDD.n2114 VDD.n2113 146.341
R3074 VDD.n2110 VDD.n2109 146.341
R3075 VDD.n2103 VDD.n2102 146.341
R3076 VDD.n2099 VDD.n2098 146.341
R3077 VDD.n2095 VDD.n2094 146.341
R3078 VDD.n2091 VDD.n2090 146.341
R3079 VDD.n2087 VDD.n2086 146.341
R3080 VDD.n1597 VDD.n1444 146.341
R3081 VDD.n1597 VDD.n1436 146.341
R3082 VDD.n1607 VDD.n1436 146.341
R3083 VDD.n1607 VDD.n1432 146.341
R3084 VDD.n1613 VDD.n1432 146.341
R3085 VDD.n1613 VDD.n1425 146.341
R3086 VDD.n1623 VDD.n1425 146.341
R3087 VDD.n1623 VDD.n1421 146.341
R3088 VDD.n1629 VDD.n1421 146.341
R3089 VDD.n1629 VDD.n1413 146.341
R3090 VDD.n1639 VDD.n1413 146.341
R3091 VDD.n1639 VDD.n1409 146.341
R3092 VDD.n1645 VDD.n1409 146.341
R3093 VDD.n1645 VDD.n1402 146.341
R3094 VDD.n1656 VDD.n1402 146.341
R3095 VDD.n1656 VDD.n1398 146.341
R3096 VDD.n1662 VDD.n1398 146.341
R3097 VDD.n1662 VDD.n1390 146.341
R3098 VDD.n1672 VDD.n1390 146.341
R3099 VDD.n1672 VDD.n1386 146.341
R3100 VDD.n1678 VDD.n1386 146.341
R3101 VDD.n1678 VDD.n1379 146.341
R3102 VDD.n1689 VDD.n1379 146.341
R3103 VDD.n1689 VDD.n1375 146.341
R3104 VDD.n1695 VDD.n1375 146.341
R3105 VDD.n1695 VDD.n1367 146.341
R3106 VDD.n1705 VDD.n1367 146.341
R3107 VDD.n1705 VDD.n1363 146.341
R3108 VDD.n1711 VDD.n1363 146.341
R3109 VDD.n1711 VDD.n1356 146.341
R3110 VDD.n1722 VDD.n1356 146.341
R3111 VDD.n1722 VDD.n1352 146.341
R3112 VDD.n1728 VDD.n1352 146.341
R3113 VDD.n1728 VDD.n1344 146.341
R3114 VDD.n1738 VDD.n1344 146.341
R3115 VDD.n1738 VDD.n1340 146.341
R3116 VDD.n1744 VDD.n1340 146.341
R3117 VDD.n1744 VDD.n1333 146.341
R3118 VDD.n1755 VDD.n1333 146.341
R3119 VDD.n1755 VDD.n1329 146.341
R3120 VDD.n1761 VDD.n1329 146.341
R3121 VDD.n1761 VDD.n1321 146.341
R3122 VDD.n1803 VDD.n1321 146.341
R3123 VDD.n1803 VDD.n1317 146.341
R3124 VDD.n1809 VDD.n1317 146.341
R3125 VDD.n1809 VDD.n1309 146.341
R3126 VDD.n1819 VDD.n1309 146.341
R3127 VDD.n1819 VDD.n1305 146.341
R3128 VDD.n1825 VDD.n1305 146.341
R3129 VDD.n1825 VDD.n1297 146.341
R3130 VDD.n1835 VDD.n1297 146.341
R3131 VDD.n1835 VDD.n1293 146.341
R3132 VDD.n1841 VDD.n1293 146.341
R3133 VDD.n1841 VDD.n1285 146.341
R3134 VDD.n1851 VDD.n1285 146.341
R3135 VDD.n1851 VDD.n1281 146.341
R3136 VDD.n1857 VDD.n1281 146.341
R3137 VDD.n1857 VDD.n1273 146.341
R3138 VDD.n1867 VDD.n1273 146.341
R3139 VDD.n1867 VDD.n1269 146.341
R3140 VDD.n1873 VDD.n1269 146.341
R3141 VDD.n1873 VDD.n1261 146.341
R3142 VDD.n1883 VDD.n1261 146.341
R3143 VDD.n1883 VDD.n1257 146.341
R3144 VDD.n1889 VDD.n1257 146.341
R3145 VDD.n1889 VDD.n1249 146.341
R3146 VDD.n1899 VDD.n1249 146.341
R3147 VDD.n1899 VDD.n1245 146.341
R3148 VDD.n1905 VDD.n1245 146.341
R3149 VDD.n1905 VDD.n1237 146.341
R3150 VDD.n1915 VDD.n1237 146.341
R3151 VDD.n1915 VDD.n1233 146.341
R3152 VDD.n1921 VDD.n1233 146.341
R3153 VDD.n1921 VDD.n1225 146.341
R3154 VDD.n1931 VDD.n1225 146.341
R3155 VDD.n1931 VDD.n1221 146.341
R3156 VDD.n1937 VDD.n1221 146.341
R3157 VDD.n1937 VDD.n1213 146.341
R3158 VDD.n1947 VDD.n1213 146.341
R3159 VDD.n1947 VDD.n1208 146.341
R3160 VDD.n1954 VDD.n1208 146.341
R3161 VDD.n1954 VDD.n1201 146.341
R3162 VDD.n1965 VDD.n1201 146.341
R3163 VDD.n1966 VDD.n1965 146.341
R3164 VDD.n1469 VDD.n1468 146.341
R3165 VDD.n1473 VDD.n1468 146.341
R3166 VDD.n1475 VDD.n1474 146.341
R3167 VDD.n1572 VDD.n1571 146.341
R3168 VDD.n1479 VDD.n1478 146.341
R3169 VDD.n1483 VDD.n1482 146.341
R3170 VDD.n1485 VDD.n1484 146.341
R3171 VDD.n1489 VDD.n1488 146.341
R3172 VDD.n1491 VDD.n1490 146.341
R3173 VDD.n1497 VDD.n1496 146.341
R3174 VDD.n1499 VDD.n1498 146.341
R3175 VDD.n1503 VDD.n1502 146.341
R3176 VDD.n1505 VDD.n1504 146.341
R3177 VDD.n1509 VDD.n1508 146.341
R3178 VDD.n1511 VDD.n1510 146.341
R3179 VDD.n1515 VDD.n1514 146.341
R3180 VDD.n1517 VDD.n1516 146.341
R3181 VDD.n1521 VDD.n1520 146.341
R3182 VDD.n1522 VDD.n1450 146.341
R3183 VDD.n1599 VDD.n1442 146.341
R3184 VDD.n1599 VDD.n1438 146.341
R3185 VDD.n1605 VDD.n1438 146.341
R3186 VDD.n1605 VDD.n1431 146.341
R3187 VDD.n1615 VDD.n1431 146.341
R3188 VDD.n1615 VDD.n1427 146.341
R3189 VDD.n1621 VDD.n1427 146.341
R3190 VDD.n1621 VDD.n1419 146.341
R3191 VDD.n1631 VDD.n1419 146.341
R3192 VDD.n1631 VDD.n1415 146.341
R3193 VDD.n1637 VDD.n1415 146.341
R3194 VDD.n1637 VDD.n1407 146.341
R3195 VDD.n1648 VDD.n1407 146.341
R3196 VDD.n1648 VDD.n1403 146.341
R3197 VDD.n1654 VDD.n1403 146.341
R3198 VDD.n1654 VDD.n1396 146.341
R3199 VDD.n1664 VDD.n1396 146.341
R3200 VDD.n1664 VDD.n1392 146.341
R3201 VDD.n1670 VDD.n1392 146.341
R3202 VDD.n1670 VDD.n1384 146.341
R3203 VDD.n1681 VDD.n1384 146.341
R3204 VDD.n1681 VDD.n1380 146.341
R3205 VDD.n1687 VDD.n1380 146.341
R3206 VDD.n1687 VDD.n1373 146.341
R3207 VDD.n1697 VDD.n1373 146.341
R3208 VDD.n1697 VDD.n1369 146.341
R3209 VDD.n1703 VDD.n1369 146.341
R3210 VDD.n1703 VDD.n1361 146.341
R3211 VDD.n1714 VDD.n1361 146.341
R3212 VDD.n1714 VDD.n1357 146.341
R3213 VDD.n1720 VDD.n1357 146.341
R3214 VDD.n1720 VDD.n1350 146.341
R3215 VDD.n1730 VDD.n1350 146.341
R3216 VDD.n1730 VDD.n1346 146.341
R3217 VDD.n1736 VDD.n1346 146.341
R3218 VDD.n1736 VDD.n1338 146.341
R3219 VDD.n1747 VDD.n1338 146.341
R3220 VDD.n1747 VDD.n1334 146.341
R3221 VDD.n1753 VDD.n1334 146.341
R3222 VDD.n1753 VDD.n1327 146.341
R3223 VDD.n1763 VDD.n1327 146.341
R3224 VDD.n1763 VDD.n1323 146.341
R3225 VDD.n1801 VDD.n1323 146.341
R3226 VDD.n1801 VDD.n1315 146.341
R3227 VDD.n1811 VDD.n1315 146.341
R3228 VDD.n1811 VDD.n1311 146.341
R3229 VDD.n1817 VDD.n1311 146.341
R3230 VDD.n1817 VDD.n1303 146.341
R3231 VDD.n1827 VDD.n1303 146.341
R3232 VDD.n1827 VDD.n1299 146.341
R3233 VDD.n1833 VDD.n1299 146.341
R3234 VDD.n1833 VDD.n1291 146.341
R3235 VDD.n1843 VDD.n1291 146.341
R3236 VDD.n1843 VDD.n1287 146.341
R3237 VDD.n1849 VDD.n1287 146.341
R3238 VDD.n1849 VDD.n1279 146.341
R3239 VDD.n1859 VDD.n1279 146.341
R3240 VDD.n1859 VDD.n1275 146.341
R3241 VDD.n1865 VDD.n1275 146.341
R3242 VDD.n1865 VDD.n1267 146.341
R3243 VDD.n1875 VDD.n1267 146.341
R3244 VDD.n1875 VDD.n1263 146.341
R3245 VDD.n1881 VDD.n1263 146.341
R3246 VDD.n1881 VDD.n1255 146.341
R3247 VDD.n1891 VDD.n1255 146.341
R3248 VDD.n1891 VDD.n1251 146.341
R3249 VDD.n1897 VDD.n1251 146.341
R3250 VDD.n1897 VDD.n1243 146.341
R3251 VDD.n1907 VDD.n1243 146.341
R3252 VDD.n1907 VDD.n1239 146.341
R3253 VDD.n1913 VDD.n1239 146.341
R3254 VDD.n1913 VDD.n1231 146.341
R3255 VDD.n1923 VDD.n1231 146.341
R3256 VDD.n1923 VDD.n1227 146.341
R3257 VDD.n1929 VDD.n1227 146.341
R3258 VDD.n1929 VDD.n1219 146.341
R3259 VDD.n1939 VDD.n1219 146.341
R3260 VDD.n1939 VDD.n1215 146.341
R3261 VDD.n1945 VDD.n1215 146.341
R3262 VDD.n1945 VDD.n1207 146.341
R3263 VDD.n1956 VDD.n1207 146.341
R3264 VDD.n1956 VDD.n1203 146.341
R3265 VDD.n1963 VDD.n1203 146.341
R3266 VDD.n1963 VDD.n1140 146.341
R3267 VDD.n9 VDD.n7 116.745
R3268 VDD.n2 VDD.n0 116.745
R3269 VDD.n9 VDD.n8 115.034
R3270 VDD.n11 VDD.n10 115.034
R3271 VDD.n13 VDD.n12 115.034
R3272 VDD.n6 VDD.n5 115.034
R3273 VDD.n4 VDD.n3 115.034
R3274 VDD.n2 VDD.n1 115.034
R3275 VDD.n1990 VDD.t6 113.427
R3276 VDD.n737 VDD.t56 113.427
R3277 VDD.n1046 VDD.t35 113.427
R3278 VDD.n748 VDD.t83 113.427
R3279 VDD.n2849 VDD.t76 113.427
R3280 VDD.n407 VDD.t43 113.427
R3281 VDD.n2725 VDD.t10 113.427
R3282 VDD.n446 VDD.t59 113.427
R3283 VDD.n3080 VDD.n2699 109.826
R3284 VDD.n3086 VDD.n705 99.5127
R3285 VDD.n3086 VDD.n695 99.5127
R3286 VDD.n3094 VDD.n695 99.5127
R3287 VDD.n3094 VDD.n693 99.5127
R3288 VDD.n3098 VDD.n693 99.5127
R3289 VDD.n3098 VDD.n684 99.5127
R3290 VDD.n3106 VDD.n684 99.5127
R3291 VDD.n3106 VDD.n682 99.5127
R3292 VDD.n3110 VDD.n682 99.5127
R3293 VDD.n3110 VDD.n672 99.5127
R3294 VDD.n3118 VDD.n672 99.5127
R3295 VDD.n3118 VDD.n670 99.5127
R3296 VDD.n3122 VDD.n670 99.5127
R3297 VDD.n3122 VDD.n659 99.5127
R3298 VDD.n3130 VDD.n659 99.5127
R3299 VDD.n3130 VDD.n657 99.5127
R3300 VDD.n3134 VDD.n657 99.5127
R3301 VDD.n3134 VDD.n648 99.5127
R3302 VDD.n3142 VDD.n648 99.5127
R3303 VDD.n3142 VDD.n646 99.5127
R3304 VDD.n3146 VDD.n646 99.5127
R3305 VDD.n3146 VDD.n636 99.5127
R3306 VDD.n3154 VDD.n636 99.5127
R3307 VDD.n3154 VDD.n634 99.5127
R3308 VDD.n3158 VDD.n634 99.5127
R3309 VDD.n3158 VDD.n623 99.5127
R3310 VDD.n3166 VDD.n623 99.5127
R3311 VDD.n3166 VDD.n621 99.5127
R3312 VDD.n3170 VDD.n621 99.5127
R3313 VDD.n3170 VDD.n612 99.5127
R3314 VDD.n3178 VDD.n612 99.5127
R3315 VDD.n3178 VDD.n610 99.5127
R3316 VDD.n3182 VDD.n610 99.5127
R3317 VDD.n3182 VDD.n600 99.5127
R3318 VDD.n3190 VDD.n600 99.5127
R3319 VDD.n3190 VDD.n598 99.5127
R3320 VDD.n3194 VDD.n598 99.5127
R3321 VDD.n3194 VDD.n587 99.5127
R3322 VDD.n3202 VDD.n587 99.5127
R3323 VDD.n3202 VDD.n585 99.5127
R3324 VDD.n3206 VDD.n585 99.5127
R3325 VDD.n3206 VDD.n576 99.5127
R3326 VDD.n3214 VDD.n576 99.5127
R3327 VDD.n3214 VDD.n574 99.5127
R3328 VDD.n3218 VDD.n574 99.5127
R3329 VDD.n3218 VDD.n564 99.5127
R3330 VDD.n3225 VDD.n564 99.5127
R3331 VDD.n3225 VDD.n562 99.5127
R3332 VDD.n3229 VDD.n562 99.5127
R3333 VDD.n3229 VDD.n552 99.5127
R3334 VDD.n3237 VDD.n552 99.5127
R3335 VDD.n3237 VDD.n550 99.5127
R3336 VDD.n3241 VDD.n550 99.5127
R3337 VDD.n3241 VDD.n539 99.5127
R3338 VDD.n3249 VDD.n539 99.5127
R3339 VDD.n3249 VDD.n537 99.5127
R3340 VDD.n3253 VDD.n537 99.5127
R3341 VDD.n3253 VDD.n528 99.5127
R3342 VDD.n3261 VDD.n528 99.5127
R3343 VDD.n3261 VDD.n526 99.5127
R3344 VDD.n3265 VDD.n526 99.5127
R3345 VDD.n3265 VDD.n516 99.5127
R3346 VDD.n3273 VDD.n516 99.5127
R3347 VDD.n3273 VDD.n514 99.5127
R3348 VDD.n3277 VDD.n514 99.5127
R3349 VDD.n3277 VDD.n503 99.5127
R3350 VDD.n3285 VDD.n503 99.5127
R3351 VDD.n3285 VDD.n501 99.5127
R3352 VDD.n3289 VDD.n501 99.5127
R3353 VDD.n3289 VDD.n492 99.5127
R3354 VDD.n3297 VDD.n492 99.5127
R3355 VDD.n3297 VDD.n490 99.5127
R3356 VDD.n3301 VDD.n490 99.5127
R3357 VDD.n3301 VDD.n480 99.5127
R3358 VDD.n3309 VDD.n480 99.5127
R3359 VDD.n3309 VDD.n478 99.5127
R3360 VDD.n3313 VDD.n478 99.5127
R3361 VDD.n3313 VDD.n468 99.5127
R3362 VDD.n3321 VDD.n468 99.5127
R3363 VDD.n3321 VDD.n466 99.5127
R3364 VDD.n3325 VDD.n466 99.5127
R3365 VDD.n3325 VDD.n455 99.5127
R3366 VDD.n3335 VDD.n455 99.5127
R3367 VDD.n3335 VDD.n453 99.5127
R3368 VDD.n3339 VDD.n453 99.5127
R3369 VDD.n3339 VDD.n420 99.5127
R3370 VDD.n3400 VDD.n420 99.5127
R3371 VDD.n3400 VDD.n417 99.5127
R3372 VDD.n3433 VDD.n417 99.5127
R3373 VDD.n3433 VDD.n418 99.5127
R3374 VDD.n3427 VDD.n3426 99.5127
R3375 VDD.n3424 VDD.n3405 99.5127
R3376 VDD.n3420 VDD.n3419 99.5127
R3377 VDD.n3417 VDD.n3408 99.5127
R3378 VDD.n3413 VDD.n3412 99.5127
R3379 VDD.n3459 VDD.n399 99.5127
R3380 VDD.n3457 VDD.n3456 99.5127
R3381 VDD.n3454 VDD.n402 99.5127
R3382 VDD.n3450 VDD.n3449 99.5127
R3383 VDD.n3447 VDD.n405 99.5127
R3384 VDD.n3442 VDD.n3441 99.5127
R3385 VDD.n3036 VDD.n703 99.5127
R3386 VDD.n3033 VDD.n703 99.5127
R3387 VDD.n3033 VDD.n697 99.5127
R3388 VDD.n3030 VDD.n697 99.5127
R3389 VDD.n3030 VDD.n691 99.5127
R3390 VDD.n3027 VDD.n691 99.5127
R3391 VDD.n3027 VDD.n685 99.5127
R3392 VDD.n2845 VDD.n685 99.5127
R3393 VDD.n2845 VDD.n680 99.5127
R3394 VDD.n2842 VDD.n680 99.5127
R3395 VDD.n2842 VDD.n674 99.5127
R3396 VDD.n2839 VDD.n674 99.5127
R3397 VDD.n2839 VDD.n668 99.5127
R3398 VDD.n2836 VDD.n668 99.5127
R3399 VDD.n2836 VDD.n661 99.5127
R3400 VDD.n2833 VDD.n661 99.5127
R3401 VDD.n2833 VDD.n655 99.5127
R3402 VDD.n2830 VDD.n655 99.5127
R3403 VDD.n2830 VDD.n650 99.5127
R3404 VDD.n2827 VDD.n650 99.5127
R3405 VDD.n2827 VDD.n644 99.5127
R3406 VDD.n2824 VDD.n644 99.5127
R3407 VDD.n2824 VDD.n638 99.5127
R3408 VDD.n2821 VDD.n638 99.5127
R3409 VDD.n2821 VDD.n632 99.5127
R3410 VDD.n2818 VDD.n632 99.5127
R3411 VDD.n2818 VDD.n625 99.5127
R3412 VDD.n2815 VDD.n625 99.5127
R3413 VDD.n2815 VDD.n619 99.5127
R3414 VDD.n2812 VDD.n619 99.5127
R3415 VDD.n2812 VDD.n614 99.5127
R3416 VDD.n2809 VDD.n614 99.5127
R3417 VDD.n2809 VDD.n608 99.5127
R3418 VDD.n2806 VDD.n608 99.5127
R3419 VDD.n2806 VDD.n602 99.5127
R3420 VDD.n2803 VDD.n602 99.5127
R3421 VDD.n2803 VDD.n596 99.5127
R3422 VDD.n2800 VDD.n596 99.5127
R3423 VDD.n2800 VDD.n589 99.5127
R3424 VDD.n2797 VDD.n589 99.5127
R3425 VDD.n2797 VDD.n583 99.5127
R3426 VDD.n2794 VDD.n583 99.5127
R3427 VDD.n2794 VDD.n578 99.5127
R3428 VDD.n2791 VDD.n578 99.5127
R3429 VDD.n2791 VDD.n573 99.5127
R3430 VDD.n2788 VDD.n573 99.5127
R3431 VDD.n2788 VDD.n566 99.5127
R3432 VDD.n2785 VDD.n566 99.5127
R3433 VDD.n2785 VDD.n560 99.5127
R3434 VDD.n2782 VDD.n560 99.5127
R3435 VDD.n2782 VDD.n554 99.5127
R3436 VDD.n2779 VDD.n554 99.5127
R3437 VDD.n2779 VDD.n548 99.5127
R3438 VDD.n2776 VDD.n548 99.5127
R3439 VDD.n2776 VDD.n541 99.5127
R3440 VDD.n2773 VDD.n541 99.5127
R3441 VDD.n2773 VDD.n535 99.5127
R3442 VDD.n2770 VDD.n535 99.5127
R3443 VDD.n2770 VDD.n530 99.5127
R3444 VDD.n2767 VDD.n530 99.5127
R3445 VDD.n2767 VDD.n524 99.5127
R3446 VDD.n2764 VDD.n524 99.5127
R3447 VDD.n2764 VDD.n518 99.5127
R3448 VDD.n2761 VDD.n518 99.5127
R3449 VDD.n2761 VDD.n512 99.5127
R3450 VDD.n2758 VDD.n512 99.5127
R3451 VDD.n2758 VDD.n505 99.5127
R3452 VDD.n2755 VDD.n505 99.5127
R3453 VDD.n2755 VDD.n499 99.5127
R3454 VDD.n2752 VDD.n499 99.5127
R3455 VDD.n2752 VDD.n494 99.5127
R3456 VDD.n2749 VDD.n494 99.5127
R3457 VDD.n2749 VDD.n488 99.5127
R3458 VDD.n2746 VDD.n488 99.5127
R3459 VDD.n2746 VDD.n482 99.5127
R3460 VDD.n2743 VDD.n482 99.5127
R3461 VDD.n2743 VDD.n476 99.5127
R3462 VDD.n2740 VDD.n476 99.5127
R3463 VDD.n2740 VDD.n470 99.5127
R3464 VDD.n2737 VDD.n470 99.5127
R3465 VDD.n2737 VDD.n464 99.5127
R3466 VDD.n2734 VDD.n464 99.5127
R3467 VDD.n2734 VDD.n457 99.5127
R3468 VDD.n2731 VDD.n457 99.5127
R3469 VDD.n2731 VDD.n451 99.5127
R3470 VDD.n2728 VDD.n451 99.5127
R3471 VDD.n2728 VDD.n422 99.5127
R3472 VDD.n422 VDD.n412 99.5127
R3473 VDD.n3435 VDD.n412 99.5127
R3474 VDD.n3435 VDD.n410 99.5127
R3475 VDD.n3079 VDD.n707 99.5127
R3476 VDD.n3079 VDD.n2723 99.5127
R3477 VDD.n3075 VDD.n3074 99.5127
R3478 VDD.n3071 VDD.n3070 99.5127
R3479 VDD.n3067 VDD.n3066 99.5127
R3480 VDD.n3063 VDD.n3062 99.5127
R3481 VDD.n3059 VDD.n3058 99.5127
R3482 VDD.n3055 VDD.n3054 99.5127
R3483 VDD.n3051 VDD.n3050 99.5127
R3484 VDD.n3047 VDD.n3046 99.5127
R3485 VDD.n3043 VDD.n3042 99.5127
R3486 VDD.n3039 VDD.n2710 99.5127
R3487 VDD.n2642 VDD.n2641 99.5127
R3488 VDD.n2638 VDD.n2637 99.5127
R3489 VDD.n2634 VDD.n2633 99.5127
R3490 VDD.n2630 VDD.n2629 99.5127
R3491 VDD.n2626 VDD.n2625 99.5127
R3492 VDD.n2622 VDD.n2621 99.5127
R3493 VDD.n2618 VDD.n2617 99.5127
R3494 VDD.n2614 VDD.n2613 99.5127
R3495 VDD.n2610 VDD.n2609 99.5127
R3496 VDD.n2606 VDD.n2605 99.5127
R3497 VDD.n2601 VDD.n2600 99.5127
R3498 VDD.n1112 VDD.n1015 99.5127
R3499 VDD.n1109 VDD.n1015 99.5127
R3500 VDD.n1109 VDD.n1009 99.5127
R3501 VDD.n1106 VDD.n1009 99.5127
R3502 VDD.n1106 VDD.n1002 99.5127
R3503 VDD.n1103 VDD.n1002 99.5127
R3504 VDD.n1103 VDD.n995 99.5127
R3505 VDD.n1100 VDD.n995 99.5127
R3506 VDD.n1100 VDD.n990 99.5127
R3507 VDD.n1097 VDD.n990 99.5127
R3508 VDD.n1097 VDD.n985 99.5127
R3509 VDD.n1094 VDD.n985 99.5127
R3510 VDD.n1094 VDD.n979 99.5127
R3511 VDD.n1091 VDD.n979 99.5127
R3512 VDD.n1091 VDD.n973 99.5127
R3513 VDD.n1088 VDD.n973 99.5127
R3514 VDD.n1088 VDD.n967 99.5127
R3515 VDD.n1085 VDD.n967 99.5127
R3516 VDD.n1085 VDD.n960 99.5127
R3517 VDD.n1082 VDD.n960 99.5127
R3518 VDD.n1082 VDD.n954 99.5127
R3519 VDD.n1079 VDD.n954 99.5127
R3520 VDD.n1079 VDD.n949 99.5127
R3521 VDD.n1076 VDD.n949 99.5127
R3522 VDD.n1076 VDD.n943 99.5127
R3523 VDD.n1073 VDD.n943 99.5127
R3524 VDD.n1073 VDD.n937 99.5127
R3525 VDD.n1070 VDD.n937 99.5127
R3526 VDD.n1070 VDD.n931 99.5127
R3527 VDD.n1067 VDD.n931 99.5127
R3528 VDD.n1067 VDD.n924 99.5127
R3529 VDD.n1064 VDD.n924 99.5127
R3530 VDD.n1064 VDD.n918 99.5127
R3531 VDD.n1061 VDD.n918 99.5127
R3532 VDD.n1061 VDD.n913 99.5127
R3533 VDD.n1058 VDD.n913 99.5127
R3534 VDD.n1058 VDD.n907 99.5127
R3535 VDD.n1055 VDD.n907 99.5127
R3536 VDD.n1055 VDD.n901 99.5127
R3537 VDD.n1052 VDD.n901 99.5127
R3538 VDD.n1052 VDD.n894 99.5127
R3539 VDD.n1049 VDD.n894 99.5127
R3540 VDD.n1049 VDD.n888 99.5127
R3541 VDD.n888 VDD.n880 99.5127
R3542 VDD.n2459 VDD.n880 99.5127
R3543 VDD.n2459 VDD.n881 99.5127
R3544 VDD.n881 VDD.n872 99.5127
R3545 VDD.n2454 VDD.n872 99.5127
R3546 VDD.n2454 VDD.n866 99.5127
R3547 VDD.n2451 VDD.n866 99.5127
R3548 VDD.n2451 VDD.n860 99.5127
R3549 VDD.n2448 VDD.n860 99.5127
R3550 VDD.n2448 VDD.n854 99.5127
R3551 VDD.n2445 VDD.n854 99.5127
R3552 VDD.n2445 VDD.n847 99.5127
R3553 VDD.n2442 VDD.n847 99.5127
R3554 VDD.n2442 VDD.n841 99.5127
R3555 VDD.n2439 VDD.n841 99.5127
R3556 VDD.n2439 VDD.n836 99.5127
R3557 VDD.n2436 VDD.n836 99.5127
R3558 VDD.n2436 VDD.n830 99.5127
R3559 VDD.n2433 VDD.n830 99.5127
R3560 VDD.n2433 VDD.n824 99.5127
R3561 VDD.n2430 VDD.n824 99.5127
R3562 VDD.n2430 VDD.n818 99.5127
R3563 VDD.n2427 VDD.n818 99.5127
R3564 VDD.n2427 VDD.n811 99.5127
R3565 VDD.n2424 VDD.n811 99.5127
R3566 VDD.n2424 VDD.n805 99.5127
R3567 VDD.n2421 VDD.n805 99.5127
R3568 VDD.n2421 VDD.n800 99.5127
R3569 VDD.n2418 VDD.n800 99.5127
R3570 VDD.n2418 VDD.n794 99.5127
R3571 VDD.n2415 VDD.n794 99.5127
R3572 VDD.n2415 VDD.n788 99.5127
R3573 VDD.n2412 VDD.n788 99.5127
R3574 VDD.n2412 VDD.n782 99.5127
R3575 VDD.n2409 VDD.n782 99.5127
R3576 VDD.n2409 VDD.n776 99.5127
R3577 VDD.n2406 VDD.n776 99.5127
R3578 VDD.n2406 VDD.n770 99.5127
R3579 VDD.n2403 VDD.n770 99.5127
R3580 VDD.n2403 VDD.n764 99.5127
R3581 VDD.n2400 VDD.n764 99.5127
R3582 VDD.n2400 VDD.n757 99.5127
R3583 VDD.n757 VDD.n750 99.5127
R3584 VDD.n2591 VDD.n750 99.5127
R3585 VDD.n2592 VDD.n2591 99.5127
R3586 VDD.n2592 VDD.n742 99.5127
R3587 VDD.n2596 VDD.n742 99.5127
R3588 VDD.n1044 VDD.n1043 99.5127
R3589 VDD.n2186 VDD.n1043 99.5127
R3590 VDD.n2184 VDD.n2183 99.5127
R3591 VDD.n2180 VDD.n2179 99.5127
R3592 VDD.n2176 VDD.n2175 99.5127
R3593 VDD.n2172 VDD.n2171 99.5127
R3594 VDD.n1135 VDD.n1134 99.5127
R3595 VDD.n1131 VDD.n1130 99.5127
R3596 VDD.n1127 VDD.n1126 99.5127
R3597 VDD.n1123 VDD.n1122 99.5127
R3598 VDD.n1119 VDD.n1118 99.5127
R3599 VDD.n1115 VDD.n1030 99.5127
R3600 VDD.n2200 VDD.n1013 99.5127
R3601 VDD.n2200 VDD.n1011 99.5127
R3602 VDD.n2204 VDD.n1011 99.5127
R3603 VDD.n2204 VDD.n1000 99.5127
R3604 VDD.n2212 VDD.n1000 99.5127
R3605 VDD.n2212 VDD.n998 99.5127
R3606 VDD.n2216 VDD.n998 99.5127
R3607 VDD.n2216 VDD.n989 99.5127
R3608 VDD.n2224 VDD.n989 99.5127
R3609 VDD.n2224 VDD.n987 99.5127
R3610 VDD.n2228 VDD.n987 99.5127
R3611 VDD.n2228 VDD.n977 99.5127
R3612 VDD.n2236 VDD.n977 99.5127
R3613 VDD.n2236 VDD.n975 99.5127
R3614 VDD.n2240 VDD.n975 99.5127
R3615 VDD.n2240 VDD.n965 99.5127
R3616 VDD.n2248 VDD.n965 99.5127
R3617 VDD.n2248 VDD.n963 99.5127
R3618 VDD.n2252 VDD.n963 99.5127
R3619 VDD.n2252 VDD.n953 99.5127
R3620 VDD.n2260 VDD.n953 99.5127
R3621 VDD.n2260 VDD.n951 99.5127
R3622 VDD.n2264 VDD.n951 99.5127
R3623 VDD.n2264 VDD.n941 99.5127
R3624 VDD.n2272 VDD.n941 99.5127
R3625 VDD.n2272 VDD.n939 99.5127
R3626 VDD.n2276 VDD.n939 99.5127
R3627 VDD.n2276 VDD.n929 99.5127
R3628 VDD.n2284 VDD.n929 99.5127
R3629 VDD.n2284 VDD.n927 99.5127
R3630 VDD.n2288 VDD.n927 99.5127
R3631 VDD.n2288 VDD.n917 99.5127
R3632 VDD.n2296 VDD.n917 99.5127
R3633 VDD.n2296 VDD.n915 99.5127
R3634 VDD.n2300 VDD.n915 99.5127
R3635 VDD.n2300 VDD.n905 99.5127
R3636 VDD.n2308 VDD.n905 99.5127
R3637 VDD.n2308 VDD.n903 99.5127
R3638 VDD.n2312 VDD.n903 99.5127
R3639 VDD.n2312 VDD.n892 99.5127
R3640 VDD.n2325 VDD.n892 99.5127
R3641 VDD.n2325 VDD.n890 99.5127
R3642 VDD.n2329 VDD.n890 99.5127
R3643 VDD.n2329 VDD.n876 99.5127
R3644 VDD.n2460 VDD.n876 99.5127
R3645 VDD.n2460 VDD.n874 99.5127
R3646 VDD.n2464 VDD.n874 99.5127
R3647 VDD.n2464 VDD.n864 99.5127
R3648 VDD.n2472 VDD.n864 99.5127
R3649 VDD.n2472 VDD.n862 99.5127
R3650 VDD.n2476 VDD.n862 99.5127
R3651 VDD.n2476 VDD.n852 99.5127
R3652 VDD.n2484 VDD.n852 99.5127
R3653 VDD.n2484 VDD.n850 99.5127
R3654 VDD.n2488 VDD.n850 99.5127
R3655 VDD.n2488 VDD.n840 99.5127
R3656 VDD.n2496 VDD.n840 99.5127
R3657 VDD.n2496 VDD.n838 99.5127
R3658 VDD.n2500 VDD.n838 99.5127
R3659 VDD.n2500 VDD.n828 99.5127
R3660 VDD.n2508 VDD.n828 99.5127
R3661 VDD.n2508 VDD.n826 99.5127
R3662 VDD.n2512 VDD.n826 99.5127
R3663 VDD.n2512 VDD.n816 99.5127
R3664 VDD.n2520 VDD.n816 99.5127
R3665 VDD.n2520 VDD.n814 99.5127
R3666 VDD.n2524 VDD.n814 99.5127
R3667 VDD.n2524 VDD.n804 99.5127
R3668 VDD.n2532 VDD.n804 99.5127
R3669 VDD.n2532 VDD.n802 99.5127
R3670 VDD.n2536 VDD.n802 99.5127
R3671 VDD.n2536 VDD.n792 99.5127
R3672 VDD.n2544 VDD.n792 99.5127
R3673 VDD.n2544 VDD.n790 99.5127
R3674 VDD.n2548 VDD.n790 99.5127
R3675 VDD.n2548 VDD.n780 99.5127
R3676 VDD.n2556 VDD.n780 99.5127
R3677 VDD.n2556 VDD.n778 99.5127
R3678 VDD.n2560 VDD.n778 99.5127
R3679 VDD.n2560 VDD.n768 99.5127
R3680 VDD.n2568 VDD.n768 99.5127
R3681 VDD.n2568 VDD.n766 99.5127
R3682 VDD.n2572 VDD.n766 99.5127
R3683 VDD.n2572 VDD.n756 99.5127
R3684 VDD.n2585 VDD.n756 99.5127
R3685 VDD.n2585 VDD.n754 99.5127
R3686 VDD.n2589 VDD.n754 99.5127
R3687 VDD.n2589 VDD.n744 99.5127
R3688 VDD.n2648 VDD.n744 99.5127
R3689 VDD.n2648 VDD.n745 99.5127
R3690 VDD.n3390 VDD.n428 99.5127
R3691 VDD.n3386 VDD.n3385 99.5127
R3692 VDD.n3383 VDD.n431 99.5127
R3693 VDD.n3379 VDD.n3378 99.5127
R3694 VDD.n3376 VDD.n434 99.5127
R3695 VDD.n3372 VDD.n3371 99.5127
R3696 VDD.n3369 VDD.n438 99.5127
R3697 VDD.n3365 VDD.n3364 99.5127
R3698 VDD.n3362 VDD.n441 99.5127
R3699 VDD.n3358 VDD.n3357 99.5127
R3700 VDD.n3355 VDD.n444 99.5127
R3701 VDD.n2899 VDD.n704 99.5127
R3702 VDD.n2902 VDD.n704 99.5127
R3703 VDD.n2902 VDD.n698 99.5127
R3704 VDD.n2905 VDD.n698 99.5127
R3705 VDD.n2905 VDD.n692 99.5127
R3706 VDD.n3025 VDD.n692 99.5127
R3707 VDD.n3025 VDD.n686 99.5127
R3708 VDD.n3021 VDD.n686 99.5127
R3709 VDD.n3021 VDD.n681 99.5127
R3710 VDD.n3018 VDD.n681 99.5127
R3711 VDD.n3018 VDD.n675 99.5127
R3712 VDD.n3015 VDD.n675 99.5127
R3713 VDD.n3015 VDD.n669 99.5127
R3714 VDD.n3012 VDD.n669 99.5127
R3715 VDD.n3012 VDD.n662 99.5127
R3716 VDD.n3009 VDD.n662 99.5127
R3717 VDD.n3009 VDD.n656 99.5127
R3718 VDD.n3006 VDD.n656 99.5127
R3719 VDD.n3006 VDD.n651 99.5127
R3720 VDD.n3003 VDD.n651 99.5127
R3721 VDD.n3003 VDD.n645 99.5127
R3722 VDD.n3000 VDD.n645 99.5127
R3723 VDD.n3000 VDD.n639 99.5127
R3724 VDD.n2997 VDD.n639 99.5127
R3725 VDD.n2997 VDD.n633 99.5127
R3726 VDD.n2994 VDD.n633 99.5127
R3727 VDD.n2994 VDD.n626 99.5127
R3728 VDD.n2991 VDD.n626 99.5127
R3729 VDD.n2991 VDD.n620 99.5127
R3730 VDD.n2988 VDD.n620 99.5127
R3731 VDD.n2988 VDD.n615 99.5127
R3732 VDD.n2985 VDD.n615 99.5127
R3733 VDD.n2985 VDD.n609 99.5127
R3734 VDD.n2982 VDD.n609 99.5127
R3735 VDD.n2982 VDD.n603 99.5127
R3736 VDD.n2979 VDD.n603 99.5127
R3737 VDD.n2979 VDD.n597 99.5127
R3738 VDD.n2976 VDD.n597 99.5127
R3739 VDD.n2976 VDD.n590 99.5127
R3740 VDD.n2973 VDD.n590 99.5127
R3741 VDD.n2973 VDD.n584 99.5127
R3742 VDD.n2970 VDD.n584 99.5127
R3743 VDD.n2970 VDD.n579 99.5127
R3744 VDD.n2967 VDD.n579 99.5127
R3745 VDD.n2967 VDD.n572 99.5127
R3746 VDD.n2964 VDD.n572 99.5127
R3747 VDD.n2964 VDD.n567 99.5127
R3748 VDD.n2961 VDD.n567 99.5127
R3749 VDD.n2961 VDD.n561 99.5127
R3750 VDD.n2958 VDD.n561 99.5127
R3751 VDD.n2958 VDD.n555 99.5127
R3752 VDD.n2955 VDD.n555 99.5127
R3753 VDD.n2955 VDD.n549 99.5127
R3754 VDD.n2952 VDD.n549 99.5127
R3755 VDD.n2952 VDD.n542 99.5127
R3756 VDD.n2949 VDD.n542 99.5127
R3757 VDD.n2949 VDD.n536 99.5127
R3758 VDD.n2946 VDD.n536 99.5127
R3759 VDD.n2946 VDD.n531 99.5127
R3760 VDD.n2943 VDD.n531 99.5127
R3761 VDD.n2943 VDD.n525 99.5127
R3762 VDD.n2940 VDD.n525 99.5127
R3763 VDD.n2940 VDD.n519 99.5127
R3764 VDD.n2937 VDD.n519 99.5127
R3765 VDD.n2937 VDD.n513 99.5127
R3766 VDD.n2934 VDD.n513 99.5127
R3767 VDD.n2934 VDD.n506 99.5127
R3768 VDD.n2931 VDD.n506 99.5127
R3769 VDD.n2931 VDD.n500 99.5127
R3770 VDD.n2928 VDD.n500 99.5127
R3771 VDD.n2928 VDD.n495 99.5127
R3772 VDD.n2925 VDD.n495 99.5127
R3773 VDD.n2925 VDD.n489 99.5127
R3774 VDD.n2922 VDD.n489 99.5127
R3775 VDD.n2922 VDD.n483 99.5127
R3776 VDD.n2919 VDD.n483 99.5127
R3777 VDD.n2919 VDD.n477 99.5127
R3778 VDD.n2916 VDD.n477 99.5127
R3779 VDD.n2916 VDD.n471 99.5127
R3780 VDD.n2913 VDD.n471 99.5127
R3781 VDD.n2913 VDD.n465 99.5127
R3782 VDD.n2910 VDD.n465 99.5127
R3783 VDD.n2910 VDD.n458 99.5127
R3784 VDD.n458 VDD.n449 99.5127
R3785 VDD.n3341 VDD.n449 99.5127
R3786 VDD.n3342 VDD.n3341 99.5127
R3787 VDD.n3342 VDD.n423 99.5127
R3788 VDD.n3345 VDD.n423 99.5127
R3789 VDD.n3345 VDD.n414 99.5127
R3790 VDD.n3350 VDD.n414 99.5127
R3791 VDD.n2854 VDD.n2853 99.5127
R3792 VDD.n2858 VDD.n2857 99.5127
R3793 VDD.n2862 VDD.n2861 99.5127
R3794 VDD.n2866 VDD.n2865 99.5127
R3795 VDD.n2870 VDD.n2869 99.5127
R3796 VDD.n2874 VDD.n2873 99.5127
R3797 VDD.n2878 VDD.n2877 99.5127
R3798 VDD.n2882 VDD.n2881 99.5127
R3799 VDD.n2886 VDD.n2885 99.5127
R3800 VDD.n2890 VDD.n2889 99.5127
R3801 VDD.n2895 VDD.n2894 99.5127
R3802 VDD.n3088 VDD.n701 99.5127
R3803 VDD.n3088 VDD.n699 99.5127
R3804 VDD.n3092 VDD.n699 99.5127
R3805 VDD.n3092 VDD.n689 99.5127
R3806 VDD.n3100 VDD.n689 99.5127
R3807 VDD.n3100 VDD.n687 99.5127
R3808 VDD.n3104 VDD.n687 99.5127
R3809 VDD.n3104 VDD.n678 99.5127
R3810 VDD.n3112 VDD.n678 99.5127
R3811 VDD.n3112 VDD.n676 99.5127
R3812 VDD.n3116 VDD.n676 99.5127
R3813 VDD.n3116 VDD.n666 99.5127
R3814 VDD.n3124 VDD.n666 99.5127
R3815 VDD.n3124 VDD.n664 99.5127
R3816 VDD.n3128 VDD.n664 99.5127
R3817 VDD.n3128 VDD.n654 99.5127
R3818 VDD.n3136 VDD.n654 99.5127
R3819 VDD.n3136 VDD.n652 99.5127
R3820 VDD.n3140 VDD.n652 99.5127
R3821 VDD.n3140 VDD.n642 99.5127
R3822 VDD.n3148 VDD.n642 99.5127
R3823 VDD.n3148 VDD.n640 99.5127
R3824 VDD.n3152 VDD.n640 99.5127
R3825 VDD.n3152 VDD.n630 99.5127
R3826 VDD.n3160 VDD.n630 99.5127
R3827 VDD.n3160 VDD.n628 99.5127
R3828 VDD.n3164 VDD.n628 99.5127
R3829 VDD.n3164 VDD.n618 99.5127
R3830 VDD.n3172 VDD.n618 99.5127
R3831 VDD.n3172 VDD.n616 99.5127
R3832 VDD.n3176 VDD.n616 99.5127
R3833 VDD.n3176 VDD.n606 99.5127
R3834 VDD.n3184 VDD.n606 99.5127
R3835 VDD.n3184 VDD.n604 99.5127
R3836 VDD.n3188 VDD.n604 99.5127
R3837 VDD.n3188 VDD.n594 99.5127
R3838 VDD.n3196 VDD.n594 99.5127
R3839 VDD.n3196 VDD.n592 99.5127
R3840 VDD.n3200 VDD.n592 99.5127
R3841 VDD.n3200 VDD.n582 99.5127
R3842 VDD.n3208 VDD.n582 99.5127
R3843 VDD.n3208 VDD.n580 99.5127
R3844 VDD.n3212 VDD.n580 99.5127
R3845 VDD.n3212 VDD.n570 99.5127
R3846 VDD.n3219 VDD.n570 99.5127
R3847 VDD.n3219 VDD.n568 99.5127
R3848 VDD.n3223 VDD.n568 99.5127
R3849 VDD.n3223 VDD.n558 99.5127
R3850 VDD.n3231 VDD.n558 99.5127
R3851 VDD.n3231 VDD.n556 99.5127
R3852 VDD.n3235 VDD.n556 99.5127
R3853 VDD.n3235 VDD.n546 99.5127
R3854 VDD.n3243 VDD.n546 99.5127
R3855 VDD.n3243 VDD.n544 99.5127
R3856 VDD.n3247 VDD.n544 99.5127
R3857 VDD.n3247 VDD.n534 99.5127
R3858 VDD.n3255 VDD.n534 99.5127
R3859 VDD.n3255 VDD.n532 99.5127
R3860 VDD.n3259 VDD.n532 99.5127
R3861 VDD.n3259 VDD.n522 99.5127
R3862 VDD.n3267 VDD.n522 99.5127
R3863 VDD.n3267 VDD.n520 99.5127
R3864 VDD.n3271 VDD.n520 99.5127
R3865 VDD.n3271 VDD.n510 99.5127
R3866 VDD.n3279 VDD.n510 99.5127
R3867 VDD.n3279 VDD.n508 99.5127
R3868 VDD.n3283 VDD.n508 99.5127
R3869 VDD.n3283 VDD.n498 99.5127
R3870 VDD.n3291 VDD.n498 99.5127
R3871 VDD.n3291 VDD.n496 99.5127
R3872 VDD.n3295 VDD.n496 99.5127
R3873 VDD.n3295 VDD.n486 99.5127
R3874 VDD.n3303 VDD.n486 99.5127
R3875 VDD.n3303 VDD.n484 99.5127
R3876 VDD.n3307 VDD.n484 99.5127
R3877 VDD.n3307 VDD.n474 99.5127
R3878 VDD.n3315 VDD.n474 99.5127
R3879 VDD.n3315 VDD.n472 99.5127
R3880 VDD.n3319 VDD.n472 99.5127
R3881 VDD.n3319 VDD.n462 99.5127
R3882 VDD.n3327 VDD.n462 99.5127
R3883 VDD.n3327 VDD.n459 99.5127
R3884 VDD.n3333 VDD.n459 99.5127
R3885 VDD.n3333 VDD.n460 99.5127
R3886 VDD.n460 VDD.n452 99.5127
R3887 VDD.n452 VDD.n424 99.5127
R3888 VDD.n3398 VDD.n424 99.5127
R3889 VDD.n3398 VDD.n425 99.5127
R3890 VDD.n425 VDD.n416 99.5127
R3891 VDD.n3393 VDD.n416 99.5127
R3892 VDD.n2698 VDD.n734 99.5127
R3893 VDD.n2694 VDD.n2693 99.5127
R3894 VDD.n2690 VDD.n2689 99.5127
R3895 VDD.n2686 VDD.n2685 99.5127
R3896 VDD.n2682 VDD.n2681 99.5127
R3897 VDD.n2678 VDD.n2677 99.5127
R3898 VDD.n2674 VDD.n2673 99.5127
R3899 VDD.n2670 VDD.n2669 99.5127
R3900 VDD.n2666 VDD.n2665 99.5127
R3901 VDD.n2662 VDD.n2661 99.5127
R3902 VDD.n2658 VDD.n2657 99.5127
R3903 VDD.n2654 VDD.n732 99.5127
R3904 VDD.n2054 VDD.n1016 99.5127
R3905 VDD.n2051 VDD.n1016 99.5127
R3906 VDD.n2051 VDD.n1010 99.5127
R3907 VDD.n2048 VDD.n1010 99.5127
R3908 VDD.n2048 VDD.n1003 99.5127
R3909 VDD.n2045 VDD.n1003 99.5127
R3910 VDD.n2045 VDD.n996 99.5127
R3911 VDD.n2042 VDD.n996 99.5127
R3912 VDD.n2042 VDD.n991 99.5127
R3913 VDD.n2039 VDD.n991 99.5127
R3914 VDD.n2039 VDD.n986 99.5127
R3915 VDD.n2036 VDD.n986 99.5127
R3916 VDD.n2036 VDD.n980 99.5127
R3917 VDD.n2033 VDD.n980 99.5127
R3918 VDD.n2033 VDD.n974 99.5127
R3919 VDD.n2030 VDD.n974 99.5127
R3920 VDD.n2030 VDD.n968 99.5127
R3921 VDD.n2027 VDD.n968 99.5127
R3922 VDD.n2027 VDD.n961 99.5127
R3923 VDD.n2024 VDD.n961 99.5127
R3924 VDD.n2024 VDD.n955 99.5127
R3925 VDD.n2021 VDD.n955 99.5127
R3926 VDD.n2021 VDD.n950 99.5127
R3927 VDD.n2018 VDD.n950 99.5127
R3928 VDD.n2018 VDD.n944 99.5127
R3929 VDD.n2015 VDD.n944 99.5127
R3930 VDD.n2015 VDD.n938 99.5127
R3931 VDD.n2012 VDD.n938 99.5127
R3932 VDD.n2012 VDD.n932 99.5127
R3933 VDD.n2009 VDD.n932 99.5127
R3934 VDD.n2009 VDD.n925 99.5127
R3935 VDD.n2006 VDD.n925 99.5127
R3936 VDD.n2006 VDD.n919 99.5127
R3937 VDD.n2003 VDD.n919 99.5127
R3938 VDD.n2003 VDD.n914 99.5127
R3939 VDD.n2000 VDD.n914 99.5127
R3940 VDD.n2000 VDD.n908 99.5127
R3941 VDD.n1997 VDD.n908 99.5127
R3942 VDD.n1997 VDD.n902 99.5127
R3943 VDD.n1994 VDD.n902 99.5127
R3944 VDD.n1994 VDD.n895 99.5127
R3945 VDD.n895 VDD.n886 99.5127
R3946 VDD.n2331 VDD.n886 99.5127
R3947 VDD.n2332 VDD.n2331 99.5127
R3948 VDD.n2332 VDD.n879 99.5127
R3949 VDD.n2335 VDD.n879 99.5127
R3950 VDD.n2335 VDD.n873 99.5127
R3951 VDD.n2338 VDD.n873 99.5127
R3952 VDD.n2338 VDD.n867 99.5127
R3953 VDD.n2341 VDD.n867 99.5127
R3954 VDD.n2341 VDD.n861 99.5127
R3955 VDD.n2344 VDD.n861 99.5127
R3956 VDD.n2344 VDD.n855 99.5127
R3957 VDD.n2347 VDD.n855 99.5127
R3958 VDD.n2347 VDD.n848 99.5127
R3959 VDD.n2350 VDD.n848 99.5127
R3960 VDD.n2350 VDD.n842 99.5127
R3961 VDD.n2353 VDD.n842 99.5127
R3962 VDD.n2353 VDD.n837 99.5127
R3963 VDD.n2356 VDD.n837 99.5127
R3964 VDD.n2356 VDD.n831 99.5127
R3965 VDD.n2359 VDD.n831 99.5127
R3966 VDD.n2359 VDD.n825 99.5127
R3967 VDD.n2362 VDD.n825 99.5127
R3968 VDD.n2362 VDD.n819 99.5127
R3969 VDD.n2365 VDD.n819 99.5127
R3970 VDD.n2365 VDD.n812 99.5127
R3971 VDD.n2368 VDD.n812 99.5127
R3972 VDD.n2368 VDD.n806 99.5127
R3973 VDD.n2371 VDD.n806 99.5127
R3974 VDD.n2371 VDD.n801 99.5127
R3975 VDD.n2374 VDD.n801 99.5127
R3976 VDD.n2374 VDD.n795 99.5127
R3977 VDD.n2377 VDD.n795 99.5127
R3978 VDD.n2377 VDD.n789 99.5127
R3979 VDD.n2380 VDD.n789 99.5127
R3980 VDD.n2380 VDD.n783 99.5127
R3981 VDD.n2383 VDD.n783 99.5127
R3982 VDD.n2383 VDD.n777 99.5127
R3983 VDD.n2386 VDD.n777 99.5127
R3984 VDD.n2386 VDD.n771 99.5127
R3985 VDD.n2389 VDD.n771 99.5127
R3986 VDD.n2389 VDD.n765 99.5127
R3987 VDD.n2398 VDD.n765 99.5127
R3988 VDD.n2398 VDD.n758 99.5127
R3989 VDD.n2394 VDD.n758 99.5127
R3990 VDD.n2394 VDD.n752 99.5127
R3991 VDD.n752 VDD.n740 99.5127
R3992 VDD.n2650 VDD.n740 99.5127
R3993 VDD.n2651 VDD.n2650 99.5127
R3994 VDD.n2194 VDD.n1019 99.5127
R3995 VDD.n1971 VDD.n1970 99.5127
R3996 VDD.n1975 VDD.n1974 99.5127
R3997 VDD.n1979 VDD.n1978 99.5127
R3998 VDD.n1983 VDD.n1982 99.5127
R3999 VDD.n1987 VDD.n1986 99.5127
R4000 VDD.n2077 VDD.n2076 99.5127
R4001 VDD.n2073 VDD.n2072 99.5127
R4002 VDD.n2069 VDD.n2068 99.5127
R4003 VDD.n2065 VDD.n2064 99.5127
R4004 VDD.n2061 VDD.n2060 99.5127
R4005 VDD.n2057 VDD.n1042 99.5127
R4006 VDD.n2198 VDD.n1017 99.5127
R4007 VDD.n2198 VDD.n1007 99.5127
R4008 VDD.n2206 VDD.n1007 99.5127
R4009 VDD.n2206 VDD.n1005 99.5127
R4010 VDD.n2210 VDD.n1005 99.5127
R4011 VDD.n2210 VDD.n994 99.5127
R4012 VDD.n2218 VDD.n994 99.5127
R4013 VDD.n2218 VDD.n992 99.5127
R4014 VDD.n2222 VDD.n992 99.5127
R4015 VDD.n2222 VDD.n983 99.5127
R4016 VDD.n2230 VDD.n983 99.5127
R4017 VDD.n2230 VDD.n981 99.5127
R4018 VDD.n2234 VDD.n981 99.5127
R4019 VDD.n2234 VDD.n971 99.5127
R4020 VDD.n2242 VDD.n971 99.5127
R4021 VDD.n2242 VDD.n969 99.5127
R4022 VDD.n2246 VDD.n969 99.5127
R4023 VDD.n2246 VDD.n958 99.5127
R4024 VDD.n2254 VDD.n958 99.5127
R4025 VDD.n2254 VDD.n956 99.5127
R4026 VDD.n2258 VDD.n956 99.5127
R4027 VDD.n2258 VDD.n947 99.5127
R4028 VDD.n2266 VDD.n947 99.5127
R4029 VDD.n2266 VDD.n945 99.5127
R4030 VDD.n2270 VDD.n945 99.5127
R4031 VDD.n2270 VDD.n935 99.5127
R4032 VDD.n2278 VDD.n935 99.5127
R4033 VDD.n2278 VDD.n933 99.5127
R4034 VDD.n2282 VDD.n933 99.5127
R4035 VDD.n2282 VDD.n922 99.5127
R4036 VDD.n2290 VDD.n922 99.5127
R4037 VDD.n2290 VDD.n920 99.5127
R4038 VDD.n2294 VDD.n920 99.5127
R4039 VDD.n2294 VDD.n911 99.5127
R4040 VDD.n2302 VDD.n911 99.5127
R4041 VDD.n2302 VDD.n909 99.5127
R4042 VDD.n2306 VDD.n909 99.5127
R4043 VDD.n2306 VDD.n899 99.5127
R4044 VDD.n2314 VDD.n899 99.5127
R4045 VDD.n2314 VDD.n896 99.5127
R4046 VDD.n2323 VDD.n896 99.5127
R4047 VDD.n2323 VDD.n897 99.5127
R4048 VDD.n897 VDD.n889 99.5127
R4049 VDD.n2318 VDD.n889 99.5127
R4050 VDD.n2318 VDD.n878 99.5127
R4051 VDD.n878 VDD.n870 99.5127
R4052 VDD.n2466 VDD.n870 99.5127
R4053 VDD.n2466 VDD.n868 99.5127
R4054 VDD.n2470 VDD.n868 99.5127
R4055 VDD.n2470 VDD.n858 99.5127
R4056 VDD.n2478 VDD.n858 99.5127
R4057 VDD.n2478 VDD.n856 99.5127
R4058 VDD.n2482 VDD.n856 99.5127
R4059 VDD.n2482 VDD.n845 99.5127
R4060 VDD.n2490 VDD.n845 99.5127
R4061 VDD.n2490 VDD.n843 99.5127
R4062 VDD.n2494 VDD.n843 99.5127
R4063 VDD.n2494 VDD.n834 99.5127
R4064 VDD.n2502 VDD.n834 99.5127
R4065 VDD.n2502 VDD.n832 99.5127
R4066 VDD.n2506 VDD.n832 99.5127
R4067 VDD.n2506 VDD.n822 99.5127
R4068 VDD.n2514 VDD.n822 99.5127
R4069 VDD.n2514 VDD.n820 99.5127
R4070 VDD.n2518 VDD.n820 99.5127
R4071 VDD.n2518 VDD.n809 99.5127
R4072 VDD.n2526 VDD.n809 99.5127
R4073 VDD.n2526 VDD.n807 99.5127
R4074 VDD.n2530 VDD.n807 99.5127
R4075 VDD.n2530 VDD.n798 99.5127
R4076 VDD.n2538 VDD.n798 99.5127
R4077 VDD.n2538 VDD.n796 99.5127
R4078 VDD.n2542 VDD.n796 99.5127
R4079 VDD.n2542 VDD.n786 99.5127
R4080 VDD.n2550 VDD.n786 99.5127
R4081 VDD.n2550 VDD.n784 99.5127
R4082 VDD.n2554 VDD.n784 99.5127
R4083 VDD.n2554 VDD.n774 99.5127
R4084 VDD.n2562 VDD.n774 99.5127
R4085 VDD.n2562 VDD.n772 99.5127
R4086 VDD.n2566 VDD.n772 99.5127
R4087 VDD.n2566 VDD.n762 99.5127
R4088 VDD.n2574 VDD.n762 99.5127
R4089 VDD.n2574 VDD.n759 99.5127
R4090 VDD.n2583 VDD.n759 99.5127
R4091 VDD.n2583 VDD.n760 99.5127
R4092 VDD.n760 VDD.n753 99.5127
R4093 VDD.n2578 VDD.n753 99.5127
R4094 VDD.n2578 VDD.n743 99.5127
R4095 VDD.n743 VDD.n733 99.5127
R4096 VDD.n1448 VDD.n1447 77.1884
R4097 VDD.n1539 VDD.n1538 77.1884
R4098 VDD.n1493 VDD.n1492 77.1884
R4099 VDD.n1574 VDD.n1573 77.1884
R4100 VDD.n2083 VDD.n2082 77.1884
R4101 VDD.n2106 VDD.n2105 77.1884
R4102 VDD.n2129 VDD.n2128 77.1884
R4103 VDD.n1169 VDD.n1168 77.1884
R4104 VDD.n3842 VDD.n3841 77.1884
R4105 VDD.n220 VDD.n219 77.1884
R4106 VDD.n3880 VDD.n3879 77.1884
R4107 VDD.n180 VDD.n179 77.1884
R4108 VDD.n3473 VDD.n3472 77.1884
R4109 VDD.n3490 VDD.n3489 77.1884
R4110 VDD.n3508 VDD.n3507 77.1884
R4111 VDD.n3524 VDD.n3523 77.1884
R4112 VDD.n1990 VDD.n1989 76.9944
R4113 VDD.n737 VDD.n736 76.9944
R4114 VDD.n1046 VDD.n1045 76.9944
R4115 VDD.n748 VDD.n747 76.9944
R4116 VDD.n2849 VDD.n2848 76.9944
R4117 VDD.n407 VDD.n406 76.9944
R4118 VDD.n2725 VDD.n2724 76.9944
R4119 VDD.n446 VDD.n445 76.9944
R4120 VDD.n3080 VDD.n2722 72.8958
R4121 VDD.n3080 VDD.n2721 72.8958
R4122 VDD.n3080 VDD.n2720 72.8958
R4123 VDD.n3080 VDD.n2719 72.8958
R4124 VDD.n3080 VDD.n2718 72.8958
R4125 VDD.n3080 VDD.n2717 72.8958
R4126 VDD.n3080 VDD.n2716 72.8958
R4127 VDD.n3080 VDD.n2715 72.8958
R4128 VDD.n3080 VDD.n2714 72.8958
R4129 VDD.n3080 VDD.n2713 72.8958
R4130 VDD.n3080 VDD.n2712 72.8958
R4131 VDD.n3080 VDD.n2711 72.8958
R4132 VDD.n3349 VDD.n400 72.8958
R4133 VDD.n3356 VDD.n400 72.8958
R4134 VDD.n443 VDD.n400 72.8958
R4135 VDD.n3363 VDD.n400 72.8958
R4136 VDD.n440 VDD.n400 72.8958
R4137 VDD.n3370 VDD.n400 72.8958
R4138 VDD.n436 VDD.n400 72.8958
R4139 VDD.n3377 VDD.n400 72.8958
R4140 VDD.n433 VDD.n400 72.8958
R4141 VDD.n3384 VDD.n400 72.8958
R4142 VDD.n430 VDD.n400 72.8958
R4143 VDD.n3391 VDD.n400 72.8958
R4144 VDD.n2193 VDD.n2192 72.8958
R4145 VDD.n2193 VDD.n1020 72.8958
R4146 VDD.n2193 VDD.n1021 72.8958
R4147 VDD.n2193 VDD.n1022 72.8958
R4148 VDD.n2193 VDD.n1023 72.8958
R4149 VDD.n2193 VDD.n1024 72.8958
R4150 VDD.n2193 VDD.n1025 72.8958
R4151 VDD.n2193 VDD.n1026 72.8958
R4152 VDD.n2193 VDD.n1027 72.8958
R4153 VDD.n2193 VDD.n1028 72.8958
R4154 VDD.n2193 VDD.n1029 72.8958
R4155 VDD.n2699 VDD.n720 72.8958
R4156 VDD.n2699 VDD.n719 72.8958
R4157 VDD.n2699 VDD.n718 72.8958
R4158 VDD.n2699 VDD.n717 72.8958
R4159 VDD.n2699 VDD.n716 72.8958
R4160 VDD.n2699 VDD.n715 72.8958
R4161 VDD.n2699 VDD.n714 72.8958
R4162 VDD.n2699 VDD.n713 72.8958
R4163 VDD.n2699 VDD.n712 72.8958
R4164 VDD.n2699 VDD.n711 72.8958
R4165 VDD.n2699 VDD.n710 72.8958
R4166 VDD.n2699 VDD.n709 72.8958
R4167 VDD.n3081 VDD.n3080 72.8958
R4168 VDD.n3080 VDD.n2700 72.8958
R4169 VDD.n3080 VDD.n2701 72.8958
R4170 VDD.n3080 VDD.n2702 72.8958
R4171 VDD.n3080 VDD.n2703 72.8958
R4172 VDD.n3080 VDD.n2704 72.8958
R4173 VDD.n3080 VDD.n2705 72.8958
R4174 VDD.n3080 VDD.n2706 72.8958
R4175 VDD.n3080 VDD.n2707 72.8958
R4176 VDD.n3080 VDD.n2708 72.8958
R4177 VDD.n3080 VDD.n2709 72.8958
R4178 VDD.n3440 VDD.n400 72.8958
R4179 VDD.n409 VDD.n400 72.8958
R4180 VDD.n3448 VDD.n400 72.8958
R4181 VDD.n404 VDD.n400 72.8958
R4182 VDD.n3455 VDD.n400 72.8958
R4183 VDD.n3458 VDD.n400 72.8958
R4184 VDD.n3411 VDD.n400 72.8958
R4185 VDD.n3410 VDD.n400 72.8958
R4186 VDD.n3418 VDD.n400 72.8958
R4187 VDD.n3407 VDD.n400 72.8958
R4188 VDD.n3425 VDD.n400 72.8958
R4189 VDD.n3428 VDD.n400 72.8958
R4190 VDD.n2699 VDD.n731 72.8958
R4191 VDD.n2699 VDD.n730 72.8958
R4192 VDD.n2699 VDD.n729 72.8958
R4193 VDD.n2699 VDD.n728 72.8958
R4194 VDD.n2699 VDD.n727 72.8958
R4195 VDD.n2699 VDD.n726 72.8958
R4196 VDD.n2699 VDD.n725 72.8958
R4197 VDD.n2699 VDD.n724 72.8958
R4198 VDD.n2699 VDD.n723 72.8958
R4199 VDD.n2699 VDD.n722 72.8958
R4200 VDD.n2699 VDD.n721 72.8958
R4201 VDD.n2193 VDD.n1031 72.8958
R4202 VDD.n2193 VDD.n1032 72.8958
R4203 VDD.n2193 VDD.n1033 72.8958
R4204 VDD.n2193 VDD.n1034 72.8958
R4205 VDD.n2193 VDD.n1035 72.8958
R4206 VDD.n2193 VDD.n1036 72.8958
R4207 VDD.n2193 VDD.n1037 72.8958
R4208 VDD.n2193 VDD.n1038 72.8958
R4209 VDD.n2193 VDD.n1039 72.8958
R4210 VDD.n2193 VDD.n1040 72.8958
R4211 VDD.n2193 VDD.n1041 72.8958
R4212 VDD.n1589 VDD.n1588 66.2847
R4213 VDD.n1589 VDD.n1451 66.2847
R4214 VDD.n1589 VDD.n1452 66.2847
R4215 VDD.n1589 VDD.n1453 66.2847
R4216 VDD.n1589 VDD.n1454 66.2847
R4217 VDD.n1589 VDD.n1455 66.2847
R4218 VDD.n1589 VDD.n1456 66.2847
R4219 VDD.n1589 VDD.n1457 66.2847
R4220 VDD.n1589 VDD.n1458 66.2847
R4221 VDD.n1589 VDD.n1459 66.2847
R4222 VDD.n1589 VDD.n1460 66.2847
R4223 VDD.n1589 VDD.n1461 66.2847
R4224 VDD.n1589 VDD.n1462 66.2847
R4225 VDD.n1589 VDD.n1463 66.2847
R4226 VDD.n1589 VDD.n1464 66.2847
R4227 VDD.n1589 VDD.n1465 66.2847
R4228 VDD.n1589 VDD.n1466 66.2847
R4229 VDD.n1589 VDD.n1467 66.2847
R4230 VDD.n1590 VDD.n1589 66.2847
R4231 VDD.n2165 VDD.n1143 66.2847
R4232 VDD.n2165 VDD.n1144 66.2847
R4233 VDD.n2165 VDD.n1145 66.2847
R4234 VDD.n2165 VDD.n1146 66.2847
R4235 VDD.n2165 VDD.n1147 66.2847
R4236 VDD.n2165 VDD.n1148 66.2847
R4237 VDD.n2165 VDD.n1149 66.2847
R4238 VDD.n2165 VDD.n1150 66.2847
R4239 VDD.n2165 VDD.n1151 66.2847
R4240 VDD.n2165 VDD.n1152 66.2847
R4241 VDD.n2165 VDD.n1153 66.2847
R4242 VDD.n2165 VDD.n1154 66.2847
R4243 VDD.n2165 VDD.n1155 66.2847
R4244 VDD.n2165 VDD.n1156 66.2847
R4245 VDD.n2165 VDD.n1157 66.2847
R4246 VDD.n2165 VDD.n1158 66.2847
R4247 VDD.n2165 VDD.n1159 66.2847
R4248 VDD.n2165 VDD.n1160 66.2847
R4249 VDD.n2165 VDD.n2164 66.2847
R4250 VDD.n3600 VDD.n394 66.2847
R4251 VDD.n3463 VDD.n394 66.2847
R4252 VDD.n3593 VDD.n394 66.2847
R4253 VDD.n3587 VDD.n394 66.2847
R4254 VDD.n3585 VDD.n394 66.2847
R4255 VDD.n3579 VDD.n394 66.2847
R4256 VDD.n3577 VDD.n394 66.2847
R4257 VDD.n3571 VDD.n394 66.2847
R4258 VDD.n3569 VDD.n394 66.2847
R4259 VDD.n3563 VDD.n394 66.2847
R4260 VDD.n3561 VDD.n394 66.2847
R4261 VDD.n3555 VDD.n394 66.2847
R4262 VDD.n3553 VDD.n394 66.2847
R4263 VDD.n3546 VDD.n394 66.2847
R4264 VDD.n3544 VDD.n394 66.2847
R4265 VDD.n3538 VDD.n394 66.2847
R4266 VDD.n3536 VDD.n394 66.2847
R4267 VDD.n3530 VDD.n394 66.2847
R4268 VDD.n3528 VDD.n394 66.2847
R4269 VDD.n3838 VDD.n166 66.2847
R4270 VDD.n3847 VDD.n166 66.2847
R4271 VDD.n234 VDD.n166 66.2847
R4272 VDD.n3854 VDD.n166 66.2847
R4273 VDD.n227 VDD.n166 66.2847
R4274 VDD.n3861 VDD.n166 66.2847
R4275 VDD.n217 VDD.n166 66.2847
R4276 VDD.n3868 VDD.n166 66.2847
R4277 VDD.n210 VDD.n166 66.2847
R4278 VDD.n3875 VDD.n166 66.2847
R4279 VDD.n203 VDD.n166 66.2847
R4280 VDD.n3885 VDD.n166 66.2847
R4281 VDD.n196 VDD.n166 66.2847
R4282 VDD.n3892 VDD.n166 66.2847
R4283 VDD.n189 VDD.n166 66.2847
R4284 VDD.n3899 VDD.n166 66.2847
R4285 VDD.n182 VDD.n166 66.2847
R4286 VDD.n3906 VDD.n166 66.2847
R4287 VDD.n173 VDD.n166 66.2847
R4288 VDD.n3908 VDD.n173 52.4337
R4289 VDD.n3906 VDD.n3905 52.4337
R4290 VDD.n3901 VDD.n182 52.4337
R4291 VDD.n3899 VDD.n3898 52.4337
R4292 VDD.n3894 VDD.n189 52.4337
R4293 VDD.n3892 VDD.n3891 52.4337
R4294 VDD.n3887 VDD.n196 52.4337
R4295 VDD.n3885 VDD.n3884 52.4337
R4296 VDD.n3877 VDD.n203 52.4337
R4297 VDD.n3875 VDD.n3874 52.4337
R4298 VDD.n3870 VDD.n210 52.4337
R4299 VDD.n3868 VDD.n3867 52.4337
R4300 VDD.n3863 VDD.n217 52.4337
R4301 VDD.n3861 VDD.n3860 52.4337
R4302 VDD.n3856 VDD.n227 52.4337
R4303 VDD.n3854 VDD.n3853 52.4337
R4304 VDD.n3849 VDD.n234 52.4337
R4305 VDD.n3847 VDD.n3846 52.4337
R4306 VDD.n3839 VDD.n3838 52.4337
R4307 VDD.n3600 VDD.n395 52.4337
R4308 VDD.n3598 VDD.n3463 52.4337
R4309 VDD.n3594 VDD.n3593 52.4337
R4310 VDD.n3587 VDD.n3468 52.4337
R4311 VDD.n3586 VDD.n3585 52.4337
R4312 VDD.n3579 VDD.n3476 52.4337
R4313 VDD.n3578 VDD.n3577 52.4337
R4314 VDD.n3571 VDD.n3482 52.4337
R4315 VDD.n3570 VDD.n3569 52.4337
R4316 VDD.n3563 VDD.n3488 52.4337
R4317 VDD.n3562 VDD.n3561 52.4337
R4318 VDD.n3555 VDD.n3497 52.4337
R4319 VDD.n3554 VDD.n3553 52.4337
R4320 VDD.n3546 VDD.n3503 52.4337
R4321 VDD.n3545 VDD.n3544 52.4337
R4322 VDD.n3538 VDD.n3511 52.4337
R4323 VDD.n3537 VDD.n3536 52.4337
R4324 VDD.n3530 VDD.n3517 52.4337
R4325 VDD.n3529 VDD.n3528 52.4337
R4326 VDD.n2164 VDD.n2163 52.4337
R4327 VDD.n2159 VDD.n1160 52.4337
R4328 VDD.n2155 VDD.n1159 52.4337
R4329 VDD.n2147 VDD.n1158 52.4337
R4330 VDD.n2145 VDD.n1157 52.4337
R4331 VDD.n2141 VDD.n1156 52.4337
R4332 VDD.n2137 VDD.n1155 52.4337
R4333 VDD.n2133 VDD.n1154 52.4337
R4334 VDD.n2126 VDD.n1153 52.4337
R4335 VDD.n2122 VDD.n1152 52.4337
R4336 VDD.n2118 VDD.n1151 52.4337
R4337 VDD.n2114 VDD.n1150 52.4337
R4338 VDD.n2110 VDD.n1149 52.4337
R4339 VDD.n2103 VDD.n1148 52.4337
R4340 VDD.n2099 VDD.n1147 52.4337
R4341 VDD.n2095 VDD.n1146 52.4337
R4342 VDD.n2091 VDD.n1145 52.4337
R4343 VDD.n2087 VDD.n1144 52.4337
R4344 VDD.n1198 VDD.n1143 52.4337
R4345 VDD.n1588 VDD.n1587 52.4337
R4346 VDD.n1473 VDD.n1451 52.4337
R4347 VDD.n1475 VDD.n1452 52.4337
R4348 VDD.n1572 VDD.n1453 52.4337
R4349 VDD.n1479 VDD.n1454 52.4337
R4350 VDD.n1483 VDD.n1455 52.4337
R4351 VDD.n1485 VDD.n1456 52.4337
R4352 VDD.n1489 VDD.n1457 52.4337
R4353 VDD.n1491 VDD.n1458 52.4337
R4354 VDD.n1497 VDD.n1459 52.4337
R4355 VDD.n1499 VDD.n1460 52.4337
R4356 VDD.n1503 VDD.n1461 52.4337
R4357 VDD.n1505 VDD.n1462 52.4337
R4358 VDD.n1509 VDD.n1463 52.4337
R4359 VDD.n1511 VDD.n1464 52.4337
R4360 VDD.n1515 VDD.n1465 52.4337
R4361 VDD.n1517 VDD.n1466 52.4337
R4362 VDD.n1521 VDD.n1467 52.4337
R4363 VDD.n1590 VDD.n1450 52.4337
R4364 VDD.n1588 VDD.n1469 52.4337
R4365 VDD.n1474 VDD.n1451 52.4337
R4366 VDD.n1571 VDD.n1452 52.4337
R4367 VDD.n1478 VDD.n1453 52.4337
R4368 VDD.n1482 VDD.n1454 52.4337
R4369 VDD.n1484 VDD.n1455 52.4337
R4370 VDD.n1488 VDD.n1456 52.4337
R4371 VDD.n1490 VDD.n1457 52.4337
R4372 VDD.n1496 VDD.n1458 52.4337
R4373 VDD.n1498 VDD.n1459 52.4337
R4374 VDD.n1502 VDD.n1460 52.4337
R4375 VDD.n1504 VDD.n1461 52.4337
R4376 VDD.n1508 VDD.n1462 52.4337
R4377 VDD.n1510 VDD.n1463 52.4337
R4378 VDD.n1514 VDD.n1464 52.4337
R4379 VDD.n1516 VDD.n1465 52.4337
R4380 VDD.n1520 VDD.n1466 52.4337
R4381 VDD.n1522 VDD.n1467 52.4337
R4382 VDD.n1591 VDD.n1590 52.4337
R4383 VDD.n2086 VDD.n1143 52.4337
R4384 VDD.n2090 VDD.n1144 52.4337
R4385 VDD.n2094 VDD.n1145 52.4337
R4386 VDD.n2098 VDD.n1146 52.4337
R4387 VDD.n2102 VDD.n1147 52.4337
R4388 VDD.n2109 VDD.n1148 52.4337
R4389 VDD.n2113 VDD.n1149 52.4337
R4390 VDD.n2117 VDD.n1150 52.4337
R4391 VDD.n2121 VDD.n1151 52.4337
R4392 VDD.n2125 VDD.n1152 52.4337
R4393 VDD.n2132 VDD.n1153 52.4337
R4394 VDD.n2136 VDD.n1154 52.4337
R4395 VDD.n2140 VDD.n1155 52.4337
R4396 VDD.n2144 VDD.n1156 52.4337
R4397 VDD.n2148 VDD.n1157 52.4337
R4398 VDD.n2154 VDD.n1158 52.4337
R4399 VDD.n2158 VDD.n1159 52.4337
R4400 VDD.n1161 VDD.n1160 52.4337
R4401 VDD.n2164 VDD.n1141 52.4337
R4402 VDD.n3601 VDD.n3600 52.4337
R4403 VDD.n3595 VDD.n3463 52.4337
R4404 VDD.n3593 VDD.n3592 52.4337
R4405 VDD.n3588 VDD.n3587 52.4337
R4406 VDD.n3585 VDD.n3584 52.4337
R4407 VDD.n3580 VDD.n3579 52.4337
R4408 VDD.n3577 VDD.n3576 52.4337
R4409 VDD.n3572 VDD.n3571 52.4337
R4410 VDD.n3569 VDD.n3568 52.4337
R4411 VDD.n3564 VDD.n3563 52.4337
R4412 VDD.n3561 VDD.n3560 52.4337
R4413 VDD.n3556 VDD.n3555 52.4337
R4414 VDD.n3553 VDD.n3552 52.4337
R4415 VDD.n3547 VDD.n3546 52.4337
R4416 VDD.n3544 VDD.n3543 52.4337
R4417 VDD.n3539 VDD.n3538 52.4337
R4418 VDD.n3536 VDD.n3535 52.4337
R4419 VDD.n3531 VDD.n3530 52.4337
R4420 VDD.n3528 VDD.n393 52.4337
R4421 VDD.n3838 VDD.n235 52.4337
R4422 VDD.n3848 VDD.n3847 52.4337
R4423 VDD.n234 VDD.n228 52.4337
R4424 VDD.n3855 VDD.n3854 52.4337
R4425 VDD.n227 VDD.n218 52.4337
R4426 VDD.n3862 VDD.n3861 52.4337
R4427 VDD.n217 VDD.n211 52.4337
R4428 VDD.n3869 VDD.n3868 52.4337
R4429 VDD.n210 VDD.n204 52.4337
R4430 VDD.n3876 VDD.n3875 52.4337
R4431 VDD.n203 VDD.n197 52.4337
R4432 VDD.n3886 VDD.n3885 52.4337
R4433 VDD.n196 VDD.n190 52.4337
R4434 VDD.n3893 VDD.n3892 52.4337
R4435 VDD.n189 VDD.n183 52.4337
R4436 VDD.n3900 VDD.n3899 52.4337
R4437 VDD.n182 VDD.n174 52.4337
R4438 VDD.n3907 VDD.n3906 52.4337
R4439 VDD.n173 VDD.n170 52.4337
R4440 VDD.n3428 VDD.n3427 39.2114
R4441 VDD.n3425 VDD.n3424 39.2114
R4442 VDD.n3420 VDD.n3407 39.2114
R4443 VDD.n3418 VDD.n3417 39.2114
R4444 VDD.n3413 VDD.n3410 39.2114
R4445 VDD.n3411 VDD.n399 39.2114
R4446 VDD.n3458 VDD.n3457 39.2114
R4447 VDD.n3455 VDD.n3454 39.2114
R4448 VDD.n3450 VDD.n404 39.2114
R4449 VDD.n3448 VDD.n3447 39.2114
R4450 VDD.n3442 VDD.n409 39.2114
R4451 VDD.n3440 VDD.n3439 39.2114
R4452 VDD.n3082 VDD.n3081 39.2114
R4453 VDD.n2723 VDD.n2700 39.2114
R4454 VDD.n3074 VDD.n2701 39.2114
R4455 VDD.n3070 VDD.n2702 39.2114
R4456 VDD.n3066 VDD.n2703 39.2114
R4457 VDD.n3062 VDD.n2704 39.2114
R4458 VDD.n3058 VDD.n2705 39.2114
R4459 VDD.n3054 VDD.n2706 39.2114
R4460 VDD.n3050 VDD.n2707 39.2114
R4461 VDD.n3046 VDD.n2708 39.2114
R4462 VDD.n3042 VDD.n2709 39.2114
R4463 VDD.n2642 VDD.n709 39.2114
R4464 VDD.n2638 VDD.n710 39.2114
R4465 VDD.n2634 VDD.n711 39.2114
R4466 VDD.n2630 VDD.n712 39.2114
R4467 VDD.n2626 VDD.n713 39.2114
R4468 VDD.n2622 VDD.n714 39.2114
R4469 VDD.n2618 VDD.n715 39.2114
R4470 VDD.n2614 VDD.n716 39.2114
R4471 VDD.n2610 VDD.n717 39.2114
R4472 VDD.n2606 VDD.n718 39.2114
R4473 VDD.n2601 VDD.n719 39.2114
R4474 VDD.n2597 VDD.n720 39.2114
R4475 VDD.n2192 VDD.n2191 39.2114
R4476 VDD.n2186 VDD.n1020 39.2114
R4477 VDD.n2183 VDD.n1021 39.2114
R4478 VDD.n2179 VDD.n1022 39.2114
R4479 VDD.n2175 VDD.n1023 39.2114
R4480 VDD.n2171 VDD.n1024 39.2114
R4481 VDD.n1134 VDD.n1025 39.2114
R4482 VDD.n1130 VDD.n1026 39.2114
R4483 VDD.n1126 VDD.n1027 39.2114
R4484 VDD.n1122 VDD.n1028 39.2114
R4485 VDD.n1118 VDD.n1029 39.2114
R4486 VDD.n3391 VDD.n3390 39.2114
R4487 VDD.n3386 VDD.n430 39.2114
R4488 VDD.n3384 VDD.n3383 39.2114
R4489 VDD.n3379 VDD.n433 39.2114
R4490 VDD.n3377 VDD.n3376 39.2114
R4491 VDD.n3372 VDD.n436 39.2114
R4492 VDD.n3370 VDD.n3369 39.2114
R4493 VDD.n3365 VDD.n440 39.2114
R4494 VDD.n3363 VDD.n3362 39.2114
R4495 VDD.n3358 VDD.n443 39.2114
R4496 VDD.n3356 VDD.n3355 39.2114
R4497 VDD.n3351 VDD.n3349 39.2114
R4498 VDD.n2850 VDD.n2722 39.2114
R4499 VDD.n2854 VDD.n2721 39.2114
R4500 VDD.n2858 VDD.n2720 39.2114
R4501 VDD.n2862 VDD.n2719 39.2114
R4502 VDD.n2866 VDD.n2718 39.2114
R4503 VDD.n2870 VDD.n2717 39.2114
R4504 VDD.n2874 VDD.n2716 39.2114
R4505 VDD.n2878 VDD.n2715 39.2114
R4506 VDD.n2882 VDD.n2714 39.2114
R4507 VDD.n2886 VDD.n2713 39.2114
R4508 VDD.n2890 VDD.n2712 39.2114
R4509 VDD.n2895 VDD.n2711 39.2114
R4510 VDD.n2853 VDD.n2722 39.2114
R4511 VDD.n2857 VDD.n2721 39.2114
R4512 VDD.n2861 VDD.n2720 39.2114
R4513 VDD.n2865 VDD.n2719 39.2114
R4514 VDD.n2869 VDD.n2718 39.2114
R4515 VDD.n2873 VDD.n2717 39.2114
R4516 VDD.n2877 VDD.n2716 39.2114
R4517 VDD.n2881 VDD.n2715 39.2114
R4518 VDD.n2885 VDD.n2714 39.2114
R4519 VDD.n2889 VDD.n2713 39.2114
R4520 VDD.n2894 VDD.n2712 39.2114
R4521 VDD.n2898 VDD.n2711 39.2114
R4522 VDD.n3349 VDD.n444 39.2114
R4523 VDD.n3357 VDD.n3356 39.2114
R4524 VDD.n443 VDD.n441 39.2114
R4525 VDD.n3364 VDD.n3363 39.2114
R4526 VDD.n440 VDD.n438 39.2114
R4527 VDD.n3371 VDD.n3370 39.2114
R4528 VDD.n436 VDD.n434 39.2114
R4529 VDD.n3378 VDD.n3377 39.2114
R4530 VDD.n433 VDD.n431 39.2114
R4531 VDD.n3385 VDD.n3384 39.2114
R4532 VDD.n430 VDD.n428 39.2114
R4533 VDD.n3392 VDD.n3391 39.2114
R4534 VDD.n2192 VDD.n1044 39.2114
R4535 VDD.n2184 VDD.n1020 39.2114
R4536 VDD.n2180 VDD.n1021 39.2114
R4537 VDD.n2176 VDD.n1022 39.2114
R4538 VDD.n2172 VDD.n1023 39.2114
R4539 VDD.n1135 VDD.n1024 39.2114
R4540 VDD.n1131 VDD.n1025 39.2114
R4541 VDD.n1127 VDD.n1026 39.2114
R4542 VDD.n1123 VDD.n1027 39.2114
R4543 VDD.n1119 VDD.n1028 39.2114
R4544 VDD.n1115 VDD.n1029 39.2114
R4545 VDD.n2600 VDD.n720 39.2114
R4546 VDD.n2605 VDD.n719 39.2114
R4547 VDD.n2609 VDD.n718 39.2114
R4548 VDD.n2613 VDD.n717 39.2114
R4549 VDD.n2617 VDD.n716 39.2114
R4550 VDD.n2621 VDD.n715 39.2114
R4551 VDD.n2625 VDD.n714 39.2114
R4552 VDD.n2629 VDD.n713 39.2114
R4553 VDD.n2633 VDD.n712 39.2114
R4554 VDD.n2637 VDD.n711 39.2114
R4555 VDD.n2641 VDD.n710 39.2114
R4556 VDD.n2644 VDD.n709 39.2114
R4557 VDD.n3081 VDD.n707 39.2114
R4558 VDD.n3075 VDD.n2700 39.2114
R4559 VDD.n3071 VDD.n2701 39.2114
R4560 VDD.n3067 VDD.n2702 39.2114
R4561 VDD.n3063 VDD.n2703 39.2114
R4562 VDD.n3059 VDD.n2704 39.2114
R4563 VDD.n3055 VDD.n2705 39.2114
R4564 VDD.n3051 VDD.n2706 39.2114
R4565 VDD.n3047 VDD.n2707 39.2114
R4566 VDD.n3043 VDD.n2708 39.2114
R4567 VDD.n3039 VDD.n2709 39.2114
R4568 VDD.n3441 VDD.n3440 39.2114
R4569 VDD.n409 VDD.n405 39.2114
R4570 VDD.n3449 VDD.n3448 39.2114
R4571 VDD.n404 VDD.n402 39.2114
R4572 VDD.n3456 VDD.n3455 39.2114
R4573 VDD.n3459 VDD.n3458 39.2114
R4574 VDD.n3412 VDD.n3411 39.2114
R4575 VDD.n3410 VDD.n3408 39.2114
R4576 VDD.n3419 VDD.n3418 39.2114
R4577 VDD.n3407 VDD.n3405 39.2114
R4578 VDD.n3426 VDD.n3425 39.2114
R4579 VDD.n3429 VDD.n3428 39.2114
R4580 VDD.n734 VDD.n721 39.2114
R4581 VDD.n2693 VDD.n722 39.2114
R4582 VDD.n2689 VDD.n723 39.2114
R4583 VDD.n2685 VDD.n724 39.2114
R4584 VDD.n2681 VDD.n725 39.2114
R4585 VDD.n2677 VDD.n726 39.2114
R4586 VDD.n2673 VDD.n727 39.2114
R4587 VDD.n2669 VDD.n728 39.2114
R4588 VDD.n2665 VDD.n729 39.2114
R4589 VDD.n2661 VDD.n730 39.2114
R4590 VDD.n2657 VDD.n731 39.2114
R4591 VDD.n1031 VDD.n1019 39.2114
R4592 VDD.n1971 VDD.n1032 39.2114
R4593 VDD.n1975 VDD.n1033 39.2114
R4594 VDD.n1979 VDD.n1034 39.2114
R4595 VDD.n1983 VDD.n1035 39.2114
R4596 VDD.n1987 VDD.n1036 39.2114
R4597 VDD.n2076 VDD.n1037 39.2114
R4598 VDD.n2072 VDD.n1038 39.2114
R4599 VDD.n2068 VDD.n1039 39.2114
R4600 VDD.n2064 VDD.n1040 39.2114
R4601 VDD.n2060 VDD.n1041 39.2114
R4602 VDD.n2654 VDD.n731 39.2114
R4603 VDD.n2658 VDD.n730 39.2114
R4604 VDD.n2662 VDD.n729 39.2114
R4605 VDD.n2666 VDD.n728 39.2114
R4606 VDD.n2670 VDD.n727 39.2114
R4607 VDD.n2674 VDD.n726 39.2114
R4608 VDD.n2678 VDD.n725 39.2114
R4609 VDD.n2682 VDD.n724 39.2114
R4610 VDD.n2686 VDD.n723 39.2114
R4611 VDD.n2690 VDD.n722 39.2114
R4612 VDD.n2694 VDD.n721 39.2114
R4613 VDD.n1970 VDD.n1031 39.2114
R4614 VDD.n1974 VDD.n1032 39.2114
R4615 VDD.n1978 VDD.n1033 39.2114
R4616 VDD.n1982 VDD.n1034 39.2114
R4617 VDD.n1986 VDD.n1035 39.2114
R4618 VDD.n2077 VDD.n1036 39.2114
R4619 VDD.n2073 VDD.n1037 39.2114
R4620 VDD.n2069 VDD.n1038 39.2114
R4621 VDD.n2065 VDD.n1039 39.2114
R4622 VDD.n2061 VDD.n1040 39.2114
R4623 VDD.n2057 VDD.n1041 39.2114
R4624 VDD.n1449 VDD.n1448 37.2369
R4625 VDD.n1540 VDD.n1539 37.2369
R4626 VDD.n1494 VDD.n1493 37.2369
R4627 VDD.n1575 VDD.n1574 37.2369
R4628 VDD.n2084 VDD.n2083 37.2369
R4629 VDD.n2107 VDD.n2106 37.2369
R4630 VDD.n2130 VDD.n2129 37.2369
R4631 VDD.n2153 VDD.n1169 37.2369
R4632 VDD.n3843 VDD.n3842 37.2369
R4633 VDD.n221 VDD.n220 37.2369
R4634 VDD.n3881 VDD.n3880 37.2369
R4635 VDD.n181 VDD.n180 37.2369
R4636 VDD.n3590 VDD.n3473 37.2369
R4637 VDD.n3491 VDD.n3490 37.2369
R4638 VDD.n3549 VDD.n3508 37.2369
R4639 VDD.n3525 VDD.n3524 37.2369
R4640 VDD.n2190 VDD.n1012 36.5273
R4641 VDD.n2646 VDD.n2645 36.5273
R4642 VDD.n2598 VDD.n2595 36.5273
R4643 VDD.n1114 VDD.n1113 36.5273
R4644 VDD.n3038 VDD.n3037 36.5273
R4645 VDD.n3438 VDD.n3437 36.5273
R4646 VDD.n3084 VDD.n3083 36.5273
R4647 VDD.n3431 VDD.n3430 36.5273
R4648 VDD.n3394 VDD.n427 36.5273
R4649 VDD.n3352 VDD.n3348 36.5273
R4650 VDD.n2900 VDD.n2897 36.5273
R4651 VDD.n2851 VDD.n700 36.5273
R4652 VDD.n2196 VDD.n2195 36.5273
R4653 VDD.n2697 VDD.n735 36.5273
R4654 VDD.n2653 VDD.n2652 36.5273
R4655 VDD.n2056 VDD.n2055 36.5273
R4656 VDD.n1991 VDD.n1990 30.449
R4657 VDD.n738 VDD.n737 30.449
R4658 VDD.n1047 VDD.n1046 30.449
R4659 VDD.n2603 VDD.n748 30.449
R4660 VDD.n2892 VDD.n2849 30.449
R4661 VDD.n3444 VDD.n407 30.449
R4662 VDD.n2726 VDD.n2725 30.449
R4663 VDD.n447 VDD.n446 30.449
R4664 VDD.n1589 VDD.n1443 28.7425
R4665 VDD.n2165 VDD.n1142 28.7425
R4666 VDD.n3608 VDD.n394 28.7425
R4667 VDD.n3916 VDD.n166 28.7425
R4668 VDD.n2193 VDD.n1014 20.4225
R4669 VDD.n2699 VDD.n708 20.4225
R4670 VDD.n3080 VDD.n702 20.4225
R4671 VDD.n415 VDD.n400 20.4225
R4672 VDD.n1596 VDD.n1445 19.3944
R4673 VDD.n1596 VDD.n1435 19.3944
R4674 VDD.n1608 VDD.n1435 19.3944
R4675 VDD.n1608 VDD.n1433 19.3944
R4676 VDD.n1612 VDD.n1433 19.3944
R4677 VDD.n1612 VDD.n1424 19.3944
R4678 VDD.n1624 VDD.n1424 19.3944
R4679 VDD.n1624 VDD.n1422 19.3944
R4680 VDD.n1628 VDD.n1422 19.3944
R4681 VDD.n1628 VDD.n1412 19.3944
R4682 VDD.n1640 VDD.n1412 19.3944
R4683 VDD.n1640 VDD.n1410 19.3944
R4684 VDD.n1644 VDD.n1410 19.3944
R4685 VDD.n1644 VDD.n1401 19.3944
R4686 VDD.n1657 VDD.n1401 19.3944
R4687 VDD.n1657 VDD.n1399 19.3944
R4688 VDD.n1661 VDD.n1399 19.3944
R4689 VDD.n1661 VDD.n1389 19.3944
R4690 VDD.n1673 VDD.n1389 19.3944
R4691 VDD.n1673 VDD.n1387 19.3944
R4692 VDD.n1677 VDD.n1387 19.3944
R4693 VDD.n1677 VDD.n1378 19.3944
R4694 VDD.n1690 VDD.n1378 19.3944
R4695 VDD.n1690 VDD.n1376 19.3944
R4696 VDD.n1694 VDD.n1376 19.3944
R4697 VDD.n1694 VDD.n1366 19.3944
R4698 VDD.n1706 VDD.n1366 19.3944
R4699 VDD.n1706 VDD.n1364 19.3944
R4700 VDD.n1710 VDD.n1364 19.3944
R4701 VDD.n1710 VDD.n1355 19.3944
R4702 VDD.n1723 VDD.n1355 19.3944
R4703 VDD.n1723 VDD.n1353 19.3944
R4704 VDD.n1727 VDD.n1353 19.3944
R4705 VDD.n1727 VDD.n1343 19.3944
R4706 VDD.n1739 VDD.n1343 19.3944
R4707 VDD.n1739 VDD.n1341 19.3944
R4708 VDD.n1743 VDD.n1341 19.3944
R4709 VDD.n1743 VDD.n1332 19.3944
R4710 VDD.n1756 VDD.n1332 19.3944
R4711 VDD.n1756 VDD.n1330 19.3944
R4712 VDD.n1760 VDD.n1330 19.3944
R4713 VDD.n1760 VDD.n1320 19.3944
R4714 VDD.n1804 VDD.n1320 19.3944
R4715 VDD.n1804 VDD.n1318 19.3944
R4716 VDD.n1808 VDD.n1318 19.3944
R4717 VDD.n1808 VDD.n1308 19.3944
R4718 VDD.n1820 VDD.n1308 19.3944
R4719 VDD.n1820 VDD.n1306 19.3944
R4720 VDD.n1824 VDD.n1306 19.3944
R4721 VDD.n1824 VDD.n1296 19.3944
R4722 VDD.n1836 VDD.n1296 19.3944
R4723 VDD.n1836 VDD.n1294 19.3944
R4724 VDD.n1840 VDD.n1294 19.3944
R4725 VDD.n1840 VDD.n1284 19.3944
R4726 VDD.n1852 VDD.n1284 19.3944
R4727 VDD.n1852 VDD.n1282 19.3944
R4728 VDD.n1856 VDD.n1282 19.3944
R4729 VDD.n1856 VDD.n1272 19.3944
R4730 VDD.n1868 VDD.n1272 19.3944
R4731 VDD.n1868 VDD.n1270 19.3944
R4732 VDD.n1872 VDD.n1270 19.3944
R4733 VDD.n1872 VDD.n1260 19.3944
R4734 VDD.n1884 VDD.n1260 19.3944
R4735 VDD.n1884 VDD.n1258 19.3944
R4736 VDD.n1888 VDD.n1258 19.3944
R4737 VDD.n1888 VDD.n1248 19.3944
R4738 VDD.n1900 VDD.n1248 19.3944
R4739 VDD.n1900 VDD.n1246 19.3944
R4740 VDD.n1904 VDD.n1246 19.3944
R4741 VDD.n1904 VDD.n1236 19.3944
R4742 VDD.n1916 VDD.n1236 19.3944
R4743 VDD.n1916 VDD.n1234 19.3944
R4744 VDD.n1920 VDD.n1234 19.3944
R4745 VDD.n1920 VDD.n1224 19.3944
R4746 VDD.n1932 VDD.n1224 19.3944
R4747 VDD.n1932 VDD.n1222 19.3944
R4748 VDD.n1936 VDD.n1222 19.3944
R4749 VDD.n1936 VDD.n1212 19.3944
R4750 VDD.n1948 VDD.n1212 19.3944
R4751 VDD.n1948 VDD.n1209 19.3944
R4752 VDD.n1953 VDD.n1209 19.3944
R4753 VDD.n1953 VDD.n1210 19.3944
R4754 VDD.n1210 VDD.n1200 19.3944
R4755 VDD.n1967 VDD.n1200 19.3944
R4756 VDD.n1537 VDD.n1512 19.3944
R4757 VDD.n1533 VDD.n1512 19.3944
R4758 VDD.n1533 VDD.n1532 19.3944
R4759 VDD.n1532 VDD.n1531 19.3944
R4760 VDD.n1531 VDD.n1518 19.3944
R4761 VDD.n1527 VDD.n1518 19.3944
R4762 VDD.n1527 VDD.n1526 19.3944
R4763 VDD.n1526 VDD.n1525 19.3944
R4764 VDD.n1525 VDD.n1523 19.3944
R4765 VDD.n1554 VDD.n1553 19.3944
R4766 VDD.n1553 VDD.n1552 19.3944
R4767 VDD.n1552 VDD.n1500 19.3944
R4768 VDD.n1548 VDD.n1500 19.3944
R4769 VDD.n1548 VDD.n1547 19.3944
R4770 VDD.n1547 VDD.n1546 19.3944
R4771 VDD.n1546 VDD.n1506 19.3944
R4772 VDD.n1542 VDD.n1506 19.3944
R4773 VDD.n1542 VDD.n1541 19.3944
R4774 VDD.n1570 VDD.n1569 19.3944
R4775 VDD.n1569 VDD.n1480 19.3944
R4776 VDD.n1565 VDD.n1480 19.3944
R4777 VDD.n1565 VDD.n1564 19.3944
R4778 VDD.n1564 VDD.n1563 19.3944
R4779 VDD.n1563 VDD.n1486 19.3944
R4780 VDD.n1559 VDD.n1486 19.3944
R4781 VDD.n1559 VDD.n1558 19.3944
R4782 VDD.n1558 VDD.n1557 19.3944
R4783 VDD.n1586 VDD.n1585 19.3944
R4784 VDD.n1585 VDD.n1471 19.3944
R4785 VDD.n1581 VDD.n1471 19.3944
R4786 VDD.n1581 VDD.n1580 19.3944
R4787 VDD.n1580 VDD.n1579 19.3944
R4788 VDD.n1579 VDD.n1476 19.3944
R4789 VDD.n2104 VDD.n2101 19.3944
R4790 VDD.n2101 VDD.n2100 19.3944
R4791 VDD.n2100 VDD.n2097 19.3944
R4792 VDD.n2097 VDD.n2096 19.3944
R4793 VDD.n2096 VDD.n2093 19.3944
R4794 VDD.n2093 VDD.n2092 19.3944
R4795 VDD.n2092 VDD.n2089 19.3944
R4796 VDD.n2089 VDD.n2088 19.3944
R4797 VDD.n2088 VDD.n2085 19.3944
R4798 VDD.n2127 VDD.n2124 19.3944
R4799 VDD.n2124 VDD.n2123 19.3944
R4800 VDD.n2123 VDD.n2120 19.3944
R4801 VDD.n2120 VDD.n2119 19.3944
R4802 VDD.n2119 VDD.n2116 19.3944
R4803 VDD.n2116 VDD.n2115 19.3944
R4804 VDD.n2115 VDD.n2112 19.3944
R4805 VDD.n2112 VDD.n2111 19.3944
R4806 VDD.n2111 VDD.n2108 19.3944
R4807 VDD.n2149 VDD.n1167 19.3944
R4808 VDD.n2149 VDD.n2146 19.3944
R4809 VDD.n2146 VDD.n2143 19.3944
R4810 VDD.n2143 VDD.n2142 19.3944
R4811 VDD.n2142 VDD.n2139 19.3944
R4812 VDD.n2139 VDD.n2138 19.3944
R4813 VDD.n2138 VDD.n2135 19.3944
R4814 VDD.n2135 VDD.n2134 19.3944
R4815 VDD.n2134 VDD.n2131 19.3944
R4816 VDD.n2167 VDD.n1139 19.3944
R4817 VDD.n2162 VDD.n1139 19.3944
R4818 VDD.n2162 VDD.n2161 19.3944
R4819 VDD.n2161 VDD.n2160 19.3944
R4820 VDD.n2160 VDD.n2157 19.3944
R4821 VDD.n2157 VDD.n2156 19.3944
R4822 VDD.n1600 VDD.n1441 19.3944
R4823 VDD.n1600 VDD.n1439 19.3944
R4824 VDD.n1604 VDD.n1439 19.3944
R4825 VDD.n1604 VDD.n1430 19.3944
R4826 VDD.n1616 VDD.n1430 19.3944
R4827 VDD.n1616 VDD.n1428 19.3944
R4828 VDD.n1620 VDD.n1428 19.3944
R4829 VDD.n1620 VDD.n1418 19.3944
R4830 VDD.n1632 VDD.n1418 19.3944
R4831 VDD.n1632 VDD.n1416 19.3944
R4832 VDD.n1636 VDD.n1416 19.3944
R4833 VDD.n1636 VDD.n1406 19.3944
R4834 VDD.n1649 VDD.n1406 19.3944
R4835 VDD.n1649 VDD.n1404 19.3944
R4836 VDD.n1653 VDD.n1404 19.3944
R4837 VDD.n1653 VDD.n1395 19.3944
R4838 VDD.n1665 VDD.n1395 19.3944
R4839 VDD.n1665 VDD.n1393 19.3944
R4840 VDD.n1669 VDD.n1393 19.3944
R4841 VDD.n1669 VDD.n1383 19.3944
R4842 VDD.n1682 VDD.n1383 19.3944
R4843 VDD.n1682 VDD.n1381 19.3944
R4844 VDD.n1686 VDD.n1381 19.3944
R4845 VDD.n1686 VDD.n1372 19.3944
R4846 VDD.n1698 VDD.n1372 19.3944
R4847 VDD.n1698 VDD.n1370 19.3944
R4848 VDD.n1702 VDD.n1370 19.3944
R4849 VDD.n1702 VDD.n1360 19.3944
R4850 VDD.n1715 VDD.n1360 19.3944
R4851 VDD.n1715 VDD.n1358 19.3944
R4852 VDD.n1719 VDD.n1358 19.3944
R4853 VDD.n1719 VDD.n1349 19.3944
R4854 VDD.n1731 VDD.n1349 19.3944
R4855 VDD.n1731 VDD.n1347 19.3944
R4856 VDD.n1735 VDD.n1347 19.3944
R4857 VDD.n1735 VDD.n1337 19.3944
R4858 VDD.n1748 VDD.n1337 19.3944
R4859 VDD.n1748 VDD.n1335 19.3944
R4860 VDD.n1752 VDD.n1335 19.3944
R4861 VDD.n1752 VDD.n1326 19.3944
R4862 VDD.n1764 VDD.n1326 19.3944
R4863 VDD.n1764 VDD.n1324 19.3944
R4864 VDD.n1800 VDD.n1324 19.3944
R4865 VDD.n1800 VDD.n1314 19.3944
R4866 VDD.n1812 VDD.n1314 19.3944
R4867 VDD.n1812 VDD.n1312 19.3944
R4868 VDD.n1816 VDD.n1312 19.3944
R4869 VDD.n1816 VDD.n1302 19.3944
R4870 VDD.n1828 VDD.n1302 19.3944
R4871 VDD.n1828 VDD.n1300 19.3944
R4872 VDD.n1832 VDD.n1300 19.3944
R4873 VDD.n1832 VDD.n1290 19.3944
R4874 VDD.n1844 VDD.n1290 19.3944
R4875 VDD.n1844 VDD.n1288 19.3944
R4876 VDD.n1848 VDD.n1288 19.3944
R4877 VDD.n1848 VDD.n1278 19.3944
R4878 VDD.n1860 VDD.n1278 19.3944
R4879 VDD.n1860 VDD.n1276 19.3944
R4880 VDD.n1864 VDD.n1276 19.3944
R4881 VDD.n1864 VDD.n1266 19.3944
R4882 VDD.n1876 VDD.n1266 19.3944
R4883 VDD.n1876 VDD.n1264 19.3944
R4884 VDD.n1880 VDD.n1264 19.3944
R4885 VDD.n1880 VDD.n1254 19.3944
R4886 VDD.n1892 VDD.n1254 19.3944
R4887 VDD.n1892 VDD.n1252 19.3944
R4888 VDD.n1896 VDD.n1252 19.3944
R4889 VDD.n1896 VDD.n1242 19.3944
R4890 VDD.n1908 VDD.n1242 19.3944
R4891 VDD.n1908 VDD.n1240 19.3944
R4892 VDD.n1912 VDD.n1240 19.3944
R4893 VDD.n1912 VDD.n1230 19.3944
R4894 VDD.n1924 VDD.n1230 19.3944
R4895 VDD.n1924 VDD.n1228 19.3944
R4896 VDD.n1928 VDD.n1228 19.3944
R4897 VDD.n1928 VDD.n1218 19.3944
R4898 VDD.n1940 VDD.n1218 19.3944
R4899 VDD.n1940 VDD.n1216 19.3944
R4900 VDD.n1944 VDD.n1216 19.3944
R4901 VDD.n1944 VDD.n1206 19.3944
R4902 VDD.n1957 VDD.n1206 19.3944
R4903 VDD.n1957 VDD.n1204 19.3944
R4904 VDD.n1962 VDD.n1204 19.3944
R4905 VDD.n1962 VDD.n1961 19.3944
R4906 VDD.n3610 VDD.n391 19.3944
R4907 VDD.n3614 VDD.n391 19.3944
R4908 VDD.n3614 VDD.n381 19.3944
R4909 VDD.n3625 VDD.n381 19.3944
R4910 VDD.n3625 VDD.n379 19.3944
R4911 VDD.n3629 VDD.n379 19.3944
R4912 VDD.n3629 VDD.n369 19.3944
R4913 VDD.n3641 VDD.n369 19.3944
R4914 VDD.n3641 VDD.n367 19.3944
R4915 VDD.n3645 VDD.n367 19.3944
R4916 VDD.n3645 VDD.n357 19.3944
R4917 VDD.n3657 VDD.n357 19.3944
R4918 VDD.n3657 VDD.n355 19.3944
R4919 VDD.n3661 VDD.n355 19.3944
R4920 VDD.n3661 VDD.n345 19.3944
R4921 VDD.n3673 VDD.n345 19.3944
R4922 VDD.n3673 VDD.n343 19.3944
R4923 VDD.n3677 VDD.n343 19.3944
R4924 VDD.n3677 VDD.n333 19.3944
R4925 VDD.n3689 VDD.n333 19.3944
R4926 VDD.n3689 VDD.n331 19.3944
R4927 VDD.n3693 VDD.n331 19.3944
R4928 VDD.n3693 VDD.n321 19.3944
R4929 VDD.n3705 VDD.n321 19.3944
R4930 VDD.n3705 VDD.n319 19.3944
R4931 VDD.n3709 VDD.n319 19.3944
R4932 VDD.n3709 VDD.n309 19.3944
R4933 VDD.n3721 VDD.n309 19.3944
R4934 VDD.n3721 VDD.n307 19.3944
R4935 VDD.n3725 VDD.n307 19.3944
R4936 VDD.n3725 VDD.n297 19.3944
R4937 VDD.n3737 VDD.n297 19.3944
R4938 VDD.n3737 VDD.n295 19.3944
R4939 VDD.n3741 VDD.n295 19.3944
R4940 VDD.n3741 VDD.n285 19.3944
R4941 VDD.n3753 VDD.n285 19.3944
R4942 VDD.n3753 VDD.n283 19.3944
R4943 VDD.n3757 VDD.n283 19.3944
R4944 VDD.n3757 VDD.n272 19.3944
R4945 VDD.n3769 VDD.n272 19.3944
R4946 VDD.n3769 VDD.n270 19.3944
R4947 VDD.n3773 VDD.n270 19.3944
R4948 VDD.n3774 VDD.n3773 19.3944
R4949 VDD.n3775 VDD.n3774 19.3944
R4950 VDD.n3775 VDD.n268 19.3944
R4951 VDD.n3779 VDD.n268 19.3944
R4952 VDD.n3780 VDD.n3779 19.3944
R4953 VDD.n3781 VDD.n3780 19.3944
R4954 VDD.n3781 VDD.n265 19.3944
R4955 VDD.n3785 VDD.n265 19.3944
R4956 VDD.n3786 VDD.n3785 19.3944
R4957 VDD.n3787 VDD.n3786 19.3944
R4958 VDD.n3787 VDD.n262 19.3944
R4959 VDD.n3791 VDD.n262 19.3944
R4960 VDD.n3792 VDD.n3791 19.3944
R4961 VDD.n3793 VDD.n3792 19.3944
R4962 VDD.n3793 VDD.n259 19.3944
R4963 VDD.n3797 VDD.n259 19.3944
R4964 VDD.n3798 VDD.n3797 19.3944
R4965 VDD.n3799 VDD.n3798 19.3944
R4966 VDD.n3799 VDD.n256 19.3944
R4967 VDD.n3803 VDD.n256 19.3944
R4968 VDD.n3804 VDD.n3803 19.3944
R4969 VDD.n3805 VDD.n3804 19.3944
R4970 VDD.n3805 VDD.n253 19.3944
R4971 VDD.n3809 VDD.n253 19.3944
R4972 VDD.n3810 VDD.n3809 19.3944
R4973 VDD.n3811 VDD.n3810 19.3944
R4974 VDD.n3811 VDD.n250 19.3944
R4975 VDD.n3815 VDD.n250 19.3944
R4976 VDD.n3816 VDD.n3815 19.3944
R4977 VDD.n3817 VDD.n3816 19.3944
R4978 VDD.n3817 VDD.n247 19.3944
R4979 VDD.n3821 VDD.n247 19.3944
R4980 VDD.n3822 VDD.n3821 19.3944
R4981 VDD.n3823 VDD.n3822 19.3944
R4982 VDD.n3823 VDD.n244 19.3944
R4983 VDD.n3827 VDD.n244 19.3944
R4984 VDD.n3828 VDD.n3827 19.3944
R4985 VDD.n3829 VDD.n3828 19.3944
R4986 VDD.n3829 VDD.n241 19.3944
R4987 VDD.n3833 VDD.n241 19.3944
R4988 VDD.n3834 VDD.n3833 19.3944
R4989 VDD.n3835 VDD.n3834 19.3944
R4990 VDD.n3859 VDD.n3858 19.3944
R4991 VDD.n3858 VDD.n3857 19.3944
R4992 VDD.n3857 VDD.n226 19.3944
R4993 VDD.n3852 VDD.n226 19.3944
R4994 VDD.n3852 VDD.n3851 19.3944
R4995 VDD.n3851 VDD.n3850 19.3944
R4996 VDD.n3850 VDD.n233 19.3944
R4997 VDD.n3845 VDD.n233 19.3944
R4998 VDD.n3845 VDD.n3844 19.3944
R4999 VDD.n3878 VDD.n202 19.3944
R5000 VDD.n3873 VDD.n202 19.3944
R5001 VDD.n3873 VDD.n3872 19.3944
R5002 VDD.n3872 VDD.n3871 19.3944
R5003 VDD.n3871 VDD.n209 19.3944
R5004 VDD.n3866 VDD.n209 19.3944
R5005 VDD.n3866 VDD.n3865 19.3944
R5006 VDD.n3865 VDD.n3864 19.3944
R5007 VDD.n3864 VDD.n216 19.3944
R5008 VDD.n3897 VDD.n3896 19.3944
R5009 VDD.n3896 VDD.n3895 19.3944
R5010 VDD.n3895 VDD.n188 19.3944
R5011 VDD.n3890 VDD.n188 19.3944
R5012 VDD.n3890 VDD.n3889 19.3944
R5013 VDD.n3889 VDD.n3888 19.3944
R5014 VDD.n3888 VDD.n195 19.3944
R5015 VDD.n3883 VDD.n195 19.3944
R5016 VDD.n3883 VDD.n3882 19.3944
R5017 VDD.n3911 VDD.n3910 19.3944
R5018 VDD.n3910 VDD.n3909 19.3944
R5019 VDD.n3909 VDD.n172 19.3944
R5020 VDD.n3904 VDD.n172 19.3944
R5021 VDD.n3904 VDD.n3903 19.3944
R5022 VDD.n3903 VDD.n3902 19.3944
R5023 VDD.n3606 VDD.n387 19.3944
R5024 VDD.n3618 VDD.n387 19.3944
R5025 VDD.n3618 VDD.n385 19.3944
R5026 VDD.n3622 VDD.n385 19.3944
R5027 VDD.n3622 VDD.n375 19.3944
R5028 VDD.n3633 VDD.n375 19.3944
R5029 VDD.n3633 VDD.n373 19.3944
R5030 VDD.n3637 VDD.n373 19.3944
R5031 VDD.n3637 VDD.n363 19.3944
R5032 VDD.n3649 VDD.n363 19.3944
R5033 VDD.n3649 VDD.n361 19.3944
R5034 VDD.n3653 VDD.n361 19.3944
R5035 VDD.n3653 VDD.n351 19.3944
R5036 VDD.n3665 VDD.n351 19.3944
R5037 VDD.n3665 VDD.n349 19.3944
R5038 VDD.n3669 VDD.n349 19.3944
R5039 VDD.n3669 VDD.n339 19.3944
R5040 VDD.n3681 VDD.n339 19.3944
R5041 VDD.n3681 VDD.n337 19.3944
R5042 VDD.n3685 VDD.n337 19.3944
R5043 VDD.n3685 VDD.n327 19.3944
R5044 VDD.n3697 VDD.n327 19.3944
R5045 VDD.n3697 VDD.n325 19.3944
R5046 VDD.n3701 VDD.n325 19.3944
R5047 VDD.n3701 VDD.n315 19.3944
R5048 VDD.n3713 VDD.n315 19.3944
R5049 VDD.n3713 VDD.n313 19.3944
R5050 VDD.n3717 VDD.n313 19.3944
R5051 VDD.n3717 VDD.n303 19.3944
R5052 VDD.n3729 VDD.n303 19.3944
R5053 VDD.n3729 VDD.n301 19.3944
R5054 VDD.n3733 VDD.n301 19.3944
R5055 VDD.n3733 VDD.n291 19.3944
R5056 VDD.n3745 VDD.n291 19.3944
R5057 VDD.n3745 VDD.n289 19.3944
R5058 VDD.n3749 VDD.n289 19.3944
R5059 VDD.n3749 VDD.n279 19.3944
R5060 VDD.n3761 VDD.n279 19.3944
R5061 VDD.n3761 VDD.n277 19.3944
R5062 VDD.n3765 VDD.n277 19.3944
R5063 VDD.n3765 VDD.n49 19.3944
R5064 VDD.n3999 VDD.n49 19.3944
R5065 VDD.n3999 VDD.n50 19.3944
R5066 VDD.n3993 VDD.n50 19.3944
R5067 VDD.n3993 VDD.n3992 19.3944
R5068 VDD.n3992 VDD.n3991 19.3944
R5069 VDD.n3991 VDD.n62 19.3944
R5070 VDD.n3985 VDD.n62 19.3944
R5071 VDD.n3985 VDD.n3984 19.3944
R5072 VDD.n3984 VDD.n3983 19.3944
R5073 VDD.n3983 VDD.n73 19.3944
R5074 VDD.n3977 VDD.n73 19.3944
R5075 VDD.n3977 VDD.n3976 19.3944
R5076 VDD.n3976 VDD.n3975 19.3944
R5077 VDD.n3975 VDD.n84 19.3944
R5078 VDD.n3969 VDD.n84 19.3944
R5079 VDD.n3969 VDD.n3968 19.3944
R5080 VDD.n3968 VDD.n3967 19.3944
R5081 VDD.n3967 VDD.n95 19.3944
R5082 VDD.n3961 VDD.n95 19.3944
R5083 VDD.n3961 VDD.n3960 19.3944
R5084 VDD.n3960 VDD.n3959 19.3944
R5085 VDD.n3959 VDD.n106 19.3944
R5086 VDD.n3953 VDD.n106 19.3944
R5087 VDD.n3953 VDD.n3952 19.3944
R5088 VDD.n3952 VDD.n3951 19.3944
R5089 VDD.n3951 VDD.n117 19.3944
R5090 VDD.n3945 VDD.n117 19.3944
R5091 VDD.n3945 VDD.n3944 19.3944
R5092 VDD.n3944 VDD.n3943 19.3944
R5093 VDD.n3943 VDD.n128 19.3944
R5094 VDD.n3937 VDD.n128 19.3944
R5095 VDD.n3937 VDD.n3936 19.3944
R5096 VDD.n3936 VDD.n3935 19.3944
R5097 VDD.n3935 VDD.n139 19.3944
R5098 VDD.n3929 VDD.n139 19.3944
R5099 VDD.n3929 VDD.n3928 19.3944
R5100 VDD.n3928 VDD.n3927 19.3944
R5101 VDD.n3927 VDD.n150 19.3944
R5102 VDD.n3922 VDD.n150 19.3944
R5103 VDD.n3922 VDD.n3921 19.3944
R5104 VDD.n3921 VDD.n3920 19.3944
R5105 VDD.n3920 VDD.n161 19.3944
R5106 VDD.n3914 VDD.n161 19.3944
R5107 VDD.n3603 VDD.n3602 19.3944
R5108 VDD.n3602 VDD.n3462 19.3944
R5109 VDD.n3597 VDD.n3462 19.3944
R5110 VDD.n3597 VDD.n3596 19.3944
R5111 VDD.n3596 VDD.n3467 19.3944
R5112 VDD.n3591 VDD.n3467 19.3944
R5113 VDD.n3589 VDD.n3475 19.3944
R5114 VDD.n3583 VDD.n3475 19.3944
R5115 VDD.n3583 VDD.n3582 19.3944
R5116 VDD.n3582 VDD.n3581 19.3944
R5117 VDD.n3581 VDD.n3481 19.3944
R5118 VDD.n3575 VDD.n3481 19.3944
R5119 VDD.n3575 VDD.n3574 19.3944
R5120 VDD.n3574 VDD.n3573 19.3944
R5121 VDD.n3573 VDD.n3487 19.3944
R5122 VDD.n3567 VDD.n3566 19.3944
R5123 VDD.n3566 VDD.n3565 19.3944
R5124 VDD.n3565 VDD.n3496 19.3944
R5125 VDD.n3559 VDD.n3496 19.3944
R5126 VDD.n3559 VDD.n3558 19.3944
R5127 VDD.n3558 VDD.n3557 19.3944
R5128 VDD.n3557 VDD.n3502 19.3944
R5129 VDD.n3551 VDD.n3502 19.3944
R5130 VDD.n3551 VDD.n3550 19.3944
R5131 VDD.n3548 VDD.n3510 19.3944
R5132 VDD.n3542 VDD.n3510 19.3944
R5133 VDD.n3542 VDD.n3541 19.3944
R5134 VDD.n3541 VDD.n3540 19.3944
R5135 VDD.n3540 VDD.n3516 19.3944
R5136 VDD.n3534 VDD.n3516 19.3944
R5137 VDD.n3534 VDD.n3533 19.3944
R5138 VDD.n3533 VDD.n3532 19.3944
R5139 VDD.n3532 VDD.n3527 19.3944
R5140 VDD.n1575 VDD.n1476 18.8126
R5141 VDD.n2156 VDD.n2153 18.8126
R5142 VDD.n3902 VDD.n181 18.8126
R5143 VDD.n3591 VDD.n3590 18.8126
R5144 VDD.n1598 VDD.n1443 15.1279
R5145 VDD.n1598 VDD.n1437 15.1279
R5146 VDD.n1606 VDD.n1437 15.1279
R5147 VDD.n1606 VDD.t17 15.1279
R5148 VDD.n1614 VDD.t17 15.1279
R5149 VDD.n1614 VDD.n1426 15.1279
R5150 VDD.n1622 VDD.n1426 15.1279
R5151 VDD.n1622 VDD.n1420 15.1279
R5152 VDD.n1630 VDD.n1420 15.1279
R5153 VDD.n1630 VDD.n1414 15.1279
R5154 VDD.n1638 VDD.n1414 15.1279
R5155 VDD.n1638 VDD.n1408 15.1279
R5156 VDD.n1647 VDD.n1408 15.1279
R5157 VDD.n1647 VDD.n1646 15.1279
R5158 VDD.n1655 VDD.n1397 15.1279
R5159 VDD.n1663 VDD.n1397 15.1279
R5160 VDD.n1663 VDD.n1391 15.1279
R5161 VDD.n1671 VDD.n1391 15.1279
R5162 VDD.n1671 VDD.n1385 15.1279
R5163 VDD.n1680 VDD.n1385 15.1279
R5164 VDD.n1680 VDD.n1679 15.1279
R5165 VDD.n1688 VDD.n1374 15.1279
R5166 VDD.n1696 VDD.n1374 15.1279
R5167 VDD.n1696 VDD.n1368 15.1279
R5168 VDD.n1704 VDD.n1368 15.1279
R5169 VDD.n1704 VDD.n1362 15.1279
R5170 VDD.n1713 VDD.n1362 15.1279
R5171 VDD.n1713 VDD.n1712 15.1279
R5172 VDD.n1721 VDD.n1351 15.1279
R5173 VDD.n1729 VDD.n1351 15.1279
R5174 VDD.n1729 VDD.n1345 15.1279
R5175 VDD.n1737 VDD.n1345 15.1279
R5176 VDD.n1737 VDD.n1339 15.1279
R5177 VDD.n1746 VDD.n1339 15.1279
R5178 VDD.n1746 VDD.n1745 15.1279
R5179 VDD.n1754 VDD.n1328 15.1279
R5180 VDD.n1762 VDD.n1328 15.1279
R5181 VDD.n1762 VDD.n1322 15.1279
R5182 VDD.n1802 VDD.n1322 15.1279
R5183 VDD.n1802 VDD.n1316 15.1279
R5184 VDD.n1810 VDD.n1316 15.1279
R5185 VDD.n1818 VDD.n1310 15.1279
R5186 VDD.n1818 VDD.n1304 15.1279
R5187 VDD.n1826 VDD.n1304 15.1279
R5188 VDD.n1826 VDD.n1298 15.1279
R5189 VDD.n1834 VDD.n1298 15.1279
R5190 VDD.n1834 VDD.n1292 15.1279
R5191 VDD.n1842 VDD.n1292 15.1279
R5192 VDD.n1850 VDD.n1286 15.1279
R5193 VDD.n1850 VDD.n1280 15.1279
R5194 VDD.n1858 VDD.n1280 15.1279
R5195 VDD.n1858 VDD.n1274 15.1279
R5196 VDD.n1866 VDD.n1274 15.1279
R5197 VDD.n1866 VDD.n1268 15.1279
R5198 VDD.n1874 VDD.n1268 15.1279
R5199 VDD.n1882 VDD.n1262 15.1279
R5200 VDD.n1882 VDD.n1256 15.1279
R5201 VDD.n1890 VDD.n1256 15.1279
R5202 VDD.n1890 VDD.n1250 15.1279
R5203 VDD.n1898 VDD.n1250 15.1279
R5204 VDD.n1898 VDD.n1244 15.1279
R5205 VDD.n1906 VDD.n1244 15.1279
R5206 VDD.n1914 VDD.n1238 15.1279
R5207 VDD.n1914 VDD.n1232 15.1279
R5208 VDD.n1922 VDD.n1232 15.1279
R5209 VDD.n1922 VDD.n1226 15.1279
R5210 VDD.n1930 VDD.n1226 15.1279
R5211 VDD.n1930 VDD.n1220 15.1279
R5212 VDD.n1938 VDD.n1220 15.1279
R5213 VDD.n1938 VDD.n1214 15.1279
R5214 VDD.n1946 VDD.n1214 15.1279
R5215 VDD.n1946 VDD.t28 15.1279
R5216 VDD.n1955 VDD.t28 15.1279
R5217 VDD.n1955 VDD.n1202 15.1279
R5218 VDD.n1964 VDD.n1202 15.1279
R5219 VDD.n1964 VDD.n1142 15.1279
R5220 VDD.n3608 VDD.n389 15.1279
R5221 VDD.n3616 VDD.n389 15.1279
R5222 VDD.n3616 VDD.n383 15.1279
R5223 VDD.t13 VDD.n383 15.1279
R5224 VDD.t13 VDD.n377 15.1279
R5225 VDD.n3631 VDD.n377 15.1279
R5226 VDD.n3631 VDD.n371 15.1279
R5227 VDD.n3639 VDD.n371 15.1279
R5228 VDD.n3639 VDD.n365 15.1279
R5229 VDD.n3647 VDD.n365 15.1279
R5230 VDD.n3647 VDD.n359 15.1279
R5231 VDD.n3655 VDD.n359 15.1279
R5232 VDD.n3655 VDD.n353 15.1279
R5233 VDD.n3663 VDD.n353 15.1279
R5234 VDD.n3671 VDD.n347 15.1279
R5235 VDD.n3671 VDD.n341 15.1279
R5236 VDD.n3679 VDD.n341 15.1279
R5237 VDD.n3679 VDD.n335 15.1279
R5238 VDD.n3687 VDD.n335 15.1279
R5239 VDD.n3687 VDD.n329 15.1279
R5240 VDD.n3695 VDD.n329 15.1279
R5241 VDD.n3703 VDD.n323 15.1279
R5242 VDD.n3703 VDD.n317 15.1279
R5243 VDD.n3711 VDD.n317 15.1279
R5244 VDD.n3711 VDD.n311 15.1279
R5245 VDD.n3719 VDD.n311 15.1279
R5246 VDD.n3719 VDD.n305 15.1279
R5247 VDD.n3727 VDD.n305 15.1279
R5248 VDD.n3735 VDD.n299 15.1279
R5249 VDD.n3735 VDD.n293 15.1279
R5250 VDD.n3743 VDD.n293 15.1279
R5251 VDD.n3743 VDD.n287 15.1279
R5252 VDD.n3751 VDD.n287 15.1279
R5253 VDD.n3751 VDD.n281 15.1279
R5254 VDD.n3759 VDD.n281 15.1279
R5255 VDD.n3767 VDD.n275 15.1279
R5256 VDD.n3767 VDD.n53 15.1279
R5257 VDD.n3997 VDD.n53 15.1279
R5258 VDD.n3997 VDD.n3996 15.1279
R5259 VDD.n3996 VDD.n3995 15.1279
R5260 VDD.n3995 VDD.n57 15.1279
R5261 VDD.n3989 VDD.n3988 15.1279
R5262 VDD.n3988 VDD.n3987 15.1279
R5263 VDD.n3987 VDD.n67 15.1279
R5264 VDD.n3981 VDD.n67 15.1279
R5265 VDD.n3981 VDD.n3980 15.1279
R5266 VDD.n3980 VDD.n3979 15.1279
R5267 VDD.n3979 VDD.n78 15.1279
R5268 VDD.n3973 VDD.n3972 15.1279
R5269 VDD.n3972 VDD.n3971 15.1279
R5270 VDD.n3971 VDD.n89 15.1279
R5271 VDD.n3965 VDD.n89 15.1279
R5272 VDD.n3965 VDD.n3964 15.1279
R5273 VDD.n3964 VDD.n3963 15.1279
R5274 VDD.n3963 VDD.n100 15.1279
R5275 VDD.n3957 VDD.n3956 15.1279
R5276 VDD.n3956 VDD.n3955 15.1279
R5277 VDD.n3955 VDD.n111 15.1279
R5278 VDD.n3949 VDD.n111 15.1279
R5279 VDD.n3949 VDD.n3948 15.1279
R5280 VDD.n3948 VDD.n3947 15.1279
R5281 VDD.n3947 VDD.n122 15.1279
R5282 VDD.n3941 VDD.n3940 15.1279
R5283 VDD.n3940 VDD.n3939 15.1279
R5284 VDD.n3939 VDD.n133 15.1279
R5285 VDD.n3933 VDD.n133 15.1279
R5286 VDD.n3933 VDD.n3932 15.1279
R5287 VDD.n3932 VDD.n3931 15.1279
R5288 VDD.n3931 VDD.n144 15.1279
R5289 VDD.n3925 VDD.n144 15.1279
R5290 VDD.n3925 VDD.n3924 15.1279
R5291 VDD.n3924 VDD.t24 15.1279
R5292 VDD.t24 VDD.n155 15.1279
R5293 VDD.n3918 VDD.n155 15.1279
R5294 VDD.n3918 VDD.n3917 15.1279
R5295 VDD.n3917 VDD.n3916 15.1279
R5296 VDD.n43 VDD.t173 14.9798
R5297 VDD.n43 VDD.t130 14.9798
R5298 VDD.n41 VDD.t170 14.9798
R5299 VDD.n41 VDD.t139 14.9798
R5300 VDD.n39 VDD.t128 14.9798
R5301 VDD.n39 VDD.t133 14.9798
R5302 VDD.n35 VDD.t141 14.9798
R5303 VDD.n35 VDD.t177 14.9798
R5304 VDD.n33 VDD.t136 14.9798
R5305 VDD.n33 VDD.t184 14.9798
R5306 VDD.n31 VDD.t131 14.9798
R5307 VDD.n31 VDD.t181 14.9798
R5308 VDD.n27 VDD.t197 14.9798
R5309 VDD.n27 VDD.t191 14.9798
R5310 VDD.n25 VDD.t172 14.9798
R5311 VDD.n25 VDD.t138 14.9798
R5312 VDD.n23 VDD.t134 14.9798
R5313 VDD.n23 VDD.t179 14.9798
R5314 VDD.n20 VDD.t151 14.9798
R5315 VDD.n20 VDD.t146 14.9798
R5316 VDD.n18 VDD.t190 14.9798
R5317 VDD.n18 VDD.t167 14.9798
R5318 VDD.n16 VDD.t162 14.9798
R5319 VDD.n16 VDD.t121 14.9798
R5320 VDD.n1789 VDD.t153 14.9798
R5321 VDD.n1789 VDD.t185 14.9798
R5322 VDD.n1791 VDD.t126 14.9798
R5323 VDD.n1791 VDD.t125 14.9798
R5324 VDD.n1793 VDD.t180 14.9798
R5325 VDD.n1793 VDD.t155 14.9798
R5326 VDD.n1781 VDD.t192 14.9798
R5327 VDD.n1781 VDD.t161 14.9798
R5328 VDD.n1783 VDD.t152 14.9798
R5329 VDD.n1783 VDD.t176 14.9798
R5330 VDD.n1785 VDD.t157 14.9798
R5331 VDD.n1785 VDD.t196 14.9798
R5332 VDD.n1773 VDD.t188 14.9798
R5333 VDD.n1773 VDD.t195 14.9798
R5334 VDD.n1775 VDD.t123 14.9798
R5335 VDD.n1775 VDD.t160 14.9798
R5336 VDD.n1777 VDD.t168 14.9798
R5337 VDD.n1777 VDD.t175 14.9798
R5338 VDD.n1766 VDD.t143 14.9798
R5339 VDD.n1766 VDD.t150 14.9798
R5340 VDD.n1768 VDD.t163 14.9798
R5341 VDD.n1768 VDD.t183 14.9798
R5342 VDD.n1770 VDD.t186 14.9798
R5343 VDD.n1770 VDD.t193 14.9798
R5344 VDD.n1754 VDD.t122 14.8253
R5345 VDD.n1810 VDD.t124 14.8253
R5346 VDD.t135 VDD.n275 14.8253
R5347 VDD.t137 VDD.n57 14.8253
R5348 VDD.n1721 VDD.t154 14.2202
R5349 VDD.n1842 VDD.t142 14.2202
R5350 VDD.t120 VDD.n299 14.2202
R5351 VDD.t140 VDD.n78 14.2202
R5352 VDD.n1688 VDD.t156 13.6151
R5353 VDD.n1874 VDD.t149 13.6151
R5354 VDD.t127 VDD.n323 13.6151
R5355 VDD.t129 VDD.n100 13.6151
R5356 VDD.n1655 VDD.t147 13.0101
R5357 VDD.n1906 VDD.t118 13.0101
R5358 VDD.t144 VDD.n347 13.0101
R5359 VDD.t158 VDD.n122 13.0101
R5360 VDD.n2201 VDD.n1012 10.6151
R5361 VDD.n2202 VDD.n2201 10.6151
R5362 VDD.n2203 VDD.n2202 10.6151
R5363 VDD.n2203 VDD.n999 10.6151
R5364 VDD.n2213 VDD.n999 10.6151
R5365 VDD.n2214 VDD.n2213 10.6151
R5366 VDD.n2215 VDD.n2214 10.6151
R5367 VDD.n2215 VDD.n988 10.6151
R5368 VDD.n2225 VDD.n988 10.6151
R5369 VDD.n2226 VDD.n2225 10.6151
R5370 VDD.n2227 VDD.n2226 10.6151
R5371 VDD.n2227 VDD.n976 10.6151
R5372 VDD.n2237 VDD.n976 10.6151
R5373 VDD.n2238 VDD.n2237 10.6151
R5374 VDD.n2239 VDD.n2238 10.6151
R5375 VDD.n2239 VDD.n964 10.6151
R5376 VDD.n2249 VDD.n964 10.6151
R5377 VDD.n2250 VDD.n2249 10.6151
R5378 VDD.n2251 VDD.n2250 10.6151
R5379 VDD.n2251 VDD.n952 10.6151
R5380 VDD.n2261 VDD.n952 10.6151
R5381 VDD.n2262 VDD.n2261 10.6151
R5382 VDD.n2263 VDD.n2262 10.6151
R5383 VDD.n2263 VDD.n940 10.6151
R5384 VDD.n2273 VDD.n940 10.6151
R5385 VDD.n2274 VDD.n2273 10.6151
R5386 VDD.n2275 VDD.n2274 10.6151
R5387 VDD.n2275 VDD.n928 10.6151
R5388 VDD.n2285 VDD.n928 10.6151
R5389 VDD.n2286 VDD.n2285 10.6151
R5390 VDD.n2287 VDD.n2286 10.6151
R5391 VDD.n2287 VDD.n916 10.6151
R5392 VDD.n2297 VDD.n916 10.6151
R5393 VDD.n2298 VDD.n2297 10.6151
R5394 VDD.n2299 VDD.n2298 10.6151
R5395 VDD.n2299 VDD.n904 10.6151
R5396 VDD.n2309 VDD.n904 10.6151
R5397 VDD.n2310 VDD.n2309 10.6151
R5398 VDD.n2311 VDD.n2310 10.6151
R5399 VDD.n2311 VDD.n891 10.6151
R5400 VDD.n2326 VDD.n891 10.6151
R5401 VDD.n2327 VDD.n2326 10.6151
R5402 VDD.n2328 VDD.n2327 10.6151
R5403 VDD.n2328 VDD.n875 10.6151
R5404 VDD.n2461 VDD.n875 10.6151
R5405 VDD.n2462 VDD.n2461 10.6151
R5406 VDD.n2463 VDD.n2462 10.6151
R5407 VDD.n2463 VDD.n863 10.6151
R5408 VDD.n2473 VDD.n863 10.6151
R5409 VDD.n2474 VDD.n2473 10.6151
R5410 VDD.n2475 VDD.n2474 10.6151
R5411 VDD.n2475 VDD.n851 10.6151
R5412 VDD.n2485 VDD.n851 10.6151
R5413 VDD.n2486 VDD.n2485 10.6151
R5414 VDD.n2487 VDD.n2486 10.6151
R5415 VDD.n2487 VDD.n839 10.6151
R5416 VDD.n2497 VDD.n839 10.6151
R5417 VDD.n2498 VDD.n2497 10.6151
R5418 VDD.n2499 VDD.n2498 10.6151
R5419 VDD.n2499 VDD.n827 10.6151
R5420 VDD.n2509 VDD.n827 10.6151
R5421 VDD.n2510 VDD.n2509 10.6151
R5422 VDD.n2511 VDD.n2510 10.6151
R5423 VDD.n2511 VDD.n815 10.6151
R5424 VDD.n2521 VDD.n815 10.6151
R5425 VDD.n2522 VDD.n2521 10.6151
R5426 VDD.n2523 VDD.n2522 10.6151
R5427 VDD.n2523 VDD.n803 10.6151
R5428 VDD.n2533 VDD.n803 10.6151
R5429 VDD.n2534 VDD.n2533 10.6151
R5430 VDD.n2535 VDD.n2534 10.6151
R5431 VDD.n2535 VDD.n791 10.6151
R5432 VDD.n2545 VDD.n791 10.6151
R5433 VDD.n2546 VDD.n2545 10.6151
R5434 VDD.n2547 VDD.n2546 10.6151
R5435 VDD.n2547 VDD.n779 10.6151
R5436 VDD.n2557 VDD.n779 10.6151
R5437 VDD.n2558 VDD.n2557 10.6151
R5438 VDD.n2559 VDD.n2558 10.6151
R5439 VDD.n2559 VDD.n767 10.6151
R5440 VDD.n2569 VDD.n767 10.6151
R5441 VDD.n2570 VDD.n2569 10.6151
R5442 VDD.n2571 VDD.n2570 10.6151
R5443 VDD.n2571 VDD.n755 10.6151
R5444 VDD.n2586 VDD.n755 10.6151
R5445 VDD.n2587 VDD.n2586 10.6151
R5446 VDD.n2588 VDD.n2587 10.6151
R5447 VDD.n2588 VDD.n746 10.6151
R5448 VDD.n2647 VDD.n746 10.6151
R5449 VDD.n2647 VDD.n2646 10.6151
R5450 VDD.n2645 VDD.n2643 10.6151
R5451 VDD.n2643 VDD.n2640 10.6151
R5452 VDD.n2640 VDD.n2639 10.6151
R5453 VDD.n2639 VDD.n2636 10.6151
R5454 VDD.n2636 VDD.n2635 10.6151
R5455 VDD.n2635 VDD.n2632 10.6151
R5456 VDD.n2632 VDD.n2631 10.6151
R5457 VDD.n2631 VDD.n2628 10.6151
R5458 VDD.n2628 VDD.n2627 10.6151
R5459 VDD.n2627 VDD.n2624 10.6151
R5460 VDD.n2624 VDD.n2623 10.6151
R5461 VDD.n2623 VDD.n2620 10.6151
R5462 VDD.n2620 VDD.n2619 10.6151
R5463 VDD.n2619 VDD.n2616 10.6151
R5464 VDD.n2616 VDD.n2615 10.6151
R5465 VDD.n2615 VDD.n2612 10.6151
R5466 VDD.n2612 VDD.n2611 10.6151
R5467 VDD.n2611 VDD.n2608 10.6151
R5468 VDD.n2608 VDD.n2607 10.6151
R5469 VDD.n2607 VDD.n2604 10.6151
R5470 VDD.n2602 VDD.n2599 10.6151
R5471 VDD.n2599 VDD.n2598 10.6151
R5472 VDD.n1113 VDD.n1111 10.6151
R5473 VDD.n1111 VDD.n1110 10.6151
R5474 VDD.n1110 VDD.n1108 10.6151
R5475 VDD.n1108 VDD.n1107 10.6151
R5476 VDD.n1107 VDD.n1105 10.6151
R5477 VDD.n1105 VDD.n1104 10.6151
R5478 VDD.n1104 VDD.n1102 10.6151
R5479 VDD.n1102 VDD.n1101 10.6151
R5480 VDD.n1101 VDD.n1099 10.6151
R5481 VDD.n1099 VDD.n1098 10.6151
R5482 VDD.n1098 VDD.n1096 10.6151
R5483 VDD.n1096 VDD.n1095 10.6151
R5484 VDD.n1095 VDD.n1093 10.6151
R5485 VDD.n1093 VDD.n1092 10.6151
R5486 VDD.n1092 VDD.n1090 10.6151
R5487 VDD.n1090 VDD.n1089 10.6151
R5488 VDD.n1089 VDD.n1087 10.6151
R5489 VDD.n1087 VDD.n1086 10.6151
R5490 VDD.n1086 VDD.n1084 10.6151
R5491 VDD.n1084 VDD.n1083 10.6151
R5492 VDD.n1083 VDD.n1081 10.6151
R5493 VDD.n1081 VDD.n1080 10.6151
R5494 VDD.n1080 VDD.n1078 10.6151
R5495 VDD.n1078 VDD.n1077 10.6151
R5496 VDD.n1077 VDD.n1075 10.6151
R5497 VDD.n1075 VDD.n1074 10.6151
R5498 VDD.n1074 VDD.n1072 10.6151
R5499 VDD.n1072 VDD.n1071 10.6151
R5500 VDD.n1071 VDD.n1069 10.6151
R5501 VDD.n1069 VDD.n1068 10.6151
R5502 VDD.n1068 VDD.n1066 10.6151
R5503 VDD.n1066 VDD.n1065 10.6151
R5504 VDD.n1065 VDD.n1063 10.6151
R5505 VDD.n1063 VDD.n1062 10.6151
R5506 VDD.n1062 VDD.n1060 10.6151
R5507 VDD.n1060 VDD.n1059 10.6151
R5508 VDD.n1059 VDD.n1057 10.6151
R5509 VDD.n1057 VDD.n1056 10.6151
R5510 VDD.n1056 VDD.n1054 10.6151
R5511 VDD.n1054 VDD.n1053 10.6151
R5512 VDD.n1053 VDD.n1051 10.6151
R5513 VDD.n1051 VDD.n1050 10.6151
R5514 VDD.n1050 VDD.n1048 10.6151
R5515 VDD.n1048 VDD.n882 10.6151
R5516 VDD.n2458 VDD.n882 10.6151
R5517 VDD.n2458 VDD.n2457 10.6151
R5518 VDD.n2457 VDD.n2456 10.6151
R5519 VDD.n2456 VDD.n2455 10.6151
R5520 VDD.n2455 VDD.n2453 10.6151
R5521 VDD.n2453 VDD.n2452 10.6151
R5522 VDD.n2452 VDD.n2450 10.6151
R5523 VDD.n2450 VDD.n2449 10.6151
R5524 VDD.n2449 VDD.n2447 10.6151
R5525 VDD.n2447 VDD.n2446 10.6151
R5526 VDD.n2446 VDD.n2444 10.6151
R5527 VDD.n2444 VDD.n2443 10.6151
R5528 VDD.n2443 VDD.n2441 10.6151
R5529 VDD.n2441 VDD.n2440 10.6151
R5530 VDD.n2440 VDD.n2438 10.6151
R5531 VDD.n2438 VDD.n2437 10.6151
R5532 VDD.n2437 VDD.n2435 10.6151
R5533 VDD.n2435 VDD.n2434 10.6151
R5534 VDD.n2434 VDD.n2432 10.6151
R5535 VDD.n2432 VDD.n2431 10.6151
R5536 VDD.n2431 VDD.n2429 10.6151
R5537 VDD.n2429 VDD.n2428 10.6151
R5538 VDD.n2428 VDD.n2426 10.6151
R5539 VDD.n2426 VDD.n2425 10.6151
R5540 VDD.n2425 VDD.n2423 10.6151
R5541 VDD.n2423 VDD.n2422 10.6151
R5542 VDD.n2422 VDD.n2420 10.6151
R5543 VDD.n2420 VDD.n2419 10.6151
R5544 VDD.n2419 VDD.n2417 10.6151
R5545 VDD.n2417 VDD.n2416 10.6151
R5546 VDD.n2416 VDD.n2414 10.6151
R5547 VDD.n2414 VDD.n2413 10.6151
R5548 VDD.n2413 VDD.n2411 10.6151
R5549 VDD.n2411 VDD.n2410 10.6151
R5550 VDD.n2410 VDD.n2408 10.6151
R5551 VDD.n2408 VDD.n2407 10.6151
R5552 VDD.n2407 VDD.n2405 10.6151
R5553 VDD.n2405 VDD.n2404 10.6151
R5554 VDD.n2404 VDD.n2402 10.6151
R5555 VDD.n2402 VDD.n2401 10.6151
R5556 VDD.n2401 VDD.n884 10.6151
R5557 VDD.n884 VDD.n883 10.6151
R5558 VDD.n883 VDD.n749 10.6151
R5559 VDD.n2593 VDD.n749 10.6151
R5560 VDD.n2594 VDD.n2593 10.6151
R5561 VDD.n2595 VDD.n2594 10.6151
R5562 VDD.n2190 VDD.n2189 10.6151
R5563 VDD.n2189 VDD.n2188 10.6151
R5564 VDD.n2188 VDD.n2187 10.6151
R5565 VDD.n2187 VDD.n2185 10.6151
R5566 VDD.n2185 VDD.n2182 10.6151
R5567 VDD.n2182 VDD.n2181 10.6151
R5568 VDD.n2181 VDD.n2178 10.6151
R5569 VDD.n2178 VDD.n2177 10.6151
R5570 VDD.n2177 VDD.n2174 10.6151
R5571 VDD.n2174 VDD.n2173 10.6151
R5572 VDD.n2173 VDD.n2170 10.6151
R5573 VDD.n1136 VDD.n1133 10.6151
R5574 VDD.n1133 VDD.n1132 10.6151
R5575 VDD.n1132 VDD.n1129 10.6151
R5576 VDD.n1129 VDD.n1128 10.6151
R5577 VDD.n1128 VDD.n1125 10.6151
R5578 VDD.n1125 VDD.n1124 10.6151
R5579 VDD.n1124 VDD.n1121 10.6151
R5580 VDD.n1121 VDD.n1120 10.6151
R5581 VDD.n1117 VDD.n1116 10.6151
R5582 VDD.n1116 VDD.n1114 10.6151
R5583 VDD.n3037 VDD.n3035 10.6151
R5584 VDD.n3035 VDD.n3034 10.6151
R5585 VDD.n3034 VDD.n3032 10.6151
R5586 VDD.n3032 VDD.n3031 10.6151
R5587 VDD.n3031 VDD.n3029 10.6151
R5588 VDD.n3029 VDD.n3028 10.6151
R5589 VDD.n3028 VDD.n2847 10.6151
R5590 VDD.n2847 VDD.n2846 10.6151
R5591 VDD.n2846 VDD.n2844 10.6151
R5592 VDD.n2844 VDD.n2843 10.6151
R5593 VDD.n2843 VDD.n2841 10.6151
R5594 VDD.n2841 VDD.n2840 10.6151
R5595 VDD.n2840 VDD.n2838 10.6151
R5596 VDD.n2838 VDD.n2837 10.6151
R5597 VDD.n2837 VDD.n2835 10.6151
R5598 VDD.n2835 VDD.n2834 10.6151
R5599 VDD.n2834 VDD.n2832 10.6151
R5600 VDD.n2832 VDD.n2831 10.6151
R5601 VDD.n2831 VDD.n2829 10.6151
R5602 VDD.n2829 VDD.n2828 10.6151
R5603 VDD.n2828 VDD.n2826 10.6151
R5604 VDD.n2826 VDD.n2825 10.6151
R5605 VDD.n2825 VDD.n2823 10.6151
R5606 VDD.n2823 VDD.n2822 10.6151
R5607 VDD.n2822 VDD.n2820 10.6151
R5608 VDD.n2820 VDD.n2819 10.6151
R5609 VDD.n2819 VDD.n2817 10.6151
R5610 VDD.n2817 VDD.n2816 10.6151
R5611 VDD.n2816 VDD.n2814 10.6151
R5612 VDD.n2814 VDD.n2813 10.6151
R5613 VDD.n2813 VDD.n2811 10.6151
R5614 VDD.n2811 VDD.n2810 10.6151
R5615 VDD.n2810 VDD.n2808 10.6151
R5616 VDD.n2808 VDD.n2807 10.6151
R5617 VDD.n2807 VDD.n2805 10.6151
R5618 VDD.n2805 VDD.n2804 10.6151
R5619 VDD.n2804 VDD.n2802 10.6151
R5620 VDD.n2802 VDD.n2801 10.6151
R5621 VDD.n2801 VDD.n2799 10.6151
R5622 VDD.n2799 VDD.n2798 10.6151
R5623 VDD.n2798 VDD.n2796 10.6151
R5624 VDD.n2796 VDD.n2795 10.6151
R5625 VDD.n2795 VDD.n2793 10.6151
R5626 VDD.n2793 VDD.n2792 10.6151
R5627 VDD.n2792 VDD.n2790 10.6151
R5628 VDD.n2790 VDD.n2789 10.6151
R5629 VDD.n2789 VDD.n2787 10.6151
R5630 VDD.n2787 VDD.n2786 10.6151
R5631 VDD.n2786 VDD.n2784 10.6151
R5632 VDD.n2784 VDD.n2783 10.6151
R5633 VDD.n2783 VDD.n2781 10.6151
R5634 VDD.n2781 VDD.n2780 10.6151
R5635 VDD.n2780 VDD.n2778 10.6151
R5636 VDD.n2778 VDD.n2777 10.6151
R5637 VDD.n2777 VDD.n2775 10.6151
R5638 VDD.n2775 VDD.n2774 10.6151
R5639 VDD.n2774 VDD.n2772 10.6151
R5640 VDD.n2772 VDD.n2771 10.6151
R5641 VDD.n2771 VDD.n2769 10.6151
R5642 VDD.n2769 VDD.n2768 10.6151
R5643 VDD.n2768 VDD.n2766 10.6151
R5644 VDD.n2766 VDD.n2765 10.6151
R5645 VDD.n2765 VDD.n2763 10.6151
R5646 VDD.n2763 VDD.n2762 10.6151
R5647 VDD.n2762 VDD.n2760 10.6151
R5648 VDD.n2760 VDD.n2759 10.6151
R5649 VDD.n2759 VDD.n2757 10.6151
R5650 VDD.n2757 VDD.n2756 10.6151
R5651 VDD.n2756 VDD.n2754 10.6151
R5652 VDD.n2754 VDD.n2753 10.6151
R5653 VDD.n2753 VDD.n2751 10.6151
R5654 VDD.n2751 VDD.n2750 10.6151
R5655 VDD.n2750 VDD.n2748 10.6151
R5656 VDD.n2748 VDD.n2747 10.6151
R5657 VDD.n2747 VDD.n2745 10.6151
R5658 VDD.n2745 VDD.n2744 10.6151
R5659 VDD.n2744 VDD.n2742 10.6151
R5660 VDD.n2742 VDD.n2741 10.6151
R5661 VDD.n2741 VDD.n2739 10.6151
R5662 VDD.n2739 VDD.n2738 10.6151
R5663 VDD.n2738 VDD.n2736 10.6151
R5664 VDD.n2736 VDD.n2735 10.6151
R5665 VDD.n2735 VDD.n2733 10.6151
R5666 VDD.n2733 VDD.n2732 10.6151
R5667 VDD.n2732 VDD.n2730 10.6151
R5668 VDD.n2730 VDD.n2729 10.6151
R5669 VDD.n2729 VDD.n2727 10.6151
R5670 VDD.n2727 VDD.n411 10.6151
R5671 VDD.n3436 VDD.n411 10.6151
R5672 VDD.n3437 VDD.n3436 10.6151
R5673 VDD.n3083 VDD.n706 10.6151
R5674 VDD.n3078 VDD.n706 10.6151
R5675 VDD.n3078 VDD.n3077 10.6151
R5676 VDD.n3077 VDD.n3076 10.6151
R5677 VDD.n3076 VDD.n3073 10.6151
R5678 VDD.n3073 VDD.n3072 10.6151
R5679 VDD.n3072 VDD.n3069 10.6151
R5680 VDD.n3069 VDD.n3068 10.6151
R5681 VDD.n3068 VDD.n3065 10.6151
R5682 VDD.n3065 VDD.n3064 10.6151
R5683 VDD.n3064 VDD.n3061 10.6151
R5684 VDD.n3061 VDD.n3060 10.6151
R5685 VDD.n3060 VDD.n3057 10.6151
R5686 VDD.n3057 VDD.n3056 10.6151
R5687 VDD.n3056 VDD.n3053 10.6151
R5688 VDD.n3053 VDD.n3052 10.6151
R5689 VDD.n3052 VDD.n3049 10.6151
R5690 VDD.n3049 VDD.n3048 10.6151
R5691 VDD.n3048 VDD.n3045 10.6151
R5692 VDD.n3045 VDD.n3044 10.6151
R5693 VDD.n3041 VDD.n3040 10.6151
R5694 VDD.n3040 VDD.n3038 10.6151
R5695 VDD.n3085 VDD.n3084 10.6151
R5696 VDD.n3085 VDD.n694 10.6151
R5697 VDD.n3095 VDD.n694 10.6151
R5698 VDD.n3096 VDD.n3095 10.6151
R5699 VDD.n3097 VDD.n3096 10.6151
R5700 VDD.n3097 VDD.n683 10.6151
R5701 VDD.n3107 VDD.n683 10.6151
R5702 VDD.n3108 VDD.n3107 10.6151
R5703 VDD.n3109 VDD.n3108 10.6151
R5704 VDD.n3109 VDD.n671 10.6151
R5705 VDD.n3119 VDD.n671 10.6151
R5706 VDD.n3120 VDD.n3119 10.6151
R5707 VDD.n3121 VDD.n3120 10.6151
R5708 VDD.n3121 VDD.n658 10.6151
R5709 VDD.n3131 VDD.n658 10.6151
R5710 VDD.n3132 VDD.n3131 10.6151
R5711 VDD.n3133 VDD.n3132 10.6151
R5712 VDD.n3133 VDD.n647 10.6151
R5713 VDD.n3143 VDD.n647 10.6151
R5714 VDD.n3144 VDD.n3143 10.6151
R5715 VDD.n3145 VDD.n3144 10.6151
R5716 VDD.n3145 VDD.n635 10.6151
R5717 VDD.n3155 VDD.n635 10.6151
R5718 VDD.n3156 VDD.n3155 10.6151
R5719 VDD.n3157 VDD.n3156 10.6151
R5720 VDD.n3157 VDD.n622 10.6151
R5721 VDD.n3167 VDD.n622 10.6151
R5722 VDD.n3168 VDD.n3167 10.6151
R5723 VDD.n3169 VDD.n3168 10.6151
R5724 VDD.n3169 VDD.n611 10.6151
R5725 VDD.n3179 VDD.n611 10.6151
R5726 VDD.n3180 VDD.n3179 10.6151
R5727 VDD.n3181 VDD.n3180 10.6151
R5728 VDD.n3181 VDD.n599 10.6151
R5729 VDD.n3191 VDD.n599 10.6151
R5730 VDD.n3192 VDD.n3191 10.6151
R5731 VDD.n3193 VDD.n3192 10.6151
R5732 VDD.n3193 VDD.n586 10.6151
R5733 VDD.n3203 VDD.n586 10.6151
R5734 VDD.n3204 VDD.n3203 10.6151
R5735 VDD.n3205 VDD.n3204 10.6151
R5736 VDD.n3205 VDD.n575 10.6151
R5737 VDD.n3215 VDD.n575 10.6151
R5738 VDD.n3216 VDD.n3215 10.6151
R5739 VDD.n3217 VDD.n3216 10.6151
R5740 VDD.n3217 VDD.n563 10.6151
R5741 VDD.n3226 VDD.n563 10.6151
R5742 VDD.n3227 VDD.n3226 10.6151
R5743 VDD.n3228 VDD.n3227 10.6151
R5744 VDD.n3228 VDD.n551 10.6151
R5745 VDD.n3238 VDD.n551 10.6151
R5746 VDD.n3239 VDD.n3238 10.6151
R5747 VDD.n3240 VDD.n3239 10.6151
R5748 VDD.n3240 VDD.n538 10.6151
R5749 VDD.n3250 VDD.n538 10.6151
R5750 VDD.n3251 VDD.n3250 10.6151
R5751 VDD.n3252 VDD.n3251 10.6151
R5752 VDD.n3252 VDD.n527 10.6151
R5753 VDD.n3262 VDD.n527 10.6151
R5754 VDD.n3263 VDD.n3262 10.6151
R5755 VDD.n3264 VDD.n3263 10.6151
R5756 VDD.n3264 VDD.n515 10.6151
R5757 VDD.n3274 VDD.n515 10.6151
R5758 VDD.n3275 VDD.n3274 10.6151
R5759 VDD.n3276 VDD.n3275 10.6151
R5760 VDD.n3276 VDD.n502 10.6151
R5761 VDD.n3286 VDD.n502 10.6151
R5762 VDD.n3287 VDD.n3286 10.6151
R5763 VDD.n3288 VDD.n3287 10.6151
R5764 VDD.n3288 VDD.n491 10.6151
R5765 VDD.n3298 VDD.n491 10.6151
R5766 VDD.n3299 VDD.n3298 10.6151
R5767 VDD.n3300 VDD.n3299 10.6151
R5768 VDD.n3300 VDD.n479 10.6151
R5769 VDD.n3310 VDD.n479 10.6151
R5770 VDD.n3311 VDD.n3310 10.6151
R5771 VDD.n3312 VDD.n3311 10.6151
R5772 VDD.n3312 VDD.n467 10.6151
R5773 VDD.n3322 VDD.n467 10.6151
R5774 VDD.n3323 VDD.n3322 10.6151
R5775 VDD.n3324 VDD.n3323 10.6151
R5776 VDD.n3324 VDD.n454 10.6151
R5777 VDD.n3336 VDD.n454 10.6151
R5778 VDD.n3337 VDD.n3336 10.6151
R5779 VDD.n3338 VDD.n3337 10.6151
R5780 VDD.n3338 VDD.n419 10.6151
R5781 VDD.n3401 VDD.n419 10.6151
R5782 VDD.n3402 VDD.n3401 10.6151
R5783 VDD.n3432 VDD.n3402 10.6151
R5784 VDD.n3432 VDD.n3431 10.6151
R5785 VDD.n3430 VDD.n3403 10.6151
R5786 VDD.n3404 VDD.n3403 10.6151
R5787 VDD.n3423 VDD.n3404 10.6151
R5788 VDD.n3423 VDD.n3422 10.6151
R5789 VDD.n3422 VDD.n3421 10.6151
R5790 VDD.n3421 VDD.n3406 10.6151
R5791 VDD.n3416 VDD.n3406 10.6151
R5792 VDD.n3416 VDD.n3415 10.6151
R5793 VDD.n3415 VDD.n3414 10.6151
R5794 VDD.n3414 VDD.n3409 10.6151
R5795 VDD.n3409 VDD.n397 10.6151
R5796 VDD.n3460 VDD.n398 10.6151
R5797 VDD.n401 VDD.n398 10.6151
R5798 VDD.n3453 VDD.n401 10.6151
R5799 VDD.n3453 VDD.n3452 10.6151
R5800 VDD.n3452 VDD.n3451 10.6151
R5801 VDD.n3451 VDD.n403 10.6151
R5802 VDD.n3446 VDD.n403 10.6151
R5803 VDD.n3446 VDD.n3445 10.6151
R5804 VDD.n3443 VDD.n408 10.6151
R5805 VDD.n3438 VDD.n408 10.6151
R5806 VDD.n3389 VDD.n427 10.6151
R5807 VDD.n3389 VDD.n3388 10.6151
R5808 VDD.n3388 VDD.n3387 10.6151
R5809 VDD.n3387 VDD.n429 10.6151
R5810 VDD.n3382 VDD.n429 10.6151
R5811 VDD.n3382 VDD.n3381 10.6151
R5812 VDD.n3381 VDD.n3380 10.6151
R5813 VDD.n3380 VDD.n432 10.6151
R5814 VDD.n3375 VDD.n432 10.6151
R5815 VDD.n3375 VDD.n3374 10.6151
R5816 VDD.n3374 VDD.n3373 10.6151
R5817 VDD.n3368 VDD.n437 10.6151
R5818 VDD.n3368 VDD.n3367 10.6151
R5819 VDD.n3367 VDD.n3366 10.6151
R5820 VDD.n3366 VDD.n439 10.6151
R5821 VDD.n3361 VDD.n439 10.6151
R5822 VDD.n3361 VDD.n3360 10.6151
R5823 VDD.n3360 VDD.n3359 10.6151
R5824 VDD.n3359 VDD.n442 10.6151
R5825 VDD.n3354 VDD.n3353 10.6151
R5826 VDD.n3353 VDD.n3352 10.6151
R5827 VDD.n2901 VDD.n2900 10.6151
R5828 VDD.n2903 VDD.n2901 10.6151
R5829 VDD.n2904 VDD.n2903 10.6151
R5830 VDD.n2906 VDD.n2904 10.6151
R5831 VDD.n2907 VDD.n2906 10.6151
R5832 VDD.n3024 VDD.n2907 10.6151
R5833 VDD.n3024 VDD.n3023 10.6151
R5834 VDD.n3023 VDD.n3022 10.6151
R5835 VDD.n3022 VDD.n3020 10.6151
R5836 VDD.n3020 VDD.n3019 10.6151
R5837 VDD.n3019 VDD.n3017 10.6151
R5838 VDD.n3017 VDD.n3016 10.6151
R5839 VDD.n3016 VDD.n3014 10.6151
R5840 VDD.n3014 VDD.n3013 10.6151
R5841 VDD.n3013 VDD.n3011 10.6151
R5842 VDD.n3011 VDD.n3010 10.6151
R5843 VDD.n3010 VDD.n3008 10.6151
R5844 VDD.n3008 VDD.n3007 10.6151
R5845 VDD.n3007 VDD.n3005 10.6151
R5846 VDD.n3005 VDD.n3004 10.6151
R5847 VDD.n3004 VDD.n3002 10.6151
R5848 VDD.n3002 VDD.n3001 10.6151
R5849 VDD.n3001 VDD.n2999 10.6151
R5850 VDD.n2999 VDD.n2998 10.6151
R5851 VDD.n2998 VDD.n2996 10.6151
R5852 VDD.n2996 VDD.n2995 10.6151
R5853 VDD.n2995 VDD.n2993 10.6151
R5854 VDD.n2993 VDD.n2992 10.6151
R5855 VDD.n2992 VDD.n2990 10.6151
R5856 VDD.n2990 VDD.n2989 10.6151
R5857 VDD.n2989 VDD.n2987 10.6151
R5858 VDD.n2987 VDD.n2986 10.6151
R5859 VDD.n2986 VDD.n2984 10.6151
R5860 VDD.n2984 VDD.n2983 10.6151
R5861 VDD.n2983 VDD.n2981 10.6151
R5862 VDD.n2981 VDD.n2980 10.6151
R5863 VDD.n2980 VDD.n2978 10.6151
R5864 VDD.n2978 VDD.n2977 10.6151
R5865 VDD.n2977 VDD.n2975 10.6151
R5866 VDD.n2975 VDD.n2974 10.6151
R5867 VDD.n2974 VDD.n2972 10.6151
R5868 VDD.n2972 VDD.n2971 10.6151
R5869 VDD.n2971 VDD.n2969 10.6151
R5870 VDD.n2969 VDD.n2968 10.6151
R5871 VDD.n2968 VDD.n2966 10.6151
R5872 VDD.n2966 VDD.n2965 10.6151
R5873 VDD.n2965 VDD.n2963 10.6151
R5874 VDD.n2963 VDD.n2962 10.6151
R5875 VDD.n2962 VDD.n2960 10.6151
R5876 VDD.n2960 VDD.n2959 10.6151
R5877 VDD.n2959 VDD.n2957 10.6151
R5878 VDD.n2957 VDD.n2956 10.6151
R5879 VDD.n2956 VDD.n2954 10.6151
R5880 VDD.n2954 VDD.n2953 10.6151
R5881 VDD.n2953 VDD.n2951 10.6151
R5882 VDD.n2951 VDD.n2950 10.6151
R5883 VDD.n2950 VDD.n2948 10.6151
R5884 VDD.n2948 VDD.n2947 10.6151
R5885 VDD.n2947 VDD.n2945 10.6151
R5886 VDD.n2945 VDD.n2944 10.6151
R5887 VDD.n2944 VDD.n2942 10.6151
R5888 VDD.n2942 VDD.n2941 10.6151
R5889 VDD.n2941 VDD.n2939 10.6151
R5890 VDD.n2939 VDD.n2938 10.6151
R5891 VDD.n2938 VDD.n2936 10.6151
R5892 VDD.n2936 VDD.n2935 10.6151
R5893 VDD.n2935 VDD.n2933 10.6151
R5894 VDD.n2933 VDD.n2932 10.6151
R5895 VDD.n2932 VDD.n2930 10.6151
R5896 VDD.n2930 VDD.n2929 10.6151
R5897 VDD.n2929 VDD.n2927 10.6151
R5898 VDD.n2927 VDD.n2926 10.6151
R5899 VDD.n2926 VDD.n2924 10.6151
R5900 VDD.n2924 VDD.n2923 10.6151
R5901 VDD.n2923 VDD.n2921 10.6151
R5902 VDD.n2921 VDD.n2920 10.6151
R5903 VDD.n2920 VDD.n2918 10.6151
R5904 VDD.n2918 VDD.n2917 10.6151
R5905 VDD.n2917 VDD.n2915 10.6151
R5906 VDD.n2915 VDD.n2914 10.6151
R5907 VDD.n2914 VDD.n2912 10.6151
R5908 VDD.n2912 VDD.n2911 10.6151
R5909 VDD.n2911 VDD.n2909 10.6151
R5910 VDD.n2909 VDD.n2908 10.6151
R5911 VDD.n2908 VDD.n448 10.6151
R5912 VDD.n3343 VDD.n448 10.6151
R5913 VDD.n3344 VDD.n3343 10.6151
R5914 VDD.n3346 VDD.n3344 10.6151
R5915 VDD.n3347 VDD.n3346 10.6151
R5916 VDD.n3348 VDD.n3347 10.6151
R5917 VDD.n2852 VDD.n2851 10.6151
R5918 VDD.n2855 VDD.n2852 10.6151
R5919 VDD.n2856 VDD.n2855 10.6151
R5920 VDD.n2859 VDD.n2856 10.6151
R5921 VDD.n2860 VDD.n2859 10.6151
R5922 VDD.n2863 VDD.n2860 10.6151
R5923 VDD.n2864 VDD.n2863 10.6151
R5924 VDD.n2867 VDD.n2864 10.6151
R5925 VDD.n2868 VDD.n2867 10.6151
R5926 VDD.n2871 VDD.n2868 10.6151
R5927 VDD.n2872 VDD.n2871 10.6151
R5928 VDD.n2875 VDD.n2872 10.6151
R5929 VDD.n2876 VDD.n2875 10.6151
R5930 VDD.n2879 VDD.n2876 10.6151
R5931 VDD.n2880 VDD.n2879 10.6151
R5932 VDD.n2883 VDD.n2880 10.6151
R5933 VDD.n2884 VDD.n2883 10.6151
R5934 VDD.n2887 VDD.n2884 10.6151
R5935 VDD.n2888 VDD.n2887 10.6151
R5936 VDD.n2891 VDD.n2888 10.6151
R5937 VDD.n2896 VDD.n2893 10.6151
R5938 VDD.n2897 VDD.n2896 10.6151
R5939 VDD.n3089 VDD.n700 10.6151
R5940 VDD.n3090 VDD.n3089 10.6151
R5941 VDD.n3091 VDD.n3090 10.6151
R5942 VDD.n3091 VDD.n688 10.6151
R5943 VDD.n3101 VDD.n688 10.6151
R5944 VDD.n3102 VDD.n3101 10.6151
R5945 VDD.n3103 VDD.n3102 10.6151
R5946 VDD.n3103 VDD.n677 10.6151
R5947 VDD.n3113 VDD.n677 10.6151
R5948 VDD.n3114 VDD.n3113 10.6151
R5949 VDD.n3115 VDD.n3114 10.6151
R5950 VDD.n3115 VDD.n665 10.6151
R5951 VDD.n3125 VDD.n665 10.6151
R5952 VDD.n3126 VDD.n3125 10.6151
R5953 VDD.n3127 VDD.n3126 10.6151
R5954 VDD.n3127 VDD.n653 10.6151
R5955 VDD.n3137 VDD.n653 10.6151
R5956 VDD.n3138 VDD.n3137 10.6151
R5957 VDD.n3139 VDD.n3138 10.6151
R5958 VDD.n3139 VDD.n641 10.6151
R5959 VDD.n3149 VDD.n641 10.6151
R5960 VDD.n3150 VDD.n3149 10.6151
R5961 VDD.n3151 VDD.n3150 10.6151
R5962 VDD.n3151 VDD.n629 10.6151
R5963 VDD.n3161 VDD.n629 10.6151
R5964 VDD.n3162 VDD.n3161 10.6151
R5965 VDD.n3163 VDD.n3162 10.6151
R5966 VDD.n3163 VDD.n617 10.6151
R5967 VDD.n3173 VDD.n617 10.6151
R5968 VDD.n3174 VDD.n3173 10.6151
R5969 VDD.n3175 VDD.n3174 10.6151
R5970 VDD.n3175 VDD.n605 10.6151
R5971 VDD.n3185 VDD.n605 10.6151
R5972 VDD.n3186 VDD.n3185 10.6151
R5973 VDD.n3187 VDD.n3186 10.6151
R5974 VDD.n3187 VDD.n593 10.6151
R5975 VDD.n3197 VDD.n593 10.6151
R5976 VDD.n3198 VDD.n3197 10.6151
R5977 VDD.n3199 VDD.n3198 10.6151
R5978 VDD.n3199 VDD.n581 10.6151
R5979 VDD.n3209 VDD.n581 10.6151
R5980 VDD.n3210 VDD.n3209 10.6151
R5981 VDD.n3211 VDD.n3210 10.6151
R5982 VDD.n3211 VDD.n569 10.6151
R5983 VDD.n3220 VDD.n569 10.6151
R5984 VDD.n3221 VDD.n3220 10.6151
R5985 VDD.n3222 VDD.n3221 10.6151
R5986 VDD.n3222 VDD.n557 10.6151
R5987 VDD.n3232 VDD.n557 10.6151
R5988 VDD.n3233 VDD.n3232 10.6151
R5989 VDD.n3234 VDD.n3233 10.6151
R5990 VDD.n3234 VDD.n545 10.6151
R5991 VDD.n3244 VDD.n545 10.6151
R5992 VDD.n3245 VDD.n3244 10.6151
R5993 VDD.n3246 VDD.n3245 10.6151
R5994 VDD.n3246 VDD.n533 10.6151
R5995 VDD.n3256 VDD.n533 10.6151
R5996 VDD.n3257 VDD.n3256 10.6151
R5997 VDD.n3258 VDD.n3257 10.6151
R5998 VDD.n3258 VDD.n521 10.6151
R5999 VDD.n3268 VDD.n521 10.6151
R6000 VDD.n3269 VDD.n3268 10.6151
R6001 VDD.n3270 VDD.n3269 10.6151
R6002 VDD.n3270 VDD.n509 10.6151
R6003 VDD.n3280 VDD.n509 10.6151
R6004 VDD.n3281 VDD.n3280 10.6151
R6005 VDD.n3282 VDD.n3281 10.6151
R6006 VDD.n3282 VDD.n497 10.6151
R6007 VDD.n3292 VDD.n497 10.6151
R6008 VDD.n3293 VDD.n3292 10.6151
R6009 VDD.n3294 VDD.n3293 10.6151
R6010 VDD.n3294 VDD.n485 10.6151
R6011 VDD.n3304 VDD.n485 10.6151
R6012 VDD.n3305 VDD.n3304 10.6151
R6013 VDD.n3306 VDD.n3305 10.6151
R6014 VDD.n3306 VDD.n473 10.6151
R6015 VDD.n3316 VDD.n473 10.6151
R6016 VDD.n3317 VDD.n3316 10.6151
R6017 VDD.n3318 VDD.n3317 10.6151
R6018 VDD.n3318 VDD.n461 10.6151
R6019 VDD.n3328 VDD.n461 10.6151
R6020 VDD.n3329 VDD.n3328 10.6151
R6021 VDD.n3332 VDD.n3329 10.6151
R6022 VDD.n3332 VDD.n3331 10.6151
R6023 VDD.n3331 VDD.n3330 10.6151
R6024 VDD.n3330 VDD.n426 10.6151
R6025 VDD.n3397 VDD.n426 10.6151
R6026 VDD.n3397 VDD.n3396 10.6151
R6027 VDD.n3396 VDD.n3395 10.6151
R6028 VDD.n3395 VDD.n3394 10.6151
R6029 VDD.n2197 VDD.n2196 10.6151
R6030 VDD.n2197 VDD.n1006 10.6151
R6031 VDD.n2207 VDD.n1006 10.6151
R6032 VDD.n2208 VDD.n2207 10.6151
R6033 VDD.n2209 VDD.n2208 10.6151
R6034 VDD.n2209 VDD.n993 10.6151
R6035 VDD.n2219 VDD.n993 10.6151
R6036 VDD.n2220 VDD.n2219 10.6151
R6037 VDD.n2221 VDD.n2220 10.6151
R6038 VDD.n2221 VDD.n982 10.6151
R6039 VDD.n2231 VDD.n982 10.6151
R6040 VDD.n2232 VDD.n2231 10.6151
R6041 VDD.n2233 VDD.n2232 10.6151
R6042 VDD.n2233 VDD.n970 10.6151
R6043 VDD.n2243 VDD.n970 10.6151
R6044 VDD.n2244 VDD.n2243 10.6151
R6045 VDD.n2245 VDD.n2244 10.6151
R6046 VDD.n2245 VDD.n957 10.6151
R6047 VDD.n2255 VDD.n957 10.6151
R6048 VDD.n2256 VDD.n2255 10.6151
R6049 VDD.n2257 VDD.n2256 10.6151
R6050 VDD.n2257 VDD.n946 10.6151
R6051 VDD.n2267 VDD.n946 10.6151
R6052 VDD.n2268 VDD.n2267 10.6151
R6053 VDD.n2269 VDD.n2268 10.6151
R6054 VDD.n2269 VDD.n934 10.6151
R6055 VDD.n2279 VDD.n934 10.6151
R6056 VDD.n2280 VDD.n2279 10.6151
R6057 VDD.n2281 VDD.n2280 10.6151
R6058 VDD.n2281 VDD.n921 10.6151
R6059 VDD.n2291 VDD.n921 10.6151
R6060 VDD.n2292 VDD.n2291 10.6151
R6061 VDD.n2293 VDD.n2292 10.6151
R6062 VDD.n2293 VDD.n910 10.6151
R6063 VDD.n2303 VDD.n910 10.6151
R6064 VDD.n2304 VDD.n2303 10.6151
R6065 VDD.n2305 VDD.n2304 10.6151
R6066 VDD.n2305 VDD.n898 10.6151
R6067 VDD.n2315 VDD.n898 10.6151
R6068 VDD.n2316 VDD.n2315 10.6151
R6069 VDD.n2322 VDD.n2316 10.6151
R6070 VDD.n2322 VDD.n2321 10.6151
R6071 VDD.n2321 VDD.n2320 10.6151
R6072 VDD.n2320 VDD.n2319 10.6151
R6073 VDD.n2319 VDD.n2317 10.6151
R6074 VDD.n2317 VDD.n869 10.6151
R6075 VDD.n2467 VDD.n869 10.6151
R6076 VDD.n2468 VDD.n2467 10.6151
R6077 VDD.n2469 VDD.n2468 10.6151
R6078 VDD.n2469 VDD.n857 10.6151
R6079 VDD.n2479 VDD.n857 10.6151
R6080 VDD.n2480 VDD.n2479 10.6151
R6081 VDD.n2481 VDD.n2480 10.6151
R6082 VDD.n2481 VDD.n844 10.6151
R6083 VDD.n2491 VDD.n844 10.6151
R6084 VDD.n2492 VDD.n2491 10.6151
R6085 VDD.n2493 VDD.n2492 10.6151
R6086 VDD.n2493 VDD.n833 10.6151
R6087 VDD.n2503 VDD.n833 10.6151
R6088 VDD.n2504 VDD.n2503 10.6151
R6089 VDD.n2505 VDD.n2504 10.6151
R6090 VDD.n2505 VDD.n821 10.6151
R6091 VDD.n2515 VDD.n821 10.6151
R6092 VDD.n2516 VDD.n2515 10.6151
R6093 VDD.n2517 VDD.n2516 10.6151
R6094 VDD.n2517 VDD.n808 10.6151
R6095 VDD.n2527 VDD.n808 10.6151
R6096 VDD.n2528 VDD.n2527 10.6151
R6097 VDD.n2529 VDD.n2528 10.6151
R6098 VDD.n2529 VDD.n797 10.6151
R6099 VDD.n2539 VDD.n797 10.6151
R6100 VDD.n2540 VDD.n2539 10.6151
R6101 VDD.n2541 VDD.n2540 10.6151
R6102 VDD.n2541 VDD.n785 10.6151
R6103 VDD.n2551 VDD.n785 10.6151
R6104 VDD.n2552 VDD.n2551 10.6151
R6105 VDD.n2553 VDD.n2552 10.6151
R6106 VDD.n2553 VDD.n773 10.6151
R6107 VDD.n2563 VDD.n773 10.6151
R6108 VDD.n2564 VDD.n2563 10.6151
R6109 VDD.n2565 VDD.n2564 10.6151
R6110 VDD.n2565 VDD.n761 10.6151
R6111 VDD.n2575 VDD.n761 10.6151
R6112 VDD.n2576 VDD.n2575 10.6151
R6113 VDD.n2582 VDD.n2576 10.6151
R6114 VDD.n2582 VDD.n2581 10.6151
R6115 VDD.n2581 VDD.n2580 10.6151
R6116 VDD.n2580 VDD.n2579 10.6151
R6117 VDD.n2579 VDD.n2577 10.6151
R6118 VDD.n2577 VDD.n735 10.6151
R6119 VDD.n2697 VDD.n2696 10.6151
R6120 VDD.n2696 VDD.n2695 10.6151
R6121 VDD.n2695 VDD.n2692 10.6151
R6122 VDD.n2692 VDD.n2691 10.6151
R6123 VDD.n2691 VDD.n2688 10.6151
R6124 VDD.n2688 VDD.n2687 10.6151
R6125 VDD.n2687 VDD.n2684 10.6151
R6126 VDD.n2684 VDD.n2683 10.6151
R6127 VDD.n2683 VDD.n2680 10.6151
R6128 VDD.n2680 VDD.n2679 10.6151
R6129 VDD.n2679 VDD.n2676 10.6151
R6130 VDD.n2676 VDD.n2675 10.6151
R6131 VDD.n2675 VDD.n2672 10.6151
R6132 VDD.n2672 VDD.n2671 10.6151
R6133 VDD.n2671 VDD.n2668 10.6151
R6134 VDD.n2668 VDD.n2667 10.6151
R6135 VDD.n2667 VDD.n2664 10.6151
R6136 VDD.n2664 VDD.n2663 10.6151
R6137 VDD.n2663 VDD.n2660 10.6151
R6138 VDD.n2660 VDD.n2659 10.6151
R6139 VDD.n2656 VDD.n2655 10.6151
R6140 VDD.n2655 VDD.n2653 10.6151
R6141 VDD.n2055 VDD.n2053 10.6151
R6142 VDD.n2053 VDD.n2052 10.6151
R6143 VDD.n2052 VDD.n2050 10.6151
R6144 VDD.n2050 VDD.n2049 10.6151
R6145 VDD.n2049 VDD.n2047 10.6151
R6146 VDD.n2047 VDD.n2046 10.6151
R6147 VDD.n2046 VDD.n2044 10.6151
R6148 VDD.n2044 VDD.n2043 10.6151
R6149 VDD.n2043 VDD.n2041 10.6151
R6150 VDD.n2041 VDD.n2040 10.6151
R6151 VDD.n2040 VDD.n2038 10.6151
R6152 VDD.n2038 VDD.n2037 10.6151
R6153 VDD.n2037 VDD.n2035 10.6151
R6154 VDD.n2035 VDD.n2034 10.6151
R6155 VDD.n2034 VDD.n2032 10.6151
R6156 VDD.n2032 VDD.n2031 10.6151
R6157 VDD.n2031 VDD.n2029 10.6151
R6158 VDD.n2029 VDD.n2028 10.6151
R6159 VDD.n2028 VDD.n2026 10.6151
R6160 VDD.n2026 VDD.n2025 10.6151
R6161 VDD.n2025 VDD.n2023 10.6151
R6162 VDD.n2023 VDD.n2022 10.6151
R6163 VDD.n2022 VDD.n2020 10.6151
R6164 VDD.n2020 VDD.n2019 10.6151
R6165 VDD.n2019 VDD.n2017 10.6151
R6166 VDD.n2017 VDD.n2016 10.6151
R6167 VDD.n2016 VDD.n2014 10.6151
R6168 VDD.n2014 VDD.n2013 10.6151
R6169 VDD.n2013 VDD.n2011 10.6151
R6170 VDD.n2011 VDD.n2010 10.6151
R6171 VDD.n2010 VDD.n2008 10.6151
R6172 VDD.n2008 VDD.n2007 10.6151
R6173 VDD.n2007 VDD.n2005 10.6151
R6174 VDD.n2005 VDD.n2004 10.6151
R6175 VDD.n2004 VDD.n2002 10.6151
R6176 VDD.n2002 VDD.n2001 10.6151
R6177 VDD.n2001 VDD.n1999 10.6151
R6178 VDD.n1999 VDD.n1998 10.6151
R6179 VDD.n1998 VDD.n1996 10.6151
R6180 VDD.n1996 VDD.n1995 10.6151
R6181 VDD.n1995 VDD.n1993 10.6151
R6182 VDD.n1993 VDD.n1992 10.6151
R6183 VDD.n1992 VDD.n885 10.6151
R6184 VDD.n2333 VDD.n885 10.6151
R6185 VDD.n2334 VDD.n2333 10.6151
R6186 VDD.n2336 VDD.n2334 10.6151
R6187 VDD.n2337 VDD.n2336 10.6151
R6188 VDD.n2339 VDD.n2337 10.6151
R6189 VDD.n2340 VDD.n2339 10.6151
R6190 VDD.n2342 VDD.n2340 10.6151
R6191 VDD.n2343 VDD.n2342 10.6151
R6192 VDD.n2345 VDD.n2343 10.6151
R6193 VDD.n2346 VDD.n2345 10.6151
R6194 VDD.n2348 VDD.n2346 10.6151
R6195 VDD.n2349 VDD.n2348 10.6151
R6196 VDD.n2351 VDD.n2349 10.6151
R6197 VDD.n2352 VDD.n2351 10.6151
R6198 VDD.n2354 VDD.n2352 10.6151
R6199 VDD.n2355 VDD.n2354 10.6151
R6200 VDD.n2357 VDD.n2355 10.6151
R6201 VDD.n2358 VDD.n2357 10.6151
R6202 VDD.n2360 VDD.n2358 10.6151
R6203 VDD.n2361 VDD.n2360 10.6151
R6204 VDD.n2363 VDD.n2361 10.6151
R6205 VDD.n2364 VDD.n2363 10.6151
R6206 VDD.n2366 VDD.n2364 10.6151
R6207 VDD.n2367 VDD.n2366 10.6151
R6208 VDD.n2369 VDD.n2367 10.6151
R6209 VDD.n2370 VDD.n2369 10.6151
R6210 VDD.n2372 VDD.n2370 10.6151
R6211 VDD.n2373 VDD.n2372 10.6151
R6212 VDD.n2375 VDD.n2373 10.6151
R6213 VDD.n2376 VDD.n2375 10.6151
R6214 VDD.n2378 VDD.n2376 10.6151
R6215 VDD.n2379 VDD.n2378 10.6151
R6216 VDD.n2381 VDD.n2379 10.6151
R6217 VDD.n2382 VDD.n2381 10.6151
R6218 VDD.n2384 VDD.n2382 10.6151
R6219 VDD.n2385 VDD.n2384 10.6151
R6220 VDD.n2387 VDD.n2385 10.6151
R6221 VDD.n2388 VDD.n2387 10.6151
R6222 VDD.n2390 VDD.n2388 10.6151
R6223 VDD.n2391 VDD.n2390 10.6151
R6224 VDD.n2397 VDD.n2391 10.6151
R6225 VDD.n2397 VDD.n2396 10.6151
R6226 VDD.n2396 VDD.n2395 10.6151
R6227 VDD.n2395 VDD.n2393 10.6151
R6228 VDD.n2393 VDD.n2392 10.6151
R6229 VDD.n2392 VDD.n739 10.6151
R6230 VDD.n2652 VDD.n739 10.6151
R6231 VDD.n2195 VDD.n1018 10.6151
R6232 VDD.n1969 VDD.n1018 10.6151
R6233 VDD.n1972 VDD.n1969 10.6151
R6234 VDD.n1973 VDD.n1972 10.6151
R6235 VDD.n1976 VDD.n1973 10.6151
R6236 VDD.n1977 VDD.n1976 10.6151
R6237 VDD.n1980 VDD.n1977 10.6151
R6238 VDD.n1981 VDD.n1980 10.6151
R6239 VDD.n1984 VDD.n1981 10.6151
R6240 VDD.n1985 VDD.n1984 10.6151
R6241 VDD.n1988 VDD.n1985 10.6151
R6242 VDD.n2078 VDD.n2075 10.6151
R6243 VDD.n2075 VDD.n2074 10.6151
R6244 VDD.n2074 VDD.n2071 10.6151
R6245 VDD.n2071 VDD.n2070 10.6151
R6246 VDD.n2070 VDD.n2067 10.6151
R6247 VDD.n2067 VDD.n2066 10.6151
R6248 VDD.n2066 VDD.n2063 10.6151
R6249 VDD.n2063 VDD.n2062 10.6151
R6250 VDD.n2059 VDD.n2058 10.6151
R6251 VDD.n2058 VDD.n2056 10.6151
R6252 VDD.n2169 VDD.n2168 10.391
R6253 VDD.n3604 VDD.n3461 10.391
R6254 VDD.n2199 VDD.n1014 10.2871
R6255 VDD.n2199 VDD.n1008 10.2871
R6256 VDD.n2205 VDD.n1008 10.2871
R6257 VDD.n2205 VDD.n1001 10.2871
R6258 VDD.n2211 VDD.n1001 10.2871
R6259 VDD.n2211 VDD.n1004 10.2871
R6260 VDD.n2217 VDD.n997 10.2871
R6261 VDD.n2223 VDD.n984 10.2871
R6262 VDD.n2229 VDD.n984 10.2871
R6263 VDD.n2229 VDD.n978 10.2871
R6264 VDD.n2235 VDD.n978 10.2871
R6265 VDD.n2235 VDD.n972 10.2871
R6266 VDD.n2241 VDD.n972 10.2871
R6267 VDD.n2241 VDD.n966 10.2871
R6268 VDD.n2247 VDD.n966 10.2871
R6269 VDD.n2247 VDD.n959 10.2871
R6270 VDD.n2253 VDD.n959 10.2871
R6271 VDD.n2253 VDD.n962 10.2871
R6272 VDD.n2265 VDD.n948 10.2871
R6273 VDD.n2265 VDD.n942 10.2871
R6274 VDD.n2271 VDD.n942 10.2871
R6275 VDD.n2271 VDD.n936 10.2871
R6276 VDD.n2277 VDD.n936 10.2871
R6277 VDD.n2277 VDD.n930 10.2871
R6278 VDD.n2283 VDD.n930 10.2871
R6279 VDD.n2283 VDD.n923 10.2871
R6280 VDD.n2289 VDD.n923 10.2871
R6281 VDD.n2289 VDD.n926 10.2871
R6282 VDD.n2301 VDD.n912 10.2871
R6283 VDD.n2301 VDD.n906 10.2871
R6284 VDD.n2307 VDD.n906 10.2871
R6285 VDD.n2307 VDD.n900 10.2871
R6286 VDD.n2313 VDD.n900 10.2871
R6287 VDD.n2313 VDD.n893 10.2871
R6288 VDD.n2324 VDD.n893 10.2871
R6289 VDD.n2324 VDD.n887 10.2871
R6290 VDD.n2330 VDD.n887 10.2871
R6291 VDD.n2330 VDD.n877 10.2871
R6292 VDD.t100 VDD.n877 10.2871
R6293 VDD.t100 VDD.n871 10.2871
R6294 VDD.n2465 VDD.n871 10.2871
R6295 VDD.n2465 VDD.n865 10.2871
R6296 VDD.n2471 VDD.n865 10.2871
R6297 VDD.n2477 VDD.n859 10.2871
R6298 VDD.n2477 VDD.n853 10.2871
R6299 VDD.n2483 VDD.n853 10.2871
R6300 VDD.n2483 VDD.n846 10.2871
R6301 VDD.n2489 VDD.n846 10.2871
R6302 VDD.n2489 VDD.n849 10.2871
R6303 VDD.n2495 VDD.n835 10.2871
R6304 VDD.n2501 VDD.n835 10.2871
R6305 VDD.n2501 VDD.n829 10.2871
R6306 VDD.n2507 VDD.n829 10.2871
R6307 VDD.n2513 VDD.n823 10.2871
R6308 VDD.n2513 VDD.n817 10.2871
R6309 VDD.n2519 VDD.n817 10.2871
R6310 VDD.n2519 VDD.n810 10.2871
R6311 VDD.n2525 VDD.n810 10.2871
R6312 VDD.n2525 VDD.n813 10.2871
R6313 VDD.n2531 VDD.n799 10.2871
R6314 VDD.n2537 VDD.n799 10.2871
R6315 VDD.n2537 VDD.n793 10.2871
R6316 VDD.n2543 VDD.n793 10.2871
R6317 VDD.n2549 VDD.n787 10.2871
R6318 VDD.n2549 VDD.n781 10.2871
R6319 VDD.n2555 VDD.n781 10.2871
R6320 VDD.n2555 VDD.n775 10.2871
R6321 VDD.n2561 VDD.n775 10.2871
R6322 VDD.n2561 VDD.n769 10.2871
R6323 VDD.n2567 VDD.n769 10.2871
R6324 VDD.n2567 VDD.n763 10.2871
R6325 VDD.n2573 VDD.n763 10.2871
R6326 VDD.n2584 VDD.n751 10.2871
R6327 VDD.n2590 VDD.n751 10.2871
R6328 VDD.n2590 VDD.n741 10.2871
R6329 VDD.n2649 VDD.n741 10.2871
R6330 VDD.n2649 VDD.n708 10.2871
R6331 VDD.n3087 VDD.n702 10.2871
R6332 VDD.n3087 VDD.n696 10.2871
R6333 VDD.n3093 VDD.n696 10.2871
R6334 VDD.n3093 VDD.n690 10.2871
R6335 VDD.n3099 VDD.n690 10.2871
R6336 VDD.n3105 VDD.n679 10.2871
R6337 VDD.n3111 VDD.n679 10.2871
R6338 VDD.n3111 VDD.n673 10.2871
R6339 VDD.n3117 VDD.n673 10.2871
R6340 VDD.n3117 VDD.n667 10.2871
R6341 VDD.n3123 VDD.n667 10.2871
R6342 VDD.n3123 VDD.n660 10.2871
R6343 VDD.n3129 VDD.n660 10.2871
R6344 VDD.n3129 VDD.n663 10.2871
R6345 VDD.n3135 VDD.n649 10.2871
R6346 VDD.n3141 VDD.n649 10.2871
R6347 VDD.n3141 VDD.n643 10.2871
R6348 VDD.n3147 VDD.n643 10.2871
R6349 VDD.n3153 VDD.n637 10.2871
R6350 VDD.n3153 VDD.n631 10.2871
R6351 VDD.n3159 VDD.n631 10.2871
R6352 VDD.n3159 VDD.n624 10.2871
R6353 VDD.n3165 VDD.n624 10.2871
R6354 VDD.n3165 VDD.n627 10.2871
R6355 VDD.n3171 VDD.n613 10.2871
R6356 VDD.n3177 VDD.n613 10.2871
R6357 VDD.n3177 VDD.n607 10.2871
R6358 VDD.n3183 VDD.n607 10.2871
R6359 VDD.n3189 VDD.n601 10.2871
R6360 VDD.n3189 VDD.n595 10.2871
R6361 VDD.n3195 VDD.n595 10.2871
R6362 VDD.n3195 VDD.n588 10.2871
R6363 VDD.n3201 VDD.n588 10.2871
R6364 VDD.n3201 VDD.n591 10.2871
R6365 VDD.n3207 VDD.n577 10.2871
R6366 VDD.n3213 VDD.n577 10.2871
R6367 VDD.n3213 VDD.n571 10.2871
R6368 VDD.t108 VDD.n571 10.2871
R6369 VDD.t108 VDD.n565 10.2871
R6370 VDD.n3224 VDD.n565 10.2871
R6371 VDD.n3224 VDD.n559 10.2871
R6372 VDD.n3230 VDD.n559 10.2871
R6373 VDD.n3230 VDD.n553 10.2871
R6374 VDD.n3236 VDD.n553 10.2871
R6375 VDD.n3236 VDD.n547 10.2871
R6376 VDD.n3242 VDD.n547 10.2871
R6377 VDD.n3242 VDD.n540 10.2871
R6378 VDD.n3248 VDD.n540 10.2871
R6379 VDD.n3248 VDD.n543 10.2871
R6380 VDD.n3260 VDD.n529 10.2871
R6381 VDD.n3260 VDD.n523 10.2871
R6382 VDD.n3266 VDD.n523 10.2871
R6383 VDD.n3266 VDD.n517 10.2871
R6384 VDD.n3272 VDD.n517 10.2871
R6385 VDD.n3272 VDD.n511 10.2871
R6386 VDD.n3278 VDD.n511 10.2871
R6387 VDD.n3278 VDD.n504 10.2871
R6388 VDD.n3284 VDD.n504 10.2871
R6389 VDD.n3284 VDD.n507 10.2871
R6390 VDD.n3296 VDD.n493 10.2871
R6391 VDD.n3296 VDD.n487 10.2871
R6392 VDD.n3302 VDD.n487 10.2871
R6393 VDD.n3302 VDD.n481 10.2871
R6394 VDD.n3308 VDD.n481 10.2871
R6395 VDD.n3308 VDD.n475 10.2871
R6396 VDD.n3314 VDD.n475 10.2871
R6397 VDD.n3314 VDD.n469 10.2871
R6398 VDD.n3320 VDD.n469 10.2871
R6399 VDD.n3320 VDD.n463 10.2871
R6400 VDD.n3326 VDD.n463 10.2871
R6401 VDD.n3334 VDD.n456 10.2871
R6402 VDD.n3340 VDD.n450 10.2871
R6403 VDD.n3340 VDD.n421 10.2871
R6404 VDD.n3399 VDD.n421 10.2871
R6405 VDD.n3399 VDD.n413 10.2871
R6406 VDD.n3434 VDD.n413 10.2871
R6407 VDD.n3434 VDD.n415 10.2871
R6408 VDD.n435 VDD.n392 10.0121
R6409 VDD.n2080 VDD.n2079 10.0121
R6410 VDD.n2193 VDD.t91 9.98458
R6411 VDD.n400 VDD.t114 9.98458
R6412 VDD.n2295 VDD.t102 9.53076
R6413 VDD.t93 VDD.n787 9.53076
R6414 VDD.n663 VDD.t109 9.53076
R6415 VDD.n3254 VDD.t84 9.53076
R6416 VDD.n1139 VDD.n1137 9.3005
R6417 VDD.n2162 VDD.n1162 9.3005
R6418 VDD.n2161 VDD.n1163 9.3005
R6419 VDD.n2160 VDD.n1164 9.3005
R6420 VDD.n2157 VDD.n1165 9.3005
R6421 VDD.n2156 VDD.n1166 9.3005
R6422 VDD.n2153 VDD.n2152 9.3005
R6423 VDD.n2151 VDD.n1167 9.3005
R6424 VDD.n2150 VDD.n2149 9.3005
R6425 VDD.n2146 VDD.n1170 9.3005
R6426 VDD.n2143 VDD.n1171 9.3005
R6427 VDD.n2142 VDD.n1172 9.3005
R6428 VDD.n2139 VDD.n1173 9.3005
R6429 VDD.n2138 VDD.n1174 9.3005
R6430 VDD.n2135 VDD.n1175 9.3005
R6431 VDD.n2134 VDD.n1176 9.3005
R6432 VDD.n2131 VDD.n1177 9.3005
R6433 VDD.n2127 VDD.n1178 9.3005
R6434 VDD.n2124 VDD.n1179 9.3005
R6435 VDD.n2123 VDD.n1180 9.3005
R6436 VDD.n2120 VDD.n1181 9.3005
R6437 VDD.n2119 VDD.n1182 9.3005
R6438 VDD.n2116 VDD.n1183 9.3005
R6439 VDD.n2115 VDD.n1184 9.3005
R6440 VDD.n2112 VDD.n1185 9.3005
R6441 VDD.n2111 VDD.n1186 9.3005
R6442 VDD.n2108 VDD.n1187 9.3005
R6443 VDD.n2104 VDD.n1188 9.3005
R6444 VDD.n2101 VDD.n1189 9.3005
R6445 VDD.n2100 VDD.n1190 9.3005
R6446 VDD.n2097 VDD.n1191 9.3005
R6447 VDD.n2096 VDD.n1192 9.3005
R6448 VDD.n2093 VDD.n1193 9.3005
R6449 VDD.n2092 VDD.n1194 9.3005
R6450 VDD.n2089 VDD.n1195 9.3005
R6451 VDD.n2088 VDD.n1196 9.3005
R6452 VDD.n2085 VDD.n1197 9.3005
R6453 VDD.n2168 VDD.n2167 9.3005
R6454 VDD.n1800 VDD.n1799 9.3005
R6455 VDD.n1314 VDD.n1313 9.3005
R6456 VDD.n1813 VDD.n1812 9.3005
R6457 VDD.n1814 VDD.n1312 9.3005
R6458 VDD.n1816 VDD.n1815 9.3005
R6459 VDD.n1302 VDD.n1301 9.3005
R6460 VDD.n1829 VDD.n1828 9.3005
R6461 VDD.n1830 VDD.n1300 9.3005
R6462 VDD.n1832 VDD.n1831 9.3005
R6463 VDD.n1290 VDD.n1289 9.3005
R6464 VDD.n1845 VDD.n1844 9.3005
R6465 VDD.n1846 VDD.n1288 9.3005
R6466 VDD.n1848 VDD.n1847 9.3005
R6467 VDD.n1278 VDD.n1277 9.3005
R6468 VDD.n1861 VDD.n1860 9.3005
R6469 VDD.n1862 VDD.n1276 9.3005
R6470 VDD.n1864 VDD.n1863 9.3005
R6471 VDD.n1266 VDD.n1265 9.3005
R6472 VDD.n1877 VDD.n1876 9.3005
R6473 VDD.n1878 VDD.n1264 9.3005
R6474 VDD.n1880 VDD.n1879 9.3005
R6475 VDD.n1254 VDD.n1253 9.3005
R6476 VDD.n1893 VDD.n1892 9.3005
R6477 VDD.n1894 VDD.n1252 9.3005
R6478 VDD.n1896 VDD.n1895 9.3005
R6479 VDD.n1242 VDD.n1241 9.3005
R6480 VDD.n1909 VDD.n1908 9.3005
R6481 VDD.n1910 VDD.n1240 9.3005
R6482 VDD.n1912 VDD.n1911 9.3005
R6483 VDD.n1230 VDD.n1229 9.3005
R6484 VDD.n1925 VDD.n1924 9.3005
R6485 VDD.n1926 VDD.n1228 9.3005
R6486 VDD.n1928 VDD.n1927 9.3005
R6487 VDD.n1218 VDD.n1217 9.3005
R6488 VDD.n1941 VDD.n1940 9.3005
R6489 VDD.n1942 VDD.n1216 9.3005
R6490 VDD.n1944 VDD.n1943 9.3005
R6491 VDD.n1206 VDD.n1205 9.3005
R6492 VDD.n1958 VDD.n1957 9.3005
R6493 VDD.n1959 VDD.n1204 9.3005
R6494 VDD.n1962 VDD.n1960 9.3005
R6495 VDD.n1961 VDD.n1138 9.3005
R6496 VDD.n3527 VDD.n3526 9.3005
R6497 VDD.n3532 VDD.n3521 9.3005
R6498 VDD.n3533 VDD.n3520 9.3005
R6499 VDD.n3534 VDD.n3519 9.3005
R6500 VDD.n3518 VDD.n3516 9.3005
R6501 VDD.n3540 VDD.n3515 9.3005
R6502 VDD.n3541 VDD.n3514 9.3005
R6503 VDD.n3542 VDD.n3513 9.3005
R6504 VDD.n3512 VDD.n3510 9.3005
R6505 VDD.n3548 VDD.n3509 9.3005
R6506 VDD.n3550 VDD.n3506 9.3005
R6507 VDD.n3551 VDD.n3505 9.3005
R6508 VDD.n3504 VDD.n3502 9.3005
R6509 VDD.n3557 VDD.n3501 9.3005
R6510 VDD.n3558 VDD.n3500 9.3005
R6511 VDD.n3559 VDD.n3499 9.3005
R6512 VDD.n3498 VDD.n3496 9.3005
R6513 VDD.n3565 VDD.n3495 9.3005
R6514 VDD.n3566 VDD.n3494 9.3005
R6515 VDD.n3567 VDD.n3493 9.3005
R6516 VDD.n3573 VDD.n3486 9.3005
R6517 VDD.n3574 VDD.n3485 9.3005
R6518 VDD.n3575 VDD.n3484 9.3005
R6519 VDD.n3483 VDD.n3481 9.3005
R6520 VDD.n3581 VDD.n3480 9.3005
R6521 VDD.n3582 VDD.n3479 9.3005
R6522 VDD.n3583 VDD.n3478 9.3005
R6523 VDD.n3477 VDD.n3475 9.3005
R6524 VDD.n3589 VDD.n3474 9.3005
R6525 VDD.n3591 VDD.n3470 9.3005
R6526 VDD.n3469 VDD.n3467 9.3005
R6527 VDD.n3596 VDD.n3466 9.3005
R6528 VDD.n3597 VDD.n3465 9.3005
R6529 VDD.n3464 VDD.n3462 9.3005
R6530 VDD.n3602 VDD.n396 9.3005
R6531 VDD.n3590 VDD.n3471 9.3005
R6532 VDD.n3492 VDD.n3487 9.3005
R6533 VDD.n3604 VDD.n3603 9.3005
R6534 VDD.n387 VDD.n386 9.3005
R6535 VDD.n3619 VDD.n3618 9.3005
R6536 VDD.n3620 VDD.n385 9.3005
R6537 VDD.n3622 VDD.n3621 9.3005
R6538 VDD.n375 VDD.n374 9.3005
R6539 VDD.n3634 VDD.n3633 9.3005
R6540 VDD.n3635 VDD.n373 9.3005
R6541 VDD.n3637 VDD.n3636 9.3005
R6542 VDD.n363 VDD.n362 9.3005
R6543 VDD.n3650 VDD.n3649 9.3005
R6544 VDD.n3651 VDD.n361 9.3005
R6545 VDD.n3653 VDD.n3652 9.3005
R6546 VDD.n351 VDD.n350 9.3005
R6547 VDD.n3666 VDD.n3665 9.3005
R6548 VDD.n3667 VDD.n349 9.3005
R6549 VDD.n3669 VDD.n3668 9.3005
R6550 VDD.n339 VDD.n338 9.3005
R6551 VDD.n3682 VDD.n3681 9.3005
R6552 VDD.n3683 VDD.n337 9.3005
R6553 VDD.n3685 VDD.n3684 9.3005
R6554 VDD.n327 VDD.n326 9.3005
R6555 VDD.n3698 VDD.n3697 9.3005
R6556 VDD.n3699 VDD.n325 9.3005
R6557 VDD.n3701 VDD.n3700 9.3005
R6558 VDD.n315 VDD.n314 9.3005
R6559 VDD.n3714 VDD.n3713 9.3005
R6560 VDD.n3715 VDD.n313 9.3005
R6561 VDD.n3717 VDD.n3716 9.3005
R6562 VDD.n303 VDD.n302 9.3005
R6563 VDD.n3730 VDD.n3729 9.3005
R6564 VDD.n3731 VDD.n301 9.3005
R6565 VDD.n3733 VDD.n3732 9.3005
R6566 VDD.n291 VDD.n290 9.3005
R6567 VDD.n3746 VDD.n3745 9.3005
R6568 VDD.n3747 VDD.n289 9.3005
R6569 VDD.n3749 VDD.n3748 9.3005
R6570 VDD.n279 VDD.n278 9.3005
R6571 VDD.n3762 VDD.n3761 9.3005
R6572 VDD.n3763 VDD.n277 9.3005
R6573 VDD.n3765 VDD.n3764 9.3005
R6574 VDD.n49 VDD.n47 9.3005
R6575 VDD.n3606 VDD.n3605 9.3005
R6576 VDD.n4000 VDD.n3999 9.3005
R6577 VDD.n50 VDD.n48 9.3005
R6578 VDD.n3993 VDD.n59 9.3005
R6579 VDD.n3992 VDD.n60 9.3005
R6580 VDD.n3991 VDD.n61 9.3005
R6581 VDD.n69 VDD.n62 9.3005
R6582 VDD.n3985 VDD.n70 9.3005
R6583 VDD.n3984 VDD.n71 9.3005
R6584 VDD.n3983 VDD.n72 9.3005
R6585 VDD.n80 VDD.n73 9.3005
R6586 VDD.n3977 VDD.n81 9.3005
R6587 VDD.n3976 VDD.n82 9.3005
R6588 VDD.n3975 VDD.n83 9.3005
R6589 VDD.n91 VDD.n84 9.3005
R6590 VDD.n3969 VDD.n92 9.3005
R6591 VDD.n3968 VDD.n93 9.3005
R6592 VDD.n3967 VDD.n94 9.3005
R6593 VDD.n102 VDD.n95 9.3005
R6594 VDD.n3961 VDD.n103 9.3005
R6595 VDD.n3960 VDD.n104 9.3005
R6596 VDD.n3959 VDD.n105 9.3005
R6597 VDD.n113 VDD.n106 9.3005
R6598 VDD.n3953 VDD.n114 9.3005
R6599 VDD.n3952 VDD.n115 9.3005
R6600 VDD.n3951 VDD.n116 9.3005
R6601 VDD.n124 VDD.n117 9.3005
R6602 VDD.n3945 VDD.n125 9.3005
R6603 VDD.n3944 VDD.n126 9.3005
R6604 VDD.n3943 VDD.n127 9.3005
R6605 VDD.n135 VDD.n128 9.3005
R6606 VDD.n3937 VDD.n136 9.3005
R6607 VDD.n3936 VDD.n137 9.3005
R6608 VDD.n3935 VDD.n138 9.3005
R6609 VDD.n146 VDD.n139 9.3005
R6610 VDD.n3929 VDD.n147 9.3005
R6611 VDD.n3928 VDD.n148 9.3005
R6612 VDD.n3927 VDD.n149 9.3005
R6613 VDD.n157 VDD.n150 9.3005
R6614 VDD.n3922 VDD.n158 9.3005
R6615 VDD.n3921 VDD.n159 9.3005
R6616 VDD.n3920 VDD.n160 9.3005
R6617 VDD.n168 VDD.n161 9.3005
R6618 VDD.n3914 VDD.n3913 9.3005
R6619 VDD.n3910 VDD.n169 9.3005
R6620 VDD.n3909 VDD.n171 9.3005
R6621 VDD.n175 VDD.n172 9.3005
R6622 VDD.n3904 VDD.n176 9.3005
R6623 VDD.n3903 VDD.n177 9.3005
R6624 VDD.n3902 VDD.n178 9.3005
R6625 VDD.n184 VDD.n181 9.3005
R6626 VDD.n3897 VDD.n185 9.3005
R6627 VDD.n3896 VDD.n186 9.3005
R6628 VDD.n3895 VDD.n187 9.3005
R6629 VDD.n191 VDD.n188 9.3005
R6630 VDD.n3890 VDD.n192 9.3005
R6631 VDD.n3889 VDD.n193 9.3005
R6632 VDD.n3888 VDD.n194 9.3005
R6633 VDD.n198 VDD.n195 9.3005
R6634 VDD.n3883 VDD.n199 9.3005
R6635 VDD.n3882 VDD.n200 9.3005
R6636 VDD.n3878 VDD.n201 9.3005
R6637 VDD.n205 VDD.n202 9.3005
R6638 VDD.n3873 VDD.n206 9.3005
R6639 VDD.n3872 VDD.n207 9.3005
R6640 VDD.n3871 VDD.n208 9.3005
R6641 VDD.n212 VDD.n209 9.3005
R6642 VDD.n3866 VDD.n213 9.3005
R6643 VDD.n3865 VDD.n214 9.3005
R6644 VDD.n3864 VDD.n215 9.3005
R6645 VDD.n222 VDD.n216 9.3005
R6646 VDD.n3859 VDD.n223 9.3005
R6647 VDD.n3858 VDD.n224 9.3005
R6648 VDD.n3857 VDD.n225 9.3005
R6649 VDD.n229 VDD.n226 9.3005
R6650 VDD.n3852 VDD.n230 9.3005
R6651 VDD.n3851 VDD.n231 9.3005
R6652 VDD.n3850 VDD.n232 9.3005
R6653 VDD.n236 VDD.n233 9.3005
R6654 VDD.n3845 VDD.n237 9.3005
R6655 VDD.n3844 VDD.n238 9.3005
R6656 VDD.n3840 VDD.n3837 9.3005
R6657 VDD.n3912 VDD.n3911 9.3005
R6658 VDD.n3612 VDD.n391 9.3005
R6659 VDD.n3614 VDD.n3613 9.3005
R6660 VDD.n381 VDD.n380 9.3005
R6661 VDD.n3626 VDD.n3625 9.3005
R6662 VDD.n3627 VDD.n379 9.3005
R6663 VDD.n3629 VDD.n3628 9.3005
R6664 VDD.n369 VDD.n368 9.3005
R6665 VDD.n3642 VDD.n3641 9.3005
R6666 VDD.n3643 VDD.n367 9.3005
R6667 VDD.n3645 VDD.n3644 9.3005
R6668 VDD.n357 VDD.n356 9.3005
R6669 VDD.n3658 VDD.n3657 9.3005
R6670 VDD.n3659 VDD.n355 9.3005
R6671 VDD.n3661 VDD.n3660 9.3005
R6672 VDD.n345 VDD.n344 9.3005
R6673 VDD.n3674 VDD.n3673 9.3005
R6674 VDD.n3675 VDD.n343 9.3005
R6675 VDD.n3677 VDD.n3676 9.3005
R6676 VDD.n333 VDD.n332 9.3005
R6677 VDD.n3690 VDD.n3689 9.3005
R6678 VDD.n3691 VDD.n331 9.3005
R6679 VDD.n3693 VDD.n3692 9.3005
R6680 VDD.n321 VDD.n320 9.3005
R6681 VDD.n3706 VDD.n3705 9.3005
R6682 VDD.n3707 VDD.n319 9.3005
R6683 VDD.n3709 VDD.n3708 9.3005
R6684 VDD.n309 VDD.n308 9.3005
R6685 VDD.n3722 VDD.n3721 9.3005
R6686 VDD.n3723 VDD.n307 9.3005
R6687 VDD.n3725 VDD.n3724 9.3005
R6688 VDD.n297 VDD.n296 9.3005
R6689 VDD.n3738 VDD.n3737 9.3005
R6690 VDD.n3739 VDD.n295 9.3005
R6691 VDD.n3741 VDD.n3740 9.3005
R6692 VDD.n285 VDD.n284 9.3005
R6693 VDD.n3754 VDD.n3753 9.3005
R6694 VDD.n3755 VDD.n283 9.3005
R6695 VDD.n3757 VDD.n3756 9.3005
R6696 VDD.n272 VDD.n271 9.3005
R6697 VDD.n3770 VDD.n3769 9.3005
R6698 VDD.n3771 VDD.n270 9.3005
R6699 VDD.n3773 VDD.n3772 9.3005
R6700 VDD.n3774 VDD.n269 9.3005
R6701 VDD.n3776 VDD.n3775 9.3005
R6702 VDD.n3777 VDD.n268 9.3005
R6703 VDD.n3779 VDD.n3778 9.3005
R6704 VDD.n3780 VDD.n266 9.3005
R6705 VDD.n3782 VDD.n3781 9.3005
R6706 VDD.n3783 VDD.n265 9.3005
R6707 VDD.n3785 VDD.n3784 9.3005
R6708 VDD.n3786 VDD.n263 9.3005
R6709 VDD.n3788 VDD.n3787 9.3005
R6710 VDD.n3789 VDD.n262 9.3005
R6711 VDD.n3791 VDD.n3790 9.3005
R6712 VDD.n3792 VDD.n260 9.3005
R6713 VDD.n3794 VDD.n3793 9.3005
R6714 VDD.n3795 VDD.n259 9.3005
R6715 VDD.n3797 VDD.n3796 9.3005
R6716 VDD.n3798 VDD.n257 9.3005
R6717 VDD.n3800 VDD.n3799 9.3005
R6718 VDD.n3801 VDD.n256 9.3005
R6719 VDD.n3803 VDD.n3802 9.3005
R6720 VDD.n3804 VDD.n254 9.3005
R6721 VDD.n3806 VDD.n3805 9.3005
R6722 VDD.n3807 VDD.n253 9.3005
R6723 VDD.n3809 VDD.n3808 9.3005
R6724 VDD.n3810 VDD.n251 9.3005
R6725 VDD.n3812 VDD.n3811 9.3005
R6726 VDD.n3813 VDD.n250 9.3005
R6727 VDD.n3815 VDD.n3814 9.3005
R6728 VDD.n3816 VDD.n248 9.3005
R6729 VDD.n3818 VDD.n3817 9.3005
R6730 VDD.n3819 VDD.n247 9.3005
R6731 VDD.n3821 VDD.n3820 9.3005
R6732 VDD.n3822 VDD.n245 9.3005
R6733 VDD.n3824 VDD.n3823 9.3005
R6734 VDD.n3825 VDD.n244 9.3005
R6735 VDD.n3827 VDD.n3826 9.3005
R6736 VDD.n3828 VDD.n242 9.3005
R6737 VDD.n3830 VDD.n3829 9.3005
R6738 VDD.n3831 VDD.n241 9.3005
R6739 VDD.n3833 VDD.n3832 9.3005
R6740 VDD.n3834 VDD.n239 9.3005
R6741 VDD.n3836 VDD.n3835 9.3005
R6742 VDD.n3611 VDD.n3610 9.3005
R6743 VDD.n3522 VDD.n392 9.3005
R6744 VDD.n2081 VDD.n2080 9.3005
R6745 VDD.n1596 VDD.n1595 9.3005
R6746 VDD.n1435 VDD.n1434 9.3005
R6747 VDD.n1609 VDD.n1608 9.3005
R6748 VDD.n1610 VDD.n1433 9.3005
R6749 VDD.n1612 VDD.n1611 9.3005
R6750 VDD.n1424 VDD.n1423 9.3005
R6751 VDD.n1625 VDD.n1624 9.3005
R6752 VDD.n1626 VDD.n1422 9.3005
R6753 VDD.n1628 VDD.n1627 9.3005
R6754 VDD.n1412 VDD.n1411 9.3005
R6755 VDD.n1641 VDD.n1640 9.3005
R6756 VDD.n1642 VDD.n1410 9.3005
R6757 VDD.n1644 VDD.n1643 9.3005
R6758 VDD.n1401 VDD.n1400 9.3005
R6759 VDD.n1658 VDD.n1657 9.3005
R6760 VDD.n1659 VDD.n1399 9.3005
R6761 VDD.n1661 VDD.n1660 9.3005
R6762 VDD.n1389 VDD.n1388 9.3005
R6763 VDD.n1674 VDD.n1673 9.3005
R6764 VDD.n1675 VDD.n1387 9.3005
R6765 VDD.n1677 VDD.n1676 9.3005
R6766 VDD.n1378 VDD.n1377 9.3005
R6767 VDD.n1691 VDD.n1690 9.3005
R6768 VDD.n1692 VDD.n1376 9.3005
R6769 VDD.n1694 VDD.n1693 9.3005
R6770 VDD.n1366 VDD.n1365 9.3005
R6771 VDD.n1707 VDD.n1706 9.3005
R6772 VDD.n1708 VDD.n1364 9.3005
R6773 VDD.n1710 VDD.n1709 9.3005
R6774 VDD.n1355 VDD.n1354 9.3005
R6775 VDD.n1724 VDD.n1723 9.3005
R6776 VDD.n1725 VDD.n1353 9.3005
R6777 VDD.n1727 VDD.n1726 9.3005
R6778 VDD.n1343 VDD.n1342 9.3005
R6779 VDD.n1740 VDD.n1739 9.3005
R6780 VDD.n1741 VDD.n1341 9.3005
R6781 VDD.n1743 VDD.n1742 9.3005
R6782 VDD.n1332 VDD.n1331 9.3005
R6783 VDD.n1757 VDD.n1756 9.3005
R6784 VDD.n1758 VDD.n1330 9.3005
R6785 VDD.n1760 VDD.n1759 9.3005
R6786 VDD.n1320 VDD.n1319 9.3005
R6787 VDD.n1805 VDD.n1804 9.3005
R6788 VDD.n1806 VDD.n1318 9.3005
R6789 VDD.n1808 VDD.n1807 9.3005
R6790 VDD.n1308 VDD.n1307 9.3005
R6791 VDD.n1821 VDD.n1820 9.3005
R6792 VDD.n1822 VDD.n1306 9.3005
R6793 VDD.n1824 VDD.n1823 9.3005
R6794 VDD.n1296 VDD.n1295 9.3005
R6795 VDD.n1837 VDD.n1836 9.3005
R6796 VDD.n1838 VDD.n1294 9.3005
R6797 VDD.n1840 VDD.n1839 9.3005
R6798 VDD.n1284 VDD.n1283 9.3005
R6799 VDD.n1853 VDD.n1852 9.3005
R6800 VDD.n1854 VDD.n1282 9.3005
R6801 VDD.n1856 VDD.n1855 9.3005
R6802 VDD.n1272 VDD.n1271 9.3005
R6803 VDD.n1869 VDD.n1868 9.3005
R6804 VDD.n1870 VDD.n1270 9.3005
R6805 VDD.n1872 VDD.n1871 9.3005
R6806 VDD.n1260 VDD.n1259 9.3005
R6807 VDD.n1885 VDD.n1884 9.3005
R6808 VDD.n1886 VDD.n1258 9.3005
R6809 VDD.n1888 VDD.n1887 9.3005
R6810 VDD.n1248 VDD.n1247 9.3005
R6811 VDD.n1901 VDD.n1900 9.3005
R6812 VDD.n1902 VDD.n1246 9.3005
R6813 VDD.n1904 VDD.n1903 9.3005
R6814 VDD.n1236 VDD.n1235 9.3005
R6815 VDD.n1917 VDD.n1916 9.3005
R6816 VDD.n1918 VDD.n1234 9.3005
R6817 VDD.n1920 VDD.n1919 9.3005
R6818 VDD.n1224 VDD.n1223 9.3005
R6819 VDD.n1933 VDD.n1932 9.3005
R6820 VDD.n1934 VDD.n1222 9.3005
R6821 VDD.n1936 VDD.n1935 9.3005
R6822 VDD.n1212 VDD.n1211 9.3005
R6823 VDD.n1949 VDD.n1948 9.3005
R6824 VDD.n1950 VDD.n1209 9.3005
R6825 VDD.n1953 VDD.n1952 9.3005
R6826 VDD.n1951 VDD.n1210 9.3005
R6827 VDD.n1200 VDD.n1199 9.3005
R6828 VDD.n1968 VDD.n1967 9.3005
R6829 VDD.n1594 VDD.n1445 9.3005
R6830 VDD.n1523 VDD.n1446 9.3005
R6831 VDD.n1525 VDD.n1524 9.3005
R6832 VDD.n1526 VDD.n1519 9.3005
R6833 VDD.n1528 VDD.n1527 9.3005
R6834 VDD.n1529 VDD.n1518 9.3005
R6835 VDD.n1531 VDD.n1530 9.3005
R6836 VDD.n1532 VDD.n1513 9.3005
R6837 VDD.n1534 VDD.n1533 9.3005
R6838 VDD.n1535 VDD.n1512 9.3005
R6839 VDD.n1537 VDD.n1536 9.3005
R6840 VDD.n1541 VDD.n1507 9.3005
R6841 VDD.n1543 VDD.n1542 9.3005
R6842 VDD.n1544 VDD.n1506 9.3005
R6843 VDD.n1546 VDD.n1545 9.3005
R6844 VDD.n1547 VDD.n1501 9.3005
R6845 VDD.n1549 VDD.n1548 9.3005
R6846 VDD.n1550 VDD.n1500 9.3005
R6847 VDD.n1552 VDD.n1551 9.3005
R6848 VDD.n1553 VDD.n1495 9.3005
R6849 VDD.n1555 VDD.n1554 9.3005
R6850 VDD.n1558 VDD.n1487 9.3005
R6851 VDD.n1560 VDD.n1559 9.3005
R6852 VDD.n1561 VDD.n1486 9.3005
R6853 VDD.n1563 VDD.n1562 9.3005
R6854 VDD.n1564 VDD.n1481 9.3005
R6855 VDD.n1566 VDD.n1565 9.3005
R6856 VDD.n1567 VDD.n1480 9.3005
R6857 VDD.n1569 VDD.n1568 9.3005
R6858 VDD.n1570 VDD.n1477 9.3005
R6859 VDD.n1577 VDD.n1476 9.3005
R6860 VDD.n1579 VDD.n1578 9.3005
R6861 VDD.n1580 VDD.n1472 9.3005
R6862 VDD.n1582 VDD.n1581 9.3005
R6863 VDD.n1583 VDD.n1471 9.3005
R6864 VDD.n1585 VDD.n1584 9.3005
R6865 VDD.n1586 VDD.n1470 9.3005
R6866 VDD.n1576 VDD.n1575 9.3005
R6867 VDD.n1557 VDD.n1556 9.3005
R6868 VDD.n1593 VDD.n1592 9.3005
R6869 VDD.n1601 VDD.n1600 9.3005
R6870 VDD.n1602 VDD.n1439 9.3005
R6871 VDD.n1604 VDD.n1603 9.3005
R6872 VDD.n1430 VDD.n1429 9.3005
R6873 VDD.n1617 VDD.n1616 9.3005
R6874 VDD.n1618 VDD.n1428 9.3005
R6875 VDD.n1620 VDD.n1619 9.3005
R6876 VDD.n1418 VDD.n1417 9.3005
R6877 VDD.n1633 VDD.n1632 9.3005
R6878 VDD.n1634 VDD.n1416 9.3005
R6879 VDD.n1636 VDD.n1635 9.3005
R6880 VDD.n1406 VDD.n1405 9.3005
R6881 VDD.n1650 VDD.n1649 9.3005
R6882 VDD.n1651 VDD.n1404 9.3005
R6883 VDD.n1653 VDD.n1652 9.3005
R6884 VDD.n1395 VDD.n1394 9.3005
R6885 VDD.n1666 VDD.n1665 9.3005
R6886 VDD.n1667 VDD.n1393 9.3005
R6887 VDD.n1669 VDD.n1668 9.3005
R6888 VDD.n1383 VDD.n1382 9.3005
R6889 VDD.n1683 VDD.n1682 9.3005
R6890 VDD.n1684 VDD.n1381 9.3005
R6891 VDD.n1686 VDD.n1685 9.3005
R6892 VDD.n1372 VDD.n1371 9.3005
R6893 VDD.n1699 VDD.n1698 9.3005
R6894 VDD.n1700 VDD.n1370 9.3005
R6895 VDD.n1702 VDD.n1701 9.3005
R6896 VDD.n1360 VDD.n1359 9.3005
R6897 VDD.n1716 VDD.n1715 9.3005
R6898 VDD.n1717 VDD.n1358 9.3005
R6899 VDD.n1719 VDD.n1718 9.3005
R6900 VDD.n1349 VDD.n1348 9.3005
R6901 VDD.n1732 VDD.n1731 9.3005
R6902 VDD.n1733 VDD.n1347 9.3005
R6903 VDD.n1735 VDD.n1734 9.3005
R6904 VDD.n1337 VDD.n1336 9.3005
R6905 VDD.n1749 VDD.n1748 9.3005
R6906 VDD.n1750 VDD.n1335 9.3005
R6907 VDD.n1752 VDD.n1751 9.3005
R6908 VDD.n1326 VDD.n1325 9.3005
R6909 VDD.n1765 VDD.n1764 9.3005
R6910 VDD.n1441 VDD.n1440 9.3005
R6911 VDD.n1798 VDD.n1324 9.3005
R6912 VDD.n2604 VDD.n2603 8.58587
R6913 VDD.n1120 VDD.n1047 8.58587
R6914 VDD.n3044 VDD.n2726 8.58587
R6915 VDD.n3445 VDD.n3444 8.58587
R6916 VDD.n447 VDD.n442 8.58587
R6917 VDD.n2892 VDD.n2891 8.58587
R6918 VDD.n2659 VDD.n738 8.58587
R6919 VDD.n2062 VDD.n1991 8.58587
R6920 VDD.n15 VDD.n14 8.31282
R6921 VDD.n4001 VDD.n4000 8.18662
R6922 VDD.n1798 VDD.n1797 8.18662
R6923 VDD.n1004 VDD.t5 7.86674
R6924 VDD.n2399 VDD.t54 7.86674
R6925 VDD.n3026 VDD.t9 7.86674
R6926 VDD.t41 VDD.n450 7.86674
R6927 VDD.n2399 VDD.t111 7.71547
R6928 VDD.n3026 VDD.t96 7.71547
R6929 VDD.n997 VDD.t88 7.41292
R6930 VDD.n2471 VDD.t86 7.41292
R6931 VDD.n3207 VDD.t200 7.41292
R6932 VDD.t202 VDD.n456 7.41292
R6933 VDD.n1575 VDD.n1570 7.17626
R6934 VDD.n2153 VDD.n1167 7.17626
R6935 VDD.n3897 VDD.n181 7.17626
R6936 VDD.n3590 VDD.n3589 7.17626
R6937 VDD.t3 VDD.n912 6.9591
R6938 VDD.n849 VDD.t95 6.9591
R6939 VDD.t90 VDD.n601 6.9591
R6940 VDD.n543 VDD.t116 6.9591
R6941 VDD.n2259 VDD.t107 6.65655
R6942 VDD.n2531 VDD.t113 6.65655
R6943 VDD.n3147 VDD.t0 6.65655
R6944 VDD.n3290 VDD.t104 6.65655
R6945 VDD.n1554 VDD.n1494 6.4005
R6946 VDD.n2130 VDD.n2127 6.4005
R6947 VDD.n3881 VDD.n3878 6.4005
R6948 VDD.n3567 VDD.n3491 6.4005
R6949 VDD.n2259 VDD.t98 6.20273
R6950 VDD.t105 VDD.n823 6.20273
R6951 VDD.n627 VDD.t1 6.20273
R6952 VDD.n3290 VDD.t198 6.20273
R6953 VDD.n7 VDD.t203 5.9105
R6954 VDD.n7 VDD.t115 5.9105
R6955 VDD.n8 VDD.t85 5.9105
R6956 VDD.n8 VDD.t199 5.9105
R6957 VDD.n10 VDD.t2 5.9105
R6958 VDD.n10 VDD.t201 5.9105
R6959 VDD.n12 VDD.t97 5.9105
R6960 VDD.n12 VDD.t110 5.9105
R6961 VDD.n5 VDD.t94 5.9105
R6962 VDD.n5 VDD.t112 5.9105
R6963 VDD.n3 VDD.t87 5.9105
R6964 VDD.n3 VDD.t106 5.9105
R6965 VDD.n1 VDD.t99 5.9105
R6966 VDD.n1 VDD.t103 5.9105
R6967 VDD.n0 VDD.t92 5.9105
R6968 VDD.n0 VDD.t89 5.9105
R6969 VDD.n30 VDD.n22 5.78929
R6970 VDD.n1780 VDD.n1772 5.78929
R6971 VDD.n4001 VDD.n46 5.69978
R6972 VDD.n1797 VDD.n1796 5.69978
R6973 VDD.n1540 VDD.n1537 5.62474
R6974 VDD.n2107 VDD.n2104 5.62474
R6975 VDD.n3859 VDD.n221 5.62474
R6976 VDD.n3549 VDD.n3548 5.62474
R6977 VDD.n2170 VDD.n2169 5.30782
R6978 VDD.n2169 VDD.n1136 5.30782
R6979 VDD.n3461 VDD.n397 5.30782
R6980 VDD.n3461 VDD.n3460 5.30782
R6981 VDD.n3373 VDD.n435 5.30782
R6982 VDD.n437 VDD.n435 5.30782
R6983 VDD.n2079 VDD.n1988 5.30782
R6984 VDD.n2079 VDD.n2078 5.30782
R6985 VDD.n1592 VDD.n1449 4.84898
R6986 VDD.n2084 VDD.n2081 4.84898
R6987 VDD.n3843 VDD.n3840 4.84898
R6988 VDD.n3525 VDD.n3522 4.84898
R6989 VDD.n46 VDD.n45 4.7074
R6990 VDD.n38 VDD.n37 4.7074
R6991 VDD.n30 VDD.n29 4.7074
R6992 VDD.n1796 VDD.n1795 4.7074
R6993 VDD.n1788 VDD.n1787 4.7074
R6994 VDD.n1780 VDD.n1779 4.7074
R6995 VDD.n962 VDD.t98 4.08489
R6996 VDD.n2507 VDD.t105 4.08489
R6997 VDD.n3171 VDD.t1 4.08489
R6998 VDD.t198 VDD.n493 4.08489
R6999 VDD.t107 VDD.n948 3.63107
R7000 VDD.n813 VDD.t113 3.63107
R7001 VDD.t0 VDD.n637 3.63107
R7002 VDD.n507 VDD.t104 3.63107
R7003 VDD.n2295 VDD.t3 3.32853
R7004 VDD.n2495 VDD.t95 3.32853
R7005 VDD.n3183 VDD.t90 3.32853
R7006 VDD.n3254 VDD.t116 3.32853
R7007 VDD.n2223 VDD.t88 2.8747
R7008 VDD.t86 VDD.n859 2.8747
R7009 VDD.n591 VDD.t200 2.8747
R7010 VDD.n3326 VDD.t202 2.8747
R7011 VDD.n2584 VDD.t111 2.57216
R7012 VDD.n3099 VDD.t96 2.57216
R7013 VDD.n2217 VDD.t5 2.42088
R7014 VDD.n2573 VDD.t54 2.42088
R7015 VDD.n3105 VDD.t9 2.42088
R7016 VDD.n3334 VDD.t41 2.42088
R7017 VDD.n4 VDD.n2 2.14921
R7018 VDD.n11 VDD.n9 2.14921
R7019 VDD.n1646 VDD.t147 2.11833
R7020 VDD.t118 VDD.n1238 2.11833
R7021 VDD.n3663 VDD.t144 2.11833
R7022 VDD.n3941 VDD.t158 2.11833
R7023 VDD.n1797 VDD.n15 2.07022
R7024 VDD VDD.n4001 2.06239
R7025 VDD.n2603 VDD.n2602 2.02977
R7026 VDD.n1117 VDD.n1047 2.02977
R7027 VDD.n3041 VDD.n2726 2.02977
R7028 VDD.n3444 VDD.n3443 2.02977
R7029 VDD.n3354 VDD.n447 2.02977
R7030 VDD.n2893 VDD.n2892 2.02977
R7031 VDD.n2656 VDD.n738 2.02977
R7032 VDD.n2059 VDD.n1991 2.02977
R7033 VDD.n1523 VDD.n1449 1.74595
R7034 VDD.n2085 VDD.n2084 1.74595
R7035 VDD.n3844 VDD.n3843 1.74595
R7036 VDD.n3527 VDD.n3525 1.74595
R7037 VDD.n42 VDD.n40 1.71602
R7038 VDD.n44 VDD.n42 1.71602
R7039 VDD.n45 VDD.n44 1.71602
R7040 VDD.n34 VDD.n32 1.71602
R7041 VDD.n36 VDD.n34 1.71602
R7042 VDD.n37 VDD.n36 1.71602
R7043 VDD.n26 VDD.n24 1.71602
R7044 VDD.n28 VDD.n26 1.71602
R7045 VDD.n29 VDD.n28 1.71602
R7046 VDD.n19 VDD.n17 1.71602
R7047 VDD.n21 VDD.n19 1.71602
R7048 VDD.n22 VDD.n21 1.71602
R7049 VDD.n1795 VDD.n1794 1.71602
R7050 VDD.n1794 VDD.n1792 1.71602
R7051 VDD.n1792 VDD.n1790 1.71602
R7052 VDD.n1787 VDD.n1786 1.71602
R7053 VDD.n1786 VDD.n1784 1.71602
R7054 VDD.n1784 VDD.n1782 1.71602
R7055 VDD.n1779 VDD.n1778 1.71602
R7056 VDD.n1778 VDD.n1776 1.71602
R7057 VDD.n1776 VDD.n1774 1.71602
R7058 VDD.n1772 VDD.n1771 1.71602
R7059 VDD.n1771 VDD.n1769 1.71602
R7060 VDD.n1769 VDD.n1767 1.71602
R7061 VDD.n6 VDD.n4 1.71171
R7062 VDD.n13 VDD.n11 1.71171
R7063 VDD.n1679 VDD.t156 1.51324
R7064 VDD.t149 VDD.n1262 1.51324
R7065 VDD.n3695 VDD.t127 1.51324
R7066 VDD.n3957 VDD.t129 1.51324
R7067 VDD.n14 VDD.n6 1.34964
R7068 VDD.n14 VDD.n13 1.34964
R7069 VDD.n46 VDD.n38 1.0824
R7070 VDD.n38 VDD.n30 1.0824
R7071 VDD.n1796 VDD.n1788 1.0824
R7072 VDD.n1788 VDD.n1780 1.0824
R7073 VDD.n1541 VDD.n1540 0.970197
R7074 VDD.n2108 VDD.n2107 0.970197
R7075 VDD.n221 VDD.n216 0.970197
R7076 VDD.n3550 VDD.n3549 0.970197
R7077 VDD.n1712 VDD.t154 0.908143
R7078 VDD.t142 VDD.n1286 0.908143
R7079 VDD.n3727 VDD.t120 0.908143
R7080 VDD.n3973 VDD.t140 0.908143
R7081 VDD.n926 VDD.t102 0.756869
R7082 VDD.n2543 VDD.t93 0.756869
R7083 VDD.n3135 VDD.t109 0.756869
R7084 VDD.t84 VDD.n529 0.756869
R7085 VDD.n3913 VDD.n3912 0.529463
R7086 VDD.n3837 VDD.n3836 0.529463
R7087 VDD.n1594 VDD.n1593 0.529463
R7088 VDD.n1470 VDD.n1440 0.529463
R7089 VDD.n1745 VDD.t122 0.303048
R7090 VDD.t124 VDD.n1310 0.303048
R7091 VDD.n3759 VDD.t135 0.303048
R7092 VDD.n3989 VDD.t137 0.303048
R7093 VDD.n2168 VDD.n1138 0.24727
R7094 VDD.n3605 VDD.n3604 0.24727
R7095 VDD.n3611 VDD.n392 0.240447
R7096 VDD.n2080 VDD.n1968 0.240447
R7097 VDD.n1557 VDD.n1494 0.194439
R7098 VDD.n2131 VDD.n2130 0.194439
R7099 VDD.n3882 VDD.n3881 0.194439
R7100 VDD.n3491 VDD.n3487 0.194439
R7101 VDD.n1162 VDD.n1137 0.152939
R7102 VDD.n1163 VDD.n1162 0.152939
R7103 VDD.n1164 VDD.n1163 0.152939
R7104 VDD.n1165 VDD.n1164 0.152939
R7105 VDD.n1166 VDD.n1165 0.152939
R7106 VDD.n2152 VDD.n1166 0.152939
R7107 VDD.n2152 VDD.n2151 0.152939
R7108 VDD.n2151 VDD.n2150 0.152939
R7109 VDD.n2150 VDD.n1170 0.152939
R7110 VDD.n1171 VDD.n1170 0.152939
R7111 VDD.n1172 VDD.n1171 0.152939
R7112 VDD.n1173 VDD.n1172 0.152939
R7113 VDD.n1174 VDD.n1173 0.152939
R7114 VDD.n1175 VDD.n1174 0.152939
R7115 VDD.n1176 VDD.n1175 0.152939
R7116 VDD.n1177 VDD.n1176 0.152939
R7117 VDD.n1178 VDD.n1177 0.152939
R7118 VDD.n1179 VDD.n1178 0.152939
R7119 VDD.n1180 VDD.n1179 0.152939
R7120 VDD.n1181 VDD.n1180 0.152939
R7121 VDD.n1182 VDD.n1181 0.152939
R7122 VDD.n1183 VDD.n1182 0.152939
R7123 VDD.n1184 VDD.n1183 0.152939
R7124 VDD.n1185 VDD.n1184 0.152939
R7125 VDD.n1186 VDD.n1185 0.152939
R7126 VDD.n1187 VDD.n1186 0.152939
R7127 VDD.n1188 VDD.n1187 0.152939
R7128 VDD.n1189 VDD.n1188 0.152939
R7129 VDD.n1190 VDD.n1189 0.152939
R7130 VDD.n1191 VDD.n1190 0.152939
R7131 VDD.n1192 VDD.n1191 0.152939
R7132 VDD.n1193 VDD.n1192 0.152939
R7133 VDD.n1194 VDD.n1193 0.152939
R7134 VDD.n1195 VDD.n1194 0.152939
R7135 VDD.n1196 VDD.n1195 0.152939
R7136 VDD.n1197 VDD.n1196 0.152939
R7137 VDD.n1799 VDD.n1313 0.152939
R7138 VDD.n1813 VDD.n1313 0.152939
R7139 VDD.n1814 VDD.n1813 0.152939
R7140 VDD.n1815 VDD.n1814 0.152939
R7141 VDD.n1815 VDD.n1301 0.152939
R7142 VDD.n1829 VDD.n1301 0.152939
R7143 VDD.n1830 VDD.n1829 0.152939
R7144 VDD.n1831 VDD.n1830 0.152939
R7145 VDD.n1831 VDD.n1289 0.152939
R7146 VDD.n1845 VDD.n1289 0.152939
R7147 VDD.n1846 VDD.n1845 0.152939
R7148 VDD.n1847 VDD.n1846 0.152939
R7149 VDD.n1847 VDD.n1277 0.152939
R7150 VDD.n1861 VDD.n1277 0.152939
R7151 VDD.n1862 VDD.n1861 0.152939
R7152 VDD.n1863 VDD.n1862 0.152939
R7153 VDD.n1863 VDD.n1265 0.152939
R7154 VDD.n1877 VDD.n1265 0.152939
R7155 VDD.n1878 VDD.n1877 0.152939
R7156 VDD.n1879 VDD.n1878 0.152939
R7157 VDD.n1879 VDD.n1253 0.152939
R7158 VDD.n1893 VDD.n1253 0.152939
R7159 VDD.n1894 VDD.n1893 0.152939
R7160 VDD.n1895 VDD.n1894 0.152939
R7161 VDD.n1895 VDD.n1241 0.152939
R7162 VDD.n1909 VDD.n1241 0.152939
R7163 VDD.n1910 VDD.n1909 0.152939
R7164 VDD.n1911 VDD.n1910 0.152939
R7165 VDD.n1911 VDD.n1229 0.152939
R7166 VDD.n1925 VDD.n1229 0.152939
R7167 VDD.n1926 VDD.n1925 0.152939
R7168 VDD.n1927 VDD.n1926 0.152939
R7169 VDD.n1927 VDD.n1217 0.152939
R7170 VDD.n1941 VDD.n1217 0.152939
R7171 VDD.n1942 VDD.n1941 0.152939
R7172 VDD.n1943 VDD.n1942 0.152939
R7173 VDD.n1943 VDD.n1205 0.152939
R7174 VDD.n1958 VDD.n1205 0.152939
R7175 VDD.n1959 VDD.n1958 0.152939
R7176 VDD.n1960 VDD.n1959 0.152939
R7177 VDD.n1960 VDD.n1138 0.152939
R7178 VDD.n3464 VDD.n396 0.152939
R7179 VDD.n3465 VDD.n3464 0.152939
R7180 VDD.n3466 VDD.n3465 0.152939
R7181 VDD.n3469 VDD.n3466 0.152939
R7182 VDD.n3470 VDD.n3469 0.152939
R7183 VDD.n3471 VDD.n3470 0.152939
R7184 VDD.n3474 VDD.n3471 0.152939
R7185 VDD.n3477 VDD.n3474 0.152939
R7186 VDD.n3478 VDD.n3477 0.152939
R7187 VDD.n3479 VDD.n3478 0.152939
R7188 VDD.n3480 VDD.n3479 0.152939
R7189 VDD.n3483 VDD.n3480 0.152939
R7190 VDD.n3484 VDD.n3483 0.152939
R7191 VDD.n3485 VDD.n3484 0.152939
R7192 VDD.n3486 VDD.n3485 0.152939
R7193 VDD.n3492 VDD.n3486 0.152939
R7194 VDD.n3493 VDD.n3492 0.152939
R7195 VDD.n3494 VDD.n3493 0.152939
R7196 VDD.n3495 VDD.n3494 0.152939
R7197 VDD.n3498 VDD.n3495 0.152939
R7198 VDD.n3499 VDD.n3498 0.152939
R7199 VDD.n3500 VDD.n3499 0.152939
R7200 VDD.n3501 VDD.n3500 0.152939
R7201 VDD.n3504 VDD.n3501 0.152939
R7202 VDD.n3505 VDD.n3504 0.152939
R7203 VDD.n3506 VDD.n3505 0.152939
R7204 VDD.n3509 VDD.n3506 0.152939
R7205 VDD.n3512 VDD.n3509 0.152939
R7206 VDD.n3513 VDD.n3512 0.152939
R7207 VDD.n3514 VDD.n3513 0.152939
R7208 VDD.n3515 VDD.n3514 0.152939
R7209 VDD.n3518 VDD.n3515 0.152939
R7210 VDD.n3519 VDD.n3518 0.152939
R7211 VDD.n3520 VDD.n3519 0.152939
R7212 VDD.n3521 VDD.n3520 0.152939
R7213 VDD.n3526 VDD.n3521 0.152939
R7214 VDD.n3605 VDD.n386 0.152939
R7215 VDD.n3619 VDD.n386 0.152939
R7216 VDD.n3620 VDD.n3619 0.152939
R7217 VDD.n3621 VDD.n3620 0.152939
R7218 VDD.n3621 VDD.n374 0.152939
R7219 VDD.n3634 VDD.n374 0.152939
R7220 VDD.n3635 VDD.n3634 0.152939
R7221 VDD.n3636 VDD.n3635 0.152939
R7222 VDD.n3636 VDD.n362 0.152939
R7223 VDD.n3650 VDD.n362 0.152939
R7224 VDD.n3651 VDD.n3650 0.152939
R7225 VDD.n3652 VDD.n3651 0.152939
R7226 VDD.n3652 VDD.n350 0.152939
R7227 VDD.n3666 VDD.n350 0.152939
R7228 VDD.n3667 VDD.n3666 0.152939
R7229 VDD.n3668 VDD.n3667 0.152939
R7230 VDD.n3668 VDD.n338 0.152939
R7231 VDD.n3682 VDD.n338 0.152939
R7232 VDD.n3683 VDD.n3682 0.152939
R7233 VDD.n3684 VDD.n3683 0.152939
R7234 VDD.n3684 VDD.n326 0.152939
R7235 VDD.n3698 VDD.n326 0.152939
R7236 VDD.n3699 VDD.n3698 0.152939
R7237 VDD.n3700 VDD.n3699 0.152939
R7238 VDD.n3700 VDD.n314 0.152939
R7239 VDD.n3714 VDD.n314 0.152939
R7240 VDD.n3715 VDD.n3714 0.152939
R7241 VDD.n3716 VDD.n3715 0.152939
R7242 VDD.n3716 VDD.n302 0.152939
R7243 VDD.n3730 VDD.n302 0.152939
R7244 VDD.n3731 VDD.n3730 0.152939
R7245 VDD.n3732 VDD.n3731 0.152939
R7246 VDD.n3732 VDD.n290 0.152939
R7247 VDD.n3746 VDD.n290 0.152939
R7248 VDD.n3747 VDD.n3746 0.152939
R7249 VDD.n3748 VDD.n3747 0.152939
R7250 VDD.n3748 VDD.n278 0.152939
R7251 VDD.n3762 VDD.n278 0.152939
R7252 VDD.n3763 VDD.n3762 0.152939
R7253 VDD.n3764 VDD.n3763 0.152939
R7254 VDD.n3764 VDD.n47 0.152939
R7255 VDD.n59 VDD.n48 0.152939
R7256 VDD.n60 VDD.n59 0.152939
R7257 VDD.n61 VDD.n60 0.152939
R7258 VDD.n69 VDD.n61 0.152939
R7259 VDD.n70 VDD.n69 0.152939
R7260 VDD.n71 VDD.n70 0.152939
R7261 VDD.n72 VDD.n71 0.152939
R7262 VDD.n80 VDD.n72 0.152939
R7263 VDD.n81 VDD.n80 0.152939
R7264 VDD.n82 VDD.n81 0.152939
R7265 VDD.n83 VDD.n82 0.152939
R7266 VDD.n91 VDD.n83 0.152939
R7267 VDD.n92 VDD.n91 0.152939
R7268 VDD.n93 VDD.n92 0.152939
R7269 VDD.n94 VDD.n93 0.152939
R7270 VDD.n102 VDD.n94 0.152939
R7271 VDD.n103 VDD.n102 0.152939
R7272 VDD.n104 VDD.n103 0.152939
R7273 VDD.n105 VDD.n104 0.152939
R7274 VDD.n113 VDD.n105 0.152939
R7275 VDD.n114 VDD.n113 0.152939
R7276 VDD.n115 VDD.n114 0.152939
R7277 VDD.n116 VDD.n115 0.152939
R7278 VDD.n124 VDD.n116 0.152939
R7279 VDD.n125 VDD.n124 0.152939
R7280 VDD.n126 VDD.n125 0.152939
R7281 VDD.n127 VDD.n126 0.152939
R7282 VDD.n135 VDD.n127 0.152939
R7283 VDD.n136 VDD.n135 0.152939
R7284 VDD.n137 VDD.n136 0.152939
R7285 VDD.n138 VDD.n137 0.152939
R7286 VDD.n146 VDD.n138 0.152939
R7287 VDD.n147 VDD.n146 0.152939
R7288 VDD.n148 VDD.n147 0.152939
R7289 VDD.n149 VDD.n148 0.152939
R7290 VDD.n157 VDD.n149 0.152939
R7291 VDD.n158 VDD.n157 0.152939
R7292 VDD.n159 VDD.n158 0.152939
R7293 VDD.n160 VDD.n159 0.152939
R7294 VDD.n168 VDD.n160 0.152939
R7295 VDD.n3913 VDD.n168 0.152939
R7296 VDD.n3912 VDD.n169 0.152939
R7297 VDD.n171 VDD.n169 0.152939
R7298 VDD.n175 VDD.n171 0.152939
R7299 VDD.n176 VDD.n175 0.152939
R7300 VDD.n177 VDD.n176 0.152939
R7301 VDD.n178 VDD.n177 0.152939
R7302 VDD.n184 VDD.n178 0.152939
R7303 VDD.n185 VDD.n184 0.152939
R7304 VDD.n186 VDD.n185 0.152939
R7305 VDD.n187 VDD.n186 0.152939
R7306 VDD.n191 VDD.n187 0.152939
R7307 VDD.n192 VDD.n191 0.152939
R7308 VDD.n193 VDD.n192 0.152939
R7309 VDD.n194 VDD.n193 0.152939
R7310 VDD.n198 VDD.n194 0.152939
R7311 VDD.n199 VDD.n198 0.152939
R7312 VDD.n200 VDD.n199 0.152939
R7313 VDD.n201 VDD.n200 0.152939
R7314 VDD.n205 VDD.n201 0.152939
R7315 VDD.n206 VDD.n205 0.152939
R7316 VDD.n207 VDD.n206 0.152939
R7317 VDD.n208 VDD.n207 0.152939
R7318 VDD.n212 VDD.n208 0.152939
R7319 VDD.n213 VDD.n212 0.152939
R7320 VDD.n214 VDD.n213 0.152939
R7321 VDD.n215 VDD.n214 0.152939
R7322 VDD.n222 VDD.n215 0.152939
R7323 VDD.n223 VDD.n222 0.152939
R7324 VDD.n224 VDD.n223 0.152939
R7325 VDD.n225 VDD.n224 0.152939
R7326 VDD.n229 VDD.n225 0.152939
R7327 VDD.n230 VDD.n229 0.152939
R7328 VDD.n231 VDD.n230 0.152939
R7329 VDD.n232 VDD.n231 0.152939
R7330 VDD.n236 VDD.n232 0.152939
R7331 VDD.n237 VDD.n236 0.152939
R7332 VDD.n238 VDD.n237 0.152939
R7333 VDD.n3837 VDD.n238 0.152939
R7334 VDD.n3612 VDD.n3611 0.152939
R7335 VDD.n3613 VDD.n3612 0.152939
R7336 VDD.n3613 VDD.n380 0.152939
R7337 VDD.n3626 VDD.n380 0.152939
R7338 VDD.n3627 VDD.n3626 0.152939
R7339 VDD.n3628 VDD.n3627 0.152939
R7340 VDD.n3628 VDD.n368 0.152939
R7341 VDD.n3642 VDD.n368 0.152939
R7342 VDD.n3643 VDD.n3642 0.152939
R7343 VDD.n3644 VDD.n3643 0.152939
R7344 VDD.n3644 VDD.n356 0.152939
R7345 VDD.n3658 VDD.n356 0.152939
R7346 VDD.n3659 VDD.n3658 0.152939
R7347 VDD.n3660 VDD.n3659 0.152939
R7348 VDD.n3660 VDD.n344 0.152939
R7349 VDD.n3674 VDD.n344 0.152939
R7350 VDD.n3675 VDD.n3674 0.152939
R7351 VDD.n3676 VDD.n3675 0.152939
R7352 VDD.n3676 VDD.n332 0.152939
R7353 VDD.n3690 VDD.n332 0.152939
R7354 VDD.n3691 VDD.n3690 0.152939
R7355 VDD.n3692 VDD.n3691 0.152939
R7356 VDD.n3692 VDD.n320 0.152939
R7357 VDD.n3706 VDD.n320 0.152939
R7358 VDD.n3707 VDD.n3706 0.152939
R7359 VDD.n3708 VDD.n3707 0.152939
R7360 VDD.n3708 VDD.n308 0.152939
R7361 VDD.n3722 VDD.n308 0.152939
R7362 VDD.n3723 VDD.n3722 0.152939
R7363 VDD.n3724 VDD.n3723 0.152939
R7364 VDD.n3724 VDD.n296 0.152939
R7365 VDD.n3738 VDD.n296 0.152939
R7366 VDD.n3739 VDD.n3738 0.152939
R7367 VDD.n3740 VDD.n3739 0.152939
R7368 VDD.n3740 VDD.n284 0.152939
R7369 VDD.n3754 VDD.n284 0.152939
R7370 VDD.n3755 VDD.n3754 0.152939
R7371 VDD.n3756 VDD.n3755 0.152939
R7372 VDD.n3756 VDD.n271 0.152939
R7373 VDD.n3770 VDD.n271 0.152939
R7374 VDD.n3771 VDD.n3770 0.152939
R7375 VDD.n3772 VDD.n3771 0.152939
R7376 VDD.n3772 VDD.n269 0.152939
R7377 VDD.n3776 VDD.n269 0.152939
R7378 VDD.n3777 VDD.n3776 0.152939
R7379 VDD.n3778 VDD.n3777 0.152939
R7380 VDD.n3778 VDD.n266 0.152939
R7381 VDD.n3782 VDD.n266 0.152939
R7382 VDD.n3783 VDD.n3782 0.152939
R7383 VDD.n3784 VDD.n3783 0.152939
R7384 VDD.n3784 VDD.n263 0.152939
R7385 VDD.n3788 VDD.n263 0.152939
R7386 VDD.n3789 VDD.n3788 0.152939
R7387 VDD.n3790 VDD.n3789 0.152939
R7388 VDD.n3790 VDD.n260 0.152939
R7389 VDD.n3794 VDD.n260 0.152939
R7390 VDD.n3795 VDD.n3794 0.152939
R7391 VDD.n3796 VDD.n3795 0.152939
R7392 VDD.n3796 VDD.n257 0.152939
R7393 VDD.n3800 VDD.n257 0.152939
R7394 VDD.n3801 VDD.n3800 0.152939
R7395 VDD.n3802 VDD.n3801 0.152939
R7396 VDD.n3802 VDD.n254 0.152939
R7397 VDD.n3806 VDD.n254 0.152939
R7398 VDD.n3807 VDD.n3806 0.152939
R7399 VDD.n3808 VDD.n3807 0.152939
R7400 VDD.n3808 VDD.n251 0.152939
R7401 VDD.n3812 VDD.n251 0.152939
R7402 VDD.n3813 VDD.n3812 0.152939
R7403 VDD.n3814 VDD.n3813 0.152939
R7404 VDD.n3814 VDD.n248 0.152939
R7405 VDD.n3818 VDD.n248 0.152939
R7406 VDD.n3819 VDD.n3818 0.152939
R7407 VDD.n3820 VDD.n3819 0.152939
R7408 VDD.n3820 VDD.n245 0.152939
R7409 VDD.n3824 VDD.n245 0.152939
R7410 VDD.n3825 VDD.n3824 0.152939
R7411 VDD.n3826 VDD.n3825 0.152939
R7412 VDD.n3826 VDD.n242 0.152939
R7413 VDD.n3830 VDD.n242 0.152939
R7414 VDD.n3831 VDD.n3830 0.152939
R7415 VDD.n3832 VDD.n3831 0.152939
R7416 VDD.n3832 VDD.n239 0.152939
R7417 VDD.n3836 VDD.n239 0.152939
R7418 VDD.n1595 VDD.n1594 0.152939
R7419 VDD.n1595 VDD.n1434 0.152939
R7420 VDD.n1609 VDD.n1434 0.152939
R7421 VDD.n1610 VDD.n1609 0.152939
R7422 VDD.n1611 VDD.n1610 0.152939
R7423 VDD.n1611 VDD.n1423 0.152939
R7424 VDD.n1625 VDD.n1423 0.152939
R7425 VDD.n1626 VDD.n1625 0.152939
R7426 VDD.n1627 VDD.n1626 0.152939
R7427 VDD.n1627 VDD.n1411 0.152939
R7428 VDD.n1641 VDD.n1411 0.152939
R7429 VDD.n1642 VDD.n1641 0.152939
R7430 VDD.n1643 VDD.n1642 0.152939
R7431 VDD.n1643 VDD.n1400 0.152939
R7432 VDD.n1658 VDD.n1400 0.152939
R7433 VDD.n1659 VDD.n1658 0.152939
R7434 VDD.n1660 VDD.n1659 0.152939
R7435 VDD.n1660 VDD.n1388 0.152939
R7436 VDD.n1674 VDD.n1388 0.152939
R7437 VDD.n1675 VDD.n1674 0.152939
R7438 VDD.n1676 VDD.n1675 0.152939
R7439 VDD.n1676 VDD.n1377 0.152939
R7440 VDD.n1691 VDD.n1377 0.152939
R7441 VDD.n1692 VDD.n1691 0.152939
R7442 VDD.n1693 VDD.n1692 0.152939
R7443 VDD.n1693 VDD.n1365 0.152939
R7444 VDD.n1707 VDD.n1365 0.152939
R7445 VDD.n1708 VDD.n1707 0.152939
R7446 VDD.n1709 VDD.n1708 0.152939
R7447 VDD.n1709 VDD.n1354 0.152939
R7448 VDD.n1724 VDD.n1354 0.152939
R7449 VDD.n1725 VDD.n1724 0.152939
R7450 VDD.n1726 VDD.n1725 0.152939
R7451 VDD.n1726 VDD.n1342 0.152939
R7452 VDD.n1740 VDD.n1342 0.152939
R7453 VDD.n1741 VDD.n1740 0.152939
R7454 VDD.n1742 VDD.n1741 0.152939
R7455 VDD.n1742 VDD.n1331 0.152939
R7456 VDD.n1757 VDD.n1331 0.152939
R7457 VDD.n1758 VDD.n1757 0.152939
R7458 VDD.n1759 VDD.n1758 0.152939
R7459 VDD.n1759 VDD.n1319 0.152939
R7460 VDD.n1805 VDD.n1319 0.152939
R7461 VDD.n1806 VDD.n1805 0.152939
R7462 VDD.n1807 VDD.n1806 0.152939
R7463 VDD.n1807 VDD.n1307 0.152939
R7464 VDD.n1821 VDD.n1307 0.152939
R7465 VDD.n1822 VDD.n1821 0.152939
R7466 VDD.n1823 VDD.n1822 0.152939
R7467 VDD.n1823 VDD.n1295 0.152939
R7468 VDD.n1837 VDD.n1295 0.152939
R7469 VDD.n1838 VDD.n1837 0.152939
R7470 VDD.n1839 VDD.n1838 0.152939
R7471 VDD.n1839 VDD.n1283 0.152939
R7472 VDD.n1853 VDD.n1283 0.152939
R7473 VDD.n1854 VDD.n1853 0.152939
R7474 VDD.n1855 VDD.n1854 0.152939
R7475 VDD.n1855 VDD.n1271 0.152939
R7476 VDD.n1869 VDD.n1271 0.152939
R7477 VDD.n1870 VDD.n1869 0.152939
R7478 VDD.n1871 VDD.n1870 0.152939
R7479 VDD.n1871 VDD.n1259 0.152939
R7480 VDD.n1885 VDD.n1259 0.152939
R7481 VDD.n1886 VDD.n1885 0.152939
R7482 VDD.n1887 VDD.n1886 0.152939
R7483 VDD.n1887 VDD.n1247 0.152939
R7484 VDD.n1901 VDD.n1247 0.152939
R7485 VDD.n1902 VDD.n1901 0.152939
R7486 VDD.n1903 VDD.n1902 0.152939
R7487 VDD.n1903 VDD.n1235 0.152939
R7488 VDD.n1917 VDD.n1235 0.152939
R7489 VDD.n1918 VDD.n1917 0.152939
R7490 VDD.n1919 VDD.n1918 0.152939
R7491 VDD.n1919 VDD.n1223 0.152939
R7492 VDD.n1933 VDD.n1223 0.152939
R7493 VDD.n1934 VDD.n1933 0.152939
R7494 VDD.n1935 VDD.n1934 0.152939
R7495 VDD.n1935 VDD.n1211 0.152939
R7496 VDD.n1949 VDD.n1211 0.152939
R7497 VDD.n1950 VDD.n1949 0.152939
R7498 VDD.n1952 VDD.n1950 0.152939
R7499 VDD.n1952 VDD.n1951 0.152939
R7500 VDD.n1951 VDD.n1199 0.152939
R7501 VDD.n1968 VDD.n1199 0.152939
R7502 VDD.n1584 VDD.n1470 0.152939
R7503 VDD.n1584 VDD.n1583 0.152939
R7504 VDD.n1583 VDD.n1582 0.152939
R7505 VDD.n1582 VDD.n1472 0.152939
R7506 VDD.n1578 VDD.n1472 0.152939
R7507 VDD.n1578 VDD.n1577 0.152939
R7508 VDD.n1577 VDD.n1576 0.152939
R7509 VDD.n1576 VDD.n1477 0.152939
R7510 VDD.n1568 VDD.n1477 0.152939
R7511 VDD.n1568 VDD.n1567 0.152939
R7512 VDD.n1567 VDD.n1566 0.152939
R7513 VDD.n1566 VDD.n1481 0.152939
R7514 VDD.n1562 VDD.n1481 0.152939
R7515 VDD.n1562 VDD.n1561 0.152939
R7516 VDD.n1561 VDD.n1560 0.152939
R7517 VDD.n1560 VDD.n1487 0.152939
R7518 VDD.n1556 VDD.n1487 0.152939
R7519 VDD.n1556 VDD.n1555 0.152939
R7520 VDD.n1555 VDD.n1495 0.152939
R7521 VDD.n1551 VDD.n1495 0.152939
R7522 VDD.n1551 VDD.n1550 0.152939
R7523 VDD.n1550 VDD.n1549 0.152939
R7524 VDD.n1549 VDD.n1501 0.152939
R7525 VDD.n1545 VDD.n1501 0.152939
R7526 VDD.n1545 VDD.n1544 0.152939
R7527 VDD.n1544 VDD.n1543 0.152939
R7528 VDD.n1543 VDD.n1507 0.152939
R7529 VDD.n1536 VDD.n1507 0.152939
R7530 VDD.n1536 VDD.n1535 0.152939
R7531 VDD.n1535 VDD.n1534 0.152939
R7532 VDD.n1534 VDD.n1513 0.152939
R7533 VDD.n1530 VDD.n1513 0.152939
R7534 VDD.n1530 VDD.n1529 0.152939
R7535 VDD.n1529 VDD.n1528 0.152939
R7536 VDD.n1528 VDD.n1519 0.152939
R7537 VDD.n1524 VDD.n1519 0.152939
R7538 VDD.n1524 VDD.n1446 0.152939
R7539 VDD.n1593 VDD.n1446 0.152939
R7540 VDD.n1601 VDD.n1440 0.152939
R7541 VDD.n1602 VDD.n1601 0.152939
R7542 VDD.n1603 VDD.n1602 0.152939
R7543 VDD.n1603 VDD.n1429 0.152939
R7544 VDD.n1617 VDD.n1429 0.152939
R7545 VDD.n1618 VDD.n1617 0.152939
R7546 VDD.n1619 VDD.n1618 0.152939
R7547 VDD.n1619 VDD.n1417 0.152939
R7548 VDD.n1633 VDD.n1417 0.152939
R7549 VDD.n1634 VDD.n1633 0.152939
R7550 VDD.n1635 VDD.n1634 0.152939
R7551 VDD.n1635 VDD.n1405 0.152939
R7552 VDD.n1650 VDD.n1405 0.152939
R7553 VDD.n1651 VDD.n1650 0.152939
R7554 VDD.n1652 VDD.n1651 0.152939
R7555 VDD.n1652 VDD.n1394 0.152939
R7556 VDD.n1666 VDD.n1394 0.152939
R7557 VDD.n1667 VDD.n1666 0.152939
R7558 VDD.n1668 VDD.n1667 0.152939
R7559 VDD.n1668 VDD.n1382 0.152939
R7560 VDD.n1683 VDD.n1382 0.152939
R7561 VDD.n1684 VDD.n1683 0.152939
R7562 VDD.n1685 VDD.n1684 0.152939
R7563 VDD.n1685 VDD.n1371 0.152939
R7564 VDD.n1699 VDD.n1371 0.152939
R7565 VDD.n1700 VDD.n1699 0.152939
R7566 VDD.n1701 VDD.n1700 0.152939
R7567 VDD.n1701 VDD.n1359 0.152939
R7568 VDD.n1716 VDD.n1359 0.152939
R7569 VDD.n1717 VDD.n1716 0.152939
R7570 VDD.n1718 VDD.n1717 0.152939
R7571 VDD.n1718 VDD.n1348 0.152939
R7572 VDD.n1732 VDD.n1348 0.152939
R7573 VDD.n1733 VDD.n1732 0.152939
R7574 VDD.n1734 VDD.n1733 0.152939
R7575 VDD.n1734 VDD.n1336 0.152939
R7576 VDD.n1749 VDD.n1336 0.152939
R7577 VDD.n1750 VDD.n1749 0.152939
R7578 VDD.n1751 VDD.n1750 0.152939
R7579 VDD.n1751 VDD.n1325 0.152939
R7580 VDD.n1765 VDD.n1325 0.152939
R7581 VDD.n1799 VDD.n1798 0.145814
R7582 VDD.n4000 VDD.n47 0.145814
R7583 VDD.n4000 VDD.n48 0.145814
R7584 VDD.n1798 VDD.n1765 0.145814
R7585 VDD.n2168 VDD.n1137 0.119402
R7586 VDD.n2080 VDD.n1197 0.119402
R7587 VDD.n3604 VDD.n396 0.119402
R7588 VDD.n3526 VDD.n392 0.119402
R7589 VDD VDD.n15 0.00833333
R7590 VOUT.n132 VOUT.n130 289.615
R7591 VOUT.n120 VOUT.n118 289.615
R7592 VOUT.n108 VOUT.n106 289.615
R7593 VOUT.n96 VOUT.n94 289.615
R7594 VOUT.n85 VOUT.n83 289.615
R7595 VOUT.n195 VOUT.n193 289.615
R7596 VOUT.n183 VOUT.n181 289.615
R7597 VOUT.n171 VOUT.n169 289.615
R7598 VOUT.n159 VOUT.n157 289.615
R7599 VOUT.n148 VOUT.n146 289.615
R7600 VOUT.n76 VOUT.n74 191.948
R7601 VOUT.n68 VOUT.n66 191.948
R7602 VOUT.n60 VOUT.n58 191.948
R7603 VOUT.n53 VOUT.n51 191.948
R7604 VOUT.n25 VOUT.n23 191.948
R7605 VOUT.n17 VOUT.n15 191.948
R7606 VOUT.n9 VOUT.n7 191.948
R7607 VOUT.n2 VOUT.n0 191.948
R7608 VOUT.n78 VOUT.n77 190.233
R7609 VOUT.n76 VOUT.n75 190.233
R7610 VOUT.n72 VOUT.n71 190.233
R7611 VOUT.n70 VOUT.n69 190.233
R7612 VOUT.n68 VOUT.n67 190.233
R7613 VOUT.n64 VOUT.n63 190.233
R7614 VOUT.n62 VOUT.n61 190.233
R7615 VOUT.n60 VOUT.n59 190.233
R7616 VOUT.n57 VOUT.n56 190.233
R7617 VOUT.n55 VOUT.n54 190.233
R7618 VOUT.n53 VOUT.n52 190.233
R7619 VOUT.n25 VOUT.n24 190.233
R7620 VOUT.n27 VOUT.n26 190.233
R7621 VOUT.n29 VOUT.n28 190.233
R7622 VOUT.n17 VOUT.n16 190.233
R7623 VOUT.n19 VOUT.n18 190.233
R7624 VOUT.n21 VOUT.n20 190.233
R7625 VOUT.n9 VOUT.n8 190.233
R7626 VOUT.n11 VOUT.n10 190.233
R7627 VOUT.n13 VOUT.n12 190.233
R7628 VOUT.n2 VOUT.n1 190.233
R7629 VOUT.n4 VOUT.n3 190.233
R7630 VOUT.n6 VOUT.n5 190.233
R7631 VOUT.n80 VOUT.n79 190.233
R7632 VOUT.n133 VOUT.n132 185
R7633 VOUT.n121 VOUT.n120 185
R7634 VOUT.n109 VOUT.n108 185
R7635 VOUT.n97 VOUT.n96 185
R7636 VOUT.n86 VOUT.n85 185
R7637 VOUT.n196 VOUT.n195 185
R7638 VOUT.n184 VOUT.n183 185
R7639 VOUT.n172 VOUT.n171 185
R7640 VOUT.n160 VOUT.n159 185
R7641 VOUT.n149 VOUT.n148 185
R7642 VOUT.t11 VOUT.n131 167.117
R7643 VOUT.t5 VOUT.n119 167.117
R7644 VOUT.t1 VOUT.n107 167.117
R7645 VOUT.t36 VOUT.n95 167.117
R7646 VOUT.t14 VOUT.n84 167.117
R7647 VOUT.t25 VOUT.n194 167.117
R7648 VOUT.t30 VOUT.n182 167.117
R7649 VOUT.t8 VOUT.n170 167.117
R7650 VOUT.t21 VOUT.n158 167.117
R7651 VOUT.t10 VOUT.n147 167.117
R7652 VOUT.n192 VOUT.n190 120.328
R7653 VOUT.n180 VOUT.n178 120.328
R7654 VOUT.n168 VOUT.n166 120.328
R7655 VOUT.n156 VOUT.n154 120.328
R7656 VOUT.n145 VOUT.n143 120.328
R7657 VOUT.n140 VOUT.n139 118.251
R7658 VOUT.n138 VOUT.n137 118.251
R7659 VOUT.n128 VOUT.n127 118.251
R7660 VOUT.n126 VOUT.n125 118.251
R7661 VOUT.n116 VOUT.n115 118.251
R7662 VOUT.n114 VOUT.n113 118.251
R7663 VOUT.n104 VOUT.n103 118.251
R7664 VOUT.n102 VOUT.n101 118.251
R7665 VOUT.n93 VOUT.n92 118.251
R7666 VOUT.n91 VOUT.n90 118.251
R7667 VOUT.n192 VOUT.n191 118.251
R7668 VOUT.n180 VOUT.n179 118.251
R7669 VOUT.n168 VOUT.n167 118.251
R7670 VOUT.n156 VOUT.n155 118.251
R7671 VOUT.n145 VOUT.n144 118.251
R7672 VOUT.n138 VOUT.n136 67.6205
R7673 VOUT.n126 VOUT.n124 67.6205
R7674 VOUT.n114 VOUT.n112 67.6205
R7675 VOUT.n102 VOUT.n100 67.6205
R7676 VOUT.n91 VOUT.n89 67.6205
R7677 VOUT.n200 VOUT.n199 65.5429
R7678 VOUT.n188 VOUT.n187 65.5429
R7679 VOUT.n176 VOUT.n175 65.5429
R7680 VOUT.n164 VOUT.n163 65.5429
R7681 VOUT.n153 VOUT.n152 65.5429
R7682 VOUT.n132 VOUT.t11 52.3082
R7683 VOUT.n120 VOUT.t5 52.3082
R7684 VOUT.n108 VOUT.t1 52.3082
R7685 VOUT.n96 VOUT.t36 52.3082
R7686 VOUT.n85 VOUT.t14 52.3082
R7687 VOUT.n195 VOUT.t25 52.3082
R7688 VOUT.n183 VOUT.t30 52.3082
R7689 VOUT.n171 VOUT.t8 52.3082
R7690 VOUT.n159 VOUT.t21 52.3082
R7691 VOUT.n148 VOUT.t10 52.3082
R7692 VOUT.n79 VOUT.t48 14.9798
R7693 VOUT.n79 VOUT.t91 14.9798
R7694 VOUT.n77 VOUT.t55 14.9798
R7695 VOUT.n77 VOUT.t82 14.9798
R7696 VOUT.n75 VOUT.t51 14.9798
R7697 VOUT.n75 VOUT.t79 14.9798
R7698 VOUT.n74 VOUT.t104 14.9798
R7699 VOUT.n74 VOUT.t77 14.9798
R7700 VOUT.n71 VOUT.t87 14.9798
R7701 VOUT.n71 VOUT.t67 14.9798
R7702 VOUT.n69 VOUT.t94 14.9798
R7703 VOUT.n69 VOUT.t56 14.9798
R7704 VOUT.n67 VOUT.t92 14.9798
R7705 VOUT.n67 VOUT.t53 14.9798
R7706 VOUT.n66 VOUT.t83 14.9798
R7707 VOUT.n66 VOUT.t49 14.9798
R7708 VOUT.n63 VOUT.t101 14.9798
R7709 VOUT.n63 VOUT.t78 14.9798
R7710 VOUT.n61 VOUT.t54 14.9798
R7711 VOUT.n61 VOUT.t107 14.9798
R7712 VOUT.n59 VOUT.t89 14.9798
R7713 VOUT.n59 VOUT.t81 14.9798
R7714 VOUT.n58 VOUT.t58 14.9798
R7715 VOUT.n58 VOUT.t52 14.9798
R7716 VOUT.n56 VOUT.t59 14.9798
R7717 VOUT.n56 VOUT.t97 14.9798
R7718 VOUT.n54 VOUT.t74 14.9798
R7719 VOUT.n54 VOUT.t62 14.9798
R7720 VOUT.n52 VOUT.t45 14.9798
R7721 VOUT.n52 VOUT.t100 14.9798
R7722 VOUT.n51 VOUT.t80 14.9798
R7723 VOUT.n51 VOUT.t73 14.9798
R7724 VOUT.n23 VOUT.t95 14.9798
R7725 VOUT.n23 VOUT.t70 14.9798
R7726 VOUT.n24 VOUT.t47 14.9798
R7727 VOUT.n24 VOUT.t64 14.9798
R7728 VOUT.n26 VOUT.t65 14.9798
R7729 VOUT.n26 VOUT.t86 14.9798
R7730 VOUT.n28 VOUT.t60 14.9798
R7731 VOUT.n28 VOUT.t90 14.9798
R7732 VOUT.n15 VOUT.t71 14.9798
R7733 VOUT.n15 VOUT.t44 14.9798
R7734 VOUT.n16 VOUT.t85 14.9798
R7735 VOUT.n16 VOUT.t102 14.9798
R7736 VOUT.n18 VOUT.t106 14.9798
R7737 VOUT.n18 VOUT.t63 14.9798
R7738 VOUT.n20 VOUT.t99 14.9798
R7739 VOUT.n20 VOUT.t66 14.9798
R7740 VOUT.n7 VOUT.t105 14.9798
R7741 VOUT.n7 VOUT.t50 14.9798
R7742 VOUT.n8 VOUT.t75 14.9798
R7743 VOUT.n8 VOUT.t98 14.9798
R7744 VOUT.n10 VOUT.t84 14.9798
R7745 VOUT.n10 VOUT.t46 14.9798
R7746 VOUT.n12 VOUT.t69 14.9798
R7747 VOUT.n12 VOUT.t76 14.9798
R7748 VOUT.n0 VOUT.t61 14.9798
R7749 VOUT.n0 VOUT.t72 14.9798
R7750 VOUT.n1 VOUT.t93 14.9798
R7751 VOUT.n1 VOUT.t57 14.9798
R7752 VOUT.n3 VOUT.t103 14.9798
R7753 VOUT.n3 VOUT.t68 14.9798
R7754 VOUT.n5 VOUT.t88 14.9798
R7755 VOUT.n5 VOUT.t96 14.9798
R7756 VOUT.n139 VOUT.t110 9.75419
R7757 VOUT.n139 VOUT.t27 9.75419
R7758 VOUT.n137 VOUT.t40 9.75419
R7759 VOUT.n137 VOUT.t24 9.75419
R7760 VOUT.n127 VOUT.t31 9.75419
R7761 VOUT.n127 VOUT.t43 9.75419
R7762 VOUT.n125 VOUT.t17 9.75419
R7763 VOUT.n125 VOUT.t19 9.75419
R7764 VOUT.n115 VOUT.t2 9.75419
R7765 VOUT.n115 VOUT.t4 9.75419
R7766 VOUT.n113 VOUT.t32 9.75419
R7767 VOUT.n113 VOUT.t28 9.75419
R7768 VOUT.n103 VOUT.t12 9.75419
R7769 VOUT.n103 VOUT.t42 9.75419
R7770 VOUT.n101 VOUT.t23 9.75419
R7771 VOUT.n101 VOUT.t37 9.75419
R7772 VOUT.n92 VOUT.t108 9.75419
R7773 VOUT.n92 VOUT.t26 9.75419
R7774 VOUT.n90 VOUT.t15 9.75419
R7775 VOUT.n90 VOUT.t33 9.75419
R7776 VOUT.n190 VOUT.t113 9.75419
R7777 VOUT.n190 VOUT.t29 9.75419
R7778 VOUT.n191 VOUT.t39 9.75419
R7779 VOUT.n191 VOUT.t13 9.75419
R7780 VOUT.n178 VOUT.t18 9.75419
R7781 VOUT.n178 VOUT.t111 9.75419
R7782 VOUT.n179 VOUT.t35 9.75419
R7783 VOUT.n179 VOUT.t6 9.75419
R7784 VOUT.n166 VOUT.t34 9.75419
R7785 VOUT.n166 VOUT.t9 9.75419
R7786 VOUT.n167 VOUT.t109 9.75419
R7787 VOUT.n167 VOUT.t16 9.75419
R7788 VOUT.n154 VOUT.t112 9.75419
R7789 VOUT.n154 VOUT.t41 9.75419
R7790 VOUT.n155 VOUT.t38 9.75419
R7791 VOUT.n155 VOUT.t0 9.75419
R7792 VOUT.n143 VOUT.t20 9.75419
R7793 VOUT.n143 VOUT.t22 9.75419
R7794 VOUT.n144 VOUT.t3 9.75419
R7795 VOUT.n144 VOUT.t7 9.75419
R7796 VOUT.n133 VOUT.n131 9.71174
R7797 VOUT.n121 VOUT.n119 9.71174
R7798 VOUT.n109 VOUT.n107 9.71174
R7799 VOUT.n97 VOUT.n95 9.71174
R7800 VOUT.n86 VOUT.n84 9.71174
R7801 VOUT.n196 VOUT.n194 9.71174
R7802 VOUT.n184 VOUT.n182 9.71174
R7803 VOUT.n172 VOUT.n170 9.71174
R7804 VOUT.n160 VOUT.n158 9.71174
R7805 VOUT.n149 VOUT.n147 9.71174
R7806 VOUT.n136 VOUT.n135 9.45567
R7807 VOUT.n124 VOUT.n123 9.45567
R7808 VOUT.n112 VOUT.n111 9.45567
R7809 VOUT.n100 VOUT.n99 9.45567
R7810 VOUT.n89 VOUT.n88 9.45567
R7811 VOUT.n199 VOUT.n198 9.45567
R7812 VOUT.n187 VOUT.n186 9.45567
R7813 VOUT.n175 VOUT.n174 9.45567
R7814 VOUT.n163 VOUT.n162 9.45567
R7815 VOUT.n152 VOUT.n151 9.45567
R7816 VOUT.n135 VOUT.n134 9.3005
R7817 VOUT.n123 VOUT.n122 9.3005
R7818 VOUT.n111 VOUT.n110 9.3005
R7819 VOUT.n99 VOUT.n98 9.3005
R7820 VOUT.n88 VOUT.n87 9.3005
R7821 VOUT.n198 VOUT.n197 9.3005
R7822 VOUT.n186 VOUT.n185 9.3005
R7823 VOUT.n174 VOUT.n173 9.3005
R7824 VOUT.n162 VOUT.n161 9.3005
R7825 VOUT.n151 VOUT.n150 9.3005
R7826 VOUT.n142 VOUT.n82 8.49284
R7827 VOUT.n136 VOUT.n130 8.14595
R7828 VOUT.n124 VOUT.n118 8.14595
R7829 VOUT.n112 VOUT.n106 8.14595
R7830 VOUT.n100 VOUT.n94 8.14595
R7831 VOUT.n89 VOUT.n83 8.14595
R7832 VOUT.n199 VOUT.n193 8.14595
R7833 VOUT.n187 VOUT.n181 8.14595
R7834 VOUT.n175 VOUT.n169 8.14595
R7835 VOUT.n163 VOUT.n157 8.14595
R7836 VOUT.n152 VOUT.n146 8.14595
R7837 VOUT.n134 VOUT.n133 7.3702
R7838 VOUT.n122 VOUT.n121 7.3702
R7839 VOUT.n110 VOUT.n109 7.3702
R7840 VOUT.n98 VOUT.n97 7.3702
R7841 VOUT.n87 VOUT.n86 7.3702
R7842 VOUT.n197 VOUT.n196 7.3702
R7843 VOUT.n185 VOUT.n184 7.3702
R7844 VOUT.n173 VOUT.n172 7.3702
R7845 VOUT.n161 VOUT.n160 7.3702
R7846 VOUT.n150 VOUT.n149 7.3702
R7847 VOUT.n105 VOUT.n93 7.05653
R7848 VOUT.n65 VOUT.n57 6.90567
R7849 VOUT.n14 VOUT.n6 6.90567
R7850 VOUT.n165 VOUT.n153 6.01774
R7851 VOUT.n141 VOUT.n140 6.00481
R7852 VOUT.n129 VOUT.n128 6.00481
R7853 VOUT.n117 VOUT.n116 6.00481
R7854 VOUT.n105 VOUT.n104 6.00481
R7855 VOUT.n81 VOUT.n80 5.82378
R7856 VOUT.n73 VOUT.n72 5.82378
R7857 VOUT.n65 VOUT.n64 5.82378
R7858 VOUT.n30 VOUT.n29 5.82378
R7859 VOUT.n22 VOUT.n21 5.82378
R7860 VOUT.n14 VOUT.n13 5.82378
R7861 VOUT.n134 VOUT.n130 5.81868
R7862 VOUT.n122 VOUT.n118 5.81868
R7863 VOUT.n110 VOUT.n106 5.81868
R7864 VOUT.n98 VOUT.n94 5.81868
R7865 VOUT.n87 VOUT.n83 5.81868
R7866 VOUT.n197 VOUT.n193 5.81868
R7867 VOUT.n185 VOUT.n181 5.81868
R7868 VOUT.n173 VOUT.n169 5.81868
R7869 VOUT.n161 VOUT.n157 5.81868
R7870 VOUT.n150 VOUT.n146 5.81868
R7871 VOUT.n82 VOUT.n81 5.76287
R7872 VOUT.n31 VOUT.n30 5.76287
R7873 VOUT.n82 VOUT.n31 5.38012
R7874 VOUT.n202 VOUT.n142 5.31714
R7875 VOUT.n142 VOUT.n141 5.00748
R7876 VOUT.n202 VOUT.n201 5.00748
R7877 VOUT.n201 VOUT.n200 4.96602
R7878 VOUT.n189 VOUT.n188 4.96602
R7879 VOUT.n177 VOUT.n176 4.96602
R7880 VOUT.n165 VOUT.n164 4.96602
R7881 VOUT.n203 VOUT.n31 4.78447
R7882 VOUT.n50 VOUT 4.02605
R7883 VOUT.n203 VOUT.n202 3.68937
R7884 VOUT.n135 VOUT.n131 3.44771
R7885 VOUT.n123 VOUT.n119 3.44771
R7886 VOUT.n111 VOUT.n107 3.44771
R7887 VOUT.n99 VOUT.n95 3.44771
R7888 VOUT.n88 VOUT.n84 3.44771
R7889 VOUT.n198 VOUT.n194 3.44771
R7890 VOUT.n186 VOUT.n182 3.44771
R7891 VOUT.n174 VOUT.n170 3.44771
R7892 VOUT.n162 VOUT.n158 3.44771
R7893 VOUT.n151 VOUT.n147 3.44771
R7894 VOUT.n140 VOUT.n138 2.07809
R7895 VOUT.n128 VOUT.n126 2.07809
R7896 VOUT.n116 VOUT.n114 2.07809
R7897 VOUT.n104 VOUT.n102 2.07809
R7898 VOUT.n93 VOUT.n91 2.07809
R7899 VOUT.n200 VOUT.n192 2.07809
R7900 VOUT.n188 VOUT.n180 2.07809
R7901 VOUT.n176 VOUT.n168 2.07809
R7902 VOUT.n164 VOUT.n156 2.07809
R7903 VOUT.n153 VOUT.n145 2.07809
R7904 VOUT.n78 VOUT.n76 1.71602
R7905 VOUT.n80 VOUT.n78 1.71602
R7906 VOUT.n70 VOUT.n68 1.71602
R7907 VOUT.n72 VOUT.n70 1.71602
R7908 VOUT.n62 VOUT.n60 1.71602
R7909 VOUT.n64 VOUT.n62 1.71602
R7910 VOUT.n55 VOUT.n53 1.71602
R7911 VOUT.n57 VOUT.n55 1.71602
R7912 VOUT.n29 VOUT.n27 1.71602
R7913 VOUT.n27 VOUT.n25 1.71602
R7914 VOUT.n21 VOUT.n19 1.71602
R7915 VOUT.n19 VOUT.n17 1.71602
R7916 VOUT.n13 VOUT.n11 1.71602
R7917 VOUT.n11 VOUT.n9 1.71602
R7918 VOUT.n6 VOUT.n4 1.71602
R7919 VOUT.n4 VOUT.n2 1.71602
R7920 VOUT.n81 VOUT.n73 1.0824
R7921 VOUT.n73 VOUT.n65 1.0824
R7922 VOUT.n30 VOUT.n22 1.0824
R7923 VOUT.n22 VOUT.n14 1.0824
R7924 VOUT.n141 VOUT.n129 1.05222
R7925 VOUT.n129 VOUT.n117 1.05222
R7926 VOUT.n117 VOUT.n105 1.05222
R7927 VOUT.n201 VOUT.n189 1.05222
R7928 VOUT.n189 VOUT.n177 1.05222
R7929 VOUT.n177 VOUT.n165 1.05222
R7930 VOUT.n50 VOUT.n49 0.397402
R7931 VOUT.n203 VOUT.n50 0.393655
R7932 VOUT.n36 VOUT.n35 0.0825984
R7933 VOUT.n42 VOUT.n41 0.0819129
R7934 VOUT.n44 VOUT.n43 0.0819129
R7935 VOUT.n39 VOUT.n38 0.0779202
R7936 VOUT.n46 VOUT.n45 0.0779202
R7937 VOUT.n48 VOUT.n47 0.0779202
R7938 VOUT.n43 VOUT.n42 0.0659614
R7939 VOUT.n35 VOUT.n32 0.0474378
R7940 VOUT.n40 VOUT.n34 0.0391444
R7941 VOUT.n37 VOUT.n33 0.0391444
R7942 VOUT.n36 VOUT.t120 0.0219306
R7943 VOUT.n39 VOUT.t121 0.0219306
R7944 VOUT.n45 VOUT.t117 0.0219306
R7945 VOUT.n47 VOUT.t116 0.0219306
R7946 VOUT.n49 VOUT.t119 0.0219306
R7947 VOUT.n38 VOUT.t120 0.0219025
R7948 VOUT.n41 VOUT.t121 0.0219025
R7949 VOUT.t117 VOUT.n44 0.0219025
R7950 VOUT.t116 VOUT.n46 0.0219025
R7951 VOUT.t119 VOUT.n48 0.0219025
R7952 VOUT.n37 VOUT.n36 0.0199893
R7953 VOUT.n40 VOUT.n39 0.0199893
R7954 VOUT.n45 VOUT.n34 0.0199893
R7955 VOUT.n47 VOUT.n33 0.0199893
R7956 VOUT.n49 VOUT.n32 0.0199893
R7957 VOUT.n38 VOUT.n37 0.0153757
R7958 VOUT.n41 VOUT.n40 0.0153757
R7959 VOUT.n44 VOUT.n34 0.0153757
R7960 VOUT.n46 VOUT.n33 0.0153757
R7961 VOUT.n48 VOUT.n32 0.0153757
R7962 VOUT.n42 VOUT.t118 0.0127855
R7963 VOUT.n43 VOUT.t115 0.0127855
R7964 VOUT.n35 VOUT.t114 0.0122127
R7965 VOUT VOUT.n203 0.0099
R7966 a_n7183_9410.n26 a_n7183_9410.n5 4.70021
R7967 a_n7183_9410.n25 a_n7183_9410.n7 4.70021
R7968 a_n7183_9410.n24 a_n7183_9410.n10 4.70021
R7969 a_n7183_9410.n23 a_n7183_9410.t18 94.727
R7970 a_n7183_9410.n22 a_n7183_9410.t20 93.0149
R7971 a_n7183_9410.n28 a_n7183_9410.t3 91.746
R7972 a_n7183_9410.n22 a_n7183_9410.t9 88.817
R7973 a_n7183_9410.n14 a_n7183_9410.t1 88.4228
R7974 a_n7183_9410.t7 a_n7183_9410.n23 87.1058
R7975 a_n7183_9410.n22 a_n7183_9410.t16 87.1058
R7976 a_n7183_9410.n23 a_n7183_9410.t11 87.1058
R7977 a_n7183_9410.n29 a_n7183_9410.n4 65.6103
R7978 a_n7183_9410.n20 a_n7183_9410.t28 69.0423
R7979 a_n7183_9410.n30 a_n7183_9410.t44 36.4153
R7980 a_n7183_9410.n31 a_n7183_9410.t35 36.4153
R7981 a_n7183_9410.n11 a_n7183_9410.t25 65.3077
R7982 a_n7183_9410.n10 a_n7183_9410.t43 69.0428
R7983 a_n7183_9410.n3 a_n7183_9410.t14 69.0427
R7984 a_n7183_9410.n4 a_n7183_9410.t6 64.7454
R7985 a_n7183_9410.n29 a_n7183_9410.t13 36.4153
R7986 a_n7183_9410.n9 a_n7183_9410.t10 64.8582
R7987 a_n7183_9410.n3 a_n7183_9410.t17 69.0428
R7988 a_n7183_9410.n19 a_n7183_9410.t12 69.0423
R7989 a_n7183_9410.n34 a_n7183_9410.t8 36.4153
R7990 a_n7183_9410.n35 a_n7183_9410.t15 36.4153
R7991 a_n7183_9410.n8 a_n7183_9410.t21 65.3077
R7992 a_n7183_9410.n7 a_n7183_9410.t19 69.0428
R7993 a_n7183_9410.n18 a_n7183_9410.t37 69.0423
R7994 a_n7183_9410.n32 a_n7183_9410.t38 36.4153
R7995 a_n7183_9410.n33 a_n7183_9410.t30 36.4153
R7996 a_n7183_9410.n6 a_n7183_9410.t33 65.3077
R7997 a_n7183_9410.n5 a_n7183_9410.t34 69.0428
R7998 a_n7183_9410.n16 a_n7183_9410.t39 69.157
R7999 a_n7183_9410.n38 a_n7183_9410.t36 36.4153
R8000 a_n7183_9410.n13 a_n7183_9410.t27 66.1425
R8001 a_n7183_9410.n0 a_n7183_9410.t24 69.1575
R8002 a_n7183_9410.n0 a_n7183_9410.t22 69.157
R8003 a_n7183_9410.n2 a_n7183_9410.t45 69.8501
R8004 a_n7183_9410.n2 a_n7183_9410.t29 65.9734
R8005 a_n7183_9410.n0 a_n7183_9410.t26 69.1575
R8006 a_n7183_9410.n17 a_n7183_9410.t46 69.157
R8007 a_n7183_9410.n37 a_n7183_9410.t31 36.4153
R8008 a_n7183_9410.n12 a_n7183_9410.t41 66.1425
R8009 a_n7183_9410.n0 a_n7183_9410.t32 69.1575
R8010 a_n7183_9410.n21 a_n7183_9410.t40 69.157
R8011 a_n7183_9410.n36 a_n7183_9410.t47 36.4153
R8012 a_n7183_9410.n1 a_n7183_9410.t23 66.1425
R8013 a_n7183_9410.n0 a_n7183_9410.t42 69.1575
R8014 a_n7183_9410.n20 a_n7183_9410.n30 64.1735
R8015 a_n7183_9410.n30 a_n7183_9410.n24 59.3274
R8016 a_n7183_9410.n24 a_n7183_9410.n31 60.8029
R8017 a_n7183_9410.n31 a_n7183_9410.n11 64.5284
R8018 a_n7183_9410.n11 a_n7183_9410.n10 4.03027
R8019 a_n7183_9410.n29 a_n7183_9410.n9 65.3935
R8020 a_n7183_9410.n9 a_n7183_9410.n3 4.966
R8021 a_n7183_9410.n34 a_n7183_9410.n19 64.1735
R8022 a_n7183_9410.n25 a_n7183_9410.n34 59.3274
R8023 a_n7183_9410.n35 a_n7183_9410.n25 60.8029
R8024 a_n7183_9410.n8 a_n7183_9410.n35 64.5284
R8025 a_n7183_9410.n7 a_n7183_9410.n8 4.03027
R8026 a_n7183_9410.n32 a_n7183_9410.n18 64.1735
R8027 a_n7183_9410.n26 a_n7183_9410.n32 59.3274
R8028 a_n7183_9410.n33 a_n7183_9410.n26 60.8029
R8029 a_n7183_9410.n6 a_n7183_9410.n33 64.5284
R8030 a_n7183_9410.n5 a_n7183_9410.n6 4.03027
R8031 a_n7183_9410.n38 a_n7183_9410.n16 63.4599
R8032 a_n7183_9410.n13 a_n7183_9410.n38 62.2672
R8033 a_n7183_9410.n37 a_n7183_9410.n17 63.4599
R8034 a_n7183_9410.n12 a_n7183_9410.n37 62.2672
R8035 a_n7183_9410.n36 a_n7183_9410.n21 63.4599
R8036 a_n7183_9410.n1 a_n7183_9410.n36 62.2672
R8037 a_n7183_9410.n14 a_n7183_9410.t2 86.7989
R8038 a_n7183_9410.n28 a_n7183_9410.t5 86.7987
R8039 a_n7183_9410.n14 a_n7183_9410.t4 84.3065
R8040 a_n7183_9410.n28 a_n7183_9410.t0 84.3062
R8041 a_n7183_9410.n0 a_n7183_9410.n1 2.32694
R8042 a_n7183_9410.n14 a_n7183_9410.n28 42.9755
R8043 a_n7183_9410.n5 a_n7183_9410.n27 14.2178
R8044 a_n7183_9410.n10 a_n7183_9410.n15 14.0133
R8045 a_n7183_9410.n4 a_n7183_9410.n3 5.19983
R8046 a_n7183_9410.n27 a_n7183_9410.n3 12.7084
R8047 a_n7183_9410.n15 a_n7183_9410.n22 11.7143
R8048 a_n7183_9410.n3 a_n7183_9410.n14 28.0748
R8049 a_n7183_9410.n15 a_n7183_9410.n0 11.0549
R8050 a_n7183_9410.n15 a_n7183_9410.n7 10.1989
R8051 a_n7183_9410.n0 a_n7183_9410.n2 10.187
R8052 a_n7183_9410.n23 a_n7183_9410.n27 10.0522
R8053 a_n7183_9410.n0 a_n7183_9410.n12 8.73495
R8054 a_n7183_9410.n0 a_n7183_9410.n27 8.34093
R8055 a_n7183_9410.n10 a_n7183_9410.n20 8.30785
R8056 a_n7183_9410.n7 a_n7183_9410.n19 8.30785
R8057 a_n7183_9410.n5 a_n7183_9410.n18 8.30785
R8058 a_n7183_9410.n0 a_n7183_9410.n21 8.25951
R8059 a_n7183_9410.n0 a_n7183_9410.n13 7.95939
R8060 a_n7183_9410.n17 a_n7183_9410.n0 7.69185
R8061 a_n7183_9410.n16 a_n7183_9410.n0 7.37442
R8062 a_n7183_9410.n7 a_n7183_9410.n5 6.90107
R8063 a_n7183_9410.n3 a_n7183_9410.n10 6.90107
R8064 a_n7261_9606.n13 a_n7261_9606.t17 122.654
R8065 a_n7261_9606.n2 a_n7261_9606.t9 121.642
R8066 a_n7261_9606.n4 a_n7261_9606.n3 115.034
R8067 a_n7261_9606.n2 a_n7261_9606.n1 115.034
R8068 a_n7261_9606.n14 a_n7261_9606.n13 115.034
R8069 a_n7261_9606.n12 a_n7261_9606.n11 115.032
R8070 a_n7261_9606.n6 a_n7261_9606.t7 94.727
R8071 a_n7261_9606.n9 a_n7261_9606.t6 93.0158
R8072 a_n7261_9606.n0 a_n7261_9606.t1 93.0158
R8073 a_n7261_9606.n0 a_n7261_9606.t5 93.0158
R8074 a_n7261_9606.n8 a_n7261_9606.n7 87.1058
R8075 a_n7261_9606.n6 a_n7261_9606.n5 87.1058
R8076 a_n7261_9606.n10 a_n7261_9606.n4 18.9058
R8077 a_n7261_9606.n12 a_n7261_9606.n10 12.7547
R8078 a_n7261_9606.n11 a_n7261_9606.t14 5.9105
R8079 a_n7261_9606.n11 a_n7261_9606.t11 5.9105
R8080 a_n7261_9606.n7 a_n7261_9606.t2 5.9105
R8081 a_n7261_9606.n7 a_n7261_9606.t4 5.9105
R8082 a_n7261_9606.n5 a_n7261_9606.t0 5.9105
R8083 a_n7261_9606.n5 a_n7261_9606.t3 5.9105
R8084 a_n7261_9606.n3 a_n7261_9606.t12 5.9105
R8085 a_n7261_9606.n3 a_n7261_9606.t10 5.9105
R8086 a_n7261_9606.n1 a_n7261_9606.t8 5.9105
R8087 a_n7261_9606.n1 a_n7261_9606.t13 5.9105
R8088 a_n7261_9606.t16 a_n7261_9606.n14 5.9105
R8089 a_n7261_9606.n14 a_n7261_9606.t15 5.9105
R8090 a_n7261_9606.n10 a_n7261_9606.n9 5.86149
R8091 a_n7261_9606.n8 a_n7261_9606.n0 2.14921
R8092 a_n7261_9606.n0 a_n7261_9606.n6 1.71171
R8093 a_n7261_9606.n9 a_n7261_9606.n8 1.71171
R8094 a_n7261_9606.n13 a_n7261_9606.n12 1.71171
R8095 a_n7261_9606.n4 a_n7261_9606.n2 0.699444
R8096 GND.n3937 GND.n3936 2183.74
R8097 GND.n4128 GND.n2152 1631.62
R8098 GND.n6919 GND.n1079 812.024
R8099 GND.n6972 GND.n6971 812.024
R8100 GND.n6110 GND.n1566 812.024
R8101 GND.n6098 GND.n1568 812.024
R8102 GND.n8462 GND.n347 759.172
R8103 GND.n8449 GND.n345 759.172
R8104 GND.n7736 GND.n659 759.172
R8105 GND.n695 GND.n651 759.172
R8106 GND.n4344 GND.n2134 759.172
R8107 GND.n6045 GND.n6044 759.172
R8108 GND.n4314 GND.n2132 759.172
R8109 GND.n1642 GND.n1609 759.172
R8110 GND.n3935 GND.n2248 723.135
R8111 GND.n3213 GND.n2965 723.135
R8112 GND.n8264 GND.n383 723.135
R8113 GND.n4127 GND.n2154 723.135
R8114 GND.n8464 GND.n342 660.672
R8115 GND.n8342 GND.n344 660.672
R8116 GND.n7738 GND.n657 660.672
R8117 GND.n7723 GND.n646 660.672
R8118 GND.n5905 GND.n1608 660.672
R8119 GND.n6047 GND.n1606 660.672
R8120 GND.n4214 GND.n2131 660.672
R8121 GND.n4346 GND.n2129 660.672
R8122 GND.n695 GND.n662 589.749
R8123 GND.n6044 GND.n1596 589.749
R8124 GND.n1642 GND.n1600 587.591
R8125 GND.n7730 GND.n659 587.591
R8126 GND.n2248 GND.n2247 585
R8127 GND.n3937 GND.n2248 585
R8128 GND.n3940 GND.n3939 585
R8129 GND.n3939 GND.n3938 585
R8130 GND.n2245 GND.n2244 585
R8131 GND.n2244 GND.n2243 585
R8132 GND.n3945 GND.n3944 585
R8133 GND.n3946 GND.n3945 585
R8134 GND.n2242 GND.n2241 585
R8135 GND.n3947 GND.n2242 585
R8136 GND.n3950 GND.n3949 585
R8137 GND.n3949 GND.n3948 585
R8138 GND.n2239 GND.n2238 585
R8139 GND.n2238 GND.n2237 585
R8140 GND.n3955 GND.n3954 585
R8141 GND.n3956 GND.n3955 585
R8142 GND.n2236 GND.n2235 585
R8143 GND.n3957 GND.n2236 585
R8144 GND.n3960 GND.n3959 585
R8145 GND.n3959 GND.n3958 585
R8146 GND.n2233 GND.n2232 585
R8147 GND.n2232 GND.n2231 585
R8148 GND.n3965 GND.n3964 585
R8149 GND.n3966 GND.n3965 585
R8150 GND.n2230 GND.n2229 585
R8151 GND.n3967 GND.n2230 585
R8152 GND.n3970 GND.n3969 585
R8153 GND.n3969 GND.n3968 585
R8154 GND.n2227 GND.n2226 585
R8155 GND.n2226 GND.n2225 585
R8156 GND.n3975 GND.n3974 585
R8157 GND.n3976 GND.n3975 585
R8158 GND.n2224 GND.n2223 585
R8159 GND.n3977 GND.n2224 585
R8160 GND.n3980 GND.n3979 585
R8161 GND.n3979 GND.n3978 585
R8162 GND.n2221 GND.n2220 585
R8163 GND.n2220 GND.n2219 585
R8164 GND.n3985 GND.n3984 585
R8165 GND.n3986 GND.n3985 585
R8166 GND.n2218 GND.n2217 585
R8167 GND.n3987 GND.n2218 585
R8168 GND.n3990 GND.n3989 585
R8169 GND.n3989 GND.n3988 585
R8170 GND.n2215 GND.n2214 585
R8171 GND.n2214 GND.n2213 585
R8172 GND.n3995 GND.n3994 585
R8173 GND.n3996 GND.n3995 585
R8174 GND.n2212 GND.n2211 585
R8175 GND.n3997 GND.n2212 585
R8176 GND.n4000 GND.n3999 585
R8177 GND.n3999 GND.n3998 585
R8178 GND.n2209 GND.n2208 585
R8179 GND.n2208 GND.n2207 585
R8180 GND.n4005 GND.n4004 585
R8181 GND.n4006 GND.n4005 585
R8182 GND.n2206 GND.n2205 585
R8183 GND.n4007 GND.n2206 585
R8184 GND.n4010 GND.n4009 585
R8185 GND.n4009 GND.n4008 585
R8186 GND.n2203 GND.n2202 585
R8187 GND.n2202 GND.n2201 585
R8188 GND.n4015 GND.n4014 585
R8189 GND.n4016 GND.n4015 585
R8190 GND.n2200 GND.n2199 585
R8191 GND.n4017 GND.n2200 585
R8192 GND.n4020 GND.n4019 585
R8193 GND.n4019 GND.n4018 585
R8194 GND.n2197 GND.n2196 585
R8195 GND.n2196 GND.n2195 585
R8196 GND.n4025 GND.n4024 585
R8197 GND.n4026 GND.n4025 585
R8198 GND.n2194 GND.n2193 585
R8199 GND.n4027 GND.n2194 585
R8200 GND.n4030 GND.n4029 585
R8201 GND.n4029 GND.n4028 585
R8202 GND.n2191 GND.n2190 585
R8203 GND.n2190 GND.n2189 585
R8204 GND.n4035 GND.n4034 585
R8205 GND.n4036 GND.n4035 585
R8206 GND.n2188 GND.n2187 585
R8207 GND.n4037 GND.n2188 585
R8208 GND.n4040 GND.n4039 585
R8209 GND.n4039 GND.n4038 585
R8210 GND.n2185 GND.n2184 585
R8211 GND.n2184 GND.n2183 585
R8212 GND.n4045 GND.n4044 585
R8213 GND.n4046 GND.n4045 585
R8214 GND.n2182 GND.n2181 585
R8215 GND.n4047 GND.n2182 585
R8216 GND.n4050 GND.n4049 585
R8217 GND.n4049 GND.n4048 585
R8218 GND.n2179 GND.n2178 585
R8219 GND.n2178 GND.n2177 585
R8220 GND.n4055 GND.n4054 585
R8221 GND.n4056 GND.n4055 585
R8222 GND.n2176 GND.n2175 585
R8223 GND.n4057 GND.n2176 585
R8224 GND.n4060 GND.n4059 585
R8225 GND.n4059 GND.n4058 585
R8226 GND.n2173 GND.n2172 585
R8227 GND.n2172 GND.n2171 585
R8228 GND.n4065 GND.n4064 585
R8229 GND.n4066 GND.n4065 585
R8230 GND.n2170 GND.n2169 585
R8231 GND.n4067 GND.n2170 585
R8232 GND.n4070 GND.n4069 585
R8233 GND.n4069 GND.n4068 585
R8234 GND.n2167 GND.n2166 585
R8235 GND.n2166 GND.n2165 585
R8236 GND.n4075 GND.n4074 585
R8237 GND.n4076 GND.n4075 585
R8238 GND.n2164 GND.n2163 585
R8239 GND.n4077 GND.n2164 585
R8240 GND.n4080 GND.n4079 585
R8241 GND.n4079 GND.n4078 585
R8242 GND.n2161 GND.n2160 585
R8243 GND.n2160 GND.n2159 585
R8244 GND.n4085 GND.n4084 585
R8245 GND.n4086 GND.n4085 585
R8246 GND.n2158 GND.n2157 585
R8247 GND.n4087 GND.n2158 585
R8248 GND.n4090 GND.n4089 585
R8249 GND.n4089 GND.n4088 585
R8250 GND.n2155 GND.n2153 585
R8251 GND.n2153 GND.n2152 585
R8252 GND.n3935 GND.n3934 585
R8253 GND.n3936 GND.n3935 585
R8254 GND.n2251 GND.n2250 585
R8255 GND.n2250 GND.n2249 585
R8256 GND.n3930 GND.n3929 585
R8257 GND.n3929 GND.n3928 585
R8258 GND.n2254 GND.n2253 585
R8259 GND.n3927 GND.n2254 585
R8260 GND.n3925 GND.n3924 585
R8261 GND.n3926 GND.n3925 585
R8262 GND.n3923 GND.n2256 585
R8263 GND.n2256 GND.n2255 585
R8264 GND.n3922 GND.n3921 585
R8265 GND.n3921 GND.n3920 585
R8266 GND.n2261 GND.n2260 585
R8267 GND.n3919 GND.n2261 585
R8268 GND.n3917 GND.n3916 585
R8269 GND.n3918 GND.n3917 585
R8270 GND.n3915 GND.n2263 585
R8271 GND.n2263 GND.n2262 585
R8272 GND.n3914 GND.n3913 585
R8273 GND.n3913 GND.n3912 585
R8274 GND.n2269 GND.n2268 585
R8275 GND.n3911 GND.n2269 585
R8276 GND.n3909 GND.n3908 585
R8277 GND.n3910 GND.n3909 585
R8278 GND.n3907 GND.n2271 585
R8279 GND.n2271 GND.n2270 585
R8280 GND.n3906 GND.n3905 585
R8281 GND.n3905 GND.n3904 585
R8282 GND.n2277 GND.n2276 585
R8283 GND.n3903 GND.n2277 585
R8284 GND.n3901 GND.n3900 585
R8285 GND.n3902 GND.n3901 585
R8286 GND.n3899 GND.n2279 585
R8287 GND.n2279 GND.n2278 585
R8288 GND.n3898 GND.n3897 585
R8289 GND.n3897 GND.n3896 585
R8290 GND.n2285 GND.n2284 585
R8291 GND.n3895 GND.n2285 585
R8292 GND.n3893 GND.n3892 585
R8293 GND.n3894 GND.n3893 585
R8294 GND.n3891 GND.n2287 585
R8295 GND.n2287 GND.n2286 585
R8296 GND.n3890 GND.n3889 585
R8297 GND.n3889 GND.n3888 585
R8298 GND.n2293 GND.n2292 585
R8299 GND.n3887 GND.n2293 585
R8300 GND.n3885 GND.n3884 585
R8301 GND.n3886 GND.n3885 585
R8302 GND.n3883 GND.n2295 585
R8303 GND.n2295 GND.n2294 585
R8304 GND.n3882 GND.n3881 585
R8305 GND.n3881 GND.n3880 585
R8306 GND.n2301 GND.n2300 585
R8307 GND.n3879 GND.n2301 585
R8308 GND.n3877 GND.n3876 585
R8309 GND.n3878 GND.n3877 585
R8310 GND.n3875 GND.n2303 585
R8311 GND.n2303 GND.n2302 585
R8312 GND.n3874 GND.n3873 585
R8313 GND.n3873 GND.n3872 585
R8314 GND.n2309 GND.n2308 585
R8315 GND.n3871 GND.n2309 585
R8316 GND.n3869 GND.n3868 585
R8317 GND.n3870 GND.n3869 585
R8318 GND.n3867 GND.n2311 585
R8319 GND.n2311 GND.n2310 585
R8320 GND.n3866 GND.n3865 585
R8321 GND.n3865 GND.n3864 585
R8322 GND.n2317 GND.n2316 585
R8323 GND.n3863 GND.n2317 585
R8324 GND.n3861 GND.n3860 585
R8325 GND.n3862 GND.n3861 585
R8326 GND.n3859 GND.n2319 585
R8327 GND.n2319 GND.n2318 585
R8328 GND.n3858 GND.n3857 585
R8329 GND.n3857 GND.n3856 585
R8330 GND.n2325 GND.n2324 585
R8331 GND.n3855 GND.n2325 585
R8332 GND.n3853 GND.n3852 585
R8333 GND.n3854 GND.n3853 585
R8334 GND.n3851 GND.n2327 585
R8335 GND.n2327 GND.n2326 585
R8336 GND.n3850 GND.n3849 585
R8337 GND.n3849 GND.n3848 585
R8338 GND.n2333 GND.n2332 585
R8339 GND.n3847 GND.n2333 585
R8340 GND.n3845 GND.n3844 585
R8341 GND.n3846 GND.n3845 585
R8342 GND.n3843 GND.n2335 585
R8343 GND.n2335 GND.n2334 585
R8344 GND.n3842 GND.n3841 585
R8345 GND.n3841 GND.n3840 585
R8346 GND.n2341 GND.n2340 585
R8347 GND.n3839 GND.n2341 585
R8348 GND.n3837 GND.n3836 585
R8349 GND.n3838 GND.n3837 585
R8350 GND.n3835 GND.n2343 585
R8351 GND.n2343 GND.n2342 585
R8352 GND.n3834 GND.n3833 585
R8353 GND.n3833 GND.n3832 585
R8354 GND.n2349 GND.n2348 585
R8355 GND.n3831 GND.n2349 585
R8356 GND.n3829 GND.n3828 585
R8357 GND.n3830 GND.n3829 585
R8358 GND.n3827 GND.n2351 585
R8359 GND.n2351 GND.n2350 585
R8360 GND.n3826 GND.n3825 585
R8361 GND.n3825 GND.n3824 585
R8362 GND.n2357 GND.n2356 585
R8363 GND.n3823 GND.n2357 585
R8364 GND.n3821 GND.n3820 585
R8365 GND.n3822 GND.n3821 585
R8366 GND.n3819 GND.n2359 585
R8367 GND.n2359 GND.n2358 585
R8368 GND.n3818 GND.n3817 585
R8369 GND.n3817 GND.n3816 585
R8370 GND.n2365 GND.n2364 585
R8371 GND.n3815 GND.n2365 585
R8372 GND.n3813 GND.n3812 585
R8373 GND.n3814 GND.n3813 585
R8374 GND.n3811 GND.n2367 585
R8375 GND.n2367 GND.n2366 585
R8376 GND.n3810 GND.n3809 585
R8377 GND.n3809 GND.n3808 585
R8378 GND.n2373 GND.n2372 585
R8379 GND.n3807 GND.n2373 585
R8380 GND.n3805 GND.n3804 585
R8381 GND.n3806 GND.n3805 585
R8382 GND.n3803 GND.n2375 585
R8383 GND.n2375 GND.n2374 585
R8384 GND.n3802 GND.n3801 585
R8385 GND.n3801 GND.n3800 585
R8386 GND.n2381 GND.n2380 585
R8387 GND.n3799 GND.n2381 585
R8388 GND.n3797 GND.n3796 585
R8389 GND.n3798 GND.n3797 585
R8390 GND.n3795 GND.n2383 585
R8391 GND.n2383 GND.n2382 585
R8392 GND.n3794 GND.n3793 585
R8393 GND.n3793 GND.n3792 585
R8394 GND.n2389 GND.n2388 585
R8395 GND.n3791 GND.n2389 585
R8396 GND.n3789 GND.n3788 585
R8397 GND.n3790 GND.n3789 585
R8398 GND.n3787 GND.n2391 585
R8399 GND.n2391 GND.n2390 585
R8400 GND.n3786 GND.n3785 585
R8401 GND.n3785 GND.n3784 585
R8402 GND.n2397 GND.n2396 585
R8403 GND.n3783 GND.n2397 585
R8404 GND.n3781 GND.n3780 585
R8405 GND.n3782 GND.n3781 585
R8406 GND.n3779 GND.n2399 585
R8407 GND.n2399 GND.n2398 585
R8408 GND.n3778 GND.n3777 585
R8409 GND.n3777 GND.n3776 585
R8410 GND.n2405 GND.n2404 585
R8411 GND.n3775 GND.n2405 585
R8412 GND.n3773 GND.n3772 585
R8413 GND.n3774 GND.n3773 585
R8414 GND.n3771 GND.n2407 585
R8415 GND.n2407 GND.n2406 585
R8416 GND.n3770 GND.n3769 585
R8417 GND.n3769 GND.n3768 585
R8418 GND.n2413 GND.n2412 585
R8419 GND.n3767 GND.n2413 585
R8420 GND.n3765 GND.n3764 585
R8421 GND.n3766 GND.n3765 585
R8422 GND.n3763 GND.n2415 585
R8423 GND.n2415 GND.n2414 585
R8424 GND.n3762 GND.n3761 585
R8425 GND.n3761 GND.n3760 585
R8426 GND.n2421 GND.n2420 585
R8427 GND.n3759 GND.n2421 585
R8428 GND.n3757 GND.n3756 585
R8429 GND.n3758 GND.n3757 585
R8430 GND.n3755 GND.n2423 585
R8431 GND.n2423 GND.n2422 585
R8432 GND.n3754 GND.n3753 585
R8433 GND.n3753 GND.n3752 585
R8434 GND.n2429 GND.n2428 585
R8435 GND.n3751 GND.n2429 585
R8436 GND.n3749 GND.n3748 585
R8437 GND.n3750 GND.n3749 585
R8438 GND.n3747 GND.n2431 585
R8439 GND.n2431 GND.n2430 585
R8440 GND.n3746 GND.n3745 585
R8441 GND.n3745 GND.n3744 585
R8442 GND.n2437 GND.n2436 585
R8443 GND.n3743 GND.n2437 585
R8444 GND.n3741 GND.n3740 585
R8445 GND.n3742 GND.n3741 585
R8446 GND.n3739 GND.n2439 585
R8447 GND.n2439 GND.n2438 585
R8448 GND.n3738 GND.n3737 585
R8449 GND.n3737 GND.n3736 585
R8450 GND.n2445 GND.n2444 585
R8451 GND.n3735 GND.n2445 585
R8452 GND.n3733 GND.n3732 585
R8453 GND.n3734 GND.n3733 585
R8454 GND.n3731 GND.n2447 585
R8455 GND.n2447 GND.n2446 585
R8456 GND.n3730 GND.n3729 585
R8457 GND.n3729 GND.n3728 585
R8458 GND.n2453 GND.n2452 585
R8459 GND.n3727 GND.n2453 585
R8460 GND.n3725 GND.n3724 585
R8461 GND.n3726 GND.n3725 585
R8462 GND.n3723 GND.n2455 585
R8463 GND.n2455 GND.n2454 585
R8464 GND.n3722 GND.n3721 585
R8465 GND.n3721 GND.n3720 585
R8466 GND.n2461 GND.n2460 585
R8467 GND.n3719 GND.n2461 585
R8468 GND.n3717 GND.n3716 585
R8469 GND.n3718 GND.n3717 585
R8470 GND.n3715 GND.n2463 585
R8471 GND.n2463 GND.n2462 585
R8472 GND.n3714 GND.n3713 585
R8473 GND.n3713 GND.n3712 585
R8474 GND.n2469 GND.n2468 585
R8475 GND.n3711 GND.n2469 585
R8476 GND.n3709 GND.n3708 585
R8477 GND.n3710 GND.n3709 585
R8478 GND.n3707 GND.n2471 585
R8479 GND.n2471 GND.n2470 585
R8480 GND.n3706 GND.n3705 585
R8481 GND.n3705 GND.n3704 585
R8482 GND.n2477 GND.n2476 585
R8483 GND.n3703 GND.n2477 585
R8484 GND.n3701 GND.n3700 585
R8485 GND.n3702 GND.n3701 585
R8486 GND.n3699 GND.n2479 585
R8487 GND.n2479 GND.n2478 585
R8488 GND.n3698 GND.n3697 585
R8489 GND.n3697 GND.n3696 585
R8490 GND.n2485 GND.n2484 585
R8491 GND.n3695 GND.n2485 585
R8492 GND.n3693 GND.n3692 585
R8493 GND.n3694 GND.n3693 585
R8494 GND.n3691 GND.n2487 585
R8495 GND.n2487 GND.n2486 585
R8496 GND.n3690 GND.n3689 585
R8497 GND.n3689 GND.n3688 585
R8498 GND.n2493 GND.n2492 585
R8499 GND.n3687 GND.n2493 585
R8500 GND.n3685 GND.n3684 585
R8501 GND.n3686 GND.n3685 585
R8502 GND.n3683 GND.n2495 585
R8503 GND.n2495 GND.n2494 585
R8504 GND.n3682 GND.n3681 585
R8505 GND.n3681 GND.n3680 585
R8506 GND.n2501 GND.n2500 585
R8507 GND.n3679 GND.n2501 585
R8508 GND.n3677 GND.n3676 585
R8509 GND.n3678 GND.n3677 585
R8510 GND.n3675 GND.n2503 585
R8511 GND.n2503 GND.n2502 585
R8512 GND.n3674 GND.n3673 585
R8513 GND.n3673 GND.n3672 585
R8514 GND.n2509 GND.n2508 585
R8515 GND.n3671 GND.n2509 585
R8516 GND.n3669 GND.n3668 585
R8517 GND.n3670 GND.n3669 585
R8518 GND.n3667 GND.n2511 585
R8519 GND.n2511 GND.n2510 585
R8520 GND.n3666 GND.n3665 585
R8521 GND.n3665 GND.n3664 585
R8522 GND.n2517 GND.n2516 585
R8523 GND.n3663 GND.n2517 585
R8524 GND.n3661 GND.n3660 585
R8525 GND.n3662 GND.n3661 585
R8526 GND.n3659 GND.n2519 585
R8527 GND.n2519 GND.n2518 585
R8528 GND.n3658 GND.n3657 585
R8529 GND.n3657 GND.n3656 585
R8530 GND.n2525 GND.n2524 585
R8531 GND.n3655 GND.n2525 585
R8532 GND.n3653 GND.n3652 585
R8533 GND.n3654 GND.n3653 585
R8534 GND.n3651 GND.n2527 585
R8535 GND.n2527 GND.n2526 585
R8536 GND.n3650 GND.n3649 585
R8537 GND.n3649 GND.n3648 585
R8538 GND.n2533 GND.n2532 585
R8539 GND.n3647 GND.n2533 585
R8540 GND.n3645 GND.n3644 585
R8541 GND.n3646 GND.n3645 585
R8542 GND.n3643 GND.n2535 585
R8543 GND.n2535 GND.n2534 585
R8544 GND.n3642 GND.n3641 585
R8545 GND.n3641 GND.n3640 585
R8546 GND.n2541 GND.n2540 585
R8547 GND.n3639 GND.n2541 585
R8548 GND.n3637 GND.n3636 585
R8549 GND.n3638 GND.n3637 585
R8550 GND.n3635 GND.n2543 585
R8551 GND.n2543 GND.n2542 585
R8552 GND.n3634 GND.n3633 585
R8553 GND.n3633 GND.n3632 585
R8554 GND.n2549 GND.n2548 585
R8555 GND.n3631 GND.n2549 585
R8556 GND.n3629 GND.n3628 585
R8557 GND.n3630 GND.n3629 585
R8558 GND.n3627 GND.n2551 585
R8559 GND.n2551 GND.n2550 585
R8560 GND.n3626 GND.n3625 585
R8561 GND.n3625 GND.n3624 585
R8562 GND.n2557 GND.n2556 585
R8563 GND.n3623 GND.n2557 585
R8564 GND.n3621 GND.n3620 585
R8565 GND.n3622 GND.n3621 585
R8566 GND.n3619 GND.n2559 585
R8567 GND.n2559 GND.n2558 585
R8568 GND.n3618 GND.n3617 585
R8569 GND.n3617 GND.n3616 585
R8570 GND.n2565 GND.n2564 585
R8571 GND.n3615 GND.n2565 585
R8572 GND.n3613 GND.n3612 585
R8573 GND.n3614 GND.n3613 585
R8574 GND.n3611 GND.n2567 585
R8575 GND.n2567 GND.n2566 585
R8576 GND.n3610 GND.n3609 585
R8577 GND.n3609 GND.n3608 585
R8578 GND.n2573 GND.n2572 585
R8579 GND.n3607 GND.n2573 585
R8580 GND.n3605 GND.n3604 585
R8581 GND.n3606 GND.n3605 585
R8582 GND.n3603 GND.n2575 585
R8583 GND.n2575 GND.n2574 585
R8584 GND.n3602 GND.n3601 585
R8585 GND.n3601 GND.n3600 585
R8586 GND.n2581 GND.n2580 585
R8587 GND.n3599 GND.n2581 585
R8588 GND.n3597 GND.n3596 585
R8589 GND.n3598 GND.n3597 585
R8590 GND.n3595 GND.n2583 585
R8591 GND.n2583 GND.n2582 585
R8592 GND.n3594 GND.n3593 585
R8593 GND.n3593 GND.n3592 585
R8594 GND.n2589 GND.n2588 585
R8595 GND.n3591 GND.n2589 585
R8596 GND.n3589 GND.n3588 585
R8597 GND.n3590 GND.n3589 585
R8598 GND.n3587 GND.n2591 585
R8599 GND.n2591 GND.n2590 585
R8600 GND.n3586 GND.n3585 585
R8601 GND.n3585 GND.n3584 585
R8602 GND.n2597 GND.n2596 585
R8603 GND.n3583 GND.n2597 585
R8604 GND.n3581 GND.n3580 585
R8605 GND.n3582 GND.n3581 585
R8606 GND.n3579 GND.n2599 585
R8607 GND.n2599 GND.n2598 585
R8608 GND.n3578 GND.n3577 585
R8609 GND.n3577 GND.n3576 585
R8610 GND.n2605 GND.n2604 585
R8611 GND.n3575 GND.n2605 585
R8612 GND.n3573 GND.n3572 585
R8613 GND.n3574 GND.n3573 585
R8614 GND.n3571 GND.n2607 585
R8615 GND.n2607 GND.n2606 585
R8616 GND.n3570 GND.n3569 585
R8617 GND.n3569 GND.n3568 585
R8618 GND.n2613 GND.n2612 585
R8619 GND.n3567 GND.n2613 585
R8620 GND.n3565 GND.n3564 585
R8621 GND.n3566 GND.n3565 585
R8622 GND.n3563 GND.n2615 585
R8623 GND.n2615 GND.n2614 585
R8624 GND.n3562 GND.n3561 585
R8625 GND.n3561 GND.n3560 585
R8626 GND.n2621 GND.n2620 585
R8627 GND.n3559 GND.n2621 585
R8628 GND.n3557 GND.n3556 585
R8629 GND.n3558 GND.n3557 585
R8630 GND.n3555 GND.n2623 585
R8631 GND.n2623 GND.n2622 585
R8632 GND.n3554 GND.n3553 585
R8633 GND.n3553 GND.n3552 585
R8634 GND.n2629 GND.n2628 585
R8635 GND.n3551 GND.n2629 585
R8636 GND.n3549 GND.n3548 585
R8637 GND.n3550 GND.n3549 585
R8638 GND.n3547 GND.n2631 585
R8639 GND.n2631 GND.n2630 585
R8640 GND.n3546 GND.n3545 585
R8641 GND.n3545 GND.n3544 585
R8642 GND.n2637 GND.n2636 585
R8643 GND.n3543 GND.n2637 585
R8644 GND.n3541 GND.n3540 585
R8645 GND.n3542 GND.n3541 585
R8646 GND.n3539 GND.n2639 585
R8647 GND.n2639 GND.n2638 585
R8648 GND.n3538 GND.n3537 585
R8649 GND.n3537 GND.n3536 585
R8650 GND.n2645 GND.n2644 585
R8651 GND.n3535 GND.n2645 585
R8652 GND.n3533 GND.n3532 585
R8653 GND.n3534 GND.n3533 585
R8654 GND.n3531 GND.n2647 585
R8655 GND.n2647 GND.n2646 585
R8656 GND.n3530 GND.n3529 585
R8657 GND.n3529 GND.n3528 585
R8658 GND.n2653 GND.n2652 585
R8659 GND.n3527 GND.n2653 585
R8660 GND.n3525 GND.n3524 585
R8661 GND.n3526 GND.n3525 585
R8662 GND.n3523 GND.n2655 585
R8663 GND.n2655 GND.n2654 585
R8664 GND.n3522 GND.n3521 585
R8665 GND.n3521 GND.n3520 585
R8666 GND.n2661 GND.n2660 585
R8667 GND.n3519 GND.n2661 585
R8668 GND.n3517 GND.n3516 585
R8669 GND.n3518 GND.n3517 585
R8670 GND.n3515 GND.n2663 585
R8671 GND.n2663 GND.n2662 585
R8672 GND.n3514 GND.n3513 585
R8673 GND.n3513 GND.n3512 585
R8674 GND.n2669 GND.n2668 585
R8675 GND.n3511 GND.n2669 585
R8676 GND.n3509 GND.n3508 585
R8677 GND.n3510 GND.n3509 585
R8678 GND.n3507 GND.n2671 585
R8679 GND.n2671 GND.n2670 585
R8680 GND.n3506 GND.n3505 585
R8681 GND.n3505 GND.n3504 585
R8682 GND.n2677 GND.n2676 585
R8683 GND.n3503 GND.n2677 585
R8684 GND.n3501 GND.n3500 585
R8685 GND.n3502 GND.n3501 585
R8686 GND.n3499 GND.n2679 585
R8687 GND.n2679 GND.n2678 585
R8688 GND.n3498 GND.n3497 585
R8689 GND.n3497 GND.n3496 585
R8690 GND.n2685 GND.n2684 585
R8691 GND.n3495 GND.n2685 585
R8692 GND.n3493 GND.n3492 585
R8693 GND.n3494 GND.n3493 585
R8694 GND.n3491 GND.n2687 585
R8695 GND.n2687 GND.n2686 585
R8696 GND.n3490 GND.n3489 585
R8697 GND.n3489 GND.n3488 585
R8698 GND.n2693 GND.n2692 585
R8699 GND.n3487 GND.n2693 585
R8700 GND.n3485 GND.n3484 585
R8701 GND.n3486 GND.n3485 585
R8702 GND.n3483 GND.n2695 585
R8703 GND.n2695 GND.n2694 585
R8704 GND.n3482 GND.n3481 585
R8705 GND.n3481 GND.n3480 585
R8706 GND.n2701 GND.n2700 585
R8707 GND.n3479 GND.n2701 585
R8708 GND.n3477 GND.n3476 585
R8709 GND.n3478 GND.n3477 585
R8710 GND.n3475 GND.n2703 585
R8711 GND.n2703 GND.n2702 585
R8712 GND.n3474 GND.n3473 585
R8713 GND.n3473 GND.n3472 585
R8714 GND.n2709 GND.n2708 585
R8715 GND.n3471 GND.n2709 585
R8716 GND.n3469 GND.n3468 585
R8717 GND.n3470 GND.n3469 585
R8718 GND.n3467 GND.n2711 585
R8719 GND.n2711 GND.n2710 585
R8720 GND.n3466 GND.n3465 585
R8721 GND.n3465 GND.n3464 585
R8722 GND.n2717 GND.n2716 585
R8723 GND.n3463 GND.n2717 585
R8724 GND.n3461 GND.n3460 585
R8725 GND.n3462 GND.n3461 585
R8726 GND.n3459 GND.n2719 585
R8727 GND.n2719 GND.n2718 585
R8728 GND.n3458 GND.n3457 585
R8729 GND.n3457 GND.n3456 585
R8730 GND.n2725 GND.n2724 585
R8731 GND.n3455 GND.n2725 585
R8732 GND.n3453 GND.n3452 585
R8733 GND.n3454 GND.n3453 585
R8734 GND.n3451 GND.n2727 585
R8735 GND.n2727 GND.n2726 585
R8736 GND.n3450 GND.n3449 585
R8737 GND.n3449 GND.n3448 585
R8738 GND.n2733 GND.n2732 585
R8739 GND.n3447 GND.n2733 585
R8740 GND.n3445 GND.n3444 585
R8741 GND.n3446 GND.n3445 585
R8742 GND.n3443 GND.n2735 585
R8743 GND.n2735 GND.n2734 585
R8744 GND.n3442 GND.n3441 585
R8745 GND.n3441 GND.n3440 585
R8746 GND.n2741 GND.n2740 585
R8747 GND.n3439 GND.n2741 585
R8748 GND.n3437 GND.n3436 585
R8749 GND.n3438 GND.n3437 585
R8750 GND.n3435 GND.n2743 585
R8751 GND.n2743 GND.n2742 585
R8752 GND.n3434 GND.n3433 585
R8753 GND.n3433 GND.n3432 585
R8754 GND.n2749 GND.n2748 585
R8755 GND.n3431 GND.n2749 585
R8756 GND.n3429 GND.n3428 585
R8757 GND.n3430 GND.n3429 585
R8758 GND.n3427 GND.n2751 585
R8759 GND.n2751 GND.n2750 585
R8760 GND.n3426 GND.n3425 585
R8761 GND.n3425 GND.n3424 585
R8762 GND.n2757 GND.n2756 585
R8763 GND.n3423 GND.n2757 585
R8764 GND.n3421 GND.n3420 585
R8765 GND.n3422 GND.n3421 585
R8766 GND.n3419 GND.n2759 585
R8767 GND.n2759 GND.n2758 585
R8768 GND.n3418 GND.n3417 585
R8769 GND.n3417 GND.n3416 585
R8770 GND.n2765 GND.n2764 585
R8771 GND.n3415 GND.n2765 585
R8772 GND.n3413 GND.n3412 585
R8773 GND.n3414 GND.n3413 585
R8774 GND.n3411 GND.n2767 585
R8775 GND.n2767 GND.n2766 585
R8776 GND.n3410 GND.n3409 585
R8777 GND.n3409 GND.n3408 585
R8778 GND.n2773 GND.n2772 585
R8779 GND.n3407 GND.n2773 585
R8780 GND.n3405 GND.n3404 585
R8781 GND.n3406 GND.n3405 585
R8782 GND.n3403 GND.n2775 585
R8783 GND.n2775 GND.n2774 585
R8784 GND.n3402 GND.n3401 585
R8785 GND.n3401 GND.n3400 585
R8786 GND.n2781 GND.n2780 585
R8787 GND.n3399 GND.n2781 585
R8788 GND.n3397 GND.n3396 585
R8789 GND.n3398 GND.n3397 585
R8790 GND.n3395 GND.n2783 585
R8791 GND.n2783 GND.n2782 585
R8792 GND.n3394 GND.n3393 585
R8793 GND.n3393 GND.n3392 585
R8794 GND.n2789 GND.n2788 585
R8795 GND.n3391 GND.n2789 585
R8796 GND.n3389 GND.n3388 585
R8797 GND.n3390 GND.n3389 585
R8798 GND.n3387 GND.n2791 585
R8799 GND.n2791 GND.n2790 585
R8800 GND.n3386 GND.n3385 585
R8801 GND.n3385 GND.n3384 585
R8802 GND.n2797 GND.n2796 585
R8803 GND.n3383 GND.n2797 585
R8804 GND.n3381 GND.n3380 585
R8805 GND.n3382 GND.n3381 585
R8806 GND.n3379 GND.n2799 585
R8807 GND.n2799 GND.n2798 585
R8808 GND.n3378 GND.n3377 585
R8809 GND.n3377 GND.n3376 585
R8810 GND.n2805 GND.n2804 585
R8811 GND.n3375 GND.n2805 585
R8812 GND.n3373 GND.n3372 585
R8813 GND.n3374 GND.n3373 585
R8814 GND.n3371 GND.n2807 585
R8815 GND.n2807 GND.n2806 585
R8816 GND.n3370 GND.n3369 585
R8817 GND.n3369 GND.n3368 585
R8818 GND.n2813 GND.n2812 585
R8819 GND.n3367 GND.n2813 585
R8820 GND.n3365 GND.n3364 585
R8821 GND.n3366 GND.n3365 585
R8822 GND.n3363 GND.n2815 585
R8823 GND.n2815 GND.n2814 585
R8824 GND.n3362 GND.n3361 585
R8825 GND.n3361 GND.n3360 585
R8826 GND.n2821 GND.n2820 585
R8827 GND.n3359 GND.n2821 585
R8828 GND.n3357 GND.n3356 585
R8829 GND.n3358 GND.n3357 585
R8830 GND.n3355 GND.n2823 585
R8831 GND.n2823 GND.n2822 585
R8832 GND.n3354 GND.n3353 585
R8833 GND.n3353 GND.n3352 585
R8834 GND.n2829 GND.n2828 585
R8835 GND.n3351 GND.n2829 585
R8836 GND.n3349 GND.n3348 585
R8837 GND.n3350 GND.n3349 585
R8838 GND.n3347 GND.n2831 585
R8839 GND.n2831 GND.n2830 585
R8840 GND.n3346 GND.n3345 585
R8841 GND.n3345 GND.n3344 585
R8842 GND.n2837 GND.n2836 585
R8843 GND.n3343 GND.n2837 585
R8844 GND.n3341 GND.n3340 585
R8845 GND.n3342 GND.n3341 585
R8846 GND.n3339 GND.n2839 585
R8847 GND.n2839 GND.n2838 585
R8848 GND.n3338 GND.n3337 585
R8849 GND.n3337 GND.n3336 585
R8850 GND.n2845 GND.n2844 585
R8851 GND.n3335 GND.n2845 585
R8852 GND.n3333 GND.n3332 585
R8853 GND.n3334 GND.n3333 585
R8854 GND.n3331 GND.n2847 585
R8855 GND.n2847 GND.n2846 585
R8856 GND.n3330 GND.n3329 585
R8857 GND.n3329 GND.n3328 585
R8858 GND.n2853 GND.n2852 585
R8859 GND.n3327 GND.n2853 585
R8860 GND.n3325 GND.n3324 585
R8861 GND.n3326 GND.n3325 585
R8862 GND.n3323 GND.n2855 585
R8863 GND.n2855 GND.n2854 585
R8864 GND.n3322 GND.n3321 585
R8865 GND.n3321 GND.n3320 585
R8866 GND.n2861 GND.n2860 585
R8867 GND.n3319 GND.n2861 585
R8868 GND.n3317 GND.n3316 585
R8869 GND.n3318 GND.n3317 585
R8870 GND.n3315 GND.n2863 585
R8871 GND.n2863 GND.n2862 585
R8872 GND.n3314 GND.n3313 585
R8873 GND.n3313 GND.n3312 585
R8874 GND.n2869 GND.n2868 585
R8875 GND.n3311 GND.n2869 585
R8876 GND.n3309 GND.n3308 585
R8877 GND.n3310 GND.n3309 585
R8878 GND.n3307 GND.n2871 585
R8879 GND.n2871 GND.n2870 585
R8880 GND.n3306 GND.n3305 585
R8881 GND.n3305 GND.n3304 585
R8882 GND.n2877 GND.n2876 585
R8883 GND.n3303 GND.n2877 585
R8884 GND.n3301 GND.n3300 585
R8885 GND.n3302 GND.n3301 585
R8886 GND.n3299 GND.n2879 585
R8887 GND.n2879 GND.n2878 585
R8888 GND.n3298 GND.n3297 585
R8889 GND.n3297 GND.n3296 585
R8890 GND.n2885 GND.n2884 585
R8891 GND.n3295 GND.n2885 585
R8892 GND.n3293 GND.n3292 585
R8893 GND.n3294 GND.n3293 585
R8894 GND.n3291 GND.n2887 585
R8895 GND.n2887 GND.n2886 585
R8896 GND.n3290 GND.n3289 585
R8897 GND.n3289 GND.n3288 585
R8898 GND.n2893 GND.n2892 585
R8899 GND.n3287 GND.n2893 585
R8900 GND.n3285 GND.n3284 585
R8901 GND.n3286 GND.n3285 585
R8902 GND.n3283 GND.n2895 585
R8903 GND.n2895 GND.n2894 585
R8904 GND.n3282 GND.n3281 585
R8905 GND.n3281 GND.n3280 585
R8906 GND.n2901 GND.n2900 585
R8907 GND.n3279 GND.n2901 585
R8908 GND.n3277 GND.n3276 585
R8909 GND.n3278 GND.n3277 585
R8910 GND.n3275 GND.n2903 585
R8911 GND.n2903 GND.n2902 585
R8912 GND.n3274 GND.n3273 585
R8913 GND.n3273 GND.n3272 585
R8914 GND.n2909 GND.n2908 585
R8915 GND.n3271 GND.n2909 585
R8916 GND.n3269 GND.n3268 585
R8917 GND.n3270 GND.n3269 585
R8918 GND.n3267 GND.n2911 585
R8919 GND.n2911 GND.n2910 585
R8920 GND.n3266 GND.n3265 585
R8921 GND.n3265 GND.n3264 585
R8922 GND.n2917 GND.n2916 585
R8923 GND.n3263 GND.n2917 585
R8924 GND.n3261 GND.n3260 585
R8925 GND.n3262 GND.n3261 585
R8926 GND.n3259 GND.n2919 585
R8927 GND.n2919 GND.n2918 585
R8928 GND.n3258 GND.n3257 585
R8929 GND.n3257 GND.n3256 585
R8930 GND.n2925 GND.n2924 585
R8931 GND.n3255 GND.n2925 585
R8932 GND.n3253 GND.n3252 585
R8933 GND.n3254 GND.n3253 585
R8934 GND.n3251 GND.n2927 585
R8935 GND.n2927 GND.n2926 585
R8936 GND.n3250 GND.n3249 585
R8937 GND.n3249 GND.n3248 585
R8938 GND.n2933 GND.n2932 585
R8939 GND.n3247 GND.n2933 585
R8940 GND.n3245 GND.n3244 585
R8941 GND.n3246 GND.n3245 585
R8942 GND.n3243 GND.n2935 585
R8943 GND.n2935 GND.n2934 585
R8944 GND.n3242 GND.n3241 585
R8945 GND.n3241 GND.n3240 585
R8946 GND.n2941 GND.n2940 585
R8947 GND.n3239 GND.n2941 585
R8948 GND.n3237 GND.n3236 585
R8949 GND.n3238 GND.n3237 585
R8950 GND.n3235 GND.n2943 585
R8951 GND.n2943 GND.n2942 585
R8952 GND.n3234 GND.n3233 585
R8953 GND.n3233 GND.n3232 585
R8954 GND.n2949 GND.n2948 585
R8955 GND.n3231 GND.n2949 585
R8956 GND.n3229 GND.n3228 585
R8957 GND.n3230 GND.n3229 585
R8958 GND.n3227 GND.n2951 585
R8959 GND.n2951 GND.n2950 585
R8960 GND.n3226 GND.n3225 585
R8961 GND.n3225 GND.n3224 585
R8962 GND.n2957 GND.n2956 585
R8963 GND.n3223 GND.n2957 585
R8964 GND.n3221 GND.n3220 585
R8965 GND.n3222 GND.n3221 585
R8966 GND.n3219 GND.n2959 585
R8967 GND.n2959 GND.n2958 585
R8968 GND.n3218 GND.n3217 585
R8969 GND.n3217 GND.n3216 585
R8970 GND.n2965 GND.n2964 585
R8971 GND.n3215 GND.n2965 585
R8972 GND.n384 GND.n382 585
R8973 GND.n382 GND.n381 585
R8974 GND.n3090 GND.n3089 585
R8975 GND.n3091 GND.n3090 585
R8976 GND.n3086 GND.n3085 585
R8977 GND.n3092 GND.n3086 585
R8978 GND.n3095 GND.n3094 585
R8979 GND.n3094 GND.n3093 585
R8980 GND.n3096 GND.n3080 585
R8981 GND.n3080 GND.n3079 585
R8982 GND.n3098 GND.n3097 585
R8983 GND.n3099 GND.n3098 585
R8984 GND.n3078 GND.n3077 585
R8985 GND.n3100 GND.n3078 585
R8986 GND.n3103 GND.n3102 585
R8987 GND.n3102 GND.n3101 585
R8988 GND.n3104 GND.n3072 585
R8989 GND.n3072 GND.n3071 585
R8990 GND.n3106 GND.n3105 585
R8991 GND.n3107 GND.n3106 585
R8992 GND.n3070 GND.n3069 585
R8993 GND.n3108 GND.n3070 585
R8994 GND.n3111 GND.n3110 585
R8995 GND.n3110 GND.n3109 585
R8996 GND.n3112 GND.n3064 585
R8997 GND.n3064 GND.n3063 585
R8998 GND.n3114 GND.n3113 585
R8999 GND.n3115 GND.n3114 585
R9000 GND.n3062 GND.n3061 585
R9001 GND.n3116 GND.n3062 585
R9002 GND.n3119 GND.n3118 585
R9003 GND.n3118 GND.n3117 585
R9004 GND.n3120 GND.n3056 585
R9005 GND.n3056 GND.n3055 585
R9006 GND.n3122 GND.n3121 585
R9007 GND.n3123 GND.n3122 585
R9008 GND.n3054 GND.n3053 585
R9009 GND.n3124 GND.n3054 585
R9010 GND.n3127 GND.n3126 585
R9011 GND.n3126 GND.n3125 585
R9012 GND.n3128 GND.n3048 585
R9013 GND.n3048 GND.n3047 585
R9014 GND.n3130 GND.n3129 585
R9015 GND.n3131 GND.n3130 585
R9016 GND.n3046 GND.n3045 585
R9017 GND.n3132 GND.n3046 585
R9018 GND.n3135 GND.n3134 585
R9019 GND.n3134 GND.n3133 585
R9020 GND.n3136 GND.n3040 585
R9021 GND.n3040 GND.n3039 585
R9022 GND.n3138 GND.n3137 585
R9023 GND.n3139 GND.n3138 585
R9024 GND.n3038 GND.n3037 585
R9025 GND.n3140 GND.n3038 585
R9026 GND.n3143 GND.n3142 585
R9027 GND.n3142 GND.n3141 585
R9028 GND.n3144 GND.n3032 585
R9029 GND.n3032 GND.n3031 585
R9030 GND.n3146 GND.n3145 585
R9031 GND.n3147 GND.n3146 585
R9032 GND.n3030 GND.n3029 585
R9033 GND.n3148 GND.n3030 585
R9034 GND.n3151 GND.n3150 585
R9035 GND.n3150 GND.n3149 585
R9036 GND.n3152 GND.n3024 585
R9037 GND.n3024 GND.n3023 585
R9038 GND.n3154 GND.n3153 585
R9039 GND.n3155 GND.n3154 585
R9040 GND.n3022 GND.n3021 585
R9041 GND.n3156 GND.n3022 585
R9042 GND.n3159 GND.n3158 585
R9043 GND.n3158 GND.n3157 585
R9044 GND.n3160 GND.n3016 585
R9045 GND.n3016 GND.n3015 585
R9046 GND.n3162 GND.n3161 585
R9047 GND.n3163 GND.n3162 585
R9048 GND.n3014 GND.n3013 585
R9049 GND.n3164 GND.n3014 585
R9050 GND.n3167 GND.n3166 585
R9051 GND.n3166 GND.n3165 585
R9052 GND.n3168 GND.n3008 585
R9053 GND.n3008 GND.n3007 585
R9054 GND.n3170 GND.n3169 585
R9055 GND.n3171 GND.n3170 585
R9056 GND.n3006 GND.n3005 585
R9057 GND.n3172 GND.n3006 585
R9058 GND.n3175 GND.n3174 585
R9059 GND.n3174 GND.n3173 585
R9060 GND.n3176 GND.n3000 585
R9061 GND.n3000 GND.n2999 585
R9062 GND.n3178 GND.n3177 585
R9063 GND.n3179 GND.n3178 585
R9064 GND.n2998 GND.n2997 585
R9065 GND.n3180 GND.n2998 585
R9066 GND.n3183 GND.n3182 585
R9067 GND.n3182 GND.n3181 585
R9068 GND.n3184 GND.n2992 585
R9069 GND.n2992 GND.n2991 585
R9070 GND.n3186 GND.n3185 585
R9071 GND.n3187 GND.n3186 585
R9072 GND.n2990 GND.n2989 585
R9073 GND.n3188 GND.n2990 585
R9074 GND.n3191 GND.n3190 585
R9075 GND.n3190 GND.n3189 585
R9076 GND.n3192 GND.n2984 585
R9077 GND.n2984 GND.n2983 585
R9078 GND.n3194 GND.n3193 585
R9079 GND.n3195 GND.n3194 585
R9080 GND.n2982 GND.n2981 585
R9081 GND.n3196 GND.n2982 585
R9082 GND.n3199 GND.n3198 585
R9083 GND.n3198 GND.n3197 585
R9084 GND.n3200 GND.n2977 585
R9085 GND.n2977 GND.n2976 585
R9086 GND.n3202 GND.n3201 585
R9087 GND.n3203 GND.n3202 585
R9088 GND.n2974 GND.n2972 585
R9089 GND.n3204 GND.n2974 585
R9090 GND.n3207 GND.n3206 585
R9091 GND.n3206 GND.n3205 585
R9092 GND.n2973 GND.n2970 585
R9093 GND.n2975 GND.n2973 585
R9094 GND.n3211 GND.n2967 585
R9095 GND.n2967 GND.n2966 585
R9096 GND.n3213 GND.n3212 585
R9097 GND.n3214 GND.n3213 585
R9098 GND.n8462 GND.n8461 585
R9099 GND.n8463 GND.n8462 585
R9100 GND.n332 GND.n331 585
R9101 GND.n8456 GND.n332 585
R9102 GND.n8471 GND.n8470 585
R9103 GND.n8470 GND.n8469 585
R9104 GND.n8472 GND.n327 585
R9105 GND.n8240 GND.n327 585
R9106 GND.n8474 GND.n8473 585
R9107 GND.n8475 GND.n8474 585
R9108 GND.n312 GND.n311 585
R9109 GND.n8246 GND.n312 585
R9110 GND.n8483 GND.n8482 585
R9111 GND.n8482 GND.n8481 585
R9112 GND.n8484 GND.n307 585
R9113 GND.n8231 GND.n307 585
R9114 GND.n8486 GND.n8485 585
R9115 GND.n8487 GND.n8486 585
R9116 GND.n291 GND.n290 585
R9117 GND.n8222 GND.n291 585
R9118 GND.n8495 GND.n8494 585
R9119 GND.n8494 GND.n8493 585
R9120 GND.n8496 GND.n286 585
R9121 GND.n8215 GND.n286 585
R9122 GND.n8498 GND.n8497 585
R9123 GND.n8499 GND.n8498 585
R9124 GND.n270 GND.n269 585
R9125 GND.n8207 GND.n270 585
R9126 GND.n8507 GND.n8506 585
R9127 GND.n8506 GND.n8505 585
R9128 GND.n8508 GND.n265 585
R9129 GND.n8200 GND.n265 585
R9130 GND.n8510 GND.n8509 585
R9131 GND.n8511 GND.n8510 585
R9132 GND.n250 GND.n249 585
R9133 GND.n8192 GND.n250 585
R9134 GND.n8519 GND.n8518 585
R9135 GND.n8518 GND.n8517 585
R9136 GND.n8520 GND.n245 585
R9137 GND.n8185 GND.n245 585
R9138 GND.n8522 GND.n8521 585
R9139 GND.n8523 GND.n8522 585
R9140 GND.n229 GND.n228 585
R9141 GND.n8177 GND.n229 585
R9142 GND.n8531 GND.n8530 585
R9143 GND.n8530 GND.n8529 585
R9144 GND.n8532 GND.n224 585
R9145 GND.n8170 GND.n224 585
R9146 GND.n8534 GND.n8533 585
R9147 GND.n8535 GND.n8534 585
R9148 GND.n208 GND.n207 585
R9149 GND.n8162 GND.n208 585
R9150 GND.n8543 GND.n8542 585
R9151 GND.n8542 GND.n8541 585
R9152 GND.n8544 GND.n203 585
R9153 GND.n8155 GND.n203 585
R9154 GND.n8546 GND.n8545 585
R9155 GND.n8547 GND.n8546 585
R9156 GND.n188 GND.n187 585
R9157 GND.n8147 GND.n188 585
R9158 GND.n8555 GND.n8554 585
R9159 GND.n8554 GND.n8553 585
R9160 GND.n8556 GND.n182 585
R9161 GND.n8140 GND.n182 585
R9162 GND.n8558 GND.n8557 585
R9163 GND.n8559 GND.n8558 585
R9164 GND.n183 GND.n181 585
R9165 GND.n8132 GND.n181 585
R9166 GND.n8127 GND.n8126 585
R9167 GND.n8126 GND.n8125 585
R9168 GND.n434 GND.n433 585
R9169 GND.n435 GND.n434 585
R9170 GND.n8029 GND.n161 585
R9171 GND.n8566 GND.n161 585
R9172 GND.n8031 GND.n8030 585
R9173 GND.n8032 GND.n8031 585
R9174 GND.n444 GND.n443 585
R9175 GND.n443 GND.n441 585
R9176 GND.n8012 GND.n452 585
R9177 GND.n8020 GND.n452 585
R9178 GND.n8014 GND.n8013 585
R9179 GND.n8015 GND.n8014 585
R9180 GND.n458 GND.n457 585
R9181 GND.n8006 GND.n457 585
R9182 GND.n7976 GND.n7975 585
R9183 GND.n7975 GND.n7974 585
R9184 GND.n7977 GND.n471 585
R9185 GND.n7991 GND.n471 585
R9186 GND.n7978 GND.n483 585
R9187 GND.n7968 GND.n483 585
R9188 GND.n7980 GND.n7979 585
R9189 GND.n7981 GND.n7980 585
R9190 GND.n484 GND.n482 585
R9191 GND.n7964 GND.n482 585
R9192 GND.n7939 GND.n7938 585
R9193 GND.n7938 GND.n7937 585
R9194 GND.n7940 GND.n498 585
R9195 GND.n7954 GND.n498 585
R9196 GND.n7941 GND.n510 585
R9197 GND.n549 GND.n510 585
R9198 GND.n7943 GND.n7942 585
R9199 GND.n7944 GND.n7943 585
R9200 GND.n511 GND.n509 585
R9201 GND.n7882 GND.n509 585
R9202 GND.n7887 GND.n530 585
R9203 GND.n7899 GND.n530 585
R9204 GND.n7888 GND.n541 585
R9205 GND.n541 GND.n526 585
R9206 GND.n7890 GND.n7889 585
R9207 GND.n7891 GND.n7890 585
R9208 GND.n542 GND.n540 585
R9209 GND.n7869 GND.n540 585
R9210 GND.n7863 GND.n7862 585
R9211 GND.n7862 GND.n7861 585
R9212 GND.n563 GND.n562 585
R9213 GND.n7846 GND.n563 585
R9214 GND.n7852 GND.n7851 585
R9215 GND.n7853 GND.n7852 585
R9216 GND.n575 GND.n574 585
R9217 GND.n7837 GND.n574 585
R9218 GND.n7822 GND.n586 585
R9219 GND.n7834 GND.n586 585
R9220 GND.n7823 GND.n597 585
R9221 GND.n7809 GND.n597 585
R9222 GND.n7825 GND.n7824 585
R9223 GND.n7826 GND.n7825 585
R9224 GND.n598 GND.n596 585
R9225 GND.n7815 GND.n596 585
R9226 GND.n7786 GND.n7785 585
R9227 GND.n7785 GND.n7784 585
R9228 GND.n7787 GND.n612 585
R9229 GND.n7801 GND.n612 585
R9230 GND.n7788 GND.n624 585
R9231 GND.n7778 GND.n624 585
R9232 GND.n7790 GND.n7789 585
R9233 GND.n7791 GND.n7790 585
R9234 GND.n625 GND.n623 585
R9235 GND.n7774 GND.n623 585
R9236 GND.n7743 GND.n7742 585
R9237 GND.n7742 GND.n7741 585
R9238 GND.n7740 GND.n640 585
R9239 GND.n7764 GND.n640 585
R9240 GND.n654 GND.n652 585
R9241 GND.n7747 GND.n652 585
R9242 GND.n7753 GND.n7752 585
R9243 GND.n7754 GND.n7753 585
R9244 GND.n653 GND.n651 585
R9245 GND.n7737 GND.n651 585
R9246 GND.n698 GND.n697 585
R9247 GND.n700 GND.n699 585
R9248 GND.n703 GND.n702 585
R9249 GND.n704 GND.n664 585
R9250 GND.n670 GND.n669 585
R9251 GND.n7728 GND.n7727 585
R9252 GND.n7729 GND.n666 585
R9253 GND.n7725 GND.n659 585
R9254 GND.n8450 GND.n8449 585
R9255 GND.n357 GND.n356 585
R9256 GND.n379 GND.n378 585
R9257 GND.n361 GND.n360 585
R9258 GND.n374 GND.n373 585
R9259 GND.n372 GND.n371 585
R9260 GND.n370 GND.n369 585
R9261 GND.n364 GND.n363 585
R9262 GND.n365 GND.n347 585
R9263 GND.n8447 GND.n347 585
R9264 GND.n8453 GND.n345 585
R9265 GND.n8463 GND.n345 585
R9266 GND.n8455 GND.n8454 585
R9267 GND.n8456 GND.n8455 585
R9268 GND.n351 GND.n335 585
R9269 GND.n8469 GND.n335 585
R9270 GND.n8242 GND.n8241 585
R9271 GND.n8241 GND.n8240 585
R9272 GND.n8243 GND.n325 585
R9273 GND.n8475 GND.n325 585
R9274 GND.n8245 GND.n8244 585
R9275 GND.n8246 GND.n8245 585
R9276 GND.n394 GND.n315 585
R9277 GND.n8481 GND.n315 585
R9278 GND.n8230 GND.n8229 585
R9279 GND.n8231 GND.n8230 585
R9280 GND.n400 GND.n305 585
R9281 GND.n8487 GND.n305 585
R9282 GND.n8224 GND.n8223 585
R9283 GND.n8223 GND.n8222 585
R9284 GND.n402 GND.n294 585
R9285 GND.n8493 GND.n294 585
R9286 GND.n8214 GND.n8213 585
R9287 GND.n8215 GND.n8214 585
R9288 GND.n404 GND.n284 585
R9289 GND.n8499 GND.n284 585
R9290 GND.n8209 GND.n8208 585
R9291 GND.n8208 GND.n8207 585
R9292 GND.n406 GND.n273 585
R9293 GND.n8505 GND.n273 585
R9294 GND.n8199 GND.n8198 585
R9295 GND.n8200 GND.n8199 585
R9296 GND.n408 GND.n263 585
R9297 GND.n8511 GND.n263 585
R9298 GND.n8194 GND.n8193 585
R9299 GND.n8193 GND.n8192 585
R9300 GND.n410 GND.n253 585
R9301 GND.n8517 GND.n253 585
R9302 GND.n8184 GND.n8183 585
R9303 GND.n8185 GND.n8184 585
R9304 GND.n413 GND.n243 585
R9305 GND.n8523 GND.n243 585
R9306 GND.n8179 GND.n8178 585
R9307 GND.n8178 GND.n8177 585
R9308 GND.n415 GND.n232 585
R9309 GND.n8529 GND.n232 585
R9310 GND.n8169 GND.n8168 585
R9311 GND.n8170 GND.n8169 585
R9312 GND.n417 GND.n222 585
R9313 GND.n8535 GND.n222 585
R9314 GND.n8164 GND.n8163 585
R9315 GND.n8163 GND.n8162 585
R9316 GND.n419 GND.n211 585
R9317 GND.n8541 GND.n211 585
R9318 GND.n8154 GND.n8153 585
R9319 GND.n8155 GND.n8154 585
R9320 GND.n421 GND.n201 585
R9321 GND.n8547 GND.n201 585
R9322 GND.n8149 GND.n8148 585
R9323 GND.n8148 GND.n8147 585
R9324 GND.n423 GND.n191 585
R9325 GND.n8553 GND.n191 585
R9326 GND.n8139 GND.n8138 585
R9327 GND.n8140 GND.n8139 585
R9328 GND.n425 GND.n179 585
R9329 GND.n8559 GND.n179 585
R9330 GND.n8134 GND.n8133 585
R9331 GND.n8133 GND.n8132 585
R9332 GND.n428 GND.n427 585
R9333 GND.n8125 GND.n428 585
R9334 GND.n157 GND.n155 585
R9335 GND.n435 GND.n157 585
R9336 GND.n8568 GND.n8567 585
R9337 GND.n8567 GND.n8566 585
R9338 GND.n156 GND.n154 585
R9339 GND.n8032 GND.n156 585
R9340 GND.n8001 GND.n8000 585
R9341 GND.n8000 GND.n441 585
R9342 GND.n8002 GND.n450 585
R9343 GND.n8020 GND.n450 585
R9344 GND.n8003 GND.n456 585
R9345 GND.n8015 GND.n456 585
R9346 GND.n8005 GND.n8004 585
R9347 GND.n8006 GND.n8005 585
R9348 GND.n464 GND.n463 585
R9349 GND.n7974 GND.n463 585
R9350 GND.n7993 GND.n7992 585
R9351 GND.n7992 GND.n7991 585
R9352 GND.n467 GND.n466 585
R9353 GND.n7968 GND.n467 585
R9354 GND.n7961 GND.n480 585
R9355 GND.n7981 GND.n480 585
R9356 GND.n7963 GND.n7962 585
R9357 GND.n7964 GND.n7963 585
R9358 GND.n491 GND.n490 585
R9359 GND.n7937 GND.n490 585
R9360 GND.n7956 GND.n7955 585
R9361 GND.n7955 GND.n7954 585
R9362 GND.n494 GND.n493 585
R9363 GND.n549 GND.n494 585
R9364 GND.n7879 GND.n507 585
R9365 GND.n7944 GND.n507 585
R9366 GND.n7881 GND.n7880 585
R9367 GND.n7882 GND.n7881 585
R9368 GND.n553 GND.n528 585
R9369 GND.n7899 GND.n528 585
R9370 GND.n7874 GND.n7873 585
R9371 GND.n7873 GND.n526 585
R9372 GND.n7872 GND.n538 585
R9373 GND.n7891 GND.n538 585
R9374 GND.n7871 GND.n7870 585
R9375 GND.n7870 GND.n7869 585
R9376 GND.n557 GND.n555 585
R9377 GND.n7861 GND.n557 585
R9378 GND.n7845 GND.n7844 585
R9379 GND.n7846 GND.n7845 585
R9380 GND.n578 GND.n572 585
R9381 GND.n7853 GND.n572 585
R9382 GND.n7839 GND.n7838 585
R9383 GND.n7838 GND.n7837 585
R9384 GND.n581 GND.n580 585
R9385 GND.n7834 GND.n581 585
R9386 GND.n7811 GND.n7810 585
R9387 GND.n7810 GND.n7809 585
R9388 GND.n7812 GND.n594 585
R9389 GND.n7826 GND.n594 585
R9390 GND.n7814 GND.n7813 585
R9391 GND.n7815 GND.n7814 585
R9392 GND.n605 GND.n604 585
R9393 GND.n7784 GND.n604 585
R9394 GND.n7803 GND.n7802 585
R9395 GND.n7802 GND.n7801 585
R9396 GND.n608 GND.n607 585
R9397 GND.n7778 GND.n608 585
R9398 GND.n7771 GND.n621 585
R9399 GND.n7791 GND.n621 585
R9400 GND.n7773 GND.n7772 585
R9401 GND.n7774 GND.n7773 585
R9402 GND.n633 GND.n632 585
R9403 GND.n7741 GND.n632 585
R9404 GND.n7766 GND.n7765 585
R9405 GND.n7765 GND.n7764 585
R9406 GND.n636 GND.n635 585
R9407 GND.n7747 GND.n636 585
R9408 GND.n7734 GND.n649 585
R9409 GND.n7754 GND.n649 585
R9410 GND.n7736 GND.n7735 585
R9411 GND.n7737 GND.n7736 585
R9412 GND.n6915 GND.n1079 585
R9413 GND.n1079 GND.n1037 585
R9414 GND.n6914 GND.n6913 585
R9415 GND.n6913 GND.n1041 585
R9416 GND.n6912 GND.n1047 585
R9417 GND.n6992 GND.n1047 585
R9418 GND.n1083 GND.n1082 585
R9419 GND.n1082 GND.n1081 585
R9420 GND.n6908 GND.n1056 585
R9421 GND.n6979 GND.n1056 585
R9422 GND.n6907 GND.n6906 585
R9423 GND.n6906 GND.n6905 585
R9424 GND.n1086 GND.n1085 585
R9425 GND.n6894 GND.n1086 585
R9426 GND.n6737 GND.n6736 585
R9427 GND.n6736 GND.n6735 585
R9428 GND.n6738 GND.n1102 585
R9429 GND.n6886 GND.n1102 585
R9430 GND.n6740 GND.n6739 585
R9431 GND.n6741 GND.n6740 585
R9432 GND.n6720 GND.n1111 585
R9433 GND.t209 GND.n1111 585
R9434 GND.n6728 GND.n6727 585
R9435 GND.n6727 GND.n6710 585
R9436 GND.n6726 GND.n1119 585
R9437 GND.n6866 GND.n1119 585
R9438 GND.n6725 GND.n6724 585
R9439 GND.n6724 GND.n1203 585
R9440 GND.n1195 GND.n1127 585
R9441 GND.n6858 GND.n1127 585
R9442 GND.n6791 GND.n6790 585
R9443 GND.n6790 GND.n6789 585
R9444 GND.n6792 GND.n1135 585
R9445 GND.n6850 GND.n1135 585
R9446 GND.n6794 GND.n6793 585
R9447 GND.t203 GND.n6794 585
R9448 GND.n1182 GND.n1143 585
R9449 GND.n6842 GND.n1143 585
R9450 GND.n6805 GND.n6804 585
R9451 GND.n6804 GND.n6803 585
R9452 GND.n6806 GND.n1151 585
R9453 GND.n6834 GND.n1151 585
R9454 GND.n6808 GND.n6807 585
R9455 GND.n6809 GND.n6808 585
R9456 GND.n1178 GND.n1159 585
R9457 GND.n6826 GND.n1159 585
R9458 GND.n6462 GND.n6461 585
R9459 GND.n6461 GND.n6460 585
R9460 GND.n6463 GND.n1167 585
R9461 GND.t213 GND.n1167 585
R9462 GND.n6465 GND.n6464 585
R9463 GND.n6464 GND.n1210 585
R9464 GND.n6466 GND.n1216 585
R9465 GND.n6672 GND.n1216 585
R9466 GND.n6468 GND.n6467 585
R9467 GND.n6467 GND.n1214 585
R9468 GND.n6469 GND.n1224 585
R9469 GND.n6664 GND.n1224 585
R9470 GND.n6471 GND.n6470 585
R9471 GND.n6470 GND.n1397 585
R9472 GND.n6472 GND.n1233 585
R9473 GND.n6647 GND.n1233 585
R9474 GND.n6474 GND.n6473 585
R9475 GND.t199 GND.n6474 585
R9476 GND.n1408 GND.n1241 585
R9477 GND.n6639 GND.n1241 585
R9478 GND.n6447 GND.n6446 585
R9479 GND.n6446 GND.n6445 585
R9480 GND.n6444 GND.n1249 585
R9481 GND.n6631 GND.n1249 585
R9482 GND.n6443 GND.n6442 585
R9483 GND.n6442 GND.n1379 585
R9484 GND.n1410 GND.n1257 585
R9485 GND.n6623 GND.n1257 585
R9486 GND.n6438 GND.n6437 585
R9487 GND.n6437 GND.n1372 585
R9488 GND.n6436 GND.n1265 585
R9489 GND.t207 GND.n1265 585
R9490 GND.n6435 GND.n6434 585
R9491 GND.n6434 GND.n1365 585
R9492 GND.n1412 GND.n1273 585
R9493 GND.n6608 GND.n1273 585
R9494 GND.n6430 GND.n6429 585
R9495 GND.n6429 GND.n1358 585
R9496 GND.n6428 GND.n1281 585
R9497 GND.n6600 GND.n1281 585
R9498 GND.n6427 GND.n6426 585
R9499 GND.n6426 GND.n1351 585
R9500 GND.n1414 GND.n1289 585
R9501 GND.n6592 GND.n1289 585
R9502 GND.n6422 GND.n6421 585
R9503 GND.n6421 GND.t201 585
R9504 GND.n6420 GND.n1297 585
R9505 GND.n6584 GND.n1297 585
R9506 GND.n6419 GND.n6418 585
R9507 GND.n6418 GND.n1339 585
R9508 GND.n1416 GND.n1305 585
R9509 GND.n6576 GND.n1305 585
R9510 GND.n6414 GND.n6413 585
R9511 GND.n6413 GND.n1335 585
R9512 GND.n6412 GND.n1312 585
R9513 GND.n6568 GND.n1312 585
R9514 GND.n6411 GND.n6410 585
R9515 GND.n6410 GND.n1329 585
R9516 GND.n1418 GND.n1320 585
R9517 GND.t211 GND.n1320 585
R9518 GND.n6406 GND.n6405 585
R9519 GND.n6405 GND.n6404 585
R9520 GND.n1421 GND.n1420 585
R9521 GND.n6245 GND.n1421 585
R9522 GND.n6234 GND.n1429 585
R9523 GND.n6394 GND.n1429 585
R9524 GND.n6236 GND.n6235 585
R9525 GND.n6237 GND.n6236 585
R9526 GND.n6206 GND.n1438 585
R9527 GND.n6384 GND.n1438 585
R9528 GND.n6229 GND.n6228 585
R9529 GND.n6228 GND.n6199 585
R9530 GND.n6227 GND.n1446 585
R9531 GND.t195 GND.n1446 585
R9532 GND.n6226 GND.n6225 585
R9533 GND.n6225 GND.n6192 585
R9534 GND.n6208 GND.n1454 585
R9535 GND.n6369 GND.n1454 585
R9536 GND.n6221 GND.n6220 585
R9537 GND.n6220 GND.n6185 585
R9538 GND.n6219 GND.n1462 585
R9539 GND.n6361 GND.n1462 585
R9540 GND.n6218 GND.n6217 585
R9541 GND.n6217 GND.n6178 585
R9542 GND.n6210 GND.n1470 585
R9543 GND.n6353 GND.n1470 585
R9544 GND.n6213 GND.n6212 585
R9545 GND.n6212 GND.t205 585
R9546 GND.n1517 GND.n1478 585
R9547 GND.n6345 GND.n1478 585
R9548 GND.n6308 GND.n6307 585
R9549 GND.n6307 GND.n6306 585
R9550 GND.n6309 GND.n1486 585
R9551 GND.n6337 GND.n1486 585
R9552 GND.n6311 GND.n6310 585
R9553 GND.n6312 GND.n6311 585
R9554 GND.n1513 GND.n1494 585
R9555 GND.n6329 GND.n1494 585
R9556 GND.n5613 GND.n5612 585
R9557 GND.n5612 GND.n5611 585
R9558 GND.n5614 GND.n1502 585
R9559 GND.t197 GND.n1502 585
R9560 GND.n5616 GND.n5615 585
R9561 GND.n5615 GND.n1531 585
R9562 GND.n5617 GND.n1537 585
R9563 GND.n6150 GND.n1537 585
R9564 GND.n5619 GND.n5618 585
R9565 GND.n5618 GND.n1535 585
R9566 GND.n5620 GND.n1545 585
R9567 GND.n6142 GND.n1545 585
R9568 GND.n5622 GND.n5621 585
R9569 GND.n5623 GND.n5622 585
R9570 GND.n5590 GND.n1554 585
R9571 GND.n6125 GND.n1554 585
R9572 GND.n5600 GND.n5599 585
R9573 GND.n5599 GND.n5598 585
R9574 GND.n5597 GND.n1561 585
R9575 GND.n6117 GND.n1561 585
R9576 GND.n5596 GND.n5593 585
R9577 GND.n5593 GND.n5200 585
R9578 GND.n5592 GND.n1568 585
R9579 GND.n6109 GND.n1568 585
R9580 GND.n6098 GND.n6097 585
R9581 GND.n6096 GND.n1587 585
R9582 GND.n6095 GND.n1586 585
R9583 GND.n6100 GND.n1586 585
R9584 GND.n6094 GND.n6093 585
R9585 GND.n6092 GND.n6091 585
R9586 GND.n6090 GND.n6089 585
R9587 GND.n6088 GND.n1594 585
R9588 GND.n6086 GND.n6053 585
R9589 GND.n6085 GND.n6054 585
R9590 GND.n6083 GND.n6055 585
R9591 GND.n6082 GND.n6056 585
R9592 GND.n6080 GND.n6057 585
R9593 GND.n6079 GND.n6058 585
R9594 GND.n6077 GND.n6059 585
R9595 GND.n6076 GND.n6060 585
R9596 GND.n6074 GND.n6061 585
R9597 GND.n6072 GND.n6064 585
R9598 GND.n6071 GND.n6070 585
R9599 GND.n6069 GND.n6066 585
R9600 GND.n6067 GND.n1566 585
R9601 GND.n6100 GND.n1566 585
R9602 GND.n6971 GND.n6970 585
R9603 GND.n6963 GND.n1067 585
R9604 GND.n6965 GND.n6964 585
R9605 GND.n6961 GND.n1068 585
R9606 GND.n6960 GND.n6959 585
R9607 GND.n6954 GND.n6953 585
R9608 GND.n6952 GND.n1070 585
R9609 GND.n6950 GND.n6949 585
R9610 GND.n6947 GND.n1071 585
R9611 GND.n6945 GND.n6944 585
R9612 GND.n6942 GND.n1072 585
R9613 GND.n6940 GND.n6939 585
R9614 GND.n6937 GND.n1073 585
R9615 GND.n6935 GND.n6934 585
R9616 GND.n6932 GND.n1074 585
R9617 GND.n6930 GND.n6929 585
R9618 GND.n1076 GND.n1075 585
R9619 GND.n6924 GND.n6923 585
R9620 GND.n6921 GND.n1078 585
R9621 GND.n6919 GND.n6918 585
R9622 GND.n6972 GND.n1065 585
R9623 GND.n6972 GND.n1037 585
R9624 GND.n6974 GND.n6973 585
R9625 GND.n6973 GND.n1041 585
R9626 GND.n6975 GND.n1048 585
R9627 GND.n6992 GND.n1048 585
R9628 GND.n6976 GND.n1059 585
R9629 GND.n1081 GND.n1059 585
R9630 GND.n6978 GND.n6977 585
R9631 GND.n6979 GND.n6978 585
R9632 GND.n1060 GND.n1058 585
R9633 GND.n6905 GND.n1058 585
R9634 GND.n6882 GND.n1095 585
R9635 GND.n6894 GND.n1095 585
R9636 GND.n6883 GND.n1105 585
R9637 GND.n6735 GND.n1105 585
R9638 GND.n6885 GND.n6884 585
R9639 GND.n6886 GND.n6885 585
R9640 GND.n1106 GND.n1104 585
R9641 GND.n6741 GND.n1104 585
R9642 GND.n6875 GND.n6874 585
R9643 GND.n6874 GND.t209 585
R9644 GND.n1109 GND.n1108 585
R9645 GND.n6710 GND.n1109 585
R9646 GND.n6865 GND.n6864 585
R9647 GND.n6866 GND.n6865 585
R9648 GND.n1122 GND.n1121 585
R9649 GND.n1203 GND.n1121 585
R9650 GND.n6860 GND.n6859 585
R9651 GND.n6859 GND.n6858 585
R9652 GND.n1125 GND.n1124 585
R9653 GND.n6789 GND.n1125 585
R9654 GND.n6849 GND.n6848 585
R9655 GND.n6850 GND.n6849 585
R9656 GND.n1138 GND.n1137 585
R9657 GND.t203 GND.n1137 585
R9658 GND.n6844 GND.n6843 585
R9659 GND.n6843 GND.n6842 585
R9660 GND.n1141 GND.n1140 585
R9661 GND.n6803 GND.n1141 585
R9662 GND.n6833 GND.n6832 585
R9663 GND.n6834 GND.n6833 585
R9664 GND.n1154 GND.n1153 585
R9665 GND.n6809 GND.n1153 585
R9666 GND.n6828 GND.n6827 585
R9667 GND.n6827 GND.n6826 585
R9668 GND.n1157 GND.n1156 585
R9669 GND.n6460 GND.n1157 585
R9670 GND.n6657 GND.n1168 585
R9671 GND.t213 GND.n1168 585
R9672 GND.n6659 GND.n6658 585
R9673 GND.n6658 GND.n1210 585
R9674 GND.n6660 GND.n1217 585
R9675 GND.n6672 GND.n1217 585
R9676 GND.n6661 GND.n1227 585
R9677 GND.n1227 GND.n1214 585
R9678 GND.n6663 GND.n6662 585
R9679 GND.n6664 GND.n6663 585
R9680 GND.n1228 GND.n1226 585
R9681 GND.n1397 GND.n1226 585
R9682 GND.n6649 GND.n6648 585
R9683 GND.n6648 GND.n6647 585
R9684 GND.n1231 GND.n1230 585
R9685 GND.t199 GND.n1231 585
R9686 GND.n6638 GND.n6637 585
R9687 GND.n6639 GND.n6638 585
R9688 GND.n1244 GND.n1243 585
R9689 GND.n6445 GND.n1243 585
R9690 GND.n6633 GND.n6632 585
R9691 GND.n6632 GND.n6631 585
R9692 GND.n1247 GND.n1246 585
R9693 GND.n1379 GND.n1247 585
R9694 GND.n6622 GND.n6621 585
R9695 GND.n6623 GND.n6622 585
R9696 GND.n1260 GND.n1259 585
R9697 GND.n1372 GND.n1259 585
R9698 GND.n6617 GND.n6616 585
R9699 GND.n6616 GND.t207 585
R9700 GND.n1263 GND.n1262 585
R9701 GND.n1365 GND.n1263 585
R9702 GND.n6607 GND.n6606 585
R9703 GND.n6608 GND.n6607 585
R9704 GND.n1276 GND.n1275 585
R9705 GND.n1358 GND.n1275 585
R9706 GND.n6602 GND.n6601 585
R9707 GND.n6601 GND.n6600 585
R9708 GND.n1279 GND.n1278 585
R9709 GND.n1351 GND.n1279 585
R9710 GND.n6591 GND.n6590 585
R9711 GND.n6592 GND.n6591 585
R9712 GND.n1292 GND.n1291 585
R9713 GND.t201 GND.n1291 585
R9714 GND.n6586 GND.n6585 585
R9715 GND.n6585 GND.n6584 585
R9716 GND.n1295 GND.n1294 585
R9717 GND.n1339 GND.n1295 585
R9718 GND.n6575 GND.n6574 585
R9719 GND.n6576 GND.n6575 585
R9720 GND.n1308 GND.n1307 585
R9721 GND.n1335 GND.n1307 585
R9722 GND.n6570 GND.n6569 585
R9723 GND.n6569 GND.n6568 585
R9724 GND.n1311 GND.n1310 585
R9725 GND.n1329 GND.n1311 585
R9726 GND.n6401 GND.n1321 585
R9727 GND.t211 GND.n1321 585
R9728 GND.n6403 GND.n6402 585
R9729 GND.n6404 GND.n6403 585
R9730 GND.n1424 GND.n1423 585
R9731 GND.n6245 GND.n1423 585
R9732 GND.n6396 GND.n6395 585
R9733 GND.n6395 GND.n6394 585
R9734 GND.n1427 GND.n1426 585
R9735 GND.n6237 GND.n1427 585
R9736 GND.n6383 GND.n6382 585
R9737 GND.n6384 GND.n6383 585
R9738 GND.n1441 GND.n1440 585
R9739 GND.n6199 GND.n1440 585
R9740 GND.n6378 GND.n6377 585
R9741 GND.n6377 GND.t195 585
R9742 GND.n1444 GND.n1443 585
R9743 GND.n6192 GND.n1444 585
R9744 GND.n6368 GND.n6367 585
R9745 GND.n6369 GND.n6368 585
R9746 GND.n1457 GND.n1456 585
R9747 GND.n6185 GND.n1456 585
R9748 GND.n6363 GND.n6362 585
R9749 GND.n6362 GND.n6361 585
R9750 GND.n1460 GND.n1459 585
R9751 GND.n6178 GND.n1460 585
R9752 GND.n6352 GND.n6351 585
R9753 GND.n6353 GND.n6352 585
R9754 GND.n1473 GND.n1472 585
R9755 GND.t205 GND.n1472 585
R9756 GND.n6347 GND.n6346 585
R9757 GND.n6346 GND.n6345 585
R9758 GND.n1476 GND.n1475 585
R9759 GND.n6306 GND.n1476 585
R9760 GND.n6336 GND.n6335 585
R9761 GND.n6337 GND.n6336 585
R9762 GND.n1489 GND.n1488 585
R9763 GND.n6312 GND.n1488 585
R9764 GND.n6331 GND.n6330 585
R9765 GND.n6330 GND.n6329 585
R9766 GND.n1492 GND.n1491 585
R9767 GND.n5611 GND.n1492 585
R9768 GND.n6135 GND.n1503 585
R9769 GND.t197 GND.n1503 585
R9770 GND.n6137 GND.n6136 585
R9771 GND.n6136 GND.n1531 585
R9772 GND.n6138 GND.n1538 585
R9773 GND.n6150 GND.n1538 585
R9774 GND.n6139 GND.n1548 585
R9775 GND.n1548 GND.n1535 585
R9776 GND.n6141 GND.n6140 585
R9777 GND.n6142 GND.n6141 585
R9778 GND.n1549 GND.n1547 585
R9779 GND.n5623 GND.n1547 585
R9780 GND.n6127 GND.n6126 585
R9781 GND.n6126 GND.n6125 585
R9782 GND.n1552 GND.n1551 585
R9783 GND.n5598 GND.n1552 585
R9784 GND.n6116 GND.n6115 585
R9785 GND.n6117 GND.n6116 585
R9786 GND.n1564 GND.n1563 585
R9787 GND.n5200 GND.n1563 585
R9788 GND.n6111 GND.n6110 585
R9789 GND.n6110 GND.n6109 585
R9790 GND.n7538 GND.n765 585
R9791 GND.n7425 GND.n765 585
R9792 GND.n7537 GND.n7536 585
R9793 GND.n7536 GND.n7535 585
R9794 GND.n797 GND.n796 585
R9795 GND.n798 GND.n797 585
R9796 GND.n7440 GND.n7439 585
R9797 GND.n7441 GND.n7440 585
R9798 GND.n7438 GND.n809 585
R9799 GND.n809 GND.n806 585
R9800 GND.n7437 GND.n7436 585
R9801 GND.n7436 GND.n7435 585
R9802 GND.n811 GND.n810 585
R9803 GND.n817 GND.n811 585
R9804 GND.n7367 GND.n7366 585
R9805 GND.n7368 GND.n7367 585
R9806 GND.n7365 GND.n819 585
R9807 GND.n7361 GND.n819 585
R9808 GND.n7364 GND.n7363 585
R9809 GND.n7363 GND.n7362 585
R9810 GND.n821 GND.n820 585
R9811 GND.t36 GND.n821 585
R9812 GND.n7340 GND.n836 585
R9813 GND.n836 GND.n830 585
R9814 GND.n7342 GND.n7341 585
R9815 GND.n7343 GND.n7342 585
R9816 GND.n7339 GND.n835 585
R9817 GND.n840 GND.n835 585
R9818 GND.n7338 GND.n7337 585
R9819 GND.n7337 GND.n7336 585
R9820 GND.n838 GND.n837 585
R9821 GND.n7313 GND.n838 585
R9822 GND.n7325 GND.n7324 585
R9823 GND.n7326 GND.n7325 585
R9824 GND.n7323 GND.n849 585
R9825 GND.n849 GND.n846 585
R9826 GND.n7322 GND.n7321 585
R9827 GND.n7321 GND.n7320 585
R9828 GND.n851 GND.n850 585
R9829 GND.n858 GND.n851 585
R9830 GND.n7307 GND.n7306 585
R9831 GND.n7308 GND.n7307 585
R9832 GND.n7305 GND.n860 585
R9833 GND.n860 GND.n857 585
R9834 GND.n7304 GND.n7303 585
R9835 GND.n7303 GND.n7302 585
R9836 GND.n862 GND.n861 585
R9837 GND.n873 GND.n862 585
R9838 GND.n7289 GND.n7288 585
R9839 GND.n7290 GND.n7289 585
R9840 GND.n7287 GND.n874 585
R9841 GND.n874 GND.n871 585
R9842 GND.n7286 GND.n7285 585
R9843 GND.n7285 GND.n7284 585
R9844 GND.n876 GND.n875 585
R9845 GND.n877 GND.n876 585
R9846 GND.n7271 GND.n7270 585
R9847 GND.n7272 GND.n7271 585
R9848 GND.n7269 GND.n884 585
R9849 GND.n7265 GND.n884 585
R9850 GND.n7268 GND.n7267 585
R9851 GND.n7267 GND.n7266 585
R9852 GND.n886 GND.n885 585
R9853 GND.n892 GND.n886 585
R9854 GND.n7258 GND.n7257 585
R9855 GND.n7259 GND.n7258 585
R9856 GND.n7256 GND.n894 585
R9857 GND.n7252 GND.n894 585
R9858 GND.n7255 GND.n7254 585
R9859 GND.n7254 GND.n7253 585
R9860 GND.n896 GND.n895 585
R9861 GND.n902 GND.n896 585
R9862 GND.n7245 GND.n7244 585
R9863 GND.n7246 GND.n7245 585
R9864 GND.n7243 GND.n904 585
R9865 GND.n904 GND.n901 585
R9866 GND.n7242 GND.n7241 585
R9867 GND.n7241 GND.n7240 585
R9868 GND.n906 GND.n905 585
R9869 GND.n916 GND.n906 585
R9870 GND.n7209 GND.n7208 585
R9871 GND.n7210 GND.n7209 585
R9872 GND.n7207 GND.n917 585
R9873 GND.n7202 GND.n917 585
R9874 GND.n7206 GND.n7205 585
R9875 GND.n7205 GND.n7204 585
R9876 GND.n919 GND.n918 585
R9877 GND.n920 GND.n919 585
R9878 GND.n7190 GND.n7189 585
R9879 GND.n7191 GND.n7190 585
R9880 GND.n7188 GND.n926 585
R9881 GND.n7184 GND.n926 585
R9882 GND.n7187 GND.n7186 585
R9883 GND.n7186 GND.n7185 585
R9884 GND.n928 GND.n927 585
R9885 GND.n934 GND.n928 585
R9886 GND.n7176 GND.n7175 585
R9887 GND.n7177 GND.n7176 585
R9888 GND.n7174 GND.n936 585
R9889 GND.n936 GND.n933 585
R9890 GND.n7173 GND.n7172 585
R9891 GND.n7172 GND.n7171 585
R9892 GND.n938 GND.n937 585
R9893 GND.n949 GND.n938 585
R9894 GND.n7149 GND.n7148 585
R9895 GND.n7150 GND.n7149 585
R9896 GND.n7147 GND.n950 585
R9897 GND.n950 GND.n947 585
R9898 GND.n7146 GND.n7145 585
R9899 GND.n7145 GND.n7144 585
R9900 GND.n952 GND.n951 585
R9901 GND.n953 GND.n952 585
R9902 GND.n7131 GND.n7130 585
R9903 GND.n7132 GND.n7131 585
R9904 GND.n7129 GND.n960 585
R9905 GND.n965 GND.n960 585
R9906 GND.n7128 GND.n7127 585
R9907 GND.n7127 GND.n7126 585
R9908 GND.n962 GND.n961 585
R9909 GND.n963 GND.n962 585
R9910 GND.n7110 GND.n7109 585
R9911 GND.n7111 GND.n7110 585
R9912 GND.n7108 GND.n975 585
R9913 GND.n975 GND.n972 585
R9914 GND.n7107 GND.n7106 585
R9915 GND.n7106 GND.n7105 585
R9916 GND.n977 GND.n976 585
R9917 GND.n984 GND.n977 585
R9918 GND.n7093 GND.n7092 585
R9919 GND.n7094 GND.n7093 585
R9920 GND.n7091 GND.n986 585
R9921 GND.n986 GND.n983 585
R9922 GND.n7090 GND.n7089 585
R9923 GND.n7089 GND.n7088 585
R9924 GND.n988 GND.n987 585
R9925 GND.n999 GND.n988 585
R9926 GND.n7075 GND.n7074 585
R9927 GND.n7076 GND.n7075 585
R9928 GND.n7073 GND.n1000 585
R9929 GND.n1000 GND.n997 585
R9930 GND.n7072 GND.n7071 585
R9931 GND.n7071 GND.n7070 585
R9932 GND.n1002 GND.n1001 585
R9933 GND.n1003 GND.n1002 585
R9934 GND.n7057 GND.n7056 585
R9935 GND.n7058 GND.n7057 585
R9936 GND.n7055 GND.n1010 585
R9937 GND.n7051 GND.n1010 585
R9938 GND.n7054 GND.n7053 585
R9939 GND.n7053 GND.n7052 585
R9940 GND.n1012 GND.n1011 585
R9941 GND.n1018 GND.n1012 585
R9942 GND.n7044 GND.n7043 585
R9943 GND.n7045 GND.n7044 585
R9944 GND.n7042 GND.n1020 585
R9945 GND.n1020 GND.n1017 585
R9946 GND.n7041 GND.n7040 585
R9947 GND.n7040 GND.n7039 585
R9948 GND.n1022 GND.n1021 585
R9949 GND.n1033 GND.n1022 585
R9950 GND.n7017 GND.n7016 585
R9951 GND.n7018 GND.n7017 585
R9952 GND.n7015 GND.n1034 585
R9953 GND.n7010 GND.n1034 585
R9954 GND.n7014 GND.n7013 585
R9955 GND.n7013 GND.n7012 585
R9956 GND.n1036 GND.n1035 585
R9957 GND.n7000 GND.n1036 585
R9958 GND.n6998 GND.n6997 585
R9959 GND.n6999 GND.n6998 585
R9960 GND.n6996 GND.n1042 585
R9961 GND.n6747 GND.n1042 585
R9962 GND.n6995 GND.n6994 585
R9963 GND.n6994 GND.n6993 585
R9964 GND.n1044 GND.n1043 585
R9965 GND.n1045 GND.n1044 585
R9966 GND.n6900 GND.n6899 585
R9967 GND.n6899 GND.n1057 585
R9968 GND.n6901 GND.n1090 585
R9969 GND.n1090 GND.n1055 585
R9970 GND.n6903 GND.n6902 585
R9971 GND.n6904 GND.n6903 585
R9972 GND.n6898 GND.n1089 585
R9973 GND.n1089 GND.n1087 585
R9974 GND.n6897 GND.n6896 585
R9975 GND.n6896 GND.n6895 585
R9976 GND.n1092 GND.n1091 585
R9977 GND.n1093 GND.n1092 585
R9978 GND.n6717 GND.n6716 585
R9979 GND.n6716 GND.n1103 585
R9980 GND.n6719 GND.n6718 585
R9981 GND.n6719 GND.n1101 585
R9982 GND.n6768 GND.n6715 585
R9983 GND.n6768 GND.n6767 585
R9984 GND.n6770 GND.n6769 585
R9985 GND.n6769 GND.n1112 585
R9986 GND.n6771 GND.n6712 585
R9987 GND.n6712 GND.n1110 585
R9988 GND.n6773 GND.n6772 585
R9989 GND.n6774 GND.n6773 585
R9990 GND.n6714 GND.n6711 585
R9991 GND.n6711 GND.n1120 585
R9992 GND.n6713 GND.n1202 585
R9993 GND.n1202 GND.n1118 585
R9994 GND.n6782 GND.n1201 585
R9995 GND.n6782 GND.n6781 585
R9996 GND.n6784 GND.n6783 585
R9997 GND.n6783 GND.n1128 585
R9998 GND.n6785 GND.n1198 585
R9999 GND.n1198 GND.n1126 585
R10000 GND.n6787 GND.n6786 585
R10001 GND.n6788 GND.n6787 585
R10002 GND.n1200 GND.n1197 585
R10003 GND.n1197 GND.n1136 585
R10004 GND.n1199 GND.n1189 585
R10005 GND.n1189 GND.n1134 585
R10006 GND.n6796 GND.n1188 585
R10007 GND.n6796 GND.n6795 585
R10008 GND.n6798 GND.n6797 585
R10009 GND.n6797 GND.n1144 585
R10010 GND.n6799 GND.n1185 585
R10011 GND.n1185 GND.n1142 585
R10012 GND.n6801 GND.n6800 585
R10013 GND.n6802 GND.n6801 585
R10014 GND.n1187 GND.n1184 585
R10015 GND.n1184 GND.n1152 585
R10016 GND.n1186 GND.n1175 585
R10017 GND.n1175 GND.n1150 585
R10018 GND.n6811 GND.n1176 585
R10019 GND.n6811 GND.n6810 585
R10020 GND.n6812 GND.n1174 585
R10021 GND.n6812 GND.n1160 585
R10022 GND.n6814 GND.n6813 585
R10023 GND.n6813 GND.n1158 585
R10024 GND.n6815 GND.n1172 585
R10025 GND.n1172 GND.n1170 585
R10026 GND.n6817 GND.n6816 585
R10027 GND.n6818 GND.n6817 585
R10028 GND.n1173 GND.n1171 585
R10029 GND.n1171 GND.n1166 585
R10030 GND.n6678 GND.n6677 585
R10031 GND.n6679 GND.n6678 585
R10032 GND.n6676 GND.n1211 585
R10033 GND.n1211 GND.n1209 585
R10034 GND.n6675 GND.n6674 585
R10035 GND.n6674 GND.n6673 585
R10036 GND.n1213 GND.n1212 585
R10037 GND.n1391 GND.n1213 585
R10038 GND.n6481 GND.n6480 585
R10039 GND.n6480 GND.n1225 585
R10040 GND.n6482 GND.n1399 585
R10041 GND.n1399 GND.n1223 585
R10042 GND.n6484 GND.n6483 585
R10043 GND.n6485 GND.n6484 585
R10044 GND.n6479 GND.n1398 585
R10045 GND.n1398 GND.n1234 585
R10046 GND.n6478 GND.n6477 585
R10047 GND.n6477 GND.n1232 585
R10048 GND.n6476 GND.n1400 585
R10049 GND.n6476 GND.n6475 585
R10050 GND.n1407 GND.n1406 585
R10051 GND.n1407 GND.n1242 585
R10052 GND.n1405 GND.n1401 585
R10053 GND.n1401 GND.n1240 585
R10054 GND.n1404 GND.n1403 585
R10055 GND.n1403 GND.n1250 585
R10056 GND.n1402 GND.n1378 585
R10057 GND.n1378 GND.n1248 585
R10058 GND.n6500 GND.n1377 585
R10059 GND.n6500 GND.n6499 585
R10060 GND.n6502 GND.n6501 585
R10061 GND.n6501 GND.n1258 585
R10062 GND.n6503 GND.n1374 585
R10063 GND.n1374 GND.n1256 585
R10064 GND.n6505 GND.n6504 585
R10065 GND.n6506 GND.n6505 585
R10066 GND.n1376 GND.n1373 585
R10067 GND.n1373 GND.n1266 585
R10068 GND.n1375 GND.n1364 585
R10069 GND.n1364 GND.n1264 585
R10070 GND.n6514 GND.n1363 585
R10071 GND.n6514 GND.n6513 585
R10072 GND.n6516 GND.n6515 585
R10073 GND.n6515 GND.n1274 585
R10074 GND.n6517 GND.n1360 585
R10075 GND.n1360 GND.n1272 585
R10076 GND.n6519 GND.n6518 585
R10077 GND.n6520 GND.n6519 585
R10078 GND.n1362 GND.n1359 585
R10079 GND.n1359 GND.n1282 585
R10080 GND.n1361 GND.n1350 585
R10081 GND.n1350 GND.n1280 585
R10082 GND.n6528 GND.n1349 585
R10083 GND.n6528 GND.n6527 585
R10084 GND.n6530 GND.n6529 585
R10085 GND.n6529 GND.n1290 585
R10086 GND.n6531 GND.n1346 585
R10087 GND.n1346 GND.n1288 585
R10088 GND.n6533 GND.n6532 585
R10089 GND.n6534 GND.n6533 585
R10090 GND.n1348 GND.n1345 585
R10091 GND.n1345 GND.n1298 585
R10092 GND.n1347 GND.n1338 585
R10093 GND.n1338 GND.n1296 585
R10094 GND.n6542 GND.n1337 585
R10095 GND.n6542 GND.n6541 585
R10096 GND.n6544 GND.n6543 585
R10097 GND.n6543 GND.n1306 585
R10098 GND.n6545 GND.n1336 585
R10099 GND.n1336 GND.n1304 585
R10100 GND.n6547 GND.n6546 585
R10101 GND.n6548 GND.n6547 585
R10102 GND.n1328 GND.n1327 585
R10103 GND.n1328 GND.n1313 585
R10104 GND.n6556 GND.n6555 585
R10105 GND.n6555 GND.n6554 585
R10106 GND.n6557 GND.n1325 585
R10107 GND.n1325 GND.n1323 585
R10108 GND.n6559 GND.n6558 585
R10109 GND.n6560 GND.n6559 585
R10110 GND.n1326 GND.n1324 585
R10111 GND.n1324 GND.n1319 585
R10112 GND.n6244 GND.n6243 585
R10113 GND.n6244 GND.n1422 585
R10114 GND.n6257 GND.n6242 585
R10115 GND.n6257 GND.n6256 585
R10116 GND.n6259 GND.n6258 585
R10117 GND.n6258 GND.n1430 585
R10118 GND.n6260 GND.n6239 585
R10119 GND.n6239 GND.n1428 585
R10120 GND.n6262 GND.n6261 585
R10121 GND.n6263 GND.n6262 585
R10122 GND.n6241 GND.n6238 585
R10123 GND.n6238 GND.n1439 585
R10124 GND.n6240 GND.n6198 585
R10125 GND.n6198 GND.n1437 585
R10126 GND.n6271 GND.n6197 585
R10127 GND.n6271 GND.n6270 585
R10128 GND.n6273 GND.n6272 585
R10129 GND.n6272 GND.n1447 585
R10130 GND.n6274 GND.n6194 585
R10131 GND.n6194 GND.n1445 585
R10132 GND.n6276 GND.n6275 585
R10133 GND.n6277 GND.n6276 585
R10134 GND.n6196 GND.n6193 585
R10135 GND.n6193 GND.n1455 585
R10136 GND.n6195 GND.n6184 585
R10137 GND.n6184 GND.n1453 585
R10138 GND.n6285 GND.n6183 585
R10139 GND.n6285 GND.n6284 585
R10140 GND.n6287 GND.n6286 585
R10141 GND.n6286 GND.n1463 585
R10142 GND.n6288 GND.n6180 585
R10143 GND.n6180 GND.n1461 585
R10144 GND.n6290 GND.n6289 585
R10145 GND.n6291 GND.n6290 585
R10146 GND.n6182 GND.n6179 585
R10147 GND.n6179 GND.n1471 585
R10148 GND.n6181 GND.n1524 585
R10149 GND.n1524 GND.n1469 585
R10150 GND.n6299 GND.n1523 585
R10151 GND.n6299 GND.n6298 585
R10152 GND.n6301 GND.n6300 585
R10153 GND.n6300 GND.n1479 585
R10154 GND.n6302 GND.n1520 585
R10155 GND.n1520 GND.n1477 585
R10156 GND.n6304 GND.n6303 585
R10157 GND.n6305 GND.n6304 585
R10158 GND.n1522 GND.n1519 585
R10159 GND.n1519 GND.n1487 585
R10160 GND.n1521 GND.n1510 585
R10161 GND.n1510 GND.n1485 585
R10162 GND.n6314 GND.n1511 585
R10163 GND.n6314 GND.n6313 585
R10164 GND.n6315 GND.n1509 585
R10165 GND.n6315 GND.n1495 585
R10166 GND.n6317 GND.n6316 585
R10167 GND.n6316 GND.n1493 585
R10168 GND.n6318 GND.n1507 585
R10169 GND.n1507 GND.n1505 585
R10170 GND.n6320 GND.n6319 585
R10171 GND.n6321 GND.n6320 585
R10172 GND.n1508 GND.n1506 585
R10173 GND.n1506 GND.n1501 585
R10174 GND.n6156 GND.n6155 585
R10175 GND.n6157 GND.n6156 585
R10176 GND.n6154 GND.n1532 585
R10177 GND.n1532 GND.n1530 585
R10178 GND.n6153 GND.n6152 585
R10179 GND.n6152 GND.n6151 585
R10180 GND.n1534 GND.n1533 585
R10181 GND.n5583 GND.n1534 585
R10182 GND.n5574 GND.n5573 585
R10183 GND.n5573 GND.n1546 585
R10184 GND.n5576 GND.n5575 585
R10185 GND.n5576 GND.n1544 585
R10186 GND.n5625 GND.n5572 585
R10187 GND.n5625 GND.n5624 585
R10188 GND.n5627 GND.n5626 585
R10189 GND.n5626 GND.n1555 585
R10190 GND.n5628 GND.n5571 585
R10191 GND.n5571 GND.n1553 585
R10192 GND.n5630 GND.n5629 585
R10193 GND.n5631 GND.n5630 585
R10194 GND.n5199 GND.n5198 585
R10195 GND.n5199 GND.n1562 585
R10196 GND.n5639 GND.n5638 585
R10197 GND.n5638 GND.n5637 585
R10198 GND.n5640 GND.n5197 585
R10199 GND.n5201 GND.n5197 585
R10200 GND.n5642 GND.n5641 585
R10201 GND.n5642 GND.n1569 585
R10202 GND.n5643 GND.n5196 585
R10203 GND.n5643 GND.n1567 585
R10204 GND.n5645 GND.n5644 585
R10205 GND.n5644 GND.n1585 585
R10206 GND.n5646 GND.n5195 585
R10207 GND.n5195 GND.n1575 585
R10208 GND.n5648 GND.n5647 585
R10209 GND.n5649 GND.n5648 585
R10210 GND.n5190 GND.n5189 585
R10211 GND.n5651 GND.n5190 585
R10212 GND.n5659 GND.n5658 585
R10213 GND.n5658 GND.n5657 585
R10214 GND.n5660 GND.n5187 585
R10215 GND.n5191 GND.n5187 585
R10216 GND.n5662 GND.n5661 585
R10217 GND.n5663 GND.n5662 585
R10218 GND.n5188 GND.n5186 585
R10219 GND.n5186 GND.n5183 585
R10220 GND.n5551 GND.n5550 585
R10221 GND.n5552 GND.n5551 585
R10222 GND.n5172 GND.n5171 585
R10223 GND.n5175 GND.n5172 585
R10224 GND.n5673 GND.n5672 585
R10225 GND.n5672 GND.n5671 585
R10226 GND.n5674 GND.n5169 585
R10227 GND.n5173 GND.n5169 585
R10228 GND.n5676 GND.n5675 585
R10229 GND.n5677 GND.n5676 585
R10230 GND.n5170 GND.n5168 585
R10231 GND.n5168 GND.n5165 585
R10232 GND.n5538 GND.n5537 585
R10233 GND.n5539 GND.n5538 585
R10234 GND.n5153 GND.n5152 585
R10235 GND.n5157 GND.n5153 585
R10236 GND.n5687 GND.n5686 585
R10237 GND.n5686 GND.n5685 585
R10238 GND.n5688 GND.n5150 585
R10239 GND.n5155 GND.n5150 585
R10240 GND.n5690 GND.n5689 585
R10241 GND.n5691 GND.n5690 585
R10242 GND.n5151 GND.n5149 585
R10243 GND.n5149 GND.n5147 585
R10244 GND.n5525 GND.n5524 585
R10245 GND.n5526 GND.n5525 585
R10246 GND.n5523 GND.n5522 585
R10247 GND.n5522 GND.n5136 585
R10248 GND.n5132 GND.n5131 585
R10249 GND.n5699 GND.n5132 585
R10250 GND.n5702 GND.n5701 585
R10251 GND.n5701 GND.n5700 585
R10252 GND.n5703 GND.n5129 585
R10253 GND.n5514 GND.n5129 585
R10254 GND.n5705 GND.n5704 585
R10255 GND.n5706 GND.n5705 585
R10256 GND.n5130 GND.n5128 585
R10257 GND.n5128 GND.n5125 585
R10258 GND.n5508 GND.n5507 585
R10259 GND.n5509 GND.n5508 585
R10260 GND.n5114 GND.n5113 585
R10261 GND.n5117 GND.n5114 585
R10262 GND.n5716 GND.n5715 585
R10263 GND.n5715 GND.n5714 585
R10264 GND.n5717 GND.n5111 585
R10265 GND.n5115 GND.n5111 585
R10266 GND.n5719 GND.n5718 585
R10267 GND.n5720 GND.n5719 585
R10268 GND.n5112 GND.n5110 585
R10269 GND.n5110 GND.n5107 585
R10270 GND.n5495 GND.n5494 585
R10271 GND.n5496 GND.n5495 585
R10272 GND.n5096 GND.n5095 585
R10273 GND.n5099 GND.n5096 585
R10274 GND.n5730 GND.n5729 585
R10275 GND.n5729 GND.n5728 585
R10276 GND.n5731 GND.n5093 585
R10277 GND.n5097 GND.n5093 585
R10278 GND.n5733 GND.n5732 585
R10279 GND.n5734 GND.n5733 585
R10280 GND.n5094 GND.n5092 585
R10281 GND.n5092 GND.n5089 585
R10282 GND.n5482 GND.n5481 585
R10283 GND.n5483 GND.n5482 585
R10284 GND.n5079 GND.n5078 585
R10285 GND.n5479 GND.n5079 585
R10286 GND.n5744 GND.n5743 585
R10287 GND.n5743 GND.n5742 585
R10288 GND.n5745 GND.n5076 585
R10289 GND.n5080 GND.n5076 585
R10290 GND.n5747 GND.n5746 585
R10291 GND.n5748 GND.n5747 585
R10292 GND.n5077 GND.n5075 585
R10293 GND.n5075 GND.n5072 585
R10294 GND.n5468 GND.n5467 585
R10295 GND.n5469 GND.n5468 585
R10296 GND.n5466 GND.n5465 585
R10297 GND.n5465 GND.n5061 585
R10298 GND.n5057 GND.n5056 585
R10299 GND.n5756 GND.n5057 585
R10300 GND.n5759 GND.n5758 585
R10301 GND.n5758 GND.n5757 585
R10302 GND.n5760 GND.n5054 585
R10303 GND.n5457 GND.n5054 585
R10304 GND.n5762 GND.n5761 585
R10305 GND.n5763 GND.n5762 585
R10306 GND.n5055 GND.n5053 585
R10307 GND.n5053 GND.n5050 585
R10308 GND.n5451 GND.n5450 585
R10309 GND.n5452 GND.n5451 585
R10310 GND.n5039 GND.n5038 585
R10311 GND.n5042 GND.n5039 585
R10312 GND.n5773 GND.n5772 585
R10313 GND.n5772 GND.n5771 585
R10314 GND.n5774 GND.n5036 585
R10315 GND.n5040 GND.n5036 585
R10316 GND.n5776 GND.n5775 585
R10317 GND.n5777 GND.n5776 585
R10318 GND.n5037 GND.n5035 585
R10319 GND.n5035 GND.n5032 585
R10320 GND.n5438 GND.n5437 585
R10321 GND.n5439 GND.n5438 585
R10322 GND.n5021 GND.n5020 585
R10323 GND.n5024 GND.n5021 585
R10324 GND.n5787 GND.n5786 585
R10325 GND.n5786 GND.n5785 585
R10326 GND.n5788 GND.n5018 585
R10327 GND.n5022 GND.n5018 585
R10328 GND.n5790 GND.n5789 585
R10329 GND.n5791 GND.n5790 585
R10330 GND.n5019 GND.n5017 585
R10331 GND.n5017 GND.n5014 585
R10332 GND.n5425 GND.n5424 585
R10333 GND.n5426 GND.n5425 585
R10334 GND.n5004 GND.n5003 585
R10335 GND.n5006 GND.n5004 585
R10336 GND.n5801 GND.n5800 585
R10337 GND.n5800 GND.n5799 585
R10338 GND.n5802 GND.n5001 585
R10339 GND.n5417 GND.n5001 585
R10340 GND.n5804 GND.n5803 585
R10341 GND.n5805 GND.n5804 585
R10342 GND.n5002 GND.n5000 585
R10343 GND.n5000 GND.n4997 585
R10344 GND.n5411 GND.n5410 585
R10345 GND.n5412 GND.n5411 585
R10346 GND.n4986 GND.n4985 585
R10347 GND.n4989 GND.n4986 585
R10348 GND.n5815 GND.n5814 585
R10349 GND.n5814 GND.n5813 585
R10350 GND.n5816 GND.n4983 585
R10351 GND.n4987 GND.n4983 585
R10352 GND.n5818 GND.n5817 585
R10353 GND.n5819 GND.n5818 585
R10354 GND.n4984 GND.n4982 585
R10355 GND.n4982 GND.n4979 585
R10356 GND.n5398 GND.n5397 585
R10357 GND.n5399 GND.n5398 585
R10358 GND.n4968 GND.n4967 585
R10359 GND.n4971 GND.n4968 585
R10360 GND.n5829 GND.n5828 585
R10361 GND.n5828 GND.n5827 585
R10362 GND.n5830 GND.n4965 585
R10363 GND.n5390 GND.n4965 585
R10364 GND.n5832 GND.n5831 585
R10365 GND.n5833 GND.n5832 585
R10366 GND.n4966 GND.n4964 585
R10367 GND.n4964 GND.n4962 585
R10368 GND.n5278 GND.n5277 585
R10369 GND.n5280 GND.n5245 585
R10370 GND.n5281 GND.n5244 585
R10371 GND.n5281 GND.n4953 585
R10372 GND.n5284 GND.n5283 585
R10373 GND.n5285 GND.n5243 585
R10374 GND.n5287 GND.n5286 585
R10375 GND.n5289 GND.n5242 585
R10376 GND.n5292 GND.n5291 585
R10377 GND.n5293 GND.n5241 585
R10378 GND.n5295 GND.n5294 585
R10379 GND.n5297 GND.n5240 585
R10380 GND.n5300 GND.n5299 585
R10381 GND.n5301 GND.n5239 585
R10382 GND.n5303 GND.n5302 585
R10383 GND.n5305 GND.n5238 585
R10384 GND.n5308 GND.n5307 585
R10385 GND.n5309 GND.n5237 585
R10386 GND.n5311 GND.n5310 585
R10387 GND.n5313 GND.n5236 585
R10388 GND.n5316 GND.n5315 585
R10389 GND.n5317 GND.n5235 585
R10390 GND.n5322 GND.n5321 585
R10391 GND.n5324 GND.n5234 585
R10392 GND.n5327 GND.n5326 585
R10393 GND.n5328 GND.n5233 585
R10394 GND.n5330 GND.n5329 585
R10395 GND.n5334 GND.n5231 585
R10396 GND.n5337 GND.n5336 585
R10397 GND.n5338 GND.n5230 585
R10398 GND.n5343 GND.n5342 585
R10399 GND.n5345 GND.n5229 585
R10400 GND.n5348 GND.n5347 585
R10401 GND.n5349 GND.n5228 585
R10402 GND.n5351 GND.n5350 585
R10403 GND.n5353 GND.n5227 585
R10404 GND.n5356 GND.n5355 585
R10405 GND.n5357 GND.n5226 585
R10406 GND.n5359 GND.n5358 585
R10407 GND.n5361 GND.n5225 585
R10408 GND.n5364 GND.n5363 585
R10409 GND.n5365 GND.n5224 585
R10410 GND.n5367 GND.n5366 585
R10411 GND.n5369 GND.n5223 585
R10412 GND.n5372 GND.n5371 585
R10413 GND.n5373 GND.n5222 585
R10414 GND.n5375 GND.n5374 585
R10415 GND.n5377 GND.n5221 585
R10416 GND.n5380 GND.n5379 585
R10417 GND.n5381 GND.n5220 585
R10418 GND.n5383 GND.n5382 585
R10419 GND.n5385 GND.n5219 585
R10420 GND.n5386 GND.n5218 585
R10421 GND.n5386 GND.n4953 585
R10422 GND.n7424 GND.n7423 585
R10423 GND.n7422 GND.n7421 585
R10424 GND.n7420 GND.n7419 585
R10425 GND.n7418 GND.n7417 585
R10426 GND.n7416 GND.n7415 585
R10427 GND.n7414 GND.n7413 585
R10428 GND.n7412 GND.n7411 585
R10429 GND.n7410 GND.n7409 585
R10430 GND.n7408 GND.n7407 585
R10431 GND.n7406 GND.n7405 585
R10432 GND.n7404 GND.n7403 585
R10433 GND.n7402 GND.n7401 585
R10434 GND.n7400 GND.n7399 585
R10435 GND.n7398 GND.n7397 585
R10436 GND.n7396 GND.n7395 585
R10437 GND.n7394 GND.n7393 585
R10438 GND.n7392 GND.n7391 585
R10439 GND.n7390 GND.n7389 585
R10440 GND.n7388 GND.n7387 585
R10441 GND.n7386 GND.n7385 585
R10442 GND.n7384 GND.n7383 585
R10443 GND.n7382 GND.n7381 585
R10444 GND.n7380 GND.n7379 585
R10445 GND.n7378 GND.n7377 585
R10446 GND.n7376 GND.n7375 585
R10447 GND.n738 GND.n735 585
R10448 GND.n7594 GND.n7593 585
R10449 GND.n7542 GND.n736 585
R10450 GND.n7544 GND.n7543 585
R10451 GND.n7546 GND.n7545 585
R10452 GND.n7548 GND.n7547 585
R10453 GND.n7551 GND.n7550 585
R10454 GND.n7553 GND.n7552 585
R10455 GND.n7555 GND.n7554 585
R10456 GND.n7557 GND.n7556 585
R10457 GND.n7559 GND.n7558 585
R10458 GND.n7561 GND.n7560 585
R10459 GND.n7563 GND.n7562 585
R10460 GND.n7565 GND.n7564 585
R10461 GND.n7567 GND.n7566 585
R10462 GND.n7569 GND.n7568 585
R10463 GND.n7571 GND.n7570 585
R10464 GND.n7573 GND.n7572 585
R10465 GND.n7575 GND.n7574 585
R10466 GND.n7577 GND.n7576 585
R10467 GND.n7579 GND.n7578 585
R10468 GND.n7581 GND.n7580 585
R10469 GND.n7583 GND.n7582 585
R10470 GND.n7585 GND.n7584 585
R10471 GND.n7587 GND.n7586 585
R10472 GND.n7589 GND.n7588 585
R10473 GND.n7590 GND.n766 585
R10474 GND.n7592 GND.n7591 585
R10475 GND.n7593 GND.n7592 585
R10476 GND.n7427 GND.n7426 585
R10477 GND.n7426 GND.n7425 585
R10478 GND.n7428 GND.n799 585
R10479 GND.n7535 GND.n799 585
R10480 GND.n7430 GND.n7429 585
R10481 GND.n7429 GND.n798 585
R10482 GND.n7431 GND.n807 585
R10483 GND.n7441 GND.n807 585
R10484 GND.n7432 GND.n814 585
R10485 GND.n814 GND.n806 585
R10486 GND.n7434 GND.n7433 585
R10487 GND.n7435 GND.n7434 585
R10488 GND.n7371 GND.n813 585
R10489 GND.n817 GND.n813 585
R10490 GND.n7370 GND.n7369 585
R10491 GND.n7369 GND.n7368 585
R10492 GND.n816 GND.n815 585
R10493 GND.n7361 GND.n816 585
R10494 GND.n7347 GND.n823 585
R10495 GND.n7362 GND.n823 585
R10496 GND.n7349 GND.n7348 585
R10497 GND.t36 GND.n7349 585
R10498 GND.n7346 GND.n831 585
R10499 GND.n831 GND.n830 585
R10500 GND.n7345 GND.n7344 585
R10501 GND.n7344 GND.n7343 585
R10502 GND.n833 GND.n832 585
R10503 GND.n840 GND.n833 585
R10504 GND.n7312 GND.n839 585
R10505 GND.n7336 GND.n839 585
R10506 GND.n7315 GND.n7314 585
R10507 GND.n7314 GND.n7313 585
R10508 GND.n7316 GND.n847 585
R10509 GND.n7326 GND.n847 585
R10510 GND.n7317 GND.n854 585
R10511 GND.n854 GND.n846 585
R10512 GND.n7319 GND.n7318 585
R10513 GND.n7320 GND.n7319 585
R10514 GND.n7311 GND.n853 585
R10515 GND.n858 GND.n853 585
R10516 GND.n7310 GND.n7309 585
R10517 GND.n7309 GND.n7308 585
R10518 GND.n856 GND.n855 585
R10519 GND.n857 GND.n856 585
R10520 GND.n7276 GND.n864 585
R10521 GND.n7302 GND.n864 585
R10522 GND.n7278 GND.n7277 585
R10523 GND.n7277 GND.n873 585
R10524 GND.n7279 GND.n872 585
R10525 GND.n7290 GND.n872 585
R10526 GND.n7280 GND.n879 585
R10527 GND.n879 GND.n871 585
R10528 GND.n7282 GND.n7281 585
R10529 GND.n7284 GND.n7282 585
R10530 GND.n7275 GND.n878 585
R10531 GND.n878 GND.n877 585
R10532 GND.n7274 GND.n7273 585
R10533 GND.n7273 GND.n7272 585
R10534 GND.n881 GND.n880 585
R10535 GND.n7265 GND.n881 585
R10536 GND.n7264 GND.n7263 585
R10537 GND.n7266 GND.n7264 585
R10538 GND.n7262 GND.n888 585
R10539 GND.n892 GND.n888 585
R10540 GND.n7261 GND.n7260 585
R10541 GND.n7260 GND.n7259 585
R10542 GND.n890 GND.n889 585
R10543 GND.n7252 GND.n890 585
R10544 GND.n7251 GND.n7250 585
R10545 GND.n7253 GND.n7251 585
R10546 GND.n7249 GND.n898 585
R10547 GND.n902 GND.n898 585
R10548 GND.n7248 GND.n7247 585
R10549 GND.n7247 GND.n7246 585
R10550 GND.n900 GND.n899 585
R10551 GND.n901 GND.n900 585
R10552 GND.n7196 GND.n908 585
R10553 GND.n7240 GND.n908 585
R10554 GND.n7198 GND.n7197 585
R10555 GND.n7197 GND.n916 585
R10556 GND.n7199 GND.n915 585
R10557 GND.n7210 GND.n915 585
R10558 GND.n7201 GND.n7200 585
R10559 GND.n7202 GND.n7201 585
R10560 GND.n7195 GND.n921 585
R10561 GND.n7204 GND.n921 585
R10562 GND.n7194 GND.n7193 585
R10563 GND.n7193 GND.n920 585
R10564 GND.n7192 GND.n922 585
R10565 GND.n7192 GND.n7191 585
R10566 GND.n7181 GND.n923 585
R10567 GND.n7184 GND.n923 585
R10568 GND.n7183 GND.n7182 585
R10569 GND.n7185 GND.n7183 585
R10570 GND.n7180 GND.n930 585
R10571 GND.n934 GND.n930 585
R10572 GND.n7179 GND.n7178 585
R10573 GND.n7178 GND.n7177 585
R10574 GND.n932 GND.n931 585
R10575 GND.n933 GND.n932 585
R10576 GND.n7136 GND.n940 585
R10577 GND.n7171 GND.n940 585
R10578 GND.n7138 GND.n7137 585
R10579 GND.n7137 GND.n949 585
R10580 GND.n7139 GND.n948 585
R10581 GND.n7150 GND.n948 585
R10582 GND.n7140 GND.n955 585
R10583 GND.n955 GND.n947 585
R10584 GND.n7142 GND.n7141 585
R10585 GND.n7144 GND.n7142 585
R10586 GND.n7135 GND.n954 585
R10587 GND.n954 GND.n953 585
R10588 GND.n7134 GND.n7133 585
R10589 GND.n7133 GND.n7132 585
R10590 GND.n957 GND.n956 585
R10591 GND.n965 GND.n957 585
R10592 GND.n7098 GND.n964 585
R10593 GND.n7126 GND.n964 585
R10594 GND.n7100 GND.n7099 585
R10595 GND.n7099 GND.n963 585
R10596 GND.n7101 GND.n973 585
R10597 GND.n7111 GND.n973 585
R10598 GND.n7102 GND.n980 585
R10599 GND.n980 GND.n972 585
R10600 GND.n7104 GND.n7103 585
R10601 GND.n7105 GND.n7104 585
R10602 GND.n7097 GND.n979 585
R10603 GND.n984 GND.n979 585
R10604 GND.n7096 GND.n7095 585
R10605 GND.n7095 GND.n7094 585
R10606 GND.n982 GND.n981 585
R10607 GND.n983 GND.n982 585
R10608 GND.n7062 GND.n990 585
R10609 GND.n7088 GND.n990 585
R10610 GND.n7064 GND.n7063 585
R10611 GND.n7063 GND.n999 585
R10612 GND.n7065 GND.n998 585
R10613 GND.n7076 GND.n998 585
R10614 GND.n7066 GND.n1005 585
R10615 GND.n1005 GND.n997 585
R10616 GND.n7068 GND.n7067 585
R10617 GND.n7070 GND.n7068 585
R10618 GND.n7061 GND.n1004 585
R10619 GND.n1004 GND.n1003 585
R10620 GND.n7060 GND.n7059 585
R10621 GND.n7059 GND.n7058 585
R10622 GND.n1007 GND.n1006 585
R10623 GND.n7051 GND.n1007 585
R10624 GND.n7050 GND.n7049 585
R10625 GND.n7052 GND.n7050 585
R10626 GND.n7048 GND.n1014 585
R10627 GND.n1018 GND.n1014 585
R10628 GND.n7047 GND.n7046 585
R10629 GND.n7046 GND.n7045 585
R10630 GND.n1016 GND.n1015 585
R10631 GND.n1017 GND.n1016 585
R10632 GND.n7004 GND.n1024 585
R10633 GND.n7039 GND.n1024 585
R10634 GND.n7006 GND.n7005 585
R10635 GND.n7005 GND.n1033 585
R10636 GND.n7007 GND.n1032 585
R10637 GND.n7018 GND.n1032 585
R10638 GND.n7009 GND.n7008 585
R10639 GND.n7010 GND.n7009 585
R10640 GND.n7003 GND.n1038 585
R10641 GND.n7012 GND.n1038 585
R10642 GND.n7002 GND.n7001 585
R10643 GND.n7001 GND.n7000 585
R10644 GND.n1040 GND.n1039 585
R10645 GND.n6999 GND.n1040 585
R10646 GND.n6749 GND.n6748 585
R10647 GND.n6748 GND.n6747 585
R10648 GND.n6750 GND.n1046 585
R10649 GND.n6993 GND.n1046 585
R10650 GND.n6752 GND.n6751 585
R10651 GND.n6752 GND.n1045 585
R10652 GND.n6753 GND.n6746 585
R10653 GND.n6753 GND.n1057 585
R10654 GND.n6755 GND.n6754 585
R10655 GND.n6754 GND.n1055 585
R10656 GND.n6756 GND.n1088 585
R10657 GND.n6904 GND.n1088 585
R10658 GND.n6758 GND.n6757 585
R10659 GND.n6757 GND.n1087 585
R10660 GND.n6759 GND.n1094 585
R10661 GND.n6895 GND.n1094 585
R10662 GND.n6761 GND.n6760 585
R10663 GND.n6761 GND.n1093 585
R10664 GND.n6763 GND.n6762 585
R10665 GND.n6762 GND.n1103 585
R10666 GND.n6764 GND.n6743 585
R10667 GND.n6743 GND.n1101 585
R10668 GND.n6766 GND.n6765 585
R10669 GND.n6767 GND.n6766 585
R10670 GND.n6745 GND.n6742 585
R10671 GND.n6742 GND.n1112 585
R10672 GND.n6744 GND.n6709 585
R10673 GND.n6709 GND.n1110 585
R10674 GND.n6775 GND.n6708 585
R10675 GND.n6775 GND.n6774 585
R10676 GND.n6777 GND.n6776 585
R10677 GND.n6776 GND.n1120 585
R10678 GND.n6778 GND.n1205 585
R10679 GND.n1205 GND.n1118 585
R10680 GND.n6780 GND.n6779 585
R10681 GND.n6781 GND.n6780 585
R10682 GND.n6707 GND.n1204 585
R10683 GND.n1204 GND.n1128 585
R10684 GND.n6706 GND.n6705 585
R10685 GND.n6705 GND.n1126 585
R10686 GND.n6704 GND.n1196 585
R10687 GND.n6788 GND.n1196 585
R10688 GND.n6703 GND.n6702 585
R10689 GND.n6702 GND.n1136 585
R10690 GND.n6701 GND.n6700 585
R10691 GND.n6701 GND.n1134 585
R10692 GND.n6699 GND.n1190 585
R10693 GND.n6795 GND.n1190 585
R10694 GND.n6698 GND.n6697 585
R10695 GND.n6697 GND.n1144 585
R10696 GND.n6696 GND.n6695 585
R10697 GND.n6696 GND.n1142 585
R10698 GND.n6694 GND.n1183 585
R10699 GND.n6802 GND.n1183 585
R10700 GND.n6693 GND.n6692 585
R10701 GND.n6692 GND.n1152 585
R10702 GND.n6691 GND.n6690 585
R10703 GND.n6691 GND.n1150 585
R10704 GND.n6689 GND.n1177 585
R10705 GND.n6810 GND.n1177 585
R10706 GND.n6688 GND.n6687 585
R10707 GND.n6687 GND.n1160 585
R10708 GND.n6686 GND.n1206 585
R10709 GND.n6686 GND.n1158 585
R10710 GND.n6685 GND.n6684 585
R10711 GND.n6685 GND.n1170 585
R10712 GND.n6683 GND.n1169 585
R10713 GND.n6818 GND.n1169 585
R10714 GND.n6682 GND.n6681 585
R10715 GND.n6681 GND.n1166 585
R10716 GND.n6680 GND.n1207 585
R10717 GND.n6680 GND.n6679 585
R10718 GND.n1388 GND.n1208 585
R10719 GND.n1209 GND.n1208 585
R10720 GND.n1389 GND.n1215 585
R10721 GND.n6673 GND.n1215 585
R10722 GND.n1392 GND.n1390 585
R10723 GND.n1392 GND.n1391 585
R10724 GND.n1394 GND.n1393 585
R10725 GND.n1393 GND.n1225 585
R10726 GND.n1395 GND.n1387 585
R10727 GND.n1387 GND.n1223 585
R10728 GND.n6486 GND.n1396 585
R10729 GND.n6486 GND.n6485 585
R10730 GND.n6487 GND.n1386 585
R10731 GND.n6487 GND.n1234 585
R10732 GND.n6489 GND.n6488 585
R10733 GND.n6488 GND.n1232 585
R10734 GND.n6490 GND.n1385 585
R10735 GND.n6475 GND.n1385 585
R10736 GND.n6492 GND.n6491 585
R10737 GND.n6492 GND.n1242 585
R10738 GND.n6493 GND.n1384 585
R10739 GND.n6493 GND.n1240 585
R10740 GND.n6495 GND.n6494 585
R10741 GND.n6494 GND.n1250 585
R10742 GND.n6496 GND.n1381 585
R10743 GND.n1381 GND.n1248 585
R10744 GND.n6498 GND.n6497 585
R10745 GND.n6499 GND.n6498 585
R10746 GND.n1383 GND.n1380 585
R10747 GND.n1380 GND.n1258 585
R10748 GND.n1382 GND.n1371 585
R10749 GND.n1371 GND.n1256 585
R10750 GND.n6507 GND.n1370 585
R10751 GND.n6507 GND.n6506 585
R10752 GND.n6509 GND.n6508 585
R10753 GND.n6508 GND.n1266 585
R10754 GND.n6510 GND.n1367 585
R10755 GND.n1367 GND.n1264 585
R10756 GND.n6512 GND.n6511 585
R10757 GND.n6513 GND.n6512 585
R10758 GND.n1369 GND.n1366 585
R10759 GND.n1366 GND.n1274 585
R10760 GND.n1368 GND.n1357 585
R10761 GND.n1357 GND.n1272 585
R10762 GND.n6521 GND.n1356 585
R10763 GND.n6521 GND.n6520 585
R10764 GND.n6523 GND.n6522 585
R10765 GND.n6522 GND.n1282 585
R10766 GND.n6524 GND.n1353 585
R10767 GND.n1353 GND.n1280 585
R10768 GND.n6526 GND.n6525 585
R10769 GND.n6527 GND.n6526 585
R10770 GND.n1355 GND.n1352 585
R10771 GND.n1352 GND.n1290 585
R10772 GND.n1354 GND.n1344 585
R10773 GND.n1344 GND.n1288 585
R10774 GND.n6535 GND.n1343 585
R10775 GND.n6535 GND.n6534 585
R10776 GND.n6537 GND.n6536 585
R10777 GND.n6536 GND.n1298 585
R10778 GND.n6538 GND.n1341 585
R10779 GND.n1341 GND.n1296 585
R10780 GND.n6540 GND.n6539 585
R10781 GND.n6541 GND.n6540 585
R10782 GND.n1342 GND.n1340 585
R10783 GND.n1340 GND.n1306 585
R10784 GND.n1334 GND.n1333 585
R10785 GND.n1334 GND.n1304 585
R10786 GND.n6550 GND.n6549 585
R10787 GND.n6549 GND.n6548 585
R10788 GND.n6551 GND.n1331 585
R10789 GND.n1331 GND.n1313 585
R10790 GND.n6553 GND.n6552 585
R10791 GND.n6554 GND.n6553 585
R10792 GND.n1332 GND.n1330 585
R10793 GND.n1330 GND.n1323 585
R10794 GND.n6250 GND.n1322 585
R10795 GND.n6560 GND.n1322 585
R10796 GND.n6252 GND.n6251 585
R10797 GND.n6251 GND.n1319 585
R10798 GND.n6253 GND.n6247 585
R10799 GND.n6247 GND.n1422 585
R10800 GND.n6255 GND.n6254 585
R10801 GND.n6256 GND.n6255 585
R10802 GND.n6249 GND.n6246 585
R10803 GND.n6246 GND.n1430 585
R10804 GND.n6248 GND.n6205 585
R10805 GND.n6205 GND.n1428 585
R10806 GND.n6264 GND.n6204 585
R10807 GND.n6264 GND.n6263 585
R10808 GND.n6266 GND.n6265 585
R10809 GND.n6265 GND.n1439 585
R10810 GND.n6267 GND.n6201 585
R10811 GND.n6201 GND.n1437 585
R10812 GND.n6269 GND.n6268 585
R10813 GND.n6270 GND.n6269 585
R10814 GND.n6203 GND.n6200 585
R10815 GND.n6200 GND.n1447 585
R10816 GND.n6202 GND.n6191 585
R10817 GND.n6191 GND.n1445 585
R10818 GND.n6278 GND.n6190 585
R10819 GND.n6278 GND.n6277 585
R10820 GND.n6280 GND.n6279 585
R10821 GND.n6279 GND.n1455 585
R10822 GND.n6281 GND.n6187 585
R10823 GND.n6187 GND.n1453 585
R10824 GND.n6283 GND.n6282 585
R10825 GND.n6284 GND.n6283 585
R10826 GND.n6189 GND.n6186 585
R10827 GND.n6186 GND.n1463 585
R10828 GND.n6188 GND.n6177 585
R10829 GND.n6177 GND.n1461 585
R10830 GND.n6292 GND.n6176 585
R10831 GND.n6292 GND.n6291 585
R10832 GND.n6294 GND.n6293 585
R10833 GND.n6293 GND.n1471 585
R10834 GND.n6295 GND.n1526 585
R10835 GND.n1526 GND.n1469 585
R10836 GND.n6297 GND.n6296 585
R10837 GND.n6298 GND.n6297 585
R10838 GND.n6175 GND.n1525 585
R10839 GND.n1525 GND.n1479 585
R10840 GND.n6174 GND.n6173 585
R10841 GND.n6173 GND.n1477 585
R10842 GND.n6172 GND.n1518 585
R10843 GND.n6305 GND.n1518 585
R10844 GND.n6171 GND.n6170 585
R10845 GND.n6170 GND.n1487 585
R10846 GND.n6169 GND.n6168 585
R10847 GND.n6169 GND.n1485 585
R10848 GND.n6167 GND.n1512 585
R10849 GND.n6313 GND.n1512 585
R10850 GND.n6166 GND.n6165 585
R10851 GND.n6165 GND.n1495 585
R10852 GND.n6164 GND.n1527 585
R10853 GND.n6164 GND.n1493 585
R10854 GND.n6163 GND.n6162 585
R10855 GND.n6163 GND.n1505 585
R10856 GND.n6161 GND.n1504 585
R10857 GND.n6321 GND.n1504 585
R10858 GND.n6160 GND.n6159 585
R10859 GND.n6159 GND.n1501 585
R10860 GND.n6158 GND.n1528 585
R10861 GND.n6158 GND.n6157 585
R10862 GND.n5580 GND.n1529 585
R10863 GND.n1530 GND.n1529 585
R10864 GND.n5581 GND.n1536 585
R10865 GND.n6151 GND.n1536 585
R10866 GND.n5584 GND.n5582 585
R10867 GND.n5584 GND.n5583 585
R10868 GND.n5586 GND.n5585 585
R10869 GND.n5585 GND.n1546 585
R10870 GND.n5587 GND.n5578 585
R10871 GND.n5578 GND.n1544 585
R10872 GND.n5589 GND.n5588 585
R10873 GND.n5624 GND.n5589 585
R10874 GND.n5579 GND.n5577 585
R10875 GND.n5577 GND.n1555 585
R10876 GND.n5570 GND.n5569 585
R10877 GND.n5570 GND.n1553 585
R10878 GND.n5633 GND.n5632 585
R10879 GND.n5632 GND.n5631 585
R10880 GND.n5634 GND.n5203 585
R10881 GND.n5203 GND.n1562 585
R10882 GND.n5636 GND.n5635 585
R10883 GND.n5637 GND.n5636 585
R10884 GND.n5568 GND.n5202 585
R10885 GND.n5202 GND.n5201 585
R10886 GND.n5567 GND.n5566 585
R10887 GND.n5566 GND.n1569 585
R10888 GND.n5565 GND.n5204 585
R10889 GND.n5565 GND.n1567 585
R10890 GND.n5564 GND.n5563 585
R10891 GND.n5564 GND.n1585 585
R10892 GND.n5562 GND.n5205 585
R10893 GND.n5205 GND.n1575 585
R10894 GND.n5561 GND.n5194 585
R10895 GND.n5649 GND.n5194 585
R10896 GND.n5560 GND.n5193 585
R10897 GND.n5651 GND.n5193 585
R10898 GND.n5559 GND.n5192 585
R10899 GND.n5657 GND.n5192 585
R10900 GND.n5558 GND.n5557 585
R10901 GND.n5557 GND.n5191 585
R10902 GND.n5556 GND.n5184 585
R10903 GND.n5663 GND.n5184 585
R10904 GND.n5555 GND.n5554 585
R10905 GND.n5554 GND.n5183 585
R10906 GND.n5553 GND.n5206 585
R10907 GND.n5553 GND.n5552 585
R10908 GND.n5548 GND.n5547 585
R10909 GND.n5548 GND.n5175 585
R10910 GND.n5546 GND.n5174 585
R10911 GND.n5671 GND.n5174 585
R10912 GND.n5545 GND.n5544 585
R10913 GND.n5544 GND.n5173 585
R10914 GND.n5543 GND.n5166 585
R10915 GND.n5677 GND.n5166 585
R10916 GND.n5542 GND.n5541 585
R10917 GND.n5541 GND.n5165 585
R10918 GND.n5540 GND.n5207 585
R10919 GND.n5540 GND.n5539 585
R10920 GND.n5535 GND.n5534 585
R10921 GND.n5535 GND.n5157 585
R10922 GND.n5533 GND.n5156 585
R10923 GND.n5685 GND.n5156 585
R10924 GND.n5532 GND.n5531 585
R10925 GND.n5531 GND.n5155 585
R10926 GND.n5530 GND.n5148 585
R10927 GND.n5691 GND.n5148 585
R10928 GND.n5529 GND.n5528 585
R10929 GND.n5528 GND.n5147 585
R10930 GND.n5527 GND.n5208 585
R10931 GND.n5527 GND.n5526 585
R10932 GND.n5520 GND.n5519 585
R10933 GND.n5520 GND.n5136 585
R10934 GND.n5518 GND.n5135 585
R10935 GND.n5699 GND.n5135 585
R10936 GND.n5517 GND.n5134 585
R10937 GND.n5700 GND.n5134 585
R10938 GND.n5516 GND.n5515 585
R10939 GND.n5515 GND.n5514 585
R10940 GND.n5513 GND.n5126 585
R10941 GND.n5706 GND.n5126 585
R10942 GND.n5512 GND.n5511 585
R10943 GND.n5511 GND.n5125 585
R10944 GND.n5510 GND.n5209 585
R10945 GND.n5510 GND.n5509 585
R10946 GND.n5505 GND.n5504 585
R10947 GND.n5505 GND.n5117 585
R10948 GND.n5503 GND.n5116 585
R10949 GND.n5714 GND.n5116 585
R10950 GND.n5502 GND.n5501 585
R10951 GND.n5501 GND.n5115 585
R10952 GND.n5500 GND.n5108 585
R10953 GND.n5720 GND.n5108 585
R10954 GND.n5499 GND.n5498 585
R10955 GND.n5498 GND.n5107 585
R10956 GND.n5497 GND.n5210 585
R10957 GND.n5497 GND.n5496 585
R10958 GND.n5492 GND.n5491 585
R10959 GND.n5492 GND.n5099 585
R10960 GND.n5490 GND.n5098 585
R10961 GND.n5728 GND.n5098 585
R10962 GND.n5489 GND.n5488 585
R10963 GND.n5488 GND.n5097 585
R10964 GND.n5487 GND.n5090 585
R10965 GND.n5734 GND.n5090 585
R10966 GND.n5486 GND.n5485 585
R10967 GND.n5485 GND.n5089 585
R10968 GND.n5484 GND.n5211 585
R10969 GND.n5484 GND.n5483 585
R10970 GND.n5478 GND.n5477 585
R10971 GND.n5479 GND.n5478 585
R10972 GND.n5476 GND.n5081 585
R10973 GND.n5742 GND.n5081 585
R10974 GND.n5475 GND.n5474 585
R10975 GND.n5474 GND.n5080 585
R10976 GND.n5473 GND.n5073 585
R10977 GND.n5748 GND.n5073 585
R10978 GND.n5472 GND.n5471 585
R10979 GND.n5471 GND.n5072 585
R10980 GND.n5470 GND.n5212 585
R10981 GND.n5470 GND.n5469 585
R10982 GND.n5463 GND.n5462 585
R10983 GND.n5463 GND.n5061 585
R10984 GND.n5461 GND.n5060 585
R10985 GND.n5756 GND.n5060 585
R10986 GND.n5460 GND.n5059 585
R10987 GND.n5757 GND.n5059 585
R10988 GND.n5459 GND.n5458 585
R10989 GND.n5458 GND.n5457 585
R10990 GND.n5456 GND.n5051 585
R10991 GND.n5763 GND.n5051 585
R10992 GND.n5455 GND.n5454 585
R10993 GND.n5454 GND.n5050 585
R10994 GND.n5453 GND.n5213 585
R10995 GND.n5453 GND.n5452 585
R10996 GND.n5448 GND.n5447 585
R10997 GND.n5448 GND.n5042 585
R10998 GND.n5446 GND.n5041 585
R10999 GND.n5771 GND.n5041 585
R11000 GND.n5445 GND.n5444 585
R11001 GND.n5444 GND.n5040 585
R11002 GND.n5443 GND.n5033 585
R11003 GND.n5777 GND.n5033 585
R11004 GND.n5442 GND.n5441 585
R11005 GND.n5441 GND.n5032 585
R11006 GND.n5440 GND.n5214 585
R11007 GND.n5440 GND.n5439 585
R11008 GND.n5435 GND.n5434 585
R11009 GND.n5435 GND.n5024 585
R11010 GND.n5433 GND.n5023 585
R11011 GND.n5785 GND.n5023 585
R11012 GND.n5432 GND.n5431 585
R11013 GND.n5431 GND.n5022 585
R11014 GND.n5430 GND.n5015 585
R11015 GND.n5791 GND.n5015 585
R11016 GND.n5429 GND.n5428 585
R11017 GND.n5428 GND.n5014 585
R11018 GND.n5427 GND.n5215 585
R11019 GND.n5427 GND.n5426 585
R11020 GND.n5422 GND.n5421 585
R11021 GND.n5422 GND.n5006 585
R11022 GND.n5420 GND.n5005 585
R11023 GND.n5799 GND.n5005 585
R11024 GND.n5419 GND.n5418 585
R11025 GND.n5418 GND.n5417 585
R11026 GND.n5416 GND.n4998 585
R11027 GND.n5805 GND.n4998 585
R11028 GND.n5415 GND.n5414 585
R11029 GND.n5414 GND.n4997 585
R11030 GND.n5413 GND.n5216 585
R11031 GND.n5413 GND.n5412 585
R11032 GND.n5408 GND.n5407 585
R11033 GND.n5408 GND.n4989 585
R11034 GND.n5406 GND.n4988 585
R11035 GND.n5813 GND.n4988 585
R11036 GND.n5405 GND.n5404 585
R11037 GND.n5404 GND.n4987 585
R11038 GND.n5403 GND.n4980 585
R11039 GND.n5819 GND.n4980 585
R11040 GND.n5402 GND.n5401 585
R11041 GND.n5401 GND.n4979 585
R11042 GND.n5400 GND.n5217 585
R11043 GND.n5400 GND.n5399 585
R11044 GND.n5395 GND.n5394 585
R11045 GND.n5395 GND.n4971 585
R11046 GND.n5393 GND.n4970 585
R11047 GND.n5827 GND.n4970 585
R11048 GND.n5392 GND.n5391 585
R11049 GND.n5391 GND.n5390 585
R11050 GND.n5389 GND.n4963 585
R11051 GND.n5833 GND.n4963 585
R11052 GND.n5388 GND.n5387 585
R11053 GND.n5387 GND.n4962 585
R11054 GND.n5902 GND.n1608 585
R11055 GND.n6046 GND.n1608 585
R11056 GND.n5901 GND.n5900 585
R11057 GND.n5900 GND.n5899 585
R11058 GND.n1675 GND.n1674 585
R11059 GND.n5869 GND.n1675 585
R11060 GND.n5889 GND.n5888 585
R11061 GND.n5890 GND.n5889 585
R11062 GND.n1687 GND.n1686 585
R11063 GND.n5864 GND.n1686 585
R11064 GND.n5883 GND.n5882 585
R11065 GND.n5882 GND.n5881 585
R11066 GND.n1690 GND.n1689 585
R11067 GND.n5861 GND.n1690 585
R11068 GND.n4928 GND.n4927 585
R11069 GND.n4929 GND.n4928 585
R11070 GND.n1714 GND.n1713 585
R11071 GND.n1713 GND.n1710 585
R11072 GND.n4923 GND.n4922 585
R11073 GND.n4922 GND.n4921 585
R11074 GND.n1717 GND.n1716 585
R11075 GND.n4912 GND.n1717 585
R11076 GND.n4890 GND.n1743 585
R11077 GND.n4872 GND.n1743 585
R11078 GND.n4892 GND.n4891 585
R11079 GND.n4893 GND.n4892 585
R11080 GND.n1744 GND.n1742 585
R11081 GND.n4869 GND.n1742 585
R11082 GND.n4885 GND.n4884 585
R11083 GND.n4884 GND.n4883 585
R11084 GND.n1747 GND.n1746 585
R11085 GND.n4866 GND.n1747 585
R11086 GND.n4853 GND.n1770 585
R11087 GND.n4835 GND.n1770 585
R11088 GND.n4855 GND.n4854 585
R11089 GND.n4856 GND.n4855 585
R11090 GND.n1771 GND.n1769 585
R11091 GND.n4832 GND.n1769 585
R11092 GND.n4848 GND.n4847 585
R11093 GND.n4847 GND.n4846 585
R11094 GND.n1774 GND.n1773 585
R11095 GND.n4798 GND.n1774 585
R11096 GND.n4785 GND.n1804 585
R11097 GND.n1804 GND.n1792 585
R11098 GND.n4787 GND.n4786 585
R11099 GND.n4788 GND.n4787 585
R11100 GND.n1805 GND.n1803 585
R11101 GND.n4763 GND.n1803 585
R11102 GND.n4780 GND.n4779 585
R11103 GND.n4779 GND.n4778 585
R11104 GND.n1808 GND.n1807 585
R11105 GND.n4760 GND.n1808 585
R11106 GND.n4747 GND.n1831 585
R11107 GND.n4729 GND.n1831 585
R11108 GND.n4749 GND.n4748 585
R11109 GND.n4750 GND.n4749 585
R11110 GND.n1832 GND.n1830 585
R11111 GND.n1847 GND.n1830 585
R11112 GND.n4742 GND.n4741 585
R11113 GND.n4741 GND.n4740 585
R11114 GND.n1835 GND.n1834 585
R11115 GND.n4704 GND.n1835 585
R11116 GND.n4691 GND.n1869 585
R11117 GND.n1869 GND.n1857 585
R11118 GND.n4693 GND.n4692 585
R11119 GND.n4694 GND.n4693 585
R11120 GND.n1870 GND.n1868 585
R11121 GND.n4660 GND.n1868 585
R11122 GND.n4656 GND.n4655 585
R11123 GND.n4657 GND.n4656 585
R11124 GND.n4654 GND.n4653 585
R11125 GND.n4653 GND.n4652 585
R11126 GND.n4638 GND.n1913 585
R11127 GND.n1923 GND.n1913 585
R11128 GND.n4640 GND.n4639 585
R11129 GND.n4641 GND.n4640 585
R11130 GND.n4637 GND.n1927 585
R11131 GND.n4637 GND.n4636 585
R11132 GND.n1926 GND.n1877 585
R11133 GND.n4633 GND.n1926 585
R11134 GND.n1881 GND.n1878 585
R11135 GND.n1931 GND.n1881 585
R11136 GND.n4687 GND.n4686 585
R11137 GND.n4686 GND.n4685 585
R11138 GND.n1880 GND.n1879 585
R11139 GND.n4624 GND.n1880 585
R11140 GND.n4620 GND.n4619 585
R11141 GND.n4621 GND.n4620 585
R11142 GND.n1943 GND.n1942 585
R11143 GND.n4597 GND.n1942 585
R11144 GND.n4615 GND.n4614 585
R11145 GND.n4614 GND.n4613 585
R11146 GND.n1946 GND.n1945 585
R11147 GND.n4605 GND.n1946 585
R11148 GND.n4588 GND.n1972 585
R11149 GND.n4570 GND.n1972 585
R11150 GND.n4590 GND.n4589 585
R11151 GND.n4591 GND.n4590 585
R11152 GND.n1973 GND.n1971 585
R11153 GND.n1988 GND.n1971 585
R11154 GND.n4583 GND.n4582 585
R11155 GND.n4582 GND.n4581 585
R11156 GND.n1976 GND.n1975 585
R11157 GND.n4481 GND.n1976 585
R11158 GND.n4513 GND.n4512 585
R11159 GND.n4514 GND.n4513 585
R11160 GND.n2007 GND.n2006 585
R11161 GND.n2006 GND.n2001 585
R11162 GND.n4508 GND.n4507 585
R11163 GND.n4507 GND.n4506 585
R11164 GND.n2010 GND.n2009 585
R11165 GND.n4494 GND.n2010 585
R11166 GND.n4470 GND.n2034 585
R11167 GND.n4452 GND.n2034 585
R11168 GND.n4472 GND.n4471 585
R11169 GND.n4473 GND.n4472 585
R11170 GND.n2035 GND.n2033 585
R11171 GND.n2050 GND.n2033 585
R11172 GND.n4465 GND.n4464 585
R11173 GND.n4464 GND.n4463 585
R11174 GND.n2038 GND.n2037 585
R11175 GND.n4399 GND.n2038 585
R11176 GND.n4431 GND.n4430 585
R11177 GND.n4432 GND.n4431 585
R11178 GND.n2069 GND.n2068 585
R11179 GND.n2068 GND.n2063 585
R11180 GND.n4426 GND.n4425 585
R11181 GND.n4425 GND.n4424 585
R11182 GND.n2072 GND.n2071 585
R11183 GND.n4412 GND.n2072 585
R11184 GND.n4388 GND.n2097 585
R11185 GND.n4370 GND.n2097 585
R11186 GND.n4390 GND.n4389 585
R11187 GND.n4391 GND.n4390 585
R11188 GND.n2098 GND.n2096 585
R11189 GND.n4367 GND.n2096 585
R11190 GND.n4383 GND.n4382 585
R11191 GND.n4382 GND.n4381 585
R11192 GND.n2101 GND.n2100 585
R11193 GND.n4364 GND.n2101 585
R11194 GND.n4352 GND.n2126 585
R11195 GND.n4334 GND.n2126 585
R11196 GND.n4354 GND.n4353 585
R11197 GND.n4355 GND.n4354 585
R11198 GND.n2127 GND.n2125 585
R11199 GND.n4331 GND.n2125 585
R11200 GND.n4347 GND.n4346 585
R11201 GND.n4346 GND.n4345 585
R11202 GND.n4158 GND.n2129 585
R11203 GND.n4311 GND.n4310 585
R11204 GND.n4309 GND.n4157 585
R11205 GND.n4313 GND.n4157 585
R11206 GND.n4308 GND.n4307 585
R11207 GND.n4306 GND.n4305 585
R11208 GND.n4304 GND.n4303 585
R11209 GND.n4302 GND.n4301 585
R11210 GND.n4300 GND.n4299 585
R11211 GND.n4298 GND.n4166 585
R11212 GND.n4297 GND.n4296 585
R11213 GND.n4295 GND.n4294 585
R11214 GND.n4293 GND.n4292 585
R11215 GND.n4291 GND.n4290 585
R11216 GND.n4289 GND.n4288 585
R11217 GND.n4287 GND.n4286 585
R11218 GND.n4285 GND.n4284 585
R11219 GND.n4283 GND.n4282 585
R11220 GND.n4281 GND.n4280 585
R11221 GND.n4278 GND.n4277 585
R11222 GND.n4276 GND.n4275 585
R11223 GND.n4274 GND.n4273 585
R11224 GND.n4272 GND.n4271 585
R11225 GND.n4270 GND.n4269 585
R11226 GND.n4268 GND.n4267 585
R11227 GND.n4266 GND.n4265 585
R11228 GND.n4264 GND.n4263 585
R11229 GND.n4262 GND.n4261 585
R11230 GND.n4260 GND.n4259 585
R11231 GND.n4258 GND.n4257 585
R11232 GND.n4256 GND.n4255 585
R11233 GND.n4254 GND.n4253 585
R11234 GND.n4252 GND.n4251 585
R11235 GND.n4250 GND.n4249 585
R11236 GND.n4248 GND.n4247 585
R11237 GND.n4246 GND.n4245 585
R11238 GND.n4244 GND.n4243 585
R11239 GND.n4242 GND.n4241 585
R11240 GND.n4240 GND.n4239 585
R11241 GND.n4238 GND.n4237 585
R11242 GND.n4236 GND.n4235 585
R11243 GND.n4234 GND.n4233 585
R11244 GND.n4232 GND.n4231 585
R11245 GND.n4230 GND.n4229 585
R11246 GND.n4228 GND.n4227 585
R11247 GND.n4226 GND.n4225 585
R11248 GND.n4224 GND.n4223 585
R11249 GND.n4222 GND.n4221 585
R11250 GND.n4220 GND.n4219 585
R11251 GND.n4215 GND.n4214 585
R11252 GND.n6002 GND.n1606 585
R11253 GND.n6003 GND.n6001 585
R11254 GND.n6004 GND.n5998 585
R11255 GND.n5996 GND.n5995 585
R11256 GND.n6008 GND.n5994 585
R11257 GND.n6009 GND.n5993 585
R11258 GND.n6010 GND.n5992 585
R11259 GND.n5990 GND.n5989 585
R11260 GND.n6014 GND.n5988 585
R11261 GND.n6015 GND.n5987 585
R11262 GND.n6016 GND.n5986 585
R11263 GND.n5984 GND.n5983 585
R11264 GND.n6020 GND.n5980 585
R11265 GND.n6021 GND.n5979 585
R11266 GND.n6022 GND.n5978 585
R11267 GND.n5976 GND.n5975 585
R11268 GND.n6026 GND.n5974 585
R11269 GND.n6027 GND.n5973 585
R11270 GND.n6028 GND.n5972 585
R11271 GND.n5970 GND.n5969 585
R11272 GND.n6032 GND.n5968 585
R11273 GND.n6033 GND.n5967 585
R11274 GND.n6034 GND.n5963 585
R11275 GND.n6035 GND.n5962 585
R11276 GND.n5961 GND.n1659 585
R11277 GND.n6040 GND.n6039 585
R11278 GND.n6042 GND.n6041 585
R11279 GND.n5957 GND.n5956 585
R11280 GND.n5955 GND.n5954 585
R11281 GND.n5953 GND.n1664 585
R11282 GND.n5950 GND.n5949 585
R11283 GND.n5948 GND.n5947 585
R11284 GND.n5946 GND.n5945 585
R11285 GND.n5939 GND.n1666 585
R11286 GND.n5941 GND.n5940 585
R11287 GND.n5938 GND.n5937 585
R11288 GND.n5936 GND.n5935 585
R11289 GND.n5929 GND.n1668 585
R11290 GND.n5931 GND.n5930 585
R11291 GND.n5928 GND.n5927 585
R11292 GND.n5926 GND.n5923 585
R11293 GND.n5917 GND.n1670 585
R11294 GND.n5919 GND.n5918 585
R11295 GND.n5916 GND.n5915 585
R11296 GND.n5914 GND.n5913 585
R11297 GND.n5907 GND.n1672 585
R11298 GND.n5909 GND.n5908 585
R11299 GND.n5906 GND.n5905 585
R11300 GND.n6048 GND.n6047 585
R11301 GND.n6047 GND.n6046 585
R11302 GND.n1605 GND.n1604 585
R11303 GND.n5899 GND.n1605 585
R11304 GND.n5868 GND.n5866 585
R11305 GND.n5869 GND.n5868 585
R11306 GND.n5875 GND.n1683 585
R11307 GND.n5890 GND.n1683 585
R11308 GND.n5876 GND.n5865 585
R11309 GND.n5865 GND.n5864 585
R11310 GND.n5877 GND.n1691 585
R11311 GND.n5881 GND.n1691 585
R11312 GND.n5863 GND.n5862 585
R11313 GND.n5862 GND.n5861 585
R11314 GND.n1701 GND.n1700 585
R11315 GND.n4929 GND.n1701 585
R11316 GND.n4916 GND.n4915 585
R11317 GND.n4915 GND.n1710 585
R11318 GND.n4917 GND.n1719 585
R11319 GND.n4921 GND.n1719 585
R11320 GND.n4914 GND.n4913 585
R11321 GND.n4913 GND.n4912 585
R11322 GND.n1731 GND.n1730 585
R11323 GND.n4872 GND.n1731 585
R11324 GND.n4877 GND.n1739 585
R11325 GND.n4893 GND.n1739 585
R11326 GND.n4878 GND.n4870 585
R11327 GND.n4870 GND.n4869 585
R11328 GND.n4879 GND.n1749 585
R11329 GND.n4883 GND.n1749 585
R11330 GND.n4868 GND.n4867 585
R11331 GND.n4867 GND.n4866 585
R11332 GND.n1759 GND.n1758 585
R11333 GND.n4835 GND.n1759 585
R11334 GND.n4840 GND.n1766 585
R11335 GND.n4856 GND.n1766 585
R11336 GND.n4841 GND.n4833 585
R11337 GND.n4833 GND.n4832 585
R11338 GND.n4842 GND.n1776 585
R11339 GND.n4846 GND.n1776 585
R11340 GND.n1793 GND.n1785 585
R11341 GND.n4798 GND.n1793 585
R11342 GND.n4766 GND.n4765 585
R11343 GND.n4765 GND.n1792 585
R11344 GND.n4772 GND.n1800 585
R11345 GND.n4788 GND.n1800 585
R11346 GND.n4773 GND.n4764 585
R11347 GND.n4764 GND.n4763 585
R11348 GND.n4774 GND.n1810 585
R11349 GND.n4778 GND.n1810 585
R11350 GND.n4762 GND.n4761 585
R11351 GND.n4761 GND.n4760 585
R11352 GND.n1820 GND.n1819 585
R11353 GND.n4729 GND.n1820 585
R11354 GND.n4734 GND.n1828 585
R11355 GND.n4750 GND.n1828 585
R11356 GND.n4735 GND.n1848 585
R11357 GND.n1848 GND.n1847 585
R11358 GND.n4736 GND.n1837 585
R11359 GND.n4740 GND.n1837 585
R11360 GND.n1858 GND.n1846 585
R11361 GND.n4704 GND.n1858 585
R11362 GND.n4667 GND.n4662 585
R11363 GND.n4662 GND.n1857 585
R11364 GND.n4668 GND.n1865 585
R11365 GND.n4694 GND.n1865 585
R11366 GND.n4669 GND.n4661 585
R11367 GND.n4661 GND.n4660 585
R11368 GND.n1908 GND.n1903 585
R11369 GND.n4657 GND.n1908 585
R11370 GND.n4673 GND.n1902 585
R11371 GND.n4652 GND.n1902 585
R11372 GND.n4674 GND.n1901 585
R11373 GND.n1923 GND.n1901 585
R11374 GND.n4675 GND.n1900 585
R11375 GND.n4641 GND.n1900 585
R11376 GND.n1929 GND.n1895 585
R11377 GND.n4636 GND.n1929 585
R11378 GND.n4679 GND.n1894 585
R11379 GND.n4633 GND.n1894 585
R11380 GND.n4680 GND.n1893 585
R11381 GND.n1931 GND.n1893 585
R11382 GND.n4681 GND.n1883 585
R11383 GND.n4685 GND.n1883 585
R11384 GND.n4623 GND.n1892 585
R11385 GND.n4624 GND.n4623 585
R11386 GND.n4622 GND.n1939 585
R11387 GND.n4622 GND.n4621 585
R11388 GND.n4608 GND.n1938 585
R11389 GND.n4597 GND.n1938 585
R11390 GND.n4609 GND.n1948 585
R11391 GND.n4613 GND.n1948 585
R11392 GND.n4607 GND.n4606 585
R11393 GND.n4606 GND.n4605 585
R11394 GND.n1960 GND.n1959 585
R11395 GND.n4570 GND.n1960 585
R11396 GND.n4575 GND.n1968 585
R11397 GND.n4591 GND.n1968 585
R11398 GND.n4576 GND.n1989 585
R11399 GND.n1989 GND.n1988 585
R11400 GND.n4577 GND.n1978 585
R11401 GND.n4581 GND.n1978 585
R11402 GND.n4480 GND.n1987 585
R11403 GND.n4481 GND.n4480 585
R11404 GND.n4500 GND.n2002 585
R11405 GND.n4514 GND.n2002 585
R11406 GND.n4501 GND.n4497 585
R11407 GND.n4497 GND.n2001 585
R11408 GND.n4502 GND.n2012 585
R11409 GND.n4506 GND.n2012 585
R11410 GND.n4496 GND.n4495 585
R11411 GND.n4495 GND.n4494 585
R11412 GND.n2022 GND.n2021 585
R11413 GND.n4452 GND.n2022 585
R11414 GND.n4457 GND.n2030 585
R11415 GND.n4473 GND.n2030 585
R11416 GND.n4458 GND.n2051 585
R11417 GND.n2051 GND.n2050 585
R11418 GND.n4459 GND.n2040 585
R11419 GND.n4463 GND.n2040 585
R11420 GND.n4398 GND.n2049 585
R11421 GND.n4399 GND.n4398 585
R11422 GND.n4418 GND.n2064 585
R11423 GND.n4432 GND.n2064 585
R11424 GND.n4419 GND.n4415 585
R11425 GND.n4415 GND.n2063 585
R11426 GND.n4420 GND.n2074 585
R11427 GND.n4424 GND.n2074 585
R11428 GND.n4414 GND.n4413 585
R11429 GND.n4413 GND.n4412 585
R11430 GND.n2084 GND.n2083 585
R11431 GND.n4370 GND.n2084 585
R11432 GND.n4375 GND.n2093 585
R11433 GND.n4391 GND.n2093 585
R11434 GND.n4376 GND.n4368 585
R11435 GND.n4368 GND.n4367 585
R11436 GND.n4377 GND.n2103 585
R11437 GND.n4381 GND.n2103 585
R11438 GND.n4366 GND.n4365 585
R11439 GND.n4365 GND.n4364 585
R11440 GND.n2113 GND.n2112 585
R11441 GND.n4334 GND.n2113 585
R11442 GND.n4339 GND.n2122 585
R11443 GND.n4355 GND.n2122 585
R11444 GND.n4340 GND.n4332 585
R11445 GND.n4332 GND.n4331 585
R11446 GND.n4341 GND.n2131 585
R11447 GND.n4345 GND.n2131 585
R11448 GND.n8465 GND.n8464 585
R11449 GND.n8464 GND.n8463 585
R11450 GND.n8466 GND.n337 585
R11451 GND.n8456 GND.n337 585
R11452 GND.n8468 GND.n8467 585
R11453 GND.n8469 GND.n8468 585
R11454 GND.n322 GND.n321 585
R11455 GND.n8240 GND.n322 585
R11456 GND.n8477 GND.n8476 585
R11457 GND.n8476 GND.n8475 585
R11458 GND.n8478 GND.n316 585
R11459 GND.n8246 GND.n316 585
R11460 GND.n8480 GND.n8479 585
R11461 GND.n8481 GND.n8480 585
R11462 GND.n302 GND.n301 585
R11463 GND.n8231 GND.n302 585
R11464 GND.n8489 GND.n8488 585
R11465 GND.n8488 GND.n8487 585
R11466 GND.n8490 GND.n296 585
R11467 GND.n8222 GND.n296 585
R11468 GND.n8492 GND.n8491 585
R11469 GND.n8493 GND.n8492 585
R11470 GND.n281 GND.n280 585
R11471 GND.n8215 GND.n281 585
R11472 GND.n8501 GND.n8500 585
R11473 GND.n8500 GND.n8499 585
R11474 GND.n8502 GND.n275 585
R11475 GND.n8207 GND.n275 585
R11476 GND.n8504 GND.n8503 585
R11477 GND.n8505 GND.n8504 585
R11478 GND.n260 GND.n259 585
R11479 GND.n8200 GND.n260 585
R11480 GND.n8513 GND.n8512 585
R11481 GND.n8512 GND.n8511 585
R11482 GND.n8514 GND.n254 585
R11483 GND.n8192 GND.n254 585
R11484 GND.n8516 GND.n8515 585
R11485 GND.n8517 GND.n8516 585
R11486 GND.n240 GND.n239 585
R11487 GND.n8185 GND.n240 585
R11488 GND.n8525 GND.n8524 585
R11489 GND.n8524 GND.n8523 585
R11490 GND.n8526 GND.n234 585
R11491 GND.n8177 GND.n234 585
R11492 GND.n8528 GND.n8527 585
R11493 GND.n8529 GND.n8528 585
R11494 GND.n219 GND.n218 585
R11495 GND.n8170 GND.n219 585
R11496 GND.n8537 GND.n8536 585
R11497 GND.n8536 GND.n8535 585
R11498 GND.n8538 GND.n213 585
R11499 GND.n8162 GND.n213 585
R11500 GND.n8540 GND.n8539 585
R11501 GND.n8541 GND.n8540 585
R11502 GND.n198 GND.n197 585
R11503 GND.n8155 GND.n198 585
R11504 GND.n8549 GND.n8548 585
R11505 GND.n8548 GND.n8547 585
R11506 GND.n8550 GND.n193 585
R11507 GND.n8147 GND.n193 585
R11508 GND.n8552 GND.n8551 585
R11509 GND.n8553 GND.n8552 585
R11510 GND.n176 GND.n174 585
R11511 GND.n8140 GND.n176 585
R11512 GND.n8561 GND.n8560 585
R11513 GND.n8560 GND.n8559 585
R11514 GND.n175 GND.n173 585
R11515 GND.n8132 GND.n175 585
R11516 GND.n8124 GND.n8123 585
R11517 GND.n8125 GND.n8124 585
R11518 GND.n165 GND.n163 585
R11519 GND.n435 GND.n163 585
R11520 GND.n8565 GND.n8564 585
R11521 GND.n8566 GND.n8565 585
R11522 GND.n164 GND.n162 585
R11523 GND.n8032 GND.n162 585
R11524 GND.n8018 GND.n8017 585
R11525 GND.n8018 GND.n441 585
R11526 GND.n8019 GND.n171 585
R11527 GND.n8020 GND.n8019 585
R11528 GND.n8016 GND.n454 585
R11529 GND.n8016 GND.n8015 585
R11530 GND.n7987 GND.n453 585
R11531 GND.n8006 GND.n453 585
R11532 GND.n7988 GND.n473 585
R11533 GND.n7974 GND.n473 585
R11534 GND.n7990 GND.n7989 585
R11535 GND.n7991 GND.n7990 585
R11536 GND.n474 GND.n472 585
R11537 GND.n7968 GND.n472 585
R11538 GND.n7983 GND.n7982 585
R11539 GND.n7982 GND.n7981 585
R11540 GND.n477 GND.n476 585
R11541 GND.n7964 GND.n477 585
R11542 GND.n7951 GND.n500 585
R11543 GND.n7937 GND.n500 585
R11544 GND.n7953 GND.n7952 585
R11545 GND.n7954 GND.n7953 585
R11546 GND.n501 GND.n499 585
R11547 GND.n549 GND.n499 585
R11548 GND.n7946 GND.n7945 585
R11549 GND.n7945 GND.n7944 585
R11550 GND.n504 GND.n503 585
R11551 GND.n7882 GND.n504 585
R11552 GND.n7898 GND.n7897 585
R11553 GND.n7899 GND.n7898 585
R11554 GND.n532 GND.n531 585
R11555 GND.n531 GND.n526 585
R11556 GND.n7893 GND.n7892 585
R11557 GND.n7892 GND.n7891 585
R11558 GND.n535 GND.n534 585
R11559 GND.n7869 GND.n535 585
R11560 GND.n7860 GND.n7859 585
R11561 GND.n7861 GND.n7860 585
R11562 GND.n566 GND.n565 585
R11563 GND.n7846 GND.n565 585
R11564 GND.n7855 GND.n7854 585
R11565 GND.n7854 GND.n7853 585
R11566 GND.n569 GND.n568 585
R11567 GND.n7837 GND.n569 585
R11568 GND.n7833 GND.n7832 585
R11569 GND.n7834 GND.n7833 585
R11570 GND.n588 GND.n587 585
R11571 GND.n7809 GND.n587 585
R11572 GND.n7828 GND.n7827 585
R11573 GND.n7827 GND.n7826 585
R11574 GND.n591 GND.n590 585
R11575 GND.n7815 GND.n591 585
R11576 GND.n7798 GND.n614 585
R11577 GND.n7784 GND.n614 585
R11578 GND.n7800 GND.n7799 585
R11579 GND.n7801 GND.n7800 585
R11580 GND.n615 GND.n613 585
R11581 GND.n7778 GND.n613 585
R11582 GND.n7793 GND.n7792 585
R11583 GND.n7792 GND.n7791 585
R11584 GND.n618 GND.n617 585
R11585 GND.n7774 GND.n618 585
R11586 GND.n7761 GND.n642 585
R11587 GND.n7741 GND.n642 585
R11588 GND.n7763 GND.n7762 585
R11589 GND.n7764 GND.n7763 585
R11590 GND.n643 GND.n641 585
R11591 GND.n7747 GND.n641 585
R11592 GND.n7756 GND.n7755 585
R11593 GND.n7755 GND.n7754 585
R11594 GND.n646 GND.n645 585
R11595 GND.n7737 GND.n646 585
R11596 GND.n7723 GND.n7722 585
R11597 GND.n7721 GND.n708 585
R11598 GND.n7720 GND.n707 585
R11599 GND.n7725 GND.n707 585
R11600 GND.n7719 GND.n7718 585
R11601 GND.n7717 GND.n7716 585
R11602 GND.n7715 GND.n7714 585
R11603 GND.n7713 GND.n7712 585
R11604 GND.n7711 GND.n7710 585
R11605 GND.n7709 GND.n717 585
R11606 GND.n7708 GND.n7707 585
R11607 GND.n7706 GND.n7705 585
R11608 GND.n7704 GND.n7703 585
R11609 GND.n7702 GND.n7701 585
R11610 GND.n7700 GND.n7699 585
R11611 GND.n7698 GND.n7697 585
R11612 GND.n7696 GND.n7695 585
R11613 GND.n7694 GND.n7693 585
R11614 GND.n7692 GND.n7691 585
R11615 GND.n7689 GND.n7688 585
R11616 GND.n7687 GND.n7686 585
R11617 GND.n7685 GND.n7684 585
R11618 GND.n7683 GND.n7682 585
R11619 GND.n7682 GND.n7597 585
R11620 GND.n7681 GND.n7680 585
R11621 GND.n7679 GND.n7678 585
R11622 GND.n7677 GND.n7676 585
R11623 GND.n7675 GND.n7674 585
R11624 GND.n7673 GND.n7672 585
R11625 GND.n7671 GND.n7670 585
R11626 GND.n7669 GND.n7668 585
R11627 GND.n7667 GND.n7666 585
R11628 GND.n7665 GND.n7664 585
R11629 GND.n7663 GND.n7662 585
R11630 GND.n7661 GND.n7660 585
R11631 GND.n7659 GND.n7658 585
R11632 GND.n7657 GND.n7656 585
R11633 GND.n7655 GND.n7654 585
R11634 GND.n7653 GND.n7652 585
R11635 GND.n7651 GND.n7650 585
R11636 GND.n7649 GND.n7648 585
R11637 GND.n7647 GND.n7646 585
R11638 GND.n7645 GND.n7644 585
R11639 GND.n7643 GND.n7642 585
R11640 GND.n7641 GND.n7640 585
R11641 GND.n7639 GND.n7638 585
R11642 GND.n7637 GND.n7636 585
R11643 GND.n7635 GND.n7634 585
R11644 GND.n7633 GND.n7632 585
R11645 GND.n7627 GND.n657 585
R11646 GND.n8343 GND.n8342 585
R11647 GND.n8349 GND.n8348 585
R11648 GND.n8351 GND.n8350 585
R11649 GND.n8353 GND.n8352 585
R11650 GND.n8355 GND.n8354 585
R11651 GND.n8357 GND.n8356 585
R11652 GND.n8359 GND.n8358 585
R11653 GND.n8361 GND.n8360 585
R11654 GND.n8363 GND.n8362 585
R11655 GND.n8366 GND.n8365 585
R11656 GND.n8364 GND.n8332 585
R11657 GND.n8371 GND.n8370 585
R11658 GND.n8373 GND.n8372 585
R11659 GND.n8375 GND.n8374 585
R11660 GND.n8377 GND.n8376 585
R11661 GND.n8379 GND.n8378 585
R11662 GND.n8381 GND.n8380 585
R11663 GND.n8383 GND.n8382 585
R11664 GND.n8385 GND.n8384 585
R11665 GND.n8388 GND.n8387 585
R11666 GND.n8386 GND.n8322 585
R11667 GND.n8393 GND.n8392 585
R11668 GND.n8395 GND.n8394 585
R11669 GND.n8397 GND.n8396 585
R11670 GND.n8399 GND.n8398 585
R11671 GND.n8401 GND.n8400 585
R11672 GND.n8403 GND.n8402 585
R11673 GND.n8405 GND.n8404 585
R11674 GND.n8407 GND.n8406 585
R11675 GND.n8409 GND.n8408 585
R11676 GND.n8411 GND.n8410 585
R11677 GND.n8416 GND.n8415 585
R11678 GND.n8418 GND.n8417 585
R11679 GND.n8420 GND.n8419 585
R11680 GND.n8422 GND.n8421 585
R11681 GND.n8424 GND.n8423 585
R11682 GND.n8426 GND.n8425 585
R11683 GND.n8428 GND.n8427 585
R11684 GND.n8430 GND.n8429 585
R11685 GND.n8304 GND.n8301 585
R11686 GND.n8434 GND.n8305 585
R11687 GND.n8436 GND.n8435 585
R11688 GND.n8438 GND.n8437 585
R11689 GND.n8440 GND.n8439 585
R11690 GND.n8442 GND.n8441 585
R11691 GND.n8443 GND.n8290 585
R11692 GND.n8445 GND.n8444 585
R11693 GND.n8291 GND.n8289 585
R11694 GND.n8292 GND.n342 585
R11695 GND.n8447 GND.n342 585
R11696 GND.n8459 GND.n344 585
R11697 GND.n8463 GND.n344 585
R11698 GND.n8458 GND.n8457 585
R11699 GND.n8457 GND.n8456 585
R11700 GND.n350 GND.n334 585
R11701 GND.n8469 GND.n334 585
R11702 GND.n8239 GND.n8238 585
R11703 GND.n8240 GND.n8239 585
R11704 GND.n8237 GND.n324 585
R11705 GND.n8475 GND.n324 585
R11706 GND.n8236 GND.n393 585
R11707 GND.n8246 GND.n393 585
R11708 GND.n8234 GND.n314 585
R11709 GND.n8481 GND.n314 585
R11710 GND.n8233 GND.n8232 585
R11711 GND.n8232 GND.n8231 585
R11712 GND.n399 GND.n304 585
R11713 GND.n8487 GND.n304 585
R11714 GND.n8221 GND.n8220 585
R11715 GND.n8222 GND.n8221 585
R11716 GND.n8218 GND.n293 585
R11717 GND.n8493 GND.n293 585
R11718 GND.n8217 GND.n8216 585
R11719 GND.n8216 GND.n8215 585
R11720 GND.n403 GND.n283 585
R11721 GND.n8499 GND.n283 585
R11722 GND.n8206 GND.n8205 585
R11723 GND.n8207 GND.n8206 585
R11724 GND.n8203 GND.n272 585
R11725 GND.n8505 GND.n272 585
R11726 GND.n8202 GND.n8201 585
R11727 GND.n8201 GND.n8200 585
R11728 GND.n407 GND.n262 585
R11729 GND.n8511 GND.n262 585
R11730 GND.n8191 GND.n8190 585
R11731 GND.n8192 GND.n8191 585
R11732 GND.n8188 GND.n252 585
R11733 GND.n8517 GND.n252 585
R11734 GND.n8187 GND.n8186 585
R11735 GND.n8186 GND.n8185 585
R11736 GND.n412 GND.n242 585
R11737 GND.n8523 GND.n242 585
R11738 GND.n8176 GND.n8175 585
R11739 GND.n8177 GND.n8176 585
R11740 GND.n8173 GND.n231 585
R11741 GND.n8529 GND.n231 585
R11742 GND.n8172 GND.n8171 585
R11743 GND.n8171 GND.n8170 585
R11744 GND.n416 GND.n221 585
R11745 GND.n8535 GND.n221 585
R11746 GND.n8161 GND.n8160 585
R11747 GND.n8162 GND.n8161 585
R11748 GND.n8158 GND.n210 585
R11749 GND.n8541 GND.n210 585
R11750 GND.n8157 GND.n8156 585
R11751 GND.n8156 GND.n8155 585
R11752 GND.n420 GND.n200 585
R11753 GND.n8547 GND.n200 585
R11754 GND.n8146 GND.n8145 585
R11755 GND.n8147 GND.n8146 585
R11756 GND.n8143 GND.n190 585
R11757 GND.n8553 GND.n190 585
R11758 GND.n8142 GND.n8141 585
R11759 GND.n8141 GND.n8140 585
R11760 GND.n424 GND.n178 585
R11761 GND.n8559 GND.n178 585
R11762 GND.n8131 GND.n8130 585
R11763 GND.n8132 GND.n8131 585
R11764 GND.n431 GND.n430 585
R11765 GND.n8125 GND.n430 585
R11766 GND.n8026 GND.n8025 585
R11767 GND.n8025 GND.n435 585
R11768 GND.n8027 GND.n159 585
R11769 GND.n8566 GND.n159 585
R11770 GND.n8024 GND.n442 585
R11771 GND.n8032 GND.n442 585
R11772 GND.n8023 GND.n8022 585
R11773 GND.n8022 GND.n441 585
R11774 GND.n8021 GND.n446 585
R11775 GND.n8021 GND.n8020 585
R11776 GND.n8009 GND.n448 585
R11777 GND.n8015 GND.n448 585
R11778 GND.n8008 GND.n8007 585
R11779 GND.n8007 GND.n8006 585
R11780 GND.n461 GND.n460 585
R11781 GND.n7974 GND.n461 585
R11782 GND.n7971 GND.n469 585
R11783 GND.n7991 GND.n469 585
R11784 GND.n7970 GND.n7969 585
R11785 GND.n7969 GND.n7968 585
R11786 GND.n7967 GND.n479 585
R11787 GND.n7981 GND.n479 585
R11788 GND.n7966 GND.n7965 585
R11789 GND.n7965 GND.n7964 585
R11790 GND.n489 GND.n487 585
R11791 GND.n7937 GND.n489 585
R11792 GND.n548 GND.n496 585
R11793 GND.n7954 GND.n496 585
R11794 GND.n551 GND.n550 585
R11795 GND.n550 GND.n549 585
R11796 GND.n552 GND.n506 585
R11797 GND.n7944 GND.n506 585
R11798 GND.n7884 GND.n7883 585
R11799 GND.n7883 GND.n7882 585
R11800 GND.n7885 GND.n527 585
R11801 GND.n7899 GND.n527 585
R11802 GND.n547 GND.n546 585
R11803 GND.n546 GND.n526 585
R11804 GND.n7866 GND.n537 585
R11805 GND.n7891 GND.n537 585
R11806 GND.n7868 GND.n7867 585
R11807 GND.n7869 GND.n7868 585
R11808 GND.n560 GND.n559 585
R11809 GND.n7861 GND.n559 585
R11810 GND.n7848 GND.n7847 585
R11811 GND.n7847 GND.n7846 585
R11812 GND.n7849 GND.n571 585
R11813 GND.n7853 GND.n571 585
R11814 GND.n7836 GND.n577 585
R11815 GND.n7837 GND.n7836 585
R11816 GND.n7835 GND.n584 585
R11817 GND.n7835 GND.n7834 585
R11818 GND.n7819 GND.n583 585
R11819 GND.n7809 GND.n583 585
R11820 GND.n7818 GND.n593 585
R11821 GND.n7826 GND.n593 585
R11822 GND.n7817 GND.n7816 585
R11823 GND.n7816 GND.n7815 585
R11824 GND.n602 GND.n600 585
R11825 GND.n7784 GND.n602 585
R11826 GND.n7781 GND.n610 585
R11827 GND.n7801 GND.n610 585
R11828 GND.n7780 GND.n7779 585
R11829 GND.n7779 GND.n7778 585
R11830 GND.n7777 GND.n620 585
R11831 GND.n7791 GND.n620 585
R11832 GND.n7776 GND.n7775 585
R11833 GND.n7775 GND.n7774 585
R11834 GND.n630 GND.n628 585
R11835 GND.n7741 GND.n630 585
R11836 GND.n7746 GND.n638 585
R11837 GND.n7764 GND.n638 585
R11838 GND.n7749 GND.n7748 585
R11839 GND.n7748 GND.n7747 585
R11840 GND.n7750 GND.n648 585
R11841 GND.n7754 GND.n648 585
R11842 GND.n7739 GND.n7738 585
R11843 GND.n7738 GND.n7737 585
R11844 GND.n4127 GND.n4126 585
R11845 GND.n4128 GND.n4127 585
R11846 GND.n8264 GND.n8263 585
R11847 GND.n8265 GND.n8264 585
R11848 GND.n8260 GND.n383 585
R11849 GND.n383 GND.n346 585
R11850 GND.n8259 GND.n8258 585
R11851 GND.n8258 GND.n343 585
R11852 GND.n8257 GND.n387 585
R11853 GND.n8257 GND.n336 585
R11854 GND.n8256 GND.n8255 585
R11855 GND.n8256 GND.n333 585
R11856 GND.n389 GND.n388 585
R11857 GND.n388 GND.n326 585
R11858 GND.n8250 GND.n8249 585
R11859 GND.n8249 GND.n323 585
R11860 GND.n8248 GND.n391 585
R11861 GND.n8248 GND.n8247 585
R11862 GND.n8077 GND.n392 585
R11863 GND.n392 GND.n313 585
R11864 GND.n8079 GND.n8078 585
R11865 GND.n8079 GND.n306 585
R11866 GND.n8081 GND.n8080 585
R11867 GND.n8080 GND.n303 585
R11868 GND.n8082 GND.n8070 585
R11869 GND.n8070 GND.n295 585
R11870 GND.n8084 GND.n8083 585
R11871 GND.n8084 GND.n292 585
R11872 GND.n8085 GND.n8069 585
R11873 GND.n8085 GND.n285 585
R11874 GND.n8087 GND.n8086 585
R11875 GND.n8086 GND.n282 585
R11876 GND.n8088 GND.n8064 585
R11877 GND.n8064 GND.n274 585
R11878 GND.n8090 GND.n8089 585
R11879 GND.n8090 GND.n271 585
R11880 GND.n8091 GND.n8063 585
R11881 GND.n8091 GND.n264 585
R11882 GND.n8093 GND.n8092 585
R11883 GND.n8092 GND.n261 585
R11884 GND.n8094 GND.n8058 585
R11885 GND.n8058 GND.n411 585
R11886 GND.n8096 GND.n8095 585
R11887 GND.n8096 GND.n251 585
R11888 GND.n8097 GND.n8057 585
R11889 GND.n8097 GND.n244 585
R11890 GND.n8099 GND.n8098 585
R11891 GND.n8098 GND.n241 585
R11892 GND.n8100 GND.n8052 585
R11893 GND.n8052 GND.n233 585
R11894 GND.n8102 GND.n8101 585
R11895 GND.n8102 GND.n230 585
R11896 GND.n8103 GND.n8051 585
R11897 GND.n8103 GND.n223 585
R11898 GND.n8105 GND.n8104 585
R11899 GND.n8104 GND.n220 585
R11900 GND.n8106 GND.n8046 585
R11901 GND.n8046 GND.n212 585
R11902 GND.n8108 GND.n8107 585
R11903 GND.n8108 GND.n209 585
R11904 GND.n8109 GND.n8045 585
R11905 GND.n8109 GND.n202 585
R11906 GND.n8111 GND.n8110 585
R11907 GND.n8110 GND.n199 585
R11908 GND.n8112 GND.n8040 585
R11909 GND.n8040 GND.n192 585
R11910 GND.n8114 GND.n8113 585
R11911 GND.n8114 GND.n189 585
R11912 GND.n8115 GND.n8039 585
R11913 GND.n8115 GND.n180 585
R11914 GND.n8117 GND.n8116 585
R11915 GND.n8116 GND.n177 585
R11916 GND.n8119 GND.n437 585
R11917 GND.n437 GND.n429 585
R11918 GND.n8121 GND.n8120 585
R11919 GND.n8122 GND.n8121 585
R11920 GND.n8037 GND.n436 585
R11921 GND.n436 GND.n160 585
R11922 GND.n8036 GND.n8035 585
R11923 GND.n8035 GND.n158 585
R11924 GND.n8034 GND.n440 585
R11925 GND.n8034 GND.n8033 585
R11926 GND.n7920 GND.n439 585
R11927 GND.n451 GND.n439 585
R11928 GND.n7923 GND.n7922 585
R11929 GND.n7923 GND.n449 585
R11930 GND.n7925 GND.n7924 585
R11931 GND.n7924 GND.n455 585
R11932 GND.n7927 GND.n7917 585
R11933 GND.n7917 GND.n462 585
R11934 GND.n7929 GND.n7928 585
R11935 GND.n7929 GND.n470 585
R11936 GND.n7930 GND.n7916 585
R11937 GND.n7930 GND.n468 585
R11938 GND.n7932 GND.n7931 585
R11939 GND.n7931 GND.n481 585
R11940 GND.n7933 GND.n517 585
R11941 GND.n517 GND.n478 585
R11942 GND.n7935 GND.n7934 585
R11943 GND.n7936 GND.n7935 585
R11944 GND.n518 GND.n516 585
R11945 GND.n516 GND.n497 585
R11946 GND.n7910 GND.n7909 585
R11947 GND.n7909 GND.n495 585
R11948 GND.n7908 GND.n520 585
R11949 GND.n7908 GND.n508 585
R11950 GND.n7907 GND.n7906 585
R11951 GND.n7907 GND.n505 585
R11952 GND.n522 GND.n521 585
R11953 GND.n529 GND.n521 585
R11954 GND.n7902 GND.n7901 585
R11955 GND.n7901 GND.n7900 585
R11956 GND.n525 GND.n524 585
R11957 GND.n539 GND.n525 585
R11958 GND.n7490 GND.n7489 585
R11959 GND.n7490 GND.n536 585
R11960 GND.n7492 GND.n7491 585
R11961 GND.n7491 GND.n558 585
R11962 GND.n7493 GND.n7483 585
R11963 GND.n7483 GND.n564 585
R11964 GND.n7495 GND.n7494 585
R11965 GND.n7495 GND.n573 585
R11966 GND.n7496 GND.n7482 585
R11967 GND.n7496 GND.n570 585
R11968 GND.n7498 GND.n7497 585
R11969 GND.n7497 GND.n582 585
R11970 GND.n7499 GND.n7477 585
R11971 GND.n7477 GND.n585 585
R11972 GND.n7501 GND.n7500 585
R11973 GND.n7501 GND.n595 585
R11974 GND.n7502 GND.n7476 585
R11975 GND.n7502 GND.n592 585
R11976 GND.n7504 GND.n7503 585
R11977 GND.n7503 GND.n603 585
R11978 GND.n7505 GND.n7471 585
R11979 GND.n7471 GND.n611 585
R11980 GND.n7507 GND.n7506 585
R11981 GND.n7507 GND.n609 585
R11982 GND.n7508 GND.n7470 585
R11983 GND.n7508 GND.n622 585
R11984 GND.n7510 GND.n7509 585
R11985 GND.n7509 GND.n619 585
R11986 GND.n7511 GND.n7465 585
R11987 GND.n7465 GND.n631 585
R11988 GND.n7513 GND.n7512 585
R11989 GND.n7513 GND.n639 585
R11990 GND.n7514 GND.n7464 585
R11991 GND.n7514 GND.n637 585
R11992 GND.n7516 GND.n7515 585
R11993 GND.n7515 GND.n650 585
R11994 GND.n7517 GND.n7459 585
R11995 GND.n7459 GND.n647 585
R11996 GND.n7519 GND.n7518 585
R11997 GND.n7519 GND.n658 585
R11998 GND.n7520 GND.n7458 585
R11999 GND.n7520 GND.n706 585
R12000 GND.n7522 GND.n7521 585
R12001 GND.n7521 GND.n671 585
R12002 GND.n7523 GND.n7453 585
R12003 GND.n7453 GND.n7452 585
R12004 GND.n7525 GND.n7524 585
R12005 GND.n7526 GND.n7525 585
R12006 GND.n7451 GND.n7450 585
R12007 GND.n7527 GND.n7451 585
R12008 GND.n7530 GND.n7529 585
R12009 GND.n7529 GND.n7528 585
R12010 GND.n7531 GND.n801 585
R12011 GND.n801 GND.n739 585
R12012 GND.n7533 GND.n7532 585
R12013 GND.n7534 GND.n7533 585
R12014 GND.n802 GND.n800 585
R12015 GND.n808 GND.n800 585
R12016 GND.n7444 GND.n7443 585
R12017 GND.n7443 GND.n7442 585
R12018 GND.n805 GND.n804 585
R12019 GND.n812 GND.n805 585
R12020 GND.n7357 GND.n825 585
R12021 GND.n825 GND.n818 585
R12022 GND.n7359 GND.n7358 585
R12023 GND.n7360 GND.n7359 585
R12024 GND.n826 GND.n824 585
R12025 GND.n824 GND.n822 585
R12026 GND.n7352 GND.n7351 585
R12027 GND.n7351 GND.n7350 585
R12028 GND.n829 GND.n828 585
R12029 GND.n834 GND.n829 585
R12030 GND.n7334 GND.n7333 585
R12031 GND.n7335 GND.n7334 585
R12032 GND.n842 GND.n841 585
R12033 GND.n848 GND.n841 585
R12034 GND.n7329 GND.n7328 585
R12035 GND.n7328 GND.n7327 585
R12036 GND.n845 GND.n844 585
R12037 GND.n852 GND.n845 585
R12038 GND.n7298 GND.n866 585
R12039 GND.n866 GND.n859 585
R12040 GND.n7300 GND.n7299 585
R12041 GND.n7301 GND.n7300 585
R12042 GND.n867 GND.n865 585
R12043 GND.n865 GND.n863 585
R12044 GND.n7293 GND.n7292 585
R12045 GND.n7292 GND.n7291 585
R12046 GND.n870 GND.n869 585
R12047 GND.n7283 GND.n870 585
R12048 GND.n7227 GND.n7226 585
R12049 GND.n7227 GND.n883 585
R12050 GND.n7229 GND.n7228 585
R12051 GND.n7228 GND.n882 585
R12052 GND.n7230 GND.n7220 585
R12053 GND.n7220 GND.n887 585
R12054 GND.n7232 GND.n7231 585
R12055 GND.n7232 GND.n893 585
R12056 GND.n7233 GND.n7219 585
R12057 GND.n7233 GND.n891 585
R12058 GND.n7235 GND.n7234 585
R12059 GND.n7234 GND.n897 585
R12060 GND.n7236 GND.n910 585
R12061 GND.n910 GND.n903 585
R12062 GND.n7238 GND.n7237 585
R12063 GND.n7239 GND.n7238 585
R12064 GND.n911 GND.n909 585
R12065 GND.n909 GND.n907 585
R12066 GND.n7213 GND.n7212 585
R12067 GND.n7212 GND.n7211 585
R12068 GND.n914 GND.n913 585
R12069 GND.n7203 GND.n914 585
R12070 GND.n7163 GND.n7162 585
R12071 GND.n7163 GND.n925 585
R12072 GND.n7164 GND.n7159 585
R12073 GND.n7164 GND.n924 585
R12074 GND.n7166 GND.n7165 585
R12075 GND.n7165 GND.n929 585
R12076 GND.n7167 GND.n942 585
R12077 GND.n942 GND.n935 585
R12078 GND.n7169 GND.n7168 585
R12079 GND.n7170 GND.n7169 585
R12080 GND.n943 GND.n941 585
R12081 GND.n941 GND.n939 585
R12082 GND.n7153 GND.n7152 585
R12083 GND.n7152 GND.n7151 585
R12084 GND.n946 GND.n945 585
R12085 GND.n7143 GND.n946 585
R12086 GND.n7121 GND.n7120 585
R12087 GND.n7120 GND.n959 585
R12088 GND.n7122 GND.n967 585
R12089 GND.n967 GND.n958 585
R12090 GND.n7124 GND.n7123 585
R12091 GND.n7125 GND.n7124 585
R12092 GND.n968 GND.n966 585
R12093 GND.n974 GND.n966 585
R12094 GND.n7114 GND.n7113 585
R12095 GND.n7113 GND.n7112 585
R12096 GND.n971 GND.n970 585
R12097 GND.n978 GND.n971 585
R12098 GND.n7084 GND.n992 585
R12099 GND.n992 GND.n985 585
R12100 GND.n7086 GND.n7085 585
R12101 GND.n7087 GND.n7086 585
R12102 GND.n993 GND.n991 585
R12103 GND.n991 GND.n989 585
R12104 GND.n7079 GND.n7078 585
R12105 GND.n7078 GND.n7077 585
R12106 GND.n996 GND.n995 585
R12107 GND.n7069 GND.n996 585
R12108 GND.n7031 GND.n7030 585
R12109 GND.n7031 GND.n1009 585
R12110 GND.n7032 GND.n7027 585
R12111 GND.n7032 GND.n1008 585
R12112 GND.n7034 GND.n7033 585
R12113 GND.n7033 GND.n1013 585
R12114 GND.n7035 GND.n1026 585
R12115 GND.n1026 GND.n1019 585
R12116 GND.n7037 GND.n7036 585
R12117 GND.n7038 GND.n7037 585
R12118 GND.n1027 GND.n1025 585
R12119 GND.n1025 GND.n1023 585
R12120 GND.n7021 GND.n7020 585
R12121 GND.n7020 GND.n7019 585
R12122 GND.n1030 GND.n1029 585
R12123 GND.n7011 GND.n1030 585
R12124 GND.n6988 GND.n6987 585
R12125 GND.n6987 GND.n1037 585
R12126 GND.n6989 GND.n1050 585
R12127 GND.n1050 GND.n1041 585
R12128 GND.n6991 GND.n6990 585
R12129 GND.n6992 GND.n6991 585
R12130 GND.n1051 GND.n1049 585
R12131 GND.n1081 GND.n1049 585
R12132 GND.n6981 GND.n6980 585
R12133 GND.n6980 GND.n6979 585
R12134 GND.n1054 GND.n1053 585
R12135 GND.n6905 GND.n1054 585
R12136 GND.n6893 GND.n6892 585
R12137 GND.n6894 GND.n6893 585
R12138 GND.n1097 GND.n1096 585
R12139 GND.n6735 GND.n1096 585
R12140 GND.n6888 GND.n6887 585
R12141 GND.n6887 GND.n6886 585
R12142 GND.n1100 GND.n1099 585
R12143 GND.n6741 GND.n1100 585
R12144 GND.n6873 GND.n6872 585
R12145 GND.t209 GND.n6873 585
R12146 GND.n1114 GND.n1113 585
R12147 GND.n6710 GND.n1113 585
R12148 GND.n6868 GND.n6867 585
R12149 GND.n6867 GND.n6866 585
R12150 GND.n1117 GND.n1116 585
R12151 GND.n1203 GND.n1117 585
R12152 GND.n6857 GND.n6856 585
R12153 GND.n6858 GND.n6857 585
R12154 GND.n1130 GND.n1129 585
R12155 GND.n6789 GND.n1129 585
R12156 GND.n6852 GND.n6851 585
R12157 GND.n6851 GND.n6850 585
R12158 GND.n1133 GND.n1132 585
R12159 GND.t203 GND.n1133 585
R12160 GND.n6841 GND.n6840 585
R12161 GND.n6842 GND.n6841 585
R12162 GND.n1146 GND.n1145 585
R12163 GND.n6803 GND.n1145 585
R12164 GND.n6836 GND.n6835 585
R12165 GND.n6835 GND.n6834 585
R12166 GND.n1149 GND.n1148 585
R12167 GND.n6809 GND.n1149 585
R12168 GND.n6825 GND.n6824 585
R12169 GND.n6826 GND.n6825 585
R12170 GND.n1162 GND.n1161 585
R12171 GND.n6460 GND.n1161 585
R12172 GND.n6820 GND.n6819 585
R12173 GND.n6819 GND.t213 585
R12174 GND.n1165 GND.n1164 585
R12175 GND.n1210 GND.n1165 585
R12176 GND.n6671 GND.n6670 585
R12177 GND.n6672 GND.n6671 585
R12178 GND.n1219 GND.n1218 585
R12179 GND.n1218 GND.n1214 585
R12180 GND.n6666 GND.n6665 585
R12181 GND.n6665 GND.n6664 585
R12182 GND.n1222 GND.n1221 585
R12183 GND.n1397 GND.n1222 585
R12184 GND.n6646 GND.n6645 585
R12185 GND.n6647 GND.n6646 585
R12186 GND.n1236 GND.n1235 585
R12187 GND.t199 GND.n1235 585
R12188 GND.n6641 GND.n6640 585
R12189 GND.n6640 GND.n6639 585
R12190 GND.n1239 GND.n1238 585
R12191 GND.n6445 GND.n1239 585
R12192 GND.n6630 GND.n6629 585
R12193 GND.n6631 GND.n6630 585
R12194 GND.n1252 GND.n1251 585
R12195 GND.n1379 GND.n1251 585
R12196 GND.n6625 GND.n6624 585
R12197 GND.n6624 GND.n6623 585
R12198 GND.n1255 GND.n1254 585
R12199 GND.n1372 GND.n1255 585
R12200 GND.n6615 GND.n6614 585
R12201 GND.t207 GND.n6615 585
R12202 GND.n1268 GND.n1267 585
R12203 GND.n1365 GND.n1267 585
R12204 GND.n6610 GND.n6609 585
R12205 GND.n6609 GND.n6608 585
R12206 GND.n1271 GND.n1270 585
R12207 GND.n1358 GND.n1271 585
R12208 GND.n6599 GND.n6598 585
R12209 GND.n6600 GND.n6599 585
R12210 GND.n1284 GND.n1283 585
R12211 GND.n1351 GND.n1283 585
R12212 GND.n6594 GND.n6593 585
R12213 GND.n6593 GND.n6592 585
R12214 GND.n1287 GND.n1286 585
R12215 GND.t201 GND.n1287 585
R12216 GND.n6583 GND.n6582 585
R12217 GND.n6584 GND.n6583 585
R12218 GND.n1300 GND.n1299 585
R12219 GND.n1339 GND.n1299 585
R12220 GND.n6578 GND.n6577 585
R12221 GND.n6577 GND.n6576 585
R12222 GND.n1303 GND.n1302 585
R12223 GND.n1335 GND.n1303 585
R12224 GND.n6567 GND.n6566 585
R12225 GND.n6568 GND.n6567 585
R12226 GND.n1315 GND.n1314 585
R12227 GND.n1329 GND.n1314 585
R12228 GND.n6562 GND.n6561 585
R12229 GND.n6561 GND.t211 585
R12230 GND.n1318 GND.n1317 585
R12231 GND.n6404 GND.n1318 585
R12232 GND.n6391 GND.n1432 585
R12233 GND.n6245 GND.n1432 585
R12234 GND.n6393 GND.n6392 585
R12235 GND.n6394 GND.n6393 585
R12236 GND.n1433 GND.n1431 585
R12237 GND.n6237 GND.n1431 585
R12238 GND.n6386 GND.n6385 585
R12239 GND.n6385 GND.n6384 585
R12240 GND.n1436 GND.n1435 585
R12241 GND.n6199 GND.n1436 585
R12242 GND.n6376 GND.n6375 585
R12243 GND.t195 GND.n6376 585
R12244 GND.n1449 GND.n1448 585
R12245 GND.n6192 GND.n1448 585
R12246 GND.n6371 GND.n6370 585
R12247 GND.n6370 GND.n6369 585
R12248 GND.n1452 GND.n1451 585
R12249 GND.n6185 GND.n1452 585
R12250 GND.n6360 GND.n6359 585
R12251 GND.n6361 GND.n6360 585
R12252 GND.n1465 GND.n1464 585
R12253 GND.n6178 GND.n1464 585
R12254 GND.n6355 GND.n6354 585
R12255 GND.n6354 GND.n6353 585
R12256 GND.n1468 GND.n1467 585
R12257 GND.t205 GND.n1468 585
R12258 GND.n6344 GND.n6343 585
R12259 GND.n6345 GND.n6344 585
R12260 GND.n1481 GND.n1480 585
R12261 GND.n6306 GND.n1480 585
R12262 GND.n6339 GND.n6338 585
R12263 GND.n6338 GND.n6337 585
R12264 GND.n1484 GND.n1483 585
R12265 GND.n6312 GND.n1484 585
R12266 GND.n6328 GND.n6327 585
R12267 GND.n6329 GND.n6328 585
R12268 GND.n1497 GND.n1496 585
R12269 GND.n5611 GND.n1496 585
R12270 GND.n6323 GND.n6322 585
R12271 GND.n6322 GND.t197 585
R12272 GND.n1500 GND.n1499 585
R12273 GND.n1531 GND.n1500 585
R12274 GND.n6149 GND.n6148 585
R12275 GND.n6150 GND.n6149 585
R12276 GND.n1540 GND.n1539 585
R12277 GND.n1539 GND.n1535 585
R12278 GND.n6144 GND.n6143 585
R12279 GND.n6143 GND.n6142 585
R12280 GND.n1543 GND.n1542 585
R12281 GND.n5623 GND.n1543 585
R12282 GND.n6124 GND.n6123 585
R12283 GND.n6125 GND.n6124 585
R12284 GND.n1557 GND.n1556 585
R12285 GND.n5598 GND.n1556 585
R12286 GND.n6119 GND.n6118 585
R12287 GND.n6118 GND.n6117 585
R12288 GND.n1560 GND.n1559 585
R12289 GND.n5200 GND.n1560 585
R12290 GND.n6108 GND.n6107 585
R12291 GND.n6109 GND.n6108 585
R12292 GND.n1571 GND.n1570 585
R12293 GND.n1584 GND.n1570 585
R12294 GND.n6103 GND.n6102 585
R12295 GND.n6102 GND.n6101 585
R12296 GND.n1574 GND.n1573 585
R12297 GND.n5650 GND.n1574 585
R12298 GND.n5655 GND.n5654 585
R12299 GND.n5656 GND.n5655 585
R12300 GND.n5182 GND.n5181 585
R12301 GND.n5185 GND.n5182 585
R12302 GND.n5666 GND.n5665 585
R12303 GND.n5665 GND.n5664 585
R12304 GND.n5667 GND.n5176 585
R12305 GND.n5549 GND.n5176 585
R12306 GND.n5669 GND.n5668 585
R12307 GND.n5670 GND.n5669 585
R12308 GND.n5164 GND.n5163 585
R12309 GND.n5167 GND.n5164 585
R12310 GND.n5680 GND.n5679 585
R12311 GND.n5679 GND.n5678 585
R12312 GND.n5681 GND.n5158 585
R12313 GND.n5536 GND.n5158 585
R12314 GND.n5683 GND.n5682 585
R12315 GND.n5684 GND.n5683 585
R12316 GND.n5146 GND.n5145 585
R12317 GND.n5154 GND.n5146 585
R12318 GND.n5694 GND.n5693 585
R12319 GND.n5693 GND.n5692 585
R12320 GND.n5695 GND.n5138 585
R12321 GND.n5521 GND.n5138 585
R12322 GND.n5697 GND.n5696 585
R12323 GND.n5698 GND.n5697 585
R12324 GND.n5139 GND.n5137 585
R12325 GND.n5137 GND.n5133 585
R12326 GND.n5124 GND.n5123 585
R12327 GND.n5127 GND.n5124 585
R12328 GND.n5709 GND.n5708 585
R12329 GND.n5708 GND.n5707 585
R12330 GND.n5710 GND.n5118 585
R12331 GND.n5506 GND.n5118 585
R12332 GND.n5712 GND.n5711 585
R12333 GND.n5713 GND.n5712 585
R12334 GND.n5106 GND.n5105 585
R12335 GND.n5109 GND.n5106 585
R12336 GND.n5723 GND.n5722 585
R12337 GND.n5722 GND.n5721 585
R12338 GND.n5724 GND.n5100 585
R12339 GND.n5493 GND.n5100 585
R12340 GND.n5726 GND.n5725 585
R12341 GND.n5727 GND.n5726 585
R12342 GND.n5088 GND.n5087 585
R12343 GND.n5091 GND.n5088 585
R12344 GND.n5737 GND.n5736 585
R12345 GND.n5736 GND.n5735 585
R12346 GND.n5738 GND.n5082 585
R12347 GND.n5480 GND.n5082 585
R12348 GND.n5740 GND.n5739 585
R12349 GND.n5741 GND.n5740 585
R12350 GND.n5071 GND.n5070 585
R12351 GND.n5074 GND.n5071 585
R12352 GND.n5751 GND.n5750 585
R12353 GND.n5750 GND.n5749 585
R12354 GND.n5752 GND.n5063 585
R12355 GND.n5464 GND.n5063 585
R12356 GND.n5754 GND.n5753 585
R12357 GND.n5755 GND.n5754 585
R12358 GND.n5064 GND.n5062 585
R12359 GND.n5062 GND.n5058 585
R12360 GND.n5049 GND.n5048 585
R12361 GND.n5052 GND.n5049 585
R12362 GND.n5766 GND.n5765 585
R12363 GND.n5765 GND.n5764 585
R12364 GND.n5767 GND.n5043 585
R12365 GND.n5449 GND.n5043 585
R12366 GND.n5769 GND.n5768 585
R12367 GND.n5770 GND.n5769 585
R12368 GND.n5031 GND.n5030 585
R12369 GND.n5034 GND.n5031 585
R12370 GND.n5780 GND.n5779 585
R12371 GND.n5779 GND.n5778 585
R12372 GND.n5781 GND.n5025 585
R12373 GND.n5436 GND.n5025 585
R12374 GND.n5783 GND.n5782 585
R12375 GND.n5784 GND.n5783 585
R12376 GND.n5013 GND.n5012 585
R12377 GND.n5016 GND.n5013 585
R12378 GND.n5794 GND.n5793 585
R12379 GND.n5793 GND.n5792 585
R12380 GND.n5795 GND.n5007 585
R12381 GND.n5423 GND.n5007 585
R12382 GND.n5797 GND.n5796 585
R12383 GND.n5798 GND.n5797 585
R12384 GND.n4996 GND.n4995 585
R12385 GND.n4999 GND.n4996 585
R12386 GND.n5808 GND.n5807 585
R12387 GND.n5807 GND.n5806 585
R12388 GND.n5809 GND.n4990 585
R12389 GND.n5409 GND.n4990 585
R12390 GND.n5811 GND.n5810 585
R12391 GND.n5812 GND.n5811 585
R12392 GND.n4978 GND.n4977 585
R12393 GND.n4981 GND.n4978 585
R12394 GND.n5822 GND.n5821 585
R12395 GND.n5821 GND.n5820 585
R12396 GND.n5823 GND.n4972 585
R12397 GND.n5396 GND.n4972 585
R12398 GND.n5825 GND.n5824 585
R12399 GND.n5826 GND.n5825 585
R12400 GND.n4960 GND.n4959 585
R12401 GND.n4969 GND.n4960 585
R12402 GND.n5836 GND.n5835 585
R12403 GND.n5835 GND.n5834 585
R12404 GND.n5837 GND.n4954 585
R12405 GND.n4961 GND.n4954 585
R12406 GND.n5839 GND.n5838 585
R12407 GND.n5840 GND.n5839 585
R12408 GND.n4951 GND.n4950 585
R12409 GND.n5841 GND.n4951 585
R12410 GND.n5844 GND.n5843 585
R12411 GND.n5843 GND.n5842 585
R12412 GND.n5845 GND.n4945 585
R12413 GND.n4952 GND.n4945 585
R12414 GND.n5847 GND.n5846 585
R12415 GND.n5847 GND.n1643 585
R12416 GND.n5848 GND.n4944 585
R12417 GND.n5848 GND.n1613 585
R12418 GND.n5850 GND.n5849 585
R12419 GND.n5849 GND.n1610 585
R12420 GND.n5851 GND.n4939 585
R12421 GND.n4939 GND.n1607 585
R12422 GND.n5853 GND.n5852 585
R12423 GND.n5853 GND.n1676 585
R12424 GND.n5854 GND.n4938 585
R12425 GND.n5854 GND.n1684 585
R12426 GND.n5856 GND.n5855 585
R12427 GND.n5855 GND.n1682 585
R12428 GND.n5857 GND.n1705 585
R12429 GND.n1705 GND.n1693 585
R12430 GND.n5859 GND.n5858 585
R12431 GND.n5860 GND.n5859 585
R12432 GND.n1706 GND.n1704 585
R12433 GND.n1704 GND.n1702 585
R12434 GND.n4932 GND.n4931 585
R12435 GND.n4931 GND.n4930 585
R12436 GND.n1709 GND.n1708 585
R12437 GND.n1721 GND.n1709 585
R12438 GND.n4818 GND.n4817 585
R12439 GND.n4818 GND.n1718 585
R12440 GND.n4819 GND.n4814 585
R12441 GND.n4819 GND.n1732 585
R12442 GND.n4821 GND.n4820 585
R12443 GND.n4820 GND.n1740 585
R12444 GND.n4822 GND.n4809 585
R12445 GND.n4809 GND.n1738 585
R12446 GND.n4824 GND.n4823 585
R12447 GND.n4824 GND.n1751 585
R12448 GND.n4825 GND.n4808 585
R12449 GND.n4825 GND.n1748 585
R12450 GND.n4827 GND.n4826 585
R12451 GND.n4826 GND.n1760 585
R12452 GND.n4828 GND.n1787 585
R12453 GND.n1787 GND.n1767 585
R12454 GND.n4830 GND.n4829 585
R12455 GND.n4831 GND.n4830 585
R12456 GND.n1788 GND.n1786 585
R12457 GND.n1786 GND.n1778 585
R12458 GND.n4802 GND.n4801 585
R12459 GND.n4801 GND.n1775 585
R12460 GND.n4800 GND.n1790 585
R12461 GND.n4800 GND.n4799 585
R12462 GND.n4719 GND.n1791 585
R12463 GND.n1801 GND.n1791 585
R12464 GND.n4721 GND.n4720 585
R12465 GND.n4721 GND.n1799 585
R12466 GND.n4722 GND.n4715 585
R12467 GND.n4722 GND.n1812 585
R12468 GND.n4724 GND.n4723 585
R12469 GND.n4723 GND.n1809 585
R12470 GND.n4725 GND.n1851 585
R12471 GND.n1851 GND.n1821 585
R12472 GND.n4727 GND.n4726 585
R12473 GND.n4728 GND.n4727 585
R12474 GND.n1852 GND.n1850 585
R12475 GND.n1850 GND.n1827 585
R12476 GND.n4709 GND.n4708 585
R12477 GND.n4708 GND.n1839 585
R12478 GND.n4707 GND.n1854 585
R12479 GND.n4707 GND.n1836 585
R12480 GND.n4706 GND.n1856 585
R12481 GND.n4706 GND.n4705 585
R12482 GND.n4543 GND.n1855 585
R12483 GND.n1866 GND.n1855 585
R12484 GND.n4545 GND.n4541 585
R12485 GND.n4541 GND.n1864 585
R12486 GND.n4547 GND.n4546 585
R12487 GND.n4547 GND.n1909 585
R12488 GND.n4548 GND.n4540 585
R12489 GND.n4548 GND.n1911 585
R12490 GND.n4550 GND.n4549 585
R12491 GND.n4549 GND.n1914 585
R12492 GND.n4552 GND.n4538 585
R12493 GND.n4538 GND.n1921 585
R12494 GND.n4554 GND.n4553 585
R12495 GND.n4554 GND.n1920 585
R12496 GND.n4555 GND.n4537 585
R12497 GND.n4555 GND.n1928 585
R12498 GND.n4557 GND.n4556 585
R12499 GND.n4556 GND.n1930 585
R12500 GND.n4559 GND.n4536 585
R12501 GND.n4536 GND.n1885 585
R12502 GND.n4560 GND.n4532 585
R12503 GND.n4532 GND.n1882 585
R12504 GND.n4562 GND.n4561 585
R12505 GND.n4562 GND.n1937 585
R12506 GND.n4563 GND.n4531 585
R12507 GND.n4563 GND.n1940 585
R12508 GND.n4565 GND.n4564 585
R12509 GND.n4564 GND.n1950 585
R12510 GND.n4566 GND.n1992 585
R12511 GND.n1992 GND.n1947 585
R12512 GND.n4568 GND.n4567 585
R12513 GND.n4569 GND.n4568 585
R12514 GND.n1993 GND.n1991 585
R12515 GND.n1991 GND.n1969 585
R12516 GND.n4525 GND.n4524 585
R12517 GND.n4524 GND.n1967 585
R12518 GND.n4523 GND.n1995 585
R12519 GND.n4523 GND.n1980 585
R12520 GND.n4522 GND.n4521 585
R12521 GND.n4522 GND.n1977 585
R12522 GND.n1997 GND.n1996 585
R12523 GND.n2004 GND.n1996 585
R12524 GND.n4517 GND.n4516 585
R12525 GND.n4516 GND.n4515 585
R12526 GND.n2000 GND.n1999 585
R12527 GND.n2014 GND.n2000 585
R12528 GND.n4448 GND.n2054 585
R12529 GND.n2054 GND.n2011 585
R12530 GND.n4450 GND.n4449 585
R12531 GND.n4451 GND.n4450 585
R12532 GND.n2055 GND.n2053 585
R12533 GND.n2053 GND.n2031 585
R12534 GND.n4443 GND.n4442 585
R12535 GND.n4442 GND.n2029 585
R12536 GND.n4441 GND.n2057 585
R12537 GND.n4441 GND.n2042 585
R12538 GND.n4440 GND.n4439 585
R12539 GND.n4440 GND.n2039 585
R12540 GND.n2059 GND.n2058 585
R12541 GND.n2066 GND.n2058 585
R12542 GND.n4435 GND.n4434 585
R12543 GND.n4434 GND.n4433 585
R12544 GND.n2062 GND.n2061 585
R12545 GND.n2076 GND.n2062 585
R12546 GND.n4108 GND.n4107 585
R12547 GND.n4108 GND.n2073 585
R12548 GND.n4110 GND.n4109 585
R12549 GND.n4109 GND.n2085 585
R12550 GND.n4111 GND.n4101 585
R12551 GND.n4101 GND.n2094 585
R12552 GND.n4113 GND.n4112 585
R12553 GND.n4113 GND.n2092 585
R12554 GND.n4114 GND.n4100 585
R12555 GND.n4114 GND.n2105 585
R12556 GND.n4116 GND.n4115 585
R12557 GND.n4115 GND.n2102 585
R12558 GND.n4117 GND.n4095 585
R12559 GND.n4095 GND.n2114 585
R12560 GND.n4119 GND.n4118 585
R12561 GND.n4119 GND.n2123 585
R12562 GND.n4120 GND.n4094 585
R12563 GND.n4120 GND.n2121 585
R12564 GND.n4122 GND.n4121 585
R12565 GND.n4121 GND.n2133 585
R12566 GND.n4123 GND.n2154 585
R12567 GND.n2154 GND.n2130 585
R12568 GND.n6045 GND.n1603 585
R12569 GND.n6046 GND.n6045 585
R12570 GND.n5871 GND.n1611 585
R12571 GND.n5899 GND.n1611 585
R12572 GND.n5872 GND.n5870 585
R12573 GND.n5870 GND.n5869 585
R12574 GND.n5867 GND.n1685 585
R12575 GND.n5890 GND.n1685 585
R12576 GND.n1697 GND.n1695 585
R12577 GND.n5864 GND.n1695 585
R12578 GND.n5880 GND.n5879 585
R12579 GND.n5881 GND.n5880 585
R12580 GND.n1696 GND.n1694 585
R12581 GND.n5861 GND.n1694 585
R12582 GND.n1727 GND.n1712 585
R12583 GND.n4929 GND.n1712 585
R12584 GND.n1725 GND.n1723 585
R12585 GND.n1723 GND.n1710 585
R12586 GND.n4920 GND.n4919 585
R12587 GND.n4921 GND.n4920 585
R12588 GND.n1724 GND.n1722 585
R12589 GND.n4912 GND.n1722 585
R12590 GND.n4874 GND.n4873 585
R12591 GND.n4873 GND.n4872 585
R12592 GND.n4871 GND.n1741 585
R12593 GND.n4893 GND.n1741 585
R12594 GND.n1755 GND.n1753 585
R12595 GND.n4869 GND.n1753 585
R12596 GND.n4882 GND.n4881 585
R12597 GND.n4883 GND.n4882 585
R12598 GND.n1754 GND.n1752 585
R12599 GND.n4866 GND.n1752 585
R12600 GND.n4837 GND.n4836 585
R12601 GND.n4836 GND.n4835 585
R12602 GND.n4834 GND.n1768 585
R12603 GND.n4856 GND.n1768 585
R12604 GND.n1782 GND.n1780 585
R12605 GND.n4832 GND.n1780 585
R12606 GND.n4845 GND.n4844 585
R12607 GND.n4846 GND.n4845 585
R12608 GND.n1781 GND.n1779 585
R12609 GND.n4798 GND.n1779 585
R12610 GND.n4769 GND.n4768 585
R12611 GND.n4768 GND.n1792 585
R12612 GND.n4767 GND.n1802 585
R12613 GND.n4788 GND.n1802 585
R12614 GND.n1816 GND.n1814 585
R12615 GND.n4763 GND.n1814 585
R12616 GND.n4777 GND.n4776 585
R12617 GND.n4778 GND.n4777 585
R12618 GND.n1815 GND.n1813 585
R12619 GND.n4760 GND.n1813 585
R12620 GND.n4731 GND.n4730 585
R12621 GND.n4730 GND.n4729 585
R12622 GND.n1849 GND.n1829 585
R12623 GND.n4750 GND.n1829 585
R12624 GND.n1843 GND.n1841 585
R12625 GND.n1847 GND.n1841 585
R12626 GND.n4739 GND.n4738 585
R12627 GND.n4740 GND.n4739 585
R12628 GND.n1842 GND.n1840 585
R12629 GND.n4704 GND.n1840 585
R12630 GND.n4665 GND.n4664 585
R12631 GND.n4664 GND.n1857 585
R12632 GND.n4663 GND.n1867 585
R12633 GND.n4694 GND.n1867 585
R12634 GND.n4659 GND.n1906 585
R12635 GND.n4660 GND.n4659 585
R12636 GND.n4658 GND.n1905 585
R12637 GND.n4658 GND.n4657 585
R12638 GND.n1910 GND.n1904 585
R12639 GND.n4652 GND.n1910 585
R12640 GND.n1924 GND.n1922 585
R12641 GND.n1924 GND.n1923 585
R12642 GND.n1925 GND.n1898 585
R12643 GND.n4641 GND.n1925 585
R12644 GND.n4635 GND.n1897 585
R12645 GND.n4636 GND.n4635 585
R12646 GND.n4634 GND.n1896 585
R12647 GND.n4634 GND.n4633 585
R12648 GND.n1889 GND.n1887 585
R12649 GND.n1931 GND.n1887 585
R12650 GND.n4684 GND.n4683 585
R12651 GND.n4685 GND.n4684 585
R12652 GND.n1888 GND.n1886 585
R12653 GND.n4624 GND.n1886 585
R12654 GND.n1956 GND.n1941 585
R12655 GND.n4621 GND.n1941 585
R12656 GND.n1954 GND.n1952 585
R12657 GND.n4597 GND.n1952 585
R12658 GND.n4612 GND.n4611 585
R12659 GND.n4613 GND.n4612 585
R12660 GND.n1953 GND.n1951 585
R12661 GND.n4605 GND.n1951 585
R12662 GND.n4572 GND.n4571 585
R12663 GND.n4571 GND.n4570 585
R12664 GND.n1990 GND.n1970 585
R12665 GND.n4591 GND.n1970 585
R12666 GND.n1984 GND.n1982 585
R12667 GND.n1988 GND.n1982 585
R12668 GND.n4580 GND.n4579 585
R12669 GND.n4581 GND.n4580 585
R12670 GND.n1983 GND.n1981 585
R12671 GND.n4481 GND.n1981 585
R12672 GND.n4498 GND.n2005 585
R12673 GND.n4514 GND.n2005 585
R12674 GND.n2018 GND.n2016 585
R12675 GND.n2016 GND.n2001 585
R12676 GND.n4505 GND.n4504 585
R12677 GND.n4506 GND.n4505 585
R12678 GND.n2017 GND.n2015 585
R12679 GND.n4494 GND.n2015 585
R12680 GND.n4454 GND.n4453 585
R12681 GND.n4453 GND.n4452 585
R12682 GND.n2052 GND.n2032 585
R12683 GND.n4473 GND.n2032 585
R12684 GND.n2046 GND.n2044 585
R12685 GND.n2050 GND.n2044 585
R12686 GND.n4462 GND.n4461 585
R12687 GND.n4463 GND.n4462 585
R12688 GND.n2045 GND.n2043 585
R12689 GND.n4399 GND.n2043 585
R12690 GND.n4416 GND.n2067 585
R12691 GND.n4432 GND.n2067 585
R12692 GND.n2080 GND.n2078 585
R12693 GND.n2078 GND.n2063 585
R12694 GND.n4423 GND.n4422 585
R12695 GND.n4424 GND.n4423 585
R12696 GND.n2079 GND.n2077 585
R12697 GND.n4412 GND.n2077 585
R12698 GND.n4372 GND.n4371 585
R12699 GND.n4371 GND.n4370 585
R12700 GND.n4369 GND.n2095 585
R12701 GND.n4391 GND.n2095 585
R12702 GND.n2109 GND.n2107 585
R12703 GND.n4367 GND.n2107 585
R12704 GND.n4380 GND.n4379 585
R12705 GND.n4381 GND.n4380 585
R12706 GND.n2108 GND.n2106 585
R12707 GND.n4364 GND.n2106 585
R12708 GND.n4336 GND.n4335 585
R12709 GND.n4335 GND.n4334 585
R12710 GND.n4333 GND.n2124 585
R12711 GND.n4355 GND.n2124 585
R12712 GND.n2136 GND.n2135 585
R12713 GND.n4331 GND.n2135 585
R12714 GND.n4344 GND.n4343 585
R12715 GND.n4345 GND.n4344 585
R12716 GND.n4327 GND.n2134 585
R12717 GND.n4326 GND.n2139 585
R12718 GND.n4325 GND.n2140 585
R12719 GND.n4153 GND.n2141 585
R12720 GND.n4321 GND.n2143 585
R12721 GND.n4320 GND.n2144 585
R12722 GND.n4319 GND.n2145 585
R12723 GND.n2151 GND.n2148 585
R12724 GND.n4315 GND.n4314 585
R12725 GND.n4314 GND.n4313 585
R12726 GND.n5896 GND.n1609 585
R12727 GND.n6046 GND.n1609 585
R12728 GND.n5898 GND.n5897 585
R12729 GND.n5899 GND.n5898 585
R12730 GND.n1678 GND.n1677 585
R12731 GND.n5869 GND.n1677 585
R12732 GND.n5892 GND.n5891 585
R12733 GND.n5891 GND.n5890 585
R12734 GND.n1681 GND.n1680 585
R12735 GND.n5864 GND.n1681 585
R12736 GND.n4904 GND.n1692 585
R12737 GND.n5881 GND.n1692 585
R12738 GND.n4905 GND.n1703 585
R12739 GND.n5861 GND.n1703 585
R12740 GND.n4906 GND.n1711 585
R12741 GND.n4929 GND.n1711 585
R12742 GND.n4908 GND.n4907 585
R12743 GND.n4907 GND.n1710 585
R12744 GND.n4909 GND.n1720 585
R12745 GND.n4921 GND.n1720 585
R12746 GND.n4911 GND.n4910 585
R12747 GND.n4912 GND.n4911 585
R12748 GND.n1734 GND.n1733 585
R12749 GND.n4872 GND.n1733 585
R12750 GND.n4895 GND.n4894 585
R12751 GND.n4894 GND.n4893 585
R12752 GND.n1737 GND.n1736 585
R12753 GND.n4869 GND.n1737 585
R12754 GND.n4863 GND.n1750 585
R12755 GND.n4883 GND.n1750 585
R12756 GND.n4865 GND.n4864 585
R12757 GND.n4866 GND.n4865 585
R12758 GND.n1762 GND.n1761 585
R12759 GND.n4835 GND.n1761 585
R12760 GND.n4858 GND.n4857 585
R12761 GND.n4857 GND.n4856 585
R12762 GND.n1765 GND.n1764 585
R12763 GND.n4832 GND.n1765 585
R12764 GND.n4795 GND.n1777 585
R12765 GND.n4846 GND.n1777 585
R12766 GND.n4797 GND.n4796 585
R12767 GND.n4798 GND.n4797 585
R12768 GND.n1795 GND.n1794 585
R12769 GND.n1794 GND.n1792 585
R12770 GND.n4790 GND.n4789 585
R12771 GND.n4789 GND.n4788 585
R12772 GND.n1798 GND.n1797 585
R12773 GND.n4763 GND.n1798 585
R12774 GND.n4757 GND.n1811 585
R12775 GND.n4778 GND.n1811 585
R12776 GND.n4759 GND.n4758 585
R12777 GND.n4760 GND.n4759 585
R12778 GND.n1823 GND.n1822 585
R12779 GND.n4729 GND.n1822 585
R12780 GND.n4752 GND.n4751 585
R12781 GND.n4751 GND.n4750 585
R12782 GND.n1826 GND.n1825 585
R12783 GND.n1847 GND.n1826 585
R12784 GND.n4701 GND.n1838 585
R12785 GND.n4740 GND.n1838 585
R12786 GND.n4703 GND.n4702 585
R12787 GND.n4704 GND.n4703 585
R12788 GND.n1860 GND.n1859 585
R12789 GND.n1859 GND.n1857 585
R12790 GND.n4696 GND.n4695 585
R12791 GND.n4695 GND.n4694 585
R12792 GND.n1863 GND.n1862 585
R12793 GND.n4660 GND.n1863 585
R12794 GND.n4649 GND.n1912 585
R12795 GND.n4657 GND.n1912 585
R12796 GND.n4651 GND.n4650 585
R12797 GND.n4652 GND.n4651 585
R12798 GND.n1916 GND.n1915 585
R12799 GND.n1923 GND.n1915 585
R12800 GND.n4643 GND.n4642 585
R12801 GND.n4642 GND.n4641 585
R12802 GND.n1919 GND.n1918 585
R12803 GND.n4636 GND.n1919 585
R12804 GND.n4632 GND.n4631 585
R12805 GND.n4633 GND.n4632 585
R12806 GND.n1933 GND.n1932 585
R12807 GND.n1932 GND.n1931 585
R12808 GND.n4627 GND.n1884 585
R12809 GND.n4685 GND.n1884 585
R12810 GND.n4626 GND.n4625 585
R12811 GND.n4625 GND.n4624 585
R12812 GND.n1936 GND.n1935 585
R12813 GND.n4621 GND.n1936 585
R12814 GND.n4599 GND.n4598 585
R12815 GND.n4598 GND.n4597 585
R12816 GND.n1963 GND.n1949 585
R12817 GND.n4613 GND.n1949 585
R12818 GND.n4604 GND.n4603 585
R12819 GND.n4605 GND.n4604 585
R12820 GND.n1962 GND.n1961 585
R12821 GND.n4570 GND.n1961 585
R12822 GND.n4593 GND.n4592 585
R12823 GND.n4592 GND.n4591 585
R12824 GND.n1966 GND.n1965 585
R12825 GND.n1988 GND.n1966 585
R12826 GND.n4483 GND.n1979 585
R12827 GND.n4581 GND.n1979 585
R12828 GND.n4486 GND.n4482 585
R12829 GND.n4482 GND.n4481 585
R12830 GND.n4487 GND.n2003 585
R12831 GND.n4514 GND.n2003 585
R12832 GND.n4488 GND.n4479 585
R12833 GND.n4479 GND.n2001 585
R12834 GND.n2025 GND.n2013 585
R12835 GND.n4506 GND.n2013 585
R12836 GND.n4493 GND.n4492 585
R12837 GND.n4494 GND.n4493 585
R12838 GND.n2024 GND.n2023 585
R12839 GND.n4452 GND.n2023 585
R12840 GND.n4475 GND.n4474 585
R12841 GND.n4474 GND.n4473 585
R12842 GND.n2028 GND.n2027 585
R12843 GND.n2050 GND.n2028 585
R12844 GND.n4401 GND.n2041 585
R12845 GND.n4463 GND.n2041 585
R12846 GND.n4404 GND.n4400 585
R12847 GND.n4400 GND.n4399 585
R12848 GND.n4405 GND.n2065 585
R12849 GND.n4432 GND.n2065 585
R12850 GND.n4406 GND.n4397 585
R12851 GND.n4397 GND.n2063 585
R12852 GND.n2088 GND.n2075 585
R12853 GND.n4424 GND.n2075 585
R12854 GND.n4411 GND.n4410 585
R12855 GND.n4412 GND.n4411 585
R12856 GND.n2087 GND.n2086 585
R12857 GND.n4370 GND.n2086 585
R12858 GND.n4393 GND.n4392 585
R12859 GND.n4392 GND.n4391 585
R12860 GND.n2091 GND.n2090 585
R12861 GND.n4367 GND.n2091 585
R12862 GND.n2117 GND.n2104 585
R12863 GND.n4381 GND.n2104 585
R12864 GND.n4363 GND.n4362 585
R12865 GND.n4364 GND.n4363 585
R12866 GND.n2116 GND.n2115 585
R12867 GND.n4334 GND.n2115 585
R12868 GND.n4357 GND.n4356 585
R12869 GND.n4356 GND.n4355 585
R12870 GND.n2120 GND.n2119 585
R12871 GND.n4331 GND.n2120 585
R12872 GND.n2149 GND.n2132 585
R12873 GND.n4345 GND.n2132 585
R12874 GND.n6042 GND.n1642 585
R12875 GND.n1641 GND.n1640 585
R12876 GND.n1636 GND.n1599 585
R12877 GND.n1635 GND.n1634 585
R12878 GND.n1632 GND.n1631 585
R12879 GND.n1630 GND.n1629 585
R12880 GND.n1627 GND.n1626 585
R12881 GND.n1625 GND.n1612 585
R12882 GND.n7592 GND.n765 521.33
R12883 GND.n7426 GND.n7424 521.33
R12884 GND.n5387 GND.n5386 521.33
R12885 GND.n5278 GND.n4964 521.33
R12886 GND.n3215 GND.n3214 422.007
R12887 GND.n8265 GND.n381 393.24
R12888 GND.n3214 GND.n2966 301.784
R12889 GND.n2975 GND.n2966 301.784
R12890 GND.n3205 GND.n2975 301.784
R12891 GND.n3205 GND.n3204 301.784
R12892 GND.n3204 GND.n3203 301.784
R12893 GND.n3203 GND.n2976 301.784
R12894 GND.n3197 GND.n2976 301.784
R12895 GND.n3197 GND.n3196 301.784
R12896 GND.n3196 GND.n3195 301.784
R12897 GND.n3195 GND.n2983 301.784
R12898 GND.n3189 GND.n2983 301.784
R12899 GND.n3189 GND.n3188 301.784
R12900 GND.n3188 GND.n3187 301.784
R12901 GND.n3187 GND.n2991 301.784
R12902 GND.n3181 GND.n2991 301.784
R12903 GND.n3181 GND.n3180 301.784
R12904 GND.n3180 GND.n3179 301.784
R12905 GND.n3179 GND.n2999 301.784
R12906 GND.n3173 GND.n2999 301.784
R12907 GND.n3173 GND.n3172 301.784
R12908 GND.n3172 GND.n3171 301.784
R12909 GND.n3171 GND.n3007 301.784
R12910 GND.n3165 GND.n3007 301.784
R12911 GND.n3165 GND.n3164 301.784
R12912 GND.n3164 GND.n3163 301.784
R12913 GND.n3163 GND.n3015 301.784
R12914 GND.n3157 GND.n3015 301.784
R12915 GND.n3157 GND.n3156 301.784
R12916 GND.n3156 GND.n3155 301.784
R12917 GND.n3155 GND.n3023 301.784
R12918 GND.n3149 GND.n3023 301.784
R12919 GND.n3149 GND.n3148 301.784
R12920 GND.n3148 GND.n3147 301.784
R12921 GND.n3147 GND.n3031 301.784
R12922 GND.n3141 GND.n3031 301.784
R12923 GND.n3141 GND.n3140 301.784
R12924 GND.n3140 GND.n3139 301.784
R12925 GND.n3139 GND.n3039 301.784
R12926 GND.n3133 GND.n3039 301.784
R12927 GND.n3133 GND.n3132 301.784
R12928 GND.n3132 GND.n3131 301.784
R12929 GND.n3131 GND.n3047 301.784
R12930 GND.n3125 GND.n3047 301.784
R12931 GND.n3125 GND.n3124 301.784
R12932 GND.n3124 GND.n3123 301.784
R12933 GND.n3123 GND.n3055 301.784
R12934 GND.n3117 GND.n3055 301.784
R12935 GND.n3117 GND.n3116 301.784
R12936 GND.n3116 GND.n3115 301.784
R12937 GND.n3115 GND.n3063 301.784
R12938 GND.n3109 GND.n3063 301.784
R12939 GND.n3109 GND.n3108 301.784
R12940 GND.n3108 GND.n3107 301.784
R12941 GND.n3107 GND.n3071 301.784
R12942 GND.n3101 GND.n3071 301.784
R12943 GND.n3101 GND.n3100 301.784
R12944 GND.n3100 GND.n3099 301.784
R12945 GND.n3099 GND.n3079 301.784
R12946 GND.n3093 GND.n3079 301.784
R12947 GND.n3093 GND.n3092 301.784
R12948 GND.n3092 GND.n3091 301.784
R12949 GND.n3091 GND.n381 301.784
R12950 GND.n13 GND.n11 289.615
R12951 GND.n24 GND.n22 289.615
R12952 GND.n36 GND.n34 289.615
R12953 GND.n48 GND.n46 289.615
R12954 GND.n60 GND.n58 289.615
R12955 GND.n2 GND.n0 289.615
R12956 GND.n86 GND.n84 289.615
R12957 GND.n97 GND.n95 289.615
R12958 GND.n109 GND.n107 289.615
R12959 GND.n121 GND.n119 289.615
R12960 GND.n133 GND.n131 289.615
R12961 GND.n145 GND.n143 289.615
R12962 GND.n5254 GND.t119 260.649
R12963 GND.n786 GND.t141 260.649
R12964 GND.n5279 GND.n4953 256.663
R12965 GND.n5282 GND.n4953 256.663
R12966 GND.n5288 GND.n4953 256.663
R12967 GND.n5290 GND.n4953 256.663
R12968 GND.n5296 GND.n4953 256.663
R12969 GND.n5298 GND.n4953 256.663
R12970 GND.n5304 GND.n4953 256.663
R12971 GND.n5306 GND.n4953 256.663
R12972 GND.n5312 GND.n4953 256.663
R12973 GND.n5314 GND.n4953 256.663
R12974 GND.n5323 GND.n4953 256.663
R12975 GND.n5325 GND.n4953 256.663
R12976 GND.n5331 GND.n4953 256.663
R12977 GND.n5332 GND.n5232 256.663
R12978 GND.n5333 GND.n4953 256.663
R12979 GND.n5335 GND.n4953 256.663
R12980 GND.n5344 GND.n4953 256.663
R12981 GND.n5346 GND.n4953 256.663
R12982 GND.n5352 GND.n4953 256.663
R12983 GND.n5354 GND.n4953 256.663
R12984 GND.n5360 GND.n4953 256.663
R12985 GND.n5362 GND.n4953 256.663
R12986 GND.n5368 GND.n4953 256.663
R12987 GND.n5370 GND.n4953 256.663
R12988 GND.n5376 GND.n4953 256.663
R12989 GND.n5378 GND.n4953 256.663
R12990 GND.n5384 GND.n4953 256.663
R12991 GND.n7593 GND.n752 256.663
R12992 GND.n7593 GND.n751 256.663
R12993 GND.n7593 GND.n750 256.663
R12994 GND.n7593 GND.n749 256.663
R12995 GND.n7593 GND.n748 256.663
R12996 GND.n7593 GND.n747 256.663
R12997 GND.n7593 GND.n746 256.663
R12998 GND.n7593 GND.n745 256.663
R12999 GND.n7593 GND.n744 256.663
R13000 GND.n7593 GND.n743 256.663
R13001 GND.n7593 GND.n742 256.663
R13002 GND.n7593 GND.n741 256.663
R13003 GND.n7593 GND.n740 256.663
R13004 GND.n7596 GND.n7595 256.663
R13005 GND.n7593 GND.n737 256.663
R13006 GND.n7593 GND.n753 256.663
R13007 GND.n7593 GND.n754 256.663
R13008 GND.n7593 GND.n755 256.663
R13009 GND.n7593 GND.n756 256.663
R13010 GND.n7593 GND.n757 256.663
R13011 GND.n7593 GND.n758 256.663
R13012 GND.n7593 GND.n759 256.663
R13013 GND.n7593 GND.n760 256.663
R13014 GND.n7593 GND.n761 256.663
R13015 GND.n7593 GND.n762 256.663
R13016 GND.n7593 GND.n763 256.663
R13017 GND.n7593 GND.n764 256.663
R13018 GND.n7725 GND.n696 242.672
R13019 GND.n7725 GND.n701 242.672
R13020 GND.n7725 GND.n705 242.672
R13021 GND.n7726 GND.n7725 242.672
R13022 GND.n8448 GND.n8447 242.672
R13023 GND.n8447 GND.n380 242.672
R13024 GND.n8447 GND.n359 242.672
R13025 GND.n8447 GND.n358 242.672
R13026 GND.n6100 GND.n6099 242.672
R13027 GND.n6100 GND.n1576 242.672
R13028 GND.n6100 GND.n1577 242.672
R13029 GND.n6100 GND.n1578 242.672
R13030 GND.n6100 GND.n1579 242.672
R13031 GND.n6100 GND.n1580 242.672
R13032 GND.n6100 GND.n1581 242.672
R13033 GND.n6100 GND.n1582 242.672
R13034 GND.n6100 GND.n1583 242.672
R13035 GND.n1066 GND.n1031 242.672
R13036 GND.n6962 GND.n1031 242.672
R13037 GND.n1069 GND.n1031 242.672
R13038 GND.n6951 GND.n1031 242.672
R13039 GND.n6943 GND.n1031 242.672
R13040 GND.n6941 GND.n1031 242.672
R13041 GND.n6933 GND.n1031 242.672
R13042 GND.n6931 GND.n1031 242.672
R13043 GND.n6922 GND.n1031 242.672
R13044 GND.n6920 GND.n1031 242.672
R13045 GND.n4313 GND.n4312 242.672
R13046 GND.n4313 GND.n4129 242.672
R13047 GND.n4313 GND.n4130 242.672
R13048 GND.n4313 GND.n4131 242.672
R13049 GND.n4313 GND.n4132 242.672
R13050 GND.n4313 GND.n4133 242.672
R13051 GND.n4313 GND.n4134 242.672
R13052 GND.n4313 GND.n4135 242.672
R13053 GND.n4313 GND.n4136 242.672
R13054 GND.n4313 GND.n4137 242.672
R13055 GND.n4313 GND.n4138 242.672
R13056 GND.n4313 GND.n4139 242.672
R13057 GND.n4313 GND.n4140 242.672
R13058 GND.n4313 GND.n4141 242.672
R13059 GND.n4313 GND.n4142 242.672
R13060 GND.n4313 GND.n4143 242.672
R13061 GND.n4313 GND.n4144 242.672
R13062 GND.n4313 GND.n4145 242.672
R13063 GND.n4313 GND.n4146 242.672
R13064 GND.n4313 GND.n4147 242.672
R13065 GND.n4313 GND.n4148 242.672
R13066 GND.n4313 GND.n4149 242.672
R13067 GND.n4313 GND.n4150 242.672
R13068 GND.n4313 GND.n4151 242.672
R13069 GND.n6042 GND.n1644 242.672
R13070 GND.n6042 GND.n1645 242.672
R13071 GND.n6042 GND.n1646 242.672
R13072 GND.n6042 GND.n1647 242.672
R13073 GND.n6042 GND.n1648 242.672
R13074 GND.n6042 GND.n1649 242.672
R13075 GND.n6042 GND.n1650 242.672
R13076 GND.n6042 GND.n1651 242.672
R13077 GND.n6042 GND.n1652 242.672
R13078 GND.n6042 GND.n1653 242.672
R13079 GND.n6042 GND.n1654 242.672
R13080 GND.n6042 GND.n1655 242.672
R13081 GND.n6042 GND.n1656 242.672
R13082 GND.n1658 GND.n1657 242.672
R13083 GND.n6042 GND.n1624 242.672
R13084 GND.n6042 GND.n1623 242.672
R13085 GND.n6042 GND.n1622 242.672
R13086 GND.n6042 GND.n1621 242.672
R13087 GND.n6042 GND.n1620 242.672
R13088 GND.n6042 GND.n1619 242.672
R13089 GND.n6042 GND.n1618 242.672
R13090 GND.n6042 GND.n1617 242.672
R13091 GND.n6042 GND.n1616 242.672
R13092 GND.n6042 GND.n1615 242.672
R13093 GND.n6042 GND.n1614 242.672
R13094 GND.n7725 GND.n7724 242.672
R13095 GND.n7725 GND.n672 242.672
R13096 GND.n7725 GND.n673 242.672
R13097 GND.n7725 GND.n674 242.672
R13098 GND.n7725 GND.n675 242.672
R13099 GND.n7725 GND.n676 242.672
R13100 GND.n7725 GND.n677 242.672
R13101 GND.n7725 GND.n678 242.672
R13102 GND.n7725 GND.n679 242.672
R13103 GND.n7725 GND.n680 242.672
R13104 GND.n7725 GND.n681 242.672
R13105 GND.n7725 GND.n682 242.672
R13106 GND.n7725 GND.n683 242.672
R13107 GND.n7725 GND.n684 242.672
R13108 GND.n7725 GND.n685 242.672
R13109 GND.n7725 GND.n686 242.672
R13110 GND.n7725 GND.n687 242.672
R13111 GND.n7725 GND.n688 242.672
R13112 GND.n7725 GND.n689 242.672
R13113 GND.n7725 GND.n690 242.672
R13114 GND.n7725 GND.n691 242.672
R13115 GND.n7725 GND.n692 242.672
R13116 GND.n7725 GND.n693 242.672
R13117 GND.n7725 GND.n694 242.672
R13118 GND.n8447 GND.n8266 242.672
R13119 GND.n8447 GND.n8267 242.672
R13120 GND.n8447 GND.n8268 242.672
R13121 GND.n8447 GND.n8269 242.672
R13122 GND.n8447 GND.n8270 242.672
R13123 GND.n8447 GND.n8271 242.672
R13124 GND.n8447 GND.n8272 242.672
R13125 GND.n8447 GND.n8273 242.672
R13126 GND.n8447 GND.n8274 242.672
R13127 GND.n8447 GND.n8275 242.672
R13128 GND.n8447 GND.n8276 242.672
R13129 GND.n8447 GND.n8277 242.672
R13130 GND.n8447 GND.n8278 242.672
R13131 GND.n8447 GND.n8279 242.672
R13132 GND.n8447 GND.n8280 242.672
R13133 GND.n8447 GND.n8281 242.672
R13134 GND.n8447 GND.n8282 242.672
R13135 GND.n8447 GND.n8283 242.672
R13136 GND.n8447 GND.n8284 242.672
R13137 GND.n8447 GND.n8285 242.672
R13138 GND.n8447 GND.n8286 242.672
R13139 GND.n8447 GND.n8287 242.672
R13140 GND.n8447 GND.n8288 242.672
R13141 GND.n8447 GND.n8446 242.672
R13142 GND.n4313 GND.n4152 242.672
R13143 GND.n4313 GND.n4154 242.672
R13144 GND.n4313 GND.n4155 242.672
R13145 GND.n4313 GND.n4156 242.672
R13146 GND.n6042 GND.n1637 242.672
R13147 GND.n6042 GND.n1633 242.672
R13148 GND.n6042 GND.n1628 242.672
R13149 GND.n6043 GND.n6042 242.672
R13150 GND.n8289 GND.n342 240.244
R13151 GND.n8445 GND.n8290 240.244
R13152 GND.n8441 GND.n8440 240.244
R13153 GND.n8437 GND.n8436 240.244
R13154 GND.n8305 GND.n8304 240.244
R13155 GND.n8429 GND.n8428 240.244
R13156 GND.n8425 GND.n8424 240.244
R13157 GND.n8421 GND.n8420 240.244
R13158 GND.n8417 GND.n8416 240.244
R13159 GND.n8410 GND.n8409 240.244
R13160 GND.n8406 GND.n8405 240.244
R13161 GND.n8402 GND.n8401 240.244
R13162 GND.n8398 GND.n8397 240.244
R13163 GND.n8394 GND.n8393 240.244
R13164 GND.n8387 GND.n8386 240.244
R13165 GND.n8384 GND.n8383 240.244
R13166 GND.n8380 GND.n8379 240.244
R13167 GND.n8376 GND.n8375 240.244
R13168 GND.n8372 GND.n8371 240.244
R13169 GND.n8365 GND.n8364 240.244
R13170 GND.n8362 GND.n8361 240.244
R13171 GND.n8358 GND.n8357 240.244
R13172 GND.n8354 GND.n8353 240.244
R13173 GND.n8350 GND.n8349 240.244
R13174 GND.n7738 GND.n648 240.244
R13175 GND.n7748 GND.n648 240.244
R13176 GND.n7748 GND.n638 240.244
R13177 GND.n638 GND.n630 240.244
R13178 GND.n7775 GND.n630 240.244
R13179 GND.n7775 GND.n620 240.244
R13180 GND.n7779 GND.n620 240.244
R13181 GND.n7779 GND.n610 240.244
R13182 GND.n610 GND.n602 240.244
R13183 GND.n7816 GND.n602 240.244
R13184 GND.n7816 GND.n593 240.244
R13185 GND.n593 GND.n583 240.244
R13186 GND.n7835 GND.n583 240.244
R13187 GND.n7836 GND.n7835 240.244
R13188 GND.n7836 GND.n571 240.244
R13189 GND.n7847 GND.n571 240.244
R13190 GND.n7847 GND.n559 240.244
R13191 GND.n7868 GND.n559 240.244
R13192 GND.n7868 GND.n537 240.244
R13193 GND.n546 GND.n537 240.244
R13194 GND.n546 GND.n527 240.244
R13195 GND.n7883 GND.n527 240.244
R13196 GND.n7883 GND.n506 240.244
R13197 GND.n550 GND.n506 240.244
R13198 GND.n550 GND.n496 240.244
R13199 GND.n496 GND.n489 240.244
R13200 GND.n7965 GND.n489 240.244
R13201 GND.n7965 GND.n479 240.244
R13202 GND.n7969 GND.n479 240.244
R13203 GND.n7969 GND.n469 240.244
R13204 GND.n469 GND.n461 240.244
R13205 GND.n8007 GND.n461 240.244
R13206 GND.n8007 GND.n448 240.244
R13207 GND.n8021 GND.n448 240.244
R13208 GND.n8022 GND.n8021 240.244
R13209 GND.n8022 GND.n442 240.244
R13210 GND.n442 GND.n159 240.244
R13211 GND.n8025 GND.n159 240.244
R13212 GND.n8025 GND.n430 240.244
R13213 GND.n8131 GND.n430 240.244
R13214 GND.n8131 GND.n178 240.244
R13215 GND.n8141 GND.n178 240.244
R13216 GND.n8141 GND.n190 240.244
R13217 GND.n8146 GND.n190 240.244
R13218 GND.n8146 GND.n200 240.244
R13219 GND.n8156 GND.n200 240.244
R13220 GND.n8156 GND.n210 240.244
R13221 GND.n8161 GND.n210 240.244
R13222 GND.n8161 GND.n221 240.244
R13223 GND.n8171 GND.n221 240.244
R13224 GND.n8171 GND.n231 240.244
R13225 GND.n8176 GND.n231 240.244
R13226 GND.n8176 GND.n242 240.244
R13227 GND.n8186 GND.n242 240.244
R13228 GND.n8186 GND.n252 240.244
R13229 GND.n8191 GND.n252 240.244
R13230 GND.n8191 GND.n262 240.244
R13231 GND.n8201 GND.n262 240.244
R13232 GND.n8201 GND.n272 240.244
R13233 GND.n8206 GND.n272 240.244
R13234 GND.n8206 GND.n283 240.244
R13235 GND.n8216 GND.n283 240.244
R13236 GND.n8216 GND.n293 240.244
R13237 GND.n8221 GND.n293 240.244
R13238 GND.n8221 GND.n304 240.244
R13239 GND.n8232 GND.n304 240.244
R13240 GND.n8232 GND.n314 240.244
R13241 GND.n393 GND.n314 240.244
R13242 GND.n393 GND.n324 240.244
R13243 GND.n8239 GND.n324 240.244
R13244 GND.n8239 GND.n334 240.244
R13245 GND.n8457 GND.n334 240.244
R13246 GND.n8457 GND.n344 240.244
R13247 GND.n708 GND.n707 240.244
R13248 GND.n7718 GND.n707 240.244
R13249 GND.n7716 GND.n7715 240.244
R13250 GND.n7712 GND.n7711 240.244
R13251 GND.n7707 GND.n717 240.244
R13252 GND.n7705 GND.n7704 240.244
R13253 GND.n7701 GND.n7700 240.244
R13254 GND.n7697 GND.n7696 240.244
R13255 GND.n7693 GND.n7692 240.244
R13256 GND.n7688 GND.n7687 240.244
R13257 GND.n7684 GND.n7683 240.244
R13258 GND.n7680 GND.n7597 240.244
R13259 GND.n7678 GND.n7677 240.244
R13260 GND.n7674 GND.n7673 240.244
R13261 GND.n7670 GND.n7669 240.244
R13262 GND.n7666 GND.n7665 240.244
R13263 GND.n7662 GND.n7661 240.244
R13264 GND.n7658 GND.n7657 240.244
R13265 GND.n7654 GND.n7653 240.244
R13266 GND.n7650 GND.n7649 240.244
R13267 GND.n7646 GND.n7645 240.244
R13268 GND.n7642 GND.n7641 240.244
R13269 GND.n7638 GND.n7637 240.244
R13270 GND.n7634 GND.n7633 240.244
R13271 GND.n7755 GND.n646 240.244
R13272 GND.n7755 GND.n641 240.244
R13273 GND.n7763 GND.n641 240.244
R13274 GND.n7763 GND.n642 240.244
R13275 GND.n642 GND.n618 240.244
R13276 GND.n7792 GND.n618 240.244
R13277 GND.n7792 GND.n613 240.244
R13278 GND.n7800 GND.n613 240.244
R13279 GND.n7800 GND.n614 240.244
R13280 GND.n614 GND.n591 240.244
R13281 GND.n7827 GND.n591 240.244
R13282 GND.n7827 GND.n587 240.244
R13283 GND.n7833 GND.n587 240.244
R13284 GND.n7833 GND.n569 240.244
R13285 GND.n7854 GND.n569 240.244
R13286 GND.n7854 GND.n565 240.244
R13287 GND.n7860 GND.n565 240.244
R13288 GND.n7860 GND.n535 240.244
R13289 GND.n7892 GND.n535 240.244
R13290 GND.n7892 GND.n531 240.244
R13291 GND.n7898 GND.n531 240.244
R13292 GND.n7898 GND.n504 240.244
R13293 GND.n7945 GND.n504 240.244
R13294 GND.n7945 GND.n499 240.244
R13295 GND.n7953 GND.n499 240.244
R13296 GND.n7953 GND.n500 240.244
R13297 GND.n500 GND.n477 240.244
R13298 GND.n7982 GND.n477 240.244
R13299 GND.n7982 GND.n472 240.244
R13300 GND.n7990 GND.n472 240.244
R13301 GND.n7990 GND.n473 240.244
R13302 GND.n473 GND.n453 240.244
R13303 GND.n8016 GND.n453 240.244
R13304 GND.n8019 GND.n8016 240.244
R13305 GND.n8019 GND.n8018 240.244
R13306 GND.n8018 GND.n162 240.244
R13307 GND.n8565 GND.n162 240.244
R13308 GND.n8565 GND.n163 240.244
R13309 GND.n8124 GND.n163 240.244
R13310 GND.n8124 GND.n175 240.244
R13311 GND.n8560 GND.n175 240.244
R13312 GND.n8560 GND.n176 240.244
R13313 GND.n8552 GND.n176 240.244
R13314 GND.n8552 GND.n193 240.244
R13315 GND.n8548 GND.n193 240.244
R13316 GND.n8548 GND.n198 240.244
R13317 GND.n8540 GND.n198 240.244
R13318 GND.n8540 GND.n213 240.244
R13319 GND.n8536 GND.n213 240.244
R13320 GND.n8536 GND.n219 240.244
R13321 GND.n8528 GND.n219 240.244
R13322 GND.n8528 GND.n234 240.244
R13323 GND.n8524 GND.n234 240.244
R13324 GND.n8524 GND.n240 240.244
R13325 GND.n8516 GND.n240 240.244
R13326 GND.n8516 GND.n254 240.244
R13327 GND.n8512 GND.n254 240.244
R13328 GND.n8512 GND.n260 240.244
R13329 GND.n8504 GND.n260 240.244
R13330 GND.n8504 GND.n275 240.244
R13331 GND.n8500 GND.n275 240.244
R13332 GND.n8500 GND.n281 240.244
R13333 GND.n8492 GND.n281 240.244
R13334 GND.n8492 GND.n296 240.244
R13335 GND.n8488 GND.n296 240.244
R13336 GND.n8488 GND.n302 240.244
R13337 GND.n8480 GND.n302 240.244
R13338 GND.n8480 GND.n316 240.244
R13339 GND.n8476 GND.n316 240.244
R13340 GND.n8476 GND.n322 240.244
R13341 GND.n8468 GND.n322 240.244
R13342 GND.n8468 GND.n337 240.244
R13343 GND.n8464 GND.n337 240.244
R13344 GND.n5908 GND.n5907 240.244
R13345 GND.n5915 GND.n5914 240.244
R13346 GND.n5918 GND.n5917 240.244
R13347 GND.n5927 GND.n5926 240.244
R13348 GND.n5930 GND.n5929 240.244
R13349 GND.n5937 GND.n5936 240.244
R13350 GND.n5940 GND.n5939 240.244
R13351 GND.n5947 GND.n5946 240.244
R13352 GND.n5949 GND.n1664 240.244
R13353 GND.n5956 GND.n5955 240.244
R13354 GND.n6041 GND.n6040 240.244
R13355 GND.n5962 GND.n5961 240.244
R13356 GND.n5967 GND.n5963 240.244
R13357 GND.n5969 GND.n5968 240.244
R13358 GND.n5973 GND.n5972 240.244
R13359 GND.n5975 GND.n5974 240.244
R13360 GND.n5979 GND.n5978 240.244
R13361 GND.n5983 GND.n5980 240.244
R13362 GND.n5987 GND.n5986 240.244
R13363 GND.n5989 GND.n5988 240.244
R13364 GND.n5993 GND.n5992 240.244
R13365 GND.n5995 GND.n5994 240.244
R13366 GND.n6001 GND.n5998 240.244
R13367 GND.n4332 GND.n2131 240.244
R13368 GND.n4332 GND.n2122 240.244
R13369 GND.n2122 GND.n2113 240.244
R13370 GND.n4365 GND.n2113 240.244
R13371 GND.n4365 GND.n2103 240.244
R13372 GND.n4368 GND.n2103 240.244
R13373 GND.n4368 GND.n2093 240.244
R13374 GND.n2093 GND.n2084 240.244
R13375 GND.n4413 GND.n2084 240.244
R13376 GND.n4413 GND.n2074 240.244
R13377 GND.n4415 GND.n2074 240.244
R13378 GND.n4415 GND.n2064 240.244
R13379 GND.n4398 GND.n2064 240.244
R13380 GND.n4398 GND.n2040 240.244
R13381 GND.n2051 GND.n2040 240.244
R13382 GND.n2051 GND.n2030 240.244
R13383 GND.n2030 GND.n2022 240.244
R13384 GND.n4495 GND.n2022 240.244
R13385 GND.n4495 GND.n2012 240.244
R13386 GND.n4497 GND.n2012 240.244
R13387 GND.n4497 GND.n2002 240.244
R13388 GND.n4480 GND.n2002 240.244
R13389 GND.n4480 GND.n1978 240.244
R13390 GND.n1989 GND.n1978 240.244
R13391 GND.n1989 GND.n1968 240.244
R13392 GND.n1968 GND.n1960 240.244
R13393 GND.n4606 GND.n1960 240.244
R13394 GND.n4606 GND.n1948 240.244
R13395 GND.n1948 GND.n1938 240.244
R13396 GND.n4622 GND.n1938 240.244
R13397 GND.n4623 GND.n4622 240.244
R13398 GND.n4623 GND.n1883 240.244
R13399 GND.n1893 GND.n1883 240.244
R13400 GND.n1894 GND.n1893 240.244
R13401 GND.n1929 GND.n1894 240.244
R13402 GND.n1929 GND.n1900 240.244
R13403 GND.n1901 GND.n1900 240.244
R13404 GND.n1902 GND.n1901 240.244
R13405 GND.n1908 GND.n1902 240.244
R13406 GND.n4661 GND.n1908 240.244
R13407 GND.n4661 GND.n1865 240.244
R13408 GND.n4662 GND.n1865 240.244
R13409 GND.n4662 GND.n1858 240.244
R13410 GND.n1858 GND.n1837 240.244
R13411 GND.n1848 GND.n1837 240.244
R13412 GND.n1848 GND.n1828 240.244
R13413 GND.n1828 GND.n1820 240.244
R13414 GND.n4761 GND.n1820 240.244
R13415 GND.n4761 GND.n1810 240.244
R13416 GND.n4764 GND.n1810 240.244
R13417 GND.n4764 GND.n1800 240.244
R13418 GND.n4765 GND.n1800 240.244
R13419 GND.n4765 GND.n1793 240.244
R13420 GND.n1793 GND.n1776 240.244
R13421 GND.n4833 GND.n1776 240.244
R13422 GND.n4833 GND.n1766 240.244
R13423 GND.n1766 GND.n1759 240.244
R13424 GND.n4867 GND.n1759 240.244
R13425 GND.n4867 GND.n1749 240.244
R13426 GND.n4870 GND.n1749 240.244
R13427 GND.n4870 GND.n1739 240.244
R13428 GND.n1739 GND.n1731 240.244
R13429 GND.n4913 GND.n1731 240.244
R13430 GND.n4913 GND.n1719 240.244
R13431 GND.n4915 GND.n1719 240.244
R13432 GND.n4915 GND.n1701 240.244
R13433 GND.n5862 GND.n1701 240.244
R13434 GND.n5862 GND.n1691 240.244
R13435 GND.n5865 GND.n1691 240.244
R13436 GND.n5865 GND.n1683 240.244
R13437 GND.n5868 GND.n1683 240.244
R13438 GND.n5868 GND.n1605 240.244
R13439 GND.n6047 GND.n1605 240.244
R13440 GND.n4311 GND.n4157 240.244
R13441 GND.n4307 GND.n4157 240.244
R13442 GND.n4305 GND.n4304 240.244
R13443 GND.n4301 GND.n4300 240.244
R13444 GND.n4296 GND.n4166 240.244
R13445 GND.n4294 GND.n4293 240.244
R13446 GND.n4290 GND.n4289 240.244
R13447 GND.n4286 GND.n4285 240.244
R13448 GND.n4282 GND.n4281 240.244
R13449 GND.n4277 GND.n4276 240.244
R13450 GND.n4273 GND.n4272 240.244
R13451 GND.n4269 GND.n4268 240.244
R13452 GND.n4265 GND.n4264 240.244
R13453 GND.n4261 GND.n4260 240.244
R13454 GND.n4257 GND.n4256 240.244
R13455 GND.n4253 GND.n4252 240.244
R13456 GND.n4249 GND.n4248 240.244
R13457 GND.n4245 GND.n4244 240.244
R13458 GND.n4241 GND.n4240 240.244
R13459 GND.n4237 GND.n4236 240.244
R13460 GND.n4233 GND.n4232 240.244
R13461 GND.n4229 GND.n4228 240.244
R13462 GND.n4225 GND.n4224 240.244
R13463 GND.n4221 GND.n4220 240.244
R13464 GND.n4346 GND.n2125 240.244
R13465 GND.n4354 GND.n2125 240.244
R13466 GND.n4354 GND.n2126 240.244
R13467 GND.n2126 GND.n2101 240.244
R13468 GND.n4382 GND.n2101 240.244
R13469 GND.n4382 GND.n2096 240.244
R13470 GND.n4390 GND.n2096 240.244
R13471 GND.n4390 GND.n2097 240.244
R13472 GND.n2097 GND.n2072 240.244
R13473 GND.n4425 GND.n2072 240.244
R13474 GND.n4425 GND.n2068 240.244
R13475 GND.n4431 GND.n2068 240.244
R13476 GND.n4431 GND.n2038 240.244
R13477 GND.n4464 GND.n2038 240.244
R13478 GND.n4464 GND.n2033 240.244
R13479 GND.n4472 GND.n2033 240.244
R13480 GND.n4472 GND.n2034 240.244
R13481 GND.n2034 GND.n2010 240.244
R13482 GND.n4507 GND.n2010 240.244
R13483 GND.n4507 GND.n2006 240.244
R13484 GND.n4513 GND.n2006 240.244
R13485 GND.n4513 GND.n1976 240.244
R13486 GND.n4582 GND.n1976 240.244
R13487 GND.n4582 GND.n1971 240.244
R13488 GND.n4590 GND.n1971 240.244
R13489 GND.n4590 GND.n1972 240.244
R13490 GND.n1972 GND.n1946 240.244
R13491 GND.n4614 GND.n1946 240.244
R13492 GND.n4614 GND.n1942 240.244
R13493 GND.n4620 GND.n1942 240.244
R13494 GND.n4620 GND.n1880 240.244
R13495 GND.n4686 GND.n1880 240.244
R13496 GND.n4686 GND.n1881 240.244
R13497 GND.n1926 GND.n1881 240.244
R13498 GND.n4637 GND.n1926 240.244
R13499 GND.n4640 GND.n4637 240.244
R13500 GND.n4640 GND.n1913 240.244
R13501 GND.n4653 GND.n1913 240.244
R13502 GND.n4656 GND.n4653 240.244
R13503 GND.n4656 GND.n1868 240.244
R13504 GND.n4693 GND.n1868 240.244
R13505 GND.n4693 GND.n1869 240.244
R13506 GND.n1869 GND.n1835 240.244
R13507 GND.n4741 GND.n1835 240.244
R13508 GND.n4741 GND.n1830 240.244
R13509 GND.n4749 GND.n1830 240.244
R13510 GND.n4749 GND.n1831 240.244
R13511 GND.n1831 GND.n1808 240.244
R13512 GND.n4779 GND.n1808 240.244
R13513 GND.n4779 GND.n1803 240.244
R13514 GND.n4787 GND.n1803 240.244
R13515 GND.n4787 GND.n1804 240.244
R13516 GND.n1804 GND.n1774 240.244
R13517 GND.n4847 GND.n1774 240.244
R13518 GND.n4847 GND.n1769 240.244
R13519 GND.n4855 GND.n1769 240.244
R13520 GND.n4855 GND.n1770 240.244
R13521 GND.n1770 GND.n1747 240.244
R13522 GND.n4884 GND.n1747 240.244
R13523 GND.n4884 GND.n1742 240.244
R13524 GND.n4892 GND.n1742 240.244
R13525 GND.n4892 GND.n1743 240.244
R13526 GND.n1743 GND.n1717 240.244
R13527 GND.n4922 GND.n1717 240.244
R13528 GND.n4922 GND.n1713 240.244
R13529 GND.n4928 GND.n1713 240.244
R13530 GND.n4928 GND.n1690 240.244
R13531 GND.n5882 GND.n1690 240.244
R13532 GND.n5882 GND.n1686 240.244
R13533 GND.n5889 GND.n1686 240.244
R13534 GND.n5889 GND.n1675 240.244
R13535 GND.n5900 GND.n1675 240.244
R13536 GND.n5900 GND.n1608 240.244
R13537 GND.n6923 GND.n6921 240.244
R13538 GND.n6930 GND.n1075 240.244
R13539 GND.n6934 GND.n6932 240.244
R13540 GND.n6940 GND.n1073 240.244
R13541 GND.n6944 GND.n6942 240.244
R13542 GND.n6950 GND.n1071 240.244
R13543 GND.n6953 GND.n6952 240.244
R13544 GND.n6961 GND.n6960 240.244
R13545 GND.n6964 GND.n6963 240.244
R13546 GND.n6110 GND.n1563 240.244
R13547 GND.n6116 GND.n1563 240.244
R13548 GND.n6116 GND.n1552 240.244
R13549 GND.n6126 GND.n1552 240.244
R13550 GND.n6126 GND.n1547 240.244
R13551 GND.n6141 GND.n1547 240.244
R13552 GND.n6141 GND.n1548 240.244
R13553 GND.n1548 GND.n1538 240.244
R13554 GND.n6136 GND.n1538 240.244
R13555 GND.n6136 GND.n1503 240.244
R13556 GND.n1503 GND.n1492 240.244
R13557 GND.n6330 GND.n1492 240.244
R13558 GND.n6330 GND.n1488 240.244
R13559 GND.n6336 GND.n1488 240.244
R13560 GND.n6336 GND.n1476 240.244
R13561 GND.n6346 GND.n1476 240.244
R13562 GND.n6346 GND.n1472 240.244
R13563 GND.n6352 GND.n1472 240.244
R13564 GND.n6352 GND.n1460 240.244
R13565 GND.n6362 GND.n1460 240.244
R13566 GND.n6362 GND.n1456 240.244
R13567 GND.n6368 GND.n1456 240.244
R13568 GND.n6368 GND.n1444 240.244
R13569 GND.n6377 GND.n1444 240.244
R13570 GND.n6377 GND.n1440 240.244
R13571 GND.n6383 GND.n1440 240.244
R13572 GND.n6383 GND.n1427 240.244
R13573 GND.n6395 GND.n1427 240.244
R13574 GND.n6395 GND.n1423 240.244
R13575 GND.n6403 GND.n1423 240.244
R13576 GND.n6403 GND.n1321 240.244
R13577 GND.n1321 GND.n1311 240.244
R13578 GND.n6569 GND.n1311 240.244
R13579 GND.n6569 GND.n1307 240.244
R13580 GND.n6575 GND.n1307 240.244
R13581 GND.n6575 GND.n1295 240.244
R13582 GND.n6585 GND.n1295 240.244
R13583 GND.n6585 GND.n1291 240.244
R13584 GND.n6591 GND.n1291 240.244
R13585 GND.n6591 GND.n1279 240.244
R13586 GND.n6601 GND.n1279 240.244
R13587 GND.n6601 GND.n1275 240.244
R13588 GND.n6607 GND.n1275 240.244
R13589 GND.n6607 GND.n1263 240.244
R13590 GND.n6616 GND.n1263 240.244
R13591 GND.n6616 GND.n1259 240.244
R13592 GND.n6622 GND.n1259 240.244
R13593 GND.n6622 GND.n1247 240.244
R13594 GND.n6632 GND.n1247 240.244
R13595 GND.n6632 GND.n1243 240.244
R13596 GND.n6638 GND.n1243 240.244
R13597 GND.n6638 GND.n1231 240.244
R13598 GND.n6648 GND.n1231 240.244
R13599 GND.n6648 GND.n1226 240.244
R13600 GND.n6663 GND.n1226 240.244
R13601 GND.n6663 GND.n1227 240.244
R13602 GND.n1227 GND.n1217 240.244
R13603 GND.n6658 GND.n1217 240.244
R13604 GND.n6658 GND.n1168 240.244
R13605 GND.n1168 GND.n1157 240.244
R13606 GND.n6827 GND.n1157 240.244
R13607 GND.n6827 GND.n1153 240.244
R13608 GND.n6833 GND.n1153 240.244
R13609 GND.n6833 GND.n1141 240.244
R13610 GND.n6843 GND.n1141 240.244
R13611 GND.n6843 GND.n1137 240.244
R13612 GND.n6849 GND.n1137 240.244
R13613 GND.n6849 GND.n1125 240.244
R13614 GND.n6859 GND.n1125 240.244
R13615 GND.n6859 GND.n1121 240.244
R13616 GND.n6865 GND.n1121 240.244
R13617 GND.n6865 GND.n1109 240.244
R13618 GND.n6874 GND.n1109 240.244
R13619 GND.n6874 GND.n1104 240.244
R13620 GND.n6885 GND.n1104 240.244
R13621 GND.n6885 GND.n1105 240.244
R13622 GND.n1105 GND.n1095 240.244
R13623 GND.n1095 GND.n1058 240.244
R13624 GND.n6978 GND.n1058 240.244
R13625 GND.n6978 GND.n1059 240.244
R13626 GND.n1059 GND.n1048 240.244
R13627 GND.n6973 GND.n1048 240.244
R13628 GND.n6973 GND.n6972 240.244
R13629 GND.n1587 GND.n1586 240.244
R13630 GND.n6093 GND.n1586 240.244
R13631 GND.n6091 GND.n6090 240.244
R13632 GND.n6053 GND.n1594 240.244
R13633 GND.n6055 GND.n6054 240.244
R13634 GND.n6057 GND.n6056 240.244
R13635 GND.n6059 GND.n6058 240.244
R13636 GND.n6061 GND.n6060 240.244
R13637 GND.n6070 GND.n6064 240.244
R13638 GND.n6066 GND.n1566 240.244
R13639 GND.n5593 GND.n1568 240.244
R13640 GND.n5593 GND.n1561 240.244
R13641 GND.n5599 GND.n1561 240.244
R13642 GND.n5599 GND.n1554 240.244
R13643 GND.n5622 GND.n1554 240.244
R13644 GND.n5622 GND.n1545 240.244
R13645 GND.n5618 GND.n1545 240.244
R13646 GND.n5618 GND.n1537 240.244
R13647 GND.n5615 GND.n1537 240.244
R13648 GND.n5615 GND.n1502 240.244
R13649 GND.n5612 GND.n1502 240.244
R13650 GND.n5612 GND.n1494 240.244
R13651 GND.n6311 GND.n1494 240.244
R13652 GND.n6311 GND.n1486 240.244
R13653 GND.n6307 GND.n1486 240.244
R13654 GND.n6307 GND.n1478 240.244
R13655 GND.n6212 GND.n1478 240.244
R13656 GND.n6212 GND.n1470 240.244
R13657 GND.n6217 GND.n1470 240.244
R13658 GND.n6217 GND.n1462 240.244
R13659 GND.n6220 GND.n1462 240.244
R13660 GND.n6220 GND.n1454 240.244
R13661 GND.n6225 GND.n1454 240.244
R13662 GND.n6225 GND.n1446 240.244
R13663 GND.n6228 GND.n1446 240.244
R13664 GND.n6228 GND.n1438 240.244
R13665 GND.n6236 GND.n1438 240.244
R13666 GND.n6236 GND.n1429 240.244
R13667 GND.n1429 GND.n1421 240.244
R13668 GND.n6405 GND.n1421 240.244
R13669 GND.n6405 GND.n1320 240.244
R13670 GND.n6410 GND.n1320 240.244
R13671 GND.n6410 GND.n1312 240.244
R13672 GND.n6413 GND.n1312 240.244
R13673 GND.n6413 GND.n1305 240.244
R13674 GND.n6418 GND.n1305 240.244
R13675 GND.n6418 GND.n1297 240.244
R13676 GND.n6421 GND.n1297 240.244
R13677 GND.n6421 GND.n1289 240.244
R13678 GND.n6426 GND.n1289 240.244
R13679 GND.n6426 GND.n1281 240.244
R13680 GND.n6429 GND.n1281 240.244
R13681 GND.n6429 GND.n1273 240.244
R13682 GND.n6434 GND.n1273 240.244
R13683 GND.n6434 GND.n1265 240.244
R13684 GND.n6437 GND.n1265 240.244
R13685 GND.n6437 GND.n1257 240.244
R13686 GND.n6442 GND.n1257 240.244
R13687 GND.n6442 GND.n1249 240.244
R13688 GND.n6446 GND.n1249 240.244
R13689 GND.n6446 GND.n1241 240.244
R13690 GND.n6474 GND.n1241 240.244
R13691 GND.n6474 GND.n1233 240.244
R13692 GND.n6470 GND.n1233 240.244
R13693 GND.n6470 GND.n1224 240.244
R13694 GND.n6467 GND.n1224 240.244
R13695 GND.n6467 GND.n1216 240.244
R13696 GND.n6464 GND.n1216 240.244
R13697 GND.n6464 GND.n1167 240.244
R13698 GND.n6461 GND.n1167 240.244
R13699 GND.n6461 GND.n1159 240.244
R13700 GND.n6808 GND.n1159 240.244
R13701 GND.n6808 GND.n1151 240.244
R13702 GND.n6804 GND.n1151 240.244
R13703 GND.n6804 GND.n1143 240.244
R13704 GND.n6794 GND.n1143 240.244
R13705 GND.n6794 GND.n1135 240.244
R13706 GND.n6790 GND.n1135 240.244
R13707 GND.n6790 GND.n1127 240.244
R13708 GND.n6724 GND.n1127 240.244
R13709 GND.n6724 GND.n1119 240.244
R13710 GND.n6727 GND.n1119 240.244
R13711 GND.n6727 GND.n1111 240.244
R13712 GND.n6740 GND.n1111 240.244
R13713 GND.n6740 GND.n1102 240.244
R13714 GND.n6736 GND.n1102 240.244
R13715 GND.n6736 GND.n1086 240.244
R13716 GND.n6906 GND.n1086 240.244
R13717 GND.n6906 GND.n1056 240.244
R13718 GND.n1082 GND.n1056 240.244
R13719 GND.n1082 GND.n1047 240.244
R13720 GND.n6913 GND.n1047 240.244
R13721 GND.n6913 GND.n1079 240.244
R13722 GND.n363 GND.n347 240.244
R13723 GND.n371 GND.n370 240.244
R13724 GND.n373 GND.n360 240.244
R13725 GND.n379 GND.n357 240.244
R13726 GND.n7736 GND.n649 240.244
R13727 GND.n649 GND.n636 240.244
R13728 GND.n7765 GND.n636 240.244
R13729 GND.n7765 GND.n632 240.244
R13730 GND.n7773 GND.n632 240.244
R13731 GND.n7773 GND.n621 240.244
R13732 GND.n621 GND.n608 240.244
R13733 GND.n7802 GND.n608 240.244
R13734 GND.n7802 GND.n604 240.244
R13735 GND.n7814 GND.n604 240.244
R13736 GND.n7814 GND.n594 240.244
R13737 GND.n7810 GND.n594 240.244
R13738 GND.n7810 GND.n581 240.244
R13739 GND.n7838 GND.n581 240.244
R13740 GND.n7838 GND.n572 240.244
R13741 GND.n7845 GND.n572 240.244
R13742 GND.n7845 GND.n557 240.244
R13743 GND.n7870 GND.n557 240.244
R13744 GND.n7870 GND.n538 240.244
R13745 GND.n7873 GND.n538 240.244
R13746 GND.n7873 GND.n528 240.244
R13747 GND.n7881 GND.n528 240.244
R13748 GND.n7881 GND.n507 240.244
R13749 GND.n507 GND.n494 240.244
R13750 GND.n7955 GND.n494 240.244
R13751 GND.n7955 GND.n490 240.244
R13752 GND.n7963 GND.n490 240.244
R13753 GND.n7963 GND.n480 240.244
R13754 GND.n480 GND.n467 240.244
R13755 GND.n7992 GND.n467 240.244
R13756 GND.n7992 GND.n463 240.244
R13757 GND.n8005 GND.n463 240.244
R13758 GND.n8005 GND.n456 240.244
R13759 GND.n456 GND.n450 240.244
R13760 GND.n8000 GND.n450 240.244
R13761 GND.n8000 GND.n156 240.244
R13762 GND.n8567 GND.n156 240.244
R13763 GND.n8567 GND.n157 240.244
R13764 GND.n428 GND.n157 240.244
R13765 GND.n8133 GND.n428 240.244
R13766 GND.n8133 GND.n179 240.244
R13767 GND.n8139 GND.n179 240.244
R13768 GND.n8139 GND.n191 240.244
R13769 GND.n8148 GND.n191 240.244
R13770 GND.n8148 GND.n201 240.244
R13771 GND.n8154 GND.n201 240.244
R13772 GND.n8154 GND.n211 240.244
R13773 GND.n8163 GND.n211 240.244
R13774 GND.n8163 GND.n222 240.244
R13775 GND.n8169 GND.n222 240.244
R13776 GND.n8169 GND.n232 240.244
R13777 GND.n8178 GND.n232 240.244
R13778 GND.n8178 GND.n243 240.244
R13779 GND.n8184 GND.n243 240.244
R13780 GND.n8184 GND.n253 240.244
R13781 GND.n8193 GND.n253 240.244
R13782 GND.n8193 GND.n263 240.244
R13783 GND.n8199 GND.n263 240.244
R13784 GND.n8199 GND.n273 240.244
R13785 GND.n8208 GND.n273 240.244
R13786 GND.n8208 GND.n284 240.244
R13787 GND.n8214 GND.n284 240.244
R13788 GND.n8214 GND.n294 240.244
R13789 GND.n8223 GND.n294 240.244
R13790 GND.n8223 GND.n305 240.244
R13791 GND.n8230 GND.n305 240.244
R13792 GND.n8230 GND.n315 240.244
R13793 GND.n8245 GND.n315 240.244
R13794 GND.n8245 GND.n325 240.244
R13795 GND.n8241 GND.n325 240.244
R13796 GND.n8241 GND.n335 240.244
R13797 GND.n8455 GND.n335 240.244
R13798 GND.n8455 GND.n345 240.244
R13799 GND.n700 GND.n697 240.244
R13800 GND.n704 GND.n703 240.244
R13801 GND.n7727 GND.n670 240.244
R13802 GND.n666 GND.n659 240.244
R13803 GND.n7753 GND.n651 240.244
R13804 GND.n7753 GND.n652 240.244
R13805 GND.n652 GND.n640 240.244
R13806 GND.n7742 GND.n640 240.244
R13807 GND.n7742 GND.n623 240.244
R13808 GND.n7790 GND.n623 240.244
R13809 GND.n7790 GND.n624 240.244
R13810 GND.n624 GND.n612 240.244
R13811 GND.n7785 GND.n612 240.244
R13812 GND.n7785 GND.n596 240.244
R13813 GND.n7825 GND.n596 240.244
R13814 GND.n7825 GND.n597 240.244
R13815 GND.n597 GND.n586 240.244
R13816 GND.n586 GND.n574 240.244
R13817 GND.n7852 GND.n574 240.244
R13818 GND.n7852 GND.n563 240.244
R13819 GND.n7862 GND.n563 240.244
R13820 GND.n7862 GND.n540 240.244
R13821 GND.n7890 GND.n540 240.244
R13822 GND.n7890 GND.n541 240.244
R13823 GND.n541 GND.n530 240.244
R13824 GND.n530 GND.n509 240.244
R13825 GND.n7943 GND.n509 240.244
R13826 GND.n7943 GND.n510 240.244
R13827 GND.n510 GND.n498 240.244
R13828 GND.n7938 GND.n498 240.244
R13829 GND.n7938 GND.n482 240.244
R13830 GND.n7980 GND.n482 240.244
R13831 GND.n7980 GND.n483 240.244
R13832 GND.n483 GND.n471 240.244
R13833 GND.n7975 GND.n471 240.244
R13834 GND.n7975 GND.n457 240.244
R13835 GND.n8014 GND.n457 240.244
R13836 GND.n8014 GND.n452 240.244
R13837 GND.n452 GND.n443 240.244
R13838 GND.n8031 GND.n443 240.244
R13839 GND.n8031 GND.n161 240.244
R13840 GND.n434 GND.n161 240.244
R13841 GND.n8126 GND.n434 240.244
R13842 GND.n8126 GND.n181 240.244
R13843 GND.n8558 GND.n181 240.244
R13844 GND.n8558 GND.n182 240.244
R13845 GND.n8554 GND.n182 240.244
R13846 GND.n8554 GND.n188 240.244
R13847 GND.n8546 GND.n188 240.244
R13848 GND.n8546 GND.n203 240.244
R13849 GND.n8542 GND.n203 240.244
R13850 GND.n8542 GND.n208 240.244
R13851 GND.n8534 GND.n208 240.244
R13852 GND.n8534 GND.n224 240.244
R13853 GND.n8530 GND.n224 240.244
R13854 GND.n8530 GND.n229 240.244
R13855 GND.n8522 GND.n229 240.244
R13856 GND.n8522 GND.n245 240.244
R13857 GND.n8518 GND.n245 240.244
R13858 GND.n8518 GND.n250 240.244
R13859 GND.n8510 GND.n250 240.244
R13860 GND.n8510 GND.n265 240.244
R13861 GND.n8506 GND.n265 240.244
R13862 GND.n8506 GND.n270 240.244
R13863 GND.n8498 GND.n270 240.244
R13864 GND.n8498 GND.n286 240.244
R13865 GND.n8494 GND.n286 240.244
R13866 GND.n8494 GND.n291 240.244
R13867 GND.n8486 GND.n291 240.244
R13868 GND.n8486 GND.n307 240.244
R13869 GND.n8482 GND.n307 240.244
R13870 GND.n8482 GND.n312 240.244
R13871 GND.n8474 GND.n312 240.244
R13872 GND.n8474 GND.n327 240.244
R13873 GND.n8470 GND.n327 240.244
R13874 GND.n8470 GND.n332 240.244
R13875 GND.n8462 GND.n332 240.244
R13876 GND.n3935 GND.n2250 240.244
R13877 GND.n3929 GND.n2250 240.244
R13878 GND.n3929 GND.n2254 240.244
R13879 GND.n3925 GND.n2254 240.244
R13880 GND.n3925 GND.n2256 240.244
R13881 GND.n3921 GND.n2256 240.244
R13882 GND.n3921 GND.n2261 240.244
R13883 GND.n3917 GND.n2261 240.244
R13884 GND.n3917 GND.n2263 240.244
R13885 GND.n3913 GND.n2263 240.244
R13886 GND.n3913 GND.n2269 240.244
R13887 GND.n3909 GND.n2269 240.244
R13888 GND.n3909 GND.n2271 240.244
R13889 GND.n3905 GND.n2271 240.244
R13890 GND.n3905 GND.n2277 240.244
R13891 GND.n3901 GND.n2277 240.244
R13892 GND.n3901 GND.n2279 240.244
R13893 GND.n3897 GND.n2279 240.244
R13894 GND.n3897 GND.n2285 240.244
R13895 GND.n3893 GND.n2285 240.244
R13896 GND.n3893 GND.n2287 240.244
R13897 GND.n3889 GND.n2287 240.244
R13898 GND.n3889 GND.n2293 240.244
R13899 GND.n3885 GND.n2293 240.244
R13900 GND.n3885 GND.n2295 240.244
R13901 GND.n3881 GND.n2295 240.244
R13902 GND.n3881 GND.n2301 240.244
R13903 GND.n3877 GND.n2301 240.244
R13904 GND.n3877 GND.n2303 240.244
R13905 GND.n3873 GND.n2303 240.244
R13906 GND.n3873 GND.n2309 240.244
R13907 GND.n3869 GND.n2309 240.244
R13908 GND.n3869 GND.n2311 240.244
R13909 GND.n3865 GND.n2311 240.244
R13910 GND.n3865 GND.n2317 240.244
R13911 GND.n3861 GND.n2317 240.244
R13912 GND.n3861 GND.n2319 240.244
R13913 GND.n3857 GND.n2319 240.244
R13914 GND.n3857 GND.n2325 240.244
R13915 GND.n3853 GND.n2325 240.244
R13916 GND.n3853 GND.n2327 240.244
R13917 GND.n3849 GND.n2327 240.244
R13918 GND.n3849 GND.n2333 240.244
R13919 GND.n3845 GND.n2333 240.244
R13920 GND.n3845 GND.n2335 240.244
R13921 GND.n3841 GND.n2335 240.244
R13922 GND.n3841 GND.n2341 240.244
R13923 GND.n3837 GND.n2341 240.244
R13924 GND.n3837 GND.n2343 240.244
R13925 GND.n3833 GND.n2343 240.244
R13926 GND.n3833 GND.n2349 240.244
R13927 GND.n3829 GND.n2349 240.244
R13928 GND.n3829 GND.n2351 240.244
R13929 GND.n3825 GND.n2351 240.244
R13930 GND.n3825 GND.n2357 240.244
R13931 GND.n3821 GND.n2357 240.244
R13932 GND.n3821 GND.n2359 240.244
R13933 GND.n3817 GND.n2359 240.244
R13934 GND.n3817 GND.n2365 240.244
R13935 GND.n3813 GND.n2365 240.244
R13936 GND.n3813 GND.n2367 240.244
R13937 GND.n3809 GND.n2367 240.244
R13938 GND.n3809 GND.n2373 240.244
R13939 GND.n3805 GND.n2373 240.244
R13940 GND.n3805 GND.n2375 240.244
R13941 GND.n3801 GND.n2375 240.244
R13942 GND.n3801 GND.n2381 240.244
R13943 GND.n3797 GND.n2381 240.244
R13944 GND.n3797 GND.n2383 240.244
R13945 GND.n3793 GND.n2383 240.244
R13946 GND.n3793 GND.n2389 240.244
R13947 GND.n3789 GND.n2389 240.244
R13948 GND.n3789 GND.n2391 240.244
R13949 GND.n3785 GND.n2391 240.244
R13950 GND.n3785 GND.n2397 240.244
R13951 GND.n3781 GND.n2397 240.244
R13952 GND.n3781 GND.n2399 240.244
R13953 GND.n3777 GND.n2399 240.244
R13954 GND.n3777 GND.n2405 240.244
R13955 GND.n3773 GND.n2405 240.244
R13956 GND.n3773 GND.n2407 240.244
R13957 GND.n3769 GND.n2407 240.244
R13958 GND.n3769 GND.n2413 240.244
R13959 GND.n3765 GND.n2413 240.244
R13960 GND.n3765 GND.n2415 240.244
R13961 GND.n3761 GND.n2415 240.244
R13962 GND.n3761 GND.n2421 240.244
R13963 GND.n3757 GND.n2421 240.244
R13964 GND.n3757 GND.n2423 240.244
R13965 GND.n3753 GND.n2423 240.244
R13966 GND.n3753 GND.n2429 240.244
R13967 GND.n3749 GND.n2429 240.244
R13968 GND.n3749 GND.n2431 240.244
R13969 GND.n3745 GND.n2431 240.244
R13970 GND.n3745 GND.n2437 240.244
R13971 GND.n3741 GND.n2437 240.244
R13972 GND.n3741 GND.n2439 240.244
R13973 GND.n3737 GND.n2439 240.244
R13974 GND.n3737 GND.n2445 240.244
R13975 GND.n3733 GND.n2445 240.244
R13976 GND.n3733 GND.n2447 240.244
R13977 GND.n3729 GND.n2447 240.244
R13978 GND.n3729 GND.n2453 240.244
R13979 GND.n3725 GND.n2453 240.244
R13980 GND.n3725 GND.n2455 240.244
R13981 GND.n3721 GND.n2455 240.244
R13982 GND.n3721 GND.n2461 240.244
R13983 GND.n3717 GND.n2461 240.244
R13984 GND.n3717 GND.n2463 240.244
R13985 GND.n3713 GND.n2463 240.244
R13986 GND.n3713 GND.n2469 240.244
R13987 GND.n3709 GND.n2469 240.244
R13988 GND.n3709 GND.n2471 240.244
R13989 GND.n3705 GND.n2471 240.244
R13990 GND.n3705 GND.n2477 240.244
R13991 GND.n3701 GND.n2477 240.244
R13992 GND.n3701 GND.n2479 240.244
R13993 GND.n3697 GND.n2479 240.244
R13994 GND.n3697 GND.n2485 240.244
R13995 GND.n3693 GND.n2485 240.244
R13996 GND.n3693 GND.n2487 240.244
R13997 GND.n3689 GND.n2487 240.244
R13998 GND.n3689 GND.n2493 240.244
R13999 GND.n3685 GND.n2493 240.244
R14000 GND.n3685 GND.n2495 240.244
R14001 GND.n3681 GND.n2495 240.244
R14002 GND.n3681 GND.n2501 240.244
R14003 GND.n3677 GND.n2501 240.244
R14004 GND.n3677 GND.n2503 240.244
R14005 GND.n3673 GND.n2503 240.244
R14006 GND.n3673 GND.n2509 240.244
R14007 GND.n3669 GND.n2509 240.244
R14008 GND.n3669 GND.n2511 240.244
R14009 GND.n3665 GND.n2511 240.244
R14010 GND.n3665 GND.n2517 240.244
R14011 GND.n3661 GND.n2517 240.244
R14012 GND.n3661 GND.n2519 240.244
R14013 GND.n3657 GND.n2519 240.244
R14014 GND.n3657 GND.n2525 240.244
R14015 GND.n3653 GND.n2525 240.244
R14016 GND.n3653 GND.n2527 240.244
R14017 GND.n3649 GND.n2527 240.244
R14018 GND.n3649 GND.n2533 240.244
R14019 GND.n3645 GND.n2533 240.244
R14020 GND.n3645 GND.n2535 240.244
R14021 GND.n3641 GND.n2535 240.244
R14022 GND.n3641 GND.n2541 240.244
R14023 GND.n3637 GND.n2541 240.244
R14024 GND.n3637 GND.n2543 240.244
R14025 GND.n3633 GND.n2543 240.244
R14026 GND.n3633 GND.n2549 240.244
R14027 GND.n3629 GND.n2549 240.244
R14028 GND.n3629 GND.n2551 240.244
R14029 GND.n3625 GND.n2551 240.244
R14030 GND.n3625 GND.n2557 240.244
R14031 GND.n3621 GND.n2557 240.244
R14032 GND.n3621 GND.n2559 240.244
R14033 GND.n3617 GND.n2559 240.244
R14034 GND.n3617 GND.n2565 240.244
R14035 GND.n3613 GND.n2565 240.244
R14036 GND.n3613 GND.n2567 240.244
R14037 GND.n3609 GND.n2567 240.244
R14038 GND.n3609 GND.n2573 240.244
R14039 GND.n3605 GND.n2573 240.244
R14040 GND.n3605 GND.n2575 240.244
R14041 GND.n3601 GND.n2575 240.244
R14042 GND.n3601 GND.n2581 240.244
R14043 GND.n3597 GND.n2581 240.244
R14044 GND.n3597 GND.n2583 240.244
R14045 GND.n3593 GND.n2583 240.244
R14046 GND.n3593 GND.n2589 240.244
R14047 GND.n3589 GND.n2589 240.244
R14048 GND.n3589 GND.n2591 240.244
R14049 GND.n3585 GND.n2591 240.244
R14050 GND.n3585 GND.n2597 240.244
R14051 GND.n3581 GND.n2597 240.244
R14052 GND.n3581 GND.n2599 240.244
R14053 GND.n3577 GND.n2599 240.244
R14054 GND.n3577 GND.n2605 240.244
R14055 GND.n3573 GND.n2605 240.244
R14056 GND.n3573 GND.n2607 240.244
R14057 GND.n3569 GND.n2607 240.244
R14058 GND.n3569 GND.n2613 240.244
R14059 GND.n3565 GND.n2613 240.244
R14060 GND.n3565 GND.n2615 240.244
R14061 GND.n3561 GND.n2615 240.244
R14062 GND.n3561 GND.n2621 240.244
R14063 GND.n3557 GND.n2621 240.244
R14064 GND.n3557 GND.n2623 240.244
R14065 GND.n3553 GND.n2623 240.244
R14066 GND.n3553 GND.n2629 240.244
R14067 GND.n3549 GND.n2629 240.244
R14068 GND.n3549 GND.n2631 240.244
R14069 GND.n3545 GND.n2631 240.244
R14070 GND.n3545 GND.n2637 240.244
R14071 GND.n3541 GND.n2637 240.244
R14072 GND.n3541 GND.n2639 240.244
R14073 GND.n3537 GND.n2639 240.244
R14074 GND.n3537 GND.n2645 240.244
R14075 GND.n3533 GND.n2645 240.244
R14076 GND.n3533 GND.n2647 240.244
R14077 GND.n3529 GND.n2647 240.244
R14078 GND.n3529 GND.n2653 240.244
R14079 GND.n3525 GND.n2653 240.244
R14080 GND.n3525 GND.n2655 240.244
R14081 GND.n3521 GND.n2655 240.244
R14082 GND.n3521 GND.n2661 240.244
R14083 GND.n3517 GND.n2661 240.244
R14084 GND.n3517 GND.n2663 240.244
R14085 GND.n3513 GND.n2663 240.244
R14086 GND.n3513 GND.n2669 240.244
R14087 GND.n3509 GND.n2669 240.244
R14088 GND.n3509 GND.n2671 240.244
R14089 GND.n3505 GND.n2671 240.244
R14090 GND.n3505 GND.n2677 240.244
R14091 GND.n3501 GND.n2677 240.244
R14092 GND.n3501 GND.n2679 240.244
R14093 GND.n3497 GND.n2679 240.244
R14094 GND.n3497 GND.n2685 240.244
R14095 GND.n3493 GND.n2685 240.244
R14096 GND.n3493 GND.n2687 240.244
R14097 GND.n3489 GND.n2687 240.244
R14098 GND.n3489 GND.n2693 240.244
R14099 GND.n3485 GND.n2693 240.244
R14100 GND.n3485 GND.n2695 240.244
R14101 GND.n3481 GND.n2695 240.244
R14102 GND.n3481 GND.n2701 240.244
R14103 GND.n3477 GND.n2701 240.244
R14104 GND.n3477 GND.n2703 240.244
R14105 GND.n3473 GND.n2703 240.244
R14106 GND.n3473 GND.n2709 240.244
R14107 GND.n3469 GND.n2709 240.244
R14108 GND.n3469 GND.n2711 240.244
R14109 GND.n3465 GND.n2711 240.244
R14110 GND.n3465 GND.n2717 240.244
R14111 GND.n3461 GND.n2717 240.244
R14112 GND.n3461 GND.n2719 240.244
R14113 GND.n3457 GND.n2719 240.244
R14114 GND.n3457 GND.n2725 240.244
R14115 GND.n3453 GND.n2725 240.244
R14116 GND.n3453 GND.n2727 240.244
R14117 GND.n3449 GND.n2727 240.244
R14118 GND.n3449 GND.n2733 240.244
R14119 GND.n3445 GND.n2733 240.244
R14120 GND.n3445 GND.n2735 240.244
R14121 GND.n3441 GND.n2735 240.244
R14122 GND.n3441 GND.n2741 240.244
R14123 GND.n3437 GND.n2741 240.244
R14124 GND.n3437 GND.n2743 240.244
R14125 GND.n3433 GND.n2743 240.244
R14126 GND.n3433 GND.n2749 240.244
R14127 GND.n3429 GND.n2749 240.244
R14128 GND.n3429 GND.n2751 240.244
R14129 GND.n3425 GND.n2751 240.244
R14130 GND.n3425 GND.n2757 240.244
R14131 GND.n3421 GND.n2757 240.244
R14132 GND.n3421 GND.n2759 240.244
R14133 GND.n3417 GND.n2759 240.244
R14134 GND.n3417 GND.n2765 240.244
R14135 GND.n3413 GND.n2765 240.244
R14136 GND.n3413 GND.n2767 240.244
R14137 GND.n3409 GND.n2767 240.244
R14138 GND.n3409 GND.n2773 240.244
R14139 GND.n3405 GND.n2773 240.244
R14140 GND.n3405 GND.n2775 240.244
R14141 GND.n3401 GND.n2775 240.244
R14142 GND.n3401 GND.n2781 240.244
R14143 GND.n3397 GND.n2781 240.244
R14144 GND.n3397 GND.n2783 240.244
R14145 GND.n3393 GND.n2783 240.244
R14146 GND.n3393 GND.n2789 240.244
R14147 GND.n3389 GND.n2789 240.244
R14148 GND.n3389 GND.n2791 240.244
R14149 GND.n3385 GND.n2791 240.244
R14150 GND.n3385 GND.n2797 240.244
R14151 GND.n3381 GND.n2797 240.244
R14152 GND.n3381 GND.n2799 240.244
R14153 GND.n3377 GND.n2799 240.244
R14154 GND.n3377 GND.n2805 240.244
R14155 GND.n3373 GND.n2805 240.244
R14156 GND.n3373 GND.n2807 240.244
R14157 GND.n3369 GND.n2807 240.244
R14158 GND.n3369 GND.n2813 240.244
R14159 GND.n3365 GND.n2813 240.244
R14160 GND.n3365 GND.n2815 240.244
R14161 GND.n3361 GND.n2815 240.244
R14162 GND.n3361 GND.n2821 240.244
R14163 GND.n3357 GND.n2821 240.244
R14164 GND.n3357 GND.n2823 240.244
R14165 GND.n3353 GND.n2823 240.244
R14166 GND.n3353 GND.n2829 240.244
R14167 GND.n3349 GND.n2829 240.244
R14168 GND.n3349 GND.n2831 240.244
R14169 GND.n3345 GND.n2831 240.244
R14170 GND.n3345 GND.n2837 240.244
R14171 GND.n3341 GND.n2837 240.244
R14172 GND.n3341 GND.n2839 240.244
R14173 GND.n3337 GND.n2839 240.244
R14174 GND.n3337 GND.n2845 240.244
R14175 GND.n3333 GND.n2845 240.244
R14176 GND.n3333 GND.n2847 240.244
R14177 GND.n3329 GND.n2847 240.244
R14178 GND.n3329 GND.n2853 240.244
R14179 GND.n3325 GND.n2853 240.244
R14180 GND.n3325 GND.n2855 240.244
R14181 GND.n3321 GND.n2855 240.244
R14182 GND.n3321 GND.n2861 240.244
R14183 GND.n3317 GND.n2861 240.244
R14184 GND.n3317 GND.n2863 240.244
R14185 GND.n3313 GND.n2863 240.244
R14186 GND.n3313 GND.n2869 240.244
R14187 GND.n3309 GND.n2869 240.244
R14188 GND.n3309 GND.n2871 240.244
R14189 GND.n3305 GND.n2871 240.244
R14190 GND.n3305 GND.n2877 240.244
R14191 GND.n3301 GND.n2877 240.244
R14192 GND.n3301 GND.n2879 240.244
R14193 GND.n3297 GND.n2879 240.244
R14194 GND.n3297 GND.n2885 240.244
R14195 GND.n3293 GND.n2885 240.244
R14196 GND.n3293 GND.n2887 240.244
R14197 GND.n3289 GND.n2887 240.244
R14198 GND.n3289 GND.n2893 240.244
R14199 GND.n3285 GND.n2893 240.244
R14200 GND.n3285 GND.n2895 240.244
R14201 GND.n3281 GND.n2895 240.244
R14202 GND.n3281 GND.n2901 240.244
R14203 GND.n3277 GND.n2901 240.244
R14204 GND.n3277 GND.n2903 240.244
R14205 GND.n3273 GND.n2903 240.244
R14206 GND.n3273 GND.n2909 240.244
R14207 GND.n3269 GND.n2909 240.244
R14208 GND.n3269 GND.n2911 240.244
R14209 GND.n3265 GND.n2911 240.244
R14210 GND.n3265 GND.n2917 240.244
R14211 GND.n3261 GND.n2917 240.244
R14212 GND.n3261 GND.n2919 240.244
R14213 GND.n3257 GND.n2919 240.244
R14214 GND.n3257 GND.n2925 240.244
R14215 GND.n3253 GND.n2925 240.244
R14216 GND.n3253 GND.n2927 240.244
R14217 GND.n3249 GND.n2927 240.244
R14218 GND.n3249 GND.n2933 240.244
R14219 GND.n3245 GND.n2933 240.244
R14220 GND.n3245 GND.n2935 240.244
R14221 GND.n3241 GND.n2935 240.244
R14222 GND.n3241 GND.n2941 240.244
R14223 GND.n3237 GND.n2941 240.244
R14224 GND.n3237 GND.n2943 240.244
R14225 GND.n3233 GND.n2943 240.244
R14226 GND.n3233 GND.n2949 240.244
R14227 GND.n3229 GND.n2949 240.244
R14228 GND.n3229 GND.n2951 240.244
R14229 GND.n3225 GND.n2951 240.244
R14230 GND.n3225 GND.n2957 240.244
R14231 GND.n3221 GND.n2957 240.244
R14232 GND.n3221 GND.n2959 240.244
R14233 GND.n3217 GND.n2959 240.244
R14234 GND.n3217 GND.n2965 240.244
R14235 GND.n3213 GND.n2967 240.244
R14236 GND.n2973 GND.n2967 240.244
R14237 GND.n3206 GND.n2973 240.244
R14238 GND.n3206 GND.n2974 240.244
R14239 GND.n3202 GND.n2974 240.244
R14240 GND.n3202 GND.n2977 240.244
R14241 GND.n3198 GND.n2977 240.244
R14242 GND.n3198 GND.n2982 240.244
R14243 GND.n3194 GND.n2982 240.244
R14244 GND.n3194 GND.n2984 240.244
R14245 GND.n3190 GND.n2984 240.244
R14246 GND.n3190 GND.n2990 240.244
R14247 GND.n3186 GND.n2990 240.244
R14248 GND.n3186 GND.n2992 240.244
R14249 GND.n3182 GND.n2992 240.244
R14250 GND.n3182 GND.n2998 240.244
R14251 GND.n3178 GND.n2998 240.244
R14252 GND.n3178 GND.n3000 240.244
R14253 GND.n3174 GND.n3000 240.244
R14254 GND.n3174 GND.n3006 240.244
R14255 GND.n3170 GND.n3006 240.244
R14256 GND.n3170 GND.n3008 240.244
R14257 GND.n3166 GND.n3008 240.244
R14258 GND.n3166 GND.n3014 240.244
R14259 GND.n3162 GND.n3014 240.244
R14260 GND.n3162 GND.n3016 240.244
R14261 GND.n3158 GND.n3016 240.244
R14262 GND.n3158 GND.n3022 240.244
R14263 GND.n3154 GND.n3022 240.244
R14264 GND.n3154 GND.n3024 240.244
R14265 GND.n3150 GND.n3024 240.244
R14266 GND.n3150 GND.n3030 240.244
R14267 GND.n3146 GND.n3030 240.244
R14268 GND.n3146 GND.n3032 240.244
R14269 GND.n3142 GND.n3032 240.244
R14270 GND.n3142 GND.n3038 240.244
R14271 GND.n3138 GND.n3038 240.244
R14272 GND.n3138 GND.n3040 240.244
R14273 GND.n3134 GND.n3040 240.244
R14274 GND.n3134 GND.n3046 240.244
R14275 GND.n3130 GND.n3046 240.244
R14276 GND.n3130 GND.n3048 240.244
R14277 GND.n3126 GND.n3048 240.244
R14278 GND.n3126 GND.n3054 240.244
R14279 GND.n3122 GND.n3054 240.244
R14280 GND.n3122 GND.n3056 240.244
R14281 GND.n3118 GND.n3056 240.244
R14282 GND.n3118 GND.n3062 240.244
R14283 GND.n3114 GND.n3062 240.244
R14284 GND.n3114 GND.n3064 240.244
R14285 GND.n3110 GND.n3064 240.244
R14286 GND.n3110 GND.n3070 240.244
R14287 GND.n3106 GND.n3070 240.244
R14288 GND.n3106 GND.n3072 240.244
R14289 GND.n3102 GND.n3072 240.244
R14290 GND.n3102 GND.n3078 240.244
R14291 GND.n3098 GND.n3078 240.244
R14292 GND.n3098 GND.n3080 240.244
R14293 GND.n3094 GND.n3080 240.244
R14294 GND.n3094 GND.n3086 240.244
R14295 GND.n3090 GND.n3086 240.244
R14296 GND.n3090 GND.n382 240.244
R14297 GND.n8264 GND.n382 240.244
R14298 GND.n4121 GND.n2154 240.244
R14299 GND.n4121 GND.n4120 240.244
R14300 GND.n4120 GND.n4119 240.244
R14301 GND.n4119 GND.n4095 240.244
R14302 GND.n4115 GND.n4095 240.244
R14303 GND.n4115 GND.n4114 240.244
R14304 GND.n4114 GND.n4113 240.244
R14305 GND.n4113 GND.n4101 240.244
R14306 GND.n4109 GND.n4101 240.244
R14307 GND.n4109 GND.n4108 240.244
R14308 GND.n4108 GND.n2062 240.244
R14309 GND.n4434 GND.n2062 240.244
R14310 GND.n4434 GND.n2058 240.244
R14311 GND.n4440 GND.n2058 240.244
R14312 GND.n4441 GND.n4440 240.244
R14313 GND.n4442 GND.n4441 240.244
R14314 GND.n4442 GND.n2053 240.244
R14315 GND.n4450 GND.n2053 240.244
R14316 GND.n4450 GND.n2054 240.244
R14317 GND.n2054 GND.n2000 240.244
R14318 GND.n4516 GND.n2000 240.244
R14319 GND.n4516 GND.n1996 240.244
R14320 GND.n4522 GND.n1996 240.244
R14321 GND.n4523 GND.n4522 240.244
R14322 GND.n4524 GND.n4523 240.244
R14323 GND.n4524 GND.n1991 240.244
R14324 GND.n4568 GND.n1991 240.244
R14325 GND.n4568 GND.n1992 240.244
R14326 GND.n4564 GND.n1992 240.244
R14327 GND.n4564 GND.n4563 240.244
R14328 GND.n4563 GND.n4562 240.244
R14329 GND.n4562 GND.n4532 240.244
R14330 GND.n4536 GND.n4532 240.244
R14331 GND.n4556 GND.n4536 240.244
R14332 GND.n4556 GND.n4555 240.244
R14333 GND.n4555 GND.n4554 240.244
R14334 GND.n4554 GND.n4538 240.244
R14335 GND.n4549 GND.n4538 240.244
R14336 GND.n4549 GND.n4548 240.244
R14337 GND.n4548 GND.n4547 240.244
R14338 GND.n4547 GND.n4541 240.244
R14339 GND.n4541 GND.n1855 240.244
R14340 GND.n4706 GND.n1855 240.244
R14341 GND.n4707 GND.n4706 240.244
R14342 GND.n4708 GND.n4707 240.244
R14343 GND.n4708 GND.n1850 240.244
R14344 GND.n4727 GND.n1850 240.244
R14345 GND.n4727 GND.n1851 240.244
R14346 GND.n4723 GND.n1851 240.244
R14347 GND.n4723 GND.n4722 240.244
R14348 GND.n4722 GND.n4721 240.244
R14349 GND.n4721 GND.n1791 240.244
R14350 GND.n4800 GND.n1791 240.244
R14351 GND.n4801 GND.n4800 240.244
R14352 GND.n4801 GND.n1786 240.244
R14353 GND.n4830 GND.n1786 240.244
R14354 GND.n4830 GND.n1787 240.244
R14355 GND.n4826 GND.n1787 240.244
R14356 GND.n4826 GND.n4825 240.244
R14357 GND.n4825 GND.n4824 240.244
R14358 GND.n4824 GND.n4809 240.244
R14359 GND.n4820 GND.n4809 240.244
R14360 GND.n4820 GND.n4819 240.244
R14361 GND.n4819 GND.n4818 240.244
R14362 GND.n4818 GND.n1709 240.244
R14363 GND.n4931 GND.n1709 240.244
R14364 GND.n4931 GND.n1704 240.244
R14365 GND.n5859 GND.n1704 240.244
R14366 GND.n5859 GND.n1705 240.244
R14367 GND.n5855 GND.n1705 240.244
R14368 GND.n5855 GND.n5854 240.244
R14369 GND.n5854 GND.n5853 240.244
R14370 GND.n5853 GND.n4939 240.244
R14371 GND.n5849 GND.n4939 240.244
R14372 GND.n5849 GND.n5848 240.244
R14373 GND.n5848 GND.n5847 240.244
R14374 GND.n5847 GND.n4945 240.244
R14375 GND.n5843 GND.n4945 240.244
R14376 GND.n5843 GND.n4951 240.244
R14377 GND.n5839 GND.n4951 240.244
R14378 GND.n5839 GND.n4954 240.244
R14379 GND.n5835 GND.n4954 240.244
R14380 GND.n5835 GND.n4960 240.244
R14381 GND.n5825 GND.n4960 240.244
R14382 GND.n5825 GND.n4972 240.244
R14383 GND.n5821 GND.n4972 240.244
R14384 GND.n5821 GND.n4978 240.244
R14385 GND.n5811 GND.n4978 240.244
R14386 GND.n5811 GND.n4990 240.244
R14387 GND.n5807 GND.n4990 240.244
R14388 GND.n5807 GND.n4996 240.244
R14389 GND.n5797 GND.n4996 240.244
R14390 GND.n5797 GND.n5007 240.244
R14391 GND.n5793 GND.n5007 240.244
R14392 GND.n5793 GND.n5013 240.244
R14393 GND.n5783 GND.n5013 240.244
R14394 GND.n5783 GND.n5025 240.244
R14395 GND.n5779 GND.n5025 240.244
R14396 GND.n5779 GND.n5031 240.244
R14397 GND.n5769 GND.n5031 240.244
R14398 GND.n5769 GND.n5043 240.244
R14399 GND.n5765 GND.n5043 240.244
R14400 GND.n5765 GND.n5049 240.244
R14401 GND.n5062 GND.n5049 240.244
R14402 GND.n5754 GND.n5062 240.244
R14403 GND.n5754 GND.n5063 240.244
R14404 GND.n5750 GND.n5063 240.244
R14405 GND.n5750 GND.n5071 240.244
R14406 GND.n5740 GND.n5071 240.244
R14407 GND.n5740 GND.n5082 240.244
R14408 GND.n5736 GND.n5082 240.244
R14409 GND.n5736 GND.n5088 240.244
R14410 GND.n5726 GND.n5088 240.244
R14411 GND.n5726 GND.n5100 240.244
R14412 GND.n5722 GND.n5100 240.244
R14413 GND.n5722 GND.n5106 240.244
R14414 GND.n5712 GND.n5106 240.244
R14415 GND.n5712 GND.n5118 240.244
R14416 GND.n5708 GND.n5118 240.244
R14417 GND.n5708 GND.n5124 240.244
R14418 GND.n5137 GND.n5124 240.244
R14419 GND.n5697 GND.n5137 240.244
R14420 GND.n5697 GND.n5138 240.244
R14421 GND.n5693 GND.n5138 240.244
R14422 GND.n5693 GND.n5146 240.244
R14423 GND.n5683 GND.n5146 240.244
R14424 GND.n5683 GND.n5158 240.244
R14425 GND.n5679 GND.n5158 240.244
R14426 GND.n5679 GND.n5164 240.244
R14427 GND.n5669 GND.n5164 240.244
R14428 GND.n5669 GND.n5176 240.244
R14429 GND.n5665 GND.n5176 240.244
R14430 GND.n5665 GND.n5182 240.244
R14431 GND.n5655 GND.n5182 240.244
R14432 GND.n5655 GND.n1574 240.244
R14433 GND.n6102 GND.n1574 240.244
R14434 GND.n6102 GND.n1570 240.244
R14435 GND.n6108 GND.n1570 240.244
R14436 GND.n6108 GND.n1560 240.244
R14437 GND.n6118 GND.n1560 240.244
R14438 GND.n6118 GND.n1556 240.244
R14439 GND.n6124 GND.n1556 240.244
R14440 GND.n6124 GND.n1543 240.244
R14441 GND.n6143 GND.n1543 240.244
R14442 GND.n6143 GND.n1539 240.244
R14443 GND.n6149 GND.n1539 240.244
R14444 GND.n6149 GND.n1500 240.244
R14445 GND.n6322 GND.n1500 240.244
R14446 GND.n6322 GND.n1496 240.244
R14447 GND.n6328 GND.n1496 240.244
R14448 GND.n6328 GND.n1484 240.244
R14449 GND.n6338 GND.n1484 240.244
R14450 GND.n6338 GND.n1480 240.244
R14451 GND.n6344 GND.n1480 240.244
R14452 GND.n6344 GND.n1468 240.244
R14453 GND.n6354 GND.n1468 240.244
R14454 GND.n6354 GND.n1464 240.244
R14455 GND.n6360 GND.n1464 240.244
R14456 GND.n6360 GND.n1452 240.244
R14457 GND.n6370 GND.n1452 240.244
R14458 GND.n6370 GND.n1448 240.244
R14459 GND.n6376 GND.n1448 240.244
R14460 GND.n6376 GND.n1436 240.244
R14461 GND.n6385 GND.n1436 240.244
R14462 GND.n6385 GND.n1431 240.244
R14463 GND.n6393 GND.n1431 240.244
R14464 GND.n6393 GND.n1432 240.244
R14465 GND.n1432 GND.n1318 240.244
R14466 GND.n6561 GND.n1318 240.244
R14467 GND.n6561 GND.n1314 240.244
R14468 GND.n6567 GND.n1314 240.244
R14469 GND.n6567 GND.n1303 240.244
R14470 GND.n6577 GND.n1303 240.244
R14471 GND.n6577 GND.n1299 240.244
R14472 GND.n6583 GND.n1299 240.244
R14473 GND.n6583 GND.n1287 240.244
R14474 GND.n6593 GND.n1287 240.244
R14475 GND.n6593 GND.n1283 240.244
R14476 GND.n6599 GND.n1283 240.244
R14477 GND.n6599 GND.n1271 240.244
R14478 GND.n6609 GND.n1271 240.244
R14479 GND.n6609 GND.n1267 240.244
R14480 GND.n6615 GND.n1267 240.244
R14481 GND.n6615 GND.n1255 240.244
R14482 GND.n6624 GND.n1255 240.244
R14483 GND.n6624 GND.n1251 240.244
R14484 GND.n6630 GND.n1251 240.244
R14485 GND.n6630 GND.n1239 240.244
R14486 GND.n6640 GND.n1239 240.244
R14487 GND.n6640 GND.n1235 240.244
R14488 GND.n6646 GND.n1235 240.244
R14489 GND.n6646 GND.n1222 240.244
R14490 GND.n6665 GND.n1222 240.244
R14491 GND.n6665 GND.n1218 240.244
R14492 GND.n6671 GND.n1218 240.244
R14493 GND.n6671 GND.n1165 240.244
R14494 GND.n6819 GND.n1165 240.244
R14495 GND.n6819 GND.n1161 240.244
R14496 GND.n6825 GND.n1161 240.244
R14497 GND.n6825 GND.n1149 240.244
R14498 GND.n6835 GND.n1149 240.244
R14499 GND.n6835 GND.n1145 240.244
R14500 GND.n6841 GND.n1145 240.244
R14501 GND.n6841 GND.n1133 240.244
R14502 GND.n6851 GND.n1133 240.244
R14503 GND.n6851 GND.n1129 240.244
R14504 GND.n6857 GND.n1129 240.244
R14505 GND.n6857 GND.n1117 240.244
R14506 GND.n6867 GND.n1117 240.244
R14507 GND.n6867 GND.n1113 240.244
R14508 GND.n6873 GND.n1113 240.244
R14509 GND.n6873 GND.n1100 240.244
R14510 GND.n6887 GND.n1100 240.244
R14511 GND.n6887 GND.n1096 240.244
R14512 GND.n6893 GND.n1096 240.244
R14513 GND.n6893 GND.n1054 240.244
R14514 GND.n6980 GND.n1054 240.244
R14515 GND.n6980 GND.n1049 240.244
R14516 GND.n6991 GND.n1049 240.244
R14517 GND.n6991 GND.n1050 240.244
R14518 GND.n6987 GND.n1050 240.244
R14519 GND.n6987 GND.n1030 240.244
R14520 GND.n7020 GND.n1030 240.244
R14521 GND.n7020 GND.n1025 240.244
R14522 GND.n7037 GND.n1025 240.244
R14523 GND.n7037 GND.n1026 240.244
R14524 GND.n7033 GND.n1026 240.244
R14525 GND.n7033 GND.n7032 240.244
R14526 GND.n7032 GND.n7031 240.244
R14527 GND.n7031 GND.n996 240.244
R14528 GND.n7078 GND.n996 240.244
R14529 GND.n7078 GND.n991 240.244
R14530 GND.n7086 GND.n991 240.244
R14531 GND.n7086 GND.n992 240.244
R14532 GND.n992 GND.n971 240.244
R14533 GND.n7113 GND.n971 240.244
R14534 GND.n7113 GND.n966 240.244
R14535 GND.n7124 GND.n966 240.244
R14536 GND.n7124 GND.n967 240.244
R14537 GND.n7120 GND.n967 240.244
R14538 GND.n7120 GND.n946 240.244
R14539 GND.n7152 GND.n946 240.244
R14540 GND.n7152 GND.n941 240.244
R14541 GND.n7169 GND.n941 240.244
R14542 GND.n7169 GND.n942 240.244
R14543 GND.n7165 GND.n942 240.244
R14544 GND.n7165 GND.n7164 240.244
R14545 GND.n7164 GND.n7163 240.244
R14546 GND.n7163 GND.n914 240.244
R14547 GND.n7212 GND.n914 240.244
R14548 GND.n7212 GND.n909 240.244
R14549 GND.n7238 GND.n909 240.244
R14550 GND.n7238 GND.n910 240.244
R14551 GND.n7234 GND.n910 240.244
R14552 GND.n7234 GND.n7233 240.244
R14553 GND.n7233 GND.n7232 240.244
R14554 GND.n7232 GND.n7220 240.244
R14555 GND.n7228 GND.n7220 240.244
R14556 GND.n7228 GND.n7227 240.244
R14557 GND.n7227 GND.n870 240.244
R14558 GND.n7292 GND.n870 240.244
R14559 GND.n7292 GND.n865 240.244
R14560 GND.n7300 GND.n865 240.244
R14561 GND.n7300 GND.n866 240.244
R14562 GND.n866 GND.n845 240.244
R14563 GND.n7328 GND.n845 240.244
R14564 GND.n7328 GND.n841 240.244
R14565 GND.n7334 GND.n841 240.244
R14566 GND.n7334 GND.n829 240.244
R14567 GND.n7351 GND.n829 240.244
R14568 GND.n7351 GND.n824 240.244
R14569 GND.n7359 GND.n824 240.244
R14570 GND.n7359 GND.n825 240.244
R14571 GND.n825 GND.n805 240.244
R14572 GND.n7443 GND.n805 240.244
R14573 GND.n7443 GND.n800 240.244
R14574 GND.n7533 GND.n800 240.244
R14575 GND.n7533 GND.n801 240.244
R14576 GND.n7529 GND.n801 240.244
R14577 GND.n7529 GND.n7451 240.244
R14578 GND.n7525 GND.n7451 240.244
R14579 GND.n7525 GND.n7453 240.244
R14580 GND.n7521 GND.n7453 240.244
R14581 GND.n7521 GND.n7520 240.244
R14582 GND.n7520 GND.n7519 240.244
R14583 GND.n7519 GND.n7459 240.244
R14584 GND.n7515 GND.n7459 240.244
R14585 GND.n7515 GND.n7514 240.244
R14586 GND.n7514 GND.n7513 240.244
R14587 GND.n7513 GND.n7465 240.244
R14588 GND.n7509 GND.n7465 240.244
R14589 GND.n7509 GND.n7508 240.244
R14590 GND.n7508 GND.n7507 240.244
R14591 GND.n7507 GND.n7471 240.244
R14592 GND.n7503 GND.n7471 240.244
R14593 GND.n7503 GND.n7502 240.244
R14594 GND.n7502 GND.n7501 240.244
R14595 GND.n7501 GND.n7477 240.244
R14596 GND.n7497 GND.n7477 240.244
R14597 GND.n7497 GND.n7496 240.244
R14598 GND.n7496 GND.n7495 240.244
R14599 GND.n7495 GND.n7483 240.244
R14600 GND.n7491 GND.n7483 240.244
R14601 GND.n7491 GND.n7490 240.244
R14602 GND.n7490 GND.n525 240.244
R14603 GND.n7901 GND.n525 240.244
R14604 GND.n7901 GND.n521 240.244
R14605 GND.n7907 GND.n521 240.244
R14606 GND.n7908 GND.n7907 240.244
R14607 GND.n7909 GND.n7908 240.244
R14608 GND.n7909 GND.n516 240.244
R14609 GND.n7935 GND.n516 240.244
R14610 GND.n7935 GND.n517 240.244
R14611 GND.n7931 GND.n517 240.244
R14612 GND.n7931 GND.n7930 240.244
R14613 GND.n7930 GND.n7929 240.244
R14614 GND.n7929 GND.n7917 240.244
R14615 GND.n7924 GND.n7917 240.244
R14616 GND.n7924 GND.n7923 240.244
R14617 GND.n7923 GND.n439 240.244
R14618 GND.n8034 GND.n439 240.244
R14619 GND.n8035 GND.n8034 240.244
R14620 GND.n8035 GND.n436 240.244
R14621 GND.n8121 GND.n436 240.244
R14622 GND.n8121 GND.n437 240.244
R14623 GND.n8116 GND.n437 240.244
R14624 GND.n8116 GND.n8115 240.244
R14625 GND.n8115 GND.n8114 240.244
R14626 GND.n8114 GND.n8040 240.244
R14627 GND.n8110 GND.n8040 240.244
R14628 GND.n8110 GND.n8109 240.244
R14629 GND.n8109 GND.n8108 240.244
R14630 GND.n8108 GND.n8046 240.244
R14631 GND.n8104 GND.n8046 240.244
R14632 GND.n8104 GND.n8103 240.244
R14633 GND.n8103 GND.n8102 240.244
R14634 GND.n8102 GND.n8052 240.244
R14635 GND.n8098 GND.n8052 240.244
R14636 GND.n8098 GND.n8097 240.244
R14637 GND.n8097 GND.n8096 240.244
R14638 GND.n8096 GND.n8058 240.244
R14639 GND.n8092 GND.n8058 240.244
R14640 GND.n8092 GND.n8091 240.244
R14641 GND.n8091 GND.n8090 240.244
R14642 GND.n8090 GND.n8064 240.244
R14643 GND.n8086 GND.n8064 240.244
R14644 GND.n8086 GND.n8085 240.244
R14645 GND.n8085 GND.n8084 240.244
R14646 GND.n8084 GND.n8070 240.244
R14647 GND.n8080 GND.n8070 240.244
R14648 GND.n8080 GND.n8079 240.244
R14649 GND.n8079 GND.n392 240.244
R14650 GND.n8248 GND.n392 240.244
R14651 GND.n8249 GND.n8248 240.244
R14652 GND.n8249 GND.n388 240.244
R14653 GND.n8256 GND.n388 240.244
R14654 GND.n8257 GND.n8256 240.244
R14655 GND.n8258 GND.n8257 240.244
R14656 GND.n8258 GND.n383 240.244
R14657 GND.n3939 GND.n2248 240.244
R14658 GND.n3939 GND.n2244 240.244
R14659 GND.n3945 GND.n2244 240.244
R14660 GND.n3945 GND.n2242 240.244
R14661 GND.n3949 GND.n2242 240.244
R14662 GND.n3949 GND.n2238 240.244
R14663 GND.n3955 GND.n2238 240.244
R14664 GND.n3955 GND.n2236 240.244
R14665 GND.n3959 GND.n2236 240.244
R14666 GND.n3959 GND.n2232 240.244
R14667 GND.n3965 GND.n2232 240.244
R14668 GND.n3965 GND.n2230 240.244
R14669 GND.n3969 GND.n2230 240.244
R14670 GND.n3969 GND.n2226 240.244
R14671 GND.n3975 GND.n2226 240.244
R14672 GND.n3975 GND.n2224 240.244
R14673 GND.n3979 GND.n2224 240.244
R14674 GND.n3979 GND.n2220 240.244
R14675 GND.n3985 GND.n2220 240.244
R14676 GND.n3985 GND.n2218 240.244
R14677 GND.n3989 GND.n2218 240.244
R14678 GND.n3989 GND.n2214 240.244
R14679 GND.n3995 GND.n2214 240.244
R14680 GND.n3995 GND.n2212 240.244
R14681 GND.n3999 GND.n2212 240.244
R14682 GND.n3999 GND.n2208 240.244
R14683 GND.n4005 GND.n2208 240.244
R14684 GND.n4005 GND.n2206 240.244
R14685 GND.n4009 GND.n2206 240.244
R14686 GND.n4009 GND.n2202 240.244
R14687 GND.n4015 GND.n2202 240.244
R14688 GND.n4015 GND.n2200 240.244
R14689 GND.n4019 GND.n2200 240.244
R14690 GND.n4019 GND.n2196 240.244
R14691 GND.n4025 GND.n2196 240.244
R14692 GND.n4025 GND.n2194 240.244
R14693 GND.n4029 GND.n2194 240.244
R14694 GND.n4029 GND.n2190 240.244
R14695 GND.n4035 GND.n2190 240.244
R14696 GND.n4035 GND.n2188 240.244
R14697 GND.n4039 GND.n2188 240.244
R14698 GND.n4039 GND.n2184 240.244
R14699 GND.n4045 GND.n2184 240.244
R14700 GND.n4045 GND.n2182 240.244
R14701 GND.n4049 GND.n2182 240.244
R14702 GND.n4049 GND.n2178 240.244
R14703 GND.n4055 GND.n2178 240.244
R14704 GND.n4055 GND.n2176 240.244
R14705 GND.n4059 GND.n2176 240.244
R14706 GND.n4059 GND.n2172 240.244
R14707 GND.n4065 GND.n2172 240.244
R14708 GND.n4065 GND.n2170 240.244
R14709 GND.n4069 GND.n2170 240.244
R14710 GND.n4069 GND.n2166 240.244
R14711 GND.n4075 GND.n2166 240.244
R14712 GND.n4075 GND.n2164 240.244
R14713 GND.n4079 GND.n2164 240.244
R14714 GND.n4079 GND.n2160 240.244
R14715 GND.n4085 GND.n2160 240.244
R14716 GND.n4085 GND.n2158 240.244
R14717 GND.n4089 GND.n2158 240.244
R14718 GND.n4089 GND.n2153 240.244
R14719 GND.n4127 GND.n2153 240.244
R14720 GND.n4344 GND.n2135 240.244
R14721 GND.n2135 GND.n2124 240.244
R14722 GND.n4335 GND.n2124 240.244
R14723 GND.n4335 GND.n2106 240.244
R14724 GND.n4380 GND.n2106 240.244
R14725 GND.n4380 GND.n2107 240.244
R14726 GND.n2107 GND.n2095 240.244
R14727 GND.n4371 GND.n2095 240.244
R14728 GND.n4371 GND.n2077 240.244
R14729 GND.n4423 GND.n2077 240.244
R14730 GND.n4423 GND.n2078 240.244
R14731 GND.n2078 GND.n2067 240.244
R14732 GND.n2067 GND.n2043 240.244
R14733 GND.n4462 GND.n2043 240.244
R14734 GND.n4462 GND.n2044 240.244
R14735 GND.n2044 GND.n2032 240.244
R14736 GND.n4453 GND.n2032 240.244
R14737 GND.n4453 GND.n2015 240.244
R14738 GND.n4505 GND.n2015 240.244
R14739 GND.n4505 GND.n2016 240.244
R14740 GND.n2016 GND.n2005 240.244
R14741 GND.n2005 GND.n1981 240.244
R14742 GND.n4580 GND.n1981 240.244
R14743 GND.n4580 GND.n1982 240.244
R14744 GND.n1982 GND.n1970 240.244
R14745 GND.n4571 GND.n1970 240.244
R14746 GND.n4571 GND.n1951 240.244
R14747 GND.n4612 GND.n1951 240.244
R14748 GND.n4612 GND.n1952 240.244
R14749 GND.n1952 GND.n1941 240.244
R14750 GND.n1941 GND.n1886 240.244
R14751 GND.n4684 GND.n1886 240.244
R14752 GND.n4684 GND.n1887 240.244
R14753 GND.n4634 GND.n1887 240.244
R14754 GND.n4635 GND.n4634 240.244
R14755 GND.n4635 GND.n1925 240.244
R14756 GND.n1925 GND.n1924 240.244
R14757 GND.n1924 GND.n1910 240.244
R14758 GND.n4658 GND.n1910 240.244
R14759 GND.n4659 GND.n4658 240.244
R14760 GND.n4659 GND.n1867 240.244
R14761 GND.n4664 GND.n1867 240.244
R14762 GND.n4664 GND.n1840 240.244
R14763 GND.n4739 GND.n1840 240.244
R14764 GND.n4739 GND.n1841 240.244
R14765 GND.n1841 GND.n1829 240.244
R14766 GND.n4730 GND.n1829 240.244
R14767 GND.n4730 GND.n1813 240.244
R14768 GND.n4777 GND.n1813 240.244
R14769 GND.n4777 GND.n1814 240.244
R14770 GND.n1814 GND.n1802 240.244
R14771 GND.n4768 GND.n1802 240.244
R14772 GND.n4768 GND.n1779 240.244
R14773 GND.n4845 GND.n1779 240.244
R14774 GND.n4845 GND.n1780 240.244
R14775 GND.n1780 GND.n1768 240.244
R14776 GND.n4836 GND.n1768 240.244
R14777 GND.n4836 GND.n1752 240.244
R14778 GND.n4882 GND.n1752 240.244
R14779 GND.n4882 GND.n1753 240.244
R14780 GND.n1753 GND.n1741 240.244
R14781 GND.n4873 GND.n1741 240.244
R14782 GND.n4873 GND.n1722 240.244
R14783 GND.n4920 GND.n1722 240.244
R14784 GND.n4920 GND.n1723 240.244
R14785 GND.n1723 GND.n1712 240.244
R14786 GND.n1712 GND.n1694 240.244
R14787 GND.n5880 GND.n1694 240.244
R14788 GND.n5880 GND.n1695 240.244
R14789 GND.n1695 GND.n1685 240.244
R14790 GND.n5870 GND.n1685 240.244
R14791 GND.n5870 GND.n1611 240.244
R14792 GND.n6045 GND.n1611 240.244
R14793 GND.n2140 GND.n2139 240.244
R14794 GND.n4153 GND.n2143 240.244
R14795 GND.n2145 GND.n2144 240.244
R14796 GND.n4314 GND.n2151 240.244
R14797 GND.n2132 GND.n2120 240.244
R14798 GND.n4356 GND.n2120 240.244
R14799 GND.n4356 GND.n2115 240.244
R14800 GND.n4363 GND.n2115 240.244
R14801 GND.n4363 GND.n2104 240.244
R14802 GND.n2104 GND.n2091 240.244
R14803 GND.n4392 GND.n2091 240.244
R14804 GND.n4392 GND.n2086 240.244
R14805 GND.n4411 GND.n2086 240.244
R14806 GND.n4411 GND.n2075 240.244
R14807 GND.n4397 GND.n2075 240.244
R14808 GND.n4397 GND.n2065 240.244
R14809 GND.n4400 GND.n2065 240.244
R14810 GND.n4400 GND.n2041 240.244
R14811 GND.n2041 GND.n2028 240.244
R14812 GND.n4474 GND.n2028 240.244
R14813 GND.n4474 GND.n2023 240.244
R14814 GND.n4493 GND.n2023 240.244
R14815 GND.n4493 GND.n2013 240.244
R14816 GND.n4479 GND.n2013 240.244
R14817 GND.n4479 GND.n2003 240.244
R14818 GND.n4482 GND.n2003 240.244
R14819 GND.n4482 GND.n1979 240.244
R14820 GND.n1979 GND.n1966 240.244
R14821 GND.n4592 GND.n1966 240.244
R14822 GND.n4592 GND.n1961 240.244
R14823 GND.n4604 GND.n1961 240.244
R14824 GND.n4604 GND.n1949 240.244
R14825 GND.n4598 GND.n1949 240.244
R14826 GND.n4598 GND.n1936 240.244
R14827 GND.n4625 GND.n1936 240.244
R14828 GND.n4625 GND.n1884 240.244
R14829 GND.n1932 GND.n1884 240.244
R14830 GND.n4632 GND.n1932 240.244
R14831 GND.n4632 GND.n1919 240.244
R14832 GND.n4642 GND.n1919 240.244
R14833 GND.n4642 GND.n1915 240.244
R14834 GND.n4651 GND.n1915 240.244
R14835 GND.n4651 GND.n1912 240.244
R14836 GND.n1912 GND.n1863 240.244
R14837 GND.n4695 GND.n1863 240.244
R14838 GND.n4695 GND.n1859 240.244
R14839 GND.n4703 GND.n1859 240.244
R14840 GND.n4703 GND.n1838 240.244
R14841 GND.n1838 GND.n1826 240.244
R14842 GND.n4751 GND.n1826 240.244
R14843 GND.n4751 GND.n1822 240.244
R14844 GND.n4759 GND.n1822 240.244
R14845 GND.n4759 GND.n1811 240.244
R14846 GND.n1811 GND.n1798 240.244
R14847 GND.n4789 GND.n1798 240.244
R14848 GND.n4789 GND.n1794 240.244
R14849 GND.n4797 GND.n1794 240.244
R14850 GND.n4797 GND.n1777 240.244
R14851 GND.n1777 GND.n1765 240.244
R14852 GND.n4857 GND.n1765 240.244
R14853 GND.n4857 GND.n1761 240.244
R14854 GND.n4865 GND.n1761 240.244
R14855 GND.n4865 GND.n1750 240.244
R14856 GND.n1750 GND.n1737 240.244
R14857 GND.n4894 GND.n1737 240.244
R14858 GND.n4894 GND.n1733 240.244
R14859 GND.n4911 GND.n1733 240.244
R14860 GND.n4911 GND.n1720 240.244
R14861 GND.n4907 GND.n1720 240.244
R14862 GND.n4907 GND.n1711 240.244
R14863 GND.n1711 GND.n1703 240.244
R14864 GND.n1703 GND.n1692 240.244
R14865 GND.n1692 GND.n1681 240.244
R14866 GND.n5891 GND.n1681 240.244
R14867 GND.n5891 GND.n1677 240.244
R14868 GND.n5898 GND.n1677 240.244
R14869 GND.n5898 GND.n1609 240.244
R14870 GND.n1627 GND.n1612 240.244
R14871 GND.n1632 GND.n1629 240.244
R14872 GND.n1636 GND.n1635 240.244
R14873 GND.n1642 GND.n1641 240.244
R14874 GND.n5256 GND.n5255 240.132
R14875 GND.n5254 GND.n5253 240.132
R14876 GND.n788 GND.n787 240.132
R14877 GND.n786 GND.n785 240.132
R14878 GND.n6062 GND.t78 237.815
R14879 GND.n6956 GND.t126 237.815
R14880 GND.n5318 GND.t136 226.552
R14881 GND.n5339 GND.t103 226.552
R14882 GND.n7372 GND.t74 226.552
R14883 GND.n7540 GND.t97 226.552
R14884 GND.n5339 GND.t106 220.841
R14885 GND.n7372 GND.t76 220.841
R14886 GND.n5318 GND.t138 220.837
R14887 GND.n7540 GND.t98 220.837
R14888 GND.n2146 GND.t159 217.078
R14889 GND.n5924 GND.t83 217.078
R14890 GND.n1661 GND.t66 217.078
R14891 GND.n5964 GND.t40 217.078
R14892 GND.n5981 GND.t167 217.078
R14893 GND.n5999 GND.t143 217.078
R14894 GND.n719 GND.t70 217.078
R14895 GND.n730 GND.t61 217.078
R14896 GND.n7604 GND.t49 217.078
R14897 GND.n7616 GND.t150 217.078
R14898 GND.n7628 GND.t93 217.078
R14899 GND.n8344 GND.t44 217.078
R14900 GND.n8333 GND.t95 217.078
R14901 GND.n8323 GND.t57 217.078
R14902 GND.n8412 GND.t134 217.078
R14903 GND.n8302 GND.t152 217.078
R14904 GND.n354 GND.t101 217.078
R14905 GND.n667 GND.t132 217.078
R14906 GND.n4168 GND.t165 217.078
R14907 GND.n4179 GND.t147 217.078
R14908 GND.n4191 GND.t125 217.078
R14909 GND.n4203 GND.t110 217.078
R14910 GND.n4216 GND.t116 217.078
R14911 GND.n1638 GND.t51 217.078
R14912 GND.n2146 GND.t157 210.106
R14913 GND.n5924 GND.t82 210.106
R14914 GND.n1661 GND.t65 210.106
R14915 GND.n5964 GND.t38 210.106
R14916 GND.n5981 GND.t166 210.106
R14917 GND.n5999 GND.t142 210.106
R14918 GND.n719 GND.t68 210.106
R14919 GND.n730 GND.t59 210.106
R14920 GND.n7604 GND.t46 210.106
R14921 GND.n7616 GND.t148 210.106
R14922 GND.n7628 GND.t91 210.106
R14923 GND.n8344 GND.t42 210.106
R14924 GND.n8333 GND.t94 210.106
R14925 GND.n8323 GND.t56 210.106
R14926 GND.n8412 GND.t133 210.106
R14927 GND.n8302 GND.t151 210.106
R14928 GND.n354 GND.t100 210.106
R14929 GND.n667 GND.t130 210.106
R14930 GND.n4168 GND.t163 210.106
R14931 GND.n4179 GND.t145 210.106
R14932 GND.n4191 GND.t123 210.106
R14933 GND.n4203 GND.t107 210.106
R14934 GND.n4216 GND.t114 210.106
R14935 GND.n1638 GND.t50 210.106
R14936 GND.n1657 GND.n1624 199.319
R14937 GND.n72 GND.t198 192.404
R14938 GND.n75 GND.t204 191.386
R14939 GND.n74 GND.t200 191.386
R14940 GND.n73 GND.t202 191.386
R14941 GND.n72 GND.t196 191.386
R14942 GND.n5257 GND.n5252 186.49
R14943 GND.n789 GND.n784 186.49
R14944 GND.n14 GND.n13 185
R14945 GND.n25 GND.n24 185
R14946 GND.n37 GND.n36 185
R14947 GND.n49 GND.n48 185
R14948 GND.n61 GND.n60 185
R14949 GND.n3 GND.n2 185
R14950 GND.n87 GND.n86 185
R14951 GND.n98 GND.n97 185
R14952 GND.n110 GND.n109 185
R14953 GND.n122 GND.n121 185
R14954 GND.n134 GND.n133 185
R14955 GND.n146 GND.n145 185
R14956 GND.t191 GND.n12 167.117
R14957 GND.t237 GND.n23 167.117
R14958 GND.t28 GND.n35 167.117
R14959 GND.t226 GND.n47 167.117
R14960 GND.t184 GND.n59 167.117
R14961 GND.t224 GND.n1 167.117
R14962 GND.t189 GND.n85 167.117
R14963 GND.t230 GND.n96 167.117
R14964 GND.t19 GND.n108 167.117
R14965 GND.t227 GND.n120 167.117
R14966 GND.t188 GND.n132 167.117
R14967 GND.t236 GND.n144 167.117
R14968 GND.n7592 GND.n766 163.367
R14969 GND.n7588 GND.n7587 163.367
R14970 GND.n7584 GND.n7583 163.367
R14971 GND.n7580 GND.n7579 163.367
R14972 GND.n7576 GND.n7575 163.367
R14973 GND.n7572 GND.n7571 163.367
R14974 GND.n7568 GND.n7567 163.367
R14975 GND.n7564 GND.n7563 163.367
R14976 GND.n7560 GND.n7559 163.367
R14977 GND.n7556 GND.n7555 163.367
R14978 GND.n7552 GND.n7551 163.367
R14979 GND.n7547 GND.n7546 163.367
R14980 GND.n7543 GND.n7542 163.367
R14981 GND.n7594 GND.n738 163.367
R14982 GND.n7377 GND.n7376 163.367
R14983 GND.n7381 GND.n7380 163.367
R14984 GND.n7385 GND.n7384 163.367
R14985 GND.n7389 GND.n7388 163.367
R14986 GND.n7393 GND.n7392 163.367
R14987 GND.n7397 GND.n7396 163.367
R14988 GND.n7401 GND.n7400 163.367
R14989 GND.n7405 GND.n7404 163.367
R14990 GND.n7409 GND.n7408 163.367
R14991 GND.n7413 GND.n7412 163.367
R14992 GND.n7417 GND.n7416 163.367
R14993 GND.n7421 GND.n7420 163.367
R14994 GND.n5387 GND.n4963 163.367
R14995 GND.n5391 GND.n4963 163.367
R14996 GND.n5391 GND.n4970 163.367
R14997 GND.n5395 GND.n4970 163.367
R14998 GND.n5400 GND.n5395 163.367
R14999 GND.n5401 GND.n5400 163.367
R15000 GND.n5401 GND.n4980 163.367
R15001 GND.n5404 GND.n4980 163.367
R15002 GND.n5404 GND.n4988 163.367
R15003 GND.n5408 GND.n4988 163.367
R15004 GND.n5413 GND.n5408 163.367
R15005 GND.n5414 GND.n5413 163.367
R15006 GND.n5414 GND.n4998 163.367
R15007 GND.n5418 GND.n4998 163.367
R15008 GND.n5418 GND.n5005 163.367
R15009 GND.n5422 GND.n5005 163.367
R15010 GND.n5427 GND.n5422 163.367
R15011 GND.n5428 GND.n5427 163.367
R15012 GND.n5428 GND.n5015 163.367
R15013 GND.n5431 GND.n5015 163.367
R15014 GND.n5431 GND.n5023 163.367
R15015 GND.n5435 GND.n5023 163.367
R15016 GND.n5440 GND.n5435 163.367
R15017 GND.n5441 GND.n5440 163.367
R15018 GND.n5441 GND.n5033 163.367
R15019 GND.n5444 GND.n5033 163.367
R15020 GND.n5444 GND.n5041 163.367
R15021 GND.n5448 GND.n5041 163.367
R15022 GND.n5453 GND.n5448 163.367
R15023 GND.n5454 GND.n5453 163.367
R15024 GND.n5454 GND.n5051 163.367
R15025 GND.n5458 GND.n5051 163.367
R15026 GND.n5458 GND.n5059 163.367
R15027 GND.n5060 GND.n5059 163.367
R15028 GND.n5463 GND.n5060 163.367
R15029 GND.n5470 GND.n5463 163.367
R15030 GND.n5471 GND.n5470 163.367
R15031 GND.n5471 GND.n5073 163.367
R15032 GND.n5474 GND.n5073 163.367
R15033 GND.n5474 GND.n5081 163.367
R15034 GND.n5478 GND.n5081 163.367
R15035 GND.n5484 GND.n5478 163.367
R15036 GND.n5485 GND.n5484 163.367
R15037 GND.n5485 GND.n5090 163.367
R15038 GND.n5488 GND.n5090 163.367
R15039 GND.n5488 GND.n5098 163.367
R15040 GND.n5492 GND.n5098 163.367
R15041 GND.n5497 GND.n5492 163.367
R15042 GND.n5498 GND.n5497 163.367
R15043 GND.n5498 GND.n5108 163.367
R15044 GND.n5501 GND.n5108 163.367
R15045 GND.n5501 GND.n5116 163.367
R15046 GND.n5505 GND.n5116 163.367
R15047 GND.n5510 GND.n5505 163.367
R15048 GND.n5511 GND.n5510 163.367
R15049 GND.n5511 GND.n5126 163.367
R15050 GND.n5515 GND.n5126 163.367
R15051 GND.n5515 GND.n5134 163.367
R15052 GND.n5135 GND.n5134 163.367
R15053 GND.n5520 GND.n5135 163.367
R15054 GND.n5527 GND.n5520 163.367
R15055 GND.n5528 GND.n5527 163.367
R15056 GND.n5528 GND.n5148 163.367
R15057 GND.n5531 GND.n5148 163.367
R15058 GND.n5531 GND.n5156 163.367
R15059 GND.n5535 GND.n5156 163.367
R15060 GND.n5540 GND.n5535 163.367
R15061 GND.n5541 GND.n5540 163.367
R15062 GND.n5541 GND.n5166 163.367
R15063 GND.n5544 GND.n5166 163.367
R15064 GND.n5544 GND.n5174 163.367
R15065 GND.n5548 GND.n5174 163.367
R15066 GND.n5553 GND.n5548 163.367
R15067 GND.n5554 GND.n5553 163.367
R15068 GND.n5554 GND.n5184 163.367
R15069 GND.n5557 GND.n5184 163.367
R15070 GND.n5557 GND.n5192 163.367
R15071 GND.n5193 GND.n5192 163.367
R15072 GND.n5194 GND.n5193 163.367
R15073 GND.n5205 GND.n5194 163.367
R15074 GND.n5564 GND.n5205 163.367
R15075 GND.n5565 GND.n5564 163.367
R15076 GND.n5566 GND.n5565 163.367
R15077 GND.n5566 GND.n5202 163.367
R15078 GND.n5636 GND.n5202 163.367
R15079 GND.n5636 GND.n5203 163.367
R15080 GND.n5632 GND.n5203 163.367
R15081 GND.n5632 GND.n5570 163.367
R15082 GND.n5577 GND.n5570 163.367
R15083 GND.n5589 GND.n5577 163.367
R15084 GND.n5589 GND.n5578 163.367
R15085 GND.n5585 GND.n5578 163.367
R15086 GND.n5585 GND.n5584 163.367
R15087 GND.n5584 GND.n1536 163.367
R15088 GND.n1536 GND.n1529 163.367
R15089 GND.n6158 GND.n1529 163.367
R15090 GND.n6159 GND.n6158 163.367
R15091 GND.n6159 GND.n1504 163.367
R15092 GND.n6163 GND.n1504 163.367
R15093 GND.n6164 GND.n6163 163.367
R15094 GND.n6165 GND.n6164 163.367
R15095 GND.n6165 GND.n1512 163.367
R15096 GND.n6169 GND.n1512 163.367
R15097 GND.n6170 GND.n6169 163.367
R15098 GND.n6170 GND.n1518 163.367
R15099 GND.n6173 GND.n1518 163.367
R15100 GND.n6173 GND.n1525 163.367
R15101 GND.n6297 GND.n1525 163.367
R15102 GND.n6297 GND.n1526 163.367
R15103 GND.n6293 GND.n1526 163.367
R15104 GND.n6293 GND.n6292 163.367
R15105 GND.n6292 GND.n6177 163.367
R15106 GND.n6186 GND.n6177 163.367
R15107 GND.n6283 GND.n6186 163.367
R15108 GND.n6283 GND.n6187 163.367
R15109 GND.n6279 GND.n6187 163.367
R15110 GND.n6279 GND.n6278 163.367
R15111 GND.n6278 GND.n6191 163.367
R15112 GND.n6200 GND.n6191 163.367
R15113 GND.n6269 GND.n6200 163.367
R15114 GND.n6269 GND.n6201 163.367
R15115 GND.n6265 GND.n6201 163.367
R15116 GND.n6265 GND.n6264 163.367
R15117 GND.n6264 GND.n6205 163.367
R15118 GND.n6246 GND.n6205 163.367
R15119 GND.n6255 GND.n6246 163.367
R15120 GND.n6255 GND.n6247 163.367
R15121 GND.n6251 GND.n6247 163.367
R15122 GND.n6251 GND.n1322 163.367
R15123 GND.n1330 GND.n1322 163.367
R15124 GND.n6553 GND.n1330 163.367
R15125 GND.n6553 GND.n1331 163.367
R15126 GND.n6549 GND.n1331 163.367
R15127 GND.n6549 GND.n1334 163.367
R15128 GND.n1340 GND.n1334 163.367
R15129 GND.n6540 GND.n1340 163.367
R15130 GND.n6540 GND.n1341 163.367
R15131 GND.n6536 GND.n1341 163.367
R15132 GND.n6536 GND.n6535 163.367
R15133 GND.n6535 GND.n1344 163.367
R15134 GND.n1352 GND.n1344 163.367
R15135 GND.n6526 GND.n1352 163.367
R15136 GND.n6526 GND.n1353 163.367
R15137 GND.n6522 GND.n1353 163.367
R15138 GND.n6522 GND.n6521 163.367
R15139 GND.n6521 GND.n1357 163.367
R15140 GND.n1366 GND.n1357 163.367
R15141 GND.n6512 GND.n1366 163.367
R15142 GND.n6512 GND.n1367 163.367
R15143 GND.n6508 GND.n1367 163.367
R15144 GND.n6508 GND.n6507 163.367
R15145 GND.n6507 GND.n1371 163.367
R15146 GND.n1380 GND.n1371 163.367
R15147 GND.n6498 GND.n1380 163.367
R15148 GND.n6498 GND.n1381 163.367
R15149 GND.n6494 GND.n1381 163.367
R15150 GND.n6494 GND.n6493 163.367
R15151 GND.n6493 GND.n6492 163.367
R15152 GND.n6492 GND.n1385 163.367
R15153 GND.n6488 GND.n1385 163.367
R15154 GND.n6488 GND.n6487 163.367
R15155 GND.n6487 GND.n6486 163.367
R15156 GND.n6486 GND.n1387 163.367
R15157 GND.n1393 GND.n1387 163.367
R15158 GND.n1393 GND.n1392 163.367
R15159 GND.n1392 GND.n1215 163.367
R15160 GND.n1215 GND.n1208 163.367
R15161 GND.n6680 GND.n1208 163.367
R15162 GND.n6681 GND.n6680 163.367
R15163 GND.n6681 GND.n1169 163.367
R15164 GND.n6685 GND.n1169 163.367
R15165 GND.n6686 GND.n6685 163.367
R15166 GND.n6687 GND.n6686 163.367
R15167 GND.n6687 GND.n1177 163.367
R15168 GND.n6691 GND.n1177 163.367
R15169 GND.n6692 GND.n6691 163.367
R15170 GND.n6692 GND.n1183 163.367
R15171 GND.n6696 GND.n1183 163.367
R15172 GND.n6697 GND.n6696 163.367
R15173 GND.n6697 GND.n1190 163.367
R15174 GND.n6701 GND.n1190 163.367
R15175 GND.n6702 GND.n6701 163.367
R15176 GND.n6702 GND.n1196 163.367
R15177 GND.n6705 GND.n1196 163.367
R15178 GND.n6705 GND.n1204 163.367
R15179 GND.n6780 GND.n1204 163.367
R15180 GND.n6780 GND.n1205 163.367
R15181 GND.n6776 GND.n1205 163.367
R15182 GND.n6776 GND.n6775 163.367
R15183 GND.n6775 GND.n6709 163.367
R15184 GND.n6742 GND.n6709 163.367
R15185 GND.n6766 GND.n6742 163.367
R15186 GND.n6766 GND.n6743 163.367
R15187 GND.n6762 GND.n6743 163.367
R15188 GND.n6762 GND.n6761 163.367
R15189 GND.n6761 GND.n1094 163.367
R15190 GND.n6757 GND.n1094 163.367
R15191 GND.n6757 GND.n1088 163.367
R15192 GND.n6754 GND.n1088 163.367
R15193 GND.n6754 GND.n6753 163.367
R15194 GND.n6753 GND.n6752 163.367
R15195 GND.n6752 GND.n1046 163.367
R15196 GND.n6748 GND.n1046 163.367
R15197 GND.n6748 GND.n1040 163.367
R15198 GND.n7001 GND.n1040 163.367
R15199 GND.n7001 GND.n1038 163.367
R15200 GND.n7009 GND.n1038 163.367
R15201 GND.n7009 GND.n1032 163.367
R15202 GND.n7005 GND.n1032 163.367
R15203 GND.n7005 GND.n1024 163.367
R15204 GND.n1024 GND.n1016 163.367
R15205 GND.n7046 GND.n1016 163.367
R15206 GND.n7046 GND.n1014 163.367
R15207 GND.n7050 GND.n1014 163.367
R15208 GND.n7050 GND.n1007 163.367
R15209 GND.n7059 GND.n1007 163.367
R15210 GND.n7059 GND.n1004 163.367
R15211 GND.n7068 GND.n1004 163.367
R15212 GND.n7068 GND.n1005 163.367
R15213 GND.n1005 GND.n998 163.367
R15214 GND.n7063 GND.n998 163.367
R15215 GND.n7063 GND.n990 163.367
R15216 GND.n990 GND.n982 163.367
R15217 GND.n7095 GND.n982 163.367
R15218 GND.n7095 GND.n979 163.367
R15219 GND.n7104 GND.n979 163.367
R15220 GND.n7104 GND.n980 163.367
R15221 GND.n980 GND.n973 163.367
R15222 GND.n7099 GND.n973 163.367
R15223 GND.n7099 GND.n964 163.367
R15224 GND.n964 GND.n957 163.367
R15225 GND.n7133 GND.n957 163.367
R15226 GND.n7133 GND.n954 163.367
R15227 GND.n7142 GND.n954 163.367
R15228 GND.n7142 GND.n955 163.367
R15229 GND.n955 GND.n948 163.367
R15230 GND.n7137 GND.n948 163.367
R15231 GND.n7137 GND.n940 163.367
R15232 GND.n940 GND.n932 163.367
R15233 GND.n7178 GND.n932 163.367
R15234 GND.n7178 GND.n930 163.367
R15235 GND.n7183 GND.n930 163.367
R15236 GND.n7183 GND.n923 163.367
R15237 GND.n7192 GND.n923 163.367
R15238 GND.n7193 GND.n7192 163.367
R15239 GND.n7193 GND.n921 163.367
R15240 GND.n7201 GND.n921 163.367
R15241 GND.n7201 GND.n915 163.367
R15242 GND.n7197 GND.n915 163.367
R15243 GND.n7197 GND.n908 163.367
R15244 GND.n908 GND.n900 163.367
R15245 GND.n7247 GND.n900 163.367
R15246 GND.n7247 GND.n898 163.367
R15247 GND.n7251 GND.n898 163.367
R15248 GND.n7251 GND.n890 163.367
R15249 GND.n7260 GND.n890 163.367
R15250 GND.n7260 GND.n888 163.367
R15251 GND.n7264 GND.n888 163.367
R15252 GND.n7264 GND.n881 163.367
R15253 GND.n7273 GND.n881 163.367
R15254 GND.n7273 GND.n878 163.367
R15255 GND.n7282 GND.n878 163.367
R15256 GND.n7282 GND.n879 163.367
R15257 GND.n879 GND.n872 163.367
R15258 GND.n7277 GND.n872 163.367
R15259 GND.n7277 GND.n864 163.367
R15260 GND.n864 GND.n856 163.367
R15261 GND.n7309 GND.n856 163.367
R15262 GND.n7309 GND.n853 163.367
R15263 GND.n7319 GND.n853 163.367
R15264 GND.n7319 GND.n854 163.367
R15265 GND.n854 GND.n847 163.367
R15266 GND.n7314 GND.n847 163.367
R15267 GND.n7314 GND.n839 163.367
R15268 GND.n839 GND.n833 163.367
R15269 GND.n7344 GND.n833 163.367
R15270 GND.n7344 GND.n831 163.367
R15271 GND.n7349 GND.n831 163.367
R15272 GND.n7349 GND.n823 163.367
R15273 GND.n823 GND.n816 163.367
R15274 GND.n7369 GND.n816 163.367
R15275 GND.n7369 GND.n813 163.367
R15276 GND.n7434 GND.n813 163.367
R15277 GND.n7434 GND.n814 163.367
R15278 GND.n814 GND.n807 163.367
R15279 GND.n7429 GND.n807 163.367
R15280 GND.n7429 GND.n799 163.367
R15281 GND.n7426 GND.n799 163.367
R15282 GND.n5281 GND.n5280 163.367
R15283 GND.n5283 GND.n5281 163.367
R15284 GND.n5287 GND.n5243 163.367
R15285 GND.n5291 GND.n5289 163.367
R15286 GND.n5295 GND.n5241 163.367
R15287 GND.n5299 GND.n5297 163.367
R15288 GND.n5303 GND.n5239 163.367
R15289 GND.n5307 GND.n5305 163.367
R15290 GND.n5311 GND.n5237 163.367
R15291 GND.n5315 GND.n5313 163.367
R15292 GND.n5322 GND.n5235 163.367
R15293 GND.n5326 GND.n5324 163.367
R15294 GND.n5330 GND.n5233 163.367
R15295 GND.n5336 GND.n5334 163.367
R15296 GND.n5343 GND.n5230 163.367
R15297 GND.n5347 GND.n5345 163.367
R15298 GND.n5351 GND.n5228 163.367
R15299 GND.n5355 GND.n5353 163.367
R15300 GND.n5359 GND.n5226 163.367
R15301 GND.n5363 GND.n5361 163.367
R15302 GND.n5367 GND.n5224 163.367
R15303 GND.n5371 GND.n5369 163.367
R15304 GND.n5375 GND.n5222 163.367
R15305 GND.n5379 GND.n5377 163.367
R15306 GND.n5383 GND.n5220 163.367
R15307 GND.n5386 GND.n5385 163.367
R15308 GND.n5832 GND.n4964 163.367
R15309 GND.n5832 GND.n4965 163.367
R15310 GND.n5828 GND.n4965 163.367
R15311 GND.n5828 GND.n4968 163.367
R15312 GND.n5398 GND.n4968 163.367
R15313 GND.n5398 GND.n4982 163.367
R15314 GND.n5818 GND.n4982 163.367
R15315 GND.n5818 GND.n4983 163.367
R15316 GND.n5814 GND.n4983 163.367
R15317 GND.n5814 GND.n4986 163.367
R15318 GND.n5411 GND.n4986 163.367
R15319 GND.n5411 GND.n5000 163.367
R15320 GND.n5804 GND.n5000 163.367
R15321 GND.n5804 GND.n5001 163.367
R15322 GND.n5800 GND.n5001 163.367
R15323 GND.n5800 GND.n5004 163.367
R15324 GND.n5425 GND.n5004 163.367
R15325 GND.n5425 GND.n5017 163.367
R15326 GND.n5790 GND.n5017 163.367
R15327 GND.n5790 GND.n5018 163.367
R15328 GND.n5786 GND.n5018 163.367
R15329 GND.n5786 GND.n5021 163.367
R15330 GND.n5438 GND.n5021 163.367
R15331 GND.n5438 GND.n5035 163.367
R15332 GND.n5776 GND.n5035 163.367
R15333 GND.n5776 GND.n5036 163.367
R15334 GND.n5772 GND.n5036 163.367
R15335 GND.n5772 GND.n5039 163.367
R15336 GND.n5451 GND.n5039 163.367
R15337 GND.n5451 GND.n5053 163.367
R15338 GND.n5762 GND.n5053 163.367
R15339 GND.n5762 GND.n5054 163.367
R15340 GND.n5758 GND.n5054 163.367
R15341 GND.n5758 GND.n5057 163.367
R15342 GND.n5465 GND.n5057 163.367
R15343 GND.n5468 GND.n5465 163.367
R15344 GND.n5468 GND.n5075 163.367
R15345 GND.n5747 GND.n5075 163.367
R15346 GND.n5747 GND.n5076 163.367
R15347 GND.n5743 GND.n5076 163.367
R15348 GND.n5743 GND.n5079 163.367
R15349 GND.n5482 GND.n5079 163.367
R15350 GND.n5482 GND.n5092 163.367
R15351 GND.n5733 GND.n5092 163.367
R15352 GND.n5733 GND.n5093 163.367
R15353 GND.n5729 GND.n5093 163.367
R15354 GND.n5729 GND.n5096 163.367
R15355 GND.n5495 GND.n5096 163.367
R15356 GND.n5495 GND.n5110 163.367
R15357 GND.n5719 GND.n5110 163.367
R15358 GND.n5719 GND.n5111 163.367
R15359 GND.n5715 GND.n5111 163.367
R15360 GND.n5715 GND.n5114 163.367
R15361 GND.n5508 GND.n5114 163.367
R15362 GND.n5508 GND.n5128 163.367
R15363 GND.n5705 GND.n5128 163.367
R15364 GND.n5705 GND.n5129 163.367
R15365 GND.n5701 GND.n5129 163.367
R15366 GND.n5701 GND.n5132 163.367
R15367 GND.n5522 GND.n5132 163.367
R15368 GND.n5525 GND.n5522 163.367
R15369 GND.n5525 GND.n5149 163.367
R15370 GND.n5690 GND.n5149 163.367
R15371 GND.n5690 GND.n5150 163.367
R15372 GND.n5686 GND.n5150 163.367
R15373 GND.n5686 GND.n5153 163.367
R15374 GND.n5538 GND.n5153 163.367
R15375 GND.n5538 GND.n5168 163.367
R15376 GND.n5676 GND.n5168 163.367
R15377 GND.n5676 GND.n5169 163.367
R15378 GND.n5672 GND.n5169 163.367
R15379 GND.n5672 GND.n5172 163.367
R15380 GND.n5551 GND.n5172 163.367
R15381 GND.n5551 GND.n5186 163.367
R15382 GND.n5662 GND.n5186 163.367
R15383 GND.n5662 GND.n5187 163.367
R15384 GND.n5658 GND.n5187 163.367
R15385 GND.n5658 GND.n5190 163.367
R15386 GND.n5648 GND.n5190 163.367
R15387 GND.n5648 GND.n5195 163.367
R15388 GND.n5644 GND.n5195 163.367
R15389 GND.n5644 GND.n5643 163.367
R15390 GND.n5643 GND.n5642 163.367
R15391 GND.n5642 GND.n5197 163.367
R15392 GND.n5638 GND.n5197 163.367
R15393 GND.n5638 GND.n5199 163.367
R15394 GND.n5630 GND.n5199 163.367
R15395 GND.n5630 GND.n5571 163.367
R15396 GND.n5626 GND.n5571 163.367
R15397 GND.n5626 GND.n5625 163.367
R15398 GND.n5625 GND.n5576 163.367
R15399 GND.n5576 GND.n5573 163.367
R15400 GND.n5573 GND.n1534 163.367
R15401 GND.n6152 GND.n1534 163.367
R15402 GND.n6152 GND.n1532 163.367
R15403 GND.n6156 GND.n1532 163.367
R15404 GND.n6156 GND.n1506 163.367
R15405 GND.n6320 GND.n1506 163.367
R15406 GND.n6320 GND.n1507 163.367
R15407 GND.n6316 GND.n1507 163.367
R15408 GND.n6316 GND.n6315 163.367
R15409 GND.n6315 GND.n6314 163.367
R15410 GND.n6314 GND.n1510 163.367
R15411 GND.n1519 GND.n1510 163.367
R15412 GND.n6304 GND.n1519 163.367
R15413 GND.n6304 GND.n1520 163.367
R15414 GND.n6300 GND.n1520 163.367
R15415 GND.n6300 GND.n6299 163.367
R15416 GND.n6299 GND.n1524 163.367
R15417 GND.n6179 GND.n1524 163.367
R15418 GND.n6290 GND.n6179 163.367
R15419 GND.n6290 GND.n6180 163.367
R15420 GND.n6286 GND.n6180 163.367
R15421 GND.n6286 GND.n6285 163.367
R15422 GND.n6285 GND.n6184 163.367
R15423 GND.n6193 GND.n6184 163.367
R15424 GND.n6276 GND.n6193 163.367
R15425 GND.n6276 GND.n6194 163.367
R15426 GND.n6272 GND.n6194 163.367
R15427 GND.n6272 GND.n6271 163.367
R15428 GND.n6271 GND.n6198 163.367
R15429 GND.n6238 GND.n6198 163.367
R15430 GND.n6262 GND.n6238 163.367
R15431 GND.n6262 GND.n6239 163.367
R15432 GND.n6258 GND.n6239 163.367
R15433 GND.n6258 GND.n6257 163.367
R15434 GND.n6257 GND.n6244 163.367
R15435 GND.n6244 GND.n1324 163.367
R15436 GND.n6559 GND.n1324 163.367
R15437 GND.n6559 GND.n1325 163.367
R15438 GND.n6555 GND.n1325 163.367
R15439 GND.n6555 GND.n1328 163.367
R15440 GND.n6547 GND.n1328 163.367
R15441 GND.n6547 GND.n1336 163.367
R15442 GND.n6543 GND.n1336 163.367
R15443 GND.n6543 GND.n6542 163.367
R15444 GND.n6542 GND.n1338 163.367
R15445 GND.n1345 GND.n1338 163.367
R15446 GND.n6533 GND.n1345 163.367
R15447 GND.n6533 GND.n1346 163.367
R15448 GND.n6529 GND.n1346 163.367
R15449 GND.n6529 GND.n6528 163.367
R15450 GND.n6528 GND.n1350 163.367
R15451 GND.n1359 GND.n1350 163.367
R15452 GND.n6519 GND.n1359 163.367
R15453 GND.n6519 GND.n1360 163.367
R15454 GND.n6515 GND.n1360 163.367
R15455 GND.n6515 GND.n6514 163.367
R15456 GND.n6514 GND.n1364 163.367
R15457 GND.n1373 GND.n1364 163.367
R15458 GND.n6505 GND.n1373 163.367
R15459 GND.n6505 GND.n1374 163.367
R15460 GND.n6501 GND.n1374 163.367
R15461 GND.n6501 GND.n6500 163.367
R15462 GND.n6500 GND.n1378 163.367
R15463 GND.n1403 GND.n1378 163.367
R15464 GND.n1403 GND.n1401 163.367
R15465 GND.n1407 GND.n1401 163.367
R15466 GND.n6476 GND.n1407 163.367
R15467 GND.n6477 GND.n6476 163.367
R15468 GND.n6477 GND.n1398 163.367
R15469 GND.n6484 GND.n1398 163.367
R15470 GND.n6484 GND.n1399 163.367
R15471 GND.n6480 GND.n1399 163.367
R15472 GND.n6480 GND.n1213 163.367
R15473 GND.n6674 GND.n1213 163.367
R15474 GND.n6674 GND.n1211 163.367
R15475 GND.n6678 GND.n1211 163.367
R15476 GND.n6678 GND.n1171 163.367
R15477 GND.n6817 GND.n1171 163.367
R15478 GND.n6817 GND.n1172 163.367
R15479 GND.n6813 GND.n1172 163.367
R15480 GND.n6813 GND.n6812 163.367
R15481 GND.n6812 GND.n6811 163.367
R15482 GND.n6811 GND.n1175 163.367
R15483 GND.n1184 GND.n1175 163.367
R15484 GND.n6801 GND.n1184 163.367
R15485 GND.n6801 GND.n1185 163.367
R15486 GND.n6797 GND.n1185 163.367
R15487 GND.n6797 GND.n6796 163.367
R15488 GND.n6796 GND.n1189 163.367
R15489 GND.n1197 GND.n1189 163.367
R15490 GND.n6787 GND.n1197 163.367
R15491 GND.n6787 GND.n1198 163.367
R15492 GND.n6783 GND.n1198 163.367
R15493 GND.n6783 GND.n6782 163.367
R15494 GND.n6782 GND.n1202 163.367
R15495 GND.n6711 GND.n1202 163.367
R15496 GND.n6773 GND.n6711 163.367
R15497 GND.n6773 GND.n6712 163.367
R15498 GND.n6769 GND.n6712 163.367
R15499 GND.n6769 GND.n6768 163.367
R15500 GND.n6768 GND.n6719 163.367
R15501 GND.n6719 GND.n6716 163.367
R15502 GND.n6716 GND.n1092 163.367
R15503 GND.n6896 GND.n1092 163.367
R15504 GND.n6896 GND.n1089 163.367
R15505 GND.n6903 GND.n1089 163.367
R15506 GND.n6903 GND.n1090 163.367
R15507 GND.n6899 GND.n1090 163.367
R15508 GND.n6899 GND.n1044 163.367
R15509 GND.n6994 GND.n1044 163.367
R15510 GND.n6994 GND.n1042 163.367
R15511 GND.n6998 GND.n1042 163.367
R15512 GND.n6998 GND.n1036 163.367
R15513 GND.n7013 GND.n1036 163.367
R15514 GND.n7013 GND.n1034 163.367
R15515 GND.n7017 GND.n1034 163.367
R15516 GND.n7017 GND.n1022 163.367
R15517 GND.n7040 GND.n1022 163.367
R15518 GND.n7040 GND.n1020 163.367
R15519 GND.n7044 GND.n1020 163.367
R15520 GND.n7044 GND.n1012 163.367
R15521 GND.n7053 GND.n1012 163.367
R15522 GND.n7053 GND.n1010 163.367
R15523 GND.n7057 GND.n1010 163.367
R15524 GND.n7057 GND.n1002 163.367
R15525 GND.n7071 GND.n1002 163.367
R15526 GND.n7071 GND.n1000 163.367
R15527 GND.n7075 GND.n1000 163.367
R15528 GND.n7075 GND.n988 163.367
R15529 GND.n7089 GND.n988 163.367
R15530 GND.n7089 GND.n986 163.367
R15531 GND.n7093 GND.n986 163.367
R15532 GND.n7093 GND.n977 163.367
R15533 GND.n7106 GND.n977 163.367
R15534 GND.n7106 GND.n975 163.367
R15535 GND.n7110 GND.n975 163.367
R15536 GND.n7110 GND.n962 163.367
R15537 GND.n7127 GND.n962 163.367
R15538 GND.n7127 GND.n960 163.367
R15539 GND.n7131 GND.n960 163.367
R15540 GND.n7131 GND.n952 163.367
R15541 GND.n7145 GND.n952 163.367
R15542 GND.n7145 GND.n950 163.367
R15543 GND.n7149 GND.n950 163.367
R15544 GND.n7149 GND.n938 163.367
R15545 GND.n7172 GND.n938 163.367
R15546 GND.n7172 GND.n936 163.367
R15547 GND.n7176 GND.n936 163.367
R15548 GND.n7176 GND.n928 163.367
R15549 GND.n7186 GND.n928 163.367
R15550 GND.n7186 GND.n926 163.367
R15551 GND.n7190 GND.n926 163.367
R15552 GND.n7190 GND.n919 163.367
R15553 GND.n7205 GND.n919 163.367
R15554 GND.n7205 GND.n917 163.367
R15555 GND.n7209 GND.n917 163.367
R15556 GND.n7209 GND.n906 163.367
R15557 GND.n7241 GND.n906 163.367
R15558 GND.n7241 GND.n904 163.367
R15559 GND.n7245 GND.n904 163.367
R15560 GND.n7245 GND.n896 163.367
R15561 GND.n7254 GND.n896 163.367
R15562 GND.n7254 GND.n894 163.367
R15563 GND.n7258 GND.n894 163.367
R15564 GND.n7258 GND.n886 163.367
R15565 GND.n7267 GND.n886 163.367
R15566 GND.n7267 GND.n884 163.367
R15567 GND.n7271 GND.n884 163.367
R15568 GND.n7271 GND.n876 163.367
R15569 GND.n7285 GND.n876 163.367
R15570 GND.n7285 GND.n874 163.367
R15571 GND.n7289 GND.n874 163.367
R15572 GND.n7289 GND.n862 163.367
R15573 GND.n7303 GND.n862 163.367
R15574 GND.n7303 GND.n860 163.367
R15575 GND.n7307 GND.n860 163.367
R15576 GND.n7307 GND.n851 163.367
R15577 GND.n7321 GND.n851 163.367
R15578 GND.n7321 GND.n849 163.367
R15579 GND.n7325 GND.n849 163.367
R15580 GND.n7325 GND.n838 163.367
R15581 GND.n7337 GND.n838 163.367
R15582 GND.n7337 GND.n835 163.367
R15583 GND.n7342 GND.n835 163.367
R15584 GND.n7342 GND.n836 163.367
R15585 GND.n836 GND.n821 163.367
R15586 GND.n7363 GND.n821 163.367
R15587 GND.n7363 GND.n819 163.367
R15588 GND.n7367 GND.n819 163.367
R15589 GND.n7367 GND.n811 163.367
R15590 GND.n7436 GND.n811 163.367
R15591 GND.n7436 GND.n809 163.367
R15592 GND.n7440 GND.n809 163.367
R15593 GND.n7440 GND.n797 163.367
R15594 GND.n7536 GND.n797 163.367
R15595 GND.n7536 GND.n765 163.367
R15596 GND.n795 GND.n794 157.237
R15597 GND.n5262 GND.n5261 152
R15598 GND.n5263 GND.n5250 152
R15599 GND.n5265 GND.n5264 152
R15600 GND.n5268 GND.n5267 152
R15601 GND.n5269 GND.n5248 152
R15602 GND.n5271 GND.n5270 152
R15603 GND.n5273 GND.n5246 152
R15604 GND.n5275 GND.n5274 152
R15605 GND.n793 GND.n767 152
R15606 GND.n783 GND.n768 152
R15607 GND.n782 GND.n781 152
R15608 GND.n780 GND.n769 152
R15609 GND.n777 GND.n770 152
R15610 GND.n776 GND.n775 152
R15611 GND.n774 GND.n771 152
R15612 GND.n772 GND.t139 149.72
R15613 GND.n5319 GND.n5318 149.528
R15614 GND.n5340 GND.n5339 149.528
R15615 GND.n7373 GND.n7372 149.528
R15616 GND.n7541 GND.n7540 149.528
R15617 GND.n7595 GND.n737 143.351
R15618 GND.n5332 GND.n5331 143.351
R15619 GND.n5333 GND.n5332 143.351
R15620 GND.n5259 GND.t71 129.018
R15621 GND.n5274 GND.t117 126.766
R15622 GND.n5272 GND.t172 126.766
R15623 GND.n5248 GND.t88 126.766
R15624 GND.n5266 GND.t120 126.766
R15625 GND.n5250 GND.t85 126.766
R15626 GND.n5260 GND.t53 126.766
R15627 GND.n773 GND.t35 126.766
R15628 GND.n775 GND.t154 126.766
R15629 GND.n779 GND.t62 126.766
R15630 GND.n781 GND.t169 126.766
R15631 GND.n792 GND.t111 126.766
R15632 GND.n794 GND.t160 126.766
R15633 GND.n6062 GND.t81 125.573
R15634 GND.n6956 GND.t128 125.573
R15635 GND.n2147 GND.t158 123.6
R15636 GND.n5925 GND.t84 123.6
R15637 GND.n1662 GND.t67 123.6
R15638 GND.n5965 GND.t41 123.6
R15639 GND.n5982 GND.t168 123.6
R15640 GND.n6000 GND.t144 123.6
R15641 GND.n720 GND.t69 123.6
R15642 GND.n731 GND.t60 123.6
R15643 GND.n7605 GND.t48 123.6
R15644 GND.n7617 GND.t149 123.6
R15645 GND.n7629 GND.t92 123.6
R15646 GND.n8345 GND.t45 123.6
R15647 GND.n8334 GND.t96 123.6
R15648 GND.n8324 GND.t58 123.6
R15649 GND.n8413 GND.t135 123.6
R15650 GND.n8303 GND.t153 123.6
R15651 GND.n355 GND.t102 123.6
R15652 GND.n668 GND.t131 123.6
R15653 GND.n4169 GND.t164 123.6
R15654 GND.n4180 GND.t146 123.6
R15655 GND.n4192 GND.t124 123.6
R15656 GND.n4204 GND.t109 123.6
R15657 GND.n4217 GND.t115 123.6
R15658 GND.n1639 GND.t52 123.6
R15659 GND.n8446 GND.n8445 99.6594
R15660 GND.n8441 GND.n8288 99.6594
R15661 GND.n8437 GND.n8287 99.6594
R15662 GND.n8305 GND.n8286 99.6594
R15663 GND.n8429 GND.n8285 99.6594
R15664 GND.n8425 GND.n8284 99.6594
R15665 GND.n8421 GND.n8283 99.6594
R15666 GND.n8417 GND.n8282 99.6594
R15667 GND.n8410 GND.n8281 99.6594
R15668 GND.n8406 GND.n8280 99.6594
R15669 GND.n8402 GND.n8279 99.6594
R15670 GND.n8398 GND.n8278 99.6594
R15671 GND.n8394 GND.n8277 99.6594
R15672 GND.n8386 GND.n8276 99.6594
R15673 GND.n8384 GND.n8275 99.6594
R15674 GND.n8380 GND.n8274 99.6594
R15675 GND.n8376 GND.n8273 99.6594
R15676 GND.n8372 GND.n8272 99.6594
R15677 GND.n8364 GND.n8271 99.6594
R15678 GND.n8362 GND.n8270 99.6594
R15679 GND.n8358 GND.n8269 99.6594
R15680 GND.n8354 GND.n8268 99.6594
R15681 GND.n8350 GND.n8267 99.6594
R15682 GND.n8342 GND.n8266 99.6594
R15683 GND.n7724 GND.n7723 99.6594
R15684 GND.n7718 GND.n672 99.6594
R15685 GND.n7715 GND.n673 99.6594
R15686 GND.n7711 GND.n674 99.6594
R15687 GND.n7707 GND.n675 99.6594
R15688 GND.n7704 GND.n676 99.6594
R15689 GND.n7700 GND.n677 99.6594
R15690 GND.n7696 GND.n678 99.6594
R15691 GND.n7692 GND.n679 99.6594
R15692 GND.n7687 GND.n680 99.6594
R15693 GND.n7683 GND.n681 99.6594
R15694 GND.n7680 GND.n682 99.6594
R15695 GND.n7677 GND.n683 99.6594
R15696 GND.n7673 GND.n684 99.6594
R15697 GND.n7669 GND.n685 99.6594
R15698 GND.n7665 GND.n686 99.6594
R15699 GND.n7661 GND.n687 99.6594
R15700 GND.n7657 GND.n688 99.6594
R15701 GND.n7653 GND.n689 99.6594
R15702 GND.n7649 GND.n690 99.6594
R15703 GND.n7645 GND.n691 99.6594
R15704 GND.n7641 GND.n692 99.6594
R15705 GND.n7637 GND.n693 99.6594
R15706 GND.n7633 GND.n694 99.6594
R15707 GND.n5908 GND.n1614 99.6594
R15708 GND.n5914 GND.n1615 99.6594
R15709 GND.n5918 GND.n1616 99.6594
R15710 GND.n5926 GND.n1617 99.6594
R15711 GND.n5930 GND.n1618 99.6594
R15712 GND.n5936 GND.n1619 99.6594
R15713 GND.n5940 GND.n1620 99.6594
R15714 GND.n5946 GND.n1621 99.6594
R15715 GND.n5949 GND.n1622 99.6594
R15716 GND.n5955 GND.n1623 99.6594
R15717 GND.n6041 GND.n1657 99.6594
R15718 GND.n5961 GND.n1656 99.6594
R15719 GND.n5963 GND.n1655 99.6594
R15720 GND.n5968 GND.n1654 99.6594
R15721 GND.n5972 GND.n1653 99.6594
R15722 GND.n5974 GND.n1652 99.6594
R15723 GND.n5978 GND.n1651 99.6594
R15724 GND.n5980 GND.n1650 99.6594
R15725 GND.n5986 GND.n1649 99.6594
R15726 GND.n5988 GND.n1648 99.6594
R15727 GND.n5992 GND.n1647 99.6594
R15728 GND.n5994 GND.n1646 99.6594
R15729 GND.n5998 GND.n1645 99.6594
R15730 GND.n1644 GND.n1606 99.6594
R15731 GND.n4312 GND.n2129 99.6594
R15732 GND.n4307 GND.n4129 99.6594
R15733 GND.n4304 GND.n4130 99.6594
R15734 GND.n4300 GND.n4131 99.6594
R15735 GND.n4296 GND.n4132 99.6594
R15736 GND.n4293 GND.n4133 99.6594
R15737 GND.n4289 GND.n4134 99.6594
R15738 GND.n4285 GND.n4135 99.6594
R15739 GND.n4281 GND.n4136 99.6594
R15740 GND.n4276 GND.n4137 99.6594
R15741 GND.n4272 GND.n4138 99.6594
R15742 GND.n4268 GND.n4139 99.6594
R15743 GND.n4264 GND.n4140 99.6594
R15744 GND.n4260 GND.n4141 99.6594
R15745 GND.n4256 GND.n4142 99.6594
R15746 GND.n4252 GND.n4143 99.6594
R15747 GND.n4248 GND.n4144 99.6594
R15748 GND.n4244 GND.n4145 99.6594
R15749 GND.n4240 GND.n4146 99.6594
R15750 GND.n4236 GND.n4147 99.6594
R15751 GND.n4232 GND.n4148 99.6594
R15752 GND.n4228 GND.n4149 99.6594
R15753 GND.n4224 GND.n4150 99.6594
R15754 GND.n4220 GND.n4151 99.6594
R15755 GND.n6921 GND.n6920 99.6594
R15756 GND.n6922 GND.n1075 99.6594
R15757 GND.n6932 GND.n6931 99.6594
R15758 GND.n6933 GND.n1073 99.6594
R15759 GND.n6942 GND.n6941 99.6594
R15760 GND.n6943 GND.n1071 99.6594
R15761 GND.n6952 GND.n6951 99.6594
R15762 GND.n6960 GND.n1069 99.6594
R15763 GND.n6964 GND.n6962 99.6594
R15764 GND.n6971 GND.n1066 99.6594
R15765 GND.n6099 GND.n6098 99.6594
R15766 GND.n6093 GND.n1576 99.6594
R15767 GND.n6090 GND.n1577 99.6594
R15768 GND.n6053 GND.n1578 99.6594
R15769 GND.n6055 GND.n1579 99.6594
R15770 GND.n6057 GND.n1580 99.6594
R15771 GND.n6059 GND.n1581 99.6594
R15772 GND.n6061 GND.n1582 99.6594
R15773 GND.n6070 GND.n1583 99.6594
R15774 GND.n370 GND.n358 99.6594
R15775 GND.n373 GND.n359 99.6594
R15776 GND.n380 GND.n379 99.6594
R15777 GND.n8449 GND.n8448 99.6594
R15778 GND.n696 GND.n695 99.6594
R15779 GND.n701 GND.n700 99.6594
R15780 GND.n705 GND.n704 99.6594
R15781 GND.n7727 GND.n7726 99.6594
R15782 GND.n697 GND.n696 99.6594
R15783 GND.n703 GND.n701 99.6594
R15784 GND.n705 GND.n670 99.6594
R15785 GND.n7726 GND.n666 99.6594
R15786 GND.n8448 GND.n357 99.6594
R15787 GND.n380 GND.n360 99.6594
R15788 GND.n371 GND.n359 99.6594
R15789 GND.n363 GND.n358 99.6594
R15790 GND.n6099 GND.n1587 99.6594
R15791 GND.n6091 GND.n1576 99.6594
R15792 GND.n1594 GND.n1577 99.6594
R15793 GND.n6054 GND.n1578 99.6594
R15794 GND.n6056 GND.n1579 99.6594
R15795 GND.n6058 GND.n1580 99.6594
R15796 GND.n6060 GND.n1581 99.6594
R15797 GND.n6064 GND.n1582 99.6594
R15798 GND.n6066 GND.n1583 99.6594
R15799 GND.n6963 GND.n1066 99.6594
R15800 GND.n6962 GND.n6961 99.6594
R15801 GND.n6953 GND.n1069 99.6594
R15802 GND.n6951 GND.n6950 99.6594
R15803 GND.n6944 GND.n6943 99.6594
R15804 GND.n6941 GND.n6940 99.6594
R15805 GND.n6934 GND.n6933 99.6594
R15806 GND.n6931 GND.n6930 99.6594
R15807 GND.n6923 GND.n6922 99.6594
R15808 GND.n6920 GND.n6919 99.6594
R15809 GND.n4312 GND.n4311 99.6594
R15810 GND.n4305 GND.n4129 99.6594
R15811 GND.n4301 GND.n4130 99.6594
R15812 GND.n4166 GND.n4131 99.6594
R15813 GND.n4294 GND.n4132 99.6594
R15814 GND.n4290 GND.n4133 99.6594
R15815 GND.n4286 GND.n4134 99.6594
R15816 GND.n4282 GND.n4135 99.6594
R15817 GND.n4277 GND.n4136 99.6594
R15818 GND.n4273 GND.n4137 99.6594
R15819 GND.n4269 GND.n4138 99.6594
R15820 GND.n4265 GND.n4139 99.6594
R15821 GND.n4261 GND.n4140 99.6594
R15822 GND.n4257 GND.n4141 99.6594
R15823 GND.n4253 GND.n4142 99.6594
R15824 GND.n4249 GND.n4143 99.6594
R15825 GND.n4245 GND.n4144 99.6594
R15826 GND.n4241 GND.n4145 99.6594
R15827 GND.n4237 GND.n4146 99.6594
R15828 GND.n4233 GND.n4147 99.6594
R15829 GND.n4229 GND.n4148 99.6594
R15830 GND.n4225 GND.n4149 99.6594
R15831 GND.n4221 GND.n4150 99.6594
R15832 GND.n4214 GND.n4151 99.6594
R15833 GND.n6001 GND.n1644 99.6594
R15834 GND.n5995 GND.n1645 99.6594
R15835 GND.n5993 GND.n1646 99.6594
R15836 GND.n5989 GND.n1647 99.6594
R15837 GND.n5987 GND.n1648 99.6594
R15838 GND.n5983 GND.n1649 99.6594
R15839 GND.n5979 GND.n1650 99.6594
R15840 GND.n5975 GND.n1651 99.6594
R15841 GND.n5973 GND.n1652 99.6594
R15842 GND.n5969 GND.n1653 99.6594
R15843 GND.n5967 GND.n1654 99.6594
R15844 GND.n5962 GND.n1655 99.6594
R15845 GND.n6040 GND.n1656 99.6594
R15846 GND.n5956 GND.n1624 99.6594
R15847 GND.n1664 GND.n1623 99.6594
R15848 GND.n5947 GND.n1622 99.6594
R15849 GND.n5939 GND.n1621 99.6594
R15850 GND.n5937 GND.n1620 99.6594
R15851 GND.n5929 GND.n1619 99.6594
R15852 GND.n5927 GND.n1618 99.6594
R15853 GND.n5917 GND.n1617 99.6594
R15854 GND.n5915 GND.n1616 99.6594
R15855 GND.n5907 GND.n1615 99.6594
R15856 GND.n5905 GND.n1614 99.6594
R15857 GND.n7724 GND.n708 99.6594
R15858 GND.n7716 GND.n672 99.6594
R15859 GND.n7712 GND.n673 99.6594
R15860 GND.n717 GND.n674 99.6594
R15861 GND.n7705 GND.n675 99.6594
R15862 GND.n7701 GND.n676 99.6594
R15863 GND.n7697 GND.n677 99.6594
R15864 GND.n7693 GND.n678 99.6594
R15865 GND.n7688 GND.n679 99.6594
R15866 GND.n7684 GND.n680 99.6594
R15867 GND.n7597 GND.n681 99.6594
R15868 GND.n7678 GND.n682 99.6594
R15869 GND.n7674 GND.n683 99.6594
R15870 GND.n7670 GND.n684 99.6594
R15871 GND.n7666 GND.n685 99.6594
R15872 GND.n7662 GND.n686 99.6594
R15873 GND.n7658 GND.n687 99.6594
R15874 GND.n7654 GND.n688 99.6594
R15875 GND.n7650 GND.n689 99.6594
R15876 GND.n7646 GND.n690 99.6594
R15877 GND.n7642 GND.n691 99.6594
R15878 GND.n7638 GND.n692 99.6594
R15879 GND.n7634 GND.n693 99.6594
R15880 GND.n694 GND.n657 99.6594
R15881 GND.n8349 GND.n8266 99.6594
R15882 GND.n8353 GND.n8267 99.6594
R15883 GND.n8357 GND.n8268 99.6594
R15884 GND.n8361 GND.n8269 99.6594
R15885 GND.n8365 GND.n8270 99.6594
R15886 GND.n8371 GND.n8271 99.6594
R15887 GND.n8375 GND.n8272 99.6594
R15888 GND.n8379 GND.n8273 99.6594
R15889 GND.n8383 GND.n8274 99.6594
R15890 GND.n8387 GND.n8275 99.6594
R15891 GND.n8393 GND.n8276 99.6594
R15892 GND.n8397 GND.n8277 99.6594
R15893 GND.n8401 GND.n8278 99.6594
R15894 GND.n8405 GND.n8279 99.6594
R15895 GND.n8409 GND.n8280 99.6594
R15896 GND.n8416 GND.n8281 99.6594
R15897 GND.n8420 GND.n8282 99.6594
R15898 GND.n8424 GND.n8283 99.6594
R15899 GND.n8428 GND.n8284 99.6594
R15900 GND.n8304 GND.n8285 99.6594
R15901 GND.n8436 GND.n8286 99.6594
R15902 GND.n8440 GND.n8287 99.6594
R15903 GND.n8290 GND.n8288 99.6594
R15904 GND.n8446 GND.n8289 99.6594
R15905 GND.n4152 GND.n2134 99.6594
R15906 GND.n4154 GND.n2140 99.6594
R15907 GND.n4155 GND.n2143 99.6594
R15908 GND.n4156 GND.n2145 99.6594
R15909 GND.n4152 GND.n2139 99.6594
R15910 GND.n4154 GND.n4153 99.6594
R15911 GND.n4155 GND.n2144 99.6594
R15912 GND.n4156 GND.n2151 99.6594
R15913 GND.n6044 GND.n6043 99.6594
R15914 GND.n1628 GND.n1627 99.6594
R15915 GND.n1633 GND.n1632 99.6594
R15916 GND.n1637 GND.n1636 99.6594
R15917 GND.n1641 GND.n1637 99.6594
R15918 GND.n1635 GND.n1633 99.6594
R15919 GND.n1629 GND.n1628 99.6594
R15920 GND.n6043 GND.n1612 99.6594
R15921 GND.n2147 GND.n2146 93.4793
R15922 GND.n5925 GND.n5924 93.4793
R15923 GND.n1662 GND.n1661 93.4793
R15924 GND.n5965 GND.n5964 93.4793
R15925 GND.n5982 GND.n5981 93.4793
R15926 GND.n6000 GND.n5999 93.4793
R15927 GND.n720 GND.n719 93.4793
R15928 GND.n731 GND.n730 93.4793
R15929 GND.n7605 GND.n7604 93.4793
R15930 GND.n7617 GND.n7616 93.4793
R15931 GND.n7629 GND.n7628 93.4793
R15932 GND.n8345 GND.n8344 93.4793
R15933 GND.n8334 GND.n8333 93.4793
R15934 GND.n8324 GND.n8323 93.4793
R15935 GND.n8413 GND.n8412 93.4793
R15936 GND.n8303 GND.n8302 93.4793
R15937 GND.n355 GND.n354 93.4793
R15938 GND.n668 GND.n667 93.4793
R15939 GND.n4169 GND.n4168 93.4793
R15940 GND.n4180 GND.n4179 93.4793
R15941 GND.n4192 GND.n4191 93.4793
R15942 GND.n4204 GND.n4203 93.4793
R15943 GND.n4217 GND.n4216 93.4793
R15944 GND.n1639 GND.n1638 93.4793
R15945 GND.n83 GND.n81 92.4005
R15946 GND.n94 GND.n92 92.4005
R15947 GND.n106 GND.n104 92.4005
R15948 GND.n118 GND.n116 92.4005
R15949 GND.n130 GND.n128 92.4005
R15950 GND.n142 GND.n140 92.4005
R15951 GND.n76 GND.t206 90.7789
R15952 GND.n19 GND.n18 90.3229
R15953 GND.n21 GND.n20 90.3229
R15954 GND.n30 GND.n29 90.3229
R15955 GND.n32 GND.n31 90.3229
R15956 GND.n42 GND.n41 90.3229
R15957 GND.n44 GND.n43 90.3229
R15958 GND.n54 GND.n53 90.3229
R15959 GND.n56 GND.n55 90.3229
R15960 GND.n66 GND.n65 90.3229
R15961 GND.n68 GND.n67 90.3229
R15962 GND.n8 GND.n7 90.3229
R15963 GND.n10 GND.n9 90.3229
R15964 GND.n83 GND.n82 90.3229
R15965 GND.n94 GND.n93 90.3229
R15966 GND.n106 GND.n105 90.3229
R15967 GND.n118 GND.n117 90.3229
R15968 GND.n130 GND.n129 90.3229
R15969 GND.n142 GND.n141 90.3229
R15970 GND.n79 GND.t210 89.7615
R15971 GND.n78 GND.t214 89.7615
R15972 GND.n77 GND.t208 89.7615
R15973 GND.n76 GND.t212 89.7615
R15974 GND.n5259 GND.n5258 83.3186
R15975 GND.n6063 GND.t80 76.7004
R15976 GND.n6957 GND.t129 76.7004
R15977 GND.n5260 GND.n5251 72.8411
R15978 GND.n5266 GND.n5249 72.8411
R15979 GND.n5272 GND.n5247 72.8411
R15980 GND.n792 GND.n791 72.8411
R15981 GND.n779 GND.n778 72.8411
R15982 GND.n7588 GND.n764 71.676
R15983 GND.n7584 GND.n763 71.676
R15984 GND.n7580 GND.n762 71.676
R15985 GND.n7576 GND.n761 71.676
R15986 GND.n7572 GND.n760 71.676
R15987 GND.n7568 GND.n759 71.676
R15988 GND.n7564 GND.n758 71.676
R15989 GND.n7560 GND.n757 71.676
R15990 GND.n7556 GND.n756 71.676
R15991 GND.n7552 GND.n755 71.676
R15992 GND.n7547 GND.n754 71.676
R15993 GND.n7543 GND.n753 71.676
R15994 GND.n7595 GND.n7594 71.676
R15995 GND.n7376 GND.n740 71.676
R15996 GND.n7380 GND.n741 71.676
R15997 GND.n7384 GND.n742 71.676
R15998 GND.n7388 GND.n743 71.676
R15999 GND.n7392 GND.n744 71.676
R16000 GND.n7396 GND.n745 71.676
R16001 GND.n7400 GND.n746 71.676
R16002 GND.n7404 GND.n747 71.676
R16003 GND.n7408 GND.n748 71.676
R16004 GND.n7412 GND.n749 71.676
R16005 GND.n7416 GND.n750 71.676
R16006 GND.n7420 GND.n751 71.676
R16007 GND.n7424 GND.n752 71.676
R16008 GND.n5279 GND.n5278 71.676
R16009 GND.n5283 GND.n5282 71.676
R16010 GND.n5288 GND.n5287 71.676
R16011 GND.n5291 GND.n5290 71.676
R16012 GND.n5296 GND.n5295 71.676
R16013 GND.n5299 GND.n5298 71.676
R16014 GND.n5304 GND.n5303 71.676
R16015 GND.n5307 GND.n5306 71.676
R16016 GND.n5312 GND.n5311 71.676
R16017 GND.n5315 GND.n5314 71.676
R16018 GND.n5323 GND.n5322 71.676
R16019 GND.n5326 GND.n5325 71.676
R16020 GND.n5331 GND.n5330 71.676
R16021 GND.n5336 GND.n5335 71.676
R16022 GND.n5344 GND.n5343 71.676
R16023 GND.n5347 GND.n5346 71.676
R16024 GND.n5352 GND.n5351 71.676
R16025 GND.n5355 GND.n5354 71.676
R16026 GND.n5360 GND.n5359 71.676
R16027 GND.n5363 GND.n5362 71.676
R16028 GND.n5368 GND.n5367 71.676
R16029 GND.n5371 GND.n5370 71.676
R16030 GND.n5376 GND.n5375 71.676
R16031 GND.n5379 GND.n5378 71.676
R16032 GND.n5384 GND.n5383 71.676
R16033 GND.n5280 GND.n5279 71.676
R16034 GND.n5282 GND.n5243 71.676
R16035 GND.n5289 GND.n5288 71.676
R16036 GND.n5290 GND.n5241 71.676
R16037 GND.n5297 GND.n5296 71.676
R16038 GND.n5298 GND.n5239 71.676
R16039 GND.n5305 GND.n5304 71.676
R16040 GND.n5306 GND.n5237 71.676
R16041 GND.n5313 GND.n5312 71.676
R16042 GND.n5314 GND.n5235 71.676
R16043 GND.n5324 GND.n5323 71.676
R16044 GND.n5325 GND.n5233 71.676
R16045 GND.n5334 GND.n5333 71.676
R16046 GND.n5335 GND.n5230 71.676
R16047 GND.n5345 GND.n5344 71.676
R16048 GND.n5346 GND.n5228 71.676
R16049 GND.n5353 GND.n5352 71.676
R16050 GND.n5354 GND.n5226 71.676
R16051 GND.n5361 GND.n5360 71.676
R16052 GND.n5362 GND.n5224 71.676
R16053 GND.n5369 GND.n5368 71.676
R16054 GND.n5370 GND.n5222 71.676
R16055 GND.n5377 GND.n5376 71.676
R16056 GND.n5378 GND.n5220 71.676
R16057 GND.n5385 GND.n5384 71.676
R16058 GND.n7421 GND.n752 71.676
R16059 GND.n7417 GND.n751 71.676
R16060 GND.n7413 GND.n750 71.676
R16061 GND.n7409 GND.n749 71.676
R16062 GND.n7405 GND.n748 71.676
R16063 GND.n7401 GND.n747 71.676
R16064 GND.n7397 GND.n746 71.676
R16065 GND.n7393 GND.n745 71.676
R16066 GND.n7389 GND.n744 71.676
R16067 GND.n7385 GND.n743 71.676
R16068 GND.n7381 GND.n742 71.676
R16069 GND.n7377 GND.n741 71.676
R16070 GND.n740 GND.n738 71.676
R16071 GND.n7542 GND.n737 71.676
R16072 GND.n7546 GND.n753 71.676
R16073 GND.n7551 GND.n754 71.676
R16074 GND.n7555 GND.n755 71.676
R16075 GND.n7559 GND.n756 71.676
R16076 GND.n7563 GND.n757 71.676
R16077 GND.n7567 GND.n758 71.676
R16078 GND.n7571 GND.n759 71.676
R16079 GND.n7575 GND.n760 71.676
R16080 GND.n7579 GND.n761 71.676
R16081 GND.n7583 GND.n762 71.676
R16082 GND.n7587 GND.n763 71.676
R16083 GND.n766 GND.n764 71.676
R16084 GND.n5340 GND.t105 71.314
R16085 GND.n7373 GND.t77 71.314
R16086 GND.n5319 GND.t137 71.3092
R16087 GND.n7541 GND.t99 71.3092
R16088 GND.n5320 GND.n5319 59.5399
R16089 GND.n5341 GND.n5340 59.5399
R16090 GND.n7374 GND.n7373 59.5399
R16091 GND.n7549 GND.n7541 59.5399
R16092 GND.n5276 GND.n5275 58.4046
R16093 GND.n5257 GND.n5256 54.358
R16094 GND.n789 GND.n788 54.358
R16095 GND.n772 GND.n771 52.3702
R16096 GND.n13 GND.t191 52.3082
R16097 GND.n24 GND.t237 52.3082
R16098 GND.n36 GND.t28 52.3082
R16099 GND.n48 GND.t226 52.3082
R16100 GND.n60 GND.t184 52.3082
R16101 GND.n2 GND.t224 52.3082
R16102 GND.n86 GND.t189 52.3082
R16103 GND.n97 GND.t230 52.3082
R16104 GND.n109 GND.t19 52.3082
R16105 GND.n121 GND.t227 52.3082
R16106 GND.n133 GND.t188 52.3082
R16107 GND.n145 GND.t236 52.3082
R16108 GND.n6063 GND.n6062 48.8732
R16109 GND.n6957 GND.n6956 48.8732
R16110 GND.n3938 GND.n3937 48.004
R16111 GND.n3938 GND.n2243 48.004
R16112 GND.n3946 GND.n2243 48.004
R16113 GND.n3947 GND.n3946 48.004
R16114 GND.n3948 GND.n3947 48.004
R16115 GND.n3948 GND.n2237 48.004
R16116 GND.n3956 GND.n2237 48.004
R16117 GND.n3957 GND.n3956 48.004
R16118 GND.n3958 GND.n3957 48.004
R16119 GND.n3958 GND.n2231 48.004
R16120 GND.n3966 GND.n2231 48.004
R16121 GND.n3967 GND.n3966 48.004
R16122 GND.n3968 GND.n3967 48.004
R16123 GND.n3968 GND.n2225 48.004
R16124 GND.n3976 GND.n2225 48.004
R16125 GND.n3977 GND.n3976 48.004
R16126 GND.n3978 GND.n3977 48.004
R16127 GND.n3978 GND.n2219 48.004
R16128 GND.n3986 GND.n2219 48.004
R16129 GND.n3987 GND.n3986 48.004
R16130 GND.n3988 GND.n3987 48.004
R16131 GND.n3988 GND.n2213 48.004
R16132 GND.n3996 GND.n2213 48.004
R16133 GND.n3997 GND.n3996 48.004
R16134 GND.n3998 GND.n3997 48.004
R16135 GND.n3998 GND.n2207 48.004
R16136 GND.n4006 GND.n2207 48.004
R16137 GND.n4007 GND.n4006 48.004
R16138 GND.n4008 GND.n4007 48.004
R16139 GND.n4008 GND.n2201 48.004
R16140 GND.n4016 GND.n2201 48.004
R16141 GND.n4017 GND.n4016 48.004
R16142 GND.n4018 GND.n4017 48.004
R16143 GND.n4018 GND.n2195 48.004
R16144 GND.n4026 GND.n2195 48.004
R16145 GND.n4027 GND.n4026 48.004
R16146 GND.n4028 GND.n4027 48.004
R16147 GND.n4028 GND.n2189 48.004
R16148 GND.n4036 GND.n2189 48.004
R16149 GND.n4037 GND.n4036 48.004
R16150 GND.n4038 GND.n4037 48.004
R16151 GND.n4038 GND.n2183 48.004
R16152 GND.n4046 GND.n2183 48.004
R16153 GND.n4047 GND.n4046 48.004
R16154 GND.n4048 GND.n4047 48.004
R16155 GND.n4048 GND.n2177 48.004
R16156 GND.n4056 GND.n2177 48.004
R16157 GND.n4057 GND.n4056 48.004
R16158 GND.n4058 GND.n4057 48.004
R16159 GND.n4058 GND.n2171 48.004
R16160 GND.n4066 GND.n2171 48.004
R16161 GND.n4067 GND.n4066 48.004
R16162 GND.n4068 GND.n4067 48.004
R16163 GND.n4068 GND.n2165 48.004
R16164 GND.n4076 GND.n2165 48.004
R16165 GND.n4077 GND.n4076 48.004
R16166 GND.n4078 GND.n4077 48.004
R16167 GND.n4078 GND.n2159 48.004
R16168 GND.n4086 GND.n2159 48.004
R16169 GND.n4087 GND.n4086 48.004
R16170 GND.n4088 GND.n4087 48.004
R16171 GND.n4088 GND.n2152 48.004
R16172 GND.n3936 GND.n2249 47.0291
R16173 GND.n3928 GND.n2249 47.0291
R16174 GND.n3928 GND.n3927 47.0291
R16175 GND.n3927 GND.n3926 47.0291
R16176 GND.n3926 GND.n2255 47.0291
R16177 GND.n3920 GND.n2255 47.0291
R16178 GND.n3920 GND.n3919 47.0291
R16179 GND.n3919 GND.n3918 47.0291
R16180 GND.n3918 GND.n2262 47.0291
R16181 GND.n3912 GND.n2262 47.0291
R16182 GND.n3912 GND.n3911 47.0291
R16183 GND.n3911 GND.n3910 47.0291
R16184 GND.n3910 GND.n2270 47.0291
R16185 GND.n3904 GND.n2270 47.0291
R16186 GND.n3904 GND.n3903 47.0291
R16187 GND.n3903 GND.n3902 47.0291
R16188 GND.n3902 GND.n2278 47.0291
R16189 GND.n3896 GND.n2278 47.0291
R16190 GND.n3896 GND.n3895 47.0291
R16191 GND.n3895 GND.n3894 47.0291
R16192 GND.n3894 GND.n2286 47.0291
R16193 GND.n3888 GND.n2286 47.0291
R16194 GND.n3888 GND.n3887 47.0291
R16195 GND.n3887 GND.n3886 47.0291
R16196 GND.n3886 GND.n2294 47.0291
R16197 GND.n3880 GND.n2294 47.0291
R16198 GND.n3880 GND.n3879 47.0291
R16199 GND.n3879 GND.n3878 47.0291
R16200 GND.n3878 GND.n2302 47.0291
R16201 GND.n3872 GND.n2302 47.0291
R16202 GND.n3872 GND.n3871 47.0291
R16203 GND.n3871 GND.n3870 47.0291
R16204 GND.n3870 GND.n2310 47.0291
R16205 GND.n3864 GND.n2310 47.0291
R16206 GND.n3864 GND.n3863 47.0291
R16207 GND.n3863 GND.n3862 47.0291
R16208 GND.n3862 GND.n2318 47.0291
R16209 GND.n3856 GND.n2318 47.0291
R16210 GND.n3856 GND.n3855 47.0291
R16211 GND.n3855 GND.n3854 47.0291
R16212 GND.n3854 GND.n2326 47.0291
R16213 GND.n3848 GND.n2326 47.0291
R16214 GND.n3848 GND.n3847 47.0291
R16215 GND.n3847 GND.n3846 47.0291
R16216 GND.n3846 GND.n2334 47.0291
R16217 GND.n3840 GND.n2334 47.0291
R16218 GND.n3840 GND.n3839 47.0291
R16219 GND.n3839 GND.n3838 47.0291
R16220 GND.n3838 GND.n2342 47.0291
R16221 GND.n3832 GND.n2342 47.0291
R16222 GND.n3832 GND.n3831 47.0291
R16223 GND.n3831 GND.n3830 47.0291
R16224 GND.n3830 GND.n2350 47.0291
R16225 GND.n3824 GND.n2350 47.0291
R16226 GND.n3824 GND.n3823 47.0291
R16227 GND.n3823 GND.n3822 47.0291
R16228 GND.n3822 GND.n2358 47.0291
R16229 GND.n3816 GND.n2358 47.0291
R16230 GND.n3816 GND.n3815 47.0291
R16231 GND.n3815 GND.n3814 47.0291
R16232 GND.n3814 GND.n2366 47.0291
R16233 GND.n3808 GND.n2366 47.0291
R16234 GND.n3808 GND.n3807 47.0291
R16235 GND.n3807 GND.n3806 47.0291
R16236 GND.n3806 GND.n2374 47.0291
R16237 GND.n3800 GND.n2374 47.0291
R16238 GND.n3800 GND.n3799 47.0291
R16239 GND.n3799 GND.n3798 47.0291
R16240 GND.n3798 GND.n2382 47.0291
R16241 GND.n3792 GND.n2382 47.0291
R16242 GND.n3792 GND.n3791 47.0291
R16243 GND.n3791 GND.n3790 47.0291
R16244 GND.n3790 GND.n2390 47.0291
R16245 GND.n3784 GND.n2390 47.0291
R16246 GND.n3784 GND.n3783 47.0291
R16247 GND.n3783 GND.n3782 47.0291
R16248 GND.n3782 GND.n2398 47.0291
R16249 GND.n3776 GND.n2398 47.0291
R16250 GND.n3776 GND.n3775 47.0291
R16251 GND.n3775 GND.n3774 47.0291
R16252 GND.n3774 GND.n2406 47.0291
R16253 GND.n3768 GND.n2406 47.0291
R16254 GND.n3768 GND.n3767 47.0291
R16255 GND.n3767 GND.n3766 47.0291
R16256 GND.n3766 GND.n2414 47.0291
R16257 GND.n3760 GND.n2414 47.0291
R16258 GND.n3760 GND.n3759 47.0291
R16259 GND.n3759 GND.n3758 47.0291
R16260 GND.n3758 GND.n2422 47.0291
R16261 GND.n3752 GND.n2422 47.0291
R16262 GND.n3752 GND.n3751 47.0291
R16263 GND.n3751 GND.n3750 47.0291
R16264 GND.n3750 GND.n2430 47.0291
R16265 GND.n3744 GND.n2430 47.0291
R16266 GND.n3744 GND.n3743 47.0291
R16267 GND.n3743 GND.n3742 47.0291
R16268 GND.n3742 GND.n2438 47.0291
R16269 GND.n3736 GND.n2438 47.0291
R16270 GND.n3736 GND.n3735 47.0291
R16271 GND.n3735 GND.n3734 47.0291
R16272 GND.n3734 GND.n2446 47.0291
R16273 GND.n3728 GND.n2446 47.0291
R16274 GND.n3728 GND.n3727 47.0291
R16275 GND.n3727 GND.n3726 47.0291
R16276 GND.n3726 GND.n2454 47.0291
R16277 GND.n3720 GND.n2454 47.0291
R16278 GND.n3720 GND.n3719 47.0291
R16279 GND.n3719 GND.n3718 47.0291
R16280 GND.n3718 GND.n2462 47.0291
R16281 GND.n3712 GND.n2462 47.0291
R16282 GND.n3712 GND.n3711 47.0291
R16283 GND.n3711 GND.n3710 47.0291
R16284 GND.n3710 GND.n2470 47.0291
R16285 GND.n3704 GND.n2470 47.0291
R16286 GND.n3704 GND.n3703 47.0291
R16287 GND.n3703 GND.n3702 47.0291
R16288 GND.n3702 GND.n2478 47.0291
R16289 GND.n3696 GND.n2478 47.0291
R16290 GND.n3696 GND.n3695 47.0291
R16291 GND.n3695 GND.n3694 47.0291
R16292 GND.n3694 GND.n2486 47.0291
R16293 GND.n3688 GND.n2486 47.0291
R16294 GND.n3688 GND.n3687 47.0291
R16295 GND.n3687 GND.n3686 47.0291
R16296 GND.n3686 GND.n2494 47.0291
R16297 GND.n3680 GND.n2494 47.0291
R16298 GND.n3680 GND.n3679 47.0291
R16299 GND.n3679 GND.n3678 47.0291
R16300 GND.n3678 GND.n2502 47.0291
R16301 GND.n3672 GND.n2502 47.0291
R16302 GND.n3672 GND.n3671 47.0291
R16303 GND.n3671 GND.n3670 47.0291
R16304 GND.n3670 GND.n2510 47.0291
R16305 GND.n3664 GND.n2510 47.0291
R16306 GND.n3664 GND.n3663 47.0291
R16307 GND.n3663 GND.n3662 47.0291
R16308 GND.n3662 GND.n2518 47.0291
R16309 GND.n3656 GND.n2518 47.0291
R16310 GND.n3656 GND.n3655 47.0291
R16311 GND.n3655 GND.n3654 47.0291
R16312 GND.n3654 GND.n2526 47.0291
R16313 GND.n3648 GND.n2526 47.0291
R16314 GND.n3648 GND.n3647 47.0291
R16315 GND.n3647 GND.n3646 47.0291
R16316 GND.n3646 GND.n2534 47.0291
R16317 GND.n3640 GND.n2534 47.0291
R16318 GND.n3640 GND.n3639 47.0291
R16319 GND.n3639 GND.n3638 47.0291
R16320 GND.n3638 GND.n2542 47.0291
R16321 GND.n3632 GND.n2542 47.0291
R16322 GND.n3632 GND.n3631 47.0291
R16323 GND.n3631 GND.n3630 47.0291
R16324 GND.n3630 GND.n2550 47.0291
R16325 GND.n3624 GND.n2550 47.0291
R16326 GND.n3624 GND.n3623 47.0291
R16327 GND.n3623 GND.n3622 47.0291
R16328 GND.n3622 GND.n2558 47.0291
R16329 GND.n3616 GND.n2558 47.0291
R16330 GND.n3616 GND.n3615 47.0291
R16331 GND.n3615 GND.n3614 47.0291
R16332 GND.n3614 GND.n2566 47.0291
R16333 GND.n3608 GND.n2566 47.0291
R16334 GND.n3608 GND.n3607 47.0291
R16335 GND.n3607 GND.n3606 47.0291
R16336 GND.n3606 GND.n2574 47.0291
R16337 GND.n3600 GND.n2574 47.0291
R16338 GND.n3600 GND.n3599 47.0291
R16339 GND.n3599 GND.n3598 47.0291
R16340 GND.n3598 GND.n2582 47.0291
R16341 GND.n3592 GND.n2582 47.0291
R16342 GND.n3592 GND.n3591 47.0291
R16343 GND.n3591 GND.n3590 47.0291
R16344 GND.n3590 GND.n2590 47.0291
R16345 GND.n3584 GND.n2590 47.0291
R16346 GND.n3584 GND.n3583 47.0291
R16347 GND.n3583 GND.n3582 47.0291
R16348 GND.n3582 GND.n2598 47.0291
R16349 GND.n3576 GND.n2598 47.0291
R16350 GND.n3576 GND.n3575 47.0291
R16351 GND.n3575 GND.n3574 47.0291
R16352 GND.n3574 GND.n2606 47.0291
R16353 GND.n3568 GND.n2606 47.0291
R16354 GND.n3568 GND.n3567 47.0291
R16355 GND.n3567 GND.n3566 47.0291
R16356 GND.n3566 GND.n2614 47.0291
R16357 GND.n3560 GND.n2614 47.0291
R16358 GND.n3560 GND.n3559 47.0291
R16359 GND.n3559 GND.n3558 47.0291
R16360 GND.n3558 GND.n2622 47.0291
R16361 GND.n3552 GND.n2622 47.0291
R16362 GND.n3552 GND.n3551 47.0291
R16363 GND.n3551 GND.n3550 47.0291
R16364 GND.n3550 GND.n2630 47.0291
R16365 GND.n3544 GND.n2630 47.0291
R16366 GND.n3544 GND.n3543 47.0291
R16367 GND.n3543 GND.n3542 47.0291
R16368 GND.n3542 GND.n2638 47.0291
R16369 GND.n3536 GND.n2638 47.0291
R16370 GND.n3536 GND.n3535 47.0291
R16371 GND.n3535 GND.n3534 47.0291
R16372 GND.n3534 GND.n2646 47.0291
R16373 GND.n3528 GND.n2646 47.0291
R16374 GND.n3528 GND.n3527 47.0291
R16375 GND.n3527 GND.n3526 47.0291
R16376 GND.n3526 GND.n2654 47.0291
R16377 GND.n3520 GND.n2654 47.0291
R16378 GND.n3520 GND.n3519 47.0291
R16379 GND.n3519 GND.n3518 47.0291
R16380 GND.n3518 GND.n2662 47.0291
R16381 GND.n3512 GND.n2662 47.0291
R16382 GND.n3512 GND.n3511 47.0291
R16383 GND.n3511 GND.n3510 47.0291
R16384 GND.n3510 GND.n2670 47.0291
R16385 GND.n3504 GND.n2670 47.0291
R16386 GND.n3504 GND.n3503 47.0291
R16387 GND.n3503 GND.n3502 47.0291
R16388 GND.n3502 GND.n2678 47.0291
R16389 GND.n3496 GND.n2678 47.0291
R16390 GND.n3496 GND.n3495 47.0291
R16391 GND.n3495 GND.n3494 47.0291
R16392 GND.n3494 GND.n2686 47.0291
R16393 GND.n3488 GND.n2686 47.0291
R16394 GND.n3488 GND.n3487 47.0291
R16395 GND.n3487 GND.n3486 47.0291
R16396 GND.n3486 GND.n2694 47.0291
R16397 GND.n3480 GND.n2694 47.0291
R16398 GND.n3480 GND.n3479 47.0291
R16399 GND.n3479 GND.n3478 47.0291
R16400 GND.n3478 GND.n2702 47.0291
R16401 GND.n3472 GND.n2702 47.0291
R16402 GND.n3472 GND.n3471 47.0291
R16403 GND.n3471 GND.n3470 47.0291
R16404 GND.n3470 GND.n2710 47.0291
R16405 GND.n3464 GND.n2710 47.0291
R16406 GND.n3464 GND.n3463 47.0291
R16407 GND.n3463 GND.n3462 47.0291
R16408 GND.n3462 GND.n2718 47.0291
R16409 GND.n3456 GND.n2718 47.0291
R16410 GND.n3456 GND.n3455 47.0291
R16411 GND.n3455 GND.n3454 47.0291
R16412 GND.n3454 GND.n2726 47.0291
R16413 GND.n3448 GND.n2726 47.0291
R16414 GND.n3448 GND.n3447 47.0291
R16415 GND.n3447 GND.n3446 47.0291
R16416 GND.n3446 GND.n2734 47.0291
R16417 GND.n3440 GND.n2734 47.0291
R16418 GND.n3440 GND.n3439 47.0291
R16419 GND.n3439 GND.n3438 47.0291
R16420 GND.n3438 GND.n2742 47.0291
R16421 GND.n3432 GND.n2742 47.0291
R16422 GND.n3432 GND.n3431 47.0291
R16423 GND.n3431 GND.n3430 47.0291
R16424 GND.n3430 GND.n2750 47.0291
R16425 GND.n3424 GND.n2750 47.0291
R16426 GND.n3424 GND.n3423 47.0291
R16427 GND.n3423 GND.n3422 47.0291
R16428 GND.n3422 GND.n2758 47.0291
R16429 GND.n3416 GND.n2758 47.0291
R16430 GND.n3416 GND.n3415 47.0291
R16431 GND.n3415 GND.n3414 47.0291
R16432 GND.n3414 GND.n2766 47.0291
R16433 GND.n3408 GND.n2766 47.0291
R16434 GND.n3408 GND.n3407 47.0291
R16435 GND.n3407 GND.n3406 47.0291
R16436 GND.n3406 GND.n2774 47.0291
R16437 GND.n3400 GND.n2774 47.0291
R16438 GND.n3400 GND.n3399 47.0291
R16439 GND.n3399 GND.n3398 47.0291
R16440 GND.n3398 GND.n2782 47.0291
R16441 GND.n3392 GND.n2782 47.0291
R16442 GND.n3392 GND.n3391 47.0291
R16443 GND.n3391 GND.n3390 47.0291
R16444 GND.n3390 GND.n2790 47.0291
R16445 GND.n3384 GND.n2790 47.0291
R16446 GND.n3384 GND.n3383 47.0291
R16447 GND.n3383 GND.n3382 47.0291
R16448 GND.n3382 GND.n2798 47.0291
R16449 GND.n3376 GND.n2798 47.0291
R16450 GND.n3376 GND.n3375 47.0291
R16451 GND.n3375 GND.n3374 47.0291
R16452 GND.n3374 GND.n2806 47.0291
R16453 GND.n3368 GND.n2806 47.0291
R16454 GND.n3368 GND.n3367 47.0291
R16455 GND.n3367 GND.n3366 47.0291
R16456 GND.n3366 GND.n2814 47.0291
R16457 GND.n3360 GND.n2814 47.0291
R16458 GND.n3360 GND.n3359 47.0291
R16459 GND.n3359 GND.n3358 47.0291
R16460 GND.n3358 GND.n2822 47.0291
R16461 GND.n3352 GND.n2822 47.0291
R16462 GND.n3352 GND.n3351 47.0291
R16463 GND.n3351 GND.n3350 47.0291
R16464 GND.n3350 GND.n2830 47.0291
R16465 GND.n3344 GND.n2830 47.0291
R16466 GND.n3344 GND.n3343 47.0291
R16467 GND.n3343 GND.n3342 47.0291
R16468 GND.n3342 GND.n2838 47.0291
R16469 GND.n3336 GND.n2838 47.0291
R16470 GND.n3336 GND.n3335 47.0291
R16471 GND.n3335 GND.n3334 47.0291
R16472 GND.n3334 GND.n2846 47.0291
R16473 GND.n3328 GND.n2846 47.0291
R16474 GND.n3328 GND.n3327 47.0291
R16475 GND.n3327 GND.n3326 47.0291
R16476 GND.n3326 GND.n2854 47.0291
R16477 GND.n3320 GND.n2854 47.0291
R16478 GND.n3320 GND.n3319 47.0291
R16479 GND.n3319 GND.n3318 47.0291
R16480 GND.n3318 GND.n2862 47.0291
R16481 GND.n3312 GND.n2862 47.0291
R16482 GND.n3312 GND.n3311 47.0291
R16483 GND.n3311 GND.n3310 47.0291
R16484 GND.n3310 GND.n2870 47.0291
R16485 GND.n3304 GND.n2870 47.0291
R16486 GND.n3304 GND.n3303 47.0291
R16487 GND.n3303 GND.n3302 47.0291
R16488 GND.n3302 GND.n2878 47.0291
R16489 GND.n3296 GND.n2878 47.0291
R16490 GND.n3296 GND.n3295 47.0291
R16491 GND.n3295 GND.n3294 47.0291
R16492 GND.n3294 GND.n2886 47.0291
R16493 GND.n3288 GND.n2886 47.0291
R16494 GND.n3288 GND.n3287 47.0291
R16495 GND.n3287 GND.n3286 47.0291
R16496 GND.n3286 GND.n2894 47.0291
R16497 GND.n3280 GND.n2894 47.0291
R16498 GND.n3280 GND.n3279 47.0291
R16499 GND.n3279 GND.n3278 47.0291
R16500 GND.n3278 GND.n2902 47.0291
R16501 GND.n3272 GND.n2902 47.0291
R16502 GND.n3272 GND.n3271 47.0291
R16503 GND.n3271 GND.n3270 47.0291
R16504 GND.n3270 GND.n2910 47.0291
R16505 GND.n3264 GND.n2910 47.0291
R16506 GND.n3264 GND.n3263 47.0291
R16507 GND.n3263 GND.n3262 47.0291
R16508 GND.n3262 GND.n2918 47.0291
R16509 GND.n3256 GND.n2918 47.0291
R16510 GND.n3256 GND.n3255 47.0291
R16511 GND.n3255 GND.n3254 47.0291
R16512 GND.n3254 GND.n2926 47.0291
R16513 GND.n3248 GND.n2926 47.0291
R16514 GND.n3248 GND.n3247 47.0291
R16515 GND.n3247 GND.n3246 47.0291
R16516 GND.n3246 GND.n2934 47.0291
R16517 GND.n3240 GND.n2934 47.0291
R16518 GND.n3240 GND.n3239 47.0291
R16519 GND.n3239 GND.n3238 47.0291
R16520 GND.n3238 GND.n2942 47.0291
R16521 GND.n3232 GND.n2942 47.0291
R16522 GND.n3232 GND.n3231 47.0291
R16523 GND.n3231 GND.n3230 47.0291
R16524 GND.n3230 GND.n2950 47.0291
R16525 GND.n3224 GND.n2950 47.0291
R16526 GND.n3224 GND.n3223 47.0291
R16527 GND.n3223 GND.n3222 47.0291
R16528 GND.n3222 GND.n2958 47.0291
R16529 GND.n3216 GND.n2958 47.0291
R16530 GND.n3216 GND.n3215 47.0291
R16531 GND.n5260 GND.n5259 45.8904
R16532 GND.n7539 GND.n795 44.3322
R16533 GND.n5273 GND.n5272 43.8187
R16534 GND.n793 GND.n792 43.8187
R16535 GND.n2148 GND.n2147 42.4732
R16536 GND.n5928 GND.n5925 42.4732
R16537 GND.n1663 GND.n1662 42.4732
R16538 GND.n6033 GND.n5965 42.4732
R16539 GND.n5984 GND.n5982 42.4732
R16540 GND.n6003 GND.n6000 42.4732
R16541 GND.n7709 GND.n720 42.4732
R16542 GND.n7690 GND.n731 42.4732
R16543 GND.n7672 GND.n7605 42.4732
R16544 GND.n7652 GND.n7617 42.4732
R16545 GND.n7632 GND.n7629 42.4732
R16546 GND.n8348 GND.n8345 42.4732
R16547 GND.n8370 GND.n8334 42.4732
R16548 GND.n8392 GND.n8324 42.4732
R16549 GND.n8414 GND.n8413 42.4732
R16550 GND.n8434 GND.n8303 42.4732
R16551 GND.n356 GND.n355 42.4732
R16552 GND.n6073 GND.n6063 42.4732
R16553 GND.n6958 GND.n6957 42.4732
R16554 GND.n7729 GND.n668 42.4732
R16555 GND.n4298 GND.n4169 42.4732
R16556 GND.n4279 GND.n4180 42.4732
R16557 GND.n4259 GND.n4192 42.4732
R16558 GND.n4239 GND.n4204 42.4732
R16559 GND.n4219 GND.n4217 42.4732
R16560 GND.n1640 GND.n1639 42.4732
R16561 GND.n5258 GND.n5257 41.6274
R16562 GND.n790 GND.n789 41.6274
R16563 GND.n19 GND.n17 39.6932
R16564 GND.n30 GND.n28 39.6932
R16565 GND.n42 GND.n40 39.6932
R16566 GND.n54 GND.n52 39.6932
R16567 GND.n66 GND.n64 39.6932
R16568 GND.n8 GND.n6 39.6932
R16569 GND.n5267 GND.n5266 37.9763
R16570 GND.n5266 GND.n5265 37.9763
R16571 GND.n779 GND.n770 37.9763
R16572 GND.n780 GND.n779 37.9763
R16573 GND.n91 GND.n90 37.6157
R16574 GND.n102 GND.n101 37.6157
R16575 GND.n114 GND.n113 37.6157
R16576 GND.n126 GND.n125 37.6157
R16577 GND.n138 GND.n137 37.6157
R16578 GND.n150 GND.n149 37.6157
R16579 GND.n4313 GND.n4128 36.8055
R16580 GND.n8447 GND.n8265 36.8055
R16581 GND.n1613 GND.n1610 36.0838
R16582 GND.n4952 GND.n1643 36.0838
R16583 GND.n5842 GND.n4952 36.0838
R16584 GND.n5842 GND.n5841 36.0838
R16585 GND.n5841 GND.n5840 36.0838
R16586 GND.n7528 GND.n7527 36.0838
R16587 GND.n7527 GND.n7526 36.0838
R16588 GND.n7526 GND.n7452 36.0838
R16589 GND.n7452 GND.n671 36.0838
R16590 GND.n706 GND.n658 36.0838
R16591 GND.n7427 GND.n7423 33.8737
R16592 GND.n5388 GND.n5218 33.8737
R16593 GND.n5272 GND.n5271 32.1338
R16594 GND.n5261 GND.n5260 32.1338
R16595 GND.n774 GND.n773 32.1338
R16596 GND.n792 GND.n768 32.1338
R16597 GND.n5232 GND.n1658 30.7205
R16598 GND.n7682 GND.n7596 30.7205
R16599 GND.n4345 GND.n2130 29.5888
R16600 GND.n4331 GND.n2133 29.5888
R16601 GND.n4355 GND.n2121 29.5888
R16602 GND.n4334 GND.n2123 29.5888
R16603 GND.n4364 GND.n2114 29.5888
R16604 GND.n4381 GND.n2102 29.5888
R16605 GND.n4391 GND.n2092 29.5888
R16606 GND.n4370 GND.n2094 29.5888
R16607 GND.n4412 GND.n2085 29.5888
R16608 GND.n4424 GND.n2073 29.5888
R16609 GND.n2076 GND.n2063 29.5888
R16610 GND.n4433 GND.n4432 29.5888
R16611 GND.n4399 GND.n2066 29.5888
R16612 GND.n4463 GND.n2039 29.5888
R16613 GND.n2050 GND.n2042 29.5888
R16614 GND.n4473 GND.n2029 29.5888
R16615 GND.n4452 GND.n2031 29.5888
R16616 GND.n4506 GND.n2011 29.5888
R16617 GND.n2014 GND.n2001 29.5888
R16618 GND.n4515 GND.n4514 29.5888
R16619 GND.n4481 GND.n2004 29.5888
R16620 GND.n4581 GND.n1977 29.5888
R16621 GND.n1988 GND.n1980 29.5888
R16622 GND.n4591 GND.n1967 29.5888
R16623 GND.n4570 GND.n1969 29.5888
R16624 GND.n4613 GND.n1947 29.5888
R16625 GND.n4597 GND.n1950 29.5888
R16626 GND.n4621 GND.n1940 29.5888
R16627 GND.n4624 GND.n1937 29.5888
R16628 GND.n4685 GND.n1882 29.5888
R16629 GND.n1931 GND.n1885 29.5888
R16630 GND.n4633 GND.n1930 29.5888
R16631 GND.n4636 GND.n1928 29.5888
R16632 GND.n4641 GND.n1920 29.5888
R16633 GND.n4652 GND.n1914 29.5888
R16634 GND.n4657 GND.n1911 29.5888
R16635 GND.n4660 GND.n1909 29.5888
R16636 GND.n4694 GND.n1864 29.5888
R16637 GND.n1866 GND.n1857 29.5888
R16638 GND.n4705 GND.n4704 29.5888
R16639 GND.n4740 GND.n1836 29.5888
R16640 GND.n1847 GND.n1839 29.5888
R16641 GND.n4750 GND.n1827 29.5888
R16642 GND.n4729 GND.n4728 29.5888
R16643 GND.n4760 GND.n1821 29.5888
R16644 GND.n4778 GND.n1809 29.5888
R16645 GND.n4763 GND.n1812 29.5888
R16646 GND.n4788 GND.n1799 29.5888
R16647 GND.n1801 GND.n1792 29.5888
R16648 GND.n4799 GND.n4798 29.5888
R16649 GND.n4846 GND.n1775 29.5888
R16650 GND.n4832 GND.n1778 29.5888
R16651 GND.n4835 GND.n1767 29.5888
R16652 GND.n4866 GND.n1760 29.5888
R16653 GND.n4883 GND.n1748 29.5888
R16654 GND.n4869 GND.n1751 29.5888
R16655 GND.n4893 GND.n1738 29.5888
R16656 GND.n4872 GND.n1740 29.5888
R16657 GND.n4912 GND.n1732 29.5888
R16658 GND.n4921 GND.n1718 29.5888
R16659 GND.n1721 GND.n1710 29.5888
R16660 GND.n4930 GND.n4929 29.5888
R16661 GND.n5861 GND.n1702 29.5888
R16662 GND.n5864 GND.n1693 29.5888
R16663 GND.n5890 GND.n1682 29.5888
R16664 GND.n5869 GND.n1684 29.5888
R16665 GND.n5899 GND.n1676 29.5888
R16666 GND.n6046 GND.n1607 29.5888
R16667 GND.n7737 GND.n647 29.5888
R16668 GND.n7754 GND.n650 29.5888
R16669 GND.n7747 GND.n637 29.5888
R16670 GND.n7764 GND.n639 29.5888
R16671 GND.n7741 GND.n631 29.5888
R16672 GND.n7791 GND.n622 29.5888
R16673 GND.n7778 GND.n609 29.5888
R16674 GND.n7801 GND.n611 29.5888
R16675 GND.n7784 GND.n603 29.5888
R16676 GND.n7815 GND.n592 29.5888
R16677 GND.n7826 GND.n595 29.5888
R16678 GND.n7809 GND.n585 29.5888
R16679 GND.n7834 GND.n582 29.5888
R16680 GND.n7837 GND.n570 29.5888
R16681 GND.n7853 GND.n573 29.5888
R16682 GND.n7846 GND.n564 29.5888
R16683 GND.n7869 GND.n536 29.5888
R16684 GND.n7891 GND.n539 29.5888
R16685 GND.n7900 GND.n526 29.5888
R16686 GND.n7899 GND.n529 29.5888
R16687 GND.n7882 GND.n505 29.5888
R16688 GND.n7944 GND.n508 29.5888
R16689 GND.n549 GND.n495 29.5888
R16690 GND.n7954 GND.n497 29.5888
R16691 GND.n7937 GND.n7936 29.5888
R16692 GND.n7964 GND.n478 29.5888
R16693 GND.n7981 GND.n481 29.5888
R16694 GND.n7968 GND.n468 29.5888
R16695 GND.n7991 GND.n470 29.5888
R16696 GND.n7974 GND.n462 29.5888
R16697 GND.n8006 GND.n455 29.5888
R16698 GND.n8015 GND.n449 29.5888
R16699 GND.n8020 GND.n451 29.5888
R16700 GND.n8033 GND.n441 29.5888
R16701 GND.n8566 GND.n160 29.5888
R16702 GND.n8122 GND.n435 29.5888
R16703 GND.n8125 GND.n429 29.5888
R16704 GND.n8132 GND.n177 29.5888
R16705 GND.n8559 GND.n180 29.5888
R16706 GND.n8140 GND.n189 29.5888
R16707 GND.n8553 GND.n192 29.5888
R16708 GND.n8147 GND.n199 29.5888
R16709 GND.n8547 GND.n202 29.5888
R16710 GND.n8541 GND.n212 29.5888
R16711 GND.n8162 GND.n220 29.5888
R16712 GND.n8535 GND.n223 29.5888
R16713 GND.n8170 GND.n230 29.5888
R16714 GND.n8529 GND.n233 29.5888
R16715 GND.n8177 GND.n241 29.5888
R16716 GND.n8523 GND.n244 29.5888
R16717 GND.n8185 GND.n251 29.5888
R16718 GND.n8192 GND.n261 29.5888
R16719 GND.n8511 GND.n264 29.5888
R16720 GND.n8200 GND.n271 29.5888
R16721 GND.n8505 GND.n274 29.5888
R16722 GND.n8207 GND.n282 29.5888
R16723 GND.n8499 GND.n285 29.5888
R16724 GND.n8215 GND.n292 29.5888
R16725 GND.n8493 GND.n295 29.5888
R16726 GND.n8222 GND.n303 29.5888
R16727 GND.n8487 GND.n306 29.5888
R16728 GND.n8231 GND.n313 29.5888
R16729 GND.n8246 GND.n323 29.5888
R16730 GND.n8475 GND.n326 29.5888
R16731 GND.n8240 GND.n333 29.5888
R16732 GND.n8469 GND.n336 29.5888
R16733 GND.n8456 GND.n343 29.5888
R16734 GND.n8463 GND.n346 29.5888
R16735 GND.n4313 GND.n2130 28.5063
R16736 GND.n8447 GND.n346 28.5063
R16737 GND.n4494 GND.t16 28.1455
R16738 GND.n8517 GND.t18 28.1455
R16739 GND.n4961 GND.n4953 27.7847
R16740 GND.n7593 GND.n739 27.7847
R16741 GND.n4569 GND.t6 24.5372
R16742 GND.n5813 GND.n4987 24.5372
R16743 GND.n5426 GND.n5014 24.5372
R16744 GND.n5785 GND.n5022 24.5372
R16745 GND.n5439 GND.n5032 24.5372
R16746 GND.n5771 GND.n5040 24.5372
R16747 GND.n5452 GND.n5050 24.5372
R16748 GND.n5757 GND.n5756 24.5372
R16749 GND.n5469 GND.n5072 24.5372
R16750 GND.n5742 GND.n5080 24.5372
R16751 GND.n5483 GND.n5089 24.5372
R16752 GND.n5728 GND.n5097 24.5372
R16753 GND.n5496 GND.n5107 24.5372
R16754 GND.n5714 GND.n5115 24.5372
R16755 GND.n5509 GND.n5125 24.5372
R16756 GND.n5700 GND.n5699 24.5372
R16757 GND.n5526 GND.n5147 24.5372
R16758 GND.n5685 GND.n5155 24.5372
R16759 GND.n5539 GND.n5165 24.5372
R16760 GND.n5671 GND.n5173 24.5372
R16761 GND.n5552 GND.n5183 24.5372
R16762 GND.n5657 GND.n5191 24.5372
R16763 GND.n5649 GND.n1575 24.5372
R16764 GND.n5201 GND.n1569 24.5372
R16765 GND.n5631 GND.n1562 24.5372
R16766 GND.n5624 GND.n1555 24.5372
R16767 GND.n5583 GND.n1546 24.5372
R16768 GND.n6157 GND.n1530 24.5372
R16769 GND.n6321 GND.n1505 24.5372
R16770 GND.n6313 GND.n1495 24.5372
R16771 GND.n6305 GND.n1487 24.5372
R16772 GND.n6291 GND.n1461 24.5372
R16773 GND.n6284 GND.n1453 24.5372
R16774 GND.n6277 GND.n1445 24.5372
R16775 GND.n6270 GND.n1437 24.5372
R16776 GND.n6263 GND.n1428 24.5372
R16777 GND.n6256 GND.n1422 24.5372
R16778 GND.n6560 GND.n1323 24.5372
R16779 GND.n6548 GND.n1304 24.5372
R16780 GND.n6541 GND.n1296 24.5372
R16781 GND.n6534 GND.n1288 24.5372
R16782 GND.n6527 GND.n1280 24.5372
R16783 GND.n6520 GND.n1272 24.5372
R16784 GND.n6513 GND.n1264 24.5372
R16785 GND.n6506 GND.n1256 24.5372
R16786 GND.n6499 GND.n1248 24.5372
R16787 GND.n6475 GND.n1242 24.5372
R16788 GND.n6485 GND.n1234 24.5372
R16789 GND.n1391 GND.n1225 24.5372
R16790 GND.n6679 GND.n1209 24.5372
R16791 GND.n6818 GND.n1170 24.5372
R16792 GND.n6810 GND.n1160 24.5372
R16793 GND.n6802 GND.n1152 24.5372
R16794 GND.n6788 GND.n1126 24.5372
R16795 GND.n6781 GND.n1118 24.5372
R16796 GND.n6774 GND.n1110 24.5372
R16797 GND.n6767 GND.n1101 24.5372
R16798 GND.n6895 GND.n1093 24.5372
R16799 GND.n6904 GND.n1055 24.5372
R16800 GND.n6993 GND.n1045 24.5372
R16801 GND.n7000 GND.n6999 24.5372
R16802 GND.n7018 GND.n1033 24.5372
R16803 GND.n7045 GND.n1017 24.5372
R16804 GND.n7052 GND.n7051 24.5372
R16805 GND.n7070 GND.n1003 24.5372
R16806 GND.n7076 GND.n999 24.5372
R16807 GND.n7094 GND.n983 24.5372
R16808 GND.n7105 GND.n972 24.5372
R16809 GND.n7126 GND.n963 24.5372
R16810 GND.n7144 GND.n953 24.5372
R16811 GND.n7150 GND.n949 24.5372
R16812 GND.n7177 GND.n933 24.5372
R16813 GND.n7185 GND.n7184 24.5372
R16814 GND.n7204 GND.n920 24.5372
R16815 GND.n7210 GND.n916 24.5372
R16816 GND.n7246 GND.n901 24.5372
R16817 GND.n7253 GND.n7252 24.5372
R16818 GND.n7266 GND.n7265 24.5372
R16819 GND.n7284 GND.n877 24.5372
R16820 GND.n7290 GND.n873 24.5372
R16821 GND.n7308 GND.n857 24.5372
R16822 GND.n7320 GND.n846 24.5372
R16823 GND.n7343 GND.n830 24.5372
R16824 GND.n7362 GND.n7361 24.5372
R16825 GND.n7435 GND.n806 24.5372
R16826 GND.n7535 GND.n798 24.5372
R16827 GND.t4 GND.n209 24.5372
R16828 GND.n5396 GND.n4979 23.8155
R16829 GND.n5819 GND.n4981 23.8155
R16830 GND.n5764 GND.n5763 23.8155
R16831 GND.n5457 GND.n5058 23.8155
R16832 GND.n5707 GND.n5706 23.8155
R16833 GND.n5514 GND.n5133 23.8155
R16834 GND.n6109 GND.n1567 23.8155
R16835 GND.n6306 GND.n1477 23.8155
R16836 GND.t205 GND.n1479 23.8155
R16837 GND.n6554 GND.n1329 23.8155
R16838 GND.n1335 GND.n1313 23.8155
R16839 GND.n6631 GND.n1250 23.8155
R16840 GND.n6639 GND.n1240 23.8155
R16841 GND.t203 GND.n1134 23.8155
R16842 GND.n6789 GND.n1136 23.8155
R16843 GND.n7012 GND.n1037 23.8155
R16844 GND.n7125 GND.n965 23.8155
R16845 GND.n7132 GND.n959 23.8155
R16846 GND.n7259 GND.n891 23.8155
R16847 GND.n892 GND.n887 23.8155
R16848 GND.n5833 GND.t173 22.3722
R16849 GND.n5827 GND.n4969 22.3722
R16850 GND.n5409 GND.n4989 22.3722
R16851 GND.n5770 GND.n5042 22.3722
R16852 GND.n5464 GND.n5061 22.3722
R16853 GND.n5713 GND.n5117 22.3722
R16854 GND.n5521 GND.n5136 22.3722
R16855 GND.n5656 GND.n5651 22.3722
R16856 GND.n6312 GND.n1485 22.3722
R16857 GND.n6178 GND.n1471 22.3722
R16858 GND.n6404 GND.n1319 22.3722
R16859 GND.n1339 GND.n1306 22.3722
R16860 GND.n6623 GND.n1258 22.3722
R16861 GND.n6647 GND.n1232 22.3722
R16862 GND.n6803 GND.n1142 22.3722
R16863 GND.n1203 GND.n1128 22.3722
R16864 GND.n7039 GND.n7038 22.3722
R16865 GND.n7112 GND.n7111 22.3722
R16866 GND.n7151 GND.n947 22.3722
R16867 GND.n903 GND.n902 22.3722
R16868 GND.n7272 GND.n883 22.3722
R16869 GND.n7350 GND.t36 22.3722
R16870 GND.n4367 GND.t108 21.6505
R16871 GND.n4831 GND.t27 21.6505
R16872 GND.n817 GND.t63 21.6505
R16873 GND.t2 GND.n558 21.6505
R16874 GND.n8481 GND.t43 21.6505
R16875 GND.n6100 GND.n1585 21.2897
R16876 GND.n7010 GND.n1031 21.2897
R16877 GND.n5276 GND.n4966 21.0737
R16878 GND.n7539 GND.n7538 21.0737
R16879 GND.n5805 GND.n4999 20.9288
R16880 GND.n5778 GND.n5777 20.9288
R16881 GND.n5748 GND.n5074 20.9288
R16882 GND.n5721 GND.n5720 20.9288
R16883 GND.n5664 GND.n5663 20.9288
R16884 GND.n6125 GND.n1553 20.9288
R16885 GND.n5611 GND.n1493 20.9288
R16886 GND.n6185 GND.n1463 20.9288
R16887 GND.n6394 GND.n1430 20.9288
R16888 GND.t201 GND.n1298 20.9288
R16889 GND.t207 GND.n1266 20.9288
R16890 GND.n6664 GND.n1223 20.9288
R16891 GND.n6809 GND.n1150 20.9288
R16892 GND.n6710 GND.n1120 20.9288
R16893 GND.n6979 GND.n1057 20.9288
R16894 GND.n1018 GND.n1013 20.9288
R16895 GND.n7171 GND.n7170 20.9288
R16896 GND.n7240 GND.n907 20.9288
R16897 GND.n7291 GND.n871 20.9288
R16898 GND.n7335 GND.n840 20.9288
R16899 GND.n7425 GND.n739 20.9288
R16900 GND.n6042 GND.n1643 20.568
R16901 GND.n7725 GND.n671 20.568
R16902 GND.n5154 GND.t235 20.2072
R16903 GND.n985 GND.t23 20.2072
R16904 GND.n5255 GND.t122 19.8005
R16905 GND.n5255 GND.t87 19.8005
R16906 GND.n5253 GND.t174 19.8005
R16907 GND.n5253 GND.t90 19.8005
R16908 GND.n5252 GND.t55 19.8005
R16909 GND.n5252 GND.t73 19.8005
R16910 GND.n784 GND.t113 19.8005
R16911 GND.n784 GND.t162 19.8005
R16912 GND.n787 GND.t64 19.8005
R16913 GND.n787 GND.t171 19.8005
R16914 GND.n785 GND.t37 19.8005
R16915 GND.n785 GND.t156 19.8005
R16916 GND.n5247 GND.n5246 19.5087
R16917 GND.n5270 GND.n5247 19.5087
R16918 GND.n5268 GND.n5249 19.5087
R16919 GND.n5264 GND.n5249 19.5087
R16920 GND.n5262 GND.n5251 19.5087
R16921 GND.n778 GND.n777 19.5087
R16922 GND.n778 GND.n769 19.5087
R16923 GND.n791 GND.n783 19.5087
R16924 GND.n5423 GND.n5006 19.4855
R16925 GND.n5784 GND.n5024 19.4855
R16926 GND.n5480 GND.n5479 19.4855
R16927 GND.n5727 GND.n5099 19.4855
R16928 GND.n5536 GND.n5157 19.4855
R16929 GND.n5670 GND.n5175 19.4855
R16930 GND.n6142 GND.n1544 19.4855
R16931 GND.n1531 GND.n1501 19.4855
R16932 GND.n6192 GND.n1455 19.4855
R16933 GND.n6384 GND.n1439 19.4855
R16934 GND.n1351 GND.n1290 19.4855
R16935 GND.n6608 GND.n1274 19.4855
R16936 GND.n6673 GND.n6672 19.4855
R16937 GND.n6460 GND.n1158 19.4855
R16938 GND.n6741 GND.n1112 19.4855
R16939 GND.n6894 GND.n1087 19.4855
R16940 GND.n7058 GND.n1009 19.4855
R16941 GND.n7088 GND.n989 19.4855
R16942 GND.n934 GND.n929 19.4855
R16943 GND.n7203 GND.n7202 19.4855
R16944 GND.n7302 GND.n7301 19.4855
R16945 GND.n7327 GND.n7326 19.4855
R16946 GND.n2149 GND.n2119 19.3944
R16947 GND.n4357 GND.n2119 19.3944
R16948 GND.n4357 GND.n2116 19.3944
R16949 GND.n4362 GND.n2116 19.3944
R16950 GND.n4362 GND.n2117 19.3944
R16951 GND.n2117 GND.n2090 19.3944
R16952 GND.n4393 GND.n2090 19.3944
R16953 GND.n4393 GND.n2087 19.3944
R16954 GND.n4410 GND.n2087 19.3944
R16955 GND.n4410 GND.n2088 19.3944
R16956 GND.n4406 GND.n2088 19.3944
R16957 GND.n4406 GND.n4405 19.3944
R16958 GND.n4405 GND.n4404 19.3944
R16959 GND.n4404 GND.n4401 19.3944
R16960 GND.n4401 GND.n2027 19.3944
R16961 GND.n4475 GND.n2027 19.3944
R16962 GND.n4475 GND.n2024 19.3944
R16963 GND.n4492 GND.n2024 19.3944
R16964 GND.n4492 GND.n2025 19.3944
R16965 GND.n4488 GND.n2025 19.3944
R16966 GND.n4488 GND.n4487 19.3944
R16967 GND.n4487 GND.n4486 19.3944
R16968 GND.n4486 GND.n4483 19.3944
R16969 GND.n4483 GND.n1965 19.3944
R16970 GND.n4593 GND.n1965 19.3944
R16971 GND.n4593 GND.n1962 19.3944
R16972 GND.n4603 GND.n1962 19.3944
R16973 GND.n4603 GND.n1963 19.3944
R16974 GND.n4599 GND.n1963 19.3944
R16975 GND.n4599 GND.n1935 19.3944
R16976 GND.n4626 GND.n1935 19.3944
R16977 GND.n4627 GND.n4626 19.3944
R16978 GND.n4627 GND.n1933 19.3944
R16979 GND.n4631 GND.n1933 19.3944
R16980 GND.n4631 GND.n1918 19.3944
R16981 GND.n4643 GND.n1918 19.3944
R16982 GND.n4643 GND.n1916 19.3944
R16983 GND.n4650 GND.n1916 19.3944
R16984 GND.n4650 GND.n4649 19.3944
R16985 GND.n4649 GND.n1862 19.3944
R16986 GND.n4696 GND.n1862 19.3944
R16987 GND.n4696 GND.n1860 19.3944
R16988 GND.n4702 GND.n1860 19.3944
R16989 GND.n4702 GND.n4701 19.3944
R16990 GND.n4701 GND.n1825 19.3944
R16991 GND.n4752 GND.n1825 19.3944
R16992 GND.n4752 GND.n1823 19.3944
R16993 GND.n4758 GND.n1823 19.3944
R16994 GND.n4758 GND.n4757 19.3944
R16995 GND.n4757 GND.n1797 19.3944
R16996 GND.n4790 GND.n1797 19.3944
R16997 GND.n4790 GND.n1795 19.3944
R16998 GND.n4796 GND.n1795 19.3944
R16999 GND.n4796 GND.n4795 19.3944
R17000 GND.n4795 GND.n1764 19.3944
R17001 GND.n4858 GND.n1764 19.3944
R17002 GND.n4858 GND.n1762 19.3944
R17003 GND.n4864 GND.n1762 19.3944
R17004 GND.n4864 GND.n4863 19.3944
R17005 GND.n4863 GND.n1736 19.3944
R17006 GND.n4895 GND.n1736 19.3944
R17007 GND.n4895 GND.n1734 19.3944
R17008 GND.n4910 GND.n1734 19.3944
R17009 GND.n4910 GND.n4909 19.3944
R17010 GND.n4909 GND.n4908 19.3944
R17011 GND.n4908 GND.n4906 19.3944
R17012 GND.n4906 GND.n4905 19.3944
R17013 GND.n4905 GND.n4904 19.3944
R17014 GND.n4904 GND.n1680 19.3944
R17015 GND.n5892 GND.n1680 19.3944
R17016 GND.n5892 GND.n1678 19.3944
R17017 GND.n5897 GND.n1678 19.3944
R17018 GND.n5897 GND.n5896 19.3944
R17019 GND.n4327 GND.n4326 19.3944
R17020 GND.n4326 GND.n4325 19.3944
R17021 GND.n4325 GND.n2141 19.3944
R17022 GND.n4321 GND.n2141 19.3944
R17023 GND.n4321 GND.n4320 19.3944
R17024 GND.n4320 GND.n4319 19.3944
R17025 GND.n4341 GND.n4340 19.3944
R17026 GND.n4340 GND.n4339 19.3944
R17027 GND.n4339 GND.n2112 19.3944
R17028 GND.n4366 GND.n2112 19.3944
R17029 GND.n4377 GND.n4366 19.3944
R17030 GND.n4377 GND.n4376 19.3944
R17031 GND.n4376 GND.n4375 19.3944
R17032 GND.n4375 GND.n2083 19.3944
R17033 GND.n4414 GND.n2083 19.3944
R17034 GND.n4420 GND.n4414 19.3944
R17035 GND.n4420 GND.n4419 19.3944
R17036 GND.n4419 GND.n4418 19.3944
R17037 GND.n4418 GND.n2049 19.3944
R17038 GND.n4459 GND.n2049 19.3944
R17039 GND.n4459 GND.n4458 19.3944
R17040 GND.n4458 GND.n4457 19.3944
R17041 GND.n4457 GND.n2021 19.3944
R17042 GND.n4496 GND.n2021 19.3944
R17043 GND.n4502 GND.n4496 19.3944
R17044 GND.n4502 GND.n4501 19.3944
R17045 GND.n4501 GND.n4500 19.3944
R17046 GND.n4500 GND.n1987 19.3944
R17047 GND.n4577 GND.n1987 19.3944
R17048 GND.n4577 GND.n4576 19.3944
R17049 GND.n4576 GND.n4575 19.3944
R17050 GND.n4575 GND.n1959 19.3944
R17051 GND.n4607 GND.n1959 19.3944
R17052 GND.n4609 GND.n4607 19.3944
R17053 GND.n4609 GND.n4608 19.3944
R17054 GND.n4608 GND.n1939 19.3944
R17055 GND.n1939 GND.n1892 19.3944
R17056 GND.n4681 GND.n1892 19.3944
R17057 GND.n4681 GND.n4680 19.3944
R17058 GND.n4680 GND.n4679 19.3944
R17059 GND.n4679 GND.n1895 19.3944
R17060 GND.n4675 GND.n1895 19.3944
R17061 GND.n4675 GND.n4674 19.3944
R17062 GND.n4674 GND.n4673 19.3944
R17063 GND.n4673 GND.n1903 19.3944
R17064 GND.n4669 GND.n1903 19.3944
R17065 GND.n4669 GND.n4668 19.3944
R17066 GND.n4668 GND.n4667 19.3944
R17067 GND.n4667 GND.n1846 19.3944
R17068 GND.n4736 GND.n1846 19.3944
R17069 GND.n4736 GND.n4735 19.3944
R17070 GND.n4735 GND.n4734 19.3944
R17071 GND.n4734 GND.n1819 19.3944
R17072 GND.n4762 GND.n1819 19.3944
R17073 GND.n4774 GND.n4762 19.3944
R17074 GND.n4774 GND.n4773 19.3944
R17075 GND.n4773 GND.n4772 19.3944
R17076 GND.n4772 GND.n4766 19.3944
R17077 GND.n4766 GND.n1785 19.3944
R17078 GND.n4842 GND.n1785 19.3944
R17079 GND.n4842 GND.n4841 19.3944
R17080 GND.n4841 GND.n4840 19.3944
R17081 GND.n4840 GND.n1758 19.3944
R17082 GND.n4868 GND.n1758 19.3944
R17083 GND.n4879 GND.n4868 19.3944
R17084 GND.n4879 GND.n4878 19.3944
R17085 GND.n4878 GND.n4877 19.3944
R17086 GND.n4877 GND.n1730 19.3944
R17087 GND.n4914 GND.n1730 19.3944
R17088 GND.n4917 GND.n4914 19.3944
R17089 GND.n4917 GND.n4916 19.3944
R17090 GND.n4916 GND.n1700 19.3944
R17091 GND.n5863 GND.n1700 19.3944
R17092 GND.n5877 GND.n5863 19.3944
R17093 GND.n5877 GND.n5876 19.3944
R17094 GND.n5876 GND.n5875 19.3944
R17095 GND.n5875 GND.n5866 19.3944
R17096 GND.n5866 GND.n1604 19.3944
R17097 GND.n6048 GND.n1604 19.3944
R17098 GND.n5909 GND.n5906 19.3944
R17099 GND.n5909 GND.n1672 19.3944
R17100 GND.n5913 GND.n1672 19.3944
R17101 GND.n5916 GND.n5913 19.3944
R17102 GND.n5919 GND.n5916 19.3944
R17103 GND.n5919 GND.n1670 19.3944
R17104 GND.n5923 GND.n1670 19.3944
R17105 GND.n5931 GND.n1668 19.3944
R17106 GND.n5935 GND.n1668 19.3944
R17107 GND.n5938 GND.n5935 19.3944
R17108 GND.n5941 GND.n5938 19.3944
R17109 GND.n5941 GND.n1666 19.3944
R17110 GND.n5945 GND.n1666 19.3944
R17111 GND.n5948 GND.n5945 19.3944
R17112 GND.n5950 GND.n5948 19.3944
R17113 GND.n5954 GND.n5953 19.3944
R17114 GND.n5957 GND.n5954 19.3944
R17115 GND.n6039 GND.n1659 19.3944
R17116 GND.n6035 GND.n1659 19.3944
R17117 GND.n6035 GND.n6034 19.3944
R17118 GND.n6032 GND.n5970 19.3944
R17119 GND.n6028 GND.n5970 19.3944
R17120 GND.n6028 GND.n6027 19.3944
R17121 GND.n6027 GND.n6026 19.3944
R17122 GND.n6026 GND.n5976 19.3944
R17123 GND.n6022 GND.n5976 19.3944
R17124 GND.n6022 GND.n6021 19.3944
R17125 GND.n6021 GND.n6020 19.3944
R17126 GND.n6016 GND.n6015 19.3944
R17127 GND.n6015 GND.n6014 19.3944
R17128 GND.n6014 GND.n5990 19.3944
R17129 GND.n6010 GND.n5990 19.3944
R17130 GND.n6010 GND.n6009 19.3944
R17131 GND.n6009 GND.n6008 19.3944
R17132 GND.n6008 GND.n5996 19.3944
R17133 GND.n6004 GND.n5996 19.3944
R17134 GND.n3212 GND.n3211 19.3944
R17135 GND.n3211 GND.n2970 19.3944
R17136 GND.n3207 GND.n2970 19.3944
R17137 GND.n3207 GND.n2972 19.3944
R17138 GND.n3201 GND.n2972 19.3944
R17139 GND.n3201 GND.n3200 19.3944
R17140 GND.n3200 GND.n3199 19.3944
R17141 GND.n3199 GND.n2981 19.3944
R17142 GND.n3193 GND.n2981 19.3944
R17143 GND.n3193 GND.n3192 19.3944
R17144 GND.n3192 GND.n3191 19.3944
R17145 GND.n3191 GND.n2989 19.3944
R17146 GND.n3185 GND.n2989 19.3944
R17147 GND.n3185 GND.n3184 19.3944
R17148 GND.n3184 GND.n3183 19.3944
R17149 GND.n3183 GND.n2997 19.3944
R17150 GND.n3177 GND.n2997 19.3944
R17151 GND.n3177 GND.n3176 19.3944
R17152 GND.n3176 GND.n3175 19.3944
R17153 GND.n3175 GND.n3005 19.3944
R17154 GND.n3169 GND.n3005 19.3944
R17155 GND.n3169 GND.n3168 19.3944
R17156 GND.n3168 GND.n3167 19.3944
R17157 GND.n3167 GND.n3013 19.3944
R17158 GND.n3161 GND.n3013 19.3944
R17159 GND.n3161 GND.n3160 19.3944
R17160 GND.n3160 GND.n3159 19.3944
R17161 GND.n3159 GND.n3021 19.3944
R17162 GND.n3153 GND.n3021 19.3944
R17163 GND.n3153 GND.n3152 19.3944
R17164 GND.n3152 GND.n3151 19.3944
R17165 GND.n3151 GND.n3029 19.3944
R17166 GND.n3145 GND.n3029 19.3944
R17167 GND.n3145 GND.n3144 19.3944
R17168 GND.n3144 GND.n3143 19.3944
R17169 GND.n3143 GND.n3037 19.3944
R17170 GND.n3137 GND.n3037 19.3944
R17171 GND.n3137 GND.n3136 19.3944
R17172 GND.n3136 GND.n3135 19.3944
R17173 GND.n3135 GND.n3045 19.3944
R17174 GND.n3129 GND.n3045 19.3944
R17175 GND.n3129 GND.n3128 19.3944
R17176 GND.n3128 GND.n3127 19.3944
R17177 GND.n3127 GND.n3053 19.3944
R17178 GND.n3121 GND.n3053 19.3944
R17179 GND.n3121 GND.n3120 19.3944
R17180 GND.n3120 GND.n3119 19.3944
R17181 GND.n3119 GND.n3061 19.3944
R17182 GND.n3113 GND.n3061 19.3944
R17183 GND.n3113 GND.n3112 19.3944
R17184 GND.n3112 GND.n3111 19.3944
R17185 GND.n3111 GND.n3069 19.3944
R17186 GND.n3105 GND.n3069 19.3944
R17187 GND.n3105 GND.n3104 19.3944
R17188 GND.n3104 GND.n3103 19.3944
R17189 GND.n3103 GND.n3077 19.3944
R17190 GND.n3097 GND.n3077 19.3944
R17191 GND.n3097 GND.n3096 19.3944
R17192 GND.n3096 GND.n3095 19.3944
R17193 GND.n3095 GND.n3085 19.3944
R17194 GND.n3089 GND.n3085 19.3944
R17195 GND.n3089 GND.n384 19.3944
R17196 GND.n8263 GND.n384 19.3944
R17197 GND.n3934 GND.n2251 19.3944
R17198 GND.n3930 GND.n2251 19.3944
R17199 GND.n3930 GND.n2253 19.3944
R17200 GND.n3924 GND.n2253 19.3944
R17201 GND.n3924 GND.n3923 19.3944
R17202 GND.n3923 GND.n3922 19.3944
R17203 GND.n3922 GND.n2260 19.3944
R17204 GND.n3916 GND.n2260 19.3944
R17205 GND.n3916 GND.n3915 19.3944
R17206 GND.n3915 GND.n3914 19.3944
R17207 GND.n3914 GND.n2268 19.3944
R17208 GND.n3908 GND.n2268 19.3944
R17209 GND.n3908 GND.n3907 19.3944
R17210 GND.n3907 GND.n3906 19.3944
R17211 GND.n3906 GND.n2276 19.3944
R17212 GND.n3900 GND.n2276 19.3944
R17213 GND.n3900 GND.n3899 19.3944
R17214 GND.n3899 GND.n3898 19.3944
R17215 GND.n3898 GND.n2284 19.3944
R17216 GND.n3892 GND.n2284 19.3944
R17217 GND.n3892 GND.n3891 19.3944
R17218 GND.n3891 GND.n3890 19.3944
R17219 GND.n3890 GND.n2292 19.3944
R17220 GND.n3884 GND.n2292 19.3944
R17221 GND.n3884 GND.n3883 19.3944
R17222 GND.n3883 GND.n3882 19.3944
R17223 GND.n3882 GND.n2300 19.3944
R17224 GND.n3876 GND.n2300 19.3944
R17225 GND.n3876 GND.n3875 19.3944
R17226 GND.n3875 GND.n3874 19.3944
R17227 GND.n3874 GND.n2308 19.3944
R17228 GND.n3868 GND.n2308 19.3944
R17229 GND.n3868 GND.n3867 19.3944
R17230 GND.n3867 GND.n3866 19.3944
R17231 GND.n3866 GND.n2316 19.3944
R17232 GND.n3860 GND.n2316 19.3944
R17233 GND.n3860 GND.n3859 19.3944
R17234 GND.n3859 GND.n3858 19.3944
R17235 GND.n3858 GND.n2324 19.3944
R17236 GND.n3852 GND.n2324 19.3944
R17237 GND.n3852 GND.n3851 19.3944
R17238 GND.n3851 GND.n3850 19.3944
R17239 GND.n3850 GND.n2332 19.3944
R17240 GND.n3844 GND.n2332 19.3944
R17241 GND.n3844 GND.n3843 19.3944
R17242 GND.n3843 GND.n3842 19.3944
R17243 GND.n3842 GND.n2340 19.3944
R17244 GND.n3836 GND.n2340 19.3944
R17245 GND.n3836 GND.n3835 19.3944
R17246 GND.n3835 GND.n3834 19.3944
R17247 GND.n3834 GND.n2348 19.3944
R17248 GND.n3828 GND.n2348 19.3944
R17249 GND.n3828 GND.n3827 19.3944
R17250 GND.n3827 GND.n3826 19.3944
R17251 GND.n3826 GND.n2356 19.3944
R17252 GND.n3820 GND.n2356 19.3944
R17253 GND.n3820 GND.n3819 19.3944
R17254 GND.n3819 GND.n3818 19.3944
R17255 GND.n3818 GND.n2364 19.3944
R17256 GND.n3812 GND.n2364 19.3944
R17257 GND.n3812 GND.n3811 19.3944
R17258 GND.n3811 GND.n3810 19.3944
R17259 GND.n3810 GND.n2372 19.3944
R17260 GND.n3804 GND.n2372 19.3944
R17261 GND.n3804 GND.n3803 19.3944
R17262 GND.n3803 GND.n3802 19.3944
R17263 GND.n3802 GND.n2380 19.3944
R17264 GND.n3796 GND.n2380 19.3944
R17265 GND.n3796 GND.n3795 19.3944
R17266 GND.n3795 GND.n3794 19.3944
R17267 GND.n3794 GND.n2388 19.3944
R17268 GND.n3788 GND.n2388 19.3944
R17269 GND.n3788 GND.n3787 19.3944
R17270 GND.n3787 GND.n3786 19.3944
R17271 GND.n3786 GND.n2396 19.3944
R17272 GND.n3780 GND.n2396 19.3944
R17273 GND.n3780 GND.n3779 19.3944
R17274 GND.n3779 GND.n3778 19.3944
R17275 GND.n3778 GND.n2404 19.3944
R17276 GND.n3772 GND.n2404 19.3944
R17277 GND.n3772 GND.n3771 19.3944
R17278 GND.n3771 GND.n3770 19.3944
R17279 GND.n3770 GND.n2412 19.3944
R17280 GND.n3764 GND.n2412 19.3944
R17281 GND.n3764 GND.n3763 19.3944
R17282 GND.n3763 GND.n3762 19.3944
R17283 GND.n3762 GND.n2420 19.3944
R17284 GND.n3756 GND.n2420 19.3944
R17285 GND.n3756 GND.n3755 19.3944
R17286 GND.n3755 GND.n3754 19.3944
R17287 GND.n3754 GND.n2428 19.3944
R17288 GND.n3748 GND.n2428 19.3944
R17289 GND.n3748 GND.n3747 19.3944
R17290 GND.n3747 GND.n3746 19.3944
R17291 GND.n3746 GND.n2436 19.3944
R17292 GND.n3740 GND.n2436 19.3944
R17293 GND.n3740 GND.n3739 19.3944
R17294 GND.n3739 GND.n3738 19.3944
R17295 GND.n3738 GND.n2444 19.3944
R17296 GND.n3732 GND.n2444 19.3944
R17297 GND.n3732 GND.n3731 19.3944
R17298 GND.n3731 GND.n3730 19.3944
R17299 GND.n3730 GND.n2452 19.3944
R17300 GND.n3724 GND.n2452 19.3944
R17301 GND.n3724 GND.n3723 19.3944
R17302 GND.n3723 GND.n3722 19.3944
R17303 GND.n3722 GND.n2460 19.3944
R17304 GND.n3716 GND.n2460 19.3944
R17305 GND.n3716 GND.n3715 19.3944
R17306 GND.n3715 GND.n3714 19.3944
R17307 GND.n3714 GND.n2468 19.3944
R17308 GND.n3708 GND.n2468 19.3944
R17309 GND.n3708 GND.n3707 19.3944
R17310 GND.n3707 GND.n3706 19.3944
R17311 GND.n3706 GND.n2476 19.3944
R17312 GND.n3700 GND.n2476 19.3944
R17313 GND.n3700 GND.n3699 19.3944
R17314 GND.n3699 GND.n3698 19.3944
R17315 GND.n3698 GND.n2484 19.3944
R17316 GND.n3692 GND.n2484 19.3944
R17317 GND.n3692 GND.n3691 19.3944
R17318 GND.n3691 GND.n3690 19.3944
R17319 GND.n3690 GND.n2492 19.3944
R17320 GND.n3684 GND.n2492 19.3944
R17321 GND.n3684 GND.n3683 19.3944
R17322 GND.n3683 GND.n3682 19.3944
R17323 GND.n3682 GND.n2500 19.3944
R17324 GND.n3676 GND.n2500 19.3944
R17325 GND.n3676 GND.n3675 19.3944
R17326 GND.n3675 GND.n3674 19.3944
R17327 GND.n3674 GND.n2508 19.3944
R17328 GND.n3668 GND.n2508 19.3944
R17329 GND.n3668 GND.n3667 19.3944
R17330 GND.n3667 GND.n3666 19.3944
R17331 GND.n3666 GND.n2516 19.3944
R17332 GND.n3660 GND.n2516 19.3944
R17333 GND.n3660 GND.n3659 19.3944
R17334 GND.n3659 GND.n3658 19.3944
R17335 GND.n3658 GND.n2524 19.3944
R17336 GND.n3652 GND.n2524 19.3944
R17337 GND.n3652 GND.n3651 19.3944
R17338 GND.n3651 GND.n3650 19.3944
R17339 GND.n3650 GND.n2532 19.3944
R17340 GND.n3644 GND.n2532 19.3944
R17341 GND.n3644 GND.n3643 19.3944
R17342 GND.n3643 GND.n3642 19.3944
R17343 GND.n3642 GND.n2540 19.3944
R17344 GND.n3636 GND.n2540 19.3944
R17345 GND.n3636 GND.n3635 19.3944
R17346 GND.n3635 GND.n3634 19.3944
R17347 GND.n3634 GND.n2548 19.3944
R17348 GND.n3628 GND.n2548 19.3944
R17349 GND.n3628 GND.n3627 19.3944
R17350 GND.n3627 GND.n3626 19.3944
R17351 GND.n3626 GND.n2556 19.3944
R17352 GND.n3620 GND.n2556 19.3944
R17353 GND.n3620 GND.n3619 19.3944
R17354 GND.n3619 GND.n3618 19.3944
R17355 GND.n3618 GND.n2564 19.3944
R17356 GND.n3612 GND.n2564 19.3944
R17357 GND.n3612 GND.n3611 19.3944
R17358 GND.n3611 GND.n3610 19.3944
R17359 GND.n3610 GND.n2572 19.3944
R17360 GND.n3604 GND.n2572 19.3944
R17361 GND.n3604 GND.n3603 19.3944
R17362 GND.n3603 GND.n3602 19.3944
R17363 GND.n3602 GND.n2580 19.3944
R17364 GND.n3596 GND.n2580 19.3944
R17365 GND.n3596 GND.n3595 19.3944
R17366 GND.n3595 GND.n3594 19.3944
R17367 GND.n3594 GND.n2588 19.3944
R17368 GND.n3588 GND.n2588 19.3944
R17369 GND.n3588 GND.n3587 19.3944
R17370 GND.n3587 GND.n3586 19.3944
R17371 GND.n3586 GND.n2596 19.3944
R17372 GND.n3580 GND.n2596 19.3944
R17373 GND.n3580 GND.n3579 19.3944
R17374 GND.n3579 GND.n3578 19.3944
R17375 GND.n3578 GND.n2604 19.3944
R17376 GND.n3572 GND.n2604 19.3944
R17377 GND.n3572 GND.n3571 19.3944
R17378 GND.n3571 GND.n3570 19.3944
R17379 GND.n3570 GND.n2612 19.3944
R17380 GND.n3564 GND.n2612 19.3944
R17381 GND.n3564 GND.n3563 19.3944
R17382 GND.n3563 GND.n3562 19.3944
R17383 GND.n3562 GND.n2620 19.3944
R17384 GND.n3556 GND.n2620 19.3944
R17385 GND.n3556 GND.n3555 19.3944
R17386 GND.n3555 GND.n3554 19.3944
R17387 GND.n3554 GND.n2628 19.3944
R17388 GND.n3548 GND.n2628 19.3944
R17389 GND.n3548 GND.n3547 19.3944
R17390 GND.n3547 GND.n3546 19.3944
R17391 GND.n3546 GND.n2636 19.3944
R17392 GND.n3540 GND.n2636 19.3944
R17393 GND.n3540 GND.n3539 19.3944
R17394 GND.n3539 GND.n3538 19.3944
R17395 GND.n3538 GND.n2644 19.3944
R17396 GND.n3532 GND.n2644 19.3944
R17397 GND.n3532 GND.n3531 19.3944
R17398 GND.n3531 GND.n3530 19.3944
R17399 GND.n3530 GND.n2652 19.3944
R17400 GND.n3524 GND.n2652 19.3944
R17401 GND.n3524 GND.n3523 19.3944
R17402 GND.n3523 GND.n3522 19.3944
R17403 GND.n3522 GND.n2660 19.3944
R17404 GND.n3516 GND.n2660 19.3944
R17405 GND.n3516 GND.n3515 19.3944
R17406 GND.n3515 GND.n3514 19.3944
R17407 GND.n3514 GND.n2668 19.3944
R17408 GND.n3508 GND.n2668 19.3944
R17409 GND.n3508 GND.n3507 19.3944
R17410 GND.n3507 GND.n3506 19.3944
R17411 GND.n3506 GND.n2676 19.3944
R17412 GND.n3500 GND.n2676 19.3944
R17413 GND.n3500 GND.n3499 19.3944
R17414 GND.n3499 GND.n3498 19.3944
R17415 GND.n3498 GND.n2684 19.3944
R17416 GND.n3492 GND.n2684 19.3944
R17417 GND.n3492 GND.n3491 19.3944
R17418 GND.n3491 GND.n3490 19.3944
R17419 GND.n3490 GND.n2692 19.3944
R17420 GND.n3484 GND.n2692 19.3944
R17421 GND.n3484 GND.n3483 19.3944
R17422 GND.n3483 GND.n3482 19.3944
R17423 GND.n3482 GND.n2700 19.3944
R17424 GND.n3476 GND.n2700 19.3944
R17425 GND.n3476 GND.n3475 19.3944
R17426 GND.n3475 GND.n3474 19.3944
R17427 GND.n3474 GND.n2708 19.3944
R17428 GND.n3468 GND.n2708 19.3944
R17429 GND.n3468 GND.n3467 19.3944
R17430 GND.n3467 GND.n3466 19.3944
R17431 GND.n3466 GND.n2716 19.3944
R17432 GND.n3460 GND.n2716 19.3944
R17433 GND.n3460 GND.n3459 19.3944
R17434 GND.n3459 GND.n3458 19.3944
R17435 GND.n3458 GND.n2724 19.3944
R17436 GND.n3452 GND.n2724 19.3944
R17437 GND.n3452 GND.n3451 19.3944
R17438 GND.n3451 GND.n3450 19.3944
R17439 GND.n3450 GND.n2732 19.3944
R17440 GND.n3444 GND.n2732 19.3944
R17441 GND.n3444 GND.n3443 19.3944
R17442 GND.n3443 GND.n3442 19.3944
R17443 GND.n3442 GND.n2740 19.3944
R17444 GND.n3436 GND.n2740 19.3944
R17445 GND.n3436 GND.n3435 19.3944
R17446 GND.n3435 GND.n3434 19.3944
R17447 GND.n3434 GND.n2748 19.3944
R17448 GND.n3428 GND.n2748 19.3944
R17449 GND.n3428 GND.n3427 19.3944
R17450 GND.n3427 GND.n3426 19.3944
R17451 GND.n3426 GND.n2756 19.3944
R17452 GND.n3420 GND.n2756 19.3944
R17453 GND.n3420 GND.n3419 19.3944
R17454 GND.n3419 GND.n3418 19.3944
R17455 GND.n3418 GND.n2764 19.3944
R17456 GND.n3412 GND.n2764 19.3944
R17457 GND.n3412 GND.n3411 19.3944
R17458 GND.n3411 GND.n3410 19.3944
R17459 GND.n3410 GND.n2772 19.3944
R17460 GND.n3404 GND.n2772 19.3944
R17461 GND.n3404 GND.n3403 19.3944
R17462 GND.n3403 GND.n3402 19.3944
R17463 GND.n3402 GND.n2780 19.3944
R17464 GND.n3396 GND.n2780 19.3944
R17465 GND.n3396 GND.n3395 19.3944
R17466 GND.n3395 GND.n3394 19.3944
R17467 GND.n3394 GND.n2788 19.3944
R17468 GND.n3388 GND.n2788 19.3944
R17469 GND.n3388 GND.n3387 19.3944
R17470 GND.n3387 GND.n3386 19.3944
R17471 GND.n3386 GND.n2796 19.3944
R17472 GND.n3380 GND.n2796 19.3944
R17473 GND.n3380 GND.n3379 19.3944
R17474 GND.n3379 GND.n3378 19.3944
R17475 GND.n3378 GND.n2804 19.3944
R17476 GND.n3372 GND.n2804 19.3944
R17477 GND.n3372 GND.n3371 19.3944
R17478 GND.n3371 GND.n3370 19.3944
R17479 GND.n3370 GND.n2812 19.3944
R17480 GND.n3364 GND.n2812 19.3944
R17481 GND.n3364 GND.n3363 19.3944
R17482 GND.n3363 GND.n3362 19.3944
R17483 GND.n3362 GND.n2820 19.3944
R17484 GND.n3356 GND.n2820 19.3944
R17485 GND.n3356 GND.n3355 19.3944
R17486 GND.n3355 GND.n3354 19.3944
R17487 GND.n3354 GND.n2828 19.3944
R17488 GND.n3348 GND.n2828 19.3944
R17489 GND.n3348 GND.n3347 19.3944
R17490 GND.n3347 GND.n3346 19.3944
R17491 GND.n3346 GND.n2836 19.3944
R17492 GND.n3340 GND.n2836 19.3944
R17493 GND.n3340 GND.n3339 19.3944
R17494 GND.n3339 GND.n3338 19.3944
R17495 GND.n3338 GND.n2844 19.3944
R17496 GND.n3332 GND.n2844 19.3944
R17497 GND.n3332 GND.n3331 19.3944
R17498 GND.n3331 GND.n3330 19.3944
R17499 GND.n3330 GND.n2852 19.3944
R17500 GND.n3324 GND.n2852 19.3944
R17501 GND.n3324 GND.n3323 19.3944
R17502 GND.n3323 GND.n3322 19.3944
R17503 GND.n3322 GND.n2860 19.3944
R17504 GND.n3316 GND.n2860 19.3944
R17505 GND.n3316 GND.n3315 19.3944
R17506 GND.n3315 GND.n3314 19.3944
R17507 GND.n3314 GND.n2868 19.3944
R17508 GND.n3308 GND.n2868 19.3944
R17509 GND.n3308 GND.n3307 19.3944
R17510 GND.n3307 GND.n3306 19.3944
R17511 GND.n3306 GND.n2876 19.3944
R17512 GND.n3300 GND.n2876 19.3944
R17513 GND.n3300 GND.n3299 19.3944
R17514 GND.n3299 GND.n3298 19.3944
R17515 GND.n3298 GND.n2884 19.3944
R17516 GND.n3292 GND.n2884 19.3944
R17517 GND.n3292 GND.n3291 19.3944
R17518 GND.n3291 GND.n3290 19.3944
R17519 GND.n3290 GND.n2892 19.3944
R17520 GND.n3284 GND.n2892 19.3944
R17521 GND.n3284 GND.n3283 19.3944
R17522 GND.n3283 GND.n3282 19.3944
R17523 GND.n3282 GND.n2900 19.3944
R17524 GND.n3276 GND.n2900 19.3944
R17525 GND.n3276 GND.n3275 19.3944
R17526 GND.n3275 GND.n3274 19.3944
R17527 GND.n3274 GND.n2908 19.3944
R17528 GND.n3268 GND.n2908 19.3944
R17529 GND.n3268 GND.n3267 19.3944
R17530 GND.n3267 GND.n3266 19.3944
R17531 GND.n3266 GND.n2916 19.3944
R17532 GND.n3260 GND.n2916 19.3944
R17533 GND.n3260 GND.n3259 19.3944
R17534 GND.n3259 GND.n3258 19.3944
R17535 GND.n3258 GND.n2924 19.3944
R17536 GND.n3252 GND.n2924 19.3944
R17537 GND.n3252 GND.n3251 19.3944
R17538 GND.n3251 GND.n3250 19.3944
R17539 GND.n3250 GND.n2932 19.3944
R17540 GND.n3244 GND.n2932 19.3944
R17541 GND.n3244 GND.n3243 19.3944
R17542 GND.n3243 GND.n3242 19.3944
R17543 GND.n3242 GND.n2940 19.3944
R17544 GND.n3236 GND.n2940 19.3944
R17545 GND.n3236 GND.n3235 19.3944
R17546 GND.n3235 GND.n3234 19.3944
R17547 GND.n3234 GND.n2948 19.3944
R17548 GND.n3228 GND.n2948 19.3944
R17549 GND.n3228 GND.n3227 19.3944
R17550 GND.n3227 GND.n3226 19.3944
R17551 GND.n3226 GND.n2956 19.3944
R17552 GND.n3220 GND.n2956 19.3944
R17553 GND.n3220 GND.n3219 19.3944
R17554 GND.n3219 GND.n3218 19.3944
R17555 GND.n3218 GND.n2964 19.3944
R17556 GND.n7722 GND.n7721 19.3944
R17557 GND.n7721 GND.n7720 19.3944
R17558 GND.n7720 GND.n7719 19.3944
R17559 GND.n7719 GND.n7717 19.3944
R17560 GND.n7717 GND.n7714 19.3944
R17561 GND.n7714 GND.n7713 19.3944
R17562 GND.n7713 GND.n7710 19.3944
R17563 GND.n7708 GND.n7706 19.3944
R17564 GND.n7706 GND.n7703 19.3944
R17565 GND.n7703 GND.n7702 19.3944
R17566 GND.n7702 GND.n7699 19.3944
R17567 GND.n7699 GND.n7698 19.3944
R17568 GND.n7698 GND.n7695 19.3944
R17569 GND.n7695 GND.n7694 19.3944
R17570 GND.n7694 GND.n7691 19.3944
R17571 GND.n7689 GND.n7686 19.3944
R17572 GND.n7686 GND.n7685 19.3944
R17573 GND.n7681 GND.n7679 19.3944
R17574 GND.n7679 GND.n7676 19.3944
R17575 GND.n7676 GND.n7675 19.3944
R17576 GND.n7671 GND.n7668 19.3944
R17577 GND.n7668 GND.n7667 19.3944
R17578 GND.n7667 GND.n7664 19.3944
R17579 GND.n7664 GND.n7663 19.3944
R17580 GND.n7663 GND.n7660 19.3944
R17581 GND.n7660 GND.n7659 19.3944
R17582 GND.n7659 GND.n7656 19.3944
R17583 GND.n7656 GND.n7655 19.3944
R17584 GND.n7651 GND.n7648 19.3944
R17585 GND.n7648 GND.n7647 19.3944
R17586 GND.n7647 GND.n7644 19.3944
R17587 GND.n7644 GND.n7643 19.3944
R17588 GND.n7643 GND.n7640 19.3944
R17589 GND.n7640 GND.n7639 19.3944
R17590 GND.n7639 GND.n7636 19.3944
R17591 GND.n7636 GND.n7635 19.3944
R17592 GND.n7750 GND.n7739 19.3944
R17593 GND.n7750 GND.n7749 19.3944
R17594 GND.n7749 GND.n7746 19.3944
R17595 GND.n7746 GND.n628 19.3944
R17596 GND.n7776 GND.n628 19.3944
R17597 GND.n7777 GND.n7776 19.3944
R17598 GND.n7780 GND.n7777 19.3944
R17599 GND.n7781 GND.n7780 19.3944
R17600 GND.n7781 GND.n600 19.3944
R17601 GND.n7817 GND.n600 19.3944
R17602 GND.n7818 GND.n7817 19.3944
R17603 GND.n7819 GND.n7818 19.3944
R17604 GND.n7819 GND.n584 19.3944
R17605 GND.n584 GND.n577 19.3944
R17606 GND.n7849 GND.n577 19.3944
R17607 GND.n7849 GND.n7848 19.3944
R17608 GND.n7848 GND.n560 19.3944
R17609 GND.n7867 GND.n560 19.3944
R17610 GND.n7867 GND.n7866 19.3944
R17611 GND.n7866 GND.n547 19.3944
R17612 GND.n7885 GND.n547 19.3944
R17613 GND.n7885 GND.n7884 19.3944
R17614 GND.n7884 GND.n552 19.3944
R17615 GND.n552 GND.n551 19.3944
R17616 GND.n551 GND.n548 19.3944
R17617 GND.n548 GND.n487 19.3944
R17618 GND.n7966 GND.n487 19.3944
R17619 GND.n7967 GND.n7966 19.3944
R17620 GND.n7970 GND.n7967 19.3944
R17621 GND.n7971 GND.n7970 19.3944
R17622 GND.n7971 GND.n460 19.3944
R17623 GND.n8008 GND.n460 19.3944
R17624 GND.n8009 GND.n8008 19.3944
R17625 GND.n8009 GND.n446 19.3944
R17626 GND.n8023 GND.n446 19.3944
R17627 GND.n8024 GND.n8023 19.3944
R17628 GND.n8027 GND.n8024 19.3944
R17629 GND.n8027 GND.n8026 19.3944
R17630 GND.n8026 GND.n431 19.3944
R17631 GND.n8130 GND.n431 19.3944
R17632 GND.n8130 GND.n424 19.3944
R17633 GND.n8142 GND.n424 19.3944
R17634 GND.n8143 GND.n8142 19.3944
R17635 GND.n8145 GND.n8143 19.3944
R17636 GND.n8145 GND.n420 19.3944
R17637 GND.n8157 GND.n420 19.3944
R17638 GND.n8158 GND.n8157 19.3944
R17639 GND.n8160 GND.n8158 19.3944
R17640 GND.n8160 GND.n416 19.3944
R17641 GND.n8172 GND.n416 19.3944
R17642 GND.n8173 GND.n8172 19.3944
R17643 GND.n8175 GND.n8173 19.3944
R17644 GND.n8175 GND.n412 19.3944
R17645 GND.n8187 GND.n412 19.3944
R17646 GND.n8188 GND.n8187 19.3944
R17647 GND.n8190 GND.n8188 19.3944
R17648 GND.n8190 GND.n407 19.3944
R17649 GND.n8202 GND.n407 19.3944
R17650 GND.n8203 GND.n8202 19.3944
R17651 GND.n8205 GND.n8203 19.3944
R17652 GND.n8205 GND.n403 19.3944
R17653 GND.n8217 GND.n403 19.3944
R17654 GND.n8218 GND.n8217 19.3944
R17655 GND.n8220 GND.n8218 19.3944
R17656 GND.n8220 GND.n399 19.3944
R17657 GND.n8233 GND.n399 19.3944
R17658 GND.n8234 GND.n8233 19.3944
R17659 GND.n8236 GND.n8234 19.3944
R17660 GND.n8237 GND.n8236 19.3944
R17661 GND.n8238 GND.n8237 19.3944
R17662 GND.n8238 GND.n350 19.3944
R17663 GND.n8458 GND.n350 19.3944
R17664 GND.n8459 GND.n8458 19.3944
R17665 GND.n7752 GND.n653 19.3944
R17666 GND.n7752 GND.n654 19.3944
R17667 GND.n7740 GND.n654 19.3944
R17668 GND.n7743 GND.n7740 19.3944
R17669 GND.n7743 GND.n625 19.3944
R17670 GND.n7789 GND.n625 19.3944
R17671 GND.n7789 GND.n7788 19.3944
R17672 GND.n7788 GND.n7787 19.3944
R17673 GND.n7787 GND.n7786 19.3944
R17674 GND.n7786 GND.n598 19.3944
R17675 GND.n7824 GND.n598 19.3944
R17676 GND.n7824 GND.n7823 19.3944
R17677 GND.n7823 GND.n7822 19.3944
R17678 GND.n7822 GND.n575 19.3944
R17679 GND.n7851 GND.n575 19.3944
R17680 GND.n7851 GND.n562 19.3944
R17681 GND.n7863 GND.n562 19.3944
R17682 GND.n7863 GND.n542 19.3944
R17683 GND.n7889 GND.n542 19.3944
R17684 GND.n7889 GND.n7888 19.3944
R17685 GND.n7888 GND.n7887 19.3944
R17686 GND.n7887 GND.n511 19.3944
R17687 GND.n7942 GND.n511 19.3944
R17688 GND.n7942 GND.n7941 19.3944
R17689 GND.n7941 GND.n7940 19.3944
R17690 GND.n7940 GND.n7939 19.3944
R17691 GND.n7939 GND.n484 19.3944
R17692 GND.n7979 GND.n484 19.3944
R17693 GND.n7979 GND.n7978 19.3944
R17694 GND.n7978 GND.n7977 19.3944
R17695 GND.n7977 GND.n7976 19.3944
R17696 GND.n7976 GND.n458 19.3944
R17697 GND.n8013 GND.n458 19.3944
R17698 GND.n8013 GND.n8012 19.3944
R17699 GND.n8012 GND.n444 19.3944
R17700 GND.n8030 GND.n444 19.3944
R17701 GND.n8030 GND.n8029 19.3944
R17702 GND.n8029 GND.n433 19.3944
R17703 GND.n8127 GND.n433 19.3944
R17704 GND.n8127 GND.n183 19.3944
R17705 GND.n8557 GND.n183 19.3944
R17706 GND.n8557 GND.n8556 19.3944
R17707 GND.n8556 GND.n8555 19.3944
R17708 GND.n8555 GND.n187 19.3944
R17709 GND.n8545 GND.n187 19.3944
R17710 GND.n8545 GND.n8544 19.3944
R17711 GND.n8544 GND.n8543 19.3944
R17712 GND.n8543 GND.n207 19.3944
R17713 GND.n8533 GND.n207 19.3944
R17714 GND.n8533 GND.n8532 19.3944
R17715 GND.n8532 GND.n8531 19.3944
R17716 GND.n8531 GND.n228 19.3944
R17717 GND.n8521 GND.n228 19.3944
R17718 GND.n8521 GND.n8520 19.3944
R17719 GND.n8520 GND.n8519 19.3944
R17720 GND.n8519 GND.n249 19.3944
R17721 GND.n8509 GND.n249 19.3944
R17722 GND.n8509 GND.n8508 19.3944
R17723 GND.n8508 GND.n8507 19.3944
R17724 GND.n8507 GND.n269 19.3944
R17725 GND.n8497 GND.n269 19.3944
R17726 GND.n8497 GND.n8496 19.3944
R17727 GND.n8496 GND.n8495 19.3944
R17728 GND.n8495 GND.n290 19.3944
R17729 GND.n8485 GND.n290 19.3944
R17730 GND.n8485 GND.n8484 19.3944
R17731 GND.n8484 GND.n8483 19.3944
R17732 GND.n8483 GND.n311 19.3944
R17733 GND.n8473 GND.n311 19.3944
R17734 GND.n8473 GND.n8472 19.3944
R17735 GND.n8472 GND.n8471 19.3944
R17736 GND.n8471 GND.n331 19.3944
R17737 GND.n8461 GND.n331 19.3944
R17738 GND.n8366 GND.n8332 19.3944
R17739 GND.n8366 GND.n8363 19.3944
R17740 GND.n8363 GND.n8360 19.3944
R17741 GND.n8360 GND.n8359 19.3944
R17742 GND.n8359 GND.n8356 19.3944
R17743 GND.n8356 GND.n8355 19.3944
R17744 GND.n8355 GND.n8352 19.3944
R17745 GND.n8352 GND.n8351 19.3944
R17746 GND.n8388 GND.n8322 19.3944
R17747 GND.n8388 GND.n8385 19.3944
R17748 GND.n8385 GND.n8382 19.3944
R17749 GND.n8382 GND.n8381 19.3944
R17750 GND.n8381 GND.n8378 19.3944
R17751 GND.n8378 GND.n8377 19.3944
R17752 GND.n8377 GND.n8374 19.3944
R17753 GND.n8374 GND.n8373 19.3944
R17754 GND.n8411 GND.n8408 19.3944
R17755 GND.n8408 GND.n8407 19.3944
R17756 GND.n8407 GND.n8404 19.3944
R17757 GND.n8404 GND.n8403 19.3944
R17758 GND.n8403 GND.n8400 19.3944
R17759 GND.n8400 GND.n8399 19.3944
R17760 GND.n8399 GND.n8396 19.3944
R17761 GND.n8396 GND.n8395 19.3944
R17762 GND.n8430 GND.n8301 19.3944
R17763 GND.n8430 GND.n8427 19.3944
R17764 GND.n8427 GND.n8426 19.3944
R17765 GND.n8426 GND.n8423 19.3944
R17766 GND.n8423 GND.n8422 19.3944
R17767 GND.n8422 GND.n8419 19.3944
R17768 GND.n8419 GND.n8418 19.3944
R17769 GND.n8418 GND.n8415 19.3944
R17770 GND.n8292 GND.n8291 19.3944
R17771 GND.n8444 GND.n8291 19.3944
R17772 GND.n8444 GND.n8443 19.3944
R17773 GND.n8443 GND.n8442 19.3944
R17774 GND.n8442 GND.n8439 19.3944
R17775 GND.n8439 GND.n8438 19.3944
R17776 GND.n8438 GND.n8435 19.3944
R17777 GND.n365 GND.n364 19.3944
R17778 GND.n369 GND.n364 19.3944
R17779 GND.n372 GND.n369 19.3944
R17780 GND.n374 GND.n372 19.3944
R17781 GND.n374 GND.n361 19.3944
R17782 GND.n378 GND.n361 19.3944
R17783 GND.n7735 GND.n7734 19.3944
R17784 GND.n7734 GND.n635 19.3944
R17785 GND.n7766 GND.n635 19.3944
R17786 GND.n7766 GND.n633 19.3944
R17787 GND.n7772 GND.n633 19.3944
R17788 GND.n7772 GND.n7771 19.3944
R17789 GND.n7771 GND.n607 19.3944
R17790 GND.n7803 GND.n607 19.3944
R17791 GND.n7803 GND.n605 19.3944
R17792 GND.n7813 GND.n605 19.3944
R17793 GND.n7813 GND.n7812 19.3944
R17794 GND.n7812 GND.n7811 19.3944
R17795 GND.n7811 GND.n580 19.3944
R17796 GND.n7839 GND.n580 19.3944
R17797 GND.n7839 GND.n578 19.3944
R17798 GND.n7844 GND.n578 19.3944
R17799 GND.n7844 GND.n555 19.3944
R17800 GND.n7871 GND.n555 19.3944
R17801 GND.n7872 GND.n7871 19.3944
R17802 GND.n7874 GND.n7872 19.3944
R17803 GND.n7874 GND.n553 19.3944
R17804 GND.n7880 GND.n553 19.3944
R17805 GND.n7880 GND.n7879 19.3944
R17806 GND.n7879 GND.n493 19.3944
R17807 GND.n7956 GND.n493 19.3944
R17808 GND.n7956 GND.n491 19.3944
R17809 GND.n7962 GND.n491 19.3944
R17810 GND.n7962 GND.n7961 19.3944
R17811 GND.n7961 GND.n466 19.3944
R17812 GND.n7993 GND.n466 19.3944
R17813 GND.n7993 GND.n464 19.3944
R17814 GND.n8004 GND.n464 19.3944
R17815 GND.n8004 GND.n8003 19.3944
R17816 GND.n8003 GND.n8002 19.3944
R17817 GND.n8002 GND.n8001 19.3944
R17818 GND.n8001 GND.n154 19.3944
R17819 GND.n8568 GND.n154 19.3944
R17820 GND.n8568 GND.n155 19.3944
R17821 GND.n427 GND.n155 19.3944
R17822 GND.n8134 GND.n427 19.3944
R17823 GND.n8134 GND.n425 19.3944
R17824 GND.n8138 GND.n425 19.3944
R17825 GND.n8138 GND.n423 19.3944
R17826 GND.n8149 GND.n423 19.3944
R17827 GND.n8149 GND.n421 19.3944
R17828 GND.n8153 GND.n421 19.3944
R17829 GND.n8153 GND.n419 19.3944
R17830 GND.n8164 GND.n419 19.3944
R17831 GND.n8164 GND.n417 19.3944
R17832 GND.n8168 GND.n417 19.3944
R17833 GND.n8168 GND.n415 19.3944
R17834 GND.n8179 GND.n415 19.3944
R17835 GND.n8179 GND.n413 19.3944
R17836 GND.n8183 GND.n413 19.3944
R17837 GND.n8183 GND.n410 19.3944
R17838 GND.n8194 GND.n410 19.3944
R17839 GND.n8194 GND.n408 19.3944
R17840 GND.n8198 GND.n408 19.3944
R17841 GND.n8198 GND.n406 19.3944
R17842 GND.n8209 GND.n406 19.3944
R17843 GND.n8209 GND.n404 19.3944
R17844 GND.n8213 GND.n404 19.3944
R17845 GND.n8213 GND.n402 19.3944
R17846 GND.n8224 GND.n402 19.3944
R17847 GND.n8224 GND.n400 19.3944
R17848 GND.n8229 GND.n400 19.3944
R17849 GND.n8229 GND.n394 19.3944
R17850 GND.n8244 GND.n394 19.3944
R17851 GND.n8244 GND.n8243 19.3944
R17852 GND.n8243 GND.n8242 19.3944
R17853 GND.n8242 GND.n351 19.3944
R17854 GND.n8454 GND.n351 19.3944
R17855 GND.n8454 GND.n8453 19.3944
R17856 GND.n6111 GND.n1564 19.3944
R17857 GND.n6115 GND.n1564 19.3944
R17858 GND.n6115 GND.n1551 19.3944
R17859 GND.n6127 GND.n1551 19.3944
R17860 GND.n6127 GND.n1549 19.3944
R17861 GND.n6140 GND.n1549 19.3944
R17862 GND.n6140 GND.n6139 19.3944
R17863 GND.n6139 GND.n6138 19.3944
R17864 GND.n6138 GND.n6137 19.3944
R17865 GND.n6137 GND.n6135 19.3944
R17866 GND.n6135 GND.n1491 19.3944
R17867 GND.n6331 GND.n1491 19.3944
R17868 GND.n6331 GND.n1489 19.3944
R17869 GND.n6335 GND.n1489 19.3944
R17870 GND.n6335 GND.n1475 19.3944
R17871 GND.n6347 GND.n1475 19.3944
R17872 GND.n6347 GND.n1473 19.3944
R17873 GND.n6351 GND.n1473 19.3944
R17874 GND.n6351 GND.n1459 19.3944
R17875 GND.n6363 GND.n1459 19.3944
R17876 GND.n6363 GND.n1457 19.3944
R17877 GND.n6367 GND.n1457 19.3944
R17878 GND.n6367 GND.n1443 19.3944
R17879 GND.n6378 GND.n1443 19.3944
R17880 GND.n6378 GND.n1441 19.3944
R17881 GND.n6382 GND.n1441 19.3944
R17882 GND.n6382 GND.n1426 19.3944
R17883 GND.n6396 GND.n1426 19.3944
R17884 GND.n6396 GND.n1424 19.3944
R17885 GND.n6402 GND.n1424 19.3944
R17886 GND.n6402 GND.n6401 19.3944
R17887 GND.n6401 GND.n1310 19.3944
R17888 GND.n6570 GND.n1310 19.3944
R17889 GND.n6570 GND.n1308 19.3944
R17890 GND.n6574 GND.n1308 19.3944
R17891 GND.n6574 GND.n1294 19.3944
R17892 GND.n6586 GND.n1294 19.3944
R17893 GND.n6586 GND.n1292 19.3944
R17894 GND.n6590 GND.n1292 19.3944
R17895 GND.n6590 GND.n1278 19.3944
R17896 GND.n6602 GND.n1278 19.3944
R17897 GND.n6602 GND.n1276 19.3944
R17898 GND.n6606 GND.n1276 19.3944
R17899 GND.n6606 GND.n1262 19.3944
R17900 GND.n6617 GND.n1262 19.3944
R17901 GND.n6617 GND.n1260 19.3944
R17902 GND.n6621 GND.n1260 19.3944
R17903 GND.n6621 GND.n1246 19.3944
R17904 GND.n6633 GND.n1246 19.3944
R17905 GND.n6633 GND.n1244 19.3944
R17906 GND.n6637 GND.n1244 19.3944
R17907 GND.n6637 GND.n1230 19.3944
R17908 GND.n6649 GND.n1230 19.3944
R17909 GND.n6649 GND.n1228 19.3944
R17910 GND.n6662 GND.n1228 19.3944
R17911 GND.n6662 GND.n6661 19.3944
R17912 GND.n6661 GND.n6660 19.3944
R17913 GND.n6660 GND.n6659 19.3944
R17914 GND.n6659 GND.n6657 19.3944
R17915 GND.n6657 GND.n1156 19.3944
R17916 GND.n6828 GND.n1156 19.3944
R17917 GND.n6828 GND.n1154 19.3944
R17918 GND.n6832 GND.n1154 19.3944
R17919 GND.n6832 GND.n1140 19.3944
R17920 GND.n6844 GND.n1140 19.3944
R17921 GND.n6844 GND.n1138 19.3944
R17922 GND.n6848 GND.n1138 19.3944
R17923 GND.n6848 GND.n1124 19.3944
R17924 GND.n6860 GND.n1124 19.3944
R17925 GND.n6860 GND.n1122 19.3944
R17926 GND.n6864 GND.n1122 19.3944
R17927 GND.n6864 GND.n1108 19.3944
R17928 GND.n6875 GND.n1108 19.3944
R17929 GND.n6875 GND.n1106 19.3944
R17930 GND.n6884 GND.n1106 19.3944
R17931 GND.n6884 GND.n6883 19.3944
R17932 GND.n6883 GND.n6882 19.3944
R17933 GND.n6882 GND.n1060 19.3944
R17934 GND.n6977 GND.n1060 19.3944
R17935 GND.n6977 GND.n6976 19.3944
R17936 GND.n6976 GND.n6975 19.3944
R17937 GND.n6975 GND.n6974 19.3944
R17938 GND.n6974 GND.n1065 19.3944
R17939 GND.n5596 GND.n5592 19.3944
R17940 GND.n5597 GND.n5596 19.3944
R17941 GND.n5600 GND.n5597 19.3944
R17942 GND.n5600 GND.n5590 19.3944
R17943 GND.n5621 GND.n5590 19.3944
R17944 GND.n5621 GND.n5620 19.3944
R17945 GND.n5620 GND.n5619 19.3944
R17946 GND.n5619 GND.n5617 19.3944
R17947 GND.n5617 GND.n5616 19.3944
R17948 GND.n5616 GND.n5614 19.3944
R17949 GND.n5614 GND.n5613 19.3944
R17950 GND.n5613 GND.n1513 19.3944
R17951 GND.n6310 GND.n1513 19.3944
R17952 GND.n6310 GND.n6309 19.3944
R17953 GND.n6309 GND.n6308 19.3944
R17954 GND.n6308 GND.n1517 19.3944
R17955 GND.n6213 GND.n1517 19.3944
R17956 GND.n6213 GND.n6210 19.3944
R17957 GND.n6218 GND.n6210 19.3944
R17958 GND.n6219 GND.n6218 19.3944
R17959 GND.n6221 GND.n6219 19.3944
R17960 GND.n6221 GND.n6208 19.3944
R17961 GND.n6226 GND.n6208 19.3944
R17962 GND.n6227 GND.n6226 19.3944
R17963 GND.n6229 GND.n6227 19.3944
R17964 GND.n6229 GND.n6206 19.3944
R17965 GND.n6235 GND.n6206 19.3944
R17966 GND.n6235 GND.n6234 19.3944
R17967 GND.n6234 GND.n1420 19.3944
R17968 GND.n6406 GND.n1420 19.3944
R17969 GND.n6406 GND.n1418 19.3944
R17970 GND.n6411 GND.n1418 19.3944
R17971 GND.n6412 GND.n6411 19.3944
R17972 GND.n6414 GND.n6412 19.3944
R17973 GND.n6414 GND.n1416 19.3944
R17974 GND.n6419 GND.n1416 19.3944
R17975 GND.n6420 GND.n6419 19.3944
R17976 GND.n6422 GND.n6420 19.3944
R17977 GND.n6422 GND.n1414 19.3944
R17978 GND.n6427 GND.n1414 19.3944
R17979 GND.n6428 GND.n6427 19.3944
R17980 GND.n6430 GND.n6428 19.3944
R17981 GND.n6430 GND.n1412 19.3944
R17982 GND.n6435 GND.n1412 19.3944
R17983 GND.n6436 GND.n6435 19.3944
R17984 GND.n6438 GND.n6436 19.3944
R17985 GND.n6438 GND.n1410 19.3944
R17986 GND.n6443 GND.n1410 19.3944
R17987 GND.n6444 GND.n6443 19.3944
R17988 GND.n6447 GND.n6444 19.3944
R17989 GND.n6447 GND.n1408 19.3944
R17990 GND.n6473 GND.n1408 19.3944
R17991 GND.n6473 GND.n6472 19.3944
R17992 GND.n6472 GND.n6471 19.3944
R17993 GND.n6471 GND.n6469 19.3944
R17994 GND.n6469 GND.n6468 19.3944
R17995 GND.n6468 GND.n6466 19.3944
R17996 GND.n6466 GND.n6465 19.3944
R17997 GND.n6465 GND.n6463 19.3944
R17998 GND.n6463 GND.n6462 19.3944
R17999 GND.n6462 GND.n1178 19.3944
R18000 GND.n6807 GND.n1178 19.3944
R18001 GND.n6807 GND.n6806 19.3944
R18002 GND.n6806 GND.n6805 19.3944
R18003 GND.n6805 GND.n1182 19.3944
R18004 GND.n6793 GND.n1182 19.3944
R18005 GND.n6793 GND.n6792 19.3944
R18006 GND.n6792 GND.n6791 19.3944
R18007 GND.n6791 GND.n1195 19.3944
R18008 GND.n6725 GND.n1195 19.3944
R18009 GND.n6726 GND.n6725 19.3944
R18010 GND.n6728 GND.n6726 19.3944
R18011 GND.n6728 GND.n6720 19.3944
R18012 GND.n6739 GND.n6720 19.3944
R18013 GND.n6739 GND.n6738 19.3944
R18014 GND.n6738 GND.n6737 19.3944
R18015 GND.n6737 GND.n1085 19.3944
R18016 GND.n6907 GND.n1085 19.3944
R18017 GND.n6908 GND.n6907 19.3944
R18018 GND.n6908 GND.n1083 19.3944
R18019 GND.n6912 GND.n1083 19.3944
R18020 GND.n6914 GND.n6912 19.3944
R18021 GND.n6915 GND.n6914 19.3944
R18022 GND.n6097 GND.n6096 19.3944
R18023 GND.n6096 GND.n6095 19.3944
R18024 GND.n6095 GND.n6094 19.3944
R18025 GND.n6094 GND.n6092 19.3944
R18026 GND.n6092 GND.n6089 19.3944
R18027 GND.n6089 GND.n6088 19.3944
R18028 GND.n6086 GND.n6085 19.3944
R18029 GND.n6083 GND.n6082 19.3944
R18030 GND.n6080 GND.n6079 19.3944
R18031 GND.n6077 GND.n6076 19.3944
R18032 GND.n6072 GND.n6071 19.3944
R18033 GND.n6071 GND.n6069 19.3944
R18034 GND.n6069 GND.n6067 19.3944
R18035 GND.n6965 GND.n1068 19.3944
R18036 GND.n6965 GND.n1067 19.3944
R18037 GND.n6970 GND.n1067 19.3944
R18038 GND.n6918 GND.n1078 19.3944
R18039 GND.n6924 GND.n1078 19.3944
R18040 GND.n6924 GND.n1076 19.3944
R18041 GND.n6929 GND.n1076 19.3944
R18042 GND.n6929 GND.n1074 19.3944
R18043 GND.n6935 GND.n1074 19.3944
R18044 GND.n6939 GND.n6937 19.3944
R18045 GND.n6945 GND.n1072 19.3944
R18046 GND.n6949 GND.n6947 19.3944
R18047 GND.n6954 GND.n1070 19.3944
R18048 GND.n699 GND.n698 19.3944
R18049 GND.n702 GND.n664 19.3944
R18050 GND.n669 GND.n664 19.3944
R18051 GND.n7756 GND.n645 19.3944
R18052 GND.n7756 GND.n643 19.3944
R18053 GND.n7762 GND.n643 19.3944
R18054 GND.n7762 GND.n7761 19.3944
R18055 GND.n7761 GND.n617 19.3944
R18056 GND.n7793 GND.n617 19.3944
R18057 GND.n7793 GND.n615 19.3944
R18058 GND.n7799 GND.n615 19.3944
R18059 GND.n7799 GND.n7798 19.3944
R18060 GND.n7798 GND.n590 19.3944
R18061 GND.n7828 GND.n590 19.3944
R18062 GND.n7828 GND.n588 19.3944
R18063 GND.n7832 GND.n588 19.3944
R18064 GND.n7832 GND.n568 19.3944
R18065 GND.n7855 GND.n568 19.3944
R18066 GND.n7855 GND.n566 19.3944
R18067 GND.n7859 GND.n566 19.3944
R18068 GND.n7859 GND.n534 19.3944
R18069 GND.n7893 GND.n534 19.3944
R18070 GND.n7893 GND.n532 19.3944
R18071 GND.n7897 GND.n532 19.3944
R18072 GND.n7897 GND.n503 19.3944
R18073 GND.n7946 GND.n503 19.3944
R18074 GND.n7946 GND.n501 19.3944
R18075 GND.n7952 GND.n501 19.3944
R18076 GND.n7952 GND.n7951 19.3944
R18077 GND.n7951 GND.n476 19.3944
R18078 GND.n7983 GND.n476 19.3944
R18079 GND.n7983 GND.n474 19.3944
R18080 GND.n7989 GND.n474 19.3944
R18081 GND.n7989 GND.n7988 19.3944
R18082 GND.n7988 GND.n7987 19.3944
R18083 GND.n454 GND.n171 19.3944
R18084 GND.n8017 GND.n171 19.3944
R18085 GND.n8564 GND.n164 19.3944
R18086 GND.n8123 GND.n165 19.3944
R18087 GND.n8561 GND.n173 19.3944
R18088 GND.n8561 GND.n174 19.3944
R18089 GND.n8551 GND.n174 19.3944
R18090 GND.n8551 GND.n8550 19.3944
R18091 GND.n8550 GND.n8549 19.3944
R18092 GND.n8549 GND.n197 19.3944
R18093 GND.n8539 GND.n197 19.3944
R18094 GND.n8539 GND.n8538 19.3944
R18095 GND.n8538 GND.n8537 19.3944
R18096 GND.n8537 GND.n218 19.3944
R18097 GND.n8527 GND.n218 19.3944
R18098 GND.n8527 GND.n8526 19.3944
R18099 GND.n8526 GND.n8525 19.3944
R18100 GND.n8525 GND.n239 19.3944
R18101 GND.n8515 GND.n239 19.3944
R18102 GND.n8515 GND.n8514 19.3944
R18103 GND.n8514 GND.n8513 19.3944
R18104 GND.n8513 GND.n259 19.3944
R18105 GND.n8503 GND.n259 19.3944
R18106 GND.n8503 GND.n8502 19.3944
R18107 GND.n8502 GND.n8501 19.3944
R18108 GND.n8501 GND.n280 19.3944
R18109 GND.n8491 GND.n280 19.3944
R18110 GND.n8491 GND.n8490 19.3944
R18111 GND.n8490 GND.n8489 19.3944
R18112 GND.n8489 GND.n301 19.3944
R18113 GND.n8479 GND.n301 19.3944
R18114 GND.n8479 GND.n8478 19.3944
R18115 GND.n8478 GND.n8477 19.3944
R18116 GND.n8477 GND.n321 19.3944
R18117 GND.n8467 GND.n321 19.3944
R18118 GND.n8467 GND.n8466 19.3944
R18119 GND.n8466 GND.n8465 19.3944
R18120 GND.n4123 GND.n4122 19.3944
R18121 GND.n4122 GND.n4094 19.3944
R18122 GND.n4118 GND.n4094 19.3944
R18123 GND.n4118 GND.n4117 19.3944
R18124 GND.n4117 GND.n4116 19.3944
R18125 GND.n4116 GND.n4100 19.3944
R18126 GND.n4112 GND.n4100 19.3944
R18127 GND.n4112 GND.n4111 19.3944
R18128 GND.n4111 GND.n4110 19.3944
R18129 GND.n4110 GND.n4107 19.3944
R18130 GND.n4107 GND.n2061 19.3944
R18131 GND.n4435 GND.n2061 19.3944
R18132 GND.n4435 GND.n2059 19.3944
R18133 GND.n4439 GND.n2059 19.3944
R18134 GND.n4439 GND.n2057 19.3944
R18135 GND.n4443 GND.n2057 19.3944
R18136 GND.n4443 GND.n2055 19.3944
R18137 GND.n4449 GND.n2055 19.3944
R18138 GND.n4449 GND.n4448 19.3944
R18139 GND.n4448 GND.n1999 19.3944
R18140 GND.n4517 GND.n1999 19.3944
R18141 GND.n4517 GND.n1997 19.3944
R18142 GND.n4521 GND.n1997 19.3944
R18143 GND.n4521 GND.n1995 19.3944
R18144 GND.n4525 GND.n1995 19.3944
R18145 GND.n4525 GND.n1993 19.3944
R18146 GND.n4567 GND.n1993 19.3944
R18147 GND.n4567 GND.n4566 19.3944
R18148 GND.n4566 GND.n4565 19.3944
R18149 GND.n4565 GND.n4531 19.3944
R18150 GND.n4561 GND.n4531 19.3944
R18151 GND.n4561 GND.n4560 19.3944
R18152 GND.n4560 GND.n4559 19.3944
R18153 GND.n4557 GND.n4537 19.3944
R18154 GND.n4553 GND.n4552 19.3944
R18155 GND.n4550 GND.n4540 19.3944
R18156 GND.n4546 GND.n4545 19.3944
R18157 GND.n4543 GND.n1856 19.3944
R18158 GND.n1856 GND.n1854 19.3944
R18159 GND.n4709 GND.n1854 19.3944
R18160 GND.n4709 GND.n1852 19.3944
R18161 GND.n4726 GND.n1852 19.3944
R18162 GND.n4726 GND.n4725 19.3944
R18163 GND.n4725 GND.n4724 19.3944
R18164 GND.n4724 GND.n4715 19.3944
R18165 GND.n4720 GND.n4715 19.3944
R18166 GND.n4720 GND.n4719 19.3944
R18167 GND.n4719 GND.n1790 19.3944
R18168 GND.n4802 GND.n1790 19.3944
R18169 GND.n4802 GND.n1788 19.3944
R18170 GND.n4829 GND.n1788 19.3944
R18171 GND.n4829 GND.n4828 19.3944
R18172 GND.n4828 GND.n4827 19.3944
R18173 GND.n4827 GND.n4808 19.3944
R18174 GND.n4823 GND.n4808 19.3944
R18175 GND.n4823 GND.n4822 19.3944
R18176 GND.n4822 GND.n4821 19.3944
R18177 GND.n4821 GND.n4814 19.3944
R18178 GND.n4817 GND.n4814 19.3944
R18179 GND.n4817 GND.n1708 19.3944
R18180 GND.n4932 GND.n1708 19.3944
R18181 GND.n4932 GND.n1706 19.3944
R18182 GND.n5858 GND.n1706 19.3944
R18183 GND.n5858 GND.n5857 19.3944
R18184 GND.n5857 GND.n5856 19.3944
R18185 GND.n5856 GND.n4938 19.3944
R18186 GND.n5852 GND.n4938 19.3944
R18187 GND.n5852 GND.n5851 19.3944
R18188 GND.n5851 GND.n5850 19.3944
R18189 GND.n5850 GND.n4944 19.3944
R18190 GND.n5846 GND.n4944 19.3944
R18191 GND.n5846 GND.n5845 19.3944
R18192 GND.n5845 GND.n5844 19.3944
R18193 GND.n5844 GND.n4950 19.3944
R18194 GND.n5838 GND.n4950 19.3944
R18195 GND.n5838 GND.n5837 19.3944
R18196 GND.n5837 GND.n5836 19.3944
R18197 GND.n5836 GND.n4959 19.3944
R18198 GND.n5824 GND.n4959 19.3944
R18199 GND.n5824 GND.n5823 19.3944
R18200 GND.n5823 GND.n5822 19.3944
R18201 GND.n5822 GND.n4977 19.3944
R18202 GND.n5810 GND.n4977 19.3944
R18203 GND.n5810 GND.n5809 19.3944
R18204 GND.n5809 GND.n5808 19.3944
R18205 GND.n5808 GND.n4995 19.3944
R18206 GND.n5796 GND.n4995 19.3944
R18207 GND.n5796 GND.n5795 19.3944
R18208 GND.n5795 GND.n5794 19.3944
R18209 GND.n5794 GND.n5012 19.3944
R18210 GND.n5782 GND.n5012 19.3944
R18211 GND.n5782 GND.n5781 19.3944
R18212 GND.n5781 GND.n5780 19.3944
R18213 GND.n5780 GND.n5030 19.3944
R18214 GND.n5768 GND.n5030 19.3944
R18215 GND.n5768 GND.n5767 19.3944
R18216 GND.n5767 GND.n5766 19.3944
R18217 GND.n5766 GND.n5048 19.3944
R18218 GND.n5064 GND.n5048 19.3944
R18219 GND.n5753 GND.n5064 19.3944
R18220 GND.n5753 GND.n5752 19.3944
R18221 GND.n5752 GND.n5751 19.3944
R18222 GND.n5751 GND.n5070 19.3944
R18223 GND.n5739 GND.n5070 19.3944
R18224 GND.n5739 GND.n5738 19.3944
R18225 GND.n5738 GND.n5737 19.3944
R18226 GND.n5737 GND.n5087 19.3944
R18227 GND.n5725 GND.n5087 19.3944
R18228 GND.n5725 GND.n5724 19.3944
R18229 GND.n5724 GND.n5723 19.3944
R18230 GND.n5723 GND.n5105 19.3944
R18231 GND.n5711 GND.n5105 19.3944
R18232 GND.n5711 GND.n5710 19.3944
R18233 GND.n5710 GND.n5709 19.3944
R18234 GND.n5709 GND.n5123 19.3944
R18235 GND.n5139 GND.n5123 19.3944
R18236 GND.n5696 GND.n5139 19.3944
R18237 GND.n5696 GND.n5695 19.3944
R18238 GND.n5695 GND.n5694 19.3944
R18239 GND.n5694 GND.n5145 19.3944
R18240 GND.n5682 GND.n5145 19.3944
R18241 GND.n5682 GND.n5681 19.3944
R18242 GND.n5681 GND.n5680 19.3944
R18243 GND.n5680 GND.n5163 19.3944
R18244 GND.n5668 GND.n5163 19.3944
R18245 GND.n5668 GND.n5667 19.3944
R18246 GND.n5667 GND.n5666 19.3944
R18247 GND.n5666 GND.n5181 19.3944
R18248 GND.n5654 GND.n5181 19.3944
R18249 GND.n5654 GND.n1573 19.3944
R18250 GND.n6103 GND.n1573 19.3944
R18251 GND.n6103 GND.n1571 19.3944
R18252 GND.n6107 GND.n1571 19.3944
R18253 GND.n6107 GND.n1559 19.3944
R18254 GND.n6119 GND.n1559 19.3944
R18255 GND.n6119 GND.n1557 19.3944
R18256 GND.n6123 GND.n1557 19.3944
R18257 GND.n6123 GND.n1542 19.3944
R18258 GND.n6144 GND.n1542 19.3944
R18259 GND.n6144 GND.n1540 19.3944
R18260 GND.n6148 GND.n1540 19.3944
R18261 GND.n6148 GND.n1499 19.3944
R18262 GND.n6323 GND.n1499 19.3944
R18263 GND.n6323 GND.n1497 19.3944
R18264 GND.n6327 GND.n1497 19.3944
R18265 GND.n6327 GND.n1483 19.3944
R18266 GND.n6339 GND.n1483 19.3944
R18267 GND.n6339 GND.n1481 19.3944
R18268 GND.n6343 GND.n1481 19.3944
R18269 GND.n6343 GND.n1467 19.3944
R18270 GND.n6355 GND.n1467 19.3944
R18271 GND.n6355 GND.n1465 19.3944
R18272 GND.n6359 GND.n1465 19.3944
R18273 GND.n6359 GND.n1451 19.3944
R18274 GND.n6371 GND.n1451 19.3944
R18275 GND.n6371 GND.n1449 19.3944
R18276 GND.n6375 GND.n1449 19.3944
R18277 GND.n6375 GND.n1435 19.3944
R18278 GND.n6386 GND.n1435 19.3944
R18279 GND.n6386 GND.n1433 19.3944
R18280 GND.n6392 GND.n1433 19.3944
R18281 GND.n6392 GND.n6391 19.3944
R18282 GND.n6391 GND.n1317 19.3944
R18283 GND.n6562 GND.n1317 19.3944
R18284 GND.n6562 GND.n1315 19.3944
R18285 GND.n6566 GND.n1315 19.3944
R18286 GND.n6566 GND.n1302 19.3944
R18287 GND.n6578 GND.n1302 19.3944
R18288 GND.n6578 GND.n1300 19.3944
R18289 GND.n6582 GND.n1300 19.3944
R18290 GND.n6582 GND.n1286 19.3944
R18291 GND.n6594 GND.n1286 19.3944
R18292 GND.n6594 GND.n1284 19.3944
R18293 GND.n6598 GND.n1284 19.3944
R18294 GND.n6598 GND.n1270 19.3944
R18295 GND.n6610 GND.n1270 19.3944
R18296 GND.n6610 GND.n1268 19.3944
R18297 GND.n6614 GND.n1268 19.3944
R18298 GND.n6614 GND.n1254 19.3944
R18299 GND.n6625 GND.n1254 19.3944
R18300 GND.n6625 GND.n1252 19.3944
R18301 GND.n6629 GND.n1252 19.3944
R18302 GND.n6629 GND.n1238 19.3944
R18303 GND.n6641 GND.n1238 19.3944
R18304 GND.n6641 GND.n1236 19.3944
R18305 GND.n6645 GND.n1236 19.3944
R18306 GND.n6645 GND.n1221 19.3944
R18307 GND.n6666 GND.n1221 19.3944
R18308 GND.n6666 GND.n1219 19.3944
R18309 GND.n6670 GND.n1219 19.3944
R18310 GND.n6670 GND.n1164 19.3944
R18311 GND.n6820 GND.n1164 19.3944
R18312 GND.n6820 GND.n1162 19.3944
R18313 GND.n6824 GND.n1162 19.3944
R18314 GND.n6824 GND.n1148 19.3944
R18315 GND.n6836 GND.n1148 19.3944
R18316 GND.n6836 GND.n1146 19.3944
R18317 GND.n6840 GND.n1146 19.3944
R18318 GND.n6840 GND.n1132 19.3944
R18319 GND.n6852 GND.n1132 19.3944
R18320 GND.n6852 GND.n1130 19.3944
R18321 GND.n6856 GND.n1130 19.3944
R18322 GND.n6856 GND.n1116 19.3944
R18323 GND.n6868 GND.n1116 19.3944
R18324 GND.n6868 GND.n1114 19.3944
R18325 GND.n6872 GND.n1114 19.3944
R18326 GND.n6872 GND.n1099 19.3944
R18327 GND.n6888 GND.n1099 19.3944
R18328 GND.n6888 GND.n1097 19.3944
R18329 GND.n6892 GND.n1097 19.3944
R18330 GND.n6892 GND.n1053 19.3944
R18331 GND.n6981 GND.n1053 19.3944
R18332 GND.n6981 GND.n1051 19.3944
R18333 GND.n6990 GND.n1051 19.3944
R18334 GND.n6990 GND.n6989 19.3944
R18335 GND.n6989 GND.n6988 19.3944
R18336 GND.n6988 GND.n1029 19.3944
R18337 GND.n7021 GND.n1029 19.3944
R18338 GND.n7021 GND.n1027 19.3944
R18339 GND.n7036 GND.n1027 19.3944
R18340 GND.n7036 GND.n7035 19.3944
R18341 GND.n7035 GND.n7034 19.3944
R18342 GND.n7034 GND.n7027 19.3944
R18343 GND.n7030 GND.n7027 19.3944
R18344 GND.n7030 GND.n995 19.3944
R18345 GND.n7079 GND.n995 19.3944
R18346 GND.n7079 GND.n993 19.3944
R18347 GND.n7085 GND.n993 19.3944
R18348 GND.n7085 GND.n7084 19.3944
R18349 GND.n7084 GND.n970 19.3944
R18350 GND.n7114 GND.n970 19.3944
R18351 GND.n7114 GND.n968 19.3944
R18352 GND.n7123 GND.n968 19.3944
R18353 GND.n7123 GND.n7122 19.3944
R18354 GND.n7122 GND.n7121 19.3944
R18355 GND.n7121 GND.n945 19.3944
R18356 GND.n7153 GND.n945 19.3944
R18357 GND.n7153 GND.n943 19.3944
R18358 GND.n7168 GND.n943 19.3944
R18359 GND.n7168 GND.n7167 19.3944
R18360 GND.n7167 GND.n7166 19.3944
R18361 GND.n7166 GND.n7159 19.3944
R18362 GND.n7162 GND.n7159 19.3944
R18363 GND.n7162 GND.n913 19.3944
R18364 GND.n7213 GND.n913 19.3944
R18365 GND.n7213 GND.n911 19.3944
R18366 GND.n7237 GND.n911 19.3944
R18367 GND.n7237 GND.n7236 19.3944
R18368 GND.n7236 GND.n7235 19.3944
R18369 GND.n7235 GND.n7219 19.3944
R18370 GND.n7231 GND.n7219 19.3944
R18371 GND.n7231 GND.n7230 19.3944
R18372 GND.n7230 GND.n7229 19.3944
R18373 GND.n7229 GND.n7226 19.3944
R18374 GND.n7226 GND.n869 19.3944
R18375 GND.n7293 GND.n869 19.3944
R18376 GND.n7293 GND.n867 19.3944
R18377 GND.n7299 GND.n867 19.3944
R18378 GND.n7299 GND.n7298 19.3944
R18379 GND.n7298 GND.n844 19.3944
R18380 GND.n7329 GND.n844 19.3944
R18381 GND.n7329 GND.n842 19.3944
R18382 GND.n7333 GND.n842 19.3944
R18383 GND.n7333 GND.n828 19.3944
R18384 GND.n7352 GND.n828 19.3944
R18385 GND.n7352 GND.n826 19.3944
R18386 GND.n7358 GND.n826 19.3944
R18387 GND.n7358 GND.n7357 19.3944
R18388 GND.n7357 GND.n804 19.3944
R18389 GND.n7444 GND.n804 19.3944
R18390 GND.n7444 GND.n802 19.3944
R18391 GND.n7532 GND.n802 19.3944
R18392 GND.n7532 GND.n7531 19.3944
R18393 GND.n7531 GND.n7530 19.3944
R18394 GND.n7530 GND.n7450 19.3944
R18395 GND.n7524 GND.n7450 19.3944
R18396 GND.n7524 GND.n7523 19.3944
R18397 GND.n7523 GND.n7522 19.3944
R18398 GND.n7522 GND.n7458 19.3944
R18399 GND.n7518 GND.n7458 19.3944
R18400 GND.n7518 GND.n7517 19.3944
R18401 GND.n7517 GND.n7516 19.3944
R18402 GND.n7516 GND.n7464 19.3944
R18403 GND.n7512 GND.n7464 19.3944
R18404 GND.n7512 GND.n7511 19.3944
R18405 GND.n7511 GND.n7510 19.3944
R18406 GND.n7510 GND.n7470 19.3944
R18407 GND.n7506 GND.n7470 19.3944
R18408 GND.n7506 GND.n7505 19.3944
R18409 GND.n7505 GND.n7504 19.3944
R18410 GND.n7504 GND.n7476 19.3944
R18411 GND.n7500 GND.n7476 19.3944
R18412 GND.n7500 GND.n7499 19.3944
R18413 GND.n7499 GND.n7498 19.3944
R18414 GND.n7498 GND.n7482 19.3944
R18415 GND.n7494 GND.n7482 19.3944
R18416 GND.n7494 GND.n7493 19.3944
R18417 GND.n7493 GND.n7492 19.3944
R18418 GND.n7492 GND.n7489 19.3944
R18419 GND.n7489 GND.n524 19.3944
R18420 GND.n7902 GND.n524 19.3944
R18421 GND.n7902 GND.n522 19.3944
R18422 GND.n7906 GND.n522 19.3944
R18423 GND.n7906 GND.n520 19.3944
R18424 GND.n7910 GND.n520 19.3944
R18425 GND.n7910 GND.n518 19.3944
R18426 GND.n7934 GND.n518 19.3944
R18427 GND.n7934 GND.n7933 19.3944
R18428 GND.n7933 GND.n7932 19.3944
R18429 GND.n7932 GND.n7916 19.3944
R18430 GND.n7928 GND.n7916 19.3944
R18431 GND.n7928 GND.n7927 19.3944
R18432 GND.n7925 GND.n7922 19.3944
R18433 GND.n7920 GND.n440 19.3944
R18434 GND.n8037 GND.n8036 19.3944
R18435 GND.n8120 GND.n8119 19.3944
R18436 GND.n8117 GND.n8039 19.3944
R18437 GND.n8113 GND.n8039 19.3944
R18438 GND.n8113 GND.n8112 19.3944
R18439 GND.n8112 GND.n8111 19.3944
R18440 GND.n8111 GND.n8045 19.3944
R18441 GND.n8107 GND.n8045 19.3944
R18442 GND.n8107 GND.n8106 19.3944
R18443 GND.n8106 GND.n8105 19.3944
R18444 GND.n8105 GND.n8051 19.3944
R18445 GND.n8101 GND.n8051 19.3944
R18446 GND.n8101 GND.n8100 19.3944
R18447 GND.n8100 GND.n8099 19.3944
R18448 GND.n8099 GND.n8057 19.3944
R18449 GND.n8095 GND.n8057 19.3944
R18450 GND.n8095 GND.n8094 19.3944
R18451 GND.n8094 GND.n8093 19.3944
R18452 GND.n8093 GND.n8063 19.3944
R18453 GND.n8089 GND.n8063 19.3944
R18454 GND.n8089 GND.n8088 19.3944
R18455 GND.n8088 GND.n8087 19.3944
R18456 GND.n8087 GND.n8069 19.3944
R18457 GND.n8083 GND.n8069 19.3944
R18458 GND.n8083 GND.n8082 19.3944
R18459 GND.n8082 GND.n8081 19.3944
R18460 GND.n8081 GND.n8078 19.3944
R18461 GND.n8078 GND.n8077 19.3944
R18462 GND.n8077 GND.n391 19.3944
R18463 GND.n8250 GND.n391 19.3944
R18464 GND.n8250 GND.n389 19.3944
R18465 GND.n8255 GND.n389 19.3944
R18466 GND.n8255 GND.n387 19.3944
R18467 GND.n8259 GND.n387 19.3944
R18468 GND.n8260 GND.n8259 19.3944
R18469 GND.n4310 GND.n4158 19.3944
R18470 GND.n4310 GND.n4309 19.3944
R18471 GND.n4309 GND.n4308 19.3944
R18472 GND.n4308 GND.n4306 19.3944
R18473 GND.n4306 GND.n4303 19.3944
R18474 GND.n4303 GND.n4302 19.3944
R18475 GND.n4302 GND.n4299 19.3944
R18476 GND.n4297 GND.n4295 19.3944
R18477 GND.n4295 GND.n4292 19.3944
R18478 GND.n4292 GND.n4291 19.3944
R18479 GND.n4291 GND.n4288 19.3944
R18480 GND.n4288 GND.n4287 19.3944
R18481 GND.n4287 GND.n4284 19.3944
R18482 GND.n4284 GND.n4283 19.3944
R18483 GND.n4283 GND.n4280 19.3944
R18484 GND.n4278 GND.n4275 19.3944
R18485 GND.n4275 GND.n4274 19.3944
R18486 GND.n4274 GND.n4271 19.3944
R18487 GND.n4271 GND.n4270 19.3944
R18488 GND.n4270 GND.n4267 19.3944
R18489 GND.n4267 GND.n4266 19.3944
R18490 GND.n4266 GND.n4263 19.3944
R18491 GND.n4263 GND.n4262 19.3944
R18492 GND.n4258 GND.n4255 19.3944
R18493 GND.n4255 GND.n4254 19.3944
R18494 GND.n4254 GND.n4251 19.3944
R18495 GND.n4251 GND.n4250 19.3944
R18496 GND.n4250 GND.n4247 19.3944
R18497 GND.n4247 GND.n4246 19.3944
R18498 GND.n4246 GND.n4243 19.3944
R18499 GND.n4243 GND.n4242 19.3944
R18500 GND.n4238 GND.n4235 19.3944
R18501 GND.n4235 GND.n4234 19.3944
R18502 GND.n4234 GND.n4231 19.3944
R18503 GND.n4231 GND.n4230 19.3944
R18504 GND.n4230 GND.n4227 19.3944
R18505 GND.n4227 GND.n4226 19.3944
R18506 GND.n4226 GND.n4223 19.3944
R18507 GND.n4223 GND.n4222 19.3944
R18508 GND.n4347 GND.n2127 19.3944
R18509 GND.n4353 GND.n2127 19.3944
R18510 GND.n4353 GND.n4352 19.3944
R18511 GND.n4352 GND.n2100 19.3944
R18512 GND.n4383 GND.n2100 19.3944
R18513 GND.n4383 GND.n2098 19.3944
R18514 GND.n4389 GND.n2098 19.3944
R18515 GND.n4389 GND.n4388 19.3944
R18516 GND.n4388 GND.n2071 19.3944
R18517 GND.n4426 GND.n2071 19.3944
R18518 GND.n4426 GND.n2069 19.3944
R18519 GND.n4430 GND.n2069 19.3944
R18520 GND.n4430 GND.n2037 19.3944
R18521 GND.n4465 GND.n2037 19.3944
R18522 GND.n4465 GND.n2035 19.3944
R18523 GND.n4471 GND.n2035 19.3944
R18524 GND.n4471 GND.n4470 19.3944
R18525 GND.n4470 GND.n2009 19.3944
R18526 GND.n4508 GND.n2009 19.3944
R18527 GND.n4508 GND.n2007 19.3944
R18528 GND.n4512 GND.n2007 19.3944
R18529 GND.n4512 GND.n1975 19.3944
R18530 GND.n4583 GND.n1975 19.3944
R18531 GND.n4583 GND.n1973 19.3944
R18532 GND.n4589 GND.n1973 19.3944
R18533 GND.n4589 GND.n4588 19.3944
R18534 GND.n4588 GND.n1945 19.3944
R18535 GND.n4615 GND.n1945 19.3944
R18536 GND.n4615 GND.n1943 19.3944
R18537 GND.n4619 GND.n1943 19.3944
R18538 GND.n4619 GND.n1879 19.3944
R18539 GND.n4687 GND.n1879 19.3944
R18540 GND.n1878 GND.n1877 19.3944
R18541 GND.n1927 GND.n1877 19.3944
R18542 GND.n4639 GND.n4638 19.3944
R18543 GND.n4655 GND.n4654 19.3944
R18544 GND.n4692 GND.n1870 19.3944
R18545 GND.n4692 GND.n4691 19.3944
R18546 GND.n4691 GND.n1834 19.3944
R18547 GND.n4742 GND.n1834 19.3944
R18548 GND.n4742 GND.n1832 19.3944
R18549 GND.n4748 GND.n1832 19.3944
R18550 GND.n4748 GND.n4747 19.3944
R18551 GND.n4747 GND.n1807 19.3944
R18552 GND.n4780 GND.n1807 19.3944
R18553 GND.n4780 GND.n1805 19.3944
R18554 GND.n4786 GND.n1805 19.3944
R18555 GND.n4786 GND.n4785 19.3944
R18556 GND.n4785 GND.n1773 19.3944
R18557 GND.n4848 GND.n1773 19.3944
R18558 GND.n4848 GND.n1771 19.3944
R18559 GND.n4854 GND.n1771 19.3944
R18560 GND.n4854 GND.n4853 19.3944
R18561 GND.n4853 GND.n1746 19.3944
R18562 GND.n4885 GND.n1746 19.3944
R18563 GND.n4885 GND.n1744 19.3944
R18564 GND.n4891 GND.n1744 19.3944
R18565 GND.n4891 GND.n4890 19.3944
R18566 GND.n4890 GND.n1716 19.3944
R18567 GND.n4923 GND.n1716 19.3944
R18568 GND.n4923 GND.n1714 19.3944
R18569 GND.n4927 GND.n1714 19.3944
R18570 GND.n4927 GND.n1689 19.3944
R18571 GND.n5883 GND.n1689 19.3944
R18572 GND.n5883 GND.n1687 19.3944
R18573 GND.n5888 GND.n1687 19.3944
R18574 GND.n5888 GND.n1674 19.3944
R18575 GND.n5901 GND.n1674 19.3944
R18576 GND.n5902 GND.n5901 19.3944
R18577 GND.n3940 GND.n2247 19.3944
R18578 GND.n3940 GND.n2245 19.3944
R18579 GND.n3944 GND.n2245 19.3944
R18580 GND.n3944 GND.n2241 19.3944
R18581 GND.n3950 GND.n2241 19.3944
R18582 GND.n3950 GND.n2239 19.3944
R18583 GND.n3954 GND.n2239 19.3944
R18584 GND.n3954 GND.n2235 19.3944
R18585 GND.n3960 GND.n2235 19.3944
R18586 GND.n3960 GND.n2233 19.3944
R18587 GND.n3964 GND.n2233 19.3944
R18588 GND.n3964 GND.n2229 19.3944
R18589 GND.n3970 GND.n2229 19.3944
R18590 GND.n3970 GND.n2227 19.3944
R18591 GND.n3974 GND.n2227 19.3944
R18592 GND.n3974 GND.n2223 19.3944
R18593 GND.n3980 GND.n2223 19.3944
R18594 GND.n3980 GND.n2221 19.3944
R18595 GND.n3984 GND.n2221 19.3944
R18596 GND.n3984 GND.n2217 19.3944
R18597 GND.n3990 GND.n2217 19.3944
R18598 GND.n3990 GND.n2215 19.3944
R18599 GND.n3994 GND.n2215 19.3944
R18600 GND.n3994 GND.n2211 19.3944
R18601 GND.n4000 GND.n2211 19.3944
R18602 GND.n4000 GND.n2209 19.3944
R18603 GND.n4004 GND.n2209 19.3944
R18604 GND.n4004 GND.n2205 19.3944
R18605 GND.n4010 GND.n2205 19.3944
R18606 GND.n4010 GND.n2203 19.3944
R18607 GND.n4014 GND.n2203 19.3944
R18608 GND.n4014 GND.n2199 19.3944
R18609 GND.n4020 GND.n2199 19.3944
R18610 GND.n4020 GND.n2197 19.3944
R18611 GND.n4024 GND.n2197 19.3944
R18612 GND.n4024 GND.n2193 19.3944
R18613 GND.n4030 GND.n2193 19.3944
R18614 GND.n4030 GND.n2191 19.3944
R18615 GND.n4034 GND.n2191 19.3944
R18616 GND.n4034 GND.n2187 19.3944
R18617 GND.n4040 GND.n2187 19.3944
R18618 GND.n4040 GND.n2185 19.3944
R18619 GND.n4044 GND.n2185 19.3944
R18620 GND.n4044 GND.n2181 19.3944
R18621 GND.n4050 GND.n2181 19.3944
R18622 GND.n4050 GND.n2179 19.3944
R18623 GND.n4054 GND.n2179 19.3944
R18624 GND.n4054 GND.n2175 19.3944
R18625 GND.n4060 GND.n2175 19.3944
R18626 GND.n4060 GND.n2173 19.3944
R18627 GND.n4064 GND.n2173 19.3944
R18628 GND.n4064 GND.n2169 19.3944
R18629 GND.n4070 GND.n2169 19.3944
R18630 GND.n4070 GND.n2167 19.3944
R18631 GND.n4074 GND.n2167 19.3944
R18632 GND.n4074 GND.n2163 19.3944
R18633 GND.n4080 GND.n2163 19.3944
R18634 GND.n4080 GND.n2161 19.3944
R18635 GND.n4084 GND.n2161 19.3944
R18636 GND.n4084 GND.n2157 19.3944
R18637 GND.n4090 GND.n2157 19.3944
R18638 GND.n4090 GND.n2155 19.3944
R18639 GND.n4126 GND.n2155 19.3944
R18640 GND.n4343 GND.n2136 19.3944
R18641 GND.n4333 GND.n2136 19.3944
R18642 GND.n4336 GND.n4333 19.3944
R18643 GND.n4336 GND.n2108 19.3944
R18644 GND.n4379 GND.n2108 19.3944
R18645 GND.n4379 GND.n2109 19.3944
R18646 GND.n4369 GND.n2109 19.3944
R18647 GND.n4372 GND.n4369 19.3944
R18648 GND.n4372 GND.n2079 19.3944
R18649 GND.n4422 GND.n2079 19.3944
R18650 GND.n4422 GND.n2080 19.3944
R18651 GND.n4416 GND.n2080 19.3944
R18652 GND.n4416 GND.n2045 19.3944
R18653 GND.n4461 GND.n2045 19.3944
R18654 GND.n4461 GND.n2046 19.3944
R18655 GND.n2052 GND.n2046 19.3944
R18656 GND.n4454 GND.n2052 19.3944
R18657 GND.n4454 GND.n2017 19.3944
R18658 GND.n4504 GND.n2017 19.3944
R18659 GND.n4504 GND.n2018 19.3944
R18660 GND.n4498 GND.n2018 19.3944
R18661 GND.n4498 GND.n1983 19.3944
R18662 GND.n4579 GND.n1983 19.3944
R18663 GND.n4579 GND.n1984 19.3944
R18664 GND.n1990 GND.n1984 19.3944
R18665 GND.n4572 GND.n1990 19.3944
R18666 GND.n4572 GND.n1953 19.3944
R18667 GND.n4611 GND.n1953 19.3944
R18668 GND.n4611 GND.n1954 19.3944
R18669 GND.n1956 GND.n1954 19.3944
R18670 GND.n1956 GND.n1888 19.3944
R18671 GND.n4683 GND.n1888 19.3944
R18672 GND.n4683 GND.n1889 19.3944
R18673 GND.n1896 GND.n1889 19.3944
R18674 GND.n1897 GND.n1896 19.3944
R18675 GND.n1898 GND.n1897 19.3944
R18676 GND.n1922 GND.n1898 19.3944
R18677 GND.n1922 GND.n1904 19.3944
R18678 GND.n1905 GND.n1904 19.3944
R18679 GND.n1906 GND.n1905 19.3944
R18680 GND.n4663 GND.n1906 19.3944
R18681 GND.n4665 GND.n4663 19.3944
R18682 GND.n4665 GND.n1842 19.3944
R18683 GND.n4738 GND.n1842 19.3944
R18684 GND.n4738 GND.n1843 19.3944
R18685 GND.n1849 GND.n1843 19.3944
R18686 GND.n4731 GND.n1849 19.3944
R18687 GND.n4731 GND.n1815 19.3944
R18688 GND.n4776 GND.n1815 19.3944
R18689 GND.n4776 GND.n1816 19.3944
R18690 GND.n4767 GND.n1816 19.3944
R18691 GND.n4769 GND.n4767 19.3944
R18692 GND.n4769 GND.n1781 19.3944
R18693 GND.n4844 GND.n1781 19.3944
R18694 GND.n4844 GND.n1782 19.3944
R18695 GND.n4834 GND.n1782 19.3944
R18696 GND.n4837 GND.n4834 19.3944
R18697 GND.n4837 GND.n1754 19.3944
R18698 GND.n4881 GND.n1754 19.3944
R18699 GND.n4881 GND.n1755 19.3944
R18700 GND.n4871 GND.n1755 19.3944
R18701 GND.n4874 GND.n4871 19.3944
R18702 GND.n4874 GND.n1724 19.3944
R18703 GND.n4919 GND.n1724 19.3944
R18704 GND.n4919 GND.n1725 19.3944
R18705 GND.n1727 GND.n1725 19.3944
R18706 GND.n1727 GND.n1696 19.3944
R18707 GND.n5879 GND.n1696 19.3944
R18708 GND.n5879 GND.n1697 19.3944
R18709 GND.n5867 GND.n1697 19.3944
R18710 GND.n5872 GND.n5867 19.3944
R18711 GND.n5872 GND.n5871 19.3944
R18712 GND.n5871 GND.n1603 19.3944
R18713 GND.n1626 GND.n1625 19.3944
R18714 GND.n1631 GND.n1630 19.3944
R18715 GND.n1634 GND.n1599 19.3944
R18716 GND.n4319 GND.n2148 18.8126
R18717 GND.n5931 GND.n5928 18.8126
R18718 GND.n7709 GND.n7708 18.8126
R18719 GND.n8434 GND.n8301 18.8126
R18720 GND.n378 GND.n356 18.8126
R18721 GND.n7729 GND.n7728 18.8126
R18722 GND.n4298 GND.n4297 18.8126
R18723 GND.n1640 GND.n1599 18.8126
R18724 GND.n5957 GND.n1658 18.6187
R18725 GND.n7685 GND.n7682 18.6187
R18726 GND.n1923 GND.t0 18.0422
R18727 GND.n5792 GND.n5791 18.0422
R18728 GND.n5791 GND.n5016 18.0422
R18729 GND.n5735 GND.n5734 18.0422
R18730 GND.n5734 GND.n5091 18.0422
R18731 GND.n5678 GND.n5677 18.0422
R18732 GND.n5677 GND.n5167 18.0422
R18733 GND.n6151 GND.n1535 18.0422
R18734 GND.n6151 GND.n6150 18.0422
R18735 GND.t195 GND.n1447 18.0422
R18736 GND.n6199 GND.n1447 18.0422
R18737 GND.n6600 GND.n1282 18.0422
R18738 GND.n1358 GND.n1282 18.0422
R18739 GND.n1210 GND.n1166 18.0422
R18740 GND.t213 GND.n1166 18.0422
R18741 GND.n6886 GND.n1103 18.0422
R18742 GND.n6735 GND.n1103 18.0422
R18743 GND.n7069 GND.n997 18.0422
R18744 GND.n7077 GND.n997 18.0422
R18745 GND.n7191 GND.n924 18.0422
R18746 GND.n7191 GND.n925 18.0422
R18747 GND.n859 GND.n858 18.0422
R18748 GND.n858 GND.n852 18.0422
R18749 GND.n8032 GND.t30 18.0422
R18750 GND.n6003 GND.n6002 18.0369
R18751 GND.n7632 GND.n7627 18.0369
R18752 GND.n8348 GND.n8343 18.0369
R18753 GND.n4219 GND.n4215 18.0369
R18754 GND.n5637 GND.t25 17.3205
R18755 GND.n6747 GND.t13 17.3205
R18756 GND.n6034 GND.n6033 17.2611
R18757 GND.n7675 GND.n7672 17.2611
R18758 GND.n8395 GND.n8392 17.2611
R18759 GND.n4262 GND.n4259 17.2611
R18760 GND.n5412 GND.t54 16.5988
R18761 GND.n5798 GND.n5006 16.5988
R18762 GND.n5436 GND.n5024 16.5988
R18763 GND.n5493 GND.n5099 16.5988
R18764 GND.n5684 GND.n5157 16.5988
R18765 GND.n5549 GND.n5175 16.5988
R18766 GND.n5623 GND.n1544 16.5988
R18767 GND.t197 GND.n1501 16.5988
R18768 GND.n6369 GND.n1455 16.5988
R18769 GND.n6237 GND.n1439 16.5988
R18770 GND.n6592 GND.n1290 16.5988
R18771 GND.n1365 GND.n1274 16.5988
R18772 GND.n6673 GND.n1214 16.5988
R18773 GND.n6826 GND.n1158 16.5988
R18774 GND.t209 GND.n1112 16.5988
R18775 GND.n6905 GND.n1087 16.5988
R18776 GND.n7058 GND.n1008 16.5988
R18777 GND.n7088 GND.n7087 16.5988
R18778 GND.n935 GND.n934 16.5988
R18779 GND.n7302 GND.n863 16.5988
R18780 GND.n7326 GND.n848 16.5988
R18781 GND.n5271 GND.n5248 16.0672
R18782 GND.n5261 GND.n5250 16.0672
R18783 GND.n775 GND.n774 16.0672
R18784 GND.n781 GND.n768 16.0672
R18785 GND.n5399 GND.t89 15.8772
R18786 GND.n5479 GND.t12 15.8772
R18787 GND.n7202 GND.t10 15.8772
R18788 GND.n6042 GND.n1613 15.5163
R18789 GND.n7725 GND.n706 15.5163
R18790 GND.n773 GND.n772 15.4533
R18791 GND.n5860 GND.t39 15.1555
R18792 GND.n5834 GND.n4962 15.1555
R18793 GND.n5806 GND.n5805 15.1555
R18794 GND.n5777 GND.n5034 15.1555
R18795 GND.n5749 GND.n5748 15.1555
R18796 GND.n5720 GND.n5109 15.1555
R18797 GND.n5692 GND.n5691 15.1555
R18798 GND.n5663 GND.n5185 15.1555
R18799 GND.n5598 GND.n1553 15.1555
R18800 GND.n6329 GND.n1493 15.1555
R18801 GND.t9 GND.n1469 15.1555
R18802 GND.n6361 GND.n1463 15.1555
R18803 GND.n6245 GND.n1430 15.1555
R18804 GND.n6584 GND.n1298 15.1555
R18805 GND.n1372 GND.n1266 15.1555
R18806 GND.n1397 GND.n1223 15.1555
R18807 GND.n6834 GND.n1150 15.1555
R18808 GND.t8 GND.n1144 15.1555
R18809 GND.n6866 GND.n1120 15.1555
R18810 GND.n1081 GND.n1057 15.1555
R18811 GND.n1019 GND.n1018 15.1555
R18812 GND.n984 GND.n978 15.1555
R18813 GND.n7171 GND.n939 15.1555
R18814 GND.n7240 GND.n7239 15.1555
R18815 GND.n7283 GND.n871 15.1555
R18816 GND.t47 GND.n619 15.1555
R18817 GND.n5881 GND.t39 14.4338
R18818 GND.t170 GND.n808 14.4338
R18819 GND.n7774 GND.t47 14.4338
R18820 GND.n5258 GND.n5251 14.2723
R18821 GND.n791 GND.n790 14.2723
R18822 GND.n5827 GND.n5826 13.7122
R18823 GND.n5812 GND.n4989 13.7122
R18824 GND.n5449 GND.n5042 13.7122
R18825 GND.n5755 GND.n5061 13.7122
R18826 GND.n5506 GND.n5117 13.7122
R18827 GND.n5698 GND.n5136 13.7122
R18828 GND.n5651 GND.n5650 13.7122
R18829 GND.n5637 GND.n5200 13.7122
R18830 GND.n6337 GND.n1485 13.7122
R18831 GND.n6353 GND.n1471 13.7122
R18832 GND.t211 GND.n1319 13.7122
R18833 GND.n6576 GND.n1306 13.7122
R18834 GND.n1379 GND.n1258 13.7122
R18835 GND.t199 GND.n1232 13.7122
R18836 GND.n6842 GND.n1142 13.7122
R18837 GND.n6858 GND.n1128 13.7122
R18838 GND.n6747 GND.n1041 13.7122
R18839 GND.n7039 GND.n1023 13.7122
R18840 GND.n7111 GND.n974 13.7122
R18841 GND.n7143 GND.n947 13.7122
R18842 GND.n902 GND.n897 13.7122
R18843 GND.n7272 GND.n882 13.7122
R18844 GND.n840 GND.t140 13.7122
R18845 GND.t36 GND.n822 13.7122
R18846 GND.n7368 GND.t155 13.7122
R18847 GND.n7442 GND.n7441 13.7122
R18848 GND.n6016 GND.n5984 13.3823
R18849 GND.n7652 GND.n7651 13.3823
R18850 GND.n8370 GND.n8332 13.3823
R18851 GND.n4239 GND.n4238 13.3823
R18852 GND.n5275 GND.n5246 13.1884
R18853 GND.n5270 GND.n5269 13.1884
R18854 GND.n5269 GND.n5268 13.1884
R18855 GND.n5264 GND.n5263 13.1884
R18856 GND.n5263 GND.n5262 13.1884
R18857 GND.n776 GND.n771 13.1884
R18858 GND.n777 GND.n776 13.1884
R18859 GND.n782 GND.n769 13.1884
R18860 GND.n783 GND.n782 13.1884
R18861 GND.n4962 GND.t118 12.9905
R18862 GND.n5799 GND.t104 12.9905
R18863 GND.n7313 GND.t75 12.9905
R18864 GND.n5277 GND.n5276 12.8005
R18865 GND.n7591 GND.n7539 12.8005
R18866 GND.n6020 GND.n5984 12.6066
R18867 GND.n7655 GND.n7652 12.6066
R18868 GND.n8373 GND.n8370 12.6066
R18869 GND.n4242 GND.n4239 12.6066
R18870 GND.n5820 GND.n4979 12.2688
R18871 GND.n5763 GND.n5052 12.2688
R18872 GND.n5457 GND.n5052 12.2688
R18873 GND.n5706 GND.n5127 12.2688
R18874 GND.n5514 GND.n5127 12.2688
R18875 GND.n1585 GND.n1584 12.2688
R18876 GND.n1584 GND.n1567 12.2688
R18877 GND.n6345 GND.n1477 12.2688
R18878 GND.n6345 GND.n1479 12.2688
R18879 GND.n6568 GND.n1313 12.2688
R18880 GND.n6445 GND.n1250 12.2688
R18881 GND.n6850 GND.n1134 12.2688
R18882 GND.n6850 GND.n1136 12.2688
R18883 GND.n7012 GND.n7011 12.2688
R18884 GND.n7011 GND.n7010 12.2688
R18885 GND.n965 GND.n958 12.2688
R18886 GND.n7132 GND.n958 12.2688
R18887 GND.n7259 GND.n893 12.2688
R18888 GND.n893 GND.n892 12.2688
R18889 GND.n7368 GND.n818 12.2688
R18890 GND.n818 GND.n817 12.2688
R18891 GND.t0 GND.n1921 11.5472
R18892 GND.n7336 GND.t75 11.5472
R18893 GND.t30 GND.n158 11.5472
R18894 GND.n5826 GND.n4971 10.8255
R18895 GND.n5452 GND.n5449 10.8255
R18896 GND.n5756 GND.n5755 10.8255
R18897 GND.n5509 GND.n5506 10.8255
R18898 GND.n5699 GND.n5698 10.8255
R18899 GND.n5650 GND.n5649 10.8255
R18900 GND.n5201 GND.n5200 10.8255
R18901 GND.n6337 GND.n1487 10.8255
R18902 GND.n6353 GND.n1469 10.8255
R18903 GND.t211 GND.n6560 10.8255
R18904 GND.n6568 GND.t11 10.8255
R18905 GND.n6576 GND.n1304 10.8255
R18906 GND.n6499 GND.n1379 10.8255
R18907 GND.n6445 GND.t24 10.8255
R18908 GND.n6475 GND.t199 10.8255
R18909 GND.n6842 GND.n1144 10.8255
R18910 GND.n6858 GND.n1126 10.8255
R18911 GND.n6999 GND.n1041 10.8255
R18912 GND.n1033 GND.n1023 10.8255
R18913 GND.n974 GND.n963 10.8255
R18914 GND.n7144 GND.n7143 10.8255
R18915 GND.n7253 GND.n897 10.8255
R18916 GND.n7265 GND.n882 10.8255
R18917 GND.n7362 GND.n822 10.8255
R18918 GND.n7442 GND.n806 10.8255
R18919 GND.n7375 GND.n735 10.6151
R18920 GND.n7378 GND.n7375 10.6151
R18921 GND.n7379 GND.n7378 10.6151
R18922 GND.n7383 GND.n7382 10.6151
R18923 GND.n7386 GND.n7383 10.6151
R18924 GND.n7387 GND.n7386 10.6151
R18925 GND.n7390 GND.n7387 10.6151
R18926 GND.n7391 GND.n7390 10.6151
R18927 GND.n7394 GND.n7391 10.6151
R18928 GND.n7395 GND.n7394 10.6151
R18929 GND.n7398 GND.n7395 10.6151
R18930 GND.n7399 GND.n7398 10.6151
R18931 GND.n7402 GND.n7399 10.6151
R18932 GND.n7403 GND.n7402 10.6151
R18933 GND.n7406 GND.n7403 10.6151
R18934 GND.n7407 GND.n7406 10.6151
R18935 GND.n7410 GND.n7407 10.6151
R18936 GND.n7411 GND.n7410 10.6151
R18937 GND.n7414 GND.n7411 10.6151
R18938 GND.n7415 GND.n7414 10.6151
R18939 GND.n7418 GND.n7415 10.6151
R18940 GND.n7419 GND.n7418 10.6151
R18941 GND.n7422 GND.n7419 10.6151
R18942 GND.n7423 GND.n7422 10.6151
R18943 GND.n5389 GND.n5388 10.6151
R18944 GND.n5392 GND.n5389 10.6151
R18945 GND.n5393 GND.n5392 10.6151
R18946 GND.n5394 GND.n5393 10.6151
R18947 GND.n5394 GND.n5217 10.6151
R18948 GND.n5402 GND.n5217 10.6151
R18949 GND.n5403 GND.n5402 10.6151
R18950 GND.n5405 GND.n5403 10.6151
R18951 GND.n5406 GND.n5405 10.6151
R18952 GND.n5407 GND.n5406 10.6151
R18953 GND.n5407 GND.n5216 10.6151
R18954 GND.n5415 GND.n5216 10.6151
R18955 GND.n5416 GND.n5415 10.6151
R18956 GND.n5419 GND.n5416 10.6151
R18957 GND.n5420 GND.n5419 10.6151
R18958 GND.n5421 GND.n5420 10.6151
R18959 GND.n5421 GND.n5215 10.6151
R18960 GND.n5429 GND.n5215 10.6151
R18961 GND.n5430 GND.n5429 10.6151
R18962 GND.n5432 GND.n5430 10.6151
R18963 GND.n5433 GND.n5432 10.6151
R18964 GND.n5434 GND.n5433 10.6151
R18965 GND.n5434 GND.n5214 10.6151
R18966 GND.n5442 GND.n5214 10.6151
R18967 GND.n5443 GND.n5442 10.6151
R18968 GND.n5445 GND.n5443 10.6151
R18969 GND.n5446 GND.n5445 10.6151
R18970 GND.n5447 GND.n5446 10.6151
R18971 GND.n5447 GND.n5213 10.6151
R18972 GND.n5455 GND.n5213 10.6151
R18973 GND.n5456 GND.n5455 10.6151
R18974 GND.n5459 GND.n5456 10.6151
R18975 GND.n5460 GND.n5459 10.6151
R18976 GND.n5461 GND.n5460 10.6151
R18977 GND.n5462 GND.n5461 10.6151
R18978 GND.n5462 GND.n5212 10.6151
R18979 GND.n5472 GND.n5212 10.6151
R18980 GND.n5473 GND.n5472 10.6151
R18981 GND.n5475 GND.n5473 10.6151
R18982 GND.n5476 GND.n5475 10.6151
R18983 GND.n5477 GND.n5476 10.6151
R18984 GND.n5477 GND.n5211 10.6151
R18985 GND.n5486 GND.n5211 10.6151
R18986 GND.n5487 GND.n5486 10.6151
R18987 GND.n5489 GND.n5487 10.6151
R18988 GND.n5490 GND.n5489 10.6151
R18989 GND.n5491 GND.n5490 10.6151
R18990 GND.n5491 GND.n5210 10.6151
R18991 GND.n5499 GND.n5210 10.6151
R18992 GND.n5500 GND.n5499 10.6151
R18993 GND.n5502 GND.n5500 10.6151
R18994 GND.n5503 GND.n5502 10.6151
R18995 GND.n5504 GND.n5503 10.6151
R18996 GND.n5504 GND.n5209 10.6151
R18997 GND.n5512 GND.n5209 10.6151
R18998 GND.n5513 GND.n5512 10.6151
R18999 GND.n5516 GND.n5513 10.6151
R19000 GND.n5517 GND.n5516 10.6151
R19001 GND.n5518 GND.n5517 10.6151
R19002 GND.n5519 GND.n5518 10.6151
R19003 GND.n5519 GND.n5208 10.6151
R19004 GND.n5529 GND.n5208 10.6151
R19005 GND.n5530 GND.n5529 10.6151
R19006 GND.n5532 GND.n5530 10.6151
R19007 GND.n5533 GND.n5532 10.6151
R19008 GND.n5534 GND.n5533 10.6151
R19009 GND.n5534 GND.n5207 10.6151
R19010 GND.n5542 GND.n5207 10.6151
R19011 GND.n5543 GND.n5542 10.6151
R19012 GND.n5545 GND.n5543 10.6151
R19013 GND.n5546 GND.n5545 10.6151
R19014 GND.n5547 GND.n5546 10.6151
R19015 GND.n5547 GND.n5206 10.6151
R19016 GND.n5555 GND.n5206 10.6151
R19017 GND.n5556 GND.n5555 10.6151
R19018 GND.n5558 GND.n5556 10.6151
R19019 GND.n5559 GND.n5558 10.6151
R19020 GND.n5560 GND.n5559 10.6151
R19021 GND.n5561 GND.n5560 10.6151
R19022 GND.n5562 GND.n5561 10.6151
R19023 GND.n5563 GND.n5562 10.6151
R19024 GND.n5563 GND.n5204 10.6151
R19025 GND.n5567 GND.n5204 10.6151
R19026 GND.n5568 GND.n5567 10.6151
R19027 GND.n5635 GND.n5568 10.6151
R19028 GND.n5635 GND.n5634 10.6151
R19029 GND.n5634 GND.n5633 10.6151
R19030 GND.n5633 GND.n5569 10.6151
R19031 GND.n5579 GND.n5569 10.6151
R19032 GND.n5588 GND.n5579 10.6151
R19033 GND.n5588 GND.n5587 10.6151
R19034 GND.n5587 GND.n5586 10.6151
R19035 GND.n5586 GND.n5582 10.6151
R19036 GND.n5582 GND.n5581 10.6151
R19037 GND.n5581 GND.n5580 10.6151
R19038 GND.n5580 GND.n1528 10.6151
R19039 GND.n6160 GND.n1528 10.6151
R19040 GND.n6161 GND.n6160 10.6151
R19041 GND.n6162 GND.n6161 10.6151
R19042 GND.n6162 GND.n1527 10.6151
R19043 GND.n6166 GND.n1527 10.6151
R19044 GND.n6167 GND.n6166 10.6151
R19045 GND.n6168 GND.n6167 10.6151
R19046 GND.n6171 GND.n6168 10.6151
R19047 GND.n6172 GND.n6171 10.6151
R19048 GND.n6174 GND.n6172 10.6151
R19049 GND.n6175 GND.n6174 10.6151
R19050 GND.n6296 GND.n6175 10.6151
R19051 GND.n6296 GND.n6295 10.6151
R19052 GND.n6295 GND.n6294 10.6151
R19053 GND.n6294 GND.n6176 10.6151
R19054 GND.n6188 GND.n6176 10.6151
R19055 GND.n6189 GND.n6188 10.6151
R19056 GND.n6282 GND.n6189 10.6151
R19057 GND.n6282 GND.n6281 10.6151
R19058 GND.n6281 GND.n6280 10.6151
R19059 GND.n6280 GND.n6190 10.6151
R19060 GND.n6202 GND.n6190 10.6151
R19061 GND.n6203 GND.n6202 10.6151
R19062 GND.n6268 GND.n6203 10.6151
R19063 GND.n6268 GND.n6267 10.6151
R19064 GND.n6267 GND.n6266 10.6151
R19065 GND.n6266 GND.n6204 10.6151
R19066 GND.n6248 GND.n6204 10.6151
R19067 GND.n6249 GND.n6248 10.6151
R19068 GND.n6254 GND.n6249 10.6151
R19069 GND.n6254 GND.n6253 10.6151
R19070 GND.n6253 GND.n6252 10.6151
R19071 GND.n6252 GND.n6250 10.6151
R19072 GND.n6250 GND.n1332 10.6151
R19073 GND.n6552 GND.n1332 10.6151
R19074 GND.n6552 GND.n6551 10.6151
R19075 GND.n6551 GND.n6550 10.6151
R19076 GND.n6550 GND.n1333 10.6151
R19077 GND.n1342 GND.n1333 10.6151
R19078 GND.n6539 GND.n1342 10.6151
R19079 GND.n6539 GND.n6538 10.6151
R19080 GND.n6538 GND.n6537 10.6151
R19081 GND.n6537 GND.n1343 10.6151
R19082 GND.n1354 GND.n1343 10.6151
R19083 GND.n1355 GND.n1354 10.6151
R19084 GND.n6525 GND.n1355 10.6151
R19085 GND.n6525 GND.n6524 10.6151
R19086 GND.n6524 GND.n6523 10.6151
R19087 GND.n6523 GND.n1356 10.6151
R19088 GND.n1368 GND.n1356 10.6151
R19089 GND.n1369 GND.n1368 10.6151
R19090 GND.n6511 GND.n1369 10.6151
R19091 GND.n6511 GND.n6510 10.6151
R19092 GND.n6510 GND.n6509 10.6151
R19093 GND.n6509 GND.n1370 10.6151
R19094 GND.n1382 GND.n1370 10.6151
R19095 GND.n1383 GND.n1382 10.6151
R19096 GND.n6497 GND.n1383 10.6151
R19097 GND.n6497 GND.n6496 10.6151
R19098 GND.n6496 GND.n6495 10.6151
R19099 GND.n6495 GND.n1384 10.6151
R19100 GND.n6491 GND.n1384 10.6151
R19101 GND.n6491 GND.n6490 10.6151
R19102 GND.n6490 GND.n6489 10.6151
R19103 GND.n6489 GND.n1386 10.6151
R19104 GND.n1396 GND.n1386 10.6151
R19105 GND.n1396 GND.n1395 10.6151
R19106 GND.n1395 GND.n1394 10.6151
R19107 GND.n1394 GND.n1390 10.6151
R19108 GND.n1390 GND.n1389 10.6151
R19109 GND.n1389 GND.n1388 10.6151
R19110 GND.n1388 GND.n1207 10.6151
R19111 GND.n6682 GND.n1207 10.6151
R19112 GND.n6683 GND.n6682 10.6151
R19113 GND.n6684 GND.n6683 10.6151
R19114 GND.n6684 GND.n1206 10.6151
R19115 GND.n6688 GND.n1206 10.6151
R19116 GND.n6689 GND.n6688 10.6151
R19117 GND.n6690 GND.n6689 10.6151
R19118 GND.n6693 GND.n6690 10.6151
R19119 GND.n6694 GND.n6693 10.6151
R19120 GND.n6695 GND.n6694 10.6151
R19121 GND.n6698 GND.n6695 10.6151
R19122 GND.n6699 GND.n6698 10.6151
R19123 GND.n6700 GND.n6699 10.6151
R19124 GND.n6703 GND.n6700 10.6151
R19125 GND.n6704 GND.n6703 10.6151
R19126 GND.n6706 GND.n6704 10.6151
R19127 GND.n6707 GND.n6706 10.6151
R19128 GND.n6779 GND.n6707 10.6151
R19129 GND.n6779 GND.n6778 10.6151
R19130 GND.n6778 GND.n6777 10.6151
R19131 GND.n6777 GND.n6708 10.6151
R19132 GND.n6744 GND.n6708 10.6151
R19133 GND.n6745 GND.n6744 10.6151
R19134 GND.n6765 GND.n6745 10.6151
R19135 GND.n6765 GND.n6764 10.6151
R19136 GND.n6764 GND.n6763 10.6151
R19137 GND.n6763 GND.n6760 10.6151
R19138 GND.n6760 GND.n6759 10.6151
R19139 GND.n6759 GND.n6758 10.6151
R19140 GND.n6758 GND.n6756 10.6151
R19141 GND.n6756 GND.n6755 10.6151
R19142 GND.n6755 GND.n6746 10.6151
R19143 GND.n6751 GND.n6746 10.6151
R19144 GND.n6751 GND.n6750 10.6151
R19145 GND.n6750 GND.n6749 10.6151
R19146 GND.n6749 GND.n1039 10.6151
R19147 GND.n7002 GND.n1039 10.6151
R19148 GND.n7003 GND.n7002 10.6151
R19149 GND.n7008 GND.n7003 10.6151
R19150 GND.n7008 GND.n7007 10.6151
R19151 GND.n7007 GND.n7006 10.6151
R19152 GND.n7006 GND.n7004 10.6151
R19153 GND.n7004 GND.n1015 10.6151
R19154 GND.n7047 GND.n1015 10.6151
R19155 GND.n7048 GND.n7047 10.6151
R19156 GND.n7049 GND.n7048 10.6151
R19157 GND.n7049 GND.n1006 10.6151
R19158 GND.n7060 GND.n1006 10.6151
R19159 GND.n7061 GND.n7060 10.6151
R19160 GND.n7067 GND.n7061 10.6151
R19161 GND.n7067 GND.n7066 10.6151
R19162 GND.n7066 GND.n7065 10.6151
R19163 GND.n7065 GND.n7064 10.6151
R19164 GND.n7064 GND.n7062 10.6151
R19165 GND.n7062 GND.n981 10.6151
R19166 GND.n7096 GND.n981 10.6151
R19167 GND.n7097 GND.n7096 10.6151
R19168 GND.n7103 GND.n7097 10.6151
R19169 GND.n7103 GND.n7102 10.6151
R19170 GND.n7102 GND.n7101 10.6151
R19171 GND.n7101 GND.n7100 10.6151
R19172 GND.n7100 GND.n7098 10.6151
R19173 GND.n7098 GND.n956 10.6151
R19174 GND.n7134 GND.n956 10.6151
R19175 GND.n7135 GND.n7134 10.6151
R19176 GND.n7141 GND.n7135 10.6151
R19177 GND.n7141 GND.n7140 10.6151
R19178 GND.n7140 GND.n7139 10.6151
R19179 GND.n7139 GND.n7138 10.6151
R19180 GND.n7138 GND.n7136 10.6151
R19181 GND.n7136 GND.n931 10.6151
R19182 GND.n7179 GND.n931 10.6151
R19183 GND.n7180 GND.n7179 10.6151
R19184 GND.n7182 GND.n7180 10.6151
R19185 GND.n7182 GND.n7181 10.6151
R19186 GND.n7181 GND.n922 10.6151
R19187 GND.n7194 GND.n922 10.6151
R19188 GND.n7195 GND.n7194 10.6151
R19189 GND.n7200 GND.n7195 10.6151
R19190 GND.n7200 GND.n7199 10.6151
R19191 GND.n7199 GND.n7198 10.6151
R19192 GND.n7198 GND.n7196 10.6151
R19193 GND.n7196 GND.n899 10.6151
R19194 GND.n7248 GND.n899 10.6151
R19195 GND.n7249 GND.n7248 10.6151
R19196 GND.n7250 GND.n7249 10.6151
R19197 GND.n7250 GND.n889 10.6151
R19198 GND.n7261 GND.n889 10.6151
R19199 GND.n7262 GND.n7261 10.6151
R19200 GND.n7263 GND.n7262 10.6151
R19201 GND.n7263 GND.n880 10.6151
R19202 GND.n7274 GND.n880 10.6151
R19203 GND.n7275 GND.n7274 10.6151
R19204 GND.n7281 GND.n7275 10.6151
R19205 GND.n7281 GND.n7280 10.6151
R19206 GND.n7280 GND.n7279 10.6151
R19207 GND.n7279 GND.n7278 10.6151
R19208 GND.n7278 GND.n7276 10.6151
R19209 GND.n7276 GND.n855 10.6151
R19210 GND.n7310 GND.n855 10.6151
R19211 GND.n7311 GND.n7310 10.6151
R19212 GND.n7318 GND.n7311 10.6151
R19213 GND.n7318 GND.n7317 10.6151
R19214 GND.n7317 GND.n7316 10.6151
R19215 GND.n7316 GND.n7315 10.6151
R19216 GND.n7315 GND.n7312 10.6151
R19217 GND.n7312 GND.n832 10.6151
R19218 GND.n7345 GND.n832 10.6151
R19219 GND.n7346 GND.n7345 10.6151
R19220 GND.n7348 GND.n7346 10.6151
R19221 GND.n7348 GND.n7347 10.6151
R19222 GND.n7347 GND.n815 10.6151
R19223 GND.n7370 GND.n815 10.6151
R19224 GND.n7371 GND.n7370 10.6151
R19225 GND.n7433 GND.n7371 10.6151
R19226 GND.n7433 GND.n7432 10.6151
R19227 GND.n7432 GND.n7431 10.6151
R19228 GND.n7431 GND.n7430 10.6151
R19229 GND.n7430 GND.n7428 10.6151
R19230 GND.n7428 GND.n7427 10.6151
R19231 GND.n5337 GND.n5231 10.6151
R19232 GND.n5338 GND.n5337 10.6151
R19233 GND.n5342 GND.n5338 10.6151
R19234 GND.n5348 GND.n5229 10.6151
R19235 GND.n5349 GND.n5348 10.6151
R19236 GND.n5350 GND.n5349 10.6151
R19237 GND.n5350 GND.n5227 10.6151
R19238 GND.n5356 GND.n5227 10.6151
R19239 GND.n5357 GND.n5356 10.6151
R19240 GND.n5358 GND.n5357 10.6151
R19241 GND.n5358 GND.n5225 10.6151
R19242 GND.n5364 GND.n5225 10.6151
R19243 GND.n5365 GND.n5364 10.6151
R19244 GND.n5366 GND.n5365 10.6151
R19245 GND.n5366 GND.n5223 10.6151
R19246 GND.n5372 GND.n5223 10.6151
R19247 GND.n5373 GND.n5372 10.6151
R19248 GND.n5374 GND.n5373 10.6151
R19249 GND.n5374 GND.n5221 10.6151
R19250 GND.n5380 GND.n5221 10.6151
R19251 GND.n5381 GND.n5380 10.6151
R19252 GND.n5382 GND.n5381 10.6151
R19253 GND.n5382 GND.n5219 10.6151
R19254 GND.n5219 GND.n5218 10.6151
R19255 GND.n5277 GND.n5245 10.6151
R19256 GND.n5245 GND.n5244 10.6151
R19257 GND.n5284 GND.n5244 10.6151
R19258 GND.n5285 GND.n5284 10.6151
R19259 GND.n5286 GND.n5285 10.6151
R19260 GND.n5286 GND.n5242 10.6151
R19261 GND.n5292 GND.n5242 10.6151
R19262 GND.n5293 GND.n5292 10.6151
R19263 GND.n5294 GND.n5293 10.6151
R19264 GND.n5294 GND.n5240 10.6151
R19265 GND.n5300 GND.n5240 10.6151
R19266 GND.n5301 GND.n5300 10.6151
R19267 GND.n5302 GND.n5301 10.6151
R19268 GND.n5302 GND.n5238 10.6151
R19269 GND.n5308 GND.n5238 10.6151
R19270 GND.n5309 GND.n5308 10.6151
R19271 GND.n5310 GND.n5309 10.6151
R19272 GND.n5310 GND.n5236 10.6151
R19273 GND.n5316 GND.n5236 10.6151
R19274 GND.n5317 GND.n5316 10.6151
R19275 GND.n5321 GND.n5317 10.6151
R19276 GND.n5327 GND.n5234 10.6151
R19277 GND.n5328 GND.n5327 10.6151
R19278 GND.n5329 GND.n5328 10.6151
R19279 GND.n7591 GND.n7590 10.6151
R19280 GND.n7590 GND.n7589 10.6151
R19281 GND.n7589 GND.n7586 10.6151
R19282 GND.n7586 GND.n7585 10.6151
R19283 GND.n7585 GND.n7582 10.6151
R19284 GND.n7582 GND.n7581 10.6151
R19285 GND.n7581 GND.n7578 10.6151
R19286 GND.n7578 GND.n7577 10.6151
R19287 GND.n7577 GND.n7574 10.6151
R19288 GND.n7574 GND.n7573 10.6151
R19289 GND.n7573 GND.n7570 10.6151
R19290 GND.n7570 GND.n7569 10.6151
R19291 GND.n7569 GND.n7566 10.6151
R19292 GND.n7566 GND.n7565 10.6151
R19293 GND.n7565 GND.n7562 10.6151
R19294 GND.n7562 GND.n7561 10.6151
R19295 GND.n7561 GND.n7558 10.6151
R19296 GND.n7558 GND.n7557 10.6151
R19297 GND.n7557 GND.n7554 10.6151
R19298 GND.n7554 GND.n7553 10.6151
R19299 GND.n7553 GND.n7550 10.6151
R19300 GND.n7548 GND.n7545 10.6151
R19301 GND.n7545 GND.n7544 10.6151
R19302 GND.n7544 GND.n736 10.6151
R19303 GND.n5831 GND.n4966 10.6151
R19304 GND.n5831 GND.n5830 10.6151
R19305 GND.n5830 GND.n5829 10.6151
R19306 GND.n5829 GND.n4967 10.6151
R19307 GND.n5397 GND.n4967 10.6151
R19308 GND.n5397 GND.n4984 10.6151
R19309 GND.n5817 GND.n4984 10.6151
R19310 GND.n5817 GND.n5816 10.6151
R19311 GND.n5816 GND.n5815 10.6151
R19312 GND.n5815 GND.n4985 10.6151
R19313 GND.n5410 GND.n4985 10.6151
R19314 GND.n5410 GND.n5002 10.6151
R19315 GND.n5803 GND.n5002 10.6151
R19316 GND.n5803 GND.n5802 10.6151
R19317 GND.n5802 GND.n5801 10.6151
R19318 GND.n5801 GND.n5003 10.6151
R19319 GND.n5424 GND.n5003 10.6151
R19320 GND.n5424 GND.n5019 10.6151
R19321 GND.n5789 GND.n5019 10.6151
R19322 GND.n5789 GND.n5788 10.6151
R19323 GND.n5788 GND.n5787 10.6151
R19324 GND.n5787 GND.n5020 10.6151
R19325 GND.n5437 GND.n5020 10.6151
R19326 GND.n5437 GND.n5037 10.6151
R19327 GND.n5775 GND.n5037 10.6151
R19328 GND.n5775 GND.n5774 10.6151
R19329 GND.n5774 GND.n5773 10.6151
R19330 GND.n5773 GND.n5038 10.6151
R19331 GND.n5450 GND.n5038 10.6151
R19332 GND.n5450 GND.n5055 10.6151
R19333 GND.n5761 GND.n5055 10.6151
R19334 GND.n5761 GND.n5760 10.6151
R19335 GND.n5760 GND.n5759 10.6151
R19336 GND.n5759 GND.n5056 10.6151
R19337 GND.n5466 GND.n5056 10.6151
R19338 GND.n5467 GND.n5466 10.6151
R19339 GND.n5467 GND.n5077 10.6151
R19340 GND.n5746 GND.n5077 10.6151
R19341 GND.n5746 GND.n5745 10.6151
R19342 GND.n5745 GND.n5744 10.6151
R19343 GND.n5744 GND.n5078 10.6151
R19344 GND.n5481 GND.n5078 10.6151
R19345 GND.n5481 GND.n5094 10.6151
R19346 GND.n5732 GND.n5094 10.6151
R19347 GND.n5732 GND.n5731 10.6151
R19348 GND.n5731 GND.n5730 10.6151
R19349 GND.n5730 GND.n5095 10.6151
R19350 GND.n5494 GND.n5095 10.6151
R19351 GND.n5494 GND.n5112 10.6151
R19352 GND.n5718 GND.n5112 10.6151
R19353 GND.n5718 GND.n5717 10.6151
R19354 GND.n5717 GND.n5716 10.6151
R19355 GND.n5716 GND.n5113 10.6151
R19356 GND.n5507 GND.n5113 10.6151
R19357 GND.n5507 GND.n5130 10.6151
R19358 GND.n5704 GND.n5130 10.6151
R19359 GND.n5704 GND.n5703 10.6151
R19360 GND.n5703 GND.n5702 10.6151
R19361 GND.n5702 GND.n5131 10.6151
R19362 GND.n5523 GND.n5131 10.6151
R19363 GND.n5524 GND.n5523 10.6151
R19364 GND.n5524 GND.n5151 10.6151
R19365 GND.n5689 GND.n5151 10.6151
R19366 GND.n5689 GND.n5688 10.6151
R19367 GND.n5688 GND.n5687 10.6151
R19368 GND.n5687 GND.n5152 10.6151
R19369 GND.n5537 GND.n5152 10.6151
R19370 GND.n5537 GND.n5170 10.6151
R19371 GND.n5675 GND.n5170 10.6151
R19372 GND.n5675 GND.n5674 10.6151
R19373 GND.n5674 GND.n5673 10.6151
R19374 GND.n5673 GND.n5171 10.6151
R19375 GND.n5550 GND.n5171 10.6151
R19376 GND.n5550 GND.n5188 10.6151
R19377 GND.n5661 GND.n5188 10.6151
R19378 GND.n5661 GND.n5660 10.6151
R19379 GND.n5660 GND.n5659 10.6151
R19380 GND.n5659 GND.n5189 10.6151
R19381 GND.n5647 GND.n5189 10.6151
R19382 GND.n5647 GND.n5646 10.6151
R19383 GND.n5646 GND.n5645 10.6151
R19384 GND.n5645 GND.n5196 10.6151
R19385 GND.n5641 GND.n5196 10.6151
R19386 GND.n5641 GND.n5640 10.6151
R19387 GND.n5640 GND.n5639 10.6151
R19388 GND.n5639 GND.n5198 10.6151
R19389 GND.n5629 GND.n5198 10.6151
R19390 GND.n5629 GND.n5628 10.6151
R19391 GND.n5628 GND.n5627 10.6151
R19392 GND.n5627 GND.n5572 10.6151
R19393 GND.n5575 GND.n5572 10.6151
R19394 GND.n5575 GND.n5574 10.6151
R19395 GND.n5574 GND.n1533 10.6151
R19396 GND.n6153 GND.n1533 10.6151
R19397 GND.n6154 GND.n6153 10.6151
R19398 GND.n6155 GND.n6154 10.6151
R19399 GND.n6155 GND.n1508 10.6151
R19400 GND.n6319 GND.n1508 10.6151
R19401 GND.n6319 GND.n6318 10.6151
R19402 GND.n6318 GND.n6317 10.6151
R19403 GND.n6317 GND.n1509 10.6151
R19404 GND.n1511 GND.n1509 10.6151
R19405 GND.n1521 GND.n1511 10.6151
R19406 GND.n1522 GND.n1521 10.6151
R19407 GND.n6303 GND.n1522 10.6151
R19408 GND.n6303 GND.n6302 10.6151
R19409 GND.n6302 GND.n6301 10.6151
R19410 GND.n6301 GND.n1523 10.6151
R19411 GND.n6181 GND.n1523 10.6151
R19412 GND.n6182 GND.n6181 10.6151
R19413 GND.n6289 GND.n6182 10.6151
R19414 GND.n6289 GND.n6288 10.6151
R19415 GND.n6288 GND.n6287 10.6151
R19416 GND.n6287 GND.n6183 10.6151
R19417 GND.n6195 GND.n6183 10.6151
R19418 GND.n6196 GND.n6195 10.6151
R19419 GND.n6275 GND.n6196 10.6151
R19420 GND.n6275 GND.n6274 10.6151
R19421 GND.n6274 GND.n6273 10.6151
R19422 GND.n6273 GND.n6197 10.6151
R19423 GND.n6240 GND.n6197 10.6151
R19424 GND.n6241 GND.n6240 10.6151
R19425 GND.n6261 GND.n6241 10.6151
R19426 GND.n6261 GND.n6260 10.6151
R19427 GND.n6260 GND.n6259 10.6151
R19428 GND.n6259 GND.n6242 10.6151
R19429 GND.n6243 GND.n6242 10.6151
R19430 GND.n6243 GND.n1326 10.6151
R19431 GND.n6558 GND.n1326 10.6151
R19432 GND.n6558 GND.n6557 10.6151
R19433 GND.n6557 GND.n6556 10.6151
R19434 GND.n6556 GND.n1327 10.6151
R19435 GND.n6546 GND.n1327 10.6151
R19436 GND.n6546 GND.n6545 10.6151
R19437 GND.n6545 GND.n6544 10.6151
R19438 GND.n6544 GND.n1337 10.6151
R19439 GND.n1347 GND.n1337 10.6151
R19440 GND.n1348 GND.n1347 10.6151
R19441 GND.n6532 GND.n1348 10.6151
R19442 GND.n6532 GND.n6531 10.6151
R19443 GND.n6531 GND.n6530 10.6151
R19444 GND.n6530 GND.n1349 10.6151
R19445 GND.n1361 GND.n1349 10.6151
R19446 GND.n1362 GND.n1361 10.6151
R19447 GND.n6518 GND.n1362 10.6151
R19448 GND.n6518 GND.n6517 10.6151
R19449 GND.n6517 GND.n6516 10.6151
R19450 GND.n6516 GND.n1363 10.6151
R19451 GND.n1375 GND.n1363 10.6151
R19452 GND.n1376 GND.n1375 10.6151
R19453 GND.n6504 GND.n1376 10.6151
R19454 GND.n6504 GND.n6503 10.6151
R19455 GND.n6503 GND.n6502 10.6151
R19456 GND.n6502 GND.n1377 10.6151
R19457 GND.n1402 GND.n1377 10.6151
R19458 GND.n1404 GND.n1402 10.6151
R19459 GND.n1405 GND.n1404 10.6151
R19460 GND.n1406 GND.n1405 10.6151
R19461 GND.n1406 GND.n1400 10.6151
R19462 GND.n6478 GND.n1400 10.6151
R19463 GND.n6479 GND.n6478 10.6151
R19464 GND.n6483 GND.n6479 10.6151
R19465 GND.n6483 GND.n6482 10.6151
R19466 GND.n6482 GND.n6481 10.6151
R19467 GND.n6481 GND.n1212 10.6151
R19468 GND.n6675 GND.n1212 10.6151
R19469 GND.n6676 GND.n6675 10.6151
R19470 GND.n6677 GND.n6676 10.6151
R19471 GND.n6677 GND.n1173 10.6151
R19472 GND.n6816 GND.n1173 10.6151
R19473 GND.n6816 GND.n6815 10.6151
R19474 GND.n6815 GND.n6814 10.6151
R19475 GND.n6814 GND.n1174 10.6151
R19476 GND.n1176 GND.n1174 10.6151
R19477 GND.n1186 GND.n1176 10.6151
R19478 GND.n1187 GND.n1186 10.6151
R19479 GND.n6800 GND.n1187 10.6151
R19480 GND.n6800 GND.n6799 10.6151
R19481 GND.n6799 GND.n6798 10.6151
R19482 GND.n6798 GND.n1188 10.6151
R19483 GND.n1199 GND.n1188 10.6151
R19484 GND.n1200 GND.n1199 10.6151
R19485 GND.n6786 GND.n1200 10.6151
R19486 GND.n6786 GND.n6785 10.6151
R19487 GND.n6785 GND.n6784 10.6151
R19488 GND.n6784 GND.n1201 10.6151
R19489 GND.n6713 GND.n1201 10.6151
R19490 GND.n6714 GND.n6713 10.6151
R19491 GND.n6772 GND.n6714 10.6151
R19492 GND.n6772 GND.n6771 10.6151
R19493 GND.n6771 GND.n6770 10.6151
R19494 GND.n6770 GND.n6715 10.6151
R19495 GND.n6718 GND.n6715 10.6151
R19496 GND.n6718 GND.n6717 10.6151
R19497 GND.n6717 GND.n1091 10.6151
R19498 GND.n6897 GND.n1091 10.6151
R19499 GND.n6898 GND.n6897 10.6151
R19500 GND.n6902 GND.n6898 10.6151
R19501 GND.n6902 GND.n6901 10.6151
R19502 GND.n6901 GND.n6900 10.6151
R19503 GND.n6900 GND.n1043 10.6151
R19504 GND.n6995 GND.n1043 10.6151
R19505 GND.n6996 GND.n6995 10.6151
R19506 GND.n6997 GND.n6996 10.6151
R19507 GND.n6997 GND.n1035 10.6151
R19508 GND.n7014 GND.n1035 10.6151
R19509 GND.n7015 GND.n7014 10.6151
R19510 GND.n7016 GND.n7015 10.6151
R19511 GND.n7016 GND.n1021 10.6151
R19512 GND.n7041 GND.n1021 10.6151
R19513 GND.n7042 GND.n7041 10.6151
R19514 GND.n7043 GND.n7042 10.6151
R19515 GND.n7043 GND.n1011 10.6151
R19516 GND.n7054 GND.n1011 10.6151
R19517 GND.n7055 GND.n7054 10.6151
R19518 GND.n7056 GND.n7055 10.6151
R19519 GND.n7056 GND.n1001 10.6151
R19520 GND.n7072 GND.n1001 10.6151
R19521 GND.n7073 GND.n7072 10.6151
R19522 GND.n7074 GND.n7073 10.6151
R19523 GND.n7074 GND.n987 10.6151
R19524 GND.n7090 GND.n987 10.6151
R19525 GND.n7091 GND.n7090 10.6151
R19526 GND.n7092 GND.n7091 10.6151
R19527 GND.n7092 GND.n976 10.6151
R19528 GND.n7107 GND.n976 10.6151
R19529 GND.n7108 GND.n7107 10.6151
R19530 GND.n7109 GND.n7108 10.6151
R19531 GND.n7109 GND.n961 10.6151
R19532 GND.n7128 GND.n961 10.6151
R19533 GND.n7129 GND.n7128 10.6151
R19534 GND.n7130 GND.n7129 10.6151
R19535 GND.n7130 GND.n951 10.6151
R19536 GND.n7146 GND.n951 10.6151
R19537 GND.n7147 GND.n7146 10.6151
R19538 GND.n7148 GND.n7147 10.6151
R19539 GND.n7148 GND.n937 10.6151
R19540 GND.n7173 GND.n937 10.6151
R19541 GND.n7174 GND.n7173 10.6151
R19542 GND.n7175 GND.n7174 10.6151
R19543 GND.n7175 GND.n927 10.6151
R19544 GND.n7187 GND.n927 10.6151
R19545 GND.n7188 GND.n7187 10.6151
R19546 GND.n7189 GND.n7188 10.6151
R19547 GND.n7189 GND.n918 10.6151
R19548 GND.n7206 GND.n918 10.6151
R19549 GND.n7207 GND.n7206 10.6151
R19550 GND.n7208 GND.n7207 10.6151
R19551 GND.n7208 GND.n905 10.6151
R19552 GND.n7242 GND.n905 10.6151
R19553 GND.n7243 GND.n7242 10.6151
R19554 GND.n7244 GND.n7243 10.6151
R19555 GND.n7244 GND.n895 10.6151
R19556 GND.n7255 GND.n895 10.6151
R19557 GND.n7256 GND.n7255 10.6151
R19558 GND.n7257 GND.n7256 10.6151
R19559 GND.n7257 GND.n885 10.6151
R19560 GND.n7268 GND.n885 10.6151
R19561 GND.n7269 GND.n7268 10.6151
R19562 GND.n7270 GND.n7269 10.6151
R19563 GND.n7270 GND.n875 10.6151
R19564 GND.n7286 GND.n875 10.6151
R19565 GND.n7287 GND.n7286 10.6151
R19566 GND.n7288 GND.n7287 10.6151
R19567 GND.n7288 GND.n861 10.6151
R19568 GND.n7304 GND.n861 10.6151
R19569 GND.n7305 GND.n7304 10.6151
R19570 GND.n7306 GND.n7305 10.6151
R19571 GND.n7306 GND.n850 10.6151
R19572 GND.n7322 GND.n850 10.6151
R19573 GND.n7323 GND.n7322 10.6151
R19574 GND.n7324 GND.n7323 10.6151
R19575 GND.n7324 GND.n837 10.6151
R19576 GND.n7338 GND.n837 10.6151
R19577 GND.n7339 GND.n7338 10.6151
R19578 GND.n7341 GND.n7339 10.6151
R19579 GND.n7341 GND.n7340 10.6151
R19580 GND.n7340 GND.n820 10.6151
R19581 GND.n7364 GND.n820 10.6151
R19582 GND.n7365 GND.n7364 10.6151
R19583 GND.n7366 GND.n7365 10.6151
R19584 GND.n7366 GND.n810 10.6151
R19585 GND.n7437 GND.n810 10.6151
R19586 GND.n7438 GND.n7437 10.6151
R19587 GND.n7439 GND.n7438 10.6151
R19588 GND.n7439 GND.n796 10.6151
R19589 GND.n7537 GND.n796 10.6151
R19590 GND.n7538 GND.n7537 10.6151
R19591 GND.n5267 GND.n5248 10.2247
R19592 GND.n5265 GND.n5250 10.2247
R19593 GND.n775 GND.n770 10.2247
R19594 GND.n781 GND.n780 10.2247
R19595 GND.n7360 GND.t155 10.1038
R19596 GND.n18 GND.t34 9.75419
R19597 GND.n18 GND.t239 9.75419
R19598 GND.n20 GND.t187 9.75419
R19599 GND.n20 GND.t223 9.75419
R19600 GND.n29 GND.t21 9.75419
R19601 GND.n29 GND.t180 9.75419
R19602 GND.n31 GND.t192 9.75419
R19603 GND.n31 GND.t218 9.75419
R19604 GND.n41 GND.t178 9.75419
R19605 GND.n41 GND.t216 9.75419
R19606 GND.n43 GND.t26 9.75419
R19607 GND.n43 GND.t233 9.75419
R19608 GND.n53 GND.t1 9.75419
R19609 GND.n53 GND.t238 9.75419
R19610 GND.n55 GND.t183 9.75419
R19611 GND.n55 GND.t222 9.75419
R19612 GND.n65 GND.t22 9.75419
R19613 GND.n65 GND.t182 9.75419
R19614 GND.n67 GND.t29 9.75419
R19615 GND.n67 GND.t7 9.75419
R19616 GND.n7 GND.t228 9.75419
R19617 GND.n7 GND.t15 9.75419
R19618 GND.n9 GND.t17 9.75419
R19619 GND.n9 GND.t229 9.75419
R19620 GND.n82 GND.t186 9.75419
R19621 GND.n82 GND.t234 9.75419
R19622 GND.n81 GND.t32 9.75419
R19623 GND.n81 GND.t225 9.75419
R19624 GND.n93 GND.t181 9.75419
R19625 GND.n93 GND.t193 9.75419
R19626 GND.n92 GND.t20 9.75419
R19627 GND.n92 GND.t179 9.75419
R19628 GND.n105 GND.t190 9.75419
R19629 GND.n105 GND.t5 9.75419
R19630 GND.n104 GND.t3 9.75419
R19631 GND.n104 GND.t194 9.75419
R19632 GND.n117 GND.t220 9.75419
R19633 GND.n117 GND.t33 9.75419
R19634 GND.n116 GND.t219 9.75419
R19635 GND.n116 GND.t185 9.75419
R19636 GND.n129 GND.t215 9.75419
R19637 GND.n129 GND.t232 9.75419
R19638 GND.n128 GND.t175 9.75419
R19639 GND.n128 GND.t177 9.75419
R19640 GND.n141 GND.t31 9.75419
R19641 GND.n141 GND.t221 9.75419
R19642 GND.n140 GND.t231 9.75419
R19643 GND.n140 GND.t217 9.75419
R19644 GND.n14 GND.n12 9.71174
R19645 GND.n25 GND.n23 9.71174
R19646 GND.n37 GND.n35 9.71174
R19647 GND.n49 GND.n47 9.71174
R19648 GND.n61 GND.n59 9.71174
R19649 GND.n3 GND.n1 9.71174
R19650 GND.n87 GND.n85 9.71174
R19651 GND.n98 GND.n96 9.71174
R19652 GND.n110 GND.n108 9.71174
R19653 GND.n122 GND.n120 9.71174
R19654 GND.n134 GND.n132 9.71174
R19655 GND.n146 GND.n144 9.71174
R19656 GND.n17 GND.n16 9.45567
R19657 GND.n28 GND.n27 9.45567
R19658 GND.n40 GND.n39 9.45567
R19659 GND.n52 GND.n51 9.45567
R19660 GND.n64 GND.n63 9.45567
R19661 GND.n6 GND.n5 9.45567
R19662 GND.n90 GND.n89 9.45567
R19663 GND.n101 GND.n100 9.45567
R19664 GND.n113 GND.n112 9.45567
R19665 GND.n125 GND.n124 9.45567
R19666 GND.n137 GND.n136 9.45567
R19667 GND.n149 GND.n148 9.45567
R19668 GND.n5834 GND.n5833 9.38216
R19669 GND.n5806 GND.n4997 9.38216
R19670 GND.n5040 GND.n5034 9.38216
R19671 GND.n5749 GND.n5072 9.38216
R19672 GND.n5115 GND.n5109 9.38216
R19673 GND.n5692 GND.n5147 9.38216
R19674 GND.n5191 GND.n5185 9.38216
R19675 GND.n6329 GND.n1495 9.38216
R19676 GND.n6298 GND.t9 9.38216
R19677 GND.n6361 GND.n1461 9.38216
R19678 GND.n6256 GND.n6245 9.38216
R19679 GND.n6584 GND.n1296 9.38216
R19680 GND.n6506 GND.n1372 9.38216
R19681 GND.n6485 GND.n1397 9.38216
R19682 GND.n6834 GND.n1152 9.38216
R19683 GND.n6795 GND.t8 9.38216
R19684 GND.n6866 GND.n1118 9.38216
R19685 GND.n7045 GND.n1019 9.38216
R19686 GND.n7105 GND.n978 9.38216
R19687 GND.n949 GND.n939 9.38216
R19688 GND.n7239 GND.n901 9.38216
R19689 GND.n7284 GND.n7283 9.38216
R19690 GND.n7343 GND.n834 9.38216
R19691 GND.n7535 GND.n7534 9.38216
R19692 GND.n7534 GND.t112 9.38216
R19693 GND.n7382 GND.n7374 9.36635
R19694 GND.n5341 GND.n5229 9.36635
R19695 GND.n5321 GND.n5320 9.36635
R19696 GND.n7550 GND.n7549 9.36635
R19697 GND.n16 GND.n15 9.3005
R19698 GND.n27 GND.n26 9.3005
R19699 GND.n39 GND.n38 9.3005
R19700 GND.n51 GND.n50 9.3005
R19701 GND.n63 GND.n62 9.3005
R19702 GND.n5 GND.n4 9.3005
R19703 GND.n4646 GND.n1916 9.3005
R19704 GND.n4650 GND.n4647 9.3005
R19705 GND.n4649 GND.n4648 9.3005
R19706 GND.n1862 GND.n1861 9.3005
R19707 GND.n4697 GND.n4696 9.3005
R19708 GND.n4698 GND.n1860 9.3005
R19709 GND.n4702 GND.n4699 9.3005
R19710 GND.n4701 GND.n4700 9.3005
R19711 GND.n1825 GND.n1824 9.3005
R19712 GND.n4753 GND.n4752 9.3005
R19713 GND.n4754 GND.n1823 9.3005
R19714 GND.n4758 GND.n4755 9.3005
R19715 GND.n4757 GND.n4756 9.3005
R19716 GND.n1797 GND.n1796 9.3005
R19717 GND.n4791 GND.n4790 9.3005
R19718 GND.n4792 GND.n1795 9.3005
R19719 GND.n4796 GND.n4793 9.3005
R19720 GND.n4795 GND.n4794 9.3005
R19721 GND.n1764 GND.n1763 9.3005
R19722 GND.n4859 GND.n4858 9.3005
R19723 GND.n4860 GND.n1762 9.3005
R19724 GND.n4864 GND.n4861 9.3005
R19725 GND.n4863 GND.n4862 9.3005
R19726 GND.n1736 GND.n1735 9.3005
R19727 GND.n4896 GND.n4895 9.3005
R19728 GND.n4897 GND.n1734 9.3005
R19729 GND.n4910 GND.n4898 9.3005
R19730 GND.n4909 GND.n4899 9.3005
R19731 GND.n4908 GND.n4900 9.3005
R19732 GND.n4906 GND.n4901 9.3005
R19733 GND.n4905 GND.n4902 9.3005
R19734 GND.n4904 GND.n4903 9.3005
R19735 GND.n1680 GND.n1679 9.3005
R19736 GND.n5893 GND.n5892 9.3005
R19737 GND.n5894 GND.n1678 9.3005
R19738 GND.n5897 GND.n5895 9.3005
R19739 GND.n5896 GND.n1595 9.3005
R19740 GND.n3934 GND.n3933 9.3005
R19741 GND.n3932 GND.n2251 9.3005
R19742 GND.n3931 GND.n3930 9.3005
R19743 GND.n2253 GND.n2252 9.3005
R19744 GND.n3924 GND.n2257 9.3005
R19745 GND.n3923 GND.n2258 9.3005
R19746 GND.n3922 GND.n2259 9.3005
R19747 GND.n2264 GND.n2260 9.3005
R19748 GND.n3916 GND.n2265 9.3005
R19749 GND.n3915 GND.n2266 9.3005
R19750 GND.n3914 GND.n2267 9.3005
R19751 GND.n2272 GND.n2268 9.3005
R19752 GND.n3908 GND.n2273 9.3005
R19753 GND.n3907 GND.n2274 9.3005
R19754 GND.n3906 GND.n2275 9.3005
R19755 GND.n2280 GND.n2276 9.3005
R19756 GND.n3900 GND.n2281 9.3005
R19757 GND.n3899 GND.n2282 9.3005
R19758 GND.n3898 GND.n2283 9.3005
R19759 GND.n2288 GND.n2284 9.3005
R19760 GND.n3892 GND.n2289 9.3005
R19761 GND.n3891 GND.n2290 9.3005
R19762 GND.n3890 GND.n2291 9.3005
R19763 GND.n2296 GND.n2292 9.3005
R19764 GND.n3884 GND.n2297 9.3005
R19765 GND.n3883 GND.n2298 9.3005
R19766 GND.n3882 GND.n2299 9.3005
R19767 GND.n2304 GND.n2300 9.3005
R19768 GND.n3876 GND.n2305 9.3005
R19769 GND.n3875 GND.n2306 9.3005
R19770 GND.n3874 GND.n2307 9.3005
R19771 GND.n2312 GND.n2308 9.3005
R19772 GND.n3868 GND.n2313 9.3005
R19773 GND.n3867 GND.n2314 9.3005
R19774 GND.n3866 GND.n2315 9.3005
R19775 GND.n2320 GND.n2316 9.3005
R19776 GND.n3860 GND.n2321 9.3005
R19777 GND.n3859 GND.n2322 9.3005
R19778 GND.n3858 GND.n2323 9.3005
R19779 GND.n2328 GND.n2324 9.3005
R19780 GND.n3852 GND.n2329 9.3005
R19781 GND.n3851 GND.n2330 9.3005
R19782 GND.n3850 GND.n2331 9.3005
R19783 GND.n2336 GND.n2332 9.3005
R19784 GND.n3844 GND.n2337 9.3005
R19785 GND.n3843 GND.n2338 9.3005
R19786 GND.n3842 GND.n2339 9.3005
R19787 GND.n2344 GND.n2340 9.3005
R19788 GND.n3836 GND.n2345 9.3005
R19789 GND.n3835 GND.n2346 9.3005
R19790 GND.n3834 GND.n2347 9.3005
R19791 GND.n2352 GND.n2348 9.3005
R19792 GND.n3828 GND.n2353 9.3005
R19793 GND.n3827 GND.n2354 9.3005
R19794 GND.n3826 GND.n2355 9.3005
R19795 GND.n2360 GND.n2356 9.3005
R19796 GND.n3820 GND.n2361 9.3005
R19797 GND.n3819 GND.n2362 9.3005
R19798 GND.n3818 GND.n2363 9.3005
R19799 GND.n2368 GND.n2364 9.3005
R19800 GND.n3812 GND.n2369 9.3005
R19801 GND.n3811 GND.n2370 9.3005
R19802 GND.n3810 GND.n2371 9.3005
R19803 GND.n2376 GND.n2372 9.3005
R19804 GND.n3804 GND.n2377 9.3005
R19805 GND.n3803 GND.n2378 9.3005
R19806 GND.n3802 GND.n2379 9.3005
R19807 GND.n2384 GND.n2380 9.3005
R19808 GND.n3796 GND.n2385 9.3005
R19809 GND.n3795 GND.n2386 9.3005
R19810 GND.n3794 GND.n2387 9.3005
R19811 GND.n2392 GND.n2388 9.3005
R19812 GND.n3788 GND.n2393 9.3005
R19813 GND.n3787 GND.n2394 9.3005
R19814 GND.n3786 GND.n2395 9.3005
R19815 GND.n2400 GND.n2396 9.3005
R19816 GND.n3780 GND.n2401 9.3005
R19817 GND.n3779 GND.n2402 9.3005
R19818 GND.n3778 GND.n2403 9.3005
R19819 GND.n2408 GND.n2404 9.3005
R19820 GND.n3772 GND.n2409 9.3005
R19821 GND.n3771 GND.n2410 9.3005
R19822 GND.n3770 GND.n2411 9.3005
R19823 GND.n2416 GND.n2412 9.3005
R19824 GND.n3764 GND.n2417 9.3005
R19825 GND.n3763 GND.n2418 9.3005
R19826 GND.n3762 GND.n2419 9.3005
R19827 GND.n2424 GND.n2420 9.3005
R19828 GND.n3756 GND.n2425 9.3005
R19829 GND.n3755 GND.n2426 9.3005
R19830 GND.n3754 GND.n2427 9.3005
R19831 GND.n2432 GND.n2428 9.3005
R19832 GND.n3748 GND.n2433 9.3005
R19833 GND.n3747 GND.n2434 9.3005
R19834 GND.n3746 GND.n2435 9.3005
R19835 GND.n2440 GND.n2436 9.3005
R19836 GND.n3740 GND.n2441 9.3005
R19837 GND.n3739 GND.n2442 9.3005
R19838 GND.n3738 GND.n2443 9.3005
R19839 GND.n2448 GND.n2444 9.3005
R19840 GND.n3732 GND.n2449 9.3005
R19841 GND.n3731 GND.n2450 9.3005
R19842 GND.n3730 GND.n2451 9.3005
R19843 GND.n2456 GND.n2452 9.3005
R19844 GND.n3724 GND.n2457 9.3005
R19845 GND.n3723 GND.n2458 9.3005
R19846 GND.n3722 GND.n2459 9.3005
R19847 GND.n2464 GND.n2460 9.3005
R19848 GND.n3716 GND.n2465 9.3005
R19849 GND.n3715 GND.n2466 9.3005
R19850 GND.n3714 GND.n2467 9.3005
R19851 GND.n2472 GND.n2468 9.3005
R19852 GND.n3708 GND.n2473 9.3005
R19853 GND.n3707 GND.n2474 9.3005
R19854 GND.n3706 GND.n2475 9.3005
R19855 GND.n2480 GND.n2476 9.3005
R19856 GND.n3700 GND.n2481 9.3005
R19857 GND.n3699 GND.n2482 9.3005
R19858 GND.n3698 GND.n2483 9.3005
R19859 GND.n2488 GND.n2484 9.3005
R19860 GND.n3692 GND.n2489 9.3005
R19861 GND.n3691 GND.n2490 9.3005
R19862 GND.n3690 GND.n2491 9.3005
R19863 GND.n2496 GND.n2492 9.3005
R19864 GND.n3684 GND.n2497 9.3005
R19865 GND.n3683 GND.n2498 9.3005
R19866 GND.n3682 GND.n2499 9.3005
R19867 GND.n2504 GND.n2500 9.3005
R19868 GND.n3676 GND.n2505 9.3005
R19869 GND.n3675 GND.n2506 9.3005
R19870 GND.n3674 GND.n2507 9.3005
R19871 GND.n2512 GND.n2508 9.3005
R19872 GND.n3668 GND.n2513 9.3005
R19873 GND.n3667 GND.n2514 9.3005
R19874 GND.n3666 GND.n2515 9.3005
R19875 GND.n2520 GND.n2516 9.3005
R19876 GND.n3660 GND.n2521 9.3005
R19877 GND.n3659 GND.n2522 9.3005
R19878 GND.n3658 GND.n2523 9.3005
R19879 GND.n2528 GND.n2524 9.3005
R19880 GND.n3652 GND.n2529 9.3005
R19881 GND.n3651 GND.n2530 9.3005
R19882 GND.n3650 GND.n2531 9.3005
R19883 GND.n2536 GND.n2532 9.3005
R19884 GND.n3644 GND.n2537 9.3005
R19885 GND.n3643 GND.n2538 9.3005
R19886 GND.n3642 GND.n2539 9.3005
R19887 GND.n2544 GND.n2540 9.3005
R19888 GND.n3636 GND.n2545 9.3005
R19889 GND.n3635 GND.n2546 9.3005
R19890 GND.n3634 GND.n2547 9.3005
R19891 GND.n2552 GND.n2548 9.3005
R19892 GND.n3628 GND.n2553 9.3005
R19893 GND.n3627 GND.n2554 9.3005
R19894 GND.n3626 GND.n2555 9.3005
R19895 GND.n2560 GND.n2556 9.3005
R19896 GND.n3620 GND.n2561 9.3005
R19897 GND.n3619 GND.n2562 9.3005
R19898 GND.n3618 GND.n2563 9.3005
R19899 GND.n2568 GND.n2564 9.3005
R19900 GND.n3612 GND.n2569 9.3005
R19901 GND.n3611 GND.n2570 9.3005
R19902 GND.n3610 GND.n2571 9.3005
R19903 GND.n2576 GND.n2572 9.3005
R19904 GND.n3604 GND.n2577 9.3005
R19905 GND.n3603 GND.n2578 9.3005
R19906 GND.n3602 GND.n2579 9.3005
R19907 GND.n2584 GND.n2580 9.3005
R19908 GND.n3596 GND.n2585 9.3005
R19909 GND.n3595 GND.n2586 9.3005
R19910 GND.n3594 GND.n2587 9.3005
R19911 GND.n2592 GND.n2588 9.3005
R19912 GND.n3588 GND.n2593 9.3005
R19913 GND.n3587 GND.n2594 9.3005
R19914 GND.n3586 GND.n2595 9.3005
R19915 GND.n2600 GND.n2596 9.3005
R19916 GND.n3580 GND.n2601 9.3005
R19917 GND.n3579 GND.n2602 9.3005
R19918 GND.n3578 GND.n2603 9.3005
R19919 GND.n2608 GND.n2604 9.3005
R19920 GND.n3572 GND.n2609 9.3005
R19921 GND.n3571 GND.n2610 9.3005
R19922 GND.n3570 GND.n2611 9.3005
R19923 GND.n2616 GND.n2612 9.3005
R19924 GND.n3564 GND.n2617 9.3005
R19925 GND.n3563 GND.n2618 9.3005
R19926 GND.n3562 GND.n2619 9.3005
R19927 GND.n2624 GND.n2620 9.3005
R19928 GND.n3556 GND.n2625 9.3005
R19929 GND.n3555 GND.n2626 9.3005
R19930 GND.n3554 GND.n2627 9.3005
R19931 GND.n2632 GND.n2628 9.3005
R19932 GND.n3548 GND.n2633 9.3005
R19933 GND.n3547 GND.n2634 9.3005
R19934 GND.n3546 GND.n2635 9.3005
R19935 GND.n2640 GND.n2636 9.3005
R19936 GND.n3540 GND.n2641 9.3005
R19937 GND.n3539 GND.n2642 9.3005
R19938 GND.n3538 GND.n2643 9.3005
R19939 GND.n2648 GND.n2644 9.3005
R19940 GND.n3532 GND.n2649 9.3005
R19941 GND.n3531 GND.n2650 9.3005
R19942 GND.n3530 GND.n2651 9.3005
R19943 GND.n2656 GND.n2652 9.3005
R19944 GND.n3524 GND.n2657 9.3005
R19945 GND.n3523 GND.n2658 9.3005
R19946 GND.n3522 GND.n2659 9.3005
R19947 GND.n2664 GND.n2660 9.3005
R19948 GND.n3516 GND.n2665 9.3005
R19949 GND.n3515 GND.n2666 9.3005
R19950 GND.n3514 GND.n2667 9.3005
R19951 GND.n2672 GND.n2668 9.3005
R19952 GND.n3508 GND.n2673 9.3005
R19953 GND.n3507 GND.n2674 9.3005
R19954 GND.n3506 GND.n2675 9.3005
R19955 GND.n2680 GND.n2676 9.3005
R19956 GND.n3500 GND.n2681 9.3005
R19957 GND.n3499 GND.n2682 9.3005
R19958 GND.n3498 GND.n2683 9.3005
R19959 GND.n2688 GND.n2684 9.3005
R19960 GND.n3492 GND.n2689 9.3005
R19961 GND.n3491 GND.n2690 9.3005
R19962 GND.n3490 GND.n2691 9.3005
R19963 GND.n2696 GND.n2692 9.3005
R19964 GND.n3484 GND.n2697 9.3005
R19965 GND.n3483 GND.n2698 9.3005
R19966 GND.n3482 GND.n2699 9.3005
R19967 GND.n2704 GND.n2700 9.3005
R19968 GND.n3476 GND.n2705 9.3005
R19969 GND.n3475 GND.n2706 9.3005
R19970 GND.n3474 GND.n2707 9.3005
R19971 GND.n2712 GND.n2708 9.3005
R19972 GND.n3468 GND.n2713 9.3005
R19973 GND.n3467 GND.n2714 9.3005
R19974 GND.n3466 GND.n2715 9.3005
R19975 GND.n2720 GND.n2716 9.3005
R19976 GND.n3460 GND.n2721 9.3005
R19977 GND.n3459 GND.n2722 9.3005
R19978 GND.n3458 GND.n2723 9.3005
R19979 GND.n2728 GND.n2724 9.3005
R19980 GND.n3452 GND.n2729 9.3005
R19981 GND.n3451 GND.n2730 9.3005
R19982 GND.n3450 GND.n2731 9.3005
R19983 GND.n2736 GND.n2732 9.3005
R19984 GND.n3444 GND.n2737 9.3005
R19985 GND.n3443 GND.n2738 9.3005
R19986 GND.n3442 GND.n2739 9.3005
R19987 GND.n2744 GND.n2740 9.3005
R19988 GND.n3436 GND.n2745 9.3005
R19989 GND.n3435 GND.n2746 9.3005
R19990 GND.n3434 GND.n2747 9.3005
R19991 GND.n2752 GND.n2748 9.3005
R19992 GND.n3428 GND.n2753 9.3005
R19993 GND.n3427 GND.n2754 9.3005
R19994 GND.n3426 GND.n2755 9.3005
R19995 GND.n2760 GND.n2756 9.3005
R19996 GND.n3420 GND.n2761 9.3005
R19997 GND.n3419 GND.n2762 9.3005
R19998 GND.n3418 GND.n2763 9.3005
R19999 GND.n2768 GND.n2764 9.3005
R20000 GND.n3412 GND.n2769 9.3005
R20001 GND.n3411 GND.n2770 9.3005
R20002 GND.n3410 GND.n2771 9.3005
R20003 GND.n2776 GND.n2772 9.3005
R20004 GND.n3404 GND.n2777 9.3005
R20005 GND.n3403 GND.n2778 9.3005
R20006 GND.n3402 GND.n2779 9.3005
R20007 GND.n2784 GND.n2780 9.3005
R20008 GND.n3396 GND.n2785 9.3005
R20009 GND.n3395 GND.n2786 9.3005
R20010 GND.n3394 GND.n2787 9.3005
R20011 GND.n2792 GND.n2788 9.3005
R20012 GND.n3388 GND.n2793 9.3005
R20013 GND.n3387 GND.n2794 9.3005
R20014 GND.n3386 GND.n2795 9.3005
R20015 GND.n2800 GND.n2796 9.3005
R20016 GND.n3380 GND.n2801 9.3005
R20017 GND.n3379 GND.n2802 9.3005
R20018 GND.n3378 GND.n2803 9.3005
R20019 GND.n2808 GND.n2804 9.3005
R20020 GND.n3372 GND.n2809 9.3005
R20021 GND.n3371 GND.n2810 9.3005
R20022 GND.n3370 GND.n2811 9.3005
R20023 GND.n2816 GND.n2812 9.3005
R20024 GND.n3364 GND.n2817 9.3005
R20025 GND.n3363 GND.n2818 9.3005
R20026 GND.n3362 GND.n2819 9.3005
R20027 GND.n2824 GND.n2820 9.3005
R20028 GND.n3356 GND.n2825 9.3005
R20029 GND.n3355 GND.n2826 9.3005
R20030 GND.n3354 GND.n2827 9.3005
R20031 GND.n2832 GND.n2828 9.3005
R20032 GND.n3348 GND.n2833 9.3005
R20033 GND.n3347 GND.n2834 9.3005
R20034 GND.n3346 GND.n2835 9.3005
R20035 GND.n2840 GND.n2836 9.3005
R20036 GND.n3340 GND.n2841 9.3005
R20037 GND.n3339 GND.n2842 9.3005
R20038 GND.n3338 GND.n2843 9.3005
R20039 GND.n2848 GND.n2844 9.3005
R20040 GND.n3332 GND.n2849 9.3005
R20041 GND.n3331 GND.n2850 9.3005
R20042 GND.n3330 GND.n2851 9.3005
R20043 GND.n2856 GND.n2852 9.3005
R20044 GND.n3324 GND.n2857 9.3005
R20045 GND.n3323 GND.n2858 9.3005
R20046 GND.n3322 GND.n2859 9.3005
R20047 GND.n2864 GND.n2860 9.3005
R20048 GND.n3316 GND.n2865 9.3005
R20049 GND.n3315 GND.n2866 9.3005
R20050 GND.n3314 GND.n2867 9.3005
R20051 GND.n2872 GND.n2868 9.3005
R20052 GND.n3308 GND.n2873 9.3005
R20053 GND.n3307 GND.n2874 9.3005
R20054 GND.n3306 GND.n2875 9.3005
R20055 GND.n2880 GND.n2876 9.3005
R20056 GND.n3300 GND.n2881 9.3005
R20057 GND.n3299 GND.n2882 9.3005
R20058 GND.n3298 GND.n2883 9.3005
R20059 GND.n2888 GND.n2884 9.3005
R20060 GND.n3292 GND.n2889 9.3005
R20061 GND.n3291 GND.n2890 9.3005
R20062 GND.n3290 GND.n2891 9.3005
R20063 GND.n2896 GND.n2892 9.3005
R20064 GND.n3284 GND.n2897 9.3005
R20065 GND.n3283 GND.n2898 9.3005
R20066 GND.n3282 GND.n2899 9.3005
R20067 GND.n2904 GND.n2900 9.3005
R20068 GND.n3276 GND.n2905 9.3005
R20069 GND.n3275 GND.n2906 9.3005
R20070 GND.n3274 GND.n2907 9.3005
R20071 GND.n2912 GND.n2908 9.3005
R20072 GND.n3268 GND.n2913 9.3005
R20073 GND.n3267 GND.n2914 9.3005
R20074 GND.n3266 GND.n2915 9.3005
R20075 GND.n2920 GND.n2916 9.3005
R20076 GND.n3260 GND.n2921 9.3005
R20077 GND.n3259 GND.n2922 9.3005
R20078 GND.n3258 GND.n2923 9.3005
R20079 GND.n2928 GND.n2924 9.3005
R20080 GND.n3252 GND.n2929 9.3005
R20081 GND.n3251 GND.n2930 9.3005
R20082 GND.n3250 GND.n2931 9.3005
R20083 GND.n2936 GND.n2932 9.3005
R20084 GND.n3244 GND.n2937 9.3005
R20085 GND.n3243 GND.n2938 9.3005
R20086 GND.n3242 GND.n2939 9.3005
R20087 GND.n2944 GND.n2940 9.3005
R20088 GND.n3236 GND.n2945 9.3005
R20089 GND.n3235 GND.n2946 9.3005
R20090 GND.n3234 GND.n2947 9.3005
R20091 GND.n2952 GND.n2948 9.3005
R20092 GND.n3228 GND.n2953 9.3005
R20093 GND.n3227 GND.n2954 9.3005
R20094 GND.n3226 GND.n2955 9.3005
R20095 GND.n2960 GND.n2956 9.3005
R20096 GND.n3220 GND.n2961 9.3005
R20097 GND.n3219 GND.n2962 9.3005
R20098 GND.n3218 GND.n2963 9.3005
R20099 GND.n2968 GND.n2964 9.3005
R20100 GND.n3211 GND.n3210 9.3005
R20101 GND.n3209 GND.n2970 9.3005
R20102 GND.n3208 GND.n3207 9.3005
R20103 GND.n2972 GND.n2971 9.3005
R20104 GND.n3201 GND.n2978 9.3005
R20105 GND.n3200 GND.n2979 9.3005
R20106 GND.n3199 GND.n2980 9.3005
R20107 GND.n2985 GND.n2981 9.3005
R20108 GND.n3193 GND.n2986 9.3005
R20109 GND.n3192 GND.n2987 9.3005
R20110 GND.n3191 GND.n2988 9.3005
R20111 GND.n2993 GND.n2989 9.3005
R20112 GND.n3185 GND.n2994 9.3005
R20113 GND.n3184 GND.n2995 9.3005
R20114 GND.n3183 GND.n2996 9.3005
R20115 GND.n3001 GND.n2997 9.3005
R20116 GND.n3177 GND.n3002 9.3005
R20117 GND.n3176 GND.n3003 9.3005
R20118 GND.n3175 GND.n3004 9.3005
R20119 GND.n3009 GND.n3005 9.3005
R20120 GND.n3169 GND.n3010 9.3005
R20121 GND.n3168 GND.n3011 9.3005
R20122 GND.n3167 GND.n3012 9.3005
R20123 GND.n3017 GND.n3013 9.3005
R20124 GND.n3161 GND.n3018 9.3005
R20125 GND.n3160 GND.n3019 9.3005
R20126 GND.n3159 GND.n3020 9.3005
R20127 GND.n3025 GND.n3021 9.3005
R20128 GND.n3153 GND.n3026 9.3005
R20129 GND.n3152 GND.n3027 9.3005
R20130 GND.n3151 GND.n3028 9.3005
R20131 GND.n3033 GND.n3029 9.3005
R20132 GND.n3145 GND.n3034 9.3005
R20133 GND.n3144 GND.n3035 9.3005
R20134 GND.n3143 GND.n3036 9.3005
R20135 GND.n3041 GND.n3037 9.3005
R20136 GND.n3137 GND.n3042 9.3005
R20137 GND.n3136 GND.n3043 9.3005
R20138 GND.n3135 GND.n3044 9.3005
R20139 GND.n3049 GND.n3045 9.3005
R20140 GND.n3129 GND.n3050 9.3005
R20141 GND.n3128 GND.n3051 9.3005
R20142 GND.n3127 GND.n3052 9.3005
R20143 GND.n3057 GND.n3053 9.3005
R20144 GND.n3121 GND.n3058 9.3005
R20145 GND.n3120 GND.n3059 9.3005
R20146 GND.n3119 GND.n3060 9.3005
R20147 GND.n3065 GND.n3061 9.3005
R20148 GND.n3113 GND.n3066 9.3005
R20149 GND.n3112 GND.n3067 9.3005
R20150 GND.n3111 GND.n3068 9.3005
R20151 GND.n3073 GND.n3069 9.3005
R20152 GND.n3105 GND.n3074 9.3005
R20153 GND.n3104 GND.n3075 9.3005
R20154 GND.n3103 GND.n3076 9.3005
R20155 GND.n3081 GND.n3077 9.3005
R20156 GND.n3097 GND.n3082 9.3005
R20157 GND.n3096 GND.n3083 9.3005
R20158 GND.n3095 GND.n3084 9.3005
R20159 GND.n3087 GND.n3085 9.3005
R20160 GND.n3089 GND.n3088 9.3005
R20161 GND.n385 GND.n384 9.3005
R20162 GND.n8263 GND.n8262 9.3005
R20163 GND.n3212 GND.n2969 9.3005
R20164 GND.n89 GND.n88 9.3005
R20165 GND.n100 GND.n99 9.3005
R20166 GND.n112 GND.n111 9.3005
R20167 GND.n124 GND.n123 9.3005
R20168 GND.n136 GND.n135 9.3005
R20169 GND.n148 GND.n147 9.3005
R20170 GND.n5596 GND.n5595 9.3005
R20171 GND.n5597 GND.n5591 9.3005
R20172 GND.n5601 GND.n5600 9.3005
R20173 GND.n5602 GND.n5590 9.3005
R20174 GND.n5621 GND.n5603 9.3005
R20175 GND.n5620 GND.n5604 9.3005
R20176 GND.n5619 GND.n5605 9.3005
R20177 GND.n5617 GND.n5606 9.3005
R20178 GND.n5616 GND.n5607 9.3005
R20179 GND.n5614 GND.n5608 9.3005
R20180 GND.n5613 GND.n5610 9.3005
R20181 GND.n5609 GND.n1513 9.3005
R20182 GND.n6310 GND.n1514 9.3005
R20183 GND.n6309 GND.n1515 9.3005
R20184 GND.n6308 GND.n1516 9.3005
R20185 GND.n6211 GND.n1517 9.3005
R20186 GND.n6214 GND.n6213 9.3005
R20187 GND.n6215 GND.n6210 9.3005
R20188 GND.n6218 GND.n6216 9.3005
R20189 GND.n6219 GND.n6209 9.3005
R20190 GND.n6222 GND.n6221 9.3005
R20191 GND.n6223 GND.n6208 9.3005
R20192 GND.n6226 GND.n6224 9.3005
R20193 GND.n6227 GND.n6207 9.3005
R20194 GND.n6230 GND.n6229 9.3005
R20195 GND.n6231 GND.n6206 9.3005
R20196 GND.n6235 GND.n6232 9.3005
R20197 GND.n6234 GND.n6233 9.3005
R20198 GND.n1420 GND.n1419 9.3005
R20199 GND.n6407 GND.n6406 9.3005
R20200 GND.n6408 GND.n1418 9.3005
R20201 GND.n6411 GND.n6409 9.3005
R20202 GND.n6412 GND.n1417 9.3005
R20203 GND.n6415 GND.n6414 9.3005
R20204 GND.n6416 GND.n1416 9.3005
R20205 GND.n6419 GND.n6417 9.3005
R20206 GND.n6420 GND.n1415 9.3005
R20207 GND.n6423 GND.n6422 9.3005
R20208 GND.n6424 GND.n1414 9.3005
R20209 GND.n6427 GND.n6425 9.3005
R20210 GND.n6428 GND.n1413 9.3005
R20211 GND.n6431 GND.n6430 9.3005
R20212 GND.n6432 GND.n1412 9.3005
R20213 GND.n6435 GND.n6433 9.3005
R20214 GND.n6436 GND.n1411 9.3005
R20215 GND.n6439 GND.n6438 9.3005
R20216 GND.n6440 GND.n1410 9.3005
R20217 GND.n6443 GND.n6441 9.3005
R20218 GND.n6444 GND.n1409 9.3005
R20219 GND.n6448 GND.n6447 9.3005
R20220 GND.n6449 GND.n1408 9.3005
R20221 GND.n6473 GND.n6450 9.3005
R20222 GND.n6472 GND.n6451 9.3005
R20223 GND.n6471 GND.n6452 9.3005
R20224 GND.n6469 GND.n6453 9.3005
R20225 GND.n6468 GND.n6454 9.3005
R20226 GND.n6466 GND.n6455 9.3005
R20227 GND.n6465 GND.n6456 9.3005
R20228 GND.n6463 GND.n6457 9.3005
R20229 GND.n6462 GND.n6459 9.3005
R20230 GND.n6458 GND.n1178 9.3005
R20231 GND.n6807 GND.n1179 9.3005
R20232 GND.n6806 GND.n1180 9.3005
R20233 GND.n6805 GND.n1181 9.3005
R20234 GND.n1191 GND.n1182 9.3005
R20235 GND.n6793 GND.n1192 9.3005
R20236 GND.n6792 GND.n1193 9.3005
R20237 GND.n6791 GND.n1194 9.3005
R20238 GND.n6722 GND.n1195 9.3005
R20239 GND.n6725 GND.n6723 9.3005
R20240 GND.n6726 GND.n6721 9.3005
R20241 GND.n6729 GND.n6728 9.3005
R20242 GND.n6730 GND.n6720 9.3005
R20243 GND.n6739 GND.n6731 9.3005
R20244 GND.n6738 GND.n6732 9.3005
R20245 GND.n6737 GND.n6734 9.3005
R20246 GND.n6733 GND.n1085 9.3005
R20247 GND.n6907 GND.n1084 9.3005
R20248 GND.n6909 GND.n6908 9.3005
R20249 GND.n6910 GND.n1083 9.3005
R20250 GND.n6912 GND.n6911 9.3005
R20251 GND.n6914 GND.n1080 9.3005
R20252 GND.n6916 GND.n6915 9.3005
R20253 GND.n5594 GND.n5592 9.3005
R20254 GND.n6089 GND.n1593 9.3005
R20255 GND.n6092 GND.n1592 9.3005
R20256 GND.n6094 GND.n1591 9.3005
R20257 GND.n6095 GND.n1590 9.3005
R20258 GND.n6096 GND.n1589 9.3005
R20259 GND.n6097 GND.n1588 9.3005
R20260 GND.n6069 GND.n6068 9.3005
R20261 GND.n6071 GND.n6065 9.3005
R20262 GND.n6067 GND.n1565 9.3005
R20263 GND.n6113 GND.n1564 9.3005
R20264 GND.n6115 GND.n6114 9.3005
R20265 GND.n1551 GND.n1550 9.3005
R20266 GND.n6128 GND.n6127 9.3005
R20267 GND.n6129 GND.n1549 9.3005
R20268 GND.n6140 GND.n6130 9.3005
R20269 GND.n6139 GND.n6131 9.3005
R20270 GND.n6138 GND.n6132 9.3005
R20271 GND.n6137 GND.n6133 9.3005
R20272 GND.n6135 GND.n6134 9.3005
R20273 GND.n1491 GND.n1490 9.3005
R20274 GND.n6332 GND.n6331 9.3005
R20275 GND.n6333 GND.n1489 9.3005
R20276 GND.n6335 GND.n6334 9.3005
R20277 GND.n1475 GND.n1474 9.3005
R20278 GND.n6348 GND.n6347 9.3005
R20279 GND.n6349 GND.n1473 9.3005
R20280 GND.n6351 GND.n6350 9.3005
R20281 GND.n1459 GND.n1458 9.3005
R20282 GND.n6364 GND.n6363 9.3005
R20283 GND.n6365 GND.n1457 9.3005
R20284 GND.n6367 GND.n6366 9.3005
R20285 GND.n1443 GND.n1442 9.3005
R20286 GND.n6379 GND.n6378 9.3005
R20287 GND.n6380 GND.n1441 9.3005
R20288 GND.n6382 GND.n6381 9.3005
R20289 GND.n1426 GND.n1425 9.3005
R20290 GND.n6397 GND.n6396 9.3005
R20291 GND.n6398 GND.n1424 9.3005
R20292 GND.n6402 GND.n6399 9.3005
R20293 GND.n6401 GND.n6400 9.3005
R20294 GND.n1310 GND.n1309 9.3005
R20295 GND.n6571 GND.n6570 9.3005
R20296 GND.n6572 GND.n1308 9.3005
R20297 GND.n6574 GND.n6573 9.3005
R20298 GND.n1294 GND.n1293 9.3005
R20299 GND.n6587 GND.n6586 9.3005
R20300 GND.n6588 GND.n1292 9.3005
R20301 GND.n6590 GND.n6589 9.3005
R20302 GND.n1278 GND.n1277 9.3005
R20303 GND.n6603 GND.n6602 9.3005
R20304 GND.n6604 GND.n1276 9.3005
R20305 GND.n6606 GND.n6605 9.3005
R20306 GND.n1262 GND.n1261 9.3005
R20307 GND.n6618 GND.n6617 9.3005
R20308 GND.n6619 GND.n1260 9.3005
R20309 GND.n6621 GND.n6620 9.3005
R20310 GND.n1246 GND.n1245 9.3005
R20311 GND.n6634 GND.n6633 9.3005
R20312 GND.n6635 GND.n1244 9.3005
R20313 GND.n6637 GND.n6636 9.3005
R20314 GND.n1230 GND.n1229 9.3005
R20315 GND.n6650 GND.n6649 9.3005
R20316 GND.n6651 GND.n1228 9.3005
R20317 GND.n6662 GND.n6652 9.3005
R20318 GND.n6661 GND.n6653 9.3005
R20319 GND.n6660 GND.n6654 9.3005
R20320 GND.n6659 GND.n6655 9.3005
R20321 GND.n6657 GND.n6656 9.3005
R20322 GND.n1156 GND.n1155 9.3005
R20323 GND.n6829 GND.n6828 9.3005
R20324 GND.n6830 GND.n1154 9.3005
R20325 GND.n6832 GND.n6831 9.3005
R20326 GND.n1140 GND.n1139 9.3005
R20327 GND.n6845 GND.n6844 9.3005
R20328 GND.n6846 GND.n1138 9.3005
R20329 GND.n6848 GND.n6847 9.3005
R20330 GND.n1124 GND.n1123 9.3005
R20331 GND.n6861 GND.n6860 9.3005
R20332 GND.n6862 GND.n1122 9.3005
R20333 GND.n6864 GND.n6863 9.3005
R20334 GND.n1108 GND.n1107 9.3005
R20335 GND.n6876 GND.n6875 9.3005
R20336 GND.n6877 GND.n1106 9.3005
R20337 GND.n6884 GND.n6878 9.3005
R20338 GND.n6883 GND.n6879 9.3005
R20339 GND.n6882 GND.n6881 9.3005
R20340 GND.n6880 GND.n1060 9.3005
R20341 GND.n6977 GND.n1061 9.3005
R20342 GND.n6976 GND.n1062 9.3005
R20343 GND.n6975 GND.n1063 9.3005
R20344 GND.n6974 GND.n1064 9.3005
R20345 GND.n6968 GND.n1065 9.3005
R20346 GND.n6112 GND.n6111 9.3005
R20347 GND.n6966 GND.n6965 9.3005
R20348 GND.n6967 GND.n1067 9.3005
R20349 GND.n6970 GND.n6969 9.3005
R20350 GND.n1078 GND.n1077 9.3005
R20351 GND.n6925 GND.n6924 9.3005
R20352 GND.n6926 GND.n1076 9.3005
R20353 GND.n6929 GND.n6928 9.3005
R20354 GND.n6927 GND.n1074 9.3005
R20355 GND.n6918 GND.n6917 9.3005
R20356 GND.n7731 GND.n664 9.3005
R20357 GND.n1068 GND.n661 9.3005
R20358 GND.n7734 GND.n7733 9.3005
R20359 GND.n635 GND.n634 9.3005
R20360 GND.n7767 GND.n7766 9.3005
R20361 GND.n7768 GND.n633 9.3005
R20362 GND.n7772 GND.n7769 9.3005
R20363 GND.n7771 GND.n7770 9.3005
R20364 GND.n607 GND.n606 9.3005
R20365 GND.n7804 GND.n7803 9.3005
R20366 GND.n7805 GND.n605 9.3005
R20367 GND.n7813 GND.n7806 9.3005
R20368 GND.n7812 GND.n7807 9.3005
R20369 GND.n7811 GND.n7808 9.3005
R20370 GND.n580 GND.n579 9.3005
R20371 GND.n7840 GND.n7839 9.3005
R20372 GND.n7841 GND.n578 9.3005
R20373 GND.n7844 GND.n7843 9.3005
R20374 GND.n7842 GND.n555 9.3005
R20375 GND.n7871 GND.n556 9.3005
R20376 GND.n7872 GND.n554 9.3005
R20377 GND.n7875 GND.n7874 9.3005
R20378 GND.n7876 GND.n553 9.3005
R20379 GND.n7880 GND.n7877 9.3005
R20380 GND.n7879 GND.n7878 9.3005
R20381 GND.n493 GND.n492 9.3005
R20382 GND.n7957 GND.n7956 9.3005
R20383 GND.n7958 GND.n491 9.3005
R20384 GND.n7962 GND.n7959 9.3005
R20385 GND.n7961 GND.n7960 9.3005
R20386 GND.n466 GND.n465 9.3005
R20387 GND.n7994 GND.n7993 9.3005
R20388 GND.n7995 GND.n464 9.3005
R20389 GND.n8004 GND.n7996 9.3005
R20390 GND.n8003 GND.n7997 9.3005
R20391 GND.n8002 GND.n7998 9.3005
R20392 GND.n8001 GND.n7999 9.3005
R20393 GND.n154 GND.n152 9.3005
R20394 GND.n7735 GND.n7732 9.3005
R20395 GND.n8569 GND.n8568 9.3005
R20396 GND.n155 GND.n153 9.3005
R20397 GND.n427 GND.n426 9.3005
R20398 GND.n8135 GND.n8134 9.3005
R20399 GND.n8136 GND.n425 9.3005
R20400 GND.n8138 GND.n8137 9.3005
R20401 GND.n423 GND.n422 9.3005
R20402 GND.n8150 GND.n8149 9.3005
R20403 GND.n8151 GND.n421 9.3005
R20404 GND.n8153 GND.n8152 9.3005
R20405 GND.n419 GND.n418 9.3005
R20406 GND.n8165 GND.n8164 9.3005
R20407 GND.n8166 GND.n417 9.3005
R20408 GND.n8168 GND.n8167 9.3005
R20409 GND.n415 GND.n414 9.3005
R20410 GND.n8180 GND.n8179 9.3005
R20411 GND.n8181 GND.n413 9.3005
R20412 GND.n8183 GND.n8182 9.3005
R20413 GND.n410 GND.n409 9.3005
R20414 GND.n8195 GND.n8194 9.3005
R20415 GND.n8196 GND.n408 9.3005
R20416 GND.n8198 GND.n8197 9.3005
R20417 GND.n406 GND.n405 9.3005
R20418 GND.n8210 GND.n8209 9.3005
R20419 GND.n8211 GND.n404 9.3005
R20420 GND.n8213 GND.n8212 9.3005
R20421 GND.n402 GND.n401 9.3005
R20422 GND.n8225 GND.n8224 9.3005
R20423 GND.n8226 GND.n400 9.3005
R20424 GND.n8229 GND.n8228 9.3005
R20425 GND.n8227 GND.n394 9.3005
R20426 GND.n8244 GND.n395 9.3005
R20427 GND.n8243 GND.n396 9.3005
R20428 GND.n8242 GND.n398 9.3005
R20429 GND.n397 GND.n351 9.3005
R20430 GND.n8454 GND.n352 9.3005
R20431 GND.n8453 GND.n8452 9.3005
R20432 GND.n367 GND.n364 9.3005
R20433 GND.n369 GND.n368 9.3005
R20434 GND.n372 GND.n362 9.3005
R20435 GND.n375 GND.n374 9.3005
R20436 GND.n376 GND.n361 9.3005
R20437 GND.n378 GND.n377 9.3005
R20438 GND.n356 GND.n353 9.3005
R20439 GND.n8451 GND.n8450 9.3005
R20440 GND.n366 GND.n365 9.3005
R20441 GND.n8294 GND.n8291 9.3005
R20442 GND.n8444 GND.n8295 9.3005
R20443 GND.n8443 GND.n8296 9.3005
R20444 GND.n8442 GND.n8297 9.3005
R20445 GND.n8439 GND.n8298 9.3005
R20446 GND.n8438 GND.n8299 9.3005
R20447 GND.n8435 GND.n8300 9.3005
R20448 GND.n8434 GND.n8433 9.3005
R20449 GND.n8432 GND.n8301 9.3005
R20450 GND.n8431 GND.n8430 9.3005
R20451 GND.n8427 GND.n8306 9.3005
R20452 GND.n8426 GND.n8307 9.3005
R20453 GND.n8423 GND.n8308 9.3005
R20454 GND.n8422 GND.n8309 9.3005
R20455 GND.n8419 GND.n8310 9.3005
R20456 GND.n8418 GND.n8311 9.3005
R20457 GND.n8415 GND.n8312 9.3005
R20458 GND.n8411 GND.n8313 9.3005
R20459 GND.n8408 GND.n8314 9.3005
R20460 GND.n8407 GND.n8315 9.3005
R20461 GND.n8404 GND.n8316 9.3005
R20462 GND.n8403 GND.n8317 9.3005
R20463 GND.n8400 GND.n8318 9.3005
R20464 GND.n8399 GND.n8319 9.3005
R20465 GND.n8396 GND.n8320 9.3005
R20466 GND.n8395 GND.n8321 9.3005
R20467 GND.n8392 GND.n8391 9.3005
R20468 GND.n8390 GND.n8322 9.3005
R20469 GND.n8389 GND.n8388 9.3005
R20470 GND.n8385 GND.n8325 9.3005
R20471 GND.n8382 GND.n8326 9.3005
R20472 GND.n8381 GND.n8327 9.3005
R20473 GND.n8378 GND.n8328 9.3005
R20474 GND.n8377 GND.n8329 9.3005
R20475 GND.n8374 GND.n8330 9.3005
R20476 GND.n8373 GND.n8331 9.3005
R20477 GND.n8370 GND.n8369 9.3005
R20478 GND.n8368 GND.n8332 9.3005
R20479 GND.n8367 GND.n8366 9.3005
R20480 GND.n8363 GND.n8335 9.3005
R20481 GND.n8360 GND.n8336 9.3005
R20482 GND.n8359 GND.n8337 9.3005
R20483 GND.n8356 GND.n8338 9.3005
R20484 GND.n8355 GND.n8339 9.3005
R20485 GND.n8352 GND.n8340 9.3005
R20486 GND.n8351 GND.n8341 9.3005
R20487 GND.n8348 GND.n8347 9.3005
R20488 GND.n8346 GND.n8343 9.3005
R20489 GND.n8293 GND.n8292 9.3005
R20490 GND.n7752 GND.n7751 9.3005
R20491 GND.n656 GND.n654 9.3005
R20492 GND.n7745 GND.n7740 9.3005
R20493 GND.n7744 GND.n7743 9.3005
R20494 GND.n629 GND.n625 9.3005
R20495 GND.n7789 GND.n626 9.3005
R20496 GND.n7788 GND.n627 9.3005
R20497 GND.n7787 GND.n7782 9.3005
R20498 GND.n7786 GND.n7783 9.3005
R20499 GND.n601 GND.n598 9.3005
R20500 GND.n7824 GND.n599 9.3005
R20501 GND.n7823 GND.n7820 9.3005
R20502 GND.n7822 GND.n7821 9.3005
R20503 GND.n576 GND.n575 9.3005
R20504 GND.n7851 GND.n7850 9.3005
R20505 GND.n562 GND.n561 9.3005
R20506 GND.n7864 GND.n7863 9.3005
R20507 GND.n7865 GND.n542 9.3005
R20508 GND.n7889 GND.n543 9.3005
R20509 GND.n7888 GND.n544 9.3005
R20510 GND.n7887 GND.n7886 9.3005
R20511 GND.n545 GND.n511 9.3005
R20512 GND.n7942 GND.n512 9.3005
R20513 GND.n7941 GND.n513 9.3005
R20514 GND.n7940 GND.n514 9.3005
R20515 GND.n7939 GND.n515 9.3005
R20516 GND.n488 GND.n484 9.3005
R20517 GND.n7979 GND.n485 9.3005
R20518 GND.n7978 GND.n486 9.3005
R20519 GND.n7977 GND.n7972 9.3005
R20520 GND.n7976 GND.n7973 9.3005
R20521 GND.n459 GND.n458 9.3005
R20522 GND.n8013 GND.n8010 9.3005
R20523 GND.n8012 GND.n8011 9.3005
R20524 GND.n447 GND.n444 9.3005
R20525 GND.n8030 GND.n445 9.3005
R20526 GND.n8029 GND.n8028 9.3005
R20527 GND.n433 GND.n432 9.3005
R20528 GND.n8128 GND.n8127 9.3005
R20529 GND.n8129 GND.n183 9.3005
R20530 GND.n8557 GND.n184 9.3005
R20531 GND.n8556 GND.n185 9.3005
R20532 GND.n8555 GND.n186 9.3005
R20533 GND.n8144 GND.n187 9.3005
R20534 GND.n8545 GND.n204 9.3005
R20535 GND.n8544 GND.n205 9.3005
R20536 GND.n8543 GND.n206 9.3005
R20537 GND.n8159 GND.n207 9.3005
R20538 GND.n8533 GND.n225 9.3005
R20539 GND.n8532 GND.n226 9.3005
R20540 GND.n8531 GND.n227 9.3005
R20541 GND.n8174 GND.n228 9.3005
R20542 GND.n8521 GND.n246 9.3005
R20543 GND.n8520 GND.n247 9.3005
R20544 GND.n8519 GND.n248 9.3005
R20545 GND.n8189 GND.n249 9.3005
R20546 GND.n8509 GND.n266 9.3005
R20547 GND.n8508 GND.n267 9.3005
R20548 GND.n8507 GND.n268 9.3005
R20549 GND.n8204 GND.n269 9.3005
R20550 GND.n8497 GND.n287 9.3005
R20551 GND.n8496 GND.n288 9.3005
R20552 GND.n8495 GND.n289 9.3005
R20553 GND.n8219 GND.n290 9.3005
R20554 GND.n8485 GND.n308 9.3005
R20555 GND.n8484 GND.n309 9.3005
R20556 GND.n8483 GND.n310 9.3005
R20557 GND.n8235 GND.n311 9.3005
R20558 GND.n8473 GND.n328 9.3005
R20559 GND.n8472 GND.n329 9.3005
R20560 GND.n8471 GND.n330 9.3005
R20561 GND.n348 GND.n331 9.3005
R20562 GND.n8461 GND.n8460 9.3005
R20563 GND.n655 GND.n653 9.3005
R20564 GND.n7751 GND.n7750 9.3005
R20565 GND.n7749 GND.n656 9.3005
R20566 GND.n7746 GND.n7745 9.3005
R20567 GND.n7744 GND.n628 9.3005
R20568 GND.n7776 GND.n629 9.3005
R20569 GND.n7777 GND.n626 9.3005
R20570 GND.n7780 GND.n627 9.3005
R20571 GND.n7782 GND.n7781 9.3005
R20572 GND.n7783 GND.n600 9.3005
R20573 GND.n7817 GND.n601 9.3005
R20574 GND.n7818 GND.n599 9.3005
R20575 GND.n7820 GND.n7819 9.3005
R20576 GND.n7821 GND.n584 9.3005
R20577 GND.n577 GND.n576 9.3005
R20578 GND.n7850 GND.n7849 9.3005
R20579 GND.n7848 GND.n561 9.3005
R20580 GND.n7864 GND.n560 9.3005
R20581 GND.n7867 GND.n7865 9.3005
R20582 GND.n7866 GND.n543 9.3005
R20583 GND.n547 GND.n544 9.3005
R20584 GND.n7886 GND.n7885 9.3005
R20585 GND.n7884 GND.n545 9.3005
R20586 GND.n552 GND.n512 9.3005
R20587 GND.n551 GND.n513 9.3005
R20588 GND.n548 GND.n514 9.3005
R20589 GND.n515 GND.n487 9.3005
R20590 GND.n7966 GND.n488 9.3005
R20591 GND.n7967 GND.n485 9.3005
R20592 GND.n7970 GND.n486 9.3005
R20593 GND.n7972 GND.n7971 9.3005
R20594 GND.n7973 GND.n460 9.3005
R20595 GND.n8008 GND.n459 9.3005
R20596 GND.n8010 GND.n8009 9.3005
R20597 GND.n8011 GND.n446 9.3005
R20598 GND.n8023 GND.n447 9.3005
R20599 GND.n8024 GND.n445 9.3005
R20600 GND.n8028 GND.n8027 9.3005
R20601 GND.n8026 GND.n432 9.3005
R20602 GND.n8128 GND.n431 9.3005
R20603 GND.n8130 GND.n8129 9.3005
R20604 GND.n424 GND.n184 9.3005
R20605 GND.n8142 GND.n185 9.3005
R20606 GND.n8143 GND.n186 9.3005
R20607 GND.n8145 GND.n8144 9.3005
R20608 GND.n420 GND.n204 9.3005
R20609 GND.n8157 GND.n205 9.3005
R20610 GND.n8158 GND.n206 9.3005
R20611 GND.n8160 GND.n8159 9.3005
R20612 GND.n416 GND.n225 9.3005
R20613 GND.n8172 GND.n226 9.3005
R20614 GND.n8173 GND.n227 9.3005
R20615 GND.n8175 GND.n8174 9.3005
R20616 GND.n412 GND.n246 9.3005
R20617 GND.n8187 GND.n247 9.3005
R20618 GND.n8188 GND.n248 9.3005
R20619 GND.n8190 GND.n8189 9.3005
R20620 GND.n407 GND.n266 9.3005
R20621 GND.n8202 GND.n267 9.3005
R20622 GND.n8203 GND.n268 9.3005
R20623 GND.n8205 GND.n8204 9.3005
R20624 GND.n403 GND.n287 9.3005
R20625 GND.n8217 GND.n288 9.3005
R20626 GND.n8218 GND.n289 9.3005
R20627 GND.n8220 GND.n8219 9.3005
R20628 GND.n399 GND.n308 9.3005
R20629 GND.n8233 GND.n309 9.3005
R20630 GND.n8234 GND.n310 9.3005
R20631 GND.n8236 GND.n8235 9.3005
R20632 GND.n8237 GND.n328 9.3005
R20633 GND.n8238 GND.n329 9.3005
R20634 GND.n350 GND.n330 9.3005
R20635 GND.n8458 GND.n348 9.3005
R20636 GND.n8460 GND.n8459 9.3005
R20637 GND.n7739 GND.n655 9.3005
R20638 GND.n7632 GND.n7631 9.3005
R20639 GND.n7635 GND.n7626 9.3005
R20640 GND.n7636 GND.n7625 9.3005
R20641 GND.n7639 GND.n7624 9.3005
R20642 GND.n7640 GND.n7623 9.3005
R20643 GND.n7643 GND.n7622 9.3005
R20644 GND.n7644 GND.n7621 9.3005
R20645 GND.n7647 GND.n7620 9.3005
R20646 GND.n7648 GND.n7619 9.3005
R20647 GND.n7651 GND.n7618 9.3005
R20648 GND.n7652 GND.n7615 9.3005
R20649 GND.n7655 GND.n7614 9.3005
R20650 GND.n7656 GND.n7613 9.3005
R20651 GND.n7659 GND.n7612 9.3005
R20652 GND.n7660 GND.n7611 9.3005
R20653 GND.n7663 GND.n7610 9.3005
R20654 GND.n7664 GND.n7609 9.3005
R20655 GND.n7667 GND.n7608 9.3005
R20656 GND.n7668 GND.n7607 9.3005
R20657 GND.n7671 GND.n7606 9.3005
R20658 GND.n7675 GND.n7602 9.3005
R20659 GND.n7676 GND.n7601 9.3005
R20660 GND.n7679 GND.n7600 9.3005
R20661 GND.n7681 GND.n7599 9.3005
R20662 GND.n7685 GND.n734 9.3005
R20663 GND.n7686 GND.n733 9.3005
R20664 GND.n7689 GND.n732 9.3005
R20665 GND.n7691 GND.n729 9.3005
R20666 GND.n7694 GND.n728 9.3005
R20667 GND.n7695 GND.n727 9.3005
R20668 GND.n7698 GND.n726 9.3005
R20669 GND.n7699 GND.n725 9.3005
R20670 GND.n7702 GND.n724 9.3005
R20671 GND.n7703 GND.n723 9.3005
R20672 GND.n7706 GND.n722 9.3005
R20673 GND.n7708 GND.n721 9.3005
R20674 GND.n7709 GND.n718 9.3005
R20675 GND.n7710 GND.n716 9.3005
R20676 GND.n7713 GND.n715 9.3005
R20677 GND.n7714 GND.n714 9.3005
R20678 GND.n7717 GND.n713 9.3005
R20679 GND.n7719 GND.n712 9.3005
R20680 GND.n7720 GND.n711 9.3005
R20681 GND.n7721 GND.n710 9.3005
R20682 GND.n7722 GND.n709 9.3005
R20683 GND.n7672 GND.n7603 9.3005
R20684 GND.n7630 GND.n7627 9.3005
R20685 GND.n7757 GND.n7756 9.3005
R20686 GND.n7758 GND.n643 9.3005
R20687 GND.n7762 GND.n7759 9.3005
R20688 GND.n7761 GND.n7760 9.3005
R20689 GND.n617 GND.n616 9.3005
R20690 GND.n7794 GND.n7793 9.3005
R20691 GND.n7795 GND.n615 9.3005
R20692 GND.n7799 GND.n7796 9.3005
R20693 GND.n7798 GND.n7797 9.3005
R20694 GND.n590 GND.n589 9.3005
R20695 GND.n7829 GND.n7828 9.3005
R20696 GND.n7830 GND.n588 9.3005
R20697 GND.n7832 GND.n7831 9.3005
R20698 GND.n568 GND.n567 9.3005
R20699 GND.n7856 GND.n7855 9.3005
R20700 GND.n7857 GND.n566 9.3005
R20701 GND.n7859 GND.n7858 9.3005
R20702 GND.n534 GND.n533 9.3005
R20703 GND.n7894 GND.n7893 9.3005
R20704 GND.n7895 GND.n532 9.3005
R20705 GND.n7897 GND.n7896 9.3005
R20706 GND.n503 GND.n502 9.3005
R20707 GND.n7947 GND.n7946 9.3005
R20708 GND.n7948 GND.n501 9.3005
R20709 GND.n7952 GND.n7949 9.3005
R20710 GND.n7951 GND.n7950 9.3005
R20711 GND.n476 GND.n475 9.3005
R20712 GND.n7984 GND.n7983 9.3005
R20713 GND.n7985 GND.n474 9.3005
R20714 GND.n7989 GND.n7986 9.3005
R20715 GND.n7988 GND.n167 9.3005
R20716 GND.n174 GND.n166 9.3005
R20717 GND.n8551 GND.n194 9.3005
R20718 GND.n8550 GND.n195 9.3005
R20719 GND.n8549 GND.n196 9.3005
R20720 GND.n214 GND.n197 9.3005
R20721 GND.n8539 GND.n215 9.3005
R20722 GND.n8538 GND.n216 9.3005
R20723 GND.n8537 GND.n217 9.3005
R20724 GND.n235 GND.n218 9.3005
R20725 GND.n8527 GND.n236 9.3005
R20726 GND.n8526 GND.n237 9.3005
R20727 GND.n8525 GND.n238 9.3005
R20728 GND.n255 GND.n239 9.3005
R20729 GND.n8515 GND.n256 9.3005
R20730 GND.n8514 GND.n257 9.3005
R20731 GND.n8513 GND.n258 9.3005
R20732 GND.n276 GND.n259 9.3005
R20733 GND.n8503 GND.n277 9.3005
R20734 GND.n8502 GND.n278 9.3005
R20735 GND.n8501 GND.n279 9.3005
R20736 GND.n297 GND.n280 9.3005
R20737 GND.n8491 GND.n298 9.3005
R20738 GND.n8490 GND.n299 9.3005
R20739 GND.n8489 GND.n300 9.3005
R20740 GND.n317 GND.n301 9.3005
R20741 GND.n8479 GND.n318 9.3005
R20742 GND.n8478 GND.n319 9.3005
R20743 GND.n8477 GND.n320 9.3005
R20744 GND.n338 GND.n321 9.3005
R20745 GND.n8467 GND.n339 9.3005
R20746 GND.n8466 GND.n340 9.3005
R20747 GND.n8465 GND.n341 9.3005
R20748 GND.n645 GND.n644 9.3005
R20749 GND.n8562 GND.n171 9.3005
R20750 GND.n8562 GND.n8561 9.3005
R20751 GND.n1872 GND.n1856 9.3005
R20752 GND.n1854 GND.n1853 9.3005
R20753 GND.n4710 GND.n4709 9.3005
R20754 GND.n4711 GND.n1852 9.3005
R20755 GND.n4726 GND.n4712 9.3005
R20756 GND.n4725 GND.n4713 9.3005
R20757 GND.n4724 GND.n4714 9.3005
R20758 GND.n4716 GND.n4715 9.3005
R20759 GND.n4720 GND.n4717 9.3005
R20760 GND.n4719 GND.n4718 9.3005
R20761 GND.n1790 GND.n1789 9.3005
R20762 GND.n4803 GND.n4802 9.3005
R20763 GND.n4804 GND.n1788 9.3005
R20764 GND.n4829 GND.n4805 9.3005
R20765 GND.n4828 GND.n4806 9.3005
R20766 GND.n4827 GND.n4807 9.3005
R20767 GND.n4810 GND.n4808 9.3005
R20768 GND.n4823 GND.n4811 9.3005
R20769 GND.n4822 GND.n4812 9.3005
R20770 GND.n4821 GND.n4813 9.3005
R20771 GND.n4815 GND.n4814 9.3005
R20772 GND.n4817 GND.n4816 9.3005
R20773 GND.n1708 GND.n1707 9.3005
R20774 GND.n4933 GND.n4932 9.3005
R20775 GND.n4934 GND.n1706 9.3005
R20776 GND.n5858 GND.n4935 9.3005
R20777 GND.n5857 GND.n4936 9.3005
R20778 GND.n5856 GND.n4937 9.3005
R20779 GND.n4940 GND.n4938 9.3005
R20780 GND.n5852 GND.n4941 9.3005
R20781 GND.n5851 GND.n4942 9.3005
R20782 GND.n5850 GND.n4943 9.3005
R20783 GND.n4946 GND.n4944 9.3005
R20784 GND.n5846 GND.n4947 9.3005
R20785 GND.n5845 GND.n4948 9.3005
R20786 GND.n5844 GND.n4949 9.3005
R20787 GND.n4955 GND.n4950 9.3005
R20788 GND.n5838 GND.n4956 9.3005
R20789 GND.n5837 GND.n4957 9.3005
R20790 GND.n5836 GND.n4958 9.3005
R20791 GND.n4973 GND.n4959 9.3005
R20792 GND.n5824 GND.n4974 9.3005
R20793 GND.n5823 GND.n4975 9.3005
R20794 GND.n5822 GND.n4976 9.3005
R20795 GND.n4991 GND.n4977 9.3005
R20796 GND.n5810 GND.n4992 9.3005
R20797 GND.n5809 GND.n4993 9.3005
R20798 GND.n5808 GND.n4994 9.3005
R20799 GND.n5008 GND.n4995 9.3005
R20800 GND.n5796 GND.n5009 9.3005
R20801 GND.n5795 GND.n5010 9.3005
R20802 GND.n5794 GND.n5011 9.3005
R20803 GND.n5026 GND.n5012 9.3005
R20804 GND.n5782 GND.n5027 9.3005
R20805 GND.n5781 GND.n5028 9.3005
R20806 GND.n5780 GND.n5029 9.3005
R20807 GND.n5044 GND.n5030 9.3005
R20808 GND.n5768 GND.n5045 9.3005
R20809 GND.n5767 GND.n5046 9.3005
R20810 GND.n5766 GND.n5047 9.3005
R20811 GND.n5065 GND.n5048 9.3005
R20812 GND.n5066 GND.n5064 9.3005
R20813 GND.n5753 GND.n5067 9.3005
R20814 GND.n5752 GND.n5068 9.3005
R20815 GND.n5751 GND.n5069 9.3005
R20816 GND.n5083 GND.n5070 9.3005
R20817 GND.n5739 GND.n5084 9.3005
R20818 GND.n5738 GND.n5085 9.3005
R20819 GND.n5737 GND.n5086 9.3005
R20820 GND.n5101 GND.n5087 9.3005
R20821 GND.n5725 GND.n5102 9.3005
R20822 GND.n5724 GND.n5103 9.3005
R20823 GND.n5723 GND.n5104 9.3005
R20824 GND.n5119 GND.n5105 9.3005
R20825 GND.n5711 GND.n5120 9.3005
R20826 GND.n5710 GND.n5121 9.3005
R20827 GND.n5709 GND.n5122 9.3005
R20828 GND.n5140 GND.n5123 9.3005
R20829 GND.n5141 GND.n5139 9.3005
R20830 GND.n5696 GND.n5142 9.3005
R20831 GND.n5695 GND.n5143 9.3005
R20832 GND.n5694 GND.n5144 9.3005
R20833 GND.n5159 GND.n5145 9.3005
R20834 GND.n5682 GND.n5160 9.3005
R20835 GND.n5681 GND.n5161 9.3005
R20836 GND.n5680 GND.n5162 9.3005
R20837 GND.n5177 GND.n5163 9.3005
R20838 GND.n5668 GND.n5178 9.3005
R20839 GND.n5667 GND.n5179 9.3005
R20840 GND.n5666 GND.n5180 9.3005
R20841 GND.n5652 GND.n5181 9.3005
R20842 GND.n5654 GND.n5653 9.3005
R20843 GND.n1573 GND.n1572 9.3005
R20844 GND.n6104 GND.n6103 9.3005
R20845 GND.n6105 GND.n1571 9.3005
R20846 GND.n6107 GND.n6106 9.3005
R20847 GND.n1559 GND.n1558 9.3005
R20848 GND.n6120 GND.n6119 9.3005
R20849 GND.n6121 GND.n1557 9.3005
R20850 GND.n6123 GND.n6122 9.3005
R20851 GND.n1542 GND.n1541 9.3005
R20852 GND.n6145 GND.n6144 9.3005
R20853 GND.n6146 GND.n1540 9.3005
R20854 GND.n6148 GND.n6147 9.3005
R20855 GND.n1499 GND.n1498 9.3005
R20856 GND.n6324 GND.n6323 9.3005
R20857 GND.n6325 GND.n1497 9.3005
R20858 GND.n6327 GND.n6326 9.3005
R20859 GND.n1483 GND.n1482 9.3005
R20860 GND.n6340 GND.n6339 9.3005
R20861 GND.n6341 GND.n1481 9.3005
R20862 GND.n6343 GND.n6342 9.3005
R20863 GND.n1467 GND.n1466 9.3005
R20864 GND.n6356 GND.n6355 9.3005
R20865 GND.n6357 GND.n1465 9.3005
R20866 GND.n6359 GND.n6358 9.3005
R20867 GND.n1451 GND.n1450 9.3005
R20868 GND.n6372 GND.n6371 9.3005
R20869 GND.n6373 GND.n1449 9.3005
R20870 GND.n6375 GND.n6374 9.3005
R20871 GND.n1435 GND.n1434 9.3005
R20872 GND.n6387 GND.n6386 9.3005
R20873 GND.n6388 GND.n1433 9.3005
R20874 GND.n6392 GND.n6389 9.3005
R20875 GND.n6391 GND.n6390 9.3005
R20876 GND.n1317 GND.n1316 9.3005
R20877 GND.n6563 GND.n6562 9.3005
R20878 GND.n6564 GND.n1315 9.3005
R20879 GND.n6566 GND.n6565 9.3005
R20880 GND.n1302 GND.n1301 9.3005
R20881 GND.n6579 GND.n6578 9.3005
R20882 GND.n6580 GND.n1300 9.3005
R20883 GND.n6582 GND.n6581 9.3005
R20884 GND.n1286 GND.n1285 9.3005
R20885 GND.n6595 GND.n6594 9.3005
R20886 GND.n6596 GND.n1284 9.3005
R20887 GND.n6598 GND.n6597 9.3005
R20888 GND.n1270 GND.n1269 9.3005
R20889 GND.n6611 GND.n6610 9.3005
R20890 GND.n6612 GND.n1268 9.3005
R20891 GND.n6614 GND.n6613 9.3005
R20892 GND.n1254 GND.n1253 9.3005
R20893 GND.n6626 GND.n6625 9.3005
R20894 GND.n6627 GND.n1252 9.3005
R20895 GND.n6629 GND.n6628 9.3005
R20896 GND.n1238 GND.n1237 9.3005
R20897 GND.n6642 GND.n6641 9.3005
R20898 GND.n6643 GND.n1236 9.3005
R20899 GND.n6645 GND.n6644 9.3005
R20900 GND.n1221 GND.n1220 9.3005
R20901 GND.n6667 GND.n6666 9.3005
R20902 GND.n6668 GND.n1219 9.3005
R20903 GND.n6670 GND.n6669 9.3005
R20904 GND.n1164 GND.n1163 9.3005
R20905 GND.n6821 GND.n6820 9.3005
R20906 GND.n6822 GND.n1162 9.3005
R20907 GND.n6824 GND.n6823 9.3005
R20908 GND.n1148 GND.n1147 9.3005
R20909 GND.n6837 GND.n6836 9.3005
R20910 GND.n6838 GND.n1146 9.3005
R20911 GND.n6840 GND.n6839 9.3005
R20912 GND.n1132 GND.n1131 9.3005
R20913 GND.n6853 GND.n6852 9.3005
R20914 GND.n6854 GND.n1130 9.3005
R20915 GND.n6856 GND.n6855 9.3005
R20916 GND.n1116 GND.n1115 9.3005
R20917 GND.n6869 GND.n6868 9.3005
R20918 GND.n6870 GND.n1114 9.3005
R20919 GND.n6872 GND.n6871 9.3005
R20920 GND.n1099 GND.n1098 9.3005
R20921 GND.n6889 GND.n6888 9.3005
R20922 GND.n6890 GND.n1097 9.3005
R20923 GND.n6892 GND.n6891 9.3005
R20924 GND.n1053 GND.n1052 9.3005
R20925 GND.n6982 GND.n6981 9.3005
R20926 GND.n6983 GND.n1051 9.3005
R20927 GND.n6990 GND.n6984 9.3005
R20928 GND.n6989 GND.n6985 9.3005
R20929 GND.n6988 GND.n6986 9.3005
R20930 GND.n1029 GND.n1028 9.3005
R20931 GND.n7022 GND.n7021 9.3005
R20932 GND.n7023 GND.n1027 9.3005
R20933 GND.n7036 GND.n7024 9.3005
R20934 GND.n7035 GND.n7025 9.3005
R20935 GND.n7034 GND.n7026 9.3005
R20936 GND.n7028 GND.n7027 9.3005
R20937 GND.n7030 GND.n7029 9.3005
R20938 GND.n995 GND.n994 9.3005
R20939 GND.n7080 GND.n7079 9.3005
R20940 GND.n7081 GND.n993 9.3005
R20941 GND.n7085 GND.n7082 9.3005
R20942 GND.n7084 GND.n7083 9.3005
R20943 GND.n970 GND.n969 9.3005
R20944 GND.n7115 GND.n7114 9.3005
R20945 GND.n7116 GND.n968 9.3005
R20946 GND.n7123 GND.n7117 9.3005
R20947 GND.n7122 GND.n7118 9.3005
R20948 GND.n7121 GND.n7119 9.3005
R20949 GND.n945 GND.n944 9.3005
R20950 GND.n7154 GND.n7153 9.3005
R20951 GND.n7155 GND.n943 9.3005
R20952 GND.n7168 GND.n7156 9.3005
R20953 GND.n7167 GND.n7157 9.3005
R20954 GND.n7166 GND.n7158 9.3005
R20955 GND.n7160 GND.n7159 9.3005
R20956 GND.n7162 GND.n7161 9.3005
R20957 GND.n913 GND.n912 9.3005
R20958 GND.n7214 GND.n7213 9.3005
R20959 GND.n7215 GND.n911 9.3005
R20960 GND.n7237 GND.n7216 9.3005
R20961 GND.n7236 GND.n7217 9.3005
R20962 GND.n7235 GND.n7218 9.3005
R20963 GND.n7221 GND.n7219 9.3005
R20964 GND.n7231 GND.n7222 9.3005
R20965 GND.n7230 GND.n7223 9.3005
R20966 GND.n7229 GND.n7224 9.3005
R20967 GND.n7226 GND.n7225 9.3005
R20968 GND.n869 GND.n868 9.3005
R20969 GND.n7294 GND.n7293 9.3005
R20970 GND.n7295 GND.n867 9.3005
R20971 GND.n7299 GND.n7296 9.3005
R20972 GND.n7298 GND.n7297 9.3005
R20973 GND.n844 GND.n843 9.3005
R20974 GND.n7330 GND.n7329 9.3005
R20975 GND.n7331 GND.n842 9.3005
R20976 GND.n7333 GND.n7332 9.3005
R20977 GND.n828 GND.n827 9.3005
R20978 GND.n7353 GND.n7352 9.3005
R20979 GND.n7354 GND.n826 9.3005
R20980 GND.n7358 GND.n7355 9.3005
R20981 GND.n7357 GND.n7356 9.3005
R20982 GND.n804 GND.n803 9.3005
R20983 GND.n7445 GND.n7444 9.3005
R20984 GND.n7446 GND.n802 9.3005
R20985 GND.n7532 GND.n7447 9.3005
R20986 GND.n7531 GND.n7448 9.3005
R20987 GND.n7530 GND.n7449 9.3005
R20988 GND.n7454 GND.n7450 9.3005
R20989 GND.n7524 GND.n7455 9.3005
R20990 GND.n7523 GND.n7456 9.3005
R20991 GND.n7522 GND.n7457 9.3005
R20992 GND.n7460 GND.n7458 9.3005
R20993 GND.n7518 GND.n7461 9.3005
R20994 GND.n7517 GND.n7462 9.3005
R20995 GND.n7516 GND.n7463 9.3005
R20996 GND.n7466 GND.n7464 9.3005
R20997 GND.n7512 GND.n7467 9.3005
R20998 GND.n7511 GND.n7468 9.3005
R20999 GND.n7510 GND.n7469 9.3005
R21000 GND.n7472 GND.n7470 9.3005
R21001 GND.n7506 GND.n7473 9.3005
R21002 GND.n7505 GND.n7474 9.3005
R21003 GND.n7504 GND.n7475 9.3005
R21004 GND.n7478 GND.n7476 9.3005
R21005 GND.n7500 GND.n7479 9.3005
R21006 GND.n7499 GND.n7480 9.3005
R21007 GND.n7498 GND.n7481 9.3005
R21008 GND.n7484 GND.n7482 9.3005
R21009 GND.n7494 GND.n7485 9.3005
R21010 GND.n7493 GND.n7486 9.3005
R21011 GND.n7492 GND.n7487 9.3005
R21012 GND.n7489 GND.n7488 9.3005
R21013 GND.n524 GND.n523 9.3005
R21014 GND.n7903 GND.n7902 9.3005
R21015 GND.n7904 GND.n522 9.3005
R21016 GND.n7906 GND.n7905 9.3005
R21017 GND.n520 GND.n519 9.3005
R21018 GND.n7911 GND.n7910 9.3005
R21019 GND.n7912 GND.n518 9.3005
R21020 GND.n7934 GND.n7913 9.3005
R21021 GND.n7933 GND.n7914 9.3005
R21022 GND.n7932 GND.n7915 9.3005
R21023 GND.n7918 GND.n7916 9.3005
R21024 GND.n7928 GND.n7919 9.3005
R21025 GND.n8041 GND.n8039 9.3005
R21026 GND.n8113 GND.n8042 9.3005
R21027 GND.n8112 GND.n8043 9.3005
R21028 GND.n8111 GND.n8044 9.3005
R21029 GND.n8047 GND.n8045 9.3005
R21030 GND.n8107 GND.n8048 9.3005
R21031 GND.n8106 GND.n8049 9.3005
R21032 GND.n8105 GND.n8050 9.3005
R21033 GND.n8053 GND.n8051 9.3005
R21034 GND.n8101 GND.n8054 9.3005
R21035 GND.n8100 GND.n8055 9.3005
R21036 GND.n8099 GND.n8056 9.3005
R21037 GND.n8059 GND.n8057 9.3005
R21038 GND.n8095 GND.n8060 9.3005
R21039 GND.n8094 GND.n8061 9.3005
R21040 GND.n8093 GND.n8062 9.3005
R21041 GND.n8065 GND.n8063 9.3005
R21042 GND.n8089 GND.n8066 9.3005
R21043 GND.n8088 GND.n8067 9.3005
R21044 GND.n8087 GND.n8068 9.3005
R21045 GND.n8071 GND.n8069 9.3005
R21046 GND.n8083 GND.n8072 9.3005
R21047 GND.n8082 GND.n8073 9.3005
R21048 GND.n8081 GND.n8074 9.3005
R21049 GND.n8078 GND.n8075 9.3005
R21050 GND.n8077 GND.n8076 9.3005
R21051 GND.n391 GND.n390 9.3005
R21052 GND.n8251 GND.n8250 9.3005
R21053 GND.n8252 GND.n389 9.3005
R21054 GND.n8255 GND.n8254 9.3005
R21055 GND.n8253 GND.n387 9.3005
R21056 GND.n8259 GND.n386 9.3005
R21057 GND.n8261 GND.n8260 9.3005
R21058 GND.n4219 GND.n4218 9.3005
R21059 GND.n4222 GND.n4213 9.3005
R21060 GND.n4223 GND.n4212 9.3005
R21061 GND.n4226 GND.n4211 9.3005
R21062 GND.n4227 GND.n4210 9.3005
R21063 GND.n4230 GND.n4209 9.3005
R21064 GND.n4231 GND.n4208 9.3005
R21065 GND.n4234 GND.n4207 9.3005
R21066 GND.n4235 GND.n4206 9.3005
R21067 GND.n4238 GND.n4205 9.3005
R21068 GND.n4239 GND.n4202 9.3005
R21069 GND.n4242 GND.n4201 9.3005
R21070 GND.n4243 GND.n4200 9.3005
R21071 GND.n4246 GND.n4199 9.3005
R21072 GND.n4247 GND.n4198 9.3005
R21073 GND.n4250 GND.n4197 9.3005
R21074 GND.n4251 GND.n4196 9.3005
R21075 GND.n4254 GND.n4195 9.3005
R21076 GND.n4255 GND.n4194 9.3005
R21077 GND.n4258 GND.n4193 9.3005
R21078 GND.n4262 GND.n4189 9.3005
R21079 GND.n4263 GND.n4188 9.3005
R21080 GND.n4266 GND.n4187 9.3005
R21081 GND.n4267 GND.n4186 9.3005
R21082 GND.n4270 GND.n4185 9.3005
R21083 GND.n4271 GND.n4184 9.3005
R21084 GND.n4274 GND.n4183 9.3005
R21085 GND.n4275 GND.n4182 9.3005
R21086 GND.n4278 GND.n4181 9.3005
R21087 GND.n4280 GND.n4178 9.3005
R21088 GND.n4283 GND.n4177 9.3005
R21089 GND.n4284 GND.n4176 9.3005
R21090 GND.n4287 GND.n4175 9.3005
R21091 GND.n4288 GND.n4174 9.3005
R21092 GND.n4291 GND.n4173 9.3005
R21093 GND.n4292 GND.n4172 9.3005
R21094 GND.n4295 GND.n4171 9.3005
R21095 GND.n4297 GND.n4170 9.3005
R21096 GND.n4298 GND.n4167 9.3005
R21097 GND.n4299 GND.n4165 9.3005
R21098 GND.n4302 GND.n4164 9.3005
R21099 GND.n4303 GND.n4163 9.3005
R21100 GND.n4306 GND.n4162 9.3005
R21101 GND.n4308 GND.n4161 9.3005
R21102 GND.n4309 GND.n4160 9.3005
R21103 GND.n4310 GND.n4159 9.3005
R21104 GND.n4158 GND.n2128 9.3005
R21105 GND.n4259 GND.n4190 9.3005
R21106 GND.n4215 GND.n2137 9.3005
R21107 GND.n4349 GND.n2127 9.3005
R21108 GND.n4353 GND.n4350 9.3005
R21109 GND.n4352 GND.n4351 9.3005
R21110 GND.n2100 GND.n2099 9.3005
R21111 GND.n4384 GND.n4383 9.3005
R21112 GND.n4385 GND.n2098 9.3005
R21113 GND.n4389 GND.n4386 9.3005
R21114 GND.n4388 GND.n4387 9.3005
R21115 GND.n2071 GND.n2070 9.3005
R21116 GND.n4427 GND.n4426 9.3005
R21117 GND.n4428 GND.n2069 9.3005
R21118 GND.n4430 GND.n4429 9.3005
R21119 GND.n2037 GND.n2036 9.3005
R21120 GND.n4466 GND.n4465 9.3005
R21121 GND.n4467 GND.n2035 9.3005
R21122 GND.n4471 GND.n4468 9.3005
R21123 GND.n4470 GND.n4469 9.3005
R21124 GND.n2009 GND.n2008 9.3005
R21125 GND.n4509 GND.n4508 9.3005
R21126 GND.n4510 GND.n2007 9.3005
R21127 GND.n4512 GND.n4511 9.3005
R21128 GND.n1975 GND.n1974 9.3005
R21129 GND.n4584 GND.n4583 9.3005
R21130 GND.n4585 GND.n1973 9.3005
R21131 GND.n4589 GND.n4586 9.3005
R21132 GND.n4588 GND.n4587 9.3005
R21133 GND.n1945 GND.n1944 9.3005
R21134 GND.n4616 GND.n4615 9.3005
R21135 GND.n4617 GND.n1943 9.3005
R21136 GND.n4619 GND.n4618 9.3005
R21137 GND.n1879 GND.n1871 9.3005
R21138 GND.n4691 GND.n4690 9.3005
R21139 GND.n1834 GND.n1833 9.3005
R21140 GND.n4743 GND.n4742 9.3005
R21141 GND.n4744 GND.n1832 9.3005
R21142 GND.n4748 GND.n4745 9.3005
R21143 GND.n4747 GND.n4746 9.3005
R21144 GND.n1807 GND.n1806 9.3005
R21145 GND.n4781 GND.n4780 9.3005
R21146 GND.n4782 GND.n1805 9.3005
R21147 GND.n4786 GND.n4783 9.3005
R21148 GND.n4785 GND.n4784 9.3005
R21149 GND.n1773 GND.n1772 9.3005
R21150 GND.n4849 GND.n4848 9.3005
R21151 GND.n4850 GND.n1771 9.3005
R21152 GND.n4854 GND.n4851 9.3005
R21153 GND.n4853 GND.n4852 9.3005
R21154 GND.n1746 GND.n1745 9.3005
R21155 GND.n4886 GND.n4885 9.3005
R21156 GND.n4887 GND.n1744 9.3005
R21157 GND.n4891 GND.n4888 9.3005
R21158 GND.n4890 GND.n4889 9.3005
R21159 GND.n1716 GND.n1715 9.3005
R21160 GND.n4924 GND.n4923 9.3005
R21161 GND.n4925 GND.n1714 9.3005
R21162 GND.n4927 GND.n4926 9.3005
R21163 GND.n1689 GND.n1688 9.3005
R21164 GND.n5884 GND.n5883 9.3005
R21165 GND.n5885 GND.n1687 9.3005
R21166 GND.n5888 GND.n5887 9.3005
R21167 GND.n5886 GND.n1674 9.3005
R21168 GND.n5901 GND.n1673 9.3005
R21169 GND.n5903 GND.n5902 9.3005
R21170 GND.n4348 GND.n4347 9.3005
R21171 GND.n4689 GND.n1877 9.3005
R21172 GND.n4692 GND.n4689 9.3005
R21173 GND.n4122 GND.n4093 9.3005
R21174 GND.n4096 GND.n4094 9.3005
R21175 GND.n4118 GND.n4097 9.3005
R21176 GND.n4117 GND.n4098 9.3005
R21177 GND.n4116 GND.n4099 9.3005
R21178 GND.n4102 GND.n4100 9.3005
R21179 GND.n4112 GND.n4103 9.3005
R21180 GND.n4111 GND.n4104 9.3005
R21181 GND.n4110 GND.n4105 9.3005
R21182 GND.n4107 GND.n4106 9.3005
R21183 GND.n2061 GND.n2060 9.3005
R21184 GND.n4436 GND.n4435 9.3005
R21185 GND.n4437 GND.n2059 9.3005
R21186 GND.n4439 GND.n4438 9.3005
R21187 GND.n2057 GND.n2056 9.3005
R21188 GND.n4444 GND.n4443 9.3005
R21189 GND.n4445 GND.n2055 9.3005
R21190 GND.n4449 GND.n4446 9.3005
R21191 GND.n4448 GND.n4447 9.3005
R21192 GND.n1999 GND.n1998 9.3005
R21193 GND.n4518 GND.n4517 9.3005
R21194 GND.n4519 GND.n1997 9.3005
R21195 GND.n4521 GND.n4520 9.3005
R21196 GND.n1995 GND.n1994 9.3005
R21197 GND.n4526 GND.n4525 9.3005
R21198 GND.n4527 GND.n1993 9.3005
R21199 GND.n4567 GND.n4528 9.3005
R21200 GND.n4566 GND.n4529 9.3005
R21201 GND.n4565 GND.n4530 9.3005
R21202 GND.n4533 GND.n4531 9.3005
R21203 GND.n4561 GND.n4534 9.3005
R21204 GND.n4560 GND.n4535 9.3005
R21205 GND.n4124 GND.n4123 9.3005
R21206 GND.n4092 GND.n2155 9.3005
R21207 GND.n4091 GND.n4090 9.3005
R21208 GND.n2157 GND.n2156 9.3005
R21209 GND.n4084 GND.n4083 9.3005
R21210 GND.n4082 GND.n2161 9.3005
R21211 GND.n4081 GND.n4080 9.3005
R21212 GND.n2163 GND.n2162 9.3005
R21213 GND.n4074 GND.n4073 9.3005
R21214 GND.n4072 GND.n2167 9.3005
R21215 GND.n4071 GND.n4070 9.3005
R21216 GND.n2169 GND.n2168 9.3005
R21217 GND.n4064 GND.n4063 9.3005
R21218 GND.n4062 GND.n2173 9.3005
R21219 GND.n4061 GND.n4060 9.3005
R21220 GND.n2175 GND.n2174 9.3005
R21221 GND.n4054 GND.n4053 9.3005
R21222 GND.n4052 GND.n2179 9.3005
R21223 GND.n4051 GND.n4050 9.3005
R21224 GND.n2181 GND.n2180 9.3005
R21225 GND.n4044 GND.n4043 9.3005
R21226 GND.n4042 GND.n2185 9.3005
R21227 GND.n4041 GND.n4040 9.3005
R21228 GND.n2187 GND.n2186 9.3005
R21229 GND.n4034 GND.n4033 9.3005
R21230 GND.n4032 GND.n2191 9.3005
R21231 GND.n4031 GND.n4030 9.3005
R21232 GND.n2193 GND.n2192 9.3005
R21233 GND.n4024 GND.n4023 9.3005
R21234 GND.n4022 GND.n2197 9.3005
R21235 GND.n4021 GND.n4020 9.3005
R21236 GND.n2199 GND.n2198 9.3005
R21237 GND.n4014 GND.n4013 9.3005
R21238 GND.n4012 GND.n2203 9.3005
R21239 GND.n4011 GND.n4010 9.3005
R21240 GND.n2205 GND.n2204 9.3005
R21241 GND.n4004 GND.n4003 9.3005
R21242 GND.n4002 GND.n2209 9.3005
R21243 GND.n4001 GND.n4000 9.3005
R21244 GND.n2211 GND.n2210 9.3005
R21245 GND.n3994 GND.n3993 9.3005
R21246 GND.n3992 GND.n2215 9.3005
R21247 GND.n3991 GND.n3990 9.3005
R21248 GND.n2217 GND.n2216 9.3005
R21249 GND.n3984 GND.n3983 9.3005
R21250 GND.n3982 GND.n2221 9.3005
R21251 GND.n3981 GND.n3980 9.3005
R21252 GND.n2223 GND.n2222 9.3005
R21253 GND.n3974 GND.n3973 9.3005
R21254 GND.n3972 GND.n2227 9.3005
R21255 GND.n3971 GND.n3970 9.3005
R21256 GND.n2229 GND.n2228 9.3005
R21257 GND.n3964 GND.n3963 9.3005
R21258 GND.n3962 GND.n2233 9.3005
R21259 GND.n3961 GND.n3960 9.3005
R21260 GND.n2235 GND.n2234 9.3005
R21261 GND.n3954 GND.n3953 9.3005
R21262 GND.n3952 GND.n2239 9.3005
R21263 GND.n3951 GND.n3950 9.3005
R21264 GND.n2241 GND.n2240 9.3005
R21265 GND.n3944 GND.n3943 9.3005
R21266 GND.n3942 GND.n2245 9.3005
R21267 GND.n3941 GND.n3940 9.3005
R21268 GND.n2247 GND.n2246 9.3005
R21269 GND.n4126 GND.n4125 9.3005
R21270 GND.n6051 GND.n1599 9.3005
R21271 GND.n6072 GND.n6052 9.3005
R21272 GND.n5958 GND.n5957 9.3005
R21273 GND.n5954 GND.n1660 9.3005
R21274 GND.n5953 GND.n5952 9.3005
R21275 GND.n5951 GND.n5950 9.3005
R21276 GND.n5948 GND.n1665 9.3005
R21277 GND.n5945 GND.n5944 9.3005
R21278 GND.n5943 GND.n1666 9.3005
R21279 GND.n5942 GND.n5941 9.3005
R21280 GND.n5938 GND.n1667 9.3005
R21281 GND.n5935 GND.n5934 9.3005
R21282 GND.n5933 GND.n1668 9.3005
R21283 GND.n5932 GND.n5931 9.3005
R21284 GND.n5928 GND.n1669 9.3005
R21285 GND.n5923 GND.n5922 9.3005
R21286 GND.n5921 GND.n1670 9.3005
R21287 GND.n5920 GND.n5919 9.3005
R21288 GND.n5916 GND.n1671 9.3005
R21289 GND.n5913 GND.n5912 9.3005
R21290 GND.n5911 GND.n1672 9.3005
R21291 GND.n5910 GND.n5909 9.3005
R21292 GND.n5906 GND.n5904 9.3005
R21293 GND.n6039 GND.n6038 9.3005
R21294 GND.n6037 GND.n1659 9.3005
R21295 GND.n6036 GND.n6035 9.3005
R21296 GND.n6034 GND.n5960 9.3005
R21297 GND.n6033 GND.n5966 9.3005
R21298 GND.n6032 GND.n6031 9.3005
R21299 GND.n6030 GND.n5970 9.3005
R21300 GND.n6029 GND.n6028 9.3005
R21301 GND.n6027 GND.n5971 9.3005
R21302 GND.n6026 GND.n6025 9.3005
R21303 GND.n6024 GND.n5976 9.3005
R21304 GND.n6023 GND.n6022 9.3005
R21305 GND.n6021 GND.n5977 9.3005
R21306 GND.n6020 GND.n6019 9.3005
R21307 GND.n6018 GND.n5984 9.3005
R21308 GND.n6017 GND.n6016 9.3005
R21309 GND.n6015 GND.n5985 9.3005
R21310 GND.n6014 GND.n6013 9.3005
R21311 GND.n6012 GND.n5990 9.3005
R21312 GND.n6011 GND.n6010 9.3005
R21313 GND.n6009 GND.n5991 9.3005
R21314 GND.n6008 GND.n6007 9.3005
R21315 GND.n6006 GND.n5996 9.3005
R21316 GND.n6005 GND.n6004 9.3005
R21317 GND.n6003 GND.n5997 9.3005
R21318 GND.n6002 GND.n1601 9.3005
R21319 GND.n4330 GND.n2136 9.3005
R21320 GND.n4338 GND.n4333 9.3005
R21321 GND.n4337 GND.n4336 9.3005
R21322 GND.n2110 GND.n2108 9.3005
R21323 GND.n4379 GND.n4378 9.3005
R21324 GND.n2111 GND.n2109 9.3005
R21325 GND.n4374 GND.n4369 9.3005
R21326 GND.n4373 GND.n4372 9.3005
R21327 GND.n2081 GND.n2079 9.3005
R21328 GND.n4422 GND.n4421 9.3005
R21329 GND.n2082 GND.n2080 9.3005
R21330 GND.n4417 GND.n4416 9.3005
R21331 GND.n2047 GND.n2045 9.3005
R21332 GND.n4461 GND.n4460 9.3005
R21333 GND.n2048 GND.n2046 9.3005
R21334 GND.n4456 GND.n2052 9.3005
R21335 GND.n4455 GND.n4454 9.3005
R21336 GND.n2019 GND.n2017 9.3005
R21337 GND.n4504 GND.n4503 9.3005
R21338 GND.n2020 GND.n2018 9.3005
R21339 GND.n4499 GND.n4498 9.3005
R21340 GND.n1985 GND.n1983 9.3005
R21341 GND.n4579 GND.n4578 9.3005
R21342 GND.n1986 GND.n1984 9.3005
R21343 GND.n4574 GND.n1990 9.3005
R21344 GND.n4573 GND.n4572 9.3005
R21345 GND.n1955 GND.n1953 9.3005
R21346 GND.n4611 GND.n4610 9.3005
R21347 GND.n1958 GND.n1954 9.3005
R21348 GND.n1957 GND.n1956 9.3005
R21349 GND.n1890 GND.n1888 9.3005
R21350 GND.n4683 GND.n4682 9.3005
R21351 GND.n1891 GND.n1889 9.3005
R21352 GND.n4678 GND.n1896 9.3005
R21353 GND.n4677 GND.n1897 9.3005
R21354 GND.n4676 GND.n1898 9.3005
R21355 GND.n1922 GND.n1899 9.3005
R21356 GND.n4672 GND.n1904 9.3005
R21357 GND.n4671 GND.n1905 9.3005
R21358 GND.n4670 GND.n1906 9.3005
R21359 GND.n4663 GND.n1907 9.3005
R21360 GND.n4666 GND.n4665 9.3005
R21361 GND.n1844 GND.n1842 9.3005
R21362 GND.n4738 GND.n4737 9.3005
R21363 GND.n1845 GND.n1843 9.3005
R21364 GND.n4733 GND.n1849 9.3005
R21365 GND.n4732 GND.n4731 9.3005
R21366 GND.n1817 GND.n1815 9.3005
R21367 GND.n4776 GND.n4775 9.3005
R21368 GND.n1818 GND.n1816 9.3005
R21369 GND.n4771 GND.n4767 9.3005
R21370 GND.n4770 GND.n4769 9.3005
R21371 GND.n1783 GND.n1781 9.3005
R21372 GND.n4844 GND.n4843 9.3005
R21373 GND.n1784 GND.n1782 9.3005
R21374 GND.n4839 GND.n4834 9.3005
R21375 GND.n4838 GND.n4837 9.3005
R21376 GND.n1756 GND.n1754 9.3005
R21377 GND.n4881 GND.n4880 9.3005
R21378 GND.n1757 GND.n1755 9.3005
R21379 GND.n4876 GND.n4871 9.3005
R21380 GND.n4875 GND.n4874 9.3005
R21381 GND.n1726 GND.n1724 9.3005
R21382 GND.n4919 GND.n4918 9.3005
R21383 GND.n1729 GND.n1725 9.3005
R21384 GND.n1728 GND.n1727 9.3005
R21385 GND.n1698 GND.n1696 9.3005
R21386 GND.n5879 GND.n5878 9.3005
R21387 GND.n1699 GND.n1697 9.3005
R21388 GND.n5874 GND.n5867 9.3005
R21389 GND.n5873 GND.n5872 9.3005
R21390 GND.n5871 GND.n1602 9.3005
R21391 GND.n6049 GND.n1603 9.3005
R21392 GND.n4343 GND.n4342 9.3005
R21393 GND.n4340 GND.n4330 9.3005
R21394 GND.n4339 GND.n4338 9.3005
R21395 GND.n4337 GND.n2112 9.3005
R21396 GND.n4366 GND.n2110 9.3005
R21397 GND.n4378 GND.n4377 9.3005
R21398 GND.n4376 GND.n2111 9.3005
R21399 GND.n4375 GND.n4374 9.3005
R21400 GND.n4373 GND.n2083 9.3005
R21401 GND.n4414 GND.n2081 9.3005
R21402 GND.n4421 GND.n4420 9.3005
R21403 GND.n4419 GND.n2082 9.3005
R21404 GND.n4418 GND.n4417 9.3005
R21405 GND.n2049 GND.n2047 9.3005
R21406 GND.n4460 GND.n4459 9.3005
R21407 GND.n4458 GND.n2048 9.3005
R21408 GND.n4457 GND.n4456 9.3005
R21409 GND.n4455 GND.n2021 9.3005
R21410 GND.n4496 GND.n2019 9.3005
R21411 GND.n4503 GND.n4502 9.3005
R21412 GND.n4501 GND.n2020 9.3005
R21413 GND.n4500 GND.n4499 9.3005
R21414 GND.n1987 GND.n1985 9.3005
R21415 GND.n4578 GND.n4577 9.3005
R21416 GND.n4576 GND.n1986 9.3005
R21417 GND.n4575 GND.n4574 9.3005
R21418 GND.n4573 GND.n1959 9.3005
R21419 GND.n4607 GND.n1955 9.3005
R21420 GND.n4610 GND.n4609 9.3005
R21421 GND.n4608 GND.n1958 9.3005
R21422 GND.n1957 GND.n1939 9.3005
R21423 GND.n1892 GND.n1890 9.3005
R21424 GND.n4682 GND.n4681 9.3005
R21425 GND.n4680 GND.n1891 9.3005
R21426 GND.n4679 GND.n4678 9.3005
R21427 GND.n4677 GND.n1895 9.3005
R21428 GND.n4676 GND.n4675 9.3005
R21429 GND.n4674 GND.n1899 9.3005
R21430 GND.n4673 GND.n4672 9.3005
R21431 GND.n4671 GND.n1903 9.3005
R21432 GND.n4670 GND.n4669 9.3005
R21433 GND.n4668 GND.n1907 9.3005
R21434 GND.n4667 GND.n4666 9.3005
R21435 GND.n1846 GND.n1844 9.3005
R21436 GND.n4737 GND.n4736 9.3005
R21437 GND.n4735 GND.n1845 9.3005
R21438 GND.n4734 GND.n4733 9.3005
R21439 GND.n4732 GND.n1819 9.3005
R21440 GND.n4762 GND.n1817 9.3005
R21441 GND.n4775 GND.n4774 9.3005
R21442 GND.n4773 GND.n1818 9.3005
R21443 GND.n4772 GND.n4771 9.3005
R21444 GND.n4770 GND.n4766 9.3005
R21445 GND.n1785 GND.n1783 9.3005
R21446 GND.n4843 GND.n4842 9.3005
R21447 GND.n4841 GND.n1784 9.3005
R21448 GND.n4840 GND.n4839 9.3005
R21449 GND.n4838 GND.n1758 9.3005
R21450 GND.n4868 GND.n1756 9.3005
R21451 GND.n4880 GND.n4879 9.3005
R21452 GND.n4878 GND.n1757 9.3005
R21453 GND.n4877 GND.n4876 9.3005
R21454 GND.n4875 GND.n1730 9.3005
R21455 GND.n4914 GND.n1726 9.3005
R21456 GND.n4918 GND.n4917 9.3005
R21457 GND.n4916 GND.n1729 9.3005
R21458 GND.n1728 GND.n1700 9.3005
R21459 GND.n5863 GND.n1698 9.3005
R21460 GND.n5878 GND.n5877 9.3005
R21461 GND.n5876 GND.n1699 9.3005
R21462 GND.n5875 GND.n5874 9.3005
R21463 GND.n5873 GND.n5866 9.3005
R21464 GND.n1604 GND.n1602 9.3005
R21465 GND.n6049 GND.n6048 9.3005
R21466 GND.n4342 GND.n4341 9.3005
R21467 GND.n4319 GND.n4318 9.3005
R21468 GND.n4320 GND.n2142 9.3005
R21469 GND.n4322 GND.n4321 9.3005
R21470 GND.n4323 GND.n2141 9.3005
R21471 GND.n4325 GND.n4324 9.3005
R21472 GND.n4326 GND.n2138 9.3005
R21473 GND.n4328 GND.n4327 9.3005
R21474 GND.n4317 GND.n2148 9.3005
R21475 GND.n4316 GND.n4315 9.3005
R21476 GND.n2119 GND.n2118 9.3005
R21477 GND.n4358 GND.n4357 9.3005
R21478 GND.n4359 GND.n2116 9.3005
R21479 GND.n4362 GND.n4361 9.3005
R21480 GND.n4360 GND.n2117 9.3005
R21481 GND.n2090 GND.n2089 9.3005
R21482 GND.n4394 GND.n4393 9.3005
R21483 GND.n4395 GND.n2087 9.3005
R21484 GND.n4410 GND.n4409 9.3005
R21485 GND.n4408 GND.n2088 9.3005
R21486 GND.n4407 GND.n4406 9.3005
R21487 GND.n4405 GND.n4396 9.3005
R21488 GND.n4404 GND.n4403 9.3005
R21489 GND.n4402 GND.n4401 9.3005
R21490 GND.n2027 GND.n2026 9.3005
R21491 GND.n4476 GND.n4475 9.3005
R21492 GND.n4477 GND.n2024 9.3005
R21493 GND.n4492 GND.n4491 9.3005
R21494 GND.n4490 GND.n2025 9.3005
R21495 GND.n4489 GND.n4488 9.3005
R21496 GND.n4487 GND.n4478 9.3005
R21497 GND.n4486 GND.n4485 9.3005
R21498 GND.n4484 GND.n4483 9.3005
R21499 GND.n1965 GND.n1964 9.3005
R21500 GND.n4594 GND.n4593 9.3005
R21501 GND.n4595 GND.n1962 9.3005
R21502 GND.n4603 GND.n4602 9.3005
R21503 GND.n4601 GND.n1963 9.3005
R21504 GND.n4600 GND.n4599 9.3005
R21505 GND.n4596 GND.n1935 9.3005
R21506 GND.n4626 GND.n1934 9.3005
R21507 GND.n4628 GND.n4627 9.3005
R21508 GND.n4629 GND.n1933 9.3005
R21509 GND.n4631 GND.n4630 9.3005
R21510 GND.n1918 GND.n1917 9.3005
R21511 GND.n4644 GND.n4643 9.3005
R21512 GND.n2150 GND.n2149 9.3005
R21513 GND.n6033 GND.n6032 8.72777
R21514 GND.n7672 GND.n7671 8.72777
R21515 GND.n8392 GND.n8322 8.72777
R21516 GND.n4259 GND.n4258 8.72777
R21517 GND.t89 GND.n4971 8.6605
R21518 GND.t72 GND.t104 8.6605
R21519 GND.n5840 GND.n4953 8.29966
R21520 GND.n8571 GND.n8570 8.17456
R21521 GND.n4645 GND.n71 8.17456
R21522 GND.n17 GND.n11 8.14595
R21523 GND.n28 GND.n22 8.14595
R21524 GND.n40 GND.n34 8.14595
R21525 GND.n52 GND.n46 8.14595
R21526 GND.n64 GND.n58 8.14595
R21527 GND.n6 GND.n0 8.14595
R21528 GND.n90 GND.n84 8.14595
R21529 GND.n101 GND.n95 8.14595
R21530 GND.n113 GND.n107 8.14595
R21531 GND.n125 GND.n119 8.14595
R21532 GND.n137 GND.n131 8.14595
R21533 GND.n149 GND.n143 8.14595
R21534 GND.n6004 GND.n6003 7.95202
R21535 GND.n795 GND.n767 7.95202
R21536 GND.n7635 GND.n7632 7.95202
R21537 GND.n8351 GND.n8348 7.95202
R21538 GND.n4222 GND.n4219 7.95202
R21539 GND.t108 GND.n2105 7.93883
R21540 GND.n4856 GND.t27 7.93883
R21541 GND.t118 GND.n4961 7.93883
R21542 GND.t54 GND.n4997 7.93883
R21543 GND.n5799 GND.n5798 7.93883
R21544 GND.n5439 GND.n5436 7.93883
R21545 GND.n5742 GND.n5741 7.93883
R21546 GND.n5496 GND.n5493 7.93883
R21547 GND.n5685 GND.n5684 7.93883
R21548 GND.n5552 GND.n5549 7.93883
R21549 GND.n5598 GND.t79 7.93883
R21550 GND.n5624 GND.n5623 7.93883
R21551 GND.t197 GND.n6321 7.93883
R21552 GND.n6369 GND.n1453 7.93883
R21553 GND.n6263 GND.n6237 7.93883
R21554 GND.n6592 GND.n1288 7.93883
R21555 GND.n6513 GND.n1365 7.93883
R21556 GND.n1391 GND.n1214 7.93883
R21557 GND.n6826 GND.n1160 7.93883
R21558 GND.t209 GND.n1110 7.93883
R21559 GND.n6905 GND.n6904 7.93883
R21560 GND.n1081 GND.t127 7.93883
R21561 GND.n7051 GND.n1008 7.93883
R21562 GND.n7087 GND.n983 7.93883
R21563 GND.n7177 GND.n935 7.93883
R21564 GND.n7211 GND.n7210 7.93883
R21565 GND.n873 GND.n863 7.93883
R21566 GND.n7313 GND.n848 7.93883
R21567 GND.n7441 GND.t170 7.93883
R21568 GND.n7861 GND.t2 7.93883
R21569 GND.n8247 GND.t43 7.93883
R21570 GND.n15 GND.n14 7.3702
R21571 GND.n26 GND.n25 7.3702
R21572 GND.n38 GND.n37 7.3702
R21573 GND.n50 GND.n49 7.3702
R21574 GND.n62 GND.n61 7.3702
R21575 GND.n4 GND.n3 7.3702
R21576 GND.n88 GND.n87 7.3702
R21577 GND.n99 GND.n98 7.3702
R21578 GND.n111 GND.n110 7.3702
R21579 GND.n123 GND.n122 7.3702
R21580 GND.n135 GND.n134 7.3702
R21581 GND.n147 GND.n146 7.3702
R21582 GND.n5820 GND.t121 7.21716
R21583 GND.n4315 GND.n2148 7.17626
R21584 GND.n5928 GND.n5923 7.17626
R21585 GND.n7710 GND.n7709 7.17626
R21586 GND.n8435 GND.n8434 7.17626
R21587 GND.n8450 GND.n356 7.17626
R21588 GND.n4299 GND.n4298 7.17626
R21589 GND.n33 GND.n21 6.79791
R21590 GND.n4345 GND.n2133 6.4955
R21591 GND.n4331 GND.n2121 6.4955
R21592 GND.n4355 GND.n2123 6.4955
R21593 GND.n4334 GND.n2114 6.4955
R21594 GND.n4364 GND.n2102 6.4955
R21595 GND.n4381 GND.n2105 6.4955
R21596 GND.n4367 GND.n2092 6.4955
R21597 GND.n4391 GND.n2094 6.4955
R21598 GND.n4370 GND.n2085 6.4955
R21599 GND.n4412 GND.n2073 6.4955
R21600 GND.n4424 GND.n2076 6.4955
R21601 GND.n4433 GND.n2063 6.4955
R21602 GND.n4432 GND.n2066 6.4955
R21603 GND.n4399 GND.n2039 6.4955
R21604 GND.n4463 GND.n2042 6.4955
R21605 GND.n2050 GND.n2029 6.4955
R21606 GND.n4473 GND.n2031 6.4955
R21607 GND.n4452 GND.n4451 6.4955
R21608 GND.n4494 GND.n2011 6.4955
R21609 GND.n4506 GND.n2014 6.4955
R21610 GND.n4515 GND.n2001 6.4955
R21611 GND.n4514 GND.n2004 6.4955
R21612 GND.n4481 GND.n1977 6.4955
R21613 GND.n4581 GND.n1980 6.4955
R21614 GND.n1988 GND.n1967 6.4955
R21615 GND.n4591 GND.n1969 6.4955
R21616 GND.n4570 GND.n4569 6.4955
R21617 GND.n4605 GND.n1947 6.4955
R21618 GND.n4613 GND.n1950 6.4955
R21619 GND.n4597 GND.n1940 6.4955
R21620 GND.n4621 GND.n1937 6.4955
R21621 GND.n4624 GND.n1882 6.4955
R21622 GND.n4685 GND.n1885 6.4955
R21623 GND.n1931 GND.n1930 6.4955
R21624 GND.n4633 GND.n1928 6.4955
R21625 GND.n4636 GND.n1920 6.4955
R21626 GND.n4641 GND.n1921 6.4955
R21627 GND.n1923 GND.n1914 6.4955
R21628 GND.n4652 GND.n1911 6.4955
R21629 GND.n4657 GND.n1909 6.4955
R21630 GND.n4660 GND.n1864 6.4955
R21631 GND.n4694 GND.n1866 6.4955
R21632 GND.n4705 GND.n1857 6.4955
R21633 GND.n4704 GND.n1836 6.4955
R21634 GND.n4740 GND.n1839 6.4955
R21635 GND.n1847 GND.n1827 6.4955
R21636 GND.n4729 GND.n1821 6.4955
R21637 GND.n4760 GND.n1809 6.4955
R21638 GND.n4778 GND.n1812 6.4955
R21639 GND.n4763 GND.n1799 6.4955
R21640 GND.n4788 GND.n1801 6.4955
R21641 GND.n4799 GND.n1792 6.4955
R21642 GND.n4798 GND.n1775 6.4955
R21643 GND.n4846 GND.n1778 6.4955
R21644 GND.n4832 GND.n4831 6.4955
R21645 GND.n4856 GND.n1767 6.4955
R21646 GND.n4835 GND.n1760 6.4955
R21647 GND.n4866 GND.n1748 6.4955
R21648 GND.n4883 GND.n1751 6.4955
R21649 GND.n4869 GND.n1738 6.4955
R21650 GND.n4893 GND.n1740 6.4955
R21651 GND.n4872 GND.n1732 6.4955
R21652 GND.n4912 GND.n1718 6.4955
R21653 GND.n4921 GND.n1721 6.4955
R21654 GND.n4930 GND.n1710 6.4955
R21655 GND.n4929 GND.n1702 6.4955
R21656 GND.n5861 GND.n5860 6.4955
R21657 GND.n5881 GND.n1693 6.4955
R21658 GND.n5864 GND.n1682 6.4955
R21659 GND.n5890 GND.n1684 6.4955
R21660 GND.n5869 GND.n1676 6.4955
R21661 GND.n5899 GND.n1607 6.4955
R21662 GND.n6046 GND.n1610 6.4955
R21663 GND.n5792 GND.n5014 6.4955
R21664 GND.n5022 GND.n5016 6.4955
R21665 GND.n5735 GND.n5089 6.4955
R21666 GND.n5097 GND.n5091 6.4955
R21667 GND.n5678 GND.n5165 6.4955
R21668 GND.n5173 GND.n5167 6.4955
R21669 GND.n5583 GND.n1535 6.4955
R21670 GND.n6150 GND.n1530 6.4955
R21671 GND.t195 GND.n1445 6.4955
R21672 GND.n6270 GND.n6199 6.4955
R21673 GND.n6600 GND.n1280 6.4955
R21674 GND.n6520 GND.n1358 6.4955
R21675 GND.n6679 GND.n1210 6.4955
R21676 GND.t213 GND.n6818 6.4955
R21677 GND.n6886 GND.n1101 6.4955
R21678 GND.n6735 GND.n1093 6.4955
R21679 GND.n7070 GND.n7069 6.4955
R21680 GND.n7077 GND.n7076 6.4955
R21681 GND.n7184 GND.n924 6.4955
R21682 GND.n925 GND.n920 6.4955
R21683 GND.n7308 GND.n859 6.4955
R21684 GND.n7320 GND.n852 6.4955
R21685 GND.n7737 GND.n658 6.4955
R21686 GND.n7754 GND.n647 6.4955
R21687 GND.n7747 GND.n650 6.4955
R21688 GND.n7764 GND.n637 6.4955
R21689 GND.n7741 GND.n639 6.4955
R21690 GND.n7774 GND.n631 6.4955
R21691 GND.n7791 GND.n619 6.4955
R21692 GND.n7778 GND.n622 6.4955
R21693 GND.n7801 GND.n609 6.4955
R21694 GND.n7784 GND.n611 6.4955
R21695 GND.n7815 GND.n603 6.4955
R21696 GND.n7826 GND.n592 6.4955
R21697 GND.n7809 GND.n595 6.4955
R21698 GND.n7834 GND.n585 6.4955
R21699 GND.n7837 GND.n582 6.4955
R21700 GND.n7853 GND.n570 6.4955
R21701 GND.n7846 GND.n573 6.4955
R21702 GND.n7861 GND.n564 6.4955
R21703 GND.n7869 GND.n558 6.4955
R21704 GND.n7891 GND.n536 6.4955
R21705 GND.n539 GND.n526 6.4955
R21706 GND.n7900 GND.n7899 6.4955
R21707 GND.n7882 GND.n529 6.4955
R21708 GND.n7944 GND.n505 6.4955
R21709 GND.n549 GND.n508 6.4955
R21710 GND.n7954 GND.n495 6.4955
R21711 GND.n7937 GND.n497 6.4955
R21712 GND.n7981 GND.n478 6.4955
R21713 GND.n7968 GND.n481 6.4955
R21714 GND.n7991 GND.n468 6.4955
R21715 GND.n7974 GND.n470 6.4955
R21716 GND.n8006 GND.n462 6.4955
R21717 GND.n8015 GND.n455 6.4955
R21718 GND.n8020 GND.n449 6.4955
R21719 GND.n451 GND.n441 6.4955
R21720 GND.n8033 GND.n8032 6.4955
R21721 GND.n8566 GND.n158 6.4955
R21722 GND.n435 GND.n160 6.4955
R21723 GND.n8125 GND.n8122 6.4955
R21724 GND.n8132 GND.n429 6.4955
R21725 GND.n8559 GND.n177 6.4955
R21726 GND.n8140 GND.n180 6.4955
R21727 GND.n8553 GND.n189 6.4955
R21728 GND.n8147 GND.n192 6.4955
R21729 GND.n8547 GND.n199 6.4955
R21730 GND.n8155 GND.n202 6.4955
R21731 GND.n8541 GND.n209 6.4955
R21732 GND.n8162 GND.n212 6.4955
R21733 GND.n8535 GND.n220 6.4955
R21734 GND.n8170 GND.n223 6.4955
R21735 GND.n8529 GND.n230 6.4955
R21736 GND.n8177 GND.n233 6.4955
R21737 GND.n8523 GND.n241 6.4955
R21738 GND.n8185 GND.n244 6.4955
R21739 GND.n8517 GND.n251 6.4955
R21740 GND.n8192 GND.n411 6.4955
R21741 GND.n8511 GND.n261 6.4955
R21742 GND.n8200 GND.n264 6.4955
R21743 GND.n8505 GND.n271 6.4955
R21744 GND.n8207 GND.n274 6.4955
R21745 GND.n8499 GND.n282 6.4955
R21746 GND.n8215 GND.n285 6.4955
R21747 GND.n8493 GND.n292 6.4955
R21748 GND.n8222 GND.n295 6.4955
R21749 GND.n8487 GND.n303 6.4955
R21750 GND.n8231 GND.n306 6.4955
R21751 GND.n8481 GND.n313 6.4955
R21752 GND.n8247 GND.n8246 6.4955
R21753 GND.n8475 GND.n323 6.4955
R21754 GND.n8240 GND.n326 6.4955
R21755 GND.n8469 GND.n333 6.4955
R21756 GND.n8456 GND.n336 6.4955
R21757 GND.n8463 GND.n343 6.4955
R21758 GND.n6074 GND.n6073 6.4005
R21759 GND.n6959 GND.n6958 6.4005
R21760 GND.n15 GND.n11 5.81868
R21761 GND.n26 GND.n22 5.81868
R21762 GND.n38 GND.n34 5.81868
R21763 GND.n50 GND.n46 5.81868
R21764 GND.n62 GND.n58 5.81868
R21765 GND.n4 GND.n0 5.81868
R21766 GND.n88 GND.n84 5.81868
R21767 GND.n99 GND.n95 5.81868
R21768 GND.n111 GND.n107 5.81868
R21769 GND.n123 GND.n119 5.81868
R21770 GND.n135 GND.n131 5.81868
R21771 GND.n147 GND.n143 5.81868
R21772 GND.n70 GND.n10 5.80869
R21773 GND.n5813 GND.t86 5.77383
R21774 GND.n7425 GND.t112 5.77383
R21775 GND.n103 GND.n91 5.75912
R21776 GND.n33 GND.n32 5.74619
R21777 GND.n45 GND.n44 5.74619
R21778 GND.n57 GND.n56 5.74619
R21779 GND.n69 GND.n68 5.74619
R21780 GND.n7593 GND.t161 5.413
R21781 GND.n71 GND.n70 5.34331
R21782 GND.n8571 GND.n151 5.34331
R21783 GND.n790 GND.n767 5.23686
R21784 GND.n4605 GND.t6 5.05216
R21785 GND.n4750 GND.t14 5.05216
R21786 GND.t121 GND.n5819 5.05216
R21787 GND.t86 GND.n5812 5.05216
R21788 GND.n5426 GND.n5423 5.05216
R21789 GND.n5785 GND.n5784 5.05216
R21790 GND.n5483 GND.n5480 5.05216
R21791 GND.n5728 GND.n5727 5.05216
R21792 GND.n5539 GND.n5536 5.05216
R21793 GND.n5671 GND.n5670 5.05216
R21794 GND.n6117 GND.t25 5.05216
R21795 GND.n6142 GND.n1546 5.05216
R21796 GND.n6157 GND.n1531 5.05216
R21797 GND.n6277 GND.n6192 5.05216
R21798 GND.n6384 GND.n1437 5.05216
R21799 GND.n6527 GND.n1351 5.05216
R21800 GND.n6608 GND.n1272 5.05216
R21801 GND.n6672 GND.n1209 5.05216
R21802 GND.n6460 GND.n1170 5.05216
R21803 GND.n6767 GND.n6741 5.05216
R21804 GND.n6895 GND.n6894 5.05216
R21805 GND.n6992 GND.t13 5.05216
R21806 GND.n1009 GND.n1003 5.05216
R21807 GND.n999 GND.n989 5.05216
R21808 GND.n7185 GND.n929 5.05216
R21809 GND.n7204 GND.n7203 5.05216
R21810 GND.n7301 GND.n857 5.05216
R21811 GND.n7327 GND.n846 5.05216
R21812 GND.n7964 GND.t176 5.05216
R21813 GND.n8155 GND.t4 5.05216
R21814 GND.n151 GND.n150 4.7699
R21815 GND.n6087 GND.n6086 4.74817
R21816 GND.n6084 GND.n6083 4.74817
R21817 GND.n6081 GND.n6080 4.74817
R21818 GND.n6078 GND.n6077 4.74817
R21819 GND.n6075 GND.n6074 4.74817
R21820 GND.n6936 GND.n6935 4.74817
R21821 GND.n6938 GND.n1072 4.74817
R21822 GND.n6947 GND.n6946 4.74817
R21823 GND.n6948 GND.n1070 4.74817
R21824 GND.n6959 GND.n6955 4.74817
R21825 GND.n699 GND.n663 4.74817
R21826 GND.n7728 GND.n665 4.74817
R21827 GND.n669 GND.n665 4.74817
R21828 GND.n702 GND.n663 4.74817
R21829 GND.n698 GND.n662 4.74817
R21830 GND.n6937 GND.n6936 4.74817
R21831 GND.n6939 GND.n6938 4.74817
R21832 GND.n6946 GND.n6945 4.74817
R21833 GND.n6949 GND.n6948 4.74817
R21834 GND.n6955 GND.n6954 4.74817
R21835 GND.n7987 GND.n172 4.74817
R21836 GND.n170 GND.n164 4.74817
R21837 GND.n8563 GND.n165 4.74817
R21838 GND.n173 GND.n169 4.74817
R21839 GND.n454 GND.n172 4.74817
R21840 GND.n8017 GND.n170 4.74817
R21841 GND.n8564 GND.n8563 4.74817
R21842 GND.n8123 GND.n169 4.74817
R21843 GND.n4559 GND.n4558 4.74817
R21844 GND.n4553 GND.n4539 4.74817
R21845 GND.n4551 GND.n4550 4.74817
R21846 GND.n4546 GND.n4542 4.74817
R21847 GND.n4544 GND.n4543 4.74817
R21848 GND.n7926 GND.n7925 4.74817
R21849 GND.n7921 GND.n7920 4.74817
R21850 GND.n8036 GND.n438 4.74817
R21851 GND.n8120 GND.n8038 4.74817
R21852 GND.n8118 GND.n8117 4.74817
R21853 GND.n7927 GND.n7926 4.74817
R21854 GND.n7922 GND.n7921 4.74817
R21855 GND.n440 GND.n438 4.74817
R21856 GND.n8038 GND.n8037 4.74817
R21857 GND.n8119 GND.n8118 4.74817
R21858 GND.n4688 GND.n4687 4.74817
R21859 GND.n4639 GND.n1876 4.74817
R21860 GND.n4654 GND.n1875 4.74817
R21861 GND.n1874 GND.n1870 4.74817
R21862 GND.n4688 GND.n1878 4.74817
R21863 GND.n1927 GND.n1876 4.74817
R21864 GND.n4638 GND.n1875 4.74817
R21865 GND.n4655 GND.n1874 4.74817
R21866 GND.n4558 GND.n4557 4.74817
R21867 GND.n4539 GND.n4537 4.74817
R21868 GND.n4552 GND.n4551 4.74817
R21869 GND.n4542 GND.n4540 4.74817
R21870 GND.n4545 GND.n4544 4.74817
R21871 GND.n1625 GND.n1596 4.74817
R21872 GND.n1626 GND.n1597 4.74817
R21873 GND.n1631 GND.n1598 4.74817
R21874 GND.n1630 GND.n1597 4.74817
R21875 GND.n1634 GND.n1598 4.74817
R21876 GND.n6076 GND.n6075 4.74817
R21877 GND.n6079 GND.n6078 4.74817
R21878 GND.n6082 GND.n6081 4.74817
R21879 GND.n6085 GND.n6084 4.74817
R21880 GND.n6088 GND.n6087 4.74817
R21881 GND.n103 GND.n102 4.7074
R21882 GND.n115 GND.n114 4.7074
R21883 GND.n127 GND.n126 4.7074
R21884 GND.n139 GND.n138 4.7074
R21885 GND.n7682 GND.n7598 4.6132
R21886 GND.n5959 GND.n1658 4.6132
R21887 GND.n5274 GND.n5273 4.38232
R21888 GND.n794 GND.n793 4.38232
R21889 GND.n80 GND.n75 4.17239
R21890 GND.n5953 GND.n1663 4.07323
R21891 GND.n7690 GND.n7689 4.07323
R21892 GND.n8414 GND.n8411 4.07323
R21893 GND.n4279 GND.n4278 4.07323
R21894 GND.n5417 GND.n4999 3.60883
R21895 GND.n5778 GND.n5032 3.60883
R21896 GND.n5080 GND.n5074 3.60883
R21897 GND.n5721 GND.n5107 3.60883
R21898 GND.n5155 GND.n5154 3.60883
R21899 GND.n5664 GND.n5183 3.60883
R21900 GND.n6125 GND.n1555 3.60883
R21901 GND.n5611 GND.n1505 3.60883
R21902 GND.n6284 GND.n6185 3.60883
R21903 GND.n6394 GND.n1428 3.60883
R21904 GND.n6534 GND.t201 3.60883
R21905 GND.t207 GND.n1264 3.60883
R21906 GND.n6664 GND.n1225 3.60883
R21907 GND.n6810 GND.n6809 3.60883
R21908 GND.n6774 GND.n6710 3.60883
R21909 GND.n6979 GND.n1055 3.60883
R21910 GND.n7052 GND.n1013 3.60883
R21911 GND.n7094 GND.n985 3.60883
R21912 GND.n7170 GND.n933 3.60883
R21913 GND.n916 GND.n907 3.60883
R21914 GND.n7291 GND.n7290 3.60883
R21915 GND.n7336 GND.n7335 3.60883
R21916 GND.n80 GND.n79 3.60163
R21917 GND.n16 GND.n12 3.44771
R21918 GND.n27 GND.n23 3.44771
R21919 GND.n39 GND.n35 3.44771
R21920 GND.n51 GND.n47 3.44771
R21921 GND.n63 GND.n59 3.44771
R21922 GND.n5 GND.n1 3.44771
R21923 GND.n89 GND.n85 3.44771
R21924 GND.n100 GND.n96 3.44771
R21925 GND.n112 GND.n108 3.44771
R21926 GND.n124 GND.n120 3.44771
R21927 GND.n136 GND.n132 3.44771
R21928 GND.n148 GND.n144 3.44771
R21929 GND.n7731 GND.n7730 3.35648
R21930 GND.n6051 GND.n1600 3.35648
R21931 GND.n5417 GND.t72 2.88717
R21932 GND.n7528 GND.t161 2.88717
R21933 GND.n7730 GND.n7729 2.59004
R21934 GND.n1640 GND.n1600 2.59004
R21935 GND.n6101 GND.n6100 2.52633
R21936 GND.n7019 GND.n1031 2.52633
R21937 GND.n5950 GND.n1663 2.52171
R21938 GND.n7691 GND.n7690 2.52171
R21939 GND.n8415 GND.n8414 2.52171
R21940 GND.n4280 GND.n4279 2.52171
R21941 GND.n7731 GND.n665 2.27742
R21942 GND.n7731 GND.n663 2.27742
R21943 GND.n7731 GND.n662 2.27742
R21944 GND.n6936 GND.n661 2.27742
R21945 GND.n6938 GND.n661 2.27742
R21946 GND.n6946 GND.n661 2.27742
R21947 GND.n6948 GND.n661 2.27742
R21948 GND.n6955 GND.n661 2.27742
R21949 GND.n8562 GND.n172 2.27742
R21950 GND.n8562 GND.n170 2.27742
R21951 GND.n8563 GND.n8562 2.27742
R21952 GND.n8562 GND.n169 2.27742
R21953 GND.n7926 GND.n168 2.27742
R21954 GND.n7921 GND.n168 2.27742
R21955 GND.n438 GND.n168 2.27742
R21956 GND.n8038 GND.n168 2.27742
R21957 GND.n8118 GND.n168 2.27742
R21958 GND.n4689 GND.n4688 2.27742
R21959 GND.n4689 GND.n1876 2.27742
R21960 GND.n4689 GND.n1875 2.27742
R21961 GND.n4689 GND.n1874 2.27742
R21962 GND.n4558 GND.n1873 2.27742
R21963 GND.n4539 GND.n1873 2.27742
R21964 GND.n4551 GND.n1873 2.27742
R21965 GND.n4542 GND.n1873 2.27742
R21966 GND.n4544 GND.n1873 2.27742
R21967 GND.n6051 GND.n1596 2.27742
R21968 GND.n6051 GND.n1597 2.27742
R21969 GND.n6051 GND.n1598 2.27742
R21970 GND.n6075 GND.n6052 2.27742
R21971 GND.n6078 GND.n6052 2.27742
R21972 GND.n6081 GND.n6052 2.27742
R21973 GND.n6084 GND.n6052 2.27742
R21974 GND.n6087 GND.n6052 2.27742
R21975 GND GND.n71 2.20449
R21976 GND.n5390 GND.t173 2.1655
R21977 GND.n5390 GND.n4969 2.1655
R21978 GND.n5412 GND.n5409 2.1655
R21979 GND.n5771 GND.n5770 2.1655
R21980 GND.n5469 GND.n5464 2.1655
R21981 GND.n5714 GND.n5713 2.1655
R21982 GND.n5526 GND.n5521 2.1655
R21983 GND.n5657 GND.n5656 2.1655
R21984 GND.n6117 GND.n1562 2.1655
R21985 GND.n6313 GND.n6312 2.1655
R21986 GND.n6291 GND.n6178 2.1655
R21987 GND.n6404 GND.n1422 2.1655
R21988 GND.n6541 GND.n1339 2.1655
R21989 GND.n6623 GND.n1256 2.1655
R21990 GND.n6647 GND.n1234 2.1655
R21991 GND.n6803 GND.n6802 2.1655
R21992 GND.n6781 GND.n1203 2.1655
R21993 GND.n6993 GND.n6992 2.1655
R21994 GND.n7038 GND.n1017 2.1655
R21995 GND.n7112 GND.n972 2.1655
R21996 GND.n7151 GND.n7150 2.1655
R21997 GND.n7246 GND.n903 2.1655
R21998 GND.n883 GND.n877 2.1655
R21999 GND.n7350 GND.n830 2.1655
R22000 GND.t63 GND.n812 2.1655
R22001 GND.n808 GND.n798 2.1655
R22002 GND.n21 GND.n19 2.07809
R22003 GND.n32 GND.n30 2.07809
R22004 GND.n44 GND.n42 2.07809
R22005 GND.n56 GND.n54 2.07809
R22006 GND.n68 GND.n66 2.07809
R22007 GND.n10 GND.n8 2.07809
R22008 GND.n91 GND.n83 2.07809
R22009 GND.n102 GND.n94 2.07809
R22010 GND.n114 GND.n106 2.07809
R22011 GND.n126 GND.n118 2.07809
R22012 GND.n138 GND.n130 2.07809
R22013 GND.n150 GND.n142 2.07809
R22014 GND.n8572 GND.n8571 1.64989
R22015 GND.n70 GND.n69 1.59317
R22016 GND.n151 GND.n139 1.59317
R22017 GND.n4451 GND.t16 1.44383
R22018 GND.n4728 GND.t14 1.44383
R22019 GND.n5631 GND.t79 1.44383
R22020 GND.n6554 GND.t11 1.44383
R22021 GND.t24 GND.n1240 1.44383
R22022 GND.t127 GND.n1045 1.44383
R22023 GND.t140 GND.n834 1.44383
R22024 GND.n7936 GND.t176 1.44383
R22025 GND.n411 GND.t18 1.44383
R22026 GND.n7379 GND.n7374 1.24928
R22027 GND.n5342 GND.n5341 1.24928
R22028 GND.n5320 GND.n5234 1.24928
R22029 GND.n7549 GND.n7548 1.24928
R22030 GND.n45 GND.n33 1.05222
R22031 GND.n57 GND.n45 1.05222
R22032 GND.n69 GND.n57 1.05222
R22033 GND.n115 GND.n103 1.05222
R22034 GND.n127 GND.n115 1.05222
R22035 GND.n139 GND.n127 1.05222
R22036 GND.n73 GND.n72 1.01794
R22037 GND.n74 GND.n73 1.01794
R22038 GND.n75 GND.n74 1.01794
R22039 GND.n77 GND.n76 1.01794
R22040 GND.n78 GND.n77 1.01794
R22041 GND.n79 GND.n78 1.01794
R22042 GND.n6039 GND.n1658 0.776258
R22043 GND.n7682 GND.n7681 0.776258
R22044 GND.n5399 GND.n5396 0.722166
R22045 GND.n4987 GND.n4981 0.722166
R22046 GND.n5764 GND.n5050 0.722166
R22047 GND.n5757 GND.n5058 0.722166
R22048 GND.n5741 GND.t12 0.722166
R22049 GND.n5707 GND.n5125 0.722166
R22050 GND.n5700 GND.n5133 0.722166
R22051 GND.n5691 GND.t235 0.722166
R22052 GND.n6101 GND.n1575 0.722166
R22053 GND.n6109 GND.n1569 0.722166
R22054 GND.n6306 GND.n6305 0.722166
R22055 GND.n6298 GND.t205 0.722166
R22056 GND.n1329 GND.n1323 0.722166
R22057 GND.n6548 GND.n1335 0.722166
R22058 GND.n6631 GND.n1248 0.722166
R22059 GND.n6639 GND.n1242 0.722166
R22060 GND.n6795 GND.t203 0.722166
R22061 GND.n6789 GND.n6788 0.722166
R22062 GND.n7000 GND.n1037 0.722166
R22063 GND.n7019 GND.n7018 0.722166
R22064 GND.t23 GND.n984 0.722166
R22065 GND.n7126 GND.n7125 0.722166
R22066 GND.n959 GND.n953 0.722166
R22067 GND.n7211 GND.t10 0.722166
R22068 GND.n7252 GND.n891 0.722166
R22069 GND.n7266 GND.n887 0.722166
R22070 GND.n7361 GND.n7360 0.722166
R22071 GND.n7435 GND.n812 0.722166
R22072 GND.n5256 GND.n5254 0.716017
R22073 GND.n788 GND.n786 0.716017
R22074 GND.n7731 GND.n661 0.683383
R22075 GND.n6052 GND.n6051 0.683383
R22076 GND.n6917 GND.n6916 0.515744
R22077 GND.n5594 GND.n1588 0.515744
R22078 GND.n6112 GND.n1565 0.515744
R22079 GND.n6969 GND.n6968 0.515744
R22080 GND.n8452 GND.n8451 0.482207
R22081 GND.n4316 GND.n2150 0.482207
R22082 GND.n3933 GND.n2246 0.459342
R22083 GND.n2969 GND.n2968 0.459342
R22084 GND.n8262 GND.n8261 0.459342
R22085 GND.n4125 GND.n4124 0.459342
R22086 GND.n8562 GND.n168 0.449125
R22087 GND.n4689 GND.n1873 0.449125
R22088 GND.n8293 GND.n341 0.419707
R22089 GND.n709 GND.n644 0.419707
R22090 GND.n5904 GND.n5903 0.419707
R22091 GND.n4348 GND.n2128 0.419707
R22092 GND.n7596 GND.n735 0.312695
R22093 GND.n5232 GND.n5231 0.312695
R22094 GND.n5329 GND.n5232 0.312695
R22095 GND.n7596 GND.n736 0.312695
R22096 GND.n366 GND.n349 0.299281
R22097 GND.n4329 GND.n4328 0.299281
R22098 GND GND.n8572 0.279758
R22099 GND.n6051 GND.n1595 0.245927
R22100 GND.n7732 GND.n7731 0.245927
R22101 GND.n8572 GND.n80 0.240827
R22102 GND.n8346 GND.n349 0.23678
R22103 GND.n7630 GND.n660 0.23678
R22104 GND.n4329 GND.n2137 0.23678
R22105 GND.n6050 GND.n1601 0.23678
R22106 GND.n7598 GND.n734 0.229039
R22107 GND.n7599 GND.n7598 0.229039
R22108 GND.n5959 GND.n5958 0.229039
R22109 GND.n6038 GND.n5959 0.229039
R22110 GND.n6073 GND.n6072 0.194439
R22111 GND.n6958 GND.n1068 0.194439
R22112 GND.n4647 GND.n4646 0.152939
R22113 GND.n4648 GND.n4647 0.152939
R22114 GND.n4648 GND.n1861 0.152939
R22115 GND.n4697 GND.n1861 0.152939
R22116 GND.n4698 GND.n4697 0.152939
R22117 GND.n4699 GND.n4698 0.152939
R22118 GND.n4700 GND.n4699 0.152939
R22119 GND.n4700 GND.n1824 0.152939
R22120 GND.n4753 GND.n1824 0.152939
R22121 GND.n4754 GND.n4753 0.152939
R22122 GND.n4755 GND.n4754 0.152939
R22123 GND.n4756 GND.n4755 0.152939
R22124 GND.n4756 GND.n1796 0.152939
R22125 GND.n4791 GND.n1796 0.152939
R22126 GND.n4792 GND.n4791 0.152939
R22127 GND.n4793 GND.n4792 0.152939
R22128 GND.n4794 GND.n4793 0.152939
R22129 GND.n4794 GND.n1763 0.152939
R22130 GND.n4859 GND.n1763 0.152939
R22131 GND.n4860 GND.n4859 0.152939
R22132 GND.n4861 GND.n4860 0.152939
R22133 GND.n4862 GND.n4861 0.152939
R22134 GND.n4862 GND.n1735 0.152939
R22135 GND.n4896 GND.n1735 0.152939
R22136 GND.n4897 GND.n4896 0.152939
R22137 GND.n4898 GND.n4897 0.152939
R22138 GND.n4899 GND.n4898 0.152939
R22139 GND.n4900 GND.n4899 0.152939
R22140 GND.n4901 GND.n4900 0.152939
R22141 GND.n4902 GND.n4901 0.152939
R22142 GND.n4903 GND.n4902 0.152939
R22143 GND.n4903 GND.n1679 0.152939
R22144 GND.n5893 GND.n1679 0.152939
R22145 GND.n5894 GND.n5893 0.152939
R22146 GND.n5895 GND.n5894 0.152939
R22147 GND.n5895 GND.n1595 0.152939
R22148 GND.n3933 GND.n3932 0.152939
R22149 GND.n3932 GND.n3931 0.152939
R22150 GND.n3931 GND.n2252 0.152939
R22151 GND.n2257 GND.n2252 0.152939
R22152 GND.n2258 GND.n2257 0.152939
R22153 GND.n2259 GND.n2258 0.152939
R22154 GND.n2264 GND.n2259 0.152939
R22155 GND.n2265 GND.n2264 0.152939
R22156 GND.n2266 GND.n2265 0.152939
R22157 GND.n2267 GND.n2266 0.152939
R22158 GND.n2272 GND.n2267 0.152939
R22159 GND.n2273 GND.n2272 0.152939
R22160 GND.n2274 GND.n2273 0.152939
R22161 GND.n2275 GND.n2274 0.152939
R22162 GND.n2280 GND.n2275 0.152939
R22163 GND.n2281 GND.n2280 0.152939
R22164 GND.n2282 GND.n2281 0.152939
R22165 GND.n2283 GND.n2282 0.152939
R22166 GND.n2288 GND.n2283 0.152939
R22167 GND.n2289 GND.n2288 0.152939
R22168 GND.n2290 GND.n2289 0.152939
R22169 GND.n2291 GND.n2290 0.152939
R22170 GND.n2296 GND.n2291 0.152939
R22171 GND.n2297 GND.n2296 0.152939
R22172 GND.n2298 GND.n2297 0.152939
R22173 GND.n2299 GND.n2298 0.152939
R22174 GND.n2304 GND.n2299 0.152939
R22175 GND.n2305 GND.n2304 0.152939
R22176 GND.n2306 GND.n2305 0.152939
R22177 GND.n2307 GND.n2306 0.152939
R22178 GND.n2312 GND.n2307 0.152939
R22179 GND.n2313 GND.n2312 0.152939
R22180 GND.n2314 GND.n2313 0.152939
R22181 GND.n2315 GND.n2314 0.152939
R22182 GND.n2320 GND.n2315 0.152939
R22183 GND.n2321 GND.n2320 0.152939
R22184 GND.n2322 GND.n2321 0.152939
R22185 GND.n2323 GND.n2322 0.152939
R22186 GND.n2328 GND.n2323 0.152939
R22187 GND.n2329 GND.n2328 0.152939
R22188 GND.n2330 GND.n2329 0.152939
R22189 GND.n2331 GND.n2330 0.152939
R22190 GND.n2336 GND.n2331 0.152939
R22191 GND.n2337 GND.n2336 0.152939
R22192 GND.n2338 GND.n2337 0.152939
R22193 GND.n2339 GND.n2338 0.152939
R22194 GND.n2344 GND.n2339 0.152939
R22195 GND.n2345 GND.n2344 0.152939
R22196 GND.n2346 GND.n2345 0.152939
R22197 GND.n2347 GND.n2346 0.152939
R22198 GND.n2352 GND.n2347 0.152939
R22199 GND.n2353 GND.n2352 0.152939
R22200 GND.n2354 GND.n2353 0.152939
R22201 GND.n2355 GND.n2354 0.152939
R22202 GND.n2360 GND.n2355 0.152939
R22203 GND.n2361 GND.n2360 0.152939
R22204 GND.n2362 GND.n2361 0.152939
R22205 GND.n2363 GND.n2362 0.152939
R22206 GND.n2368 GND.n2363 0.152939
R22207 GND.n2369 GND.n2368 0.152939
R22208 GND.n2370 GND.n2369 0.152939
R22209 GND.n2371 GND.n2370 0.152939
R22210 GND.n2376 GND.n2371 0.152939
R22211 GND.n2377 GND.n2376 0.152939
R22212 GND.n2378 GND.n2377 0.152939
R22213 GND.n2379 GND.n2378 0.152939
R22214 GND.n2384 GND.n2379 0.152939
R22215 GND.n2385 GND.n2384 0.152939
R22216 GND.n2386 GND.n2385 0.152939
R22217 GND.n2387 GND.n2386 0.152939
R22218 GND.n2392 GND.n2387 0.152939
R22219 GND.n2393 GND.n2392 0.152939
R22220 GND.n2394 GND.n2393 0.152939
R22221 GND.n2395 GND.n2394 0.152939
R22222 GND.n2400 GND.n2395 0.152939
R22223 GND.n2401 GND.n2400 0.152939
R22224 GND.n2402 GND.n2401 0.152939
R22225 GND.n2403 GND.n2402 0.152939
R22226 GND.n2408 GND.n2403 0.152939
R22227 GND.n2409 GND.n2408 0.152939
R22228 GND.n2410 GND.n2409 0.152939
R22229 GND.n2411 GND.n2410 0.152939
R22230 GND.n2416 GND.n2411 0.152939
R22231 GND.n2417 GND.n2416 0.152939
R22232 GND.n2418 GND.n2417 0.152939
R22233 GND.n2419 GND.n2418 0.152939
R22234 GND.n2424 GND.n2419 0.152939
R22235 GND.n2425 GND.n2424 0.152939
R22236 GND.n2426 GND.n2425 0.152939
R22237 GND.n2427 GND.n2426 0.152939
R22238 GND.n2432 GND.n2427 0.152939
R22239 GND.n2433 GND.n2432 0.152939
R22240 GND.n2434 GND.n2433 0.152939
R22241 GND.n2435 GND.n2434 0.152939
R22242 GND.n2440 GND.n2435 0.152939
R22243 GND.n2441 GND.n2440 0.152939
R22244 GND.n2442 GND.n2441 0.152939
R22245 GND.n2443 GND.n2442 0.152939
R22246 GND.n2448 GND.n2443 0.152939
R22247 GND.n2449 GND.n2448 0.152939
R22248 GND.n2450 GND.n2449 0.152939
R22249 GND.n2451 GND.n2450 0.152939
R22250 GND.n2456 GND.n2451 0.152939
R22251 GND.n2457 GND.n2456 0.152939
R22252 GND.n2458 GND.n2457 0.152939
R22253 GND.n2459 GND.n2458 0.152939
R22254 GND.n2464 GND.n2459 0.152939
R22255 GND.n2465 GND.n2464 0.152939
R22256 GND.n2466 GND.n2465 0.152939
R22257 GND.n2467 GND.n2466 0.152939
R22258 GND.n2472 GND.n2467 0.152939
R22259 GND.n2473 GND.n2472 0.152939
R22260 GND.n2474 GND.n2473 0.152939
R22261 GND.n2475 GND.n2474 0.152939
R22262 GND.n2480 GND.n2475 0.152939
R22263 GND.n2481 GND.n2480 0.152939
R22264 GND.n2482 GND.n2481 0.152939
R22265 GND.n2483 GND.n2482 0.152939
R22266 GND.n2488 GND.n2483 0.152939
R22267 GND.n2489 GND.n2488 0.152939
R22268 GND.n2490 GND.n2489 0.152939
R22269 GND.n2491 GND.n2490 0.152939
R22270 GND.n2496 GND.n2491 0.152939
R22271 GND.n2497 GND.n2496 0.152939
R22272 GND.n2498 GND.n2497 0.152939
R22273 GND.n2499 GND.n2498 0.152939
R22274 GND.n2504 GND.n2499 0.152939
R22275 GND.n2505 GND.n2504 0.152939
R22276 GND.n2506 GND.n2505 0.152939
R22277 GND.n2507 GND.n2506 0.152939
R22278 GND.n2512 GND.n2507 0.152939
R22279 GND.n2513 GND.n2512 0.152939
R22280 GND.n2514 GND.n2513 0.152939
R22281 GND.n2515 GND.n2514 0.152939
R22282 GND.n2520 GND.n2515 0.152939
R22283 GND.n2521 GND.n2520 0.152939
R22284 GND.n2522 GND.n2521 0.152939
R22285 GND.n2523 GND.n2522 0.152939
R22286 GND.n2528 GND.n2523 0.152939
R22287 GND.n2529 GND.n2528 0.152939
R22288 GND.n2530 GND.n2529 0.152939
R22289 GND.n2531 GND.n2530 0.152939
R22290 GND.n2536 GND.n2531 0.152939
R22291 GND.n2537 GND.n2536 0.152939
R22292 GND.n2538 GND.n2537 0.152939
R22293 GND.n2539 GND.n2538 0.152939
R22294 GND.n2544 GND.n2539 0.152939
R22295 GND.n2545 GND.n2544 0.152939
R22296 GND.n2546 GND.n2545 0.152939
R22297 GND.n2547 GND.n2546 0.152939
R22298 GND.n2552 GND.n2547 0.152939
R22299 GND.n2553 GND.n2552 0.152939
R22300 GND.n2554 GND.n2553 0.152939
R22301 GND.n2555 GND.n2554 0.152939
R22302 GND.n2560 GND.n2555 0.152939
R22303 GND.n2561 GND.n2560 0.152939
R22304 GND.n2562 GND.n2561 0.152939
R22305 GND.n2563 GND.n2562 0.152939
R22306 GND.n2568 GND.n2563 0.152939
R22307 GND.n2569 GND.n2568 0.152939
R22308 GND.n2570 GND.n2569 0.152939
R22309 GND.n2571 GND.n2570 0.152939
R22310 GND.n2576 GND.n2571 0.152939
R22311 GND.n2577 GND.n2576 0.152939
R22312 GND.n2578 GND.n2577 0.152939
R22313 GND.n2579 GND.n2578 0.152939
R22314 GND.n2584 GND.n2579 0.152939
R22315 GND.n2585 GND.n2584 0.152939
R22316 GND.n2586 GND.n2585 0.152939
R22317 GND.n2587 GND.n2586 0.152939
R22318 GND.n2592 GND.n2587 0.152939
R22319 GND.n2593 GND.n2592 0.152939
R22320 GND.n2594 GND.n2593 0.152939
R22321 GND.n2595 GND.n2594 0.152939
R22322 GND.n2600 GND.n2595 0.152939
R22323 GND.n2601 GND.n2600 0.152939
R22324 GND.n2602 GND.n2601 0.152939
R22325 GND.n2603 GND.n2602 0.152939
R22326 GND.n2608 GND.n2603 0.152939
R22327 GND.n2609 GND.n2608 0.152939
R22328 GND.n2610 GND.n2609 0.152939
R22329 GND.n2611 GND.n2610 0.152939
R22330 GND.n2616 GND.n2611 0.152939
R22331 GND.n2617 GND.n2616 0.152939
R22332 GND.n2618 GND.n2617 0.152939
R22333 GND.n2619 GND.n2618 0.152939
R22334 GND.n2624 GND.n2619 0.152939
R22335 GND.n2625 GND.n2624 0.152939
R22336 GND.n2626 GND.n2625 0.152939
R22337 GND.n2627 GND.n2626 0.152939
R22338 GND.n2632 GND.n2627 0.152939
R22339 GND.n2633 GND.n2632 0.152939
R22340 GND.n2634 GND.n2633 0.152939
R22341 GND.n2635 GND.n2634 0.152939
R22342 GND.n2640 GND.n2635 0.152939
R22343 GND.n2641 GND.n2640 0.152939
R22344 GND.n2642 GND.n2641 0.152939
R22345 GND.n2643 GND.n2642 0.152939
R22346 GND.n2648 GND.n2643 0.152939
R22347 GND.n2649 GND.n2648 0.152939
R22348 GND.n2650 GND.n2649 0.152939
R22349 GND.n2651 GND.n2650 0.152939
R22350 GND.n2656 GND.n2651 0.152939
R22351 GND.n2657 GND.n2656 0.152939
R22352 GND.n2658 GND.n2657 0.152939
R22353 GND.n2659 GND.n2658 0.152939
R22354 GND.n2664 GND.n2659 0.152939
R22355 GND.n2665 GND.n2664 0.152939
R22356 GND.n2666 GND.n2665 0.152939
R22357 GND.n2667 GND.n2666 0.152939
R22358 GND.n2672 GND.n2667 0.152939
R22359 GND.n2673 GND.n2672 0.152939
R22360 GND.n2674 GND.n2673 0.152939
R22361 GND.n2675 GND.n2674 0.152939
R22362 GND.n2680 GND.n2675 0.152939
R22363 GND.n2681 GND.n2680 0.152939
R22364 GND.n2682 GND.n2681 0.152939
R22365 GND.n2683 GND.n2682 0.152939
R22366 GND.n2688 GND.n2683 0.152939
R22367 GND.n2689 GND.n2688 0.152939
R22368 GND.n2690 GND.n2689 0.152939
R22369 GND.n2691 GND.n2690 0.152939
R22370 GND.n2696 GND.n2691 0.152939
R22371 GND.n2697 GND.n2696 0.152939
R22372 GND.n2698 GND.n2697 0.152939
R22373 GND.n2699 GND.n2698 0.152939
R22374 GND.n2704 GND.n2699 0.152939
R22375 GND.n2705 GND.n2704 0.152939
R22376 GND.n2706 GND.n2705 0.152939
R22377 GND.n2707 GND.n2706 0.152939
R22378 GND.n2712 GND.n2707 0.152939
R22379 GND.n2713 GND.n2712 0.152939
R22380 GND.n2714 GND.n2713 0.152939
R22381 GND.n2715 GND.n2714 0.152939
R22382 GND.n2720 GND.n2715 0.152939
R22383 GND.n2721 GND.n2720 0.152939
R22384 GND.n2722 GND.n2721 0.152939
R22385 GND.n2723 GND.n2722 0.152939
R22386 GND.n2728 GND.n2723 0.152939
R22387 GND.n2729 GND.n2728 0.152939
R22388 GND.n2730 GND.n2729 0.152939
R22389 GND.n2731 GND.n2730 0.152939
R22390 GND.n2736 GND.n2731 0.152939
R22391 GND.n2737 GND.n2736 0.152939
R22392 GND.n2738 GND.n2737 0.152939
R22393 GND.n2739 GND.n2738 0.152939
R22394 GND.n2744 GND.n2739 0.152939
R22395 GND.n2745 GND.n2744 0.152939
R22396 GND.n2746 GND.n2745 0.152939
R22397 GND.n2747 GND.n2746 0.152939
R22398 GND.n2752 GND.n2747 0.152939
R22399 GND.n2753 GND.n2752 0.152939
R22400 GND.n2754 GND.n2753 0.152939
R22401 GND.n2755 GND.n2754 0.152939
R22402 GND.n2760 GND.n2755 0.152939
R22403 GND.n2761 GND.n2760 0.152939
R22404 GND.n2762 GND.n2761 0.152939
R22405 GND.n2763 GND.n2762 0.152939
R22406 GND.n2768 GND.n2763 0.152939
R22407 GND.n2769 GND.n2768 0.152939
R22408 GND.n2770 GND.n2769 0.152939
R22409 GND.n2771 GND.n2770 0.152939
R22410 GND.n2776 GND.n2771 0.152939
R22411 GND.n2777 GND.n2776 0.152939
R22412 GND.n2778 GND.n2777 0.152939
R22413 GND.n2779 GND.n2778 0.152939
R22414 GND.n2784 GND.n2779 0.152939
R22415 GND.n2785 GND.n2784 0.152939
R22416 GND.n2786 GND.n2785 0.152939
R22417 GND.n2787 GND.n2786 0.152939
R22418 GND.n2792 GND.n2787 0.152939
R22419 GND.n2793 GND.n2792 0.152939
R22420 GND.n2794 GND.n2793 0.152939
R22421 GND.n2795 GND.n2794 0.152939
R22422 GND.n2800 GND.n2795 0.152939
R22423 GND.n2801 GND.n2800 0.152939
R22424 GND.n2802 GND.n2801 0.152939
R22425 GND.n2803 GND.n2802 0.152939
R22426 GND.n2808 GND.n2803 0.152939
R22427 GND.n2809 GND.n2808 0.152939
R22428 GND.n2810 GND.n2809 0.152939
R22429 GND.n2811 GND.n2810 0.152939
R22430 GND.n2816 GND.n2811 0.152939
R22431 GND.n2817 GND.n2816 0.152939
R22432 GND.n2818 GND.n2817 0.152939
R22433 GND.n2819 GND.n2818 0.152939
R22434 GND.n2824 GND.n2819 0.152939
R22435 GND.n2825 GND.n2824 0.152939
R22436 GND.n2826 GND.n2825 0.152939
R22437 GND.n2827 GND.n2826 0.152939
R22438 GND.n2832 GND.n2827 0.152939
R22439 GND.n2833 GND.n2832 0.152939
R22440 GND.n2834 GND.n2833 0.152939
R22441 GND.n2835 GND.n2834 0.152939
R22442 GND.n2840 GND.n2835 0.152939
R22443 GND.n2841 GND.n2840 0.152939
R22444 GND.n2842 GND.n2841 0.152939
R22445 GND.n2843 GND.n2842 0.152939
R22446 GND.n2848 GND.n2843 0.152939
R22447 GND.n2849 GND.n2848 0.152939
R22448 GND.n2850 GND.n2849 0.152939
R22449 GND.n2851 GND.n2850 0.152939
R22450 GND.n2856 GND.n2851 0.152939
R22451 GND.n2857 GND.n2856 0.152939
R22452 GND.n2858 GND.n2857 0.152939
R22453 GND.n2859 GND.n2858 0.152939
R22454 GND.n2864 GND.n2859 0.152939
R22455 GND.n2865 GND.n2864 0.152939
R22456 GND.n2866 GND.n2865 0.152939
R22457 GND.n2867 GND.n2866 0.152939
R22458 GND.n2872 GND.n2867 0.152939
R22459 GND.n2873 GND.n2872 0.152939
R22460 GND.n2874 GND.n2873 0.152939
R22461 GND.n2875 GND.n2874 0.152939
R22462 GND.n2880 GND.n2875 0.152939
R22463 GND.n2881 GND.n2880 0.152939
R22464 GND.n2882 GND.n2881 0.152939
R22465 GND.n2883 GND.n2882 0.152939
R22466 GND.n2888 GND.n2883 0.152939
R22467 GND.n2889 GND.n2888 0.152939
R22468 GND.n2890 GND.n2889 0.152939
R22469 GND.n2891 GND.n2890 0.152939
R22470 GND.n2896 GND.n2891 0.152939
R22471 GND.n2897 GND.n2896 0.152939
R22472 GND.n2898 GND.n2897 0.152939
R22473 GND.n2899 GND.n2898 0.152939
R22474 GND.n2904 GND.n2899 0.152939
R22475 GND.n2905 GND.n2904 0.152939
R22476 GND.n2906 GND.n2905 0.152939
R22477 GND.n2907 GND.n2906 0.152939
R22478 GND.n2912 GND.n2907 0.152939
R22479 GND.n2913 GND.n2912 0.152939
R22480 GND.n2914 GND.n2913 0.152939
R22481 GND.n2915 GND.n2914 0.152939
R22482 GND.n2920 GND.n2915 0.152939
R22483 GND.n2921 GND.n2920 0.152939
R22484 GND.n2922 GND.n2921 0.152939
R22485 GND.n2923 GND.n2922 0.152939
R22486 GND.n2928 GND.n2923 0.152939
R22487 GND.n2929 GND.n2928 0.152939
R22488 GND.n2930 GND.n2929 0.152939
R22489 GND.n2931 GND.n2930 0.152939
R22490 GND.n2936 GND.n2931 0.152939
R22491 GND.n2937 GND.n2936 0.152939
R22492 GND.n2938 GND.n2937 0.152939
R22493 GND.n2939 GND.n2938 0.152939
R22494 GND.n2944 GND.n2939 0.152939
R22495 GND.n2945 GND.n2944 0.152939
R22496 GND.n2946 GND.n2945 0.152939
R22497 GND.n2947 GND.n2946 0.152939
R22498 GND.n2952 GND.n2947 0.152939
R22499 GND.n2953 GND.n2952 0.152939
R22500 GND.n2954 GND.n2953 0.152939
R22501 GND.n2955 GND.n2954 0.152939
R22502 GND.n2960 GND.n2955 0.152939
R22503 GND.n2961 GND.n2960 0.152939
R22504 GND.n2962 GND.n2961 0.152939
R22505 GND.n2963 GND.n2962 0.152939
R22506 GND.n2968 GND.n2963 0.152939
R22507 GND.n3210 GND.n2969 0.152939
R22508 GND.n3210 GND.n3209 0.152939
R22509 GND.n3209 GND.n3208 0.152939
R22510 GND.n3208 GND.n2971 0.152939
R22511 GND.n2978 GND.n2971 0.152939
R22512 GND.n2979 GND.n2978 0.152939
R22513 GND.n2980 GND.n2979 0.152939
R22514 GND.n2985 GND.n2980 0.152939
R22515 GND.n2986 GND.n2985 0.152939
R22516 GND.n2987 GND.n2986 0.152939
R22517 GND.n2988 GND.n2987 0.152939
R22518 GND.n2993 GND.n2988 0.152939
R22519 GND.n2994 GND.n2993 0.152939
R22520 GND.n2995 GND.n2994 0.152939
R22521 GND.n2996 GND.n2995 0.152939
R22522 GND.n3001 GND.n2996 0.152939
R22523 GND.n3002 GND.n3001 0.152939
R22524 GND.n3003 GND.n3002 0.152939
R22525 GND.n3004 GND.n3003 0.152939
R22526 GND.n3009 GND.n3004 0.152939
R22527 GND.n3010 GND.n3009 0.152939
R22528 GND.n3011 GND.n3010 0.152939
R22529 GND.n3012 GND.n3011 0.152939
R22530 GND.n3017 GND.n3012 0.152939
R22531 GND.n3018 GND.n3017 0.152939
R22532 GND.n3019 GND.n3018 0.152939
R22533 GND.n3020 GND.n3019 0.152939
R22534 GND.n3025 GND.n3020 0.152939
R22535 GND.n3026 GND.n3025 0.152939
R22536 GND.n3027 GND.n3026 0.152939
R22537 GND.n3028 GND.n3027 0.152939
R22538 GND.n3033 GND.n3028 0.152939
R22539 GND.n3034 GND.n3033 0.152939
R22540 GND.n3035 GND.n3034 0.152939
R22541 GND.n3036 GND.n3035 0.152939
R22542 GND.n3041 GND.n3036 0.152939
R22543 GND.n3042 GND.n3041 0.152939
R22544 GND.n3043 GND.n3042 0.152939
R22545 GND.n3044 GND.n3043 0.152939
R22546 GND.n3049 GND.n3044 0.152939
R22547 GND.n3050 GND.n3049 0.152939
R22548 GND.n3051 GND.n3050 0.152939
R22549 GND.n3052 GND.n3051 0.152939
R22550 GND.n3057 GND.n3052 0.152939
R22551 GND.n3058 GND.n3057 0.152939
R22552 GND.n3059 GND.n3058 0.152939
R22553 GND.n3060 GND.n3059 0.152939
R22554 GND.n3065 GND.n3060 0.152939
R22555 GND.n3066 GND.n3065 0.152939
R22556 GND.n3067 GND.n3066 0.152939
R22557 GND.n3068 GND.n3067 0.152939
R22558 GND.n3073 GND.n3068 0.152939
R22559 GND.n3074 GND.n3073 0.152939
R22560 GND.n3075 GND.n3074 0.152939
R22561 GND.n3076 GND.n3075 0.152939
R22562 GND.n3081 GND.n3076 0.152939
R22563 GND.n3082 GND.n3081 0.152939
R22564 GND.n3083 GND.n3082 0.152939
R22565 GND.n3084 GND.n3083 0.152939
R22566 GND.n3087 GND.n3084 0.152939
R22567 GND.n3088 GND.n3087 0.152939
R22568 GND.n3088 GND.n385 0.152939
R22569 GND.n8262 GND.n385 0.152939
R22570 GND.n8042 GND.n8041 0.152939
R22571 GND.n8043 GND.n8042 0.152939
R22572 GND.n8044 GND.n8043 0.152939
R22573 GND.n8047 GND.n8044 0.152939
R22574 GND.n8048 GND.n8047 0.152939
R22575 GND.n8049 GND.n8048 0.152939
R22576 GND.n8050 GND.n8049 0.152939
R22577 GND.n8053 GND.n8050 0.152939
R22578 GND.n8054 GND.n8053 0.152939
R22579 GND.n8055 GND.n8054 0.152939
R22580 GND.n8056 GND.n8055 0.152939
R22581 GND.n8059 GND.n8056 0.152939
R22582 GND.n8060 GND.n8059 0.152939
R22583 GND.n8061 GND.n8060 0.152939
R22584 GND.n8062 GND.n8061 0.152939
R22585 GND.n8065 GND.n8062 0.152939
R22586 GND.n8066 GND.n8065 0.152939
R22587 GND.n8067 GND.n8066 0.152939
R22588 GND.n8068 GND.n8067 0.152939
R22589 GND.n8071 GND.n8068 0.152939
R22590 GND.n8072 GND.n8071 0.152939
R22591 GND.n8073 GND.n8072 0.152939
R22592 GND.n8074 GND.n8073 0.152939
R22593 GND.n8075 GND.n8074 0.152939
R22594 GND.n8076 GND.n8075 0.152939
R22595 GND.n8076 GND.n390 0.152939
R22596 GND.n8251 GND.n390 0.152939
R22597 GND.n8252 GND.n8251 0.152939
R22598 GND.n8254 GND.n8252 0.152939
R22599 GND.n8254 GND.n8253 0.152939
R22600 GND.n8253 GND.n386 0.152939
R22601 GND.n8261 GND.n386 0.152939
R22602 GND.n194 GND.n166 0.152939
R22603 GND.n195 GND.n194 0.152939
R22604 GND.n196 GND.n195 0.152939
R22605 GND.n214 GND.n196 0.152939
R22606 GND.n215 GND.n214 0.152939
R22607 GND.n216 GND.n215 0.152939
R22608 GND.n217 GND.n216 0.152939
R22609 GND.n235 GND.n217 0.152939
R22610 GND.n236 GND.n235 0.152939
R22611 GND.n237 GND.n236 0.152939
R22612 GND.n238 GND.n237 0.152939
R22613 GND.n255 GND.n238 0.152939
R22614 GND.n256 GND.n255 0.152939
R22615 GND.n257 GND.n256 0.152939
R22616 GND.n258 GND.n257 0.152939
R22617 GND.n276 GND.n258 0.152939
R22618 GND.n277 GND.n276 0.152939
R22619 GND.n278 GND.n277 0.152939
R22620 GND.n279 GND.n278 0.152939
R22621 GND.n297 GND.n279 0.152939
R22622 GND.n298 GND.n297 0.152939
R22623 GND.n299 GND.n298 0.152939
R22624 GND.n300 GND.n299 0.152939
R22625 GND.n317 GND.n300 0.152939
R22626 GND.n318 GND.n317 0.152939
R22627 GND.n319 GND.n318 0.152939
R22628 GND.n320 GND.n319 0.152939
R22629 GND.n338 GND.n320 0.152939
R22630 GND.n339 GND.n338 0.152939
R22631 GND.n340 GND.n339 0.152939
R22632 GND.n341 GND.n340 0.152939
R22633 GND.n6917 GND.n1077 0.152939
R22634 GND.n6925 GND.n1077 0.152939
R22635 GND.n6926 GND.n6925 0.152939
R22636 GND.n6928 GND.n6926 0.152939
R22637 GND.n6928 GND.n6927 0.152939
R22638 GND.n5595 GND.n5594 0.152939
R22639 GND.n5595 GND.n5591 0.152939
R22640 GND.n5601 GND.n5591 0.152939
R22641 GND.n5602 GND.n5601 0.152939
R22642 GND.n5603 GND.n5602 0.152939
R22643 GND.n5604 GND.n5603 0.152939
R22644 GND.n5605 GND.n5604 0.152939
R22645 GND.n5606 GND.n5605 0.152939
R22646 GND.n5607 GND.n5606 0.152939
R22647 GND.n5608 GND.n5607 0.152939
R22648 GND.n5610 GND.n5608 0.152939
R22649 GND.n5610 GND.n5609 0.152939
R22650 GND.n5609 GND.n1514 0.152939
R22651 GND.n1515 GND.n1514 0.152939
R22652 GND.n1516 GND.n1515 0.152939
R22653 GND.n6211 GND.n1516 0.152939
R22654 GND.n6214 GND.n6211 0.152939
R22655 GND.n6215 GND.n6214 0.152939
R22656 GND.n6216 GND.n6215 0.152939
R22657 GND.n6216 GND.n6209 0.152939
R22658 GND.n6222 GND.n6209 0.152939
R22659 GND.n6223 GND.n6222 0.152939
R22660 GND.n6224 GND.n6223 0.152939
R22661 GND.n6224 GND.n6207 0.152939
R22662 GND.n6230 GND.n6207 0.152939
R22663 GND.n6231 GND.n6230 0.152939
R22664 GND.n6232 GND.n6231 0.152939
R22665 GND.n6233 GND.n6232 0.152939
R22666 GND.n6233 GND.n1419 0.152939
R22667 GND.n6407 GND.n1419 0.152939
R22668 GND.n6408 GND.n6407 0.152939
R22669 GND.n6409 GND.n6408 0.152939
R22670 GND.n6409 GND.n1417 0.152939
R22671 GND.n6415 GND.n1417 0.152939
R22672 GND.n6416 GND.n6415 0.152939
R22673 GND.n6417 GND.n6416 0.152939
R22674 GND.n6417 GND.n1415 0.152939
R22675 GND.n6423 GND.n1415 0.152939
R22676 GND.n6424 GND.n6423 0.152939
R22677 GND.n6425 GND.n6424 0.152939
R22678 GND.n6425 GND.n1413 0.152939
R22679 GND.n6431 GND.n1413 0.152939
R22680 GND.n6432 GND.n6431 0.152939
R22681 GND.n6433 GND.n6432 0.152939
R22682 GND.n6433 GND.n1411 0.152939
R22683 GND.n6439 GND.n1411 0.152939
R22684 GND.n6440 GND.n6439 0.152939
R22685 GND.n6441 GND.n6440 0.152939
R22686 GND.n6441 GND.n1409 0.152939
R22687 GND.n6448 GND.n1409 0.152939
R22688 GND.n6449 GND.n6448 0.152939
R22689 GND.n6450 GND.n6449 0.152939
R22690 GND.n6451 GND.n6450 0.152939
R22691 GND.n6452 GND.n6451 0.152939
R22692 GND.n6453 GND.n6452 0.152939
R22693 GND.n6454 GND.n6453 0.152939
R22694 GND.n6455 GND.n6454 0.152939
R22695 GND.n6456 GND.n6455 0.152939
R22696 GND.n6457 GND.n6456 0.152939
R22697 GND.n6459 GND.n6457 0.152939
R22698 GND.n6459 GND.n6458 0.152939
R22699 GND.n6458 GND.n1179 0.152939
R22700 GND.n1180 GND.n1179 0.152939
R22701 GND.n1181 GND.n1180 0.152939
R22702 GND.n1191 GND.n1181 0.152939
R22703 GND.n1192 GND.n1191 0.152939
R22704 GND.n1193 GND.n1192 0.152939
R22705 GND.n1194 GND.n1193 0.152939
R22706 GND.n6722 GND.n1194 0.152939
R22707 GND.n6723 GND.n6722 0.152939
R22708 GND.n6723 GND.n6721 0.152939
R22709 GND.n6729 GND.n6721 0.152939
R22710 GND.n6730 GND.n6729 0.152939
R22711 GND.n6731 GND.n6730 0.152939
R22712 GND.n6732 GND.n6731 0.152939
R22713 GND.n6734 GND.n6732 0.152939
R22714 GND.n6734 GND.n6733 0.152939
R22715 GND.n6733 GND.n1084 0.152939
R22716 GND.n6909 GND.n1084 0.152939
R22717 GND.n6910 GND.n6909 0.152939
R22718 GND.n6911 GND.n6910 0.152939
R22719 GND.n6911 GND.n1080 0.152939
R22720 GND.n6916 GND.n1080 0.152939
R22721 GND.n1589 GND.n1588 0.152939
R22722 GND.n1590 GND.n1589 0.152939
R22723 GND.n1591 GND.n1590 0.152939
R22724 GND.n1592 GND.n1591 0.152939
R22725 GND.n1593 GND.n1592 0.152939
R22726 GND.n6068 GND.n6065 0.152939
R22727 GND.n6068 GND.n1565 0.152939
R22728 GND.n6113 GND.n6112 0.152939
R22729 GND.n6114 GND.n6113 0.152939
R22730 GND.n6114 GND.n1550 0.152939
R22731 GND.n6128 GND.n1550 0.152939
R22732 GND.n6129 GND.n6128 0.152939
R22733 GND.n6130 GND.n6129 0.152939
R22734 GND.n6131 GND.n6130 0.152939
R22735 GND.n6132 GND.n6131 0.152939
R22736 GND.n6133 GND.n6132 0.152939
R22737 GND.n6134 GND.n6133 0.152939
R22738 GND.n6134 GND.n1490 0.152939
R22739 GND.n6332 GND.n1490 0.152939
R22740 GND.n6333 GND.n6332 0.152939
R22741 GND.n6334 GND.n6333 0.152939
R22742 GND.n6334 GND.n1474 0.152939
R22743 GND.n6348 GND.n1474 0.152939
R22744 GND.n6349 GND.n6348 0.152939
R22745 GND.n6350 GND.n6349 0.152939
R22746 GND.n6350 GND.n1458 0.152939
R22747 GND.n6364 GND.n1458 0.152939
R22748 GND.n6365 GND.n6364 0.152939
R22749 GND.n6366 GND.n6365 0.152939
R22750 GND.n6366 GND.n1442 0.152939
R22751 GND.n6379 GND.n1442 0.152939
R22752 GND.n6380 GND.n6379 0.152939
R22753 GND.n6381 GND.n6380 0.152939
R22754 GND.n6381 GND.n1425 0.152939
R22755 GND.n6397 GND.n1425 0.152939
R22756 GND.n6398 GND.n6397 0.152939
R22757 GND.n6399 GND.n6398 0.152939
R22758 GND.n6400 GND.n6399 0.152939
R22759 GND.n6400 GND.n1309 0.152939
R22760 GND.n6571 GND.n1309 0.152939
R22761 GND.n6572 GND.n6571 0.152939
R22762 GND.n6573 GND.n6572 0.152939
R22763 GND.n6573 GND.n1293 0.152939
R22764 GND.n6587 GND.n1293 0.152939
R22765 GND.n6588 GND.n6587 0.152939
R22766 GND.n6589 GND.n6588 0.152939
R22767 GND.n6589 GND.n1277 0.152939
R22768 GND.n6603 GND.n1277 0.152939
R22769 GND.n6604 GND.n6603 0.152939
R22770 GND.n6605 GND.n6604 0.152939
R22771 GND.n6605 GND.n1261 0.152939
R22772 GND.n6618 GND.n1261 0.152939
R22773 GND.n6619 GND.n6618 0.152939
R22774 GND.n6620 GND.n6619 0.152939
R22775 GND.n6620 GND.n1245 0.152939
R22776 GND.n6634 GND.n1245 0.152939
R22777 GND.n6635 GND.n6634 0.152939
R22778 GND.n6636 GND.n6635 0.152939
R22779 GND.n6636 GND.n1229 0.152939
R22780 GND.n6650 GND.n1229 0.152939
R22781 GND.n6651 GND.n6650 0.152939
R22782 GND.n6652 GND.n6651 0.152939
R22783 GND.n6653 GND.n6652 0.152939
R22784 GND.n6654 GND.n6653 0.152939
R22785 GND.n6655 GND.n6654 0.152939
R22786 GND.n6656 GND.n6655 0.152939
R22787 GND.n6656 GND.n1155 0.152939
R22788 GND.n6829 GND.n1155 0.152939
R22789 GND.n6830 GND.n6829 0.152939
R22790 GND.n6831 GND.n6830 0.152939
R22791 GND.n6831 GND.n1139 0.152939
R22792 GND.n6845 GND.n1139 0.152939
R22793 GND.n6846 GND.n6845 0.152939
R22794 GND.n6847 GND.n6846 0.152939
R22795 GND.n6847 GND.n1123 0.152939
R22796 GND.n6861 GND.n1123 0.152939
R22797 GND.n6862 GND.n6861 0.152939
R22798 GND.n6863 GND.n6862 0.152939
R22799 GND.n6863 GND.n1107 0.152939
R22800 GND.n6876 GND.n1107 0.152939
R22801 GND.n6877 GND.n6876 0.152939
R22802 GND.n6878 GND.n6877 0.152939
R22803 GND.n6879 GND.n6878 0.152939
R22804 GND.n6881 GND.n6879 0.152939
R22805 GND.n6881 GND.n6880 0.152939
R22806 GND.n6880 GND.n1061 0.152939
R22807 GND.n1062 GND.n1061 0.152939
R22808 GND.n1063 GND.n1062 0.152939
R22809 GND.n1064 GND.n1063 0.152939
R22810 GND.n6968 GND.n1064 0.152939
R22811 GND.n6967 GND.n6966 0.152939
R22812 GND.n6969 GND.n6967 0.152939
R22813 GND.n7733 GND.n7732 0.152939
R22814 GND.n7733 GND.n634 0.152939
R22815 GND.n7767 GND.n634 0.152939
R22816 GND.n7768 GND.n7767 0.152939
R22817 GND.n7769 GND.n7768 0.152939
R22818 GND.n7770 GND.n7769 0.152939
R22819 GND.n7770 GND.n606 0.152939
R22820 GND.n7804 GND.n606 0.152939
R22821 GND.n7805 GND.n7804 0.152939
R22822 GND.n7806 GND.n7805 0.152939
R22823 GND.n7807 GND.n7806 0.152939
R22824 GND.n7808 GND.n7807 0.152939
R22825 GND.n7808 GND.n579 0.152939
R22826 GND.n7840 GND.n579 0.152939
R22827 GND.n7841 GND.n7840 0.152939
R22828 GND.n7843 GND.n7841 0.152939
R22829 GND.n7843 GND.n7842 0.152939
R22830 GND.n7842 GND.n556 0.152939
R22831 GND.n556 GND.n554 0.152939
R22832 GND.n7875 GND.n554 0.152939
R22833 GND.n7876 GND.n7875 0.152939
R22834 GND.n7877 GND.n7876 0.152939
R22835 GND.n7878 GND.n7877 0.152939
R22836 GND.n7878 GND.n492 0.152939
R22837 GND.n7957 GND.n492 0.152939
R22838 GND.n7958 GND.n7957 0.152939
R22839 GND.n7959 GND.n7958 0.152939
R22840 GND.n7960 GND.n7959 0.152939
R22841 GND.n7960 GND.n465 0.152939
R22842 GND.n7994 GND.n465 0.152939
R22843 GND.n7995 GND.n7994 0.152939
R22844 GND.n7996 GND.n7995 0.152939
R22845 GND.n7997 GND.n7996 0.152939
R22846 GND.n7998 GND.n7997 0.152939
R22847 GND.n7999 GND.n7998 0.152939
R22848 GND.n7999 GND.n152 0.152939
R22849 GND.n8569 GND.n153 0.152939
R22850 GND.n426 GND.n153 0.152939
R22851 GND.n8135 GND.n426 0.152939
R22852 GND.n8136 GND.n8135 0.152939
R22853 GND.n8137 GND.n8136 0.152939
R22854 GND.n8137 GND.n422 0.152939
R22855 GND.n8150 GND.n422 0.152939
R22856 GND.n8151 GND.n8150 0.152939
R22857 GND.n8152 GND.n8151 0.152939
R22858 GND.n8152 GND.n418 0.152939
R22859 GND.n8165 GND.n418 0.152939
R22860 GND.n8166 GND.n8165 0.152939
R22861 GND.n8167 GND.n8166 0.152939
R22862 GND.n8167 GND.n414 0.152939
R22863 GND.n8180 GND.n414 0.152939
R22864 GND.n8181 GND.n8180 0.152939
R22865 GND.n8182 GND.n8181 0.152939
R22866 GND.n8182 GND.n409 0.152939
R22867 GND.n8195 GND.n409 0.152939
R22868 GND.n8196 GND.n8195 0.152939
R22869 GND.n8197 GND.n8196 0.152939
R22870 GND.n8197 GND.n405 0.152939
R22871 GND.n8210 GND.n405 0.152939
R22872 GND.n8211 GND.n8210 0.152939
R22873 GND.n8212 GND.n8211 0.152939
R22874 GND.n8212 GND.n401 0.152939
R22875 GND.n8225 GND.n401 0.152939
R22876 GND.n8226 GND.n8225 0.152939
R22877 GND.n8228 GND.n8226 0.152939
R22878 GND.n8228 GND.n8227 0.152939
R22879 GND.n8227 GND.n395 0.152939
R22880 GND.n396 GND.n395 0.152939
R22881 GND.n398 GND.n396 0.152939
R22882 GND.n398 GND.n397 0.152939
R22883 GND.n397 GND.n352 0.152939
R22884 GND.n8452 GND.n352 0.152939
R22885 GND.n367 GND.n366 0.152939
R22886 GND.n368 GND.n367 0.152939
R22887 GND.n368 GND.n362 0.152939
R22888 GND.n375 GND.n362 0.152939
R22889 GND.n376 GND.n375 0.152939
R22890 GND.n377 GND.n376 0.152939
R22891 GND.n377 GND.n353 0.152939
R22892 GND.n8451 GND.n353 0.152939
R22893 GND.n8294 GND.n8293 0.152939
R22894 GND.n8295 GND.n8294 0.152939
R22895 GND.n8296 GND.n8295 0.152939
R22896 GND.n8297 GND.n8296 0.152939
R22897 GND.n8298 GND.n8297 0.152939
R22898 GND.n8299 GND.n8298 0.152939
R22899 GND.n8300 GND.n8299 0.152939
R22900 GND.n8433 GND.n8300 0.152939
R22901 GND.n8433 GND.n8432 0.152939
R22902 GND.n8432 GND.n8431 0.152939
R22903 GND.n8431 GND.n8306 0.152939
R22904 GND.n8307 GND.n8306 0.152939
R22905 GND.n8308 GND.n8307 0.152939
R22906 GND.n8309 GND.n8308 0.152939
R22907 GND.n8310 GND.n8309 0.152939
R22908 GND.n8311 GND.n8310 0.152939
R22909 GND.n8312 GND.n8311 0.152939
R22910 GND.n8313 GND.n8312 0.152939
R22911 GND.n8314 GND.n8313 0.152939
R22912 GND.n8315 GND.n8314 0.152939
R22913 GND.n8316 GND.n8315 0.152939
R22914 GND.n8317 GND.n8316 0.152939
R22915 GND.n8318 GND.n8317 0.152939
R22916 GND.n8319 GND.n8318 0.152939
R22917 GND.n8320 GND.n8319 0.152939
R22918 GND.n8321 GND.n8320 0.152939
R22919 GND.n8391 GND.n8321 0.152939
R22920 GND.n8391 GND.n8390 0.152939
R22921 GND.n8390 GND.n8389 0.152939
R22922 GND.n8389 GND.n8325 0.152939
R22923 GND.n8326 GND.n8325 0.152939
R22924 GND.n8327 GND.n8326 0.152939
R22925 GND.n8328 GND.n8327 0.152939
R22926 GND.n8329 GND.n8328 0.152939
R22927 GND.n8330 GND.n8329 0.152939
R22928 GND.n8331 GND.n8330 0.152939
R22929 GND.n8369 GND.n8331 0.152939
R22930 GND.n8369 GND.n8368 0.152939
R22931 GND.n8368 GND.n8367 0.152939
R22932 GND.n8367 GND.n8335 0.152939
R22933 GND.n8336 GND.n8335 0.152939
R22934 GND.n8337 GND.n8336 0.152939
R22935 GND.n8338 GND.n8337 0.152939
R22936 GND.n8339 GND.n8338 0.152939
R22937 GND.n8340 GND.n8339 0.152939
R22938 GND.n8341 GND.n8340 0.152939
R22939 GND.n8347 GND.n8341 0.152939
R22940 GND.n8347 GND.n8346 0.152939
R22941 GND.n710 GND.n709 0.152939
R22942 GND.n711 GND.n710 0.152939
R22943 GND.n712 GND.n711 0.152939
R22944 GND.n713 GND.n712 0.152939
R22945 GND.n714 GND.n713 0.152939
R22946 GND.n715 GND.n714 0.152939
R22947 GND.n716 GND.n715 0.152939
R22948 GND.n718 GND.n716 0.152939
R22949 GND.n721 GND.n718 0.152939
R22950 GND.n722 GND.n721 0.152939
R22951 GND.n723 GND.n722 0.152939
R22952 GND.n724 GND.n723 0.152939
R22953 GND.n725 GND.n724 0.152939
R22954 GND.n726 GND.n725 0.152939
R22955 GND.n727 GND.n726 0.152939
R22956 GND.n728 GND.n727 0.152939
R22957 GND.n729 GND.n728 0.152939
R22958 GND.n732 GND.n729 0.152939
R22959 GND.n733 GND.n732 0.152939
R22960 GND.n734 GND.n733 0.152939
R22961 GND.n7600 GND.n7599 0.152939
R22962 GND.n7601 GND.n7600 0.152939
R22963 GND.n7602 GND.n7601 0.152939
R22964 GND.n7603 GND.n7602 0.152939
R22965 GND.n7606 GND.n7603 0.152939
R22966 GND.n7607 GND.n7606 0.152939
R22967 GND.n7608 GND.n7607 0.152939
R22968 GND.n7609 GND.n7608 0.152939
R22969 GND.n7610 GND.n7609 0.152939
R22970 GND.n7611 GND.n7610 0.152939
R22971 GND.n7612 GND.n7611 0.152939
R22972 GND.n7613 GND.n7612 0.152939
R22973 GND.n7614 GND.n7613 0.152939
R22974 GND.n7615 GND.n7614 0.152939
R22975 GND.n7618 GND.n7615 0.152939
R22976 GND.n7619 GND.n7618 0.152939
R22977 GND.n7620 GND.n7619 0.152939
R22978 GND.n7621 GND.n7620 0.152939
R22979 GND.n7622 GND.n7621 0.152939
R22980 GND.n7623 GND.n7622 0.152939
R22981 GND.n7624 GND.n7623 0.152939
R22982 GND.n7625 GND.n7624 0.152939
R22983 GND.n7626 GND.n7625 0.152939
R22984 GND.n7631 GND.n7626 0.152939
R22985 GND.n7631 GND.n7630 0.152939
R22986 GND.n7757 GND.n644 0.152939
R22987 GND.n7758 GND.n7757 0.152939
R22988 GND.n7759 GND.n7758 0.152939
R22989 GND.n7760 GND.n7759 0.152939
R22990 GND.n7760 GND.n616 0.152939
R22991 GND.n7794 GND.n616 0.152939
R22992 GND.n7795 GND.n7794 0.152939
R22993 GND.n7796 GND.n7795 0.152939
R22994 GND.n7797 GND.n7796 0.152939
R22995 GND.n7797 GND.n589 0.152939
R22996 GND.n7829 GND.n589 0.152939
R22997 GND.n7830 GND.n7829 0.152939
R22998 GND.n7831 GND.n7830 0.152939
R22999 GND.n7831 GND.n567 0.152939
R23000 GND.n7856 GND.n567 0.152939
R23001 GND.n7857 GND.n7856 0.152939
R23002 GND.n7858 GND.n7857 0.152939
R23003 GND.n7858 GND.n533 0.152939
R23004 GND.n7894 GND.n533 0.152939
R23005 GND.n7895 GND.n7894 0.152939
R23006 GND.n7896 GND.n7895 0.152939
R23007 GND.n7896 GND.n502 0.152939
R23008 GND.n7947 GND.n502 0.152939
R23009 GND.n7948 GND.n7947 0.152939
R23010 GND.n7949 GND.n7948 0.152939
R23011 GND.n7950 GND.n7949 0.152939
R23012 GND.n7950 GND.n475 0.152939
R23013 GND.n7984 GND.n475 0.152939
R23014 GND.n7985 GND.n7984 0.152939
R23015 GND.n7986 GND.n7985 0.152939
R23016 GND.n7986 GND.n167 0.152939
R23017 GND.n1872 GND.n1853 0.152939
R23018 GND.n4710 GND.n1853 0.152939
R23019 GND.n4711 GND.n4710 0.152939
R23020 GND.n4712 GND.n4711 0.152939
R23021 GND.n4713 GND.n4712 0.152939
R23022 GND.n4714 GND.n4713 0.152939
R23023 GND.n4716 GND.n4714 0.152939
R23024 GND.n4717 GND.n4716 0.152939
R23025 GND.n4718 GND.n4717 0.152939
R23026 GND.n4718 GND.n1789 0.152939
R23027 GND.n4803 GND.n1789 0.152939
R23028 GND.n4804 GND.n4803 0.152939
R23029 GND.n4805 GND.n4804 0.152939
R23030 GND.n4806 GND.n4805 0.152939
R23031 GND.n4807 GND.n4806 0.152939
R23032 GND.n4810 GND.n4807 0.152939
R23033 GND.n4811 GND.n4810 0.152939
R23034 GND.n4812 GND.n4811 0.152939
R23035 GND.n4813 GND.n4812 0.152939
R23036 GND.n4815 GND.n4813 0.152939
R23037 GND.n4816 GND.n4815 0.152939
R23038 GND.n4816 GND.n1707 0.152939
R23039 GND.n4933 GND.n1707 0.152939
R23040 GND.n4934 GND.n4933 0.152939
R23041 GND.n4935 GND.n4934 0.152939
R23042 GND.n4936 GND.n4935 0.152939
R23043 GND.n4937 GND.n4936 0.152939
R23044 GND.n4940 GND.n4937 0.152939
R23045 GND.n4941 GND.n4940 0.152939
R23046 GND.n4942 GND.n4941 0.152939
R23047 GND.n4943 GND.n4942 0.152939
R23048 GND.n4946 GND.n4943 0.152939
R23049 GND.n4947 GND.n4946 0.152939
R23050 GND.n4948 GND.n4947 0.152939
R23051 GND.n4949 GND.n4948 0.152939
R23052 GND.n4955 GND.n4949 0.152939
R23053 GND.n4956 GND.n4955 0.152939
R23054 GND.n4957 GND.n4956 0.152939
R23055 GND.n4958 GND.n4957 0.152939
R23056 GND.n4973 GND.n4958 0.152939
R23057 GND.n4974 GND.n4973 0.152939
R23058 GND.n4975 GND.n4974 0.152939
R23059 GND.n4976 GND.n4975 0.152939
R23060 GND.n4991 GND.n4976 0.152939
R23061 GND.n4992 GND.n4991 0.152939
R23062 GND.n4993 GND.n4992 0.152939
R23063 GND.n4994 GND.n4993 0.152939
R23064 GND.n5008 GND.n4994 0.152939
R23065 GND.n5009 GND.n5008 0.152939
R23066 GND.n5010 GND.n5009 0.152939
R23067 GND.n5011 GND.n5010 0.152939
R23068 GND.n5026 GND.n5011 0.152939
R23069 GND.n5027 GND.n5026 0.152939
R23070 GND.n5028 GND.n5027 0.152939
R23071 GND.n5029 GND.n5028 0.152939
R23072 GND.n5044 GND.n5029 0.152939
R23073 GND.n5045 GND.n5044 0.152939
R23074 GND.n5046 GND.n5045 0.152939
R23075 GND.n5047 GND.n5046 0.152939
R23076 GND.n5065 GND.n5047 0.152939
R23077 GND.n5066 GND.n5065 0.152939
R23078 GND.n5067 GND.n5066 0.152939
R23079 GND.n5068 GND.n5067 0.152939
R23080 GND.n5069 GND.n5068 0.152939
R23081 GND.n5083 GND.n5069 0.152939
R23082 GND.n5084 GND.n5083 0.152939
R23083 GND.n5085 GND.n5084 0.152939
R23084 GND.n5086 GND.n5085 0.152939
R23085 GND.n5101 GND.n5086 0.152939
R23086 GND.n5102 GND.n5101 0.152939
R23087 GND.n5103 GND.n5102 0.152939
R23088 GND.n5104 GND.n5103 0.152939
R23089 GND.n5119 GND.n5104 0.152939
R23090 GND.n5120 GND.n5119 0.152939
R23091 GND.n5121 GND.n5120 0.152939
R23092 GND.n5122 GND.n5121 0.152939
R23093 GND.n5140 GND.n5122 0.152939
R23094 GND.n5141 GND.n5140 0.152939
R23095 GND.n5142 GND.n5141 0.152939
R23096 GND.n5143 GND.n5142 0.152939
R23097 GND.n5144 GND.n5143 0.152939
R23098 GND.n5159 GND.n5144 0.152939
R23099 GND.n5160 GND.n5159 0.152939
R23100 GND.n5161 GND.n5160 0.152939
R23101 GND.n5162 GND.n5161 0.152939
R23102 GND.n5177 GND.n5162 0.152939
R23103 GND.n5178 GND.n5177 0.152939
R23104 GND.n5179 GND.n5178 0.152939
R23105 GND.n5180 GND.n5179 0.152939
R23106 GND.n5652 GND.n5180 0.152939
R23107 GND.n5653 GND.n5652 0.152939
R23108 GND.n5653 GND.n1572 0.152939
R23109 GND.n6104 GND.n1572 0.152939
R23110 GND.n6105 GND.n6104 0.152939
R23111 GND.n6106 GND.n6105 0.152939
R23112 GND.n6106 GND.n1558 0.152939
R23113 GND.n6120 GND.n1558 0.152939
R23114 GND.n6121 GND.n6120 0.152939
R23115 GND.n6122 GND.n6121 0.152939
R23116 GND.n6122 GND.n1541 0.152939
R23117 GND.n6145 GND.n1541 0.152939
R23118 GND.n6146 GND.n6145 0.152939
R23119 GND.n6147 GND.n6146 0.152939
R23120 GND.n6147 GND.n1498 0.152939
R23121 GND.n6324 GND.n1498 0.152939
R23122 GND.n6325 GND.n6324 0.152939
R23123 GND.n6326 GND.n6325 0.152939
R23124 GND.n6326 GND.n1482 0.152939
R23125 GND.n6340 GND.n1482 0.152939
R23126 GND.n6341 GND.n6340 0.152939
R23127 GND.n6342 GND.n6341 0.152939
R23128 GND.n6342 GND.n1466 0.152939
R23129 GND.n6356 GND.n1466 0.152939
R23130 GND.n6357 GND.n6356 0.152939
R23131 GND.n6358 GND.n6357 0.152939
R23132 GND.n6358 GND.n1450 0.152939
R23133 GND.n6372 GND.n1450 0.152939
R23134 GND.n6373 GND.n6372 0.152939
R23135 GND.n6374 GND.n6373 0.152939
R23136 GND.n6374 GND.n1434 0.152939
R23137 GND.n6387 GND.n1434 0.152939
R23138 GND.n6388 GND.n6387 0.152939
R23139 GND.n6389 GND.n6388 0.152939
R23140 GND.n6390 GND.n6389 0.152939
R23141 GND.n6390 GND.n1316 0.152939
R23142 GND.n6563 GND.n1316 0.152939
R23143 GND.n6564 GND.n6563 0.152939
R23144 GND.n6565 GND.n6564 0.152939
R23145 GND.n6565 GND.n1301 0.152939
R23146 GND.n6579 GND.n1301 0.152939
R23147 GND.n6580 GND.n6579 0.152939
R23148 GND.n6581 GND.n6580 0.152939
R23149 GND.n6581 GND.n1285 0.152939
R23150 GND.n6595 GND.n1285 0.152939
R23151 GND.n6596 GND.n6595 0.152939
R23152 GND.n6597 GND.n6596 0.152939
R23153 GND.n6597 GND.n1269 0.152939
R23154 GND.n6611 GND.n1269 0.152939
R23155 GND.n6612 GND.n6611 0.152939
R23156 GND.n6613 GND.n6612 0.152939
R23157 GND.n6613 GND.n1253 0.152939
R23158 GND.n6626 GND.n1253 0.152939
R23159 GND.n6627 GND.n6626 0.152939
R23160 GND.n6628 GND.n6627 0.152939
R23161 GND.n6628 GND.n1237 0.152939
R23162 GND.n6642 GND.n1237 0.152939
R23163 GND.n6643 GND.n6642 0.152939
R23164 GND.n6644 GND.n6643 0.152939
R23165 GND.n6644 GND.n1220 0.152939
R23166 GND.n6667 GND.n1220 0.152939
R23167 GND.n6668 GND.n6667 0.152939
R23168 GND.n6669 GND.n6668 0.152939
R23169 GND.n6669 GND.n1163 0.152939
R23170 GND.n6821 GND.n1163 0.152939
R23171 GND.n6822 GND.n6821 0.152939
R23172 GND.n6823 GND.n6822 0.152939
R23173 GND.n6823 GND.n1147 0.152939
R23174 GND.n6837 GND.n1147 0.152939
R23175 GND.n6838 GND.n6837 0.152939
R23176 GND.n6839 GND.n6838 0.152939
R23177 GND.n6839 GND.n1131 0.152939
R23178 GND.n6853 GND.n1131 0.152939
R23179 GND.n6854 GND.n6853 0.152939
R23180 GND.n6855 GND.n6854 0.152939
R23181 GND.n6855 GND.n1115 0.152939
R23182 GND.n6869 GND.n1115 0.152939
R23183 GND.n6870 GND.n6869 0.152939
R23184 GND.n6871 GND.n6870 0.152939
R23185 GND.n6871 GND.n1098 0.152939
R23186 GND.n6889 GND.n1098 0.152939
R23187 GND.n6890 GND.n6889 0.152939
R23188 GND.n6891 GND.n6890 0.152939
R23189 GND.n6891 GND.n1052 0.152939
R23190 GND.n6982 GND.n1052 0.152939
R23191 GND.n6983 GND.n6982 0.152939
R23192 GND.n6984 GND.n6983 0.152939
R23193 GND.n6985 GND.n6984 0.152939
R23194 GND.n6986 GND.n6985 0.152939
R23195 GND.n6986 GND.n1028 0.152939
R23196 GND.n7022 GND.n1028 0.152939
R23197 GND.n7023 GND.n7022 0.152939
R23198 GND.n7024 GND.n7023 0.152939
R23199 GND.n7025 GND.n7024 0.152939
R23200 GND.n7026 GND.n7025 0.152939
R23201 GND.n7028 GND.n7026 0.152939
R23202 GND.n7029 GND.n7028 0.152939
R23203 GND.n7029 GND.n994 0.152939
R23204 GND.n7080 GND.n994 0.152939
R23205 GND.n7081 GND.n7080 0.152939
R23206 GND.n7082 GND.n7081 0.152939
R23207 GND.n7083 GND.n7082 0.152939
R23208 GND.n7083 GND.n969 0.152939
R23209 GND.n7115 GND.n969 0.152939
R23210 GND.n7116 GND.n7115 0.152939
R23211 GND.n7117 GND.n7116 0.152939
R23212 GND.n7118 GND.n7117 0.152939
R23213 GND.n7119 GND.n7118 0.152939
R23214 GND.n7119 GND.n944 0.152939
R23215 GND.n7154 GND.n944 0.152939
R23216 GND.n7155 GND.n7154 0.152939
R23217 GND.n7156 GND.n7155 0.152939
R23218 GND.n7157 GND.n7156 0.152939
R23219 GND.n7158 GND.n7157 0.152939
R23220 GND.n7160 GND.n7158 0.152939
R23221 GND.n7161 GND.n7160 0.152939
R23222 GND.n7161 GND.n912 0.152939
R23223 GND.n7214 GND.n912 0.152939
R23224 GND.n7215 GND.n7214 0.152939
R23225 GND.n7216 GND.n7215 0.152939
R23226 GND.n7217 GND.n7216 0.152939
R23227 GND.n7218 GND.n7217 0.152939
R23228 GND.n7221 GND.n7218 0.152939
R23229 GND.n7222 GND.n7221 0.152939
R23230 GND.n7223 GND.n7222 0.152939
R23231 GND.n7224 GND.n7223 0.152939
R23232 GND.n7225 GND.n7224 0.152939
R23233 GND.n7225 GND.n868 0.152939
R23234 GND.n7294 GND.n868 0.152939
R23235 GND.n7295 GND.n7294 0.152939
R23236 GND.n7296 GND.n7295 0.152939
R23237 GND.n7297 GND.n7296 0.152939
R23238 GND.n7297 GND.n843 0.152939
R23239 GND.n7330 GND.n843 0.152939
R23240 GND.n7331 GND.n7330 0.152939
R23241 GND.n7332 GND.n7331 0.152939
R23242 GND.n7332 GND.n827 0.152939
R23243 GND.n7353 GND.n827 0.152939
R23244 GND.n7354 GND.n7353 0.152939
R23245 GND.n7355 GND.n7354 0.152939
R23246 GND.n7356 GND.n7355 0.152939
R23247 GND.n7356 GND.n803 0.152939
R23248 GND.n7445 GND.n803 0.152939
R23249 GND.n7446 GND.n7445 0.152939
R23250 GND.n7447 GND.n7446 0.152939
R23251 GND.n7448 GND.n7447 0.152939
R23252 GND.n7449 GND.n7448 0.152939
R23253 GND.n7454 GND.n7449 0.152939
R23254 GND.n7455 GND.n7454 0.152939
R23255 GND.n7456 GND.n7455 0.152939
R23256 GND.n7457 GND.n7456 0.152939
R23257 GND.n7460 GND.n7457 0.152939
R23258 GND.n7461 GND.n7460 0.152939
R23259 GND.n7462 GND.n7461 0.152939
R23260 GND.n7463 GND.n7462 0.152939
R23261 GND.n7466 GND.n7463 0.152939
R23262 GND.n7467 GND.n7466 0.152939
R23263 GND.n7468 GND.n7467 0.152939
R23264 GND.n7469 GND.n7468 0.152939
R23265 GND.n7472 GND.n7469 0.152939
R23266 GND.n7473 GND.n7472 0.152939
R23267 GND.n7474 GND.n7473 0.152939
R23268 GND.n7475 GND.n7474 0.152939
R23269 GND.n7478 GND.n7475 0.152939
R23270 GND.n7479 GND.n7478 0.152939
R23271 GND.n7480 GND.n7479 0.152939
R23272 GND.n7481 GND.n7480 0.152939
R23273 GND.n7484 GND.n7481 0.152939
R23274 GND.n7485 GND.n7484 0.152939
R23275 GND.n7486 GND.n7485 0.152939
R23276 GND.n7487 GND.n7486 0.152939
R23277 GND.n7488 GND.n7487 0.152939
R23278 GND.n7488 GND.n523 0.152939
R23279 GND.n7903 GND.n523 0.152939
R23280 GND.n7904 GND.n7903 0.152939
R23281 GND.n7905 GND.n7904 0.152939
R23282 GND.n7905 GND.n519 0.152939
R23283 GND.n7911 GND.n519 0.152939
R23284 GND.n7912 GND.n7911 0.152939
R23285 GND.n7913 GND.n7912 0.152939
R23286 GND.n7914 GND.n7913 0.152939
R23287 GND.n7915 GND.n7914 0.152939
R23288 GND.n7918 GND.n7915 0.152939
R23289 GND.n7919 GND.n7918 0.152939
R23290 GND.n4690 GND.n1833 0.152939
R23291 GND.n4743 GND.n1833 0.152939
R23292 GND.n4744 GND.n4743 0.152939
R23293 GND.n4745 GND.n4744 0.152939
R23294 GND.n4746 GND.n4745 0.152939
R23295 GND.n4746 GND.n1806 0.152939
R23296 GND.n4781 GND.n1806 0.152939
R23297 GND.n4782 GND.n4781 0.152939
R23298 GND.n4783 GND.n4782 0.152939
R23299 GND.n4784 GND.n4783 0.152939
R23300 GND.n4784 GND.n1772 0.152939
R23301 GND.n4849 GND.n1772 0.152939
R23302 GND.n4850 GND.n4849 0.152939
R23303 GND.n4851 GND.n4850 0.152939
R23304 GND.n4852 GND.n4851 0.152939
R23305 GND.n4852 GND.n1745 0.152939
R23306 GND.n4886 GND.n1745 0.152939
R23307 GND.n4887 GND.n4886 0.152939
R23308 GND.n4888 GND.n4887 0.152939
R23309 GND.n4889 GND.n4888 0.152939
R23310 GND.n4889 GND.n1715 0.152939
R23311 GND.n4924 GND.n1715 0.152939
R23312 GND.n4925 GND.n4924 0.152939
R23313 GND.n4926 GND.n4925 0.152939
R23314 GND.n4926 GND.n1688 0.152939
R23315 GND.n5884 GND.n1688 0.152939
R23316 GND.n5885 GND.n5884 0.152939
R23317 GND.n5887 GND.n5885 0.152939
R23318 GND.n5887 GND.n5886 0.152939
R23319 GND.n5886 GND.n1673 0.152939
R23320 GND.n5903 GND.n1673 0.152939
R23321 GND.n4159 GND.n2128 0.152939
R23322 GND.n4160 GND.n4159 0.152939
R23323 GND.n4161 GND.n4160 0.152939
R23324 GND.n4162 GND.n4161 0.152939
R23325 GND.n4163 GND.n4162 0.152939
R23326 GND.n4164 GND.n4163 0.152939
R23327 GND.n4165 GND.n4164 0.152939
R23328 GND.n4167 GND.n4165 0.152939
R23329 GND.n4170 GND.n4167 0.152939
R23330 GND.n4171 GND.n4170 0.152939
R23331 GND.n4172 GND.n4171 0.152939
R23332 GND.n4173 GND.n4172 0.152939
R23333 GND.n4174 GND.n4173 0.152939
R23334 GND.n4175 GND.n4174 0.152939
R23335 GND.n4176 GND.n4175 0.152939
R23336 GND.n4177 GND.n4176 0.152939
R23337 GND.n4178 GND.n4177 0.152939
R23338 GND.n4181 GND.n4178 0.152939
R23339 GND.n4182 GND.n4181 0.152939
R23340 GND.n4183 GND.n4182 0.152939
R23341 GND.n4184 GND.n4183 0.152939
R23342 GND.n4185 GND.n4184 0.152939
R23343 GND.n4186 GND.n4185 0.152939
R23344 GND.n4187 GND.n4186 0.152939
R23345 GND.n4188 GND.n4187 0.152939
R23346 GND.n4189 GND.n4188 0.152939
R23347 GND.n4190 GND.n4189 0.152939
R23348 GND.n4193 GND.n4190 0.152939
R23349 GND.n4194 GND.n4193 0.152939
R23350 GND.n4195 GND.n4194 0.152939
R23351 GND.n4196 GND.n4195 0.152939
R23352 GND.n4197 GND.n4196 0.152939
R23353 GND.n4198 GND.n4197 0.152939
R23354 GND.n4199 GND.n4198 0.152939
R23355 GND.n4200 GND.n4199 0.152939
R23356 GND.n4201 GND.n4200 0.152939
R23357 GND.n4202 GND.n4201 0.152939
R23358 GND.n4205 GND.n4202 0.152939
R23359 GND.n4206 GND.n4205 0.152939
R23360 GND.n4207 GND.n4206 0.152939
R23361 GND.n4208 GND.n4207 0.152939
R23362 GND.n4209 GND.n4208 0.152939
R23363 GND.n4210 GND.n4209 0.152939
R23364 GND.n4211 GND.n4210 0.152939
R23365 GND.n4212 GND.n4211 0.152939
R23366 GND.n4213 GND.n4212 0.152939
R23367 GND.n4218 GND.n4213 0.152939
R23368 GND.n4218 GND.n2137 0.152939
R23369 GND.n4349 GND.n4348 0.152939
R23370 GND.n4350 GND.n4349 0.152939
R23371 GND.n4351 GND.n4350 0.152939
R23372 GND.n4351 GND.n2099 0.152939
R23373 GND.n4384 GND.n2099 0.152939
R23374 GND.n4385 GND.n4384 0.152939
R23375 GND.n4386 GND.n4385 0.152939
R23376 GND.n4387 GND.n4386 0.152939
R23377 GND.n4387 GND.n2070 0.152939
R23378 GND.n4427 GND.n2070 0.152939
R23379 GND.n4428 GND.n4427 0.152939
R23380 GND.n4429 GND.n4428 0.152939
R23381 GND.n4429 GND.n2036 0.152939
R23382 GND.n4466 GND.n2036 0.152939
R23383 GND.n4467 GND.n4466 0.152939
R23384 GND.n4468 GND.n4467 0.152939
R23385 GND.n4469 GND.n4468 0.152939
R23386 GND.n4469 GND.n2008 0.152939
R23387 GND.n4509 GND.n2008 0.152939
R23388 GND.n4510 GND.n4509 0.152939
R23389 GND.n4511 GND.n4510 0.152939
R23390 GND.n4511 GND.n1974 0.152939
R23391 GND.n4584 GND.n1974 0.152939
R23392 GND.n4585 GND.n4584 0.152939
R23393 GND.n4586 GND.n4585 0.152939
R23394 GND.n4587 GND.n4586 0.152939
R23395 GND.n4587 GND.n1944 0.152939
R23396 GND.n4616 GND.n1944 0.152939
R23397 GND.n4617 GND.n4616 0.152939
R23398 GND.n4618 GND.n4617 0.152939
R23399 GND.n4618 GND.n1871 0.152939
R23400 GND.n4124 GND.n4093 0.152939
R23401 GND.n4096 GND.n4093 0.152939
R23402 GND.n4097 GND.n4096 0.152939
R23403 GND.n4098 GND.n4097 0.152939
R23404 GND.n4099 GND.n4098 0.152939
R23405 GND.n4102 GND.n4099 0.152939
R23406 GND.n4103 GND.n4102 0.152939
R23407 GND.n4104 GND.n4103 0.152939
R23408 GND.n4105 GND.n4104 0.152939
R23409 GND.n4106 GND.n4105 0.152939
R23410 GND.n4106 GND.n2060 0.152939
R23411 GND.n4436 GND.n2060 0.152939
R23412 GND.n4437 GND.n4436 0.152939
R23413 GND.n4438 GND.n4437 0.152939
R23414 GND.n4438 GND.n2056 0.152939
R23415 GND.n4444 GND.n2056 0.152939
R23416 GND.n4445 GND.n4444 0.152939
R23417 GND.n4446 GND.n4445 0.152939
R23418 GND.n4447 GND.n4446 0.152939
R23419 GND.n4447 GND.n1998 0.152939
R23420 GND.n4518 GND.n1998 0.152939
R23421 GND.n4519 GND.n4518 0.152939
R23422 GND.n4520 GND.n4519 0.152939
R23423 GND.n4520 GND.n1994 0.152939
R23424 GND.n4526 GND.n1994 0.152939
R23425 GND.n4527 GND.n4526 0.152939
R23426 GND.n4528 GND.n4527 0.152939
R23427 GND.n4529 GND.n4528 0.152939
R23428 GND.n4530 GND.n4529 0.152939
R23429 GND.n4533 GND.n4530 0.152939
R23430 GND.n4534 GND.n4533 0.152939
R23431 GND.n4535 GND.n4534 0.152939
R23432 GND.n3941 GND.n2246 0.152939
R23433 GND.n3942 GND.n3941 0.152939
R23434 GND.n3943 GND.n3942 0.152939
R23435 GND.n3943 GND.n2240 0.152939
R23436 GND.n3951 GND.n2240 0.152939
R23437 GND.n3952 GND.n3951 0.152939
R23438 GND.n3953 GND.n3952 0.152939
R23439 GND.n3953 GND.n2234 0.152939
R23440 GND.n3961 GND.n2234 0.152939
R23441 GND.n3962 GND.n3961 0.152939
R23442 GND.n3963 GND.n3962 0.152939
R23443 GND.n3963 GND.n2228 0.152939
R23444 GND.n3971 GND.n2228 0.152939
R23445 GND.n3972 GND.n3971 0.152939
R23446 GND.n3973 GND.n3972 0.152939
R23447 GND.n3973 GND.n2222 0.152939
R23448 GND.n3981 GND.n2222 0.152939
R23449 GND.n3982 GND.n3981 0.152939
R23450 GND.n3983 GND.n3982 0.152939
R23451 GND.n3983 GND.n2216 0.152939
R23452 GND.n3991 GND.n2216 0.152939
R23453 GND.n3992 GND.n3991 0.152939
R23454 GND.n3993 GND.n3992 0.152939
R23455 GND.n3993 GND.n2210 0.152939
R23456 GND.n4001 GND.n2210 0.152939
R23457 GND.n4002 GND.n4001 0.152939
R23458 GND.n4003 GND.n4002 0.152939
R23459 GND.n4003 GND.n2204 0.152939
R23460 GND.n4011 GND.n2204 0.152939
R23461 GND.n4012 GND.n4011 0.152939
R23462 GND.n4013 GND.n4012 0.152939
R23463 GND.n4013 GND.n2198 0.152939
R23464 GND.n4021 GND.n2198 0.152939
R23465 GND.n4022 GND.n4021 0.152939
R23466 GND.n4023 GND.n4022 0.152939
R23467 GND.n4023 GND.n2192 0.152939
R23468 GND.n4031 GND.n2192 0.152939
R23469 GND.n4032 GND.n4031 0.152939
R23470 GND.n4033 GND.n4032 0.152939
R23471 GND.n4033 GND.n2186 0.152939
R23472 GND.n4041 GND.n2186 0.152939
R23473 GND.n4042 GND.n4041 0.152939
R23474 GND.n4043 GND.n4042 0.152939
R23475 GND.n4043 GND.n2180 0.152939
R23476 GND.n4051 GND.n2180 0.152939
R23477 GND.n4052 GND.n4051 0.152939
R23478 GND.n4053 GND.n4052 0.152939
R23479 GND.n4053 GND.n2174 0.152939
R23480 GND.n4061 GND.n2174 0.152939
R23481 GND.n4062 GND.n4061 0.152939
R23482 GND.n4063 GND.n4062 0.152939
R23483 GND.n4063 GND.n2168 0.152939
R23484 GND.n4071 GND.n2168 0.152939
R23485 GND.n4072 GND.n4071 0.152939
R23486 GND.n4073 GND.n4072 0.152939
R23487 GND.n4073 GND.n2162 0.152939
R23488 GND.n4081 GND.n2162 0.152939
R23489 GND.n4082 GND.n4081 0.152939
R23490 GND.n4083 GND.n4082 0.152939
R23491 GND.n4083 GND.n2156 0.152939
R23492 GND.n4091 GND.n2156 0.152939
R23493 GND.n4092 GND.n4091 0.152939
R23494 GND.n4125 GND.n4092 0.152939
R23495 GND.n5910 GND.n5904 0.152939
R23496 GND.n5911 GND.n5910 0.152939
R23497 GND.n5912 GND.n5911 0.152939
R23498 GND.n5912 GND.n1671 0.152939
R23499 GND.n5920 GND.n1671 0.152939
R23500 GND.n5921 GND.n5920 0.152939
R23501 GND.n5922 GND.n5921 0.152939
R23502 GND.n5922 GND.n1669 0.152939
R23503 GND.n5932 GND.n1669 0.152939
R23504 GND.n5933 GND.n5932 0.152939
R23505 GND.n5934 GND.n5933 0.152939
R23506 GND.n5934 GND.n1667 0.152939
R23507 GND.n5942 GND.n1667 0.152939
R23508 GND.n5943 GND.n5942 0.152939
R23509 GND.n5944 GND.n5943 0.152939
R23510 GND.n5944 GND.n1665 0.152939
R23511 GND.n5951 GND.n1665 0.152939
R23512 GND.n5952 GND.n5951 0.152939
R23513 GND.n5952 GND.n1660 0.152939
R23514 GND.n5958 GND.n1660 0.152939
R23515 GND.n6038 GND.n6037 0.152939
R23516 GND.n6037 GND.n6036 0.152939
R23517 GND.n6036 GND.n5960 0.152939
R23518 GND.n5966 GND.n5960 0.152939
R23519 GND.n6031 GND.n5966 0.152939
R23520 GND.n6031 GND.n6030 0.152939
R23521 GND.n6030 GND.n6029 0.152939
R23522 GND.n6029 GND.n5971 0.152939
R23523 GND.n6025 GND.n5971 0.152939
R23524 GND.n6025 GND.n6024 0.152939
R23525 GND.n6024 GND.n6023 0.152939
R23526 GND.n6023 GND.n5977 0.152939
R23527 GND.n6019 GND.n5977 0.152939
R23528 GND.n6019 GND.n6018 0.152939
R23529 GND.n6018 GND.n6017 0.152939
R23530 GND.n6017 GND.n5985 0.152939
R23531 GND.n6013 GND.n5985 0.152939
R23532 GND.n6013 GND.n6012 0.152939
R23533 GND.n6012 GND.n6011 0.152939
R23534 GND.n6011 GND.n5991 0.152939
R23535 GND.n6007 GND.n5991 0.152939
R23536 GND.n6007 GND.n6006 0.152939
R23537 GND.n6006 GND.n6005 0.152939
R23538 GND.n6005 GND.n5997 0.152939
R23539 GND.n5997 GND.n1601 0.152939
R23540 GND.n4328 GND.n2138 0.152939
R23541 GND.n4324 GND.n2138 0.152939
R23542 GND.n4324 GND.n4323 0.152939
R23543 GND.n4323 GND.n4322 0.152939
R23544 GND.n4322 GND.n2142 0.152939
R23545 GND.n4318 GND.n2142 0.152939
R23546 GND.n4318 GND.n4317 0.152939
R23547 GND.n4317 GND.n4316 0.152939
R23548 GND.n2150 GND.n2118 0.152939
R23549 GND.n4358 GND.n2118 0.152939
R23550 GND.n4359 GND.n4358 0.152939
R23551 GND.n4361 GND.n4359 0.152939
R23552 GND.n4361 GND.n4360 0.152939
R23553 GND.n4360 GND.n2089 0.152939
R23554 GND.n4394 GND.n2089 0.152939
R23555 GND.n4395 GND.n4394 0.152939
R23556 GND.n4409 GND.n4395 0.152939
R23557 GND.n4409 GND.n4408 0.152939
R23558 GND.n4408 GND.n4407 0.152939
R23559 GND.n4407 GND.n4396 0.152939
R23560 GND.n4403 GND.n4396 0.152939
R23561 GND.n4403 GND.n4402 0.152939
R23562 GND.n4402 GND.n2026 0.152939
R23563 GND.n4476 GND.n2026 0.152939
R23564 GND.n4477 GND.n4476 0.152939
R23565 GND.n4491 GND.n4477 0.152939
R23566 GND.n4491 GND.n4490 0.152939
R23567 GND.n4490 GND.n4489 0.152939
R23568 GND.n4489 GND.n4478 0.152939
R23569 GND.n4485 GND.n4478 0.152939
R23570 GND.n4485 GND.n4484 0.152939
R23571 GND.n4484 GND.n1964 0.152939
R23572 GND.n4594 GND.n1964 0.152939
R23573 GND.n4595 GND.n4594 0.152939
R23574 GND.n4602 GND.n4595 0.152939
R23575 GND.n4602 GND.n4601 0.152939
R23576 GND.n4601 GND.n4600 0.152939
R23577 GND.n4600 GND.n4596 0.152939
R23578 GND.n4596 GND.n1934 0.152939
R23579 GND.n4628 GND.n1934 0.152939
R23580 GND.n4629 GND.n4628 0.152939
R23581 GND.n4630 GND.n4629 0.152939
R23582 GND.n4630 GND.n1917 0.152939
R23583 GND.n4644 GND.n1917 0.152939
R23584 GND.n6927 GND.n661 0.127024
R23585 GND.n6052 GND.n1593 0.127024
R23586 GND.n1873 GND.n1872 0.104159
R23587 GND.n7919 GND.n168 0.104159
R23588 GND.n8562 GND.n166 0.0767195
R23589 GND.n8562 GND.n167 0.0767195
R23590 GND.n4690 GND.n4689 0.0767195
R23591 GND.n4689 GND.n1871 0.0767195
R23592 GND.n4646 GND.n4645 0.0695946
R23593 GND.n8570 GND.n152 0.0695946
R23594 GND.n8570 GND.n8569 0.0695946
R23595 GND.n4645 GND.n4644 0.0695946
R23596 GND.n7731 GND.n660 0.063
R23597 GND.n6051 GND.n6050 0.063
R23598 GND.n8041 GND.n168 0.0492805
R23599 GND.n4535 GND.n1873 0.0492805
R23600 GND.n660 GND.n655 0.0412609
R23601 GND.n8460 GND.n349 0.0412609
R23602 GND.n4342 GND.n4329 0.0412609
R23603 GND.n6050 GND.n6049 0.0412609
R23604 GND.n7751 GND.n655 0.0344674
R23605 GND.n7751 GND.n656 0.0344674
R23606 GND.n7745 GND.n656 0.0344674
R23607 GND.n7745 GND.n7744 0.0344674
R23608 GND.n7744 GND.n629 0.0344674
R23609 GND.n629 GND.n626 0.0344674
R23610 GND.n627 GND.n626 0.0344674
R23611 GND.n7782 GND.n627 0.0344674
R23612 GND.n7783 GND.n7782 0.0344674
R23613 GND.n7783 GND.n601 0.0344674
R23614 GND.n601 GND.n599 0.0344674
R23615 GND.n7820 GND.n599 0.0344674
R23616 GND.n7821 GND.n7820 0.0344674
R23617 GND.n7821 GND.n576 0.0344674
R23618 GND.n7850 GND.n576 0.0344674
R23619 GND.n7850 GND.n561 0.0344674
R23620 GND.n7864 GND.n561 0.0344674
R23621 GND.n7865 GND.n7864 0.0344674
R23622 GND.n7865 GND.n543 0.0344674
R23623 GND.n544 GND.n543 0.0344674
R23624 GND.n7886 GND.n544 0.0344674
R23625 GND.n7886 GND.n545 0.0344674
R23626 GND.n545 GND.n512 0.0344674
R23627 GND.n513 GND.n512 0.0344674
R23628 GND.n514 GND.n513 0.0344674
R23629 GND.n515 GND.n514 0.0344674
R23630 GND.n515 GND.n488 0.0344674
R23631 GND.n488 GND.n485 0.0344674
R23632 GND.n486 GND.n485 0.0344674
R23633 GND.n7972 GND.n486 0.0344674
R23634 GND.n7973 GND.n7972 0.0344674
R23635 GND.n7973 GND.n459 0.0344674
R23636 GND.n8010 GND.n459 0.0344674
R23637 GND.n8011 GND.n8010 0.0344674
R23638 GND.n8011 GND.n447 0.0344674
R23639 GND.n447 GND.n445 0.0344674
R23640 GND.n8028 GND.n445 0.0344674
R23641 GND.n8028 GND.n432 0.0344674
R23642 GND.n8128 GND.n432 0.0344674
R23643 GND.n8129 GND.n8128 0.0344674
R23644 GND.n8129 GND.n184 0.0344674
R23645 GND.n185 GND.n184 0.0344674
R23646 GND.n186 GND.n185 0.0344674
R23647 GND.n8144 GND.n186 0.0344674
R23648 GND.n8144 GND.n204 0.0344674
R23649 GND.n205 GND.n204 0.0344674
R23650 GND.n206 GND.n205 0.0344674
R23651 GND.n8159 GND.n206 0.0344674
R23652 GND.n8159 GND.n225 0.0344674
R23653 GND.n226 GND.n225 0.0344674
R23654 GND.n227 GND.n226 0.0344674
R23655 GND.n8174 GND.n227 0.0344674
R23656 GND.n8174 GND.n246 0.0344674
R23657 GND.n247 GND.n246 0.0344674
R23658 GND.n248 GND.n247 0.0344674
R23659 GND.n8189 GND.n248 0.0344674
R23660 GND.n8189 GND.n266 0.0344674
R23661 GND.n267 GND.n266 0.0344674
R23662 GND.n268 GND.n267 0.0344674
R23663 GND.n8204 GND.n268 0.0344674
R23664 GND.n8204 GND.n287 0.0344674
R23665 GND.n288 GND.n287 0.0344674
R23666 GND.n289 GND.n288 0.0344674
R23667 GND.n8219 GND.n289 0.0344674
R23668 GND.n8219 GND.n308 0.0344674
R23669 GND.n309 GND.n308 0.0344674
R23670 GND.n310 GND.n309 0.0344674
R23671 GND.n8235 GND.n310 0.0344674
R23672 GND.n8235 GND.n328 0.0344674
R23673 GND.n329 GND.n328 0.0344674
R23674 GND.n330 GND.n329 0.0344674
R23675 GND.n348 GND.n330 0.0344674
R23676 GND.n8460 GND.n348 0.0344674
R23677 GND.n4342 GND.n4330 0.0344674
R23678 GND.n4338 GND.n4330 0.0344674
R23679 GND.n4338 GND.n4337 0.0344674
R23680 GND.n4337 GND.n2110 0.0344674
R23681 GND.n4378 GND.n2110 0.0344674
R23682 GND.n4378 GND.n2111 0.0344674
R23683 GND.n4374 GND.n2111 0.0344674
R23684 GND.n4374 GND.n4373 0.0344674
R23685 GND.n4373 GND.n2081 0.0344674
R23686 GND.n4421 GND.n2081 0.0344674
R23687 GND.n4421 GND.n2082 0.0344674
R23688 GND.n4417 GND.n2082 0.0344674
R23689 GND.n4417 GND.n2047 0.0344674
R23690 GND.n4460 GND.n2047 0.0344674
R23691 GND.n4460 GND.n2048 0.0344674
R23692 GND.n4456 GND.n2048 0.0344674
R23693 GND.n4456 GND.n4455 0.0344674
R23694 GND.n4455 GND.n2019 0.0344674
R23695 GND.n4503 GND.n2019 0.0344674
R23696 GND.n4503 GND.n2020 0.0344674
R23697 GND.n4499 GND.n2020 0.0344674
R23698 GND.n4499 GND.n1985 0.0344674
R23699 GND.n4578 GND.n1985 0.0344674
R23700 GND.n4578 GND.n1986 0.0344674
R23701 GND.n4574 GND.n1986 0.0344674
R23702 GND.n4574 GND.n4573 0.0344674
R23703 GND.n4573 GND.n1955 0.0344674
R23704 GND.n4610 GND.n1955 0.0344674
R23705 GND.n4610 GND.n1958 0.0344674
R23706 GND.n1958 GND.n1957 0.0344674
R23707 GND.n1957 GND.n1890 0.0344674
R23708 GND.n4682 GND.n1890 0.0344674
R23709 GND.n4682 GND.n1891 0.0344674
R23710 GND.n4678 GND.n1891 0.0344674
R23711 GND.n4678 GND.n4677 0.0344674
R23712 GND.n4677 GND.n4676 0.0344674
R23713 GND.n4676 GND.n1899 0.0344674
R23714 GND.n4672 GND.n1899 0.0344674
R23715 GND.n4672 GND.n4671 0.0344674
R23716 GND.n4671 GND.n4670 0.0344674
R23717 GND.n4670 GND.n1907 0.0344674
R23718 GND.n4666 GND.n1907 0.0344674
R23719 GND.n4666 GND.n1844 0.0344674
R23720 GND.n4737 GND.n1844 0.0344674
R23721 GND.n4737 GND.n1845 0.0344674
R23722 GND.n4733 GND.n1845 0.0344674
R23723 GND.n4733 GND.n4732 0.0344674
R23724 GND.n4732 GND.n1817 0.0344674
R23725 GND.n4775 GND.n1817 0.0344674
R23726 GND.n4775 GND.n1818 0.0344674
R23727 GND.n4771 GND.n1818 0.0344674
R23728 GND.n4771 GND.n4770 0.0344674
R23729 GND.n4770 GND.n1783 0.0344674
R23730 GND.n4843 GND.n1783 0.0344674
R23731 GND.n4843 GND.n1784 0.0344674
R23732 GND.n4839 GND.n1784 0.0344674
R23733 GND.n4839 GND.n4838 0.0344674
R23734 GND.n4838 GND.n1756 0.0344674
R23735 GND.n4880 GND.n1756 0.0344674
R23736 GND.n4880 GND.n1757 0.0344674
R23737 GND.n4876 GND.n1757 0.0344674
R23738 GND.n4876 GND.n4875 0.0344674
R23739 GND.n4875 GND.n1726 0.0344674
R23740 GND.n4918 GND.n1726 0.0344674
R23741 GND.n4918 GND.n1729 0.0344674
R23742 GND.n1729 GND.n1728 0.0344674
R23743 GND.n1728 GND.n1698 0.0344674
R23744 GND.n5878 GND.n1698 0.0344674
R23745 GND.n5878 GND.n1699 0.0344674
R23746 GND.n5874 GND.n1699 0.0344674
R23747 GND.n5874 GND.n5873 0.0344674
R23748 GND.n5873 GND.n1602 0.0344674
R23749 GND.n6049 GND.n1602 0.0344674
R23750 GND.n6065 GND.n6052 0.0111707
R23751 GND.n6966 GND.n661 0.0111707
R23752 VN.n198 VN.t1 243.97
R23753 VN.n198 VN.n197 223.454
R23754 VN.n200 VN.n199 223.454
R23755 VN.n202 VN.n201 223.454
R23756 VN.n194 VN.n193 161.3
R23757 VN.n192 VN.n99 161.3
R23758 VN.n191 VN.n190 161.3
R23759 VN.n189 VN.n100 161.3
R23760 VN.n188 VN.n187 161.3
R23761 VN.n186 VN.n101 161.3
R23762 VN.n185 VN.n184 161.3
R23763 VN.n183 VN.n102 161.3
R23764 VN.n182 VN.n181 161.3
R23765 VN.n180 VN.n103 161.3
R23766 VN.n179 VN.n178 161.3
R23767 VN.n177 VN.n104 161.3
R23768 VN.n176 VN.n175 161.3
R23769 VN.n174 VN.n105 161.3
R23770 VN.n173 VN.n172 161.3
R23771 VN.n171 VN.n106 161.3
R23772 VN.n170 VN.n169 161.3
R23773 VN.n167 VN.n107 161.3
R23774 VN.n166 VN.n165 161.3
R23775 VN.n164 VN.n108 161.3
R23776 VN.n163 VN.n162 161.3
R23777 VN.n161 VN.n109 161.3
R23778 VN.n160 VN.n159 161.3
R23779 VN.n158 VN.n110 161.3
R23780 VN.n157 VN.n156 161.3
R23781 VN.n155 VN.n111 161.3
R23782 VN.n154 VN.n153 161.3
R23783 VN.n152 VN.n112 161.3
R23784 VN.n151 VN.n150 161.3
R23785 VN.n149 VN.n113 161.3
R23786 VN.n148 VN.n147 161.3
R23787 VN.n146 VN.n145 161.3
R23788 VN.n144 VN.n115 161.3
R23789 VN.n143 VN.n142 161.3
R23790 VN.n141 VN.n116 161.3
R23791 VN.n140 VN.n139 161.3
R23792 VN.n138 VN.n117 161.3
R23793 VN.n137 VN.n136 161.3
R23794 VN.n135 VN.n118 161.3
R23795 VN.n134 VN.n133 161.3
R23796 VN.n132 VN.n119 161.3
R23797 VN.n131 VN.n130 161.3
R23798 VN.n129 VN.n120 161.3
R23799 VN.n128 VN.n127 161.3
R23800 VN.n126 VN.n121 161.3
R23801 VN.n125 VN.n124 161.3
R23802 VN.n28 VN.n27 161.3
R23803 VN.n29 VN.n24 161.3
R23804 VN.n31 VN.n30 161.3
R23805 VN.n32 VN.n23 161.3
R23806 VN.n34 VN.n33 161.3
R23807 VN.n35 VN.n22 161.3
R23808 VN.n37 VN.n36 161.3
R23809 VN.n38 VN.n21 161.3
R23810 VN.n40 VN.n39 161.3
R23811 VN.n41 VN.n20 161.3
R23812 VN.n43 VN.n42 161.3
R23813 VN.n44 VN.n19 161.3
R23814 VN.n46 VN.n45 161.3
R23815 VN.n47 VN.n18 161.3
R23816 VN.n49 VN.n48 161.3
R23817 VN.n51 VN.n50 161.3
R23818 VN.n52 VN.n16 161.3
R23819 VN.n54 VN.n53 161.3
R23820 VN.n55 VN.n15 161.3
R23821 VN.n57 VN.n56 161.3
R23822 VN.n58 VN.n14 161.3
R23823 VN.n60 VN.n59 161.3
R23824 VN.n61 VN.n13 161.3
R23825 VN.n63 VN.n62 161.3
R23826 VN.n64 VN.n12 161.3
R23827 VN.n66 VN.n65 161.3
R23828 VN.n67 VN.n11 161.3
R23829 VN.n69 VN.n68 161.3
R23830 VN.n70 VN.n9 161.3
R23831 VN.n72 VN.n71 161.3
R23832 VN.n73 VN.n8 161.3
R23833 VN.n75 VN.n74 161.3
R23834 VN.n76 VN.n7 161.3
R23835 VN.n78 VN.n77 161.3
R23836 VN.n79 VN.n6 161.3
R23837 VN.n81 VN.n80 161.3
R23838 VN.n82 VN.n5 161.3
R23839 VN.n84 VN.n83 161.3
R23840 VN.n85 VN.n4 161.3
R23841 VN.n87 VN.n86 161.3
R23842 VN.n88 VN.n3 161.3
R23843 VN.n90 VN.n89 161.3
R23844 VN.n91 VN.n2 161.3
R23845 VN.n93 VN.n92 161.3
R23846 VN.n94 VN.n1 161.3
R23847 VN.n96 VN.n95 161.3
R23848 VN.n195 VN.n98 68.3014
R23849 VN.n97 VN.n0 68.3014
R23850 VN.n196 VN.n195 60.5217
R23851 VN.n181 VN.n102 56.5193
R23852 VN.n83 VN.n4 56.5193
R23853 VN.n123 VN.n122 53.4399
R23854 VN.n26 VN.n25 53.4399
R23855 VN.n133 VN.n118 50.6917
R23856 VN.n160 VN.n110 50.6917
R23857 VN.n63 VN.n13 50.6917
R23858 VN.n36 VN.n21 50.6917
R23859 VN.n123 VN.t12 49.7746
R23860 VN.n26 VN.t13 49.7743
R23861 VN.n137 VN.n118 30.2951
R23862 VN.n156 VN.n110 30.2951
R23863 VN.n59 VN.n13 30.2951
R23864 VN.n40 VN.n21 30.2951
R23865 VN.n126 VN.n125 24.4675
R23866 VN.n127 VN.n126 24.4675
R23867 VN.n127 VN.n120 24.4675
R23868 VN.n131 VN.n120 24.4675
R23869 VN.n132 VN.n131 24.4675
R23870 VN.n133 VN.n132 24.4675
R23871 VN.n138 VN.n137 24.4675
R23872 VN.n139 VN.n138 24.4675
R23873 VN.n139 VN.n116 24.4675
R23874 VN.n143 VN.n116 24.4675
R23875 VN.n144 VN.n143 24.4675
R23876 VN.n145 VN.n144 24.4675
R23877 VN.n149 VN.n148 24.4675
R23878 VN.n150 VN.n149 24.4675
R23879 VN.n150 VN.n112 24.4675
R23880 VN.n154 VN.n112 24.4675
R23881 VN.n155 VN.n154 24.4675
R23882 VN.n156 VN.n155 24.4675
R23883 VN.n161 VN.n160 24.4675
R23884 VN.n162 VN.n161 24.4675
R23885 VN.n162 VN.n108 24.4675
R23886 VN.n166 VN.n108 24.4675
R23887 VN.n167 VN.n166 24.4675
R23888 VN.n169 VN.n167 24.4675
R23889 VN.n173 VN.n106 24.4675
R23890 VN.n174 VN.n173 24.4675
R23891 VN.n175 VN.n174 24.4675
R23892 VN.n175 VN.n104 24.4675
R23893 VN.n179 VN.n104 24.4675
R23894 VN.n180 VN.n179 24.4675
R23895 VN.n181 VN.n180 24.4675
R23896 VN.n185 VN.n102 24.4675
R23897 VN.n186 VN.n185 24.4675
R23898 VN.n187 VN.n186 24.4675
R23899 VN.n187 VN.n100 24.4675
R23900 VN.n191 VN.n100 24.4675
R23901 VN.n192 VN.n191 24.4675
R23902 VN.n193 VN.n192 24.4675
R23903 VN.n95 VN.n94 24.4675
R23904 VN.n94 VN.n93 24.4675
R23905 VN.n93 VN.n2 24.4675
R23906 VN.n89 VN.n2 24.4675
R23907 VN.n89 VN.n88 24.4675
R23908 VN.n88 VN.n87 24.4675
R23909 VN.n87 VN.n4 24.4675
R23910 VN.n83 VN.n82 24.4675
R23911 VN.n82 VN.n81 24.4675
R23912 VN.n81 VN.n6 24.4675
R23913 VN.n77 VN.n6 24.4675
R23914 VN.n77 VN.n76 24.4675
R23915 VN.n76 VN.n75 24.4675
R23916 VN.n75 VN.n8 24.4675
R23917 VN.n71 VN.n70 24.4675
R23918 VN.n70 VN.n69 24.4675
R23919 VN.n69 VN.n11 24.4675
R23920 VN.n65 VN.n11 24.4675
R23921 VN.n65 VN.n64 24.4675
R23922 VN.n64 VN.n63 24.4675
R23923 VN.n59 VN.n58 24.4675
R23924 VN.n58 VN.n57 24.4675
R23925 VN.n57 VN.n15 24.4675
R23926 VN.n53 VN.n15 24.4675
R23927 VN.n53 VN.n52 24.4675
R23928 VN.n52 VN.n51 24.4675
R23929 VN.n48 VN.n47 24.4675
R23930 VN.n47 VN.n46 24.4675
R23931 VN.n46 VN.n19 24.4675
R23932 VN.n42 VN.n19 24.4675
R23933 VN.n42 VN.n41 24.4675
R23934 VN.n41 VN.n40 24.4675
R23935 VN.n36 VN.n35 24.4675
R23936 VN.n35 VN.n34 24.4675
R23937 VN.n34 VN.n23 24.4675
R23938 VN.n30 VN.n23 24.4675
R23939 VN.n30 VN.n29 24.4675
R23940 VN.n29 VN.n28 24.4675
R23941 VN.n125 VN.n122 22.5101
R23942 VN.n169 VN.n168 22.5101
R23943 VN.n71 VN.n10 22.5101
R23944 VN.n28 VN.n25 22.5101
R23945 VN.n197 VN.t2 19.8005
R23946 VN.n197 VN.t0 19.8005
R23947 VN.n199 VN.t3 19.8005
R23948 VN.n199 VN.t5 19.8005
R23949 VN.n201 VN.t4 19.8005
R23950 VN.n201 VN.t6 19.8005
R23951 VN VN.n203 19.0806
R23952 VN.n122 VN.t16 15.708
R23953 VN.n114 VN.t15 15.708
R23954 VN.n168 VN.t8 15.708
R23955 VN.n98 VN.t7 15.708
R23956 VN.n0 VN.t14 15.708
R23957 VN.n10 VN.t10 15.708
R23958 VN.n17 VN.t11 15.708
R23959 VN.n25 VN.t9 15.708
R23960 VN.n196 VN.n97 14.3171
R23961 VN.n145 VN.n114 12.234
R23962 VN.n148 VN.n114 12.234
R23963 VN.n51 VN.n17 12.234
R23964 VN.n48 VN.n17 12.234
R23965 VN.n193 VN.n98 8.31928
R23966 VN.n95 VN.n0 8.31928
R23967 VN.n203 VN.n202 5.40567
R23968 VN.n168 VN.n106 1.95786
R23969 VN.n10 VN.n8 1.95786
R23970 VN.n203 VN.n196 1.188
R23971 VN.n202 VN.n200 0.716017
R23972 VN.n200 VN.n198 0.716017
R23973 VN.n124 VN.n123 0.690479
R23974 VN.n27 VN.n26 0.690478
R23975 VN.n195 VN.n194 0.529113
R23976 VN.n97 VN.n96 0.529113
R23977 VN.n124 VN.n121 0.189894
R23978 VN.n128 VN.n121 0.189894
R23979 VN.n129 VN.n128 0.189894
R23980 VN.n130 VN.n129 0.189894
R23981 VN.n130 VN.n119 0.189894
R23982 VN.n134 VN.n119 0.189894
R23983 VN.n135 VN.n134 0.189894
R23984 VN.n136 VN.n135 0.189894
R23985 VN.n136 VN.n117 0.189894
R23986 VN.n140 VN.n117 0.189894
R23987 VN.n141 VN.n140 0.189894
R23988 VN.n142 VN.n141 0.189894
R23989 VN.n142 VN.n115 0.189894
R23990 VN.n146 VN.n115 0.189894
R23991 VN.n147 VN.n146 0.189894
R23992 VN.n147 VN.n113 0.189894
R23993 VN.n151 VN.n113 0.189894
R23994 VN.n152 VN.n151 0.189894
R23995 VN.n153 VN.n152 0.189894
R23996 VN.n153 VN.n111 0.189894
R23997 VN.n157 VN.n111 0.189894
R23998 VN.n158 VN.n157 0.189894
R23999 VN.n159 VN.n158 0.189894
R24000 VN.n159 VN.n109 0.189894
R24001 VN.n163 VN.n109 0.189894
R24002 VN.n164 VN.n163 0.189894
R24003 VN.n165 VN.n164 0.189894
R24004 VN.n165 VN.n107 0.189894
R24005 VN.n170 VN.n107 0.189894
R24006 VN.n171 VN.n170 0.189894
R24007 VN.n172 VN.n171 0.189894
R24008 VN.n172 VN.n105 0.189894
R24009 VN.n176 VN.n105 0.189894
R24010 VN.n177 VN.n176 0.189894
R24011 VN.n178 VN.n177 0.189894
R24012 VN.n178 VN.n103 0.189894
R24013 VN.n182 VN.n103 0.189894
R24014 VN.n183 VN.n182 0.189894
R24015 VN.n184 VN.n183 0.189894
R24016 VN.n184 VN.n101 0.189894
R24017 VN.n188 VN.n101 0.189894
R24018 VN.n189 VN.n188 0.189894
R24019 VN.n190 VN.n189 0.189894
R24020 VN.n190 VN.n99 0.189894
R24021 VN.n194 VN.n99 0.189894
R24022 VN.n96 VN.n1 0.189894
R24023 VN.n92 VN.n1 0.189894
R24024 VN.n92 VN.n91 0.189894
R24025 VN.n91 VN.n90 0.189894
R24026 VN.n90 VN.n3 0.189894
R24027 VN.n86 VN.n3 0.189894
R24028 VN.n86 VN.n85 0.189894
R24029 VN.n85 VN.n84 0.189894
R24030 VN.n84 VN.n5 0.189894
R24031 VN.n80 VN.n5 0.189894
R24032 VN.n80 VN.n79 0.189894
R24033 VN.n79 VN.n78 0.189894
R24034 VN.n78 VN.n7 0.189894
R24035 VN.n74 VN.n7 0.189894
R24036 VN.n74 VN.n73 0.189894
R24037 VN.n73 VN.n72 0.189894
R24038 VN.n72 VN.n9 0.189894
R24039 VN.n68 VN.n9 0.189894
R24040 VN.n68 VN.n67 0.189894
R24041 VN.n67 VN.n66 0.189894
R24042 VN.n66 VN.n12 0.189894
R24043 VN.n62 VN.n12 0.189894
R24044 VN.n62 VN.n61 0.189894
R24045 VN.n61 VN.n60 0.189894
R24046 VN.n60 VN.n14 0.189894
R24047 VN.n56 VN.n14 0.189894
R24048 VN.n56 VN.n55 0.189894
R24049 VN.n55 VN.n54 0.189894
R24050 VN.n54 VN.n16 0.189894
R24051 VN.n50 VN.n16 0.189894
R24052 VN.n50 VN.n49 0.189894
R24053 VN.n49 VN.n18 0.189894
R24054 VN.n45 VN.n18 0.189894
R24055 VN.n45 VN.n44 0.189894
R24056 VN.n44 VN.n43 0.189894
R24057 VN.n43 VN.n20 0.189894
R24058 VN.n39 VN.n20 0.189894
R24059 VN.n39 VN.n38 0.189894
R24060 VN.n38 VN.n37 0.189894
R24061 VN.n37 VN.n22 0.189894
R24062 VN.n33 VN.n22 0.189894
R24063 VN.n33 VN.n32 0.189894
R24064 VN.n32 VN.n31 0.189894
R24065 VN.n31 VN.n24 0.189894
R24066 VN.n27 VN.n24 0.189894
R24067 VP.n202 VP.t5 243.255
R24068 VP.n199 VP.n197 224.169
R24069 VP.n201 VP.n200 223.454
R24070 VP.n199 VP.n198 223.454
R24071 VP.n126 VP.n125 161.3
R24072 VP.n127 VP.n122 161.3
R24073 VP.n129 VP.n128 161.3
R24074 VP.n130 VP.n121 161.3
R24075 VP.n132 VP.n131 161.3
R24076 VP.n133 VP.n120 161.3
R24077 VP.n135 VP.n134 161.3
R24078 VP.n136 VP.n119 161.3
R24079 VP.n138 VP.n137 161.3
R24080 VP.n139 VP.n118 161.3
R24081 VP.n141 VP.n140 161.3
R24082 VP.n142 VP.n117 161.3
R24083 VP.n144 VP.n143 161.3
R24084 VP.n145 VP.n116 161.3
R24085 VP.n147 VP.n146 161.3
R24086 VP.n149 VP.n148 161.3
R24087 VP.n150 VP.n114 161.3
R24088 VP.n152 VP.n151 161.3
R24089 VP.n153 VP.n113 161.3
R24090 VP.n155 VP.n154 161.3
R24091 VP.n156 VP.n112 161.3
R24092 VP.n158 VP.n157 161.3
R24093 VP.n159 VP.n111 161.3
R24094 VP.n161 VP.n160 161.3
R24095 VP.n162 VP.n110 161.3
R24096 VP.n164 VP.n163 161.3
R24097 VP.n165 VP.n109 161.3
R24098 VP.n167 VP.n166 161.3
R24099 VP.n168 VP.n107 161.3
R24100 VP.n170 VP.n169 161.3
R24101 VP.n171 VP.n106 161.3
R24102 VP.n173 VP.n172 161.3
R24103 VP.n174 VP.n105 161.3
R24104 VP.n176 VP.n175 161.3
R24105 VP.n177 VP.n104 161.3
R24106 VP.n179 VP.n178 161.3
R24107 VP.n180 VP.n103 161.3
R24108 VP.n182 VP.n181 161.3
R24109 VP.n183 VP.n102 161.3
R24110 VP.n185 VP.n184 161.3
R24111 VP.n186 VP.n101 161.3
R24112 VP.n188 VP.n187 161.3
R24113 VP.n189 VP.n100 161.3
R24114 VP.n191 VP.n190 161.3
R24115 VP.n192 VP.n99 161.3
R24116 VP.n194 VP.n193 161.3
R24117 VP.n96 VP.n95 161.3
R24118 VP.n94 VP.n1 161.3
R24119 VP.n93 VP.n92 161.3
R24120 VP.n91 VP.n2 161.3
R24121 VP.n90 VP.n89 161.3
R24122 VP.n88 VP.n3 161.3
R24123 VP.n87 VP.n86 161.3
R24124 VP.n85 VP.n4 161.3
R24125 VP.n84 VP.n83 161.3
R24126 VP.n82 VP.n5 161.3
R24127 VP.n81 VP.n80 161.3
R24128 VP.n79 VP.n6 161.3
R24129 VP.n78 VP.n77 161.3
R24130 VP.n76 VP.n7 161.3
R24131 VP.n75 VP.n74 161.3
R24132 VP.n73 VP.n8 161.3
R24133 VP.n72 VP.n71 161.3
R24134 VP.n69 VP.n9 161.3
R24135 VP.n68 VP.n67 161.3
R24136 VP.n66 VP.n10 161.3
R24137 VP.n65 VP.n64 161.3
R24138 VP.n63 VP.n11 161.3
R24139 VP.n62 VP.n61 161.3
R24140 VP.n60 VP.n12 161.3
R24141 VP.n59 VP.n58 161.3
R24142 VP.n57 VP.n13 161.3
R24143 VP.n56 VP.n55 161.3
R24144 VP.n54 VP.n14 161.3
R24145 VP.n53 VP.n52 161.3
R24146 VP.n51 VP.n15 161.3
R24147 VP.n50 VP.n49 161.3
R24148 VP.n48 VP.n47 161.3
R24149 VP.n46 VP.n17 161.3
R24150 VP.n45 VP.n44 161.3
R24151 VP.n43 VP.n18 161.3
R24152 VP.n42 VP.n41 161.3
R24153 VP.n40 VP.n19 161.3
R24154 VP.n39 VP.n38 161.3
R24155 VP.n37 VP.n20 161.3
R24156 VP.n36 VP.n35 161.3
R24157 VP.n34 VP.n21 161.3
R24158 VP.n33 VP.n32 161.3
R24159 VP.n31 VP.n22 161.3
R24160 VP.n30 VP.n29 161.3
R24161 VP.n28 VP.n23 161.3
R24162 VP.n27 VP.n26 161.3
R24163 VP.n195 VP.n98 68.3014
R24164 VP.n97 VP.n0 68.3014
R24165 VP.n196 VP.n195 60.7376
R24166 VP.n181 VP.n102 56.5193
R24167 VP.n83 VP.n4 56.5193
R24168 VP.n124 VP.n123 53.4399
R24169 VP.n25 VP.n24 53.4399
R24170 VP.n161 VP.n111 50.6917
R24171 VP.n134 VP.n119 50.6917
R24172 VP.n35 VP.n20 50.6917
R24173 VP.n62 VP.n12 50.6917
R24174 VP.n25 VP.t14 49.7746
R24175 VP.n124 VP.t12 49.7743
R24176 VP.n157 VP.n111 30.2951
R24177 VP.n138 VP.n119 30.2951
R24178 VP.n39 VP.n20 30.2951
R24179 VP.n58 VP.n12 30.2951
R24180 VP.n193 VP.n192 24.4675
R24181 VP.n192 VP.n191 24.4675
R24182 VP.n191 VP.n100 24.4675
R24183 VP.n187 VP.n100 24.4675
R24184 VP.n187 VP.n186 24.4675
R24185 VP.n186 VP.n185 24.4675
R24186 VP.n185 VP.n102 24.4675
R24187 VP.n181 VP.n180 24.4675
R24188 VP.n180 VP.n179 24.4675
R24189 VP.n179 VP.n104 24.4675
R24190 VP.n175 VP.n104 24.4675
R24191 VP.n175 VP.n174 24.4675
R24192 VP.n174 VP.n173 24.4675
R24193 VP.n173 VP.n106 24.4675
R24194 VP.n169 VP.n168 24.4675
R24195 VP.n168 VP.n167 24.4675
R24196 VP.n167 VP.n109 24.4675
R24197 VP.n163 VP.n109 24.4675
R24198 VP.n163 VP.n162 24.4675
R24199 VP.n162 VP.n161 24.4675
R24200 VP.n157 VP.n156 24.4675
R24201 VP.n156 VP.n155 24.4675
R24202 VP.n155 VP.n113 24.4675
R24203 VP.n151 VP.n113 24.4675
R24204 VP.n151 VP.n150 24.4675
R24205 VP.n150 VP.n149 24.4675
R24206 VP.n146 VP.n145 24.4675
R24207 VP.n145 VP.n144 24.4675
R24208 VP.n144 VP.n117 24.4675
R24209 VP.n140 VP.n117 24.4675
R24210 VP.n140 VP.n139 24.4675
R24211 VP.n139 VP.n138 24.4675
R24212 VP.n134 VP.n133 24.4675
R24213 VP.n133 VP.n132 24.4675
R24214 VP.n132 VP.n121 24.4675
R24215 VP.n128 VP.n121 24.4675
R24216 VP.n128 VP.n127 24.4675
R24217 VP.n127 VP.n126 24.4675
R24218 VP.n28 VP.n27 24.4675
R24219 VP.n29 VP.n28 24.4675
R24220 VP.n29 VP.n22 24.4675
R24221 VP.n33 VP.n22 24.4675
R24222 VP.n34 VP.n33 24.4675
R24223 VP.n35 VP.n34 24.4675
R24224 VP.n40 VP.n39 24.4675
R24225 VP.n41 VP.n40 24.4675
R24226 VP.n41 VP.n18 24.4675
R24227 VP.n45 VP.n18 24.4675
R24228 VP.n46 VP.n45 24.4675
R24229 VP.n47 VP.n46 24.4675
R24230 VP.n51 VP.n50 24.4675
R24231 VP.n52 VP.n51 24.4675
R24232 VP.n52 VP.n14 24.4675
R24233 VP.n56 VP.n14 24.4675
R24234 VP.n57 VP.n56 24.4675
R24235 VP.n58 VP.n57 24.4675
R24236 VP.n63 VP.n62 24.4675
R24237 VP.n64 VP.n63 24.4675
R24238 VP.n64 VP.n10 24.4675
R24239 VP.n68 VP.n10 24.4675
R24240 VP.n69 VP.n68 24.4675
R24241 VP.n71 VP.n69 24.4675
R24242 VP.n75 VP.n8 24.4675
R24243 VP.n76 VP.n75 24.4675
R24244 VP.n77 VP.n76 24.4675
R24245 VP.n77 VP.n6 24.4675
R24246 VP.n81 VP.n6 24.4675
R24247 VP.n82 VP.n81 24.4675
R24248 VP.n83 VP.n82 24.4675
R24249 VP.n87 VP.n4 24.4675
R24250 VP.n88 VP.n87 24.4675
R24251 VP.n89 VP.n88 24.4675
R24252 VP.n89 VP.n2 24.4675
R24253 VP.n93 VP.n2 24.4675
R24254 VP.n94 VP.n93 24.4675
R24255 VP.n95 VP.n94 24.4675
R24256 VP.n169 VP.n108 22.5101
R24257 VP.n126 VP.n123 22.5101
R24258 VP.n27 VP.n24 22.5101
R24259 VP.n71 VP.n70 22.5101
R24260 VP.n200 VP.t6 19.8005
R24261 VP.n200 VP.t2 19.8005
R24262 VP.n198 VP.t4 19.8005
R24263 VP.n198 VP.t1 19.8005
R24264 VP.n197 VP.t3 19.8005
R24265 VP.n197 VP.t0 19.8005
R24266 VP.n98 VP.t13 15.708
R24267 VP.n108 VP.t8 15.708
R24268 VP.n115 VP.t9 15.708
R24269 VP.n123 VP.t7 15.708
R24270 VP.n24 VP.t15 15.708
R24271 VP.n16 VP.t16 15.708
R24272 VP.n70 VP.t11 15.708
R24273 VP.n0 VP.t10 15.708
R24274 VP.n196 VP.n97 14.533
R24275 VP.n149 VP.n115 12.234
R24276 VP.n146 VP.n115 12.234
R24277 VP.n47 VP.n16 12.234
R24278 VP.n50 VP.n16 12.234
R24279 VP VP.n203 11.8096
R24280 VP.n193 VP.n98 8.31928
R24281 VP.n95 VP.n0 8.31928
R24282 VP.n203 VP.n202 4.80222
R24283 VP.n108 VP.n106 1.95786
R24284 VP.n70 VP.n8 1.95786
R24285 VP.n203 VP.n196 0.972091
R24286 VP.n201 VP.n199 0.716017
R24287 VP.n202 VP.n201 0.716017
R24288 VP.n26 VP.n25 0.690479
R24289 VP.n125 VP.n124 0.690478
R24290 VP.n195 VP.n194 0.529113
R24291 VP.n97 VP.n96 0.529113
R24292 VP.n194 VP.n99 0.189894
R24293 VP.n190 VP.n99 0.189894
R24294 VP.n190 VP.n189 0.189894
R24295 VP.n189 VP.n188 0.189894
R24296 VP.n188 VP.n101 0.189894
R24297 VP.n184 VP.n101 0.189894
R24298 VP.n184 VP.n183 0.189894
R24299 VP.n183 VP.n182 0.189894
R24300 VP.n182 VP.n103 0.189894
R24301 VP.n178 VP.n103 0.189894
R24302 VP.n178 VP.n177 0.189894
R24303 VP.n177 VP.n176 0.189894
R24304 VP.n176 VP.n105 0.189894
R24305 VP.n172 VP.n105 0.189894
R24306 VP.n172 VP.n171 0.189894
R24307 VP.n171 VP.n170 0.189894
R24308 VP.n170 VP.n107 0.189894
R24309 VP.n166 VP.n107 0.189894
R24310 VP.n166 VP.n165 0.189894
R24311 VP.n165 VP.n164 0.189894
R24312 VP.n164 VP.n110 0.189894
R24313 VP.n160 VP.n110 0.189894
R24314 VP.n160 VP.n159 0.189894
R24315 VP.n159 VP.n158 0.189894
R24316 VP.n158 VP.n112 0.189894
R24317 VP.n154 VP.n112 0.189894
R24318 VP.n154 VP.n153 0.189894
R24319 VP.n153 VP.n152 0.189894
R24320 VP.n152 VP.n114 0.189894
R24321 VP.n148 VP.n114 0.189894
R24322 VP.n148 VP.n147 0.189894
R24323 VP.n147 VP.n116 0.189894
R24324 VP.n143 VP.n116 0.189894
R24325 VP.n143 VP.n142 0.189894
R24326 VP.n142 VP.n141 0.189894
R24327 VP.n141 VP.n118 0.189894
R24328 VP.n137 VP.n118 0.189894
R24329 VP.n137 VP.n136 0.189894
R24330 VP.n136 VP.n135 0.189894
R24331 VP.n135 VP.n120 0.189894
R24332 VP.n131 VP.n120 0.189894
R24333 VP.n131 VP.n130 0.189894
R24334 VP.n130 VP.n129 0.189894
R24335 VP.n129 VP.n122 0.189894
R24336 VP.n125 VP.n122 0.189894
R24337 VP.n26 VP.n23 0.189894
R24338 VP.n30 VP.n23 0.189894
R24339 VP.n31 VP.n30 0.189894
R24340 VP.n32 VP.n31 0.189894
R24341 VP.n32 VP.n21 0.189894
R24342 VP.n36 VP.n21 0.189894
R24343 VP.n37 VP.n36 0.189894
R24344 VP.n38 VP.n37 0.189894
R24345 VP.n38 VP.n19 0.189894
R24346 VP.n42 VP.n19 0.189894
R24347 VP.n43 VP.n42 0.189894
R24348 VP.n44 VP.n43 0.189894
R24349 VP.n44 VP.n17 0.189894
R24350 VP.n48 VP.n17 0.189894
R24351 VP.n49 VP.n48 0.189894
R24352 VP.n49 VP.n15 0.189894
R24353 VP.n53 VP.n15 0.189894
R24354 VP.n54 VP.n53 0.189894
R24355 VP.n55 VP.n54 0.189894
R24356 VP.n55 VP.n13 0.189894
R24357 VP.n59 VP.n13 0.189894
R24358 VP.n60 VP.n59 0.189894
R24359 VP.n61 VP.n60 0.189894
R24360 VP.n61 VP.n11 0.189894
R24361 VP.n65 VP.n11 0.189894
R24362 VP.n66 VP.n65 0.189894
R24363 VP.n67 VP.n66 0.189894
R24364 VP.n67 VP.n9 0.189894
R24365 VP.n72 VP.n9 0.189894
R24366 VP.n73 VP.n72 0.189894
R24367 VP.n74 VP.n73 0.189894
R24368 VP.n74 VP.n7 0.189894
R24369 VP.n78 VP.n7 0.189894
R24370 VP.n79 VP.n78 0.189894
R24371 VP.n80 VP.n79 0.189894
R24372 VP.n80 VP.n5 0.189894
R24373 VP.n84 VP.n5 0.189894
R24374 VP.n85 VP.n84 0.189894
R24375 VP.n86 VP.n85 0.189894
R24376 VP.n86 VP.n3 0.189894
R24377 VP.n90 VP.n3 0.189894
R24378 VP.n91 VP.n90 0.189894
R24379 VP.n92 VP.n91 0.189894
R24380 VP.n92 VP.n1 0.189894
R24381 VP.n96 VP.n1 0.189894
R24382 CS_BIAS.n75 CS_BIAS.n73 289.615
R24383 CS_BIAS.n406 CS_BIAS.n404 289.615
R24384 CS_BIAS.n76 CS_BIAS.n75 185
R24385 CS_BIAS.n407 CS_BIAS.n406 185
R24386 CS_BIAS.t1 CS_BIAS.n74 167.117
R24387 CS_BIAS.t11 CS_BIAS.n405 167.117
R24388 CS_BIAS.n390 CS_BIAS.n330 161.3
R24389 CS_BIAS.n389 CS_BIAS.n388 161.3
R24390 CS_BIAS.n387 CS_BIAS.n331 161.3
R24391 CS_BIAS.n386 CS_BIAS.n385 161.3
R24392 CS_BIAS.n384 CS_BIAS.n332 161.3
R24393 CS_BIAS.n383 CS_BIAS.n382 161.3
R24394 CS_BIAS.n381 CS_BIAS.n333 161.3
R24395 CS_BIAS.n380 CS_BIAS.n379 161.3
R24396 CS_BIAS.n378 CS_BIAS.n334 161.3
R24397 CS_BIAS.n377 CS_BIAS.n376 161.3
R24398 CS_BIAS.n375 CS_BIAS.n374 161.3
R24399 CS_BIAS.n373 CS_BIAS.n336 161.3
R24400 CS_BIAS.n372 CS_BIAS.n371 161.3
R24401 CS_BIAS.n370 CS_BIAS.n337 161.3
R24402 CS_BIAS.n369 CS_BIAS.n368 161.3
R24403 CS_BIAS.n367 CS_BIAS.n338 161.3
R24404 CS_BIAS.n366 CS_BIAS.n365 161.3
R24405 CS_BIAS.n364 CS_BIAS.n339 161.3
R24406 CS_BIAS.n363 CS_BIAS.n362 161.3
R24407 CS_BIAS.n361 CS_BIAS.n340 161.3
R24408 CS_BIAS.n360 CS_BIAS.n359 161.3
R24409 CS_BIAS.n358 CS_BIAS.n341 161.3
R24410 CS_BIAS.n357 CS_BIAS.n356 161.3
R24411 CS_BIAS.n355 CS_BIAS.n342 161.3
R24412 CS_BIAS.n354 CS_BIAS.n353 161.3
R24413 CS_BIAS.n352 CS_BIAS.n343 161.3
R24414 CS_BIAS.n351 CS_BIAS.n350 161.3
R24415 CS_BIAS.n349 CS_BIAS.n344 161.3
R24416 CS_BIAS.n348 CS_BIAS.n347 161.3
R24417 CS_BIAS.n284 CS_BIAS.n283 161.3
R24418 CS_BIAS.n285 CS_BIAS.n280 161.3
R24419 CS_BIAS.n287 CS_BIAS.n286 161.3
R24420 CS_BIAS.n288 CS_BIAS.n279 161.3
R24421 CS_BIAS.n290 CS_BIAS.n289 161.3
R24422 CS_BIAS.n291 CS_BIAS.n278 161.3
R24423 CS_BIAS.n293 CS_BIAS.n292 161.3
R24424 CS_BIAS.n294 CS_BIAS.n277 161.3
R24425 CS_BIAS.n296 CS_BIAS.n295 161.3
R24426 CS_BIAS.n297 CS_BIAS.n276 161.3
R24427 CS_BIAS.n299 CS_BIAS.n298 161.3
R24428 CS_BIAS.n300 CS_BIAS.n275 161.3
R24429 CS_BIAS.n302 CS_BIAS.n301 161.3
R24430 CS_BIAS.n303 CS_BIAS.n274 161.3
R24431 CS_BIAS.n305 CS_BIAS.n304 161.3
R24432 CS_BIAS.n306 CS_BIAS.n273 161.3
R24433 CS_BIAS.n308 CS_BIAS.n307 161.3
R24434 CS_BIAS.n309 CS_BIAS.n272 161.3
R24435 CS_BIAS.n311 CS_BIAS.n310 161.3
R24436 CS_BIAS.n313 CS_BIAS.n312 161.3
R24437 CS_BIAS.n314 CS_BIAS.n270 161.3
R24438 CS_BIAS.n316 CS_BIAS.n315 161.3
R24439 CS_BIAS.n317 CS_BIAS.n269 161.3
R24440 CS_BIAS.n319 CS_BIAS.n318 161.3
R24441 CS_BIAS.n320 CS_BIAS.n268 161.3
R24442 CS_BIAS.n322 CS_BIAS.n321 161.3
R24443 CS_BIAS.n323 CS_BIAS.n267 161.3
R24444 CS_BIAS.n325 CS_BIAS.n324 161.3
R24445 CS_BIAS.n326 CS_BIAS.n266 161.3
R24446 CS_BIAS.n220 CS_BIAS.n219 161.3
R24447 CS_BIAS.n221 CS_BIAS.n216 161.3
R24448 CS_BIAS.n223 CS_BIAS.n222 161.3
R24449 CS_BIAS.n224 CS_BIAS.n215 161.3
R24450 CS_BIAS.n226 CS_BIAS.n225 161.3
R24451 CS_BIAS.n227 CS_BIAS.n214 161.3
R24452 CS_BIAS.n229 CS_BIAS.n228 161.3
R24453 CS_BIAS.n230 CS_BIAS.n213 161.3
R24454 CS_BIAS.n232 CS_BIAS.n231 161.3
R24455 CS_BIAS.n233 CS_BIAS.n212 161.3
R24456 CS_BIAS.n235 CS_BIAS.n234 161.3
R24457 CS_BIAS.n236 CS_BIAS.n211 161.3
R24458 CS_BIAS.n238 CS_BIAS.n237 161.3
R24459 CS_BIAS.n239 CS_BIAS.n210 161.3
R24460 CS_BIAS.n241 CS_BIAS.n240 161.3
R24461 CS_BIAS.n242 CS_BIAS.n209 161.3
R24462 CS_BIAS.n244 CS_BIAS.n243 161.3
R24463 CS_BIAS.n245 CS_BIAS.n208 161.3
R24464 CS_BIAS.n247 CS_BIAS.n246 161.3
R24465 CS_BIAS.n249 CS_BIAS.n248 161.3
R24466 CS_BIAS.n250 CS_BIAS.n206 161.3
R24467 CS_BIAS.n252 CS_BIAS.n251 161.3
R24468 CS_BIAS.n253 CS_BIAS.n205 161.3
R24469 CS_BIAS.n255 CS_BIAS.n254 161.3
R24470 CS_BIAS.n256 CS_BIAS.n204 161.3
R24471 CS_BIAS.n258 CS_BIAS.n257 161.3
R24472 CS_BIAS.n259 CS_BIAS.n203 161.3
R24473 CS_BIAS.n261 CS_BIAS.n260 161.3
R24474 CS_BIAS.n262 CS_BIAS.n202 161.3
R24475 CS_BIAS.n156 CS_BIAS.n155 161.3
R24476 CS_BIAS.n157 CS_BIAS.n152 161.3
R24477 CS_BIAS.n159 CS_BIAS.n158 161.3
R24478 CS_BIAS.n160 CS_BIAS.n151 161.3
R24479 CS_BIAS.n162 CS_BIAS.n161 161.3
R24480 CS_BIAS.n163 CS_BIAS.n150 161.3
R24481 CS_BIAS.n165 CS_BIAS.n164 161.3
R24482 CS_BIAS.n166 CS_BIAS.n149 161.3
R24483 CS_BIAS.n168 CS_BIAS.n167 161.3
R24484 CS_BIAS.n169 CS_BIAS.n148 161.3
R24485 CS_BIAS.n171 CS_BIAS.n170 161.3
R24486 CS_BIAS.n172 CS_BIAS.n147 161.3
R24487 CS_BIAS.n174 CS_BIAS.n173 161.3
R24488 CS_BIAS.n175 CS_BIAS.n146 161.3
R24489 CS_BIAS.n177 CS_BIAS.n176 161.3
R24490 CS_BIAS.n178 CS_BIAS.n145 161.3
R24491 CS_BIAS.n180 CS_BIAS.n179 161.3
R24492 CS_BIAS.n181 CS_BIAS.n144 161.3
R24493 CS_BIAS.n183 CS_BIAS.n182 161.3
R24494 CS_BIAS.n185 CS_BIAS.n184 161.3
R24495 CS_BIAS.n186 CS_BIAS.n142 161.3
R24496 CS_BIAS.n188 CS_BIAS.n187 161.3
R24497 CS_BIAS.n189 CS_BIAS.n141 161.3
R24498 CS_BIAS.n191 CS_BIAS.n190 161.3
R24499 CS_BIAS.n192 CS_BIAS.n140 161.3
R24500 CS_BIAS.n194 CS_BIAS.n193 161.3
R24501 CS_BIAS.n195 CS_BIAS.n139 161.3
R24502 CS_BIAS.n197 CS_BIAS.n196 161.3
R24503 CS_BIAS.n198 CS_BIAS.n138 161.3
R24504 CS_BIAS.n28 CS_BIAS.n27 161.3
R24505 CS_BIAS.n29 CS_BIAS.n24 161.3
R24506 CS_BIAS.n31 CS_BIAS.n30 161.3
R24507 CS_BIAS.n32 CS_BIAS.n23 161.3
R24508 CS_BIAS.n34 CS_BIAS.n33 161.3
R24509 CS_BIAS.n35 CS_BIAS.n22 161.3
R24510 CS_BIAS.n37 CS_BIAS.n36 161.3
R24511 CS_BIAS.n38 CS_BIAS.n21 161.3
R24512 CS_BIAS.n40 CS_BIAS.n39 161.3
R24513 CS_BIAS.n41 CS_BIAS.n20 161.3
R24514 CS_BIAS.n43 CS_BIAS.n42 161.3
R24515 CS_BIAS.n44 CS_BIAS.n19 161.3
R24516 CS_BIAS.n46 CS_BIAS.n45 161.3
R24517 CS_BIAS.n47 CS_BIAS.n18 161.3
R24518 CS_BIAS.n49 CS_BIAS.n48 161.3
R24519 CS_BIAS.n50 CS_BIAS.n17 161.3
R24520 CS_BIAS.n52 CS_BIAS.n51 161.3
R24521 CS_BIAS.n53 CS_BIAS.n16 161.3
R24522 CS_BIAS.n55 CS_BIAS.n54 161.3
R24523 CS_BIAS.n57 CS_BIAS.n56 161.3
R24524 CS_BIAS.n58 CS_BIAS.n14 161.3
R24525 CS_BIAS.n60 CS_BIAS.n59 161.3
R24526 CS_BIAS.n61 CS_BIAS.n13 161.3
R24527 CS_BIAS.n63 CS_BIAS.n62 161.3
R24528 CS_BIAS.n64 CS_BIAS.n12 161.3
R24529 CS_BIAS.n66 CS_BIAS.n65 161.3
R24530 CS_BIAS.n67 CS_BIAS.n11 161.3
R24531 CS_BIAS.n69 CS_BIAS.n68 161.3
R24532 CS_BIAS.n70 CS_BIAS.n10 161.3
R24533 CS_BIAS.n93 CS_BIAS.n92 161.3
R24534 CS_BIAS.n94 CS_BIAS.n89 161.3
R24535 CS_BIAS.n96 CS_BIAS.n95 161.3
R24536 CS_BIAS.n97 CS_BIAS.n88 161.3
R24537 CS_BIAS.n99 CS_BIAS.n98 161.3
R24538 CS_BIAS.n100 CS_BIAS.n87 161.3
R24539 CS_BIAS.n102 CS_BIAS.n101 161.3
R24540 CS_BIAS.n103 CS_BIAS.n86 161.3
R24541 CS_BIAS.n105 CS_BIAS.n104 161.3
R24542 CS_BIAS.n106 CS_BIAS.n85 161.3
R24543 CS_BIAS.n108 CS_BIAS.n107 161.3
R24544 CS_BIAS.n109 CS_BIAS.n9 161.3
R24545 CS_BIAS.n111 CS_BIAS.n110 161.3
R24546 CS_BIAS.n112 CS_BIAS.n8 161.3
R24547 CS_BIAS.n114 CS_BIAS.n113 161.3
R24548 CS_BIAS.n115 CS_BIAS.n7 161.3
R24549 CS_BIAS.n117 CS_BIAS.n116 161.3
R24550 CS_BIAS.n118 CS_BIAS.n6 161.3
R24551 CS_BIAS.n120 CS_BIAS.n119 161.3
R24552 CS_BIAS.n122 CS_BIAS.n121 161.3
R24553 CS_BIAS.n123 CS_BIAS.n4 161.3
R24554 CS_BIAS.n125 CS_BIAS.n124 161.3
R24555 CS_BIAS.n126 CS_BIAS.n3 161.3
R24556 CS_BIAS.n128 CS_BIAS.n127 161.3
R24557 CS_BIAS.n129 CS_BIAS.n2 161.3
R24558 CS_BIAS.n131 CS_BIAS.n130 161.3
R24559 CS_BIAS.n132 CS_BIAS.n1 161.3
R24560 CS_BIAS.n134 CS_BIAS.n133 161.3
R24561 CS_BIAS.n135 CS_BIAS.n0 161.3
R24562 CS_BIAS.n784 CS_BIAS.n724 161.3
R24563 CS_BIAS.n783 CS_BIAS.n782 161.3
R24564 CS_BIAS.n781 CS_BIAS.n725 161.3
R24565 CS_BIAS.n780 CS_BIAS.n779 161.3
R24566 CS_BIAS.n778 CS_BIAS.n726 161.3
R24567 CS_BIAS.n777 CS_BIAS.n776 161.3
R24568 CS_BIAS.n775 CS_BIAS.n727 161.3
R24569 CS_BIAS.n774 CS_BIAS.n773 161.3
R24570 CS_BIAS.n772 CS_BIAS.n728 161.3
R24571 CS_BIAS.n771 CS_BIAS.n770 161.3
R24572 CS_BIAS.n769 CS_BIAS.n768 161.3
R24573 CS_BIAS.n767 CS_BIAS.n730 161.3
R24574 CS_BIAS.n766 CS_BIAS.n765 161.3
R24575 CS_BIAS.n764 CS_BIAS.n731 161.3
R24576 CS_BIAS.n763 CS_BIAS.n762 161.3
R24577 CS_BIAS.n761 CS_BIAS.n732 161.3
R24578 CS_BIAS.n760 CS_BIAS.n759 161.3
R24579 CS_BIAS.n758 CS_BIAS.n733 161.3
R24580 CS_BIAS.n757 CS_BIAS.n756 161.3
R24581 CS_BIAS.n755 CS_BIAS.n734 161.3
R24582 CS_BIAS.n754 CS_BIAS.n753 161.3
R24583 CS_BIAS.n752 CS_BIAS.n735 161.3
R24584 CS_BIAS.n751 CS_BIAS.n750 161.3
R24585 CS_BIAS.n749 CS_BIAS.n736 161.3
R24586 CS_BIAS.n748 CS_BIAS.n747 161.3
R24587 CS_BIAS.n746 CS_BIAS.n737 161.3
R24588 CS_BIAS.n745 CS_BIAS.n744 161.3
R24589 CS_BIAS.n743 CS_BIAS.n738 161.3
R24590 CS_BIAS.n742 CS_BIAS.n741 161.3
R24591 CS_BIAS.n720 CS_BIAS.n660 161.3
R24592 CS_BIAS.n719 CS_BIAS.n718 161.3
R24593 CS_BIAS.n717 CS_BIAS.n661 161.3
R24594 CS_BIAS.n716 CS_BIAS.n715 161.3
R24595 CS_BIAS.n714 CS_BIAS.n662 161.3
R24596 CS_BIAS.n713 CS_BIAS.n712 161.3
R24597 CS_BIAS.n711 CS_BIAS.n663 161.3
R24598 CS_BIAS.n710 CS_BIAS.n709 161.3
R24599 CS_BIAS.n708 CS_BIAS.n664 161.3
R24600 CS_BIAS.n707 CS_BIAS.n706 161.3
R24601 CS_BIAS.n705 CS_BIAS.n704 161.3
R24602 CS_BIAS.n703 CS_BIAS.n666 161.3
R24603 CS_BIAS.n702 CS_BIAS.n701 161.3
R24604 CS_BIAS.n700 CS_BIAS.n667 161.3
R24605 CS_BIAS.n699 CS_BIAS.n698 161.3
R24606 CS_BIAS.n697 CS_BIAS.n668 161.3
R24607 CS_BIAS.n696 CS_BIAS.n695 161.3
R24608 CS_BIAS.n694 CS_BIAS.n669 161.3
R24609 CS_BIAS.n693 CS_BIAS.n692 161.3
R24610 CS_BIAS.n691 CS_BIAS.n670 161.3
R24611 CS_BIAS.n690 CS_BIAS.n689 161.3
R24612 CS_BIAS.n688 CS_BIAS.n671 161.3
R24613 CS_BIAS.n687 CS_BIAS.n686 161.3
R24614 CS_BIAS.n685 CS_BIAS.n672 161.3
R24615 CS_BIAS.n684 CS_BIAS.n683 161.3
R24616 CS_BIAS.n682 CS_BIAS.n673 161.3
R24617 CS_BIAS.n681 CS_BIAS.n680 161.3
R24618 CS_BIAS.n679 CS_BIAS.n674 161.3
R24619 CS_BIAS.n678 CS_BIAS.n677 161.3
R24620 CS_BIAS.n656 CS_BIAS.n596 161.3
R24621 CS_BIAS.n655 CS_BIAS.n654 161.3
R24622 CS_BIAS.n653 CS_BIAS.n597 161.3
R24623 CS_BIAS.n652 CS_BIAS.n651 161.3
R24624 CS_BIAS.n650 CS_BIAS.n598 161.3
R24625 CS_BIAS.n649 CS_BIAS.n648 161.3
R24626 CS_BIAS.n647 CS_BIAS.n599 161.3
R24627 CS_BIAS.n646 CS_BIAS.n645 161.3
R24628 CS_BIAS.n644 CS_BIAS.n600 161.3
R24629 CS_BIAS.n643 CS_BIAS.n642 161.3
R24630 CS_BIAS.n641 CS_BIAS.n640 161.3
R24631 CS_BIAS.n639 CS_BIAS.n602 161.3
R24632 CS_BIAS.n638 CS_BIAS.n637 161.3
R24633 CS_BIAS.n636 CS_BIAS.n603 161.3
R24634 CS_BIAS.n635 CS_BIAS.n634 161.3
R24635 CS_BIAS.n633 CS_BIAS.n604 161.3
R24636 CS_BIAS.n632 CS_BIAS.n631 161.3
R24637 CS_BIAS.n630 CS_BIAS.n605 161.3
R24638 CS_BIAS.n629 CS_BIAS.n628 161.3
R24639 CS_BIAS.n627 CS_BIAS.n606 161.3
R24640 CS_BIAS.n626 CS_BIAS.n625 161.3
R24641 CS_BIAS.n624 CS_BIAS.n607 161.3
R24642 CS_BIAS.n623 CS_BIAS.n622 161.3
R24643 CS_BIAS.n621 CS_BIAS.n608 161.3
R24644 CS_BIAS.n620 CS_BIAS.n619 161.3
R24645 CS_BIAS.n618 CS_BIAS.n609 161.3
R24646 CS_BIAS.n617 CS_BIAS.n616 161.3
R24647 CS_BIAS.n615 CS_BIAS.n610 161.3
R24648 CS_BIAS.n614 CS_BIAS.n613 161.3
R24649 CS_BIAS.n592 CS_BIAS.n532 161.3
R24650 CS_BIAS.n591 CS_BIAS.n590 161.3
R24651 CS_BIAS.n589 CS_BIAS.n533 161.3
R24652 CS_BIAS.n588 CS_BIAS.n587 161.3
R24653 CS_BIAS.n586 CS_BIAS.n534 161.3
R24654 CS_BIAS.n585 CS_BIAS.n584 161.3
R24655 CS_BIAS.n583 CS_BIAS.n535 161.3
R24656 CS_BIAS.n582 CS_BIAS.n581 161.3
R24657 CS_BIAS.n580 CS_BIAS.n536 161.3
R24658 CS_BIAS.n579 CS_BIAS.n578 161.3
R24659 CS_BIAS.n577 CS_BIAS.n576 161.3
R24660 CS_BIAS.n575 CS_BIAS.n538 161.3
R24661 CS_BIAS.n574 CS_BIAS.n573 161.3
R24662 CS_BIAS.n572 CS_BIAS.n539 161.3
R24663 CS_BIAS.n571 CS_BIAS.n570 161.3
R24664 CS_BIAS.n569 CS_BIAS.n540 161.3
R24665 CS_BIAS.n568 CS_BIAS.n567 161.3
R24666 CS_BIAS.n566 CS_BIAS.n541 161.3
R24667 CS_BIAS.n565 CS_BIAS.n564 161.3
R24668 CS_BIAS.n563 CS_BIAS.n542 161.3
R24669 CS_BIAS.n562 CS_BIAS.n561 161.3
R24670 CS_BIAS.n560 CS_BIAS.n543 161.3
R24671 CS_BIAS.n559 CS_BIAS.n558 161.3
R24672 CS_BIAS.n557 CS_BIAS.n544 161.3
R24673 CS_BIAS.n556 CS_BIAS.n555 161.3
R24674 CS_BIAS.n554 CS_BIAS.n545 161.3
R24675 CS_BIAS.n553 CS_BIAS.n552 161.3
R24676 CS_BIAS.n551 CS_BIAS.n546 161.3
R24677 CS_BIAS.n550 CS_BIAS.n549 161.3
R24678 CS_BIAS.n473 CS_BIAS.n413 161.3
R24679 CS_BIAS.n472 CS_BIAS.n471 161.3
R24680 CS_BIAS.n470 CS_BIAS.n414 161.3
R24681 CS_BIAS.n469 CS_BIAS.n468 161.3
R24682 CS_BIAS.n467 CS_BIAS.n415 161.3
R24683 CS_BIAS.n466 CS_BIAS.n465 161.3
R24684 CS_BIAS.n464 CS_BIAS.n416 161.3
R24685 CS_BIAS.n463 CS_BIAS.n462 161.3
R24686 CS_BIAS.n461 CS_BIAS.n417 161.3
R24687 CS_BIAS.n460 CS_BIAS.n459 161.3
R24688 CS_BIAS.n458 CS_BIAS.n457 161.3
R24689 CS_BIAS.n456 CS_BIAS.n419 161.3
R24690 CS_BIAS.n455 CS_BIAS.n454 161.3
R24691 CS_BIAS.n453 CS_BIAS.n420 161.3
R24692 CS_BIAS.n452 CS_BIAS.n451 161.3
R24693 CS_BIAS.n450 CS_BIAS.n421 161.3
R24694 CS_BIAS.n449 CS_BIAS.n448 161.3
R24695 CS_BIAS.n447 CS_BIAS.n422 161.3
R24696 CS_BIAS.n446 CS_BIAS.n445 161.3
R24697 CS_BIAS.n444 CS_BIAS.n423 161.3
R24698 CS_BIAS.n443 CS_BIAS.n442 161.3
R24699 CS_BIAS.n441 CS_BIAS.n424 161.3
R24700 CS_BIAS.n440 CS_BIAS.n439 161.3
R24701 CS_BIAS.n438 CS_BIAS.n425 161.3
R24702 CS_BIAS.n437 CS_BIAS.n436 161.3
R24703 CS_BIAS.n435 CS_BIAS.n426 161.3
R24704 CS_BIAS.n434 CS_BIAS.n433 161.3
R24705 CS_BIAS.n432 CS_BIAS.n427 161.3
R24706 CS_BIAS.n431 CS_BIAS.n430 161.3
R24707 CS_BIAS.n499 CS_BIAS.n498 161.3
R24708 CS_BIAS.n497 CS_BIAS.n480 161.3
R24709 CS_BIAS.n496 CS_BIAS.n495 161.3
R24710 CS_BIAS.n494 CS_BIAS.n481 161.3
R24711 CS_BIAS.n493 CS_BIAS.n492 161.3
R24712 CS_BIAS.n491 CS_BIAS.n482 161.3
R24713 CS_BIAS.n490 CS_BIAS.n489 161.3
R24714 CS_BIAS.n488 CS_BIAS.n483 161.3
R24715 CS_BIAS.n487 CS_BIAS.n486 161.3
R24716 CS_BIAS.n500 CS_BIAS.n479 161.3
R24717 CS_BIAS.n529 CS_BIAS.n394 161.3
R24718 CS_BIAS.n528 CS_BIAS.n527 161.3
R24719 CS_BIAS.n526 CS_BIAS.n395 161.3
R24720 CS_BIAS.n525 CS_BIAS.n524 161.3
R24721 CS_BIAS.n523 CS_BIAS.n396 161.3
R24722 CS_BIAS.n522 CS_BIAS.n521 161.3
R24723 CS_BIAS.n520 CS_BIAS.n397 161.3
R24724 CS_BIAS.n519 CS_BIAS.n518 161.3
R24725 CS_BIAS.n517 CS_BIAS.n398 161.3
R24726 CS_BIAS.n516 CS_BIAS.n515 161.3
R24727 CS_BIAS.n514 CS_BIAS.n513 161.3
R24728 CS_BIAS.n512 CS_BIAS.n400 161.3
R24729 CS_BIAS.n511 CS_BIAS.n510 161.3
R24730 CS_BIAS.n509 CS_BIAS.n401 161.3
R24731 CS_BIAS.n508 CS_BIAS.n507 161.3
R24732 CS_BIAS.n506 CS_BIAS.n402 161.3
R24733 CS_BIAS.n505 CS_BIAS.n504 161.3
R24734 CS_BIAS.n503 CS_BIAS.n403 161.3
R24735 CS_BIAS.n502 CS_BIAS.n501 161.3
R24736 CS_BIAS.n84 CS_BIAS.n83 119.808
R24737 CS_BIAS.n82 CS_BIAS.n81 118.251
R24738 CS_BIAS.n477 CS_BIAS.n476 118.251
R24739 CS_BIAS.n412 CS_BIAS.n411 118.251
R24740 CS_BIAS.n392 CS_BIAS.n391 75.331
R24741 CS_BIAS.n328 CS_BIAS.n327 75.331
R24742 CS_BIAS.n264 CS_BIAS.n263 75.331
R24743 CS_BIAS.n200 CS_BIAS.n199 75.331
R24744 CS_BIAS.n72 CS_BIAS.n71 75.331
R24745 CS_BIAS.n137 CS_BIAS.n136 75.331
R24746 CS_BIAS.n786 CS_BIAS.n785 75.331
R24747 CS_BIAS.n722 CS_BIAS.n721 75.331
R24748 CS_BIAS.n658 CS_BIAS.n657 75.331
R24749 CS_BIAS.n594 CS_BIAS.n593 75.331
R24750 CS_BIAS.n475 CS_BIAS.n474 75.331
R24751 CS_BIAS.n531 CS_BIAS.n530 75.331
R24752 CS_BIAS.n412 CS_BIAS.n410 67.6205
R24753 CS_BIAS.n80 CS_BIAS.n79 65.5429
R24754 CS_BIAS.n282 CS_BIAS.n281 59.7098
R24755 CS_BIAS.n218 CS_BIAS.n217 59.7098
R24756 CS_BIAS.n154 CS_BIAS.n153 59.7098
R24757 CS_BIAS.n26 CS_BIAS.n25 59.7098
R24758 CS_BIAS.n91 CS_BIAS.n90 59.7098
R24759 CS_BIAS.n346 CS_BIAS.n345 59.7098
R24760 CS_BIAS.n740 CS_BIAS.n739 59.7098
R24761 CS_BIAS.n676 CS_BIAS.n675 59.7098
R24762 CS_BIAS.n612 CS_BIAS.n611 59.7098
R24763 CS_BIAS.n548 CS_BIAS.n547 59.7098
R24764 CS_BIAS.n429 CS_BIAS.n428 59.7098
R24765 CS_BIAS.n485 CS_BIAS.n484 59.7098
R24766 CS_BIAS.n384 CS_BIAS.n383 56.5193
R24767 CS_BIAS.n320 CS_BIAS.n319 56.5193
R24768 CS_BIAS.n256 CS_BIAS.n255 56.5193
R24769 CS_BIAS.n192 CS_BIAS.n191 56.5193
R24770 CS_BIAS.n64 CS_BIAS.n63 56.5193
R24771 CS_BIAS.n129 CS_BIAS.n128 56.5193
R24772 CS_BIAS.n778 CS_BIAS.n777 56.5193
R24773 CS_BIAS.n714 CS_BIAS.n713 56.5193
R24774 CS_BIAS.n650 CS_BIAS.n649 56.5193
R24775 CS_BIAS.n586 CS_BIAS.n585 56.5193
R24776 CS_BIAS.n467 CS_BIAS.n466 56.5193
R24777 CS_BIAS.n523 CS_BIAS.n522 56.5193
R24778 CS_BIAS.n75 CS_BIAS.t1 52.3082
R24779 CS_BIAS.n406 CS_BIAS.t11 52.3082
R24780 CS_BIAS.n355 CS_BIAS.n354 49.2348
R24781 CS_BIAS.n368 CS_BIAS.n367 49.2348
R24782 CS_BIAS.n304 CS_BIAS.n303 49.2348
R24783 CS_BIAS.n291 CS_BIAS.n290 49.2348
R24784 CS_BIAS.n240 CS_BIAS.n239 49.2348
R24785 CS_BIAS.n227 CS_BIAS.n226 49.2348
R24786 CS_BIAS.n176 CS_BIAS.n175 49.2348
R24787 CS_BIAS.n163 CS_BIAS.n162 49.2348
R24788 CS_BIAS.n48 CS_BIAS.n47 49.2348
R24789 CS_BIAS.n35 CS_BIAS.n34 49.2348
R24790 CS_BIAS.n113 CS_BIAS.n112 49.2348
R24791 CS_BIAS.n100 CS_BIAS.n99 49.2348
R24792 CS_BIAS.n749 CS_BIAS.n748 49.2348
R24793 CS_BIAS.n762 CS_BIAS.n761 49.2348
R24794 CS_BIAS.n685 CS_BIAS.n684 49.2348
R24795 CS_BIAS.n698 CS_BIAS.n697 49.2348
R24796 CS_BIAS.n621 CS_BIAS.n620 49.2348
R24797 CS_BIAS.n634 CS_BIAS.n633 49.2348
R24798 CS_BIAS.n557 CS_BIAS.n556 49.2348
R24799 CS_BIAS.n570 CS_BIAS.n569 49.2348
R24800 CS_BIAS.n438 CS_BIAS.n437 49.2348
R24801 CS_BIAS.n451 CS_BIAS.n450 49.2348
R24802 CS_BIAS.n507 CS_BIAS.n506 49.2348
R24803 CS_BIAS.n494 CS_BIAS.n493 49.2348
R24804 CS_BIAS.n346 CS_BIAS.t51 43.9145
R24805 CS_BIAS.n740 CS_BIAS.t44 43.9145
R24806 CS_BIAS.n676 CS_BIAS.t52 43.9145
R24807 CS_BIAS.n612 CS_BIAS.t35 43.9145
R24808 CS_BIAS.n548 CS_BIAS.t65 43.9145
R24809 CS_BIAS.n429 CS_BIAS.t10 43.9145
R24810 CS_BIAS.n485 CS_BIAS.t56 43.9145
R24811 CS_BIAS.n282 CS_BIAS.t59 43.9142
R24812 CS_BIAS.n218 CS_BIAS.t62 43.9142
R24813 CS_BIAS.n154 CS_BIAS.t21 43.9142
R24814 CS_BIAS.n26 CS_BIAS.t4 43.9142
R24815 CS_BIAS.n91 CS_BIAS.t22 43.9142
R24816 CS_BIAS.n354 CS_BIAS.n343 31.752
R24817 CS_BIAS.n368 CS_BIAS.n337 31.752
R24818 CS_BIAS.n304 CS_BIAS.n273 31.752
R24819 CS_BIAS.n290 CS_BIAS.n279 31.752
R24820 CS_BIAS.n240 CS_BIAS.n209 31.752
R24821 CS_BIAS.n226 CS_BIAS.n215 31.752
R24822 CS_BIAS.n176 CS_BIAS.n145 31.752
R24823 CS_BIAS.n162 CS_BIAS.n151 31.752
R24824 CS_BIAS.n48 CS_BIAS.n17 31.752
R24825 CS_BIAS.n34 CS_BIAS.n23 31.752
R24826 CS_BIAS.n113 CS_BIAS.n7 31.752
R24827 CS_BIAS.n99 CS_BIAS.n88 31.752
R24828 CS_BIAS.n748 CS_BIAS.n737 31.752
R24829 CS_BIAS.n762 CS_BIAS.n731 31.752
R24830 CS_BIAS.n684 CS_BIAS.n673 31.752
R24831 CS_BIAS.n698 CS_BIAS.n667 31.752
R24832 CS_BIAS.n620 CS_BIAS.n609 31.752
R24833 CS_BIAS.n634 CS_BIAS.n603 31.752
R24834 CS_BIAS.n556 CS_BIAS.n545 31.752
R24835 CS_BIAS.n570 CS_BIAS.n539 31.752
R24836 CS_BIAS.n437 CS_BIAS.n426 31.752
R24837 CS_BIAS.n451 CS_BIAS.n420 31.752
R24838 CS_BIAS.n507 CS_BIAS.n401 31.752
R24839 CS_BIAS.n493 CS_BIAS.n482 31.752
R24840 CS_BIAS.n350 CS_BIAS.n343 24.4675
R24841 CS_BIAS.n350 CS_BIAS.n349 24.4675
R24842 CS_BIAS.n349 CS_BIAS.n348 24.4675
R24843 CS_BIAS.n367 CS_BIAS.n366 24.4675
R24844 CS_BIAS.n366 CS_BIAS.n339 24.4675
R24845 CS_BIAS.n362 CS_BIAS.n339 24.4675
R24846 CS_BIAS.n362 CS_BIAS.n361 24.4675
R24847 CS_BIAS.n361 CS_BIAS.n360 24.4675
R24848 CS_BIAS.n360 CS_BIAS.n341 24.4675
R24849 CS_BIAS.n356 CS_BIAS.n341 24.4675
R24850 CS_BIAS.n356 CS_BIAS.n355 24.4675
R24851 CS_BIAS.n383 CS_BIAS.n333 24.4675
R24852 CS_BIAS.n379 CS_BIAS.n333 24.4675
R24853 CS_BIAS.n379 CS_BIAS.n378 24.4675
R24854 CS_BIAS.n378 CS_BIAS.n377 24.4675
R24855 CS_BIAS.n374 CS_BIAS.n373 24.4675
R24856 CS_BIAS.n373 CS_BIAS.n372 24.4675
R24857 CS_BIAS.n372 CS_BIAS.n337 24.4675
R24858 CS_BIAS.n390 CS_BIAS.n389 24.4675
R24859 CS_BIAS.n389 CS_BIAS.n331 24.4675
R24860 CS_BIAS.n385 CS_BIAS.n331 24.4675
R24861 CS_BIAS.n385 CS_BIAS.n384 24.4675
R24862 CS_BIAS.n326 CS_BIAS.n325 24.4675
R24863 CS_BIAS.n325 CS_BIAS.n267 24.4675
R24864 CS_BIAS.n321 CS_BIAS.n267 24.4675
R24865 CS_BIAS.n321 CS_BIAS.n320 24.4675
R24866 CS_BIAS.n319 CS_BIAS.n269 24.4675
R24867 CS_BIAS.n315 CS_BIAS.n269 24.4675
R24868 CS_BIAS.n315 CS_BIAS.n314 24.4675
R24869 CS_BIAS.n314 CS_BIAS.n313 24.4675
R24870 CS_BIAS.n310 CS_BIAS.n309 24.4675
R24871 CS_BIAS.n309 CS_BIAS.n308 24.4675
R24872 CS_BIAS.n308 CS_BIAS.n273 24.4675
R24873 CS_BIAS.n303 CS_BIAS.n302 24.4675
R24874 CS_BIAS.n302 CS_BIAS.n275 24.4675
R24875 CS_BIAS.n298 CS_BIAS.n275 24.4675
R24876 CS_BIAS.n298 CS_BIAS.n297 24.4675
R24877 CS_BIAS.n297 CS_BIAS.n296 24.4675
R24878 CS_BIAS.n296 CS_BIAS.n277 24.4675
R24879 CS_BIAS.n292 CS_BIAS.n277 24.4675
R24880 CS_BIAS.n292 CS_BIAS.n291 24.4675
R24881 CS_BIAS.n286 CS_BIAS.n279 24.4675
R24882 CS_BIAS.n286 CS_BIAS.n285 24.4675
R24883 CS_BIAS.n285 CS_BIAS.n284 24.4675
R24884 CS_BIAS.n262 CS_BIAS.n261 24.4675
R24885 CS_BIAS.n261 CS_BIAS.n203 24.4675
R24886 CS_BIAS.n257 CS_BIAS.n203 24.4675
R24887 CS_BIAS.n257 CS_BIAS.n256 24.4675
R24888 CS_BIAS.n255 CS_BIAS.n205 24.4675
R24889 CS_BIAS.n251 CS_BIAS.n205 24.4675
R24890 CS_BIAS.n251 CS_BIAS.n250 24.4675
R24891 CS_BIAS.n250 CS_BIAS.n249 24.4675
R24892 CS_BIAS.n246 CS_BIAS.n245 24.4675
R24893 CS_BIAS.n245 CS_BIAS.n244 24.4675
R24894 CS_BIAS.n244 CS_BIAS.n209 24.4675
R24895 CS_BIAS.n239 CS_BIAS.n238 24.4675
R24896 CS_BIAS.n238 CS_BIAS.n211 24.4675
R24897 CS_BIAS.n234 CS_BIAS.n211 24.4675
R24898 CS_BIAS.n234 CS_BIAS.n233 24.4675
R24899 CS_BIAS.n233 CS_BIAS.n232 24.4675
R24900 CS_BIAS.n232 CS_BIAS.n213 24.4675
R24901 CS_BIAS.n228 CS_BIAS.n213 24.4675
R24902 CS_BIAS.n228 CS_BIAS.n227 24.4675
R24903 CS_BIAS.n222 CS_BIAS.n215 24.4675
R24904 CS_BIAS.n222 CS_BIAS.n221 24.4675
R24905 CS_BIAS.n221 CS_BIAS.n220 24.4675
R24906 CS_BIAS.n198 CS_BIAS.n197 24.4675
R24907 CS_BIAS.n197 CS_BIAS.n139 24.4675
R24908 CS_BIAS.n193 CS_BIAS.n139 24.4675
R24909 CS_BIAS.n193 CS_BIAS.n192 24.4675
R24910 CS_BIAS.n191 CS_BIAS.n141 24.4675
R24911 CS_BIAS.n187 CS_BIAS.n141 24.4675
R24912 CS_BIAS.n187 CS_BIAS.n186 24.4675
R24913 CS_BIAS.n186 CS_BIAS.n185 24.4675
R24914 CS_BIAS.n182 CS_BIAS.n181 24.4675
R24915 CS_BIAS.n181 CS_BIAS.n180 24.4675
R24916 CS_BIAS.n180 CS_BIAS.n145 24.4675
R24917 CS_BIAS.n175 CS_BIAS.n174 24.4675
R24918 CS_BIAS.n174 CS_BIAS.n147 24.4675
R24919 CS_BIAS.n170 CS_BIAS.n147 24.4675
R24920 CS_BIAS.n170 CS_BIAS.n169 24.4675
R24921 CS_BIAS.n169 CS_BIAS.n168 24.4675
R24922 CS_BIAS.n168 CS_BIAS.n149 24.4675
R24923 CS_BIAS.n164 CS_BIAS.n149 24.4675
R24924 CS_BIAS.n164 CS_BIAS.n163 24.4675
R24925 CS_BIAS.n158 CS_BIAS.n151 24.4675
R24926 CS_BIAS.n158 CS_BIAS.n157 24.4675
R24927 CS_BIAS.n157 CS_BIAS.n156 24.4675
R24928 CS_BIAS.n70 CS_BIAS.n69 24.4675
R24929 CS_BIAS.n69 CS_BIAS.n11 24.4675
R24930 CS_BIAS.n65 CS_BIAS.n11 24.4675
R24931 CS_BIAS.n65 CS_BIAS.n64 24.4675
R24932 CS_BIAS.n63 CS_BIAS.n13 24.4675
R24933 CS_BIAS.n59 CS_BIAS.n13 24.4675
R24934 CS_BIAS.n59 CS_BIAS.n58 24.4675
R24935 CS_BIAS.n58 CS_BIAS.n57 24.4675
R24936 CS_BIAS.n54 CS_BIAS.n53 24.4675
R24937 CS_BIAS.n53 CS_BIAS.n52 24.4675
R24938 CS_BIAS.n52 CS_BIAS.n17 24.4675
R24939 CS_BIAS.n47 CS_BIAS.n46 24.4675
R24940 CS_BIAS.n46 CS_BIAS.n19 24.4675
R24941 CS_BIAS.n42 CS_BIAS.n19 24.4675
R24942 CS_BIAS.n42 CS_BIAS.n41 24.4675
R24943 CS_BIAS.n41 CS_BIAS.n40 24.4675
R24944 CS_BIAS.n40 CS_BIAS.n21 24.4675
R24945 CS_BIAS.n36 CS_BIAS.n21 24.4675
R24946 CS_BIAS.n36 CS_BIAS.n35 24.4675
R24947 CS_BIAS.n30 CS_BIAS.n23 24.4675
R24948 CS_BIAS.n30 CS_BIAS.n29 24.4675
R24949 CS_BIAS.n29 CS_BIAS.n28 24.4675
R24950 CS_BIAS.n135 CS_BIAS.n134 24.4675
R24951 CS_BIAS.n134 CS_BIAS.n1 24.4675
R24952 CS_BIAS.n130 CS_BIAS.n1 24.4675
R24953 CS_BIAS.n130 CS_BIAS.n129 24.4675
R24954 CS_BIAS.n128 CS_BIAS.n3 24.4675
R24955 CS_BIAS.n124 CS_BIAS.n3 24.4675
R24956 CS_BIAS.n124 CS_BIAS.n123 24.4675
R24957 CS_BIAS.n123 CS_BIAS.n122 24.4675
R24958 CS_BIAS.n119 CS_BIAS.n118 24.4675
R24959 CS_BIAS.n118 CS_BIAS.n117 24.4675
R24960 CS_BIAS.n117 CS_BIAS.n7 24.4675
R24961 CS_BIAS.n112 CS_BIAS.n111 24.4675
R24962 CS_BIAS.n111 CS_BIAS.n9 24.4675
R24963 CS_BIAS.n107 CS_BIAS.n9 24.4675
R24964 CS_BIAS.n107 CS_BIAS.n106 24.4675
R24965 CS_BIAS.n106 CS_BIAS.n105 24.4675
R24966 CS_BIAS.n105 CS_BIAS.n86 24.4675
R24967 CS_BIAS.n101 CS_BIAS.n86 24.4675
R24968 CS_BIAS.n101 CS_BIAS.n100 24.4675
R24969 CS_BIAS.n95 CS_BIAS.n88 24.4675
R24970 CS_BIAS.n95 CS_BIAS.n94 24.4675
R24971 CS_BIAS.n94 CS_BIAS.n93 24.4675
R24972 CS_BIAS.n743 CS_BIAS.n742 24.4675
R24973 CS_BIAS.n744 CS_BIAS.n743 24.4675
R24974 CS_BIAS.n744 CS_BIAS.n737 24.4675
R24975 CS_BIAS.n750 CS_BIAS.n749 24.4675
R24976 CS_BIAS.n750 CS_BIAS.n735 24.4675
R24977 CS_BIAS.n754 CS_BIAS.n735 24.4675
R24978 CS_BIAS.n755 CS_BIAS.n754 24.4675
R24979 CS_BIAS.n756 CS_BIAS.n755 24.4675
R24980 CS_BIAS.n756 CS_BIAS.n733 24.4675
R24981 CS_BIAS.n760 CS_BIAS.n733 24.4675
R24982 CS_BIAS.n761 CS_BIAS.n760 24.4675
R24983 CS_BIAS.n766 CS_BIAS.n731 24.4675
R24984 CS_BIAS.n767 CS_BIAS.n766 24.4675
R24985 CS_BIAS.n768 CS_BIAS.n767 24.4675
R24986 CS_BIAS.n772 CS_BIAS.n771 24.4675
R24987 CS_BIAS.n773 CS_BIAS.n772 24.4675
R24988 CS_BIAS.n773 CS_BIAS.n727 24.4675
R24989 CS_BIAS.n777 CS_BIAS.n727 24.4675
R24990 CS_BIAS.n779 CS_BIAS.n778 24.4675
R24991 CS_BIAS.n779 CS_BIAS.n725 24.4675
R24992 CS_BIAS.n783 CS_BIAS.n725 24.4675
R24993 CS_BIAS.n784 CS_BIAS.n783 24.4675
R24994 CS_BIAS.n679 CS_BIAS.n678 24.4675
R24995 CS_BIAS.n680 CS_BIAS.n679 24.4675
R24996 CS_BIAS.n680 CS_BIAS.n673 24.4675
R24997 CS_BIAS.n686 CS_BIAS.n685 24.4675
R24998 CS_BIAS.n686 CS_BIAS.n671 24.4675
R24999 CS_BIAS.n690 CS_BIAS.n671 24.4675
R25000 CS_BIAS.n691 CS_BIAS.n690 24.4675
R25001 CS_BIAS.n692 CS_BIAS.n691 24.4675
R25002 CS_BIAS.n692 CS_BIAS.n669 24.4675
R25003 CS_BIAS.n696 CS_BIAS.n669 24.4675
R25004 CS_BIAS.n697 CS_BIAS.n696 24.4675
R25005 CS_BIAS.n702 CS_BIAS.n667 24.4675
R25006 CS_BIAS.n703 CS_BIAS.n702 24.4675
R25007 CS_BIAS.n704 CS_BIAS.n703 24.4675
R25008 CS_BIAS.n708 CS_BIAS.n707 24.4675
R25009 CS_BIAS.n709 CS_BIAS.n708 24.4675
R25010 CS_BIAS.n709 CS_BIAS.n663 24.4675
R25011 CS_BIAS.n713 CS_BIAS.n663 24.4675
R25012 CS_BIAS.n715 CS_BIAS.n714 24.4675
R25013 CS_BIAS.n715 CS_BIAS.n661 24.4675
R25014 CS_BIAS.n719 CS_BIAS.n661 24.4675
R25015 CS_BIAS.n720 CS_BIAS.n719 24.4675
R25016 CS_BIAS.n615 CS_BIAS.n614 24.4675
R25017 CS_BIAS.n616 CS_BIAS.n615 24.4675
R25018 CS_BIAS.n616 CS_BIAS.n609 24.4675
R25019 CS_BIAS.n622 CS_BIAS.n621 24.4675
R25020 CS_BIAS.n622 CS_BIAS.n607 24.4675
R25021 CS_BIAS.n626 CS_BIAS.n607 24.4675
R25022 CS_BIAS.n627 CS_BIAS.n626 24.4675
R25023 CS_BIAS.n628 CS_BIAS.n627 24.4675
R25024 CS_BIAS.n628 CS_BIAS.n605 24.4675
R25025 CS_BIAS.n632 CS_BIAS.n605 24.4675
R25026 CS_BIAS.n633 CS_BIAS.n632 24.4675
R25027 CS_BIAS.n638 CS_BIAS.n603 24.4675
R25028 CS_BIAS.n639 CS_BIAS.n638 24.4675
R25029 CS_BIAS.n640 CS_BIAS.n639 24.4675
R25030 CS_BIAS.n644 CS_BIAS.n643 24.4675
R25031 CS_BIAS.n645 CS_BIAS.n644 24.4675
R25032 CS_BIAS.n645 CS_BIAS.n599 24.4675
R25033 CS_BIAS.n649 CS_BIAS.n599 24.4675
R25034 CS_BIAS.n651 CS_BIAS.n650 24.4675
R25035 CS_BIAS.n651 CS_BIAS.n597 24.4675
R25036 CS_BIAS.n655 CS_BIAS.n597 24.4675
R25037 CS_BIAS.n656 CS_BIAS.n655 24.4675
R25038 CS_BIAS.n551 CS_BIAS.n550 24.4675
R25039 CS_BIAS.n552 CS_BIAS.n551 24.4675
R25040 CS_BIAS.n552 CS_BIAS.n545 24.4675
R25041 CS_BIAS.n558 CS_BIAS.n557 24.4675
R25042 CS_BIAS.n558 CS_BIAS.n543 24.4675
R25043 CS_BIAS.n562 CS_BIAS.n543 24.4675
R25044 CS_BIAS.n563 CS_BIAS.n562 24.4675
R25045 CS_BIAS.n564 CS_BIAS.n563 24.4675
R25046 CS_BIAS.n564 CS_BIAS.n541 24.4675
R25047 CS_BIAS.n568 CS_BIAS.n541 24.4675
R25048 CS_BIAS.n569 CS_BIAS.n568 24.4675
R25049 CS_BIAS.n574 CS_BIAS.n539 24.4675
R25050 CS_BIAS.n575 CS_BIAS.n574 24.4675
R25051 CS_BIAS.n576 CS_BIAS.n575 24.4675
R25052 CS_BIAS.n580 CS_BIAS.n579 24.4675
R25053 CS_BIAS.n581 CS_BIAS.n580 24.4675
R25054 CS_BIAS.n581 CS_BIAS.n535 24.4675
R25055 CS_BIAS.n585 CS_BIAS.n535 24.4675
R25056 CS_BIAS.n587 CS_BIAS.n586 24.4675
R25057 CS_BIAS.n587 CS_BIAS.n533 24.4675
R25058 CS_BIAS.n591 CS_BIAS.n533 24.4675
R25059 CS_BIAS.n592 CS_BIAS.n591 24.4675
R25060 CS_BIAS.n432 CS_BIAS.n431 24.4675
R25061 CS_BIAS.n433 CS_BIAS.n432 24.4675
R25062 CS_BIAS.n433 CS_BIAS.n426 24.4675
R25063 CS_BIAS.n439 CS_BIAS.n438 24.4675
R25064 CS_BIAS.n439 CS_BIAS.n424 24.4675
R25065 CS_BIAS.n443 CS_BIAS.n424 24.4675
R25066 CS_BIAS.n444 CS_BIAS.n443 24.4675
R25067 CS_BIAS.n445 CS_BIAS.n444 24.4675
R25068 CS_BIAS.n445 CS_BIAS.n422 24.4675
R25069 CS_BIAS.n449 CS_BIAS.n422 24.4675
R25070 CS_BIAS.n450 CS_BIAS.n449 24.4675
R25071 CS_BIAS.n455 CS_BIAS.n420 24.4675
R25072 CS_BIAS.n456 CS_BIAS.n455 24.4675
R25073 CS_BIAS.n457 CS_BIAS.n456 24.4675
R25074 CS_BIAS.n461 CS_BIAS.n460 24.4675
R25075 CS_BIAS.n462 CS_BIAS.n461 24.4675
R25076 CS_BIAS.n462 CS_BIAS.n416 24.4675
R25077 CS_BIAS.n466 CS_BIAS.n416 24.4675
R25078 CS_BIAS.n468 CS_BIAS.n467 24.4675
R25079 CS_BIAS.n468 CS_BIAS.n414 24.4675
R25080 CS_BIAS.n472 CS_BIAS.n414 24.4675
R25081 CS_BIAS.n473 CS_BIAS.n472 24.4675
R25082 CS_BIAS.n524 CS_BIAS.n523 24.4675
R25083 CS_BIAS.n524 CS_BIAS.n395 24.4675
R25084 CS_BIAS.n528 CS_BIAS.n395 24.4675
R25085 CS_BIAS.n529 CS_BIAS.n528 24.4675
R25086 CS_BIAS.n511 CS_BIAS.n401 24.4675
R25087 CS_BIAS.n512 CS_BIAS.n511 24.4675
R25088 CS_BIAS.n513 CS_BIAS.n512 24.4675
R25089 CS_BIAS.n517 CS_BIAS.n516 24.4675
R25090 CS_BIAS.n518 CS_BIAS.n517 24.4675
R25091 CS_BIAS.n518 CS_BIAS.n397 24.4675
R25092 CS_BIAS.n522 CS_BIAS.n397 24.4675
R25093 CS_BIAS.n488 CS_BIAS.n487 24.4675
R25094 CS_BIAS.n489 CS_BIAS.n488 24.4675
R25095 CS_BIAS.n489 CS_BIAS.n482 24.4675
R25096 CS_BIAS.n495 CS_BIAS.n494 24.4675
R25097 CS_BIAS.n495 CS_BIAS.n480 24.4675
R25098 CS_BIAS.n499 CS_BIAS.n480 24.4675
R25099 CS_BIAS.n500 CS_BIAS.n499 24.4675
R25100 CS_BIAS.n501 CS_BIAS.n500 24.4675
R25101 CS_BIAS.n501 CS_BIAS.n403 24.4675
R25102 CS_BIAS.n505 CS_BIAS.n403 24.4675
R25103 CS_BIAS.n506 CS_BIAS.n505 24.4675
R25104 CS_BIAS.n348 CS_BIAS.n345 15.6594
R25105 CS_BIAS.n374 CS_BIAS.n335 15.6594
R25106 CS_BIAS.n310 CS_BIAS.n271 15.6594
R25107 CS_BIAS.n284 CS_BIAS.n281 15.6594
R25108 CS_BIAS.n246 CS_BIAS.n207 15.6594
R25109 CS_BIAS.n220 CS_BIAS.n217 15.6594
R25110 CS_BIAS.n182 CS_BIAS.n143 15.6594
R25111 CS_BIAS.n156 CS_BIAS.n153 15.6594
R25112 CS_BIAS.n54 CS_BIAS.n15 15.6594
R25113 CS_BIAS.n28 CS_BIAS.n25 15.6594
R25114 CS_BIAS.n119 CS_BIAS.n5 15.6594
R25115 CS_BIAS.n93 CS_BIAS.n90 15.6594
R25116 CS_BIAS.n742 CS_BIAS.n739 15.6594
R25117 CS_BIAS.n768 CS_BIAS.n729 15.6594
R25118 CS_BIAS.n678 CS_BIAS.n675 15.6594
R25119 CS_BIAS.n704 CS_BIAS.n665 15.6594
R25120 CS_BIAS.n614 CS_BIAS.n611 15.6594
R25121 CS_BIAS.n640 CS_BIAS.n601 15.6594
R25122 CS_BIAS.n550 CS_BIAS.n547 15.6594
R25123 CS_BIAS.n576 CS_BIAS.n537 15.6594
R25124 CS_BIAS.n431 CS_BIAS.n428 15.6594
R25125 CS_BIAS.n457 CS_BIAS.n418 15.6594
R25126 CS_BIAS.n513 CS_BIAS.n399 15.6594
R25127 CS_BIAS.n487 CS_BIAS.n484 15.6594
R25128 CS_BIAS.n477 CS_BIAS.n475 12.3512
R25129 CS_BIAS.n80 CS_BIAS.n72 11.3124
R25130 CS_BIAS.n361 CS_BIAS.t68 10.8965
R25131 CS_BIAS.n345 CS_BIAS.t32 10.8965
R25132 CS_BIAS.n335 CS_BIAS.t48 10.8965
R25133 CS_BIAS.n391 CS_BIAS.t31 10.8965
R25134 CS_BIAS.n297 CS_BIAS.t23 10.8965
R25135 CS_BIAS.n327 CS_BIAS.t36 10.8965
R25136 CS_BIAS.n271 CS_BIAS.t57 10.8965
R25137 CS_BIAS.n281 CS_BIAS.t38 10.8965
R25138 CS_BIAS.n233 CS_BIAS.t26 10.8965
R25139 CS_BIAS.n263 CS_BIAS.t41 10.8965
R25140 CS_BIAS.n207 CS_BIAS.t67 10.8965
R25141 CS_BIAS.n217 CS_BIAS.t49 10.8965
R25142 CS_BIAS.n169 CS_BIAS.t34 10.8965
R25143 CS_BIAS.n199 CS_BIAS.t53 10.8965
R25144 CS_BIAS.n143 CS_BIAS.t20 10.8965
R25145 CS_BIAS.n153 CS_BIAS.t55 10.8965
R25146 CS_BIAS.n41 CS_BIAS.t2 10.8965
R25147 CS_BIAS.n71 CS_BIAS.t0 10.8965
R25148 CS_BIAS.n15 CS_BIAS.t8 10.8965
R25149 CS_BIAS.n25 CS_BIAS.t12 10.8965
R25150 CS_BIAS.n106 CS_BIAS.t24 10.8965
R25151 CS_BIAS.n136 CS_BIAS.t27 10.8965
R25152 CS_BIAS.n5 CS_BIAS.t58 10.8965
R25153 CS_BIAS.n90 CS_BIAS.t47 10.8965
R25154 CS_BIAS.n755 CS_BIAS.t63 10.8965
R25155 CS_BIAS.n739 CS_BIAS.t28 10.8965
R25156 CS_BIAS.n729 CS_BIAS.t43 10.8965
R25157 CS_BIAS.n785 CS_BIAS.t40 10.8965
R25158 CS_BIAS.n691 CS_BIAS.t69 10.8965
R25159 CS_BIAS.n675 CS_BIAS.t33 10.8965
R25160 CS_BIAS.n665 CS_BIAS.t50 10.8965
R25161 CS_BIAS.n721 CS_BIAS.t42 10.8965
R25162 CS_BIAS.n627 CS_BIAS.t54 10.8965
R25163 CS_BIAS.n611 CS_BIAS.t25 10.8965
R25164 CS_BIAS.n601 CS_BIAS.t39 10.8965
R25165 CS_BIAS.n657 CS_BIAS.t66 10.8965
R25166 CS_BIAS.n563 CS_BIAS.t29 10.8965
R25167 CS_BIAS.n547 CS_BIAS.t45 10.8965
R25168 CS_BIAS.n537 CS_BIAS.t64 10.8965
R25169 CS_BIAS.n593 CS_BIAS.t61 10.8965
R25170 CS_BIAS.n444 CS_BIAS.t6 10.8965
R25171 CS_BIAS.n428 CS_BIAS.t18 10.8965
R25172 CS_BIAS.n418 CS_BIAS.t16 10.8965
R25173 CS_BIAS.n474 CS_BIAS.t14 10.8965
R25174 CS_BIAS.n500 CS_BIAS.t60 10.8965
R25175 CS_BIAS.n530 CS_BIAS.t46 10.8965
R25176 CS_BIAS.n399 CS_BIAS.t37 10.8965
R25177 CS_BIAS.n484 CS_BIAS.t30 10.8965
R25178 CS_BIAS.n788 CS_BIAS.n393 10.4074
R25179 CS_BIAS.n83 CS_BIAS.t13 9.75419
R25180 CS_BIAS.n83 CS_BIAS.t5 9.75419
R25181 CS_BIAS.n81 CS_BIAS.t9 9.75419
R25182 CS_BIAS.n81 CS_BIAS.t3 9.75419
R25183 CS_BIAS.n476 CS_BIAS.t17 9.75419
R25184 CS_BIAS.n476 CS_BIAS.t15 9.75419
R25185 CS_BIAS.n411 CS_BIAS.t19 9.75419
R25186 CS_BIAS.n411 CS_BIAS.t7 9.75419
R25187 CS_BIAS.n76 CS_BIAS.n74 9.71174
R25188 CS_BIAS.n407 CS_BIAS.n405 9.71174
R25189 CS_BIAS.n85 CS_BIAS.n84 9.50363
R25190 CS_BIAS.n479 CS_BIAS.n478 9.50363
R25191 CS_BIAS.n79 CS_BIAS.n78 9.45567
R25192 CS_BIAS.n410 CS_BIAS.n409 9.45567
R25193 CS_BIAS.n78 CS_BIAS.n77 9.3005
R25194 CS_BIAS.n409 CS_BIAS.n408 9.3005
R25195 CS_BIAS.n377 CS_BIAS.n335 8.80862
R25196 CS_BIAS.n313 CS_BIAS.n271 8.80862
R25197 CS_BIAS.n249 CS_BIAS.n207 8.80862
R25198 CS_BIAS.n185 CS_BIAS.n143 8.80862
R25199 CS_BIAS.n57 CS_BIAS.n15 8.80862
R25200 CS_BIAS.n122 CS_BIAS.n5 8.80862
R25201 CS_BIAS.n771 CS_BIAS.n729 8.80862
R25202 CS_BIAS.n707 CS_BIAS.n665 8.80862
R25203 CS_BIAS.n643 CS_BIAS.n601 8.80862
R25204 CS_BIAS.n579 CS_BIAS.n537 8.80862
R25205 CS_BIAS.n460 CS_BIAS.n418 8.80862
R25206 CS_BIAS.n516 CS_BIAS.n399 8.80862
R25207 CS_BIAS.n79 CS_BIAS.n73 8.14595
R25208 CS_BIAS.n410 CS_BIAS.n404 8.14595
R25209 CS_BIAS.n77 CS_BIAS.n76 7.3702
R25210 CS_BIAS.n408 CS_BIAS.n407 7.3702
R25211 CS_BIAS.n201 CS_BIAS.n137 7.08937
R25212 CS_BIAS.n595 CS_BIAS.n531 7.08937
R25213 CS_BIAS.n391 CS_BIAS.n390 6.85126
R25214 CS_BIAS.n327 CS_BIAS.n326 6.85126
R25215 CS_BIAS.n263 CS_BIAS.n262 6.85126
R25216 CS_BIAS.n199 CS_BIAS.n198 6.85126
R25217 CS_BIAS.n71 CS_BIAS.n70 6.85126
R25218 CS_BIAS.n136 CS_BIAS.n135 6.85126
R25219 CS_BIAS.n785 CS_BIAS.n784 6.85126
R25220 CS_BIAS.n721 CS_BIAS.n720 6.85126
R25221 CS_BIAS.n657 CS_BIAS.n656 6.85126
R25222 CS_BIAS.n593 CS_BIAS.n592 6.85126
R25223 CS_BIAS.n474 CS_BIAS.n473 6.85126
R25224 CS_BIAS.n530 CS_BIAS.n529 6.85126
R25225 CS_BIAS.n788 CS_BIAS.n787 6.71164
R25226 CS_BIAS.n77 CS_BIAS.n73 5.81868
R25227 CS_BIAS.n408 CS_BIAS.n404 5.81868
R25228 CS_BIAS.n393 CS_BIAS.n392 5.27876
R25229 CS_BIAS.n329 CS_BIAS.n328 5.27876
R25230 CS_BIAS.n265 CS_BIAS.n264 5.27876
R25231 CS_BIAS.n201 CS_BIAS.n200 5.27876
R25232 CS_BIAS.n787 CS_BIAS.n786 5.27876
R25233 CS_BIAS.n723 CS_BIAS.n722 5.27876
R25234 CS_BIAS.n659 CS_BIAS.n658 5.27876
R25235 CS_BIAS.n595 CS_BIAS.n594 5.27876
R25236 CS_BIAS CS_BIAS.n788 4.04825
R25237 CS_BIAS.n78 CS_BIAS.n74 3.44771
R25238 CS_BIAS.n409 CS_BIAS.n405 3.44771
R25239 CS_BIAS.n82 CS_BIAS.n80 2.07809
R25240 CS_BIAS.n265 CS_BIAS.n201 1.81111
R25241 CS_BIAS.n329 CS_BIAS.n265 1.81111
R25242 CS_BIAS.n393 CS_BIAS.n329 1.81111
R25243 CS_BIAS.n659 CS_BIAS.n595 1.81111
R25244 CS_BIAS.n723 CS_BIAS.n659 1.81111
R25245 CS_BIAS.n787 CS_BIAS.n723 1.81111
R25246 CS_BIAS.n347 CS_BIAS.n346 1.75081
R25247 CS_BIAS.n741 CS_BIAS.n740 1.75081
R25248 CS_BIAS.n677 CS_BIAS.n676 1.75081
R25249 CS_BIAS.n613 CS_BIAS.n612 1.75081
R25250 CS_BIAS.n549 CS_BIAS.n548 1.75081
R25251 CS_BIAS.n430 CS_BIAS.n429 1.75081
R25252 CS_BIAS.n486 CS_BIAS.n485 1.75081
R25253 CS_BIAS.n283 CS_BIAS.n282 1.7508
R25254 CS_BIAS.n219 CS_BIAS.n218 1.7508
R25255 CS_BIAS.n155 CS_BIAS.n154 1.7508
R25256 CS_BIAS.n27 CS_BIAS.n26 1.7508
R25257 CS_BIAS.n92 CS_BIAS.n91 1.7508
R25258 CS_BIAS.n478 CS_BIAS.n477 1.55869
R25259 CS_BIAS.n84 CS_BIAS.n82 0.519897
R25260 CS_BIAS.n478 CS_BIAS.n412 0.519897
R25261 CS_BIAS.n392 CS_BIAS.n330 0.417535
R25262 CS_BIAS.n328 CS_BIAS.n266 0.417535
R25263 CS_BIAS.n264 CS_BIAS.n202 0.417535
R25264 CS_BIAS.n200 CS_BIAS.n138 0.417535
R25265 CS_BIAS.n72 CS_BIAS.n10 0.417535
R25266 CS_BIAS.n137 CS_BIAS.n0 0.417535
R25267 CS_BIAS.n786 CS_BIAS.n724 0.417535
R25268 CS_BIAS.n722 CS_BIAS.n660 0.417535
R25269 CS_BIAS.n658 CS_BIAS.n596 0.417535
R25270 CS_BIAS.n594 CS_BIAS.n532 0.417535
R25271 CS_BIAS.n475 CS_BIAS.n413 0.417535
R25272 CS_BIAS.n531 CS_BIAS.n394 0.417535
R25273 CS_BIAS.n388 CS_BIAS.n330 0.189894
R25274 CS_BIAS.n388 CS_BIAS.n387 0.189894
R25275 CS_BIAS.n387 CS_BIAS.n386 0.189894
R25276 CS_BIAS.n386 CS_BIAS.n332 0.189894
R25277 CS_BIAS.n382 CS_BIAS.n332 0.189894
R25278 CS_BIAS.n382 CS_BIAS.n381 0.189894
R25279 CS_BIAS.n381 CS_BIAS.n380 0.189894
R25280 CS_BIAS.n380 CS_BIAS.n334 0.189894
R25281 CS_BIAS.n376 CS_BIAS.n334 0.189894
R25282 CS_BIAS.n376 CS_BIAS.n375 0.189894
R25283 CS_BIAS.n375 CS_BIAS.n336 0.189894
R25284 CS_BIAS.n371 CS_BIAS.n336 0.189894
R25285 CS_BIAS.n371 CS_BIAS.n370 0.189894
R25286 CS_BIAS.n370 CS_BIAS.n369 0.189894
R25287 CS_BIAS.n369 CS_BIAS.n338 0.189894
R25288 CS_BIAS.n365 CS_BIAS.n338 0.189894
R25289 CS_BIAS.n365 CS_BIAS.n364 0.189894
R25290 CS_BIAS.n364 CS_BIAS.n363 0.189894
R25291 CS_BIAS.n363 CS_BIAS.n340 0.189894
R25292 CS_BIAS.n359 CS_BIAS.n340 0.189894
R25293 CS_BIAS.n359 CS_BIAS.n358 0.189894
R25294 CS_BIAS.n358 CS_BIAS.n357 0.189894
R25295 CS_BIAS.n357 CS_BIAS.n342 0.189894
R25296 CS_BIAS.n353 CS_BIAS.n342 0.189894
R25297 CS_BIAS.n353 CS_BIAS.n352 0.189894
R25298 CS_BIAS.n352 CS_BIAS.n351 0.189894
R25299 CS_BIAS.n351 CS_BIAS.n344 0.189894
R25300 CS_BIAS.n347 CS_BIAS.n344 0.189894
R25301 CS_BIAS.n324 CS_BIAS.n266 0.189894
R25302 CS_BIAS.n324 CS_BIAS.n323 0.189894
R25303 CS_BIAS.n323 CS_BIAS.n322 0.189894
R25304 CS_BIAS.n322 CS_BIAS.n268 0.189894
R25305 CS_BIAS.n318 CS_BIAS.n268 0.189894
R25306 CS_BIAS.n318 CS_BIAS.n317 0.189894
R25307 CS_BIAS.n317 CS_BIAS.n316 0.189894
R25308 CS_BIAS.n316 CS_BIAS.n270 0.189894
R25309 CS_BIAS.n312 CS_BIAS.n270 0.189894
R25310 CS_BIAS.n312 CS_BIAS.n311 0.189894
R25311 CS_BIAS.n311 CS_BIAS.n272 0.189894
R25312 CS_BIAS.n307 CS_BIAS.n272 0.189894
R25313 CS_BIAS.n307 CS_BIAS.n306 0.189894
R25314 CS_BIAS.n306 CS_BIAS.n305 0.189894
R25315 CS_BIAS.n305 CS_BIAS.n274 0.189894
R25316 CS_BIAS.n301 CS_BIAS.n274 0.189894
R25317 CS_BIAS.n301 CS_BIAS.n300 0.189894
R25318 CS_BIAS.n300 CS_BIAS.n299 0.189894
R25319 CS_BIAS.n299 CS_BIAS.n276 0.189894
R25320 CS_BIAS.n295 CS_BIAS.n276 0.189894
R25321 CS_BIAS.n295 CS_BIAS.n294 0.189894
R25322 CS_BIAS.n294 CS_BIAS.n293 0.189894
R25323 CS_BIAS.n293 CS_BIAS.n278 0.189894
R25324 CS_BIAS.n289 CS_BIAS.n278 0.189894
R25325 CS_BIAS.n289 CS_BIAS.n288 0.189894
R25326 CS_BIAS.n288 CS_BIAS.n287 0.189894
R25327 CS_BIAS.n287 CS_BIAS.n280 0.189894
R25328 CS_BIAS.n283 CS_BIAS.n280 0.189894
R25329 CS_BIAS.n260 CS_BIAS.n202 0.189894
R25330 CS_BIAS.n260 CS_BIAS.n259 0.189894
R25331 CS_BIAS.n259 CS_BIAS.n258 0.189894
R25332 CS_BIAS.n258 CS_BIAS.n204 0.189894
R25333 CS_BIAS.n254 CS_BIAS.n204 0.189894
R25334 CS_BIAS.n254 CS_BIAS.n253 0.189894
R25335 CS_BIAS.n253 CS_BIAS.n252 0.189894
R25336 CS_BIAS.n252 CS_BIAS.n206 0.189894
R25337 CS_BIAS.n248 CS_BIAS.n206 0.189894
R25338 CS_BIAS.n248 CS_BIAS.n247 0.189894
R25339 CS_BIAS.n247 CS_BIAS.n208 0.189894
R25340 CS_BIAS.n243 CS_BIAS.n208 0.189894
R25341 CS_BIAS.n243 CS_BIAS.n242 0.189894
R25342 CS_BIAS.n242 CS_BIAS.n241 0.189894
R25343 CS_BIAS.n241 CS_BIAS.n210 0.189894
R25344 CS_BIAS.n237 CS_BIAS.n210 0.189894
R25345 CS_BIAS.n237 CS_BIAS.n236 0.189894
R25346 CS_BIAS.n236 CS_BIAS.n235 0.189894
R25347 CS_BIAS.n235 CS_BIAS.n212 0.189894
R25348 CS_BIAS.n231 CS_BIAS.n212 0.189894
R25349 CS_BIAS.n231 CS_BIAS.n230 0.189894
R25350 CS_BIAS.n230 CS_BIAS.n229 0.189894
R25351 CS_BIAS.n229 CS_BIAS.n214 0.189894
R25352 CS_BIAS.n225 CS_BIAS.n214 0.189894
R25353 CS_BIAS.n225 CS_BIAS.n224 0.189894
R25354 CS_BIAS.n224 CS_BIAS.n223 0.189894
R25355 CS_BIAS.n223 CS_BIAS.n216 0.189894
R25356 CS_BIAS.n219 CS_BIAS.n216 0.189894
R25357 CS_BIAS.n196 CS_BIAS.n138 0.189894
R25358 CS_BIAS.n196 CS_BIAS.n195 0.189894
R25359 CS_BIAS.n195 CS_BIAS.n194 0.189894
R25360 CS_BIAS.n194 CS_BIAS.n140 0.189894
R25361 CS_BIAS.n190 CS_BIAS.n140 0.189894
R25362 CS_BIAS.n190 CS_BIAS.n189 0.189894
R25363 CS_BIAS.n189 CS_BIAS.n188 0.189894
R25364 CS_BIAS.n188 CS_BIAS.n142 0.189894
R25365 CS_BIAS.n184 CS_BIAS.n142 0.189894
R25366 CS_BIAS.n184 CS_BIAS.n183 0.189894
R25367 CS_BIAS.n183 CS_BIAS.n144 0.189894
R25368 CS_BIAS.n179 CS_BIAS.n144 0.189894
R25369 CS_BIAS.n179 CS_BIAS.n178 0.189894
R25370 CS_BIAS.n178 CS_BIAS.n177 0.189894
R25371 CS_BIAS.n177 CS_BIAS.n146 0.189894
R25372 CS_BIAS.n173 CS_BIAS.n146 0.189894
R25373 CS_BIAS.n173 CS_BIAS.n172 0.189894
R25374 CS_BIAS.n172 CS_BIAS.n171 0.189894
R25375 CS_BIAS.n171 CS_BIAS.n148 0.189894
R25376 CS_BIAS.n167 CS_BIAS.n148 0.189894
R25377 CS_BIAS.n167 CS_BIAS.n166 0.189894
R25378 CS_BIAS.n166 CS_BIAS.n165 0.189894
R25379 CS_BIAS.n165 CS_BIAS.n150 0.189894
R25380 CS_BIAS.n161 CS_BIAS.n150 0.189894
R25381 CS_BIAS.n161 CS_BIAS.n160 0.189894
R25382 CS_BIAS.n160 CS_BIAS.n159 0.189894
R25383 CS_BIAS.n159 CS_BIAS.n152 0.189894
R25384 CS_BIAS.n155 CS_BIAS.n152 0.189894
R25385 CS_BIAS.n68 CS_BIAS.n10 0.189894
R25386 CS_BIAS.n68 CS_BIAS.n67 0.189894
R25387 CS_BIAS.n67 CS_BIAS.n66 0.189894
R25388 CS_BIAS.n66 CS_BIAS.n12 0.189894
R25389 CS_BIAS.n62 CS_BIAS.n12 0.189894
R25390 CS_BIAS.n62 CS_BIAS.n61 0.189894
R25391 CS_BIAS.n61 CS_BIAS.n60 0.189894
R25392 CS_BIAS.n60 CS_BIAS.n14 0.189894
R25393 CS_BIAS.n56 CS_BIAS.n14 0.189894
R25394 CS_BIAS.n56 CS_BIAS.n55 0.189894
R25395 CS_BIAS.n55 CS_BIAS.n16 0.189894
R25396 CS_BIAS.n51 CS_BIAS.n16 0.189894
R25397 CS_BIAS.n51 CS_BIAS.n50 0.189894
R25398 CS_BIAS.n50 CS_BIAS.n49 0.189894
R25399 CS_BIAS.n49 CS_BIAS.n18 0.189894
R25400 CS_BIAS.n45 CS_BIAS.n18 0.189894
R25401 CS_BIAS.n45 CS_BIAS.n44 0.189894
R25402 CS_BIAS.n44 CS_BIAS.n43 0.189894
R25403 CS_BIAS.n43 CS_BIAS.n20 0.189894
R25404 CS_BIAS.n39 CS_BIAS.n20 0.189894
R25405 CS_BIAS.n39 CS_BIAS.n38 0.189894
R25406 CS_BIAS.n38 CS_BIAS.n37 0.189894
R25407 CS_BIAS.n37 CS_BIAS.n22 0.189894
R25408 CS_BIAS.n33 CS_BIAS.n22 0.189894
R25409 CS_BIAS.n33 CS_BIAS.n32 0.189894
R25410 CS_BIAS.n32 CS_BIAS.n31 0.189894
R25411 CS_BIAS.n31 CS_BIAS.n24 0.189894
R25412 CS_BIAS.n27 CS_BIAS.n24 0.189894
R25413 CS_BIAS.n104 CS_BIAS.n103 0.189894
R25414 CS_BIAS.n103 CS_BIAS.n102 0.189894
R25415 CS_BIAS.n102 CS_BIAS.n87 0.189894
R25416 CS_BIAS.n98 CS_BIAS.n87 0.189894
R25417 CS_BIAS.n98 CS_BIAS.n97 0.189894
R25418 CS_BIAS.n97 CS_BIAS.n96 0.189894
R25419 CS_BIAS.n96 CS_BIAS.n89 0.189894
R25420 CS_BIAS.n92 CS_BIAS.n89 0.189894
R25421 CS_BIAS.n133 CS_BIAS.n0 0.189894
R25422 CS_BIAS.n133 CS_BIAS.n132 0.189894
R25423 CS_BIAS.n132 CS_BIAS.n131 0.189894
R25424 CS_BIAS.n131 CS_BIAS.n2 0.189894
R25425 CS_BIAS.n127 CS_BIAS.n2 0.189894
R25426 CS_BIAS.n127 CS_BIAS.n126 0.189894
R25427 CS_BIAS.n126 CS_BIAS.n125 0.189894
R25428 CS_BIAS.n125 CS_BIAS.n4 0.189894
R25429 CS_BIAS.n121 CS_BIAS.n4 0.189894
R25430 CS_BIAS.n121 CS_BIAS.n120 0.189894
R25431 CS_BIAS.n120 CS_BIAS.n6 0.189894
R25432 CS_BIAS.n116 CS_BIAS.n6 0.189894
R25433 CS_BIAS.n116 CS_BIAS.n115 0.189894
R25434 CS_BIAS.n115 CS_BIAS.n114 0.189894
R25435 CS_BIAS.n114 CS_BIAS.n8 0.189894
R25436 CS_BIAS.n110 CS_BIAS.n8 0.189894
R25437 CS_BIAS.n110 CS_BIAS.n109 0.189894
R25438 CS_BIAS.n109 CS_BIAS.n108 0.189894
R25439 CS_BIAS.n741 CS_BIAS.n738 0.189894
R25440 CS_BIAS.n745 CS_BIAS.n738 0.189894
R25441 CS_BIAS.n746 CS_BIAS.n745 0.189894
R25442 CS_BIAS.n747 CS_BIAS.n746 0.189894
R25443 CS_BIAS.n747 CS_BIAS.n736 0.189894
R25444 CS_BIAS.n751 CS_BIAS.n736 0.189894
R25445 CS_BIAS.n752 CS_BIAS.n751 0.189894
R25446 CS_BIAS.n753 CS_BIAS.n752 0.189894
R25447 CS_BIAS.n753 CS_BIAS.n734 0.189894
R25448 CS_BIAS.n757 CS_BIAS.n734 0.189894
R25449 CS_BIAS.n758 CS_BIAS.n757 0.189894
R25450 CS_BIAS.n759 CS_BIAS.n758 0.189894
R25451 CS_BIAS.n759 CS_BIAS.n732 0.189894
R25452 CS_BIAS.n763 CS_BIAS.n732 0.189894
R25453 CS_BIAS.n764 CS_BIAS.n763 0.189894
R25454 CS_BIAS.n765 CS_BIAS.n764 0.189894
R25455 CS_BIAS.n765 CS_BIAS.n730 0.189894
R25456 CS_BIAS.n769 CS_BIAS.n730 0.189894
R25457 CS_BIAS.n770 CS_BIAS.n769 0.189894
R25458 CS_BIAS.n770 CS_BIAS.n728 0.189894
R25459 CS_BIAS.n774 CS_BIAS.n728 0.189894
R25460 CS_BIAS.n775 CS_BIAS.n774 0.189894
R25461 CS_BIAS.n776 CS_BIAS.n775 0.189894
R25462 CS_BIAS.n776 CS_BIAS.n726 0.189894
R25463 CS_BIAS.n780 CS_BIAS.n726 0.189894
R25464 CS_BIAS.n781 CS_BIAS.n780 0.189894
R25465 CS_BIAS.n782 CS_BIAS.n781 0.189894
R25466 CS_BIAS.n782 CS_BIAS.n724 0.189894
R25467 CS_BIAS.n677 CS_BIAS.n674 0.189894
R25468 CS_BIAS.n681 CS_BIAS.n674 0.189894
R25469 CS_BIAS.n682 CS_BIAS.n681 0.189894
R25470 CS_BIAS.n683 CS_BIAS.n682 0.189894
R25471 CS_BIAS.n683 CS_BIAS.n672 0.189894
R25472 CS_BIAS.n687 CS_BIAS.n672 0.189894
R25473 CS_BIAS.n688 CS_BIAS.n687 0.189894
R25474 CS_BIAS.n689 CS_BIAS.n688 0.189894
R25475 CS_BIAS.n689 CS_BIAS.n670 0.189894
R25476 CS_BIAS.n693 CS_BIAS.n670 0.189894
R25477 CS_BIAS.n694 CS_BIAS.n693 0.189894
R25478 CS_BIAS.n695 CS_BIAS.n694 0.189894
R25479 CS_BIAS.n695 CS_BIAS.n668 0.189894
R25480 CS_BIAS.n699 CS_BIAS.n668 0.189894
R25481 CS_BIAS.n700 CS_BIAS.n699 0.189894
R25482 CS_BIAS.n701 CS_BIAS.n700 0.189894
R25483 CS_BIAS.n701 CS_BIAS.n666 0.189894
R25484 CS_BIAS.n705 CS_BIAS.n666 0.189894
R25485 CS_BIAS.n706 CS_BIAS.n705 0.189894
R25486 CS_BIAS.n706 CS_BIAS.n664 0.189894
R25487 CS_BIAS.n710 CS_BIAS.n664 0.189894
R25488 CS_BIAS.n711 CS_BIAS.n710 0.189894
R25489 CS_BIAS.n712 CS_BIAS.n711 0.189894
R25490 CS_BIAS.n712 CS_BIAS.n662 0.189894
R25491 CS_BIAS.n716 CS_BIAS.n662 0.189894
R25492 CS_BIAS.n717 CS_BIAS.n716 0.189894
R25493 CS_BIAS.n718 CS_BIAS.n717 0.189894
R25494 CS_BIAS.n718 CS_BIAS.n660 0.189894
R25495 CS_BIAS.n613 CS_BIAS.n610 0.189894
R25496 CS_BIAS.n617 CS_BIAS.n610 0.189894
R25497 CS_BIAS.n618 CS_BIAS.n617 0.189894
R25498 CS_BIAS.n619 CS_BIAS.n618 0.189894
R25499 CS_BIAS.n619 CS_BIAS.n608 0.189894
R25500 CS_BIAS.n623 CS_BIAS.n608 0.189894
R25501 CS_BIAS.n624 CS_BIAS.n623 0.189894
R25502 CS_BIAS.n625 CS_BIAS.n624 0.189894
R25503 CS_BIAS.n625 CS_BIAS.n606 0.189894
R25504 CS_BIAS.n629 CS_BIAS.n606 0.189894
R25505 CS_BIAS.n630 CS_BIAS.n629 0.189894
R25506 CS_BIAS.n631 CS_BIAS.n630 0.189894
R25507 CS_BIAS.n631 CS_BIAS.n604 0.189894
R25508 CS_BIAS.n635 CS_BIAS.n604 0.189894
R25509 CS_BIAS.n636 CS_BIAS.n635 0.189894
R25510 CS_BIAS.n637 CS_BIAS.n636 0.189894
R25511 CS_BIAS.n637 CS_BIAS.n602 0.189894
R25512 CS_BIAS.n641 CS_BIAS.n602 0.189894
R25513 CS_BIAS.n642 CS_BIAS.n641 0.189894
R25514 CS_BIAS.n642 CS_BIAS.n600 0.189894
R25515 CS_BIAS.n646 CS_BIAS.n600 0.189894
R25516 CS_BIAS.n647 CS_BIAS.n646 0.189894
R25517 CS_BIAS.n648 CS_BIAS.n647 0.189894
R25518 CS_BIAS.n648 CS_BIAS.n598 0.189894
R25519 CS_BIAS.n652 CS_BIAS.n598 0.189894
R25520 CS_BIAS.n653 CS_BIAS.n652 0.189894
R25521 CS_BIAS.n654 CS_BIAS.n653 0.189894
R25522 CS_BIAS.n654 CS_BIAS.n596 0.189894
R25523 CS_BIAS.n549 CS_BIAS.n546 0.189894
R25524 CS_BIAS.n553 CS_BIAS.n546 0.189894
R25525 CS_BIAS.n554 CS_BIAS.n553 0.189894
R25526 CS_BIAS.n555 CS_BIAS.n554 0.189894
R25527 CS_BIAS.n555 CS_BIAS.n544 0.189894
R25528 CS_BIAS.n559 CS_BIAS.n544 0.189894
R25529 CS_BIAS.n560 CS_BIAS.n559 0.189894
R25530 CS_BIAS.n561 CS_BIAS.n560 0.189894
R25531 CS_BIAS.n561 CS_BIAS.n542 0.189894
R25532 CS_BIAS.n565 CS_BIAS.n542 0.189894
R25533 CS_BIAS.n566 CS_BIAS.n565 0.189894
R25534 CS_BIAS.n567 CS_BIAS.n566 0.189894
R25535 CS_BIAS.n567 CS_BIAS.n540 0.189894
R25536 CS_BIAS.n571 CS_BIAS.n540 0.189894
R25537 CS_BIAS.n572 CS_BIAS.n571 0.189894
R25538 CS_BIAS.n573 CS_BIAS.n572 0.189894
R25539 CS_BIAS.n573 CS_BIAS.n538 0.189894
R25540 CS_BIAS.n577 CS_BIAS.n538 0.189894
R25541 CS_BIAS.n578 CS_BIAS.n577 0.189894
R25542 CS_BIAS.n578 CS_BIAS.n536 0.189894
R25543 CS_BIAS.n582 CS_BIAS.n536 0.189894
R25544 CS_BIAS.n583 CS_BIAS.n582 0.189894
R25545 CS_BIAS.n584 CS_BIAS.n583 0.189894
R25546 CS_BIAS.n584 CS_BIAS.n534 0.189894
R25547 CS_BIAS.n588 CS_BIAS.n534 0.189894
R25548 CS_BIAS.n589 CS_BIAS.n588 0.189894
R25549 CS_BIAS.n590 CS_BIAS.n589 0.189894
R25550 CS_BIAS.n590 CS_BIAS.n532 0.189894
R25551 CS_BIAS.n430 CS_BIAS.n427 0.189894
R25552 CS_BIAS.n434 CS_BIAS.n427 0.189894
R25553 CS_BIAS.n435 CS_BIAS.n434 0.189894
R25554 CS_BIAS.n436 CS_BIAS.n435 0.189894
R25555 CS_BIAS.n436 CS_BIAS.n425 0.189894
R25556 CS_BIAS.n440 CS_BIAS.n425 0.189894
R25557 CS_BIAS.n441 CS_BIAS.n440 0.189894
R25558 CS_BIAS.n442 CS_BIAS.n441 0.189894
R25559 CS_BIAS.n442 CS_BIAS.n423 0.189894
R25560 CS_BIAS.n446 CS_BIAS.n423 0.189894
R25561 CS_BIAS.n447 CS_BIAS.n446 0.189894
R25562 CS_BIAS.n448 CS_BIAS.n447 0.189894
R25563 CS_BIAS.n448 CS_BIAS.n421 0.189894
R25564 CS_BIAS.n452 CS_BIAS.n421 0.189894
R25565 CS_BIAS.n453 CS_BIAS.n452 0.189894
R25566 CS_BIAS.n454 CS_BIAS.n453 0.189894
R25567 CS_BIAS.n454 CS_BIAS.n419 0.189894
R25568 CS_BIAS.n458 CS_BIAS.n419 0.189894
R25569 CS_BIAS.n459 CS_BIAS.n458 0.189894
R25570 CS_BIAS.n459 CS_BIAS.n417 0.189894
R25571 CS_BIAS.n463 CS_BIAS.n417 0.189894
R25572 CS_BIAS.n464 CS_BIAS.n463 0.189894
R25573 CS_BIAS.n465 CS_BIAS.n464 0.189894
R25574 CS_BIAS.n465 CS_BIAS.n415 0.189894
R25575 CS_BIAS.n469 CS_BIAS.n415 0.189894
R25576 CS_BIAS.n470 CS_BIAS.n469 0.189894
R25577 CS_BIAS.n471 CS_BIAS.n470 0.189894
R25578 CS_BIAS.n471 CS_BIAS.n413 0.189894
R25579 CS_BIAS.n486 CS_BIAS.n483 0.189894
R25580 CS_BIAS.n490 CS_BIAS.n483 0.189894
R25581 CS_BIAS.n491 CS_BIAS.n490 0.189894
R25582 CS_BIAS.n492 CS_BIAS.n491 0.189894
R25583 CS_BIAS.n492 CS_BIAS.n481 0.189894
R25584 CS_BIAS.n496 CS_BIAS.n481 0.189894
R25585 CS_BIAS.n497 CS_BIAS.n496 0.189894
R25586 CS_BIAS.n498 CS_BIAS.n497 0.189894
R25587 CS_BIAS.n503 CS_BIAS.n502 0.189894
R25588 CS_BIAS.n504 CS_BIAS.n503 0.189894
R25589 CS_BIAS.n504 CS_BIAS.n402 0.189894
R25590 CS_BIAS.n508 CS_BIAS.n402 0.189894
R25591 CS_BIAS.n509 CS_BIAS.n508 0.189894
R25592 CS_BIAS.n510 CS_BIAS.n509 0.189894
R25593 CS_BIAS.n510 CS_BIAS.n400 0.189894
R25594 CS_BIAS.n514 CS_BIAS.n400 0.189894
R25595 CS_BIAS.n515 CS_BIAS.n514 0.189894
R25596 CS_BIAS.n515 CS_BIAS.n398 0.189894
R25597 CS_BIAS.n519 CS_BIAS.n398 0.189894
R25598 CS_BIAS.n520 CS_BIAS.n519 0.189894
R25599 CS_BIAS.n521 CS_BIAS.n520 0.189894
R25600 CS_BIAS.n521 CS_BIAS.n396 0.189894
R25601 CS_BIAS.n525 CS_BIAS.n396 0.189894
R25602 CS_BIAS.n526 CS_BIAS.n525 0.189894
R25603 CS_BIAS.n527 CS_BIAS.n526 0.189894
R25604 CS_BIAS.n527 CS_BIAS.n394 0.189894
R25605 CS_BIAS.n104 CS_BIAS.n85 0.170955
R25606 CS_BIAS.n108 CS_BIAS.n85 0.170955
R25607 CS_BIAS.n498 CS_BIAS.n479 0.170955
R25608 CS_BIAS.n502 CS_BIAS.n479 0.170955
R25609 a_n7864_n440.n0 a_n7864_n440.t24 235.603
R25610 a_n7864_n440.n0 a_n7864_n440.t22 235.603
R25611 a_n7864_n440.n1 a_n7864_n440.t23 235.603
R25612 a_n7864_n440.n1 a_n7864_n440.t20 235.603
R25613 a_n7864_n440.n4 a_n7864_n440.t21 235.603
R25614 a_n7864_n440.n22 a_n7864_n440.t4 60.4955
R25615 a_n7864_n440.n17 a_n7864_n440.t19 60.4955
R25616 a_n7864_n440.n15 a_n7864_n440.t6 60.4955
R25617 a_n7864_n440.n10 a_n7864_n440.t13 60.4955
R25618 a_n7864_n440.n19 a_n7864_n440.n18 56.3792
R25619 a_n7864_n440.n21 a_n7864_n440.n20 56.3792
R25620 a_n7864_n440.n3 a_n7864_n440.n2 56.3792
R25621 a_n7864_n440.n24 a_n7864_n440.n23 56.3791
R25622 a_n7864_n440.n14 a_n7864_n440.n13 56.379
R25623 a_n7864_n440.n12 a_n7864_n440.n11 56.379
R25624 a_n7864_n440.n9 a_n7864_n440.n8 56.379
R25625 a_n7864_n440.n7 a_n7864_n440.n6 56.379
R25626 a_n7864_n440.n5 a_n7864_n440.n3 13.6408
R25627 a_n7864_n440.n17 a_n7864_n440.n16 11.9791
R25628 a_n7864_n440.n7 a_n7864_n440.n5 8.22033
R25629 a_n7864_n440.n16 a_n7864_n440.n0 7.43194
R25630 a_n7864_n440.n16 a_n7864_n440.n15 6.55869
R25631 a_n7864_n440.n5 a_n7864_n440.n4 6.55694
R25632 a_n7864_n440.n18 a_n7864_n440.t11 4.11692
R25633 a_n7864_n440.n18 a_n7864_n440.t18 4.11692
R25634 a_n7864_n440.n20 a_n7864_n440.t14 4.11692
R25635 a_n7864_n440.n20 a_n7864_n440.t10 4.11692
R25636 a_n7864_n440.n2 a_n7864_n440.t3 4.11692
R25637 a_n7864_n440.n2 a_n7864_n440.t8 4.11692
R25638 a_n7864_n440.n13 a_n7864_n440.t0 4.11692
R25639 a_n7864_n440.n13 a_n7864_n440.t5 4.11692
R25640 a_n7864_n440.n11 a_n7864_n440.t2 4.11692
R25641 a_n7864_n440.n11 a_n7864_n440.t1 4.11692
R25642 a_n7864_n440.n8 a_n7864_n440.t15 4.11692
R25643 a_n7864_n440.n8 a_n7864_n440.t17 4.11692
R25644 a_n7864_n440.n6 a_n7864_n440.t12 4.11692
R25645 a_n7864_n440.n6 a_n7864_n440.t16 4.11692
R25646 a_n7864_n440.n24 a_n7864_n440.t7 4.11692
R25647 a_n7864_n440.t9 a_n7864_n440.n24 4.11692
R25648 a_n7864_n440.n9 a_n7864_n440.n7 3.32378
R25649 a_n7864_n440.n10 a_n7864_n440.n9 3.32378
R25650 a_n7864_n440.n14 a_n7864_n440.n12 3.32378
R25651 a_n7864_n440.n15 a_n7864_n440.n14 3.32378
R25652 a_n7864_n440.n23 a_n7864_n440.n3 3.32378
R25653 a_n7864_n440.n23 a_n7864_n440.n22 3.32378
R25654 a_n7864_n440.n21 a_n7864_n440.n19 3.32378
R25655 a_n7864_n440.n19 a_n7864_n440.n17 3.32378
R25656 a_n7864_n440.n1 a_n7864_n440.n0 2.03538
R25657 a_n7864_n440.n4 a_n7864_n440.n1 2.03538
R25658 a_n7864_n440.n12 a_n7864_n440.n10 1.89705
R25659 a_n7864_n440.n22 a_n7864_n440.n21 1.89705
R25660 a_n5588_7572.n13 a_n5588_7572.t10 94.727
R25661 a_n5588_7572.n7 a_n5588_7572.t6 94.727
R25662 a_n5588_7572.n2 a_n5588_7572.t14 94.7261
R25663 a_n5588_7572.n0 a_n5588_7572.t2 93.0158
R25664 a_n5588_7572.n0 a_n5588_7572.t3 93.0158
R25665 a_n5588_7572.n10 a_n5588_7572.t5 93.0158
R25666 a_n5588_7572.n13 a_n5588_7572.n12 87.1058
R25667 a_n5588_7572.n2 a_n5588_7572.n1 87.1058
R25668 a_n5588_7572.n4 a_n5588_7572.n3 87.1058
R25669 a_n5588_7572.n7 a_n5588_7572.n6 87.1058
R25670 a_n5588_7572.n9 a_n5588_7572.n8 87.1058
R25671 a_n5588_7572.n15 a_n5588_7572.n14 87.1058
R25672 a_n5588_7572.n14 a_n5588_7572.n11 28.6713
R25673 a_n5588_7572.n5 a_n5588_7572.t0 23.7194
R25674 a_n5588_7572.n5 a_n5588_7572.n4 8.5199
R25675 a_n5588_7572.n12 a_n5588_7572.t13 5.9105
R25676 a_n5588_7572.n12 a_n5588_7572.t18 5.9105
R25677 a_n5588_7572.n1 a_n5588_7572.t16 5.9105
R25678 a_n5588_7572.n1 a_n5588_7572.t15 5.9105
R25679 a_n5588_7572.n3 a_n5588_7572.t12 5.9105
R25680 a_n5588_7572.n3 a_n5588_7572.t11 5.9105
R25681 a_n5588_7572.n6 a_n5588_7572.t7 5.9105
R25682 a_n5588_7572.n6 a_n5588_7572.t4 5.9105
R25683 a_n5588_7572.n8 a_n5588_7572.t1 5.9105
R25684 a_n5588_7572.n8 a_n5588_7572.t8 5.9105
R25685 a_n5588_7572.t17 a_n5588_7572.n15 5.9105
R25686 a_n5588_7572.n15 a_n5588_7572.t9 5.9105
R25687 a_n5588_7572.n11 a_n5588_7572.n10 5.86149
R25688 a_n5588_7572.n11 a_n5588_7572.n5 4.01944
R25689 a_n5588_7572.n9 a_n5588_7572.n0 2.14921
R25690 a_n5588_7572.n4 a_n5588_7572.n2 1.71171
R25691 a_n5588_7572.n10 a_n5588_7572.n9 1.71171
R25692 a_n5588_7572.n0 a_n5588_7572.n7 1.71171
R25693 a_n5588_7572.n14 a_n5588_7572.n13 1.71171
R25694 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t5 134.996
R25695 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t1 133.98
R25696 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.t7 133.98
R25697 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.t3 133.98
R25698 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t9 133.98
R25699 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t10 133.05
R25700 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.t11 131.014
R25701 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.t14 131.014
R25702 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.t13 131.014
R25703 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t12 131.014
R25704 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.t4 90.6488
R25705 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.t0 88.6123
R25706 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.t6 88.6123
R25707 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.t2 88.6123
R25708 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.t8 88.6123
R25709 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 5.29232
R25710 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n4 4.34865
R25711 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n9 4.31215
R25712 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 2.03707
R25713 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 2.03707
R25714 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n5 2.03707
R25715 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n10 2.03704
R25716 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n11 2.03704
R25717 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n0 1.38231
R25718 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.n3 1.01794
R25719 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 1.01794
R25720 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 1.01794
R25721 DIFFPAIR_BIAS DIFFPAIR_BIAS.n13 0.684875
R25722 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n12 0.364533
C0 VDD VOUT 64.347305f
C1 VOUT VP 3.01986f
C2 VDD VN 0.14228f
C3 a_n8273_9606# VDD 1.45673f
C4 VOUT VN 1.27492f
C5 VP VN 17.7169f
C6 VOUT CS_BIAS 35.070602f
C7 VP CS_BIAS 0.593309f
C8 VP DIFFPAIR_BIAS 5.56e-19
C9 VN CS_BIAS 0.497337f
C10 VN DIFFPAIR_BIAS 0.001654f
C11 a_7389_9606# VDD 1.45673f
C12 DIFFPAIR_BIAS GND 36.1585f
C13 CS_BIAS GND 0.181673p
C14 VN GND 68.355545f
C15 VP GND 52.32566f
C16 VOUT GND 0.107159p
C17 VDD GND 0.689529p
C18 a_7389_9606# GND 0.466341f
C19 a_n8273_9606# GND 0.466341f
C20 a_n5588_7572.n0 GND 0.879122f
C21 a_n5588_7572.t0 GND 0.21498p
C22 a_n5588_7572.t9 GND 0.041533f
C23 a_n5588_7572.t14 GND 0.356358f
C24 a_n5588_7572.t16 GND 0.041533f
C25 a_n5588_7572.t15 GND 0.041533f
C26 a_n5588_7572.n1 GND 0.256861f
C27 a_n5588_7572.n2 GND 0.961829f
C28 a_n5588_7572.t12 GND 0.041533f
C29 a_n5588_7572.t11 GND 0.041533f
C30 a_n5588_7572.n3 GND 0.256861f
C31 a_n5588_7572.n4 GND 1.12737f
C32 a_n5588_7572.n5 GND 1.82143f
C33 a_n5588_7572.t6 GND 0.35636f
C34 a_n5588_7572.t7 GND 0.041533f
C35 a_n5588_7572.t4 GND 0.041533f
C36 a_n5588_7572.n6 GND 0.256861f
C37 a_n5588_7572.n7 GND 0.961827f
C38 a_n5588_7572.t2 GND 0.349253f
C39 a_n5588_7572.t3 GND 0.349253f
C40 a_n5588_7572.t1 GND 0.041533f
C41 a_n5588_7572.t8 GND 0.041533f
C42 a_n5588_7572.n8 GND 0.256861f
C43 a_n5588_7572.n9 GND 0.575559f
C44 a_n5588_7572.t5 GND 0.349253f
C45 a_n5588_7572.n10 GND 0.690769f
C46 a_n5588_7572.n11 GND 1.91489f
C47 a_n5588_7572.t10 GND 0.35636f
C48 a_n5588_7572.t13 GND 0.041533f
C49 a_n5588_7572.t18 GND 0.041533f
C50 a_n5588_7572.n12 GND 0.256861f
C51 a_n5588_7572.n13 GND 0.961827f
C52 a_n5588_7572.n14 GND 1.96937f
C53 a_n5588_7572.n15 GND 0.256861f
C54 a_n5588_7572.t17 GND 0.041533f
C55 a_n7864_n440.n0 GND 5.0054f
C56 a_n7864_n440.n1 GND 2.26937f
C57 a_n7864_n440.t7 GND 0.061304f
C58 a_n7864_n440.t3 GND 0.061304f
C59 a_n7864_n440.t8 GND 0.061304f
C60 a_n7864_n440.n2 GND 0.471051f
C61 a_n7864_n440.n3 GND 2.32754f
C62 a_n7864_n440.t24 GND 0.484983f
C63 a_n7864_n440.t22 GND 0.484983f
C64 a_n7864_n440.t23 GND 0.484983f
C65 a_n7864_n440.t20 GND 0.484983f
C66 a_n7864_n440.t21 GND 0.484983f
C67 a_n7864_n440.n4 GND 3.44474f
C68 a_n7864_n440.n5 GND 2.87778f
C69 a_n7864_n440.t12 GND 0.061304f
C70 a_n7864_n440.t16 GND 0.061304f
C71 a_n7864_n440.n6 GND 0.471049f
C72 a_n7864_n440.n7 GND 2.03673f
C73 a_n7864_n440.t15 GND 0.061304f
C74 a_n7864_n440.t17 GND 0.061304f
C75 a_n7864_n440.n8 GND 0.471049f
C76 a_n7864_n440.n9 GND 1.52042f
C77 a_n7864_n440.t13 GND 0.598981f
C78 a_n7864_n440.n10 GND 1.2631f
C79 a_n7864_n440.t2 GND 0.061304f
C80 a_n7864_n440.t1 GND 0.061304f
C81 a_n7864_n440.n11 GND 0.471049f
C82 a_n7864_n440.n12 GND 1.22384f
C83 a_n7864_n440.t0 GND 0.061304f
C84 a_n7864_n440.t5 GND 0.061304f
C85 a_n7864_n440.n13 GND 0.471049f
C86 a_n7864_n440.n14 GND 1.52042f
C87 a_n7864_n440.t6 GND 0.598981f
C88 a_n7864_n440.n15 GND 1.60349f
C89 a_n7864_n440.n16 GND 2.8734f
C90 a_n7864_n440.t19 GND 0.598981f
C91 a_n7864_n440.n17 GND 1.83586f
C92 a_n7864_n440.t11 GND 0.061304f
C93 a_n7864_n440.t18 GND 0.061304f
C94 a_n7864_n440.n18 GND 0.471051f
C95 a_n7864_n440.n19 GND 1.52042f
C96 a_n7864_n440.t14 GND 0.061304f
C97 a_n7864_n440.t10 GND 0.061304f
C98 a_n7864_n440.n20 GND 0.471051f
C99 a_n7864_n440.n21 GND 1.22384f
C100 a_n7864_n440.t4 GND 0.598985f
C101 a_n7864_n440.n22 GND 1.2631f
C102 a_n7864_n440.n23 GND 1.52042f
C103 a_n7864_n440.n24 GND 0.471052f
C104 a_n7864_n440.t9 GND 0.061304f
C105 CS_BIAS.n0 GND 0.013254f
C106 CS_BIAS.t27 GND 0.150431f
C107 CS_BIAS.n1 GND 0.013132f
C108 CS_BIAS.n2 GND 0.007046f
C109 CS_BIAS.n3 GND 0.013132f
C110 CS_BIAS.n4 GND 0.007046f
C111 CS_BIAS.t58 GND 0.150431f
C112 CS_BIAS.n5 GND 0.066478f
C113 CS_BIAS.n6 GND 0.007046f
C114 CS_BIAS.n7 GND 0.014173f
C115 CS_BIAS.n8 GND 0.007046f
C116 CS_BIAS.n9 GND 0.013132f
C117 CS_BIAS.n10 GND 0.013254f
C118 CS_BIAS.t0 GND 0.150431f
C119 CS_BIAS.n11 GND 0.013132f
C120 CS_BIAS.n12 GND 0.007046f
C121 CS_BIAS.n13 GND 0.013132f
C122 CS_BIAS.n14 GND 0.007046f
C123 CS_BIAS.t8 GND 0.150431f
C124 CS_BIAS.n15 GND 0.066478f
C125 CS_BIAS.n16 GND 0.007046f
C126 CS_BIAS.n17 GND 0.014173f
C127 CS_BIAS.n18 GND 0.007046f
C128 CS_BIAS.n19 GND 0.013132f
C129 CS_BIAS.n20 GND 0.007046f
C130 CS_BIAS.t2 GND 0.150431f
C131 CS_BIAS.n21 GND 0.013132f
C132 CS_BIAS.n22 GND 0.007046f
C133 CS_BIAS.n23 GND 0.014173f
C134 CS_BIAS.n24 GND 0.007046f
C135 CS_BIAS.t12 GND 0.150431f
C136 CS_BIAS.n25 GND 0.094199f
C137 CS_BIAS.t4 GND 0.24518f
C138 CS_BIAS.n26 GND 0.124966f
C139 CS_BIAS.n27 GND 0.096935f
C140 CS_BIAS.n28 GND 0.010798f
C141 CS_BIAS.n29 GND 0.013132f
C142 CS_BIAS.n30 GND 0.013132f
C143 CS_BIAS.n31 GND 0.007046f
C144 CS_BIAS.n32 GND 0.007046f
C145 CS_BIAS.n33 GND 0.007046f
C146 CS_BIAS.n34 GND 0.006465f
C147 CS_BIAS.n35 GND 0.013066f
C148 CS_BIAS.n36 GND 0.013132f
C149 CS_BIAS.n37 GND 0.007046f
C150 CS_BIAS.n38 GND 0.007046f
C151 CS_BIAS.n39 GND 0.007046f
C152 CS_BIAS.n40 GND 0.013132f
C153 CS_BIAS.n41 GND 0.073127f
C154 CS_BIAS.n42 GND 0.013132f
C155 CS_BIAS.n43 GND 0.007046f
C156 CS_BIAS.n44 GND 0.007046f
C157 CS_BIAS.n45 GND 0.007046f
C158 CS_BIAS.n46 GND 0.013132f
C159 CS_BIAS.n47 GND 0.013066f
C160 CS_BIAS.n48 GND 0.006465f
C161 CS_BIAS.n49 GND 0.007046f
C162 CS_BIAS.n50 GND 0.007046f
C163 CS_BIAS.n51 GND 0.007046f
C164 CS_BIAS.n52 GND 0.013132f
C165 CS_BIAS.n53 GND 0.013132f
C166 CS_BIAS.n54 GND 0.010798f
C167 CS_BIAS.n55 GND 0.007046f
C168 CS_BIAS.n56 GND 0.007046f
C169 CS_BIAS.n57 GND 0.008983f
C170 CS_BIAS.n58 GND 0.013132f
C171 CS_BIAS.n59 GND 0.013132f
C172 CS_BIAS.n60 GND 0.007046f
C173 CS_BIAS.n61 GND 0.007046f
C174 CS_BIAS.n62 GND 0.007046f
C175 CS_BIAS.n63 GND 0.009893f
C176 CS_BIAS.n64 GND 0.010679f
C177 CS_BIAS.n65 GND 0.013132f
C178 CS_BIAS.n66 GND 0.007046f
C179 CS_BIAS.n67 GND 0.007046f
C180 CS_BIAS.n68 GND 0.007046f
C181 CS_BIAS.n69 GND 0.013132f
C182 CS_BIAS.n70 GND 0.008464f
C183 CS_BIAS.n71 GND 0.094465f
C184 CS_BIAS.n72 GND 0.082592f
C185 CS_BIAS.n73 GND 0.004068f
C186 CS_BIAS.n74 GND 0.008981f
C187 CS_BIAS.t1 GND 0.006732f
C188 CS_BIAS.n75 GND 0.007046f
C189 CS_BIAS.n76 GND 0.00224f
C190 CS_BIAS.n77 GND 0.001477f
C191 CS_BIAS.n78 GND 0.019904f
C192 CS_BIAS.n79 GND 0.00827f
C193 CS_BIAS.n80 GND 0.115089f
C194 CS_BIAS.t9 GND 0.004409f
C195 CS_BIAS.t3 GND 0.004409f
C196 CS_BIAS.n81 GND 0.031231f
C197 CS_BIAS.n82 GND 0.113505f
C198 CS_BIAS.t13 GND 0.004409f
C199 CS_BIAS.t5 GND 0.004409f
C200 CS_BIAS.n83 GND 0.033215f
C201 CS_BIAS.n84 GND 0.266267f
C202 CS_BIAS.n85 GND 0.050936f
C203 CS_BIAS.t24 GND 0.150431f
C204 CS_BIAS.n86 GND 0.013132f
C205 CS_BIAS.n87 GND 0.007046f
C206 CS_BIAS.n88 GND 0.014173f
C207 CS_BIAS.n89 GND 0.007046f
C208 CS_BIAS.t47 GND 0.150431f
C209 CS_BIAS.n90 GND 0.094199f
C210 CS_BIAS.t22 GND 0.24518f
C211 CS_BIAS.n91 GND 0.124966f
C212 CS_BIAS.n92 GND 0.096935f
C213 CS_BIAS.n93 GND 0.010798f
C214 CS_BIAS.n94 GND 0.013132f
C215 CS_BIAS.n95 GND 0.013132f
C216 CS_BIAS.n96 GND 0.007046f
C217 CS_BIAS.n97 GND 0.007046f
C218 CS_BIAS.n98 GND 0.007046f
C219 CS_BIAS.n99 GND 0.006465f
C220 CS_BIAS.n100 GND 0.013066f
C221 CS_BIAS.n101 GND 0.013132f
C222 CS_BIAS.n102 GND 0.007046f
C223 CS_BIAS.n103 GND 0.007046f
C224 CS_BIAS.n104 GND 0.007012f
C225 CS_BIAS.n105 GND 0.013132f
C226 CS_BIAS.n106 GND 0.073127f
C227 CS_BIAS.n107 GND 0.013132f
C228 CS_BIAS.n108 GND 0.007012f
C229 CS_BIAS.n109 GND 0.007046f
C230 CS_BIAS.n110 GND 0.007046f
C231 CS_BIAS.n111 GND 0.013132f
C232 CS_BIAS.n112 GND 0.013066f
C233 CS_BIAS.n113 GND 0.006465f
C234 CS_BIAS.n114 GND 0.007046f
C235 CS_BIAS.n115 GND 0.007046f
C236 CS_BIAS.n116 GND 0.007046f
C237 CS_BIAS.n117 GND 0.013132f
C238 CS_BIAS.n118 GND 0.013132f
C239 CS_BIAS.n119 GND 0.010798f
C240 CS_BIAS.n120 GND 0.007046f
C241 CS_BIAS.n121 GND 0.007046f
C242 CS_BIAS.n122 GND 0.008983f
C243 CS_BIAS.n123 GND 0.013132f
C244 CS_BIAS.n124 GND 0.013132f
C245 CS_BIAS.n125 GND 0.007046f
C246 CS_BIAS.n126 GND 0.007046f
C247 CS_BIAS.n127 GND 0.007046f
C248 CS_BIAS.n128 GND 0.009893f
C249 CS_BIAS.n129 GND 0.010679f
C250 CS_BIAS.n130 GND 0.013132f
C251 CS_BIAS.n131 GND 0.007046f
C252 CS_BIAS.n132 GND 0.007046f
C253 CS_BIAS.n133 GND 0.007046f
C254 CS_BIAS.n134 GND 0.013132f
C255 CS_BIAS.n135 GND 0.008464f
C256 CS_BIAS.n136 GND 0.094465f
C257 CS_BIAS.n137 GND 0.063508f
C258 CS_BIAS.n138 GND 0.013254f
C259 CS_BIAS.t53 GND 0.150431f
C260 CS_BIAS.n139 GND 0.013132f
C261 CS_BIAS.n140 GND 0.007046f
C262 CS_BIAS.n141 GND 0.013132f
C263 CS_BIAS.n142 GND 0.007046f
C264 CS_BIAS.t20 GND 0.150431f
C265 CS_BIAS.n143 GND 0.066478f
C266 CS_BIAS.n144 GND 0.007046f
C267 CS_BIAS.n145 GND 0.014173f
C268 CS_BIAS.n146 GND 0.007046f
C269 CS_BIAS.n147 GND 0.013132f
C270 CS_BIAS.n148 GND 0.007046f
C271 CS_BIAS.t34 GND 0.150431f
C272 CS_BIAS.n149 GND 0.013132f
C273 CS_BIAS.n150 GND 0.007046f
C274 CS_BIAS.n151 GND 0.014173f
C275 CS_BIAS.n152 GND 0.007046f
C276 CS_BIAS.t55 GND 0.150431f
C277 CS_BIAS.n153 GND 0.094199f
C278 CS_BIAS.t21 GND 0.24518f
C279 CS_BIAS.n154 GND 0.124966f
C280 CS_BIAS.n155 GND 0.096935f
C281 CS_BIAS.n156 GND 0.010798f
C282 CS_BIAS.n157 GND 0.013132f
C283 CS_BIAS.n158 GND 0.013132f
C284 CS_BIAS.n159 GND 0.007046f
C285 CS_BIAS.n160 GND 0.007046f
C286 CS_BIAS.n161 GND 0.007046f
C287 CS_BIAS.n162 GND 0.006465f
C288 CS_BIAS.n163 GND 0.013066f
C289 CS_BIAS.n164 GND 0.013132f
C290 CS_BIAS.n165 GND 0.007046f
C291 CS_BIAS.n166 GND 0.007046f
C292 CS_BIAS.n167 GND 0.007046f
C293 CS_BIAS.n168 GND 0.013132f
C294 CS_BIAS.n169 GND 0.073127f
C295 CS_BIAS.n170 GND 0.013132f
C296 CS_BIAS.n171 GND 0.007046f
C297 CS_BIAS.n172 GND 0.007046f
C298 CS_BIAS.n173 GND 0.007046f
C299 CS_BIAS.n174 GND 0.013132f
C300 CS_BIAS.n175 GND 0.013066f
C301 CS_BIAS.n176 GND 0.006465f
C302 CS_BIAS.n177 GND 0.007046f
C303 CS_BIAS.n178 GND 0.007046f
C304 CS_BIAS.n179 GND 0.007046f
C305 CS_BIAS.n180 GND 0.013132f
C306 CS_BIAS.n181 GND 0.013132f
C307 CS_BIAS.n182 GND 0.010798f
C308 CS_BIAS.n183 GND 0.007046f
C309 CS_BIAS.n184 GND 0.007046f
C310 CS_BIAS.n185 GND 0.008983f
C311 CS_BIAS.n186 GND 0.013132f
C312 CS_BIAS.n187 GND 0.013132f
C313 CS_BIAS.n188 GND 0.007046f
C314 CS_BIAS.n189 GND 0.007046f
C315 CS_BIAS.n190 GND 0.007046f
C316 CS_BIAS.n191 GND 0.009893f
C317 CS_BIAS.n192 GND 0.010679f
C318 CS_BIAS.n193 GND 0.013132f
C319 CS_BIAS.n194 GND 0.007046f
C320 CS_BIAS.n195 GND 0.007046f
C321 CS_BIAS.n196 GND 0.007046f
C322 CS_BIAS.n197 GND 0.013132f
C323 CS_BIAS.n198 GND 0.008464f
C324 CS_BIAS.n199 GND 0.094465f
C325 CS_BIAS.n200 GND 0.056596f
C326 CS_BIAS.n201 GND 0.066547f
C327 CS_BIAS.n202 GND 0.013254f
C328 CS_BIAS.t41 GND 0.150431f
C329 CS_BIAS.n203 GND 0.013132f
C330 CS_BIAS.n204 GND 0.007046f
C331 CS_BIAS.n205 GND 0.013132f
C332 CS_BIAS.n206 GND 0.007046f
C333 CS_BIAS.t67 GND 0.150431f
C334 CS_BIAS.n207 GND 0.066478f
C335 CS_BIAS.n208 GND 0.007046f
C336 CS_BIAS.n209 GND 0.014173f
C337 CS_BIAS.n210 GND 0.007046f
C338 CS_BIAS.n211 GND 0.013132f
C339 CS_BIAS.n212 GND 0.007046f
C340 CS_BIAS.t26 GND 0.150431f
C341 CS_BIAS.n213 GND 0.013132f
C342 CS_BIAS.n214 GND 0.007046f
C343 CS_BIAS.n215 GND 0.014173f
C344 CS_BIAS.n216 GND 0.007046f
C345 CS_BIAS.t49 GND 0.150431f
C346 CS_BIAS.n217 GND 0.094199f
C347 CS_BIAS.t62 GND 0.24518f
C348 CS_BIAS.n218 GND 0.124966f
C349 CS_BIAS.n219 GND 0.096935f
C350 CS_BIAS.n220 GND 0.010798f
C351 CS_BIAS.n221 GND 0.013132f
C352 CS_BIAS.n222 GND 0.013132f
C353 CS_BIAS.n223 GND 0.007046f
C354 CS_BIAS.n224 GND 0.007046f
C355 CS_BIAS.n225 GND 0.007046f
C356 CS_BIAS.n226 GND 0.006465f
C357 CS_BIAS.n227 GND 0.013066f
C358 CS_BIAS.n228 GND 0.013132f
C359 CS_BIAS.n229 GND 0.007046f
C360 CS_BIAS.n230 GND 0.007046f
C361 CS_BIAS.n231 GND 0.007046f
C362 CS_BIAS.n232 GND 0.013132f
C363 CS_BIAS.n233 GND 0.073127f
C364 CS_BIAS.n234 GND 0.013132f
C365 CS_BIAS.n235 GND 0.007046f
C366 CS_BIAS.n236 GND 0.007046f
C367 CS_BIAS.n237 GND 0.007046f
C368 CS_BIAS.n238 GND 0.013132f
C369 CS_BIAS.n239 GND 0.013066f
C370 CS_BIAS.n240 GND 0.006465f
C371 CS_BIAS.n241 GND 0.007046f
C372 CS_BIAS.n242 GND 0.007046f
C373 CS_BIAS.n243 GND 0.007046f
C374 CS_BIAS.n244 GND 0.013132f
C375 CS_BIAS.n245 GND 0.013132f
C376 CS_BIAS.n246 GND 0.010798f
C377 CS_BIAS.n247 GND 0.007046f
C378 CS_BIAS.n248 GND 0.007046f
C379 CS_BIAS.n249 GND 0.008983f
C380 CS_BIAS.n250 GND 0.013132f
C381 CS_BIAS.n251 GND 0.013132f
C382 CS_BIAS.n252 GND 0.007046f
C383 CS_BIAS.n253 GND 0.007046f
C384 CS_BIAS.n254 GND 0.007046f
C385 CS_BIAS.n255 GND 0.009893f
C386 CS_BIAS.n256 GND 0.010679f
C387 CS_BIAS.n257 GND 0.013132f
C388 CS_BIAS.n258 GND 0.007046f
C389 CS_BIAS.n259 GND 0.007046f
C390 CS_BIAS.n260 GND 0.007046f
C391 CS_BIAS.n261 GND 0.013132f
C392 CS_BIAS.n262 GND 0.008464f
C393 CS_BIAS.n263 GND 0.094465f
C394 CS_BIAS.n264 GND 0.056596f
C395 CS_BIAS.n265 GND 0.046396f
C396 CS_BIAS.n266 GND 0.013254f
C397 CS_BIAS.t36 GND 0.150431f
C398 CS_BIAS.n267 GND 0.013132f
C399 CS_BIAS.n268 GND 0.007046f
C400 CS_BIAS.n269 GND 0.013132f
C401 CS_BIAS.n270 GND 0.007046f
C402 CS_BIAS.t57 GND 0.150431f
C403 CS_BIAS.n271 GND 0.066478f
C404 CS_BIAS.n272 GND 0.007046f
C405 CS_BIAS.n273 GND 0.014173f
C406 CS_BIAS.n274 GND 0.007046f
C407 CS_BIAS.n275 GND 0.013132f
C408 CS_BIAS.n276 GND 0.007046f
C409 CS_BIAS.t23 GND 0.150431f
C410 CS_BIAS.n277 GND 0.013132f
C411 CS_BIAS.n278 GND 0.007046f
C412 CS_BIAS.n279 GND 0.014173f
C413 CS_BIAS.n280 GND 0.007046f
C414 CS_BIAS.t38 GND 0.150431f
C415 CS_BIAS.n281 GND 0.094199f
C416 CS_BIAS.t59 GND 0.24518f
C417 CS_BIAS.n282 GND 0.124966f
C418 CS_BIAS.n283 GND 0.096935f
C419 CS_BIAS.n284 GND 0.010798f
C420 CS_BIAS.n285 GND 0.013132f
C421 CS_BIAS.n286 GND 0.013132f
C422 CS_BIAS.n287 GND 0.007046f
C423 CS_BIAS.n288 GND 0.007046f
C424 CS_BIAS.n289 GND 0.007046f
C425 CS_BIAS.n290 GND 0.006465f
C426 CS_BIAS.n291 GND 0.013066f
C427 CS_BIAS.n292 GND 0.013132f
C428 CS_BIAS.n293 GND 0.007046f
C429 CS_BIAS.n294 GND 0.007046f
C430 CS_BIAS.n295 GND 0.007046f
C431 CS_BIAS.n296 GND 0.013132f
C432 CS_BIAS.n297 GND 0.073127f
C433 CS_BIAS.n298 GND 0.013132f
C434 CS_BIAS.n299 GND 0.007046f
C435 CS_BIAS.n300 GND 0.007046f
C436 CS_BIAS.n301 GND 0.007046f
C437 CS_BIAS.n302 GND 0.013132f
C438 CS_BIAS.n303 GND 0.013066f
C439 CS_BIAS.n304 GND 0.006465f
C440 CS_BIAS.n305 GND 0.007046f
C441 CS_BIAS.n306 GND 0.007046f
C442 CS_BIAS.n307 GND 0.007046f
C443 CS_BIAS.n308 GND 0.013132f
C444 CS_BIAS.n309 GND 0.013132f
C445 CS_BIAS.n310 GND 0.010798f
C446 CS_BIAS.n311 GND 0.007046f
C447 CS_BIAS.n312 GND 0.007046f
C448 CS_BIAS.n313 GND 0.008983f
C449 CS_BIAS.n314 GND 0.013132f
C450 CS_BIAS.n315 GND 0.013132f
C451 CS_BIAS.n316 GND 0.007046f
C452 CS_BIAS.n317 GND 0.007046f
C453 CS_BIAS.n318 GND 0.007046f
C454 CS_BIAS.n319 GND 0.009893f
C455 CS_BIAS.n320 GND 0.010679f
C456 CS_BIAS.n321 GND 0.013132f
C457 CS_BIAS.n322 GND 0.007046f
C458 CS_BIAS.n323 GND 0.007046f
C459 CS_BIAS.n324 GND 0.007046f
C460 CS_BIAS.n325 GND 0.013132f
C461 CS_BIAS.n326 GND 0.008464f
C462 CS_BIAS.n327 GND 0.094465f
C463 CS_BIAS.n328 GND 0.056596f
C464 CS_BIAS.n329 GND 0.046396f
C465 CS_BIAS.n330 GND 0.013254f
C466 CS_BIAS.t31 GND 0.150431f
C467 CS_BIAS.n331 GND 0.013132f
C468 CS_BIAS.n332 GND 0.007046f
C469 CS_BIAS.n333 GND 0.013132f
C470 CS_BIAS.n334 GND 0.007046f
C471 CS_BIAS.t48 GND 0.150431f
C472 CS_BIAS.n335 GND 0.066478f
C473 CS_BIAS.n336 GND 0.007046f
C474 CS_BIAS.n337 GND 0.014173f
C475 CS_BIAS.n338 GND 0.007046f
C476 CS_BIAS.n339 GND 0.013132f
C477 CS_BIAS.n340 GND 0.007046f
C478 CS_BIAS.t68 GND 0.150431f
C479 CS_BIAS.n341 GND 0.013132f
C480 CS_BIAS.n342 GND 0.007046f
C481 CS_BIAS.n343 GND 0.014173f
C482 CS_BIAS.n344 GND 0.007046f
C483 CS_BIAS.t32 GND 0.150431f
C484 CS_BIAS.n345 GND 0.094199f
C485 CS_BIAS.t51 GND 0.245181f
C486 CS_BIAS.n346 GND 0.124966f
C487 CS_BIAS.n347 GND 0.096934f
C488 CS_BIAS.n348 GND 0.010798f
C489 CS_BIAS.n349 GND 0.013132f
C490 CS_BIAS.n350 GND 0.013132f
C491 CS_BIAS.n351 GND 0.007046f
C492 CS_BIAS.n352 GND 0.007046f
C493 CS_BIAS.n353 GND 0.007046f
C494 CS_BIAS.n354 GND 0.006465f
C495 CS_BIAS.n355 GND 0.013066f
C496 CS_BIAS.n356 GND 0.013132f
C497 CS_BIAS.n357 GND 0.007046f
C498 CS_BIAS.n358 GND 0.007046f
C499 CS_BIAS.n359 GND 0.007046f
C500 CS_BIAS.n360 GND 0.013132f
C501 CS_BIAS.n361 GND 0.073127f
C502 CS_BIAS.n362 GND 0.013132f
C503 CS_BIAS.n363 GND 0.007046f
C504 CS_BIAS.n364 GND 0.007046f
C505 CS_BIAS.n365 GND 0.007046f
C506 CS_BIAS.n366 GND 0.013132f
C507 CS_BIAS.n367 GND 0.013066f
C508 CS_BIAS.n368 GND 0.006465f
C509 CS_BIAS.n369 GND 0.007046f
C510 CS_BIAS.n370 GND 0.007046f
C511 CS_BIAS.n371 GND 0.007046f
C512 CS_BIAS.n372 GND 0.013132f
C513 CS_BIAS.n373 GND 0.013132f
C514 CS_BIAS.n374 GND 0.010798f
C515 CS_BIAS.n375 GND 0.007046f
C516 CS_BIAS.n376 GND 0.007046f
C517 CS_BIAS.n377 GND 0.008983f
C518 CS_BIAS.n378 GND 0.013132f
C519 CS_BIAS.n379 GND 0.013132f
C520 CS_BIAS.n380 GND 0.007046f
C521 CS_BIAS.n381 GND 0.007046f
C522 CS_BIAS.n382 GND 0.007046f
C523 CS_BIAS.n383 GND 0.009893f
C524 CS_BIAS.n384 GND 0.010679f
C525 CS_BIAS.n385 GND 0.013132f
C526 CS_BIAS.n386 GND 0.007046f
C527 CS_BIAS.n387 GND 0.007046f
C528 CS_BIAS.n388 GND 0.007046f
C529 CS_BIAS.n389 GND 0.013132f
C530 CS_BIAS.n390 GND 0.008464f
C531 CS_BIAS.n391 GND 0.094465f
C532 CS_BIAS.n392 GND 0.056596f
C533 CS_BIAS.n393 GND 0.966542f
C534 CS_BIAS.n394 GND 0.013254f
C535 CS_BIAS.t46 GND 0.150431f
C536 CS_BIAS.n395 GND 0.013132f
C537 CS_BIAS.n396 GND 0.007046f
C538 CS_BIAS.n397 GND 0.013132f
C539 CS_BIAS.n398 GND 0.007046f
C540 CS_BIAS.t37 GND 0.150431f
C541 CS_BIAS.n399 GND 0.066478f
C542 CS_BIAS.n400 GND 0.007046f
C543 CS_BIAS.n401 GND 0.014173f
C544 CS_BIAS.n402 GND 0.007046f
C545 CS_BIAS.n403 GND 0.013132f
C546 CS_BIAS.n404 GND 0.004068f
C547 CS_BIAS.n405 GND 0.008981f
C548 CS_BIAS.t11 GND 0.006732f
C549 CS_BIAS.n406 GND 0.007046f
C550 CS_BIAS.n407 GND 0.00224f
C551 CS_BIAS.n408 GND 0.001477f
C552 CS_BIAS.n409 GND 0.019904f
C553 CS_BIAS.n410 GND 0.010785f
C554 CS_BIAS.t19 GND 0.004409f
C555 CS_BIAS.t7 GND 0.004409f
C556 CS_BIAS.n411 GND 0.031231f
C557 CS_BIAS.n412 GND 0.192849f
C558 CS_BIAS.n413 GND 0.013254f
C559 CS_BIAS.t14 GND 0.150431f
C560 CS_BIAS.n414 GND 0.013132f
C561 CS_BIAS.n415 GND 0.007046f
C562 CS_BIAS.n416 GND 0.013132f
C563 CS_BIAS.n417 GND 0.007046f
C564 CS_BIAS.t16 GND 0.150431f
C565 CS_BIAS.n418 GND 0.066478f
C566 CS_BIAS.n419 GND 0.007046f
C567 CS_BIAS.n420 GND 0.014173f
C568 CS_BIAS.n421 GND 0.007046f
C569 CS_BIAS.n422 GND 0.013132f
C570 CS_BIAS.n423 GND 0.007046f
C571 CS_BIAS.t6 GND 0.150431f
C572 CS_BIAS.n424 GND 0.013132f
C573 CS_BIAS.n425 GND 0.007046f
C574 CS_BIAS.n426 GND 0.014173f
C575 CS_BIAS.n427 GND 0.007046f
C576 CS_BIAS.t18 GND 0.150431f
C577 CS_BIAS.n428 GND 0.094199f
C578 CS_BIAS.t10 GND 0.245181f
C579 CS_BIAS.n429 GND 0.124966f
C580 CS_BIAS.n430 GND 0.096934f
C581 CS_BIAS.n431 GND 0.010798f
C582 CS_BIAS.n432 GND 0.013132f
C583 CS_BIAS.n433 GND 0.013132f
C584 CS_BIAS.n434 GND 0.007046f
C585 CS_BIAS.n435 GND 0.007046f
C586 CS_BIAS.n436 GND 0.007046f
C587 CS_BIAS.n437 GND 0.006465f
C588 CS_BIAS.n438 GND 0.013066f
C589 CS_BIAS.n439 GND 0.013132f
C590 CS_BIAS.n440 GND 0.007046f
C591 CS_BIAS.n441 GND 0.007046f
C592 CS_BIAS.n442 GND 0.007046f
C593 CS_BIAS.n443 GND 0.013132f
C594 CS_BIAS.n444 GND 0.073127f
C595 CS_BIAS.n445 GND 0.013132f
C596 CS_BIAS.n446 GND 0.007046f
C597 CS_BIAS.n447 GND 0.007046f
C598 CS_BIAS.n448 GND 0.007046f
C599 CS_BIAS.n449 GND 0.013132f
C600 CS_BIAS.n450 GND 0.013066f
C601 CS_BIAS.n451 GND 0.006465f
C602 CS_BIAS.n452 GND 0.007046f
C603 CS_BIAS.n453 GND 0.007046f
C604 CS_BIAS.n454 GND 0.007046f
C605 CS_BIAS.n455 GND 0.013132f
C606 CS_BIAS.n456 GND 0.013132f
C607 CS_BIAS.n457 GND 0.010798f
C608 CS_BIAS.n458 GND 0.007046f
C609 CS_BIAS.n459 GND 0.007046f
C610 CS_BIAS.n460 GND 0.008983f
C611 CS_BIAS.n461 GND 0.013132f
C612 CS_BIAS.n462 GND 0.013132f
C613 CS_BIAS.n463 GND 0.007046f
C614 CS_BIAS.n464 GND 0.007046f
C615 CS_BIAS.n465 GND 0.007046f
C616 CS_BIAS.n466 GND 0.009893f
C617 CS_BIAS.n467 GND 0.010679f
C618 CS_BIAS.n468 GND 0.013132f
C619 CS_BIAS.n469 GND 0.007046f
C620 CS_BIAS.n470 GND 0.007046f
C621 CS_BIAS.n471 GND 0.007046f
C622 CS_BIAS.n472 GND 0.013132f
C623 CS_BIAS.n473 GND 0.008464f
C624 CS_BIAS.n474 GND 0.094465f
C625 CS_BIAS.n475 GND 0.088669f
C626 CS_BIAS.t17 GND 0.004409f
C627 CS_BIAS.t15 GND 0.004409f
C628 CS_BIAS.n476 GND 0.031231f
C629 CS_BIAS.n477 GND 0.179676f
C630 CS_BIAS.n478 GND 0.115728f
C631 CS_BIAS.n479 GND 0.050936f
C632 CS_BIAS.t60 GND 0.150431f
C633 CS_BIAS.n480 GND 0.013132f
C634 CS_BIAS.n481 GND 0.007046f
C635 CS_BIAS.n482 GND 0.014173f
C636 CS_BIAS.n483 GND 0.007046f
C637 CS_BIAS.t30 GND 0.150431f
C638 CS_BIAS.n484 GND 0.094199f
C639 CS_BIAS.t56 GND 0.245181f
C640 CS_BIAS.n485 GND 0.124966f
C641 CS_BIAS.n486 GND 0.096934f
C642 CS_BIAS.n487 GND 0.010798f
C643 CS_BIAS.n488 GND 0.013132f
C644 CS_BIAS.n489 GND 0.013132f
C645 CS_BIAS.n490 GND 0.007046f
C646 CS_BIAS.n491 GND 0.007046f
C647 CS_BIAS.n492 GND 0.007046f
C648 CS_BIAS.n493 GND 0.006465f
C649 CS_BIAS.n494 GND 0.013066f
C650 CS_BIAS.n495 GND 0.013132f
C651 CS_BIAS.n496 GND 0.007046f
C652 CS_BIAS.n497 GND 0.007046f
C653 CS_BIAS.n498 GND 0.007012f
C654 CS_BIAS.n499 GND 0.013132f
C655 CS_BIAS.n500 GND 0.073127f
C656 CS_BIAS.n501 GND 0.013132f
C657 CS_BIAS.n502 GND 0.007012f
C658 CS_BIAS.n503 GND 0.007046f
C659 CS_BIAS.n504 GND 0.007046f
C660 CS_BIAS.n505 GND 0.013132f
C661 CS_BIAS.n506 GND 0.013066f
C662 CS_BIAS.n507 GND 0.006465f
C663 CS_BIAS.n508 GND 0.007046f
C664 CS_BIAS.n509 GND 0.007046f
C665 CS_BIAS.n510 GND 0.007046f
C666 CS_BIAS.n511 GND 0.013132f
C667 CS_BIAS.n512 GND 0.013132f
C668 CS_BIAS.n513 GND 0.010798f
C669 CS_BIAS.n514 GND 0.007046f
C670 CS_BIAS.n515 GND 0.007046f
C671 CS_BIAS.n516 GND 0.008983f
C672 CS_BIAS.n517 GND 0.013132f
C673 CS_BIAS.n518 GND 0.013132f
C674 CS_BIAS.n519 GND 0.007046f
C675 CS_BIAS.n520 GND 0.007046f
C676 CS_BIAS.n521 GND 0.007046f
C677 CS_BIAS.n522 GND 0.009893f
C678 CS_BIAS.n523 GND 0.010679f
C679 CS_BIAS.n524 GND 0.013132f
C680 CS_BIAS.n525 GND 0.007046f
C681 CS_BIAS.n526 GND 0.007046f
C682 CS_BIAS.n527 GND 0.007046f
C683 CS_BIAS.n528 GND 0.013132f
C684 CS_BIAS.n529 GND 0.008464f
C685 CS_BIAS.n530 GND 0.094465f
C686 CS_BIAS.n531 GND 0.063508f
C687 CS_BIAS.n532 GND 0.013254f
C688 CS_BIAS.t61 GND 0.150431f
C689 CS_BIAS.n533 GND 0.013132f
C690 CS_BIAS.n534 GND 0.007046f
C691 CS_BIAS.n535 GND 0.013132f
C692 CS_BIAS.n536 GND 0.007046f
C693 CS_BIAS.t64 GND 0.150431f
C694 CS_BIAS.n537 GND 0.066478f
C695 CS_BIAS.n538 GND 0.007046f
C696 CS_BIAS.n539 GND 0.014173f
C697 CS_BIAS.n540 GND 0.007046f
C698 CS_BIAS.n541 GND 0.013132f
C699 CS_BIAS.n542 GND 0.007046f
C700 CS_BIAS.t29 GND 0.150431f
C701 CS_BIAS.n543 GND 0.013132f
C702 CS_BIAS.n544 GND 0.007046f
C703 CS_BIAS.n545 GND 0.014173f
C704 CS_BIAS.n546 GND 0.007046f
C705 CS_BIAS.t45 GND 0.150431f
C706 CS_BIAS.n547 GND 0.094199f
C707 CS_BIAS.t65 GND 0.245181f
C708 CS_BIAS.n548 GND 0.124966f
C709 CS_BIAS.n549 GND 0.096934f
C710 CS_BIAS.n550 GND 0.010798f
C711 CS_BIAS.n551 GND 0.013132f
C712 CS_BIAS.n552 GND 0.013132f
C713 CS_BIAS.n553 GND 0.007046f
C714 CS_BIAS.n554 GND 0.007046f
C715 CS_BIAS.n555 GND 0.007046f
C716 CS_BIAS.n556 GND 0.006465f
C717 CS_BIAS.n557 GND 0.013066f
C718 CS_BIAS.n558 GND 0.013132f
C719 CS_BIAS.n559 GND 0.007046f
C720 CS_BIAS.n560 GND 0.007046f
C721 CS_BIAS.n561 GND 0.007046f
C722 CS_BIAS.n562 GND 0.013132f
C723 CS_BIAS.n563 GND 0.073127f
C724 CS_BIAS.n564 GND 0.013132f
C725 CS_BIAS.n565 GND 0.007046f
C726 CS_BIAS.n566 GND 0.007046f
C727 CS_BIAS.n567 GND 0.007046f
C728 CS_BIAS.n568 GND 0.013132f
C729 CS_BIAS.n569 GND 0.013066f
C730 CS_BIAS.n570 GND 0.006465f
C731 CS_BIAS.n571 GND 0.007046f
C732 CS_BIAS.n572 GND 0.007046f
C733 CS_BIAS.n573 GND 0.007046f
C734 CS_BIAS.n574 GND 0.013132f
C735 CS_BIAS.n575 GND 0.013132f
C736 CS_BIAS.n576 GND 0.010798f
C737 CS_BIAS.n577 GND 0.007046f
C738 CS_BIAS.n578 GND 0.007046f
C739 CS_BIAS.n579 GND 0.008983f
C740 CS_BIAS.n580 GND 0.013132f
C741 CS_BIAS.n581 GND 0.013132f
C742 CS_BIAS.n582 GND 0.007046f
C743 CS_BIAS.n583 GND 0.007046f
C744 CS_BIAS.n584 GND 0.007046f
C745 CS_BIAS.n585 GND 0.009893f
C746 CS_BIAS.n586 GND 0.010679f
C747 CS_BIAS.n587 GND 0.013132f
C748 CS_BIAS.n588 GND 0.007046f
C749 CS_BIAS.n589 GND 0.007046f
C750 CS_BIAS.n590 GND 0.007046f
C751 CS_BIAS.n591 GND 0.013132f
C752 CS_BIAS.n592 GND 0.008464f
C753 CS_BIAS.n593 GND 0.094465f
C754 CS_BIAS.n594 GND 0.056596f
C755 CS_BIAS.n595 GND 0.066547f
C756 CS_BIAS.n596 GND 0.013254f
C757 CS_BIAS.t66 GND 0.150431f
C758 CS_BIAS.n597 GND 0.013132f
C759 CS_BIAS.n598 GND 0.007046f
C760 CS_BIAS.n599 GND 0.013132f
C761 CS_BIAS.n600 GND 0.007046f
C762 CS_BIAS.t39 GND 0.150431f
C763 CS_BIAS.n601 GND 0.066478f
C764 CS_BIAS.n602 GND 0.007046f
C765 CS_BIAS.n603 GND 0.014173f
C766 CS_BIAS.n604 GND 0.007046f
C767 CS_BIAS.n605 GND 0.013132f
C768 CS_BIAS.n606 GND 0.007046f
C769 CS_BIAS.t54 GND 0.150431f
C770 CS_BIAS.n607 GND 0.013132f
C771 CS_BIAS.n608 GND 0.007046f
C772 CS_BIAS.n609 GND 0.014173f
C773 CS_BIAS.n610 GND 0.007046f
C774 CS_BIAS.t25 GND 0.150431f
C775 CS_BIAS.n611 GND 0.094199f
C776 CS_BIAS.t35 GND 0.245181f
C777 CS_BIAS.n612 GND 0.124966f
C778 CS_BIAS.n613 GND 0.096934f
C779 CS_BIAS.n614 GND 0.010798f
C780 CS_BIAS.n615 GND 0.013132f
C781 CS_BIAS.n616 GND 0.013132f
C782 CS_BIAS.n617 GND 0.007046f
C783 CS_BIAS.n618 GND 0.007046f
C784 CS_BIAS.n619 GND 0.007046f
C785 CS_BIAS.n620 GND 0.006465f
C786 CS_BIAS.n621 GND 0.013066f
C787 CS_BIAS.n622 GND 0.013132f
C788 CS_BIAS.n623 GND 0.007046f
C789 CS_BIAS.n624 GND 0.007046f
C790 CS_BIAS.n625 GND 0.007046f
C791 CS_BIAS.n626 GND 0.013132f
C792 CS_BIAS.n627 GND 0.073127f
C793 CS_BIAS.n628 GND 0.013132f
C794 CS_BIAS.n629 GND 0.007046f
C795 CS_BIAS.n630 GND 0.007046f
C796 CS_BIAS.n631 GND 0.007046f
C797 CS_BIAS.n632 GND 0.013132f
C798 CS_BIAS.n633 GND 0.013066f
C799 CS_BIAS.n634 GND 0.006465f
C800 CS_BIAS.n635 GND 0.007046f
C801 CS_BIAS.n636 GND 0.007046f
C802 CS_BIAS.n637 GND 0.007046f
C803 CS_BIAS.n638 GND 0.013132f
C804 CS_BIAS.n639 GND 0.013132f
C805 CS_BIAS.n640 GND 0.010798f
C806 CS_BIAS.n641 GND 0.007046f
C807 CS_BIAS.n642 GND 0.007046f
C808 CS_BIAS.n643 GND 0.008983f
C809 CS_BIAS.n644 GND 0.013132f
C810 CS_BIAS.n645 GND 0.013132f
C811 CS_BIAS.n646 GND 0.007046f
C812 CS_BIAS.n647 GND 0.007046f
C813 CS_BIAS.n648 GND 0.007046f
C814 CS_BIAS.n649 GND 0.009893f
C815 CS_BIAS.n650 GND 0.010679f
C816 CS_BIAS.n651 GND 0.013132f
C817 CS_BIAS.n652 GND 0.007046f
C818 CS_BIAS.n653 GND 0.007046f
C819 CS_BIAS.n654 GND 0.007046f
C820 CS_BIAS.n655 GND 0.013132f
C821 CS_BIAS.n656 GND 0.008464f
C822 CS_BIAS.n657 GND 0.094465f
C823 CS_BIAS.n658 GND 0.056596f
C824 CS_BIAS.n659 GND 0.046396f
C825 CS_BIAS.n660 GND 0.013254f
C826 CS_BIAS.t42 GND 0.150431f
C827 CS_BIAS.n661 GND 0.013132f
C828 CS_BIAS.n662 GND 0.007046f
C829 CS_BIAS.n663 GND 0.013132f
C830 CS_BIAS.n664 GND 0.007046f
C831 CS_BIAS.t50 GND 0.150431f
C832 CS_BIAS.n665 GND 0.066478f
C833 CS_BIAS.n666 GND 0.007046f
C834 CS_BIAS.n667 GND 0.014173f
C835 CS_BIAS.n668 GND 0.007046f
C836 CS_BIAS.n669 GND 0.013132f
C837 CS_BIAS.n670 GND 0.007046f
C838 CS_BIAS.t69 GND 0.150431f
C839 CS_BIAS.n671 GND 0.013132f
C840 CS_BIAS.n672 GND 0.007046f
C841 CS_BIAS.n673 GND 0.014173f
C842 CS_BIAS.n674 GND 0.007046f
C843 CS_BIAS.t33 GND 0.150431f
C844 CS_BIAS.n675 GND 0.094199f
C845 CS_BIAS.t52 GND 0.245181f
C846 CS_BIAS.n676 GND 0.124966f
C847 CS_BIAS.n677 GND 0.096934f
C848 CS_BIAS.n678 GND 0.010798f
C849 CS_BIAS.n679 GND 0.013132f
C850 CS_BIAS.n680 GND 0.013132f
C851 CS_BIAS.n681 GND 0.007046f
C852 CS_BIAS.n682 GND 0.007046f
C853 CS_BIAS.n683 GND 0.007046f
C854 CS_BIAS.n684 GND 0.006465f
C855 CS_BIAS.n685 GND 0.013066f
C856 CS_BIAS.n686 GND 0.013132f
C857 CS_BIAS.n687 GND 0.007046f
C858 CS_BIAS.n688 GND 0.007046f
C859 CS_BIAS.n689 GND 0.007046f
C860 CS_BIAS.n690 GND 0.013132f
C861 CS_BIAS.n691 GND 0.073127f
C862 CS_BIAS.n692 GND 0.013132f
C863 CS_BIAS.n693 GND 0.007046f
C864 CS_BIAS.n694 GND 0.007046f
C865 CS_BIAS.n695 GND 0.007046f
C866 CS_BIAS.n696 GND 0.013132f
C867 CS_BIAS.n697 GND 0.013066f
C868 CS_BIAS.n698 GND 0.006465f
C869 CS_BIAS.n699 GND 0.007046f
C870 CS_BIAS.n700 GND 0.007046f
C871 CS_BIAS.n701 GND 0.007046f
C872 CS_BIAS.n702 GND 0.013132f
C873 CS_BIAS.n703 GND 0.013132f
C874 CS_BIAS.n704 GND 0.010798f
C875 CS_BIAS.n705 GND 0.007046f
C876 CS_BIAS.n706 GND 0.007046f
C877 CS_BIAS.n707 GND 0.008983f
C878 CS_BIAS.n708 GND 0.013132f
C879 CS_BIAS.n709 GND 0.013132f
C880 CS_BIAS.n710 GND 0.007046f
C881 CS_BIAS.n711 GND 0.007046f
C882 CS_BIAS.n712 GND 0.007046f
C883 CS_BIAS.n713 GND 0.009893f
C884 CS_BIAS.n714 GND 0.010679f
C885 CS_BIAS.n715 GND 0.013132f
C886 CS_BIAS.n716 GND 0.007046f
C887 CS_BIAS.n717 GND 0.007046f
C888 CS_BIAS.n718 GND 0.007046f
C889 CS_BIAS.n719 GND 0.013132f
C890 CS_BIAS.n720 GND 0.008464f
C891 CS_BIAS.n721 GND 0.094465f
C892 CS_BIAS.n722 GND 0.056596f
C893 CS_BIAS.n723 GND 0.046396f
C894 CS_BIAS.n724 GND 0.013254f
C895 CS_BIAS.t40 GND 0.150431f
C896 CS_BIAS.n725 GND 0.013132f
C897 CS_BIAS.n726 GND 0.007046f
C898 CS_BIAS.n727 GND 0.013132f
C899 CS_BIAS.n728 GND 0.007046f
C900 CS_BIAS.t43 GND 0.150431f
C901 CS_BIAS.n729 GND 0.066478f
C902 CS_BIAS.n730 GND 0.007046f
C903 CS_BIAS.n731 GND 0.014173f
C904 CS_BIAS.n732 GND 0.007046f
C905 CS_BIAS.n733 GND 0.013132f
C906 CS_BIAS.n734 GND 0.007046f
C907 CS_BIAS.t63 GND 0.150431f
C908 CS_BIAS.n735 GND 0.013132f
C909 CS_BIAS.n736 GND 0.007046f
C910 CS_BIAS.n737 GND 0.014173f
C911 CS_BIAS.n738 GND 0.007046f
C912 CS_BIAS.t28 GND 0.150431f
C913 CS_BIAS.n739 GND 0.094199f
C914 CS_BIAS.t44 GND 0.245181f
C915 CS_BIAS.n740 GND 0.124966f
C916 CS_BIAS.n741 GND 0.096934f
C917 CS_BIAS.n742 GND 0.010798f
C918 CS_BIAS.n743 GND 0.013132f
C919 CS_BIAS.n744 GND 0.013132f
C920 CS_BIAS.n745 GND 0.007046f
C921 CS_BIAS.n746 GND 0.007046f
C922 CS_BIAS.n747 GND 0.007046f
C923 CS_BIAS.n748 GND 0.006465f
C924 CS_BIAS.n749 GND 0.013066f
C925 CS_BIAS.n750 GND 0.013132f
C926 CS_BIAS.n751 GND 0.007046f
C927 CS_BIAS.n752 GND 0.007046f
C928 CS_BIAS.n753 GND 0.007046f
C929 CS_BIAS.n754 GND 0.013132f
C930 CS_BIAS.n755 GND 0.073127f
C931 CS_BIAS.n756 GND 0.013132f
C932 CS_BIAS.n757 GND 0.007046f
C933 CS_BIAS.n758 GND 0.007046f
C934 CS_BIAS.n759 GND 0.007046f
C935 CS_BIAS.n760 GND 0.013132f
C936 CS_BIAS.n761 GND 0.013066f
C937 CS_BIAS.n762 GND 0.006465f
C938 CS_BIAS.n763 GND 0.007046f
C939 CS_BIAS.n764 GND 0.007046f
C940 CS_BIAS.n765 GND 0.007046f
C941 CS_BIAS.n766 GND 0.013132f
C942 CS_BIAS.n767 GND 0.013132f
C943 CS_BIAS.n768 GND 0.010798f
C944 CS_BIAS.n769 GND 0.007046f
C945 CS_BIAS.n770 GND 0.007046f
C946 CS_BIAS.n771 GND 0.008983f
C947 CS_BIAS.n772 GND 0.013132f
C948 CS_BIAS.n773 GND 0.013132f
C949 CS_BIAS.n774 GND 0.007046f
C950 CS_BIAS.n775 GND 0.007046f
C951 CS_BIAS.n776 GND 0.007046f
C952 CS_BIAS.n777 GND 0.009893f
C953 CS_BIAS.n778 GND 0.010679f
C954 CS_BIAS.n779 GND 0.013132f
C955 CS_BIAS.n780 GND 0.007046f
C956 CS_BIAS.n781 GND 0.007046f
C957 CS_BIAS.n782 GND 0.007046f
C958 CS_BIAS.n783 GND 0.013132f
C959 CS_BIAS.n784 GND 0.008464f
C960 CS_BIAS.n785 GND 0.094465f
C961 CS_BIAS.n786 GND 0.056596f
C962 CS_BIAS.n787 GND 0.112226f
C963 CS_BIAS.n788 GND 5.64941f
C964 VP.t10 GND 1.45835f
C965 VP.n0 GND 0.602832f
C966 VP.n1 GND 0.015751f
C967 VP.n2 GND 0.029356f
C968 VP.n3 GND 0.015751f
C969 VP.n4 GND 0.020142f
C970 VP.n5 GND 0.015751f
C971 VP.n6 GND 0.029356f
C972 VP.n7 GND 0.015751f
C973 VP.n8 GND 0.016022f
C974 VP.n9 GND 0.015751f
C975 VP.n10 GND 0.029356f
C976 VP.n11 GND 0.015751f
C977 VP.n12 GND 0.015115f
C978 VP.n13 GND 0.015751f
C979 VP.n14 GND 0.029356f
C980 VP.n15 GND 0.015751f
C981 VP.t16 GND 1.45835f
C982 VP.n16 GND 0.536808f
C983 VP.n17 GND 0.015751f
C984 VP.n18 GND 0.029356f
C985 VP.n19 GND 0.015751f
C986 VP.n20 GND 0.015115f
C987 VP.n21 GND 0.015751f
C988 VP.n22 GND 0.029356f
C989 VP.n23 GND 0.015751f
C990 VP.t15 GND 1.45835f
C991 VP.n24 GND 0.610287f
C992 VP.t14 GND 1.94171f
C993 VP.n25 GND 0.878652f
C994 VP.n26 GND 0.122502f
C995 VP.n27 GND 0.028197f
C996 VP.n28 GND 0.029356f
C997 VP.n29 GND 0.029356f
C998 VP.n30 GND 0.015751f
C999 VP.n31 GND 0.015751f
C1000 VP.n32 GND 0.015751f
C1001 VP.n33 GND 0.029356f
C1002 VP.n34 GND 0.029356f
C1003 VP.n35 GND 0.028756f
C1004 VP.n36 GND 0.015751f
C1005 VP.n37 GND 0.015751f
C1006 VP.n38 GND 0.015751f
C1007 VP.n39 GND 0.031475f
C1008 VP.n40 GND 0.029356f
C1009 VP.n41 GND 0.029356f
C1010 VP.n42 GND 0.015751f
C1011 VP.n43 GND 0.015751f
C1012 VP.n44 GND 0.015751f
C1013 VP.n45 GND 0.029356f
C1014 VP.n46 GND 0.029356f
C1015 VP.n47 GND 0.02211f
C1016 VP.n48 GND 0.015751f
C1017 VP.n49 GND 0.015751f
C1018 VP.n50 GND 0.02211f
C1019 VP.n51 GND 0.029356f
C1020 VP.n52 GND 0.029356f
C1021 VP.n53 GND 0.015751f
C1022 VP.n54 GND 0.015751f
C1023 VP.n55 GND 0.015751f
C1024 VP.n56 GND 0.029356f
C1025 VP.n57 GND 0.029356f
C1026 VP.n58 GND 0.031475f
C1027 VP.n59 GND 0.015751f
C1028 VP.n60 GND 0.015751f
C1029 VP.n61 GND 0.015751f
C1030 VP.n62 GND 0.028756f
C1031 VP.n63 GND 0.029356f
C1032 VP.n64 GND 0.029356f
C1033 VP.n65 GND 0.015751f
C1034 VP.n66 GND 0.015751f
C1035 VP.n67 GND 0.015751f
C1036 VP.n68 GND 0.029356f
C1037 VP.n69 GND 0.029356f
C1038 VP.t11 GND 1.45835f
C1039 VP.n70 GND 0.536808f
C1040 VP.n71 GND 0.028197f
C1041 VP.n72 GND 0.015751f
C1042 VP.n73 GND 0.015751f
C1043 VP.n74 GND 0.015751f
C1044 VP.n75 GND 0.029356f
C1045 VP.n76 GND 0.029356f
C1046 VP.n77 GND 0.029356f
C1047 VP.n78 GND 0.015751f
C1048 VP.n79 GND 0.015751f
C1049 VP.n80 GND 0.015751f
C1050 VP.n81 GND 0.029356f
C1051 VP.n82 GND 0.029356f
C1052 VP.n83 GND 0.025848f
C1053 VP.n84 GND 0.015751f
C1054 VP.n85 GND 0.015751f
C1055 VP.n86 GND 0.015751f
C1056 VP.n87 GND 0.029356f
C1057 VP.n88 GND 0.029356f
C1058 VP.n89 GND 0.029356f
C1059 VP.n90 GND 0.015751f
C1060 VP.n91 GND 0.015751f
C1061 VP.n92 GND 0.015751f
C1062 VP.n93 GND 0.029356f
C1063 VP.n94 GND 0.029356f
C1064 VP.n95 GND 0.019791f
C1065 VP.n96 GND 0.03918f
C1066 VP.n97 GND 0.447141f
C1067 VP.t13 GND 1.45835f
C1068 VP.n98 GND 0.602832f
C1069 VP.n99 GND 0.015751f
C1070 VP.n100 GND 0.029356f
C1071 VP.n101 GND 0.015751f
C1072 VP.n102 GND 0.020142f
C1073 VP.n103 GND 0.015751f
C1074 VP.n104 GND 0.029356f
C1075 VP.n105 GND 0.015751f
C1076 VP.n106 GND 0.016022f
C1077 VP.n107 GND 0.015751f
C1078 VP.t8 GND 1.45835f
C1079 VP.n108 GND 0.536808f
C1080 VP.n109 GND 0.029356f
C1081 VP.n110 GND 0.015751f
C1082 VP.n111 GND 0.015115f
C1083 VP.n112 GND 0.015751f
C1084 VP.n113 GND 0.029356f
C1085 VP.n114 GND 0.015751f
C1086 VP.t9 GND 1.45835f
C1087 VP.n115 GND 0.536808f
C1088 VP.n116 GND 0.015751f
C1089 VP.n117 GND 0.029356f
C1090 VP.n118 GND 0.015751f
C1091 VP.n119 GND 0.015115f
C1092 VP.n120 GND 0.015751f
C1093 VP.n121 GND 0.029356f
C1094 VP.n122 GND 0.015751f
C1095 VP.t7 GND 1.45835f
C1096 VP.n123 GND 0.610287f
C1097 VP.t12 GND 1.94171f
C1098 VP.n124 GND 0.878655f
C1099 VP.n125 GND 0.122501f
C1100 VP.n126 GND 0.028197f
C1101 VP.n127 GND 0.029356f
C1102 VP.n128 GND 0.029356f
C1103 VP.n129 GND 0.015751f
C1104 VP.n130 GND 0.015751f
C1105 VP.n131 GND 0.015751f
C1106 VP.n132 GND 0.029356f
C1107 VP.n133 GND 0.029356f
C1108 VP.n134 GND 0.028756f
C1109 VP.n135 GND 0.015751f
C1110 VP.n136 GND 0.015751f
C1111 VP.n137 GND 0.015751f
C1112 VP.n138 GND 0.031475f
C1113 VP.n139 GND 0.029356f
C1114 VP.n140 GND 0.029356f
C1115 VP.n141 GND 0.015751f
C1116 VP.n142 GND 0.015751f
C1117 VP.n143 GND 0.015751f
C1118 VP.n144 GND 0.029356f
C1119 VP.n145 GND 0.029356f
C1120 VP.n146 GND 0.02211f
C1121 VP.n147 GND 0.015751f
C1122 VP.n148 GND 0.015751f
C1123 VP.n149 GND 0.02211f
C1124 VP.n150 GND 0.029356f
C1125 VP.n151 GND 0.029356f
C1126 VP.n152 GND 0.015751f
C1127 VP.n153 GND 0.015751f
C1128 VP.n154 GND 0.015751f
C1129 VP.n155 GND 0.029356f
C1130 VP.n156 GND 0.029356f
C1131 VP.n157 GND 0.031475f
C1132 VP.n158 GND 0.015751f
C1133 VP.n159 GND 0.015751f
C1134 VP.n160 GND 0.015751f
C1135 VP.n161 GND 0.028756f
C1136 VP.n162 GND 0.029356f
C1137 VP.n163 GND 0.029356f
C1138 VP.n164 GND 0.015751f
C1139 VP.n165 GND 0.015751f
C1140 VP.n166 GND 0.015751f
C1141 VP.n167 GND 0.029356f
C1142 VP.n168 GND 0.029356f
C1143 VP.n169 GND 0.028197f
C1144 VP.n170 GND 0.015751f
C1145 VP.n171 GND 0.015751f
C1146 VP.n172 GND 0.015751f
C1147 VP.n173 GND 0.029356f
C1148 VP.n174 GND 0.029356f
C1149 VP.n175 GND 0.029356f
C1150 VP.n176 GND 0.015751f
C1151 VP.n177 GND 0.015751f
C1152 VP.n178 GND 0.015751f
C1153 VP.n179 GND 0.029356f
C1154 VP.n180 GND 0.029356f
C1155 VP.n181 GND 0.025848f
C1156 VP.n182 GND 0.015751f
C1157 VP.n183 GND 0.015751f
C1158 VP.n184 GND 0.015751f
C1159 VP.n185 GND 0.029356f
C1160 VP.n186 GND 0.029356f
C1161 VP.n187 GND 0.029356f
C1162 VP.n188 GND 0.015751f
C1163 VP.n189 GND 0.015751f
C1164 VP.n190 GND 0.015751f
C1165 VP.n191 GND 0.029356f
C1166 VP.n192 GND 0.029356f
C1167 VP.n193 GND 0.019791f
C1168 VP.n194 GND 0.03918f
C1169 VP.n195 GND 1.37411f
C1170 VP.n196 GND 1.54429f
C1171 VP.t3 GND 0.004856f
C1172 VP.t0 GND 0.004856f
C1173 VP.n197 GND 0.015966f
C1174 VP.t4 GND 0.004856f
C1175 VP.t1 GND 0.004856f
C1176 VP.n198 GND 0.015748f
C1177 VP.n199 GND 0.134398f
C1178 VP.t6 GND 0.004856f
C1179 VP.t2 GND 0.004856f
C1180 VP.n200 GND 0.015748f
C1181 VP.n201 GND 0.066071f
C1182 VP.t5 GND 0.027026f
C1183 VP.n202 GND 0.07334f
C1184 VP.n203 GND 1.08403f
C1185 VN.t14 GND 1.05248f
C1186 VN.n0 GND 0.43506f
C1187 VN.n1 GND 0.011368f
C1188 VN.n2 GND 0.021186f
C1189 VN.n3 GND 0.011368f
C1190 VN.n4 GND 0.014537f
C1191 VN.n5 GND 0.011368f
C1192 VN.n6 GND 0.021186f
C1193 VN.n7 GND 0.011368f
C1194 VN.n8 GND 0.011563f
C1195 VN.n9 GND 0.011368f
C1196 VN.t10 GND 1.05248f
C1197 VN.n10 GND 0.387411f
C1198 VN.n11 GND 0.021186f
C1199 VN.n12 GND 0.011368f
C1200 VN.n13 GND 0.010909f
C1201 VN.n14 GND 0.011368f
C1202 VN.n15 GND 0.021186f
C1203 VN.n16 GND 0.011368f
C1204 VN.t11 GND 1.05248f
C1205 VN.n17 GND 0.387411f
C1206 VN.n18 GND 0.011368f
C1207 VN.n19 GND 0.021186f
C1208 VN.n20 GND 0.011368f
C1209 VN.n21 GND 0.010909f
C1210 VN.n22 GND 0.011368f
C1211 VN.n23 GND 0.021186f
C1212 VN.n24 GND 0.011368f
C1213 VN.t9 GND 1.05248f
C1214 VN.n25 GND 0.44044f
C1215 VN.t13 GND 1.40132f
C1216 VN.n26 GND 0.634119f
C1217 VN.n27 GND 0.088408f
C1218 VN.n28 GND 0.020349f
C1219 VN.n29 GND 0.021186f
C1220 VN.n30 GND 0.021186f
C1221 VN.n31 GND 0.011368f
C1222 VN.n32 GND 0.011368f
C1223 VN.n33 GND 0.011368f
C1224 VN.n34 GND 0.021186f
C1225 VN.n35 GND 0.021186f
C1226 VN.n36 GND 0.020753f
C1227 VN.n37 GND 0.011368f
C1228 VN.n38 GND 0.011368f
C1229 VN.n39 GND 0.011368f
C1230 VN.n40 GND 0.022715f
C1231 VN.n41 GND 0.021186f
C1232 VN.n42 GND 0.021186f
C1233 VN.n43 GND 0.011368f
C1234 VN.n44 GND 0.011368f
C1235 VN.n45 GND 0.011368f
C1236 VN.n46 GND 0.021186f
C1237 VN.n47 GND 0.021186f
C1238 VN.n48 GND 0.015956f
C1239 VN.n49 GND 0.011368f
C1240 VN.n50 GND 0.011368f
C1241 VN.n51 GND 0.015956f
C1242 VN.n52 GND 0.021186f
C1243 VN.n53 GND 0.021186f
C1244 VN.n54 GND 0.011368f
C1245 VN.n55 GND 0.011368f
C1246 VN.n56 GND 0.011368f
C1247 VN.n57 GND 0.021186f
C1248 VN.n58 GND 0.021186f
C1249 VN.n59 GND 0.022715f
C1250 VN.n60 GND 0.011368f
C1251 VN.n61 GND 0.011368f
C1252 VN.n62 GND 0.011368f
C1253 VN.n63 GND 0.020753f
C1254 VN.n64 GND 0.021186f
C1255 VN.n65 GND 0.021186f
C1256 VN.n66 GND 0.011368f
C1257 VN.n67 GND 0.011368f
C1258 VN.n68 GND 0.011368f
C1259 VN.n69 GND 0.021186f
C1260 VN.n70 GND 0.021186f
C1261 VN.n71 GND 0.020349f
C1262 VN.n72 GND 0.011368f
C1263 VN.n73 GND 0.011368f
C1264 VN.n74 GND 0.011368f
C1265 VN.n75 GND 0.021186f
C1266 VN.n76 GND 0.021186f
C1267 VN.n77 GND 0.021186f
C1268 VN.n78 GND 0.011368f
C1269 VN.n79 GND 0.011368f
C1270 VN.n80 GND 0.011368f
C1271 VN.n81 GND 0.021186f
C1272 VN.n82 GND 0.021186f
C1273 VN.n83 GND 0.018654f
C1274 VN.n84 GND 0.011368f
C1275 VN.n85 GND 0.011368f
C1276 VN.n86 GND 0.011368f
C1277 VN.n87 GND 0.021186f
C1278 VN.n88 GND 0.021186f
C1279 VN.n89 GND 0.021186f
C1280 VN.n90 GND 0.011368f
C1281 VN.n91 GND 0.011368f
C1282 VN.n92 GND 0.011368f
C1283 VN.n93 GND 0.021186f
C1284 VN.n94 GND 0.021186f
C1285 VN.n95 GND 0.014283f
C1286 VN.n96 GND 0.028276f
C1287 VN.n97 GND 0.319928f
C1288 VN.t7 GND 1.05248f
C1289 VN.n98 GND 0.43506f
C1290 VN.n99 GND 0.011368f
C1291 VN.n100 GND 0.021186f
C1292 VN.n101 GND 0.011368f
C1293 VN.n102 GND 0.014537f
C1294 VN.n103 GND 0.011368f
C1295 VN.n104 GND 0.021186f
C1296 VN.n105 GND 0.011368f
C1297 VN.n106 GND 0.011563f
C1298 VN.n107 GND 0.011368f
C1299 VN.n108 GND 0.021186f
C1300 VN.n109 GND 0.011368f
C1301 VN.n110 GND 0.010909f
C1302 VN.n111 GND 0.011368f
C1303 VN.n112 GND 0.021186f
C1304 VN.n113 GND 0.011368f
C1305 VN.t15 GND 1.05248f
C1306 VN.n114 GND 0.387411f
C1307 VN.n115 GND 0.011368f
C1308 VN.n116 GND 0.021186f
C1309 VN.n117 GND 0.011368f
C1310 VN.n118 GND 0.010909f
C1311 VN.n119 GND 0.011368f
C1312 VN.n120 GND 0.021186f
C1313 VN.n121 GND 0.011368f
C1314 VN.t16 GND 1.05248f
C1315 VN.n122 GND 0.44044f
C1316 VN.t12 GND 1.40132f
C1317 VN.n123 GND 0.634117f
C1318 VN.n124 GND 0.088408f
C1319 VN.n125 GND 0.020349f
C1320 VN.n126 GND 0.021186f
C1321 VN.n127 GND 0.021186f
C1322 VN.n128 GND 0.011368f
C1323 VN.n129 GND 0.011368f
C1324 VN.n130 GND 0.011368f
C1325 VN.n131 GND 0.021186f
C1326 VN.n132 GND 0.021186f
C1327 VN.n133 GND 0.020753f
C1328 VN.n134 GND 0.011368f
C1329 VN.n135 GND 0.011368f
C1330 VN.n136 GND 0.011368f
C1331 VN.n137 GND 0.022715f
C1332 VN.n138 GND 0.021186f
C1333 VN.n139 GND 0.021186f
C1334 VN.n140 GND 0.011368f
C1335 VN.n141 GND 0.011368f
C1336 VN.n142 GND 0.011368f
C1337 VN.n143 GND 0.021186f
C1338 VN.n144 GND 0.021186f
C1339 VN.n145 GND 0.015956f
C1340 VN.n146 GND 0.011368f
C1341 VN.n147 GND 0.011368f
C1342 VN.n148 GND 0.015956f
C1343 VN.n149 GND 0.021186f
C1344 VN.n150 GND 0.021186f
C1345 VN.n151 GND 0.011368f
C1346 VN.n152 GND 0.011368f
C1347 VN.n153 GND 0.011368f
C1348 VN.n154 GND 0.021186f
C1349 VN.n155 GND 0.021186f
C1350 VN.n156 GND 0.022715f
C1351 VN.n157 GND 0.011368f
C1352 VN.n158 GND 0.011368f
C1353 VN.n159 GND 0.011368f
C1354 VN.n160 GND 0.020753f
C1355 VN.n161 GND 0.021186f
C1356 VN.n162 GND 0.021186f
C1357 VN.n163 GND 0.011368f
C1358 VN.n164 GND 0.011368f
C1359 VN.n165 GND 0.011368f
C1360 VN.n166 GND 0.021186f
C1361 VN.n167 GND 0.021186f
C1362 VN.t8 GND 1.05248f
C1363 VN.n168 GND 0.387411f
C1364 VN.n169 GND 0.020349f
C1365 VN.n170 GND 0.011368f
C1366 VN.n171 GND 0.011368f
C1367 VN.n172 GND 0.011368f
C1368 VN.n173 GND 0.021186f
C1369 VN.n174 GND 0.021186f
C1370 VN.n175 GND 0.021186f
C1371 VN.n176 GND 0.011368f
C1372 VN.n177 GND 0.011368f
C1373 VN.n178 GND 0.011368f
C1374 VN.n179 GND 0.021186f
C1375 VN.n180 GND 0.021186f
C1376 VN.n181 GND 0.018654f
C1377 VN.n182 GND 0.011368f
C1378 VN.n183 GND 0.011368f
C1379 VN.n184 GND 0.011368f
C1380 VN.n185 GND 0.021186f
C1381 VN.n186 GND 0.021186f
C1382 VN.n187 GND 0.021186f
C1383 VN.n188 GND 0.011368f
C1384 VN.n189 GND 0.011368f
C1385 VN.n190 GND 0.011368f
C1386 VN.n191 GND 0.021186f
C1387 VN.n192 GND 0.021186f
C1388 VN.n193 GND 0.014283f
C1389 VN.n194 GND 0.028276f
C1390 VN.n195 GND 0.987316f
C1391 VN.n196 GND 1.10966f
C1392 VN.t1 GND 0.019623f
C1393 VN.t2 GND 0.003504f
C1394 VN.t0 GND 0.003504f
C1395 VN.n197 GND 0.011365f
C1396 VN.n198 GND 0.088227f
C1397 VN.t3 GND 0.003504f
C1398 VN.t5 GND 0.003504f
C1399 VN.n199 GND 0.011365f
C1400 VN.n200 GND 0.047683f
C1401 VN.t4 GND 0.003504f
C1402 VN.t6 GND 0.003504f
C1403 VN.n201 GND 0.011365f
C1404 VN.n202 GND 0.066225f
C1405 VN.n203 GND 3.26216f
C1406 a_n7261_9606.n0 GND 2.44118f
C1407 a_n7261_9606.t15 GND 0.11533f
C1408 a_n7261_9606.t17 GND 1.10633f
C1409 a_n7261_9606.t9 GND 1.10292f
C1410 a_n7261_9606.t8 GND 0.11533f
C1411 a_n7261_9606.t13 GND 0.11533f
C1412 a_n7261_9606.n1 GND 0.827588f
C1413 a_n7261_9606.n2 GND 5.13771f
C1414 a_n7261_9606.t12 GND 0.11533f
C1415 a_n7261_9606.t10 GND 0.11533f
C1416 a_n7261_9606.n3 GND 0.827588f
C1417 a_n7261_9606.n4 GND 8.48639f
C1418 a_n7261_9606.t7 GND 0.989554f
C1419 a_n7261_9606.t0 GND 0.11533f
C1420 a_n7261_9606.t3 GND 0.11533f
C1421 a_n7261_9606.n5 GND 0.713262f
C1422 a_n7261_9606.n6 GND 2.67084f
C1423 a_n7261_9606.t5 GND 0.969821f
C1424 a_n7261_9606.t1 GND 0.969821f
C1425 a_n7261_9606.t2 GND 0.11533f
C1426 a_n7261_9606.t4 GND 0.11533f
C1427 a_n7261_9606.n7 GND 0.713262f
C1428 a_n7261_9606.n8 GND 1.59824f
C1429 a_n7261_9606.t6 GND 0.969821f
C1430 a_n7261_9606.n9 GND 1.91816f
C1431 a_n7261_9606.n10 GND 4.3007f
C1432 a_n7261_9606.t14 GND 0.11533f
C1433 a_n7261_9606.t11 GND 0.11533f
C1434 a_n7261_9606.n11 GND 0.827584f
C1435 a_n7261_9606.n12 GND 3.45717f
C1436 a_n7261_9606.n13 GND 2.56052f
C1437 a_n7261_9606.n14 GND 0.827588f
C1438 a_n7261_9606.t16 GND 0.11533f
C1439 a_n7183_9410.n0 GND 8.4972f
C1440 a_n7183_9410.n1 GND 0.662914f
C1441 a_n7183_9410.n2 GND 1.09669f
C1442 a_n7183_9410.n3 GND 5.0631f
C1443 a_n7183_9410.n4 GND 0.665023f
C1444 a_n7183_9410.t11 GND 0.443346f
C1445 a_n7183_9410.t16 GND 0.443346f
C1446 a_n7183_9410.t9 GND 0.458003f
C1447 a_n7183_9410.t7 GND 0.443346f
C1448 a_n7183_9410.n5 GND 2.84854f
C1449 a_n7183_9410.n6 GND 0.664153f
C1450 a_n7183_9410.n7 GND 2.73806f
C1451 a_n7183_9410.n8 GND 0.664153f
C1452 a_n7183_9410.n9 GND 0.664834f
C1453 a_n7183_9410.n10 GND 2.84155f
C1454 a_n7183_9410.n11 GND 0.664153f
C1455 a_n7183_9410.n12 GND 0.662914f
C1456 a_n7183_9410.n13 GND 0.662914f
C1457 a_n7183_9410.n14 GND 7.74294f
C1458 a_n7183_9410.t2 GND 0.530793f
C1459 a_n7183_9410.t4 GND 0.500997f
C1460 a_n7183_9410.t5 GND 0.530792f
C1461 a_n7183_9410.t0 GND 0.500996f
C1462 a_n7183_9410.n15 GND 1.50646f
C1463 a_n7183_9410.n16 GND 0.653429f
C1464 a_n7183_9410.n17 GND 0.653429f
C1465 a_n7183_9410.n18 GND 0.653937f
C1466 a_n7183_9410.n19 GND 0.653937f
C1467 a_n7183_9410.n20 GND 0.653937f
C1468 a_n7183_9410.n21 GND 0.653429f
C1469 a_n7183_9410.n22 GND 2.85932f
C1470 a_n7183_9410.n23 GND 2.68598f
C1471 a_n7183_9410.n24 GND 0.206448f
C1472 a_n7183_9410.n25 GND 0.206448f
C1473 a_n7183_9410.n26 GND 0.206448f
C1474 a_n7183_9410.n27 GND 1.35001f
C1475 a_n7183_9410.n28 GND 6.09383f
C1476 a_n7183_9410.t14 GND 2.0904f
C1477 a_n7183_9410.t6 GND 2.05239f
C1478 a_n7183_9410.t13 GND 1.68385f
C1479 a_n7183_9410.n29 GND 0.865686f
C1480 a_n7183_9410.t10 GND 2.05321f
C1481 a_n7183_9410.t28 GND 2.09039f
C1482 a_n7183_9410.t44 GND 1.68385f
C1483 a_n7183_9410.n30 GND 0.842234f
C1484 a_n7183_9410.t35 GND 1.68385f
C1485 a_n7183_9410.n31 GND 0.847986f
C1486 a_n7183_9410.t25 GND 2.05646f
C1487 a_n7183_9410.t20 GND 0.455508f
C1488 a_n7183_9410.t19 GND 2.0904f
C1489 a_n7183_9410.t34 GND 2.0904f
C1490 a_n7183_9410.t37 GND 2.09039f
C1491 a_n7183_9410.t38 GND 1.68385f
C1492 a_n7183_9410.n32 GND 0.842234f
C1493 a_n7183_9410.t30 GND 1.68385f
C1494 a_n7183_9410.n33 GND 0.847986f
C1495 a_n7183_9410.t33 GND 2.05646f
C1496 a_n7183_9410.t12 GND 2.09039f
C1497 a_n7183_9410.t8 GND 1.68385f
C1498 a_n7183_9410.n34 GND 0.842234f
C1499 a_n7183_9410.t15 GND 1.68385f
C1500 a_n7183_9410.n35 GND 0.847986f
C1501 a_n7183_9410.t21 GND 2.05646f
C1502 a_n7183_9410.t24 GND 2.09142f
C1503 a_n7183_9410.t26 GND 2.09142f
C1504 a_n7183_9410.t32 GND 2.09142f
C1505 a_n7183_9410.t42 GND 2.09142f
C1506 a_n7183_9410.t40 GND 2.09141f
C1507 a_n7183_9410.t47 GND 1.68385f
C1508 a_n7183_9410.n36 GND 0.849629f
C1509 a_n7183_9410.t23 GND 2.06243f
C1510 a_n7183_9410.t46 GND 2.09141f
C1511 a_n7183_9410.t31 GND 1.68385f
C1512 a_n7183_9410.n37 GND 0.849629f
C1513 a_n7183_9410.t41 GND 2.06243f
C1514 a_n7183_9410.t22 GND 2.09141f
C1515 a_n7183_9410.t45 GND 2.09762f
C1516 a_n7183_9410.t29 GND 2.06452f
C1517 a_n7183_9410.t39 GND 2.09141f
C1518 a_n7183_9410.t36 GND 1.68385f
C1519 a_n7183_9410.n38 GND 0.849629f
C1520 a_n7183_9410.t27 GND 2.06243f
C1521 a_n7183_9410.t43 GND 2.0904f
C1522 a_n7183_9410.t17 GND 2.0904f
C1523 a_n7183_9410.t3 GND 0.536632f
C1524 a_n7183_9410.t1 GND 0.512728f
C1525 a_n7183_9410.t18 GND 0.464779f
C1526 VOUT.t61 GND 0.010105f
C1527 VOUT.t72 GND 0.010105f
C1528 VOUT.n0 GND 0.055666f
C1529 VOUT.t93 GND 0.010105f
C1530 VOUT.t57 GND 0.010105f
C1531 VOUT.n1 GND 0.0527f
C1532 VOUT.n2 GND 0.656054f
C1533 VOUT.t103 GND 0.010105f
C1534 VOUT.t68 GND 0.010105f
C1535 VOUT.n3 GND 0.0527f
C1536 VOUT.n4 GND 0.327136f
C1537 VOUT.t88 GND 0.010105f
C1538 VOUT.t96 GND 0.010105f
C1539 VOUT.n5 GND 0.0527f
C1540 VOUT.n6 GND 0.398256f
C1541 VOUT.t105 GND 0.010105f
C1542 VOUT.t50 GND 0.010105f
C1543 VOUT.n7 GND 0.055666f
C1544 VOUT.t75 GND 0.010105f
C1545 VOUT.t98 GND 0.010105f
C1546 VOUT.n8 GND 0.0527f
C1547 VOUT.n9 GND 0.656054f
C1548 VOUT.t84 GND 0.010105f
C1549 VOUT.t46 GND 0.010105f
C1550 VOUT.n10 GND 0.0527f
C1551 VOUT.n11 GND 0.327136f
C1552 VOUT.t69 GND 0.010105f
C1553 VOUT.t76 GND 0.010105f
C1554 VOUT.n12 GND 0.0527f
C1555 VOUT.n13 GND 0.38045f
C1556 VOUT.n14 GND 0.284621f
C1557 VOUT.t71 GND 0.010105f
C1558 VOUT.t44 GND 0.010105f
C1559 VOUT.n15 GND 0.055666f
C1560 VOUT.t85 GND 0.010105f
C1561 VOUT.t102 GND 0.010105f
C1562 VOUT.n16 GND 0.0527f
C1563 VOUT.n17 GND 0.656054f
C1564 VOUT.t106 GND 0.010105f
C1565 VOUT.t63 GND 0.010105f
C1566 VOUT.n18 GND 0.0527f
C1567 VOUT.n19 GND 0.327136f
C1568 VOUT.t99 GND 0.010105f
C1569 VOUT.t66 GND 0.010105f
C1570 VOUT.n20 GND 0.0527f
C1571 VOUT.n21 GND 0.38045f
C1572 VOUT.n22 GND 0.18878f
C1573 VOUT.t95 GND 0.010105f
C1574 VOUT.t70 GND 0.010105f
C1575 VOUT.n23 GND 0.055666f
C1576 VOUT.t47 GND 0.010105f
C1577 VOUT.t64 GND 0.010105f
C1578 VOUT.n24 GND 0.0527f
C1579 VOUT.n25 GND 0.656054f
C1580 VOUT.t65 GND 0.010105f
C1581 VOUT.t86 GND 0.010105f
C1582 VOUT.n26 GND 0.0527f
C1583 VOUT.n27 GND 0.327136f
C1584 VOUT.t60 GND 0.010105f
C1585 VOUT.t90 GND 0.010105f
C1586 VOUT.n28 GND 0.0527f
C1587 VOUT.n29 GND 0.38045f
C1588 VOUT.n30 GND 0.460831f
C1589 VOUT.n31 GND 8.741871f
C1590 VOUT.n32 GND 6.27947f
C1591 VOUT.n33 GND 4.9244f
C1592 VOUT.n34 GND 4.9244f
C1593 VOUT.t118 GND 17.1455f
C1594 VOUT.t121 GND 15.109599f
C1595 VOUT.t120 GND 15.109599f
C1596 VOUT.t114 GND 17.648699f
C1597 VOUT.n35 GND 10.9614f
C1598 VOUT.n36 GND 5.76356f
C1599 VOUT.n37 GND 4.9244f
C1600 VOUT.n38 GND 4.92797f
C1601 VOUT.n39 GND 5.48275f
C1602 VOUT.n40 GND 4.9244f
C1603 VOUT.n41 GND 5.22377f
C1604 VOUT.n42 GND 13.051701f
C1605 VOUT.t115 GND 17.1455f
C1606 VOUT.n43 GND 13.051701f
C1607 VOUT.n44 GND 5.22377f
C1608 VOUT.t117 GND 15.109599f
C1609 VOUT.n45 GND 5.48275f
C1610 VOUT.n46 GND 4.92797f
C1611 VOUT.t116 GND 15.109599f
C1612 VOUT.n47 GND 5.48275f
C1613 VOUT.n48 GND 4.92797f
C1614 VOUT.t119 GND 15.109599f
C1615 VOUT.n49 GND 6.93577f
C1616 VOUT.n50 GND 2.03402f
C1617 VOUT.t80 GND 0.010105f
C1618 VOUT.t73 GND 0.010105f
C1619 VOUT.n51 GND 0.055666f
C1620 VOUT.t45 GND 0.010105f
C1621 VOUT.t100 GND 0.010105f
C1622 VOUT.n52 GND 0.0527f
C1623 VOUT.n53 GND 0.656054f
C1624 VOUT.t74 GND 0.010105f
C1625 VOUT.t62 GND 0.010105f
C1626 VOUT.n54 GND 0.0527f
C1627 VOUT.n55 GND 0.327136f
C1628 VOUT.t59 GND 0.010105f
C1629 VOUT.t97 GND 0.010105f
C1630 VOUT.n56 GND 0.0527f
C1631 VOUT.n57 GND 0.398256f
C1632 VOUT.t58 GND 0.010105f
C1633 VOUT.t52 GND 0.010105f
C1634 VOUT.n58 GND 0.055666f
C1635 VOUT.t89 GND 0.010105f
C1636 VOUT.t81 GND 0.010105f
C1637 VOUT.n59 GND 0.0527f
C1638 VOUT.n60 GND 0.656054f
C1639 VOUT.t54 GND 0.010105f
C1640 VOUT.t107 GND 0.010105f
C1641 VOUT.n61 GND 0.0527f
C1642 VOUT.n62 GND 0.327136f
C1643 VOUT.t101 GND 0.010105f
C1644 VOUT.t78 GND 0.010105f
C1645 VOUT.n63 GND 0.0527f
C1646 VOUT.n64 GND 0.38045f
C1647 VOUT.n65 GND 0.284621f
C1648 VOUT.t83 GND 0.010105f
C1649 VOUT.t49 GND 0.010105f
C1650 VOUT.n66 GND 0.055666f
C1651 VOUT.t92 GND 0.010105f
C1652 VOUT.t53 GND 0.010105f
C1653 VOUT.n67 GND 0.0527f
C1654 VOUT.n68 GND 0.656054f
C1655 VOUT.t94 GND 0.010105f
C1656 VOUT.t56 GND 0.010105f
C1657 VOUT.n69 GND 0.0527f
C1658 VOUT.n70 GND 0.327136f
C1659 VOUT.t87 GND 0.010105f
C1660 VOUT.t67 GND 0.010105f
C1661 VOUT.n71 GND 0.0527f
C1662 VOUT.n72 GND 0.38045f
C1663 VOUT.n73 GND 0.18878f
C1664 VOUT.t104 GND 0.010105f
C1665 VOUT.t77 GND 0.010105f
C1666 VOUT.n74 GND 0.055666f
C1667 VOUT.t51 GND 0.010105f
C1668 VOUT.t79 GND 0.010105f
C1669 VOUT.n75 GND 0.0527f
C1670 VOUT.n76 GND 0.656054f
C1671 VOUT.t55 GND 0.010105f
C1672 VOUT.t82 GND 0.010105f
C1673 VOUT.n77 GND 0.0527f
C1674 VOUT.n78 GND 0.327136f
C1675 VOUT.t48 GND 0.010105f
C1676 VOUT.t91 GND 0.010105f
C1677 VOUT.n79 GND 0.0527f
C1678 VOUT.n80 GND 0.38045f
C1679 VOUT.n81 GND 0.460831f
C1680 VOUT.n82 GND 10.9058f
C1681 VOUT.n83 GND 0.00872f
C1682 VOUT.n84 GND 0.019253f
C1683 VOUT.t14 GND 0.014431f
C1684 VOUT.n85 GND 0.015105f
C1685 VOUT.n86 GND 0.004801f
C1686 VOUT.n87 GND 0.003167f
C1687 VOUT.n88 GND 0.042671f
C1688 VOUT.n89 GND 0.02312f
C1689 VOUT.t15 GND 0.009453f
C1690 VOUT.t33 GND 0.009453f
C1691 VOUT.n90 GND 0.066953f
C1692 VOUT.n91 GND 0.531776f
C1693 VOUT.t108 GND 0.009453f
C1694 VOUT.t26 GND 0.009453f
C1695 VOUT.n92 GND 0.066953f
C1696 VOUT.n93 GND 0.426527f
C1697 VOUT.n94 GND 0.00872f
C1698 VOUT.n95 GND 0.019253f
C1699 VOUT.t36 GND 0.014431f
C1700 VOUT.n96 GND 0.015105f
C1701 VOUT.n97 GND 0.004801f
C1702 VOUT.n98 GND 0.003167f
C1703 VOUT.n99 GND 0.042671f
C1704 VOUT.n100 GND 0.02312f
C1705 VOUT.t23 GND 0.009453f
C1706 VOUT.t37 GND 0.009453f
C1707 VOUT.n101 GND 0.066953f
C1708 VOUT.n102 GND 0.531776f
C1709 VOUT.t12 GND 0.009453f
C1710 VOUT.t42 GND 0.009453f
C1711 VOUT.n103 GND 0.066953f
C1712 VOUT.n104 GND 0.409043f
C1713 VOUT.n105 GND 0.289969f
C1714 VOUT.n106 GND 0.00872f
C1715 VOUT.n107 GND 0.019253f
C1716 VOUT.t1 GND 0.014431f
C1717 VOUT.n108 GND 0.015105f
C1718 VOUT.n109 GND 0.004801f
C1719 VOUT.n110 GND 0.003167f
C1720 VOUT.n111 GND 0.042671f
C1721 VOUT.n112 GND 0.02312f
C1722 VOUT.t32 GND 0.009453f
C1723 VOUT.t28 GND 0.009453f
C1724 VOUT.n113 GND 0.066953f
C1725 VOUT.n114 GND 0.531776f
C1726 VOUT.t2 GND 0.009453f
C1727 VOUT.t4 GND 0.009453f
C1728 VOUT.n115 GND 0.066953f
C1729 VOUT.n116 GND 0.409043f
C1730 VOUT.n117 GND 0.190147f
C1731 VOUT.n118 GND 0.00872f
C1732 VOUT.n119 GND 0.019253f
C1733 VOUT.t5 GND 0.014431f
C1734 VOUT.n120 GND 0.015105f
C1735 VOUT.n121 GND 0.004801f
C1736 VOUT.n122 GND 0.003167f
C1737 VOUT.n123 GND 0.042671f
C1738 VOUT.n124 GND 0.02312f
C1739 VOUT.t17 GND 0.009453f
C1740 VOUT.t19 GND 0.009453f
C1741 VOUT.n125 GND 0.066953f
C1742 VOUT.n126 GND 0.531776f
C1743 VOUT.t31 GND 0.009453f
C1744 VOUT.t43 GND 0.009453f
C1745 VOUT.n127 GND 0.066953f
C1746 VOUT.n128 GND 0.409043f
C1747 VOUT.n129 GND 0.190147f
C1748 VOUT.n130 GND 0.00872f
C1749 VOUT.n131 GND 0.019253f
C1750 VOUT.t11 GND 0.014431f
C1751 VOUT.n132 GND 0.015105f
C1752 VOUT.n133 GND 0.004801f
C1753 VOUT.n134 GND 0.003167f
C1754 VOUT.n135 GND 0.042671f
C1755 VOUT.n136 GND 0.02312f
C1756 VOUT.t40 GND 0.009453f
C1757 VOUT.t24 GND 0.009453f
C1758 VOUT.n137 GND 0.066953f
C1759 VOUT.n138 GND 0.531776f
C1760 VOUT.t110 GND 0.009453f
C1761 VOUT.t27 GND 0.009453f
C1762 VOUT.n139 GND 0.066953f
C1763 VOUT.n140 GND 0.409043f
C1764 VOUT.n141 GND 0.39453f
C1765 VOUT.n142 GND 10.8347f
C1766 VOUT.t20 GND 0.009453f
C1767 VOUT.t22 GND 0.009453f
C1768 VOUT.n143 GND 0.07328f
C1769 VOUT.t3 GND 0.009453f
C1770 VOUT.t7 GND 0.009453f
C1771 VOUT.n144 GND 0.066953f
C1772 VOUT.n145 GND 0.721779f
C1773 VOUT.n146 GND 0.00872f
C1774 VOUT.n147 GND 0.019253f
C1775 VOUT.t10 GND 0.014431f
C1776 VOUT.n148 GND 0.015105f
C1777 VOUT.n149 GND 0.004801f
C1778 VOUT.n150 GND 0.003167f
C1779 VOUT.n151 GND 0.042671f
C1780 VOUT.n152 GND 0.017728f
C1781 VOUT.n153 GND 0.260405f
C1782 VOUT.t112 GND 0.009453f
C1783 VOUT.t41 GND 0.009453f
C1784 VOUT.n154 GND 0.07328f
C1785 VOUT.t38 GND 0.009453f
C1786 VOUT.t0 GND 0.009453f
C1787 VOUT.n155 GND 0.066953f
C1788 VOUT.n156 GND 0.721779f
C1789 VOUT.n157 GND 0.00872f
C1790 VOUT.n158 GND 0.019253f
C1791 VOUT.t21 GND 0.014431f
C1792 VOUT.n159 GND 0.015105f
C1793 VOUT.n160 GND 0.004801f
C1794 VOUT.n161 GND 0.003167f
C1795 VOUT.n162 GND 0.042671f
C1796 VOUT.n163 GND 0.017728f
C1797 VOUT.n164 GND 0.244518f
C1798 VOUT.n165 GND 0.238739f
C1799 VOUT.t34 GND 0.009453f
C1800 VOUT.t9 GND 0.009453f
C1801 VOUT.n166 GND 0.07328f
C1802 VOUT.t109 GND 0.009453f
C1803 VOUT.t16 GND 0.009453f
C1804 VOUT.n167 GND 0.066953f
C1805 VOUT.n168 GND 0.721779f
C1806 VOUT.n169 GND 0.00872f
C1807 VOUT.n170 GND 0.019253f
C1808 VOUT.t8 GND 0.014431f
C1809 VOUT.n171 GND 0.015105f
C1810 VOUT.n172 GND 0.004801f
C1811 VOUT.n173 GND 0.003167f
C1812 VOUT.n174 GND 0.042671f
C1813 VOUT.n175 GND 0.017728f
C1814 VOUT.n176 GND 0.244518f
C1815 VOUT.n177 GND 0.163733f
C1816 VOUT.t18 GND 0.009453f
C1817 VOUT.t111 GND 0.009453f
C1818 VOUT.n178 GND 0.07328f
C1819 VOUT.t35 GND 0.009453f
C1820 VOUT.t6 GND 0.009453f
C1821 VOUT.n179 GND 0.066953f
C1822 VOUT.n180 GND 0.721779f
C1823 VOUT.n181 GND 0.00872f
C1824 VOUT.n182 GND 0.019253f
C1825 VOUT.t30 GND 0.014431f
C1826 VOUT.n183 GND 0.015105f
C1827 VOUT.n184 GND 0.004801f
C1828 VOUT.n185 GND 0.003167f
C1829 VOUT.n186 GND 0.042671f
C1830 VOUT.n187 GND 0.017728f
C1831 VOUT.n188 GND 0.244518f
C1832 VOUT.n189 GND 0.163733f
C1833 VOUT.t113 GND 0.009453f
C1834 VOUT.t29 GND 0.009453f
C1835 VOUT.n190 GND 0.07328f
C1836 VOUT.t39 GND 0.009453f
C1837 VOUT.t13 GND 0.009453f
C1838 VOUT.n191 GND 0.066953f
C1839 VOUT.n192 GND 0.721779f
C1840 VOUT.n193 GND 0.00872f
C1841 VOUT.n194 GND 0.019253f
C1842 VOUT.t25 GND 0.014431f
C1843 VOUT.n195 GND 0.015105f
C1844 VOUT.n196 GND 0.004801f
C1845 VOUT.n197 GND 0.003167f
C1846 VOUT.n198 GND 0.042671f
C1847 VOUT.n199 GND 0.017728f
C1848 VOUT.n200 GND 0.244518f
C1849 VOUT.n201 GND 0.368116f
C1850 VOUT.n202 GND 8.042621f
C1851 VOUT.n203 GND 5.08486f
C1852 VDD.t92 GND 0.017183f
C1853 VDD.t89 GND 0.017183f
C1854 VDD.n0 GND 0.126722f
C1855 VDD.t99 GND 0.017183f
C1856 VDD.t103 GND 0.017183f
C1857 VDD.n1 GND 0.123303f
C1858 VDD.n2 GND 0.482232f
C1859 VDD.t87 GND 0.017183f
C1860 VDD.t106 GND 0.017183f
C1861 VDD.n3 GND 0.123303f
C1862 VDD.n4 GND 0.25238f
C1863 VDD.t94 GND 0.017183f
C1864 VDD.t112 GND 0.017183f
C1865 VDD.n5 GND 0.123303f
C1866 VDD.n6 GND 0.211637f
C1867 VDD.t203 GND 0.017183f
C1868 VDD.t115 GND 0.017183f
C1869 VDD.n7 GND 0.126722f
C1870 VDD.t85 GND 0.017183f
C1871 VDD.t199 GND 0.017183f
C1872 VDD.n8 GND 0.123303f
C1873 VDD.n9 GND 0.482232f
C1874 VDD.t2 GND 0.017183f
C1875 VDD.t201 GND 0.017183f
C1876 VDD.n10 GND 0.123303f
C1877 VDD.n11 GND 0.25238f
C1878 VDD.t97 GND 0.017183f
C1879 VDD.t110 GND 0.017183f
C1880 VDD.n12 GND 0.123303f
C1881 VDD.n13 GND 0.211637f
C1882 VDD.n14 GND 0.16077f
C1883 VDD.n15 GND 2.87462f
C1884 VDD.t171 GND 0.044552f
C1885 VDD.t162 GND 0.006779f
C1886 VDD.t121 GND 0.006779f
C1887 VDD.n16 GND 0.028116f
C1888 VDD.n17 GND 0.353268f
C1889 VDD.t190 GND 0.006779f
C1890 VDD.t167 GND 0.006779f
C1891 VDD.n18 GND 0.028116f
C1892 VDD.n19 GND 0.217723f
C1893 VDD.t151 GND 0.006779f
C1894 VDD.t146 GND 0.006779f
C1895 VDD.n20 GND 0.028116f
C1896 VDD.n21 GND 0.217723f
C1897 VDD.t187 GND 0.043241f
C1898 VDD.n22 GND 0.17012f
C1899 VDD.t145 GND 0.044552f
C1900 VDD.t134 GND 0.006779f
C1901 VDD.t179 GND 0.006779f
C1902 VDD.n23 GND 0.028116f
C1903 VDD.n24 GND 0.353268f
C1904 VDD.t172 GND 0.006779f
C1905 VDD.t138 GND 0.006779f
C1906 VDD.n25 GND 0.028116f
C1907 VDD.n26 GND 0.217723f
C1908 VDD.t197 GND 0.006779f
C1909 VDD.t191 GND 0.006779f
C1910 VDD.n27 GND 0.028116f
C1911 VDD.n28 GND 0.217723f
C1912 VDD.t169 GND 0.043241f
C1913 VDD.n29 GND 0.158808f
C1914 VDD.n30 GND 0.160142f
C1915 VDD.t174 GND 0.044552f
C1916 VDD.t131 GND 0.006779f
C1917 VDD.t181 GND 0.006779f
C1918 VDD.n31 GND 0.028116f
C1919 VDD.n32 GND 0.353268f
C1920 VDD.t136 GND 0.006779f
C1921 VDD.t184 GND 0.006779f
C1922 VDD.n33 GND 0.028116f
C1923 VDD.n34 GND 0.217723f
C1924 VDD.t141 GND 0.006779f
C1925 VDD.t177 GND 0.006779f
C1926 VDD.n35 GND 0.028116f
C1927 VDD.n36 GND 0.217723f
C1928 VDD.t159 GND 0.043241f
C1929 VDD.n37 GND 0.158808f
C1930 VDD.n38 GND 0.11093f
C1931 VDD.t194 GND 0.044552f
C1932 VDD.t128 GND 0.006779f
C1933 VDD.t133 GND 0.006779f
C1934 VDD.n39 GND 0.028116f
C1935 VDD.n40 GND 0.353268f
C1936 VDD.t170 GND 0.006779f
C1937 VDD.t139 GND 0.006779f
C1938 VDD.n41 GND 0.028116f
C1939 VDD.n42 GND 0.217723f
C1940 VDD.t173 GND 0.006779f
C1941 VDD.t130 GND 0.006779f
C1942 VDD.n43 GND 0.028116f
C1943 VDD.n44 GND 0.217723f
C1944 VDD.t182 GND 0.043241f
C1945 VDD.n45 GND 0.158808f
C1946 VDD.n46 GND 0.308941f
C1947 VDD.n47 GND 0.007736f
C1948 VDD.n48 GND 0.007736f
C1949 VDD.n49 GND 0.006248f
C1950 VDD.n50 GND 0.006248f
C1951 VDD.n51 GND 0.007763f
C1952 VDD.n52 GND 0.007763f
C1953 VDD.n53 GND 0.594542f
C1954 VDD.n54 GND 0.007763f
C1955 VDD.n55 GND 0.007763f
C1956 VDD.n56 GND 0.007763f
C1957 VDD.n57 GND 0.588597f
C1958 VDD.n58 GND 0.007763f
C1959 VDD.n59 GND 0.007763f
C1960 VDD.n60 GND 0.007763f
C1961 VDD.n61 GND 0.007763f
C1962 VDD.n62 GND 0.006248f
C1963 VDD.n63 GND 0.007763f
C1964 VDD.t137 GND 0.297271f
C1965 VDD.n64 GND 0.007763f
C1966 VDD.n65 GND 0.007763f
C1967 VDD.n66 GND 0.007763f
C1968 VDD.n67 GND 0.594542f
C1969 VDD.n68 GND 0.007763f
C1970 VDD.n69 GND 0.007763f
C1971 VDD.n70 GND 0.007763f
C1972 VDD.n71 GND 0.007763f
C1973 VDD.n72 GND 0.007763f
C1974 VDD.n73 GND 0.006248f
C1975 VDD.n74 GND 0.007763f
C1976 VDD.n75 GND 0.007763f
C1977 VDD.n76 GND 0.007763f
C1978 VDD.n77 GND 0.007763f
C1979 VDD.n78 GND 0.576706f
C1980 VDD.n79 GND 0.007763f
C1981 VDD.n80 GND 0.007763f
C1982 VDD.n81 GND 0.007763f
C1983 VDD.n82 GND 0.007763f
C1984 VDD.n83 GND 0.007763f
C1985 VDD.n84 GND 0.006248f
C1986 VDD.n85 GND 0.007763f
C1987 VDD.t140 GND 0.297271f
C1988 VDD.n86 GND 0.007763f
C1989 VDD.n87 GND 0.007763f
C1990 VDD.n88 GND 0.007763f
C1991 VDD.n89 GND 0.594542f
C1992 VDD.n90 GND 0.007763f
C1993 VDD.n91 GND 0.007763f
C1994 VDD.n92 GND 0.007763f
C1995 VDD.n93 GND 0.007763f
C1996 VDD.n94 GND 0.007763f
C1997 VDD.n95 GND 0.006248f
C1998 VDD.n96 GND 0.007763f
C1999 VDD.n97 GND 0.007763f
C2000 VDD.n98 GND 0.007763f
C2001 VDD.n99 GND 0.007763f
C2002 VDD.n100 GND 0.564815f
C2003 VDD.n101 GND 0.007763f
C2004 VDD.n102 GND 0.007763f
C2005 VDD.n103 GND 0.007763f
C2006 VDD.n104 GND 0.007763f
C2007 VDD.n105 GND 0.007763f
C2008 VDD.n106 GND 0.006248f
C2009 VDD.n107 GND 0.007763f
C2010 VDD.t129 GND 0.297271f
C2011 VDD.n108 GND 0.007763f
C2012 VDD.n109 GND 0.007763f
C2013 VDD.n110 GND 0.007763f
C2014 VDD.n111 GND 0.594542f
C2015 VDD.n112 GND 0.007763f
C2016 VDD.n113 GND 0.007763f
C2017 VDD.n114 GND 0.007763f
C2018 VDD.n115 GND 0.007763f
C2019 VDD.n116 GND 0.007763f
C2020 VDD.n117 GND 0.006248f
C2021 VDD.n118 GND 0.007763f
C2022 VDD.n119 GND 0.007763f
C2023 VDD.n120 GND 0.007763f
C2024 VDD.n121 GND 0.007763f
C2025 VDD.n122 GND 0.552924f
C2026 VDD.n123 GND 0.007763f
C2027 VDD.n124 GND 0.007763f
C2028 VDD.n125 GND 0.007763f
C2029 VDD.n126 GND 0.007763f
C2030 VDD.n127 GND 0.007763f
C2031 VDD.n128 GND 0.006248f
C2032 VDD.n129 GND 0.007763f
C2033 VDD.t158 GND 0.297271f
C2034 VDD.n130 GND 0.007763f
C2035 VDD.n131 GND 0.007763f
C2036 VDD.n132 GND 0.007763f
C2037 VDD.n133 GND 0.594542f
C2038 VDD.n134 GND 0.007763f
C2039 VDD.n135 GND 0.007763f
C2040 VDD.n136 GND 0.007763f
C2041 VDD.n137 GND 0.007763f
C2042 VDD.n138 GND 0.007763f
C2043 VDD.n139 GND 0.006248f
C2044 VDD.n140 GND 0.007763f
C2045 VDD.n141 GND 0.007763f
C2046 VDD.n142 GND 0.007763f
C2047 VDD.n143 GND 0.007763f
C2048 VDD.n144 GND 0.594542f
C2049 VDD.n145 GND 0.007763f
C2050 VDD.n146 GND 0.007763f
C2051 VDD.n147 GND 0.007763f
C2052 VDD.n148 GND 0.007763f
C2053 VDD.n149 GND 0.007763f
C2054 VDD.n150 GND 0.006248f
C2055 VDD.n151 GND 0.007763f
C2056 VDD.n152 GND 0.007763f
C2057 VDD.n153 GND 0.007763f
C2058 VDD.n154 GND 0.007763f
C2059 VDD.n155 GND 0.594542f
C2060 VDD.n156 GND 0.007763f
C2061 VDD.n157 GND 0.007763f
C2062 VDD.n158 GND 0.007763f
C2063 VDD.n159 GND 0.007763f
C2064 VDD.n160 GND 0.007763f
C2065 VDD.n161 GND 0.006248f
C2066 VDD.n162 GND 0.007763f
C2067 VDD.n163 GND 0.007763f
C2068 VDD.n164 GND 0.007763f
C2069 VDD.n165 GND 0.018791f
C2070 VDD.n166 GND 1.39123f
C2071 VDD.n167 GND 0.019093f
C2072 VDD.n168 GND 0.007763f
C2073 VDD.n169 GND 0.007763f
C2074 VDD.n170 GND 0.007763f
C2075 VDD.n171 GND 0.007763f
C2076 VDD.n172 GND 0.006248f
C2077 VDD.n174 GND 0.007763f
C2078 VDD.n175 GND 0.007763f
C2079 VDD.n176 GND 0.007763f
C2080 VDD.n177 GND 0.007763f
C2081 VDD.n178 GND 0.007763f
C2082 VDD.t26 GND 0.035989f
C2083 VDD.t25 GND 0.048603f
C2084 VDD.t23 GND 0.295093f
C2085 VDD.n179 GND 0.062024f
C2086 VDD.n180 GND 0.044734f
C2087 VDD.n181 GND 0.012747f
C2088 VDD.n183 GND 0.007763f
C2089 VDD.n184 GND 0.007763f
C2090 VDD.n185 GND 0.007763f
C2091 VDD.n186 GND 0.007763f
C2092 VDD.n187 GND 0.007763f
C2093 VDD.n188 GND 0.006248f
C2094 VDD.n190 GND 0.007763f
C2095 VDD.n191 GND 0.007763f
C2096 VDD.n192 GND 0.007763f
C2097 VDD.n193 GND 0.007763f
C2098 VDD.n194 GND 0.007763f
C2099 VDD.n195 GND 0.006248f
C2100 VDD.n197 GND 0.007763f
C2101 VDD.n198 GND 0.007763f
C2102 VDD.n199 GND 0.007763f
C2103 VDD.n200 GND 0.007763f
C2104 VDD.n201 GND 0.007763f
C2105 VDD.n202 GND 0.006248f
C2106 VDD.n204 GND 0.007763f
C2107 VDD.n205 GND 0.007763f
C2108 VDD.n206 GND 0.007763f
C2109 VDD.n207 GND 0.007763f
C2110 VDD.n208 GND 0.007763f
C2111 VDD.n209 GND 0.006248f
C2112 VDD.n211 GND 0.007763f
C2113 VDD.n212 GND 0.007763f
C2114 VDD.n213 GND 0.007763f
C2115 VDD.n214 GND 0.007763f
C2116 VDD.n215 GND 0.007763f
C2117 VDD.n216 GND 0.00328f
C2118 VDD.n218 GND 0.007763f
C2119 VDD.t80 GND 0.035989f
C2120 VDD.t79 GND 0.048603f
C2121 VDD.t78 GND 0.295093f
C2122 VDD.n219 GND 0.062024f
C2123 VDD.n220 GND 0.044734f
C2124 VDD.n221 GND 0.009623f
C2125 VDD.n222 GND 0.007763f
C2126 VDD.n223 GND 0.007763f
C2127 VDD.n224 GND 0.007763f
C2128 VDD.n225 GND 0.007763f
C2129 VDD.n226 GND 0.006248f
C2130 VDD.n228 GND 0.007763f
C2131 VDD.n229 GND 0.007763f
C2132 VDD.n230 GND 0.007763f
C2133 VDD.n231 GND 0.007763f
C2134 VDD.n232 GND 0.007763f
C2135 VDD.n233 GND 0.006248f
C2136 VDD.n235 GND 0.007763f
C2137 VDD.n236 GND 0.007763f
C2138 VDD.n237 GND 0.007763f
C2139 VDD.n238 GND 0.007763f
C2140 VDD.n239 GND 0.007763f
C2141 VDD.n240 GND 0.007763f
C2142 VDD.n241 GND 0.006248f
C2143 VDD.n242 GND 0.007763f
C2144 VDD.n243 GND 0.007763f
C2145 VDD.n244 GND 0.006248f
C2146 VDD.n245 GND 0.007763f
C2147 VDD.n246 GND 0.007763f
C2148 VDD.n247 GND 0.006248f
C2149 VDD.n248 GND 0.007763f
C2150 VDD.n249 GND 0.007763f
C2151 VDD.n250 GND 0.006248f
C2152 VDD.n251 GND 0.007763f
C2153 VDD.n252 GND 0.007763f
C2154 VDD.n253 GND 0.006248f
C2155 VDD.n254 GND 0.007763f
C2156 VDD.n255 GND 0.007763f
C2157 VDD.n256 GND 0.006248f
C2158 VDD.n257 GND 0.007763f
C2159 VDD.n258 GND 0.007763f
C2160 VDD.n259 GND 0.006248f
C2161 VDD.n260 GND 0.007763f
C2162 VDD.n261 GND 0.007763f
C2163 VDD.n262 GND 0.006248f
C2164 VDD.n263 GND 0.007763f
C2165 VDD.n264 GND 0.007763f
C2166 VDD.n265 GND 0.006248f
C2167 VDD.n266 GND 0.007763f
C2168 VDD.n267 GND 0.007763f
C2169 VDD.n268 GND 0.006248f
C2170 VDD.n269 GND 0.007763f
C2171 VDD.n270 GND 0.006248f
C2172 VDD.n271 GND 0.007763f
C2173 VDD.n272 GND 0.006248f
C2174 VDD.n273 GND 0.007763f
C2175 VDD.n274 GND 0.007763f
C2176 VDD.n275 GND 0.588597f
C2177 VDD.n276 GND 0.007763f
C2178 VDD.n277 GND 0.006248f
C2179 VDD.n278 GND 0.007763f
C2180 VDD.n279 GND 0.006248f
C2181 VDD.n280 GND 0.007763f
C2182 VDD.n281 GND 0.594542f
C2183 VDD.n282 GND 0.007763f
C2184 VDD.n283 GND 0.006248f
C2185 VDD.n284 GND 0.007763f
C2186 VDD.n285 GND 0.006248f
C2187 VDD.n286 GND 0.007763f
C2188 VDD.n287 GND 0.594542f
C2189 VDD.n288 GND 0.007763f
C2190 VDD.n289 GND 0.006248f
C2191 VDD.n290 GND 0.007763f
C2192 VDD.n291 GND 0.006248f
C2193 VDD.n292 GND 0.007763f
C2194 VDD.n293 GND 0.594542f
C2195 VDD.n294 GND 0.007763f
C2196 VDD.n295 GND 0.006248f
C2197 VDD.n296 GND 0.007763f
C2198 VDD.n297 GND 0.006248f
C2199 VDD.n298 GND 0.007763f
C2200 VDD.n299 GND 0.576706f
C2201 VDD.n300 GND 0.007763f
C2202 VDD.n301 GND 0.006248f
C2203 VDD.n302 GND 0.007763f
C2204 VDD.n303 GND 0.006248f
C2205 VDD.n304 GND 0.007763f
C2206 VDD.n305 GND 0.594542f
C2207 VDD.n306 GND 0.007763f
C2208 VDD.n307 GND 0.006248f
C2209 VDD.n308 GND 0.007763f
C2210 VDD.n309 GND 0.006248f
C2211 VDD.n310 GND 0.007763f
C2212 VDD.n311 GND 0.594542f
C2213 VDD.n312 GND 0.007763f
C2214 VDD.n313 GND 0.006248f
C2215 VDD.n314 GND 0.007763f
C2216 VDD.n315 GND 0.006248f
C2217 VDD.n316 GND 0.007763f
C2218 VDD.n317 GND 0.594542f
C2219 VDD.n318 GND 0.007763f
C2220 VDD.n319 GND 0.006248f
C2221 VDD.n320 GND 0.007763f
C2222 VDD.n321 GND 0.006248f
C2223 VDD.n322 GND 0.007763f
C2224 VDD.n323 GND 0.564815f
C2225 VDD.n324 GND 0.007763f
C2226 VDD.n325 GND 0.006248f
C2227 VDD.n326 GND 0.007763f
C2228 VDD.n327 GND 0.006248f
C2229 VDD.n328 GND 0.007763f
C2230 VDD.n329 GND 0.594542f
C2231 VDD.n330 GND 0.007763f
C2232 VDD.n331 GND 0.006248f
C2233 VDD.n332 GND 0.007763f
C2234 VDD.n333 GND 0.006248f
C2235 VDD.n334 GND 0.007763f
C2236 VDD.n335 GND 0.594542f
C2237 VDD.n336 GND 0.007763f
C2238 VDD.n337 GND 0.006248f
C2239 VDD.n338 GND 0.007763f
C2240 VDD.n339 GND 0.006248f
C2241 VDD.n340 GND 0.007763f
C2242 VDD.n341 GND 0.594542f
C2243 VDD.n342 GND 0.007763f
C2244 VDD.n343 GND 0.006248f
C2245 VDD.n344 GND 0.007763f
C2246 VDD.n345 GND 0.006248f
C2247 VDD.n346 GND 0.007763f
C2248 VDD.n347 GND 0.552924f
C2249 VDD.n348 GND 0.007763f
C2250 VDD.n349 GND 0.006248f
C2251 VDD.n350 GND 0.007763f
C2252 VDD.n351 GND 0.006248f
C2253 VDD.n352 GND 0.007763f
C2254 VDD.n353 GND 0.594542f
C2255 VDD.n354 GND 0.007763f
C2256 VDD.n355 GND 0.006248f
C2257 VDD.n356 GND 0.007763f
C2258 VDD.n357 GND 0.006248f
C2259 VDD.n358 GND 0.007763f
C2260 VDD.n359 GND 0.594542f
C2261 VDD.n360 GND 0.007763f
C2262 VDD.n361 GND 0.006248f
C2263 VDD.n362 GND 0.007763f
C2264 VDD.n363 GND 0.006248f
C2265 VDD.n364 GND 0.007763f
C2266 VDD.n365 GND 0.594542f
C2267 VDD.n366 GND 0.007763f
C2268 VDD.n367 GND 0.006248f
C2269 VDD.n368 GND 0.007763f
C2270 VDD.n369 GND 0.006248f
C2271 VDD.n370 GND 0.007763f
C2272 VDD.n371 GND 0.594542f
C2273 VDD.n372 GND 0.007763f
C2274 VDD.n373 GND 0.006248f
C2275 VDD.n374 GND 0.007763f
C2276 VDD.n375 GND 0.006248f
C2277 VDD.n376 GND 0.007763f
C2278 VDD.n377 GND 0.594542f
C2279 VDD.n378 GND 0.007763f
C2280 VDD.n379 GND 0.006248f
C2281 VDD.n380 GND 0.007763f
C2282 VDD.n381 GND 0.006248f
C2283 VDD.n382 GND 0.007763f
C2284 VDD.n383 GND 0.594542f
C2285 VDD.n384 GND 0.007763f
C2286 VDD.n385 GND 0.006248f
C2287 VDD.n386 GND 0.007763f
C2288 VDD.n387 GND 0.006248f
C2289 VDD.n388 GND 0.007763f
C2290 VDD.n389 GND 0.594542f
C2291 VDD.n390 GND 0.007763f
C2292 VDD.n391 GND 0.006248f
C2293 VDD.n392 GND 0.856726f
C2294 VDD.n393 GND 0.019093f
C2295 VDD.n394 GND 4.25098f
C2296 VDD.n395 GND 0.019093f
C2297 VDD.n396 GND 0.006909f
C2298 VDD.n397 GND 0.003959f
C2299 VDD.n398 GND 0.005279f
C2300 VDD.n399 GND 0.005279f
C2301 VDD.t101 GND 6.69455f
C2302 VDD.t114 GND 3.20458f
C2303 VDD.n400 GND 0.597515f
C2304 VDD.n401 GND 0.005279f
C2305 VDD.n402 GND 0.005279f
C2306 VDD.n403 GND 0.005279f
C2307 VDD.n405 GND 0.005279f
C2308 VDD.t43 GND 0.118717f
C2309 VDD.t42 GND 0.138462f
C2310 VDD.t40 GND 0.726908f
C2311 VDD.n406 GND 0.089246f
C2312 VDD.n407 GND 0.051676f
C2313 VDD.n408 GND 0.005279f
C2314 VDD.n410 GND 0.013069f
C2315 VDD.n411 GND 0.005279f
C2316 VDD.n412 GND 0.005279f
C2317 VDD.n413 GND 0.404289f
C2318 VDD.n414 GND 0.005279f
C2319 VDD.n415 GND 0.603461f
C2320 VDD.n416 GND 0.005279f
C2321 VDD.n417 GND 0.005279f
C2322 VDD.n418 GND 0.013069f
C2323 VDD.n419 GND 0.005279f
C2324 VDD.n420 GND 0.005279f
C2325 VDD.n421 GND 0.404289f
C2326 VDD.n422 GND 0.005279f
C2327 VDD.n423 GND 0.005279f
C2328 VDD.n424 GND 0.005279f
C2329 VDD.n425 GND 0.005279f
C2330 VDD.n426 GND 0.005279f
C2331 VDD.n427 GND 0.013559f
C2332 VDD.n428 GND 0.005279f
C2333 VDD.n429 GND 0.005279f
C2334 VDD.n431 GND 0.005279f
C2335 VDD.n432 GND 0.005279f
C2336 VDD.n434 GND 0.005279f
C2337 VDD.n435 GND 0.031803f
C2338 VDD.n437 GND 0.003959f
C2339 VDD.n438 GND 0.005279f
C2340 VDD.n439 GND 0.005279f
C2341 VDD.n441 GND 0.005279f
C2342 VDD.n442 GND 0.004774f
C2343 VDD.n444 GND 0.005279f
C2344 VDD.t59 GND 0.118717f
C2345 VDD.t58 GND 0.138462f
C2346 VDD.t57 GND 0.726908f
C2347 VDD.n445 GND 0.089246f
C2348 VDD.n446 GND 0.051676f
C2349 VDD.n447 GND 0.007544f
C2350 VDD.n448 GND 0.005279f
C2351 VDD.n449 GND 0.005279f
C2352 VDD.n450 GND 0.356725f
C2353 VDD.n451 GND 0.005279f
C2354 VDD.n452 GND 0.005279f
C2355 VDD.n453 GND 0.005279f
C2356 VDD.n454 GND 0.005279f
C2357 VDD.n455 GND 0.005279f
C2358 VDD.n456 GND 0.347807f
C2359 VDD.n457 GND 0.005279f
C2360 VDD.n458 GND 0.005279f
C2361 VDD.t41 GND 0.202144f
C2362 VDD.n459 GND 0.005279f
C2363 VDD.n460 GND 0.005279f
C2364 VDD.n461 GND 0.005279f
C2365 VDD.n462 GND 0.005279f
C2366 VDD.n463 GND 0.404289f
C2367 VDD.n464 GND 0.005279f
C2368 VDD.n465 GND 0.005279f
C2369 VDD.t202 GND 0.202144f
C2370 VDD.n466 GND 0.005279f
C2371 VDD.n467 GND 0.005279f
C2372 VDD.n468 GND 0.005279f
C2373 VDD.n469 GND 0.404289f
C2374 VDD.n470 GND 0.005279f
C2375 VDD.n471 GND 0.005279f
C2376 VDD.n472 GND 0.005279f
C2377 VDD.n473 GND 0.005279f
C2378 VDD.n474 GND 0.005279f
C2379 VDD.n475 GND 0.404289f
C2380 VDD.n476 GND 0.005279f
C2381 VDD.n477 GND 0.005279f
C2382 VDD.n478 GND 0.005279f
C2383 VDD.n479 GND 0.005279f
C2384 VDD.n480 GND 0.005279f
C2385 VDD.n481 GND 0.404289f
C2386 VDD.n482 GND 0.005279f
C2387 VDD.n483 GND 0.005279f
C2388 VDD.n484 GND 0.005279f
C2389 VDD.n485 GND 0.005279f
C2390 VDD.n486 GND 0.005279f
C2391 VDD.n487 GND 0.404289f
C2392 VDD.n488 GND 0.005279f
C2393 VDD.n489 GND 0.005279f
C2394 VDD.n490 GND 0.005279f
C2395 VDD.n491 GND 0.005279f
C2396 VDD.n492 GND 0.005279f
C2397 VDD.n493 GND 0.282408f
C2398 VDD.n494 GND 0.005279f
C2399 VDD.n495 GND 0.005279f
C2400 VDD.n496 GND 0.005279f
C2401 VDD.n497 GND 0.005279f
C2402 VDD.n498 GND 0.005279f
C2403 VDD.t104 GND 0.202144f
C2404 VDD.n499 GND 0.005279f
C2405 VDD.n500 GND 0.005279f
C2406 VDD.t198 GND 0.202144f
C2407 VDD.n501 GND 0.005279f
C2408 VDD.n502 GND 0.005279f
C2409 VDD.n503 GND 0.005279f
C2410 VDD.n504 GND 0.404289f
C2411 VDD.n505 GND 0.005279f
C2412 VDD.n506 GND 0.005279f
C2413 VDD.n507 GND 0.27349f
C2414 VDD.n508 GND 0.005279f
C2415 VDD.n509 GND 0.005279f
C2416 VDD.n510 GND 0.005279f
C2417 VDD.n511 GND 0.404289f
C2418 VDD.n512 GND 0.005279f
C2419 VDD.n513 GND 0.005279f
C2420 VDD.n514 GND 0.005279f
C2421 VDD.n515 GND 0.005279f
C2422 VDD.n516 GND 0.005279f
C2423 VDD.n517 GND 0.404289f
C2424 VDD.n518 GND 0.005279f
C2425 VDD.n519 GND 0.005279f
C2426 VDD.n520 GND 0.005279f
C2427 VDD.n521 GND 0.005279f
C2428 VDD.n522 GND 0.005279f
C2429 VDD.n523 GND 0.404289f
C2430 VDD.n524 GND 0.005279f
C2431 VDD.n525 GND 0.005279f
C2432 VDD.n526 GND 0.005279f
C2433 VDD.n527 GND 0.005279f
C2434 VDD.n528 GND 0.005279f
C2435 VDD.n529 GND 0.217008f
C2436 VDD.n530 GND 0.005279f
C2437 VDD.n531 GND 0.005279f
C2438 VDD.n532 GND 0.005279f
C2439 VDD.n533 GND 0.005279f
C2440 VDD.n534 GND 0.005279f
C2441 VDD.t116 GND 0.202144f
C2442 VDD.n535 GND 0.005279f
C2443 VDD.n536 GND 0.005279f
C2444 VDD.t84 GND 0.202144f
C2445 VDD.n537 GND 0.005279f
C2446 VDD.n538 GND 0.005279f
C2447 VDD.n539 GND 0.005279f
C2448 VDD.n540 GND 0.404289f
C2449 VDD.n541 GND 0.005279f
C2450 VDD.n542 GND 0.005279f
C2451 VDD.n543 GND 0.338889f
C2452 VDD.n544 GND 0.005279f
C2453 VDD.n545 GND 0.005279f
C2454 VDD.n546 GND 0.005279f
C2455 VDD.n547 GND 0.404289f
C2456 VDD.n548 GND 0.005279f
C2457 VDD.n549 GND 0.005279f
C2458 VDD.n550 GND 0.005279f
C2459 VDD.n551 GND 0.005279f
C2460 VDD.n552 GND 0.005279f
C2461 VDD.n553 GND 0.404289f
C2462 VDD.n554 GND 0.005279f
C2463 VDD.n555 GND 0.005279f
C2464 VDD.n556 GND 0.005279f
C2465 VDD.n557 GND 0.005279f
C2466 VDD.n558 GND 0.005279f
C2467 VDD.n559 GND 0.404289f
C2468 VDD.n560 GND 0.005279f
C2469 VDD.n561 GND 0.005279f
C2470 VDD.n562 GND 0.005279f
C2471 VDD.n563 GND 0.005279f
C2472 VDD.n564 GND 0.005279f
C2473 VDD.n565 GND 0.404289f
C2474 VDD.n566 GND 0.005279f
C2475 VDD.n567 GND 0.005279f
C2476 VDD.n568 GND 0.005279f
C2477 VDD.n569 GND 0.005279f
C2478 VDD.n570 GND 0.005279f
C2479 VDD.n571 GND 0.404289f
C2480 VDD.n572 GND 0.005279f
C2481 VDD.n573 GND 0.005279f
C2482 VDD.n574 GND 0.005279f
C2483 VDD.n575 GND 0.005279f
C2484 VDD.n576 GND 0.005279f
C2485 VDD.n577 GND 0.404289f
C2486 VDD.n578 GND 0.005279f
C2487 VDD.n579 GND 0.005279f
C2488 VDD.n580 GND 0.005279f
C2489 VDD.n581 GND 0.005279f
C2490 VDD.n582 GND 0.005279f
C2491 VDD.t200 GND 0.202144f
C2492 VDD.n583 GND 0.005279f
C2493 VDD.n584 GND 0.005279f
C2494 VDD.n585 GND 0.005279f
C2495 VDD.n586 GND 0.005279f
C2496 VDD.n587 GND 0.005279f
C2497 VDD.n588 GND 0.404289f
C2498 VDD.n589 GND 0.005279f
C2499 VDD.n590 GND 0.005279f
C2500 VDD.n591 GND 0.258626f
C2501 VDD.n592 GND 0.005279f
C2502 VDD.n593 GND 0.005279f
C2503 VDD.n594 GND 0.005279f
C2504 VDD.n595 GND 0.404289f
C2505 VDD.n596 GND 0.005279f
C2506 VDD.n597 GND 0.005279f
C2507 VDD.n598 GND 0.005279f
C2508 VDD.n599 GND 0.005279f
C2509 VDD.n600 GND 0.005279f
C2510 VDD.n601 GND 0.338889f
C2511 VDD.n602 GND 0.005279f
C2512 VDD.n603 GND 0.005279f
C2513 VDD.n604 GND 0.005279f
C2514 VDD.n605 GND 0.005279f
C2515 VDD.n606 GND 0.005279f
C2516 VDD.n607 GND 0.404289f
C2517 VDD.n608 GND 0.005279f
C2518 VDD.n609 GND 0.005279f
C2519 VDD.t90 GND 0.202144f
C2520 VDD.n610 GND 0.005279f
C2521 VDD.n611 GND 0.005279f
C2522 VDD.n612 GND 0.005279f
C2523 VDD.n613 GND 0.404289f
C2524 VDD.n614 GND 0.005279f
C2525 VDD.n615 GND 0.005279f
C2526 VDD.n616 GND 0.005279f
C2527 VDD.n617 GND 0.005279f
C2528 VDD.n618 GND 0.005279f
C2529 VDD.t1 GND 0.202144f
C2530 VDD.n619 GND 0.005279f
C2531 VDD.n620 GND 0.005279f
C2532 VDD.n621 GND 0.005279f
C2533 VDD.n622 GND 0.005279f
C2534 VDD.n623 GND 0.005279f
C2535 VDD.n624 GND 0.404289f
C2536 VDD.n625 GND 0.005279f
C2537 VDD.n626 GND 0.005279f
C2538 VDD.n627 GND 0.324026f
C2539 VDD.n628 GND 0.005279f
C2540 VDD.n629 GND 0.005279f
C2541 VDD.n630 GND 0.005279f
C2542 VDD.n631 GND 0.404289f
C2543 VDD.n632 GND 0.005279f
C2544 VDD.n633 GND 0.005279f
C2545 VDD.n634 GND 0.005279f
C2546 VDD.n635 GND 0.005279f
C2547 VDD.n636 GND 0.005279f
C2548 VDD.n637 GND 0.27349f
C2549 VDD.n638 GND 0.005279f
C2550 VDD.n639 GND 0.005279f
C2551 VDD.n640 GND 0.005279f
C2552 VDD.n641 GND 0.005279f
C2553 VDD.n642 GND 0.005279f
C2554 VDD.n643 GND 0.404289f
C2555 VDD.n644 GND 0.005279f
C2556 VDD.n645 GND 0.005279f
C2557 VDD.t0 GND 0.202144f
C2558 VDD.n646 GND 0.005279f
C2559 VDD.n647 GND 0.005279f
C2560 VDD.n648 GND 0.005279f
C2561 VDD.n649 GND 0.404289f
C2562 VDD.n650 GND 0.005279f
C2563 VDD.n651 GND 0.005279f
C2564 VDD.n652 GND 0.005279f
C2565 VDD.n653 GND 0.005279f
C2566 VDD.n654 GND 0.005279f
C2567 VDD.t109 GND 0.202144f
C2568 VDD.n655 GND 0.005279f
C2569 VDD.n656 GND 0.005279f
C2570 VDD.n657 GND 0.005279f
C2571 VDD.n658 GND 0.005279f
C2572 VDD.n659 GND 0.005279f
C2573 VDD.n660 GND 0.404289f
C2574 VDD.n661 GND 0.005279f
C2575 VDD.n662 GND 0.005279f
C2576 VDD.n663 GND 0.389425f
C2577 VDD.n664 GND 0.005279f
C2578 VDD.n665 GND 0.005279f
C2579 VDD.n666 GND 0.005279f
C2580 VDD.n667 GND 0.404289f
C2581 VDD.n668 GND 0.005279f
C2582 VDD.n669 GND 0.005279f
C2583 VDD.n670 GND 0.005279f
C2584 VDD.n671 GND 0.005279f
C2585 VDD.n672 GND 0.005279f
C2586 VDD.n673 GND 0.404289f
C2587 VDD.n674 GND 0.005279f
C2588 VDD.n675 GND 0.005279f
C2589 VDD.n676 GND 0.005279f
C2590 VDD.n677 GND 0.005279f
C2591 VDD.n678 GND 0.005279f
C2592 VDD.n679 GND 0.404289f
C2593 VDD.n680 GND 0.005279f
C2594 VDD.n681 GND 0.005279f
C2595 VDD.n682 GND 0.005279f
C2596 VDD.n683 GND 0.005279f
C2597 VDD.n684 GND 0.005279f
C2598 VDD.t9 GND 0.202144f
C2599 VDD.n685 GND 0.005279f
C2600 VDD.n686 GND 0.005279f
C2601 VDD.n687 GND 0.005279f
C2602 VDD.n688 GND 0.005279f
C2603 VDD.n689 GND 0.005279f
C2604 VDD.n690 GND 0.404289f
C2605 VDD.n691 GND 0.005279f
C2606 VDD.n692 GND 0.005279f
C2607 VDD.t96 GND 0.202144f
C2608 VDD.n693 GND 0.005279f
C2609 VDD.n694 GND 0.005279f
C2610 VDD.n695 GND 0.005279f
C2611 VDD.n696 GND 0.404289f
C2612 VDD.n697 GND 0.005279f
C2613 VDD.n698 GND 0.005279f
C2614 VDD.n699 GND 0.005279f
C2615 VDD.n700 GND 0.013069f
C2616 VDD.n701 GND 0.013069f
C2617 VDD.n702 GND 0.603461f
C2618 VDD.n703 GND 0.005279f
C2619 VDD.n704 GND 0.005279f
C2620 VDD.n705 GND 0.013069f
C2621 VDD.n706 GND 0.005279f
C2622 VDD.n707 GND 0.005279f
C2623 VDD.n708 GND 0.603461f
C2624 VDD.n732 GND 0.013559f
C2625 VDD.n733 GND 0.013069f
C2626 VDD.n734 GND 0.005279f
C2627 VDD.n735 GND 0.013069f
C2628 VDD.t56 GND 0.118717f
C2629 VDD.t55 GND 0.138462f
C2630 VDD.t53 GND 0.726908f
C2631 VDD.n736 GND 0.089246f
C2632 VDD.n737 GND 0.051676f
C2633 VDD.n738 GND 0.007544f
C2634 VDD.n739 GND 0.005279f
C2635 VDD.n740 GND 0.005279f
C2636 VDD.n741 GND 0.404289f
C2637 VDD.n742 GND 0.005279f
C2638 VDD.n743 GND 0.005279f
C2639 VDD.n744 GND 0.005279f
C2640 VDD.n745 GND 0.013069f
C2641 VDD.n746 GND 0.005279f
C2642 VDD.t83 GND 0.118717f
C2643 VDD.t82 GND 0.138462f
C2644 VDD.t81 GND 0.726908f
C2645 VDD.n747 GND 0.089246f
C2646 VDD.n748 GND 0.051676f
C2647 VDD.n749 GND 0.005279f
C2648 VDD.n750 GND 0.005279f
C2649 VDD.n751 GND 0.404289f
C2650 VDD.n752 GND 0.005279f
C2651 VDD.n753 GND 0.005279f
C2652 VDD.n754 GND 0.005279f
C2653 VDD.n755 GND 0.005279f
C2654 VDD.n756 GND 0.005279f
C2655 VDD.t111 GND 0.202144f
C2656 VDD.n757 GND 0.005279f
C2657 VDD.n758 GND 0.005279f
C2658 VDD.n759 GND 0.005279f
C2659 VDD.n760 GND 0.005279f
C2660 VDD.n761 GND 0.005279f
C2661 VDD.n762 GND 0.005279f
C2662 VDD.n763 GND 0.404289f
C2663 VDD.n764 GND 0.005279f
C2664 VDD.n765 GND 0.005279f
C2665 VDD.t54 GND 0.202144f
C2666 VDD.n766 GND 0.005279f
C2667 VDD.n767 GND 0.005279f
C2668 VDD.n768 GND 0.005279f
C2669 VDD.n769 GND 0.404289f
C2670 VDD.n770 GND 0.005279f
C2671 VDD.n771 GND 0.005279f
C2672 VDD.n772 GND 0.005279f
C2673 VDD.n773 GND 0.005279f
C2674 VDD.n774 GND 0.005279f
C2675 VDD.n775 GND 0.404289f
C2676 VDD.n776 GND 0.005279f
C2677 VDD.n777 GND 0.005279f
C2678 VDD.n778 GND 0.005279f
C2679 VDD.n779 GND 0.005279f
C2680 VDD.n780 GND 0.005279f
C2681 VDD.n781 GND 0.404289f
C2682 VDD.n782 GND 0.005279f
C2683 VDD.n783 GND 0.005279f
C2684 VDD.n784 GND 0.005279f
C2685 VDD.n785 GND 0.005279f
C2686 VDD.n786 GND 0.005279f
C2687 VDD.n787 GND 0.389425f
C2688 VDD.n788 GND 0.005279f
C2689 VDD.n789 GND 0.005279f
C2690 VDD.n790 GND 0.005279f
C2691 VDD.n791 GND 0.005279f
C2692 VDD.n792 GND 0.005279f
C2693 VDD.n793 GND 0.404289f
C2694 VDD.n794 GND 0.005279f
C2695 VDD.n795 GND 0.005279f
C2696 VDD.t93 GND 0.202144f
C2697 VDD.n796 GND 0.005279f
C2698 VDD.n797 GND 0.005279f
C2699 VDD.n798 GND 0.005279f
C2700 VDD.n799 GND 0.404289f
C2701 VDD.n800 GND 0.005279f
C2702 VDD.n801 GND 0.005279f
C2703 VDD.n802 GND 0.005279f
C2704 VDD.n803 GND 0.005279f
C2705 VDD.n804 GND 0.005279f
C2706 VDD.t113 GND 0.202144f
C2707 VDD.n805 GND 0.005279f
C2708 VDD.n806 GND 0.005279f
C2709 VDD.n807 GND 0.005279f
C2710 VDD.n808 GND 0.005279f
C2711 VDD.n809 GND 0.005279f
C2712 VDD.n810 GND 0.404289f
C2713 VDD.n811 GND 0.005279f
C2714 VDD.n812 GND 0.005279f
C2715 VDD.n813 GND 0.27349f
C2716 VDD.n814 GND 0.005279f
C2717 VDD.n815 GND 0.005279f
C2718 VDD.n816 GND 0.005279f
C2719 VDD.n817 GND 0.404289f
C2720 VDD.n818 GND 0.005279f
C2721 VDD.n819 GND 0.005279f
C2722 VDD.n820 GND 0.005279f
C2723 VDD.n821 GND 0.005279f
C2724 VDD.n822 GND 0.005279f
C2725 VDD.n823 GND 0.324026f
C2726 VDD.n824 GND 0.005279f
C2727 VDD.n825 GND 0.005279f
C2728 VDD.n826 GND 0.005279f
C2729 VDD.n827 GND 0.005279f
C2730 VDD.n828 GND 0.005279f
C2731 VDD.n829 GND 0.404289f
C2732 VDD.n830 GND 0.005279f
C2733 VDD.n831 GND 0.005279f
C2734 VDD.t105 GND 0.202144f
C2735 VDD.n832 GND 0.005279f
C2736 VDD.n833 GND 0.005279f
C2737 VDD.n834 GND 0.005279f
C2738 VDD.n835 GND 0.404289f
C2739 VDD.n836 GND 0.005279f
C2740 VDD.n837 GND 0.005279f
C2741 VDD.n838 GND 0.005279f
C2742 VDD.n839 GND 0.005279f
C2743 VDD.n840 GND 0.005279f
C2744 VDD.t95 GND 0.202144f
C2745 VDD.n841 GND 0.005279f
C2746 VDD.n842 GND 0.005279f
C2747 VDD.n843 GND 0.005279f
C2748 VDD.n844 GND 0.005279f
C2749 VDD.n845 GND 0.005279f
C2750 VDD.n846 GND 0.404289f
C2751 VDD.n847 GND 0.005279f
C2752 VDD.n848 GND 0.005279f
C2753 VDD.n849 GND 0.338889f
C2754 VDD.n850 GND 0.005279f
C2755 VDD.n851 GND 0.005279f
C2756 VDD.n852 GND 0.005279f
C2757 VDD.n853 GND 0.404289f
C2758 VDD.n854 GND 0.005279f
C2759 VDD.n855 GND 0.005279f
C2760 VDD.n856 GND 0.005279f
C2761 VDD.n857 GND 0.005279f
C2762 VDD.n858 GND 0.005279f
C2763 VDD.n859 GND 0.258626f
C2764 VDD.n860 GND 0.005279f
C2765 VDD.n861 GND 0.005279f
C2766 VDD.n862 GND 0.005279f
C2767 VDD.n863 GND 0.005279f
C2768 VDD.n864 GND 0.005279f
C2769 VDD.n865 GND 0.404289f
C2770 VDD.n866 GND 0.005279f
C2771 VDD.n867 GND 0.005279f
C2772 VDD.t86 GND 0.202144f
C2773 VDD.n868 GND 0.005279f
C2774 VDD.n869 GND 0.005279f
C2775 VDD.n870 GND 0.005279f
C2776 VDD.n871 GND 0.404289f
C2777 VDD.n872 GND 0.005279f
C2778 VDD.n873 GND 0.005279f
C2779 VDD.n874 GND 0.005279f
C2780 VDD.n875 GND 0.005279f
C2781 VDD.n876 GND 0.005279f
C2782 VDD.n877 GND 0.404289f
C2783 VDD.n878 GND 0.005279f
C2784 VDD.n879 GND 0.005279f
C2785 VDD.n880 GND 0.005279f
C2786 VDD.n881 GND 0.005279f
C2787 VDD.n882 GND 0.005279f
C2788 VDD.n883 GND 0.005279f
C2789 VDD.n884 GND 0.005279f
C2790 VDD.n885 GND 0.005279f
C2791 VDD.n886 GND 0.005279f
C2792 VDD.n887 GND 0.404289f
C2793 VDD.n888 GND 0.005279f
C2794 VDD.n889 GND 0.005279f
C2795 VDD.n890 GND 0.005279f
C2796 VDD.n891 GND 0.005279f
C2797 VDD.n892 GND 0.005279f
C2798 VDD.n893 GND 0.404289f
C2799 VDD.n894 GND 0.005279f
C2800 VDD.n895 GND 0.005279f
C2801 VDD.n896 GND 0.005279f
C2802 VDD.n897 GND 0.005279f
C2803 VDD.n898 GND 0.005279f
C2804 VDD.n899 GND 0.005279f
C2805 VDD.n900 GND 0.404289f
C2806 VDD.n901 GND 0.005279f
C2807 VDD.n902 GND 0.005279f
C2808 VDD.n903 GND 0.005279f
C2809 VDD.n904 GND 0.005279f
C2810 VDD.n905 GND 0.005279f
C2811 VDD.n906 GND 0.404289f
C2812 VDD.n907 GND 0.005279f
C2813 VDD.n908 GND 0.005279f
C2814 VDD.n909 GND 0.005279f
C2815 VDD.n910 GND 0.005279f
C2816 VDD.n911 GND 0.005279f
C2817 VDD.n912 GND 0.338889f
C2818 VDD.n913 GND 0.005279f
C2819 VDD.n914 GND 0.005279f
C2820 VDD.n915 GND 0.005279f
C2821 VDD.n916 GND 0.005279f
C2822 VDD.n917 GND 0.005279f
C2823 VDD.t102 GND 0.202144f
C2824 VDD.n918 GND 0.005279f
C2825 VDD.n919 GND 0.005279f
C2826 VDD.t3 GND 0.202144f
C2827 VDD.n920 GND 0.005279f
C2828 VDD.n921 GND 0.005279f
C2829 VDD.n922 GND 0.005279f
C2830 VDD.n923 GND 0.404289f
C2831 VDD.n924 GND 0.005279f
C2832 VDD.n925 GND 0.005279f
C2833 VDD.n926 GND 0.217008f
C2834 VDD.n927 GND 0.005279f
C2835 VDD.n928 GND 0.005279f
C2836 VDD.n929 GND 0.005279f
C2837 VDD.n930 GND 0.404289f
C2838 VDD.n931 GND 0.005279f
C2839 VDD.n932 GND 0.005279f
C2840 VDD.n933 GND 0.005279f
C2841 VDD.n934 GND 0.005279f
C2842 VDD.n935 GND 0.005279f
C2843 VDD.n936 GND 0.404289f
C2844 VDD.n937 GND 0.005279f
C2845 VDD.n938 GND 0.005279f
C2846 VDD.n939 GND 0.005279f
C2847 VDD.n940 GND 0.005279f
C2848 VDD.n941 GND 0.005279f
C2849 VDD.n942 GND 0.404289f
C2850 VDD.n943 GND 0.005279f
C2851 VDD.n944 GND 0.005279f
C2852 VDD.n945 GND 0.005279f
C2853 VDD.n946 GND 0.005279f
C2854 VDD.n947 GND 0.005279f
C2855 VDD.n948 GND 0.27349f
C2856 VDD.n949 GND 0.005279f
C2857 VDD.n950 GND 0.005279f
C2858 VDD.n951 GND 0.005279f
C2859 VDD.n952 GND 0.005279f
C2860 VDD.n953 GND 0.005279f
C2861 VDD.t98 GND 0.202144f
C2862 VDD.n954 GND 0.005279f
C2863 VDD.n955 GND 0.005279f
C2864 VDD.t107 GND 0.202144f
C2865 VDD.n956 GND 0.005279f
C2866 VDD.n957 GND 0.005279f
C2867 VDD.n958 GND 0.005279f
C2868 VDD.n959 GND 0.404289f
C2869 VDD.n960 GND 0.005279f
C2870 VDD.n961 GND 0.005279f
C2871 VDD.n962 GND 0.282408f
C2872 VDD.n963 GND 0.005279f
C2873 VDD.n964 GND 0.005279f
C2874 VDD.n965 GND 0.005279f
C2875 VDD.n966 GND 0.404289f
C2876 VDD.n967 GND 0.005279f
C2877 VDD.n968 GND 0.005279f
C2878 VDD.n969 GND 0.005279f
C2879 VDD.n970 GND 0.005279f
C2880 VDD.n971 GND 0.005279f
C2881 VDD.n972 GND 0.404289f
C2882 VDD.n973 GND 0.005279f
C2883 VDD.n974 GND 0.005279f
C2884 VDD.n975 GND 0.005279f
C2885 VDD.n976 GND 0.005279f
C2886 VDD.n977 GND 0.005279f
C2887 VDD.n978 GND 0.404289f
C2888 VDD.n979 GND 0.005279f
C2889 VDD.n980 GND 0.005279f
C2890 VDD.n981 GND 0.005279f
C2891 VDD.n982 GND 0.005279f
C2892 VDD.n983 GND 0.005279f
C2893 VDD.n984 GND 0.404289f
C2894 VDD.n985 GND 0.005279f
C2895 VDD.n986 GND 0.005279f
C2896 VDD.n987 GND 0.005279f
C2897 VDD.n988 GND 0.005279f
C2898 VDD.n989 GND 0.005279f
C2899 VDD.t88 GND 0.202144f
C2900 VDD.n990 GND 0.005279f
C2901 VDD.n991 GND 0.005279f
C2902 VDD.n992 GND 0.005279f
C2903 VDD.n993 GND 0.005279f
C2904 VDD.n994 GND 0.005279f
C2905 VDD.t5 GND 0.202144f
C2906 VDD.n995 GND 0.005279f
C2907 VDD.n996 GND 0.005279f
C2908 VDD.n997 GND 0.347807f
C2909 VDD.n998 GND 0.005279f
C2910 VDD.n999 GND 0.005279f
C2911 VDD.n1000 GND 0.005279f
C2912 VDD.n1001 GND 0.404289f
C2913 VDD.n1002 GND 0.005279f
C2914 VDD.n1003 GND 0.005279f
C2915 VDD.n1004 GND 0.356725f
C2916 VDD.n1005 GND 0.005279f
C2917 VDD.n1006 GND 0.005279f
C2918 VDD.n1007 GND 0.005279f
C2919 VDD.n1008 GND 0.404289f
C2920 VDD.n1009 GND 0.005279f
C2921 VDD.n1010 GND 0.005279f
C2922 VDD.n1011 GND 0.005279f
C2923 VDD.n1012 GND 0.013069f
C2924 VDD.n1013 GND 0.013069f
C2925 VDD.n1014 GND 0.603461f
C2926 VDD.n1015 GND 0.005279f
C2927 VDD.n1016 GND 0.005279f
C2928 VDD.n1017 GND 0.013069f
C2929 VDD.n1018 GND 0.005279f
C2930 VDD.n1019 GND 0.005279f
C2931 VDD.t91 GND 3.20458f
C2932 VDD.n1030 GND 0.013559f
C2933 VDD.n1042 GND 0.013559f
C2934 VDD.n1043 GND 0.005279f
C2935 VDD.n1044 GND 0.005279f
C2936 VDD.t35 GND 0.118717f
C2937 VDD.t36 GND 0.138462f
C2938 VDD.t34 GND 0.726908f
C2939 VDD.n1045 GND 0.089246f
C2940 VDD.n1046 GND 0.051676f
C2941 VDD.n1047 GND 0.007544f
C2942 VDD.n1048 GND 0.005279f
C2943 VDD.n1049 GND 0.005279f
C2944 VDD.n1050 GND 0.005279f
C2945 VDD.n1051 GND 0.005279f
C2946 VDD.n1052 GND 0.005279f
C2947 VDD.n1053 GND 0.005279f
C2948 VDD.n1054 GND 0.005279f
C2949 VDD.n1055 GND 0.005279f
C2950 VDD.n1056 GND 0.005279f
C2951 VDD.n1057 GND 0.005279f
C2952 VDD.n1058 GND 0.005279f
C2953 VDD.n1059 GND 0.005279f
C2954 VDD.n1060 GND 0.005279f
C2955 VDD.n1061 GND 0.005279f
C2956 VDD.n1062 GND 0.005279f
C2957 VDD.n1063 GND 0.005279f
C2958 VDD.n1064 GND 0.005279f
C2959 VDD.n1065 GND 0.005279f
C2960 VDD.n1066 GND 0.005279f
C2961 VDD.n1067 GND 0.005279f
C2962 VDD.n1068 GND 0.005279f
C2963 VDD.n1069 GND 0.005279f
C2964 VDD.n1070 GND 0.005279f
C2965 VDD.n1071 GND 0.005279f
C2966 VDD.n1072 GND 0.005279f
C2967 VDD.n1073 GND 0.005279f
C2968 VDD.n1074 GND 0.005279f
C2969 VDD.n1075 GND 0.005279f
C2970 VDD.n1076 GND 0.005279f
C2971 VDD.n1077 GND 0.005279f
C2972 VDD.n1078 GND 0.005279f
C2973 VDD.n1079 GND 0.005279f
C2974 VDD.n1080 GND 0.005279f
C2975 VDD.n1081 GND 0.005279f
C2976 VDD.n1082 GND 0.005279f
C2977 VDD.n1083 GND 0.005279f
C2978 VDD.n1084 GND 0.005279f
C2979 VDD.n1085 GND 0.005279f
C2980 VDD.n1086 GND 0.005279f
C2981 VDD.n1087 GND 0.005279f
C2982 VDD.n1088 GND 0.005279f
C2983 VDD.n1089 GND 0.005279f
C2984 VDD.n1090 GND 0.005279f
C2985 VDD.n1091 GND 0.005279f
C2986 VDD.n1092 GND 0.005279f
C2987 VDD.n1093 GND 0.005279f
C2988 VDD.n1094 GND 0.005279f
C2989 VDD.n1095 GND 0.005279f
C2990 VDD.n1096 GND 0.005279f
C2991 VDD.n1097 GND 0.005279f
C2992 VDD.n1098 GND 0.005279f
C2993 VDD.n1099 GND 0.005279f
C2994 VDD.n1100 GND 0.005279f
C2995 VDD.n1101 GND 0.005279f
C2996 VDD.n1102 GND 0.005279f
C2997 VDD.n1103 GND 0.005279f
C2998 VDD.n1104 GND 0.005279f
C2999 VDD.n1105 GND 0.005279f
C3000 VDD.n1106 GND 0.005279f
C3001 VDD.n1107 GND 0.005279f
C3002 VDD.n1108 GND 0.005279f
C3003 VDD.n1109 GND 0.005279f
C3004 VDD.n1110 GND 0.005279f
C3005 VDD.n1111 GND 0.005279f
C3006 VDD.n1112 GND 0.013069f
C3007 VDD.n1113 GND 0.013069f
C3008 VDD.n1114 GND 0.013559f
C3009 VDD.n1115 GND 0.005279f
C3010 VDD.n1116 GND 0.005279f
C3011 VDD.n1117 GND 0.003144f
C3012 VDD.n1118 GND 0.005279f
C3013 VDD.n1119 GND 0.005279f
C3014 VDD.n1120 GND 0.004774f
C3015 VDD.n1121 GND 0.005279f
C3016 VDD.n1122 GND 0.005279f
C3017 VDD.n1123 GND 0.005279f
C3018 VDD.n1124 GND 0.005279f
C3019 VDD.n1125 GND 0.005279f
C3020 VDD.n1126 GND 0.005279f
C3021 VDD.n1127 GND 0.005279f
C3022 VDD.n1128 GND 0.005279f
C3023 VDD.n1129 GND 0.005279f
C3024 VDD.n1130 GND 0.005279f
C3025 VDD.n1131 GND 0.005279f
C3026 VDD.n1132 GND 0.005279f
C3027 VDD.n1133 GND 0.005279f
C3028 VDD.n1134 GND 0.005279f
C3029 VDD.n1135 GND 0.005279f
C3030 VDD.n1136 GND 0.003959f
C3031 VDD.n1137 GND 0.006909f
C3032 VDD.n1138 GND 0.010528f
C3033 VDD.n1139 GND 0.006248f
C3034 VDD.n1140 GND 0.018791f
C3035 VDD.n1141 GND 0.007763f
C3036 VDD.n1142 GND 0.862087f
C3037 VDD.t117 GND 6.69455f
C3038 VDD.n1161 GND 0.007763f
C3039 VDD.n1162 GND 0.007763f
C3040 VDD.n1163 GND 0.007763f
C3041 VDD.n1164 GND 0.007763f
C3042 VDD.n1165 GND 0.007763f
C3043 VDD.n1166 GND 0.007763f
C3044 VDD.n1167 GND 0.00428f
C3045 VDD.t30 GND 0.035989f
C3046 VDD.t29 GND 0.048603f
C3047 VDD.t27 GND 0.295093f
C3048 VDD.n1168 GND 0.062024f
C3049 VDD.n1169 GND 0.044734f
C3050 VDD.n1170 GND 0.007763f
C3051 VDD.n1171 GND 0.007763f
C3052 VDD.n1172 GND 0.007763f
C3053 VDD.n1173 GND 0.007763f
C3054 VDD.n1174 GND 0.007763f
C3055 VDD.n1175 GND 0.007763f
C3056 VDD.n1176 GND 0.007763f
C3057 VDD.n1177 GND 0.007763f
C3058 VDD.n1178 GND 0.007763f
C3059 VDD.n1179 GND 0.007763f
C3060 VDD.n1180 GND 0.007763f
C3061 VDD.n1181 GND 0.007763f
C3062 VDD.n1182 GND 0.007763f
C3063 VDD.n1183 GND 0.007763f
C3064 VDD.n1184 GND 0.007763f
C3065 VDD.n1185 GND 0.007763f
C3066 VDD.n1186 GND 0.007763f
C3067 VDD.n1187 GND 0.007763f
C3068 VDD.n1188 GND 0.007763f
C3069 VDD.n1189 GND 0.007763f
C3070 VDD.n1190 GND 0.007763f
C3071 VDD.n1191 GND 0.007763f
C3072 VDD.n1192 GND 0.007763f
C3073 VDD.n1193 GND 0.007763f
C3074 VDD.n1194 GND 0.007763f
C3075 VDD.n1195 GND 0.007763f
C3076 VDD.n1196 GND 0.007763f
C3077 VDD.n1197 GND 0.006909f
C3078 VDD.n1198 GND 0.019093f
C3079 VDD.n1199 GND 0.007763f
C3080 VDD.n1200 GND 0.006248f
C3081 VDD.n1201 GND 0.007763f
C3082 VDD.n1202 GND 0.594542f
C3083 VDD.n1203 GND 0.007763f
C3084 VDD.n1204 GND 0.006248f
C3085 VDD.n1205 GND 0.007763f
C3086 VDD.n1206 GND 0.006248f
C3087 VDD.n1207 GND 0.007763f
C3088 VDD.t28 GND 0.594542f
C3089 VDD.n1208 GND 0.007763f
C3090 VDD.n1209 GND 0.006248f
C3091 VDD.n1210 GND 0.006248f
C3092 VDD.n1211 GND 0.007763f
C3093 VDD.n1212 GND 0.006248f
C3094 VDD.n1213 GND 0.007763f
C3095 VDD.n1214 GND 0.594542f
C3096 VDD.n1215 GND 0.007763f
C3097 VDD.n1216 GND 0.006248f
C3098 VDD.n1217 GND 0.007763f
C3099 VDD.n1218 GND 0.006248f
C3100 VDD.n1219 GND 0.007763f
C3101 VDD.n1220 GND 0.594542f
C3102 VDD.n1221 GND 0.007763f
C3103 VDD.n1222 GND 0.006248f
C3104 VDD.n1223 GND 0.007763f
C3105 VDD.n1224 GND 0.006248f
C3106 VDD.n1225 GND 0.007763f
C3107 VDD.n1226 GND 0.594542f
C3108 VDD.n1227 GND 0.007763f
C3109 VDD.n1228 GND 0.006248f
C3110 VDD.n1229 GND 0.007763f
C3111 VDD.n1230 GND 0.006248f
C3112 VDD.n1231 GND 0.007763f
C3113 VDD.n1232 GND 0.594542f
C3114 VDD.n1233 GND 0.007763f
C3115 VDD.n1234 GND 0.006248f
C3116 VDD.n1235 GND 0.007763f
C3117 VDD.n1236 GND 0.006248f
C3118 VDD.n1237 GND 0.007763f
C3119 VDD.n1238 GND 0.338889f
C3120 VDD.n1239 GND 0.007763f
C3121 VDD.n1240 GND 0.006248f
C3122 VDD.n1241 GND 0.007763f
C3123 VDD.n1242 GND 0.006248f
C3124 VDD.n1243 GND 0.007763f
C3125 VDD.n1244 GND 0.594542f
C3126 VDD.n1245 GND 0.007763f
C3127 VDD.n1246 GND 0.006248f
C3128 VDD.n1247 GND 0.007763f
C3129 VDD.n1248 GND 0.006248f
C3130 VDD.n1249 GND 0.007763f
C3131 VDD.n1250 GND 0.594542f
C3132 VDD.n1251 GND 0.007763f
C3133 VDD.n1252 GND 0.006248f
C3134 VDD.n1253 GND 0.007763f
C3135 VDD.n1254 GND 0.006248f
C3136 VDD.n1255 GND 0.007763f
C3137 VDD.n1256 GND 0.594542f
C3138 VDD.n1257 GND 0.007763f
C3139 VDD.n1258 GND 0.006248f
C3140 VDD.n1259 GND 0.007763f
C3141 VDD.n1260 GND 0.006248f
C3142 VDD.n1261 GND 0.007763f
C3143 VDD.n1262 GND 0.326998f
C3144 VDD.n1263 GND 0.007763f
C3145 VDD.n1264 GND 0.006248f
C3146 VDD.n1265 GND 0.007763f
C3147 VDD.n1266 GND 0.006248f
C3148 VDD.n1267 GND 0.007763f
C3149 VDD.n1268 GND 0.594542f
C3150 VDD.n1269 GND 0.007763f
C3151 VDD.n1270 GND 0.006248f
C3152 VDD.n1271 GND 0.007763f
C3153 VDD.n1272 GND 0.006248f
C3154 VDD.n1273 GND 0.007763f
C3155 VDD.n1274 GND 0.594542f
C3156 VDD.n1275 GND 0.007763f
C3157 VDD.n1276 GND 0.006248f
C3158 VDD.n1277 GND 0.007763f
C3159 VDD.n1278 GND 0.006248f
C3160 VDD.n1279 GND 0.007763f
C3161 VDD.n1280 GND 0.594542f
C3162 VDD.n1281 GND 0.007763f
C3163 VDD.n1282 GND 0.006248f
C3164 VDD.n1283 GND 0.007763f
C3165 VDD.n1284 GND 0.006248f
C3166 VDD.n1285 GND 0.007763f
C3167 VDD.n1286 GND 0.315107f
C3168 VDD.n1287 GND 0.007763f
C3169 VDD.n1288 GND 0.006248f
C3170 VDD.n1289 GND 0.007763f
C3171 VDD.n1290 GND 0.006248f
C3172 VDD.n1291 GND 0.007763f
C3173 VDD.n1292 GND 0.594542f
C3174 VDD.n1293 GND 0.007763f
C3175 VDD.n1294 GND 0.006248f
C3176 VDD.n1295 GND 0.007763f
C3177 VDD.n1296 GND 0.006248f
C3178 VDD.n1297 GND 0.007763f
C3179 VDD.n1298 GND 0.594542f
C3180 VDD.n1299 GND 0.007763f
C3181 VDD.n1300 GND 0.006248f
C3182 VDD.n1301 GND 0.007763f
C3183 VDD.n1302 GND 0.006248f
C3184 VDD.n1303 GND 0.007763f
C3185 VDD.n1304 GND 0.594542f
C3186 VDD.n1305 GND 0.007763f
C3187 VDD.n1306 GND 0.006248f
C3188 VDD.n1307 GND 0.007763f
C3189 VDD.n1308 GND 0.006248f
C3190 VDD.n1309 GND 0.007763f
C3191 VDD.n1310 GND 0.303217f
C3192 VDD.n1311 GND 0.007763f
C3193 VDD.n1312 GND 0.006248f
C3194 VDD.n1313 GND 0.007763f
C3195 VDD.n1314 GND 0.006248f
C3196 VDD.n1315 GND 0.007763f
C3197 VDD.n1316 GND 0.594542f
C3198 VDD.n1317 GND 0.007763f
C3199 VDD.n1318 GND 0.006248f
C3200 VDD.n1319 GND 0.007763f
C3201 VDD.n1320 GND 0.006248f
C3202 VDD.n1321 GND 0.007763f
C3203 VDD.n1322 GND 0.594542f
C3204 VDD.n1323 GND 0.007763f
C3205 VDD.n1324 GND 0.006248f
C3206 VDD.n1325 GND 0.007763f
C3207 VDD.n1326 GND 0.006248f
C3208 VDD.n1327 GND 0.007763f
C3209 VDD.n1328 GND 0.594542f
C3210 VDD.n1329 GND 0.007763f
C3211 VDD.n1330 GND 0.006248f
C3212 VDD.n1331 GND 0.007763f
C3213 VDD.n1332 GND 0.006248f
C3214 VDD.n1333 GND 0.007763f
C3215 VDD.t122 GND 0.297271f
C3216 VDD.n1334 GND 0.007763f
C3217 VDD.n1335 GND 0.006248f
C3218 VDD.n1336 GND 0.007763f
C3219 VDD.n1337 GND 0.006248f
C3220 VDD.n1338 GND 0.007763f
C3221 VDD.n1339 GND 0.594542f
C3222 VDD.n1340 GND 0.007763f
C3223 VDD.n1341 GND 0.006248f
C3224 VDD.n1342 GND 0.007763f
C3225 VDD.n1343 GND 0.006248f
C3226 VDD.n1344 GND 0.007763f
C3227 VDD.n1345 GND 0.594542f
C3228 VDD.n1346 GND 0.007763f
C3229 VDD.n1347 GND 0.006248f
C3230 VDD.n1348 GND 0.007763f
C3231 VDD.n1349 GND 0.006248f
C3232 VDD.n1350 GND 0.007763f
C3233 VDD.n1351 GND 0.594542f
C3234 VDD.n1352 GND 0.007763f
C3235 VDD.n1353 GND 0.006248f
C3236 VDD.n1354 GND 0.007763f
C3237 VDD.n1355 GND 0.006248f
C3238 VDD.n1356 GND 0.007763f
C3239 VDD.t154 GND 0.297271f
C3240 VDD.n1357 GND 0.007763f
C3241 VDD.n1358 GND 0.006248f
C3242 VDD.n1359 GND 0.007763f
C3243 VDD.n1360 GND 0.006248f
C3244 VDD.n1361 GND 0.007763f
C3245 VDD.n1362 GND 0.594542f
C3246 VDD.n1363 GND 0.007763f
C3247 VDD.n1364 GND 0.006248f
C3248 VDD.n1365 GND 0.007763f
C3249 VDD.n1366 GND 0.006248f
C3250 VDD.n1367 GND 0.007763f
C3251 VDD.n1368 GND 0.594542f
C3252 VDD.n1369 GND 0.007763f
C3253 VDD.n1370 GND 0.006248f
C3254 VDD.n1371 GND 0.007763f
C3255 VDD.n1372 GND 0.006248f
C3256 VDD.n1373 GND 0.007763f
C3257 VDD.n1374 GND 0.594542f
C3258 VDD.n1375 GND 0.007763f
C3259 VDD.n1376 GND 0.006248f
C3260 VDD.n1377 GND 0.007763f
C3261 VDD.n1378 GND 0.006248f
C3262 VDD.n1379 GND 0.007763f
C3263 VDD.t156 GND 0.297271f
C3264 VDD.n1380 GND 0.007763f
C3265 VDD.n1381 GND 0.006248f
C3266 VDD.n1382 GND 0.007763f
C3267 VDD.n1383 GND 0.006248f
C3268 VDD.n1384 GND 0.007763f
C3269 VDD.n1385 GND 0.594542f
C3270 VDD.n1386 GND 0.007763f
C3271 VDD.n1387 GND 0.006248f
C3272 VDD.n1388 GND 0.007763f
C3273 VDD.n1389 GND 0.006248f
C3274 VDD.n1390 GND 0.007763f
C3275 VDD.n1391 GND 0.594542f
C3276 VDD.n1392 GND 0.007763f
C3277 VDD.n1393 GND 0.006248f
C3278 VDD.n1394 GND 0.007763f
C3279 VDD.n1395 GND 0.006248f
C3280 VDD.n1396 GND 0.007763f
C3281 VDD.n1397 GND 0.594542f
C3282 VDD.n1398 GND 0.007763f
C3283 VDD.n1399 GND 0.006248f
C3284 VDD.n1400 GND 0.007763f
C3285 VDD.n1401 GND 0.006248f
C3286 VDD.n1402 GND 0.007763f
C3287 VDD.t147 GND 0.297271f
C3288 VDD.n1403 GND 0.007763f
C3289 VDD.n1404 GND 0.006248f
C3290 VDD.n1405 GND 0.007763f
C3291 VDD.n1406 GND 0.006248f
C3292 VDD.n1407 GND 0.007763f
C3293 VDD.n1408 GND 0.594542f
C3294 VDD.n1409 GND 0.007763f
C3295 VDD.n1410 GND 0.006248f
C3296 VDD.n1411 GND 0.007763f
C3297 VDD.n1412 GND 0.006248f
C3298 VDD.n1413 GND 0.007763f
C3299 VDD.n1414 GND 0.594542f
C3300 VDD.n1415 GND 0.007763f
C3301 VDD.n1416 GND 0.006248f
C3302 VDD.n1417 GND 0.007763f
C3303 VDD.n1418 GND 0.006248f
C3304 VDD.n1419 GND 0.007763f
C3305 VDD.n1420 GND 0.594542f
C3306 VDD.n1421 GND 0.007763f
C3307 VDD.n1422 GND 0.006248f
C3308 VDD.n1423 GND 0.007763f
C3309 VDD.n1424 GND 0.006248f
C3310 VDD.n1425 GND 0.007763f
C3311 VDD.n1426 GND 0.594542f
C3312 VDD.n1427 GND 0.007763f
C3313 VDD.n1428 GND 0.006248f
C3314 VDD.n1429 GND 0.007763f
C3315 VDD.n1430 GND 0.006248f
C3316 VDD.n1431 GND 0.007763f
C3317 VDD.t17 GND 0.594542f
C3318 VDD.n1432 GND 0.007763f
C3319 VDD.n1433 GND 0.006248f
C3320 VDD.n1434 GND 0.007763f
C3321 VDD.n1435 GND 0.006248f
C3322 VDD.n1436 GND 0.007763f
C3323 VDD.n1437 GND 0.594542f
C3324 VDD.n1438 GND 0.007763f
C3325 VDD.n1439 GND 0.006248f
C3326 VDD.n1440 GND 0.018791f
C3327 VDD.n1441 GND 0.005186f
C3328 VDD.n1442 GND 0.018791f
C3329 VDD.n1443 GND 0.862087f
C3330 VDD.n1444 GND 0.018791f
C3331 VDD.n1445 GND 0.005186f
C3332 VDD.n1446 GND 0.007763f
C3333 VDD.t18 GND 0.035989f
C3334 VDD.t19 GND 0.048603f
C3335 VDD.t16 GND 0.295093f
C3336 VDD.n1447 GND 0.062024f
C3337 VDD.n1448 GND 0.044734f
C3338 VDD.n1449 GND 0.009623f
C3339 VDD.n1450 GND 0.007763f
C3340 VDD.n1468 GND 0.007763f
C3341 VDD.n1469 GND 0.007763f
C3342 VDD.n1470 GND 0.019093f
C3343 VDD.n1471 GND 0.006248f
C3344 VDD.n1472 GND 0.007763f
C3345 VDD.n1473 GND 0.007763f
C3346 VDD.n1474 GND 0.007763f
C3347 VDD.n1475 GND 0.007763f
C3348 VDD.n1476 GND 0.006155f
C3349 VDD.n1477 GND 0.007763f
C3350 VDD.n1478 GND 0.007763f
C3351 VDD.n1479 GND 0.007763f
C3352 VDD.n1480 GND 0.006248f
C3353 VDD.n1481 GND 0.007763f
C3354 VDD.n1482 GND 0.007763f
C3355 VDD.n1483 GND 0.007763f
C3356 VDD.n1484 GND 0.007763f
C3357 VDD.n1485 GND 0.007763f
C3358 VDD.n1486 GND 0.006248f
C3359 VDD.n1487 GND 0.007763f
C3360 VDD.n1488 GND 0.007763f
C3361 VDD.n1489 GND 0.007763f
C3362 VDD.n1490 GND 0.007763f
C3363 VDD.n1491 GND 0.007763f
C3364 VDD.t38 GND 0.035989f
C3365 VDD.t39 GND 0.048603f
C3366 VDD.t37 GND 0.295093f
C3367 VDD.n1492 GND 0.062024f
C3368 VDD.n1493 GND 0.044734f
C3369 VDD.n1494 GND 0.009623f
C3370 VDD.n1495 GND 0.007763f
C3371 VDD.n1496 GND 0.007763f
C3372 VDD.n1497 GND 0.007763f
C3373 VDD.n1498 GND 0.007763f
C3374 VDD.n1499 GND 0.007763f
C3375 VDD.n1500 GND 0.006248f
C3376 VDD.n1501 GND 0.007763f
C3377 VDD.n1502 GND 0.007763f
C3378 VDD.n1503 GND 0.007763f
C3379 VDD.n1504 GND 0.007763f
C3380 VDD.n1505 GND 0.007763f
C3381 VDD.n1506 GND 0.006248f
C3382 VDD.n1507 GND 0.007763f
C3383 VDD.n1508 GND 0.007763f
C3384 VDD.n1509 GND 0.007763f
C3385 VDD.n1510 GND 0.007763f
C3386 VDD.n1511 GND 0.007763f
C3387 VDD.n1512 GND 0.006248f
C3388 VDD.n1513 GND 0.007763f
C3389 VDD.n1514 GND 0.007763f
C3390 VDD.n1515 GND 0.007763f
C3391 VDD.n1516 GND 0.007763f
C3392 VDD.n1517 GND 0.007763f
C3393 VDD.n1518 GND 0.006248f
C3394 VDD.n1519 GND 0.007763f
C3395 VDD.n1520 GND 0.007763f
C3396 VDD.n1521 GND 0.007763f
C3397 VDD.n1522 GND 0.007763f
C3398 VDD.n1523 GND 0.003405f
C3399 VDD.n1524 GND 0.007763f
C3400 VDD.n1525 GND 0.006248f
C3401 VDD.n1526 GND 0.006248f
C3402 VDD.n1527 GND 0.006248f
C3403 VDD.n1528 GND 0.007763f
C3404 VDD.n1529 GND 0.007763f
C3405 VDD.n1530 GND 0.007763f
C3406 VDD.n1531 GND 0.006248f
C3407 VDD.n1532 GND 0.006248f
C3408 VDD.n1533 GND 0.006248f
C3409 VDD.n1534 GND 0.007763f
C3410 VDD.n1535 GND 0.007763f
C3411 VDD.n1536 GND 0.007763f
C3412 VDD.n1537 GND 0.00403f
C3413 VDD.t61 GND 0.035989f
C3414 VDD.t62 GND 0.048603f
C3415 VDD.t60 GND 0.295093f
C3416 VDD.n1538 GND 0.062024f
C3417 VDD.n1539 GND 0.044734f
C3418 VDD.n1540 GND 0.009623f
C3419 VDD.n1541 GND 0.00328f
C3420 VDD.n1542 GND 0.006248f
C3421 VDD.n1543 GND 0.007763f
C3422 VDD.n1544 GND 0.007763f
C3423 VDD.n1545 GND 0.007763f
C3424 VDD.n1546 GND 0.006248f
C3425 VDD.n1547 GND 0.006248f
C3426 VDD.n1548 GND 0.006248f
C3427 VDD.n1549 GND 0.007763f
C3428 VDD.n1550 GND 0.007763f
C3429 VDD.n1551 GND 0.007763f
C3430 VDD.n1552 GND 0.006248f
C3431 VDD.n1553 GND 0.006248f
C3432 VDD.n1554 GND 0.004155f
C3433 VDD.n1555 GND 0.007763f
C3434 VDD.n1556 GND 0.007763f
C3435 VDD.n1557 GND 0.003155f
C3436 VDD.n1558 GND 0.006248f
C3437 VDD.n1559 GND 0.006248f
C3438 VDD.n1560 GND 0.007763f
C3439 VDD.n1561 GND 0.007763f
C3440 VDD.n1562 GND 0.007763f
C3441 VDD.n1563 GND 0.006248f
C3442 VDD.n1564 GND 0.006248f
C3443 VDD.n1565 GND 0.006248f
C3444 VDD.n1566 GND 0.007763f
C3445 VDD.n1567 GND 0.007763f
C3446 VDD.n1568 GND 0.007763f
C3447 VDD.n1569 GND 0.006248f
C3448 VDD.n1570 GND 0.00428f
C3449 VDD.n1571 GND 0.007763f
C3450 VDD.n1572 GND 0.007763f
C3451 VDD.t51 GND 0.035989f
C3452 VDD.t52 GND 0.048603f
C3453 VDD.t50 GND 0.295093f
C3454 VDD.n1573 GND 0.062024f
C3455 VDD.n1574 GND 0.044734f
C3456 VDD.n1575 GND 0.012747f
C3457 VDD.n1576 GND 0.007763f
C3458 VDD.n1577 GND 0.007763f
C3459 VDD.n1578 GND 0.007763f
C3460 VDD.n1579 GND 0.006248f
C3461 VDD.n1580 GND 0.006248f
C3462 VDD.n1581 GND 0.006248f
C3463 VDD.n1582 GND 0.007763f
C3464 VDD.n1583 GND 0.007763f
C3465 VDD.n1584 GND 0.007763f
C3466 VDD.n1585 GND 0.006248f
C3467 VDD.n1586 GND 0.005186f
C3468 VDD.n1587 GND 0.019093f
C3469 VDD.n1589 GND 1.39123f
C3470 VDD.n1591 GND 0.019093f
C3471 VDD.n1592 GND 0.002843f
C3472 VDD.n1593 GND 0.019093f
C3473 VDD.n1594 GND 0.018791f
C3474 VDD.n1595 GND 0.007763f
C3475 VDD.n1596 GND 0.006248f
C3476 VDD.n1597 GND 0.007763f
C3477 VDD.n1598 GND 0.594542f
C3478 VDD.n1599 GND 0.007763f
C3479 VDD.n1600 GND 0.006248f
C3480 VDD.n1601 GND 0.007763f
C3481 VDD.n1602 GND 0.007763f
C3482 VDD.n1603 GND 0.007763f
C3483 VDD.n1604 GND 0.006248f
C3484 VDD.n1605 GND 0.007763f
C3485 VDD.n1606 GND 0.594542f
C3486 VDD.n1607 GND 0.007763f
C3487 VDD.n1608 GND 0.006248f
C3488 VDD.n1609 GND 0.007763f
C3489 VDD.n1610 GND 0.007763f
C3490 VDD.n1611 GND 0.007763f
C3491 VDD.n1612 GND 0.006248f
C3492 VDD.n1613 GND 0.007763f
C3493 VDD.n1614 GND 0.594542f
C3494 VDD.n1615 GND 0.007763f
C3495 VDD.n1616 GND 0.006248f
C3496 VDD.n1617 GND 0.007763f
C3497 VDD.n1618 GND 0.007763f
C3498 VDD.n1619 GND 0.007763f
C3499 VDD.n1620 GND 0.006248f
C3500 VDD.n1621 GND 0.007763f
C3501 VDD.n1622 GND 0.594542f
C3502 VDD.n1623 GND 0.007763f
C3503 VDD.n1624 GND 0.006248f
C3504 VDD.n1625 GND 0.007763f
C3505 VDD.n1626 GND 0.007763f
C3506 VDD.n1627 GND 0.007763f
C3507 VDD.n1628 GND 0.006248f
C3508 VDD.n1629 GND 0.007763f
C3509 VDD.n1630 GND 0.594542f
C3510 VDD.n1631 GND 0.007763f
C3511 VDD.n1632 GND 0.006248f
C3512 VDD.n1633 GND 0.007763f
C3513 VDD.n1634 GND 0.007763f
C3514 VDD.n1635 GND 0.007763f
C3515 VDD.n1636 GND 0.006248f
C3516 VDD.n1637 GND 0.007763f
C3517 VDD.n1638 GND 0.594542f
C3518 VDD.n1639 GND 0.007763f
C3519 VDD.n1640 GND 0.006248f
C3520 VDD.n1641 GND 0.007763f
C3521 VDD.n1642 GND 0.007763f
C3522 VDD.n1643 GND 0.007763f
C3523 VDD.n1644 GND 0.006248f
C3524 VDD.n1645 GND 0.007763f
C3525 VDD.n1646 GND 0.338889f
C3526 VDD.n1647 GND 0.594542f
C3527 VDD.n1648 GND 0.007763f
C3528 VDD.n1649 GND 0.006248f
C3529 VDD.n1650 GND 0.007763f
C3530 VDD.n1651 GND 0.007763f
C3531 VDD.n1652 GND 0.007763f
C3532 VDD.n1653 GND 0.006248f
C3533 VDD.n1654 GND 0.007763f
C3534 VDD.n1655 GND 0.552924f
C3535 VDD.n1656 GND 0.007763f
C3536 VDD.n1657 GND 0.006248f
C3537 VDD.n1658 GND 0.007763f
C3538 VDD.n1659 GND 0.007763f
C3539 VDD.n1660 GND 0.007763f
C3540 VDD.n1661 GND 0.006248f
C3541 VDD.n1662 GND 0.007763f
C3542 VDD.n1663 GND 0.594542f
C3543 VDD.n1664 GND 0.007763f
C3544 VDD.n1665 GND 0.006248f
C3545 VDD.n1666 GND 0.007763f
C3546 VDD.n1667 GND 0.007763f
C3547 VDD.n1668 GND 0.007763f
C3548 VDD.n1669 GND 0.006248f
C3549 VDD.n1670 GND 0.007763f
C3550 VDD.n1671 GND 0.594542f
C3551 VDD.n1672 GND 0.007763f
C3552 VDD.n1673 GND 0.006248f
C3553 VDD.n1674 GND 0.007763f
C3554 VDD.n1675 GND 0.007763f
C3555 VDD.n1676 GND 0.007763f
C3556 VDD.n1677 GND 0.006248f
C3557 VDD.n1678 GND 0.007763f
C3558 VDD.n1679 GND 0.326998f
C3559 VDD.n1680 GND 0.594542f
C3560 VDD.n1681 GND 0.007763f
C3561 VDD.n1682 GND 0.006248f
C3562 VDD.n1683 GND 0.007763f
C3563 VDD.n1684 GND 0.007763f
C3564 VDD.n1685 GND 0.007763f
C3565 VDD.n1686 GND 0.006248f
C3566 VDD.n1687 GND 0.007763f
C3567 VDD.n1688 GND 0.564815f
C3568 VDD.n1689 GND 0.007763f
C3569 VDD.n1690 GND 0.006248f
C3570 VDD.n1691 GND 0.007763f
C3571 VDD.n1692 GND 0.007763f
C3572 VDD.n1693 GND 0.007763f
C3573 VDD.n1694 GND 0.006248f
C3574 VDD.n1695 GND 0.007763f
C3575 VDD.n1696 GND 0.594542f
C3576 VDD.n1697 GND 0.007763f
C3577 VDD.n1698 GND 0.006248f
C3578 VDD.n1699 GND 0.007763f
C3579 VDD.n1700 GND 0.007763f
C3580 VDD.n1701 GND 0.007763f
C3581 VDD.n1702 GND 0.006248f
C3582 VDD.n1703 GND 0.007763f
C3583 VDD.n1704 GND 0.594542f
C3584 VDD.n1705 GND 0.007763f
C3585 VDD.n1706 GND 0.006248f
C3586 VDD.n1707 GND 0.007763f
C3587 VDD.n1708 GND 0.007763f
C3588 VDD.n1709 GND 0.007763f
C3589 VDD.n1710 GND 0.006248f
C3590 VDD.n1711 GND 0.007763f
C3591 VDD.n1712 GND 0.315107f
C3592 VDD.n1713 GND 0.594542f
C3593 VDD.n1714 GND 0.007763f
C3594 VDD.n1715 GND 0.006248f
C3595 VDD.n1716 GND 0.007763f
C3596 VDD.n1717 GND 0.007763f
C3597 VDD.n1718 GND 0.007763f
C3598 VDD.n1719 GND 0.006248f
C3599 VDD.n1720 GND 0.007763f
C3600 VDD.n1721 GND 0.576706f
C3601 VDD.n1722 GND 0.007763f
C3602 VDD.n1723 GND 0.006248f
C3603 VDD.n1724 GND 0.007763f
C3604 VDD.n1725 GND 0.007763f
C3605 VDD.n1726 GND 0.007763f
C3606 VDD.n1727 GND 0.006248f
C3607 VDD.n1728 GND 0.007763f
C3608 VDD.n1729 GND 0.594542f
C3609 VDD.n1730 GND 0.007763f
C3610 VDD.n1731 GND 0.006248f
C3611 VDD.n1732 GND 0.007763f
C3612 VDD.n1733 GND 0.007763f
C3613 VDD.n1734 GND 0.007763f
C3614 VDD.n1735 GND 0.006248f
C3615 VDD.n1736 GND 0.007763f
C3616 VDD.n1737 GND 0.594542f
C3617 VDD.n1738 GND 0.007763f
C3618 VDD.n1739 GND 0.006248f
C3619 VDD.n1740 GND 0.007763f
C3620 VDD.n1741 GND 0.007763f
C3621 VDD.n1742 GND 0.007763f
C3622 VDD.n1743 GND 0.006248f
C3623 VDD.n1744 GND 0.007763f
C3624 VDD.n1745 GND 0.303217f
C3625 VDD.n1746 GND 0.594542f
C3626 VDD.n1747 GND 0.007763f
C3627 VDD.n1748 GND 0.006248f
C3628 VDD.n1749 GND 0.007763f
C3629 VDD.n1750 GND 0.007763f
C3630 VDD.n1751 GND 0.007763f
C3631 VDD.n1752 GND 0.006248f
C3632 VDD.n1753 GND 0.007763f
C3633 VDD.n1754 GND 0.588597f
C3634 VDD.n1755 GND 0.007763f
C3635 VDD.n1756 GND 0.006248f
C3636 VDD.n1757 GND 0.007763f
C3637 VDD.n1758 GND 0.007763f
C3638 VDD.n1759 GND 0.007763f
C3639 VDD.n1760 GND 0.006248f
C3640 VDD.n1761 GND 0.007763f
C3641 VDD.n1762 GND 0.594542f
C3642 VDD.n1763 GND 0.007763f
C3643 VDD.n1764 GND 0.006248f
C3644 VDD.n1765 GND 0.007736f
C3645 VDD.t166 GND 0.044552f
C3646 VDD.t143 GND 0.006779f
C3647 VDD.t150 GND 0.006779f
C3648 VDD.n1766 GND 0.028116f
C3649 VDD.n1767 GND 0.353268f
C3650 VDD.t163 GND 0.006779f
C3651 VDD.t183 GND 0.006779f
C3652 VDD.n1768 GND 0.028116f
C3653 VDD.n1769 GND 0.217723f
C3654 VDD.t186 GND 0.006779f
C3655 VDD.t193 GND 0.006779f
C3656 VDD.n1770 GND 0.028116f
C3657 VDD.n1771 GND 0.217723f
C3658 VDD.t178 GND 0.043241f
C3659 VDD.n1772 GND 0.17012f
C3660 VDD.t132 GND 0.044552f
C3661 VDD.t188 GND 0.006779f
C3662 VDD.t195 GND 0.006779f
C3663 VDD.n1773 GND 0.028116f
C3664 VDD.n1774 GND 0.353268f
C3665 VDD.t123 GND 0.006779f
C3666 VDD.t160 GND 0.006779f
C3667 VDD.n1775 GND 0.028116f
C3668 VDD.n1776 GND 0.217723f
C3669 VDD.t168 GND 0.006779f
C3670 VDD.t175 GND 0.006779f
C3671 VDD.n1777 GND 0.028116f
C3672 VDD.n1778 GND 0.217723f
C3673 VDD.t164 GND 0.043241f
C3674 VDD.n1779 GND 0.158808f
C3675 VDD.n1780 GND 0.160142f
C3676 VDD.t119 GND 0.044552f
C3677 VDD.t192 GND 0.006779f
C3678 VDD.t161 GND 0.006779f
C3679 VDD.n1781 GND 0.028116f
C3680 VDD.n1782 GND 0.353268f
C3681 VDD.t152 GND 0.006779f
C3682 VDD.t176 GND 0.006779f
C3683 VDD.n1783 GND 0.028116f
C3684 VDD.n1784 GND 0.217723f
C3685 VDD.t157 GND 0.006779f
C3686 VDD.t196 GND 0.006779f
C3687 VDD.n1785 GND 0.028116f
C3688 VDD.n1786 GND 0.217723f
C3689 VDD.t189 GND 0.043241f
C3690 VDD.n1787 GND 0.158808f
C3691 VDD.n1788 GND 0.11093f
C3692 VDD.t165 GND 0.044552f
C3693 VDD.t153 GND 0.006779f
C3694 VDD.t185 GND 0.006779f
C3695 VDD.n1789 GND 0.028116f
C3696 VDD.n1790 GND 0.353268f
C3697 VDD.t126 GND 0.006779f
C3698 VDD.t125 GND 0.006779f
C3699 VDD.n1791 GND 0.028116f
C3700 VDD.n1792 GND 0.217723f
C3701 VDD.t180 GND 0.006779f
C3702 VDD.t155 GND 0.006779f
C3703 VDD.n1793 GND 0.028116f
C3704 VDD.n1794 GND 0.217723f
C3705 VDD.t148 GND 0.043241f
C3706 VDD.n1795 GND 0.158808f
C3707 VDD.n1796 GND 0.308941f
C3708 VDD.n1797 GND 3.56029f
C3709 VDD.n1798 GND 0.542227f
C3710 VDD.n1799 GND 0.007736f
C3711 VDD.n1800 GND 0.006248f
C3712 VDD.n1801 GND 0.007763f
C3713 VDD.n1802 GND 0.594542f
C3714 VDD.n1803 GND 0.007763f
C3715 VDD.n1804 GND 0.006248f
C3716 VDD.n1805 GND 0.007763f
C3717 VDD.n1806 GND 0.007763f
C3718 VDD.n1807 GND 0.007763f
C3719 VDD.n1808 GND 0.006248f
C3720 VDD.n1809 GND 0.007763f
C3721 VDD.t124 GND 0.297271f
C3722 VDD.n1810 GND 0.588597f
C3723 VDD.n1811 GND 0.007763f
C3724 VDD.n1812 GND 0.006248f
C3725 VDD.n1813 GND 0.007763f
C3726 VDD.n1814 GND 0.007763f
C3727 VDD.n1815 GND 0.007763f
C3728 VDD.n1816 GND 0.006248f
C3729 VDD.n1817 GND 0.007763f
C3730 VDD.n1818 GND 0.594542f
C3731 VDD.n1819 GND 0.007763f
C3732 VDD.n1820 GND 0.006248f
C3733 VDD.n1821 GND 0.007763f
C3734 VDD.n1822 GND 0.007763f
C3735 VDD.n1823 GND 0.007763f
C3736 VDD.n1824 GND 0.006248f
C3737 VDD.n1825 GND 0.007763f
C3738 VDD.n1826 GND 0.594542f
C3739 VDD.n1827 GND 0.007763f
C3740 VDD.n1828 GND 0.006248f
C3741 VDD.n1829 GND 0.007763f
C3742 VDD.n1830 GND 0.007763f
C3743 VDD.n1831 GND 0.007763f
C3744 VDD.n1832 GND 0.006248f
C3745 VDD.n1833 GND 0.007763f
C3746 VDD.n1834 GND 0.594542f
C3747 VDD.n1835 GND 0.007763f
C3748 VDD.n1836 GND 0.006248f
C3749 VDD.n1837 GND 0.007763f
C3750 VDD.n1838 GND 0.007763f
C3751 VDD.n1839 GND 0.007763f
C3752 VDD.n1840 GND 0.006248f
C3753 VDD.n1841 GND 0.007763f
C3754 VDD.t142 GND 0.297271f
C3755 VDD.n1842 GND 0.576706f
C3756 VDD.n1843 GND 0.007763f
C3757 VDD.n1844 GND 0.006248f
C3758 VDD.n1845 GND 0.007763f
C3759 VDD.n1846 GND 0.007763f
C3760 VDD.n1847 GND 0.007763f
C3761 VDD.n1848 GND 0.006248f
C3762 VDD.n1849 GND 0.007763f
C3763 VDD.n1850 GND 0.594542f
C3764 VDD.n1851 GND 0.007763f
C3765 VDD.n1852 GND 0.006248f
C3766 VDD.n1853 GND 0.007763f
C3767 VDD.n1854 GND 0.007763f
C3768 VDD.n1855 GND 0.007763f
C3769 VDD.n1856 GND 0.006248f
C3770 VDD.n1857 GND 0.007763f
C3771 VDD.n1858 GND 0.594542f
C3772 VDD.n1859 GND 0.007763f
C3773 VDD.n1860 GND 0.006248f
C3774 VDD.n1861 GND 0.007763f
C3775 VDD.n1862 GND 0.007763f
C3776 VDD.n1863 GND 0.007763f
C3777 VDD.n1864 GND 0.006248f
C3778 VDD.n1865 GND 0.007763f
C3779 VDD.n1866 GND 0.594542f
C3780 VDD.n1867 GND 0.007763f
C3781 VDD.n1868 GND 0.006248f
C3782 VDD.n1869 GND 0.007763f
C3783 VDD.n1870 GND 0.007763f
C3784 VDD.n1871 GND 0.007763f
C3785 VDD.n1872 GND 0.006248f
C3786 VDD.n1873 GND 0.007763f
C3787 VDD.t149 GND 0.297271f
C3788 VDD.n1874 GND 0.564815f
C3789 VDD.n1875 GND 0.007763f
C3790 VDD.n1876 GND 0.006248f
C3791 VDD.n1877 GND 0.007763f
C3792 VDD.n1878 GND 0.007763f
C3793 VDD.n1879 GND 0.007763f
C3794 VDD.n1880 GND 0.006248f
C3795 VDD.n1881 GND 0.007763f
C3796 VDD.n1882 GND 0.594542f
C3797 VDD.n1883 GND 0.007763f
C3798 VDD.n1884 GND 0.006248f
C3799 VDD.n1885 GND 0.007763f
C3800 VDD.n1886 GND 0.007763f
C3801 VDD.n1887 GND 0.007763f
C3802 VDD.n1888 GND 0.006248f
C3803 VDD.n1889 GND 0.007763f
C3804 VDD.n1890 GND 0.594542f
C3805 VDD.n1891 GND 0.007763f
C3806 VDD.n1892 GND 0.006248f
C3807 VDD.n1893 GND 0.007763f
C3808 VDD.n1894 GND 0.007763f
C3809 VDD.n1895 GND 0.007763f
C3810 VDD.n1896 GND 0.006248f
C3811 VDD.n1897 GND 0.007763f
C3812 VDD.n1898 GND 0.594542f
C3813 VDD.n1899 GND 0.007763f
C3814 VDD.n1900 GND 0.006248f
C3815 VDD.n1901 GND 0.007763f
C3816 VDD.n1902 GND 0.007763f
C3817 VDD.n1903 GND 0.007763f
C3818 VDD.n1904 GND 0.006248f
C3819 VDD.n1905 GND 0.007763f
C3820 VDD.t118 GND 0.297271f
C3821 VDD.n1906 GND 0.552924f
C3822 VDD.n1907 GND 0.007763f
C3823 VDD.n1908 GND 0.006248f
C3824 VDD.n1909 GND 0.007763f
C3825 VDD.n1910 GND 0.007763f
C3826 VDD.n1911 GND 0.007763f
C3827 VDD.n1912 GND 0.006248f
C3828 VDD.n1913 GND 0.007763f
C3829 VDD.n1914 GND 0.594542f
C3830 VDD.n1915 GND 0.007763f
C3831 VDD.n1916 GND 0.006248f
C3832 VDD.n1917 GND 0.007763f
C3833 VDD.n1918 GND 0.007763f
C3834 VDD.n1919 GND 0.007763f
C3835 VDD.n1920 GND 0.006248f
C3836 VDD.n1921 GND 0.007763f
C3837 VDD.n1922 GND 0.594542f
C3838 VDD.n1923 GND 0.007763f
C3839 VDD.n1924 GND 0.006248f
C3840 VDD.n1925 GND 0.007763f
C3841 VDD.n1926 GND 0.007763f
C3842 VDD.n1927 GND 0.007763f
C3843 VDD.n1928 GND 0.006248f
C3844 VDD.n1929 GND 0.007763f
C3845 VDD.n1930 GND 0.594542f
C3846 VDD.n1931 GND 0.007763f
C3847 VDD.n1932 GND 0.006248f
C3848 VDD.n1933 GND 0.007763f
C3849 VDD.n1934 GND 0.007763f
C3850 VDD.n1935 GND 0.007763f
C3851 VDD.n1936 GND 0.006248f
C3852 VDD.n1937 GND 0.007763f
C3853 VDD.n1938 GND 0.594542f
C3854 VDD.n1939 GND 0.007763f
C3855 VDD.n1940 GND 0.006248f
C3856 VDD.n1941 GND 0.007763f
C3857 VDD.n1942 GND 0.007763f
C3858 VDD.n1943 GND 0.007763f
C3859 VDD.n1944 GND 0.006248f
C3860 VDD.n1945 GND 0.007763f
C3861 VDD.n1946 GND 0.594542f
C3862 VDD.n1947 GND 0.007763f
C3863 VDD.n1948 GND 0.006248f
C3864 VDD.n1949 GND 0.007763f
C3865 VDD.n1950 GND 0.007763f
C3866 VDD.n1951 GND 0.007763f
C3867 VDD.n1952 GND 0.007763f
C3868 VDD.n1953 GND 0.006248f
C3869 VDD.n1954 GND 0.007763f
C3870 VDD.n1955 GND 0.594542f
C3871 VDD.n1956 GND 0.007763f
C3872 VDD.n1957 GND 0.006248f
C3873 VDD.n1958 GND 0.007763f
C3874 VDD.n1959 GND 0.007763f
C3875 VDD.n1960 GND 0.007763f
C3876 VDD.n1961 GND 0.005186f
C3877 VDD.n1962 GND 0.006248f
C3878 VDD.n1963 GND 0.007763f
C3879 VDD.n1964 GND 0.594542f
C3880 VDD.n1965 GND 0.007763f
C3881 VDD.n1966 GND 0.018791f
C3882 VDD.n1967 GND 0.005186f
C3883 VDD.n1968 GND 0.010389f
C3884 VDD.n1969 GND 0.005279f
C3885 VDD.n1970 GND 0.005279f
C3886 VDD.n1971 GND 0.005279f
C3887 VDD.n1972 GND 0.005279f
C3888 VDD.n1973 GND 0.005279f
C3889 VDD.n1974 GND 0.005279f
C3890 VDD.n1975 GND 0.005279f
C3891 VDD.n1976 GND 0.005279f
C3892 VDD.n1977 GND 0.005279f
C3893 VDD.n1978 GND 0.005279f
C3894 VDD.n1979 GND 0.005279f
C3895 VDD.n1980 GND 0.005279f
C3896 VDD.n1981 GND 0.005279f
C3897 VDD.n1982 GND 0.005279f
C3898 VDD.n1983 GND 0.005279f
C3899 VDD.n1984 GND 0.005279f
C3900 VDD.n1985 GND 0.005279f
C3901 VDD.n1986 GND 0.005279f
C3902 VDD.n1987 GND 0.005279f
C3903 VDD.n1988 GND 0.003959f
C3904 VDD.t6 GND 0.118717f
C3905 VDD.t7 GND 0.138462f
C3906 VDD.t4 GND 0.726908f
C3907 VDD.n1989 GND 0.089246f
C3908 VDD.n1990 GND 0.051676f
C3909 VDD.n1991 GND 0.007544f
C3910 VDD.n1992 GND 0.005279f
C3911 VDD.n1993 GND 0.005279f
C3912 VDD.n1994 GND 0.005279f
C3913 VDD.n1995 GND 0.005279f
C3914 VDD.n1996 GND 0.005279f
C3915 VDD.n1997 GND 0.005279f
C3916 VDD.n1998 GND 0.005279f
C3917 VDD.n1999 GND 0.005279f
C3918 VDD.n2000 GND 0.005279f
C3919 VDD.n2001 GND 0.005279f
C3920 VDD.n2002 GND 0.005279f
C3921 VDD.n2003 GND 0.005279f
C3922 VDD.n2004 GND 0.005279f
C3923 VDD.n2005 GND 0.005279f
C3924 VDD.n2006 GND 0.005279f
C3925 VDD.n2007 GND 0.005279f
C3926 VDD.n2008 GND 0.005279f
C3927 VDD.n2009 GND 0.005279f
C3928 VDD.n2010 GND 0.005279f
C3929 VDD.n2011 GND 0.005279f
C3930 VDD.n2012 GND 0.005279f
C3931 VDD.n2013 GND 0.005279f
C3932 VDD.n2014 GND 0.005279f
C3933 VDD.n2015 GND 0.005279f
C3934 VDD.n2016 GND 0.005279f
C3935 VDD.n2017 GND 0.005279f
C3936 VDD.n2018 GND 0.005279f
C3937 VDD.n2019 GND 0.005279f
C3938 VDD.n2020 GND 0.005279f
C3939 VDD.n2021 GND 0.005279f
C3940 VDD.n2022 GND 0.005279f
C3941 VDD.n2023 GND 0.005279f
C3942 VDD.n2024 GND 0.005279f
C3943 VDD.n2025 GND 0.005279f
C3944 VDD.n2026 GND 0.005279f
C3945 VDD.n2027 GND 0.005279f
C3946 VDD.n2028 GND 0.005279f
C3947 VDD.n2029 GND 0.005279f
C3948 VDD.n2030 GND 0.005279f
C3949 VDD.n2031 GND 0.005279f
C3950 VDD.n2032 GND 0.005279f
C3951 VDD.n2033 GND 0.005279f
C3952 VDD.n2034 GND 0.005279f
C3953 VDD.n2035 GND 0.005279f
C3954 VDD.n2036 GND 0.005279f
C3955 VDD.n2037 GND 0.005279f
C3956 VDD.n2038 GND 0.005279f
C3957 VDD.n2039 GND 0.005279f
C3958 VDD.n2040 GND 0.005279f
C3959 VDD.n2041 GND 0.005279f
C3960 VDD.n2042 GND 0.005279f
C3961 VDD.n2043 GND 0.005279f
C3962 VDD.n2044 GND 0.005279f
C3963 VDD.n2045 GND 0.005279f
C3964 VDD.n2046 GND 0.005279f
C3965 VDD.n2047 GND 0.005279f
C3966 VDD.n2048 GND 0.005279f
C3967 VDD.n2049 GND 0.005279f
C3968 VDD.n2050 GND 0.005279f
C3969 VDD.n2051 GND 0.005279f
C3970 VDD.n2052 GND 0.005279f
C3971 VDD.n2053 GND 0.005279f
C3972 VDD.n2054 GND 0.013069f
C3973 VDD.n2055 GND 0.013069f
C3974 VDD.n2056 GND 0.013559f
C3975 VDD.n2057 GND 0.005279f
C3976 VDD.n2058 GND 0.005279f
C3977 VDD.n2059 GND 0.003144f
C3978 VDD.n2060 GND 0.005279f
C3979 VDD.n2061 GND 0.005279f
C3980 VDD.n2062 GND 0.004774f
C3981 VDD.n2063 GND 0.005279f
C3982 VDD.n2064 GND 0.005279f
C3983 VDD.n2065 GND 0.005279f
C3984 VDD.n2066 GND 0.005279f
C3985 VDD.n2067 GND 0.005279f
C3986 VDD.n2068 GND 0.005279f
C3987 VDD.n2069 GND 0.005279f
C3988 VDD.n2070 GND 0.005279f
C3989 VDD.n2071 GND 0.005279f
C3990 VDD.n2072 GND 0.005279f
C3991 VDD.n2073 GND 0.005279f
C3992 VDD.n2074 GND 0.005279f
C3993 VDD.n2075 GND 0.005279f
C3994 VDD.n2076 GND 0.005279f
C3995 VDD.n2077 GND 0.005279f
C3996 VDD.n2078 GND 0.003959f
C3997 VDD.n2079 GND 0.034761f
C3998 VDD.n2080 GND 0.853768f
C3999 VDD.n2081 GND 0.002843f
C4000 VDD.t71 GND 0.035989f
C4001 VDD.t70 GND 0.048603f
C4002 VDD.t69 GND 0.295093f
C4003 VDD.n2082 GND 0.062024f
C4004 VDD.n2083 GND 0.044734f
C4005 VDD.n2084 GND 0.009623f
C4006 VDD.n2085 GND 0.003405f
C4007 VDD.n2086 GND 0.007763f
C4008 VDD.n2087 GND 0.007763f
C4009 VDD.n2088 GND 0.006248f
C4010 VDD.n2089 GND 0.006248f
C4011 VDD.n2090 GND 0.007763f
C4012 VDD.n2091 GND 0.007763f
C4013 VDD.n2092 GND 0.006248f
C4014 VDD.n2093 GND 0.006248f
C4015 VDD.n2094 GND 0.007763f
C4016 VDD.n2095 GND 0.007763f
C4017 VDD.n2096 GND 0.006248f
C4018 VDD.n2097 GND 0.006248f
C4019 VDD.n2098 GND 0.007763f
C4020 VDD.n2099 GND 0.007763f
C4021 VDD.n2100 GND 0.006248f
C4022 VDD.n2101 GND 0.006248f
C4023 VDD.n2102 GND 0.007763f
C4024 VDD.n2103 GND 0.007763f
C4025 VDD.n2104 GND 0.00403f
C4026 VDD.t49 GND 0.035989f
C4027 VDD.t48 GND 0.048603f
C4028 VDD.t47 GND 0.295093f
C4029 VDD.n2105 GND 0.062024f
C4030 VDD.n2106 GND 0.044734f
C4031 VDD.n2107 GND 0.009623f
C4032 VDD.n2108 GND 0.00328f
C4033 VDD.n2109 GND 0.007763f
C4034 VDD.n2110 GND 0.007763f
C4035 VDD.n2111 GND 0.006248f
C4036 VDD.n2112 GND 0.006248f
C4037 VDD.n2113 GND 0.007763f
C4038 VDD.n2114 GND 0.007763f
C4039 VDD.n2115 GND 0.006248f
C4040 VDD.n2116 GND 0.006248f
C4041 VDD.n2117 GND 0.007763f
C4042 VDD.n2118 GND 0.007763f
C4043 VDD.n2119 GND 0.006248f
C4044 VDD.n2120 GND 0.006248f
C4045 VDD.n2121 GND 0.007763f
C4046 VDD.n2122 GND 0.007763f
C4047 VDD.n2123 GND 0.006248f
C4048 VDD.n2124 GND 0.006248f
C4049 VDD.n2125 GND 0.007763f
C4050 VDD.n2126 GND 0.007763f
C4051 VDD.n2127 GND 0.004155f
C4052 VDD.t74 GND 0.035989f
C4053 VDD.t73 GND 0.048603f
C4054 VDD.t72 GND 0.295093f
C4055 VDD.n2128 GND 0.062024f
C4056 VDD.n2129 GND 0.044734f
C4057 VDD.n2130 GND 0.009623f
C4058 VDD.n2131 GND 0.003155f
C4059 VDD.n2132 GND 0.007763f
C4060 VDD.n2133 GND 0.007763f
C4061 VDD.n2134 GND 0.006248f
C4062 VDD.n2135 GND 0.006248f
C4063 VDD.n2136 GND 0.007763f
C4064 VDD.n2137 GND 0.007763f
C4065 VDD.n2138 GND 0.006248f
C4066 VDD.n2139 GND 0.006248f
C4067 VDD.n2140 GND 0.007763f
C4068 VDD.n2141 GND 0.007763f
C4069 VDD.n2142 GND 0.006248f
C4070 VDD.n2143 GND 0.006248f
C4071 VDD.n2144 GND 0.007763f
C4072 VDD.n2145 GND 0.007763f
C4073 VDD.n2146 GND 0.006248f
C4074 VDD.n2147 GND 0.007763f
C4075 VDD.n2148 GND 0.007763f
C4076 VDD.n2149 GND 0.006248f
C4077 VDD.n2150 GND 0.007763f
C4078 VDD.n2151 GND 0.007763f
C4079 VDD.n2152 GND 0.007763f
C4080 VDD.n2153 GND 0.012747f
C4081 VDD.n2154 GND 0.007763f
C4082 VDD.n2155 GND 0.007763f
C4083 VDD.n2156 GND 0.006155f
C4084 VDD.n2157 GND 0.006248f
C4085 VDD.n2158 GND 0.007763f
C4086 VDD.n2159 GND 0.007763f
C4087 VDD.n2160 GND 0.006248f
C4088 VDD.n2161 GND 0.006248f
C4089 VDD.n2162 GND 0.006248f
C4090 VDD.n2163 GND 0.007763f
C4091 VDD.n2165 GND 4.25098f
C4092 VDD.n2166 GND 0.019093f
C4093 VDD.n2167 GND 0.005186f
C4094 VDD.n2168 GND 0.265852f
C4095 VDD.n2169 GND 0.017859f
C4096 VDD.n2170 GND 0.003959f
C4097 VDD.n2171 GND 0.005279f
C4098 VDD.n2172 GND 0.005279f
C4099 VDD.n2173 GND 0.005279f
C4100 VDD.n2174 GND 0.005279f
C4101 VDD.n2175 GND 0.005279f
C4102 VDD.n2176 GND 0.005279f
C4103 VDD.n2177 GND 0.005279f
C4104 VDD.n2178 GND 0.005279f
C4105 VDD.n2179 GND 0.005279f
C4106 VDD.n2180 GND 0.005279f
C4107 VDD.n2181 GND 0.005279f
C4108 VDD.n2182 GND 0.005279f
C4109 VDD.n2183 GND 0.005279f
C4110 VDD.n2184 GND 0.005279f
C4111 VDD.n2185 GND 0.005279f
C4112 VDD.n2186 GND 0.005279f
C4113 VDD.n2187 GND 0.005279f
C4114 VDD.n2188 GND 0.005279f
C4115 VDD.n2189 GND 0.005279f
C4116 VDD.n2190 GND 0.013559f
C4117 VDD.n2191 GND 0.013559f
C4118 VDD.n2193 GND 0.597515f
C4119 VDD.n2194 GND 0.013559f
C4120 VDD.n2195 GND 0.013559f
C4121 VDD.n2196 GND 0.013069f
C4122 VDD.n2197 GND 0.005279f
C4123 VDD.n2198 GND 0.005279f
C4124 VDD.n2199 GND 0.404289f
C4125 VDD.n2200 GND 0.005279f
C4126 VDD.n2201 GND 0.005279f
C4127 VDD.n2202 GND 0.005279f
C4128 VDD.n2203 GND 0.005279f
C4129 VDD.n2204 GND 0.005279f
C4130 VDD.n2205 GND 0.404289f
C4131 VDD.n2206 GND 0.005279f
C4132 VDD.n2207 GND 0.005279f
C4133 VDD.n2208 GND 0.005279f
C4134 VDD.n2209 GND 0.005279f
C4135 VDD.n2210 GND 0.005279f
C4136 VDD.n2211 GND 0.404289f
C4137 VDD.n2212 GND 0.005279f
C4138 VDD.n2213 GND 0.005279f
C4139 VDD.n2214 GND 0.005279f
C4140 VDD.n2215 GND 0.005279f
C4141 VDD.n2216 GND 0.005279f
C4142 VDD.n2217 GND 0.249708f
C4143 VDD.n2218 GND 0.005279f
C4144 VDD.n2219 GND 0.005279f
C4145 VDD.n2220 GND 0.005279f
C4146 VDD.n2221 GND 0.005279f
C4147 VDD.n2222 GND 0.005279f
C4148 VDD.n2223 GND 0.258626f
C4149 VDD.n2224 GND 0.005279f
C4150 VDD.n2225 GND 0.005279f
C4151 VDD.n2226 GND 0.005279f
C4152 VDD.n2227 GND 0.005279f
C4153 VDD.n2228 GND 0.005279f
C4154 VDD.n2229 GND 0.404289f
C4155 VDD.n2230 GND 0.005279f
C4156 VDD.n2231 GND 0.005279f
C4157 VDD.n2232 GND 0.005279f
C4158 VDD.n2233 GND 0.005279f
C4159 VDD.n2234 GND 0.005279f
C4160 VDD.n2235 GND 0.404289f
C4161 VDD.n2236 GND 0.005279f
C4162 VDD.n2237 GND 0.005279f
C4163 VDD.n2238 GND 0.005279f
C4164 VDD.n2239 GND 0.005279f
C4165 VDD.n2240 GND 0.005279f
C4166 VDD.n2241 GND 0.404289f
C4167 VDD.n2242 GND 0.005279f
C4168 VDD.n2243 GND 0.005279f
C4169 VDD.n2244 GND 0.005279f
C4170 VDD.n2245 GND 0.005279f
C4171 VDD.n2246 GND 0.005279f
C4172 VDD.n2247 GND 0.404289f
C4173 VDD.n2248 GND 0.005279f
C4174 VDD.n2249 GND 0.005279f
C4175 VDD.n2250 GND 0.005279f
C4176 VDD.n2251 GND 0.005279f
C4177 VDD.n2252 GND 0.005279f
C4178 VDD.n2253 GND 0.404289f
C4179 VDD.n2254 GND 0.005279f
C4180 VDD.n2255 GND 0.005279f
C4181 VDD.n2256 GND 0.005279f
C4182 VDD.n2257 GND 0.005279f
C4183 VDD.n2258 GND 0.005279f
C4184 VDD.n2259 GND 0.252681f
C4185 VDD.n2260 GND 0.005279f
C4186 VDD.n2261 GND 0.005279f
C4187 VDD.n2262 GND 0.005279f
C4188 VDD.n2263 GND 0.005279f
C4189 VDD.n2264 GND 0.005279f
C4190 VDD.n2265 GND 0.404289f
C4191 VDD.n2266 GND 0.005279f
C4192 VDD.n2267 GND 0.005279f
C4193 VDD.n2268 GND 0.005279f
C4194 VDD.n2269 GND 0.005279f
C4195 VDD.n2270 GND 0.005279f
C4196 VDD.n2271 GND 0.404289f
C4197 VDD.n2272 GND 0.005279f
C4198 VDD.n2273 GND 0.005279f
C4199 VDD.n2274 GND 0.005279f
C4200 VDD.n2275 GND 0.005279f
C4201 VDD.n2276 GND 0.005279f
C4202 VDD.n2277 GND 0.404289f
C4203 VDD.n2278 GND 0.005279f
C4204 VDD.n2279 GND 0.005279f
C4205 VDD.n2280 GND 0.005279f
C4206 VDD.n2281 GND 0.005279f
C4207 VDD.n2282 GND 0.005279f
C4208 VDD.n2283 GND 0.404289f
C4209 VDD.n2284 GND 0.005279f
C4210 VDD.n2285 GND 0.005279f
C4211 VDD.n2286 GND 0.005279f
C4212 VDD.n2287 GND 0.005279f
C4213 VDD.n2288 GND 0.005279f
C4214 VDD.n2289 GND 0.404289f
C4215 VDD.n2290 GND 0.005279f
C4216 VDD.n2291 GND 0.005279f
C4217 VDD.n2292 GND 0.005279f
C4218 VDD.n2293 GND 0.005279f
C4219 VDD.n2294 GND 0.005279f
C4220 VDD.n2295 GND 0.252681f
C4221 VDD.n2296 GND 0.005279f
C4222 VDD.n2297 GND 0.005279f
C4223 VDD.n2298 GND 0.005279f
C4224 VDD.n2299 GND 0.005279f
C4225 VDD.n2300 GND 0.005279f
C4226 VDD.n2301 GND 0.404289f
C4227 VDD.n2302 GND 0.005279f
C4228 VDD.n2303 GND 0.005279f
C4229 VDD.n2304 GND 0.005279f
C4230 VDD.n2305 GND 0.005279f
C4231 VDD.n2306 GND 0.005279f
C4232 VDD.n2307 GND 0.404289f
C4233 VDD.n2308 GND 0.005279f
C4234 VDD.n2309 GND 0.005279f
C4235 VDD.n2310 GND 0.005279f
C4236 VDD.n2311 GND 0.005279f
C4237 VDD.n2312 GND 0.005279f
C4238 VDD.n2313 GND 0.404289f
C4239 VDD.n2314 GND 0.005279f
C4240 VDD.n2315 GND 0.005279f
C4241 VDD.n2316 GND 0.005279f
C4242 VDD.n2317 GND 0.005279f
C4243 VDD.n2318 GND 0.005279f
C4244 VDD.n2319 GND 0.005279f
C4245 VDD.n2320 GND 0.005279f
C4246 VDD.n2321 GND 0.005279f
C4247 VDD.n2322 GND 0.005279f
C4248 VDD.n2323 GND 0.005279f
C4249 VDD.n2324 GND 0.404289f
C4250 VDD.n2325 GND 0.005279f
C4251 VDD.n2326 GND 0.005279f
C4252 VDD.n2327 GND 0.005279f
C4253 VDD.n2328 GND 0.005279f
C4254 VDD.n2329 GND 0.005279f
C4255 VDD.n2330 GND 0.404289f
C4256 VDD.n2331 GND 0.005279f
C4257 VDD.n2332 GND 0.005279f
C4258 VDD.n2333 GND 0.005279f
C4259 VDD.n2334 GND 0.005279f
C4260 VDD.n2335 GND 0.005279f
C4261 VDD.n2336 GND 0.005279f
C4262 VDD.n2337 GND 0.005279f
C4263 VDD.n2338 GND 0.005279f
C4264 VDD.n2339 GND 0.005279f
C4265 VDD.n2340 GND 0.005279f
C4266 VDD.n2341 GND 0.005279f
C4267 VDD.n2342 GND 0.005279f
C4268 VDD.n2343 GND 0.005279f
C4269 VDD.n2344 GND 0.005279f
C4270 VDD.n2345 GND 0.005279f
C4271 VDD.n2346 GND 0.005279f
C4272 VDD.n2347 GND 0.005279f
C4273 VDD.n2348 GND 0.005279f
C4274 VDD.n2349 GND 0.005279f
C4275 VDD.n2350 GND 0.005279f
C4276 VDD.n2351 GND 0.005279f
C4277 VDD.n2352 GND 0.005279f
C4278 VDD.n2353 GND 0.005279f
C4279 VDD.n2354 GND 0.005279f
C4280 VDD.n2355 GND 0.005279f
C4281 VDD.n2356 GND 0.005279f
C4282 VDD.n2357 GND 0.005279f
C4283 VDD.n2358 GND 0.005279f
C4284 VDD.n2359 GND 0.005279f
C4285 VDD.n2360 GND 0.005279f
C4286 VDD.n2361 GND 0.005279f
C4287 VDD.n2362 GND 0.005279f
C4288 VDD.n2363 GND 0.005279f
C4289 VDD.n2364 GND 0.005279f
C4290 VDD.n2365 GND 0.005279f
C4291 VDD.n2366 GND 0.005279f
C4292 VDD.n2367 GND 0.005279f
C4293 VDD.n2368 GND 0.005279f
C4294 VDD.n2369 GND 0.005279f
C4295 VDD.n2370 GND 0.005279f
C4296 VDD.n2371 GND 0.005279f
C4297 VDD.n2372 GND 0.005279f
C4298 VDD.n2373 GND 0.005279f
C4299 VDD.n2374 GND 0.005279f
C4300 VDD.n2375 GND 0.005279f
C4301 VDD.n2376 GND 0.005279f
C4302 VDD.n2377 GND 0.005279f
C4303 VDD.n2378 GND 0.005279f
C4304 VDD.n2379 GND 0.005279f
C4305 VDD.n2380 GND 0.005279f
C4306 VDD.n2381 GND 0.005279f
C4307 VDD.n2382 GND 0.005279f
C4308 VDD.n2383 GND 0.005279f
C4309 VDD.n2384 GND 0.005279f
C4310 VDD.n2385 GND 0.005279f
C4311 VDD.n2386 GND 0.005279f
C4312 VDD.n2387 GND 0.005279f
C4313 VDD.n2388 GND 0.005279f
C4314 VDD.n2389 GND 0.005279f
C4315 VDD.n2390 GND 0.005279f
C4316 VDD.n2391 GND 0.005279f
C4317 VDD.n2392 GND 0.005279f
C4318 VDD.n2393 GND 0.005279f
C4319 VDD.n2394 GND 0.005279f
C4320 VDD.n2395 GND 0.005279f
C4321 VDD.n2396 GND 0.005279f
C4322 VDD.n2397 GND 0.005279f
C4323 VDD.n2398 GND 0.005279f
C4324 VDD.n2399 GND 0.306189f
C4325 VDD.n2400 GND 0.005279f
C4326 VDD.n2401 GND 0.005279f
C4327 VDD.n2402 GND 0.005279f
C4328 VDD.n2403 GND 0.005279f
C4329 VDD.n2404 GND 0.005279f
C4330 VDD.n2405 GND 0.005279f
C4331 VDD.n2406 GND 0.005279f
C4332 VDD.n2407 GND 0.005279f
C4333 VDD.n2408 GND 0.005279f
C4334 VDD.n2409 GND 0.005279f
C4335 VDD.n2410 GND 0.005279f
C4336 VDD.n2411 GND 0.005279f
C4337 VDD.n2412 GND 0.005279f
C4338 VDD.n2413 GND 0.005279f
C4339 VDD.n2414 GND 0.005279f
C4340 VDD.n2415 GND 0.005279f
C4341 VDD.n2416 GND 0.005279f
C4342 VDD.n2417 GND 0.005279f
C4343 VDD.n2418 GND 0.005279f
C4344 VDD.n2419 GND 0.005279f
C4345 VDD.n2420 GND 0.005279f
C4346 VDD.n2421 GND 0.005279f
C4347 VDD.n2422 GND 0.005279f
C4348 VDD.n2423 GND 0.005279f
C4349 VDD.n2424 GND 0.005279f
C4350 VDD.n2425 GND 0.005279f
C4351 VDD.n2426 GND 0.005279f
C4352 VDD.n2427 GND 0.005279f
C4353 VDD.n2428 GND 0.005279f
C4354 VDD.n2429 GND 0.005279f
C4355 VDD.n2430 GND 0.005279f
C4356 VDD.n2431 GND 0.005279f
C4357 VDD.n2432 GND 0.005279f
C4358 VDD.n2433 GND 0.005279f
C4359 VDD.n2434 GND 0.005279f
C4360 VDD.n2435 GND 0.005279f
C4361 VDD.n2436 GND 0.005279f
C4362 VDD.n2437 GND 0.005279f
C4363 VDD.n2438 GND 0.005279f
C4364 VDD.n2439 GND 0.005279f
C4365 VDD.n2440 GND 0.005279f
C4366 VDD.n2441 GND 0.005279f
C4367 VDD.n2442 GND 0.005279f
C4368 VDD.n2443 GND 0.005279f
C4369 VDD.n2444 GND 0.005279f
C4370 VDD.n2445 GND 0.005279f
C4371 VDD.n2446 GND 0.005279f
C4372 VDD.n2447 GND 0.005279f
C4373 VDD.n2448 GND 0.005279f
C4374 VDD.n2449 GND 0.005279f
C4375 VDD.n2450 GND 0.005279f
C4376 VDD.n2451 GND 0.005279f
C4377 VDD.n2452 GND 0.005279f
C4378 VDD.n2453 GND 0.005279f
C4379 VDD.n2454 GND 0.005279f
C4380 VDD.n2455 GND 0.005279f
C4381 VDD.n2456 GND 0.005279f
C4382 VDD.n2457 GND 0.005279f
C4383 VDD.n2458 GND 0.005279f
C4384 VDD.n2459 GND 0.005279f
C4385 VDD.t100 GND 0.404289f
C4386 VDD.n2460 GND 0.005279f
C4387 VDD.n2461 GND 0.005279f
C4388 VDD.n2462 GND 0.005279f
C4389 VDD.n2463 GND 0.005279f
C4390 VDD.n2464 GND 0.005279f
C4391 VDD.n2465 GND 0.404289f
C4392 VDD.n2466 GND 0.005279f
C4393 VDD.n2467 GND 0.005279f
C4394 VDD.n2468 GND 0.005279f
C4395 VDD.n2469 GND 0.005279f
C4396 VDD.n2470 GND 0.005279f
C4397 VDD.n2471 GND 0.347807f
C4398 VDD.n2472 GND 0.005279f
C4399 VDD.n2473 GND 0.005279f
C4400 VDD.n2474 GND 0.005279f
C4401 VDD.n2475 GND 0.005279f
C4402 VDD.n2476 GND 0.005279f
C4403 VDD.n2477 GND 0.404289f
C4404 VDD.n2478 GND 0.005279f
C4405 VDD.n2479 GND 0.005279f
C4406 VDD.n2480 GND 0.005279f
C4407 VDD.n2481 GND 0.005279f
C4408 VDD.n2482 GND 0.005279f
C4409 VDD.n2483 GND 0.404289f
C4410 VDD.n2484 GND 0.005279f
C4411 VDD.n2485 GND 0.005279f
C4412 VDD.n2486 GND 0.005279f
C4413 VDD.n2487 GND 0.005279f
C4414 VDD.n2488 GND 0.005279f
C4415 VDD.n2489 GND 0.404289f
C4416 VDD.n2490 GND 0.005279f
C4417 VDD.n2491 GND 0.005279f
C4418 VDD.n2492 GND 0.005279f
C4419 VDD.n2493 GND 0.005279f
C4420 VDD.n2494 GND 0.005279f
C4421 VDD.n2495 GND 0.267544f
C4422 VDD.n2496 GND 0.005279f
C4423 VDD.n2497 GND 0.005279f
C4424 VDD.n2498 GND 0.005279f
C4425 VDD.n2499 GND 0.005279f
C4426 VDD.n2500 GND 0.005279f
C4427 VDD.n2501 GND 0.404289f
C4428 VDD.n2502 GND 0.005279f
C4429 VDD.n2503 GND 0.005279f
C4430 VDD.n2504 GND 0.005279f
C4431 VDD.n2505 GND 0.005279f
C4432 VDD.n2506 GND 0.005279f
C4433 VDD.n2507 GND 0.282408f
C4434 VDD.n2508 GND 0.005279f
C4435 VDD.n2509 GND 0.005279f
C4436 VDD.n2510 GND 0.005279f
C4437 VDD.n2511 GND 0.005279f
C4438 VDD.n2512 GND 0.005279f
C4439 VDD.n2513 GND 0.404289f
C4440 VDD.n2514 GND 0.005279f
C4441 VDD.n2515 GND 0.005279f
C4442 VDD.n2516 GND 0.005279f
C4443 VDD.n2517 GND 0.005279f
C4444 VDD.n2518 GND 0.005279f
C4445 VDD.n2519 GND 0.404289f
C4446 VDD.n2520 GND 0.005279f
C4447 VDD.n2521 GND 0.005279f
C4448 VDD.n2522 GND 0.005279f
C4449 VDD.n2523 GND 0.005279f
C4450 VDD.n2524 GND 0.005279f
C4451 VDD.n2525 GND 0.404289f
C4452 VDD.n2526 GND 0.005279f
C4453 VDD.n2527 GND 0.005279f
C4454 VDD.n2528 GND 0.005279f
C4455 VDD.n2529 GND 0.005279f
C4456 VDD.n2530 GND 0.005279f
C4457 VDD.n2531 GND 0.332944f
C4458 VDD.n2532 GND 0.005279f
C4459 VDD.n2533 GND 0.005279f
C4460 VDD.n2534 GND 0.005279f
C4461 VDD.n2535 GND 0.005279f
C4462 VDD.n2536 GND 0.005279f
C4463 VDD.n2537 GND 0.404289f
C4464 VDD.n2538 GND 0.005279f
C4465 VDD.n2539 GND 0.005279f
C4466 VDD.n2540 GND 0.005279f
C4467 VDD.n2541 GND 0.005279f
C4468 VDD.n2542 GND 0.005279f
C4469 VDD.n2543 GND 0.217008f
C4470 VDD.n2544 GND 0.005279f
C4471 VDD.n2545 GND 0.005279f
C4472 VDD.n2546 GND 0.005279f
C4473 VDD.n2547 GND 0.005279f
C4474 VDD.n2548 GND 0.005279f
C4475 VDD.n2549 GND 0.404289f
C4476 VDD.n2550 GND 0.005279f
C4477 VDD.n2551 GND 0.005279f
C4478 VDD.n2552 GND 0.005279f
C4479 VDD.n2553 GND 0.005279f
C4480 VDD.n2554 GND 0.005279f
C4481 VDD.n2555 GND 0.404289f
C4482 VDD.n2556 GND 0.005279f
C4483 VDD.n2557 GND 0.005279f
C4484 VDD.n2558 GND 0.005279f
C4485 VDD.n2559 GND 0.005279f
C4486 VDD.n2560 GND 0.005279f
C4487 VDD.n2561 GND 0.404289f
C4488 VDD.n2562 GND 0.005279f
C4489 VDD.n2563 GND 0.005279f
C4490 VDD.n2564 GND 0.005279f
C4491 VDD.n2565 GND 0.005279f
C4492 VDD.n2566 GND 0.005279f
C4493 VDD.n2567 GND 0.404289f
C4494 VDD.n2568 GND 0.005279f
C4495 VDD.n2569 GND 0.005279f
C4496 VDD.n2570 GND 0.005279f
C4497 VDD.n2571 GND 0.005279f
C4498 VDD.n2572 GND 0.005279f
C4499 VDD.n2573 GND 0.249708f
C4500 VDD.n2574 GND 0.005279f
C4501 VDD.n2575 GND 0.005279f
C4502 VDD.n2576 GND 0.005279f
C4503 VDD.n2577 GND 0.005279f
C4504 VDD.n2578 GND 0.005279f
C4505 VDD.n2579 GND 0.005279f
C4506 VDD.n2580 GND 0.005279f
C4507 VDD.n2581 GND 0.005279f
C4508 VDD.n2582 GND 0.005279f
C4509 VDD.n2583 GND 0.005279f
C4510 VDD.n2584 GND 0.252681f
C4511 VDD.n2585 GND 0.005279f
C4512 VDD.n2586 GND 0.005279f
C4513 VDD.n2587 GND 0.005279f
C4514 VDD.n2588 GND 0.005279f
C4515 VDD.n2589 GND 0.005279f
C4516 VDD.n2590 GND 0.404289f
C4517 VDD.n2591 GND 0.005279f
C4518 VDD.n2592 GND 0.005279f
C4519 VDD.n2593 GND 0.005279f
C4520 VDD.n2594 GND 0.005279f
C4521 VDD.n2595 GND 0.013627f
C4522 VDD.n2596 GND 0.013069f
C4523 VDD.n2597 GND 0.013559f
C4524 VDD.n2598 GND 0.013001f
C4525 VDD.n2599 GND 0.005279f
C4526 VDD.n2600 GND 0.005279f
C4527 VDD.n2601 GND 0.005279f
C4528 VDD.n2602 GND 0.003144f
C4529 VDD.n2603 GND 0.007544f
C4530 VDD.n2604 GND 0.004774f
C4531 VDD.n2605 GND 0.005279f
C4532 VDD.n2606 GND 0.005279f
C4533 VDD.n2607 GND 0.005279f
C4534 VDD.n2608 GND 0.005279f
C4535 VDD.n2609 GND 0.005279f
C4536 VDD.n2610 GND 0.005279f
C4537 VDD.n2611 GND 0.005279f
C4538 VDD.n2612 GND 0.005279f
C4539 VDD.n2613 GND 0.005279f
C4540 VDD.n2614 GND 0.005279f
C4541 VDD.n2615 GND 0.005279f
C4542 VDD.n2616 GND 0.005279f
C4543 VDD.n2617 GND 0.005279f
C4544 VDD.n2618 GND 0.005279f
C4545 VDD.n2619 GND 0.005279f
C4546 VDD.n2620 GND 0.005279f
C4547 VDD.n2621 GND 0.005279f
C4548 VDD.n2622 GND 0.005279f
C4549 VDD.n2623 GND 0.005279f
C4550 VDD.n2624 GND 0.005279f
C4551 VDD.n2625 GND 0.005279f
C4552 VDD.n2626 GND 0.005279f
C4553 VDD.n2627 GND 0.005279f
C4554 VDD.n2628 GND 0.005279f
C4555 VDD.n2629 GND 0.005279f
C4556 VDD.n2630 GND 0.005279f
C4557 VDD.n2631 GND 0.005279f
C4558 VDD.n2632 GND 0.005279f
C4559 VDD.n2633 GND 0.005279f
C4560 VDD.n2634 GND 0.005279f
C4561 VDD.n2635 GND 0.005279f
C4562 VDD.n2636 GND 0.005279f
C4563 VDD.n2637 GND 0.005279f
C4564 VDD.n2638 GND 0.005279f
C4565 VDD.n2639 GND 0.005279f
C4566 VDD.n2640 GND 0.005279f
C4567 VDD.n2641 GND 0.005279f
C4568 VDD.n2642 GND 0.005279f
C4569 VDD.n2643 GND 0.005279f
C4570 VDD.n2644 GND 0.013559f
C4571 VDD.n2645 GND 0.013559f
C4572 VDD.n2646 GND 0.013069f
C4573 VDD.n2647 GND 0.005279f
C4574 VDD.n2648 GND 0.005279f
C4575 VDD.n2649 GND 0.404289f
C4576 VDD.n2650 GND 0.005279f
C4577 VDD.n2651 GND 0.013069f
C4578 VDD.n2652 GND 0.013627f
C4579 VDD.n2653 GND 0.013001f
C4580 VDD.n2654 GND 0.005279f
C4581 VDD.n2655 GND 0.005279f
C4582 VDD.n2656 GND 0.003144f
C4583 VDD.n2657 GND 0.005279f
C4584 VDD.n2658 GND 0.005279f
C4585 VDD.n2659 GND 0.004774f
C4586 VDD.n2660 GND 0.005279f
C4587 VDD.n2661 GND 0.005279f
C4588 VDD.n2662 GND 0.005279f
C4589 VDD.n2663 GND 0.005279f
C4590 VDD.n2664 GND 0.005279f
C4591 VDD.n2665 GND 0.005279f
C4592 VDD.n2666 GND 0.005279f
C4593 VDD.n2667 GND 0.005279f
C4594 VDD.n2668 GND 0.005279f
C4595 VDD.n2669 GND 0.005279f
C4596 VDD.n2670 GND 0.005279f
C4597 VDD.n2671 GND 0.005279f
C4598 VDD.n2672 GND 0.005279f
C4599 VDD.n2673 GND 0.005279f
C4600 VDD.n2674 GND 0.005279f
C4601 VDD.n2675 GND 0.005279f
C4602 VDD.n2676 GND 0.005279f
C4603 VDD.n2677 GND 0.005279f
C4604 VDD.n2678 GND 0.005279f
C4605 VDD.n2679 GND 0.005279f
C4606 VDD.n2680 GND 0.005279f
C4607 VDD.n2681 GND 0.005279f
C4608 VDD.n2682 GND 0.005279f
C4609 VDD.n2683 GND 0.005279f
C4610 VDD.n2684 GND 0.005279f
C4611 VDD.n2685 GND 0.005279f
C4612 VDD.n2686 GND 0.005279f
C4613 VDD.n2687 GND 0.005279f
C4614 VDD.n2688 GND 0.005279f
C4615 VDD.n2689 GND 0.005279f
C4616 VDD.n2690 GND 0.005279f
C4617 VDD.n2691 GND 0.005279f
C4618 VDD.n2692 GND 0.005279f
C4619 VDD.n2693 GND 0.005279f
C4620 VDD.n2694 GND 0.005279f
C4621 VDD.n2695 GND 0.005279f
C4622 VDD.n2696 GND 0.005279f
C4623 VDD.n2697 GND 0.013559f
C4624 VDD.n2698 GND 0.013559f
C4625 VDD.n2699 GND 2.55951f
C4626 VDD.n2710 GND 0.013559f
C4627 VDD.n2723 GND 0.005279f
C4628 VDD.t10 GND 0.118717f
C4629 VDD.t11 GND 0.138462f
C4630 VDD.t8 GND 0.726908f
C4631 VDD.n2724 GND 0.089246f
C4632 VDD.n2725 GND 0.051676f
C4633 VDD.n2726 GND 0.007544f
C4634 VDD.n2727 GND 0.005279f
C4635 VDD.n2728 GND 0.005279f
C4636 VDD.n2729 GND 0.005279f
C4637 VDD.n2730 GND 0.005279f
C4638 VDD.n2731 GND 0.005279f
C4639 VDD.n2732 GND 0.005279f
C4640 VDD.n2733 GND 0.005279f
C4641 VDD.n2734 GND 0.005279f
C4642 VDD.n2735 GND 0.005279f
C4643 VDD.n2736 GND 0.005279f
C4644 VDD.n2737 GND 0.005279f
C4645 VDD.n2738 GND 0.005279f
C4646 VDD.n2739 GND 0.005279f
C4647 VDD.n2740 GND 0.005279f
C4648 VDD.n2741 GND 0.005279f
C4649 VDD.n2742 GND 0.005279f
C4650 VDD.n2743 GND 0.005279f
C4651 VDD.n2744 GND 0.005279f
C4652 VDD.n2745 GND 0.005279f
C4653 VDD.n2746 GND 0.005279f
C4654 VDD.n2747 GND 0.005279f
C4655 VDD.n2748 GND 0.005279f
C4656 VDD.n2749 GND 0.005279f
C4657 VDD.n2750 GND 0.005279f
C4658 VDD.n2751 GND 0.005279f
C4659 VDD.n2752 GND 0.005279f
C4660 VDD.n2753 GND 0.005279f
C4661 VDD.n2754 GND 0.005279f
C4662 VDD.n2755 GND 0.005279f
C4663 VDD.n2756 GND 0.005279f
C4664 VDD.n2757 GND 0.005279f
C4665 VDD.n2758 GND 0.005279f
C4666 VDD.n2759 GND 0.005279f
C4667 VDD.n2760 GND 0.005279f
C4668 VDD.n2761 GND 0.005279f
C4669 VDD.n2762 GND 0.005279f
C4670 VDD.n2763 GND 0.005279f
C4671 VDD.n2764 GND 0.005279f
C4672 VDD.n2765 GND 0.005279f
C4673 VDD.n2766 GND 0.005279f
C4674 VDD.n2767 GND 0.005279f
C4675 VDD.n2768 GND 0.005279f
C4676 VDD.n2769 GND 0.005279f
C4677 VDD.n2770 GND 0.005279f
C4678 VDD.n2771 GND 0.005279f
C4679 VDD.n2772 GND 0.005279f
C4680 VDD.n2773 GND 0.005279f
C4681 VDD.n2774 GND 0.005279f
C4682 VDD.n2775 GND 0.005279f
C4683 VDD.n2776 GND 0.005279f
C4684 VDD.n2777 GND 0.005279f
C4685 VDD.n2778 GND 0.005279f
C4686 VDD.n2779 GND 0.005279f
C4687 VDD.n2780 GND 0.005279f
C4688 VDD.n2781 GND 0.005279f
C4689 VDD.n2782 GND 0.005279f
C4690 VDD.n2783 GND 0.005279f
C4691 VDD.n2784 GND 0.005279f
C4692 VDD.n2785 GND 0.005279f
C4693 VDD.n2786 GND 0.005279f
C4694 VDD.n2787 GND 0.005279f
C4695 VDD.n2788 GND 0.005279f
C4696 VDD.n2789 GND 0.005279f
C4697 VDD.n2790 GND 0.005279f
C4698 VDD.n2791 GND 0.005279f
C4699 VDD.n2792 GND 0.005279f
C4700 VDD.n2793 GND 0.005279f
C4701 VDD.n2794 GND 0.005279f
C4702 VDD.n2795 GND 0.005279f
C4703 VDD.n2796 GND 0.005279f
C4704 VDD.n2797 GND 0.005279f
C4705 VDD.n2798 GND 0.005279f
C4706 VDD.n2799 GND 0.005279f
C4707 VDD.n2800 GND 0.005279f
C4708 VDD.n2801 GND 0.005279f
C4709 VDD.n2802 GND 0.005279f
C4710 VDD.n2803 GND 0.005279f
C4711 VDD.n2804 GND 0.005279f
C4712 VDD.n2805 GND 0.005279f
C4713 VDD.n2806 GND 0.005279f
C4714 VDD.n2807 GND 0.005279f
C4715 VDD.n2808 GND 0.005279f
C4716 VDD.n2809 GND 0.005279f
C4717 VDD.n2810 GND 0.005279f
C4718 VDD.n2811 GND 0.005279f
C4719 VDD.n2812 GND 0.005279f
C4720 VDD.n2813 GND 0.005279f
C4721 VDD.n2814 GND 0.005279f
C4722 VDD.n2815 GND 0.005279f
C4723 VDD.n2816 GND 0.005279f
C4724 VDD.n2817 GND 0.005279f
C4725 VDD.n2818 GND 0.005279f
C4726 VDD.n2819 GND 0.005279f
C4727 VDD.n2820 GND 0.005279f
C4728 VDD.n2821 GND 0.005279f
C4729 VDD.n2822 GND 0.005279f
C4730 VDD.n2823 GND 0.005279f
C4731 VDD.n2824 GND 0.005279f
C4732 VDD.n2825 GND 0.005279f
C4733 VDD.n2826 GND 0.005279f
C4734 VDD.n2827 GND 0.005279f
C4735 VDD.n2828 GND 0.005279f
C4736 VDD.n2829 GND 0.005279f
C4737 VDD.n2830 GND 0.005279f
C4738 VDD.n2831 GND 0.005279f
C4739 VDD.n2832 GND 0.005279f
C4740 VDD.n2833 GND 0.005279f
C4741 VDD.n2834 GND 0.005279f
C4742 VDD.n2835 GND 0.005279f
C4743 VDD.n2836 GND 0.005279f
C4744 VDD.n2837 GND 0.005279f
C4745 VDD.n2838 GND 0.005279f
C4746 VDD.n2839 GND 0.005279f
C4747 VDD.n2840 GND 0.005279f
C4748 VDD.n2841 GND 0.005279f
C4749 VDD.n2842 GND 0.005279f
C4750 VDD.n2843 GND 0.005279f
C4751 VDD.n2844 GND 0.005279f
C4752 VDD.n2845 GND 0.005279f
C4753 VDD.n2846 GND 0.005279f
C4754 VDD.n2847 GND 0.005279f
C4755 VDD.t76 GND 0.118717f
C4756 VDD.t77 GND 0.138462f
C4757 VDD.t75 GND 0.726908f
C4758 VDD.n2848 GND 0.089246f
C4759 VDD.n2849 GND 0.051676f
C4760 VDD.n2850 GND 0.013559f
C4761 VDD.n2851 GND 0.013559f
C4762 VDD.n2852 GND 0.005279f
C4763 VDD.n2853 GND 0.005279f
C4764 VDD.n2854 GND 0.005279f
C4765 VDD.n2855 GND 0.005279f
C4766 VDD.n2856 GND 0.005279f
C4767 VDD.n2857 GND 0.005279f
C4768 VDD.n2858 GND 0.005279f
C4769 VDD.n2859 GND 0.005279f
C4770 VDD.n2860 GND 0.005279f
C4771 VDD.n2861 GND 0.005279f
C4772 VDD.n2862 GND 0.005279f
C4773 VDD.n2863 GND 0.005279f
C4774 VDD.n2864 GND 0.005279f
C4775 VDD.n2865 GND 0.005279f
C4776 VDD.n2866 GND 0.005279f
C4777 VDD.n2867 GND 0.005279f
C4778 VDD.n2868 GND 0.005279f
C4779 VDD.n2869 GND 0.005279f
C4780 VDD.n2870 GND 0.005279f
C4781 VDD.n2871 GND 0.005279f
C4782 VDD.n2872 GND 0.005279f
C4783 VDD.n2873 GND 0.005279f
C4784 VDD.n2874 GND 0.005279f
C4785 VDD.n2875 GND 0.005279f
C4786 VDD.n2876 GND 0.005279f
C4787 VDD.n2877 GND 0.005279f
C4788 VDD.n2878 GND 0.005279f
C4789 VDD.n2879 GND 0.005279f
C4790 VDD.n2880 GND 0.005279f
C4791 VDD.n2881 GND 0.005279f
C4792 VDD.n2882 GND 0.005279f
C4793 VDD.n2883 GND 0.005279f
C4794 VDD.n2884 GND 0.005279f
C4795 VDD.n2885 GND 0.005279f
C4796 VDD.n2886 GND 0.005279f
C4797 VDD.n2887 GND 0.005279f
C4798 VDD.n2888 GND 0.005279f
C4799 VDD.n2889 GND 0.005279f
C4800 VDD.n2890 GND 0.005279f
C4801 VDD.n2891 GND 0.004774f
C4802 VDD.n2892 GND 0.007544f
C4803 VDD.n2893 GND 0.003144f
C4804 VDD.n2894 GND 0.005279f
C4805 VDD.n2895 GND 0.005279f
C4806 VDD.n2896 GND 0.005279f
C4807 VDD.n2897 GND 0.013559f
C4808 VDD.n2898 GND 0.013559f
C4809 VDD.n2899 GND 0.013069f
C4810 VDD.n2900 GND 0.013069f
C4811 VDD.n2901 GND 0.005279f
C4812 VDD.n2902 GND 0.005279f
C4813 VDD.n2903 GND 0.005279f
C4814 VDD.n2904 GND 0.005279f
C4815 VDD.n2905 GND 0.005279f
C4816 VDD.n2906 GND 0.005279f
C4817 VDD.n2907 GND 0.005279f
C4818 VDD.n2908 GND 0.005279f
C4819 VDD.n2909 GND 0.005279f
C4820 VDD.n2910 GND 0.005279f
C4821 VDD.n2911 GND 0.005279f
C4822 VDD.n2912 GND 0.005279f
C4823 VDD.n2913 GND 0.005279f
C4824 VDD.n2914 GND 0.005279f
C4825 VDD.n2915 GND 0.005279f
C4826 VDD.n2916 GND 0.005279f
C4827 VDD.n2917 GND 0.005279f
C4828 VDD.n2918 GND 0.005279f
C4829 VDD.n2919 GND 0.005279f
C4830 VDD.n2920 GND 0.005279f
C4831 VDD.n2921 GND 0.005279f
C4832 VDD.n2922 GND 0.005279f
C4833 VDD.n2923 GND 0.005279f
C4834 VDD.n2924 GND 0.005279f
C4835 VDD.n2925 GND 0.005279f
C4836 VDD.n2926 GND 0.005279f
C4837 VDD.n2927 GND 0.005279f
C4838 VDD.n2928 GND 0.005279f
C4839 VDD.n2929 GND 0.005279f
C4840 VDD.n2930 GND 0.005279f
C4841 VDD.n2931 GND 0.005279f
C4842 VDD.n2932 GND 0.005279f
C4843 VDD.n2933 GND 0.005279f
C4844 VDD.n2934 GND 0.005279f
C4845 VDD.n2935 GND 0.005279f
C4846 VDD.n2936 GND 0.005279f
C4847 VDD.n2937 GND 0.005279f
C4848 VDD.n2938 GND 0.005279f
C4849 VDD.n2939 GND 0.005279f
C4850 VDD.n2940 GND 0.005279f
C4851 VDD.n2941 GND 0.005279f
C4852 VDD.n2942 GND 0.005279f
C4853 VDD.n2943 GND 0.005279f
C4854 VDD.n2944 GND 0.005279f
C4855 VDD.n2945 GND 0.005279f
C4856 VDD.n2946 GND 0.005279f
C4857 VDD.n2947 GND 0.005279f
C4858 VDD.n2948 GND 0.005279f
C4859 VDD.n2949 GND 0.005279f
C4860 VDD.n2950 GND 0.005279f
C4861 VDD.n2951 GND 0.005279f
C4862 VDD.n2952 GND 0.005279f
C4863 VDD.n2953 GND 0.005279f
C4864 VDD.n2954 GND 0.005279f
C4865 VDD.n2955 GND 0.005279f
C4866 VDD.n2956 GND 0.005279f
C4867 VDD.n2957 GND 0.005279f
C4868 VDD.n2958 GND 0.005279f
C4869 VDD.n2959 GND 0.005279f
C4870 VDD.n2960 GND 0.005279f
C4871 VDD.n2961 GND 0.005279f
C4872 VDD.n2962 GND 0.005279f
C4873 VDD.n2963 GND 0.005279f
C4874 VDD.n2964 GND 0.005279f
C4875 VDD.n2965 GND 0.005279f
C4876 VDD.n2966 GND 0.005279f
C4877 VDD.n2967 GND 0.005279f
C4878 VDD.n2968 GND 0.005279f
C4879 VDD.n2969 GND 0.005279f
C4880 VDD.n2970 GND 0.005279f
C4881 VDD.n2971 GND 0.005279f
C4882 VDD.n2972 GND 0.005279f
C4883 VDD.n2973 GND 0.005279f
C4884 VDD.n2974 GND 0.005279f
C4885 VDD.n2975 GND 0.005279f
C4886 VDD.n2976 GND 0.005279f
C4887 VDD.n2977 GND 0.005279f
C4888 VDD.n2978 GND 0.005279f
C4889 VDD.n2979 GND 0.005279f
C4890 VDD.n2980 GND 0.005279f
C4891 VDD.n2981 GND 0.005279f
C4892 VDD.n2982 GND 0.005279f
C4893 VDD.n2983 GND 0.005279f
C4894 VDD.n2984 GND 0.005279f
C4895 VDD.n2985 GND 0.005279f
C4896 VDD.n2986 GND 0.005279f
C4897 VDD.n2987 GND 0.005279f
C4898 VDD.n2988 GND 0.005279f
C4899 VDD.n2989 GND 0.005279f
C4900 VDD.n2990 GND 0.005279f
C4901 VDD.n2991 GND 0.005279f
C4902 VDD.n2992 GND 0.005279f
C4903 VDD.n2993 GND 0.005279f
C4904 VDD.n2994 GND 0.005279f
C4905 VDD.n2995 GND 0.005279f
C4906 VDD.n2996 GND 0.005279f
C4907 VDD.n2997 GND 0.005279f
C4908 VDD.n2998 GND 0.005279f
C4909 VDD.n2999 GND 0.005279f
C4910 VDD.n3000 GND 0.005279f
C4911 VDD.n3001 GND 0.005279f
C4912 VDD.n3002 GND 0.005279f
C4913 VDD.n3003 GND 0.005279f
C4914 VDD.n3004 GND 0.005279f
C4915 VDD.n3005 GND 0.005279f
C4916 VDD.n3006 GND 0.005279f
C4917 VDD.n3007 GND 0.005279f
C4918 VDD.n3008 GND 0.005279f
C4919 VDD.n3009 GND 0.005279f
C4920 VDD.n3010 GND 0.005279f
C4921 VDD.n3011 GND 0.005279f
C4922 VDD.n3012 GND 0.005279f
C4923 VDD.n3013 GND 0.005279f
C4924 VDD.n3014 GND 0.005279f
C4925 VDD.n3015 GND 0.005279f
C4926 VDD.n3016 GND 0.005279f
C4927 VDD.n3017 GND 0.005279f
C4928 VDD.n3018 GND 0.005279f
C4929 VDD.n3019 GND 0.005279f
C4930 VDD.n3020 GND 0.005279f
C4931 VDD.n3021 GND 0.005279f
C4932 VDD.n3022 GND 0.005279f
C4933 VDD.n3023 GND 0.005279f
C4934 VDD.n3024 GND 0.005279f
C4935 VDD.n3025 GND 0.005279f
C4936 VDD.n3026 GND 0.306189f
C4937 VDD.n3027 GND 0.005279f
C4938 VDD.n3028 GND 0.005279f
C4939 VDD.n3029 GND 0.005279f
C4940 VDD.n3030 GND 0.005279f
C4941 VDD.n3031 GND 0.005279f
C4942 VDD.n3032 GND 0.005279f
C4943 VDD.n3033 GND 0.005279f
C4944 VDD.n3034 GND 0.005279f
C4945 VDD.n3035 GND 0.005279f
C4946 VDD.n3036 GND 0.013069f
C4947 VDD.n3037 GND 0.013069f
C4948 VDD.n3038 GND 0.013559f
C4949 VDD.n3039 GND 0.005279f
C4950 VDD.n3040 GND 0.005279f
C4951 VDD.n3041 GND 0.003144f
C4952 VDD.n3042 GND 0.005279f
C4953 VDD.n3043 GND 0.005279f
C4954 VDD.n3044 GND 0.004774f
C4955 VDD.n3045 GND 0.005279f
C4956 VDD.n3046 GND 0.005279f
C4957 VDD.n3047 GND 0.005279f
C4958 VDD.n3048 GND 0.005279f
C4959 VDD.n3049 GND 0.005279f
C4960 VDD.n3050 GND 0.005279f
C4961 VDD.n3051 GND 0.005279f
C4962 VDD.n3052 GND 0.005279f
C4963 VDD.n3053 GND 0.005279f
C4964 VDD.n3054 GND 0.005279f
C4965 VDD.n3055 GND 0.005279f
C4966 VDD.n3056 GND 0.005279f
C4967 VDD.n3057 GND 0.005279f
C4968 VDD.n3058 GND 0.005279f
C4969 VDD.n3059 GND 0.005279f
C4970 VDD.n3060 GND 0.005279f
C4971 VDD.n3061 GND 0.005279f
C4972 VDD.n3062 GND 0.005279f
C4973 VDD.n3063 GND 0.005279f
C4974 VDD.n3064 GND 0.005279f
C4975 VDD.n3065 GND 0.005279f
C4976 VDD.n3066 GND 0.005279f
C4977 VDD.n3067 GND 0.005279f
C4978 VDD.n3068 GND 0.005279f
C4979 VDD.n3069 GND 0.005279f
C4980 VDD.n3070 GND 0.005279f
C4981 VDD.n3071 GND 0.005279f
C4982 VDD.n3072 GND 0.005279f
C4983 VDD.n3073 GND 0.005279f
C4984 VDD.n3074 GND 0.005279f
C4985 VDD.n3075 GND 0.005279f
C4986 VDD.n3076 GND 0.005279f
C4987 VDD.n3077 GND 0.005279f
C4988 VDD.n3078 GND 0.005279f
C4989 VDD.n3079 GND 0.005279f
C4990 VDD.n3080 GND 2.55951f
C4991 VDD.n3082 GND 0.013559f
C4992 VDD.n3083 GND 0.013559f
C4993 VDD.n3084 GND 0.013069f
C4994 VDD.n3085 GND 0.005279f
C4995 VDD.n3086 GND 0.005279f
C4996 VDD.n3087 GND 0.404289f
C4997 VDD.n3088 GND 0.005279f
C4998 VDD.n3089 GND 0.005279f
C4999 VDD.n3090 GND 0.005279f
C5000 VDD.n3091 GND 0.005279f
C5001 VDD.n3092 GND 0.005279f
C5002 VDD.n3093 GND 0.404289f
C5003 VDD.n3094 GND 0.005279f
C5004 VDD.n3095 GND 0.005279f
C5005 VDD.n3096 GND 0.005279f
C5006 VDD.n3097 GND 0.005279f
C5007 VDD.n3098 GND 0.005279f
C5008 VDD.n3099 GND 0.252681f
C5009 VDD.n3100 GND 0.005279f
C5010 VDD.n3101 GND 0.005279f
C5011 VDD.n3102 GND 0.005279f
C5012 VDD.n3103 GND 0.005279f
C5013 VDD.n3104 GND 0.005279f
C5014 VDD.n3105 GND 0.249708f
C5015 VDD.n3106 GND 0.005279f
C5016 VDD.n3107 GND 0.005279f
C5017 VDD.n3108 GND 0.005279f
C5018 VDD.n3109 GND 0.005279f
C5019 VDD.n3110 GND 0.005279f
C5020 VDD.n3111 GND 0.404289f
C5021 VDD.n3112 GND 0.005279f
C5022 VDD.n3113 GND 0.005279f
C5023 VDD.n3114 GND 0.005279f
C5024 VDD.n3115 GND 0.005279f
C5025 VDD.n3116 GND 0.005279f
C5026 VDD.n3117 GND 0.404289f
C5027 VDD.n3118 GND 0.005279f
C5028 VDD.n3119 GND 0.005279f
C5029 VDD.n3120 GND 0.005279f
C5030 VDD.n3121 GND 0.005279f
C5031 VDD.n3122 GND 0.005279f
C5032 VDD.n3123 GND 0.404289f
C5033 VDD.n3124 GND 0.005279f
C5034 VDD.n3125 GND 0.005279f
C5035 VDD.n3126 GND 0.005279f
C5036 VDD.n3127 GND 0.005279f
C5037 VDD.n3128 GND 0.005279f
C5038 VDD.n3129 GND 0.404289f
C5039 VDD.n3130 GND 0.005279f
C5040 VDD.n3131 GND 0.005279f
C5041 VDD.n3132 GND 0.005279f
C5042 VDD.n3133 GND 0.005279f
C5043 VDD.n3134 GND 0.005279f
C5044 VDD.n3135 GND 0.217008f
C5045 VDD.n3136 GND 0.005279f
C5046 VDD.n3137 GND 0.005279f
C5047 VDD.n3138 GND 0.005279f
C5048 VDD.n3139 GND 0.005279f
C5049 VDD.n3140 GND 0.005279f
C5050 VDD.n3141 GND 0.404289f
C5051 VDD.n3142 GND 0.005279f
C5052 VDD.n3143 GND 0.005279f
C5053 VDD.n3144 GND 0.005279f
C5054 VDD.n3145 GND 0.005279f
C5055 VDD.n3146 GND 0.005279f
C5056 VDD.n3147 GND 0.332944f
C5057 VDD.n3148 GND 0.005279f
C5058 VDD.n3149 GND 0.005279f
C5059 VDD.n3150 GND 0.005279f
C5060 VDD.n3151 GND 0.005279f
C5061 VDD.n3152 GND 0.005279f
C5062 VDD.n3153 GND 0.404289f
C5063 VDD.n3154 GND 0.005279f
C5064 VDD.n3155 GND 0.005279f
C5065 VDD.n3156 GND 0.005279f
C5066 VDD.n3157 GND 0.005279f
C5067 VDD.n3158 GND 0.005279f
C5068 VDD.n3159 GND 0.404289f
C5069 VDD.n3160 GND 0.005279f
C5070 VDD.n3161 GND 0.005279f
C5071 VDD.n3162 GND 0.005279f
C5072 VDD.n3163 GND 0.005279f
C5073 VDD.n3164 GND 0.005279f
C5074 VDD.n3165 GND 0.404289f
C5075 VDD.n3166 GND 0.005279f
C5076 VDD.n3167 GND 0.005279f
C5077 VDD.n3168 GND 0.005279f
C5078 VDD.n3169 GND 0.005279f
C5079 VDD.n3170 GND 0.005279f
C5080 VDD.n3171 GND 0.282408f
C5081 VDD.n3172 GND 0.005279f
C5082 VDD.n3173 GND 0.005279f
C5083 VDD.n3174 GND 0.005279f
C5084 VDD.n3175 GND 0.005279f
C5085 VDD.n3176 GND 0.005279f
C5086 VDD.n3177 GND 0.404289f
C5087 VDD.n3178 GND 0.005279f
C5088 VDD.n3179 GND 0.005279f
C5089 VDD.n3180 GND 0.005279f
C5090 VDD.n3181 GND 0.005279f
C5091 VDD.n3182 GND 0.005279f
C5092 VDD.n3183 GND 0.267544f
C5093 VDD.n3184 GND 0.005279f
C5094 VDD.n3185 GND 0.005279f
C5095 VDD.n3186 GND 0.005279f
C5096 VDD.n3187 GND 0.005279f
C5097 VDD.n3188 GND 0.005279f
C5098 VDD.n3189 GND 0.404289f
C5099 VDD.n3190 GND 0.005279f
C5100 VDD.n3191 GND 0.005279f
C5101 VDD.n3192 GND 0.005279f
C5102 VDD.n3193 GND 0.005279f
C5103 VDD.n3194 GND 0.005279f
C5104 VDD.n3195 GND 0.404289f
C5105 VDD.n3196 GND 0.005279f
C5106 VDD.n3197 GND 0.005279f
C5107 VDD.n3198 GND 0.005279f
C5108 VDD.n3199 GND 0.005279f
C5109 VDD.n3200 GND 0.005279f
C5110 VDD.n3201 GND 0.404289f
C5111 VDD.n3202 GND 0.005279f
C5112 VDD.n3203 GND 0.005279f
C5113 VDD.n3204 GND 0.005279f
C5114 VDD.n3205 GND 0.005279f
C5115 VDD.n3206 GND 0.005279f
C5116 VDD.n3207 GND 0.347807f
C5117 VDD.n3208 GND 0.005279f
C5118 VDD.n3209 GND 0.005279f
C5119 VDD.n3210 GND 0.005279f
C5120 VDD.n3211 GND 0.005279f
C5121 VDD.n3212 GND 0.005279f
C5122 VDD.n3213 GND 0.404289f
C5123 VDD.n3214 GND 0.005279f
C5124 VDD.n3215 GND 0.005279f
C5125 VDD.n3216 GND 0.005279f
C5126 VDD.n3217 GND 0.005279f
C5127 VDD.n3218 GND 0.005279f
C5128 VDD.t108 GND 0.404289f
C5129 VDD.n3219 GND 0.005279f
C5130 VDD.n3220 GND 0.005279f
C5131 VDD.n3221 GND 0.005279f
C5132 VDD.n3222 GND 0.005279f
C5133 VDD.n3223 GND 0.005279f
C5134 VDD.n3224 GND 0.404289f
C5135 VDD.n3225 GND 0.005279f
C5136 VDD.n3226 GND 0.005279f
C5137 VDD.n3227 GND 0.005279f
C5138 VDD.n3228 GND 0.005279f
C5139 VDD.n3229 GND 0.005279f
C5140 VDD.n3230 GND 0.404289f
C5141 VDD.n3231 GND 0.005279f
C5142 VDD.n3232 GND 0.005279f
C5143 VDD.n3233 GND 0.005279f
C5144 VDD.n3234 GND 0.005279f
C5145 VDD.n3235 GND 0.005279f
C5146 VDD.n3236 GND 0.404289f
C5147 VDD.n3237 GND 0.005279f
C5148 VDD.n3238 GND 0.005279f
C5149 VDD.n3239 GND 0.005279f
C5150 VDD.n3240 GND 0.005279f
C5151 VDD.n3241 GND 0.005279f
C5152 VDD.n3242 GND 0.404289f
C5153 VDD.n3243 GND 0.005279f
C5154 VDD.n3244 GND 0.005279f
C5155 VDD.n3245 GND 0.005279f
C5156 VDD.n3246 GND 0.005279f
C5157 VDD.n3247 GND 0.005279f
C5158 VDD.n3248 GND 0.404289f
C5159 VDD.n3249 GND 0.005279f
C5160 VDD.n3250 GND 0.005279f
C5161 VDD.n3251 GND 0.005279f
C5162 VDD.n3252 GND 0.005279f
C5163 VDD.n3253 GND 0.005279f
C5164 VDD.n3254 GND 0.252681f
C5165 VDD.n3255 GND 0.005279f
C5166 VDD.n3256 GND 0.005279f
C5167 VDD.n3257 GND 0.005279f
C5168 VDD.n3258 GND 0.005279f
C5169 VDD.n3259 GND 0.005279f
C5170 VDD.n3260 GND 0.404289f
C5171 VDD.n3261 GND 0.005279f
C5172 VDD.n3262 GND 0.005279f
C5173 VDD.n3263 GND 0.005279f
C5174 VDD.n3264 GND 0.005279f
C5175 VDD.n3265 GND 0.005279f
C5176 VDD.n3266 GND 0.404289f
C5177 VDD.n3267 GND 0.005279f
C5178 VDD.n3268 GND 0.005279f
C5179 VDD.n3269 GND 0.005279f
C5180 VDD.n3270 GND 0.005279f
C5181 VDD.n3271 GND 0.005279f
C5182 VDD.n3272 GND 0.404289f
C5183 VDD.n3273 GND 0.005279f
C5184 VDD.n3274 GND 0.005279f
C5185 VDD.n3275 GND 0.005279f
C5186 VDD.n3276 GND 0.005279f
C5187 VDD.n3277 GND 0.005279f
C5188 VDD.n3278 GND 0.404289f
C5189 VDD.n3279 GND 0.005279f
C5190 VDD.n3280 GND 0.005279f
C5191 VDD.n3281 GND 0.005279f
C5192 VDD.n3282 GND 0.005279f
C5193 VDD.n3283 GND 0.005279f
C5194 VDD.n3284 GND 0.404289f
C5195 VDD.n3285 GND 0.005279f
C5196 VDD.n3286 GND 0.005279f
C5197 VDD.n3287 GND 0.005279f
C5198 VDD.n3288 GND 0.005279f
C5199 VDD.n3289 GND 0.005279f
C5200 VDD.n3290 GND 0.252681f
C5201 VDD.n3291 GND 0.005279f
C5202 VDD.n3292 GND 0.005279f
C5203 VDD.n3293 GND 0.005279f
C5204 VDD.n3294 GND 0.005279f
C5205 VDD.n3295 GND 0.005279f
C5206 VDD.n3296 GND 0.404289f
C5207 VDD.n3297 GND 0.005279f
C5208 VDD.n3298 GND 0.005279f
C5209 VDD.n3299 GND 0.005279f
C5210 VDD.n3300 GND 0.005279f
C5211 VDD.n3301 GND 0.005279f
C5212 VDD.n3302 GND 0.404289f
C5213 VDD.n3303 GND 0.005279f
C5214 VDD.n3304 GND 0.005279f
C5215 VDD.n3305 GND 0.005279f
C5216 VDD.n3306 GND 0.005279f
C5217 VDD.n3307 GND 0.005279f
C5218 VDD.n3308 GND 0.404289f
C5219 VDD.n3309 GND 0.005279f
C5220 VDD.n3310 GND 0.005279f
C5221 VDD.n3311 GND 0.005279f
C5222 VDD.n3312 GND 0.005279f
C5223 VDD.n3313 GND 0.005279f
C5224 VDD.n3314 GND 0.404289f
C5225 VDD.n3315 GND 0.005279f
C5226 VDD.n3316 GND 0.005279f
C5227 VDD.n3317 GND 0.005279f
C5228 VDD.n3318 GND 0.005279f
C5229 VDD.n3319 GND 0.005279f
C5230 VDD.n3320 GND 0.404289f
C5231 VDD.n3321 GND 0.005279f
C5232 VDD.n3322 GND 0.005279f
C5233 VDD.n3323 GND 0.005279f
C5234 VDD.n3324 GND 0.005279f
C5235 VDD.n3325 GND 0.005279f
C5236 VDD.n3326 GND 0.258626f
C5237 VDD.n3327 GND 0.005279f
C5238 VDD.n3328 GND 0.005279f
C5239 VDD.n3329 GND 0.005279f
C5240 VDD.n3330 GND 0.005279f
C5241 VDD.n3331 GND 0.005279f
C5242 VDD.n3332 GND 0.005279f
C5243 VDD.n3333 GND 0.005279f
C5244 VDD.n3334 GND 0.249708f
C5245 VDD.n3335 GND 0.005279f
C5246 VDD.n3336 GND 0.005279f
C5247 VDD.n3337 GND 0.005279f
C5248 VDD.n3338 GND 0.005279f
C5249 VDD.n3339 GND 0.005279f
C5250 VDD.n3340 GND 0.404289f
C5251 VDD.n3341 GND 0.005279f
C5252 VDD.n3342 GND 0.005279f
C5253 VDD.n3343 GND 0.005279f
C5254 VDD.n3344 GND 0.005279f
C5255 VDD.n3345 GND 0.005279f
C5256 VDD.n3346 GND 0.005279f
C5257 VDD.n3347 GND 0.005279f
C5258 VDD.n3348 GND 0.013627f
C5259 VDD.n3350 GND 0.013069f
C5260 VDD.n3351 GND 0.013559f
C5261 VDD.n3352 GND 0.013001f
C5262 VDD.n3353 GND 0.005279f
C5263 VDD.n3354 GND 0.003144f
C5264 VDD.n3355 GND 0.005279f
C5265 VDD.n3357 GND 0.005279f
C5266 VDD.n3358 GND 0.005279f
C5267 VDD.n3359 GND 0.005279f
C5268 VDD.n3360 GND 0.005279f
C5269 VDD.n3361 GND 0.005279f
C5270 VDD.n3362 GND 0.005279f
C5271 VDD.n3364 GND 0.005279f
C5272 VDD.n3365 GND 0.005279f
C5273 VDD.n3366 GND 0.005279f
C5274 VDD.n3367 GND 0.005279f
C5275 VDD.n3368 GND 0.005279f
C5276 VDD.n3369 GND 0.005279f
C5277 VDD.n3371 GND 0.005279f
C5278 VDD.n3372 GND 0.005279f
C5279 VDD.n3373 GND 0.003959f
C5280 VDD.n3374 GND 0.005279f
C5281 VDD.n3375 GND 0.005279f
C5282 VDD.n3376 GND 0.005279f
C5283 VDD.n3378 GND 0.005279f
C5284 VDD.n3379 GND 0.005279f
C5285 VDD.n3380 GND 0.005279f
C5286 VDD.n3381 GND 0.005279f
C5287 VDD.n3382 GND 0.005279f
C5288 VDD.n3383 GND 0.005279f
C5289 VDD.n3385 GND 0.005279f
C5290 VDD.n3386 GND 0.005279f
C5291 VDD.n3387 GND 0.005279f
C5292 VDD.n3388 GND 0.005279f
C5293 VDD.n3389 GND 0.005279f
C5294 VDD.n3390 GND 0.005279f
C5295 VDD.n3392 GND 0.013559f
C5296 VDD.n3393 GND 0.013069f
C5297 VDD.n3394 GND 0.013069f
C5298 VDD.n3395 GND 0.005279f
C5299 VDD.n3396 GND 0.005279f
C5300 VDD.n3397 GND 0.005279f
C5301 VDD.n3398 GND 0.005279f
C5302 VDD.n3399 GND 0.404289f
C5303 VDD.n3400 GND 0.005279f
C5304 VDD.n3401 GND 0.005279f
C5305 VDD.n3402 GND 0.005279f
C5306 VDD.n3403 GND 0.005279f
C5307 VDD.n3404 GND 0.005279f
C5308 VDD.n3405 GND 0.005279f
C5309 VDD.n3406 GND 0.005279f
C5310 VDD.n3408 GND 0.005279f
C5311 VDD.n3409 GND 0.005279f
C5312 VDD.n3412 GND 0.005279f
C5313 VDD.n3413 GND 0.005279f
C5314 VDD.n3414 GND 0.005279f
C5315 VDD.n3415 GND 0.005279f
C5316 VDD.n3416 GND 0.005279f
C5317 VDD.n3417 GND 0.005279f
C5318 VDD.n3419 GND 0.005279f
C5319 VDD.n3420 GND 0.005279f
C5320 VDD.n3421 GND 0.005279f
C5321 VDD.n3422 GND 0.005279f
C5322 VDD.n3423 GND 0.005279f
C5323 VDD.n3424 GND 0.005279f
C5324 VDD.n3426 GND 0.005279f
C5325 VDD.n3427 GND 0.005279f
C5326 VDD.n3429 GND 0.013559f
C5327 VDD.n3430 GND 0.013559f
C5328 VDD.n3431 GND 0.013069f
C5329 VDD.n3432 GND 0.005279f
C5330 VDD.n3433 GND 0.005279f
C5331 VDD.n3434 GND 0.404289f
C5332 VDD.n3435 GND 0.005279f
C5333 VDD.n3436 GND 0.005279f
C5334 VDD.n3437 GND 0.013627f
C5335 VDD.n3438 GND 0.013001f
C5336 VDD.n3439 GND 0.013559f
C5337 VDD.n3441 GND 0.005279f
C5338 VDD.n3442 GND 0.005279f
C5339 VDD.n3443 GND 0.003144f
C5340 VDD.n3444 GND 0.007544f
C5341 VDD.n3445 GND 0.004774f
C5342 VDD.n3446 GND 0.005279f
C5343 VDD.n3447 GND 0.005279f
C5344 VDD.n3449 GND 0.005279f
C5345 VDD.n3450 GND 0.005279f
C5346 VDD.n3451 GND 0.005279f
C5347 VDD.n3452 GND 0.005279f
C5348 VDD.n3453 GND 0.005279f
C5349 VDD.n3454 GND 0.005279f
C5350 VDD.n3456 GND 0.005279f
C5351 VDD.n3457 GND 0.005279f
C5352 VDD.n3459 GND 0.005279f
C5353 VDD.n3460 GND 0.003959f
C5354 VDD.n3461 GND 0.015022f
C5355 VDD.n3462 GND 0.006248f
C5356 VDD.n3464 GND 0.007763f
C5357 VDD.n3465 GND 0.007763f
C5358 VDD.n3466 GND 0.007763f
C5359 VDD.n3467 GND 0.006248f
C5360 VDD.n3468 GND 0.007763f
C5361 VDD.n3469 GND 0.007763f
C5362 VDD.n3470 GND 0.007763f
C5363 VDD.n3471 GND 0.007763f
C5364 VDD.t45 GND 0.035989f
C5365 VDD.t46 GND 0.048603f
C5366 VDD.t44 GND 0.295093f
C5367 VDD.n3472 GND 0.062024f
C5368 VDD.n3473 GND 0.044734f
C5369 VDD.n3474 GND 0.007763f
C5370 VDD.n3475 GND 0.006248f
C5371 VDD.n3476 GND 0.007763f
C5372 VDD.n3477 GND 0.007763f
C5373 VDD.n3478 GND 0.007763f
C5374 VDD.n3479 GND 0.007763f
C5375 VDD.n3480 GND 0.007763f
C5376 VDD.n3481 GND 0.006248f
C5377 VDD.n3482 GND 0.007763f
C5378 VDD.n3483 GND 0.007763f
C5379 VDD.n3484 GND 0.007763f
C5380 VDD.n3485 GND 0.007763f
C5381 VDD.n3486 GND 0.007763f
C5382 VDD.n3487 GND 0.003155f
C5383 VDD.n3488 GND 0.007763f
C5384 VDD.t14 GND 0.035989f
C5385 VDD.t15 GND 0.048603f
C5386 VDD.t12 GND 0.295093f
C5387 VDD.n3489 GND 0.062024f
C5388 VDD.n3490 GND 0.044734f
C5389 VDD.n3491 GND 0.009623f
C5390 VDD.n3492 GND 0.007763f
C5391 VDD.n3493 GND 0.007763f
C5392 VDD.n3494 GND 0.007763f
C5393 VDD.n3495 GND 0.007763f
C5394 VDD.n3496 GND 0.006248f
C5395 VDD.n3497 GND 0.007763f
C5396 VDD.n3498 GND 0.007763f
C5397 VDD.n3499 GND 0.007763f
C5398 VDD.n3500 GND 0.007763f
C5399 VDD.n3501 GND 0.007763f
C5400 VDD.n3502 GND 0.006248f
C5401 VDD.n3503 GND 0.007763f
C5402 VDD.n3504 GND 0.007763f
C5403 VDD.n3505 GND 0.007763f
C5404 VDD.n3506 GND 0.007763f
C5405 VDD.t64 GND 0.035989f
C5406 VDD.t65 GND 0.048603f
C5407 VDD.t63 GND 0.295093f
C5408 VDD.n3507 GND 0.062024f
C5409 VDD.n3508 GND 0.044734f
C5410 VDD.n3509 GND 0.007763f
C5411 VDD.n3510 GND 0.006248f
C5412 VDD.n3511 GND 0.007763f
C5413 VDD.n3512 GND 0.007763f
C5414 VDD.n3513 GND 0.007763f
C5415 VDD.n3514 GND 0.007763f
C5416 VDD.n3515 GND 0.007763f
C5417 VDD.n3516 GND 0.006248f
C5418 VDD.n3517 GND 0.007763f
C5419 VDD.n3518 GND 0.007763f
C5420 VDD.n3519 GND 0.007763f
C5421 VDD.n3520 GND 0.007763f
C5422 VDD.n3521 GND 0.007763f
C5423 VDD.n3522 GND 0.002843f
C5424 VDD.t21 GND 0.035989f
C5425 VDD.t22 GND 0.048603f
C5426 VDD.t20 GND 0.295093f
C5427 VDD.n3523 GND 0.062024f
C5428 VDD.n3524 GND 0.044734f
C5429 VDD.n3525 GND 0.009623f
C5430 VDD.n3526 GND 0.006909f
C5431 VDD.n3527 GND 0.003405f
C5432 VDD.n3529 GND 0.007763f
C5433 VDD.n3531 GND 0.007763f
C5434 VDD.n3532 GND 0.006248f
C5435 VDD.n3533 GND 0.006248f
C5436 VDD.n3534 GND 0.006248f
C5437 VDD.n3535 GND 0.007763f
C5438 VDD.n3537 GND 0.007763f
C5439 VDD.n3539 GND 0.007763f
C5440 VDD.n3540 GND 0.006248f
C5441 VDD.n3541 GND 0.006248f
C5442 VDD.n3542 GND 0.006248f
C5443 VDD.n3543 GND 0.007763f
C5444 VDD.n3545 GND 0.007763f
C5445 VDD.n3547 GND 0.007763f
C5446 VDD.n3548 GND 0.00403f
C5447 VDD.n3549 GND 0.009623f
C5448 VDD.n3550 GND 0.00328f
C5449 VDD.n3551 GND 0.006248f
C5450 VDD.n3552 GND 0.007763f
C5451 VDD.n3554 GND 0.007763f
C5452 VDD.n3556 GND 0.007763f
C5453 VDD.n3557 GND 0.006248f
C5454 VDD.n3558 GND 0.006248f
C5455 VDD.n3559 GND 0.006248f
C5456 VDD.n3560 GND 0.007763f
C5457 VDD.n3562 GND 0.007763f
C5458 VDD.n3564 GND 0.007763f
C5459 VDD.n3565 GND 0.006248f
C5460 VDD.n3566 GND 0.006248f
C5461 VDD.n3567 GND 0.004155f
C5462 VDD.n3568 GND 0.007763f
C5463 VDD.n3570 GND 0.007763f
C5464 VDD.n3572 GND 0.007763f
C5465 VDD.n3573 GND 0.006248f
C5466 VDD.n3574 GND 0.006248f
C5467 VDD.n3575 GND 0.006248f
C5468 VDD.n3576 GND 0.007763f
C5469 VDD.n3578 GND 0.007763f
C5470 VDD.n3580 GND 0.007763f
C5471 VDD.n3581 GND 0.006248f
C5472 VDD.n3582 GND 0.006248f
C5473 VDD.n3583 GND 0.006248f
C5474 VDD.n3584 GND 0.007763f
C5475 VDD.n3586 GND 0.007763f
C5476 VDD.n3588 GND 0.007763f
C5477 VDD.n3589 GND 0.00428f
C5478 VDD.n3590 GND 0.012747f
C5479 VDD.n3591 GND 0.006155f
C5480 VDD.n3592 GND 0.007763f
C5481 VDD.n3594 GND 0.007763f
C5482 VDD.n3595 GND 0.007763f
C5483 VDD.n3596 GND 0.006248f
C5484 VDD.n3597 GND 0.006248f
C5485 VDD.n3598 GND 0.007763f
C5486 VDD.n3599 GND 0.007763f
C5487 VDD.n3601 GND 0.007763f
C5488 VDD.n3602 GND 0.006248f
C5489 VDD.n3603 GND 0.005186f
C5490 VDD.n3604 GND 0.268688f
C5491 VDD.n3605 GND 0.010528f
C5492 VDD.n3606 GND 0.005186f
C5493 VDD.n3607 GND 0.018791f
C5494 VDD.n3608 GND 0.862087f
C5495 VDD.n3609 GND 0.018791f
C5496 VDD.n3610 GND 0.005186f
C5497 VDD.n3611 GND 0.010389f
C5498 VDD.n3612 GND 0.007763f
C5499 VDD.n3613 GND 0.007763f
C5500 VDD.n3614 GND 0.006248f
C5501 VDD.n3615 GND 0.007763f
C5502 VDD.n3616 GND 0.594542f
C5503 VDD.n3617 GND 0.007763f
C5504 VDD.n3618 GND 0.006248f
C5505 VDD.n3619 GND 0.007763f
C5506 VDD.n3620 GND 0.007763f
C5507 VDD.n3621 GND 0.007763f
C5508 VDD.n3622 GND 0.006248f
C5509 VDD.n3623 GND 0.007763f
C5510 VDD.t13 GND 0.594542f
C5511 VDD.n3624 GND 0.007763f
C5512 VDD.n3625 GND 0.006248f
C5513 VDD.n3626 GND 0.007763f
C5514 VDD.n3627 GND 0.007763f
C5515 VDD.n3628 GND 0.007763f
C5516 VDD.n3629 GND 0.006248f
C5517 VDD.n3630 GND 0.007763f
C5518 VDD.n3631 GND 0.594542f
C5519 VDD.n3632 GND 0.007763f
C5520 VDD.n3633 GND 0.006248f
C5521 VDD.n3634 GND 0.007763f
C5522 VDD.n3635 GND 0.007763f
C5523 VDD.n3636 GND 0.007763f
C5524 VDD.n3637 GND 0.006248f
C5525 VDD.n3638 GND 0.007763f
C5526 VDD.n3639 GND 0.594542f
C5527 VDD.n3640 GND 0.007763f
C5528 VDD.n3641 GND 0.006248f
C5529 VDD.n3642 GND 0.007763f
C5530 VDD.n3643 GND 0.007763f
C5531 VDD.n3644 GND 0.007763f
C5532 VDD.n3645 GND 0.006248f
C5533 VDD.n3646 GND 0.007763f
C5534 VDD.n3647 GND 0.594542f
C5535 VDD.n3648 GND 0.007763f
C5536 VDD.n3649 GND 0.006248f
C5537 VDD.n3650 GND 0.007763f
C5538 VDD.n3651 GND 0.007763f
C5539 VDD.n3652 GND 0.007763f
C5540 VDD.n3653 GND 0.006248f
C5541 VDD.n3654 GND 0.007763f
C5542 VDD.n3655 GND 0.594542f
C5543 VDD.n3656 GND 0.007763f
C5544 VDD.n3657 GND 0.006248f
C5545 VDD.n3658 GND 0.007763f
C5546 VDD.n3659 GND 0.007763f
C5547 VDD.n3660 GND 0.007763f
C5548 VDD.n3661 GND 0.006248f
C5549 VDD.n3662 GND 0.007763f
C5550 VDD.t144 GND 0.297271f
C5551 VDD.n3663 GND 0.338889f
C5552 VDD.n3664 GND 0.007763f
C5553 VDD.n3665 GND 0.006248f
C5554 VDD.n3666 GND 0.007763f
C5555 VDD.n3667 GND 0.007763f
C5556 VDD.n3668 GND 0.007763f
C5557 VDD.n3669 GND 0.006248f
C5558 VDD.n3670 GND 0.007763f
C5559 VDD.n3671 GND 0.594542f
C5560 VDD.n3672 GND 0.007763f
C5561 VDD.n3673 GND 0.006248f
C5562 VDD.n3674 GND 0.007763f
C5563 VDD.n3675 GND 0.007763f
C5564 VDD.n3676 GND 0.007763f
C5565 VDD.n3677 GND 0.006248f
C5566 VDD.n3678 GND 0.007763f
C5567 VDD.n3679 GND 0.594542f
C5568 VDD.n3680 GND 0.007763f
C5569 VDD.n3681 GND 0.006248f
C5570 VDD.n3682 GND 0.007763f
C5571 VDD.n3683 GND 0.007763f
C5572 VDD.n3684 GND 0.007763f
C5573 VDD.n3685 GND 0.006248f
C5574 VDD.n3686 GND 0.007763f
C5575 VDD.n3687 GND 0.594542f
C5576 VDD.n3688 GND 0.007763f
C5577 VDD.n3689 GND 0.006248f
C5578 VDD.n3690 GND 0.007763f
C5579 VDD.n3691 GND 0.007763f
C5580 VDD.n3692 GND 0.007763f
C5581 VDD.n3693 GND 0.006248f
C5582 VDD.n3694 GND 0.007763f
C5583 VDD.t127 GND 0.297271f
C5584 VDD.n3695 GND 0.326998f
C5585 VDD.n3696 GND 0.007763f
C5586 VDD.n3697 GND 0.006248f
C5587 VDD.n3698 GND 0.007763f
C5588 VDD.n3699 GND 0.007763f
C5589 VDD.n3700 GND 0.007763f
C5590 VDD.n3701 GND 0.006248f
C5591 VDD.n3702 GND 0.007763f
C5592 VDD.n3703 GND 0.594542f
C5593 VDD.n3704 GND 0.007763f
C5594 VDD.n3705 GND 0.006248f
C5595 VDD.n3706 GND 0.007763f
C5596 VDD.n3707 GND 0.007763f
C5597 VDD.n3708 GND 0.007763f
C5598 VDD.n3709 GND 0.006248f
C5599 VDD.n3710 GND 0.007763f
C5600 VDD.n3711 GND 0.594542f
C5601 VDD.n3712 GND 0.007763f
C5602 VDD.n3713 GND 0.006248f
C5603 VDD.n3714 GND 0.007763f
C5604 VDD.n3715 GND 0.007763f
C5605 VDD.n3716 GND 0.007763f
C5606 VDD.n3717 GND 0.006248f
C5607 VDD.n3718 GND 0.007763f
C5608 VDD.n3719 GND 0.594542f
C5609 VDD.n3720 GND 0.007763f
C5610 VDD.n3721 GND 0.006248f
C5611 VDD.n3722 GND 0.007763f
C5612 VDD.n3723 GND 0.007763f
C5613 VDD.n3724 GND 0.007763f
C5614 VDD.n3725 GND 0.006248f
C5615 VDD.n3726 GND 0.007763f
C5616 VDD.t120 GND 0.297271f
C5617 VDD.n3727 GND 0.315107f
C5618 VDD.n3728 GND 0.007763f
C5619 VDD.n3729 GND 0.006248f
C5620 VDD.n3730 GND 0.007763f
C5621 VDD.n3731 GND 0.007763f
C5622 VDD.n3732 GND 0.007763f
C5623 VDD.n3733 GND 0.006248f
C5624 VDD.n3734 GND 0.007763f
C5625 VDD.n3735 GND 0.594542f
C5626 VDD.n3736 GND 0.007763f
C5627 VDD.n3737 GND 0.006248f
C5628 VDD.n3738 GND 0.007763f
C5629 VDD.n3739 GND 0.007763f
C5630 VDD.n3740 GND 0.007763f
C5631 VDD.n3741 GND 0.006248f
C5632 VDD.n3742 GND 0.007763f
C5633 VDD.n3743 GND 0.594542f
C5634 VDD.n3744 GND 0.007763f
C5635 VDD.n3745 GND 0.006248f
C5636 VDD.n3746 GND 0.007763f
C5637 VDD.n3747 GND 0.007763f
C5638 VDD.n3748 GND 0.007763f
C5639 VDD.n3749 GND 0.006248f
C5640 VDD.n3750 GND 0.007763f
C5641 VDD.n3751 GND 0.594542f
C5642 VDD.n3752 GND 0.007763f
C5643 VDD.n3753 GND 0.006248f
C5644 VDD.n3754 GND 0.007763f
C5645 VDD.n3755 GND 0.007763f
C5646 VDD.n3756 GND 0.007763f
C5647 VDD.n3757 GND 0.006248f
C5648 VDD.n3758 GND 0.007763f
C5649 VDD.t135 GND 0.297271f
C5650 VDD.n3759 GND 0.303217f
C5651 VDD.n3760 GND 0.007763f
C5652 VDD.n3761 GND 0.006248f
C5653 VDD.n3762 GND 0.007763f
C5654 VDD.n3763 GND 0.007763f
C5655 VDD.n3764 GND 0.007763f
C5656 VDD.n3765 GND 0.006248f
C5657 VDD.n3766 GND 0.007763f
C5658 VDD.n3767 GND 0.594542f
C5659 VDD.n3768 GND 0.007763f
C5660 VDD.n3769 GND 0.006248f
C5661 VDD.n3770 GND 0.007763f
C5662 VDD.n3771 GND 0.007763f
C5663 VDD.n3772 GND 0.007763f
C5664 VDD.n3773 GND 0.006248f
C5665 VDD.n3774 GND 0.006248f
C5666 VDD.n3775 GND 0.006248f
C5667 VDD.n3776 GND 0.007763f
C5668 VDD.n3777 GND 0.007763f
C5669 VDD.n3778 GND 0.007763f
C5670 VDD.n3779 GND 0.006248f
C5671 VDD.n3780 GND 0.006248f
C5672 VDD.n3781 GND 0.006248f
C5673 VDD.n3782 GND 0.007763f
C5674 VDD.n3783 GND 0.007763f
C5675 VDD.n3784 GND 0.007763f
C5676 VDD.n3785 GND 0.006248f
C5677 VDD.n3786 GND 0.006248f
C5678 VDD.n3787 GND 0.006248f
C5679 VDD.n3788 GND 0.007763f
C5680 VDD.n3789 GND 0.007763f
C5681 VDD.n3790 GND 0.007763f
C5682 VDD.n3791 GND 0.006248f
C5683 VDD.n3792 GND 0.006248f
C5684 VDD.n3793 GND 0.006248f
C5685 VDD.n3794 GND 0.007763f
C5686 VDD.n3795 GND 0.007763f
C5687 VDD.n3796 GND 0.007763f
C5688 VDD.n3797 GND 0.006248f
C5689 VDD.n3798 GND 0.006248f
C5690 VDD.n3799 GND 0.006248f
C5691 VDD.n3800 GND 0.007763f
C5692 VDD.n3801 GND 0.007763f
C5693 VDD.n3802 GND 0.007763f
C5694 VDD.n3803 GND 0.006248f
C5695 VDD.n3804 GND 0.006248f
C5696 VDD.n3805 GND 0.006248f
C5697 VDD.n3806 GND 0.007763f
C5698 VDD.n3807 GND 0.007763f
C5699 VDD.n3808 GND 0.007763f
C5700 VDD.n3809 GND 0.006248f
C5701 VDD.n3810 GND 0.006248f
C5702 VDD.n3811 GND 0.006248f
C5703 VDD.n3812 GND 0.007763f
C5704 VDD.n3813 GND 0.007763f
C5705 VDD.n3814 GND 0.007763f
C5706 VDD.n3815 GND 0.006248f
C5707 VDD.n3816 GND 0.006248f
C5708 VDD.n3817 GND 0.006248f
C5709 VDD.n3818 GND 0.007763f
C5710 VDD.n3819 GND 0.007763f
C5711 VDD.n3820 GND 0.007763f
C5712 VDD.n3821 GND 0.006248f
C5713 VDD.n3822 GND 0.006248f
C5714 VDD.n3823 GND 0.006248f
C5715 VDD.n3824 GND 0.007763f
C5716 VDD.n3825 GND 0.007763f
C5717 VDD.n3826 GND 0.007763f
C5718 VDD.n3827 GND 0.006248f
C5719 VDD.n3828 GND 0.006248f
C5720 VDD.n3829 GND 0.006248f
C5721 VDD.n3830 GND 0.007763f
C5722 VDD.n3831 GND 0.007763f
C5723 VDD.n3832 GND 0.007763f
C5724 VDD.n3833 GND 0.006248f
C5725 VDD.n3834 GND 0.006248f
C5726 VDD.n3835 GND 0.005186f
C5727 VDD.n3836 GND 0.018791f
C5728 VDD.n3837 GND 0.019093f
C5729 VDD.n3839 GND 0.019093f
C5730 VDD.n3840 GND 0.002843f
C5731 VDD.t33 GND 0.035989f
C5732 VDD.t32 GND 0.048603f
C5733 VDD.t31 GND 0.295093f
C5734 VDD.n3841 GND 0.062024f
C5735 VDD.n3842 GND 0.044734f
C5736 VDD.n3843 GND 0.009623f
C5737 VDD.n3844 GND 0.003405f
C5738 VDD.n3845 GND 0.006248f
C5739 VDD.n3846 GND 0.007763f
C5740 VDD.n3848 GND 0.007763f
C5741 VDD.n3849 GND 0.007763f
C5742 VDD.n3850 GND 0.006248f
C5743 VDD.n3851 GND 0.006248f
C5744 VDD.n3852 GND 0.006248f
C5745 VDD.n3853 GND 0.007763f
C5746 VDD.n3855 GND 0.007763f
C5747 VDD.n3856 GND 0.007763f
C5748 VDD.n3857 GND 0.006248f
C5749 VDD.n3858 GND 0.006248f
C5750 VDD.n3859 GND 0.00403f
C5751 VDD.n3860 GND 0.007763f
C5752 VDD.n3862 GND 0.007763f
C5753 VDD.n3863 GND 0.007763f
C5754 VDD.n3864 GND 0.006248f
C5755 VDD.n3865 GND 0.006248f
C5756 VDD.n3866 GND 0.006248f
C5757 VDD.n3867 GND 0.007763f
C5758 VDD.n3869 GND 0.007763f
C5759 VDD.n3870 GND 0.007763f
C5760 VDD.n3871 GND 0.006248f
C5761 VDD.n3872 GND 0.006248f
C5762 VDD.n3873 GND 0.006248f
C5763 VDD.n3874 GND 0.007763f
C5764 VDD.n3876 GND 0.007763f
C5765 VDD.n3877 GND 0.007763f
C5766 VDD.n3878 GND 0.004155f
C5767 VDD.t68 GND 0.035989f
C5768 VDD.t67 GND 0.048603f
C5769 VDD.t66 GND 0.295093f
C5770 VDD.n3879 GND 0.062024f
C5771 VDD.n3880 GND 0.044734f
C5772 VDD.n3881 GND 0.009623f
C5773 VDD.n3882 GND 0.003155f
C5774 VDD.n3883 GND 0.006248f
C5775 VDD.n3884 GND 0.007763f
C5776 VDD.n3886 GND 0.007763f
C5777 VDD.n3887 GND 0.007763f
C5778 VDD.n3888 GND 0.006248f
C5779 VDD.n3889 GND 0.006248f
C5780 VDD.n3890 GND 0.006248f
C5781 VDD.n3891 GND 0.007763f
C5782 VDD.n3893 GND 0.007763f
C5783 VDD.n3894 GND 0.007763f
C5784 VDD.n3895 GND 0.006248f
C5785 VDD.n3896 GND 0.006248f
C5786 VDD.n3897 GND 0.00428f
C5787 VDD.n3898 GND 0.007763f
C5788 VDD.n3900 GND 0.007763f
C5789 VDD.n3901 GND 0.007763f
C5790 VDD.n3902 GND 0.006155f
C5791 VDD.n3903 GND 0.006248f
C5792 VDD.n3904 GND 0.006248f
C5793 VDD.n3905 GND 0.007763f
C5794 VDD.n3907 GND 0.007763f
C5795 VDD.n3908 GND 0.007763f
C5796 VDD.n3909 GND 0.006248f
C5797 VDD.n3910 GND 0.006248f
C5798 VDD.n3911 GND 0.005186f
C5799 VDD.n3912 GND 0.019093f
C5800 VDD.n3913 GND 0.018791f
C5801 VDD.n3914 GND 0.005186f
C5802 VDD.n3915 GND 0.018791f
C5803 VDD.n3916 GND 0.862087f
C5804 VDD.n3917 GND 0.594542f
C5805 VDD.n3918 GND 0.594542f
C5806 VDD.n3919 GND 0.007763f
C5807 VDD.n3920 GND 0.006248f
C5808 VDD.n3921 GND 0.006248f
C5809 VDD.n3922 GND 0.006248f
C5810 VDD.n3923 GND 0.007763f
C5811 VDD.t24 GND 0.594542f
C5812 VDD.n3924 GND 0.594542f
C5813 VDD.n3925 GND 0.594542f
C5814 VDD.n3926 GND 0.007763f
C5815 VDD.n3927 GND 0.006248f
C5816 VDD.n3928 GND 0.006248f
C5817 VDD.n3929 GND 0.006248f
C5818 VDD.n3930 GND 0.007763f
C5819 VDD.n3931 GND 0.594542f
C5820 VDD.n3932 GND 0.594542f
C5821 VDD.n3933 GND 0.594542f
C5822 VDD.n3934 GND 0.007763f
C5823 VDD.n3935 GND 0.006248f
C5824 VDD.n3936 GND 0.006248f
C5825 VDD.n3937 GND 0.006248f
C5826 VDD.n3938 GND 0.007763f
C5827 VDD.n3939 GND 0.594542f
C5828 VDD.n3940 GND 0.594542f
C5829 VDD.n3941 GND 0.338889f
C5830 VDD.n3942 GND 0.007763f
C5831 VDD.n3943 GND 0.006248f
C5832 VDD.n3944 GND 0.006248f
C5833 VDD.n3945 GND 0.006248f
C5834 VDD.n3946 GND 0.007763f
C5835 VDD.n3947 GND 0.594542f
C5836 VDD.n3948 GND 0.594542f
C5837 VDD.n3949 GND 0.594542f
C5838 VDD.n3950 GND 0.007763f
C5839 VDD.n3951 GND 0.006248f
C5840 VDD.n3952 GND 0.006248f
C5841 VDD.n3953 GND 0.006248f
C5842 VDD.n3954 GND 0.007763f
C5843 VDD.n3955 GND 0.594542f
C5844 VDD.n3956 GND 0.594542f
C5845 VDD.n3957 GND 0.326998f
C5846 VDD.n3958 GND 0.007763f
C5847 VDD.n3959 GND 0.006248f
C5848 VDD.n3960 GND 0.006248f
C5849 VDD.n3961 GND 0.006248f
C5850 VDD.n3962 GND 0.007763f
C5851 VDD.n3963 GND 0.594542f
C5852 VDD.n3964 GND 0.594542f
C5853 VDD.n3965 GND 0.594542f
C5854 VDD.n3966 GND 0.007763f
C5855 VDD.n3967 GND 0.006248f
C5856 VDD.n3968 GND 0.006248f
C5857 VDD.n3969 GND 0.006248f
C5858 VDD.n3970 GND 0.007763f
C5859 VDD.n3971 GND 0.594542f
C5860 VDD.n3972 GND 0.594542f
C5861 VDD.n3973 GND 0.315107f
C5862 VDD.n3974 GND 0.007763f
C5863 VDD.n3975 GND 0.006248f
C5864 VDD.n3976 GND 0.006248f
C5865 VDD.n3977 GND 0.006248f
C5866 VDD.n3978 GND 0.007763f
C5867 VDD.n3979 GND 0.594542f
C5868 VDD.n3980 GND 0.594542f
C5869 VDD.n3981 GND 0.594542f
C5870 VDD.n3982 GND 0.007763f
C5871 VDD.n3983 GND 0.006248f
C5872 VDD.n3984 GND 0.006248f
C5873 VDD.n3985 GND 0.006248f
C5874 VDD.n3986 GND 0.007763f
C5875 VDD.n3987 GND 0.594542f
C5876 VDD.n3988 GND 0.594542f
C5877 VDD.n3989 GND 0.303217f
C5878 VDD.n3990 GND 0.007763f
C5879 VDD.n3991 GND 0.006248f
C5880 VDD.n3992 GND 0.006248f
C5881 VDD.n3993 GND 0.006248f
C5882 VDD.n3994 GND 0.007763f
C5883 VDD.n3995 GND 0.594542f
C5884 VDD.n3996 GND 0.594542f
C5885 VDD.n3997 GND 0.594542f
C5886 VDD.n3998 GND 0.007763f
C5887 VDD.n3999 GND 0.006248f
C5888 VDD.n4000 GND 0.542227f
C5889 VDD.n4001 GND 3.55247f
C5890 a_n16612_8244.t6 GND 0.62975f
C5891 a_n16612_8244.t8 GND 0.62975f
C5892 a_n16612_8244.t9 GND 0.643404f
C5893 a_n16612_8244.t1 GND 0.62975f
C5894 a_n16612_8244.n0 GND 5.23295f
C5895 a_n16612_8244.n1 GND 9.81401f
C5896 a_n16612_8244.n2 GND 3.20334f
C5897 a_n16612_8244.n3 GND 0.263649f
C5898 a_n16612_8244.n4 GND 0.263649f
C5899 a_n16612_8244.n5 GND 0.263649f
C5900 a_n16612_8244.n6 GND 3.24396f
C5901 a_n16612_8244.n7 GND 0.263649f
C5902 a_n16612_8244.n8 GND 1.47399f
C5903 a_n16612_8244.n9 GND 1.72935f
C5904 a_n16612_8244.n10 GND 0.263608f
C5905 a_n16612_8244.n11 GND 1.47399f
C5906 a_n16612_8244.n12 GND 0.263608f
C5907 a_n16612_8244.n13 GND 1.47399f
C5908 a_n16612_8244.n14 GND 0.263608f
C5909 a_n16612_8244.n15 GND 1.47399f
C5910 a_n16612_8244.n16 GND 1.76998f
C5911 a_n16612_8244.n17 GND 0.263608f
C5912 a_n16612_8244.n18 GND 0.263475f
C5913 a_n16612_8244.n19 GND 0.263475f
C5914 a_n16612_8244.n20 GND 0.263475f
C5915 a_n16612_8244.n21 GND 0.263475f
C5916 a_n16612_8244.t3 GND 0.634758f
C5917 a_n16612_8244.t5 GND 0.634758f
C5918 a_n16612_8244.t2 GND 0.672508f
C5919 a_n16612_8244.t10 GND 0.634757f
C5920 a_n16612_8244.n22 GND 24.437199f
C5921 a_n16612_8244.n23 GND 7.94048f
C5922 a_n16612_8244.n24 GND 0.4525f
C5923 a_n16612_8244.n25 GND 0.4525f
C5924 a_n16612_8244.n26 GND 0.4525f
C5925 a_n16612_8244.n27 GND 0.4525f
C5926 a_n16612_8244.n28 GND 0.454471f
C5927 a_n16612_8244.n29 GND 0.454471f
C5928 a_n16612_8244.n30 GND 0.454471f
C5929 a_n16612_8244.n31 GND 0.454471f
C5930 a_n16612_8244.n32 GND 0.449952f
C5931 a_n16612_8244.n33 GND 0.449952f
C5932 a_n16612_8244.n34 GND 0.449952f
C5933 a_n16612_8244.n35 GND 0.449952f
C5934 a_n16612_8244.n36 GND 5.74739f
C5935 a_n16612_8244.n37 GND 4.15476f
C5936 a_n16612_8244.n38 GND 0.263606f
C5937 a_n16612_8244.n39 GND 0.263606f
C5938 a_n16612_8244.n40 GND 0.263606f
C5939 a_n16612_8244.n41 GND 0.263606f
C5940 a_n16612_8244.n42 GND 0.263606f
C5941 a_n16612_8244.n43 GND 0.263606f
C5942 a_n16612_8244.n44 GND 0.263606f
C5943 a_n16612_8244.n45 GND 0.263606f
C5944 a_n16612_8244.n46 GND 0.263651f
C5945 a_n16612_8244.n47 GND 0.263477f
C5946 a_n16612_8244.n48 GND 0.263651f
C5947 a_n16612_8244.n49 GND 0.263477f
C5948 a_n16612_8244.n50 GND 0.263651f
C5949 a_n16612_8244.n51 GND 0.263477f
C5950 a_n16612_8244.n52 GND 0.263651f
C5951 a_n16612_8244.n53 GND 0.263477f
C5952 a_n16612_8244.n54 GND 0.449953f
C5953 a_n16612_8244.n55 GND 0.449953f
C5954 a_n16612_8244.n56 GND 0.449953f
C5955 a_n16612_8244.n57 GND 0.449953f
C5956 a_n16612_8244.n58 GND 7.91413f
C5957 a_n16612_8244.n59 GND 0.191956f
C5958 a_n16612_8244.n60 GND 0.194075f
C5959 a_n16612_8244.n61 GND 0.191956f
C5960 a_n16612_8244.n62 GND 0.194075f
C5961 a_n16612_8244.n63 GND 0.191956f
C5962 a_n16612_8244.n64 GND 0.194075f
C5963 a_n16612_8244.n65 GND 0.191956f
C5964 a_n16612_8244.n66 GND 0.194075f
C5965 a_n16612_8244.t11 GND 0.649804f
C5966 a_n16612_8244.t7 GND 0.67991f
C5967 a_n16612_8244.t4 GND 0.679908f
C5968 a_n16612_8244.t49 GND 1.20081f
C5969 a_n16612_8244.t29 GND 1.1688f
C5970 a_n16612_8244.t59 GND 1.21224f
C5971 a_n16612_8244.t54 GND 0.760483f
C5972 a_n16612_8244.n67 GND 0.618098f
C5973 a_n16612_8244.t33 GND 0.760483f
C5974 a_n16612_8244.n68 GND 0.603881f
C5975 a_n16612_8244.t72 GND 0.760483f
C5976 a_n16612_8244.n69 GND 0.603881f
C5977 a_n16612_8244.t55 GND 0.760483f
C5978 a_n16612_8244.n70 GND 0.603966f
C5979 a_n16612_8244.t24 GND 0.760483f
C5980 a_n16612_8244.n71 GND 0.611778f
C5981 a_n16612_8244.t75 GND 1.20081f
C5982 a_n16612_8244.t53 GND 1.1688f
C5983 a_n16612_8244.t20 GND 1.21224f
C5984 a_n16612_8244.t13 GND 0.760483f
C5985 a_n16612_8244.n72 GND 0.618098f
C5986 a_n16612_8244.t56 GND 0.760483f
C5987 a_n16612_8244.n73 GND 0.603881f
C5988 a_n16612_8244.t34 GND 0.760483f
C5989 a_n16612_8244.n74 GND 0.603881f
C5990 a_n16612_8244.t17 GND 0.760483f
C5991 a_n16612_8244.n75 GND 0.603966f
C5992 a_n16612_8244.t48 GND 0.760483f
C5993 a_n16612_8244.n76 GND 0.611778f
C5994 a_n16612_8244.t69 GND 1.20081f
C5995 a_n16612_8244.t43 GND 1.1688f
C5996 a_n16612_8244.t50 GND 1.21224f
C5997 a_n16612_8244.t35 GND 0.760483f
C5998 a_n16612_8244.n77 GND 0.618098f
C5999 a_n16612_8244.t73 GND 0.760483f
C6000 a_n16612_8244.n78 GND 0.603881f
C6001 a_n16612_8244.t44 GND 0.760483f
C6002 a_n16612_8244.n79 GND 0.603881f
C6003 a_n16612_8244.t21 GND 0.760483f
C6004 a_n16612_8244.n80 GND 0.603966f
C6005 a_n16612_8244.t14 GND 0.760483f
C6006 a_n16612_8244.n81 GND 0.611778f
C6007 a_n16612_8244.t47 GND 1.20081f
C6008 a_n16612_8244.t23 GND 1.1688f
C6009 a_n16612_8244.t31 GND 1.21224f
C6010 a_n16612_8244.t16 GND 0.760483f
C6011 a_n16612_8244.n82 GND 0.618098f
C6012 a_n16612_8244.t51 GND 0.760483f
C6013 a_n16612_8244.n83 GND 0.603881f
C6014 a_n16612_8244.t26 GND 0.760483f
C6015 a_n16612_8244.n84 GND 0.603881f
C6016 a_n16612_8244.t62 GND 0.760483f
C6017 a_n16612_8244.n85 GND 0.603966f
C6018 a_n16612_8244.t58 GND 0.760483f
C6019 a_n16612_8244.n86 GND 0.611778f
C6020 a_n16612_8244.t15 GND 1.20081f
C6021 a_n16612_8244.t42 GND 0.760483f
C6022 a_n16612_8244.n87 GND 0.611776f
C6023 a_n16612_8244.t68 GND 0.760483f
C6024 a_n16612_8244.n88 GND 0.603964f
C6025 a_n16612_8244.t40 GND 0.760483f
C6026 a_n16612_8244.n89 GND 0.603879f
C6027 a_n16612_8244.t64 GND 0.760483f
C6028 a_n16612_8244.n90 GND 0.543328f
C6029 a_n16612_8244.t37 GND 0.760483f
C6030 a_n16612_8244.n91 GND 0.550915f
C6031 a_n16612_8244.t28 GND 1.21224f
C6032 a_n16612_8244.t71 GND 1.17214f
C6033 a_n16612_8244.t36 GND 1.20081f
C6034 a_n16612_8244.t70 GND 0.760483f
C6035 a_n16612_8244.n92 GND 0.611776f
C6036 a_n16612_8244.t27 GND 0.760483f
C6037 a_n16612_8244.n93 GND 0.603964f
C6038 a_n16612_8244.t66 GND 0.760483f
C6039 a_n16612_8244.n94 GND 0.603879f
C6040 a_n16612_8244.t25 GND 0.760483f
C6041 a_n16612_8244.n95 GND 0.543328f
C6042 a_n16612_8244.t63 GND 0.760483f
C6043 a_n16612_8244.n96 GND 0.550915f
C6044 a_n16612_8244.t52 GND 1.21224f
C6045 a_n16612_8244.t32 GND 1.17214f
C6046 a_n16612_8244.t61 GND 1.20081f
C6047 a_n16612_8244.t67 GND 0.760483f
C6048 a_n16612_8244.n97 GND 0.611776f
C6049 a_n16612_8244.t30 GND 0.760483f
C6050 a_n16612_8244.n98 GND 0.603964f
C6051 a_n16612_8244.t38 GND 0.760483f
C6052 a_n16612_8244.n99 GND 0.603879f
C6053 a_n16612_8244.t65 GND 0.760483f
C6054 a_n16612_8244.n100 GND 0.543328f
C6055 a_n16612_8244.t12 GND 0.760483f
C6056 a_n16612_8244.n101 GND 0.550915f
C6057 a_n16612_8244.t41 GND 1.21224f
C6058 a_n16612_8244.t18 GND 1.17214f
C6059 a_n16612_8244.t39 GND 1.20081f
C6060 a_n16612_8244.t46 GND 0.760483f
C6061 a_n16612_8244.n102 GND 0.611776f
C6062 a_n16612_8244.t74 GND 0.760483f
C6063 a_n16612_8244.n103 GND 0.603964f
C6064 a_n16612_8244.t19 GND 0.760483f
C6065 a_n16612_8244.n104 GND 0.603879f
C6066 a_n16612_8244.t45 GND 0.760483f
C6067 a_n16612_8244.n105 GND 0.543328f
C6068 a_n16612_8244.t57 GND 0.760483f
C6069 a_n16612_8244.n106 GND 0.550915f
C6070 a_n16612_8244.t22 GND 1.21224f
C6071 a_n16612_8244.t60 GND 1.17214f
C6072 a_n16612_8244.n107 GND 7.77775f
C6073 a_n16612_8244.t0 GND 0.658361f
.ends

