* NGSPICE file created from diff_pair_sample_1759.ext - technology: sky130A

.subckt diff_pair_sample_1759 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n2634_n1792# sky130_fd_pr__pfet_01v8 ad=1.6068 pd=9.02 as=1.6068 ps=9.02 w=4.12 l=3.83
X1 B.t11 B.t9 B.t10 w_n2634_n1792# sky130_fd_pr__pfet_01v8 ad=1.6068 pd=9.02 as=0 ps=0 w=4.12 l=3.83
X2 VDD2.t1 VN.t0 VTAIL.t1 w_n2634_n1792# sky130_fd_pr__pfet_01v8 ad=1.6068 pd=9.02 as=1.6068 ps=9.02 w=4.12 l=3.83
X3 B.t8 B.t6 B.t7 w_n2634_n1792# sky130_fd_pr__pfet_01v8 ad=1.6068 pd=9.02 as=0 ps=0 w=4.12 l=3.83
X4 VDD1.t0 VP.t1 VTAIL.t2 w_n2634_n1792# sky130_fd_pr__pfet_01v8 ad=1.6068 pd=9.02 as=1.6068 ps=9.02 w=4.12 l=3.83
X5 VDD2.t0 VN.t1 VTAIL.t0 w_n2634_n1792# sky130_fd_pr__pfet_01v8 ad=1.6068 pd=9.02 as=1.6068 ps=9.02 w=4.12 l=3.83
X6 B.t5 B.t3 B.t4 w_n2634_n1792# sky130_fd_pr__pfet_01v8 ad=1.6068 pd=9.02 as=0 ps=0 w=4.12 l=3.83
X7 B.t2 B.t0 B.t1 w_n2634_n1792# sky130_fd_pr__pfet_01v8 ad=1.6068 pd=9.02 as=0 ps=0 w=4.12 l=3.83
R0 VP.n0 VP.t0 102.966
R1 VP.n0 VP.t1 61.0169
R2 VP VP.n0 0.62124
R3 VTAIL.n1 VTAIL.t0 98.0459
R4 VTAIL.n3 VTAIL.t1 98.0457
R5 VTAIL.n0 VTAIL.t2 98.0457
R6 VTAIL.n2 VTAIL.t3 98.0457
R7 VTAIL.n1 VTAIL.n0 23.091
R8 VTAIL.n3 VTAIL.n2 19.5048
R9 VTAIL.n2 VTAIL.n1 2.26343
R10 VTAIL VTAIL.n0 1.42507
R11 VTAIL VTAIL.n3 0.838862
R12 VDD1 VDD1.t0 150.53
R13 VDD1 VDD1.t1 115.68
R14 B.n238 B.n237 585
R15 B.n236 B.n79 585
R16 B.n235 B.n234 585
R17 B.n233 B.n80 585
R18 B.n232 B.n231 585
R19 B.n230 B.n81 585
R20 B.n229 B.n228 585
R21 B.n227 B.n82 585
R22 B.n226 B.n225 585
R23 B.n224 B.n83 585
R24 B.n223 B.n222 585
R25 B.n221 B.n84 585
R26 B.n220 B.n219 585
R27 B.n218 B.n85 585
R28 B.n217 B.n216 585
R29 B.n215 B.n86 585
R30 B.n214 B.n213 585
R31 B.n212 B.n87 585
R32 B.n210 B.n209 585
R33 B.n208 B.n90 585
R34 B.n207 B.n206 585
R35 B.n205 B.n91 585
R36 B.n204 B.n203 585
R37 B.n202 B.n92 585
R38 B.n201 B.n200 585
R39 B.n199 B.n93 585
R40 B.n198 B.n197 585
R41 B.n196 B.n94 585
R42 B.n195 B.n194 585
R43 B.n190 B.n95 585
R44 B.n189 B.n188 585
R45 B.n187 B.n96 585
R46 B.n186 B.n185 585
R47 B.n184 B.n97 585
R48 B.n183 B.n182 585
R49 B.n181 B.n98 585
R50 B.n180 B.n179 585
R51 B.n178 B.n99 585
R52 B.n177 B.n176 585
R53 B.n175 B.n100 585
R54 B.n174 B.n173 585
R55 B.n172 B.n101 585
R56 B.n171 B.n170 585
R57 B.n169 B.n102 585
R58 B.n168 B.n167 585
R59 B.n166 B.n103 585
R60 B.n239 B.n78 585
R61 B.n241 B.n240 585
R62 B.n242 B.n77 585
R63 B.n244 B.n243 585
R64 B.n245 B.n76 585
R65 B.n247 B.n246 585
R66 B.n248 B.n75 585
R67 B.n250 B.n249 585
R68 B.n251 B.n74 585
R69 B.n253 B.n252 585
R70 B.n254 B.n73 585
R71 B.n256 B.n255 585
R72 B.n257 B.n72 585
R73 B.n259 B.n258 585
R74 B.n260 B.n71 585
R75 B.n262 B.n261 585
R76 B.n263 B.n70 585
R77 B.n265 B.n264 585
R78 B.n266 B.n69 585
R79 B.n268 B.n267 585
R80 B.n269 B.n68 585
R81 B.n271 B.n270 585
R82 B.n272 B.n67 585
R83 B.n274 B.n273 585
R84 B.n275 B.n66 585
R85 B.n277 B.n276 585
R86 B.n278 B.n65 585
R87 B.n280 B.n279 585
R88 B.n281 B.n64 585
R89 B.n283 B.n282 585
R90 B.n284 B.n63 585
R91 B.n286 B.n285 585
R92 B.n287 B.n62 585
R93 B.n289 B.n288 585
R94 B.n290 B.n61 585
R95 B.n292 B.n291 585
R96 B.n293 B.n60 585
R97 B.n295 B.n294 585
R98 B.n296 B.n59 585
R99 B.n298 B.n297 585
R100 B.n299 B.n58 585
R101 B.n301 B.n300 585
R102 B.n302 B.n57 585
R103 B.n304 B.n303 585
R104 B.n305 B.n56 585
R105 B.n307 B.n306 585
R106 B.n308 B.n55 585
R107 B.n310 B.n309 585
R108 B.n311 B.n54 585
R109 B.n313 B.n312 585
R110 B.n314 B.n53 585
R111 B.n316 B.n315 585
R112 B.n317 B.n52 585
R113 B.n319 B.n318 585
R114 B.n320 B.n51 585
R115 B.n322 B.n321 585
R116 B.n323 B.n50 585
R117 B.n325 B.n324 585
R118 B.n326 B.n49 585
R119 B.n328 B.n327 585
R120 B.n329 B.n48 585
R121 B.n331 B.n330 585
R122 B.n332 B.n47 585
R123 B.n334 B.n333 585
R124 B.n335 B.n46 585
R125 B.n337 B.n336 585
R126 B.n407 B.n18 585
R127 B.n406 B.n405 585
R128 B.n404 B.n19 585
R129 B.n403 B.n402 585
R130 B.n401 B.n20 585
R131 B.n400 B.n399 585
R132 B.n398 B.n21 585
R133 B.n397 B.n396 585
R134 B.n395 B.n22 585
R135 B.n394 B.n393 585
R136 B.n392 B.n23 585
R137 B.n391 B.n390 585
R138 B.n389 B.n24 585
R139 B.n388 B.n387 585
R140 B.n386 B.n25 585
R141 B.n385 B.n384 585
R142 B.n383 B.n26 585
R143 B.n382 B.n381 585
R144 B.n379 B.n27 585
R145 B.n378 B.n377 585
R146 B.n376 B.n30 585
R147 B.n375 B.n374 585
R148 B.n373 B.n31 585
R149 B.n372 B.n371 585
R150 B.n370 B.n32 585
R151 B.n369 B.n368 585
R152 B.n367 B.n33 585
R153 B.n366 B.n365 585
R154 B.n364 B.n363 585
R155 B.n362 B.n37 585
R156 B.n361 B.n360 585
R157 B.n359 B.n38 585
R158 B.n358 B.n357 585
R159 B.n356 B.n39 585
R160 B.n355 B.n354 585
R161 B.n353 B.n40 585
R162 B.n352 B.n351 585
R163 B.n350 B.n41 585
R164 B.n349 B.n348 585
R165 B.n347 B.n42 585
R166 B.n346 B.n345 585
R167 B.n344 B.n43 585
R168 B.n343 B.n342 585
R169 B.n341 B.n44 585
R170 B.n340 B.n339 585
R171 B.n338 B.n45 585
R172 B.n409 B.n408 585
R173 B.n410 B.n17 585
R174 B.n412 B.n411 585
R175 B.n413 B.n16 585
R176 B.n415 B.n414 585
R177 B.n416 B.n15 585
R178 B.n418 B.n417 585
R179 B.n419 B.n14 585
R180 B.n421 B.n420 585
R181 B.n422 B.n13 585
R182 B.n424 B.n423 585
R183 B.n425 B.n12 585
R184 B.n427 B.n426 585
R185 B.n428 B.n11 585
R186 B.n430 B.n429 585
R187 B.n431 B.n10 585
R188 B.n433 B.n432 585
R189 B.n434 B.n9 585
R190 B.n436 B.n435 585
R191 B.n437 B.n8 585
R192 B.n439 B.n438 585
R193 B.n440 B.n7 585
R194 B.n442 B.n441 585
R195 B.n443 B.n6 585
R196 B.n445 B.n444 585
R197 B.n446 B.n5 585
R198 B.n448 B.n447 585
R199 B.n449 B.n4 585
R200 B.n451 B.n450 585
R201 B.n452 B.n3 585
R202 B.n454 B.n453 585
R203 B.n455 B.n0 585
R204 B.n2 B.n1 585
R205 B.n120 B.n119 585
R206 B.n121 B.n118 585
R207 B.n123 B.n122 585
R208 B.n124 B.n117 585
R209 B.n126 B.n125 585
R210 B.n127 B.n116 585
R211 B.n129 B.n128 585
R212 B.n130 B.n115 585
R213 B.n132 B.n131 585
R214 B.n133 B.n114 585
R215 B.n135 B.n134 585
R216 B.n136 B.n113 585
R217 B.n138 B.n137 585
R218 B.n139 B.n112 585
R219 B.n141 B.n140 585
R220 B.n142 B.n111 585
R221 B.n144 B.n143 585
R222 B.n145 B.n110 585
R223 B.n147 B.n146 585
R224 B.n148 B.n109 585
R225 B.n150 B.n149 585
R226 B.n151 B.n108 585
R227 B.n153 B.n152 585
R228 B.n154 B.n107 585
R229 B.n156 B.n155 585
R230 B.n157 B.n106 585
R231 B.n159 B.n158 585
R232 B.n160 B.n105 585
R233 B.n162 B.n161 585
R234 B.n163 B.n104 585
R235 B.n165 B.n164 585
R236 B.n164 B.n103 550.159
R237 B.n239 B.n238 550.159
R238 B.n336 B.n45 550.159
R239 B.n408 B.n407 550.159
R240 B.n457 B.n456 256.663
R241 B.n191 B.t3 235.292
R242 B.n88 B.t0 235.292
R243 B.n34 B.t9 235.292
R244 B.n28 B.t6 235.292
R245 B.n456 B.n455 235.042
R246 B.n456 B.n2 235.042
R247 B.n88 B.t1 200.469
R248 B.n34 B.t11 200.469
R249 B.n191 B.t4 200.464
R250 B.n28 B.t8 200.464
R251 B.n168 B.n103 163.367
R252 B.n169 B.n168 163.367
R253 B.n170 B.n169 163.367
R254 B.n170 B.n101 163.367
R255 B.n174 B.n101 163.367
R256 B.n175 B.n174 163.367
R257 B.n176 B.n175 163.367
R258 B.n176 B.n99 163.367
R259 B.n180 B.n99 163.367
R260 B.n181 B.n180 163.367
R261 B.n182 B.n181 163.367
R262 B.n182 B.n97 163.367
R263 B.n186 B.n97 163.367
R264 B.n187 B.n186 163.367
R265 B.n188 B.n187 163.367
R266 B.n188 B.n95 163.367
R267 B.n195 B.n95 163.367
R268 B.n196 B.n195 163.367
R269 B.n197 B.n196 163.367
R270 B.n197 B.n93 163.367
R271 B.n201 B.n93 163.367
R272 B.n202 B.n201 163.367
R273 B.n203 B.n202 163.367
R274 B.n203 B.n91 163.367
R275 B.n207 B.n91 163.367
R276 B.n208 B.n207 163.367
R277 B.n209 B.n208 163.367
R278 B.n209 B.n87 163.367
R279 B.n214 B.n87 163.367
R280 B.n215 B.n214 163.367
R281 B.n216 B.n215 163.367
R282 B.n216 B.n85 163.367
R283 B.n220 B.n85 163.367
R284 B.n221 B.n220 163.367
R285 B.n222 B.n221 163.367
R286 B.n222 B.n83 163.367
R287 B.n226 B.n83 163.367
R288 B.n227 B.n226 163.367
R289 B.n228 B.n227 163.367
R290 B.n228 B.n81 163.367
R291 B.n232 B.n81 163.367
R292 B.n233 B.n232 163.367
R293 B.n234 B.n233 163.367
R294 B.n234 B.n79 163.367
R295 B.n238 B.n79 163.367
R296 B.n336 B.n335 163.367
R297 B.n335 B.n334 163.367
R298 B.n334 B.n47 163.367
R299 B.n330 B.n47 163.367
R300 B.n330 B.n329 163.367
R301 B.n329 B.n328 163.367
R302 B.n328 B.n49 163.367
R303 B.n324 B.n49 163.367
R304 B.n324 B.n323 163.367
R305 B.n323 B.n322 163.367
R306 B.n322 B.n51 163.367
R307 B.n318 B.n51 163.367
R308 B.n318 B.n317 163.367
R309 B.n317 B.n316 163.367
R310 B.n316 B.n53 163.367
R311 B.n312 B.n53 163.367
R312 B.n312 B.n311 163.367
R313 B.n311 B.n310 163.367
R314 B.n310 B.n55 163.367
R315 B.n306 B.n55 163.367
R316 B.n306 B.n305 163.367
R317 B.n305 B.n304 163.367
R318 B.n304 B.n57 163.367
R319 B.n300 B.n57 163.367
R320 B.n300 B.n299 163.367
R321 B.n299 B.n298 163.367
R322 B.n298 B.n59 163.367
R323 B.n294 B.n59 163.367
R324 B.n294 B.n293 163.367
R325 B.n293 B.n292 163.367
R326 B.n292 B.n61 163.367
R327 B.n288 B.n61 163.367
R328 B.n288 B.n287 163.367
R329 B.n287 B.n286 163.367
R330 B.n286 B.n63 163.367
R331 B.n282 B.n63 163.367
R332 B.n282 B.n281 163.367
R333 B.n281 B.n280 163.367
R334 B.n280 B.n65 163.367
R335 B.n276 B.n65 163.367
R336 B.n276 B.n275 163.367
R337 B.n275 B.n274 163.367
R338 B.n274 B.n67 163.367
R339 B.n270 B.n67 163.367
R340 B.n270 B.n269 163.367
R341 B.n269 B.n268 163.367
R342 B.n268 B.n69 163.367
R343 B.n264 B.n69 163.367
R344 B.n264 B.n263 163.367
R345 B.n263 B.n262 163.367
R346 B.n262 B.n71 163.367
R347 B.n258 B.n71 163.367
R348 B.n258 B.n257 163.367
R349 B.n257 B.n256 163.367
R350 B.n256 B.n73 163.367
R351 B.n252 B.n73 163.367
R352 B.n252 B.n251 163.367
R353 B.n251 B.n250 163.367
R354 B.n250 B.n75 163.367
R355 B.n246 B.n75 163.367
R356 B.n246 B.n245 163.367
R357 B.n245 B.n244 163.367
R358 B.n244 B.n77 163.367
R359 B.n240 B.n77 163.367
R360 B.n240 B.n239 163.367
R361 B.n407 B.n406 163.367
R362 B.n406 B.n19 163.367
R363 B.n402 B.n19 163.367
R364 B.n402 B.n401 163.367
R365 B.n401 B.n400 163.367
R366 B.n400 B.n21 163.367
R367 B.n396 B.n21 163.367
R368 B.n396 B.n395 163.367
R369 B.n395 B.n394 163.367
R370 B.n394 B.n23 163.367
R371 B.n390 B.n23 163.367
R372 B.n390 B.n389 163.367
R373 B.n389 B.n388 163.367
R374 B.n388 B.n25 163.367
R375 B.n384 B.n25 163.367
R376 B.n384 B.n383 163.367
R377 B.n383 B.n382 163.367
R378 B.n382 B.n27 163.367
R379 B.n377 B.n27 163.367
R380 B.n377 B.n376 163.367
R381 B.n376 B.n375 163.367
R382 B.n375 B.n31 163.367
R383 B.n371 B.n31 163.367
R384 B.n371 B.n370 163.367
R385 B.n370 B.n369 163.367
R386 B.n369 B.n33 163.367
R387 B.n365 B.n33 163.367
R388 B.n365 B.n364 163.367
R389 B.n364 B.n37 163.367
R390 B.n360 B.n37 163.367
R391 B.n360 B.n359 163.367
R392 B.n359 B.n358 163.367
R393 B.n358 B.n39 163.367
R394 B.n354 B.n39 163.367
R395 B.n354 B.n353 163.367
R396 B.n353 B.n352 163.367
R397 B.n352 B.n41 163.367
R398 B.n348 B.n41 163.367
R399 B.n348 B.n347 163.367
R400 B.n347 B.n346 163.367
R401 B.n346 B.n43 163.367
R402 B.n342 B.n43 163.367
R403 B.n342 B.n341 163.367
R404 B.n341 B.n340 163.367
R405 B.n340 B.n45 163.367
R406 B.n408 B.n17 163.367
R407 B.n412 B.n17 163.367
R408 B.n413 B.n412 163.367
R409 B.n414 B.n413 163.367
R410 B.n414 B.n15 163.367
R411 B.n418 B.n15 163.367
R412 B.n419 B.n418 163.367
R413 B.n420 B.n419 163.367
R414 B.n420 B.n13 163.367
R415 B.n424 B.n13 163.367
R416 B.n425 B.n424 163.367
R417 B.n426 B.n425 163.367
R418 B.n426 B.n11 163.367
R419 B.n430 B.n11 163.367
R420 B.n431 B.n430 163.367
R421 B.n432 B.n431 163.367
R422 B.n432 B.n9 163.367
R423 B.n436 B.n9 163.367
R424 B.n437 B.n436 163.367
R425 B.n438 B.n437 163.367
R426 B.n438 B.n7 163.367
R427 B.n442 B.n7 163.367
R428 B.n443 B.n442 163.367
R429 B.n444 B.n443 163.367
R430 B.n444 B.n5 163.367
R431 B.n448 B.n5 163.367
R432 B.n449 B.n448 163.367
R433 B.n450 B.n449 163.367
R434 B.n450 B.n3 163.367
R435 B.n454 B.n3 163.367
R436 B.n455 B.n454 163.367
R437 B.n120 B.n2 163.367
R438 B.n121 B.n120 163.367
R439 B.n122 B.n121 163.367
R440 B.n122 B.n117 163.367
R441 B.n126 B.n117 163.367
R442 B.n127 B.n126 163.367
R443 B.n128 B.n127 163.367
R444 B.n128 B.n115 163.367
R445 B.n132 B.n115 163.367
R446 B.n133 B.n132 163.367
R447 B.n134 B.n133 163.367
R448 B.n134 B.n113 163.367
R449 B.n138 B.n113 163.367
R450 B.n139 B.n138 163.367
R451 B.n140 B.n139 163.367
R452 B.n140 B.n111 163.367
R453 B.n144 B.n111 163.367
R454 B.n145 B.n144 163.367
R455 B.n146 B.n145 163.367
R456 B.n146 B.n109 163.367
R457 B.n150 B.n109 163.367
R458 B.n151 B.n150 163.367
R459 B.n152 B.n151 163.367
R460 B.n152 B.n107 163.367
R461 B.n156 B.n107 163.367
R462 B.n157 B.n156 163.367
R463 B.n158 B.n157 163.367
R464 B.n158 B.n105 163.367
R465 B.n162 B.n105 163.367
R466 B.n163 B.n162 163.367
R467 B.n164 B.n163 163.367
R468 B.n89 B.t2 119.79
R469 B.n35 B.t10 119.79
R470 B.n192 B.t5 119.785
R471 B.n29 B.t7 119.785
R472 B.n192 B.n191 80.6793
R473 B.n89 B.n88 80.6793
R474 B.n35 B.n34 80.6793
R475 B.n29 B.n28 80.6793
R476 B.n193 B.n192 59.5399
R477 B.n211 B.n89 59.5399
R478 B.n36 B.n35 59.5399
R479 B.n380 B.n29 59.5399
R480 B.n409 B.n18 35.7468
R481 B.n338 B.n337 35.7468
R482 B.n166 B.n165 35.7468
R483 B.n237 B.n78 35.7468
R484 B B.n457 18.0485
R485 B.n410 B.n409 10.6151
R486 B.n411 B.n410 10.6151
R487 B.n411 B.n16 10.6151
R488 B.n415 B.n16 10.6151
R489 B.n416 B.n415 10.6151
R490 B.n417 B.n416 10.6151
R491 B.n417 B.n14 10.6151
R492 B.n421 B.n14 10.6151
R493 B.n422 B.n421 10.6151
R494 B.n423 B.n422 10.6151
R495 B.n423 B.n12 10.6151
R496 B.n427 B.n12 10.6151
R497 B.n428 B.n427 10.6151
R498 B.n429 B.n428 10.6151
R499 B.n429 B.n10 10.6151
R500 B.n433 B.n10 10.6151
R501 B.n434 B.n433 10.6151
R502 B.n435 B.n434 10.6151
R503 B.n435 B.n8 10.6151
R504 B.n439 B.n8 10.6151
R505 B.n440 B.n439 10.6151
R506 B.n441 B.n440 10.6151
R507 B.n441 B.n6 10.6151
R508 B.n445 B.n6 10.6151
R509 B.n446 B.n445 10.6151
R510 B.n447 B.n446 10.6151
R511 B.n447 B.n4 10.6151
R512 B.n451 B.n4 10.6151
R513 B.n452 B.n451 10.6151
R514 B.n453 B.n452 10.6151
R515 B.n453 B.n0 10.6151
R516 B.n405 B.n18 10.6151
R517 B.n405 B.n404 10.6151
R518 B.n404 B.n403 10.6151
R519 B.n403 B.n20 10.6151
R520 B.n399 B.n20 10.6151
R521 B.n399 B.n398 10.6151
R522 B.n398 B.n397 10.6151
R523 B.n397 B.n22 10.6151
R524 B.n393 B.n22 10.6151
R525 B.n393 B.n392 10.6151
R526 B.n392 B.n391 10.6151
R527 B.n391 B.n24 10.6151
R528 B.n387 B.n24 10.6151
R529 B.n387 B.n386 10.6151
R530 B.n386 B.n385 10.6151
R531 B.n385 B.n26 10.6151
R532 B.n381 B.n26 10.6151
R533 B.n379 B.n378 10.6151
R534 B.n378 B.n30 10.6151
R535 B.n374 B.n30 10.6151
R536 B.n374 B.n373 10.6151
R537 B.n373 B.n372 10.6151
R538 B.n372 B.n32 10.6151
R539 B.n368 B.n32 10.6151
R540 B.n368 B.n367 10.6151
R541 B.n367 B.n366 10.6151
R542 B.n363 B.n362 10.6151
R543 B.n362 B.n361 10.6151
R544 B.n361 B.n38 10.6151
R545 B.n357 B.n38 10.6151
R546 B.n357 B.n356 10.6151
R547 B.n356 B.n355 10.6151
R548 B.n355 B.n40 10.6151
R549 B.n351 B.n40 10.6151
R550 B.n351 B.n350 10.6151
R551 B.n350 B.n349 10.6151
R552 B.n349 B.n42 10.6151
R553 B.n345 B.n42 10.6151
R554 B.n345 B.n344 10.6151
R555 B.n344 B.n343 10.6151
R556 B.n343 B.n44 10.6151
R557 B.n339 B.n44 10.6151
R558 B.n339 B.n338 10.6151
R559 B.n337 B.n46 10.6151
R560 B.n333 B.n46 10.6151
R561 B.n333 B.n332 10.6151
R562 B.n332 B.n331 10.6151
R563 B.n331 B.n48 10.6151
R564 B.n327 B.n48 10.6151
R565 B.n327 B.n326 10.6151
R566 B.n326 B.n325 10.6151
R567 B.n325 B.n50 10.6151
R568 B.n321 B.n50 10.6151
R569 B.n321 B.n320 10.6151
R570 B.n320 B.n319 10.6151
R571 B.n319 B.n52 10.6151
R572 B.n315 B.n52 10.6151
R573 B.n315 B.n314 10.6151
R574 B.n314 B.n313 10.6151
R575 B.n313 B.n54 10.6151
R576 B.n309 B.n54 10.6151
R577 B.n309 B.n308 10.6151
R578 B.n308 B.n307 10.6151
R579 B.n307 B.n56 10.6151
R580 B.n303 B.n56 10.6151
R581 B.n303 B.n302 10.6151
R582 B.n302 B.n301 10.6151
R583 B.n301 B.n58 10.6151
R584 B.n297 B.n58 10.6151
R585 B.n297 B.n296 10.6151
R586 B.n296 B.n295 10.6151
R587 B.n295 B.n60 10.6151
R588 B.n291 B.n60 10.6151
R589 B.n291 B.n290 10.6151
R590 B.n290 B.n289 10.6151
R591 B.n289 B.n62 10.6151
R592 B.n285 B.n62 10.6151
R593 B.n285 B.n284 10.6151
R594 B.n284 B.n283 10.6151
R595 B.n283 B.n64 10.6151
R596 B.n279 B.n64 10.6151
R597 B.n279 B.n278 10.6151
R598 B.n278 B.n277 10.6151
R599 B.n277 B.n66 10.6151
R600 B.n273 B.n66 10.6151
R601 B.n273 B.n272 10.6151
R602 B.n272 B.n271 10.6151
R603 B.n271 B.n68 10.6151
R604 B.n267 B.n68 10.6151
R605 B.n267 B.n266 10.6151
R606 B.n266 B.n265 10.6151
R607 B.n265 B.n70 10.6151
R608 B.n261 B.n70 10.6151
R609 B.n261 B.n260 10.6151
R610 B.n260 B.n259 10.6151
R611 B.n259 B.n72 10.6151
R612 B.n255 B.n72 10.6151
R613 B.n255 B.n254 10.6151
R614 B.n254 B.n253 10.6151
R615 B.n253 B.n74 10.6151
R616 B.n249 B.n74 10.6151
R617 B.n249 B.n248 10.6151
R618 B.n248 B.n247 10.6151
R619 B.n247 B.n76 10.6151
R620 B.n243 B.n76 10.6151
R621 B.n243 B.n242 10.6151
R622 B.n242 B.n241 10.6151
R623 B.n241 B.n78 10.6151
R624 B.n119 B.n1 10.6151
R625 B.n119 B.n118 10.6151
R626 B.n123 B.n118 10.6151
R627 B.n124 B.n123 10.6151
R628 B.n125 B.n124 10.6151
R629 B.n125 B.n116 10.6151
R630 B.n129 B.n116 10.6151
R631 B.n130 B.n129 10.6151
R632 B.n131 B.n130 10.6151
R633 B.n131 B.n114 10.6151
R634 B.n135 B.n114 10.6151
R635 B.n136 B.n135 10.6151
R636 B.n137 B.n136 10.6151
R637 B.n137 B.n112 10.6151
R638 B.n141 B.n112 10.6151
R639 B.n142 B.n141 10.6151
R640 B.n143 B.n142 10.6151
R641 B.n143 B.n110 10.6151
R642 B.n147 B.n110 10.6151
R643 B.n148 B.n147 10.6151
R644 B.n149 B.n148 10.6151
R645 B.n149 B.n108 10.6151
R646 B.n153 B.n108 10.6151
R647 B.n154 B.n153 10.6151
R648 B.n155 B.n154 10.6151
R649 B.n155 B.n106 10.6151
R650 B.n159 B.n106 10.6151
R651 B.n160 B.n159 10.6151
R652 B.n161 B.n160 10.6151
R653 B.n161 B.n104 10.6151
R654 B.n165 B.n104 10.6151
R655 B.n167 B.n166 10.6151
R656 B.n167 B.n102 10.6151
R657 B.n171 B.n102 10.6151
R658 B.n172 B.n171 10.6151
R659 B.n173 B.n172 10.6151
R660 B.n173 B.n100 10.6151
R661 B.n177 B.n100 10.6151
R662 B.n178 B.n177 10.6151
R663 B.n179 B.n178 10.6151
R664 B.n179 B.n98 10.6151
R665 B.n183 B.n98 10.6151
R666 B.n184 B.n183 10.6151
R667 B.n185 B.n184 10.6151
R668 B.n185 B.n96 10.6151
R669 B.n189 B.n96 10.6151
R670 B.n190 B.n189 10.6151
R671 B.n194 B.n190 10.6151
R672 B.n198 B.n94 10.6151
R673 B.n199 B.n198 10.6151
R674 B.n200 B.n199 10.6151
R675 B.n200 B.n92 10.6151
R676 B.n204 B.n92 10.6151
R677 B.n205 B.n204 10.6151
R678 B.n206 B.n205 10.6151
R679 B.n206 B.n90 10.6151
R680 B.n210 B.n90 10.6151
R681 B.n213 B.n212 10.6151
R682 B.n213 B.n86 10.6151
R683 B.n217 B.n86 10.6151
R684 B.n218 B.n217 10.6151
R685 B.n219 B.n218 10.6151
R686 B.n219 B.n84 10.6151
R687 B.n223 B.n84 10.6151
R688 B.n224 B.n223 10.6151
R689 B.n225 B.n224 10.6151
R690 B.n225 B.n82 10.6151
R691 B.n229 B.n82 10.6151
R692 B.n230 B.n229 10.6151
R693 B.n231 B.n230 10.6151
R694 B.n231 B.n80 10.6151
R695 B.n235 B.n80 10.6151
R696 B.n236 B.n235 10.6151
R697 B.n237 B.n236 10.6151
R698 B.n381 B.n380 9.36635
R699 B.n363 B.n36 9.36635
R700 B.n194 B.n193 9.36635
R701 B.n212 B.n211 9.36635
R702 B.n457 B.n0 8.11757
R703 B.n457 B.n1 8.11757
R704 B.n380 B.n379 1.24928
R705 B.n366 B.n36 1.24928
R706 B.n193 B.n94 1.24928
R707 B.n211 B.n210 1.24928
R708 VN VN.t1 102.778
R709 VN VN.t0 61.6376
R710 VDD2.n0 VDD2.t1 149.108
R711 VDD2.n0 VDD2.t0 114.725
R712 VDD2 VDD2.n0 0.955241
C0 VDD1 VDD2 0.811165f
C1 VDD1 VN 0.153196f
C2 VDD1 VTAIL 3.35987f
C3 VDD2 VN 1.17596f
C4 VTAIL VDD2 3.42092f
C5 B w_n2634_n1792# 7.95272f
C6 VTAIL VN 1.44182f
C7 VP w_n2634_n1792# 3.9399f
C8 VDD1 w_n2634_n1792# 1.37963f
C9 B VP 1.72216f
C10 w_n2634_n1792# VDD2 1.4203f
C11 w_n2634_n1792# VN 3.60246f
C12 VTAIL w_n2634_n1792# 1.70159f
C13 VDD1 B 1.2299f
C14 B VDD2 1.27123f
C15 B VN 1.16143f
C16 VTAIL B 2.16824f
C17 VDD1 VP 1.41045f
C18 VP VDD2 0.389034f
C19 VP VN 4.57722f
C20 VTAIL VP 1.45616f
C21 VDD2 VSUBS 0.724464f
C22 VDD1 VSUBS 3.202942f
C23 VTAIL VSUBS 0.520826f
C24 VN VSUBS 5.98472f
C25 VP VSUBS 1.604712f
C26 B VSUBS 3.926878f
C27 w_n2634_n1792# VSUBS 59.391396f
C28 VDD2.t1 VSUBS 0.662733f
C29 VDD2.t0 VSUBS 0.429143f
C30 VDD2.n0 VSUBS 2.16361f
C31 VN.t0 VSUBS 1.92292f
C32 VN.t1 VSUBS 2.78819f
C33 B.n0 VSUBS 0.007759f
C34 B.n1 VSUBS 0.007759f
C35 B.n2 VSUBS 0.011475f
C36 B.n3 VSUBS 0.008794f
C37 B.n4 VSUBS 0.008794f
C38 B.n5 VSUBS 0.008794f
C39 B.n6 VSUBS 0.008794f
C40 B.n7 VSUBS 0.008794f
C41 B.n8 VSUBS 0.008794f
C42 B.n9 VSUBS 0.008794f
C43 B.n10 VSUBS 0.008794f
C44 B.n11 VSUBS 0.008794f
C45 B.n12 VSUBS 0.008794f
C46 B.n13 VSUBS 0.008794f
C47 B.n14 VSUBS 0.008794f
C48 B.n15 VSUBS 0.008794f
C49 B.n16 VSUBS 0.008794f
C50 B.n17 VSUBS 0.008794f
C51 B.n18 VSUBS 0.022191f
C52 B.n19 VSUBS 0.008794f
C53 B.n20 VSUBS 0.008794f
C54 B.n21 VSUBS 0.008794f
C55 B.n22 VSUBS 0.008794f
C56 B.n23 VSUBS 0.008794f
C57 B.n24 VSUBS 0.008794f
C58 B.n25 VSUBS 0.008794f
C59 B.n26 VSUBS 0.008794f
C60 B.n27 VSUBS 0.008794f
C61 B.t7 VSUBS 0.137348f
C62 B.t8 VSUBS 0.169572f
C63 B.t6 VSUBS 0.964718f
C64 B.n28 VSUBS 0.128703f
C65 B.n29 VSUBS 0.09261f
C66 B.n30 VSUBS 0.008794f
C67 B.n31 VSUBS 0.008794f
C68 B.n32 VSUBS 0.008794f
C69 B.n33 VSUBS 0.008794f
C70 B.t10 VSUBS 0.137348f
C71 B.t11 VSUBS 0.169571f
C72 B.t9 VSUBS 0.964718f
C73 B.n34 VSUBS 0.128703f
C74 B.n35 VSUBS 0.092609f
C75 B.n36 VSUBS 0.020374f
C76 B.n37 VSUBS 0.008794f
C77 B.n38 VSUBS 0.008794f
C78 B.n39 VSUBS 0.008794f
C79 B.n40 VSUBS 0.008794f
C80 B.n41 VSUBS 0.008794f
C81 B.n42 VSUBS 0.008794f
C82 B.n43 VSUBS 0.008794f
C83 B.n44 VSUBS 0.008794f
C84 B.n45 VSUBS 0.022191f
C85 B.n46 VSUBS 0.008794f
C86 B.n47 VSUBS 0.008794f
C87 B.n48 VSUBS 0.008794f
C88 B.n49 VSUBS 0.008794f
C89 B.n50 VSUBS 0.008794f
C90 B.n51 VSUBS 0.008794f
C91 B.n52 VSUBS 0.008794f
C92 B.n53 VSUBS 0.008794f
C93 B.n54 VSUBS 0.008794f
C94 B.n55 VSUBS 0.008794f
C95 B.n56 VSUBS 0.008794f
C96 B.n57 VSUBS 0.008794f
C97 B.n58 VSUBS 0.008794f
C98 B.n59 VSUBS 0.008794f
C99 B.n60 VSUBS 0.008794f
C100 B.n61 VSUBS 0.008794f
C101 B.n62 VSUBS 0.008794f
C102 B.n63 VSUBS 0.008794f
C103 B.n64 VSUBS 0.008794f
C104 B.n65 VSUBS 0.008794f
C105 B.n66 VSUBS 0.008794f
C106 B.n67 VSUBS 0.008794f
C107 B.n68 VSUBS 0.008794f
C108 B.n69 VSUBS 0.008794f
C109 B.n70 VSUBS 0.008794f
C110 B.n71 VSUBS 0.008794f
C111 B.n72 VSUBS 0.008794f
C112 B.n73 VSUBS 0.008794f
C113 B.n74 VSUBS 0.008794f
C114 B.n75 VSUBS 0.008794f
C115 B.n76 VSUBS 0.008794f
C116 B.n77 VSUBS 0.008794f
C117 B.n78 VSUBS 0.022468f
C118 B.n79 VSUBS 0.008794f
C119 B.n80 VSUBS 0.008794f
C120 B.n81 VSUBS 0.008794f
C121 B.n82 VSUBS 0.008794f
C122 B.n83 VSUBS 0.008794f
C123 B.n84 VSUBS 0.008794f
C124 B.n85 VSUBS 0.008794f
C125 B.n86 VSUBS 0.008794f
C126 B.n87 VSUBS 0.008794f
C127 B.t2 VSUBS 0.137348f
C128 B.t1 VSUBS 0.169571f
C129 B.t0 VSUBS 0.964718f
C130 B.n88 VSUBS 0.128703f
C131 B.n89 VSUBS 0.092609f
C132 B.n90 VSUBS 0.008794f
C133 B.n91 VSUBS 0.008794f
C134 B.n92 VSUBS 0.008794f
C135 B.n93 VSUBS 0.008794f
C136 B.n94 VSUBS 0.004914f
C137 B.n95 VSUBS 0.008794f
C138 B.n96 VSUBS 0.008794f
C139 B.n97 VSUBS 0.008794f
C140 B.n98 VSUBS 0.008794f
C141 B.n99 VSUBS 0.008794f
C142 B.n100 VSUBS 0.008794f
C143 B.n101 VSUBS 0.008794f
C144 B.n102 VSUBS 0.008794f
C145 B.n103 VSUBS 0.022191f
C146 B.n104 VSUBS 0.008794f
C147 B.n105 VSUBS 0.008794f
C148 B.n106 VSUBS 0.008794f
C149 B.n107 VSUBS 0.008794f
C150 B.n108 VSUBS 0.008794f
C151 B.n109 VSUBS 0.008794f
C152 B.n110 VSUBS 0.008794f
C153 B.n111 VSUBS 0.008794f
C154 B.n112 VSUBS 0.008794f
C155 B.n113 VSUBS 0.008794f
C156 B.n114 VSUBS 0.008794f
C157 B.n115 VSUBS 0.008794f
C158 B.n116 VSUBS 0.008794f
C159 B.n117 VSUBS 0.008794f
C160 B.n118 VSUBS 0.008794f
C161 B.n119 VSUBS 0.008794f
C162 B.n120 VSUBS 0.008794f
C163 B.n121 VSUBS 0.008794f
C164 B.n122 VSUBS 0.008794f
C165 B.n123 VSUBS 0.008794f
C166 B.n124 VSUBS 0.008794f
C167 B.n125 VSUBS 0.008794f
C168 B.n126 VSUBS 0.008794f
C169 B.n127 VSUBS 0.008794f
C170 B.n128 VSUBS 0.008794f
C171 B.n129 VSUBS 0.008794f
C172 B.n130 VSUBS 0.008794f
C173 B.n131 VSUBS 0.008794f
C174 B.n132 VSUBS 0.008794f
C175 B.n133 VSUBS 0.008794f
C176 B.n134 VSUBS 0.008794f
C177 B.n135 VSUBS 0.008794f
C178 B.n136 VSUBS 0.008794f
C179 B.n137 VSUBS 0.008794f
C180 B.n138 VSUBS 0.008794f
C181 B.n139 VSUBS 0.008794f
C182 B.n140 VSUBS 0.008794f
C183 B.n141 VSUBS 0.008794f
C184 B.n142 VSUBS 0.008794f
C185 B.n143 VSUBS 0.008794f
C186 B.n144 VSUBS 0.008794f
C187 B.n145 VSUBS 0.008794f
C188 B.n146 VSUBS 0.008794f
C189 B.n147 VSUBS 0.008794f
C190 B.n148 VSUBS 0.008794f
C191 B.n149 VSUBS 0.008794f
C192 B.n150 VSUBS 0.008794f
C193 B.n151 VSUBS 0.008794f
C194 B.n152 VSUBS 0.008794f
C195 B.n153 VSUBS 0.008794f
C196 B.n154 VSUBS 0.008794f
C197 B.n155 VSUBS 0.008794f
C198 B.n156 VSUBS 0.008794f
C199 B.n157 VSUBS 0.008794f
C200 B.n158 VSUBS 0.008794f
C201 B.n159 VSUBS 0.008794f
C202 B.n160 VSUBS 0.008794f
C203 B.n161 VSUBS 0.008794f
C204 B.n162 VSUBS 0.008794f
C205 B.n163 VSUBS 0.008794f
C206 B.n164 VSUBS 0.021519f
C207 B.n165 VSUBS 0.021519f
C208 B.n166 VSUBS 0.022191f
C209 B.n167 VSUBS 0.008794f
C210 B.n168 VSUBS 0.008794f
C211 B.n169 VSUBS 0.008794f
C212 B.n170 VSUBS 0.008794f
C213 B.n171 VSUBS 0.008794f
C214 B.n172 VSUBS 0.008794f
C215 B.n173 VSUBS 0.008794f
C216 B.n174 VSUBS 0.008794f
C217 B.n175 VSUBS 0.008794f
C218 B.n176 VSUBS 0.008794f
C219 B.n177 VSUBS 0.008794f
C220 B.n178 VSUBS 0.008794f
C221 B.n179 VSUBS 0.008794f
C222 B.n180 VSUBS 0.008794f
C223 B.n181 VSUBS 0.008794f
C224 B.n182 VSUBS 0.008794f
C225 B.n183 VSUBS 0.008794f
C226 B.n184 VSUBS 0.008794f
C227 B.n185 VSUBS 0.008794f
C228 B.n186 VSUBS 0.008794f
C229 B.n187 VSUBS 0.008794f
C230 B.n188 VSUBS 0.008794f
C231 B.n189 VSUBS 0.008794f
C232 B.n190 VSUBS 0.008794f
C233 B.t5 VSUBS 0.137348f
C234 B.t4 VSUBS 0.169572f
C235 B.t3 VSUBS 0.964718f
C236 B.n191 VSUBS 0.128703f
C237 B.n192 VSUBS 0.09261f
C238 B.n193 VSUBS 0.020374f
C239 B.n194 VSUBS 0.008276f
C240 B.n195 VSUBS 0.008794f
C241 B.n196 VSUBS 0.008794f
C242 B.n197 VSUBS 0.008794f
C243 B.n198 VSUBS 0.008794f
C244 B.n199 VSUBS 0.008794f
C245 B.n200 VSUBS 0.008794f
C246 B.n201 VSUBS 0.008794f
C247 B.n202 VSUBS 0.008794f
C248 B.n203 VSUBS 0.008794f
C249 B.n204 VSUBS 0.008794f
C250 B.n205 VSUBS 0.008794f
C251 B.n206 VSUBS 0.008794f
C252 B.n207 VSUBS 0.008794f
C253 B.n208 VSUBS 0.008794f
C254 B.n209 VSUBS 0.008794f
C255 B.n210 VSUBS 0.004914f
C256 B.n211 VSUBS 0.020374f
C257 B.n212 VSUBS 0.008276f
C258 B.n213 VSUBS 0.008794f
C259 B.n214 VSUBS 0.008794f
C260 B.n215 VSUBS 0.008794f
C261 B.n216 VSUBS 0.008794f
C262 B.n217 VSUBS 0.008794f
C263 B.n218 VSUBS 0.008794f
C264 B.n219 VSUBS 0.008794f
C265 B.n220 VSUBS 0.008794f
C266 B.n221 VSUBS 0.008794f
C267 B.n222 VSUBS 0.008794f
C268 B.n223 VSUBS 0.008794f
C269 B.n224 VSUBS 0.008794f
C270 B.n225 VSUBS 0.008794f
C271 B.n226 VSUBS 0.008794f
C272 B.n227 VSUBS 0.008794f
C273 B.n228 VSUBS 0.008794f
C274 B.n229 VSUBS 0.008794f
C275 B.n230 VSUBS 0.008794f
C276 B.n231 VSUBS 0.008794f
C277 B.n232 VSUBS 0.008794f
C278 B.n233 VSUBS 0.008794f
C279 B.n234 VSUBS 0.008794f
C280 B.n235 VSUBS 0.008794f
C281 B.n236 VSUBS 0.008794f
C282 B.n237 VSUBS 0.021241f
C283 B.n238 VSUBS 0.022191f
C284 B.n239 VSUBS 0.021519f
C285 B.n240 VSUBS 0.008794f
C286 B.n241 VSUBS 0.008794f
C287 B.n242 VSUBS 0.008794f
C288 B.n243 VSUBS 0.008794f
C289 B.n244 VSUBS 0.008794f
C290 B.n245 VSUBS 0.008794f
C291 B.n246 VSUBS 0.008794f
C292 B.n247 VSUBS 0.008794f
C293 B.n248 VSUBS 0.008794f
C294 B.n249 VSUBS 0.008794f
C295 B.n250 VSUBS 0.008794f
C296 B.n251 VSUBS 0.008794f
C297 B.n252 VSUBS 0.008794f
C298 B.n253 VSUBS 0.008794f
C299 B.n254 VSUBS 0.008794f
C300 B.n255 VSUBS 0.008794f
C301 B.n256 VSUBS 0.008794f
C302 B.n257 VSUBS 0.008794f
C303 B.n258 VSUBS 0.008794f
C304 B.n259 VSUBS 0.008794f
C305 B.n260 VSUBS 0.008794f
C306 B.n261 VSUBS 0.008794f
C307 B.n262 VSUBS 0.008794f
C308 B.n263 VSUBS 0.008794f
C309 B.n264 VSUBS 0.008794f
C310 B.n265 VSUBS 0.008794f
C311 B.n266 VSUBS 0.008794f
C312 B.n267 VSUBS 0.008794f
C313 B.n268 VSUBS 0.008794f
C314 B.n269 VSUBS 0.008794f
C315 B.n270 VSUBS 0.008794f
C316 B.n271 VSUBS 0.008794f
C317 B.n272 VSUBS 0.008794f
C318 B.n273 VSUBS 0.008794f
C319 B.n274 VSUBS 0.008794f
C320 B.n275 VSUBS 0.008794f
C321 B.n276 VSUBS 0.008794f
C322 B.n277 VSUBS 0.008794f
C323 B.n278 VSUBS 0.008794f
C324 B.n279 VSUBS 0.008794f
C325 B.n280 VSUBS 0.008794f
C326 B.n281 VSUBS 0.008794f
C327 B.n282 VSUBS 0.008794f
C328 B.n283 VSUBS 0.008794f
C329 B.n284 VSUBS 0.008794f
C330 B.n285 VSUBS 0.008794f
C331 B.n286 VSUBS 0.008794f
C332 B.n287 VSUBS 0.008794f
C333 B.n288 VSUBS 0.008794f
C334 B.n289 VSUBS 0.008794f
C335 B.n290 VSUBS 0.008794f
C336 B.n291 VSUBS 0.008794f
C337 B.n292 VSUBS 0.008794f
C338 B.n293 VSUBS 0.008794f
C339 B.n294 VSUBS 0.008794f
C340 B.n295 VSUBS 0.008794f
C341 B.n296 VSUBS 0.008794f
C342 B.n297 VSUBS 0.008794f
C343 B.n298 VSUBS 0.008794f
C344 B.n299 VSUBS 0.008794f
C345 B.n300 VSUBS 0.008794f
C346 B.n301 VSUBS 0.008794f
C347 B.n302 VSUBS 0.008794f
C348 B.n303 VSUBS 0.008794f
C349 B.n304 VSUBS 0.008794f
C350 B.n305 VSUBS 0.008794f
C351 B.n306 VSUBS 0.008794f
C352 B.n307 VSUBS 0.008794f
C353 B.n308 VSUBS 0.008794f
C354 B.n309 VSUBS 0.008794f
C355 B.n310 VSUBS 0.008794f
C356 B.n311 VSUBS 0.008794f
C357 B.n312 VSUBS 0.008794f
C358 B.n313 VSUBS 0.008794f
C359 B.n314 VSUBS 0.008794f
C360 B.n315 VSUBS 0.008794f
C361 B.n316 VSUBS 0.008794f
C362 B.n317 VSUBS 0.008794f
C363 B.n318 VSUBS 0.008794f
C364 B.n319 VSUBS 0.008794f
C365 B.n320 VSUBS 0.008794f
C366 B.n321 VSUBS 0.008794f
C367 B.n322 VSUBS 0.008794f
C368 B.n323 VSUBS 0.008794f
C369 B.n324 VSUBS 0.008794f
C370 B.n325 VSUBS 0.008794f
C371 B.n326 VSUBS 0.008794f
C372 B.n327 VSUBS 0.008794f
C373 B.n328 VSUBS 0.008794f
C374 B.n329 VSUBS 0.008794f
C375 B.n330 VSUBS 0.008794f
C376 B.n331 VSUBS 0.008794f
C377 B.n332 VSUBS 0.008794f
C378 B.n333 VSUBS 0.008794f
C379 B.n334 VSUBS 0.008794f
C380 B.n335 VSUBS 0.008794f
C381 B.n336 VSUBS 0.021519f
C382 B.n337 VSUBS 0.021519f
C383 B.n338 VSUBS 0.022191f
C384 B.n339 VSUBS 0.008794f
C385 B.n340 VSUBS 0.008794f
C386 B.n341 VSUBS 0.008794f
C387 B.n342 VSUBS 0.008794f
C388 B.n343 VSUBS 0.008794f
C389 B.n344 VSUBS 0.008794f
C390 B.n345 VSUBS 0.008794f
C391 B.n346 VSUBS 0.008794f
C392 B.n347 VSUBS 0.008794f
C393 B.n348 VSUBS 0.008794f
C394 B.n349 VSUBS 0.008794f
C395 B.n350 VSUBS 0.008794f
C396 B.n351 VSUBS 0.008794f
C397 B.n352 VSUBS 0.008794f
C398 B.n353 VSUBS 0.008794f
C399 B.n354 VSUBS 0.008794f
C400 B.n355 VSUBS 0.008794f
C401 B.n356 VSUBS 0.008794f
C402 B.n357 VSUBS 0.008794f
C403 B.n358 VSUBS 0.008794f
C404 B.n359 VSUBS 0.008794f
C405 B.n360 VSUBS 0.008794f
C406 B.n361 VSUBS 0.008794f
C407 B.n362 VSUBS 0.008794f
C408 B.n363 VSUBS 0.008276f
C409 B.n364 VSUBS 0.008794f
C410 B.n365 VSUBS 0.008794f
C411 B.n366 VSUBS 0.004914f
C412 B.n367 VSUBS 0.008794f
C413 B.n368 VSUBS 0.008794f
C414 B.n369 VSUBS 0.008794f
C415 B.n370 VSUBS 0.008794f
C416 B.n371 VSUBS 0.008794f
C417 B.n372 VSUBS 0.008794f
C418 B.n373 VSUBS 0.008794f
C419 B.n374 VSUBS 0.008794f
C420 B.n375 VSUBS 0.008794f
C421 B.n376 VSUBS 0.008794f
C422 B.n377 VSUBS 0.008794f
C423 B.n378 VSUBS 0.008794f
C424 B.n379 VSUBS 0.004914f
C425 B.n380 VSUBS 0.020374f
C426 B.n381 VSUBS 0.008276f
C427 B.n382 VSUBS 0.008794f
C428 B.n383 VSUBS 0.008794f
C429 B.n384 VSUBS 0.008794f
C430 B.n385 VSUBS 0.008794f
C431 B.n386 VSUBS 0.008794f
C432 B.n387 VSUBS 0.008794f
C433 B.n388 VSUBS 0.008794f
C434 B.n389 VSUBS 0.008794f
C435 B.n390 VSUBS 0.008794f
C436 B.n391 VSUBS 0.008794f
C437 B.n392 VSUBS 0.008794f
C438 B.n393 VSUBS 0.008794f
C439 B.n394 VSUBS 0.008794f
C440 B.n395 VSUBS 0.008794f
C441 B.n396 VSUBS 0.008794f
C442 B.n397 VSUBS 0.008794f
C443 B.n398 VSUBS 0.008794f
C444 B.n399 VSUBS 0.008794f
C445 B.n400 VSUBS 0.008794f
C446 B.n401 VSUBS 0.008794f
C447 B.n402 VSUBS 0.008794f
C448 B.n403 VSUBS 0.008794f
C449 B.n404 VSUBS 0.008794f
C450 B.n405 VSUBS 0.008794f
C451 B.n406 VSUBS 0.008794f
C452 B.n407 VSUBS 0.022191f
C453 B.n408 VSUBS 0.021519f
C454 B.n409 VSUBS 0.021519f
C455 B.n410 VSUBS 0.008794f
C456 B.n411 VSUBS 0.008794f
C457 B.n412 VSUBS 0.008794f
C458 B.n413 VSUBS 0.008794f
C459 B.n414 VSUBS 0.008794f
C460 B.n415 VSUBS 0.008794f
C461 B.n416 VSUBS 0.008794f
C462 B.n417 VSUBS 0.008794f
C463 B.n418 VSUBS 0.008794f
C464 B.n419 VSUBS 0.008794f
C465 B.n420 VSUBS 0.008794f
C466 B.n421 VSUBS 0.008794f
C467 B.n422 VSUBS 0.008794f
C468 B.n423 VSUBS 0.008794f
C469 B.n424 VSUBS 0.008794f
C470 B.n425 VSUBS 0.008794f
C471 B.n426 VSUBS 0.008794f
C472 B.n427 VSUBS 0.008794f
C473 B.n428 VSUBS 0.008794f
C474 B.n429 VSUBS 0.008794f
C475 B.n430 VSUBS 0.008794f
C476 B.n431 VSUBS 0.008794f
C477 B.n432 VSUBS 0.008794f
C478 B.n433 VSUBS 0.008794f
C479 B.n434 VSUBS 0.008794f
C480 B.n435 VSUBS 0.008794f
C481 B.n436 VSUBS 0.008794f
C482 B.n437 VSUBS 0.008794f
C483 B.n438 VSUBS 0.008794f
C484 B.n439 VSUBS 0.008794f
C485 B.n440 VSUBS 0.008794f
C486 B.n441 VSUBS 0.008794f
C487 B.n442 VSUBS 0.008794f
C488 B.n443 VSUBS 0.008794f
C489 B.n444 VSUBS 0.008794f
C490 B.n445 VSUBS 0.008794f
C491 B.n446 VSUBS 0.008794f
C492 B.n447 VSUBS 0.008794f
C493 B.n448 VSUBS 0.008794f
C494 B.n449 VSUBS 0.008794f
C495 B.n450 VSUBS 0.008794f
C496 B.n451 VSUBS 0.008794f
C497 B.n452 VSUBS 0.008794f
C498 B.n453 VSUBS 0.008794f
C499 B.n454 VSUBS 0.008794f
C500 B.n455 VSUBS 0.011475f
C501 B.n456 VSUBS 0.012224f
C502 B.n457 VSUBS 0.024309f
C503 VDD1.t1 VSUBS 0.424263f
C504 VDD1.t0 VSUBS 0.672708f
C505 VTAIL.t2 VSUBS 0.587471f
C506 VTAIL.n0 VSUBS 1.73885f
C507 VTAIL.t0 VSUBS 0.587473f
C508 VTAIL.n1 VSUBS 1.80586f
C509 VTAIL.t3 VSUBS 0.587471f
C510 VTAIL.n2 VSUBS 1.51919f
C511 VTAIL.t1 VSUBS 0.587471f
C512 VTAIL.n3 VSUBS 1.40532f
C513 VP.t0 VSUBS 2.9094f
C514 VP.t1 VSUBS 1.99859f
C515 VP.n0 VSUBS 3.43435f
.ends

