* NGSPICE file created from diff_pair_sample_1530.ext - technology: sky130A

.subckt diff_pair_sample_1530 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1270_n2568# sky130_fd_pr__pfet_01v8 ad=3.1122 pd=16.74 as=0 ps=0 w=7.98 l=0.42
X1 B.t8 B.t6 B.t7 w_n1270_n2568# sky130_fd_pr__pfet_01v8 ad=3.1122 pd=16.74 as=0 ps=0 w=7.98 l=0.42
X2 VDD1.t1 VP.t0 VTAIL.t2 w_n1270_n2568# sky130_fd_pr__pfet_01v8 ad=3.1122 pd=16.74 as=3.1122 ps=16.74 w=7.98 l=0.42
X3 B.t5 B.t3 B.t4 w_n1270_n2568# sky130_fd_pr__pfet_01v8 ad=3.1122 pd=16.74 as=0 ps=0 w=7.98 l=0.42
X4 VDD2.t1 VN.t0 VTAIL.t1 w_n1270_n2568# sky130_fd_pr__pfet_01v8 ad=3.1122 pd=16.74 as=3.1122 ps=16.74 w=7.98 l=0.42
X5 B.t2 B.t0 B.t1 w_n1270_n2568# sky130_fd_pr__pfet_01v8 ad=3.1122 pd=16.74 as=0 ps=0 w=7.98 l=0.42
X6 VDD1.t0 VP.t1 VTAIL.t3 w_n1270_n2568# sky130_fd_pr__pfet_01v8 ad=3.1122 pd=16.74 as=3.1122 ps=16.74 w=7.98 l=0.42
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n1270_n2568# sky130_fd_pr__pfet_01v8 ad=3.1122 pd=16.74 as=3.1122 ps=16.74 w=7.98 l=0.42
R0 B.n80 B.t0 666.604
R1 B.n176 B.t3 666.604
R2 B.n30 B.t9 666.604
R3 B.n24 B.t6 666.604
R4 B.n225 B.n224 585
R5 B.n223 B.n60 585
R6 B.n222 B.n221 585
R7 B.n220 B.n61 585
R8 B.n219 B.n218 585
R9 B.n217 B.n62 585
R10 B.n216 B.n215 585
R11 B.n214 B.n63 585
R12 B.n213 B.n212 585
R13 B.n211 B.n64 585
R14 B.n210 B.n209 585
R15 B.n208 B.n65 585
R16 B.n207 B.n206 585
R17 B.n205 B.n66 585
R18 B.n204 B.n203 585
R19 B.n202 B.n67 585
R20 B.n201 B.n200 585
R21 B.n199 B.n68 585
R22 B.n198 B.n197 585
R23 B.n196 B.n69 585
R24 B.n195 B.n194 585
R25 B.n193 B.n70 585
R26 B.n192 B.n191 585
R27 B.n190 B.n71 585
R28 B.n189 B.n188 585
R29 B.n187 B.n72 585
R30 B.n186 B.n185 585
R31 B.n184 B.n73 585
R32 B.n183 B.n182 585
R33 B.n181 B.n74 585
R34 B.n180 B.n179 585
R35 B.n175 B.n75 585
R36 B.n174 B.n173 585
R37 B.n172 B.n76 585
R38 B.n171 B.n170 585
R39 B.n169 B.n77 585
R40 B.n168 B.n167 585
R41 B.n166 B.n78 585
R42 B.n165 B.n164 585
R43 B.n162 B.n79 585
R44 B.n161 B.n160 585
R45 B.n159 B.n82 585
R46 B.n158 B.n157 585
R47 B.n156 B.n83 585
R48 B.n155 B.n154 585
R49 B.n153 B.n84 585
R50 B.n152 B.n151 585
R51 B.n150 B.n85 585
R52 B.n149 B.n148 585
R53 B.n147 B.n86 585
R54 B.n146 B.n145 585
R55 B.n144 B.n87 585
R56 B.n143 B.n142 585
R57 B.n141 B.n88 585
R58 B.n140 B.n139 585
R59 B.n138 B.n89 585
R60 B.n137 B.n136 585
R61 B.n135 B.n90 585
R62 B.n134 B.n133 585
R63 B.n132 B.n91 585
R64 B.n131 B.n130 585
R65 B.n129 B.n92 585
R66 B.n128 B.n127 585
R67 B.n126 B.n93 585
R68 B.n125 B.n124 585
R69 B.n123 B.n94 585
R70 B.n122 B.n121 585
R71 B.n120 B.n95 585
R72 B.n119 B.n118 585
R73 B.n226 B.n59 585
R74 B.n228 B.n227 585
R75 B.n229 B.n58 585
R76 B.n231 B.n230 585
R77 B.n232 B.n57 585
R78 B.n234 B.n233 585
R79 B.n235 B.n56 585
R80 B.n237 B.n236 585
R81 B.n238 B.n55 585
R82 B.n240 B.n239 585
R83 B.n241 B.n54 585
R84 B.n243 B.n242 585
R85 B.n244 B.n53 585
R86 B.n246 B.n245 585
R87 B.n247 B.n52 585
R88 B.n249 B.n248 585
R89 B.n250 B.n51 585
R90 B.n252 B.n251 585
R91 B.n253 B.n50 585
R92 B.n255 B.n254 585
R93 B.n256 B.n49 585
R94 B.n258 B.n257 585
R95 B.n259 B.n48 585
R96 B.n261 B.n260 585
R97 B.n262 B.n47 585
R98 B.n264 B.n263 585
R99 B.n369 B.n8 585
R100 B.n368 B.n367 585
R101 B.n366 B.n9 585
R102 B.n365 B.n364 585
R103 B.n363 B.n10 585
R104 B.n362 B.n361 585
R105 B.n360 B.n11 585
R106 B.n359 B.n358 585
R107 B.n357 B.n12 585
R108 B.n356 B.n355 585
R109 B.n354 B.n13 585
R110 B.n353 B.n352 585
R111 B.n351 B.n14 585
R112 B.n350 B.n349 585
R113 B.n348 B.n15 585
R114 B.n347 B.n346 585
R115 B.n345 B.n16 585
R116 B.n344 B.n343 585
R117 B.n342 B.n17 585
R118 B.n341 B.n340 585
R119 B.n339 B.n18 585
R120 B.n338 B.n337 585
R121 B.n336 B.n19 585
R122 B.n335 B.n334 585
R123 B.n333 B.n20 585
R124 B.n332 B.n331 585
R125 B.n330 B.n21 585
R126 B.n329 B.n328 585
R127 B.n327 B.n22 585
R128 B.n326 B.n325 585
R129 B.n323 B.n23 585
R130 B.n322 B.n321 585
R131 B.n320 B.n26 585
R132 B.n319 B.n318 585
R133 B.n317 B.n27 585
R134 B.n316 B.n315 585
R135 B.n314 B.n28 585
R136 B.n313 B.n312 585
R137 B.n311 B.n29 585
R138 B.n309 B.n308 585
R139 B.n307 B.n32 585
R140 B.n306 B.n305 585
R141 B.n304 B.n33 585
R142 B.n303 B.n302 585
R143 B.n301 B.n34 585
R144 B.n300 B.n299 585
R145 B.n298 B.n35 585
R146 B.n297 B.n296 585
R147 B.n295 B.n36 585
R148 B.n294 B.n293 585
R149 B.n292 B.n37 585
R150 B.n291 B.n290 585
R151 B.n289 B.n38 585
R152 B.n288 B.n287 585
R153 B.n286 B.n39 585
R154 B.n285 B.n284 585
R155 B.n283 B.n40 585
R156 B.n282 B.n281 585
R157 B.n280 B.n41 585
R158 B.n279 B.n278 585
R159 B.n277 B.n42 585
R160 B.n276 B.n275 585
R161 B.n274 B.n43 585
R162 B.n273 B.n272 585
R163 B.n271 B.n44 585
R164 B.n270 B.n269 585
R165 B.n268 B.n45 585
R166 B.n267 B.n266 585
R167 B.n265 B.n46 585
R168 B.n371 B.n370 585
R169 B.n372 B.n7 585
R170 B.n374 B.n373 585
R171 B.n375 B.n6 585
R172 B.n377 B.n376 585
R173 B.n378 B.n5 585
R174 B.n380 B.n379 585
R175 B.n381 B.n4 585
R176 B.n383 B.n382 585
R177 B.n384 B.n3 585
R178 B.n386 B.n385 585
R179 B.n387 B.n0 585
R180 B.n2 B.n1 585
R181 B.n102 B.n101 585
R182 B.n104 B.n103 585
R183 B.n105 B.n100 585
R184 B.n107 B.n106 585
R185 B.n108 B.n99 585
R186 B.n110 B.n109 585
R187 B.n111 B.n98 585
R188 B.n113 B.n112 585
R189 B.n114 B.n97 585
R190 B.n116 B.n115 585
R191 B.n117 B.n96 585
R192 B.n118 B.n117 526.135
R193 B.n224 B.n59 526.135
R194 B.n265 B.n264 526.135
R195 B.n370 B.n369 526.135
R196 B.n176 B.t4 317.848
R197 B.n30 B.t11 317.848
R198 B.n80 B.t1 317.848
R199 B.n24 B.t8 317.848
R200 B.n177 B.t5 303.303
R201 B.n31 B.t10 303.303
R202 B.n81 B.t2 303.303
R203 B.n25 B.t7 303.303
R204 B.n389 B.n388 256.663
R205 B.n388 B.n387 235.042
R206 B.n388 B.n2 235.042
R207 B.n118 B.n95 163.367
R208 B.n122 B.n95 163.367
R209 B.n123 B.n122 163.367
R210 B.n124 B.n123 163.367
R211 B.n124 B.n93 163.367
R212 B.n128 B.n93 163.367
R213 B.n129 B.n128 163.367
R214 B.n130 B.n129 163.367
R215 B.n130 B.n91 163.367
R216 B.n134 B.n91 163.367
R217 B.n135 B.n134 163.367
R218 B.n136 B.n135 163.367
R219 B.n136 B.n89 163.367
R220 B.n140 B.n89 163.367
R221 B.n141 B.n140 163.367
R222 B.n142 B.n141 163.367
R223 B.n142 B.n87 163.367
R224 B.n146 B.n87 163.367
R225 B.n147 B.n146 163.367
R226 B.n148 B.n147 163.367
R227 B.n148 B.n85 163.367
R228 B.n152 B.n85 163.367
R229 B.n153 B.n152 163.367
R230 B.n154 B.n153 163.367
R231 B.n154 B.n83 163.367
R232 B.n158 B.n83 163.367
R233 B.n159 B.n158 163.367
R234 B.n160 B.n159 163.367
R235 B.n160 B.n79 163.367
R236 B.n165 B.n79 163.367
R237 B.n166 B.n165 163.367
R238 B.n167 B.n166 163.367
R239 B.n167 B.n77 163.367
R240 B.n171 B.n77 163.367
R241 B.n172 B.n171 163.367
R242 B.n173 B.n172 163.367
R243 B.n173 B.n75 163.367
R244 B.n180 B.n75 163.367
R245 B.n181 B.n180 163.367
R246 B.n182 B.n181 163.367
R247 B.n182 B.n73 163.367
R248 B.n186 B.n73 163.367
R249 B.n187 B.n186 163.367
R250 B.n188 B.n187 163.367
R251 B.n188 B.n71 163.367
R252 B.n192 B.n71 163.367
R253 B.n193 B.n192 163.367
R254 B.n194 B.n193 163.367
R255 B.n194 B.n69 163.367
R256 B.n198 B.n69 163.367
R257 B.n199 B.n198 163.367
R258 B.n200 B.n199 163.367
R259 B.n200 B.n67 163.367
R260 B.n204 B.n67 163.367
R261 B.n205 B.n204 163.367
R262 B.n206 B.n205 163.367
R263 B.n206 B.n65 163.367
R264 B.n210 B.n65 163.367
R265 B.n211 B.n210 163.367
R266 B.n212 B.n211 163.367
R267 B.n212 B.n63 163.367
R268 B.n216 B.n63 163.367
R269 B.n217 B.n216 163.367
R270 B.n218 B.n217 163.367
R271 B.n218 B.n61 163.367
R272 B.n222 B.n61 163.367
R273 B.n223 B.n222 163.367
R274 B.n224 B.n223 163.367
R275 B.n264 B.n47 163.367
R276 B.n260 B.n47 163.367
R277 B.n260 B.n259 163.367
R278 B.n259 B.n258 163.367
R279 B.n258 B.n49 163.367
R280 B.n254 B.n49 163.367
R281 B.n254 B.n253 163.367
R282 B.n253 B.n252 163.367
R283 B.n252 B.n51 163.367
R284 B.n248 B.n51 163.367
R285 B.n248 B.n247 163.367
R286 B.n247 B.n246 163.367
R287 B.n246 B.n53 163.367
R288 B.n242 B.n53 163.367
R289 B.n242 B.n241 163.367
R290 B.n241 B.n240 163.367
R291 B.n240 B.n55 163.367
R292 B.n236 B.n55 163.367
R293 B.n236 B.n235 163.367
R294 B.n235 B.n234 163.367
R295 B.n234 B.n57 163.367
R296 B.n230 B.n57 163.367
R297 B.n230 B.n229 163.367
R298 B.n229 B.n228 163.367
R299 B.n228 B.n59 163.367
R300 B.n369 B.n368 163.367
R301 B.n368 B.n9 163.367
R302 B.n364 B.n9 163.367
R303 B.n364 B.n363 163.367
R304 B.n363 B.n362 163.367
R305 B.n362 B.n11 163.367
R306 B.n358 B.n11 163.367
R307 B.n358 B.n357 163.367
R308 B.n357 B.n356 163.367
R309 B.n356 B.n13 163.367
R310 B.n352 B.n13 163.367
R311 B.n352 B.n351 163.367
R312 B.n351 B.n350 163.367
R313 B.n350 B.n15 163.367
R314 B.n346 B.n15 163.367
R315 B.n346 B.n345 163.367
R316 B.n345 B.n344 163.367
R317 B.n344 B.n17 163.367
R318 B.n340 B.n17 163.367
R319 B.n340 B.n339 163.367
R320 B.n339 B.n338 163.367
R321 B.n338 B.n19 163.367
R322 B.n334 B.n19 163.367
R323 B.n334 B.n333 163.367
R324 B.n333 B.n332 163.367
R325 B.n332 B.n21 163.367
R326 B.n328 B.n21 163.367
R327 B.n328 B.n327 163.367
R328 B.n327 B.n326 163.367
R329 B.n326 B.n23 163.367
R330 B.n321 B.n23 163.367
R331 B.n321 B.n320 163.367
R332 B.n320 B.n319 163.367
R333 B.n319 B.n27 163.367
R334 B.n315 B.n27 163.367
R335 B.n315 B.n314 163.367
R336 B.n314 B.n313 163.367
R337 B.n313 B.n29 163.367
R338 B.n308 B.n29 163.367
R339 B.n308 B.n307 163.367
R340 B.n307 B.n306 163.367
R341 B.n306 B.n33 163.367
R342 B.n302 B.n33 163.367
R343 B.n302 B.n301 163.367
R344 B.n301 B.n300 163.367
R345 B.n300 B.n35 163.367
R346 B.n296 B.n35 163.367
R347 B.n296 B.n295 163.367
R348 B.n295 B.n294 163.367
R349 B.n294 B.n37 163.367
R350 B.n290 B.n37 163.367
R351 B.n290 B.n289 163.367
R352 B.n289 B.n288 163.367
R353 B.n288 B.n39 163.367
R354 B.n284 B.n39 163.367
R355 B.n284 B.n283 163.367
R356 B.n283 B.n282 163.367
R357 B.n282 B.n41 163.367
R358 B.n278 B.n41 163.367
R359 B.n278 B.n277 163.367
R360 B.n277 B.n276 163.367
R361 B.n276 B.n43 163.367
R362 B.n272 B.n43 163.367
R363 B.n272 B.n271 163.367
R364 B.n271 B.n270 163.367
R365 B.n270 B.n45 163.367
R366 B.n266 B.n45 163.367
R367 B.n266 B.n265 163.367
R368 B.n370 B.n7 163.367
R369 B.n374 B.n7 163.367
R370 B.n375 B.n374 163.367
R371 B.n376 B.n375 163.367
R372 B.n376 B.n5 163.367
R373 B.n380 B.n5 163.367
R374 B.n381 B.n380 163.367
R375 B.n382 B.n381 163.367
R376 B.n382 B.n3 163.367
R377 B.n386 B.n3 163.367
R378 B.n387 B.n386 163.367
R379 B.n101 B.n2 163.367
R380 B.n104 B.n101 163.367
R381 B.n105 B.n104 163.367
R382 B.n106 B.n105 163.367
R383 B.n106 B.n99 163.367
R384 B.n110 B.n99 163.367
R385 B.n111 B.n110 163.367
R386 B.n112 B.n111 163.367
R387 B.n112 B.n97 163.367
R388 B.n116 B.n97 163.367
R389 B.n117 B.n116 163.367
R390 B.n163 B.n81 59.5399
R391 B.n178 B.n177 59.5399
R392 B.n310 B.n31 59.5399
R393 B.n324 B.n25 59.5399
R394 B.n371 B.n8 34.1859
R395 B.n263 B.n46 34.1859
R396 B.n226 B.n225 34.1859
R397 B.n119 B.n96 34.1859
R398 B B.n389 18.0485
R399 B.n81 B.n80 14.546
R400 B.n177 B.n176 14.546
R401 B.n31 B.n30 14.546
R402 B.n25 B.n24 14.546
R403 B.n372 B.n371 10.6151
R404 B.n373 B.n372 10.6151
R405 B.n373 B.n6 10.6151
R406 B.n377 B.n6 10.6151
R407 B.n378 B.n377 10.6151
R408 B.n379 B.n378 10.6151
R409 B.n379 B.n4 10.6151
R410 B.n383 B.n4 10.6151
R411 B.n384 B.n383 10.6151
R412 B.n385 B.n384 10.6151
R413 B.n385 B.n0 10.6151
R414 B.n367 B.n8 10.6151
R415 B.n367 B.n366 10.6151
R416 B.n366 B.n365 10.6151
R417 B.n365 B.n10 10.6151
R418 B.n361 B.n10 10.6151
R419 B.n361 B.n360 10.6151
R420 B.n360 B.n359 10.6151
R421 B.n359 B.n12 10.6151
R422 B.n355 B.n12 10.6151
R423 B.n355 B.n354 10.6151
R424 B.n354 B.n353 10.6151
R425 B.n353 B.n14 10.6151
R426 B.n349 B.n14 10.6151
R427 B.n349 B.n348 10.6151
R428 B.n348 B.n347 10.6151
R429 B.n347 B.n16 10.6151
R430 B.n343 B.n16 10.6151
R431 B.n343 B.n342 10.6151
R432 B.n342 B.n341 10.6151
R433 B.n341 B.n18 10.6151
R434 B.n337 B.n18 10.6151
R435 B.n337 B.n336 10.6151
R436 B.n336 B.n335 10.6151
R437 B.n335 B.n20 10.6151
R438 B.n331 B.n20 10.6151
R439 B.n331 B.n330 10.6151
R440 B.n330 B.n329 10.6151
R441 B.n329 B.n22 10.6151
R442 B.n325 B.n22 10.6151
R443 B.n323 B.n322 10.6151
R444 B.n322 B.n26 10.6151
R445 B.n318 B.n26 10.6151
R446 B.n318 B.n317 10.6151
R447 B.n317 B.n316 10.6151
R448 B.n316 B.n28 10.6151
R449 B.n312 B.n28 10.6151
R450 B.n312 B.n311 10.6151
R451 B.n309 B.n32 10.6151
R452 B.n305 B.n32 10.6151
R453 B.n305 B.n304 10.6151
R454 B.n304 B.n303 10.6151
R455 B.n303 B.n34 10.6151
R456 B.n299 B.n34 10.6151
R457 B.n299 B.n298 10.6151
R458 B.n298 B.n297 10.6151
R459 B.n297 B.n36 10.6151
R460 B.n293 B.n36 10.6151
R461 B.n293 B.n292 10.6151
R462 B.n292 B.n291 10.6151
R463 B.n291 B.n38 10.6151
R464 B.n287 B.n38 10.6151
R465 B.n287 B.n286 10.6151
R466 B.n286 B.n285 10.6151
R467 B.n285 B.n40 10.6151
R468 B.n281 B.n40 10.6151
R469 B.n281 B.n280 10.6151
R470 B.n280 B.n279 10.6151
R471 B.n279 B.n42 10.6151
R472 B.n275 B.n42 10.6151
R473 B.n275 B.n274 10.6151
R474 B.n274 B.n273 10.6151
R475 B.n273 B.n44 10.6151
R476 B.n269 B.n44 10.6151
R477 B.n269 B.n268 10.6151
R478 B.n268 B.n267 10.6151
R479 B.n267 B.n46 10.6151
R480 B.n263 B.n262 10.6151
R481 B.n262 B.n261 10.6151
R482 B.n261 B.n48 10.6151
R483 B.n257 B.n48 10.6151
R484 B.n257 B.n256 10.6151
R485 B.n256 B.n255 10.6151
R486 B.n255 B.n50 10.6151
R487 B.n251 B.n50 10.6151
R488 B.n251 B.n250 10.6151
R489 B.n250 B.n249 10.6151
R490 B.n249 B.n52 10.6151
R491 B.n245 B.n52 10.6151
R492 B.n245 B.n244 10.6151
R493 B.n244 B.n243 10.6151
R494 B.n243 B.n54 10.6151
R495 B.n239 B.n54 10.6151
R496 B.n239 B.n238 10.6151
R497 B.n238 B.n237 10.6151
R498 B.n237 B.n56 10.6151
R499 B.n233 B.n56 10.6151
R500 B.n233 B.n232 10.6151
R501 B.n232 B.n231 10.6151
R502 B.n231 B.n58 10.6151
R503 B.n227 B.n58 10.6151
R504 B.n227 B.n226 10.6151
R505 B.n102 B.n1 10.6151
R506 B.n103 B.n102 10.6151
R507 B.n103 B.n100 10.6151
R508 B.n107 B.n100 10.6151
R509 B.n108 B.n107 10.6151
R510 B.n109 B.n108 10.6151
R511 B.n109 B.n98 10.6151
R512 B.n113 B.n98 10.6151
R513 B.n114 B.n113 10.6151
R514 B.n115 B.n114 10.6151
R515 B.n115 B.n96 10.6151
R516 B.n120 B.n119 10.6151
R517 B.n121 B.n120 10.6151
R518 B.n121 B.n94 10.6151
R519 B.n125 B.n94 10.6151
R520 B.n126 B.n125 10.6151
R521 B.n127 B.n126 10.6151
R522 B.n127 B.n92 10.6151
R523 B.n131 B.n92 10.6151
R524 B.n132 B.n131 10.6151
R525 B.n133 B.n132 10.6151
R526 B.n133 B.n90 10.6151
R527 B.n137 B.n90 10.6151
R528 B.n138 B.n137 10.6151
R529 B.n139 B.n138 10.6151
R530 B.n139 B.n88 10.6151
R531 B.n143 B.n88 10.6151
R532 B.n144 B.n143 10.6151
R533 B.n145 B.n144 10.6151
R534 B.n145 B.n86 10.6151
R535 B.n149 B.n86 10.6151
R536 B.n150 B.n149 10.6151
R537 B.n151 B.n150 10.6151
R538 B.n151 B.n84 10.6151
R539 B.n155 B.n84 10.6151
R540 B.n156 B.n155 10.6151
R541 B.n157 B.n156 10.6151
R542 B.n157 B.n82 10.6151
R543 B.n161 B.n82 10.6151
R544 B.n162 B.n161 10.6151
R545 B.n164 B.n78 10.6151
R546 B.n168 B.n78 10.6151
R547 B.n169 B.n168 10.6151
R548 B.n170 B.n169 10.6151
R549 B.n170 B.n76 10.6151
R550 B.n174 B.n76 10.6151
R551 B.n175 B.n174 10.6151
R552 B.n179 B.n175 10.6151
R553 B.n183 B.n74 10.6151
R554 B.n184 B.n183 10.6151
R555 B.n185 B.n184 10.6151
R556 B.n185 B.n72 10.6151
R557 B.n189 B.n72 10.6151
R558 B.n190 B.n189 10.6151
R559 B.n191 B.n190 10.6151
R560 B.n191 B.n70 10.6151
R561 B.n195 B.n70 10.6151
R562 B.n196 B.n195 10.6151
R563 B.n197 B.n196 10.6151
R564 B.n197 B.n68 10.6151
R565 B.n201 B.n68 10.6151
R566 B.n202 B.n201 10.6151
R567 B.n203 B.n202 10.6151
R568 B.n203 B.n66 10.6151
R569 B.n207 B.n66 10.6151
R570 B.n208 B.n207 10.6151
R571 B.n209 B.n208 10.6151
R572 B.n209 B.n64 10.6151
R573 B.n213 B.n64 10.6151
R574 B.n214 B.n213 10.6151
R575 B.n215 B.n214 10.6151
R576 B.n215 B.n62 10.6151
R577 B.n219 B.n62 10.6151
R578 B.n220 B.n219 10.6151
R579 B.n221 B.n220 10.6151
R580 B.n221 B.n60 10.6151
R581 B.n225 B.n60 10.6151
R582 B.n389 B.n0 8.11757
R583 B.n389 B.n1 8.11757
R584 B.n324 B.n323 7.18099
R585 B.n311 B.n310 7.18099
R586 B.n164 B.n163 7.18099
R587 B.n179 B.n178 7.18099
R588 B.n325 B.n324 3.43465
R589 B.n310 B.n309 3.43465
R590 B.n163 B.n162 3.43465
R591 B.n178 B.n74 3.43465
R592 VP.n0 VP.t1 749.723
R593 VP.n0 VP.t0 713.88
R594 VP VP.n0 0.0516364
R595 VTAIL.n162 VTAIL.n126 756.745
R596 VTAIL.n36 VTAIL.n0 756.745
R597 VTAIL.n120 VTAIL.n84 756.745
R598 VTAIL.n78 VTAIL.n42 756.745
R599 VTAIL.n138 VTAIL.n137 585
R600 VTAIL.n143 VTAIL.n142 585
R601 VTAIL.n145 VTAIL.n144 585
R602 VTAIL.n134 VTAIL.n133 585
R603 VTAIL.n151 VTAIL.n150 585
R604 VTAIL.n153 VTAIL.n152 585
R605 VTAIL.n130 VTAIL.n129 585
R606 VTAIL.n160 VTAIL.n159 585
R607 VTAIL.n161 VTAIL.n128 585
R608 VTAIL.n163 VTAIL.n162 585
R609 VTAIL.n12 VTAIL.n11 585
R610 VTAIL.n17 VTAIL.n16 585
R611 VTAIL.n19 VTAIL.n18 585
R612 VTAIL.n8 VTAIL.n7 585
R613 VTAIL.n25 VTAIL.n24 585
R614 VTAIL.n27 VTAIL.n26 585
R615 VTAIL.n4 VTAIL.n3 585
R616 VTAIL.n34 VTAIL.n33 585
R617 VTAIL.n35 VTAIL.n2 585
R618 VTAIL.n37 VTAIL.n36 585
R619 VTAIL.n121 VTAIL.n120 585
R620 VTAIL.n119 VTAIL.n86 585
R621 VTAIL.n118 VTAIL.n117 585
R622 VTAIL.n89 VTAIL.n87 585
R623 VTAIL.n112 VTAIL.n111 585
R624 VTAIL.n110 VTAIL.n109 585
R625 VTAIL.n93 VTAIL.n92 585
R626 VTAIL.n104 VTAIL.n103 585
R627 VTAIL.n102 VTAIL.n101 585
R628 VTAIL.n97 VTAIL.n96 585
R629 VTAIL.n79 VTAIL.n78 585
R630 VTAIL.n77 VTAIL.n44 585
R631 VTAIL.n76 VTAIL.n75 585
R632 VTAIL.n47 VTAIL.n45 585
R633 VTAIL.n70 VTAIL.n69 585
R634 VTAIL.n68 VTAIL.n67 585
R635 VTAIL.n51 VTAIL.n50 585
R636 VTAIL.n62 VTAIL.n61 585
R637 VTAIL.n60 VTAIL.n59 585
R638 VTAIL.n55 VTAIL.n54 585
R639 VTAIL.n139 VTAIL.t1 329.043
R640 VTAIL.n13 VTAIL.t2 329.043
R641 VTAIL.n98 VTAIL.t3 329.043
R642 VTAIL.n56 VTAIL.t0 329.043
R643 VTAIL.n143 VTAIL.n137 171.744
R644 VTAIL.n144 VTAIL.n143 171.744
R645 VTAIL.n144 VTAIL.n133 171.744
R646 VTAIL.n151 VTAIL.n133 171.744
R647 VTAIL.n152 VTAIL.n151 171.744
R648 VTAIL.n152 VTAIL.n129 171.744
R649 VTAIL.n160 VTAIL.n129 171.744
R650 VTAIL.n161 VTAIL.n160 171.744
R651 VTAIL.n162 VTAIL.n161 171.744
R652 VTAIL.n17 VTAIL.n11 171.744
R653 VTAIL.n18 VTAIL.n17 171.744
R654 VTAIL.n18 VTAIL.n7 171.744
R655 VTAIL.n25 VTAIL.n7 171.744
R656 VTAIL.n26 VTAIL.n25 171.744
R657 VTAIL.n26 VTAIL.n3 171.744
R658 VTAIL.n34 VTAIL.n3 171.744
R659 VTAIL.n35 VTAIL.n34 171.744
R660 VTAIL.n36 VTAIL.n35 171.744
R661 VTAIL.n120 VTAIL.n119 171.744
R662 VTAIL.n119 VTAIL.n118 171.744
R663 VTAIL.n118 VTAIL.n87 171.744
R664 VTAIL.n111 VTAIL.n87 171.744
R665 VTAIL.n111 VTAIL.n110 171.744
R666 VTAIL.n110 VTAIL.n92 171.744
R667 VTAIL.n103 VTAIL.n92 171.744
R668 VTAIL.n103 VTAIL.n102 171.744
R669 VTAIL.n102 VTAIL.n96 171.744
R670 VTAIL.n78 VTAIL.n77 171.744
R671 VTAIL.n77 VTAIL.n76 171.744
R672 VTAIL.n76 VTAIL.n45 171.744
R673 VTAIL.n69 VTAIL.n45 171.744
R674 VTAIL.n69 VTAIL.n68 171.744
R675 VTAIL.n68 VTAIL.n50 171.744
R676 VTAIL.n61 VTAIL.n50 171.744
R677 VTAIL.n61 VTAIL.n60 171.744
R678 VTAIL.n60 VTAIL.n54 171.744
R679 VTAIL.t1 VTAIL.n137 85.8723
R680 VTAIL.t2 VTAIL.n11 85.8723
R681 VTAIL.t3 VTAIL.n96 85.8723
R682 VTAIL.t0 VTAIL.n54 85.8723
R683 VTAIL.n167 VTAIL.n166 35.6763
R684 VTAIL.n41 VTAIL.n40 35.6763
R685 VTAIL.n125 VTAIL.n124 35.6763
R686 VTAIL.n83 VTAIL.n82 35.6763
R687 VTAIL.n83 VTAIL.n41 20.5565
R688 VTAIL.n167 VTAIL.n125 19.91
R689 VTAIL.n163 VTAIL.n128 13.1884
R690 VTAIL.n37 VTAIL.n2 13.1884
R691 VTAIL.n121 VTAIL.n86 13.1884
R692 VTAIL.n79 VTAIL.n44 13.1884
R693 VTAIL.n159 VTAIL.n158 12.8005
R694 VTAIL.n164 VTAIL.n126 12.8005
R695 VTAIL.n33 VTAIL.n32 12.8005
R696 VTAIL.n38 VTAIL.n0 12.8005
R697 VTAIL.n122 VTAIL.n84 12.8005
R698 VTAIL.n117 VTAIL.n88 12.8005
R699 VTAIL.n80 VTAIL.n42 12.8005
R700 VTAIL.n75 VTAIL.n46 12.8005
R701 VTAIL.n157 VTAIL.n130 12.0247
R702 VTAIL.n31 VTAIL.n4 12.0247
R703 VTAIL.n116 VTAIL.n89 12.0247
R704 VTAIL.n74 VTAIL.n47 12.0247
R705 VTAIL.n154 VTAIL.n153 11.249
R706 VTAIL.n28 VTAIL.n27 11.249
R707 VTAIL.n113 VTAIL.n112 11.249
R708 VTAIL.n71 VTAIL.n70 11.249
R709 VTAIL.n139 VTAIL.n138 10.7238
R710 VTAIL.n13 VTAIL.n12 10.7238
R711 VTAIL.n98 VTAIL.n97 10.7238
R712 VTAIL.n56 VTAIL.n55 10.7238
R713 VTAIL.n150 VTAIL.n132 10.4732
R714 VTAIL.n24 VTAIL.n6 10.4732
R715 VTAIL.n109 VTAIL.n91 10.4732
R716 VTAIL.n67 VTAIL.n49 10.4732
R717 VTAIL.n149 VTAIL.n134 9.69747
R718 VTAIL.n23 VTAIL.n8 9.69747
R719 VTAIL.n108 VTAIL.n93 9.69747
R720 VTAIL.n66 VTAIL.n51 9.69747
R721 VTAIL.n166 VTAIL.n165 9.45567
R722 VTAIL.n40 VTAIL.n39 9.45567
R723 VTAIL.n124 VTAIL.n123 9.45567
R724 VTAIL.n82 VTAIL.n81 9.45567
R725 VTAIL.n165 VTAIL.n164 9.3005
R726 VTAIL.n141 VTAIL.n140 9.3005
R727 VTAIL.n136 VTAIL.n135 9.3005
R728 VTAIL.n147 VTAIL.n146 9.3005
R729 VTAIL.n149 VTAIL.n148 9.3005
R730 VTAIL.n132 VTAIL.n131 9.3005
R731 VTAIL.n155 VTAIL.n154 9.3005
R732 VTAIL.n157 VTAIL.n156 9.3005
R733 VTAIL.n158 VTAIL.n127 9.3005
R734 VTAIL.n39 VTAIL.n38 9.3005
R735 VTAIL.n15 VTAIL.n14 9.3005
R736 VTAIL.n10 VTAIL.n9 9.3005
R737 VTAIL.n21 VTAIL.n20 9.3005
R738 VTAIL.n23 VTAIL.n22 9.3005
R739 VTAIL.n6 VTAIL.n5 9.3005
R740 VTAIL.n29 VTAIL.n28 9.3005
R741 VTAIL.n31 VTAIL.n30 9.3005
R742 VTAIL.n32 VTAIL.n1 9.3005
R743 VTAIL.n100 VTAIL.n99 9.3005
R744 VTAIL.n95 VTAIL.n94 9.3005
R745 VTAIL.n106 VTAIL.n105 9.3005
R746 VTAIL.n108 VTAIL.n107 9.3005
R747 VTAIL.n91 VTAIL.n90 9.3005
R748 VTAIL.n114 VTAIL.n113 9.3005
R749 VTAIL.n116 VTAIL.n115 9.3005
R750 VTAIL.n88 VTAIL.n85 9.3005
R751 VTAIL.n123 VTAIL.n122 9.3005
R752 VTAIL.n58 VTAIL.n57 9.3005
R753 VTAIL.n53 VTAIL.n52 9.3005
R754 VTAIL.n64 VTAIL.n63 9.3005
R755 VTAIL.n66 VTAIL.n65 9.3005
R756 VTAIL.n49 VTAIL.n48 9.3005
R757 VTAIL.n72 VTAIL.n71 9.3005
R758 VTAIL.n74 VTAIL.n73 9.3005
R759 VTAIL.n46 VTAIL.n43 9.3005
R760 VTAIL.n81 VTAIL.n80 9.3005
R761 VTAIL.n146 VTAIL.n145 8.92171
R762 VTAIL.n20 VTAIL.n19 8.92171
R763 VTAIL.n105 VTAIL.n104 8.92171
R764 VTAIL.n63 VTAIL.n62 8.92171
R765 VTAIL.n142 VTAIL.n136 8.14595
R766 VTAIL.n16 VTAIL.n10 8.14595
R767 VTAIL.n101 VTAIL.n95 8.14595
R768 VTAIL.n59 VTAIL.n53 8.14595
R769 VTAIL.n141 VTAIL.n138 7.3702
R770 VTAIL.n15 VTAIL.n12 7.3702
R771 VTAIL.n100 VTAIL.n97 7.3702
R772 VTAIL.n58 VTAIL.n55 7.3702
R773 VTAIL.n142 VTAIL.n141 5.81868
R774 VTAIL.n16 VTAIL.n15 5.81868
R775 VTAIL.n101 VTAIL.n100 5.81868
R776 VTAIL.n59 VTAIL.n58 5.81868
R777 VTAIL.n145 VTAIL.n136 5.04292
R778 VTAIL.n19 VTAIL.n10 5.04292
R779 VTAIL.n104 VTAIL.n95 5.04292
R780 VTAIL.n62 VTAIL.n53 5.04292
R781 VTAIL.n146 VTAIL.n134 4.26717
R782 VTAIL.n20 VTAIL.n8 4.26717
R783 VTAIL.n105 VTAIL.n93 4.26717
R784 VTAIL.n63 VTAIL.n51 4.26717
R785 VTAIL.n150 VTAIL.n149 3.49141
R786 VTAIL.n24 VTAIL.n23 3.49141
R787 VTAIL.n109 VTAIL.n108 3.49141
R788 VTAIL.n67 VTAIL.n66 3.49141
R789 VTAIL.n153 VTAIL.n132 2.71565
R790 VTAIL.n27 VTAIL.n6 2.71565
R791 VTAIL.n112 VTAIL.n91 2.71565
R792 VTAIL.n70 VTAIL.n49 2.71565
R793 VTAIL.n140 VTAIL.n139 2.4129
R794 VTAIL.n14 VTAIL.n13 2.4129
R795 VTAIL.n99 VTAIL.n98 2.4129
R796 VTAIL.n57 VTAIL.n56 2.4129
R797 VTAIL.n154 VTAIL.n130 1.93989
R798 VTAIL.n28 VTAIL.n4 1.93989
R799 VTAIL.n113 VTAIL.n89 1.93989
R800 VTAIL.n71 VTAIL.n47 1.93989
R801 VTAIL.n159 VTAIL.n157 1.16414
R802 VTAIL.n166 VTAIL.n126 1.16414
R803 VTAIL.n33 VTAIL.n31 1.16414
R804 VTAIL.n40 VTAIL.n0 1.16414
R805 VTAIL.n124 VTAIL.n84 1.16414
R806 VTAIL.n117 VTAIL.n116 1.16414
R807 VTAIL.n82 VTAIL.n42 1.16414
R808 VTAIL.n75 VTAIL.n74 1.16414
R809 VTAIL.n125 VTAIL.n83 0.793603
R810 VTAIL VTAIL.n41 0.690155
R811 VTAIL.n158 VTAIL.n128 0.388379
R812 VTAIL.n164 VTAIL.n163 0.388379
R813 VTAIL.n32 VTAIL.n2 0.388379
R814 VTAIL.n38 VTAIL.n37 0.388379
R815 VTAIL.n122 VTAIL.n121 0.388379
R816 VTAIL.n88 VTAIL.n86 0.388379
R817 VTAIL.n80 VTAIL.n79 0.388379
R818 VTAIL.n46 VTAIL.n44 0.388379
R819 VTAIL.n140 VTAIL.n135 0.155672
R820 VTAIL.n147 VTAIL.n135 0.155672
R821 VTAIL.n148 VTAIL.n147 0.155672
R822 VTAIL.n148 VTAIL.n131 0.155672
R823 VTAIL.n155 VTAIL.n131 0.155672
R824 VTAIL.n156 VTAIL.n155 0.155672
R825 VTAIL.n156 VTAIL.n127 0.155672
R826 VTAIL.n165 VTAIL.n127 0.155672
R827 VTAIL.n14 VTAIL.n9 0.155672
R828 VTAIL.n21 VTAIL.n9 0.155672
R829 VTAIL.n22 VTAIL.n21 0.155672
R830 VTAIL.n22 VTAIL.n5 0.155672
R831 VTAIL.n29 VTAIL.n5 0.155672
R832 VTAIL.n30 VTAIL.n29 0.155672
R833 VTAIL.n30 VTAIL.n1 0.155672
R834 VTAIL.n39 VTAIL.n1 0.155672
R835 VTAIL.n123 VTAIL.n85 0.155672
R836 VTAIL.n115 VTAIL.n85 0.155672
R837 VTAIL.n115 VTAIL.n114 0.155672
R838 VTAIL.n114 VTAIL.n90 0.155672
R839 VTAIL.n107 VTAIL.n90 0.155672
R840 VTAIL.n107 VTAIL.n106 0.155672
R841 VTAIL.n106 VTAIL.n94 0.155672
R842 VTAIL.n99 VTAIL.n94 0.155672
R843 VTAIL.n81 VTAIL.n43 0.155672
R844 VTAIL.n73 VTAIL.n43 0.155672
R845 VTAIL.n73 VTAIL.n72 0.155672
R846 VTAIL.n72 VTAIL.n48 0.155672
R847 VTAIL.n65 VTAIL.n48 0.155672
R848 VTAIL.n65 VTAIL.n64 0.155672
R849 VTAIL.n64 VTAIL.n52 0.155672
R850 VTAIL.n57 VTAIL.n52 0.155672
R851 VTAIL VTAIL.n167 0.103948
R852 VDD1.n36 VDD1.n0 756.745
R853 VDD1.n77 VDD1.n41 756.745
R854 VDD1.n37 VDD1.n36 585
R855 VDD1.n35 VDD1.n2 585
R856 VDD1.n34 VDD1.n33 585
R857 VDD1.n5 VDD1.n3 585
R858 VDD1.n28 VDD1.n27 585
R859 VDD1.n26 VDD1.n25 585
R860 VDD1.n9 VDD1.n8 585
R861 VDD1.n20 VDD1.n19 585
R862 VDD1.n18 VDD1.n17 585
R863 VDD1.n13 VDD1.n12 585
R864 VDD1.n53 VDD1.n52 585
R865 VDD1.n58 VDD1.n57 585
R866 VDD1.n60 VDD1.n59 585
R867 VDD1.n49 VDD1.n48 585
R868 VDD1.n66 VDD1.n65 585
R869 VDD1.n68 VDD1.n67 585
R870 VDD1.n45 VDD1.n44 585
R871 VDD1.n75 VDD1.n74 585
R872 VDD1.n76 VDD1.n43 585
R873 VDD1.n78 VDD1.n77 585
R874 VDD1.n14 VDD1.t0 329.043
R875 VDD1.n54 VDD1.t1 329.043
R876 VDD1.n36 VDD1.n35 171.744
R877 VDD1.n35 VDD1.n34 171.744
R878 VDD1.n34 VDD1.n3 171.744
R879 VDD1.n27 VDD1.n3 171.744
R880 VDD1.n27 VDD1.n26 171.744
R881 VDD1.n26 VDD1.n8 171.744
R882 VDD1.n19 VDD1.n8 171.744
R883 VDD1.n19 VDD1.n18 171.744
R884 VDD1.n18 VDD1.n12 171.744
R885 VDD1.n58 VDD1.n52 171.744
R886 VDD1.n59 VDD1.n58 171.744
R887 VDD1.n59 VDD1.n48 171.744
R888 VDD1.n66 VDD1.n48 171.744
R889 VDD1.n67 VDD1.n66 171.744
R890 VDD1.n67 VDD1.n44 171.744
R891 VDD1.n75 VDD1.n44 171.744
R892 VDD1.n76 VDD1.n75 171.744
R893 VDD1.n77 VDD1.n76 171.744
R894 VDD1.t0 VDD1.n12 85.8723
R895 VDD1.t1 VDD1.n52 85.8723
R896 VDD1 VDD1.n81 84.8906
R897 VDD1 VDD1.n40 52.5749
R898 VDD1.n37 VDD1.n2 13.1884
R899 VDD1.n78 VDD1.n43 13.1884
R900 VDD1.n38 VDD1.n0 12.8005
R901 VDD1.n33 VDD1.n4 12.8005
R902 VDD1.n74 VDD1.n73 12.8005
R903 VDD1.n79 VDD1.n41 12.8005
R904 VDD1.n32 VDD1.n5 12.0247
R905 VDD1.n72 VDD1.n45 12.0247
R906 VDD1.n29 VDD1.n28 11.249
R907 VDD1.n69 VDD1.n68 11.249
R908 VDD1.n14 VDD1.n13 10.7238
R909 VDD1.n54 VDD1.n53 10.7238
R910 VDD1.n25 VDD1.n7 10.4732
R911 VDD1.n65 VDD1.n47 10.4732
R912 VDD1.n24 VDD1.n9 9.69747
R913 VDD1.n64 VDD1.n49 9.69747
R914 VDD1.n40 VDD1.n39 9.45567
R915 VDD1.n81 VDD1.n80 9.45567
R916 VDD1.n16 VDD1.n15 9.3005
R917 VDD1.n11 VDD1.n10 9.3005
R918 VDD1.n22 VDD1.n21 9.3005
R919 VDD1.n24 VDD1.n23 9.3005
R920 VDD1.n7 VDD1.n6 9.3005
R921 VDD1.n30 VDD1.n29 9.3005
R922 VDD1.n32 VDD1.n31 9.3005
R923 VDD1.n4 VDD1.n1 9.3005
R924 VDD1.n39 VDD1.n38 9.3005
R925 VDD1.n80 VDD1.n79 9.3005
R926 VDD1.n56 VDD1.n55 9.3005
R927 VDD1.n51 VDD1.n50 9.3005
R928 VDD1.n62 VDD1.n61 9.3005
R929 VDD1.n64 VDD1.n63 9.3005
R930 VDD1.n47 VDD1.n46 9.3005
R931 VDD1.n70 VDD1.n69 9.3005
R932 VDD1.n72 VDD1.n71 9.3005
R933 VDD1.n73 VDD1.n42 9.3005
R934 VDD1.n21 VDD1.n20 8.92171
R935 VDD1.n61 VDD1.n60 8.92171
R936 VDD1.n17 VDD1.n11 8.14595
R937 VDD1.n57 VDD1.n51 8.14595
R938 VDD1.n16 VDD1.n13 7.3702
R939 VDD1.n56 VDD1.n53 7.3702
R940 VDD1.n17 VDD1.n16 5.81868
R941 VDD1.n57 VDD1.n56 5.81868
R942 VDD1.n20 VDD1.n11 5.04292
R943 VDD1.n60 VDD1.n51 5.04292
R944 VDD1.n21 VDD1.n9 4.26717
R945 VDD1.n61 VDD1.n49 4.26717
R946 VDD1.n25 VDD1.n24 3.49141
R947 VDD1.n65 VDD1.n64 3.49141
R948 VDD1.n28 VDD1.n7 2.71565
R949 VDD1.n68 VDD1.n47 2.71565
R950 VDD1.n15 VDD1.n14 2.4129
R951 VDD1.n55 VDD1.n54 2.4129
R952 VDD1.n29 VDD1.n5 1.93989
R953 VDD1.n69 VDD1.n45 1.93989
R954 VDD1.n40 VDD1.n0 1.16414
R955 VDD1.n33 VDD1.n32 1.16414
R956 VDD1.n74 VDD1.n72 1.16414
R957 VDD1.n81 VDD1.n41 1.16414
R958 VDD1.n38 VDD1.n37 0.388379
R959 VDD1.n4 VDD1.n2 0.388379
R960 VDD1.n73 VDD1.n43 0.388379
R961 VDD1.n79 VDD1.n78 0.388379
R962 VDD1.n39 VDD1.n1 0.155672
R963 VDD1.n31 VDD1.n1 0.155672
R964 VDD1.n31 VDD1.n30 0.155672
R965 VDD1.n30 VDD1.n6 0.155672
R966 VDD1.n23 VDD1.n6 0.155672
R967 VDD1.n23 VDD1.n22 0.155672
R968 VDD1.n22 VDD1.n10 0.155672
R969 VDD1.n15 VDD1.n10 0.155672
R970 VDD1.n55 VDD1.n50 0.155672
R971 VDD1.n62 VDD1.n50 0.155672
R972 VDD1.n63 VDD1.n62 0.155672
R973 VDD1.n63 VDD1.n46 0.155672
R974 VDD1.n70 VDD1.n46 0.155672
R975 VDD1.n71 VDD1.n70 0.155672
R976 VDD1.n71 VDD1.n42 0.155672
R977 VDD1.n80 VDD1.n42 0.155672
R978 VN VN.t1 750.105
R979 VN VN.t0 713.931
R980 VDD2.n77 VDD2.n41 756.745
R981 VDD2.n36 VDD2.n0 756.745
R982 VDD2.n78 VDD2.n77 585
R983 VDD2.n76 VDD2.n43 585
R984 VDD2.n75 VDD2.n74 585
R985 VDD2.n46 VDD2.n44 585
R986 VDD2.n69 VDD2.n68 585
R987 VDD2.n67 VDD2.n66 585
R988 VDD2.n50 VDD2.n49 585
R989 VDD2.n61 VDD2.n60 585
R990 VDD2.n59 VDD2.n58 585
R991 VDD2.n54 VDD2.n53 585
R992 VDD2.n12 VDD2.n11 585
R993 VDD2.n17 VDD2.n16 585
R994 VDD2.n19 VDD2.n18 585
R995 VDD2.n8 VDD2.n7 585
R996 VDD2.n25 VDD2.n24 585
R997 VDD2.n27 VDD2.n26 585
R998 VDD2.n4 VDD2.n3 585
R999 VDD2.n34 VDD2.n33 585
R1000 VDD2.n35 VDD2.n2 585
R1001 VDD2.n37 VDD2.n36 585
R1002 VDD2.n55 VDD2.t0 329.043
R1003 VDD2.n13 VDD2.t1 329.043
R1004 VDD2.n77 VDD2.n76 171.744
R1005 VDD2.n76 VDD2.n75 171.744
R1006 VDD2.n75 VDD2.n44 171.744
R1007 VDD2.n68 VDD2.n44 171.744
R1008 VDD2.n68 VDD2.n67 171.744
R1009 VDD2.n67 VDD2.n49 171.744
R1010 VDD2.n60 VDD2.n49 171.744
R1011 VDD2.n60 VDD2.n59 171.744
R1012 VDD2.n59 VDD2.n53 171.744
R1013 VDD2.n17 VDD2.n11 171.744
R1014 VDD2.n18 VDD2.n17 171.744
R1015 VDD2.n18 VDD2.n7 171.744
R1016 VDD2.n25 VDD2.n7 171.744
R1017 VDD2.n26 VDD2.n25 171.744
R1018 VDD2.n26 VDD2.n3 171.744
R1019 VDD2.n34 VDD2.n3 171.744
R1020 VDD2.n35 VDD2.n34 171.744
R1021 VDD2.n36 VDD2.n35 171.744
R1022 VDD2.t0 VDD2.n53 85.8723
R1023 VDD2.t1 VDD2.n11 85.8723
R1024 VDD2.n82 VDD2.n40 84.2042
R1025 VDD2.n82 VDD2.n81 52.355
R1026 VDD2.n78 VDD2.n43 13.1884
R1027 VDD2.n37 VDD2.n2 13.1884
R1028 VDD2.n79 VDD2.n41 12.8005
R1029 VDD2.n74 VDD2.n45 12.8005
R1030 VDD2.n33 VDD2.n32 12.8005
R1031 VDD2.n38 VDD2.n0 12.8005
R1032 VDD2.n73 VDD2.n46 12.0247
R1033 VDD2.n31 VDD2.n4 12.0247
R1034 VDD2.n70 VDD2.n69 11.249
R1035 VDD2.n28 VDD2.n27 11.249
R1036 VDD2.n55 VDD2.n54 10.7238
R1037 VDD2.n13 VDD2.n12 10.7238
R1038 VDD2.n66 VDD2.n48 10.4732
R1039 VDD2.n24 VDD2.n6 10.4732
R1040 VDD2.n65 VDD2.n50 9.69747
R1041 VDD2.n23 VDD2.n8 9.69747
R1042 VDD2.n81 VDD2.n80 9.45567
R1043 VDD2.n40 VDD2.n39 9.45567
R1044 VDD2.n57 VDD2.n56 9.3005
R1045 VDD2.n52 VDD2.n51 9.3005
R1046 VDD2.n63 VDD2.n62 9.3005
R1047 VDD2.n65 VDD2.n64 9.3005
R1048 VDD2.n48 VDD2.n47 9.3005
R1049 VDD2.n71 VDD2.n70 9.3005
R1050 VDD2.n73 VDD2.n72 9.3005
R1051 VDD2.n45 VDD2.n42 9.3005
R1052 VDD2.n80 VDD2.n79 9.3005
R1053 VDD2.n39 VDD2.n38 9.3005
R1054 VDD2.n15 VDD2.n14 9.3005
R1055 VDD2.n10 VDD2.n9 9.3005
R1056 VDD2.n21 VDD2.n20 9.3005
R1057 VDD2.n23 VDD2.n22 9.3005
R1058 VDD2.n6 VDD2.n5 9.3005
R1059 VDD2.n29 VDD2.n28 9.3005
R1060 VDD2.n31 VDD2.n30 9.3005
R1061 VDD2.n32 VDD2.n1 9.3005
R1062 VDD2.n62 VDD2.n61 8.92171
R1063 VDD2.n20 VDD2.n19 8.92171
R1064 VDD2.n58 VDD2.n52 8.14595
R1065 VDD2.n16 VDD2.n10 8.14595
R1066 VDD2.n57 VDD2.n54 7.3702
R1067 VDD2.n15 VDD2.n12 7.3702
R1068 VDD2.n58 VDD2.n57 5.81868
R1069 VDD2.n16 VDD2.n15 5.81868
R1070 VDD2.n61 VDD2.n52 5.04292
R1071 VDD2.n19 VDD2.n10 5.04292
R1072 VDD2.n62 VDD2.n50 4.26717
R1073 VDD2.n20 VDD2.n8 4.26717
R1074 VDD2.n66 VDD2.n65 3.49141
R1075 VDD2.n24 VDD2.n23 3.49141
R1076 VDD2.n69 VDD2.n48 2.71565
R1077 VDD2.n27 VDD2.n6 2.71565
R1078 VDD2.n56 VDD2.n55 2.4129
R1079 VDD2.n14 VDD2.n13 2.4129
R1080 VDD2.n70 VDD2.n46 1.93989
R1081 VDD2.n28 VDD2.n4 1.93989
R1082 VDD2.n81 VDD2.n41 1.16414
R1083 VDD2.n74 VDD2.n73 1.16414
R1084 VDD2.n33 VDD2.n31 1.16414
R1085 VDD2.n40 VDD2.n0 1.16414
R1086 VDD2.n79 VDD2.n78 0.388379
R1087 VDD2.n45 VDD2.n43 0.388379
R1088 VDD2.n32 VDD2.n2 0.388379
R1089 VDD2.n38 VDD2.n37 0.388379
R1090 VDD2 VDD2.n82 0.220328
R1091 VDD2.n80 VDD2.n42 0.155672
R1092 VDD2.n72 VDD2.n42 0.155672
R1093 VDD2.n72 VDD2.n71 0.155672
R1094 VDD2.n71 VDD2.n47 0.155672
R1095 VDD2.n64 VDD2.n47 0.155672
R1096 VDD2.n64 VDD2.n63 0.155672
R1097 VDD2.n63 VDD2.n51 0.155672
R1098 VDD2.n56 VDD2.n51 0.155672
R1099 VDD2.n14 VDD2.n9 0.155672
R1100 VDD2.n21 VDD2.n9 0.155672
R1101 VDD2.n22 VDD2.n21 0.155672
R1102 VDD2.n22 VDD2.n5 0.155672
R1103 VDD2.n29 VDD2.n5 0.155672
R1104 VDD2.n30 VDD2.n29 0.155672
R1105 VDD2.n30 VDD2.n1 0.155672
R1106 VDD2.n39 VDD2.n1 0.155672
C0 B VDD2 1.08985f
C1 VP VDD1 1.25643f
C2 VN VDD2 1.16546f
C3 w_n1270_n2568# VDD1 1.24169f
C4 VP B 0.879095f
C5 B w_n1270_n2568# 5.32972f
C6 VDD1 VTAIL 4.62247f
C7 VP VN 3.69259f
C8 B VTAIL 1.85971f
C9 w_n1270_n2568# VN 1.50361f
C10 VP VDD2 0.242373f
C11 VN VTAIL 0.794437f
C12 w_n1270_n2568# VDD2 1.24354f
C13 VTAIL VDD2 4.65584f
C14 B VDD1 1.0772f
C15 VP w_n1270_n2568# 1.66069f
C16 VN VDD1 0.148128f
C17 VP VTAIL 0.808944f
C18 B VN 0.629605f
C19 w_n1270_n2568# VTAIL 2.2901f
C20 VDD1 VDD2 0.435415f
C21 VDD2 VSUBS 0.588078f
C22 VDD1 VSUBS 2.3f
C23 VTAIL VSUBS 0.229674f
C24 VN VSUBS 4.1535f
C25 VP VSUBS 0.877402f
C26 B VSUBS 1.94979f
C27 w_n1270_n2568# VSUBS 40.462196f
C28 VDD2.n0 VSUBS 0.019137f
C29 VDD2.n1 VSUBS 0.017899f
C30 VDD2.n2 VSUBS 0.009901f
C31 VDD2.n3 VSUBS 0.022734f
C32 VDD2.n4 VSUBS 0.010184f
C33 VDD2.n5 VSUBS 0.017899f
C34 VDD2.n6 VSUBS 0.009618f
C35 VDD2.n7 VSUBS 0.022734f
C36 VDD2.n8 VSUBS 0.010184f
C37 VDD2.n9 VSUBS 0.017899f
C38 VDD2.n10 VSUBS 0.009618f
C39 VDD2.n11 VSUBS 0.017051f
C40 VDD2.n12 VSUBS 0.017102f
C41 VDD2.t1 VSUBS 0.048837f
C42 VDD2.n13 VSUBS 0.108509f
C43 VDD2.n14 VSUBS 0.564004f
C44 VDD2.n15 VSUBS 0.009618f
C45 VDD2.n16 VSUBS 0.010184f
C46 VDD2.n17 VSUBS 0.022734f
C47 VDD2.n18 VSUBS 0.022734f
C48 VDD2.n19 VSUBS 0.010184f
C49 VDD2.n20 VSUBS 0.009618f
C50 VDD2.n21 VSUBS 0.017899f
C51 VDD2.n22 VSUBS 0.017899f
C52 VDD2.n23 VSUBS 0.009618f
C53 VDD2.n24 VSUBS 0.010184f
C54 VDD2.n25 VSUBS 0.022734f
C55 VDD2.n26 VSUBS 0.022734f
C56 VDD2.n27 VSUBS 0.010184f
C57 VDD2.n28 VSUBS 0.009618f
C58 VDD2.n29 VSUBS 0.017899f
C59 VDD2.n30 VSUBS 0.017899f
C60 VDD2.n31 VSUBS 0.009618f
C61 VDD2.n32 VSUBS 0.009618f
C62 VDD2.n33 VSUBS 0.010184f
C63 VDD2.n34 VSUBS 0.022734f
C64 VDD2.n35 VSUBS 0.022734f
C65 VDD2.n36 VSUBS 0.053231f
C66 VDD2.n37 VSUBS 0.009901f
C67 VDD2.n38 VSUBS 0.009618f
C68 VDD2.n39 VSUBS 0.045775f
C69 VDD2.n40 VSUBS 0.324707f
C70 VDD2.n41 VSUBS 0.019137f
C71 VDD2.n42 VSUBS 0.017899f
C72 VDD2.n43 VSUBS 0.009901f
C73 VDD2.n44 VSUBS 0.022734f
C74 VDD2.n45 VSUBS 0.009618f
C75 VDD2.n46 VSUBS 0.010184f
C76 VDD2.n47 VSUBS 0.017899f
C77 VDD2.n48 VSUBS 0.009618f
C78 VDD2.n49 VSUBS 0.022734f
C79 VDD2.n50 VSUBS 0.010184f
C80 VDD2.n51 VSUBS 0.017899f
C81 VDD2.n52 VSUBS 0.009618f
C82 VDD2.n53 VSUBS 0.017051f
C83 VDD2.n54 VSUBS 0.017102f
C84 VDD2.t0 VSUBS 0.048837f
C85 VDD2.n55 VSUBS 0.108509f
C86 VDD2.n56 VSUBS 0.564004f
C87 VDD2.n57 VSUBS 0.009618f
C88 VDD2.n58 VSUBS 0.010184f
C89 VDD2.n59 VSUBS 0.022734f
C90 VDD2.n60 VSUBS 0.022734f
C91 VDD2.n61 VSUBS 0.010184f
C92 VDD2.n62 VSUBS 0.009618f
C93 VDD2.n63 VSUBS 0.017899f
C94 VDD2.n64 VSUBS 0.017899f
C95 VDD2.n65 VSUBS 0.009618f
C96 VDD2.n66 VSUBS 0.010184f
C97 VDD2.n67 VSUBS 0.022734f
C98 VDD2.n68 VSUBS 0.022734f
C99 VDD2.n69 VSUBS 0.010184f
C100 VDD2.n70 VSUBS 0.009618f
C101 VDD2.n71 VSUBS 0.017899f
C102 VDD2.n72 VSUBS 0.017899f
C103 VDD2.n73 VSUBS 0.009618f
C104 VDD2.n74 VSUBS 0.010184f
C105 VDD2.n75 VSUBS 0.022734f
C106 VDD2.n76 VSUBS 0.022734f
C107 VDD2.n77 VSUBS 0.053231f
C108 VDD2.n78 VSUBS 0.009901f
C109 VDD2.n79 VSUBS 0.009618f
C110 VDD2.n80 VSUBS 0.045775f
C111 VDD2.n81 VSUBS 0.039147f
C112 VDD2.n82 VSUBS 1.58738f
C113 VN.t0 VSUBS 0.424469f
C114 VN.t1 VSUBS 0.492245f
C115 VDD1.n0 VSUBS 0.018471f
C116 VDD1.n1 VSUBS 0.017275f
C117 VDD1.n2 VSUBS 0.009556f
C118 VDD1.n3 VSUBS 0.021942f
C119 VDD1.n4 VSUBS 0.009283f
C120 VDD1.n5 VSUBS 0.009829f
C121 VDD1.n6 VSUBS 0.017275f
C122 VDD1.n7 VSUBS 0.009283f
C123 VDD1.n8 VSUBS 0.021942f
C124 VDD1.n9 VSUBS 0.009829f
C125 VDD1.n10 VSUBS 0.017275f
C126 VDD1.n11 VSUBS 0.009283f
C127 VDD1.n12 VSUBS 0.016456f
C128 VDD1.n13 VSUBS 0.016506f
C129 VDD1.t0 VSUBS 0.047135f
C130 VDD1.n14 VSUBS 0.104727f
C131 VDD1.n15 VSUBS 0.544347f
C132 VDD1.n16 VSUBS 0.009283f
C133 VDD1.n17 VSUBS 0.009829f
C134 VDD1.n18 VSUBS 0.021942f
C135 VDD1.n19 VSUBS 0.021942f
C136 VDD1.n20 VSUBS 0.009829f
C137 VDD1.n21 VSUBS 0.009283f
C138 VDD1.n22 VSUBS 0.017275f
C139 VDD1.n23 VSUBS 0.017275f
C140 VDD1.n24 VSUBS 0.009283f
C141 VDD1.n25 VSUBS 0.009829f
C142 VDD1.n26 VSUBS 0.021942f
C143 VDD1.n27 VSUBS 0.021942f
C144 VDD1.n28 VSUBS 0.009829f
C145 VDD1.n29 VSUBS 0.009283f
C146 VDD1.n30 VSUBS 0.017275f
C147 VDD1.n31 VSUBS 0.017275f
C148 VDD1.n32 VSUBS 0.009283f
C149 VDD1.n33 VSUBS 0.009829f
C150 VDD1.n34 VSUBS 0.021942f
C151 VDD1.n35 VSUBS 0.021942f
C152 VDD1.n36 VSUBS 0.051376f
C153 VDD1.n37 VSUBS 0.009556f
C154 VDD1.n38 VSUBS 0.009283f
C155 VDD1.n39 VSUBS 0.04418f
C156 VDD1.n40 VSUBS 0.037983f
C157 VDD1.n41 VSUBS 0.018471f
C158 VDD1.n42 VSUBS 0.017275f
C159 VDD1.n43 VSUBS 0.009556f
C160 VDD1.n44 VSUBS 0.021942f
C161 VDD1.n45 VSUBS 0.009829f
C162 VDD1.n46 VSUBS 0.017275f
C163 VDD1.n47 VSUBS 0.009283f
C164 VDD1.n48 VSUBS 0.021942f
C165 VDD1.n49 VSUBS 0.009829f
C166 VDD1.n50 VSUBS 0.017275f
C167 VDD1.n51 VSUBS 0.009283f
C168 VDD1.n52 VSUBS 0.016456f
C169 VDD1.n53 VSUBS 0.016506f
C170 VDD1.t1 VSUBS 0.047135f
C171 VDD1.n54 VSUBS 0.104727f
C172 VDD1.n55 VSUBS 0.544347f
C173 VDD1.n56 VSUBS 0.009283f
C174 VDD1.n57 VSUBS 0.009829f
C175 VDD1.n58 VSUBS 0.021942f
C176 VDD1.n59 VSUBS 0.021942f
C177 VDD1.n60 VSUBS 0.009829f
C178 VDD1.n61 VSUBS 0.009283f
C179 VDD1.n62 VSUBS 0.017275f
C180 VDD1.n63 VSUBS 0.017275f
C181 VDD1.n64 VSUBS 0.009283f
C182 VDD1.n65 VSUBS 0.009829f
C183 VDD1.n66 VSUBS 0.021942f
C184 VDD1.n67 VSUBS 0.021942f
C185 VDD1.n68 VSUBS 0.009829f
C186 VDD1.n69 VSUBS 0.009283f
C187 VDD1.n70 VSUBS 0.017275f
C188 VDD1.n71 VSUBS 0.017275f
C189 VDD1.n72 VSUBS 0.009283f
C190 VDD1.n73 VSUBS 0.009283f
C191 VDD1.n74 VSUBS 0.009829f
C192 VDD1.n75 VSUBS 0.021942f
C193 VDD1.n76 VSUBS 0.021942f
C194 VDD1.n77 VSUBS 0.051376f
C195 VDD1.n78 VSUBS 0.009556f
C196 VDD1.n79 VSUBS 0.009283f
C197 VDD1.n80 VSUBS 0.04418f
C198 VDD1.n81 VSUBS 0.332693f
C199 VTAIL.n0 VSUBS 0.025866f
C200 VTAIL.n1 VSUBS 0.024192f
C201 VTAIL.n2 VSUBS 0.013382f
C202 VTAIL.n3 VSUBS 0.030727f
C203 VTAIL.n4 VSUBS 0.013765f
C204 VTAIL.n5 VSUBS 0.024192f
C205 VTAIL.n6 VSUBS 0.013f
C206 VTAIL.n7 VSUBS 0.030727f
C207 VTAIL.n8 VSUBS 0.013765f
C208 VTAIL.n9 VSUBS 0.024192f
C209 VTAIL.n10 VSUBS 0.013f
C210 VTAIL.n11 VSUBS 0.023045f
C211 VTAIL.n12 VSUBS 0.023114f
C212 VTAIL.t2 VSUBS 0.066007f
C213 VTAIL.n13 VSUBS 0.146657f
C214 VTAIL.n14 VSUBS 0.762291f
C215 VTAIL.n15 VSUBS 0.013f
C216 VTAIL.n16 VSUBS 0.013765f
C217 VTAIL.n17 VSUBS 0.030727f
C218 VTAIL.n18 VSUBS 0.030727f
C219 VTAIL.n19 VSUBS 0.013765f
C220 VTAIL.n20 VSUBS 0.013f
C221 VTAIL.n21 VSUBS 0.024192f
C222 VTAIL.n22 VSUBS 0.024192f
C223 VTAIL.n23 VSUBS 0.013f
C224 VTAIL.n24 VSUBS 0.013765f
C225 VTAIL.n25 VSUBS 0.030727f
C226 VTAIL.n26 VSUBS 0.030727f
C227 VTAIL.n27 VSUBS 0.013765f
C228 VTAIL.n28 VSUBS 0.013f
C229 VTAIL.n29 VSUBS 0.024192f
C230 VTAIL.n30 VSUBS 0.024192f
C231 VTAIL.n31 VSUBS 0.013f
C232 VTAIL.n32 VSUBS 0.013f
C233 VTAIL.n33 VSUBS 0.013765f
C234 VTAIL.n34 VSUBS 0.030727f
C235 VTAIL.n35 VSUBS 0.030727f
C236 VTAIL.n36 VSUBS 0.071946f
C237 VTAIL.n37 VSUBS 0.013382f
C238 VTAIL.n38 VSUBS 0.013f
C239 VTAIL.n39 VSUBS 0.061868f
C240 VTAIL.n40 VSUBS 0.036247f
C241 VTAIL.n41 VSUBS 1.04482f
C242 VTAIL.n42 VSUBS 0.025866f
C243 VTAIL.n43 VSUBS 0.024192f
C244 VTAIL.n44 VSUBS 0.013382f
C245 VTAIL.n45 VSUBS 0.030727f
C246 VTAIL.n46 VSUBS 0.013f
C247 VTAIL.n47 VSUBS 0.013765f
C248 VTAIL.n48 VSUBS 0.024192f
C249 VTAIL.n49 VSUBS 0.013f
C250 VTAIL.n50 VSUBS 0.030727f
C251 VTAIL.n51 VSUBS 0.013765f
C252 VTAIL.n52 VSUBS 0.024192f
C253 VTAIL.n53 VSUBS 0.013f
C254 VTAIL.n54 VSUBS 0.023045f
C255 VTAIL.n55 VSUBS 0.023114f
C256 VTAIL.t0 VSUBS 0.066007f
C257 VTAIL.n56 VSUBS 0.146657f
C258 VTAIL.n57 VSUBS 0.762291f
C259 VTAIL.n58 VSUBS 0.013f
C260 VTAIL.n59 VSUBS 0.013765f
C261 VTAIL.n60 VSUBS 0.030727f
C262 VTAIL.n61 VSUBS 0.030727f
C263 VTAIL.n62 VSUBS 0.013765f
C264 VTAIL.n63 VSUBS 0.013f
C265 VTAIL.n64 VSUBS 0.024192f
C266 VTAIL.n65 VSUBS 0.024192f
C267 VTAIL.n66 VSUBS 0.013f
C268 VTAIL.n67 VSUBS 0.013765f
C269 VTAIL.n68 VSUBS 0.030727f
C270 VTAIL.n69 VSUBS 0.030727f
C271 VTAIL.n70 VSUBS 0.013765f
C272 VTAIL.n71 VSUBS 0.013f
C273 VTAIL.n72 VSUBS 0.024192f
C274 VTAIL.n73 VSUBS 0.024192f
C275 VTAIL.n74 VSUBS 0.013f
C276 VTAIL.n75 VSUBS 0.013765f
C277 VTAIL.n76 VSUBS 0.030727f
C278 VTAIL.n77 VSUBS 0.030727f
C279 VTAIL.n78 VSUBS 0.071946f
C280 VTAIL.n79 VSUBS 0.013382f
C281 VTAIL.n80 VSUBS 0.013f
C282 VTAIL.n81 VSUBS 0.061868f
C283 VTAIL.n82 VSUBS 0.036247f
C284 VTAIL.n83 VSUBS 1.05288f
C285 VTAIL.n84 VSUBS 0.025866f
C286 VTAIL.n85 VSUBS 0.024192f
C287 VTAIL.n86 VSUBS 0.013382f
C288 VTAIL.n87 VSUBS 0.030727f
C289 VTAIL.n88 VSUBS 0.013f
C290 VTAIL.n89 VSUBS 0.013765f
C291 VTAIL.n90 VSUBS 0.024192f
C292 VTAIL.n91 VSUBS 0.013f
C293 VTAIL.n92 VSUBS 0.030727f
C294 VTAIL.n93 VSUBS 0.013765f
C295 VTAIL.n94 VSUBS 0.024192f
C296 VTAIL.n95 VSUBS 0.013f
C297 VTAIL.n96 VSUBS 0.023045f
C298 VTAIL.n97 VSUBS 0.023114f
C299 VTAIL.t3 VSUBS 0.066007f
C300 VTAIL.n98 VSUBS 0.146657f
C301 VTAIL.n99 VSUBS 0.762291f
C302 VTAIL.n100 VSUBS 0.013f
C303 VTAIL.n101 VSUBS 0.013765f
C304 VTAIL.n102 VSUBS 0.030727f
C305 VTAIL.n103 VSUBS 0.030727f
C306 VTAIL.n104 VSUBS 0.013765f
C307 VTAIL.n105 VSUBS 0.013f
C308 VTAIL.n106 VSUBS 0.024192f
C309 VTAIL.n107 VSUBS 0.024192f
C310 VTAIL.n108 VSUBS 0.013f
C311 VTAIL.n109 VSUBS 0.013765f
C312 VTAIL.n110 VSUBS 0.030727f
C313 VTAIL.n111 VSUBS 0.030727f
C314 VTAIL.n112 VSUBS 0.013765f
C315 VTAIL.n113 VSUBS 0.013f
C316 VTAIL.n114 VSUBS 0.024192f
C317 VTAIL.n115 VSUBS 0.024192f
C318 VTAIL.n116 VSUBS 0.013f
C319 VTAIL.n117 VSUBS 0.013765f
C320 VTAIL.n118 VSUBS 0.030727f
C321 VTAIL.n119 VSUBS 0.030727f
C322 VTAIL.n120 VSUBS 0.071946f
C323 VTAIL.n121 VSUBS 0.013382f
C324 VTAIL.n122 VSUBS 0.013f
C325 VTAIL.n123 VSUBS 0.061868f
C326 VTAIL.n124 VSUBS 0.036247f
C327 VTAIL.n125 VSUBS 1.00248f
C328 VTAIL.n126 VSUBS 0.025866f
C329 VTAIL.n127 VSUBS 0.024192f
C330 VTAIL.n128 VSUBS 0.013382f
C331 VTAIL.n129 VSUBS 0.030727f
C332 VTAIL.n130 VSUBS 0.013765f
C333 VTAIL.n131 VSUBS 0.024192f
C334 VTAIL.n132 VSUBS 0.013f
C335 VTAIL.n133 VSUBS 0.030727f
C336 VTAIL.n134 VSUBS 0.013765f
C337 VTAIL.n135 VSUBS 0.024192f
C338 VTAIL.n136 VSUBS 0.013f
C339 VTAIL.n137 VSUBS 0.023045f
C340 VTAIL.n138 VSUBS 0.023114f
C341 VTAIL.t1 VSUBS 0.066007f
C342 VTAIL.n139 VSUBS 0.146657f
C343 VTAIL.n140 VSUBS 0.762291f
C344 VTAIL.n141 VSUBS 0.013f
C345 VTAIL.n142 VSUBS 0.013765f
C346 VTAIL.n143 VSUBS 0.030727f
C347 VTAIL.n144 VSUBS 0.030727f
C348 VTAIL.n145 VSUBS 0.013765f
C349 VTAIL.n146 VSUBS 0.013f
C350 VTAIL.n147 VSUBS 0.024192f
C351 VTAIL.n148 VSUBS 0.024192f
C352 VTAIL.n149 VSUBS 0.013f
C353 VTAIL.n150 VSUBS 0.013765f
C354 VTAIL.n151 VSUBS 0.030727f
C355 VTAIL.n152 VSUBS 0.030727f
C356 VTAIL.n153 VSUBS 0.013765f
C357 VTAIL.n154 VSUBS 0.013f
C358 VTAIL.n155 VSUBS 0.024192f
C359 VTAIL.n156 VSUBS 0.024192f
C360 VTAIL.n157 VSUBS 0.013f
C361 VTAIL.n158 VSUBS 0.013f
C362 VTAIL.n159 VSUBS 0.013765f
C363 VTAIL.n160 VSUBS 0.030727f
C364 VTAIL.n161 VSUBS 0.030727f
C365 VTAIL.n162 VSUBS 0.071946f
C366 VTAIL.n163 VSUBS 0.013382f
C367 VTAIL.n164 VSUBS 0.013f
C368 VTAIL.n165 VSUBS 0.061868f
C369 VTAIL.n166 VSUBS 0.036247f
C370 VTAIL.n167 VSUBS 0.948721f
C371 VP.t1 VSUBS 0.497892f
C372 VP.t0 VSUBS 0.431037f
C373 VP.n0 VSUBS 2.7639f
C374 B.n0 VSUBS 0.005429f
C375 B.n1 VSUBS 0.005429f
C376 B.n2 VSUBS 0.00803f
C377 B.n3 VSUBS 0.006153f
C378 B.n4 VSUBS 0.006153f
C379 B.n5 VSUBS 0.006153f
C380 B.n6 VSUBS 0.006153f
C381 B.n7 VSUBS 0.006153f
C382 B.n8 VSUBS 0.015103f
C383 B.n9 VSUBS 0.006153f
C384 B.n10 VSUBS 0.006153f
C385 B.n11 VSUBS 0.006153f
C386 B.n12 VSUBS 0.006153f
C387 B.n13 VSUBS 0.006153f
C388 B.n14 VSUBS 0.006153f
C389 B.n15 VSUBS 0.006153f
C390 B.n16 VSUBS 0.006153f
C391 B.n17 VSUBS 0.006153f
C392 B.n18 VSUBS 0.006153f
C393 B.n19 VSUBS 0.006153f
C394 B.n20 VSUBS 0.006153f
C395 B.n21 VSUBS 0.006153f
C396 B.n22 VSUBS 0.006153f
C397 B.n23 VSUBS 0.006153f
C398 B.t7 VSUBS 0.110947f
C399 B.t8 VSUBS 0.117878f
C400 B.t6 VSUBS 0.120391f
C401 B.n24 VSUBS 0.182329f
C402 B.n25 VSUBS 0.160218f
C403 B.n26 VSUBS 0.006153f
C404 B.n27 VSUBS 0.006153f
C405 B.n28 VSUBS 0.006153f
C406 B.n29 VSUBS 0.006153f
C407 B.t10 VSUBS 0.110949f
C408 B.t11 VSUBS 0.11788f
C409 B.t9 VSUBS 0.120391f
C410 B.n30 VSUBS 0.182327f
C411 B.n31 VSUBS 0.160216f
C412 B.n32 VSUBS 0.006153f
C413 B.n33 VSUBS 0.006153f
C414 B.n34 VSUBS 0.006153f
C415 B.n35 VSUBS 0.006153f
C416 B.n36 VSUBS 0.006153f
C417 B.n37 VSUBS 0.006153f
C418 B.n38 VSUBS 0.006153f
C419 B.n39 VSUBS 0.006153f
C420 B.n40 VSUBS 0.006153f
C421 B.n41 VSUBS 0.006153f
C422 B.n42 VSUBS 0.006153f
C423 B.n43 VSUBS 0.006153f
C424 B.n44 VSUBS 0.006153f
C425 B.n45 VSUBS 0.006153f
C426 B.n46 VSUBS 0.015103f
C427 B.n47 VSUBS 0.006153f
C428 B.n48 VSUBS 0.006153f
C429 B.n49 VSUBS 0.006153f
C430 B.n50 VSUBS 0.006153f
C431 B.n51 VSUBS 0.006153f
C432 B.n52 VSUBS 0.006153f
C433 B.n53 VSUBS 0.006153f
C434 B.n54 VSUBS 0.006153f
C435 B.n55 VSUBS 0.006153f
C436 B.n56 VSUBS 0.006153f
C437 B.n57 VSUBS 0.006153f
C438 B.n58 VSUBS 0.006153f
C439 B.n59 VSUBS 0.014577f
C440 B.n60 VSUBS 0.006153f
C441 B.n61 VSUBS 0.006153f
C442 B.n62 VSUBS 0.006153f
C443 B.n63 VSUBS 0.006153f
C444 B.n64 VSUBS 0.006153f
C445 B.n65 VSUBS 0.006153f
C446 B.n66 VSUBS 0.006153f
C447 B.n67 VSUBS 0.006153f
C448 B.n68 VSUBS 0.006153f
C449 B.n69 VSUBS 0.006153f
C450 B.n70 VSUBS 0.006153f
C451 B.n71 VSUBS 0.006153f
C452 B.n72 VSUBS 0.006153f
C453 B.n73 VSUBS 0.006153f
C454 B.n74 VSUBS 0.004072f
C455 B.n75 VSUBS 0.006153f
C456 B.n76 VSUBS 0.006153f
C457 B.n77 VSUBS 0.006153f
C458 B.n78 VSUBS 0.006153f
C459 B.n79 VSUBS 0.006153f
C460 B.t2 VSUBS 0.110947f
C461 B.t1 VSUBS 0.117878f
C462 B.t0 VSUBS 0.120391f
C463 B.n80 VSUBS 0.182329f
C464 B.n81 VSUBS 0.160218f
C465 B.n82 VSUBS 0.006153f
C466 B.n83 VSUBS 0.006153f
C467 B.n84 VSUBS 0.006153f
C468 B.n85 VSUBS 0.006153f
C469 B.n86 VSUBS 0.006153f
C470 B.n87 VSUBS 0.006153f
C471 B.n88 VSUBS 0.006153f
C472 B.n89 VSUBS 0.006153f
C473 B.n90 VSUBS 0.006153f
C474 B.n91 VSUBS 0.006153f
C475 B.n92 VSUBS 0.006153f
C476 B.n93 VSUBS 0.006153f
C477 B.n94 VSUBS 0.006153f
C478 B.n95 VSUBS 0.006153f
C479 B.n96 VSUBS 0.014577f
C480 B.n97 VSUBS 0.006153f
C481 B.n98 VSUBS 0.006153f
C482 B.n99 VSUBS 0.006153f
C483 B.n100 VSUBS 0.006153f
C484 B.n101 VSUBS 0.006153f
C485 B.n102 VSUBS 0.006153f
C486 B.n103 VSUBS 0.006153f
C487 B.n104 VSUBS 0.006153f
C488 B.n105 VSUBS 0.006153f
C489 B.n106 VSUBS 0.006153f
C490 B.n107 VSUBS 0.006153f
C491 B.n108 VSUBS 0.006153f
C492 B.n109 VSUBS 0.006153f
C493 B.n110 VSUBS 0.006153f
C494 B.n111 VSUBS 0.006153f
C495 B.n112 VSUBS 0.006153f
C496 B.n113 VSUBS 0.006153f
C497 B.n114 VSUBS 0.006153f
C498 B.n115 VSUBS 0.006153f
C499 B.n116 VSUBS 0.006153f
C500 B.n117 VSUBS 0.014577f
C501 B.n118 VSUBS 0.015103f
C502 B.n119 VSUBS 0.015103f
C503 B.n120 VSUBS 0.006153f
C504 B.n121 VSUBS 0.006153f
C505 B.n122 VSUBS 0.006153f
C506 B.n123 VSUBS 0.006153f
C507 B.n124 VSUBS 0.006153f
C508 B.n125 VSUBS 0.006153f
C509 B.n126 VSUBS 0.006153f
C510 B.n127 VSUBS 0.006153f
C511 B.n128 VSUBS 0.006153f
C512 B.n129 VSUBS 0.006153f
C513 B.n130 VSUBS 0.006153f
C514 B.n131 VSUBS 0.006153f
C515 B.n132 VSUBS 0.006153f
C516 B.n133 VSUBS 0.006153f
C517 B.n134 VSUBS 0.006153f
C518 B.n135 VSUBS 0.006153f
C519 B.n136 VSUBS 0.006153f
C520 B.n137 VSUBS 0.006153f
C521 B.n138 VSUBS 0.006153f
C522 B.n139 VSUBS 0.006153f
C523 B.n140 VSUBS 0.006153f
C524 B.n141 VSUBS 0.006153f
C525 B.n142 VSUBS 0.006153f
C526 B.n143 VSUBS 0.006153f
C527 B.n144 VSUBS 0.006153f
C528 B.n145 VSUBS 0.006153f
C529 B.n146 VSUBS 0.006153f
C530 B.n147 VSUBS 0.006153f
C531 B.n148 VSUBS 0.006153f
C532 B.n149 VSUBS 0.006153f
C533 B.n150 VSUBS 0.006153f
C534 B.n151 VSUBS 0.006153f
C535 B.n152 VSUBS 0.006153f
C536 B.n153 VSUBS 0.006153f
C537 B.n154 VSUBS 0.006153f
C538 B.n155 VSUBS 0.006153f
C539 B.n156 VSUBS 0.006153f
C540 B.n157 VSUBS 0.006153f
C541 B.n158 VSUBS 0.006153f
C542 B.n159 VSUBS 0.006153f
C543 B.n160 VSUBS 0.006153f
C544 B.n161 VSUBS 0.006153f
C545 B.n162 VSUBS 0.004072f
C546 B.n163 VSUBS 0.014256f
C547 B.n164 VSUBS 0.005158f
C548 B.n165 VSUBS 0.006153f
C549 B.n166 VSUBS 0.006153f
C550 B.n167 VSUBS 0.006153f
C551 B.n168 VSUBS 0.006153f
C552 B.n169 VSUBS 0.006153f
C553 B.n170 VSUBS 0.006153f
C554 B.n171 VSUBS 0.006153f
C555 B.n172 VSUBS 0.006153f
C556 B.n173 VSUBS 0.006153f
C557 B.n174 VSUBS 0.006153f
C558 B.n175 VSUBS 0.006153f
C559 B.t5 VSUBS 0.110949f
C560 B.t4 VSUBS 0.11788f
C561 B.t3 VSUBS 0.120391f
C562 B.n176 VSUBS 0.182327f
C563 B.n177 VSUBS 0.160216f
C564 B.n178 VSUBS 0.014256f
C565 B.n179 VSUBS 0.005158f
C566 B.n180 VSUBS 0.006153f
C567 B.n181 VSUBS 0.006153f
C568 B.n182 VSUBS 0.006153f
C569 B.n183 VSUBS 0.006153f
C570 B.n184 VSUBS 0.006153f
C571 B.n185 VSUBS 0.006153f
C572 B.n186 VSUBS 0.006153f
C573 B.n187 VSUBS 0.006153f
C574 B.n188 VSUBS 0.006153f
C575 B.n189 VSUBS 0.006153f
C576 B.n190 VSUBS 0.006153f
C577 B.n191 VSUBS 0.006153f
C578 B.n192 VSUBS 0.006153f
C579 B.n193 VSUBS 0.006153f
C580 B.n194 VSUBS 0.006153f
C581 B.n195 VSUBS 0.006153f
C582 B.n196 VSUBS 0.006153f
C583 B.n197 VSUBS 0.006153f
C584 B.n198 VSUBS 0.006153f
C585 B.n199 VSUBS 0.006153f
C586 B.n200 VSUBS 0.006153f
C587 B.n201 VSUBS 0.006153f
C588 B.n202 VSUBS 0.006153f
C589 B.n203 VSUBS 0.006153f
C590 B.n204 VSUBS 0.006153f
C591 B.n205 VSUBS 0.006153f
C592 B.n206 VSUBS 0.006153f
C593 B.n207 VSUBS 0.006153f
C594 B.n208 VSUBS 0.006153f
C595 B.n209 VSUBS 0.006153f
C596 B.n210 VSUBS 0.006153f
C597 B.n211 VSUBS 0.006153f
C598 B.n212 VSUBS 0.006153f
C599 B.n213 VSUBS 0.006153f
C600 B.n214 VSUBS 0.006153f
C601 B.n215 VSUBS 0.006153f
C602 B.n216 VSUBS 0.006153f
C603 B.n217 VSUBS 0.006153f
C604 B.n218 VSUBS 0.006153f
C605 B.n219 VSUBS 0.006153f
C606 B.n220 VSUBS 0.006153f
C607 B.n221 VSUBS 0.006153f
C608 B.n222 VSUBS 0.006153f
C609 B.n223 VSUBS 0.006153f
C610 B.n224 VSUBS 0.015103f
C611 B.n225 VSUBS 0.014408f
C612 B.n226 VSUBS 0.015272f
C613 B.n227 VSUBS 0.006153f
C614 B.n228 VSUBS 0.006153f
C615 B.n229 VSUBS 0.006153f
C616 B.n230 VSUBS 0.006153f
C617 B.n231 VSUBS 0.006153f
C618 B.n232 VSUBS 0.006153f
C619 B.n233 VSUBS 0.006153f
C620 B.n234 VSUBS 0.006153f
C621 B.n235 VSUBS 0.006153f
C622 B.n236 VSUBS 0.006153f
C623 B.n237 VSUBS 0.006153f
C624 B.n238 VSUBS 0.006153f
C625 B.n239 VSUBS 0.006153f
C626 B.n240 VSUBS 0.006153f
C627 B.n241 VSUBS 0.006153f
C628 B.n242 VSUBS 0.006153f
C629 B.n243 VSUBS 0.006153f
C630 B.n244 VSUBS 0.006153f
C631 B.n245 VSUBS 0.006153f
C632 B.n246 VSUBS 0.006153f
C633 B.n247 VSUBS 0.006153f
C634 B.n248 VSUBS 0.006153f
C635 B.n249 VSUBS 0.006153f
C636 B.n250 VSUBS 0.006153f
C637 B.n251 VSUBS 0.006153f
C638 B.n252 VSUBS 0.006153f
C639 B.n253 VSUBS 0.006153f
C640 B.n254 VSUBS 0.006153f
C641 B.n255 VSUBS 0.006153f
C642 B.n256 VSUBS 0.006153f
C643 B.n257 VSUBS 0.006153f
C644 B.n258 VSUBS 0.006153f
C645 B.n259 VSUBS 0.006153f
C646 B.n260 VSUBS 0.006153f
C647 B.n261 VSUBS 0.006153f
C648 B.n262 VSUBS 0.006153f
C649 B.n263 VSUBS 0.014577f
C650 B.n264 VSUBS 0.014577f
C651 B.n265 VSUBS 0.015103f
C652 B.n266 VSUBS 0.006153f
C653 B.n267 VSUBS 0.006153f
C654 B.n268 VSUBS 0.006153f
C655 B.n269 VSUBS 0.006153f
C656 B.n270 VSUBS 0.006153f
C657 B.n271 VSUBS 0.006153f
C658 B.n272 VSUBS 0.006153f
C659 B.n273 VSUBS 0.006153f
C660 B.n274 VSUBS 0.006153f
C661 B.n275 VSUBS 0.006153f
C662 B.n276 VSUBS 0.006153f
C663 B.n277 VSUBS 0.006153f
C664 B.n278 VSUBS 0.006153f
C665 B.n279 VSUBS 0.006153f
C666 B.n280 VSUBS 0.006153f
C667 B.n281 VSUBS 0.006153f
C668 B.n282 VSUBS 0.006153f
C669 B.n283 VSUBS 0.006153f
C670 B.n284 VSUBS 0.006153f
C671 B.n285 VSUBS 0.006153f
C672 B.n286 VSUBS 0.006153f
C673 B.n287 VSUBS 0.006153f
C674 B.n288 VSUBS 0.006153f
C675 B.n289 VSUBS 0.006153f
C676 B.n290 VSUBS 0.006153f
C677 B.n291 VSUBS 0.006153f
C678 B.n292 VSUBS 0.006153f
C679 B.n293 VSUBS 0.006153f
C680 B.n294 VSUBS 0.006153f
C681 B.n295 VSUBS 0.006153f
C682 B.n296 VSUBS 0.006153f
C683 B.n297 VSUBS 0.006153f
C684 B.n298 VSUBS 0.006153f
C685 B.n299 VSUBS 0.006153f
C686 B.n300 VSUBS 0.006153f
C687 B.n301 VSUBS 0.006153f
C688 B.n302 VSUBS 0.006153f
C689 B.n303 VSUBS 0.006153f
C690 B.n304 VSUBS 0.006153f
C691 B.n305 VSUBS 0.006153f
C692 B.n306 VSUBS 0.006153f
C693 B.n307 VSUBS 0.006153f
C694 B.n308 VSUBS 0.006153f
C695 B.n309 VSUBS 0.004072f
C696 B.n310 VSUBS 0.014256f
C697 B.n311 VSUBS 0.005158f
C698 B.n312 VSUBS 0.006153f
C699 B.n313 VSUBS 0.006153f
C700 B.n314 VSUBS 0.006153f
C701 B.n315 VSUBS 0.006153f
C702 B.n316 VSUBS 0.006153f
C703 B.n317 VSUBS 0.006153f
C704 B.n318 VSUBS 0.006153f
C705 B.n319 VSUBS 0.006153f
C706 B.n320 VSUBS 0.006153f
C707 B.n321 VSUBS 0.006153f
C708 B.n322 VSUBS 0.006153f
C709 B.n323 VSUBS 0.005158f
C710 B.n324 VSUBS 0.014256f
C711 B.n325 VSUBS 0.004072f
C712 B.n326 VSUBS 0.006153f
C713 B.n327 VSUBS 0.006153f
C714 B.n328 VSUBS 0.006153f
C715 B.n329 VSUBS 0.006153f
C716 B.n330 VSUBS 0.006153f
C717 B.n331 VSUBS 0.006153f
C718 B.n332 VSUBS 0.006153f
C719 B.n333 VSUBS 0.006153f
C720 B.n334 VSUBS 0.006153f
C721 B.n335 VSUBS 0.006153f
C722 B.n336 VSUBS 0.006153f
C723 B.n337 VSUBS 0.006153f
C724 B.n338 VSUBS 0.006153f
C725 B.n339 VSUBS 0.006153f
C726 B.n340 VSUBS 0.006153f
C727 B.n341 VSUBS 0.006153f
C728 B.n342 VSUBS 0.006153f
C729 B.n343 VSUBS 0.006153f
C730 B.n344 VSUBS 0.006153f
C731 B.n345 VSUBS 0.006153f
C732 B.n346 VSUBS 0.006153f
C733 B.n347 VSUBS 0.006153f
C734 B.n348 VSUBS 0.006153f
C735 B.n349 VSUBS 0.006153f
C736 B.n350 VSUBS 0.006153f
C737 B.n351 VSUBS 0.006153f
C738 B.n352 VSUBS 0.006153f
C739 B.n353 VSUBS 0.006153f
C740 B.n354 VSUBS 0.006153f
C741 B.n355 VSUBS 0.006153f
C742 B.n356 VSUBS 0.006153f
C743 B.n357 VSUBS 0.006153f
C744 B.n358 VSUBS 0.006153f
C745 B.n359 VSUBS 0.006153f
C746 B.n360 VSUBS 0.006153f
C747 B.n361 VSUBS 0.006153f
C748 B.n362 VSUBS 0.006153f
C749 B.n363 VSUBS 0.006153f
C750 B.n364 VSUBS 0.006153f
C751 B.n365 VSUBS 0.006153f
C752 B.n366 VSUBS 0.006153f
C753 B.n367 VSUBS 0.006153f
C754 B.n368 VSUBS 0.006153f
C755 B.n369 VSUBS 0.015103f
C756 B.n370 VSUBS 0.014577f
C757 B.n371 VSUBS 0.014577f
C758 B.n372 VSUBS 0.006153f
C759 B.n373 VSUBS 0.006153f
C760 B.n374 VSUBS 0.006153f
C761 B.n375 VSUBS 0.006153f
C762 B.n376 VSUBS 0.006153f
C763 B.n377 VSUBS 0.006153f
C764 B.n378 VSUBS 0.006153f
C765 B.n379 VSUBS 0.006153f
C766 B.n380 VSUBS 0.006153f
C767 B.n381 VSUBS 0.006153f
C768 B.n382 VSUBS 0.006153f
C769 B.n383 VSUBS 0.006153f
C770 B.n384 VSUBS 0.006153f
C771 B.n385 VSUBS 0.006153f
C772 B.n386 VSUBS 0.006153f
C773 B.n387 VSUBS 0.00803f
C774 B.n388 VSUBS 0.008554f
C775 B.n389 VSUBS 0.01701f
.ends

