* NGSPICE file created from diff_pair_sample_0339.ext - technology: sky130A

.subckt diff_pair_sample_0339 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3283 pd=12.72 as=0 ps=0 w=5.97 l=3.02
X1 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3283 pd=12.72 as=2.3283 ps=12.72 w=5.97 l=3.02
X2 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3283 pd=12.72 as=0 ps=0 w=5.97 l=3.02
X3 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3283 pd=12.72 as=2.3283 ps=12.72 w=5.97 l=3.02
X4 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3283 pd=12.72 as=2.3283 ps=12.72 w=5.97 l=3.02
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.3283 pd=12.72 as=0 ps=0 w=5.97 l=3.02
X6 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3283 pd=12.72 as=2.3283 ps=12.72 w=5.97 l=3.02
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3283 pd=12.72 as=0 ps=0 w=5.97 l=3.02
R0 B.n522 B.n521 585
R1 B.n523 B.n522 585
R2 B.n198 B.n83 585
R3 B.n197 B.n196 585
R4 B.n195 B.n194 585
R5 B.n193 B.n192 585
R6 B.n191 B.n190 585
R7 B.n189 B.n188 585
R8 B.n187 B.n186 585
R9 B.n185 B.n184 585
R10 B.n183 B.n182 585
R11 B.n181 B.n180 585
R12 B.n179 B.n178 585
R13 B.n177 B.n176 585
R14 B.n175 B.n174 585
R15 B.n173 B.n172 585
R16 B.n171 B.n170 585
R17 B.n169 B.n168 585
R18 B.n167 B.n166 585
R19 B.n165 B.n164 585
R20 B.n163 B.n162 585
R21 B.n161 B.n160 585
R22 B.n159 B.n158 585
R23 B.n157 B.n156 585
R24 B.n155 B.n154 585
R25 B.n152 B.n151 585
R26 B.n150 B.n149 585
R27 B.n148 B.n147 585
R28 B.n146 B.n145 585
R29 B.n144 B.n143 585
R30 B.n142 B.n141 585
R31 B.n140 B.n139 585
R32 B.n138 B.n137 585
R33 B.n136 B.n135 585
R34 B.n134 B.n133 585
R35 B.n132 B.n131 585
R36 B.n130 B.n129 585
R37 B.n128 B.n127 585
R38 B.n126 B.n125 585
R39 B.n124 B.n123 585
R40 B.n122 B.n121 585
R41 B.n120 B.n119 585
R42 B.n118 B.n117 585
R43 B.n116 B.n115 585
R44 B.n114 B.n113 585
R45 B.n112 B.n111 585
R46 B.n110 B.n109 585
R47 B.n108 B.n107 585
R48 B.n106 B.n105 585
R49 B.n104 B.n103 585
R50 B.n102 B.n101 585
R51 B.n100 B.n99 585
R52 B.n98 B.n97 585
R53 B.n96 B.n95 585
R54 B.n94 B.n93 585
R55 B.n92 B.n91 585
R56 B.n90 B.n89 585
R57 B.n53 B.n52 585
R58 B.n520 B.n54 585
R59 B.n524 B.n54 585
R60 B.n519 B.n518 585
R61 B.n518 B.n50 585
R62 B.n517 B.n49 585
R63 B.n530 B.n49 585
R64 B.n516 B.n48 585
R65 B.n531 B.n48 585
R66 B.n515 B.n47 585
R67 B.n532 B.n47 585
R68 B.n514 B.n513 585
R69 B.n513 B.n43 585
R70 B.n512 B.n42 585
R71 B.n538 B.n42 585
R72 B.n511 B.n41 585
R73 B.n539 B.n41 585
R74 B.n510 B.n40 585
R75 B.n540 B.n40 585
R76 B.n509 B.n508 585
R77 B.n508 B.n36 585
R78 B.n507 B.n35 585
R79 B.n546 B.n35 585
R80 B.n506 B.n34 585
R81 B.n547 B.n34 585
R82 B.n505 B.n33 585
R83 B.n548 B.n33 585
R84 B.n504 B.n503 585
R85 B.n503 B.n29 585
R86 B.n502 B.n28 585
R87 B.n554 B.n28 585
R88 B.n501 B.n27 585
R89 B.n555 B.n27 585
R90 B.n500 B.n26 585
R91 B.n556 B.n26 585
R92 B.n499 B.n498 585
R93 B.n498 B.n22 585
R94 B.n497 B.n21 585
R95 B.n562 B.n21 585
R96 B.n496 B.n20 585
R97 B.n563 B.n20 585
R98 B.n495 B.n19 585
R99 B.n564 B.n19 585
R100 B.n494 B.n493 585
R101 B.n493 B.n18 585
R102 B.n492 B.n14 585
R103 B.n570 B.n14 585
R104 B.n491 B.n13 585
R105 B.n571 B.n13 585
R106 B.n490 B.n12 585
R107 B.n572 B.n12 585
R108 B.n489 B.n488 585
R109 B.n488 B.n8 585
R110 B.n487 B.n7 585
R111 B.n578 B.n7 585
R112 B.n486 B.n6 585
R113 B.n579 B.n6 585
R114 B.n485 B.n5 585
R115 B.n580 B.n5 585
R116 B.n484 B.n483 585
R117 B.n483 B.n4 585
R118 B.n482 B.n199 585
R119 B.n482 B.n481 585
R120 B.n472 B.n200 585
R121 B.n201 B.n200 585
R122 B.n474 B.n473 585
R123 B.n475 B.n474 585
R124 B.n471 B.n206 585
R125 B.n206 B.n205 585
R126 B.n470 B.n469 585
R127 B.n469 B.n468 585
R128 B.n208 B.n207 585
R129 B.n461 B.n208 585
R130 B.n460 B.n459 585
R131 B.n462 B.n460 585
R132 B.n458 B.n213 585
R133 B.n213 B.n212 585
R134 B.n457 B.n456 585
R135 B.n456 B.n455 585
R136 B.n215 B.n214 585
R137 B.n216 B.n215 585
R138 B.n448 B.n447 585
R139 B.n449 B.n448 585
R140 B.n446 B.n221 585
R141 B.n221 B.n220 585
R142 B.n445 B.n444 585
R143 B.n444 B.n443 585
R144 B.n223 B.n222 585
R145 B.n224 B.n223 585
R146 B.n436 B.n435 585
R147 B.n437 B.n436 585
R148 B.n434 B.n229 585
R149 B.n229 B.n228 585
R150 B.n433 B.n432 585
R151 B.n432 B.n431 585
R152 B.n231 B.n230 585
R153 B.n232 B.n231 585
R154 B.n424 B.n423 585
R155 B.n425 B.n424 585
R156 B.n422 B.n237 585
R157 B.n237 B.n236 585
R158 B.n421 B.n420 585
R159 B.n420 B.n419 585
R160 B.n239 B.n238 585
R161 B.n240 B.n239 585
R162 B.n412 B.n411 585
R163 B.n413 B.n412 585
R164 B.n410 B.n245 585
R165 B.n245 B.n244 585
R166 B.n409 B.n408 585
R167 B.n408 B.n407 585
R168 B.n247 B.n246 585
R169 B.n248 B.n247 585
R170 B.n400 B.n399 585
R171 B.n401 B.n400 585
R172 B.n251 B.n250 585
R173 B.n287 B.n285 585
R174 B.n288 B.n284 585
R175 B.n288 B.n252 585
R176 B.n291 B.n290 585
R177 B.n292 B.n283 585
R178 B.n294 B.n293 585
R179 B.n296 B.n282 585
R180 B.n299 B.n298 585
R181 B.n300 B.n281 585
R182 B.n302 B.n301 585
R183 B.n304 B.n280 585
R184 B.n307 B.n306 585
R185 B.n308 B.n279 585
R186 B.n310 B.n309 585
R187 B.n312 B.n278 585
R188 B.n315 B.n314 585
R189 B.n316 B.n277 585
R190 B.n318 B.n317 585
R191 B.n320 B.n276 585
R192 B.n323 B.n322 585
R193 B.n324 B.n275 585
R194 B.n326 B.n325 585
R195 B.n328 B.n274 585
R196 B.n331 B.n330 585
R197 B.n333 B.n271 585
R198 B.n335 B.n334 585
R199 B.n337 B.n270 585
R200 B.n340 B.n339 585
R201 B.n341 B.n269 585
R202 B.n343 B.n342 585
R203 B.n345 B.n268 585
R204 B.n348 B.n347 585
R205 B.n349 B.n265 585
R206 B.n352 B.n351 585
R207 B.n354 B.n264 585
R208 B.n357 B.n356 585
R209 B.n358 B.n263 585
R210 B.n360 B.n359 585
R211 B.n362 B.n262 585
R212 B.n365 B.n364 585
R213 B.n366 B.n261 585
R214 B.n368 B.n367 585
R215 B.n370 B.n260 585
R216 B.n373 B.n372 585
R217 B.n374 B.n259 585
R218 B.n376 B.n375 585
R219 B.n378 B.n258 585
R220 B.n381 B.n380 585
R221 B.n382 B.n257 585
R222 B.n384 B.n383 585
R223 B.n386 B.n256 585
R224 B.n389 B.n388 585
R225 B.n390 B.n255 585
R226 B.n392 B.n391 585
R227 B.n394 B.n254 585
R228 B.n397 B.n396 585
R229 B.n398 B.n253 585
R230 B.n403 B.n402 585
R231 B.n402 B.n401 585
R232 B.n404 B.n249 585
R233 B.n249 B.n248 585
R234 B.n406 B.n405 585
R235 B.n407 B.n406 585
R236 B.n243 B.n242 585
R237 B.n244 B.n243 585
R238 B.n415 B.n414 585
R239 B.n414 B.n413 585
R240 B.n416 B.n241 585
R241 B.n241 B.n240 585
R242 B.n418 B.n417 585
R243 B.n419 B.n418 585
R244 B.n235 B.n234 585
R245 B.n236 B.n235 585
R246 B.n427 B.n426 585
R247 B.n426 B.n425 585
R248 B.n428 B.n233 585
R249 B.n233 B.n232 585
R250 B.n430 B.n429 585
R251 B.n431 B.n430 585
R252 B.n227 B.n226 585
R253 B.n228 B.n227 585
R254 B.n439 B.n438 585
R255 B.n438 B.n437 585
R256 B.n440 B.n225 585
R257 B.n225 B.n224 585
R258 B.n442 B.n441 585
R259 B.n443 B.n442 585
R260 B.n219 B.n218 585
R261 B.n220 B.n219 585
R262 B.n451 B.n450 585
R263 B.n450 B.n449 585
R264 B.n452 B.n217 585
R265 B.n217 B.n216 585
R266 B.n454 B.n453 585
R267 B.n455 B.n454 585
R268 B.n211 B.n210 585
R269 B.n212 B.n211 585
R270 B.n464 B.n463 585
R271 B.n463 B.n462 585
R272 B.n465 B.n209 585
R273 B.n461 B.n209 585
R274 B.n467 B.n466 585
R275 B.n468 B.n467 585
R276 B.n204 B.n203 585
R277 B.n205 B.n204 585
R278 B.n477 B.n476 585
R279 B.n476 B.n475 585
R280 B.n478 B.n202 585
R281 B.n202 B.n201 585
R282 B.n480 B.n479 585
R283 B.n481 B.n480 585
R284 B.n2 B.n0 585
R285 B.n4 B.n2 585
R286 B.n3 B.n1 585
R287 B.n579 B.n3 585
R288 B.n577 B.n576 585
R289 B.n578 B.n577 585
R290 B.n575 B.n9 585
R291 B.n9 B.n8 585
R292 B.n574 B.n573 585
R293 B.n573 B.n572 585
R294 B.n11 B.n10 585
R295 B.n571 B.n11 585
R296 B.n569 B.n568 585
R297 B.n570 B.n569 585
R298 B.n567 B.n15 585
R299 B.n18 B.n15 585
R300 B.n566 B.n565 585
R301 B.n565 B.n564 585
R302 B.n17 B.n16 585
R303 B.n563 B.n17 585
R304 B.n561 B.n560 585
R305 B.n562 B.n561 585
R306 B.n559 B.n23 585
R307 B.n23 B.n22 585
R308 B.n558 B.n557 585
R309 B.n557 B.n556 585
R310 B.n25 B.n24 585
R311 B.n555 B.n25 585
R312 B.n553 B.n552 585
R313 B.n554 B.n553 585
R314 B.n551 B.n30 585
R315 B.n30 B.n29 585
R316 B.n550 B.n549 585
R317 B.n549 B.n548 585
R318 B.n32 B.n31 585
R319 B.n547 B.n32 585
R320 B.n545 B.n544 585
R321 B.n546 B.n545 585
R322 B.n543 B.n37 585
R323 B.n37 B.n36 585
R324 B.n542 B.n541 585
R325 B.n541 B.n540 585
R326 B.n39 B.n38 585
R327 B.n539 B.n39 585
R328 B.n537 B.n536 585
R329 B.n538 B.n537 585
R330 B.n535 B.n44 585
R331 B.n44 B.n43 585
R332 B.n534 B.n533 585
R333 B.n533 B.n532 585
R334 B.n46 B.n45 585
R335 B.n531 B.n46 585
R336 B.n529 B.n528 585
R337 B.n530 B.n529 585
R338 B.n527 B.n51 585
R339 B.n51 B.n50 585
R340 B.n526 B.n525 585
R341 B.n525 B.n524 585
R342 B.n582 B.n581 585
R343 B.n581 B.n580 585
R344 B.n402 B.n251 497.305
R345 B.n525 B.n53 497.305
R346 B.n400 B.n253 497.305
R347 B.n522 B.n54 497.305
R348 B.n523 B.n82 256.663
R349 B.n523 B.n81 256.663
R350 B.n523 B.n80 256.663
R351 B.n523 B.n79 256.663
R352 B.n523 B.n78 256.663
R353 B.n523 B.n77 256.663
R354 B.n523 B.n76 256.663
R355 B.n523 B.n75 256.663
R356 B.n523 B.n74 256.663
R357 B.n523 B.n73 256.663
R358 B.n523 B.n72 256.663
R359 B.n523 B.n71 256.663
R360 B.n523 B.n70 256.663
R361 B.n523 B.n69 256.663
R362 B.n523 B.n68 256.663
R363 B.n523 B.n67 256.663
R364 B.n523 B.n66 256.663
R365 B.n523 B.n65 256.663
R366 B.n523 B.n64 256.663
R367 B.n523 B.n63 256.663
R368 B.n523 B.n62 256.663
R369 B.n523 B.n61 256.663
R370 B.n523 B.n60 256.663
R371 B.n523 B.n59 256.663
R372 B.n523 B.n58 256.663
R373 B.n523 B.n57 256.663
R374 B.n523 B.n56 256.663
R375 B.n523 B.n55 256.663
R376 B.n286 B.n252 256.663
R377 B.n289 B.n252 256.663
R378 B.n295 B.n252 256.663
R379 B.n297 B.n252 256.663
R380 B.n303 B.n252 256.663
R381 B.n305 B.n252 256.663
R382 B.n311 B.n252 256.663
R383 B.n313 B.n252 256.663
R384 B.n319 B.n252 256.663
R385 B.n321 B.n252 256.663
R386 B.n327 B.n252 256.663
R387 B.n329 B.n252 256.663
R388 B.n336 B.n252 256.663
R389 B.n338 B.n252 256.663
R390 B.n344 B.n252 256.663
R391 B.n346 B.n252 256.663
R392 B.n353 B.n252 256.663
R393 B.n355 B.n252 256.663
R394 B.n361 B.n252 256.663
R395 B.n363 B.n252 256.663
R396 B.n369 B.n252 256.663
R397 B.n371 B.n252 256.663
R398 B.n377 B.n252 256.663
R399 B.n379 B.n252 256.663
R400 B.n385 B.n252 256.663
R401 B.n387 B.n252 256.663
R402 B.n393 B.n252 256.663
R403 B.n395 B.n252 256.663
R404 B.n266 B.t10 256.245
R405 B.n272 B.t2 256.245
R406 B.n86 B.t6 256.245
R407 B.n84 B.t13 256.245
R408 B.n266 B.t12 243.375
R409 B.n84 B.t14 243.375
R410 B.n272 B.t5 243.375
R411 B.n86 B.t8 243.375
R412 B.n267 B.t11 178.405
R413 B.n85 B.t15 178.405
R414 B.n273 B.t4 178.405
R415 B.n87 B.t9 178.405
R416 B.n402 B.n249 163.367
R417 B.n406 B.n249 163.367
R418 B.n406 B.n243 163.367
R419 B.n414 B.n243 163.367
R420 B.n414 B.n241 163.367
R421 B.n418 B.n241 163.367
R422 B.n418 B.n235 163.367
R423 B.n426 B.n235 163.367
R424 B.n426 B.n233 163.367
R425 B.n430 B.n233 163.367
R426 B.n430 B.n227 163.367
R427 B.n438 B.n227 163.367
R428 B.n438 B.n225 163.367
R429 B.n442 B.n225 163.367
R430 B.n442 B.n219 163.367
R431 B.n450 B.n219 163.367
R432 B.n450 B.n217 163.367
R433 B.n454 B.n217 163.367
R434 B.n454 B.n211 163.367
R435 B.n463 B.n211 163.367
R436 B.n463 B.n209 163.367
R437 B.n467 B.n209 163.367
R438 B.n467 B.n204 163.367
R439 B.n476 B.n204 163.367
R440 B.n476 B.n202 163.367
R441 B.n480 B.n202 163.367
R442 B.n480 B.n2 163.367
R443 B.n581 B.n2 163.367
R444 B.n581 B.n3 163.367
R445 B.n577 B.n3 163.367
R446 B.n577 B.n9 163.367
R447 B.n573 B.n9 163.367
R448 B.n573 B.n11 163.367
R449 B.n569 B.n11 163.367
R450 B.n569 B.n15 163.367
R451 B.n565 B.n15 163.367
R452 B.n565 B.n17 163.367
R453 B.n561 B.n17 163.367
R454 B.n561 B.n23 163.367
R455 B.n557 B.n23 163.367
R456 B.n557 B.n25 163.367
R457 B.n553 B.n25 163.367
R458 B.n553 B.n30 163.367
R459 B.n549 B.n30 163.367
R460 B.n549 B.n32 163.367
R461 B.n545 B.n32 163.367
R462 B.n545 B.n37 163.367
R463 B.n541 B.n37 163.367
R464 B.n541 B.n39 163.367
R465 B.n537 B.n39 163.367
R466 B.n537 B.n44 163.367
R467 B.n533 B.n44 163.367
R468 B.n533 B.n46 163.367
R469 B.n529 B.n46 163.367
R470 B.n529 B.n51 163.367
R471 B.n525 B.n51 163.367
R472 B.n288 B.n287 163.367
R473 B.n290 B.n288 163.367
R474 B.n294 B.n283 163.367
R475 B.n298 B.n296 163.367
R476 B.n302 B.n281 163.367
R477 B.n306 B.n304 163.367
R478 B.n310 B.n279 163.367
R479 B.n314 B.n312 163.367
R480 B.n318 B.n277 163.367
R481 B.n322 B.n320 163.367
R482 B.n326 B.n275 163.367
R483 B.n330 B.n328 163.367
R484 B.n335 B.n271 163.367
R485 B.n339 B.n337 163.367
R486 B.n343 B.n269 163.367
R487 B.n347 B.n345 163.367
R488 B.n352 B.n265 163.367
R489 B.n356 B.n354 163.367
R490 B.n360 B.n263 163.367
R491 B.n364 B.n362 163.367
R492 B.n368 B.n261 163.367
R493 B.n372 B.n370 163.367
R494 B.n376 B.n259 163.367
R495 B.n380 B.n378 163.367
R496 B.n384 B.n257 163.367
R497 B.n388 B.n386 163.367
R498 B.n392 B.n255 163.367
R499 B.n396 B.n394 163.367
R500 B.n400 B.n247 163.367
R501 B.n408 B.n247 163.367
R502 B.n408 B.n245 163.367
R503 B.n412 B.n245 163.367
R504 B.n412 B.n239 163.367
R505 B.n420 B.n239 163.367
R506 B.n420 B.n237 163.367
R507 B.n424 B.n237 163.367
R508 B.n424 B.n231 163.367
R509 B.n432 B.n231 163.367
R510 B.n432 B.n229 163.367
R511 B.n436 B.n229 163.367
R512 B.n436 B.n223 163.367
R513 B.n444 B.n223 163.367
R514 B.n444 B.n221 163.367
R515 B.n448 B.n221 163.367
R516 B.n448 B.n215 163.367
R517 B.n456 B.n215 163.367
R518 B.n456 B.n213 163.367
R519 B.n460 B.n213 163.367
R520 B.n460 B.n208 163.367
R521 B.n469 B.n208 163.367
R522 B.n469 B.n206 163.367
R523 B.n474 B.n206 163.367
R524 B.n474 B.n200 163.367
R525 B.n482 B.n200 163.367
R526 B.n483 B.n482 163.367
R527 B.n483 B.n5 163.367
R528 B.n6 B.n5 163.367
R529 B.n7 B.n6 163.367
R530 B.n488 B.n7 163.367
R531 B.n488 B.n12 163.367
R532 B.n13 B.n12 163.367
R533 B.n14 B.n13 163.367
R534 B.n493 B.n14 163.367
R535 B.n493 B.n19 163.367
R536 B.n20 B.n19 163.367
R537 B.n21 B.n20 163.367
R538 B.n498 B.n21 163.367
R539 B.n498 B.n26 163.367
R540 B.n27 B.n26 163.367
R541 B.n28 B.n27 163.367
R542 B.n503 B.n28 163.367
R543 B.n503 B.n33 163.367
R544 B.n34 B.n33 163.367
R545 B.n35 B.n34 163.367
R546 B.n508 B.n35 163.367
R547 B.n508 B.n40 163.367
R548 B.n41 B.n40 163.367
R549 B.n42 B.n41 163.367
R550 B.n513 B.n42 163.367
R551 B.n513 B.n47 163.367
R552 B.n48 B.n47 163.367
R553 B.n49 B.n48 163.367
R554 B.n518 B.n49 163.367
R555 B.n518 B.n54 163.367
R556 B.n91 B.n90 163.367
R557 B.n95 B.n94 163.367
R558 B.n99 B.n98 163.367
R559 B.n103 B.n102 163.367
R560 B.n107 B.n106 163.367
R561 B.n111 B.n110 163.367
R562 B.n115 B.n114 163.367
R563 B.n119 B.n118 163.367
R564 B.n123 B.n122 163.367
R565 B.n127 B.n126 163.367
R566 B.n131 B.n130 163.367
R567 B.n135 B.n134 163.367
R568 B.n139 B.n138 163.367
R569 B.n143 B.n142 163.367
R570 B.n147 B.n146 163.367
R571 B.n151 B.n150 163.367
R572 B.n156 B.n155 163.367
R573 B.n160 B.n159 163.367
R574 B.n164 B.n163 163.367
R575 B.n168 B.n167 163.367
R576 B.n172 B.n171 163.367
R577 B.n176 B.n175 163.367
R578 B.n180 B.n179 163.367
R579 B.n184 B.n183 163.367
R580 B.n188 B.n187 163.367
R581 B.n192 B.n191 163.367
R582 B.n196 B.n195 163.367
R583 B.n522 B.n83 163.367
R584 B.n401 B.n252 108.582
R585 B.n524 B.n523 108.582
R586 B.n286 B.n251 71.676
R587 B.n290 B.n289 71.676
R588 B.n295 B.n294 71.676
R589 B.n298 B.n297 71.676
R590 B.n303 B.n302 71.676
R591 B.n306 B.n305 71.676
R592 B.n311 B.n310 71.676
R593 B.n314 B.n313 71.676
R594 B.n319 B.n318 71.676
R595 B.n322 B.n321 71.676
R596 B.n327 B.n326 71.676
R597 B.n330 B.n329 71.676
R598 B.n336 B.n335 71.676
R599 B.n339 B.n338 71.676
R600 B.n344 B.n343 71.676
R601 B.n347 B.n346 71.676
R602 B.n353 B.n352 71.676
R603 B.n356 B.n355 71.676
R604 B.n361 B.n360 71.676
R605 B.n364 B.n363 71.676
R606 B.n369 B.n368 71.676
R607 B.n372 B.n371 71.676
R608 B.n377 B.n376 71.676
R609 B.n380 B.n379 71.676
R610 B.n385 B.n384 71.676
R611 B.n388 B.n387 71.676
R612 B.n393 B.n392 71.676
R613 B.n396 B.n395 71.676
R614 B.n55 B.n53 71.676
R615 B.n91 B.n56 71.676
R616 B.n95 B.n57 71.676
R617 B.n99 B.n58 71.676
R618 B.n103 B.n59 71.676
R619 B.n107 B.n60 71.676
R620 B.n111 B.n61 71.676
R621 B.n115 B.n62 71.676
R622 B.n119 B.n63 71.676
R623 B.n123 B.n64 71.676
R624 B.n127 B.n65 71.676
R625 B.n131 B.n66 71.676
R626 B.n135 B.n67 71.676
R627 B.n139 B.n68 71.676
R628 B.n143 B.n69 71.676
R629 B.n147 B.n70 71.676
R630 B.n151 B.n71 71.676
R631 B.n156 B.n72 71.676
R632 B.n160 B.n73 71.676
R633 B.n164 B.n74 71.676
R634 B.n168 B.n75 71.676
R635 B.n172 B.n76 71.676
R636 B.n176 B.n77 71.676
R637 B.n180 B.n78 71.676
R638 B.n184 B.n79 71.676
R639 B.n188 B.n80 71.676
R640 B.n192 B.n81 71.676
R641 B.n196 B.n82 71.676
R642 B.n83 B.n82 71.676
R643 B.n195 B.n81 71.676
R644 B.n191 B.n80 71.676
R645 B.n187 B.n79 71.676
R646 B.n183 B.n78 71.676
R647 B.n179 B.n77 71.676
R648 B.n175 B.n76 71.676
R649 B.n171 B.n75 71.676
R650 B.n167 B.n74 71.676
R651 B.n163 B.n73 71.676
R652 B.n159 B.n72 71.676
R653 B.n155 B.n71 71.676
R654 B.n150 B.n70 71.676
R655 B.n146 B.n69 71.676
R656 B.n142 B.n68 71.676
R657 B.n138 B.n67 71.676
R658 B.n134 B.n66 71.676
R659 B.n130 B.n65 71.676
R660 B.n126 B.n64 71.676
R661 B.n122 B.n63 71.676
R662 B.n118 B.n62 71.676
R663 B.n114 B.n61 71.676
R664 B.n110 B.n60 71.676
R665 B.n106 B.n59 71.676
R666 B.n102 B.n58 71.676
R667 B.n98 B.n57 71.676
R668 B.n94 B.n56 71.676
R669 B.n90 B.n55 71.676
R670 B.n287 B.n286 71.676
R671 B.n289 B.n283 71.676
R672 B.n296 B.n295 71.676
R673 B.n297 B.n281 71.676
R674 B.n304 B.n303 71.676
R675 B.n305 B.n279 71.676
R676 B.n312 B.n311 71.676
R677 B.n313 B.n277 71.676
R678 B.n320 B.n319 71.676
R679 B.n321 B.n275 71.676
R680 B.n328 B.n327 71.676
R681 B.n329 B.n271 71.676
R682 B.n337 B.n336 71.676
R683 B.n338 B.n269 71.676
R684 B.n345 B.n344 71.676
R685 B.n346 B.n265 71.676
R686 B.n354 B.n353 71.676
R687 B.n355 B.n263 71.676
R688 B.n362 B.n361 71.676
R689 B.n363 B.n261 71.676
R690 B.n370 B.n369 71.676
R691 B.n371 B.n259 71.676
R692 B.n378 B.n377 71.676
R693 B.n379 B.n257 71.676
R694 B.n386 B.n385 71.676
R695 B.n387 B.n255 71.676
R696 B.n394 B.n393 71.676
R697 B.n395 B.n253 71.676
R698 B.n401 B.n248 66.519
R699 B.n407 B.n248 66.519
R700 B.n407 B.n244 66.519
R701 B.n413 B.n244 66.519
R702 B.n413 B.n240 66.519
R703 B.n419 B.n240 66.519
R704 B.n419 B.n236 66.519
R705 B.n425 B.n236 66.519
R706 B.n431 B.n232 66.519
R707 B.n431 B.n228 66.519
R708 B.n437 B.n228 66.519
R709 B.n437 B.n224 66.519
R710 B.n443 B.n224 66.519
R711 B.n443 B.n220 66.519
R712 B.n449 B.n220 66.519
R713 B.n449 B.n216 66.519
R714 B.n455 B.n216 66.519
R715 B.n455 B.n212 66.519
R716 B.n462 B.n212 66.519
R717 B.n462 B.n461 66.519
R718 B.n468 B.n205 66.519
R719 B.n475 B.n205 66.519
R720 B.n475 B.n201 66.519
R721 B.n481 B.n201 66.519
R722 B.n481 B.n4 66.519
R723 B.n580 B.n4 66.519
R724 B.n580 B.n579 66.519
R725 B.n579 B.n578 66.519
R726 B.n578 B.n8 66.519
R727 B.n572 B.n8 66.519
R728 B.n572 B.n571 66.519
R729 B.n571 B.n570 66.519
R730 B.n564 B.n18 66.519
R731 B.n564 B.n563 66.519
R732 B.n563 B.n562 66.519
R733 B.n562 B.n22 66.519
R734 B.n556 B.n22 66.519
R735 B.n556 B.n555 66.519
R736 B.n555 B.n554 66.519
R737 B.n554 B.n29 66.519
R738 B.n548 B.n29 66.519
R739 B.n548 B.n547 66.519
R740 B.n547 B.n546 66.519
R741 B.n546 B.n36 66.519
R742 B.n540 B.n539 66.519
R743 B.n539 B.n538 66.519
R744 B.n538 B.n43 66.519
R745 B.n532 B.n43 66.519
R746 B.n532 B.n531 66.519
R747 B.n531 B.n530 66.519
R748 B.n530 B.n50 66.519
R749 B.n524 B.n50 66.519
R750 B.n267 B.n266 64.9702
R751 B.n273 B.n272 64.9702
R752 B.n87 B.n86 64.9702
R753 B.n85 B.n84 64.9702
R754 B.n350 B.n267 59.5399
R755 B.n332 B.n273 59.5399
R756 B.n88 B.n87 59.5399
R757 B.n153 B.n85 59.5399
R758 B.t3 B.n232 39.129
R759 B.t7 B.n36 39.129
R760 B.n468 B.t0 35.2162
R761 B.n570 B.t1 35.2162
R762 B.n526 B.n52 32.3127
R763 B.n521 B.n520 32.3127
R764 B.n399 B.n398 32.3127
R765 B.n403 B.n250 32.3127
R766 B.n461 B.t0 31.3033
R767 B.n18 B.t1 31.3033
R768 B.n425 B.t3 27.3905
R769 B.n540 B.t7 27.3905
R770 B B.n582 18.0485
R771 B.n89 B.n52 10.6151
R772 B.n92 B.n89 10.6151
R773 B.n93 B.n92 10.6151
R774 B.n96 B.n93 10.6151
R775 B.n97 B.n96 10.6151
R776 B.n100 B.n97 10.6151
R777 B.n101 B.n100 10.6151
R778 B.n104 B.n101 10.6151
R779 B.n105 B.n104 10.6151
R780 B.n108 B.n105 10.6151
R781 B.n109 B.n108 10.6151
R782 B.n112 B.n109 10.6151
R783 B.n113 B.n112 10.6151
R784 B.n116 B.n113 10.6151
R785 B.n117 B.n116 10.6151
R786 B.n120 B.n117 10.6151
R787 B.n121 B.n120 10.6151
R788 B.n124 B.n121 10.6151
R789 B.n125 B.n124 10.6151
R790 B.n128 B.n125 10.6151
R791 B.n129 B.n128 10.6151
R792 B.n132 B.n129 10.6151
R793 B.n133 B.n132 10.6151
R794 B.n137 B.n136 10.6151
R795 B.n140 B.n137 10.6151
R796 B.n141 B.n140 10.6151
R797 B.n144 B.n141 10.6151
R798 B.n145 B.n144 10.6151
R799 B.n148 B.n145 10.6151
R800 B.n149 B.n148 10.6151
R801 B.n152 B.n149 10.6151
R802 B.n157 B.n154 10.6151
R803 B.n158 B.n157 10.6151
R804 B.n161 B.n158 10.6151
R805 B.n162 B.n161 10.6151
R806 B.n165 B.n162 10.6151
R807 B.n166 B.n165 10.6151
R808 B.n169 B.n166 10.6151
R809 B.n170 B.n169 10.6151
R810 B.n173 B.n170 10.6151
R811 B.n174 B.n173 10.6151
R812 B.n177 B.n174 10.6151
R813 B.n178 B.n177 10.6151
R814 B.n181 B.n178 10.6151
R815 B.n182 B.n181 10.6151
R816 B.n185 B.n182 10.6151
R817 B.n186 B.n185 10.6151
R818 B.n189 B.n186 10.6151
R819 B.n190 B.n189 10.6151
R820 B.n193 B.n190 10.6151
R821 B.n194 B.n193 10.6151
R822 B.n197 B.n194 10.6151
R823 B.n198 B.n197 10.6151
R824 B.n521 B.n198 10.6151
R825 B.n399 B.n246 10.6151
R826 B.n409 B.n246 10.6151
R827 B.n410 B.n409 10.6151
R828 B.n411 B.n410 10.6151
R829 B.n411 B.n238 10.6151
R830 B.n421 B.n238 10.6151
R831 B.n422 B.n421 10.6151
R832 B.n423 B.n422 10.6151
R833 B.n423 B.n230 10.6151
R834 B.n433 B.n230 10.6151
R835 B.n434 B.n433 10.6151
R836 B.n435 B.n434 10.6151
R837 B.n435 B.n222 10.6151
R838 B.n445 B.n222 10.6151
R839 B.n446 B.n445 10.6151
R840 B.n447 B.n446 10.6151
R841 B.n447 B.n214 10.6151
R842 B.n457 B.n214 10.6151
R843 B.n458 B.n457 10.6151
R844 B.n459 B.n458 10.6151
R845 B.n459 B.n207 10.6151
R846 B.n470 B.n207 10.6151
R847 B.n471 B.n470 10.6151
R848 B.n473 B.n471 10.6151
R849 B.n473 B.n472 10.6151
R850 B.n472 B.n199 10.6151
R851 B.n484 B.n199 10.6151
R852 B.n485 B.n484 10.6151
R853 B.n486 B.n485 10.6151
R854 B.n487 B.n486 10.6151
R855 B.n489 B.n487 10.6151
R856 B.n490 B.n489 10.6151
R857 B.n491 B.n490 10.6151
R858 B.n492 B.n491 10.6151
R859 B.n494 B.n492 10.6151
R860 B.n495 B.n494 10.6151
R861 B.n496 B.n495 10.6151
R862 B.n497 B.n496 10.6151
R863 B.n499 B.n497 10.6151
R864 B.n500 B.n499 10.6151
R865 B.n501 B.n500 10.6151
R866 B.n502 B.n501 10.6151
R867 B.n504 B.n502 10.6151
R868 B.n505 B.n504 10.6151
R869 B.n506 B.n505 10.6151
R870 B.n507 B.n506 10.6151
R871 B.n509 B.n507 10.6151
R872 B.n510 B.n509 10.6151
R873 B.n511 B.n510 10.6151
R874 B.n512 B.n511 10.6151
R875 B.n514 B.n512 10.6151
R876 B.n515 B.n514 10.6151
R877 B.n516 B.n515 10.6151
R878 B.n517 B.n516 10.6151
R879 B.n519 B.n517 10.6151
R880 B.n520 B.n519 10.6151
R881 B.n285 B.n250 10.6151
R882 B.n285 B.n284 10.6151
R883 B.n291 B.n284 10.6151
R884 B.n292 B.n291 10.6151
R885 B.n293 B.n292 10.6151
R886 B.n293 B.n282 10.6151
R887 B.n299 B.n282 10.6151
R888 B.n300 B.n299 10.6151
R889 B.n301 B.n300 10.6151
R890 B.n301 B.n280 10.6151
R891 B.n307 B.n280 10.6151
R892 B.n308 B.n307 10.6151
R893 B.n309 B.n308 10.6151
R894 B.n309 B.n278 10.6151
R895 B.n315 B.n278 10.6151
R896 B.n316 B.n315 10.6151
R897 B.n317 B.n316 10.6151
R898 B.n317 B.n276 10.6151
R899 B.n323 B.n276 10.6151
R900 B.n324 B.n323 10.6151
R901 B.n325 B.n324 10.6151
R902 B.n325 B.n274 10.6151
R903 B.n331 B.n274 10.6151
R904 B.n334 B.n333 10.6151
R905 B.n334 B.n270 10.6151
R906 B.n340 B.n270 10.6151
R907 B.n341 B.n340 10.6151
R908 B.n342 B.n341 10.6151
R909 B.n342 B.n268 10.6151
R910 B.n348 B.n268 10.6151
R911 B.n349 B.n348 10.6151
R912 B.n351 B.n264 10.6151
R913 B.n357 B.n264 10.6151
R914 B.n358 B.n357 10.6151
R915 B.n359 B.n358 10.6151
R916 B.n359 B.n262 10.6151
R917 B.n365 B.n262 10.6151
R918 B.n366 B.n365 10.6151
R919 B.n367 B.n366 10.6151
R920 B.n367 B.n260 10.6151
R921 B.n373 B.n260 10.6151
R922 B.n374 B.n373 10.6151
R923 B.n375 B.n374 10.6151
R924 B.n375 B.n258 10.6151
R925 B.n381 B.n258 10.6151
R926 B.n382 B.n381 10.6151
R927 B.n383 B.n382 10.6151
R928 B.n383 B.n256 10.6151
R929 B.n389 B.n256 10.6151
R930 B.n390 B.n389 10.6151
R931 B.n391 B.n390 10.6151
R932 B.n391 B.n254 10.6151
R933 B.n397 B.n254 10.6151
R934 B.n398 B.n397 10.6151
R935 B.n404 B.n403 10.6151
R936 B.n405 B.n404 10.6151
R937 B.n405 B.n242 10.6151
R938 B.n415 B.n242 10.6151
R939 B.n416 B.n415 10.6151
R940 B.n417 B.n416 10.6151
R941 B.n417 B.n234 10.6151
R942 B.n427 B.n234 10.6151
R943 B.n428 B.n427 10.6151
R944 B.n429 B.n428 10.6151
R945 B.n429 B.n226 10.6151
R946 B.n439 B.n226 10.6151
R947 B.n440 B.n439 10.6151
R948 B.n441 B.n440 10.6151
R949 B.n441 B.n218 10.6151
R950 B.n451 B.n218 10.6151
R951 B.n452 B.n451 10.6151
R952 B.n453 B.n452 10.6151
R953 B.n453 B.n210 10.6151
R954 B.n464 B.n210 10.6151
R955 B.n465 B.n464 10.6151
R956 B.n466 B.n465 10.6151
R957 B.n466 B.n203 10.6151
R958 B.n477 B.n203 10.6151
R959 B.n478 B.n477 10.6151
R960 B.n479 B.n478 10.6151
R961 B.n479 B.n0 10.6151
R962 B.n576 B.n1 10.6151
R963 B.n576 B.n575 10.6151
R964 B.n575 B.n574 10.6151
R965 B.n574 B.n10 10.6151
R966 B.n568 B.n10 10.6151
R967 B.n568 B.n567 10.6151
R968 B.n567 B.n566 10.6151
R969 B.n566 B.n16 10.6151
R970 B.n560 B.n16 10.6151
R971 B.n560 B.n559 10.6151
R972 B.n559 B.n558 10.6151
R973 B.n558 B.n24 10.6151
R974 B.n552 B.n24 10.6151
R975 B.n552 B.n551 10.6151
R976 B.n551 B.n550 10.6151
R977 B.n550 B.n31 10.6151
R978 B.n544 B.n31 10.6151
R979 B.n544 B.n543 10.6151
R980 B.n543 B.n542 10.6151
R981 B.n542 B.n38 10.6151
R982 B.n536 B.n38 10.6151
R983 B.n536 B.n535 10.6151
R984 B.n535 B.n534 10.6151
R985 B.n534 B.n45 10.6151
R986 B.n528 B.n45 10.6151
R987 B.n528 B.n527 10.6151
R988 B.n527 B.n526 10.6151
R989 B.n136 B.n88 6.5566
R990 B.n153 B.n152 6.5566
R991 B.n333 B.n332 6.5566
R992 B.n350 B.n349 6.5566
R993 B.n133 B.n88 4.05904
R994 B.n154 B.n153 4.05904
R995 B.n332 B.n331 4.05904
R996 B.n351 B.n350 4.05904
R997 B.n582 B.n0 2.81026
R998 B.n582 B.n1 2.81026
R999 VN VN.t1 129.941
R1000 VN VN.t0 89.1689
R1001 VTAIL.n122 VTAIL.n96 289.615
R1002 VTAIL.n26 VTAIL.n0 289.615
R1003 VTAIL.n90 VTAIL.n64 289.615
R1004 VTAIL.n58 VTAIL.n32 289.615
R1005 VTAIL.n107 VTAIL.n106 185
R1006 VTAIL.n104 VTAIL.n103 185
R1007 VTAIL.n113 VTAIL.n112 185
R1008 VTAIL.n115 VTAIL.n114 185
R1009 VTAIL.n100 VTAIL.n99 185
R1010 VTAIL.n121 VTAIL.n120 185
R1011 VTAIL.n123 VTAIL.n122 185
R1012 VTAIL.n11 VTAIL.n10 185
R1013 VTAIL.n8 VTAIL.n7 185
R1014 VTAIL.n17 VTAIL.n16 185
R1015 VTAIL.n19 VTAIL.n18 185
R1016 VTAIL.n4 VTAIL.n3 185
R1017 VTAIL.n25 VTAIL.n24 185
R1018 VTAIL.n27 VTAIL.n26 185
R1019 VTAIL.n91 VTAIL.n90 185
R1020 VTAIL.n89 VTAIL.n88 185
R1021 VTAIL.n68 VTAIL.n67 185
R1022 VTAIL.n83 VTAIL.n82 185
R1023 VTAIL.n81 VTAIL.n80 185
R1024 VTAIL.n72 VTAIL.n71 185
R1025 VTAIL.n75 VTAIL.n74 185
R1026 VTAIL.n59 VTAIL.n58 185
R1027 VTAIL.n57 VTAIL.n56 185
R1028 VTAIL.n36 VTAIL.n35 185
R1029 VTAIL.n51 VTAIL.n50 185
R1030 VTAIL.n49 VTAIL.n48 185
R1031 VTAIL.n40 VTAIL.n39 185
R1032 VTAIL.n43 VTAIL.n42 185
R1033 VTAIL.t3 VTAIL.n105 147.661
R1034 VTAIL.t0 VTAIL.n9 147.661
R1035 VTAIL.t1 VTAIL.n73 147.661
R1036 VTAIL.t2 VTAIL.n41 147.661
R1037 VTAIL.n106 VTAIL.n103 104.615
R1038 VTAIL.n113 VTAIL.n103 104.615
R1039 VTAIL.n114 VTAIL.n113 104.615
R1040 VTAIL.n114 VTAIL.n99 104.615
R1041 VTAIL.n121 VTAIL.n99 104.615
R1042 VTAIL.n122 VTAIL.n121 104.615
R1043 VTAIL.n10 VTAIL.n7 104.615
R1044 VTAIL.n17 VTAIL.n7 104.615
R1045 VTAIL.n18 VTAIL.n17 104.615
R1046 VTAIL.n18 VTAIL.n3 104.615
R1047 VTAIL.n25 VTAIL.n3 104.615
R1048 VTAIL.n26 VTAIL.n25 104.615
R1049 VTAIL.n90 VTAIL.n89 104.615
R1050 VTAIL.n89 VTAIL.n67 104.615
R1051 VTAIL.n82 VTAIL.n67 104.615
R1052 VTAIL.n82 VTAIL.n81 104.615
R1053 VTAIL.n81 VTAIL.n71 104.615
R1054 VTAIL.n74 VTAIL.n71 104.615
R1055 VTAIL.n58 VTAIL.n57 104.615
R1056 VTAIL.n57 VTAIL.n35 104.615
R1057 VTAIL.n50 VTAIL.n35 104.615
R1058 VTAIL.n50 VTAIL.n49 104.615
R1059 VTAIL.n49 VTAIL.n39 104.615
R1060 VTAIL.n42 VTAIL.n39 104.615
R1061 VTAIL.n106 VTAIL.t3 52.3082
R1062 VTAIL.n10 VTAIL.t0 52.3082
R1063 VTAIL.n74 VTAIL.t1 52.3082
R1064 VTAIL.n42 VTAIL.t2 52.3082
R1065 VTAIL.n127 VTAIL.n126 31.6035
R1066 VTAIL.n31 VTAIL.n30 31.6035
R1067 VTAIL.n95 VTAIL.n94 31.6035
R1068 VTAIL.n63 VTAIL.n62 31.6035
R1069 VTAIL.n63 VTAIL.n31 23.2893
R1070 VTAIL.n127 VTAIL.n95 20.4014
R1071 VTAIL.n107 VTAIL.n105 15.6674
R1072 VTAIL.n11 VTAIL.n9 15.6674
R1073 VTAIL.n75 VTAIL.n73 15.6674
R1074 VTAIL.n43 VTAIL.n41 15.6674
R1075 VTAIL.n108 VTAIL.n104 12.8005
R1076 VTAIL.n12 VTAIL.n8 12.8005
R1077 VTAIL.n76 VTAIL.n72 12.8005
R1078 VTAIL.n44 VTAIL.n40 12.8005
R1079 VTAIL.n112 VTAIL.n111 12.0247
R1080 VTAIL.n16 VTAIL.n15 12.0247
R1081 VTAIL.n80 VTAIL.n79 12.0247
R1082 VTAIL.n48 VTAIL.n47 12.0247
R1083 VTAIL.n115 VTAIL.n102 11.249
R1084 VTAIL.n19 VTAIL.n6 11.249
R1085 VTAIL.n83 VTAIL.n70 11.249
R1086 VTAIL.n51 VTAIL.n38 11.249
R1087 VTAIL.n116 VTAIL.n100 10.4732
R1088 VTAIL.n20 VTAIL.n4 10.4732
R1089 VTAIL.n84 VTAIL.n68 10.4732
R1090 VTAIL.n52 VTAIL.n36 10.4732
R1091 VTAIL.n120 VTAIL.n119 9.69747
R1092 VTAIL.n24 VTAIL.n23 9.69747
R1093 VTAIL.n88 VTAIL.n87 9.69747
R1094 VTAIL.n56 VTAIL.n55 9.69747
R1095 VTAIL.n126 VTAIL.n125 9.45567
R1096 VTAIL.n30 VTAIL.n29 9.45567
R1097 VTAIL.n94 VTAIL.n93 9.45567
R1098 VTAIL.n62 VTAIL.n61 9.45567
R1099 VTAIL.n125 VTAIL.n124 9.3005
R1100 VTAIL.n98 VTAIL.n97 9.3005
R1101 VTAIL.n119 VTAIL.n118 9.3005
R1102 VTAIL.n117 VTAIL.n116 9.3005
R1103 VTAIL.n102 VTAIL.n101 9.3005
R1104 VTAIL.n111 VTAIL.n110 9.3005
R1105 VTAIL.n109 VTAIL.n108 9.3005
R1106 VTAIL.n29 VTAIL.n28 9.3005
R1107 VTAIL.n2 VTAIL.n1 9.3005
R1108 VTAIL.n23 VTAIL.n22 9.3005
R1109 VTAIL.n21 VTAIL.n20 9.3005
R1110 VTAIL.n6 VTAIL.n5 9.3005
R1111 VTAIL.n15 VTAIL.n14 9.3005
R1112 VTAIL.n13 VTAIL.n12 9.3005
R1113 VTAIL.n93 VTAIL.n92 9.3005
R1114 VTAIL.n66 VTAIL.n65 9.3005
R1115 VTAIL.n87 VTAIL.n86 9.3005
R1116 VTAIL.n85 VTAIL.n84 9.3005
R1117 VTAIL.n70 VTAIL.n69 9.3005
R1118 VTAIL.n79 VTAIL.n78 9.3005
R1119 VTAIL.n77 VTAIL.n76 9.3005
R1120 VTAIL.n61 VTAIL.n60 9.3005
R1121 VTAIL.n34 VTAIL.n33 9.3005
R1122 VTAIL.n55 VTAIL.n54 9.3005
R1123 VTAIL.n53 VTAIL.n52 9.3005
R1124 VTAIL.n38 VTAIL.n37 9.3005
R1125 VTAIL.n47 VTAIL.n46 9.3005
R1126 VTAIL.n45 VTAIL.n44 9.3005
R1127 VTAIL.n123 VTAIL.n98 8.92171
R1128 VTAIL.n27 VTAIL.n2 8.92171
R1129 VTAIL.n91 VTAIL.n66 8.92171
R1130 VTAIL.n59 VTAIL.n34 8.92171
R1131 VTAIL.n124 VTAIL.n96 8.14595
R1132 VTAIL.n28 VTAIL.n0 8.14595
R1133 VTAIL.n92 VTAIL.n64 8.14595
R1134 VTAIL.n60 VTAIL.n32 8.14595
R1135 VTAIL.n126 VTAIL.n96 5.81868
R1136 VTAIL.n30 VTAIL.n0 5.81868
R1137 VTAIL.n94 VTAIL.n64 5.81868
R1138 VTAIL.n62 VTAIL.n32 5.81868
R1139 VTAIL.n124 VTAIL.n123 5.04292
R1140 VTAIL.n28 VTAIL.n27 5.04292
R1141 VTAIL.n92 VTAIL.n91 5.04292
R1142 VTAIL.n60 VTAIL.n59 5.04292
R1143 VTAIL.n109 VTAIL.n105 4.38594
R1144 VTAIL.n13 VTAIL.n9 4.38594
R1145 VTAIL.n77 VTAIL.n73 4.38594
R1146 VTAIL.n45 VTAIL.n41 4.38594
R1147 VTAIL.n120 VTAIL.n98 4.26717
R1148 VTAIL.n24 VTAIL.n2 4.26717
R1149 VTAIL.n88 VTAIL.n66 4.26717
R1150 VTAIL.n56 VTAIL.n34 4.26717
R1151 VTAIL.n119 VTAIL.n100 3.49141
R1152 VTAIL.n23 VTAIL.n4 3.49141
R1153 VTAIL.n87 VTAIL.n68 3.49141
R1154 VTAIL.n55 VTAIL.n36 3.49141
R1155 VTAIL.n116 VTAIL.n115 2.71565
R1156 VTAIL.n20 VTAIL.n19 2.71565
R1157 VTAIL.n84 VTAIL.n83 2.71565
R1158 VTAIL.n52 VTAIL.n51 2.71565
R1159 VTAIL.n112 VTAIL.n102 1.93989
R1160 VTAIL.n16 VTAIL.n6 1.93989
R1161 VTAIL.n80 VTAIL.n70 1.93989
R1162 VTAIL.n48 VTAIL.n38 1.93989
R1163 VTAIL.n95 VTAIL.n63 1.91429
R1164 VTAIL VTAIL.n31 1.2505
R1165 VTAIL.n111 VTAIL.n104 1.16414
R1166 VTAIL.n15 VTAIL.n8 1.16414
R1167 VTAIL.n79 VTAIL.n72 1.16414
R1168 VTAIL.n47 VTAIL.n40 1.16414
R1169 VTAIL VTAIL.n127 0.664293
R1170 VTAIL.n108 VTAIL.n107 0.388379
R1171 VTAIL.n12 VTAIL.n11 0.388379
R1172 VTAIL.n76 VTAIL.n75 0.388379
R1173 VTAIL.n44 VTAIL.n43 0.388379
R1174 VTAIL.n110 VTAIL.n109 0.155672
R1175 VTAIL.n110 VTAIL.n101 0.155672
R1176 VTAIL.n117 VTAIL.n101 0.155672
R1177 VTAIL.n118 VTAIL.n117 0.155672
R1178 VTAIL.n118 VTAIL.n97 0.155672
R1179 VTAIL.n125 VTAIL.n97 0.155672
R1180 VTAIL.n14 VTAIL.n13 0.155672
R1181 VTAIL.n14 VTAIL.n5 0.155672
R1182 VTAIL.n21 VTAIL.n5 0.155672
R1183 VTAIL.n22 VTAIL.n21 0.155672
R1184 VTAIL.n22 VTAIL.n1 0.155672
R1185 VTAIL.n29 VTAIL.n1 0.155672
R1186 VTAIL.n93 VTAIL.n65 0.155672
R1187 VTAIL.n86 VTAIL.n65 0.155672
R1188 VTAIL.n86 VTAIL.n85 0.155672
R1189 VTAIL.n85 VTAIL.n69 0.155672
R1190 VTAIL.n78 VTAIL.n69 0.155672
R1191 VTAIL.n78 VTAIL.n77 0.155672
R1192 VTAIL.n61 VTAIL.n33 0.155672
R1193 VTAIL.n54 VTAIL.n33 0.155672
R1194 VTAIL.n54 VTAIL.n53 0.155672
R1195 VTAIL.n53 VTAIL.n37 0.155672
R1196 VTAIL.n46 VTAIL.n37 0.155672
R1197 VTAIL.n46 VTAIL.n45 0.155672
R1198 VDD2.n57 VDD2.n31 289.615
R1199 VDD2.n26 VDD2.n0 289.615
R1200 VDD2.n58 VDD2.n57 185
R1201 VDD2.n56 VDD2.n55 185
R1202 VDD2.n35 VDD2.n34 185
R1203 VDD2.n50 VDD2.n49 185
R1204 VDD2.n48 VDD2.n47 185
R1205 VDD2.n39 VDD2.n38 185
R1206 VDD2.n42 VDD2.n41 185
R1207 VDD2.n11 VDD2.n10 185
R1208 VDD2.n8 VDD2.n7 185
R1209 VDD2.n17 VDD2.n16 185
R1210 VDD2.n19 VDD2.n18 185
R1211 VDD2.n4 VDD2.n3 185
R1212 VDD2.n25 VDD2.n24 185
R1213 VDD2.n27 VDD2.n26 185
R1214 VDD2.t0 VDD2.n40 147.661
R1215 VDD2.t1 VDD2.n9 147.661
R1216 VDD2.n57 VDD2.n56 104.615
R1217 VDD2.n56 VDD2.n34 104.615
R1218 VDD2.n49 VDD2.n34 104.615
R1219 VDD2.n49 VDD2.n48 104.615
R1220 VDD2.n48 VDD2.n38 104.615
R1221 VDD2.n41 VDD2.n38 104.615
R1222 VDD2.n10 VDD2.n7 104.615
R1223 VDD2.n17 VDD2.n7 104.615
R1224 VDD2.n18 VDD2.n17 104.615
R1225 VDD2.n18 VDD2.n3 104.615
R1226 VDD2.n25 VDD2.n3 104.615
R1227 VDD2.n26 VDD2.n25 104.615
R1228 VDD2.n62 VDD2.n30 82.8642
R1229 VDD2.n41 VDD2.t0 52.3082
R1230 VDD2.n10 VDD2.t1 52.3082
R1231 VDD2.n62 VDD2.n61 48.2823
R1232 VDD2.n42 VDD2.n40 15.6674
R1233 VDD2.n11 VDD2.n9 15.6674
R1234 VDD2.n43 VDD2.n39 12.8005
R1235 VDD2.n12 VDD2.n8 12.8005
R1236 VDD2.n47 VDD2.n46 12.0247
R1237 VDD2.n16 VDD2.n15 12.0247
R1238 VDD2.n50 VDD2.n37 11.249
R1239 VDD2.n19 VDD2.n6 11.249
R1240 VDD2.n51 VDD2.n35 10.4732
R1241 VDD2.n20 VDD2.n4 10.4732
R1242 VDD2.n55 VDD2.n54 9.69747
R1243 VDD2.n24 VDD2.n23 9.69747
R1244 VDD2.n61 VDD2.n60 9.45567
R1245 VDD2.n30 VDD2.n29 9.45567
R1246 VDD2.n60 VDD2.n59 9.3005
R1247 VDD2.n33 VDD2.n32 9.3005
R1248 VDD2.n54 VDD2.n53 9.3005
R1249 VDD2.n52 VDD2.n51 9.3005
R1250 VDD2.n37 VDD2.n36 9.3005
R1251 VDD2.n46 VDD2.n45 9.3005
R1252 VDD2.n44 VDD2.n43 9.3005
R1253 VDD2.n29 VDD2.n28 9.3005
R1254 VDD2.n2 VDD2.n1 9.3005
R1255 VDD2.n23 VDD2.n22 9.3005
R1256 VDD2.n21 VDD2.n20 9.3005
R1257 VDD2.n6 VDD2.n5 9.3005
R1258 VDD2.n15 VDD2.n14 9.3005
R1259 VDD2.n13 VDD2.n12 9.3005
R1260 VDD2.n58 VDD2.n33 8.92171
R1261 VDD2.n27 VDD2.n2 8.92171
R1262 VDD2.n59 VDD2.n31 8.14595
R1263 VDD2.n28 VDD2.n0 8.14595
R1264 VDD2.n61 VDD2.n31 5.81868
R1265 VDD2.n30 VDD2.n0 5.81868
R1266 VDD2.n59 VDD2.n58 5.04292
R1267 VDD2.n28 VDD2.n27 5.04292
R1268 VDD2.n44 VDD2.n40 4.38594
R1269 VDD2.n13 VDD2.n9 4.38594
R1270 VDD2.n55 VDD2.n33 4.26717
R1271 VDD2.n24 VDD2.n2 4.26717
R1272 VDD2.n54 VDD2.n35 3.49141
R1273 VDD2.n23 VDD2.n4 3.49141
R1274 VDD2.n51 VDD2.n50 2.71565
R1275 VDD2.n20 VDD2.n19 2.71565
R1276 VDD2.n47 VDD2.n37 1.93989
R1277 VDD2.n16 VDD2.n6 1.93989
R1278 VDD2.n46 VDD2.n39 1.16414
R1279 VDD2.n15 VDD2.n8 1.16414
R1280 VDD2 VDD2.n62 0.780672
R1281 VDD2.n43 VDD2.n42 0.388379
R1282 VDD2.n12 VDD2.n11 0.388379
R1283 VDD2.n60 VDD2.n32 0.155672
R1284 VDD2.n53 VDD2.n32 0.155672
R1285 VDD2.n53 VDD2.n52 0.155672
R1286 VDD2.n52 VDD2.n36 0.155672
R1287 VDD2.n45 VDD2.n36 0.155672
R1288 VDD2.n45 VDD2.n44 0.155672
R1289 VDD2.n14 VDD2.n13 0.155672
R1290 VDD2.n14 VDD2.n5 0.155672
R1291 VDD2.n21 VDD2.n5 0.155672
R1292 VDD2.n22 VDD2.n21 0.155672
R1293 VDD2.n22 VDD2.n1 0.155672
R1294 VDD2.n29 VDD2.n1 0.155672
R1295 VP.n0 VP.t0 129.94
R1296 VP.n0 VP.t1 88.7376
R1297 VP VP.n0 0.431811
R1298 VDD1.n26 VDD1.n0 289.615
R1299 VDD1.n57 VDD1.n31 289.615
R1300 VDD1.n27 VDD1.n26 185
R1301 VDD1.n25 VDD1.n24 185
R1302 VDD1.n4 VDD1.n3 185
R1303 VDD1.n19 VDD1.n18 185
R1304 VDD1.n17 VDD1.n16 185
R1305 VDD1.n8 VDD1.n7 185
R1306 VDD1.n11 VDD1.n10 185
R1307 VDD1.n42 VDD1.n41 185
R1308 VDD1.n39 VDD1.n38 185
R1309 VDD1.n48 VDD1.n47 185
R1310 VDD1.n50 VDD1.n49 185
R1311 VDD1.n35 VDD1.n34 185
R1312 VDD1.n56 VDD1.n55 185
R1313 VDD1.n58 VDD1.n57 185
R1314 VDD1.t1 VDD1.n9 147.661
R1315 VDD1.t0 VDD1.n40 147.661
R1316 VDD1.n26 VDD1.n25 104.615
R1317 VDD1.n25 VDD1.n3 104.615
R1318 VDD1.n18 VDD1.n3 104.615
R1319 VDD1.n18 VDD1.n17 104.615
R1320 VDD1.n17 VDD1.n7 104.615
R1321 VDD1.n10 VDD1.n7 104.615
R1322 VDD1.n41 VDD1.n38 104.615
R1323 VDD1.n48 VDD1.n38 104.615
R1324 VDD1.n49 VDD1.n48 104.615
R1325 VDD1.n49 VDD1.n34 104.615
R1326 VDD1.n56 VDD1.n34 104.615
R1327 VDD1.n57 VDD1.n56 104.615
R1328 VDD1 VDD1.n61 84.111
R1329 VDD1.n10 VDD1.t1 52.3082
R1330 VDD1.n41 VDD1.t0 52.3082
R1331 VDD1 VDD1.n30 49.0625
R1332 VDD1.n11 VDD1.n9 15.6674
R1333 VDD1.n42 VDD1.n40 15.6674
R1334 VDD1.n12 VDD1.n8 12.8005
R1335 VDD1.n43 VDD1.n39 12.8005
R1336 VDD1.n16 VDD1.n15 12.0247
R1337 VDD1.n47 VDD1.n46 12.0247
R1338 VDD1.n19 VDD1.n6 11.249
R1339 VDD1.n50 VDD1.n37 11.249
R1340 VDD1.n20 VDD1.n4 10.4732
R1341 VDD1.n51 VDD1.n35 10.4732
R1342 VDD1.n24 VDD1.n23 9.69747
R1343 VDD1.n55 VDD1.n54 9.69747
R1344 VDD1.n30 VDD1.n29 9.45567
R1345 VDD1.n61 VDD1.n60 9.45567
R1346 VDD1.n29 VDD1.n28 9.3005
R1347 VDD1.n2 VDD1.n1 9.3005
R1348 VDD1.n23 VDD1.n22 9.3005
R1349 VDD1.n21 VDD1.n20 9.3005
R1350 VDD1.n6 VDD1.n5 9.3005
R1351 VDD1.n15 VDD1.n14 9.3005
R1352 VDD1.n13 VDD1.n12 9.3005
R1353 VDD1.n60 VDD1.n59 9.3005
R1354 VDD1.n33 VDD1.n32 9.3005
R1355 VDD1.n54 VDD1.n53 9.3005
R1356 VDD1.n52 VDD1.n51 9.3005
R1357 VDD1.n37 VDD1.n36 9.3005
R1358 VDD1.n46 VDD1.n45 9.3005
R1359 VDD1.n44 VDD1.n43 9.3005
R1360 VDD1.n27 VDD1.n2 8.92171
R1361 VDD1.n58 VDD1.n33 8.92171
R1362 VDD1.n28 VDD1.n0 8.14595
R1363 VDD1.n59 VDD1.n31 8.14595
R1364 VDD1.n30 VDD1.n0 5.81868
R1365 VDD1.n61 VDD1.n31 5.81868
R1366 VDD1.n28 VDD1.n27 5.04292
R1367 VDD1.n59 VDD1.n58 5.04292
R1368 VDD1.n13 VDD1.n9 4.38594
R1369 VDD1.n44 VDD1.n40 4.38594
R1370 VDD1.n24 VDD1.n2 4.26717
R1371 VDD1.n55 VDD1.n33 4.26717
R1372 VDD1.n23 VDD1.n4 3.49141
R1373 VDD1.n54 VDD1.n35 3.49141
R1374 VDD1.n20 VDD1.n19 2.71565
R1375 VDD1.n51 VDD1.n50 2.71565
R1376 VDD1.n16 VDD1.n6 1.93989
R1377 VDD1.n47 VDD1.n37 1.93989
R1378 VDD1.n15 VDD1.n8 1.16414
R1379 VDD1.n46 VDD1.n39 1.16414
R1380 VDD1.n12 VDD1.n11 0.388379
R1381 VDD1.n43 VDD1.n42 0.388379
R1382 VDD1.n29 VDD1.n1 0.155672
R1383 VDD1.n22 VDD1.n1 0.155672
R1384 VDD1.n22 VDD1.n21 0.155672
R1385 VDD1.n21 VDD1.n5 0.155672
R1386 VDD1.n14 VDD1.n5 0.155672
R1387 VDD1.n14 VDD1.n13 0.155672
R1388 VDD1.n45 VDD1.n44 0.155672
R1389 VDD1.n45 VDD1.n36 0.155672
R1390 VDD1.n52 VDD1.n36 0.155672
R1391 VDD1.n53 VDD1.n52 0.155672
R1392 VDD1.n53 VDD1.n32 0.155672
R1393 VDD1.n60 VDD1.n32 0.155672
C0 VDD2 VTAIL 3.63855f
C1 VN VDD2 1.54311f
C2 VP VDD2 0.350277f
C3 VTAIL VDD1 3.58351f
C4 VN VDD1 0.148315f
C5 VP VDD1 1.74366f
C6 VN VTAIL 1.61208f
C7 VP VTAIL 1.62626f
C8 VDD2 VDD1 0.724981f
C9 VP VN 4.53424f
C10 VDD2 B 3.449193f
C11 VDD1 B 5.1338f
C12 VTAIL B 4.854207f
C13 VN B 8.34511f
C14 VP B 6.363067f
C15 VDD1.n0 B 0.020061f
C16 VDD1.n1 B 0.014481f
C17 VDD1.n2 B 0.007781f
C18 VDD1.n3 B 0.018392f
C19 VDD1.n4 B 0.008239f
C20 VDD1.n5 B 0.014481f
C21 VDD1.n6 B 0.007781f
C22 VDD1.n7 B 0.018392f
C23 VDD1.n8 B 0.008239f
C24 VDD1.n9 B 0.061847f
C25 VDD1.t1 B 0.02997f
C26 VDD1.n10 B 0.013794f
C27 VDD1.n11 B 0.010864f
C28 VDD1.n12 B 0.007781f
C29 VDD1.n13 B 0.342584f
C30 VDD1.n14 B 0.014481f
C31 VDD1.n15 B 0.007781f
C32 VDD1.n16 B 0.008239f
C33 VDD1.n17 B 0.018392f
C34 VDD1.n18 B 0.018392f
C35 VDD1.n19 B 0.008239f
C36 VDD1.n20 B 0.007781f
C37 VDD1.n21 B 0.014481f
C38 VDD1.n22 B 0.014481f
C39 VDD1.n23 B 0.007781f
C40 VDD1.n24 B 0.008239f
C41 VDD1.n25 B 0.018392f
C42 VDD1.n26 B 0.039298f
C43 VDD1.n27 B 0.008239f
C44 VDD1.n28 B 0.007781f
C45 VDD1.n29 B 0.032878f
C46 VDD1.n30 B 0.032938f
C47 VDD1.n31 B 0.020061f
C48 VDD1.n32 B 0.014481f
C49 VDD1.n33 B 0.007781f
C50 VDD1.n34 B 0.018392f
C51 VDD1.n35 B 0.008239f
C52 VDD1.n36 B 0.014481f
C53 VDD1.n37 B 0.007781f
C54 VDD1.n38 B 0.018392f
C55 VDD1.n39 B 0.008239f
C56 VDD1.n40 B 0.061847f
C57 VDD1.t0 B 0.02997f
C58 VDD1.n41 B 0.013794f
C59 VDD1.n42 B 0.010864f
C60 VDD1.n43 B 0.007781f
C61 VDD1.n44 B 0.342584f
C62 VDD1.n45 B 0.014481f
C63 VDD1.n46 B 0.007781f
C64 VDD1.n47 B 0.008239f
C65 VDD1.n48 B 0.018392f
C66 VDD1.n49 B 0.018392f
C67 VDD1.n50 B 0.008239f
C68 VDD1.n51 B 0.007781f
C69 VDD1.n52 B 0.014481f
C70 VDD1.n53 B 0.014481f
C71 VDD1.n54 B 0.007781f
C72 VDD1.n55 B 0.008239f
C73 VDD1.n56 B 0.018392f
C74 VDD1.n57 B 0.039298f
C75 VDD1.n58 B 0.008239f
C76 VDD1.n59 B 0.007781f
C77 VDD1.n60 B 0.032878f
C78 VDD1.n61 B 0.352573f
C79 VP.t1 B 1.12207f
C80 VP.t0 B 1.47712f
C81 VP.n0 B 1.84416f
C82 VDD2.n0 B 0.020364f
C83 VDD2.n1 B 0.014699f
C84 VDD2.n2 B 0.007899f
C85 VDD2.n3 B 0.01867f
C86 VDD2.n4 B 0.008363f
C87 VDD2.n5 B 0.014699f
C88 VDD2.n6 B 0.007899f
C89 VDD2.n7 B 0.01867f
C90 VDD2.n8 B 0.008363f
C91 VDD2.n9 B 0.06278f
C92 VDD2.t1 B 0.030422f
C93 VDD2.n10 B 0.014002f
C94 VDD2.n11 B 0.011028f
C95 VDD2.n12 B 0.007899f
C96 VDD2.n13 B 0.347751f
C97 VDD2.n14 B 0.014699f
C98 VDD2.n15 B 0.007899f
C99 VDD2.n16 B 0.008363f
C100 VDD2.n17 B 0.01867f
C101 VDD2.n18 B 0.01867f
C102 VDD2.n19 B 0.008363f
C103 VDD2.n20 B 0.007899f
C104 VDD2.n21 B 0.014699f
C105 VDD2.n22 B 0.014699f
C106 VDD2.n23 B 0.007899f
C107 VDD2.n24 B 0.008363f
C108 VDD2.n25 B 0.01867f
C109 VDD2.n26 B 0.039891f
C110 VDD2.n27 B 0.008363f
C111 VDD2.n28 B 0.007899f
C112 VDD2.n29 B 0.033374f
C113 VDD2.n30 B 0.330205f
C114 VDD2.n31 B 0.020364f
C115 VDD2.n32 B 0.014699f
C116 VDD2.n33 B 0.007899f
C117 VDD2.n34 B 0.01867f
C118 VDD2.n35 B 0.008363f
C119 VDD2.n36 B 0.014699f
C120 VDD2.n37 B 0.007899f
C121 VDD2.n38 B 0.01867f
C122 VDD2.n39 B 0.008363f
C123 VDD2.n40 B 0.06278f
C124 VDD2.t0 B 0.030422f
C125 VDD2.n41 B 0.014002f
C126 VDD2.n42 B 0.011028f
C127 VDD2.n43 B 0.007899f
C128 VDD2.n44 B 0.347751f
C129 VDD2.n45 B 0.014699f
C130 VDD2.n46 B 0.007899f
C131 VDD2.n47 B 0.008363f
C132 VDD2.n48 B 0.01867f
C133 VDD2.n49 B 0.01867f
C134 VDD2.n50 B 0.008363f
C135 VDD2.n51 B 0.007899f
C136 VDD2.n52 B 0.014699f
C137 VDD2.n53 B 0.014699f
C138 VDD2.n54 B 0.007899f
C139 VDD2.n55 B 0.008363f
C140 VDD2.n56 B 0.01867f
C141 VDD2.n57 B 0.039891f
C142 VDD2.n58 B 0.008363f
C143 VDD2.n59 B 0.007899f
C144 VDD2.n60 B 0.033374f
C145 VDD2.n61 B 0.032402f
C146 VDD2.n62 B 1.46778f
C147 VTAIL.n0 B 0.022828f
C148 VTAIL.n1 B 0.016478f
C149 VTAIL.n2 B 0.008855f
C150 VTAIL.n3 B 0.02093f
C151 VTAIL.n4 B 0.009376f
C152 VTAIL.n5 B 0.016478f
C153 VTAIL.n6 B 0.008855f
C154 VTAIL.n7 B 0.02093f
C155 VTAIL.n8 B 0.009376f
C156 VTAIL.n9 B 0.070379f
C157 VTAIL.t0 B 0.034104f
C158 VTAIL.n10 B 0.015697f
C159 VTAIL.n11 B 0.012363f
C160 VTAIL.n12 B 0.008855f
C161 VTAIL.n13 B 0.389844f
C162 VTAIL.n14 B 0.016478f
C163 VTAIL.n15 B 0.008855f
C164 VTAIL.n16 B 0.009376f
C165 VTAIL.n17 B 0.02093f
C166 VTAIL.n18 B 0.02093f
C167 VTAIL.n19 B 0.009376f
C168 VTAIL.n20 B 0.008855f
C169 VTAIL.n21 B 0.016478f
C170 VTAIL.n22 B 0.016478f
C171 VTAIL.n23 B 0.008855f
C172 VTAIL.n24 B 0.009376f
C173 VTAIL.n25 B 0.02093f
C174 VTAIL.n26 B 0.044719f
C175 VTAIL.n27 B 0.009376f
C176 VTAIL.n28 B 0.008855f
C177 VTAIL.n29 B 0.037414f
C178 VTAIL.n30 B 0.024941f
C179 VTAIL.n31 B 0.883857f
C180 VTAIL.n32 B 0.022828f
C181 VTAIL.n33 B 0.016478f
C182 VTAIL.n34 B 0.008855f
C183 VTAIL.n35 B 0.02093f
C184 VTAIL.n36 B 0.009376f
C185 VTAIL.n37 B 0.016478f
C186 VTAIL.n38 B 0.008855f
C187 VTAIL.n39 B 0.02093f
C188 VTAIL.n40 B 0.009376f
C189 VTAIL.n41 B 0.070379f
C190 VTAIL.t2 B 0.034104f
C191 VTAIL.n42 B 0.015697f
C192 VTAIL.n43 B 0.012363f
C193 VTAIL.n44 B 0.008855f
C194 VTAIL.n45 B 0.389844f
C195 VTAIL.n46 B 0.016478f
C196 VTAIL.n47 B 0.008855f
C197 VTAIL.n48 B 0.009376f
C198 VTAIL.n49 B 0.02093f
C199 VTAIL.n50 B 0.02093f
C200 VTAIL.n51 B 0.009376f
C201 VTAIL.n52 B 0.008855f
C202 VTAIL.n53 B 0.016478f
C203 VTAIL.n54 B 0.016478f
C204 VTAIL.n55 B 0.008855f
C205 VTAIL.n56 B 0.009376f
C206 VTAIL.n57 B 0.02093f
C207 VTAIL.n58 B 0.044719f
C208 VTAIL.n59 B 0.009376f
C209 VTAIL.n60 B 0.008855f
C210 VTAIL.n61 B 0.037414f
C211 VTAIL.n62 B 0.024941f
C212 VTAIL.n63 B 0.919103f
C213 VTAIL.n64 B 0.022828f
C214 VTAIL.n65 B 0.016478f
C215 VTAIL.n66 B 0.008855f
C216 VTAIL.n67 B 0.02093f
C217 VTAIL.n68 B 0.009376f
C218 VTAIL.n69 B 0.016478f
C219 VTAIL.n70 B 0.008855f
C220 VTAIL.n71 B 0.02093f
C221 VTAIL.n72 B 0.009376f
C222 VTAIL.n73 B 0.070379f
C223 VTAIL.t1 B 0.034104f
C224 VTAIL.n74 B 0.015697f
C225 VTAIL.n75 B 0.012363f
C226 VTAIL.n76 B 0.008855f
C227 VTAIL.n77 B 0.389844f
C228 VTAIL.n78 B 0.016478f
C229 VTAIL.n79 B 0.008855f
C230 VTAIL.n80 B 0.009376f
C231 VTAIL.n81 B 0.02093f
C232 VTAIL.n82 B 0.02093f
C233 VTAIL.n83 B 0.009376f
C234 VTAIL.n84 B 0.008855f
C235 VTAIL.n85 B 0.016478f
C236 VTAIL.n86 B 0.016478f
C237 VTAIL.n87 B 0.008855f
C238 VTAIL.n88 B 0.009376f
C239 VTAIL.n89 B 0.02093f
C240 VTAIL.n90 B 0.044719f
C241 VTAIL.n91 B 0.009376f
C242 VTAIL.n92 B 0.008855f
C243 VTAIL.n93 B 0.037414f
C244 VTAIL.n94 B 0.024941f
C245 VTAIL.n95 B 0.765761f
C246 VTAIL.n96 B 0.022828f
C247 VTAIL.n97 B 0.016478f
C248 VTAIL.n98 B 0.008855f
C249 VTAIL.n99 B 0.02093f
C250 VTAIL.n100 B 0.009376f
C251 VTAIL.n101 B 0.016478f
C252 VTAIL.n102 B 0.008855f
C253 VTAIL.n103 B 0.02093f
C254 VTAIL.n104 B 0.009376f
C255 VTAIL.n105 B 0.070379f
C256 VTAIL.t3 B 0.034104f
C257 VTAIL.n106 B 0.015697f
C258 VTAIL.n107 B 0.012363f
C259 VTAIL.n108 B 0.008855f
C260 VTAIL.n109 B 0.389844f
C261 VTAIL.n110 B 0.016478f
C262 VTAIL.n111 B 0.008855f
C263 VTAIL.n112 B 0.009376f
C264 VTAIL.n113 B 0.02093f
C265 VTAIL.n114 B 0.02093f
C266 VTAIL.n115 B 0.009376f
C267 VTAIL.n116 B 0.008855f
C268 VTAIL.n117 B 0.016478f
C269 VTAIL.n118 B 0.016478f
C270 VTAIL.n119 B 0.008855f
C271 VTAIL.n120 B 0.009376f
C272 VTAIL.n121 B 0.02093f
C273 VTAIL.n122 B 0.044719f
C274 VTAIL.n123 B 0.009376f
C275 VTAIL.n124 B 0.008855f
C276 VTAIL.n125 B 0.037414f
C277 VTAIL.n126 B 0.024941f
C278 VTAIL.n127 B 0.699389f
C279 VN.t0 B 1.11721f
C280 VN.t1 B 1.47006f
.ends

