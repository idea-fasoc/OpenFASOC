* NGSPICE file created from diff_pair_sample_1021.ext - technology: sky130A

.subckt diff_pair_sample_1021 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n2250_n4604# sky130_fd_pr__pfet_01v8 ad=7.0902 pd=37.14 as=7.0902 ps=37.14 w=18.18 l=2.87
X1 VDD1.t0 VP.t1 VTAIL.t2 w_n2250_n4604# sky130_fd_pr__pfet_01v8 ad=7.0902 pd=37.14 as=7.0902 ps=37.14 w=18.18 l=2.87
X2 VDD2.t1 VN.t0 VTAIL.t1 w_n2250_n4604# sky130_fd_pr__pfet_01v8 ad=7.0902 pd=37.14 as=7.0902 ps=37.14 w=18.18 l=2.87
X3 B.t11 B.t9 B.t10 w_n2250_n4604# sky130_fd_pr__pfet_01v8 ad=7.0902 pd=37.14 as=0 ps=0 w=18.18 l=2.87
X4 VDD2.t0 VN.t1 VTAIL.t0 w_n2250_n4604# sky130_fd_pr__pfet_01v8 ad=7.0902 pd=37.14 as=7.0902 ps=37.14 w=18.18 l=2.87
X5 B.t8 B.t6 B.t7 w_n2250_n4604# sky130_fd_pr__pfet_01v8 ad=7.0902 pd=37.14 as=0 ps=0 w=18.18 l=2.87
X6 B.t5 B.t3 B.t4 w_n2250_n4604# sky130_fd_pr__pfet_01v8 ad=7.0902 pd=37.14 as=0 ps=0 w=18.18 l=2.87
X7 B.t2 B.t0 B.t1 w_n2250_n4604# sky130_fd_pr__pfet_01v8 ad=7.0902 pd=37.14 as=0 ps=0 w=18.18 l=2.87
R0 VP.n0 VP.t0 243.855
R1 VP.n0 VP.t1 193.799
R2 VP VP.n0 0.431812
R3 VTAIL.n402 VTAIL.n306 756.745
R4 VTAIL.n96 VTAIL.n0 756.745
R5 VTAIL.n300 VTAIL.n204 756.745
R6 VTAIL.n198 VTAIL.n102 756.745
R7 VTAIL.n338 VTAIL.n337 585
R8 VTAIL.n343 VTAIL.n342 585
R9 VTAIL.n345 VTAIL.n344 585
R10 VTAIL.n334 VTAIL.n333 585
R11 VTAIL.n351 VTAIL.n350 585
R12 VTAIL.n353 VTAIL.n352 585
R13 VTAIL.n330 VTAIL.n329 585
R14 VTAIL.n359 VTAIL.n358 585
R15 VTAIL.n361 VTAIL.n360 585
R16 VTAIL.n326 VTAIL.n325 585
R17 VTAIL.n367 VTAIL.n366 585
R18 VTAIL.n369 VTAIL.n368 585
R19 VTAIL.n322 VTAIL.n321 585
R20 VTAIL.n375 VTAIL.n374 585
R21 VTAIL.n377 VTAIL.n376 585
R22 VTAIL.n318 VTAIL.n317 585
R23 VTAIL.n384 VTAIL.n383 585
R24 VTAIL.n385 VTAIL.n316 585
R25 VTAIL.n387 VTAIL.n386 585
R26 VTAIL.n314 VTAIL.n313 585
R27 VTAIL.n393 VTAIL.n392 585
R28 VTAIL.n395 VTAIL.n394 585
R29 VTAIL.n310 VTAIL.n309 585
R30 VTAIL.n401 VTAIL.n400 585
R31 VTAIL.n403 VTAIL.n402 585
R32 VTAIL.n32 VTAIL.n31 585
R33 VTAIL.n37 VTAIL.n36 585
R34 VTAIL.n39 VTAIL.n38 585
R35 VTAIL.n28 VTAIL.n27 585
R36 VTAIL.n45 VTAIL.n44 585
R37 VTAIL.n47 VTAIL.n46 585
R38 VTAIL.n24 VTAIL.n23 585
R39 VTAIL.n53 VTAIL.n52 585
R40 VTAIL.n55 VTAIL.n54 585
R41 VTAIL.n20 VTAIL.n19 585
R42 VTAIL.n61 VTAIL.n60 585
R43 VTAIL.n63 VTAIL.n62 585
R44 VTAIL.n16 VTAIL.n15 585
R45 VTAIL.n69 VTAIL.n68 585
R46 VTAIL.n71 VTAIL.n70 585
R47 VTAIL.n12 VTAIL.n11 585
R48 VTAIL.n78 VTAIL.n77 585
R49 VTAIL.n79 VTAIL.n10 585
R50 VTAIL.n81 VTAIL.n80 585
R51 VTAIL.n8 VTAIL.n7 585
R52 VTAIL.n87 VTAIL.n86 585
R53 VTAIL.n89 VTAIL.n88 585
R54 VTAIL.n4 VTAIL.n3 585
R55 VTAIL.n95 VTAIL.n94 585
R56 VTAIL.n97 VTAIL.n96 585
R57 VTAIL.n301 VTAIL.n300 585
R58 VTAIL.n299 VTAIL.n298 585
R59 VTAIL.n208 VTAIL.n207 585
R60 VTAIL.n293 VTAIL.n292 585
R61 VTAIL.n291 VTAIL.n290 585
R62 VTAIL.n212 VTAIL.n211 585
R63 VTAIL.n285 VTAIL.n284 585
R64 VTAIL.n283 VTAIL.n214 585
R65 VTAIL.n282 VTAIL.n281 585
R66 VTAIL.n217 VTAIL.n215 585
R67 VTAIL.n276 VTAIL.n275 585
R68 VTAIL.n274 VTAIL.n273 585
R69 VTAIL.n221 VTAIL.n220 585
R70 VTAIL.n268 VTAIL.n267 585
R71 VTAIL.n266 VTAIL.n265 585
R72 VTAIL.n225 VTAIL.n224 585
R73 VTAIL.n260 VTAIL.n259 585
R74 VTAIL.n258 VTAIL.n257 585
R75 VTAIL.n229 VTAIL.n228 585
R76 VTAIL.n252 VTAIL.n251 585
R77 VTAIL.n250 VTAIL.n249 585
R78 VTAIL.n233 VTAIL.n232 585
R79 VTAIL.n244 VTAIL.n243 585
R80 VTAIL.n242 VTAIL.n241 585
R81 VTAIL.n237 VTAIL.n236 585
R82 VTAIL.n199 VTAIL.n198 585
R83 VTAIL.n197 VTAIL.n196 585
R84 VTAIL.n106 VTAIL.n105 585
R85 VTAIL.n191 VTAIL.n190 585
R86 VTAIL.n189 VTAIL.n188 585
R87 VTAIL.n110 VTAIL.n109 585
R88 VTAIL.n183 VTAIL.n182 585
R89 VTAIL.n181 VTAIL.n112 585
R90 VTAIL.n180 VTAIL.n179 585
R91 VTAIL.n115 VTAIL.n113 585
R92 VTAIL.n174 VTAIL.n173 585
R93 VTAIL.n172 VTAIL.n171 585
R94 VTAIL.n119 VTAIL.n118 585
R95 VTAIL.n166 VTAIL.n165 585
R96 VTAIL.n164 VTAIL.n163 585
R97 VTAIL.n123 VTAIL.n122 585
R98 VTAIL.n158 VTAIL.n157 585
R99 VTAIL.n156 VTAIL.n155 585
R100 VTAIL.n127 VTAIL.n126 585
R101 VTAIL.n150 VTAIL.n149 585
R102 VTAIL.n148 VTAIL.n147 585
R103 VTAIL.n131 VTAIL.n130 585
R104 VTAIL.n142 VTAIL.n141 585
R105 VTAIL.n140 VTAIL.n139 585
R106 VTAIL.n135 VTAIL.n134 585
R107 VTAIL.n339 VTAIL.t0 327.466
R108 VTAIL.n33 VTAIL.t2 327.466
R109 VTAIL.n238 VTAIL.t3 327.466
R110 VTAIL.n136 VTAIL.t1 327.466
R111 VTAIL.n343 VTAIL.n337 171.744
R112 VTAIL.n344 VTAIL.n343 171.744
R113 VTAIL.n344 VTAIL.n333 171.744
R114 VTAIL.n351 VTAIL.n333 171.744
R115 VTAIL.n352 VTAIL.n351 171.744
R116 VTAIL.n352 VTAIL.n329 171.744
R117 VTAIL.n359 VTAIL.n329 171.744
R118 VTAIL.n360 VTAIL.n359 171.744
R119 VTAIL.n360 VTAIL.n325 171.744
R120 VTAIL.n367 VTAIL.n325 171.744
R121 VTAIL.n368 VTAIL.n367 171.744
R122 VTAIL.n368 VTAIL.n321 171.744
R123 VTAIL.n375 VTAIL.n321 171.744
R124 VTAIL.n376 VTAIL.n375 171.744
R125 VTAIL.n376 VTAIL.n317 171.744
R126 VTAIL.n384 VTAIL.n317 171.744
R127 VTAIL.n385 VTAIL.n384 171.744
R128 VTAIL.n386 VTAIL.n385 171.744
R129 VTAIL.n386 VTAIL.n313 171.744
R130 VTAIL.n393 VTAIL.n313 171.744
R131 VTAIL.n394 VTAIL.n393 171.744
R132 VTAIL.n394 VTAIL.n309 171.744
R133 VTAIL.n401 VTAIL.n309 171.744
R134 VTAIL.n402 VTAIL.n401 171.744
R135 VTAIL.n37 VTAIL.n31 171.744
R136 VTAIL.n38 VTAIL.n37 171.744
R137 VTAIL.n38 VTAIL.n27 171.744
R138 VTAIL.n45 VTAIL.n27 171.744
R139 VTAIL.n46 VTAIL.n45 171.744
R140 VTAIL.n46 VTAIL.n23 171.744
R141 VTAIL.n53 VTAIL.n23 171.744
R142 VTAIL.n54 VTAIL.n53 171.744
R143 VTAIL.n54 VTAIL.n19 171.744
R144 VTAIL.n61 VTAIL.n19 171.744
R145 VTAIL.n62 VTAIL.n61 171.744
R146 VTAIL.n62 VTAIL.n15 171.744
R147 VTAIL.n69 VTAIL.n15 171.744
R148 VTAIL.n70 VTAIL.n69 171.744
R149 VTAIL.n70 VTAIL.n11 171.744
R150 VTAIL.n78 VTAIL.n11 171.744
R151 VTAIL.n79 VTAIL.n78 171.744
R152 VTAIL.n80 VTAIL.n79 171.744
R153 VTAIL.n80 VTAIL.n7 171.744
R154 VTAIL.n87 VTAIL.n7 171.744
R155 VTAIL.n88 VTAIL.n87 171.744
R156 VTAIL.n88 VTAIL.n3 171.744
R157 VTAIL.n95 VTAIL.n3 171.744
R158 VTAIL.n96 VTAIL.n95 171.744
R159 VTAIL.n300 VTAIL.n299 171.744
R160 VTAIL.n299 VTAIL.n207 171.744
R161 VTAIL.n292 VTAIL.n207 171.744
R162 VTAIL.n292 VTAIL.n291 171.744
R163 VTAIL.n291 VTAIL.n211 171.744
R164 VTAIL.n284 VTAIL.n211 171.744
R165 VTAIL.n284 VTAIL.n283 171.744
R166 VTAIL.n283 VTAIL.n282 171.744
R167 VTAIL.n282 VTAIL.n215 171.744
R168 VTAIL.n275 VTAIL.n215 171.744
R169 VTAIL.n275 VTAIL.n274 171.744
R170 VTAIL.n274 VTAIL.n220 171.744
R171 VTAIL.n267 VTAIL.n220 171.744
R172 VTAIL.n267 VTAIL.n266 171.744
R173 VTAIL.n266 VTAIL.n224 171.744
R174 VTAIL.n259 VTAIL.n224 171.744
R175 VTAIL.n259 VTAIL.n258 171.744
R176 VTAIL.n258 VTAIL.n228 171.744
R177 VTAIL.n251 VTAIL.n228 171.744
R178 VTAIL.n251 VTAIL.n250 171.744
R179 VTAIL.n250 VTAIL.n232 171.744
R180 VTAIL.n243 VTAIL.n232 171.744
R181 VTAIL.n243 VTAIL.n242 171.744
R182 VTAIL.n242 VTAIL.n236 171.744
R183 VTAIL.n198 VTAIL.n197 171.744
R184 VTAIL.n197 VTAIL.n105 171.744
R185 VTAIL.n190 VTAIL.n105 171.744
R186 VTAIL.n190 VTAIL.n189 171.744
R187 VTAIL.n189 VTAIL.n109 171.744
R188 VTAIL.n182 VTAIL.n109 171.744
R189 VTAIL.n182 VTAIL.n181 171.744
R190 VTAIL.n181 VTAIL.n180 171.744
R191 VTAIL.n180 VTAIL.n113 171.744
R192 VTAIL.n173 VTAIL.n113 171.744
R193 VTAIL.n173 VTAIL.n172 171.744
R194 VTAIL.n172 VTAIL.n118 171.744
R195 VTAIL.n165 VTAIL.n118 171.744
R196 VTAIL.n165 VTAIL.n164 171.744
R197 VTAIL.n164 VTAIL.n122 171.744
R198 VTAIL.n157 VTAIL.n122 171.744
R199 VTAIL.n157 VTAIL.n156 171.744
R200 VTAIL.n156 VTAIL.n126 171.744
R201 VTAIL.n149 VTAIL.n126 171.744
R202 VTAIL.n149 VTAIL.n148 171.744
R203 VTAIL.n148 VTAIL.n130 171.744
R204 VTAIL.n141 VTAIL.n130 171.744
R205 VTAIL.n141 VTAIL.n140 171.744
R206 VTAIL.n140 VTAIL.n134 171.744
R207 VTAIL.t0 VTAIL.n337 85.8723
R208 VTAIL.t2 VTAIL.n31 85.8723
R209 VTAIL.t3 VTAIL.n236 85.8723
R210 VTAIL.t1 VTAIL.n134 85.8723
R211 VTAIL.n203 VTAIL.n101 33.5565
R212 VTAIL.n407 VTAIL.n406 31.0217
R213 VTAIL.n101 VTAIL.n100 31.0217
R214 VTAIL.n305 VTAIL.n304 31.0217
R215 VTAIL.n203 VTAIL.n202 31.0217
R216 VTAIL.n407 VTAIL.n305 30.7979
R217 VTAIL.n339 VTAIL.n338 16.3895
R218 VTAIL.n33 VTAIL.n32 16.3895
R219 VTAIL.n238 VTAIL.n237 16.3895
R220 VTAIL.n136 VTAIL.n135 16.3895
R221 VTAIL.n387 VTAIL.n316 13.1884
R222 VTAIL.n81 VTAIL.n10 13.1884
R223 VTAIL.n285 VTAIL.n214 13.1884
R224 VTAIL.n183 VTAIL.n112 13.1884
R225 VTAIL.n342 VTAIL.n341 12.8005
R226 VTAIL.n383 VTAIL.n382 12.8005
R227 VTAIL.n388 VTAIL.n314 12.8005
R228 VTAIL.n36 VTAIL.n35 12.8005
R229 VTAIL.n77 VTAIL.n76 12.8005
R230 VTAIL.n82 VTAIL.n8 12.8005
R231 VTAIL.n286 VTAIL.n212 12.8005
R232 VTAIL.n281 VTAIL.n216 12.8005
R233 VTAIL.n241 VTAIL.n240 12.8005
R234 VTAIL.n184 VTAIL.n110 12.8005
R235 VTAIL.n179 VTAIL.n114 12.8005
R236 VTAIL.n139 VTAIL.n138 12.8005
R237 VTAIL.n345 VTAIL.n336 12.0247
R238 VTAIL.n381 VTAIL.n318 12.0247
R239 VTAIL.n392 VTAIL.n391 12.0247
R240 VTAIL.n39 VTAIL.n30 12.0247
R241 VTAIL.n75 VTAIL.n12 12.0247
R242 VTAIL.n86 VTAIL.n85 12.0247
R243 VTAIL.n290 VTAIL.n289 12.0247
R244 VTAIL.n280 VTAIL.n217 12.0247
R245 VTAIL.n244 VTAIL.n235 12.0247
R246 VTAIL.n188 VTAIL.n187 12.0247
R247 VTAIL.n178 VTAIL.n115 12.0247
R248 VTAIL.n142 VTAIL.n133 12.0247
R249 VTAIL.n346 VTAIL.n334 11.249
R250 VTAIL.n378 VTAIL.n377 11.249
R251 VTAIL.n395 VTAIL.n312 11.249
R252 VTAIL.n40 VTAIL.n28 11.249
R253 VTAIL.n72 VTAIL.n71 11.249
R254 VTAIL.n89 VTAIL.n6 11.249
R255 VTAIL.n293 VTAIL.n210 11.249
R256 VTAIL.n277 VTAIL.n276 11.249
R257 VTAIL.n245 VTAIL.n233 11.249
R258 VTAIL.n191 VTAIL.n108 11.249
R259 VTAIL.n175 VTAIL.n174 11.249
R260 VTAIL.n143 VTAIL.n131 11.249
R261 VTAIL.n350 VTAIL.n349 10.4732
R262 VTAIL.n374 VTAIL.n320 10.4732
R263 VTAIL.n396 VTAIL.n310 10.4732
R264 VTAIL.n44 VTAIL.n43 10.4732
R265 VTAIL.n68 VTAIL.n14 10.4732
R266 VTAIL.n90 VTAIL.n4 10.4732
R267 VTAIL.n294 VTAIL.n208 10.4732
R268 VTAIL.n273 VTAIL.n219 10.4732
R269 VTAIL.n249 VTAIL.n248 10.4732
R270 VTAIL.n192 VTAIL.n106 10.4732
R271 VTAIL.n171 VTAIL.n117 10.4732
R272 VTAIL.n147 VTAIL.n146 10.4732
R273 VTAIL.n353 VTAIL.n332 9.69747
R274 VTAIL.n373 VTAIL.n322 9.69747
R275 VTAIL.n400 VTAIL.n399 9.69747
R276 VTAIL.n47 VTAIL.n26 9.69747
R277 VTAIL.n67 VTAIL.n16 9.69747
R278 VTAIL.n94 VTAIL.n93 9.69747
R279 VTAIL.n298 VTAIL.n297 9.69747
R280 VTAIL.n272 VTAIL.n221 9.69747
R281 VTAIL.n252 VTAIL.n231 9.69747
R282 VTAIL.n196 VTAIL.n195 9.69747
R283 VTAIL.n170 VTAIL.n119 9.69747
R284 VTAIL.n150 VTAIL.n129 9.69747
R285 VTAIL.n406 VTAIL.n405 9.45567
R286 VTAIL.n100 VTAIL.n99 9.45567
R287 VTAIL.n304 VTAIL.n303 9.45567
R288 VTAIL.n202 VTAIL.n201 9.45567
R289 VTAIL.n405 VTAIL.n404 9.3005
R290 VTAIL.n308 VTAIL.n307 9.3005
R291 VTAIL.n399 VTAIL.n398 9.3005
R292 VTAIL.n397 VTAIL.n396 9.3005
R293 VTAIL.n312 VTAIL.n311 9.3005
R294 VTAIL.n391 VTAIL.n390 9.3005
R295 VTAIL.n389 VTAIL.n388 9.3005
R296 VTAIL.n328 VTAIL.n327 9.3005
R297 VTAIL.n357 VTAIL.n356 9.3005
R298 VTAIL.n355 VTAIL.n354 9.3005
R299 VTAIL.n332 VTAIL.n331 9.3005
R300 VTAIL.n349 VTAIL.n348 9.3005
R301 VTAIL.n347 VTAIL.n346 9.3005
R302 VTAIL.n336 VTAIL.n335 9.3005
R303 VTAIL.n341 VTAIL.n340 9.3005
R304 VTAIL.n363 VTAIL.n362 9.3005
R305 VTAIL.n365 VTAIL.n364 9.3005
R306 VTAIL.n324 VTAIL.n323 9.3005
R307 VTAIL.n371 VTAIL.n370 9.3005
R308 VTAIL.n373 VTAIL.n372 9.3005
R309 VTAIL.n320 VTAIL.n319 9.3005
R310 VTAIL.n379 VTAIL.n378 9.3005
R311 VTAIL.n381 VTAIL.n380 9.3005
R312 VTAIL.n382 VTAIL.n315 9.3005
R313 VTAIL.n99 VTAIL.n98 9.3005
R314 VTAIL.n2 VTAIL.n1 9.3005
R315 VTAIL.n93 VTAIL.n92 9.3005
R316 VTAIL.n91 VTAIL.n90 9.3005
R317 VTAIL.n6 VTAIL.n5 9.3005
R318 VTAIL.n85 VTAIL.n84 9.3005
R319 VTAIL.n83 VTAIL.n82 9.3005
R320 VTAIL.n22 VTAIL.n21 9.3005
R321 VTAIL.n51 VTAIL.n50 9.3005
R322 VTAIL.n49 VTAIL.n48 9.3005
R323 VTAIL.n26 VTAIL.n25 9.3005
R324 VTAIL.n43 VTAIL.n42 9.3005
R325 VTAIL.n41 VTAIL.n40 9.3005
R326 VTAIL.n30 VTAIL.n29 9.3005
R327 VTAIL.n35 VTAIL.n34 9.3005
R328 VTAIL.n57 VTAIL.n56 9.3005
R329 VTAIL.n59 VTAIL.n58 9.3005
R330 VTAIL.n18 VTAIL.n17 9.3005
R331 VTAIL.n65 VTAIL.n64 9.3005
R332 VTAIL.n67 VTAIL.n66 9.3005
R333 VTAIL.n14 VTAIL.n13 9.3005
R334 VTAIL.n73 VTAIL.n72 9.3005
R335 VTAIL.n75 VTAIL.n74 9.3005
R336 VTAIL.n76 VTAIL.n9 9.3005
R337 VTAIL.n264 VTAIL.n263 9.3005
R338 VTAIL.n223 VTAIL.n222 9.3005
R339 VTAIL.n270 VTAIL.n269 9.3005
R340 VTAIL.n272 VTAIL.n271 9.3005
R341 VTAIL.n219 VTAIL.n218 9.3005
R342 VTAIL.n278 VTAIL.n277 9.3005
R343 VTAIL.n280 VTAIL.n279 9.3005
R344 VTAIL.n216 VTAIL.n213 9.3005
R345 VTAIL.n303 VTAIL.n302 9.3005
R346 VTAIL.n206 VTAIL.n205 9.3005
R347 VTAIL.n297 VTAIL.n296 9.3005
R348 VTAIL.n295 VTAIL.n294 9.3005
R349 VTAIL.n210 VTAIL.n209 9.3005
R350 VTAIL.n289 VTAIL.n288 9.3005
R351 VTAIL.n287 VTAIL.n286 9.3005
R352 VTAIL.n262 VTAIL.n261 9.3005
R353 VTAIL.n227 VTAIL.n226 9.3005
R354 VTAIL.n256 VTAIL.n255 9.3005
R355 VTAIL.n254 VTAIL.n253 9.3005
R356 VTAIL.n231 VTAIL.n230 9.3005
R357 VTAIL.n248 VTAIL.n247 9.3005
R358 VTAIL.n246 VTAIL.n245 9.3005
R359 VTAIL.n235 VTAIL.n234 9.3005
R360 VTAIL.n240 VTAIL.n239 9.3005
R361 VTAIL.n162 VTAIL.n161 9.3005
R362 VTAIL.n121 VTAIL.n120 9.3005
R363 VTAIL.n168 VTAIL.n167 9.3005
R364 VTAIL.n170 VTAIL.n169 9.3005
R365 VTAIL.n117 VTAIL.n116 9.3005
R366 VTAIL.n176 VTAIL.n175 9.3005
R367 VTAIL.n178 VTAIL.n177 9.3005
R368 VTAIL.n114 VTAIL.n111 9.3005
R369 VTAIL.n201 VTAIL.n200 9.3005
R370 VTAIL.n104 VTAIL.n103 9.3005
R371 VTAIL.n195 VTAIL.n194 9.3005
R372 VTAIL.n193 VTAIL.n192 9.3005
R373 VTAIL.n108 VTAIL.n107 9.3005
R374 VTAIL.n187 VTAIL.n186 9.3005
R375 VTAIL.n185 VTAIL.n184 9.3005
R376 VTAIL.n160 VTAIL.n159 9.3005
R377 VTAIL.n125 VTAIL.n124 9.3005
R378 VTAIL.n154 VTAIL.n153 9.3005
R379 VTAIL.n152 VTAIL.n151 9.3005
R380 VTAIL.n129 VTAIL.n128 9.3005
R381 VTAIL.n146 VTAIL.n145 9.3005
R382 VTAIL.n144 VTAIL.n143 9.3005
R383 VTAIL.n133 VTAIL.n132 9.3005
R384 VTAIL.n138 VTAIL.n137 9.3005
R385 VTAIL.n354 VTAIL.n330 8.92171
R386 VTAIL.n370 VTAIL.n369 8.92171
R387 VTAIL.n403 VTAIL.n308 8.92171
R388 VTAIL.n48 VTAIL.n24 8.92171
R389 VTAIL.n64 VTAIL.n63 8.92171
R390 VTAIL.n97 VTAIL.n2 8.92171
R391 VTAIL.n301 VTAIL.n206 8.92171
R392 VTAIL.n269 VTAIL.n268 8.92171
R393 VTAIL.n253 VTAIL.n229 8.92171
R394 VTAIL.n199 VTAIL.n104 8.92171
R395 VTAIL.n167 VTAIL.n166 8.92171
R396 VTAIL.n151 VTAIL.n127 8.92171
R397 VTAIL.n358 VTAIL.n357 8.14595
R398 VTAIL.n366 VTAIL.n324 8.14595
R399 VTAIL.n404 VTAIL.n306 8.14595
R400 VTAIL.n52 VTAIL.n51 8.14595
R401 VTAIL.n60 VTAIL.n18 8.14595
R402 VTAIL.n98 VTAIL.n0 8.14595
R403 VTAIL.n302 VTAIL.n204 8.14595
R404 VTAIL.n265 VTAIL.n223 8.14595
R405 VTAIL.n257 VTAIL.n256 8.14595
R406 VTAIL.n200 VTAIL.n102 8.14595
R407 VTAIL.n163 VTAIL.n121 8.14595
R408 VTAIL.n155 VTAIL.n154 8.14595
R409 VTAIL.n361 VTAIL.n328 7.3702
R410 VTAIL.n365 VTAIL.n326 7.3702
R411 VTAIL.n55 VTAIL.n22 7.3702
R412 VTAIL.n59 VTAIL.n20 7.3702
R413 VTAIL.n264 VTAIL.n225 7.3702
R414 VTAIL.n260 VTAIL.n227 7.3702
R415 VTAIL.n162 VTAIL.n123 7.3702
R416 VTAIL.n158 VTAIL.n125 7.3702
R417 VTAIL.n362 VTAIL.n361 6.59444
R418 VTAIL.n362 VTAIL.n326 6.59444
R419 VTAIL.n56 VTAIL.n55 6.59444
R420 VTAIL.n56 VTAIL.n20 6.59444
R421 VTAIL.n261 VTAIL.n225 6.59444
R422 VTAIL.n261 VTAIL.n260 6.59444
R423 VTAIL.n159 VTAIL.n123 6.59444
R424 VTAIL.n159 VTAIL.n158 6.59444
R425 VTAIL.n358 VTAIL.n328 5.81868
R426 VTAIL.n366 VTAIL.n365 5.81868
R427 VTAIL.n406 VTAIL.n306 5.81868
R428 VTAIL.n52 VTAIL.n22 5.81868
R429 VTAIL.n60 VTAIL.n59 5.81868
R430 VTAIL.n100 VTAIL.n0 5.81868
R431 VTAIL.n304 VTAIL.n204 5.81868
R432 VTAIL.n265 VTAIL.n264 5.81868
R433 VTAIL.n257 VTAIL.n227 5.81868
R434 VTAIL.n202 VTAIL.n102 5.81868
R435 VTAIL.n163 VTAIL.n162 5.81868
R436 VTAIL.n155 VTAIL.n125 5.81868
R437 VTAIL.n357 VTAIL.n330 5.04292
R438 VTAIL.n369 VTAIL.n324 5.04292
R439 VTAIL.n404 VTAIL.n403 5.04292
R440 VTAIL.n51 VTAIL.n24 5.04292
R441 VTAIL.n63 VTAIL.n18 5.04292
R442 VTAIL.n98 VTAIL.n97 5.04292
R443 VTAIL.n302 VTAIL.n301 5.04292
R444 VTAIL.n268 VTAIL.n223 5.04292
R445 VTAIL.n256 VTAIL.n229 5.04292
R446 VTAIL.n200 VTAIL.n199 5.04292
R447 VTAIL.n166 VTAIL.n121 5.04292
R448 VTAIL.n154 VTAIL.n127 5.04292
R449 VTAIL.n354 VTAIL.n353 4.26717
R450 VTAIL.n370 VTAIL.n322 4.26717
R451 VTAIL.n400 VTAIL.n308 4.26717
R452 VTAIL.n48 VTAIL.n47 4.26717
R453 VTAIL.n64 VTAIL.n16 4.26717
R454 VTAIL.n94 VTAIL.n2 4.26717
R455 VTAIL.n298 VTAIL.n206 4.26717
R456 VTAIL.n269 VTAIL.n221 4.26717
R457 VTAIL.n253 VTAIL.n252 4.26717
R458 VTAIL.n196 VTAIL.n104 4.26717
R459 VTAIL.n167 VTAIL.n119 4.26717
R460 VTAIL.n151 VTAIL.n150 4.26717
R461 VTAIL.n340 VTAIL.n339 3.70982
R462 VTAIL.n34 VTAIL.n33 3.70982
R463 VTAIL.n239 VTAIL.n238 3.70982
R464 VTAIL.n137 VTAIL.n136 3.70982
R465 VTAIL.n350 VTAIL.n332 3.49141
R466 VTAIL.n374 VTAIL.n373 3.49141
R467 VTAIL.n399 VTAIL.n310 3.49141
R468 VTAIL.n44 VTAIL.n26 3.49141
R469 VTAIL.n68 VTAIL.n67 3.49141
R470 VTAIL.n93 VTAIL.n4 3.49141
R471 VTAIL.n297 VTAIL.n208 3.49141
R472 VTAIL.n273 VTAIL.n272 3.49141
R473 VTAIL.n249 VTAIL.n231 3.49141
R474 VTAIL.n195 VTAIL.n106 3.49141
R475 VTAIL.n171 VTAIL.n170 3.49141
R476 VTAIL.n147 VTAIL.n129 3.49141
R477 VTAIL.n349 VTAIL.n334 2.71565
R478 VTAIL.n377 VTAIL.n320 2.71565
R479 VTAIL.n396 VTAIL.n395 2.71565
R480 VTAIL.n43 VTAIL.n28 2.71565
R481 VTAIL.n71 VTAIL.n14 2.71565
R482 VTAIL.n90 VTAIL.n89 2.71565
R483 VTAIL.n294 VTAIL.n293 2.71565
R484 VTAIL.n276 VTAIL.n219 2.71565
R485 VTAIL.n248 VTAIL.n233 2.71565
R486 VTAIL.n192 VTAIL.n191 2.71565
R487 VTAIL.n174 VTAIL.n117 2.71565
R488 VTAIL.n146 VTAIL.n131 2.71565
R489 VTAIL.n346 VTAIL.n345 1.93989
R490 VTAIL.n378 VTAIL.n318 1.93989
R491 VTAIL.n392 VTAIL.n312 1.93989
R492 VTAIL.n40 VTAIL.n39 1.93989
R493 VTAIL.n72 VTAIL.n12 1.93989
R494 VTAIL.n86 VTAIL.n6 1.93989
R495 VTAIL.n290 VTAIL.n210 1.93989
R496 VTAIL.n277 VTAIL.n217 1.93989
R497 VTAIL.n245 VTAIL.n244 1.93989
R498 VTAIL.n188 VTAIL.n108 1.93989
R499 VTAIL.n175 VTAIL.n115 1.93989
R500 VTAIL.n143 VTAIL.n142 1.93989
R501 VTAIL.n305 VTAIL.n203 1.84964
R502 VTAIL VTAIL.n101 1.21817
R503 VTAIL.n342 VTAIL.n336 1.16414
R504 VTAIL.n383 VTAIL.n381 1.16414
R505 VTAIL.n391 VTAIL.n314 1.16414
R506 VTAIL.n36 VTAIL.n30 1.16414
R507 VTAIL.n77 VTAIL.n75 1.16414
R508 VTAIL.n85 VTAIL.n8 1.16414
R509 VTAIL.n289 VTAIL.n212 1.16414
R510 VTAIL.n281 VTAIL.n280 1.16414
R511 VTAIL.n241 VTAIL.n235 1.16414
R512 VTAIL.n187 VTAIL.n110 1.16414
R513 VTAIL.n179 VTAIL.n178 1.16414
R514 VTAIL.n139 VTAIL.n133 1.16414
R515 VTAIL VTAIL.n407 0.631965
R516 VTAIL.n341 VTAIL.n338 0.388379
R517 VTAIL.n382 VTAIL.n316 0.388379
R518 VTAIL.n388 VTAIL.n387 0.388379
R519 VTAIL.n35 VTAIL.n32 0.388379
R520 VTAIL.n76 VTAIL.n10 0.388379
R521 VTAIL.n82 VTAIL.n81 0.388379
R522 VTAIL.n286 VTAIL.n285 0.388379
R523 VTAIL.n216 VTAIL.n214 0.388379
R524 VTAIL.n240 VTAIL.n237 0.388379
R525 VTAIL.n184 VTAIL.n183 0.388379
R526 VTAIL.n114 VTAIL.n112 0.388379
R527 VTAIL.n138 VTAIL.n135 0.388379
R528 VTAIL.n340 VTAIL.n335 0.155672
R529 VTAIL.n347 VTAIL.n335 0.155672
R530 VTAIL.n348 VTAIL.n347 0.155672
R531 VTAIL.n348 VTAIL.n331 0.155672
R532 VTAIL.n355 VTAIL.n331 0.155672
R533 VTAIL.n356 VTAIL.n355 0.155672
R534 VTAIL.n356 VTAIL.n327 0.155672
R535 VTAIL.n363 VTAIL.n327 0.155672
R536 VTAIL.n364 VTAIL.n363 0.155672
R537 VTAIL.n364 VTAIL.n323 0.155672
R538 VTAIL.n371 VTAIL.n323 0.155672
R539 VTAIL.n372 VTAIL.n371 0.155672
R540 VTAIL.n372 VTAIL.n319 0.155672
R541 VTAIL.n379 VTAIL.n319 0.155672
R542 VTAIL.n380 VTAIL.n379 0.155672
R543 VTAIL.n380 VTAIL.n315 0.155672
R544 VTAIL.n389 VTAIL.n315 0.155672
R545 VTAIL.n390 VTAIL.n389 0.155672
R546 VTAIL.n390 VTAIL.n311 0.155672
R547 VTAIL.n397 VTAIL.n311 0.155672
R548 VTAIL.n398 VTAIL.n397 0.155672
R549 VTAIL.n398 VTAIL.n307 0.155672
R550 VTAIL.n405 VTAIL.n307 0.155672
R551 VTAIL.n34 VTAIL.n29 0.155672
R552 VTAIL.n41 VTAIL.n29 0.155672
R553 VTAIL.n42 VTAIL.n41 0.155672
R554 VTAIL.n42 VTAIL.n25 0.155672
R555 VTAIL.n49 VTAIL.n25 0.155672
R556 VTAIL.n50 VTAIL.n49 0.155672
R557 VTAIL.n50 VTAIL.n21 0.155672
R558 VTAIL.n57 VTAIL.n21 0.155672
R559 VTAIL.n58 VTAIL.n57 0.155672
R560 VTAIL.n58 VTAIL.n17 0.155672
R561 VTAIL.n65 VTAIL.n17 0.155672
R562 VTAIL.n66 VTAIL.n65 0.155672
R563 VTAIL.n66 VTAIL.n13 0.155672
R564 VTAIL.n73 VTAIL.n13 0.155672
R565 VTAIL.n74 VTAIL.n73 0.155672
R566 VTAIL.n74 VTAIL.n9 0.155672
R567 VTAIL.n83 VTAIL.n9 0.155672
R568 VTAIL.n84 VTAIL.n83 0.155672
R569 VTAIL.n84 VTAIL.n5 0.155672
R570 VTAIL.n91 VTAIL.n5 0.155672
R571 VTAIL.n92 VTAIL.n91 0.155672
R572 VTAIL.n92 VTAIL.n1 0.155672
R573 VTAIL.n99 VTAIL.n1 0.155672
R574 VTAIL.n303 VTAIL.n205 0.155672
R575 VTAIL.n296 VTAIL.n205 0.155672
R576 VTAIL.n296 VTAIL.n295 0.155672
R577 VTAIL.n295 VTAIL.n209 0.155672
R578 VTAIL.n288 VTAIL.n209 0.155672
R579 VTAIL.n288 VTAIL.n287 0.155672
R580 VTAIL.n287 VTAIL.n213 0.155672
R581 VTAIL.n279 VTAIL.n213 0.155672
R582 VTAIL.n279 VTAIL.n278 0.155672
R583 VTAIL.n278 VTAIL.n218 0.155672
R584 VTAIL.n271 VTAIL.n218 0.155672
R585 VTAIL.n271 VTAIL.n270 0.155672
R586 VTAIL.n270 VTAIL.n222 0.155672
R587 VTAIL.n263 VTAIL.n222 0.155672
R588 VTAIL.n263 VTAIL.n262 0.155672
R589 VTAIL.n262 VTAIL.n226 0.155672
R590 VTAIL.n255 VTAIL.n226 0.155672
R591 VTAIL.n255 VTAIL.n254 0.155672
R592 VTAIL.n254 VTAIL.n230 0.155672
R593 VTAIL.n247 VTAIL.n230 0.155672
R594 VTAIL.n247 VTAIL.n246 0.155672
R595 VTAIL.n246 VTAIL.n234 0.155672
R596 VTAIL.n239 VTAIL.n234 0.155672
R597 VTAIL.n201 VTAIL.n103 0.155672
R598 VTAIL.n194 VTAIL.n103 0.155672
R599 VTAIL.n194 VTAIL.n193 0.155672
R600 VTAIL.n193 VTAIL.n107 0.155672
R601 VTAIL.n186 VTAIL.n107 0.155672
R602 VTAIL.n186 VTAIL.n185 0.155672
R603 VTAIL.n185 VTAIL.n111 0.155672
R604 VTAIL.n177 VTAIL.n111 0.155672
R605 VTAIL.n177 VTAIL.n176 0.155672
R606 VTAIL.n176 VTAIL.n116 0.155672
R607 VTAIL.n169 VTAIL.n116 0.155672
R608 VTAIL.n169 VTAIL.n168 0.155672
R609 VTAIL.n168 VTAIL.n120 0.155672
R610 VTAIL.n161 VTAIL.n120 0.155672
R611 VTAIL.n161 VTAIL.n160 0.155672
R612 VTAIL.n160 VTAIL.n124 0.155672
R613 VTAIL.n153 VTAIL.n124 0.155672
R614 VTAIL.n153 VTAIL.n152 0.155672
R615 VTAIL.n152 VTAIL.n128 0.155672
R616 VTAIL.n145 VTAIL.n128 0.155672
R617 VTAIL.n145 VTAIL.n144 0.155672
R618 VTAIL.n144 VTAIL.n132 0.155672
R619 VTAIL.n137 VTAIL.n132 0.155672
R620 VDD1.n96 VDD1.n0 756.745
R621 VDD1.n197 VDD1.n101 756.745
R622 VDD1.n97 VDD1.n96 585
R623 VDD1.n95 VDD1.n94 585
R624 VDD1.n4 VDD1.n3 585
R625 VDD1.n89 VDD1.n88 585
R626 VDD1.n87 VDD1.n86 585
R627 VDD1.n8 VDD1.n7 585
R628 VDD1.n81 VDD1.n80 585
R629 VDD1.n79 VDD1.n10 585
R630 VDD1.n78 VDD1.n77 585
R631 VDD1.n13 VDD1.n11 585
R632 VDD1.n72 VDD1.n71 585
R633 VDD1.n70 VDD1.n69 585
R634 VDD1.n17 VDD1.n16 585
R635 VDD1.n64 VDD1.n63 585
R636 VDD1.n62 VDD1.n61 585
R637 VDD1.n21 VDD1.n20 585
R638 VDD1.n56 VDD1.n55 585
R639 VDD1.n54 VDD1.n53 585
R640 VDD1.n25 VDD1.n24 585
R641 VDD1.n48 VDD1.n47 585
R642 VDD1.n46 VDD1.n45 585
R643 VDD1.n29 VDD1.n28 585
R644 VDD1.n40 VDD1.n39 585
R645 VDD1.n38 VDD1.n37 585
R646 VDD1.n33 VDD1.n32 585
R647 VDD1.n133 VDD1.n132 585
R648 VDD1.n138 VDD1.n137 585
R649 VDD1.n140 VDD1.n139 585
R650 VDD1.n129 VDD1.n128 585
R651 VDD1.n146 VDD1.n145 585
R652 VDD1.n148 VDD1.n147 585
R653 VDD1.n125 VDD1.n124 585
R654 VDD1.n154 VDD1.n153 585
R655 VDD1.n156 VDD1.n155 585
R656 VDD1.n121 VDD1.n120 585
R657 VDD1.n162 VDD1.n161 585
R658 VDD1.n164 VDD1.n163 585
R659 VDD1.n117 VDD1.n116 585
R660 VDD1.n170 VDD1.n169 585
R661 VDD1.n172 VDD1.n171 585
R662 VDD1.n113 VDD1.n112 585
R663 VDD1.n179 VDD1.n178 585
R664 VDD1.n180 VDD1.n111 585
R665 VDD1.n182 VDD1.n181 585
R666 VDD1.n109 VDD1.n108 585
R667 VDD1.n188 VDD1.n187 585
R668 VDD1.n190 VDD1.n189 585
R669 VDD1.n105 VDD1.n104 585
R670 VDD1.n196 VDD1.n195 585
R671 VDD1.n198 VDD1.n197 585
R672 VDD1.n34 VDD1.t1 327.466
R673 VDD1.n134 VDD1.t0 327.466
R674 VDD1.n96 VDD1.n95 171.744
R675 VDD1.n95 VDD1.n3 171.744
R676 VDD1.n88 VDD1.n3 171.744
R677 VDD1.n88 VDD1.n87 171.744
R678 VDD1.n87 VDD1.n7 171.744
R679 VDD1.n80 VDD1.n7 171.744
R680 VDD1.n80 VDD1.n79 171.744
R681 VDD1.n79 VDD1.n78 171.744
R682 VDD1.n78 VDD1.n11 171.744
R683 VDD1.n71 VDD1.n11 171.744
R684 VDD1.n71 VDD1.n70 171.744
R685 VDD1.n70 VDD1.n16 171.744
R686 VDD1.n63 VDD1.n16 171.744
R687 VDD1.n63 VDD1.n62 171.744
R688 VDD1.n62 VDD1.n20 171.744
R689 VDD1.n55 VDD1.n20 171.744
R690 VDD1.n55 VDD1.n54 171.744
R691 VDD1.n54 VDD1.n24 171.744
R692 VDD1.n47 VDD1.n24 171.744
R693 VDD1.n47 VDD1.n46 171.744
R694 VDD1.n46 VDD1.n28 171.744
R695 VDD1.n39 VDD1.n28 171.744
R696 VDD1.n39 VDD1.n38 171.744
R697 VDD1.n38 VDD1.n32 171.744
R698 VDD1.n138 VDD1.n132 171.744
R699 VDD1.n139 VDD1.n138 171.744
R700 VDD1.n139 VDD1.n128 171.744
R701 VDD1.n146 VDD1.n128 171.744
R702 VDD1.n147 VDD1.n146 171.744
R703 VDD1.n147 VDD1.n124 171.744
R704 VDD1.n154 VDD1.n124 171.744
R705 VDD1.n155 VDD1.n154 171.744
R706 VDD1.n155 VDD1.n120 171.744
R707 VDD1.n162 VDD1.n120 171.744
R708 VDD1.n163 VDD1.n162 171.744
R709 VDD1.n163 VDD1.n116 171.744
R710 VDD1.n170 VDD1.n116 171.744
R711 VDD1.n171 VDD1.n170 171.744
R712 VDD1.n171 VDD1.n112 171.744
R713 VDD1.n179 VDD1.n112 171.744
R714 VDD1.n180 VDD1.n179 171.744
R715 VDD1.n181 VDD1.n180 171.744
R716 VDD1.n181 VDD1.n108 171.744
R717 VDD1.n188 VDD1.n108 171.744
R718 VDD1.n189 VDD1.n188 171.744
R719 VDD1.n189 VDD1.n104 171.744
R720 VDD1.n196 VDD1.n104 171.744
R721 VDD1.n197 VDD1.n196 171.744
R722 VDD1 VDD1.n201 93.7641
R723 VDD1.t1 VDD1.n32 85.8723
R724 VDD1.t0 VDD1.n132 85.8723
R725 VDD1 VDD1.n100 48.4483
R726 VDD1.n34 VDD1.n33 16.3895
R727 VDD1.n134 VDD1.n133 16.3895
R728 VDD1.n81 VDD1.n10 13.1884
R729 VDD1.n182 VDD1.n111 13.1884
R730 VDD1.n82 VDD1.n8 12.8005
R731 VDD1.n77 VDD1.n12 12.8005
R732 VDD1.n37 VDD1.n36 12.8005
R733 VDD1.n137 VDD1.n136 12.8005
R734 VDD1.n178 VDD1.n177 12.8005
R735 VDD1.n183 VDD1.n109 12.8005
R736 VDD1.n86 VDD1.n85 12.0247
R737 VDD1.n76 VDD1.n13 12.0247
R738 VDD1.n40 VDD1.n31 12.0247
R739 VDD1.n140 VDD1.n131 12.0247
R740 VDD1.n176 VDD1.n113 12.0247
R741 VDD1.n187 VDD1.n186 12.0247
R742 VDD1.n89 VDD1.n6 11.249
R743 VDD1.n73 VDD1.n72 11.249
R744 VDD1.n41 VDD1.n29 11.249
R745 VDD1.n141 VDD1.n129 11.249
R746 VDD1.n173 VDD1.n172 11.249
R747 VDD1.n190 VDD1.n107 11.249
R748 VDD1.n90 VDD1.n4 10.4732
R749 VDD1.n69 VDD1.n15 10.4732
R750 VDD1.n45 VDD1.n44 10.4732
R751 VDD1.n145 VDD1.n144 10.4732
R752 VDD1.n169 VDD1.n115 10.4732
R753 VDD1.n191 VDD1.n105 10.4732
R754 VDD1.n94 VDD1.n93 9.69747
R755 VDD1.n68 VDD1.n17 9.69747
R756 VDD1.n48 VDD1.n27 9.69747
R757 VDD1.n148 VDD1.n127 9.69747
R758 VDD1.n168 VDD1.n117 9.69747
R759 VDD1.n195 VDD1.n194 9.69747
R760 VDD1.n100 VDD1.n99 9.45567
R761 VDD1.n201 VDD1.n200 9.45567
R762 VDD1.n60 VDD1.n59 9.3005
R763 VDD1.n19 VDD1.n18 9.3005
R764 VDD1.n66 VDD1.n65 9.3005
R765 VDD1.n68 VDD1.n67 9.3005
R766 VDD1.n15 VDD1.n14 9.3005
R767 VDD1.n74 VDD1.n73 9.3005
R768 VDD1.n76 VDD1.n75 9.3005
R769 VDD1.n12 VDD1.n9 9.3005
R770 VDD1.n99 VDD1.n98 9.3005
R771 VDD1.n2 VDD1.n1 9.3005
R772 VDD1.n93 VDD1.n92 9.3005
R773 VDD1.n91 VDD1.n90 9.3005
R774 VDD1.n6 VDD1.n5 9.3005
R775 VDD1.n85 VDD1.n84 9.3005
R776 VDD1.n83 VDD1.n82 9.3005
R777 VDD1.n58 VDD1.n57 9.3005
R778 VDD1.n23 VDD1.n22 9.3005
R779 VDD1.n52 VDD1.n51 9.3005
R780 VDD1.n50 VDD1.n49 9.3005
R781 VDD1.n27 VDD1.n26 9.3005
R782 VDD1.n44 VDD1.n43 9.3005
R783 VDD1.n42 VDD1.n41 9.3005
R784 VDD1.n31 VDD1.n30 9.3005
R785 VDD1.n36 VDD1.n35 9.3005
R786 VDD1.n200 VDD1.n199 9.3005
R787 VDD1.n103 VDD1.n102 9.3005
R788 VDD1.n194 VDD1.n193 9.3005
R789 VDD1.n192 VDD1.n191 9.3005
R790 VDD1.n107 VDD1.n106 9.3005
R791 VDD1.n186 VDD1.n185 9.3005
R792 VDD1.n184 VDD1.n183 9.3005
R793 VDD1.n123 VDD1.n122 9.3005
R794 VDD1.n152 VDD1.n151 9.3005
R795 VDD1.n150 VDD1.n149 9.3005
R796 VDD1.n127 VDD1.n126 9.3005
R797 VDD1.n144 VDD1.n143 9.3005
R798 VDD1.n142 VDD1.n141 9.3005
R799 VDD1.n131 VDD1.n130 9.3005
R800 VDD1.n136 VDD1.n135 9.3005
R801 VDD1.n158 VDD1.n157 9.3005
R802 VDD1.n160 VDD1.n159 9.3005
R803 VDD1.n119 VDD1.n118 9.3005
R804 VDD1.n166 VDD1.n165 9.3005
R805 VDD1.n168 VDD1.n167 9.3005
R806 VDD1.n115 VDD1.n114 9.3005
R807 VDD1.n174 VDD1.n173 9.3005
R808 VDD1.n176 VDD1.n175 9.3005
R809 VDD1.n177 VDD1.n110 9.3005
R810 VDD1.n97 VDD1.n2 8.92171
R811 VDD1.n65 VDD1.n64 8.92171
R812 VDD1.n49 VDD1.n25 8.92171
R813 VDD1.n149 VDD1.n125 8.92171
R814 VDD1.n165 VDD1.n164 8.92171
R815 VDD1.n198 VDD1.n103 8.92171
R816 VDD1.n98 VDD1.n0 8.14595
R817 VDD1.n61 VDD1.n19 8.14595
R818 VDD1.n53 VDD1.n52 8.14595
R819 VDD1.n153 VDD1.n152 8.14595
R820 VDD1.n161 VDD1.n119 8.14595
R821 VDD1.n199 VDD1.n101 8.14595
R822 VDD1.n60 VDD1.n21 7.3702
R823 VDD1.n56 VDD1.n23 7.3702
R824 VDD1.n156 VDD1.n123 7.3702
R825 VDD1.n160 VDD1.n121 7.3702
R826 VDD1.n57 VDD1.n21 6.59444
R827 VDD1.n57 VDD1.n56 6.59444
R828 VDD1.n157 VDD1.n156 6.59444
R829 VDD1.n157 VDD1.n121 6.59444
R830 VDD1.n100 VDD1.n0 5.81868
R831 VDD1.n61 VDD1.n60 5.81868
R832 VDD1.n53 VDD1.n23 5.81868
R833 VDD1.n153 VDD1.n123 5.81868
R834 VDD1.n161 VDD1.n160 5.81868
R835 VDD1.n201 VDD1.n101 5.81868
R836 VDD1.n98 VDD1.n97 5.04292
R837 VDD1.n64 VDD1.n19 5.04292
R838 VDD1.n52 VDD1.n25 5.04292
R839 VDD1.n152 VDD1.n125 5.04292
R840 VDD1.n164 VDD1.n119 5.04292
R841 VDD1.n199 VDD1.n198 5.04292
R842 VDD1.n94 VDD1.n2 4.26717
R843 VDD1.n65 VDD1.n17 4.26717
R844 VDD1.n49 VDD1.n48 4.26717
R845 VDD1.n149 VDD1.n148 4.26717
R846 VDD1.n165 VDD1.n117 4.26717
R847 VDD1.n195 VDD1.n103 4.26717
R848 VDD1.n35 VDD1.n34 3.70982
R849 VDD1.n135 VDD1.n134 3.70982
R850 VDD1.n93 VDD1.n4 3.49141
R851 VDD1.n69 VDD1.n68 3.49141
R852 VDD1.n45 VDD1.n27 3.49141
R853 VDD1.n145 VDD1.n127 3.49141
R854 VDD1.n169 VDD1.n168 3.49141
R855 VDD1.n194 VDD1.n105 3.49141
R856 VDD1.n90 VDD1.n89 2.71565
R857 VDD1.n72 VDD1.n15 2.71565
R858 VDD1.n44 VDD1.n29 2.71565
R859 VDD1.n144 VDD1.n129 2.71565
R860 VDD1.n172 VDD1.n115 2.71565
R861 VDD1.n191 VDD1.n190 2.71565
R862 VDD1.n86 VDD1.n6 1.93989
R863 VDD1.n73 VDD1.n13 1.93989
R864 VDD1.n41 VDD1.n40 1.93989
R865 VDD1.n141 VDD1.n140 1.93989
R866 VDD1.n173 VDD1.n113 1.93989
R867 VDD1.n187 VDD1.n107 1.93989
R868 VDD1.n85 VDD1.n8 1.16414
R869 VDD1.n77 VDD1.n76 1.16414
R870 VDD1.n37 VDD1.n31 1.16414
R871 VDD1.n137 VDD1.n131 1.16414
R872 VDD1.n178 VDD1.n176 1.16414
R873 VDD1.n186 VDD1.n109 1.16414
R874 VDD1.n82 VDD1.n81 0.388379
R875 VDD1.n12 VDD1.n10 0.388379
R876 VDD1.n36 VDD1.n33 0.388379
R877 VDD1.n136 VDD1.n133 0.388379
R878 VDD1.n177 VDD1.n111 0.388379
R879 VDD1.n183 VDD1.n182 0.388379
R880 VDD1.n99 VDD1.n1 0.155672
R881 VDD1.n92 VDD1.n1 0.155672
R882 VDD1.n92 VDD1.n91 0.155672
R883 VDD1.n91 VDD1.n5 0.155672
R884 VDD1.n84 VDD1.n5 0.155672
R885 VDD1.n84 VDD1.n83 0.155672
R886 VDD1.n83 VDD1.n9 0.155672
R887 VDD1.n75 VDD1.n9 0.155672
R888 VDD1.n75 VDD1.n74 0.155672
R889 VDD1.n74 VDD1.n14 0.155672
R890 VDD1.n67 VDD1.n14 0.155672
R891 VDD1.n67 VDD1.n66 0.155672
R892 VDD1.n66 VDD1.n18 0.155672
R893 VDD1.n59 VDD1.n18 0.155672
R894 VDD1.n59 VDD1.n58 0.155672
R895 VDD1.n58 VDD1.n22 0.155672
R896 VDD1.n51 VDD1.n22 0.155672
R897 VDD1.n51 VDD1.n50 0.155672
R898 VDD1.n50 VDD1.n26 0.155672
R899 VDD1.n43 VDD1.n26 0.155672
R900 VDD1.n43 VDD1.n42 0.155672
R901 VDD1.n42 VDD1.n30 0.155672
R902 VDD1.n35 VDD1.n30 0.155672
R903 VDD1.n135 VDD1.n130 0.155672
R904 VDD1.n142 VDD1.n130 0.155672
R905 VDD1.n143 VDD1.n142 0.155672
R906 VDD1.n143 VDD1.n126 0.155672
R907 VDD1.n150 VDD1.n126 0.155672
R908 VDD1.n151 VDD1.n150 0.155672
R909 VDD1.n151 VDD1.n122 0.155672
R910 VDD1.n158 VDD1.n122 0.155672
R911 VDD1.n159 VDD1.n158 0.155672
R912 VDD1.n159 VDD1.n118 0.155672
R913 VDD1.n166 VDD1.n118 0.155672
R914 VDD1.n167 VDD1.n166 0.155672
R915 VDD1.n167 VDD1.n114 0.155672
R916 VDD1.n174 VDD1.n114 0.155672
R917 VDD1.n175 VDD1.n174 0.155672
R918 VDD1.n175 VDD1.n110 0.155672
R919 VDD1.n184 VDD1.n110 0.155672
R920 VDD1.n185 VDD1.n184 0.155672
R921 VDD1.n185 VDD1.n106 0.155672
R922 VDD1.n192 VDD1.n106 0.155672
R923 VDD1.n193 VDD1.n192 0.155672
R924 VDD1.n193 VDD1.n102 0.155672
R925 VDD1.n200 VDD1.n102 0.155672
R926 VN VN.t0 243.856
R927 VN VN.t1 194.231
R928 VDD2.n197 VDD2.n101 756.745
R929 VDD2.n96 VDD2.n0 756.745
R930 VDD2.n198 VDD2.n197 585
R931 VDD2.n196 VDD2.n195 585
R932 VDD2.n105 VDD2.n104 585
R933 VDD2.n190 VDD2.n189 585
R934 VDD2.n188 VDD2.n187 585
R935 VDD2.n109 VDD2.n108 585
R936 VDD2.n182 VDD2.n181 585
R937 VDD2.n180 VDD2.n111 585
R938 VDD2.n179 VDD2.n178 585
R939 VDD2.n114 VDD2.n112 585
R940 VDD2.n173 VDD2.n172 585
R941 VDD2.n171 VDD2.n170 585
R942 VDD2.n118 VDD2.n117 585
R943 VDD2.n165 VDD2.n164 585
R944 VDD2.n163 VDD2.n162 585
R945 VDD2.n122 VDD2.n121 585
R946 VDD2.n157 VDD2.n156 585
R947 VDD2.n155 VDD2.n154 585
R948 VDD2.n126 VDD2.n125 585
R949 VDD2.n149 VDD2.n148 585
R950 VDD2.n147 VDD2.n146 585
R951 VDD2.n130 VDD2.n129 585
R952 VDD2.n141 VDD2.n140 585
R953 VDD2.n139 VDD2.n138 585
R954 VDD2.n134 VDD2.n133 585
R955 VDD2.n32 VDD2.n31 585
R956 VDD2.n37 VDD2.n36 585
R957 VDD2.n39 VDD2.n38 585
R958 VDD2.n28 VDD2.n27 585
R959 VDD2.n45 VDD2.n44 585
R960 VDD2.n47 VDD2.n46 585
R961 VDD2.n24 VDD2.n23 585
R962 VDD2.n53 VDD2.n52 585
R963 VDD2.n55 VDD2.n54 585
R964 VDD2.n20 VDD2.n19 585
R965 VDD2.n61 VDD2.n60 585
R966 VDD2.n63 VDD2.n62 585
R967 VDD2.n16 VDD2.n15 585
R968 VDD2.n69 VDD2.n68 585
R969 VDD2.n71 VDD2.n70 585
R970 VDD2.n12 VDD2.n11 585
R971 VDD2.n78 VDD2.n77 585
R972 VDD2.n79 VDD2.n10 585
R973 VDD2.n81 VDD2.n80 585
R974 VDD2.n8 VDD2.n7 585
R975 VDD2.n87 VDD2.n86 585
R976 VDD2.n89 VDD2.n88 585
R977 VDD2.n4 VDD2.n3 585
R978 VDD2.n95 VDD2.n94 585
R979 VDD2.n97 VDD2.n96 585
R980 VDD2.n135 VDD2.t1 327.466
R981 VDD2.n33 VDD2.t0 327.466
R982 VDD2.n197 VDD2.n196 171.744
R983 VDD2.n196 VDD2.n104 171.744
R984 VDD2.n189 VDD2.n104 171.744
R985 VDD2.n189 VDD2.n188 171.744
R986 VDD2.n188 VDD2.n108 171.744
R987 VDD2.n181 VDD2.n108 171.744
R988 VDD2.n181 VDD2.n180 171.744
R989 VDD2.n180 VDD2.n179 171.744
R990 VDD2.n179 VDD2.n112 171.744
R991 VDD2.n172 VDD2.n112 171.744
R992 VDD2.n172 VDD2.n171 171.744
R993 VDD2.n171 VDD2.n117 171.744
R994 VDD2.n164 VDD2.n117 171.744
R995 VDD2.n164 VDD2.n163 171.744
R996 VDD2.n163 VDD2.n121 171.744
R997 VDD2.n156 VDD2.n121 171.744
R998 VDD2.n156 VDD2.n155 171.744
R999 VDD2.n155 VDD2.n125 171.744
R1000 VDD2.n148 VDD2.n125 171.744
R1001 VDD2.n148 VDD2.n147 171.744
R1002 VDD2.n147 VDD2.n129 171.744
R1003 VDD2.n140 VDD2.n129 171.744
R1004 VDD2.n140 VDD2.n139 171.744
R1005 VDD2.n139 VDD2.n133 171.744
R1006 VDD2.n37 VDD2.n31 171.744
R1007 VDD2.n38 VDD2.n37 171.744
R1008 VDD2.n38 VDD2.n27 171.744
R1009 VDD2.n45 VDD2.n27 171.744
R1010 VDD2.n46 VDD2.n45 171.744
R1011 VDD2.n46 VDD2.n23 171.744
R1012 VDD2.n53 VDD2.n23 171.744
R1013 VDD2.n54 VDD2.n53 171.744
R1014 VDD2.n54 VDD2.n19 171.744
R1015 VDD2.n61 VDD2.n19 171.744
R1016 VDD2.n62 VDD2.n61 171.744
R1017 VDD2.n62 VDD2.n15 171.744
R1018 VDD2.n69 VDD2.n15 171.744
R1019 VDD2.n70 VDD2.n69 171.744
R1020 VDD2.n70 VDD2.n11 171.744
R1021 VDD2.n78 VDD2.n11 171.744
R1022 VDD2.n79 VDD2.n78 171.744
R1023 VDD2.n80 VDD2.n79 171.744
R1024 VDD2.n80 VDD2.n7 171.744
R1025 VDD2.n87 VDD2.n7 171.744
R1026 VDD2.n88 VDD2.n87 171.744
R1027 VDD2.n88 VDD2.n3 171.744
R1028 VDD2.n95 VDD2.n3 171.744
R1029 VDD2.n96 VDD2.n95 171.744
R1030 VDD2.n202 VDD2.n100 92.5496
R1031 VDD2.t1 VDD2.n133 85.8723
R1032 VDD2.t0 VDD2.n31 85.8723
R1033 VDD2.n202 VDD2.n201 47.7005
R1034 VDD2.n135 VDD2.n134 16.3895
R1035 VDD2.n33 VDD2.n32 16.3895
R1036 VDD2.n182 VDD2.n111 13.1884
R1037 VDD2.n81 VDD2.n10 13.1884
R1038 VDD2.n183 VDD2.n109 12.8005
R1039 VDD2.n178 VDD2.n113 12.8005
R1040 VDD2.n138 VDD2.n137 12.8005
R1041 VDD2.n36 VDD2.n35 12.8005
R1042 VDD2.n77 VDD2.n76 12.8005
R1043 VDD2.n82 VDD2.n8 12.8005
R1044 VDD2.n187 VDD2.n186 12.0247
R1045 VDD2.n177 VDD2.n114 12.0247
R1046 VDD2.n141 VDD2.n132 12.0247
R1047 VDD2.n39 VDD2.n30 12.0247
R1048 VDD2.n75 VDD2.n12 12.0247
R1049 VDD2.n86 VDD2.n85 12.0247
R1050 VDD2.n190 VDD2.n107 11.249
R1051 VDD2.n174 VDD2.n173 11.249
R1052 VDD2.n142 VDD2.n130 11.249
R1053 VDD2.n40 VDD2.n28 11.249
R1054 VDD2.n72 VDD2.n71 11.249
R1055 VDD2.n89 VDD2.n6 11.249
R1056 VDD2.n191 VDD2.n105 10.4732
R1057 VDD2.n170 VDD2.n116 10.4732
R1058 VDD2.n146 VDD2.n145 10.4732
R1059 VDD2.n44 VDD2.n43 10.4732
R1060 VDD2.n68 VDD2.n14 10.4732
R1061 VDD2.n90 VDD2.n4 10.4732
R1062 VDD2.n195 VDD2.n194 9.69747
R1063 VDD2.n169 VDD2.n118 9.69747
R1064 VDD2.n149 VDD2.n128 9.69747
R1065 VDD2.n47 VDD2.n26 9.69747
R1066 VDD2.n67 VDD2.n16 9.69747
R1067 VDD2.n94 VDD2.n93 9.69747
R1068 VDD2.n201 VDD2.n200 9.45567
R1069 VDD2.n100 VDD2.n99 9.45567
R1070 VDD2.n161 VDD2.n160 9.3005
R1071 VDD2.n120 VDD2.n119 9.3005
R1072 VDD2.n167 VDD2.n166 9.3005
R1073 VDD2.n169 VDD2.n168 9.3005
R1074 VDD2.n116 VDD2.n115 9.3005
R1075 VDD2.n175 VDD2.n174 9.3005
R1076 VDD2.n177 VDD2.n176 9.3005
R1077 VDD2.n113 VDD2.n110 9.3005
R1078 VDD2.n200 VDD2.n199 9.3005
R1079 VDD2.n103 VDD2.n102 9.3005
R1080 VDD2.n194 VDD2.n193 9.3005
R1081 VDD2.n192 VDD2.n191 9.3005
R1082 VDD2.n107 VDD2.n106 9.3005
R1083 VDD2.n186 VDD2.n185 9.3005
R1084 VDD2.n184 VDD2.n183 9.3005
R1085 VDD2.n159 VDD2.n158 9.3005
R1086 VDD2.n124 VDD2.n123 9.3005
R1087 VDD2.n153 VDD2.n152 9.3005
R1088 VDD2.n151 VDD2.n150 9.3005
R1089 VDD2.n128 VDD2.n127 9.3005
R1090 VDD2.n145 VDD2.n144 9.3005
R1091 VDD2.n143 VDD2.n142 9.3005
R1092 VDD2.n132 VDD2.n131 9.3005
R1093 VDD2.n137 VDD2.n136 9.3005
R1094 VDD2.n99 VDD2.n98 9.3005
R1095 VDD2.n2 VDD2.n1 9.3005
R1096 VDD2.n93 VDD2.n92 9.3005
R1097 VDD2.n91 VDD2.n90 9.3005
R1098 VDD2.n6 VDD2.n5 9.3005
R1099 VDD2.n85 VDD2.n84 9.3005
R1100 VDD2.n83 VDD2.n82 9.3005
R1101 VDD2.n22 VDD2.n21 9.3005
R1102 VDD2.n51 VDD2.n50 9.3005
R1103 VDD2.n49 VDD2.n48 9.3005
R1104 VDD2.n26 VDD2.n25 9.3005
R1105 VDD2.n43 VDD2.n42 9.3005
R1106 VDD2.n41 VDD2.n40 9.3005
R1107 VDD2.n30 VDD2.n29 9.3005
R1108 VDD2.n35 VDD2.n34 9.3005
R1109 VDD2.n57 VDD2.n56 9.3005
R1110 VDD2.n59 VDD2.n58 9.3005
R1111 VDD2.n18 VDD2.n17 9.3005
R1112 VDD2.n65 VDD2.n64 9.3005
R1113 VDD2.n67 VDD2.n66 9.3005
R1114 VDD2.n14 VDD2.n13 9.3005
R1115 VDD2.n73 VDD2.n72 9.3005
R1116 VDD2.n75 VDD2.n74 9.3005
R1117 VDD2.n76 VDD2.n9 9.3005
R1118 VDD2.n198 VDD2.n103 8.92171
R1119 VDD2.n166 VDD2.n165 8.92171
R1120 VDD2.n150 VDD2.n126 8.92171
R1121 VDD2.n48 VDD2.n24 8.92171
R1122 VDD2.n64 VDD2.n63 8.92171
R1123 VDD2.n97 VDD2.n2 8.92171
R1124 VDD2.n199 VDD2.n101 8.14595
R1125 VDD2.n162 VDD2.n120 8.14595
R1126 VDD2.n154 VDD2.n153 8.14595
R1127 VDD2.n52 VDD2.n51 8.14595
R1128 VDD2.n60 VDD2.n18 8.14595
R1129 VDD2.n98 VDD2.n0 8.14595
R1130 VDD2.n161 VDD2.n122 7.3702
R1131 VDD2.n157 VDD2.n124 7.3702
R1132 VDD2.n55 VDD2.n22 7.3702
R1133 VDD2.n59 VDD2.n20 7.3702
R1134 VDD2.n158 VDD2.n122 6.59444
R1135 VDD2.n158 VDD2.n157 6.59444
R1136 VDD2.n56 VDD2.n55 6.59444
R1137 VDD2.n56 VDD2.n20 6.59444
R1138 VDD2.n201 VDD2.n101 5.81868
R1139 VDD2.n162 VDD2.n161 5.81868
R1140 VDD2.n154 VDD2.n124 5.81868
R1141 VDD2.n52 VDD2.n22 5.81868
R1142 VDD2.n60 VDD2.n59 5.81868
R1143 VDD2.n100 VDD2.n0 5.81868
R1144 VDD2.n199 VDD2.n198 5.04292
R1145 VDD2.n165 VDD2.n120 5.04292
R1146 VDD2.n153 VDD2.n126 5.04292
R1147 VDD2.n51 VDD2.n24 5.04292
R1148 VDD2.n63 VDD2.n18 5.04292
R1149 VDD2.n98 VDD2.n97 5.04292
R1150 VDD2.n195 VDD2.n103 4.26717
R1151 VDD2.n166 VDD2.n118 4.26717
R1152 VDD2.n150 VDD2.n149 4.26717
R1153 VDD2.n48 VDD2.n47 4.26717
R1154 VDD2.n64 VDD2.n16 4.26717
R1155 VDD2.n94 VDD2.n2 4.26717
R1156 VDD2.n136 VDD2.n135 3.70982
R1157 VDD2.n34 VDD2.n33 3.70982
R1158 VDD2.n194 VDD2.n105 3.49141
R1159 VDD2.n170 VDD2.n169 3.49141
R1160 VDD2.n146 VDD2.n128 3.49141
R1161 VDD2.n44 VDD2.n26 3.49141
R1162 VDD2.n68 VDD2.n67 3.49141
R1163 VDD2.n93 VDD2.n4 3.49141
R1164 VDD2.n191 VDD2.n190 2.71565
R1165 VDD2.n173 VDD2.n116 2.71565
R1166 VDD2.n145 VDD2.n130 2.71565
R1167 VDD2.n43 VDD2.n28 2.71565
R1168 VDD2.n71 VDD2.n14 2.71565
R1169 VDD2.n90 VDD2.n89 2.71565
R1170 VDD2.n187 VDD2.n107 1.93989
R1171 VDD2.n174 VDD2.n114 1.93989
R1172 VDD2.n142 VDD2.n141 1.93989
R1173 VDD2.n40 VDD2.n39 1.93989
R1174 VDD2.n72 VDD2.n12 1.93989
R1175 VDD2.n86 VDD2.n6 1.93989
R1176 VDD2.n186 VDD2.n109 1.16414
R1177 VDD2.n178 VDD2.n177 1.16414
R1178 VDD2.n138 VDD2.n132 1.16414
R1179 VDD2.n36 VDD2.n30 1.16414
R1180 VDD2.n77 VDD2.n75 1.16414
R1181 VDD2.n85 VDD2.n8 1.16414
R1182 VDD2 VDD2.n202 0.748345
R1183 VDD2.n183 VDD2.n182 0.388379
R1184 VDD2.n113 VDD2.n111 0.388379
R1185 VDD2.n137 VDD2.n134 0.388379
R1186 VDD2.n35 VDD2.n32 0.388379
R1187 VDD2.n76 VDD2.n10 0.388379
R1188 VDD2.n82 VDD2.n81 0.388379
R1189 VDD2.n200 VDD2.n102 0.155672
R1190 VDD2.n193 VDD2.n102 0.155672
R1191 VDD2.n193 VDD2.n192 0.155672
R1192 VDD2.n192 VDD2.n106 0.155672
R1193 VDD2.n185 VDD2.n106 0.155672
R1194 VDD2.n185 VDD2.n184 0.155672
R1195 VDD2.n184 VDD2.n110 0.155672
R1196 VDD2.n176 VDD2.n110 0.155672
R1197 VDD2.n176 VDD2.n175 0.155672
R1198 VDD2.n175 VDD2.n115 0.155672
R1199 VDD2.n168 VDD2.n115 0.155672
R1200 VDD2.n168 VDD2.n167 0.155672
R1201 VDD2.n167 VDD2.n119 0.155672
R1202 VDD2.n160 VDD2.n119 0.155672
R1203 VDD2.n160 VDD2.n159 0.155672
R1204 VDD2.n159 VDD2.n123 0.155672
R1205 VDD2.n152 VDD2.n123 0.155672
R1206 VDD2.n152 VDD2.n151 0.155672
R1207 VDD2.n151 VDD2.n127 0.155672
R1208 VDD2.n144 VDD2.n127 0.155672
R1209 VDD2.n144 VDD2.n143 0.155672
R1210 VDD2.n143 VDD2.n131 0.155672
R1211 VDD2.n136 VDD2.n131 0.155672
R1212 VDD2.n34 VDD2.n29 0.155672
R1213 VDD2.n41 VDD2.n29 0.155672
R1214 VDD2.n42 VDD2.n41 0.155672
R1215 VDD2.n42 VDD2.n25 0.155672
R1216 VDD2.n49 VDD2.n25 0.155672
R1217 VDD2.n50 VDD2.n49 0.155672
R1218 VDD2.n50 VDD2.n21 0.155672
R1219 VDD2.n57 VDD2.n21 0.155672
R1220 VDD2.n58 VDD2.n57 0.155672
R1221 VDD2.n58 VDD2.n17 0.155672
R1222 VDD2.n65 VDD2.n17 0.155672
R1223 VDD2.n66 VDD2.n65 0.155672
R1224 VDD2.n66 VDD2.n13 0.155672
R1225 VDD2.n73 VDD2.n13 0.155672
R1226 VDD2.n74 VDD2.n73 0.155672
R1227 VDD2.n74 VDD2.n9 0.155672
R1228 VDD2.n83 VDD2.n9 0.155672
R1229 VDD2.n84 VDD2.n83 0.155672
R1230 VDD2.n84 VDD2.n5 0.155672
R1231 VDD2.n91 VDD2.n5 0.155672
R1232 VDD2.n92 VDD2.n91 0.155672
R1233 VDD2.n92 VDD2.n1 0.155672
R1234 VDD2.n99 VDD2.n1 0.155672
R1235 B.n511 B.n84 585
R1236 B.n513 B.n512 585
R1237 B.n514 B.n83 585
R1238 B.n516 B.n515 585
R1239 B.n517 B.n82 585
R1240 B.n519 B.n518 585
R1241 B.n520 B.n81 585
R1242 B.n522 B.n521 585
R1243 B.n523 B.n80 585
R1244 B.n525 B.n524 585
R1245 B.n526 B.n79 585
R1246 B.n528 B.n527 585
R1247 B.n529 B.n78 585
R1248 B.n531 B.n530 585
R1249 B.n532 B.n77 585
R1250 B.n534 B.n533 585
R1251 B.n535 B.n76 585
R1252 B.n537 B.n536 585
R1253 B.n538 B.n75 585
R1254 B.n540 B.n539 585
R1255 B.n541 B.n74 585
R1256 B.n543 B.n542 585
R1257 B.n544 B.n73 585
R1258 B.n546 B.n545 585
R1259 B.n547 B.n72 585
R1260 B.n549 B.n548 585
R1261 B.n550 B.n71 585
R1262 B.n552 B.n551 585
R1263 B.n553 B.n70 585
R1264 B.n555 B.n554 585
R1265 B.n556 B.n69 585
R1266 B.n558 B.n557 585
R1267 B.n559 B.n68 585
R1268 B.n561 B.n560 585
R1269 B.n562 B.n67 585
R1270 B.n564 B.n563 585
R1271 B.n565 B.n66 585
R1272 B.n567 B.n566 585
R1273 B.n568 B.n65 585
R1274 B.n570 B.n569 585
R1275 B.n571 B.n64 585
R1276 B.n573 B.n572 585
R1277 B.n574 B.n63 585
R1278 B.n576 B.n575 585
R1279 B.n577 B.n62 585
R1280 B.n579 B.n578 585
R1281 B.n580 B.n61 585
R1282 B.n582 B.n581 585
R1283 B.n583 B.n60 585
R1284 B.n585 B.n584 585
R1285 B.n586 B.n59 585
R1286 B.n588 B.n587 585
R1287 B.n589 B.n58 585
R1288 B.n591 B.n590 585
R1289 B.n592 B.n57 585
R1290 B.n594 B.n593 585
R1291 B.n595 B.n56 585
R1292 B.n597 B.n596 585
R1293 B.n598 B.n55 585
R1294 B.n600 B.n599 585
R1295 B.n602 B.n601 585
R1296 B.n603 B.n51 585
R1297 B.n605 B.n604 585
R1298 B.n606 B.n50 585
R1299 B.n608 B.n607 585
R1300 B.n609 B.n49 585
R1301 B.n611 B.n610 585
R1302 B.n612 B.n48 585
R1303 B.n614 B.n613 585
R1304 B.n616 B.n45 585
R1305 B.n618 B.n617 585
R1306 B.n619 B.n44 585
R1307 B.n621 B.n620 585
R1308 B.n622 B.n43 585
R1309 B.n624 B.n623 585
R1310 B.n625 B.n42 585
R1311 B.n627 B.n626 585
R1312 B.n628 B.n41 585
R1313 B.n630 B.n629 585
R1314 B.n631 B.n40 585
R1315 B.n633 B.n632 585
R1316 B.n634 B.n39 585
R1317 B.n636 B.n635 585
R1318 B.n637 B.n38 585
R1319 B.n639 B.n638 585
R1320 B.n640 B.n37 585
R1321 B.n642 B.n641 585
R1322 B.n643 B.n36 585
R1323 B.n645 B.n644 585
R1324 B.n646 B.n35 585
R1325 B.n648 B.n647 585
R1326 B.n649 B.n34 585
R1327 B.n651 B.n650 585
R1328 B.n652 B.n33 585
R1329 B.n654 B.n653 585
R1330 B.n655 B.n32 585
R1331 B.n657 B.n656 585
R1332 B.n658 B.n31 585
R1333 B.n660 B.n659 585
R1334 B.n661 B.n30 585
R1335 B.n663 B.n662 585
R1336 B.n664 B.n29 585
R1337 B.n666 B.n665 585
R1338 B.n667 B.n28 585
R1339 B.n669 B.n668 585
R1340 B.n670 B.n27 585
R1341 B.n672 B.n671 585
R1342 B.n673 B.n26 585
R1343 B.n675 B.n674 585
R1344 B.n676 B.n25 585
R1345 B.n678 B.n677 585
R1346 B.n679 B.n24 585
R1347 B.n681 B.n680 585
R1348 B.n682 B.n23 585
R1349 B.n684 B.n683 585
R1350 B.n685 B.n22 585
R1351 B.n687 B.n686 585
R1352 B.n688 B.n21 585
R1353 B.n690 B.n689 585
R1354 B.n691 B.n20 585
R1355 B.n693 B.n692 585
R1356 B.n694 B.n19 585
R1357 B.n696 B.n695 585
R1358 B.n697 B.n18 585
R1359 B.n699 B.n698 585
R1360 B.n700 B.n17 585
R1361 B.n702 B.n701 585
R1362 B.n703 B.n16 585
R1363 B.n705 B.n704 585
R1364 B.n510 B.n509 585
R1365 B.n508 B.n85 585
R1366 B.n507 B.n506 585
R1367 B.n505 B.n86 585
R1368 B.n504 B.n503 585
R1369 B.n502 B.n87 585
R1370 B.n501 B.n500 585
R1371 B.n499 B.n88 585
R1372 B.n498 B.n497 585
R1373 B.n496 B.n89 585
R1374 B.n495 B.n494 585
R1375 B.n493 B.n90 585
R1376 B.n492 B.n491 585
R1377 B.n490 B.n91 585
R1378 B.n489 B.n488 585
R1379 B.n487 B.n92 585
R1380 B.n486 B.n485 585
R1381 B.n484 B.n93 585
R1382 B.n483 B.n482 585
R1383 B.n481 B.n94 585
R1384 B.n480 B.n479 585
R1385 B.n478 B.n95 585
R1386 B.n477 B.n476 585
R1387 B.n475 B.n96 585
R1388 B.n474 B.n473 585
R1389 B.n472 B.n97 585
R1390 B.n471 B.n470 585
R1391 B.n469 B.n98 585
R1392 B.n468 B.n467 585
R1393 B.n466 B.n99 585
R1394 B.n465 B.n464 585
R1395 B.n463 B.n100 585
R1396 B.n462 B.n461 585
R1397 B.n460 B.n101 585
R1398 B.n459 B.n458 585
R1399 B.n457 B.n102 585
R1400 B.n456 B.n455 585
R1401 B.n454 B.n103 585
R1402 B.n453 B.n452 585
R1403 B.n451 B.n104 585
R1404 B.n450 B.n449 585
R1405 B.n448 B.n105 585
R1406 B.n447 B.n446 585
R1407 B.n445 B.n106 585
R1408 B.n444 B.n443 585
R1409 B.n442 B.n107 585
R1410 B.n441 B.n440 585
R1411 B.n439 B.n108 585
R1412 B.n438 B.n437 585
R1413 B.n436 B.n109 585
R1414 B.n435 B.n434 585
R1415 B.n433 B.n110 585
R1416 B.n432 B.n431 585
R1417 B.n430 B.n111 585
R1418 B.n429 B.n428 585
R1419 B.n234 B.n233 585
R1420 B.n235 B.n180 585
R1421 B.n237 B.n236 585
R1422 B.n238 B.n179 585
R1423 B.n240 B.n239 585
R1424 B.n241 B.n178 585
R1425 B.n243 B.n242 585
R1426 B.n244 B.n177 585
R1427 B.n246 B.n245 585
R1428 B.n247 B.n176 585
R1429 B.n249 B.n248 585
R1430 B.n250 B.n175 585
R1431 B.n252 B.n251 585
R1432 B.n253 B.n174 585
R1433 B.n255 B.n254 585
R1434 B.n256 B.n173 585
R1435 B.n258 B.n257 585
R1436 B.n259 B.n172 585
R1437 B.n261 B.n260 585
R1438 B.n262 B.n171 585
R1439 B.n264 B.n263 585
R1440 B.n265 B.n170 585
R1441 B.n267 B.n266 585
R1442 B.n268 B.n169 585
R1443 B.n270 B.n269 585
R1444 B.n271 B.n168 585
R1445 B.n273 B.n272 585
R1446 B.n274 B.n167 585
R1447 B.n276 B.n275 585
R1448 B.n277 B.n166 585
R1449 B.n279 B.n278 585
R1450 B.n280 B.n165 585
R1451 B.n282 B.n281 585
R1452 B.n283 B.n164 585
R1453 B.n285 B.n284 585
R1454 B.n286 B.n163 585
R1455 B.n288 B.n287 585
R1456 B.n289 B.n162 585
R1457 B.n291 B.n290 585
R1458 B.n292 B.n161 585
R1459 B.n294 B.n293 585
R1460 B.n295 B.n160 585
R1461 B.n297 B.n296 585
R1462 B.n298 B.n159 585
R1463 B.n300 B.n299 585
R1464 B.n301 B.n158 585
R1465 B.n303 B.n302 585
R1466 B.n304 B.n157 585
R1467 B.n306 B.n305 585
R1468 B.n307 B.n156 585
R1469 B.n309 B.n308 585
R1470 B.n310 B.n155 585
R1471 B.n312 B.n311 585
R1472 B.n313 B.n154 585
R1473 B.n315 B.n314 585
R1474 B.n316 B.n153 585
R1475 B.n318 B.n317 585
R1476 B.n319 B.n152 585
R1477 B.n321 B.n320 585
R1478 B.n322 B.n149 585
R1479 B.n325 B.n324 585
R1480 B.n326 B.n148 585
R1481 B.n328 B.n327 585
R1482 B.n329 B.n147 585
R1483 B.n331 B.n330 585
R1484 B.n332 B.n146 585
R1485 B.n334 B.n333 585
R1486 B.n335 B.n145 585
R1487 B.n337 B.n336 585
R1488 B.n339 B.n338 585
R1489 B.n340 B.n141 585
R1490 B.n342 B.n341 585
R1491 B.n343 B.n140 585
R1492 B.n345 B.n344 585
R1493 B.n346 B.n139 585
R1494 B.n348 B.n347 585
R1495 B.n349 B.n138 585
R1496 B.n351 B.n350 585
R1497 B.n352 B.n137 585
R1498 B.n354 B.n353 585
R1499 B.n355 B.n136 585
R1500 B.n357 B.n356 585
R1501 B.n358 B.n135 585
R1502 B.n360 B.n359 585
R1503 B.n361 B.n134 585
R1504 B.n363 B.n362 585
R1505 B.n364 B.n133 585
R1506 B.n366 B.n365 585
R1507 B.n367 B.n132 585
R1508 B.n369 B.n368 585
R1509 B.n370 B.n131 585
R1510 B.n372 B.n371 585
R1511 B.n373 B.n130 585
R1512 B.n375 B.n374 585
R1513 B.n376 B.n129 585
R1514 B.n378 B.n377 585
R1515 B.n379 B.n128 585
R1516 B.n381 B.n380 585
R1517 B.n382 B.n127 585
R1518 B.n384 B.n383 585
R1519 B.n385 B.n126 585
R1520 B.n387 B.n386 585
R1521 B.n388 B.n125 585
R1522 B.n390 B.n389 585
R1523 B.n391 B.n124 585
R1524 B.n393 B.n392 585
R1525 B.n394 B.n123 585
R1526 B.n396 B.n395 585
R1527 B.n397 B.n122 585
R1528 B.n399 B.n398 585
R1529 B.n400 B.n121 585
R1530 B.n402 B.n401 585
R1531 B.n403 B.n120 585
R1532 B.n405 B.n404 585
R1533 B.n406 B.n119 585
R1534 B.n408 B.n407 585
R1535 B.n409 B.n118 585
R1536 B.n411 B.n410 585
R1537 B.n412 B.n117 585
R1538 B.n414 B.n413 585
R1539 B.n415 B.n116 585
R1540 B.n417 B.n416 585
R1541 B.n418 B.n115 585
R1542 B.n420 B.n419 585
R1543 B.n421 B.n114 585
R1544 B.n423 B.n422 585
R1545 B.n424 B.n113 585
R1546 B.n426 B.n425 585
R1547 B.n427 B.n112 585
R1548 B.n232 B.n181 585
R1549 B.n231 B.n230 585
R1550 B.n229 B.n182 585
R1551 B.n228 B.n227 585
R1552 B.n226 B.n183 585
R1553 B.n225 B.n224 585
R1554 B.n223 B.n184 585
R1555 B.n222 B.n221 585
R1556 B.n220 B.n185 585
R1557 B.n219 B.n218 585
R1558 B.n217 B.n186 585
R1559 B.n216 B.n215 585
R1560 B.n214 B.n187 585
R1561 B.n213 B.n212 585
R1562 B.n211 B.n188 585
R1563 B.n210 B.n209 585
R1564 B.n208 B.n189 585
R1565 B.n207 B.n206 585
R1566 B.n205 B.n190 585
R1567 B.n204 B.n203 585
R1568 B.n202 B.n191 585
R1569 B.n201 B.n200 585
R1570 B.n199 B.n192 585
R1571 B.n198 B.n197 585
R1572 B.n196 B.n193 585
R1573 B.n195 B.n194 585
R1574 B.n2 B.n0 585
R1575 B.n745 B.n1 585
R1576 B.n744 B.n743 585
R1577 B.n742 B.n3 585
R1578 B.n741 B.n740 585
R1579 B.n739 B.n4 585
R1580 B.n738 B.n737 585
R1581 B.n736 B.n5 585
R1582 B.n735 B.n734 585
R1583 B.n733 B.n6 585
R1584 B.n732 B.n731 585
R1585 B.n730 B.n7 585
R1586 B.n729 B.n728 585
R1587 B.n727 B.n8 585
R1588 B.n726 B.n725 585
R1589 B.n724 B.n9 585
R1590 B.n723 B.n722 585
R1591 B.n721 B.n10 585
R1592 B.n720 B.n719 585
R1593 B.n718 B.n11 585
R1594 B.n717 B.n716 585
R1595 B.n715 B.n12 585
R1596 B.n714 B.n713 585
R1597 B.n712 B.n13 585
R1598 B.n711 B.n710 585
R1599 B.n709 B.n14 585
R1600 B.n708 B.n707 585
R1601 B.n706 B.n15 585
R1602 B.n747 B.n746 585
R1603 B.n142 B.t5 548.986
R1604 B.n52 B.t1 548.986
R1605 B.n150 B.t11 548.986
R1606 B.n46 B.t7 548.986
R1607 B.n234 B.n181 502.111
R1608 B.n704 B.n15 502.111
R1609 B.n428 B.n427 502.111
R1610 B.n511 B.n510 502.111
R1611 B.n143 B.t4 486.925
R1612 B.n53 B.t2 486.925
R1613 B.n151 B.t10 486.925
R1614 B.n47 B.t8 486.925
R1615 B.n142 B.t3 361.082
R1616 B.n150 B.t9 361.082
R1617 B.n46 B.t6 361.082
R1618 B.n52 B.t0 361.082
R1619 B.n230 B.n181 163.367
R1620 B.n230 B.n229 163.367
R1621 B.n229 B.n228 163.367
R1622 B.n228 B.n183 163.367
R1623 B.n224 B.n183 163.367
R1624 B.n224 B.n223 163.367
R1625 B.n223 B.n222 163.367
R1626 B.n222 B.n185 163.367
R1627 B.n218 B.n185 163.367
R1628 B.n218 B.n217 163.367
R1629 B.n217 B.n216 163.367
R1630 B.n216 B.n187 163.367
R1631 B.n212 B.n187 163.367
R1632 B.n212 B.n211 163.367
R1633 B.n211 B.n210 163.367
R1634 B.n210 B.n189 163.367
R1635 B.n206 B.n189 163.367
R1636 B.n206 B.n205 163.367
R1637 B.n205 B.n204 163.367
R1638 B.n204 B.n191 163.367
R1639 B.n200 B.n191 163.367
R1640 B.n200 B.n199 163.367
R1641 B.n199 B.n198 163.367
R1642 B.n198 B.n193 163.367
R1643 B.n194 B.n193 163.367
R1644 B.n194 B.n2 163.367
R1645 B.n746 B.n2 163.367
R1646 B.n746 B.n745 163.367
R1647 B.n745 B.n744 163.367
R1648 B.n744 B.n3 163.367
R1649 B.n740 B.n3 163.367
R1650 B.n740 B.n739 163.367
R1651 B.n739 B.n738 163.367
R1652 B.n738 B.n5 163.367
R1653 B.n734 B.n5 163.367
R1654 B.n734 B.n733 163.367
R1655 B.n733 B.n732 163.367
R1656 B.n732 B.n7 163.367
R1657 B.n728 B.n7 163.367
R1658 B.n728 B.n727 163.367
R1659 B.n727 B.n726 163.367
R1660 B.n726 B.n9 163.367
R1661 B.n722 B.n9 163.367
R1662 B.n722 B.n721 163.367
R1663 B.n721 B.n720 163.367
R1664 B.n720 B.n11 163.367
R1665 B.n716 B.n11 163.367
R1666 B.n716 B.n715 163.367
R1667 B.n715 B.n714 163.367
R1668 B.n714 B.n13 163.367
R1669 B.n710 B.n13 163.367
R1670 B.n710 B.n709 163.367
R1671 B.n709 B.n708 163.367
R1672 B.n708 B.n15 163.367
R1673 B.n235 B.n234 163.367
R1674 B.n236 B.n235 163.367
R1675 B.n236 B.n179 163.367
R1676 B.n240 B.n179 163.367
R1677 B.n241 B.n240 163.367
R1678 B.n242 B.n241 163.367
R1679 B.n242 B.n177 163.367
R1680 B.n246 B.n177 163.367
R1681 B.n247 B.n246 163.367
R1682 B.n248 B.n247 163.367
R1683 B.n248 B.n175 163.367
R1684 B.n252 B.n175 163.367
R1685 B.n253 B.n252 163.367
R1686 B.n254 B.n253 163.367
R1687 B.n254 B.n173 163.367
R1688 B.n258 B.n173 163.367
R1689 B.n259 B.n258 163.367
R1690 B.n260 B.n259 163.367
R1691 B.n260 B.n171 163.367
R1692 B.n264 B.n171 163.367
R1693 B.n265 B.n264 163.367
R1694 B.n266 B.n265 163.367
R1695 B.n266 B.n169 163.367
R1696 B.n270 B.n169 163.367
R1697 B.n271 B.n270 163.367
R1698 B.n272 B.n271 163.367
R1699 B.n272 B.n167 163.367
R1700 B.n276 B.n167 163.367
R1701 B.n277 B.n276 163.367
R1702 B.n278 B.n277 163.367
R1703 B.n278 B.n165 163.367
R1704 B.n282 B.n165 163.367
R1705 B.n283 B.n282 163.367
R1706 B.n284 B.n283 163.367
R1707 B.n284 B.n163 163.367
R1708 B.n288 B.n163 163.367
R1709 B.n289 B.n288 163.367
R1710 B.n290 B.n289 163.367
R1711 B.n290 B.n161 163.367
R1712 B.n294 B.n161 163.367
R1713 B.n295 B.n294 163.367
R1714 B.n296 B.n295 163.367
R1715 B.n296 B.n159 163.367
R1716 B.n300 B.n159 163.367
R1717 B.n301 B.n300 163.367
R1718 B.n302 B.n301 163.367
R1719 B.n302 B.n157 163.367
R1720 B.n306 B.n157 163.367
R1721 B.n307 B.n306 163.367
R1722 B.n308 B.n307 163.367
R1723 B.n308 B.n155 163.367
R1724 B.n312 B.n155 163.367
R1725 B.n313 B.n312 163.367
R1726 B.n314 B.n313 163.367
R1727 B.n314 B.n153 163.367
R1728 B.n318 B.n153 163.367
R1729 B.n319 B.n318 163.367
R1730 B.n320 B.n319 163.367
R1731 B.n320 B.n149 163.367
R1732 B.n325 B.n149 163.367
R1733 B.n326 B.n325 163.367
R1734 B.n327 B.n326 163.367
R1735 B.n327 B.n147 163.367
R1736 B.n331 B.n147 163.367
R1737 B.n332 B.n331 163.367
R1738 B.n333 B.n332 163.367
R1739 B.n333 B.n145 163.367
R1740 B.n337 B.n145 163.367
R1741 B.n338 B.n337 163.367
R1742 B.n338 B.n141 163.367
R1743 B.n342 B.n141 163.367
R1744 B.n343 B.n342 163.367
R1745 B.n344 B.n343 163.367
R1746 B.n344 B.n139 163.367
R1747 B.n348 B.n139 163.367
R1748 B.n349 B.n348 163.367
R1749 B.n350 B.n349 163.367
R1750 B.n350 B.n137 163.367
R1751 B.n354 B.n137 163.367
R1752 B.n355 B.n354 163.367
R1753 B.n356 B.n355 163.367
R1754 B.n356 B.n135 163.367
R1755 B.n360 B.n135 163.367
R1756 B.n361 B.n360 163.367
R1757 B.n362 B.n361 163.367
R1758 B.n362 B.n133 163.367
R1759 B.n366 B.n133 163.367
R1760 B.n367 B.n366 163.367
R1761 B.n368 B.n367 163.367
R1762 B.n368 B.n131 163.367
R1763 B.n372 B.n131 163.367
R1764 B.n373 B.n372 163.367
R1765 B.n374 B.n373 163.367
R1766 B.n374 B.n129 163.367
R1767 B.n378 B.n129 163.367
R1768 B.n379 B.n378 163.367
R1769 B.n380 B.n379 163.367
R1770 B.n380 B.n127 163.367
R1771 B.n384 B.n127 163.367
R1772 B.n385 B.n384 163.367
R1773 B.n386 B.n385 163.367
R1774 B.n386 B.n125 163.367
R1775 B.n390 B.n125 163.367
R1776 B.n391 B.n390 163.367
R1777 B.n392 B.n391 163.367
R1778 B.n392 B.n123 163.367
R1779 B.n396 B.n123 163.367
R1780 B.n397 B.n396 163.367
R1781 B.n398 B.n397 163.367
R1782 B.n398 B.n121 163.367
R1783 B.n402 B.n121 163.367
R1784 B.n403 B.n402 163.367
R1785 B.n404 B.n403 163.367
R1786 B.n404 B.n119 163.367
R1787 B.n408 B.n119 163.367
R1788 B.n409 B.n408 163.367
R1789 B.n410 B.n409 163.367
R1790 B.n410 B.n117 163.367
R1791 B.n414 B.n117 163.367
R1792 B.n415 B.n414 163.367
R1793 B.n416 B.n415 163.367
R1794 B.n416 B.n115 163.367
R1795 B.n420 B.n115 163.367
R1796 B.n421 B.n420 163.367
R1797 B.n422 B.n421 163.367
R1798 B.n422 B.n113 163.367
R1799 B.n426 B.n113 163.367
R1800 B.n427 B.n426 163.367
R1801 B.n428 B.n111 163.367
R1802 B.n432 B.n111 163.367
R1803 B.n433 B.n432 163.367
R1804 B.n434 B.n433 163.367
R1805 B.n434 B.n109 163.367
R1806 B.n438 B.n109 163.367
R1807 B.n439 B.n438 163.367
R1808 B.n440 B.n439 163.367
R1809 B.n440 B.n107 163.367
R1810 B.n444 B.n107 163.367
R1811 B.n445 B.n444 163.367
R1812 B.n446 B.n445 163.367
R1813 B.n446 B.n105 163.367
R1814 B.n450 B.n105 163.367
R1815 B.n451 B.n450 163.367
R1816 B.n452 B.n451 163.367
R1817 B.n452 B.n103 163.367
R1818 B.n456 B.n103 163.367
R1819 B.n457 B.n456 163.367
R1820 B.n458 B.n457 163.367
R1821 B.n458 B.n101 163.367
R1822 B.n462 B.n101 163.367
R1823 B.n463 B.n462 163.367
R1824 B.n464 B.n463 163.367
R1825 B.n464 B.n99 163.367
R1826 B.n468 B.n99 163.367
R1827 B.n469 B.n468 163.367
R1828 B.n470 B.n469 163.367
R1829 B.n470 B.n97 163.367
R1830 B.n474 B.n97 163.367
R1831 B.n475 B.n474 163.367
R1832 B.n476 B.n475 163.367
R1833 B.n476 B.n95 163.367
R1834 B.n480 B.n95 163.367
R1835 B.n481 B.n480 163.367
R1836 B.n482 B.n481 163.367
R1837 B.n482 B.n93 163.367
R1838 B.n486 B.n93 163.367
R1839 B.n487 B.n486 163.367
R1840 B.n488 B.n487 163.367
R1841 B.n488 B.n91 163.367
R1842 B.n492 B.n91 163.367
R1843 B.n493 B.n492 163.367
R1844 B.n494 B.n493 163.367
R1845 B.n494 B.n89 163.367
R1846 B.n498 B.n89 163.367
R1847 B.n499 B.n498 163.367
R1848 B.n500 B.n499 163.367
R1849 B.n500 B.n87 163.367
R1850 B.n504 B.n87 163.367
R1851 B.n505 B.n504 163.367
R1852 B.n506 B.n505 163.367
R1853 B.n506 B.n85 163.367
R1854 B.n510 B.n85 163.367
R1855 B.n704 B.n703 163.367
R1856 B.n703 B.n702 163.367
R1857 B.n702 B.n17 163.367
R1858 B.n698 B.n17 163.367
R1859 B.n698 B.n697 163.367
R1860 B.n697 B.n696 163.367
R1861 B.n696 B.n19 163.367
R1862 B.n692 B.n19 163.367
R1863 B.n692 B.n691 163.367
R1864 B.n691 B.n690 163.367
R1865 B.n690 B.n21 163.367
R1866 B.n686 B.n21 163.367
R1867 B.n686 B.n685 163.367
R1868 B.n685 B.n684 163.367
R1869 B.n684 B.n23 163.367
R1870 B.n680 B.n23 163.367
R1871 B.n680 B.n679 163.367
R1872 B.n679 B.n678 163.367
R1873 B.n678 B.n25 163.367
R1874 B.n674 B.n25 163.367
R1875 B.n674 B.n673 163.367
R1876 B.n673 B.n672 163.367
R1877 B.n672 B.n27 163.367
R1878 B.n668 B.n27 163.367
R1879 B.n668 B.n667 163.367
R1880 B.n667 B.n666 163.367
R1881 B.n666 B.n29 163.367
R1882 B.n662 B.n29 163.367
R1883 B.n662 B.n661 163.367
R1884 B.n661 B.n660 163.367
R1885 B.n660 B.n31 163.367
R1886 B.n656 B.n31 163.367
R1887 B.n656 B.n655 163.367
R1888 B.n655 B.n654 163.367
R1889 B.n654 B.n33 163.367
R1890 B.n650 B.n33 163.367
R1891 B.n650 B.n649 163.367
R1892 B.n649 B.n648 163.367
R1893 B.n648 B.n35 163.367
R1894 B.n644 B.n35 163.367
R1895 B.n644 B.n643 163.367
R1896 B.n643 B.n642 163.367
R1897 B.n642 B.n37 163.367
R1898 B.n638 B.n37 163.367
R1899 B.n638 B.n637 163.367
R1900 B.n637 B.n636 163.367
R1901 B.n636 B.n39 163.367
R1902 B.n632 B.n39 163.367
R1903 B.n632 B.n631 163.367
R1904 B.n631 B.n630 163.367
R1905 B.n630 B.n41 163.367
R1906 B.n626 B.n41 163.367
R1907 B.n626 B.n625 163.367
R1908 B.n625 B.n624 163.367
R1909 B.n624 B.n43 163.367
R1910 B.n620 B.n43 163.367
R1911 B.n620 B.n619 163.367
R1912 B.n619 B.n618 163.367
R1913 B.n618 B.n45 163.367
R1914 B.n613 B.n45 163.367
R1915 B.n613 B.n612 163.367
R1916 B.n612 B.n611 163.367
R1917 B.n611 B.n49 163.367
R1918 B.n607 B.n49 163.367
R1919 B.n607 B.n606 163.367
R1920 B.n606 B.n605 163.367
R1921 B.n605 B.n51 163.367
R1922 B.n601 B.n51 163.367
R1923 B.n601 B.n600 163.367
R1924 B.n600 B.n55 163.367
R1925 B.n596 B.n55 163.367
R1926 B.n596 B.n595 163.367
R1927 B.n595 B.n594 163.367
R1928 B.n594 B.n57 163.367
R1929 B.n590 B.n57 163.367
R1930 B.n590 B.n589 163.367
R1931 B.n589 B.n588 163.367
R1932 B.n588 B.n59 163.367
R1933 B.n584 B.n59 163.367
R1934 B.n584 B.n583 163.367
R1935 B.n583 B.n582 163.367
R1936 B.n582 B.n61 163.367
R1937 B.n578 B.n61 163.367
R1938 B.n578 B.n577 163.367
R1939 B.n577 B.n576 163.367
R1940 B.n576 B.n63 163.367
R1941 B.n572 B.n63 163.367
R1942 B.n572 B.n571 163.367
R1943 B.n571 B.n570 163.367
R1944 B.n570 B.n65 163.367
R1945 B.n566 B.n65 163.367
R1946 B.n566 B.n565 163.367
R1947 B.n565 B.n564 163.367
R1948 B.n564 B.n67 163.367
R1949 B.n560 B.n67 163.367
R1950 B.n560 B.n559 163.367
R1951 B.n559 B.n558 163.367
R1952 B.n558 B.n69 163.367
R1953 B.n554 B.n69 163.367
R1954 B.n554 B.n553 163.367
R1955 B.n553 B.n552 163.367
R1956 B.n552 B.n71 163.367
R1957 B.n548 B.n71 163.367
R1958 B.n548 B.n547 163.367
R1959 B.n547 B.n546 163.367
R1960 B.n546 B.n73 163.367
R1961 B.n542 B.n73 163.367
R1962 B.n542 B.n541 163.367
R1963 B.n541 B.n540 163.367
R1964 B.n540 B.n75 163.367
R1965 B.n536 B.n75 163.367
R1966 B.n536 B.n535 163.367
R1967 B.n535 B.n534 163.367
R1968 B.n534 B.n77 163.367
R1969 B.n530 B.n77 163.367
R1970 B.n530 B.n529 163.367
R1971 B.n529 B.n528 163.367
R1972 B.n528 B.n79 163.367
R1973 B.n524 B.n79 163.367
R1974 B.n524 B.n523 163.367
R1975 B.n523 B.n522 163.367
R1976 B.n522 B.n81 163.367
R1977 B.n518 B.n81 163.367
R1978 B.n518 B.n517 163.367
R1979 B.n517 B.n516 163.367
R1980 B.n516 B.n83 163.367
R1981 B.n512 B.n83 163.367
R1982 B.n512 B.n511 163.367
R1983 B.n143 B.n142 62.0611
R1984 B.n151 B.n150 62.0611
R1985 B.n47 B.n46 62.0611
R1986 B.n53 B.n52 62.0611
R1987 B.n144 B.n143 59.5399
R1988 B.n323 B.n151 59.5399
R1989 B.n615 B.n47 59.5399
R1990 B.n54 B.n53 59.5399
R1991 B.n706 B.n705 32.6249
R1992 B.n509 B.n84 32.6249
R1993 B.n429 B.n112 32.6249
R1994 B.n233 B.n232 32.6249
R1995 B B.n747 18.0485
R1996 B.n705 B.n16 10.6151
R1997 B.n701 B.n16 10.6151
R1998 B.n701 B.n700 10.6151
R1999 B.n700 B.n699 10.6151
R2000 B.n699 B.n18 10.6151
R2001 B.n695 B.n18 10.6151
R2002 B.n695 B.n694 10.6151
R2003 B.n694 B.n693 10.6151
R2004 B.n693 B.n20 10.6151
R2005 B.n689 B.n20 10.6151
R2006 B.n689 B.n688 10.6151
R2007 B.n688 B.n687 10.6151
R2008 B.n687 B.n22 10.6151
R2009 B.n683 B.n22 10.6151
R2010 B.n683 B.n682 10.6151
R2011 B.n682 B.n681 10.6151
R2012 B.n681 B.n24 10.6151
R2013 B.n677 B.n24 10.6151
R2014 B.n677 B.n676 10.6151
R2015 B.n676 B.n675 10.6151
R2016 B.n675 B.n26 10.6151
R2017 B.n671 B.n26 10.6151
R2018 B.n671 B.n670 10.6151
R2019 B.n670 B.n669 10.6151
R2020 B.n669 B.n28 10.6151
R2021 B.n665 B.n28 10.6151
R2022 B.n665 B.n664 10.6151
R2023 B.n664 B.n663 10.6151
R2024 B.n663 B.n30 10.6151
R2025 B.n659 B.n30 10.6151
R2026 B.n659 B.n658 10.6151
R2027 B.n658 B.n657 10.6151
R2028 B.n657 B.n32 10.6151
R2029 B.n653 B.n32 10.6151
R2030 B.n653 B.n652 10.6151
R2031 B.n652 B.n651 10.6151
R2032 B.n651 B.n34 10.6151
R2033 B.n647 B.n34 10.6151
R2034 B.n647 B.n646 10.6151
R2035 B.n646 B.n645 10.6151
R2036 B.n645 B.n36 10.6151
R2037 B.n641 B.n36 10.6151
R2038 B.n641 B.n640 10.6151
R2039 B.n640 B.n639 10.6151
R2040 B.n639 B.n38 10.6151
R2041 B.n635 B.n38 10.6151
R2042 B.n635 B.n634 10.6151
R2043 B.n634 B.n633 10.6151
R2044 B.n633 B.n40 10.6151
R2045 B.n629 B.n40 10.6151
R2046 B.n629 B.n628 10.6151
R2047 B.n628 B.n627 10.6151
R2048 B.n627 B.n42 10.6151
R2049 B.n623 B.n42 10.6151
R2050 B.n623 B.n622 10.6151
R2051 B.n622 B.n621 10.6151
R2052 B.n621 B.n44 10.6151
R2053 B.n617 B.n44 10.6151
R2054 B.n617 B.n616 10.6151
R2055 B.n614 B.n48 10.6151
R2056 B.n610 B.n48 10.6151
R2057 B.n610 B.n609 10.6151
R2058 B.n609 B.n608 10.6151
R2059 B.n608 B.n50 10.6151
R2060 B.n604 B.n50 10.6151
R2061 B.n604 B.n603 10.6151
R2062 B.n603 B.n602 10.6151
R2063 B.n599 B.n598 10.6151
R2064 B.n598 B.n597 10.6151
R2065 B.n597 B.n56 10.6151
R2066 B.n593 B.n56 10.6151
R2067 B.n593 B.n592 10.6151
R2068 B.n592 B.n591 10.6151
R2069 B.n591 B.n58 10.6151
R2070 B.n587 B.n58 10.6151
R2071 B.n587 B.n586 10.6151
R2072 B.n586 B.n585 10.6151
R2073 B.n585 B.n60 10.6151
R2074 B.n581 B.n60 10.6151
R2075 B.n581 B.n580 10.6151
R2076 B.n580 B.n579 10.6151
R2077 B.n579 B.n62 10.6151
R2078 B.n575 B.n62 10.6151
R2079 B.n575 B.n574 10.6151
R2080 B.n574 B.n573 10.6151
R2081 B.n573 B.n64 10.6151
R2082 B.n569 B.n64 10.6151
R2083 B.n569 B.n568 10.6151
R2084 B.n568 B.n567 10.6151
R2085 B.n567 B.n66 10.6151
R2086 B.n563 B.n66 10.6151
R2087 B.n563 B.n562 10.6151
R2088 B.n562 B.n561 10.6151
R2089 B.n561 B.n68 10.6151
R2090 B.n557 B.n68 10.6151
R2091 B.n557 B.n556 10.6151
R2092 B.n556 B.n555 10.6151
R2093 B.n555 B.n70 10.6151
R2094 B.n551 B.n70 10.6151
R2095 B.n551 B.n550 10.6151
R2096 B.n550 B.n549 10.6151
R2097 B.n549 B.n72 10.6151
R2098 B.n545 B.n72 10.6151
R2099 B.n545 B.n544 10.6151
R2100 B.n544 B.n543 10.6151
R2101 B.n543 B.n74 10.6151
R2102 B.n539 B.n74 10.6151
R2103 B.n539 B.n538 10.6151
R2104 B.n538 B.n537 10.6151
R2105 B.n537 B.n76 10.6151
R2106 B.n533 B.n76 10.6151
R2107 B.n533 B.n532 10.6151
R2108 B.n532 B.n531 10.6151
R2109 B.n531 B.n78 10.6151
R2110 B.n527 B.n78 10.6151
R2111 B.n527 B.n526 10.6151
R2112 B.n526 B.n525 10.6151
R2113 B.n525 B.n80 10.6151
R2114 B.n521 B.n80 10.6151
R2115 B.n521 B.n520 10.6151
R2116 B.n520 B.n519 10.6151
R2117 B.n519 B.n82 10.6151
R2118 B.n515 B.n82 10.6151
R2119 B.n515 B.n514 10.6151
R2120 B.n514 B.n513 10.6151
R2121 B.n513 B.n84 10.6151
R2122 B.n430 B.n429 10.6151
R2123 B.n431 B.n430 10.6151
R2124 B.n431 B.n110 10.6151
R2125 B.n435 B.n110 10.6151
R2126 B.n436 B.n435 10.6151
R2127 B.n437 B.n436 10.6151
R2128 B.n437 B.n108 10.6151
R2129 B.n441 B.n108 10.6151
R2130 B.n442 B.n441 10.6151
R2131 B.n443 B.n442 10.6151
R2132 B.n443 B.n106 10.6151
R2133 B.n447 B.n106 10.6151
R2134 B.n448 B.n447 10.6151
R2135 B.n449 B.n448 10.6151
R2136 B.n449 B.n104 10.6151
R2137 B.n453 B.n104 10.6151
R2138 B.n454 B.n453 10.6151
R2139 B.n455 B.n454 10.6151
R2140 B.n455 B.n102 10.6151
R2141 B.n459 B.n102 10.6151
R2142 B.n460 B.n459 10.6151
R2143 B.n461 B.n460 10.6151
R2144 B.n461 B.n100 10.6151
R2145 B.n465 B.n100 10.6151
R2146 B.n466 B.n465 10.6151
R2147 B.n467 B.n466 10.6151
R2148 B.n467 B.n98 10.6151
R2149 B.n471 B.n98 10.6151
R2150 B.n472 B.n471 10.6151
R2151 B.n473 B.n472 10.6151
R2152 B.n473 B.n96 10.6151
R2153 B.n477 B.n96 10.6151
R2154 B.n478 B.n477 10.6151
R2155 B.n479 B.n478 10.6151
R2156 B.n479 B.n94 10.6151
R2157 B.n483 B.n94 10.6151
R2158 B.n484 B.n483 10.6151
R2159 B.n485 B.n484 10.6151
R2160 B.n485 B.n92 10.6151
R2161 B.n489 B.n92 10.6151
R2162 B.n490 B.n489 10.6151
R2163 B.n491 B.n490 10.6151
R2164 B.n491 B.n90 10.6151
R2165 B.n495 B.n90 10.6151
R2166 B.n496 B.n495 10.6151
R2167 B.n497 B.n496 10.6151
R2168 B.n497 B.n88 10.6151
R2169 B.n501 B.n88 10.6151
R2170 B.n502 B.n501 10.6151
R2171 B.n503 B.n502 10.6151
R2172 B.n503 B.n86 10.6151
R2173 B.n507 B.n86 10.6151
R2174 B.n508 B.n507 10.6151
R2175 B.n509 B.n508 10.6151
R2176 B.n233 B.n180 10.6151
R2177 B.n237 B.n180 10.6151
R2178 B.n238 B.n237 10.6151
R2179 B.n239 B.n238 10.6151
R2180 B.n239 B.n178 10.6151
R2181 B.n243 B.n178 10.6151
R2182 B.n244 B.n243 10.6151
R2183 B.n245 B.n244 10.6151
R2184 B.n245 B.n176 10.6151
R2185 B.n249 B.n176 10.6151
R2186 B.n250 B.n249 10.6151
R2187 B.n251 B.n250 10.6151
R2188 B.n251 B.n174 10.6151
R2189 B.n255 B.n174 10.6151
R2190 B.n256 B.n255 10.6151
R2191 B.n257 B.n256 10.6151
R2192 B.n257 B.n172 10.6151
R2193 B.n261 B.n172 10.6151
R2194 B.n262 B.n261 10.6151
R2195 B.n263 B.n262 10.6151
R2196 B.n263 B.n170 10.6151
R2197 B.n267 B.n170 10.6151
R2198 B.n268 B.n267 10.6151
R2199 B.n269 B.n268 10.6151
R2200 B.n269 B.n168 10.6151
R2201 B.n273 B.n168 10.6151
R2202 B.n274 B.n273 10.6151
R2203 B.n275 B.n274 10.6151
R2204 B.n275 B.n166 10.6151
R2205 B.n279 B.n166 10.6151
R2206 B.n280 B.n279 10.6151
R2207 B.n281 B.n280 10.6151
R2208 B.n281 B.n164 10.6151
R2209 B.n285 B.n164 10.6151
R2210 B.n286 B.n285 10.6151
R2211 B.n287 B.n286 10.6151
R2212 B.n287 B.n162 10.6151
R2213 B.n291 B.n162 10.6151
R2214 B.n292 B.n291 10.6151
R2215 B.n293 B.n292 10.6151
R2216 B.n293 B.n160 10.6151
R2217 B.n297 B.n160 10.6151
R2218 B.n298 B.n297 10.6151
R2219 B.n299 B.n298 10.6151
R2220 B.n299 B.n158 10.6151
R2221 B.n303 B.n158 10.6151
R2222 B.n304 B.n303 10.6151
R2223 B.n305 B.n304 10.6151
R2224 B.n305 B.n156 10.6151
R2225 B.n309 B.n156 10.6151
R2226 B.n310 B.n309 10.6151
R2227 B.n311 B.n310 10.6151
R2228 B.n311 B.n154 10.6151
R2229 B.n315 B.n154 10.6151
R2230 B.n316 B.n315 10.6151
R2231 B.n317 B.n316 10.6151
R2232 B.n317 B.n152 10.6151
R2233 B.n321 B.n152 10.6151
R2234 B.n322 B.n321 10.6151
R2235 B.n324 B.n148 10.6151
R2236 B.n328 B.n148 10.6151
R2237 B.n329 B.n328 10.6151
R2238 B.n330 B.n329 10.6151
R2239 B.n330 B.n146 10.6151
R2240 B.n334 B.n146 10.6151
R2241 B.n335 B.n334 10.6151
R2242 B.n336 B.n335 10.6151
R2243 B.n340 B.n339 10.6151
R2244 B.n341 B.n340 10.6151
R2245 B.n341 B.n140 10.6151
R2246 B.n345 B.n140 10.6151
R2247 B.n346 B.n345 10.6151
R2248 B.n347 B.n346 10.6151
R2249 B.n347 B.n138 10.6151
R2250 B.n351 B.n138 10.6151
R2251 B.n352 B.n351 10.6151
R2252 B.n353 B.n352 10.6151
R2253 B.n353 B.n136 10.6151
R2254 B.n357 B.n136 10.6151
R2255 B.n358 B.n357 10.6151
R2256 B.n359 B.n358 10.6151
R2257 B.n359 B.n134 10.6151
R2258 B.n363 B.n134 10.6151
R2259 B.n364 B.n363 10.6151
R2260 B.n365 B.n364 10.6151
R2261 B.n365 B.n132 10.6151
R2262 B.n369 B.n132 10.6151
R2263 B.n370 B.n369 10.6151
R2264 B.n371 B.n370 10.6151
R2265 B.n371 B.n130 10.6151
R2266 B.n375 B.n130 10.6151
R2267 B.n376 B.n375 10.6151
R2268 B.n377 B.n376 10.6151
R2269 B.n377 B.n128 10.6151
R2270 B.n381 B.n128 10.6151
R2271 B.n382 B.n381 10.6151
R2272 B.n383 B.n382 10.6151
R2273 B.n383 B.n126 10.6151
R2274 B.n387 B.n126 10.6151
R2275 B.n388 B.n387 10.6151
R2276 B.n389 B.n388 10.6151
R2277 B.n389 B.n124 10.6151
R2278 B.n393 B.n124 10.6151
R2279 B.n394 B.n393 10.6151
R2280 B.n395 B.n394 10.6151
R2281 B.n395 B.n122 10.6151
R2282 B.n399 B.n122 10.6151
R2283 B.n400 B.n399 10.6151
R2284 B.n401 B.n400 10.6151
R2285 B.n401 B.n120 10.6151
R2286 B.n405 B.n120 10.6151
R2287 B.n406 B.n405 10.6151
R2288 B.n407 B.n406 10.6151
R2289 B.n407 B.n118 10.6151
R2290 B.n411 B.n118 10.6151
R2291 B.n412 B.n411 10.6151
R2292 B.n413 B.n412 10.6151
R2293 B.n413 B.n116 10.6151
R2294 B.n417 B.n116 10.6151
R2295 B.n418 B.n417 10.6151
R2296 B.n419 B.n418 10.6151
R2297 B.n419 B.n114 10.6151
R2298 B.n423 B.n114 10.6151
R2299 B.n424 B.n423 10.6151
R2300 B.n425 B.n424 10.6151
R2301 B.n425 B.n112 10.6151
R2302 B.n232 B.n231 10.6151
R2303 B.n231 B.n182 10.6151
R2304 B.n227 B.n182 10.6151
R2305 B.n227 B.n226 10.6151
R2306 B.n226 B.n225 10.6151
R2307 B.n225 B.n184 10.6151
R2308 B.n221 B.n184 10.6151
R2309 B.n221 B.n220 10.6151
R2310 B.n220 B.n219 10.6151
R2311 B.n219 B.n186 10.6151
R2312 B.n215 B.n186 10.6151
R2313 B.n215 B.n214 10.6151
R2314 B.n214 B.n213 10.6151
R2315 B.n213 B.n188 10.6151
R2316 B.n209 B.n188 10.6151
R2317 B.n209 B.n208 10.6151
R2318 B.n208 B.n207 10.6151
R2319 B.n207 B.n190 10.6151
R2320 B.n203 B.n190 10.6151
R2321 B.n203 B.n202 10.6151
R2322 B.n202 B.n201 10.6151
R2323 B.n201 B.n192 10.6151
R2324 B.n197 B.n192 10.6151
R2325 B.n197 B.n196 10.6151
R2326 B.n196 B.n195 10.6151
R2327 B.n195 B.n0 10.6151
R2328 B.n743 B.n1 10.6151
R2329 B.n743 B.n742 10.6151
R2330 B.n742 B.n741 10.6151
R2331 B.n741 B.n4 10.6151
R2332 B.n737 B.n4 10.6151
R2333 B.n737 B.n736 10.6151
R2334 B.n736 B.n735 10.6151
R2335 B.n735 B.n6 10.6151
R2336 B.n731 B.n6 10.6151
R2337 B.n731 B.n730 10.6151
R2338 B.n730 B.n729 10.6151
R2339 B.n729 B.n8 10.6151
R2340 B.n725 B.n8 10.6151
R2341 B.n725 B.n724 10.6151
R2342 B.n724 B.n723 10.6151
R2343 B.n723 B.n10 10.6151
R2344 B.n719 B.n10 10.6151
R2345 B.n719 B.n718 10.6151
R2346 B.n718 B.n717 10.6151
R2347 B.n717 B.n12 10.6151
R2348 B.n713 B.n12 10.6151
R2349 B.n713 B.n712 10.6151
R2350 B.n712 B.n711 10.6151
R2351 B.n711 B.n14 10.6151
R2352 B.n707 B.n14 10.6151
R2353 B.n707 B.n706 10.6151
R2354 B.n615 B.n614 6.5566
R2355 B.n602 B.n54 6.5566
R2356 B.n324 B.n323 6.5566
R2357 B.n336 B.n144 6.5566
R2358 B.n616 B.n615 4.05904
R2359 B.n599 B.n54 4.05904
R2360 B.n323 B.n322 4.05904
R2361 B.n339 B.n144 4.05904
R2362 B.n747 B.n0 2.81026
R2363 B.n747 B.n1 2.81026
C0 VDD2 VN 4.14438f
C1 VTAIL B 5.17216f
C2 VN B 1.17193f
C3 VDD2 B 2.2658f
C4 VDD1 w_n2250_n4604# 2.2385f
C5 VP w_n2250_n4604# 3.53731f
C6 VTAIL w_n2250_n4604# 3.59893f
C7 VN w_n2250_n4604# 3.25012f
C8 VDD2 w_n2250_n4604# 2.26772f
C9 w_n2250_n4604# B 10.8331f
C10 VP VDD1 4.33759f
C11 VTAIL VDD1 6.71366f
C12 VN VDD1 0.14858f
C13 VP VTAIL 3.56942f
C14 VP VN 6.72417f
C15 VDD2 VDD1 0.707944f
C16 VN VTAIL 3.55507f
C17 VDD1 B 2.23332f
C18 VDD2 VP 0.345194f
C19 VDD2 VTAIL 6.76505f
C20 VP B 1.64517f
C21 VDD2 VSUBS 1.156699f
C22 VDD1 VSUBS 5.621799f
C23 VTAIL VSUBS 1.285435f
C24 VN VSUBS 9.20429f
C25 VP VSUBS 1.988155f
C26 B VSUBS 4.630575f
C27 w_n2250_n4604# VSUBS 0.126657p
C28 B.n0 VSUBS 0.004234f
C29 B.n1 VSUBS 0.004234f
C30 B.n2 VSUBS 0.006695f
C31 B.n3 VSUBS 0.006695f
C32 B.n4 VSUBS 0.006695f
C33 B.n5 VSUBS 0.006695f
C34 B.n6 VSUBS 0.006695f
C35 B.n7 VSUBS 0.006695f
C36 B.n8 VSUBS 0.006695f
C37 B.n9 VSUBS 0.006695f
C38 B.n10 VSUBS 0.006695f
C39 B.n11 VSUBS 0.006695f
C40 B.n12 VSUBS 0.006695f
C41 B.n13 VSUBS 0.006695f
C42 B.n14 VSUBS 0.006695f
C43 B.n15 VSUBS 0.015375f
C44 B.n16 VSUBS 0.006695f
C45 B.n17 VSUBS 0.006695f
C46 B.n18 VSUBS 0.006695f
C47 B.n19 VSUBS 0.006695f
C48 B.n20 VSUBS 0.006695f
C49 B.n21 VSUBS 0.006695f
C50 B.n22 VSUBS 0.006695f
C51 B.n23 VSUBS 0.006695f
C52 B.n24 VSUBS 0.006695f
C53 B.n25 VSUBS 0.006695f
C54 B.n26 VSUBS 0.006695f
C55 B.n27 VSUBS 0.006695f
C56 B.n28 VSUBS 0.006695f
C57 B.n29 VSUBS 0.006695f
C58 B.n30 VSUBS 0.006695f
C59 B.n31 VSUBS 0.006695f
C60 B.n32 VSUBS 0.006695f
C61 B.n33 VSUBS 0.006695f
C62 B.n34 VSUBS 0.006695f
C63 B.n35 VSUBS 0.006695f
C64 B.n36 VSUBS 0.006695f
C65 B.n37 VSUBS 0.006695f
C66 B.n38 VSUBS 0.006695f
C67 B.n39 VSUBS 0.006695f
C68 B.n40 VSUBS 0.006695f
C69 B.n41 VSUBS 0.006695f
C70 B.n42 VSUBS 0.006695f
C71 B.n43 VSUBS 0.006695f
C72 B.n44 VSUBS 0.006695f
C73 B.n45 VSUBS 0.006695f
C74 B.t8 VSUBS 0.339943f
C75 B.t7 VSUBS 0.374762f
C76 B.t6 VSUBS 2.2284f
C77 B.n46 VSUBS 0.581397f
C78 B.n47 VSUBS 0.317552f
C79 B.n48 VSUBS 0.006695f
C80 B.n49 VSUBS 0.006695f
C81 B.n50 VSUBS 0.006695f
C82 B.n51 VSUBS 0.006695f
C83 B.t2 VSUBS 0.339947f
C84 B.t1 VSUBS 0.374765f
C85 B.t0 VSUBS 2.2284f
C86 B.n52 VSUBS 0.581394f
C87 B.n53 VSUBS 0.317549f
C88 B.n54 VSUBS 0.015512f
C89 B.n55 VSUBS 0.006695f
C90 B.n56 VSUBS 0.006695f
C91 B.n57 VSUBS 0.006695f
C92 B.n58 VSUBS 0.006695f
C93 B.n59 VSUBS 0.006695f
C94 B.n60 VSUBS 0.006695f
C95 B.n61 VSUBS 0.006695f
C96 B.n62 VSUBS 0.006695f
C97 B.n63 VSUBS 0.006695f
C98 B.n64 VSUBS 0.006695f
C99 B.n65 VSUBS 0.006695f
C100 B.n66 VSUBS 0.006695f
C101 B.n67 VSUBS 0.006695f
C102 B.n68 VSUBS 0.006695f
C103 B.n69 VSUBS 0.006695f
C104 B.n70 VSUBS 0.006695f
C105 B.n71 VSUBS 0.006695f
C106 B.n72 VSUBS 0.006695f
C107 B.n73 VSUBS 0.006695f
C108 B.n74 VSUBS 0.006695f
C109 B.n75 VSUBS 0.006695f
C110 B.n76 VSUBS 0.006695f
C111 B.n77 VSUBS 0.006695f
C112 B.n78 VSUBS 0.006695f
C113 B.n79 VSUBS 0.006695f
C114 B.n80 VSUBS 0.006695f
C115 B.n81 VSUBS 0.006695f
C116 B.n82 VSUBS 0.006695f
C117 B.n83 VSUBS 0.006695f
C118 B.n84 VSUBS 0.015143f
C119 B.n85 VSUBS 0.006695f
C120 B.n86 VSUBS 0.006695f
C121 B.n87 VSUBS 0.006695f
C122 B.n88 VSUBS 0.006695f
C123 B.n89 VSUBS 0.006695f
C124 B.n90 VSUBS 0.006695f
C125 B.n91 VSUBS 0.006695f
C126 B.n92 VSUBS 0.006695f
C127 B.n93 VSUBS 0.006695f
C128 B.n94 VSUBS 0.006695f
C129 B.n95 VSUBS 0.006695f
C130 B.n96 VSUBS 0.006695f
C131 B.n97 VSUBS 0.006695f
C132 B.n98 VSUBS 0.006695f
C133 B.n99 VSUBS 0.006695f
C134 B.n100 VSUBS 0.006695f
C135 B.n101 VSUBS 0.006695f
C136 B.n102 VSUBS 0.006695f
C137 B.n103 VSUBS 0.006695f
C138 B.n104 VSUBS 0.006695f
C139 B.n105 VSUBS 0.006695f
C140 B.n106 VSUBS 0.006695f
C141 B.n107 VSUBS 0.006695f
C142 B.n108 VSUBS 0.006695f
C143 B.n109 VSUBS 0.006695f
C144 B.n110 VSUBS 0.006695f
C145 B.n111 VSUBS 0.006695f
C146 B.n112 VSUBS 0.015935f
C147 B.n113 VSUBS 0.006695f
C148 B.n114 VSUBS 0.006695f
C149 B.n115 VSUBS 0.006695f
C150 B.n116 VSUBS 0.006695f
C151 B.n117 VSUBS 0.006695f
C152 B.n118 VSUBS 0.006695f
C153 B.n119 VSUBS 0.006695f
C154 B.n120 VSUBS 0.006695f
C155 B.n121 VSUBS 0.006695f
C156 B.n122 VSUBS 0.006695f
C157 B.n123 VSUBS 0.006695f
C158 B.n124 VSUBS 0.006695f
C159 B.n125 VSUBS 0.006695f
C160 B.n126 VSUBS 0.006695f
C161 B.n127 VSUBS 0.006695f
C162 B.n128 VSUBS 0.006695f
C163 B.n129 VSUBS 0.006695f
C164 B.n130 VSUBS 0.006695f
C165 B.n131 VSUBS 0.006695f
C166 B.n132 VSUBS 0.006695f
C167 B.n133 VSUBS 0.006695f
C168 B.n134 VSUBS 0.006695f
C169 B.n135 VSUBS 0.006695f
C170 B.n136 VSUBS 0.006695f
C171 B.n137 VSUBS 0.006695f
C172 B.n138 VSUBS 0.006695f
C173 B.n139 VSUBS 0.006695f
C174 B.n140 VSUBS 0.006695f
C175 B.n141 VSUBS 0.006695f
C176 B.t4 VSUBS 0.339947f
C177 B.t5 VSUBS 0.374765f
C178 B.t3 VSUBS 2.2284f
C179 B.n142 VSUBS 0.581394f
C180 B.n143 VSUBS 0.317549f
C181 B.n144 VSUBS 0.015512f
C182 B.n145 VSUBS 0.006695f
C183 B.n146 VSUBS 0.006695f
C184 B.n147 VSUBS 0.006695f
C185 B.n148 VSUBS 0.006695f
C186 B.n149 VSUBS 0.006695f
C187 B.t10 VSUBS 0.339943f
C188 B.t11 VSUBS 0.374762f
C189 B.t9 VSUBS 2.2284f
C190 B.n150 VSUBS 0.581397f
C191 B.n151 VSUBS 0.317552f
C192 B.n152 VSUBS 0.006695f
C193 B.n153 VSUBS 0.006695f
C194 B.n154 VSUBS 0.006695f
C195 B.n155 VSUBS 0.006695f
C196 B.n156 VSUBS 0.006695f
C197 B.n157 VSUBS 0.006695f
C198 B.n158 VSUBS 0.006695f
C199 B.n159 VSUBS 0.006695f
C200 B.n160 VSUBS 0.006695f
C201 B.n161 VSUBS 0.006695f
C202 B.n162 VSUBS 0.006695f
C203 B.n163 VSUBS 0.006695f
C204 B.n164 VSUBS 0.006695f
C205 B.n165 VSUBS 0.006695f
C206 B.n166 VSUBS 0.006695f
C207 B.n167 VSUBS 0.006695f
C208 B.n168 VSUBS 0.006695f
C209 B.n169 VSUBS 0.006695f
C210 B.n170 VSUBS 0.006695f
C211 B.n171 VSUBS 0.006695f
C212 B.n172 VSUBS 0.006695f
C213 B.n173 VSUBS 0.006695f
C214 B.n174 VSUBS 0.006695f
C215 B.n175 VSUBS 0.006695f
C216 B.n176 VSUBS 0.006695f
C217 B.n177 VSUBS 0.006695f
C218 B.n178 VSUBS 0.006695f
C219 B.n179 VSUBS 0.006695f
C220 B.n180 VSUBS 0.006695f
C221 B.n181 VSUBS 0.015375f
C222 B.n182 VSUBS 0.006695f
C223 B.n183 VSUBS 0.006695f
C224 B.n184 VSUBS 0.006695f
C225 B.n185 VSUBS 0.006695f
C226 B.n186 VSUBS 0.006695f
C227 B.n187 VSUBS 0.006695f
C228 B.n188 VSUBS 0.006695f
C229 B.n189 VSUBS 0.006695f
C230 B.n190 VSUBS 0.006695f
C231 B.n191 VSUBS 0.006695f
C232 B.n192 VSUBS 0.006695f
C233 B.n193 VSUBS 0.006695f
C234 B.n194 VSUBS 0.006695f
C235 B.n195 VSUBS 0.006695f
C236 B.n196 VSUBS 0.006695f
C237 B.n197 VSUBS 0.006695f
C238 B.n198 VSUBS 0.006695f
C239 B.n199 VSUBS 0.006695f
C240 B.n200 VSUBS 0.006695f
C241 B.n201 VSUBS 0.006695f
C242 B.n202 VSUBS 0.006695f
C243 B.n203 VSUBS 0.006695f
C244 B.n204 VSUBS 0.006695f
C245 B.n205 VSUBS 0.006695f
C246 B.n206 VSUBS 0.006695f
C247 B.n207 VSUBS 0.006695f
C248 B.n208 VSUBS 0.006695f
C249 B.n209 VSUBS 0.006695f
C250 B.n210 VSUBS 0.006695f
C251 B.n211 VSUBS 0.006695f
C252 B.n212 VSUBS 0.006695f
C253 B.n213 VSUBS 0.006695f
C254 B.n214 VSUBS 0.006695f
C255 B.n215 VSUBS 0.006695f
C256 B.n216 VSUBS 0.006695f
C257 B.n217 VSUBS 0.006695f
C258 B.n218 VSUBS 0.006695f
C259 B.n219 VSUBS 0.006695f
C260 B.n220 VSUBS 0.006695f
C261 B.n221 VSUBS 0.006695f
C262 B.n222 VSUBS 0.006695f
C263 B.n223 VSUBS 0.006695f
C264 B.n224 VSUBS 0.006695f
C265 B.n225 VSUBS 0.006695f
C266 B.n226 VSUBS 0.006695f
C267 B.n227 VSUBS 0.006695f
C268 B.n228 VSUBS 0.006695f
C269 B.n229 VSUBS 0.006695f
C270 B.n230 VSUBS 0.006695f
C271 B.n231 VSUBS 0.006695f
C272 B.n232 VSUBS 0.015375f
C273 B.n233 VSUBS 0.015935f
C274 B.n234 VSUBS 0.015935f
C275 B.n235 VSUBS 0.006695f
C276 B.n236 VSUBS 0.006695f
C277 B.n237 VSUBS 0.006695f
C278 B.n238 VSUBS 0.006695f
C279 B.n239 VSUBS 0.006695f
C280 B.n240 VSUBS 0.006695f
C281 B.n241 VSUBS 0.006695f
C282 B.n242 VSUBS 0.006695f
C283 B.n243 VSUBS 0.006695f
C284 B.n244 VSUBS 0.006695f
C285 B.n245 VSUBS 0.006695f
C286 B.n246 VSUBS 0.006695f
C287 B.n247 VSUBS 0.006695f
C288 B.n248 VSUBS 0.006695f
C289 B.n249 VSUBS 0.006695f
C290 B.n250 VSUBS 0.006695f
C291 B.n251 VSUBS 0.006695f
C292 B.n252 VSUBS 0.006695f
C293 B.n253 VSUBS 0.006695f
C294 B.n254 VSUBS 0.006695f
C295 B.n255 VSUBS 0.006695f
C296 B.n256 VSUBS 0.006695f
C297 B.n257 VSUBS 0.006695f
C298 B.n258 VSUBS 0.006695f
C299 B.n259 VSUBS 0.006695f
C300 B.n260 VSUBS 0.006695f
C301 B.n261 VSUBS 0.006695f
C302 B.n262 VSUBS 0.006695f
C303 B.n263 VSUBS 0.006695f
C304 B.n264 VSUBS 0.006695f
C305 B.n265 VSUBS 0.006695f
C306 B.n266 VSUBS 0.006695f
C307 B.n267 VSUBS 0.006695f
C308 B.n268 VSUBS 0.006695f
C309 B.n269 VSUBS 0.006695f
C310 B.n270 VSUBS 0.006695f
C311 B.n271 VSUBS 0.006695f
C312 B.n272 VSUBS 0.006695f
C313 B.n273 VSUBS 0.006695f
C314 B.n274 VSUBS 0.006695f
C315 B.n275 VSUBS 0.006695f
C316 B.n276 VSUBS 0.006695f
C317 B.n277 VSUBS 0.006695f
C318 B.n278 VSUBS 0.006695f
C319 B.n279 VSUBS 0.006695f
C320 B.n280 VSUBS 0.006695f
C321 B.n281 VSUBS 0.006695f
C322 B.n282 VSUBS 0.006695f
C323 B.n283 VSUBS 0.006695f
C324 B.n284 VSUBS 0.006695f
C325 B.n285 VSUBS 0.006695f
C326 B.n286 VSUBS 0.006695f
C327 B.n287 VSUBS 0.006695f
C328 B.n288 VSUBS 0.006695f
C329 B.n289 VSUBS 0.006695f
C330 B.n290 VSUBS 0.006695f
C331 B.n291 VSUBS 0.006695f
C332 B.n292 VSUBS 0.006695f
C333 B.n293 VSUBS 0.006695f
C334 B.n294 VSUBS 0.006695f
C335 B.n295 VSUBS 0.006695f
C336 B.n296 VSUBS 0.006695f
C337 B.n297 VSUBS 0.006695f
C338 B.n298 VSUBS 0.006695f
C339 B.n299 VSUBS 0.006695f
C340 B.n300 VSUBS 0.006695f
C341 B.n301 VSUBS 0.006695f
C342 B.n302 VSUBS 0.006695f
C343 B.n303 VSUBS 0.006695f
C344 B.n304 VSUBS 0.006695f
C345 B.n305 VSUBS 0.006695f
C346 B.n306 VSUBS 0.006695f
C347 B.n307 VSUBS 0.006695f
C348 B.n308 VSUBS 0.006695f
C349 B.n309 VSUBS 0.006695f
C350 B.n310 VSUBS 0.006695f
C351 B.n311 VSUBS 0.006695f
C352 B.n312 VSUBS 0.006695f
C353 B.n313 VSUBS 0.006695f
C354 B.n314 VSUBS 0.006695f
C355 B.n315 VSUBS 0.006695f
C356 B.n316 VSUBS 0.006695f
C357 B.n317 VSUBS 0.006695f
C358 B.n318 VSUBS 0.006695f
C359 B.n319 VSUBS 0.006695f
C360 B.n320 VSUBS 0.006695f
C361 B.n321 VSUBS 0.006695f
C362 B.n322 VSUBS 0.004628f
C363 B.n323 VSUBS 0.015512f
C364 B.n324 VSUBS 0.005415f
C365 B.n325 VSUBS 0.006695f
C366 B.n326 VSUBS 0.006695f
C367 B.n327 VSUBS 0.006695f
C368 B.n328 VSUBS 0.006695f
C369 B.n329 VSUBS 0.006695f
C370 B.n330 VSUBS 0.006695f
C371 B.n331 VSUBS 0.006695f
C372 B.n332 VSUBS 0.006695f
C373 B.n333 VSUBS 0.006695f
C374 B.n334 VSUBS 0.006695f
C375 B.n335 VSUBS 0.006695f
C376 B.n336 VSUBS 0.005415f
C377 B.n337 VSUBS 0.006695f
C378 B.n338 VSUBS 0.006695f
C379 B.n339 VSUBS 0.004628f
C380 B.n340 VSUBS 0.006695f
C381 B.n341 VSUBS 0.006695f
C382 B.n342 VSUBS 0.006695f
C383 B.n343 VSUBS 0.006695f
C384 B.n344 VSUBS 0.006695f
C385 B.n345 VSUBS 0.006695f
C386 B.n346 VSUBS 0.006695f
C387 B.n347 VSUBS 0.006695f
C388 B.n348 VSUBS 0.006695f
C389 B.n349 VSUBS 0.006695f
C390 B.n350 VSUBS 0.006695f
C391 B.n351 VSUBS 0.006695f
C392 B.n352 VSUBS 0.006695f
C393 B.n353 VSUBS 0.006695f
C394 B.n354 VSUBS 0.006695f
C395 B.n355 VSUBS 0.006695f
C396 B.n356 VSUBS 0.006695f
C397 B.n357 VSUBS 0.006695f
C398 B.n358 VSUBS 0.006695f
C399 B.n359 VSUBS 0.006695f
C400 B.n360 VSUBS 0.006695f
C401 B.n361 VSUBS 0.006695f
C402 B.n362 VSUBS 0.006695f
C403 B.n363 VSUBS 0.006695f
C404 B.n364 VSUBS 0.006695f
C405 B.n365 VSUBS 0.006695f
C406 B.n366 VSUBS 0.006695f
C407 B.n367 VSUBS 0.006695f
C408 B.n368 VSUBS 0.006695f
C409 B.n369 VSUBS 0.006695f
C410 B.n370 VSUBS 0.006695f
C411 B.n371 VSUBS 0.006695f
C412 B.n372 VSUBS 0.006695f
C413 B.n373 VSUBS 0.006695f
C414 B.n374 VSUBS 0.006695f
C415 B.n375 VSUBS 0.006695f
C416 B.n376 VSUBS 0.006695f
C417 B.n377 VSUBS 0.006695f
C418 B.n378 VSUBS 0.006695f
C419 B.n379 VSUBS 0.006695f
C420 B.n380 VSUBS 0.006695f
C421 B.n381 VSUBS 0.006695f
C422 B.n382 VSUBS 0.006695f
C423 B.n383 VSUBS 0.006695f
C424 B.n384 VSUBS 0.006695f
C425 B.n385 VSUBS 0.006695f
C426 B.n386 VSUBS 0.006695f
C427 B.n387 VSUBS 0.006695f
C428 B.n388 VSUBS 0.006695f
C429 B.n389 VSUBS 0.006695f
C430 B.n390 VSUBS 0.006695f
C431 B.n391 VSUBS 0.006695f
C432 B.n392 VSUBS 0.006695f
C433 B.n393 VSUBS 0.006695f
C434 B.n394 VSUBS 0.006695f
C435 B.n395 VSUBS 0.006695f
C436 B.n396 VSUBS 0.006695f
C437 B.n397 VSUBS 0.006695f
C438 B.n398 VSUBS 0.006695f
C439 B.n399 VSUBS 0.006695f
C440 B.n400 VSUBS 0.006695f
C441 B.n401 VSUBS 0.006695f
C442 B.n402 VSUBS 0.006695f
C443 B.n403 VSUBS 0.006695f
C444 B.n404 VSUBS 0.006695f
C445 B.n405 VSUBS 0.006695f
C446 B.n406 VSUBS 0.006695f
C447 B.n407 VSUBS 0.006695f
C448 B.n408 VSUBS 0.006695f
C449 B.n409 VSUBS 0.006695f
C450 B.n410 VSUBS 0.006695f
C451 B.n411 VSUBS 0.006695f
C452 B.n412 VSUBS 0.006695f
C453 B.n413 VSUBS 0.006695f
C454 B.n414 VSUBS 0.006695f
C455 B.n415 VSUBS 0.006695f
C456 B.n416 VSUBS 0.006695f
C457 B.n417 VSUBS 0.006695f
C458 B.n418 VSUBS 0.006695f
C459 B.n419 VSUBS 0.006695f
C460 B.n420 VSUBS 0.006695f
C461 B.n421 VSUBS 0.006695f
C462 B.n422 VSUBS 0.006695f
C463 B.n423 VSUBS 0.006695f
C464 B.n424 VSUBS 0.006695f
C465 B.n425 VSUBS 0.006695f
C466 B.n426 VSUBS 0.006695f
C467 B.n427 VSUBS 0.015935f
C468 B.n428 VSUBS 0.015375f
C469 B.n429 VSUBS 0.015375f
C470 B.n430 VSUBS 0.006695f
C471 B.n431 VSUBS 0.006695f
C472 B.n432 VSUBS 0.006695f
C473 B.n433 VSUBS 0.006695f
C474 B.n434 VSUBS 0.006695f
C475 B.n435 VSUBS 0.006695f
C476 B.n436 VSUBS 0.006695f
C477 B.n437 VSUBS 0.006695f
C478 B.n438 VSUBS 0.006695f
C479 B.n439 VSUBS 0.006695f
C480 B.n440 VSUBS 0.006695f
C481 B.n441 VSUBS 0.006695f
C482 B.n442 VSUBS 0.006695f
C483 B.n443 VSUBS 0.006695f
C484 B.n444 VSUBS 0.006695f
C485 B.n445 VSUBS 0.006695f
C486 B.n446 VSUBS 0.006695f
C487 B.n447 VSUBS 0.006695f
C488 B.n448 VSUBS 0.006695f
C489 B.n449 VSUBS 0.006695f
C490 B.n450 VSUBS 0.006695f
C491 B.n451 VSUBS 0.006695f
C492 B.n452 VSUBS 0.006695f
C493 B.n453 VSUBS 0.006695f
C494 B.n454 VSUBS 0.006695f
C495 B.n455 VSUBS 0.006695f
C496 B.n456 VSUBS 0.006695f
C497 B.n457 VSUBS 0.006695f
C498 B.n458 VSUBS 0.006695f
C499 B.n459 VSUBS 0.006695f
C500 B.n460 VSUBS 0.006695f
C501 B.n461 VSUBS 0.006695f
C502 B.n462 VSUBS 0.006695f
C503 B.n463 VSUBS 0.006695f
C504 B.n464 VSUBS 0.006695f
C505 B.n465 VSUBS 0.006695f
C506 B.n466 VSUBS 0.006695f
C507 B.n467 VSUBS 0.006695f
C508 B.n468 VSUBS 0.006695f
C509 B.n469 VSUBS 0.006695f
C510 B.n470 VSUBS 0.006695f
C511 B.n471 VSUBS 0.006695f
C512 B.n472 VSUBS 0.006695f
C513 B.n473 VSUBS 0.006695f
C514 B.n474 VSUBS 0.006695f
C515 B.n475 VSUBS 0.006695f
C516 B.n476 VSUBS 0.006695f
C517 B.n477 VSUBS 0.006695f
C518 B.n478 VSUBS 0.006695f
C519 B.n479 VSUBS 0.006695f
C520 B.n480 VSUBS 0.006695f
C521 B.n481 VSUBS 0.006695f
C522 B.n482 VSUBS 0.006695f
C523 B.n483 VSUBS 0.006695f
C524 B.n484 VSUBS 0.006695f
C525 B.n485 VSUBS 0.006695f
C526 B.n486 VSUBS 0.006695f
C527 B.n487 VSUBS 0.006695f
C528 B.n488 VSUBS 0.006695f
C529 B.n489 VSUBS 0.006695f
C530 B.n490 VSUBS 0.006695f
C531 B.n491 VSUBS 0.006695f
C532 B.n492 VSUBS 0.006695f
C533 B.n493 VSUBS 0.006695f
C534 B.n494 VSUBS 0.006695f
C535 B.n495 VSUBS 0.006695f
C536 B.n496 VSUBS 0.006695f
C537 B.n497 VSUBS 0.006695f
C538 B.n498 VSUBS 0.006695f
C539 B.n499 VSUBS 0.006695f
C540 B.n500 VSUBS 0.006695f
C541 B.n501 VSUBS 0.006695f
C542 B.n502 VSUBS 0.006695f
C543 B.n503 VSUBS 0.006695f
C544 B.n504 VSUBS 0.006695f
C545 B.n505 VSUBS 0.006695f
C546 B.n506 VSUBS 0.006695f
C547 B.n507 VSUBS 0.006695f
C548 B.n508 VSUBS 0.006695f
C549 B.n509 VSUBS 0.016167f
C550 B.n510 VSUBS 0.015375f
C551 B.n511 VSUBS 0.015935f
C552 B.n512 VSUBS 0.006695f
C553 B.n513 VSUBS 0.006695f
C554 B.n514 VSUBS 0.006695f
C555 B.n515 VSUBS 0.006695f
C556 B.n516 VSUBS 0.006695f
C557 B.n517 VSUBS 0.006695f
C558 B.n518 VSUBS 0.006695f
C559 B.n519 VSUBS 0.006695f
C560 B.n520 VSUBS 0.006695f
C561 B.n521 VSUBS 0.006695f
C562 B.n522 VSUBS 0.006695f
C563 B.n523 VSUBS 0.006695f
C564 B.n524 VSUBS 0.006695f
C565 B.n525 VSUBS 0.006695f
C566 B.n526 VSUBS 0.006695f
C567 B.n527 VSUBS 0.006695f
C568 B.n528 VSUBS 0.006695f
C569 B.n529 VSUBS 0.006695f
C570 B.n530 VSUBS 0.006695f
C571 B.n531 VSUBS 0.006695f
C572 B.n532 VSUBS 0.006695f
C573 B.n533 VSUBS 0.006695f
C574 B.n534 VSUBS 0.006695f
C575 B.n535 VSUBS 0.006695f
C576 B.n536 VSUBS 0.006695f
C577 B.n537 VSUBS 0.006695f
C578 B.n538 VSUBS 0.006695f
C579 B.n539 VSUBS 0.006695f
C580 B.n540 VSUBS 0.006695f
C581 B.n541 VSUBS 0.006695f
C582 B.n542 VSUBS 0.006695f
C583 B.n543 VSUBS 0.006695f
C584 B.n544 VSUBS 0.006695f
C585 B.n545 VSUBS 0.006695f
C586 B.n546 VSUBS 0.006695f
C587 B.n547 VSUBS 0.006695f
C588 B.n548 VSUBS 0.006695f
C589 B.n549 VSUBS 0.006695f
C590 B.n550 VSUBS 0.006695f
C591 B.n551 VSUBS 0.006695f
C592 B.n552 VSUBS 0.006695f
C593 B.n553 VSUBS 0.006695f
C594 B.n554 VSUBS 0.006695f
C595 B.n555 VSUBS 0.006695f
C596 B.n556 VSUBS 0.006695f
C597 B.n557 VSUBS 0.006695f
C598 B.n558 VSUBS 0.006695f
C599 B.n559 VSUBS 0.006695f
C600 B.n560 VSUBS 0.006695f
C601 B.n561 VSUBS 0.006695f
C602 B.n562 VSUBS 0.006695f
C603 B.n563 VSUBS 0.006695f
C604 B.n564 VSUBS 0.006695f
C605 B.n565 VSUBS 0.006695f
C606 B.n566 VSUBS 0.006695f
C607 B.n567 VSUBS 0.006695f
C608 B.n568 VSUBS 0.006695f
C609 B.n569 VSUBS 0.006695f
C610 B.n570 VSUBS 0.006695f
C611 B.n571 VSUBS 0.006695f
C612 B.n572 VSUBS 0.006695f
C613 B.n573 VSUBS 0.006695f
C614 B.n574 VSUBS 0.006695f
C615 B.n575 VSUBS 0.006695f
C616 B.n576 VSUBS 0.006695f
C617 B.n577 VSUBS 0.006695f
C618 B.n578 VSUBS 0.006695f
C619 B.n579 VSUBS 0.006695f
C620 B.n580 VSUBS 0.006695f
C621 B.n581 VSUBS 0.006695f
C622 B.n582 VSUBS 0.006695f
C623 B.n583 VSUBS 0.006695f
C624 B.n584 VSUBS 0.006695f
C625 B.n585 VSUBS 0.006695f
C626 B.n586 VSUBS 0.006695f
C627 B.n587 VSUBS 0.006695f
C628 B.n588 VSUBS 0.006695f
C629 B.n589 VSUBS 0.006695f
C630 B.n590 VSUBS 0.006695f
C631 B.n591 VSUBS 0.006695f
C632 B.n592 VSUBS 0.006695f
C633 B.n593 VSUBS 0.006695f
C634 B.n594 VSUBS 0.006695f
C635 B.n595 VSUBS 0.006695f
C636 B.n596 VSUBS 0.006695f
C637 B.n597 VSUBS 0.006695f
C638 B.n598 VSUBS 0.006695f
C639 B.n599 VSUBS 0.004628f
C640 B.n600 VSUBS 0.006695f
C641 B.n601 VSUBS 0.006695f
C642 B.n602 VSUBS 0.005415f
C643 B.n603 VSUBS 0.006695f
C644 B.n604 VSUBS 0.006695f
C645 B.n605 VSUBS 0.006695f
C646 B.n606 VSUBS 0.006695f
C647 B.n607 VSUBS 0.006695f
C648 B.n608 VSUBS 0.006695f
C649 B.n609 VSUBS 0.006695f
C650 B.n610 VSUBS 0.006695f
C651 B.n611 VSUBS 0.006695f
C652 B.n612 VSUBS 0.006695f
C653 B.n613 VSUBS 0.006695f
C654 B.n614 VSUBS 0.005415f
C655 B.n615 VSUBS 0.015512f
C656 B.n616 VSUBS 0.004628f
C657 B.n617 VSUBS 0.006695f
C658 B.n618 VSUBS 0.006695f
C659 B.n619 VSUBS 0.006695f
C660 B.n620 VSUBS 0.006695f
C661 B.n621 VSUBS 0.006695f
C662 B.n622 VSUBS 0.006695f
C663 B.n623 VSUBS 0.006695f
C664 B.n624 VSUBS 0.006695f
C665 B.n625 VSUBS 0.006695f
C666 B.n626 VSUBS 0.006695f
C667 B.n627 VSUBS 0.006695f
C668 B.n628 VSUBS 0.006695f
C669 B.n629 VSUBS 0.006695f
C670 B.n630 VSUBS 0.006695f
C671 B.n631 VSUBS 0.006695f
C672 B.n632 VSUBS 0.006695f
C673 B.n633 VSUBS 0.006695f
C674 B.n634 VSUBS 0.006695f
C675 B.n635 VSUBS 0.006695f
C676 B.n636 VSUBS 0.006695f
C677 B.n637 VSUBS 0.006695f
C678 B.n638 VSUBS 0.006695f
C679 B.n639 VSUBS 0.006695f
C680 B.n640 VSUBS 0.006695f
C681 B.n641 VSUBS 0.006695f
C682 B.n642 VSUBS 0.006695f
C683 B.n643 VSUBS 0.006695f
C684 B.n644 VSUBS 0.006695f
C685 B.n645 VSUBS 0.006695f
C686 B.n646 VSUBS 0.006695f
C687 B.n647 VSUBS 0.006695f
C688 B.n648 VSUBS 0.006695f
C689 B.n649 VSUBS 0.006695f
C690 B.n650 VSUBS 0.006695f
C691 B.n651 VSUBS 0.006695f
C692 B.n652 VSUBS 0.006695f
C693 B.n653 VSUBS 0.006695f
C694 B.n654 VSUBS 0.006695f
C695 B.n655 VSUBS 0.006695f
C696 B.n656 VSUBS 0.006695f
C697 B.n657 VSUBS 0.006695f
C698 B.n658 VSUBS 0.006695f
C699 B.n659 VSUBS 0.006695f
C700 B.n660 VSUBS 0.006695f
C701 B.n661 VSUBS 0.006695f
C702 B.n662 VSUBS 0.006695f
C703 B.n663 VSUBS 0.006695f
C704 B.n664 VSUBS 0.006695f
C705 B.n665 VSUBS 0.006695f
C706 B.n666 VSUBS 0.006695f
C707 B.n667 VSUBS 0.006695f
C708 B.n668 VSUBS 0.006695f
C709 B.n669 VSUBS 0.006695f
C710 B.n670 VSUBS 0.006695f
C711 B.n671 VSUBS 0.006695f
C712 B.n672 VSUBS 0.006695f
C713 B.n673 VSUBS 0.006695f
C714 B.n674 VSUBS 0.006695f
C715 B.n675 VSUBS 0.006695f
C716 B.n676 VSUBS 0.006695f
C717 B.n677 VSUBS 0.006695f
C718 B.n678 VSUBS 0.006695f
C719 B.n679 VSUBS 0.006695f
C720 B.n680 VSUBS 0.006695f
C721 B.n681 VSUBS 0.006695f
C722 B.n682 VSUBS 0.006695f
C723 B.n683 VSUBS 0.006695f
C724 B.n684 VSUBS 0.006695f
C725 B.n685 VSUBS 0.006695f
C726 B.n686 VSUBS 0.006695f
C727 B.n687 VSUBS 0.006695f
C728 B.n688 VSUBS 0.006695f
C729 B.n689 VSUBS 0.006695f
C730 B.n690 VSUBS 0.006695f
C731 B.n691 VSUBS 0.006695f
C732 B.n692 VSUBS 0.006695f
C733 B.n693 VSUBS 0.006695f
C734 B.n694 VSUBS 0.006695f
C735 B.n695 VSUBS 0.006695f
C736 B.n696 VSUBS 0.006695f
C737 B.n697 VSUBS 0.006695f
C738 B.n698 VSUBS 0.006695f
C739 B.n699 VSUBS 0.006695f
C740 B.n700 VSUBS 0.006695f
C741 B.n701 VSUBS 0.006695f
C742 B.n702 VSUBS 0.006695f
C743 B.n703 VSUBS 0.006695f
C744 B.n704 VSUBS 0.015935f
C745 B.n705 VSUBS 0.015935f
C746 B.n706 VSUBS 0.015375f
C747 B.n707 VSUBS 0.006695f
C748 B.n708 VSUBS 0.006695f
C749 B.n709 VSUBS 0.006695f
C750 B.n710 VSUBS 0.006695f
C751 B.n711 VSUBS 0.006695f
C752 B.n712 VSUBS 0.006695f
C753 B.n713 VSUBS 0.006695f
C754 B.n714 VSUBS 0.006695f
C755 B.n715 VSUBS 0.006695f
C756 B.n716 VSUBS 0.006695f
C757 B.n717 VSUBS 0.006695f
C758 B.n718 VSUBS 0.006695f
C759 B.n719 VSUBS 0.006695f
C760 B.n720 VSUBS 0.006695f
C761 B.n721 VSUBS 0.006695f
C762 B.n722 VSUBS 0.006695f
C763 B.n723 VSUBS 0.006695f
C764 B.n724 VSUBS 0.006695f
C765 B.n725 VSUBS 0.006695f
C766 B.n726 VSUBS 0.006695f
C767 B.n727 VSUBS 0.006695f
C768 B.n728 VSUBS 0.006695f
C769 B.n729 VSUBS 0.006695f
C770 B.n730 VSUBS 0.006695f
C771 B.n731 VSUBS 0.006695f
C772 B.n732 VSUBS 0.006695f
C773 B.n733 VSUBS 0.006695f
C774 B.n734 VSUBS 0.006695f
C775 B.n735 VSUBS 0.006695f
C776 B.n736 VSUBS 0.006695f
C777 B.n737 VSUBS 0.006695f
C778 B.n738 VSUBS 0.006695f
C779 B.n739 VSUBS 0.006695f
C780 B.n740 VSUBS 0.006695f
C781 B.n741 VSUBS 0.006695f
C782 B.n742 VSUBS 0.006695f
C783 B.n743 VSUBS 0.006695f
C784 B.n744 VSUBS 0.006695f
C785 B.n745 VSUBS 0.006695f
C786 B.n746 VSUBS 0.006695f
C787 B.n747 VSUBS 0.015161f
C788 VDD2.n0 VSUBS 0.03029f
C789 VDD2.n1 VSUBS 0.02833f
C790 VDD2.n2 VSUBS 0.015223f
C791 VDD2.n3 VSUBS 0.035983f
C792 VDD2.n4 VSUBS 0.016119f
C793 VDD2.n5 VSUBS 0.02833f
C794 VDD2.n6 VSUBS 0.015223f
C795 VDD2.n7 VSUBS 0.035983f
C796 VDD2.n8 VSUBS 0.016119f
C797 VDD2.n9 VSUBS 0.02833f
C798 VDD2.n10 VSUBS 0.015671f
C799 VDD2.n11 VSUBS 0.035983f
C800 VDD2.n12 VSUBS 0.016119f
C801 VDD2.n13 VSUBS 0.02833f
C802 VDD2.n14 VSUBS 0.015223f
C803 VDD2.n15 VSUBS 0.035983f
C804 VDD2.n16 VSUBS 0.016119f
C805 VDD2.n17 VSUBS 0.02833f
C806 VDD2.n18 VSUBS 0.015223f
C807 VDD2.n19 VSUBS 0.035983f
C808 VDD2.n20 VSUBS 0.016119f
C809 VDD2.n21 VSUBS 0.02833f
C810 VDD2.n22 VSUBS 0.015223f
C811 VDD2.n23 VSUBS 0.035983f
C812 VDD2.n24 VSUBS 0.016119f
C813 VDD2.n25 VSUBS 0.02833f
C814 VDD2.n26 VSUBS 0.015223f
C815 VDD2.n27 VSUBS 0.035983f
C816 VDD2.n28 VSUBS 0.016119f
C817 VDD2.n29 VSUBS 0.02833f
C818 VDD2.n30 VSUBS 0.015223f
C819 VDD2.n31 VSUBS 0.026987f
C820 VDD2.n32 VSUBS 0.022891f
C821 VDD2.t0 VSUBS 0.077256f
C822 VDD2.n33 VSUBS 0.226277f
C823 VDD2.n34 VSUBS 2.21794f
C824 VDD2.n35 VSUBS 0.015223f
C825 VDD2.n36 VSUBS 0.016119f
C826 VDD2.n37 VSUBS 0.035983f
C827 VDD2.n38 VSUBS 0.035983f
C828 VDD2.n39 VSUBS 0.016119f
C829 VDD2.n40 VSUBS 0.015223f
C830 VDD2.n41 VSUBS 0.02833f
C831 VDD2.n42 VSUBS 0.02833f
C832 VDD2.n43 VSUBS 0.015223f
C833 VDD2.n44 VSUBS 0.016119f
C834 VDD2.n45 VSUBS 0.035983f
C835 VDD2.n46 VSUBS 0.035983f
C836 VDD2.n47 VSUBS 0.016119f
C837 VDD2.n48 VSUBS 0.015223f
C838 VDD2.n49 VSUBS 0.02833f
C839 VDD2.n50 VSUBS 0.02833f
C840 VDD2.n51 VSUBS 0.015223f
C841 VDD2.n52 VSUBS 0.016119f
C842 VDD2.n53 VSUBS 0.035983f
C843 VDD2.n54 VSUBS 0.035983f
C844 VDD2.n55 VSUBS 0.016119f
C845 VDD2.n56 VSUBS 0.015223f
C846 VDD2.n57 VSUBS 0.02833f
C847 VDD2.n58 VSUBS 0.02833f
C848 VDD2.n59 VSUBS 0.015223f
C849 VDD2.n60 VSUBS 0.016119f
C850 VDD2.n61 VSUBS 0.035983f
C851 VDD2.n62 VSUBS 0.035983f
C852 VDD2.n63 VSUBS 0.016119f
C853 VDD2.n64 VSUBS 0.015223f
C854 VDD2.n65 VSUBS 0.02833f
C855 VDD2.n66 VSUBS 0.02833f
C856 VDD2.n67 VSUBS 0.015223f
C857 VDD2.n68 VSUBS 0.016119f
C858 VDD2.n69 VSUBS 0.035983f
C859 VDD2.n70 VSUBS 0.035983f
C860 VDD2.n71 VSUBS 0.016119f
C861 VDD2.n72 VSUBS 0.015223f
C862 VDD2.n73 VSUBS 0.02833f
C863 VDD2.n74 VSUBS 0.02833f
C864 VDD2.n75 VSUBS 0.015223f
C865 VDD2.n76 VSUBS 0.015223f
C866 VDD2.n77 VSUBS 0.016119f
C867 VDD2.n78 VSUBS 0.035983f
C868 VDD2.n79 VSUBS 0.035983f
C869 VDD2.n80 VSUBS 0.035983f
C870 VDD2.n81 VSUBS 0.015671f
C871 VDD2.n82 VSUBS 0.015223f
C872 VDD2.n83 VSUBS 0.02833f
C873 VDD2.n84 VSUBS 0.02833f
C874 VDD2.n85 VSUBS 0.015223f
C875 VDD2.n86 VSUBS 0.016119f
C876 VDD2.n87 VSUBS 0.035983f
C877 VDD2.n88 VSUBS 0.035983f
C878 VDD2.n89 VSUBS 0.016119f
C879 VDD2.n90 VSUBS 0.015223f
C880 VDD2.n91 VSUBS 0.02833f
C881 VDD2.n92 VSUBS 0.02833f
C882 VDD2.n93 VSUBS 0.015223f
C883 VDD2.n94 VSUBS 0.016119f
C884 VDD2.n95 VSUBS 0.035983f
C885 VDD2.n96 VSUBS 0.084253f
C886 VDD2.n97 VSUBS 0.016119f
C887 VDD2.n98 VSUBS 0.015223f
C888 VDD2.n99 VSUBS 0.063162f
C889 VDD2.n100 VSUBS 1.12797f
C890 VDD2.n101 VSUBS 0.03029f
C891 VDD2.n102 VSUBS 0.02833f
C892 VDD2.n103 VSUBS 0.015223f
C893 VDD2.n104 VSUBS 0.035983f
C894 VDD2.n105 VSUBS 0.016119f
C895 VDD2.n106 VSUBS 0.02833f
C896 VDD2.n107 VSUBS 0.015223f
C897 VDD2.n108 VSUBS 0.035983f
C898 VDD2.n109 VSUBS 0.016119f
C899 VDD2.n110 VSUBS 0.02833f
C900 VDD2.n111 VSUBS 0.015671f
C901 VDD2.n112 VSUBS 0.035983f
C902 VDD2.n113 VSUBS 0.015223f
C903 VDD2.n114 VSUBS 0.016119f
C904 VDD2.n115 VSUBS 0.02833f
C905 VDD2.n116 VSUBS 0.015223f
C906 VDD2.n117 VSUBS 0.035983f
C907 VDD2.n118 VSUBS 0.016119f
C908 VDD2.n119 VSUBS 0.02833f
C909 VDD2.n120 VSUBS 0.015223f
C910 VDD2.n121 VSUBS 0.035983f
C911 VDD2.n122 VSUBS 0.016119f
C912 VDD2.n123 VSUBS 0.02833f
C913 VDD2.n124 VSUBS 0.015223f
C914 VDD2.n125 VSUBS 0.035983f
C915 VDD2.n126 VSUBS 0.016119f
C916 VDD2.n127 VSUBS 0.02833f
C917 VDD2.n128 VSUBS 0.015223f
C918 VDD2.n129 VSUBS 0.035983f
C919 VDD2.n130 VSUBS 0.016119f
C920 VDD2.n131 VSUBS 0.02833f
C921 VDD2.n132 VSUBS 0.015223f
C922 VDD2.n133 VSUBS 0.026987f
C923 VDD2.n134 VSUBS 0.022891f
C924 VDD2.t1 VSUBS 0.077256f
C925 VDD2.n135 VSUBS 0.226277f
C926 VDD2.n136 VSUBS 2.21794f
C927 VDD2.n137 VSUBS 0.015223f
C928 VDD2.n138 VSUBS 0.016119f
C929 VDD2.n139 VSUBS 0.035983f
C930 VDD2.n140 VSUBS 0.035983f
C931 VDD2.n141 VSUBS 0.016119f
C932 VDD2.n142 VSUBS 0.015223f
C933 VDD2.n143 VSUBS 0.02833f
C934 VDD2.n144 VSUBS 0.02833f
C935 VDD2.n145 VSUBS 0.015223f
C936 VDD2.n146 VSUBS 0.016119f
C937 VDD2.n147 VSUBS 0.035983f
C938 VDD2.n148 VSUBS 0.035983f
C939 VDD2.n149 VSUBS 0.016119f
C940 VDD2.n150 VSUBS 0.015223f
C941 VDD2.n151 VSUBS 0.02833f
C942 VDD2.n152 VSUBS 0.02833f
C943 VDD2.n153 VSUBS 0.015223f
C944 VDD2.n154 VSUBS 0.016119f
C945 VDD2.n155 VSUBS 0.035983f
C946 VDD2.n156 VSUBS 0.035983f
C947 VDD2.n157 VSUBS 0.016119f
C948 VDD2.n158 VSUBS 0.015223f
C949 VDD2.n159 VSUBS 0.02833f
C950 VDD2.n160 VSUBS 0.02833f
C951 VDD2.n161 VSUBS 0.015223f
C952 VDD2.n162 VSUBS 0.016119f
C953 VDD2.n163 VSUBS 0.035983f
C954 VDD2.n164 VSUBS 0.035983f
C955 VDD2.n165 VSUBS 0.016119f
C956 VDD2.n166 VSUBS 0.015223f
C957 VDD2.n167 VSUBS 0.02833f
C958 VDD2.n168 VSUBS 0.02833f
C959 VDD2.n169 VSUBS 0.015223f
C960 VDD2.n170 VSUBS 0.016119f
C961 VDD2.n171 VSUBS 0.035983f
C962 VDD2.n172 VSUBS 0.035983f
C963 VDD2.n173 VSUBS 0.016119f
C964 VDD2.n174 VSUBS 0.015223f
C965 VDD2.n175 VSUBS 0.02833f
C966 VDD2.n176 VSUBS 0.02833f
C967 VDD2.n177 VSUBS 0.015223f
C968 VDD2.n178 VSUBS 0.016119f
C969 VDD2.n179 VSUBS 0.035983f
C970 VDD2.n180 VSUBS 0.035983f
C971 VDD2.n181 VSUBS 0.035983f
C972 VDD2.n182 VSUBS 0.015671f
C973 VDD2.n183 VSUBS 0.015223f
C974 VDD2.n184 VSUBS 0.02833f
C975 VDD2.n185 VSUBS 0.02833f
C976 VDD2.n186 VSUBS 0.015223f
C977 VDD2.n187 VSUBS 0.016119f
C978 VDD2.n188 VSUBS 0.035983f
C979 VDD2.n189 VSUBS 0.035983f
C980 VDD2.n190 VSUBS 0.016119f
C981 VDD2.n191 VSUBS 0.015223f
C982 VDD2.n192 VSUBS 0.02833f
C983 VDD2.n193 VSUBS 0.02833f
C984 VDD2.n194 VSUBS 0.015223f
C985 VDD2.n195 VSUBS 0.016119f
C986 VDD2.n196 VSUBS 0.035983f
C987 VDD2.n197 VSUBS 0.084253f
C988 VDD2.n198 VSUBS 0.016119f
C989 VDD2.n199 VSUBS 0.015223f
C990 VDD2.n200 VSUBS 0.063162f
C991 VDD2.n201 VSUBS 0.061751f
C992 VDD2.n202 VSUBS 4.21281f
C993 VN.t1 VSUBS 5.27204f
C994 VN.t0 VSUBS 5.99766f
C995 VDD1.n0 VSUBS 0.029893f
C996 VDD1.n1 VSUBS 0.027959f
C997 VDD1.n2 VSUBS 0.015024f
C998 VDD1.n3 VSUBS 0.035511f
C999 VDD1.n4 VSUBS 0.015908f
C1000 VDD1.n5 VSUBS 0.027959f
C1001 VDD1.n6 VSUBS 0.015024f
C1002 VDD1.n7 VSUBS 0.035511f
C1003 VDD1.n8 VSUBS 0.015908f
C1004 VDD1.n9 VSUBS 0.027959f
C1005 VDD1.n10 VSUBS 0.015466f
C1006 VDD1.n11 VSUBS 0.035511f
C1007 VDD1.n12 VSUBS 0.015024f
C1008 VDD1.n13 VSUBS 0.015908f
C1009 VDD1.n14 VSUBS 0.027959f
C1010 VDD1.n15 VSUBS 0.015024f
C1011 VDD1.n16 VSUBS 0.035511f
C1012 VDD1.n17 VSUBS 0.015908f
C1013 VDD1.n18 VSUBS 0.027959f
C1014 VDD1.n19 VSUBS 0.015024f
C1015 VDD1.n20 VSUBS 0.035511f
C1016 VDD1.n21 VSUBS 0.015908f
C1017 VDD1.n22 VSUBS 0.027959f
C1018 VDD1.n23 VSUBS 0.015024f
C1019 VDD1.n24 VSUBS 0.035511f
C1020 VDD1.n25 VSUBS 0.015908f
C1021 VDD1.n26 VSUBS 0.027959f
C1022 VDD1.n27 VSUBS 0.015024f
C1023 VDD1.n28 VSUBS 0.035511f
C1024 VDD1.n29 VSUBS 0.015908f
C1025 VDD1.n30 VSUBS 0.027959f
C1026 VDD1.n31 VSUBS 0.015024f
C1027 VDD1.n32 VSUBS 0.026633f
C1028 VDD1.n33 VSUBS 0.02259f
C1029 VDD1.t1 VSUBS 0.076243f
C1030 VDD1.n34 VSUBS 0.22331f
C1031 VDD1.n35 VSUBS 2.18885f
C1032 VDD1.n36 VSUBS 0.015024f
C1033 VDD1.n37 VSUBS 0.015908f
C1034 VDD1.n38 VSUBS 0.035511f
C1035 VDD1.n39 VSUBS 0.035511f
C1036 VDD1.n40 VSUBS 0.015908f
C1037 VDD1.n41 VSUBS 0.015024f
C1038 VDD1.n42 VSUBS 0.027959f
C1039 VDD1.n43 VSUBS 0.027959f
C1040 VDD1.n44 VSUBS 0.015024f
C1041 VDD1.n45 VSUBS 0.015908f
C1042 VDD1.n46 VSUBS 0.035511f
C1043 VDD1.n47 VSUBS 0.035511f
C1044 VDD1.n48 VSUBS 0.015908f
C1045 VDD1.n49 VSUBS 0.015024f
C1046 VDD1.n50 VSUBS 0.027959f
C1047 VDD1.n51 VSUBS 0.027959f
C1048 VDD1.n52 VSUBS 0.015024f
C1049 VDD1.n53 VSUBS 0.015908f
C1050 VDD1.n54 VSUBS 0.035511f
C1051 VDD1.n55 VSUBS 0.035511f
C1052 VDD1.n56 VSUBS 0.015908f
C1053 VDD1.n57 VSUBS 0.015024f
C1054 VDD1.n58 VSUBS 0.027959f
C1055 VDD1.n59 VSUBS 0.027959f
C1056 VDD1.n60 VSUBS 0.015024f
C1057 VDD1.n61 VSUBS 0.015908f
C1058 VDD1.n62 VSUBS 0.035511f
C1059 VDD1.n63 VSUBS 0.035511f
C1060 VDD1.n64 VSUBS 0.015908f
C1061 VDD1.n65 VSUBS 0.015024f
C1062 VDD1.n66 VSUBS 0.027959f
C1063 VDD1.n67 VSUBS 0.027959f
C1064 VDD1.n68 VSUBS 0.015024f
C1065 VDD1.n69 VSUBS 0.015908f
C1066 VDD1.n70 VSUBS 0.035511f
C1067 VDD1.n71 VSUBS 0.035511f
C1068 VDD1.n72 VSUBS 0.015908f
C1069 VDD1.n73 VSUBS 0.015024f
C1070 VDD1.n74 VSUBS 0.027959f
C1071 VDD1.n75 VSUBS 0.027959f
C1072 VDD1.n76 VSUBS 0.015024f
C1073 VDD1.n77 VSUBS 0.015908f
C1074 VDD1.n78 VSUBS 0.035511f
C1075 VDD1.n79 VSUBS 0.035511f
C1076 VDD1.n80 VSUBS 0.035511f
C1077 VDD1.n81 VSUBS 0.015466f
C1078 VDD1.n82 VSUBS 0.015024f
C1079 VDD1.n83 VSUBS 0.027959f
C1080 VDD1.n84 VSUBS 0.027959f
C1081 VDD1.n85 VSUBS 0.015024f
C1082 VDD1.n86 VSUBS 0.015908f
C1083 VDD1.n87 VSUBS 0.035511f
C1084 VDD1.n88 VSUBS 0.035511f
C1085 VDD1.n89 VSUBS 0.015908f
C1086 VDD1.n90 VSUBS 0.015024f
C1087 VDD1.n91 VSUBS 0.027959f
C1088 VDD1.n92 VSUBS 0.027959f
C1089 VDD1.n93 VSUBS 0.015024f
C1090 VDD1.n94 VSUBS 0.015908f
C1091 VDD1.n95 VSUBS 0.035511f
C1092 VDD1.n96 VSUBS 0.083148f
C1093 VDD1.n97 VSUBS 0.015908f
C1094 VDD1.n98 VSUBS 0.015024f
C1095 VDD1.n99 VSUBS 0.062334f
C1096 VDD1.n100 VSUBS 0.062792f
C1097 VDD1.n101 VSUBS 0.029893f
C1098 VDD1.n102 VSUBS 0.027959f
C1099 VDD1.n103 VSUBS 0.015024f
C1100 VDD1.n104 VSUBS 0.035511f
C1101 VDD1.n105 VSUBS 0.015908f
C1102 VDD1.n106 VSUBS 0.027959f
C1103 VDD1.n107 VSUBS 0.015024f
C1104 VDD1.n108 VSUBS 0.035511f
C1105 VDD1.n109 VSUBS 0.015908f
C1106 VDD1.n110 VSUBS 0.027959f
C1107 VDD1.n111 VSUBS 0.015466f
C1108 VDD1.n112 VSUBS 0.035511f
C1109 VDD1.n113 VSUBS 0.015908f
C1110 VDD1.n114 VSUBS 0.027959f
C1111 VDD1.n115 VSUBS 0.015024f
C1112 VDD1.n116 VSUBS 0.035511f
C1113 VDD1.n117 VSUBS 0.015908f
C1114 VDD1.n118 VSUBS 0.027959f
C1115 VDD1.n119 VSUBS 0.015024f
C1116 VDD1.n120 VSUBS 0.035511f
C1117 VDD1.n121 VSUBS 0.015908f
C1118 VDD1.n122 VSUBS 0.027959f
C1119 VDD1.n123 VSUBS 0.015024f
C1120 VDD1.n124 VSUBS 0.035511f
C1121 VDD1.n125 VSUBS 0.015908f
C1122 VDD1.n126 VSUBS 0.027959f
C1123 VDD1.n127 VSUBS 0.015024f
C1124 VDD1.n128 VSUBS 0.035511f
C1125 VDD1.n129 VSUBS 0.015908f
C1126 VDD1.n130 VSUBS 0.027959f
C1127 VDD1.n131 VSUBS 0.015024f
C1128 VDD1.n132 VSUBS 0.026633f
C1129 VDD1.n133 VSUBS 0.02259f
C1130 VDD1.t0 VSUBS 0.076243f
C1131 VDD1.n134 VSUBS 0.22331f
C1132 VDD1.n135 VSUBS 2.18885f
C1133 VDD1.n136 VSUBS 0.015024f
C1134 VDD1.n137 VSUBS 0.015908f
C1135 VDD1.n138 VSUBS 0.035511f
C1136 VDD1.n139 VSUBS 0.035511f
C1137 VDD1.n140 VSUBS 0.015908f
C1138 VDD1.n141 VSUBS 0.015024f
C1139 VDD1.n142 VSUBS 0.027959f
C1140 VDD1.n143 VSUBS 0.027959f
C1141 VDD1.n144 VSUBS 0.015024f
C1142 VDD1.n145 VSUBS 0.015908f
C1143 VDD1.n146 VSUBS 0.035511f
C1144 VDD1.n147 VSUBS 0.035511f
C1145 VDD1.n148 VSUBS 0.015908f
C1146 VDD1.n149 VSUBS 0.015024f
C1147 VDD1.n150 VSUBS 0.027959f
C1148 VDD1.n151 VSUBS 0.027959f
C1149 VDD1.n152 VSUBS 0.015024f
C1150 VDD1.n153 VSUBS 0.015908f
C1151 VDD1.n154 VSUBS 0.035511f
C1152 VDD1.n155 VSUBS 0.035511f
C1153 VDD1.n156 VSUBS 0.015908f
C1154 VDD1.n157 VSUBS 0.015024f
C1155 VDD1.n158 VSUBS 0.027959f
C1156 VDD1.n159 VSUBS 0.027959f
C1157 VDD1.n160 VSUBS 0.015024f
C1158 VDD1.n161 VSUBS 0.015908f
C1159 VDD1.n162 VSUBS 0.035511f
C1160 VDD1.n163 VSUBS 0.035511f
C1161 VDD1.n164 VSUBS 0.015908f
C1162 VDD1.n165 VSUBS 0.015024f
C1163 VDD1.n166 VSUBS 0.027959f
C1164 VDD1.n167 VSUBS 0.027959f
C1165 VDD1.n168 VSUBS 0.015024f
C1166 VDD1.n169 VSUBS 0.015908f
C1167 VDD1.n170 VSUBS 0.035511f
C1168 VDD1.n171 VSUBS 0.035511f
C1169 VDD1.n172 VSUBS 0.015908f
C1170 VDD1.n173 VSUBS 0.015024f
C1171 VDD1.n174 VSUBS 0.027959f
C1172 VDD1.n175 VSUBS 0.027959f
C1173 VDD1.n176 VSUBS 0.015024f
C1174 VDD1.n177 VSUBS 0.015024f
C1175 VDD1.n178 VSUBS 0.015908f
C1176 VDD1.n179 VSUBS 0.035511f
C1177 VDD1.n180 VSUBS 0.035511f
C1178 VDD1.n181 VSUBS 0.035511f
C1179 VDD1.n182 VSUBS 0.015466f
C1180 VDD1.n183 VSUBS 0.015024f
C1181 VDD1.n184 VSUBS 0.027959f
C1182 VDD1.n185 VSUBS 0.027959f
C1183 VDD1.n186 VSUBS 0.015024f
C1184 VDD1.n187 VSUBS 0.015908f
C1185 VDD1.n188 VSUBS 0.035511f
C1186 VDD1.n189 VSUBS 0.035511f
C1187 VDD1.n190 VSUBS 0.015908f
C1188 VDD1.n191 VSUBS 0.015024f
C1189 VDD1.n192 VSUBS 0.027959f
C1190 VDD1.n193 VSUBS 0.027959f
C1191 VDD1.n194 VSUBS 0.015024f
C1192 VDD1.n195 VSUBS 0.015908f
C1193 VDD1.n196 VSUBS 0.035511f
C1194 VDD1.n197 VSUBS 0.083148f
C1195 VDD1.n198 VSUBS 0.015908f
C1196 VDD1.n199 VSUBS 0.015024f
C1197 VDD1.n200 VSUBS 0.062334f
C1198 VDD1.n201 VSUBS 1.17696f
C1199 VTAIL.n0 VSUBS 0.030276f
C1200 VTAIL.n1 VSUBS 0.028317f
C1201 VTAIL.n2 VSUBS 0.015217f
C1202 VTAIL.n3 VSUBS 0.035966f
C1203 VTAIL.n4 VSUBS 0.016112f
C1204 VTAIL.n5 VSUBS 0.028317f
C1205 VTAIL.n6 VSUBS 0.015217f
C1206 VTAIL.n7 VSUBS 0.035966f
C1207 VTAIL.n8 VSUBS 0.016112f
C1208 VTAIL.n9 VSUBS 0.028317f
C1209 VTAIL.n10 VSUBS 0.015664f
C1210 VTAIL.n11 VSUBS 0.035966f
C1211 VTAIL.n12 VSUBS 0.016112f
C1212 VTAIL.n13 VSUBS 0.028317f
C1213 VTAIL.n14 VSUBS 0.015217f
C1214 VTAIL.n15 VSUBS 0.035966f
C1215 VTAIL.n16 VSUBS 0.016112f
C1216 VTAIL.n17 VSUBS 0.028317f
C1217 VTAIL.n18 VSUBS 0.015217f
C1218 VTAIL.n19 VSUBS 0.035966f
C1219 VTAIL.n20 VSUBS 0.016112f
C1220 VTAIL.n21 VSUBS 0.028317f
C1221 VTAIL.n22 VSUBS 0.015217f
C1222 VTAIL.n23 VSUBS 0.035966f
C1223 VTAIL.n24 VSUBS 0.016112f
C1224 VTAIL.n25 VSUBS 0.028317f
C1225 VTAIL.n26 VSUBS 0.015217f
C1226 VTAIL.n27 VSUBS 0.035966f
C1227 VTAIL.n28 VSUBS 0.016112f
C1228 VTAIL.n29 VSUBS 0.028317f
C1229 VTAIL.n30 VSUBS 0.015217f
C1230 VTAIL.n31 VSUBS 0.026975f
C1231 VTAIL.n32 VSUBS 0.02288f
C1232 VTAIL.t2 VSUBS 0.077221f
C1233 VTAIL.n33 VSUBS 0.226174f
C1234 VTAIL.n34 VSUBS 2.21693f
C1235 VTAIL.n35 VSUBS 0.015217f
C1236 VTAIL.n36 VSUBS 0.016112f
C1237 VTAIL.n37 VSUBS 0.035966f
C1238 VTAIL.n38 VSUBS 0.035966f
C1239 VTAIL.n39 VSUBS 0.016112f
C1240 VTAIL.n40 VSUBS 0.015217f
C1241 VTAIL.n41 VSUBS 0.028317f
C1242 VTAIL.n42 VSUBS 0.028317f
C1243 VTAIL.n43 VSUBS 0.015217f
C1244 VTAIL.n44 VSUBS 0.016112f
C1245 VTAIL.n45 VSUBS 0.035966f
C1246 VTAIL.n46 VSUBS 0.035966f
C1247 VTAIL.n47 VSUBS 0.016112f
C1248 VTAIL.n48 VSUBS 0.015217f
C1249 VTAIL.n49 VSUBS 0.028317f
C1250 VTAIL.n50 VSUBS 0.028317f
C1251 VTAIL.n51 VSUBS 0.015217f
C1252 VTAIL.n52 VSUBS 0.016112f
C1253 VTAIL.n53 VSUBS 0.035966f
C1254 VTAIL.n54 VSUBS 0.035966f
C1255 VTAIL.n55 VSUBS 0.016112f
C1256 VTAIL.n56 VSUBS 0.015217f
C1257 VTAIL.n57 VSUBS 0.028317f
C1258 VTAIL.n58 VSUBS 0.028317f
C1259 VTAIL.n59 VSUBS 0.015217f
C1260 VTAIL.n60 VSUBS 0.016112f
C1261 VTAIL.n61 VSUBS 0.035966f
C1262 VTAIL.n62 VSUBS 0.035966f
C1263 VTAIL.n63 VSUBS 0.016112f
C1264 VTAIL.n64 VSUBS 0.015217f
C1265 VTAIL.n65 VSUBS 0.028317f
C1266 VTAIL.n66 VSUBS 0.028317f
C1267 VTAIL.n67 VSUBS 0.015217f
C1268 VTAIL.n68 VSUBS 0.016112f
C1269 VTAIL.n69 VSUBS 0.035966f
C1270 VTAIL.n70 VSUBS 0.035966f
C1271 VTAIL.n71 VSUBS 0.016112f
C1272 VTAIL.n72 VSUBS 0.015217f
C1273 VTAIL.n73 VSUBS 0.028317f
C1274 VTAIL.n74 VSUBS 0.028317f
C1275 VTAIL.n75 VSUBS 0.015217f
C1276 VTAIL.n76 VSUBS 0.015217f
C1277 VTAIL.n77 VSUBS 0.016112f
C1278 VTAIL.n78 VSUBS 0.035966f
C1279 VTAIL.n79 VSUBS 0.035966f
C1280 VTAIL.n80 VSUBS 0.035966f
C1281 VTAIL.n81 VSUBS 0.015664f
C1282 VTAIL.n82 VSUBS 0.015217f
C1283 VTAIL.n83 VSUBS 0.028317f
C1284 VTAIL.n84 VSUBS 0.028317f
C1285 VTAIL.n85 VSUBS 0.015217f
C1286 VTAIL.n86 VSUBS 0.016112f
C1287 VTAIL.n87 VSUBS 0.035966f
C1288 VTAIL.n88 VSUBS 0.035966f
C1289 VTAIL.n89 VSUBS 0.016112f
C1290 VTAIL.n90 VSUBS 0.015217f
C1291 VTAIL.n91 VSUBS 0.028317f
C1292 VTAIL.n92 VSUBS 0.028317f
C1293 VTAIL.n93 VSUBS 0.015217f
C1294 VTAIL.n94 VSUBS 0.016112f
C1295 VTAIL.n95 VSUBS 0.035966f
C1296 VTAIL.n96 VSUBS 0.084214f
C1297 VTAIL.n97 VSUBS 0.016112f
C1298 VTAIL.n98 VSUBS 0.015217f
C1299 VTAIL.n99 VSUBS 0.063133f
C1300 VTAIL.n100 VSUBS 0.042151f
C1301 VTAIL.n101 VSUBS 2.45209f
C1302 VTAIL.n102 VSUBS 0.030276f
C1303 VTAIL.n103 VSUBS 0.028317f
C1304 VTAIL.n104 VSUBS 0.015217f
C1305 VTAIL.n105 VSUBS 0.035966f
C1306 VTAIL.n106 VSUBS 0.016112f
C1307 VTAIL.n107 VSUBS 0.028317f
C1308 VTAIL.n108 VSUBS 0.015217f
C1309 VTAIL.n109 VSUBS 0.035966f
C1310 VTAIL.n110 VSUBS 0.016112f
C1311 VTAIL.n111 VSUBS 0.028317f
C1312 VTAIL.n112 VSUBS 0.015664f
C1313 VTAIL.n113 VSUBS 0.035966f
C1314 VTAIL.n114 VSUBS 0.015217f
C1315 VTAIL.n115 VSUBS 0.016112f
C1316 VTAIL.n116 VSUBS 0.028317f
C1317 VTAIL.n117 VSUBS 0.015217f
C1318 VTAIL.n118 VSUBS 0.035966f
C1319 VTAIL.n119 VSUBS 0.016112f
C1320 VTAIL.n120 VSUBS 0.028317f
C1321 VTAIL.n121 VSUBS 0.015217f
C1322 VTAIL.n122 VSUBS 0.035966f
C1323 VTAIL.n123 VSUBS 0.016112f
C1324 VTAIL.n124 VSUBS 0.028317f
C1325 VTAIL.n125 VSUBS 0.015217f
C1326 VTAIL.n126 VSUBS 0.035966f
C1327 VTAIL.n127 VSUBS 0.016112f
C1328 VTAIL.n128 VSUBS 0.028317f
C1329 VTAIL.n129 VSUBS 0.015217f
C1330 VTAIL.n130 VSUBS 0.035966f
C1331 VTAIL.n131 VSUBS 0.016112f
C1332 VTAIL.n132 VSUBS 0.028317f
C1333 VTAIL.n133 VSUBS 0.015217f
C1334 VTAIL.n134 VSUBS 0.026975f
C1335 VTAIL.n135 VSUBS 0.02288f
C1336 VTAIL.t1 VSUBS 0.077221f
C1337 VTAIL.n136 VSUBS 0.226174f
C1338 VTAIL.n137 VSUBS 2.21692f
C1339 VTAIL.n138 VSUBS 0.015217f
C1340 VTAIL.n139 VSUBS 0.016112f
C1341 VTAIL.n140 VSUBS 0.035966f
C1342 VTAIL.n141 VSUBS 0.035966f
C1343 VTAIL.n142 VSUBS 0.016112f
C1344 VTAIL.n143 VSUBS 0.015217f
C1345 VTAIL.n144 VSUBS 0.028317f
C1346 VTAIL.n145 VSUBS 0.028317f
C1347 VTAIL.n146 VSUBS 0.015217f
C1348 VTAIL.n147 VSUBS 0.016112f
C1349 VTAIL.n148 VSUBS 0.035966f
C1350 VTAIL.n149 VSUBS 0.035966f
C1351 VTAIL.n150 VSUBS 0.016112f
C1352 VTAIL.n151 VSUBS 0.015217f
C1353 VTAIL.n152 VSUBS 0.028317f
C1354 VTAIL.n153 VSUBS 0.028317f
C1355 VTAIL.n154 VSUBS 0.015217f
C1356 VTAIL.n155 VSUBS 0.016112f
C1357 VTAIL.n156 VSUBS 0.035966f
C1358 VTAIL.n157 VSUBS 0.035966f
C1359 VTAIL.n158 VSUBS 0.016112f
C1360 VTAIL.n159 VSUBS 0.015217f
C1361 VTAIL.n160 VSUBS 0.028317f
C1362 VTAIL.n161 VSUBS 0.028317f
C1363 VTAIL.n162 VSUBS 0.015217f
C1364 VTAIL.n163 VSUBS 0.016112f
C1365 VTAIL.n164 VSUBS 0.035966f
C1366 VTAIL.n165 VSUBS 0.035966f
C1367 VTAIL.n166 VSUBS 0.016112f
C1368 VTAIL.n167 VSUBS 0.015217f
C1369 VTAIL.n168 VSUBS 0.028317f
C1370 VTAIL.n169 VSUBS 0.028317f
C1371 VTAIL.n170 VSUBS 0.015217f
C1372 VTAIL.n171 VSUBS 0.016112f
C1373 VTAIL.n172 VSUBS 0.035966f
C1374 VTAIL.n173 VSUBS 0.035966f
C1375 VTAIL.n174 VSUBS 0.016112f
C1376 VTAIL.n175 VSUBS 0.015217f
C1377 VTAIL.n176 VSUBS 0.028317f
C1378 VTAIL.n177 VSUBS 0.028317f
C1379 VTAIL.n178 VSUBS 0.015217f
C1380 VTAIL.n179 VSUBS 0.016112f
C1381 VTAIL.n180 VSUBS 0.035966f
C1382 VTAIL.n181 VSUBS 0.035966f
C1383 VTAIL.n182 VSUBS 0.035966f
C1384 VTAIL.n183 VSUBS 0.015664f
C1385 VTAIL.n184 VSUBS 0.015217f
C1386 VTAIL.n185 VSUBS 0.028317f
C1387 VTAIL.n186 VSUBS 0.028317f
C1388 VTAIL.n187 VSUBS 0.015217f
C1389 VTAIL.n188 VSUBS 0.016112f
C1390 VTAIL.n189 VSUBS 0.035966f
C1391 VTAIL.n190 VSUBS 0.035966f
C1392 VTAIL.n191 VSUBS 0.016112f
C1393 VTAIL.n192 VSUBS 0.015217f
C1394 VTAIL.n193 VSUBS 0.028317f
C1395 VTAIL.n194 VSUBS 0.028317f
C1396 VTAIL.n195 VSUBS 0.015217f
C1397 VTAIL.n196 VSUBS 0.016112f
C1398 VTAIL.n197 VSUBS 0.035966f
C1399 VTAIL.n198 VSUBS 0.084214f
C1400 VTAIL.n199 VSUBS 0.016112f
C1401 VTAIL.n200 VSUBS 0.015217f
C1402 VTAIL.n201 VSUBS 0.063133f
C1403 VTAIL.n202 VSUBS 0.042151f
C1404 VTAIL.n203 VSUBS 2.50971f
C1405 VTAIL.n204 VSUBS 0.030276f
C1406 VTAIL.n205 VSUBS 0.028317f
C1407 VTAIL.n206 VSUBS 0.015217f
C1408 VTAIL.n207 VSUBS 0.035966f
C1409 VTAIL.n208 VSUBS 0.016112f
C1410 VTAIL.n209 VSUBS 0.028317f
C1411 VTAIL.n210 VSUBS 0.015217f
C1412 VTAIL.n211 VSUBS 0.035966f
C1413 VTAIL.n212 VSUBS 0.016112f
C1414 VTAIL.n213 VSUBS 0.028317f
C1415 VTAIL.n214 VSUBS 0.015664f
C1416 VTAIL.n215 VSUBS 0.035966f
C1417 VTAIL.n216 VSUBS 0.015217f
C1418 VTAIL.n217 VSUBS 0.016112f
C1419 VTAIL.n218 VSUBS 0.028317f
C1420 VTAIL.n219 VSUBS 0.015217f
C1421 VTAIL.n220 VSUBS 0.035966f
C1422 VTAIL.n221 VSUBS 0.016112f
C1423 VTAIL.n222 VSUBS 0.028317f
C1424 VTAIL.n223 VSUBS 0.015217f
C1425 VTAIL.n224 VSUBS 0.035966f
C1426 VTAIL.n225 VSUBS 0.016112f
C1427 VTAIL.n226 VSUBS 0.028317f
C1428 VTAIL.n227 VSUBS 0.015217f
C1429 VTAIL.n228 VSUBS 0.035966f
C1430 VTAIL.n229 VSUBS 0.016112f
C1431 VTAIL.n230 VSUBS 0.028317f
C1432 VTAIL.n231 VSUBS 0.015217f
C1433 VTAIL.n232 VSUBS 0.035966f
C1434 VTAIL.n233 VSUBS 0.016112f
C1435 VTAIL.n234 VSUBS 0.028317f
C1436 VTAIL.n235 VSUBS 0.015217f
C1437 VTAIL.n236 VSUBS 0.026975f
C1438 VTAIL.n237 VSUBS 0.02288f
C1439 VTAIL.t3 VSUBS 0.077221f
C1440 VTAIL.n238 VSUBS 0.226174f
C1441 VTAIL.n239 VSUBS 2.21692f
C1442 VTAIL.n240 VSUBS 0.015217f
C1443 VTAIL.n241 VSUBS 0.016112f
C1444 VTAIL.n242 VSUBS 0.035966f
C1445 VTAIL.n243 VSUBS 0.035966f
C1446 VTAIL.n244 VSUBS 0.016112f
C1447 VTAIL.n245 VSUBS 0.015217f
C1448 VTAIL.n246 VSUBS 0.028317f
C1449 VTAIL.n247 VSUBS 0.028317f
C1450 VTAIL.n248 VSUBS 0.015217f
C1451 VTAIL.n249 VSUBS 0.016112f
C1452 VTAIL.n250 VSUBS 0.035966f
C1453 VTAIL.n251 VSUBS 0.035966f
C1454 VTAIL.n252 VSUBS 0.016112f
C1455 VTAIL.n253 VSUBS 0.015217f
C1456 VTAIL.n254 VSUBS 0.028317f
C1457 VTAIL.n255 VSUBS 0.028317f
C1458 VTAIL.n256 VSUBS 0.015217f
C1459 VTAIL.n257 VSUBS 0.016112f
C1460 VTAIL.n258 VSUBS 0.035966f
C1461 VTAIL.n259 VSUBS 0.035966f
C1462 VTAIL.n260 VSUBS 0.016112f
C1463 VTAIL.n261 VSUBS 0.015217f
C1464 VTAIL.n262 VSUBS 0.028317f
C1465 VTAIL.n263 VSUBS 0.028317f
C1466 VTAIL.n264 VSUBS 0.015217f
C1467 VTAIL.n265 VSUBS 0.016112f
C1468 VTAIL.n266 VSUBS 0.035966f
C1469 VTAIL.n267 VSUBS 0.035966f
C1470 VTAIL.n268 VSUBS 0.016112f
C1471 VTAIL.n269 VSUBS 0.015217f
C1472 VTAIL.n270 VSUBS 0.028317f
C1473 VTAIL.n271 VSUBS 0.028317f
C1474 VTAIL.n272 VSUBS 0.015217f
C1475 VTAIL.n273 VSUBS 0.016112f
C1476 VTAIL.n274 VSUBS 0.035966f
C1477 VTAIL.n275 VSUBS 0.035966f
C1478 VTAIL.n276 VSUBS 0.016112f
C1479 VTAIL.n277 VSUBS 0.015217f
C1480 VTAIL.n278 VSUBS 0.028317f
C1481 VTAIL.n279 VSUBS 0.028317f
C1482 VTAIL.n280 VSUBS 0.015217f
C1483 VTAIL.n281 VSUBS 0.016112f
C1484 VTAIL.n282 VSUBS 0.035966f
C1485 VTAIL.n283 VSUBS 0.035966f
C1486 VTAIL.n284 VSUBS 0.035966f
C1487 VTAIL.n285 VSUBS 0.015664f
C1488 VTAIL.n286 VSUBS 0.015217f
C1489 VTAIL.n287 VSUBS 0.028317f
C1490 VTAIL.n288 VSUBS 0.028317f
C1491 VTAIL.n289 VSUBS 0.015217f
C1492 VTAIL.n290 VSUBS 0.016112f
C1493 VTAIL.n291 VSUBS 0.035966f
C1494 VTAIL.n292 VSUBS 0.035966f
C1495 VTAIL.n293 VSUBS 0.016112f
C1496 VTAIL.n294 VSUBS 0.015217f
C1497 VTAIL.n295 VSUBS 0.028317f
C1498 VTAIL.n296 VSUBS 0.028317f
C1499 VTAIL.n297 VSUBS 0.015217f
C1500 VTAIL.n298 VSUBS 0.016112f
C1501 VTAIL.n299 VSUBS 0.035966f
C1502 VTAIL.n300 VSUBS 0.084214f
C1503 VTAIL.n301 VSUBS 0.016112f
C1504 VTAIL.n302 VSUBS 0.015217f
C1505 VTAIL.n303 VSUBS 0.063133f
C1506 VTAIL.n304 VSUBS 0.042151f
C1507 VTAIL.n305 VSUBS 2.258f
C1508 VTAIL.n306 VSUBS 0.030276f
C1509 VTAIL.n307 VSUBS 0.028317f
C1510 VTAIL.n308 VSUBS 0.015217f
C1511 VTAIL.n309 VSUBS 0.035966f
C1512 VTAIL.n310 VSUBS 0.016112f
C1513 VTAIL.n311 VSUBS 0.028317f
C1514 VTAIL.n312 VSUBS 0.015217f
C1515 VTAIL.n313 VSUBS 0.035966f
C1516 VTAIL.n314 VSUBS 0.016112f
C1517 VTAIL.n315 VSUBS 0.028317f
C1518 VTAIL.n316 VSUBS 0.015664f
C1519 VTAIL.n317 VSUBS 0.035966f
C1520 VTAIL.n318 VSUBS 0.016112f
C1521 VTAIL.n319 VSUBS 0.028317f
C1522 VTAIL.n320 VSUBS 0.015217f
C1523 VTAIL.n321 VSUBS 0.035966f
C1524 VTAIL.n322 VSUBS 0.016112f
C1525 VTAIL.n323 VSUBS 0.028317f
C1526 VTAIL.n324 VSUBS 0.015217f
C1527 VTAIL.n325 VSUBS 0.035966f
C1528 VTAIL.n326 VSUBS 0.016112f
C1529 VTAIL.n327 VSUBS 0.028317f
C1530 VTAIL.n328 VSUBS 0.015217f
C1531 VTAIL.n329 VSUBS 0.035966f
C1532 VTAIL.n330 VSUBS 0.016112f
C1533 VTAIL.n331 VSUBS 0.028317f
C1534 VTAIL.n332 VSUBS 0.015217f
C1535 VTAIL.n333 VSUBS 0.035966f
C1536 VTAIL.n334 VSUBS 0.016112f
C1537 VTAIL.n335 VSUBS 0.028317f
C1538 VTAIL.n336 VSUBS 0.015217f
C1539 VTAIL.n337 VSUBS 0.026975f
C1540 VTAIL.n338 VSUBS 0.02288f
C1541 VTAIL.t0 VSUBS 0.077221f
C1542 VTAIL.n339 VSUBS 0.226174f
C1543 VTAIL.n340 VSUBS 2.21693f
C1544 VTAIL.n341 VSUBS 0.015217f
C1545 VTAIL.n342 VSUBS 0.016112f
C1546 VTAIL.n343 VSUBS 0.035966f
C1547 VTAIL.n344 VSUBS 0.035966f
C1548 VTAIL.n345 VSUBS 0.016112f
C1549 VTAIL.n346 VSUBS 0.015217f
C1550 VTAIL.n347 VSUBS 0.028317f
C1551 VTAIL.n348 VSUBS 0.028317f
C1552 VTAIL.n349 VSUBS 0.015217f
C1553 VTAIL.n350 VSUBS 0.016112f
C1554 VTAIL.n351 VSUBS 0.035966f
C1555 VTAIL.n352 VSUBS 0.035966f
C1556 VTAIL.n353 VSUBS 0.016112f
C1557 VTAIL.n354 VSUBS 0.015217f
C1558 VTAIL.n355 VSUBS 0.028317f
C1559 VTAIL.n356 VSUBS 0.028317f
C1560 VTAIL.n357 VSUBS 0.015217f
C1561 VTAIL.n358 VSUBS 0.016112f
C1562 VTAIL.n359 VSUBS 0.035966f
C1563 VTAIL.n360 VSUBS 0.035966f
C1564 VTAIL.n361 VSUBS 0.016112f
C1565 VTAIL.n362 VSUBS 0.015217f
C1566 VTAIL.n363 VSUBS 0.028317f
C1567 VTAIL.n364 VSUBS 0.028317f
C1568 VTAIL.n365 VSUBS 0.015217f
C1569 VTAIL.n366 VSUBS 0.016112f
C1570 VTAIL.n367 VSUBS 0.035966f
C1571 VTAIL.n368 VSUBS 0.035966f
C1572 VTAIL.n369 VSUBS 0.016112f
C1573 VTAIL.n370 VSUBS 0.015217f
C1574 VTAIL.n371 VSUBS 0.028317f
C1575 VTAIL.n372 VSUBS 0.028317f
C1576 VTAIL.n373 VSUBS 0.015217f
C1577 VTAIL.n374 VSUBS 0.016112f
C1578 VTAIL.n375 VSUBS 0.035966f
C1579 VTAIL.n376 VSUBS 0.035966f
C1580 VTAIL.n377 VSUBS 0.016112f
C1581 VTAIL.n378 VSUBS 0.015217f
C1582 VTAIL.n379 VSUBS 0.028317f
C1583 VTAIL.n380 VSUBS 0.028317f
C1584 VTAIL.n381 VSUBS 0.015217f
C1585 VTAIL.n382 VSUBS 0.015217f
C1586 VTAIL.n383 VSUBS 0.016112f
C1587 VTAIL.n384 VSUBS 0.035966f
C1588 VTAIL.n385 VSUBS 0.035966f
C1589 VTAIL.n386 VSUBS 0.035966f
C1590 VTAIL.n387 VSUBS 0.015664f
C1591 VTAIL.n388 VSUBS 0.015217f
C1592 VTAIL.n389 VSUBS 0.028317f
C1593 VTAIL.n390 VSUBS 0.028317f
C1594 VTAIL.n391 VSUBS 0.015217f
C1595 VTAIL.n392 VSUBS 0.016112f
C1596 VTAIL.n393 VSUBS 0.035966f
C1597 VTAIL.n394 VSUBS 0.035966f
C1598 VTAIL.n395 VSUBS 0.016112f
C1599 VTAIL.n396 VSUBS 0.015217f
C1600 VTAIL.n397 VSUBS 0.028317f
C1601 VTAIL.n398 VSUBS 0.028317f
C1602 VTAIL.n399 VSUBS 0.015217f
C1603 VTAIL.n400 VSUBS 0.016112f
C1604 VTAIL.n401 VSUBS 0.035966f
C1605 VTAIL.n402 VSUBS 0.084214f
C1606 VTAIL.n403 VSUBS 0.016112f
C1607 VTAIL.n404 VSUBS 0.015217f
C1608 VTAIL.n405 VSUBS 0.063133f
C1609 VTAIL.n406 VSUBS 0.042151f
C1610 VTAIL.n407 VSUBS 2.1469f
C1611 VP.t1 VSUBS 5.40187f
C1612 VP.t0 VSUBS 6.14814f
C1613 VP.n0 VSUBS 6.4513f
.ends

