* NGSPICE file created from diff_pair_sample_0001.ext - technology: sky130A

.subckt diff_pair_sample_0001 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n2194_n3464# sky130_fd_pr__pfet_01v8 ad=4.8672 pd=25.74 as=4.8672 ps=25.74 w=12.48 l=2.73
X1 VDD2.t1 VN.t0 VTAIL.t0 w_n2194_n3464# sky130_fd_pr__pfet_01v8 ad=4.8672 pd=25.74 as=4.8672 ps=25.74 w=12.48 l=2.73
X2 B.t11 B.t9 B.t10 w_n2194_n3464# sky130_fd_pr__pfet_01v8 ad=4.8672 pd=25.74 as=0 ps=0 w=12.48 l=2.73
X3 VDD2.t0 VN.t1 VTAIL.t1 w_n2194_n3464# sky130_fd_pr__pfet_01v8 ad=4.8672 pd=25.74 as=4.8672 ps=25.74 w=12.48 l=2.73
X4 B.t8 B.t6 B.t7 w_n2194_n3464# sky130_fd_pr__pfet_01v8 ad=4.8672 pd=25.74 as=0 ps=0 w=12.48 l=2.73
X5 VDD1.t0 VP.t1 VTAIL.t3 w_n2194_n3464# sky130_fd_pr__pfet_01v8 ad=4.8672 pd=25.74 as=4.8672 ps=25.74 w=12.48 l=2.73
X6 B.t5 B.t3 B.t4 w_n2194_n3464# sky130_fd_pr__pfet_01v8 ad=4.8672 pd=25.74 as=0 ps=0 w=12.48 l=2.73
X7 B.t2 B.t0 B.t1 w_n2194_n3464# sky130_fd_pr__pfet_01v8 ad=4.8672 pd=25.74 as=0 ps=0 w=12.48 l=2.73
R0 VP.n0 VP.t1 196.591
R1 VP.n0 VP.t0 151.226
R2 VP VP.n0 0.43181
R3 VTAIL.n1 VTAIL.t1 59.3375
R4 VTAIL.n3 VTAIL.t0 59.3373
R5 VTAIL.n0 VTAIL.t2 59.3373
R6 VTAIL.n2 VTAIL.t3 59.3373
R7 VTAIL.n1 VTAIL.n0 28.4014
R8 VTAIL.n3 VTAIL.n2 25.7634
R9 VTAIL.n2 VTAIL.n1 1.78929
R10 VTAIL VTAIL.n0 1.188
R11 VTAIL VTAIL.n3 0.601793
R12 VDD1 VDD1.t1 116.894
R13 VDD1 VDD1.t0 76.7338
R14 VN VN.t1 196.593
R15 VN VN.t0 151.657
R16 VDD2.n0 VDD2.t1 115.71
R17 VDD2.n0 VDD2.t0 76.0161
R18 VDD2 VDD2.n0 0.718172
R19 B.n423 B.n422 585
R20 B.n424 B.n67 585
R21 B.n426 B.n425 585
R22 B.n427 B.n66 585
R23 B.n429 B.n428 585
R24 B.n430 B.n65 585
R25 B.n432 B.n431 585
R26 B.n433 B.n64 585
R27 B.n435 B.n434 585
R28 B.n436 B.n63 585
R29 B.n438 B.n437 585
R30 B.n439 B.n62 585
R31 B.n441 B.n440 585
R32 B.n442 B.n61 585
R33 B.n444 B.n443 585
R34 B.n445 B.n60 585
R35 B.n447 B.n446 585
R36 B.n448 B.n59 585
R37 B.n450 B.n449 585
R38 B.n451 B.n58 585
R39 B.n453 B.n452 585
R40 B.n454 B.n57 585
R41 B.n456 B.n455 585
R42 B.n457 B.n56 585
R43 B.n459 B.n458 585
R44 B.n460 B.n55 585
R45 B.n462 B.n461 585
R46 B.n463 B.n54 585
R47 B.n465 B.n464 585
R48 B.n466 B.n53 585
R49 B.n468 B.n467 585
R50 B.n469 B.n52 585
R51 B.n471 B.n470 585
R52 B.n472 B.n51 585
R53 B.n474 B.n473 585
R54 B.n475 B.n50 585
R55 B.n477 B.n476 585
R56 B.n478 B.n49 585
R57 B.n480 B.n479 585
R58 B.n481 B.n48 585
R59 B.n483 B.n482 585
R60 B.n484 B.n47 585
R61 B.n486 B.n485 585
R62 B.n488 B.n44 585
R63 B.n490 B.n489 585
R64 B.n491 B.n43 585
R65 B.n493 B.n492 585
R66 B.n494 B.n42 585
R67 B.n496 B.n495 585
R68 B.n497 B.n41 585
R69 B.n499 B.n498 585
R70 B.n500 B.n37 585
R71 B.n502 B.n501 585
R72 B.n503 B.n36 585
R73 B.n505 B.n504 585
R74 B.n506 B.n35 585
R75 B.n508 B.n507 585
R76 B.n509 B.n34 585
R77 B.n511 B.n510 585
R78 B.n512 B.n33 585
R79 B.n514 B.n513 585
R80 B.n515 B.n32 585
R81 B.n517 B.n516 585
R82 B.n518 B.n31 585
R83 B.n520 B.n519 585
R84 B.n521 B.n30 585
R85 B.n523 B.n522 585
R86 B.n524 B.n29 585
R87 B.n526 B.n525 585
R88 B.n527 B.n28 585
R89 B.n529 B.n528 585
R90 B.n530 B.n27 585
R91 B.n532 B.n531 585
R92 B.n533 B.n26 585
R93 B.n535 B.n534 585
R94 B.n536 B.n25 585
R95 B.n538 B.n537 585
R96 B.n539 B.n24 585
R97 B.n541 B.n540 585
R98 B.n542 B.n23 585
R99 B.n544 B.n543 585
R100 B.n545 B.n22 585
R101 B.n547 B.n546 585
R102 B.n548 B.n21 585
R103 B.n550 B.n549 585
R104 B.n551 B.n20 585
R105 B.n553 B.n552 585
R106 B.n554 B.n19 585
R107 B.n556 B.n555 585
R108 B.n557 B.n18 585
R109 B.n559 B.n558 585
R110 B.n560 B.n17 585
R111 B.n562 B.n561 585
R112 B.n563 B.n16 585
R113 B.n565 B.n564 585
R114 B.n566 B.n15 585
R115 B.n421 B.n68 585
R116 B.n420 B.n419 585
R117 B.n418 B.n69 585
R118 B.n417 B.n416 585
R119 B.n415 B.n70 585
R120 B.n414 B.n413 585
R121 B.n412 B.n71 585
R122 B.n411 B.n410 585
R123 B.n409 B.n72 585
R124 B.n408 B.n407 585
R125 B.n406 B.n73 585
R126 B.n405 B.n404 585
R127 B.n403 B.n74 585
R128 B.n402 B.n401 585
R129 B.n400 B.n75 585
R130 B.n399 B.n398 585
R131 B.n397 B.n76 585
R132 B.n396 B.n395 585
R133 B.n394 B.n77 585
R134 B.n393 B.n392 585
R135 B.n391 B.n78 585
R136 B.n390 B.n389 585
R137 B.n388 B.n79 585
R138 B.n387 B.n386 585
R139 B.n385 B.n80 585
R140 B.n384 B.n383 585
R141 B.n382 B.n81 585
R142 B.n381 B.n380 585
R143 B.n379 B.n82 585
R144 B.n378 B.n377 585
R145 B.n376 B.n83 585
R146 B.n375 B.n374 585
R147 B.n373 B.n84 585
R148 B.n372 B.n371 585
R149 B.n370 B.n85 585
R150 B.n369 B.n368 585
R151 B.n367 B.n86 585
R152 B.n366 B.n365 585
R153 B.n364 B.n87 585
R154 B.n363 B.n362 585
R155 B.n361 B.n88 585
R156 B.n360 B.n359 585
R157 B.n358 B.n89 585
R158 B.n357 B.n356 585
R159 B.n355 B.n90 585
R160 B.n354 B.n353 585
R161 B.n352 B.n91 585
R162 B.n351 B.n350 585
R163 B.n349 B.n92 585
R164 B.n348 B.n347 585
R165 B.n346 B.n93 585
R166 B.n345 B.n344 585
R167 B.n343 B.n94 585
R168 B.n198 B.n197 585
R169 B.n199 B.n146 585
R170 B.n201 B.n200 585
R171 B.n202 B.n145 585
R172 B.n204 B.n203 585
R173 B.n205 B.n144 585
R174 B.n207 B.n206 585
R175 B.n208 B.n143 585
R176 B.n210 B.n209 585
R177 B.n211 B.n142 585
R178 B.n213 B.n212 585
R179 B.n214 B.n141 585
R180 B.n216 B.n215 585
R181 B.n217 B.n140 585
R182 B.n219 B.n218 585
R183 B.n220 B.n139 585
R184 B.n222 B.n221 585
R185 B.n223 B.n138 585
R186 B.n225 B.n224 585
R187 B.n226 B.n137 585
R188 B.n228 B.n227 585
R189 B.n229 B.n136 585
R190 B.n231 B.n230 585
R191 B.n232 B.n135 585
R192 B.n234 B.n233 585
R193 B.n235 B.n134 585
R194 B.n237 B.n236 585
R195 B.n238 B.n133 585
R196 B.n240 B.n239 585
R197 B.n241 B.n132 585
R198 B.n243 B.n242 585
R199 B.n244 B.n131 585
R200 B.n246 B.n245 585
R201 B.n247 B.n130 585
R202 B.n249 B.n248 585
R203 B.n250 B.n129 585
R204 B.n252 B.n251 585
R205 B.n253 B.n128 585
R206 B.n255 B.n254 585
R207 B.n256 B.n127 585
R208 B.n258 B.n257 585
R209 B.n259 B.n126 585
R210 B.n261 B.n260 585
R211 B.n263 B.n262 585
R212 B.n264 B.n122 585
R213 B.n266 B.n265 585
R214 B.n267 B.n121 585
R215 B.n269 B.n268 585
R216 B.n270 B.n120 585
R217 B.n272 B.n271 585
R218 B.n273 B.n119 585
R219 B.n275 B.n274 585
R220 B.n276 B.n116 585
R221 B.n279 B.n278 585
R222 B.n280 B.n115 585
R223 B.n282 B.n281 585
R224 B.n283 B.n114 585
R225 B.n285 B.n284 585
R226 B.n286 B.n113 585
R227 B.n288 B.n287 585
R228 B.n289 B.n112 585
R229 B.n291 B.n290 585
R230 B.n292 B.n111 585
R231 B.n294 B.n293 585
R232 B.n295 B.n110 585
R233 B.n297 B.n296 585
R234 B.n298 B.n109 585
R235 B.n300 B.n299 585
R236 B.n301 B.n108 585
R237 B.n303 B.n302 585
R238 B.n304 B.n107 585
R239 B.n306 B.n305 585
R240 B.n307 B.n106 585
R241 B.n309 B.n308 585
R242 B.n310 B.n105 585
R243 B.n312 B.n311 585
R244 B.n313 B.n104 585
R245 B.n315 B.n314 585
R246 B.n316 B.n103 585
R247 B.n318 B.n317 585
R248 B.n319 B.n102 585
R249 B.n321 B.n320 585
R250 B.n322 B.n101 585
R251 B.n324 B.n323 585
R252 B.n325 B.n100 585
R253 B.n327 B.n326 585
R254 B.n328 B.n99 585
R255 B.n330 B.n329 585
R256 B.n331 B.n98 585
R257 B.n333 B.n332 585
R258 B.n334 B.n97 585
R259 B.n336 B.n335 585
R260 B.n337 B.n96 585
R261 B.n339 B.n338 585
R262 B.n340 B.n95 585
R263 B.n342 B.n341 585
R264 B.n196 B.n147 585
R265 B.n195 B.n194 585
R266 B.n193 B.n148 585
R267 B.n192 B.n191 585
R268 B.n190 B.n149 585
R269 B.n189 B.n188 585
R270 B.n187 B.n150 585
R271 B.n186 B.n185 585
R272 B.n184 B.n151 585
R273 B.n183 B.n182 585
R274 B.n181 B.n152 585
R275 B.n180 B.n179 585
R276 B.n178 B.n153 585
R277 B.n177 B.n176 585
R278 B.n175 B.n154 585
R279 B.n174 B.n173 585
R280 B.n172 B.n155 585
R281 B.n171 B.n170 585
R282 B.n169 B.n156 585
R283 B.n168 B.n167 585
R284 B.n166 B.n157 585
R285 B.n165 B.n164 585
R286 B.n163 B.n158 585
R287 B.n162 B.n161 585
R288 B.n160 B.n159 585
R289 B.n2 B.n0 585
R290 B.n605 B.n1 585
R291 B.n604 B.n603 585
R292 B.n602 B.n3 585
R293 B.n601 B.n600 585
R294 B.n599 B.n4 585
R295 B.n598 B.n597 585
R296 B.n596 B.n5 585
R297 B.n595 B.n594 585
R298 B.n593 B.n6 585
R299 B.n592 B.n591 585
R300 B.n590 B.n7 585
R301 B.n589 B.n588 585
R302 B.n587 B.n8 585
R303 B.n586 B.n585 585
R304 B.n584 B.n9 585
R305 B.n583 B.n582 585
R306 B.n581 B.n10 585
R307 B.n580 B.n579 585
R308 B.n578 B.n11 585
R309 B.n577 B.n576 585
R310 B.n575 B.n12 585
R311 B.n574 B.n573 585
R312 B.n572 B.n13 585
R313 B.n571 B.n570 585
R314 B.n569 B.n14 585
R315 B.n568 B.n567 585
R316 B.n607 B.n606 585
R317 B.n197 B.n196 487.695
R318 B.n568 B.n15 487.695
R319 B.n341 B.n94 487.695
R320 B.n423 B.n68 487.695
R321 B.n117 B.t6 318.406
R322 B.n123 B.t9 318.406
R323 B.n38 B.t3 318.406
R324 B.n45 B.t0 318.406
R325 B.n117 B.t8 171
R326 B.n45 B.t1 171
R327 B.n123 B.t11 170.984
R328 B.n38 B.t4 170.984
R329 B.n196 B.n195 163.367
R330 B.n195 B.n148 163.367
R331 B.n191 B.n148 163.367
R332 B.n191 B.n190 163.367
R333 B.n190 B.n189 163.367
R334 B.n189 B.n150 163.367
R335 B.n185 B.n150 163.367
R336 B.n185 B.n184 163.367
R337 B.n184 B.n183 163.367
R338 B.n183 B.n152 163.367
R339 B.n179 B.n152 163.367
R340 B.n179 B.n178 163.367
R341 B.n178 B.n177 163.367
R342 B.n177 B.n154 163.367
R343 B.n173 B.n154 163.367
R344 B.n173 B.n172 163.367
R345 B.n172 B.n171 163.367
R346 B.n171 B.n156 163.367
R347 B.n167 B.n156 163.367
R348 B.n167 B.n166 163.367
R349 B.n166 B.n165 163.367
R350 B.n165 B.n158 163.367
R351 B.n161 B.n158 163.367
R352 B.n161 B.n160 163.367
R353 B.n160 B.n2 163.367
R354 B.n606 B.n2 163.367
R355 B.n606 B.n605 163.367
R356 B.n605 B.n604 163.367
R357 B.n604 B.n3 163.367
R358 B.n600 B.n3 163.367
R359 B.n600 B.n599 163.367
R360 B.n599 B.n598 163.367
R361 B.n598 B.n5 163.367
R362 B.n594 B.n5 163.367
R363 B.n594 B.n593 163.367
R364 B.n593 B.n592 163.367
R365 B.n592 B.n7 163.367
R366 B.n588 B.n7 163.367
R367 B.n588 B.n587 163.367
R368 B.n587 B.n586 163.367
R369 B.n586 B.n9 163.367
R370 B.n582 B.n9 163.367
R371 B.n582 B.n581 163.367
R372 B.n581 B.n580 163.367
R373 B.n580 B.n11 163.367
R374 B.n576 B.n11 163.367
R375 B.n576 B.n575 163.367
R376 B.n575 B.n574 163.367
R377 B.n574 B.n13 163.367
R378 B.n570 B.n13 163.367
R379 B.n570 B.n569 163.367
R380 B.n569 B.n568 163.367
R381 B.n197 B.n146 163.367
R382 B.n201 B.n146 163.367
R383 B.n202 B.n201 163.367
R384 B.n203 B.n202 163.367
R385 B.n203 B.n144 163.367
R386 B.n207 B.n144 163.367
R387 B.n208 B.n207 163.367
R388 B.n209 B.n208 163.367
R389 B.n209 B.n142 163.367
R390 B.n213 B.n142 163.367
R391 B.n214 B.n213 163.367
R392 B.n215 B.n214 163.367
R393 B.n215 B.n140 163.367
R394 B.n219 B.n140 163.367
R395 B.n220 B.n219 163.367
R396 B.n221 B.n220 163.367
R397 B.n221 B.n138 163.367
R398 B.n225 B.n138 163.367
R399 B.n226 B.n225 163.367
R400 B.n227 B.n226 163.367
R401 B.n227 B.n136 163.367
R402 B.n231 B.n136 163.367
R403 B.n232 B.n231 163.367
R404 B.n233 B.n232 163.367
R405 B.n233 B.n134 163.367
R406 B.n237 B.n134 163.367
R407 B.n238 B.n237 163.367
R408 B.n239 B.n238 163.367
R409 B.n239 B.n132 163.367
R410 B.n243 B.n132 163.367
R411 B.n244 B.n243 163.367
R412 B.n245 B.n244 163.367
R413 B.n245 B.n130 163.367
R414 B.n249 B.n130 163.367
R415 B.n250 B.n249 163.367
R416 B.n251 B.n250 163.367
R417 B.n251 B.n128 163.367
R418 B.n255 B.n128 163.367
R419 B.n256 B.n255 163.367
R420 B.n257 B.n256 163.367
R421 B.n257 B.n126 163.367
R422 B.n261 B.n126 163.367
R423 B.n262 B.n261 163.367
R424 B.n262 B.n122 163.367
R425 B.n266 B.n122 163.367
R426 B.n267 B.n266 163.367
R427 B.n268 B.n267 163.367
R428 B.n268 B.n120 163.367
R429 B.n272 B.n120 163.367
R430 B.n273 B.n272 163.367
R431 B.n274 B.n273 163.367
R432 B.n274 B.n116 163.367
R433 B.n279 B.n116 163.367
R434 B.n280 B.n279 163.367
R435 B.n281 B.n280 163.367
R436 B.n281 B.n114 163.367
R437 B.n285 B.n114 163.367
R438 B.n286 B.n285 163.367
R439 B.n287 B.n286 163.367
R440 B.n287 B.n112 163.367
R441 B.n291 B.n112 163.367
R442 B.n292 B.n291 163.367
R443 B.n293 B.n292 163.367
R444 B.n293 B.n110 163.367
R445 B.n297 B.n110 163.367
R446 B.n298 B.n297 163.367
R447 B.n299 B.n298 163.367
R448 B.n299 B.n108 163.367
R449 B.n303 B.n108 163.367
R450 B.n304 B.n303 163.367
R451 B.n305 B.n304 163.367
R452 B.n305 B.n106 163.367
R453 B.n309 B.n106 163.367
R454 B.n310 B.n309 163.367
R455 B.n311 B.n310 163.367
R456 B.n311 B.n104 163.367
R457 B.n315 B.n104 163.367
R458 B.n316 B.n315 163.367
R459 B.n317 B.n316 163.367
R460 B.n317 B.n102 163.367
R461 B.n321 B.n102 163.367
R462 B.n322 B.n321 163.367
R463 B.n323 B.n322 163.367
R464 B.n323 B.n100 163.367
R465 B.n327 B.n100 163.367
R466 B.n328 B.n327 163.367
R467 B.n329 B.n328 163.367
R468 B.n329 B.n98 163.367
R469 B.n333 B.n98 163.367
R470 B.n334 B.n333 163.367
R471 B.n335 B.n334 163.367
R472 B.n335 B.n96 163.367
R473 B.n339 B.n96 163.367
R474 B.n340 B.n339 163.367
R475 B.n341 B.n340 163.367
R476 B.n345 B.n94 163.367
R477 B.n346 B.n345 163.367
R478 B.n347 B.n346 163.367
R479 B.n347 B.n92 163.367
R480 B.n351 B.n92 163.367
R481 B.n352 B.n351 163.367
R482 B.n353 B.n352 163.367
R483 B.n353 B.n90 163.367
R484 B.n357 B.n90 163.367
R485 B.n358 B.n357 163.367
R486 B.n359 B.n358 163.367
R487 B.n359 B.n88 163.367
R488 B.n363 B.n88 163.367
R489 B.n364 B.n363 163.367
R490 B.n365 B.n364 163.367
R491 B.n365 B.n86 163.367
R492 B.n369 B.n86 163.367
R493 B.n370 B.n369 163.367
R494 B.n371 B.n370 163.367
R495 B.n371 B.n84 163.367
R496 B.n375 B.n84 163.367
R497 B.n376 B.n375 163.367
R498 B.n377 B.n376 163.367
R499 B.n377 B.n82 163.367
R500 B.n381 B.n82 163.367
R501 B.n382 B.n381 163.367
R502 B.n383 B.n382 163.367
R503 B.n383 B.n80 163.367
R504 B.n387 B.n80 163.367
R505 B.n388 B.n387 163.367
R506 B.n389 B.n388 163.367
R507 B.n389 B.n78 163.367
R508 B.n393 B.n78 163.367
R509 B.n394 B.n393 163.367
R510 B.n395 B.n394 163.367
R511 B.n395 B.n76 163.367
R512 B.n399 B.n76 163.367
R513 B.n400 B.n399 163.367
R514 B.n401 B.n400 163.367
R515 B.n401 B.n74 163.367
R516 B.n405 B.n74 163.367
R517 B.n406 B.n405 163.367
R518 B.n407 B.n406 163.367
R519 B.n407 B.n72 163.367
R520 B.n411 B.n72 163.367
R521 B.n412 B.n411 163.367
R522 B.n413 B.n412 163.367
R523 B.n413 B.n70 163.367
R524 B.n417 B.n70 163.367
R525 B.n418 B.n417 163.367
R526 B.n419 B.n418 163.367
R527 B.n419 B.n68 163.367
R528 B.n564 B.n15 163.367
R529 B.n564 B.n563 163.367
R530 B.n563 B.n562 163.367
R531 B.n562 B.n17 163.367
R532 B.n558 B.n17 163.367
R533 B.n558 B.n557 163.367
R534 B.n557 B.n556 163.367
R535 B.n556 B.n19 163.367
R536 B.n552 B.n19 163.367
R537 B.n552 B.n551 163.367
R538 B.n551 B.n550 163.367
R539 B.n550 B.n21 163.367
R540 B.n546 B.n21 163.367
R541 B.n546 B.n545 163.367
R542 B.n545 B.n544 163.367
R543 B.n544 B.n23 163.367
R544 B.n540 B.n23 163.367
R545 B.n540 B.n539 163.367
R546 B.n539 B.n538 163.367
R547 B.n538 B.n25 163.367
R548 B.n534 B.n25 163.367
R549 B.n534 B.n533 163.367
R550 B.n533 B.n532 163.367
R551 B.n532 B.n27 163.367
R552 B.n528 B.n27 163.367
R553 B.n528 B.n527 163.367
R554 B.n527 B.n526 163.367
R555 B.n526 B.n29 163.367
R556 B.n522 B.n29 163.367
R557 B.n522 B.n521 163.367
R558 B.n521 B.n520 163.367
R559 B.n520 B.n31 163.367
R560 B.n516 B.n31 163.367
R561 B.n516 B.n515 163.367
R562 B.n515 B.n514 163.367
R563 B.n514 B.n33 163.367
R564 B.n510 B.n33 163.367
R565 B.n510 B.n509 163.367
R566 B.n509 B.n508 163.367
R567 B.n508 B.n35 163.367
R568 B.n504 B.n35 163.367
R569 B.n504 B.n503 163.367
R570 B.n503 B.n502 163.367
R571 B.n502 B.n37 163.367
R572 B.n498 B.n37 163.367
R573 B.n498 B.n497 163.367
R574 B.n497 B.n496 163.367
R575 B.n496 B.n42 163.367
R576 B.n492 B.n42 163.367
R577 B.n492 B.n491 163.367
R578 B.n491 B.n490 163.367
R579 B.n490 B.n44 163.367
R580 B.n485 B.n44 163.367
R581 B.n485 B.n484 163.367
R582 B.n484 B.n483 163.367
R583 B.n483 B.n48 163.367
R584 B.n479 B.n48 163.367
R585 B.n479 B.n478 163.367
R586 B.n478 B.n477 163.367
R587 B.n477 B.n50 163.367
R588 B.n473 B.n50 163.367
R589 B.n473 B.n472 163.367
R590 B.n472 B.n471 163.367
R591 B.n471 B.n52 163.367
R592 B.n467 B.n52 163.367
R593 B.n467 B.n466 163.367
R594 B.n466 B.n465 163.367
R595 B.n465 B.n54 163.367
R596 B.n461 B.n54 163.367
R597 B.n461 B.n460 163.367
R598 B.n460 B.n459 163.367
R599 B.n459 B.n56 163.367
R600 B.n455 B.n56 163.367
R601 B.n455 B.n454 163.367
R602 B.n454 B.n453 163.367
R603 B.n453 B.n58 163.367
R604 B.n449 B.n58 163.367
R605 B.n449 B.n448 163.367
R606 B.n448 B.n447 163.367
R607 B.n447 B.n60 163.367
R608 B.n443 B.n60 163.367
R609 B.n443 B.n442 163.367
R610 B.n442 B.n441 163.367
R611 B.n441 B.n62 163.367
R612 B.n437 B.n62 163.367
R613 B.n437 B.n436 163.367
R614 B.n436 B.n435 163.367
R615 B.n435 B.n64 163.367
R616 B.n431 B.n64 163.367
R617 B.n431 B.n430 163.367
R618 B.n430 B.n429 163.367
R619 B.n429 B.n66 163.367
R620 B.n425 B.n66 163.367
R621 B.n425 B.n424 163.367
R622 B.n424 B.n423 163.367
R623 B.n118 B.t7 111.653
R624 B.n46 B.t2 111.653
R625 B.n124 B.t10 111.638
R626 B.n39 B.t5 111.638
R627 B.n277 B.n118 59.5399
R628 B.n125 B.n124 59.5399
R629 B.n40 B.n39 59.5399
R630 B.n487 B.n46 59.5399
R631 B.n118 B.n117 59.346
R632 B.n124 B.n123 59.346
R633 B.n39 B.n38 59.346
R634 B.n46 B.n45 59.346
R635 B.n567 B.n566 31.6883
R636 B.n422 B.n421 31.6883
R637 B.n343 B.n342 31.6883
R638 B.n198 B.n147 31.6883
R639 B B.n607 18.0485
R640 B.n566 B.n565 10.6151
R641 B.n565 B.n16 10.6151
R642 B.n561 B.n16 10.6151
R643 B.n561 B.n560 10.6151
R644 B.n560 B.n559 10.6151
R645 B.n559 B.n18 10.6151
R646 B.n555 B.n18 10.6151
R647 B.n555 B.n554 10.6151
R648 B.n554 B.n553 10.6151
R649 B.n553 B.n20 10.6151
R650 B.n549 B.n20 10.6151
R651 B.n549 B.n548 10.6151
R652 B.n548 B.n547 10.6151
R653 B.n547 B.n22 10.6151
R654 B.n543 B.n22 10.6151
R655 B.n543 B.n542 10.6151
R656 B.n542 B.n541 10.6151
R657 B.n541 B.n24 10.6151
R658 B.n537 B.n24 10.6151
R659 B.n537 B.n536 10.6151
R660 B.n536 B.n535 10.6151
R661 B.n535 B.n26 10.6151
R662 B.n531 B.n26 10.6151
R663 B.n531 B.n530 10.6151
R664 B.n530 B.n529 10.6151
R665 B.n529 B.n28 10.6151
R666 B.n525 B.n28 10.6151
R667 B.n525 B.n524 10.6151
R668 B.n524 B.n523 10.6151
R669 B.n523 B.n30 10.6151
R670 B.n519 B.n30 10.6151
R671 B.n519 B.n518 10.6151
R672 B.n518 B.n517 10.6151
R673 B.n517 B.n32 10.6151
R674 B.n513 B.n32 10.6151
R675 B.n513 B.n512 10.6151
R676 B.n512 B.n511 10.6151
R677 B.n511 B.n34 10.6151
R678 B.n507 B.n34 10.6151
R679 B.n507 B.n506 10.6151
R680 B.n506 B.n505 10.6151
R681 B.n505 B.n36 10.6151
R682 B.n501 B.n500 10.6151
R683 B.n500 B.n499 10.6151
R684 B.n499 B.n41 10.6151
R685 B.n495 B.n41 10.6151
R686 B.n495 B.n494 10.6151
R687 B.n494 B.n493 10.6151
R688 B.n493 B.n43 10.6151
R689 B.n489 B.n43 10.6151
R690 B.n489 B.n488 10.6151
R691 B.n486 B.n47 10.6151
R692 B.n482 B.n47 10.6151
R693 B.n482 B.n481 10.6151
R694 B.n481 B.n480 10.6151
R695 B.n480 B.n49 10.6151
R696 B.n476 B.n49 10.6151
R697 B.n476 B.n475 10.6151
R698 B.n475 B.n474 10.6151
R699 B.n474 B.n51 10.6151
R700 B.n470 B.n51 10.6151
R701 B.n470 B.n469 10.6151
R702 B.n469 B.n468 10.6151
R703 B.n468 B.n53 10.6151
R704 B.n464 B.n53 10.6151
R705 B.n464 B.n463 10.6151
R706 B.n463 B.n462 10.6151
R707 B.n462 B.n55 10.6151
R708 B.n458 B.n55 10.6151
R709 B.n458 B.n457 10.6151
R710 B.n457 B.n456 10.6151
R711 B.n456 B.n57 10.6151
R712 B.n452 B.n57 10.6151
R713 B.n452 B.n451 10.6151
R714 B.n451 B.n450 10.6151
R715 B.n450 B.n59 10.6151
R716 B.n446 B.n59 10.6151
R717 B.n446 B.n445 10.6151
R718 B.n445 B.n444 10.6151
R719 B.n444 B.n61 10.6151
R720 B.n440 B.n61 10.6151
R721 B.n440 B.n439 10.6151
R722 B.n439 B.n438 10.6151
R723 B.n438 B.n63 10.6151
R724 B.n434 B.n63 10.6151
R725 B.n434 B.n433 10.6151
R726 B.n433 B.n432 10.6151
R727 B.n432 B.n65 10.6151
R728 B.n428 B.n65 10.6151
R729 B.n428 B.n427 10.6151
R730 B.n427 B.n426 10.6151
R731 B.n426 B.n67 10.6151
R732 B.n422 B.n67 10.6151
R733 B.n344 B.n343 10.6151
R734 B.n344 B.n93 10.6151
R735 B.n348 B.n93 10.6151
R736 B.n349 B.n348 10.6151
R737 B.n350 B.n349 10.6151
R738 B.n350 B.n91 10.6151
R739 B.n354 B.n91 10.6151
R740 B.n355 B.n354 10.6151
R741 B.n356 B.n355 10.6151
R742 B.n356 B.n89 10.6151
R743 B.n360 B.n89 10.6151
R744 B.n361 B.n360 10.6151
R745 B.n362 B.n361 10.6151
R746 B.n362 B.n87 10.6151
R747 B.n366 B.n87 10.6151
R748 B.n367 B.n366 10.6151
R749 B.n368 B.n367 10.6151
R750 B.n368 B.n85 10.6151
R751 B.n372 B.n85 10.6151
R752 B.n373 B.n372 10.6151
R753 B.n374 B.n373 10.6151
R754 B.n374 B.n83 10.6151
R755 B.n378 B.n83 10.6151
R756 B.n379 B.n378 10.6151
R757 B.n380 B.n379 10.6151
R758 B.n380 B.n81 10.6151
R759 B.n384 B.n81 10.6151
R760 B.n385 B.n384 10.6151
R761 B.n386 B.n385 10.6151
R762 B.n386 B.n79 10.6151
R763 B.n390 B.n79 10.6151
R764 B.n391 B.n390 10.6151
R765 B.n392 B.n391 10.6151
R766 B.n392 B.n77 10.6151
R767 B.n396 B.n77 10.6151
R768 B.n397 B.n396 10.6151
R769 B.n398 B.n397 10.6151
R770 B.n398 B.n75 10.6151
R771 B.n402 B.n75 10.6151
R772 B.n403 B.n402 10.6151
R773 B.n404 B.n403 10.6151
R774 B.n404 B.n73 10.6151
R775 B.n408 B.n73 10.6151
R776 B.n409 B.n408 10.6151
R777 B.n410 B.n409 10.6151
R778 B.n410 B.n71 10.6151
R779 B.n414 B.n71 10.6151
R780 B.n415 B.n414 10.6151
R781 B.n416 B.n415 10.6151
R782 B.n416 B.n69 10.6151
R783 B.n420 B.n69 10.6151
R784 B.n421 B.n420 10.6151
R785 B.n199 B.n198 10.6151
R786 B.n200 B.n199 10.6151
R787 B.n200 B.n145 10.6151
R788 B.n204 B.n145 10.6151
R789 B.n205 B.n204 10.6151
R790 B.n206 B.n205 10.6151
R791 B.n206 B.n143 10.6151
R792 B.n210 B.n143 10.6151
R793 B.n211 B.n210 10.6151
R794 B.n212 B.n211 10.6151
R795 B.n212 B.n141 10.6151
R796 B.n216 B.n141 10.6151
R797 B.n217 B.n216 10.6151
R798 B.n218 B.n217 10.6151
R799 B.n218 B.n139 10.6151
R800 B.n222 B.n139 10.6151
R801 B.n223 B.n222 10.6151
R802 B.n224 B.n223 10.6151
R803 B.n224 B.n137 10.6151
R804 B.n228 B.n137 10.6151
R805 B.n229 B.n228 10.6151
R806 B.n230 B.n229 10.6151
R807 B.n230 B.n135 10.6151
R808 B.n234 B.n135 10.6151
R809 B.n235 B.n234 10.6151
R810 B.n236 B.n235 10.6151
R811 B.n236 B.n133 10.6151
R812 B.n240 B.n133 10.6151
R813 B.n241 B.n240 10.6151
R814 B.n242 B.n241 10.6151
R815 B.n242 B.n131 10.6151
R816 B.n246 B.n131 10.6151
R817 B.n247 B.n246 10.6151
R818 B.n248 B.n247 10.6151
R819 B.n248 B.n129 10.6151
R820 B.n252 B.n129 10.6151
R821 B.n253 B.n252 10.6151
R822 B.n254 B.n253 10.6151
R823 B.n254 B.n127 10.6151
R824 B.n258 B.n127 10.6151
R825 B.n259 B.n258 10.6151
R826 B.n260 B.n259 10.6151
R827 B.n264 B.n263 10.6151
R828 B.n265 B.n264 10.6151
R829 B.n265 B.n121 10.6151
R830 B.n269 B.n121 10.6151
R831 B.n270 B.n269 10.6151
R832 B.n271 B.n270 10.6151
R833 B.n271 B.n119 10.6151
R834 B.n275 B.n119 10.6151
R835 B.n276 B.n275 10.6151
R836 B.n278 B.n115 10.6151
R837 B.n282 B.n115 10.6151
R838 B.n283 B.n282 10.6151
R839 B.n284 B.n283 10.6151
R840 B.n284 B.n113 10.6151
R841 B.n288 B.n113 10.6151
R842 B.n289 B.n288 10.6151
R843 B.n290 B.n289 10.6151
R844 B.n290 B.n111 10.6151
R845 B.n294 B.n111 10.6151
R846 B.n295 B.n294 10.6151
R847 B.n296 B.n295 10.6151
R848 B.n296 B.n109 10.6151
R849 B.n300 B.n109 10.6151
R850 B.n301 B.n300 10.6151
R851 B.n302 B.n301 10.6151
R852 B.n302 B.n107 10.6151
R853 B.n306 B.n107 10.6151
R854 B.n307 B.n306 10.6151
R855 B.n308 B.n307 10.6151
R856 B.n308 B.n105 10.6151
R857 B.n312 B.n105 10.6151
R858 B.n313 B.n312 10.6151
R859 B.n314 B.n313 10.6151
R860 B.n314 B.n103 10.6151
R861 B.n318 B.n103 10.6151
R862 B.n319 B.n318 10.6151
R863 B.n320 B.n319 10.6151
R864 B.n320 B.n101 10.6151
R865 B.n324 B.n101 10.6151
R866 B.n325 B.n324 10.6151
R867 B.n326 B.n325 10.6151
R868 B.n326 B.n99 10.6151
R869 B.n330 B.n99 10.6151
R870 B.n331 B.n330 10.6151
R871 B.n332 B.n331 10.6151
R872 B.n332 B.n97 10.6151
R873 B.n336 B.n97 10.6151
R874 B.n337 B.n336 10.6151
R875 B.n338 B.n337 10.6151
R876 B.n338 B.n95 10.6151
R877 B.n342 B.n95 10.6151
R878 B.n194 B.n147 10.6151
R879 B.n194 B.n193 10.6151
R880 B.n193 B.n192 10.6151
R881 B.n192 B.n149 10.6151
R882 B.n188 B.n149 10.6151
R883 B.n188 B.n187 10.6151
R884 B.n187 B.n186 10.6151
R885 B.n186 B.n151 10.6151
R886 B.n182 B.n151 10.6151
R887 B.n182 B.n181 10.6151
R888 B.n181 B.n180 10.6151
R889 B.n180 B.n153 10.6151
R890 B.n176 B.n153 10.6151
R891 B.n176 B.n175 10.6151
R892 B.n175 B.n174 10.6151
R893 B.n174 B.n155 10.6151
R894 B.n170 B.n155 10.6151
R895 B.n170 B.n169 10.6151
R896 B.n169 B.n168 10.6151
R897 B.n168 B.n157 10.6151
R898 B.n164 B.n157 10.6151
R899 B.n164 B.n163 10.6151
R900 B.n163 B.n162 10.6151
R901 B.n162 B.n159 10.6151
R902 B.n159 B.n0 10.6151
R903 B.n603 B.n1 10.6151
R904 B.n603 B.n602 10.6151
R905 B.n602 B.n601 10.6151
R906 B.n601 B.n4 10.6151
R907 B.n597 B.n4 10.6151
R908 B.n597 B.n596 10.6151
R909 B.n596 B.n595 10.6151
R910 B.n595 B.n6 10.6151
R911 B.n591 B.n6 10.6151
R912 B.n591 B.n590 10.6151
R913 B.n590 B.n589 10.6151
R914 B.n589 B.n8 10.6151
R915 B.n585 B.n8 10.6151
R916 B.n585 B.n584 10.6151
R917 B.n584 B.n583 10.6151
R918 B.n583 B.n10 10.6151
R919 B.n579 B.n10 10.6151
R920 B.n579 B.n578 10.6151
R921 B.n578 B.n577 10.6151
R922 B.n577 B.n12 10.6151
R923 B.n573 B.n12 10.6151
R924 B.n573 B.n572 10.6151
R925 B.n572 B.n571 10.6151
R926 B.n571 B.n14 10.6151
R927 B.n567 B.n14 10.6151
R928 B.n40 B.n36 9.36635
R929 B.n487 B.n486 9.36635
R930 B.n260 B.n125 9.36635
R931 B.n278 B.n277 9.36635
R932 B.n607 B.n0 2.81026
R933 B.n607 B.n1 2.81026
R934 B.n501 B.n40 1.24928
R935 B.n488 B.n487 1.24928
R936 B.n263 B.n125 1.24928
R937 B.n277 B.n276 1.24928
C0 VN w_n2194_n3464# 3.06514f
C1 VP VTAIL 2.5723f
C2 VDD2 w_n2194_n3464# 1.85643f
C3 VN VDD2 2.90254f
C4 B w_n2194_n3464# 9.083691f
C5 VN B 1.07356f
C6 w_n2194_n3464# VDD1 1.82894f
C7 B VDD2 1.79244f
C8 VN VDD1 0.147848f
C9 VDD2 VDD1 0.690357f
C10 VP w_n2194_n3464# 3.34489f
C11 VN VP 5.61146f
C12 VP VDD2 0.338226f
C13 w_n2194_n3464# VTAIL 2.80905f
C14 VN VTAIL 2.55801f
C15 VDD2 VTAIL 5.26344f
C16 B VDD1 1.76121f
C17 VP B 1.53401f
C18 VP VDD1 3.09037f
C19 B VTAIL 3.8175f
C20 VDD1 VTAIL 5.21193f
C21 VDD2 VSUBS 0.914107f
C22 VDD1 VSUBS 4.59804f
C23 VTAIL VSUBS 1.033836f
C24 VN VSUBS 8.05488f
C25 VP VSUBS 1.746813f
C26 B VSUBS 4.044565f
C27 w_n2194_n3464# VSUBS 93.49071f
C28 B.n0 VSUBS 0.003768f
C29 B.n1 VSUBS 0.003768f
C30 B.n2 VSUBS 0.005959f
C31 B.n3 VSUBS 0.005959f
C32 B.n4 VSUBS 0.005959f
C33 B.n5 VSUBS 0.005959f
C34 B.n6 VSUBS 0.005959f
C35 B.n7 VSUBS 0.005959f
C36 B.n8 VSUBS 0.005959f
C37 B.n9 VSUBS 0.005959f
C38 B.n10 VSUBS 0.005959f
C39 B.n11 VSUBS 0.005959f
C40 B.n12 VSUBS 0.005959f
C41 B.n13 VSUBS 0.005959f
C42 B.n14 VSUBS 0.005959f
C43 B.n15 VSUBS 0.014193f
C44 B.n16 VSUBS 0.005959f
C45 B.n17 VSUBS 0.005959f
C46 B.n18 VSUBS 0.005959f
C47 B.n19 VSUBS 0.005959f
C48 B.n20 VSUBS 0.005959f
C49 B.n21 VSUBS 0.005959f
C50 B.n22 VSUBS 0.005959f
C51 B.n23 VSUBS 0.005959f
C52 B.n24 VSUBS 0.005959f
C53 B.n25 VSUBS 0.005959f
C54 B.n26 VSUBS 0.005959f
C55 B.n27 VSUBS 0.005959f
C56 B.n28 VSUBS 0.005959f
C57 B.n29 VSUBS 0.005959f
C58 B.n30 VSUBS 0.005959f
C59 B.n31 VSUBS 0.005959f
C60 B.n32 VSUBS 0.005959f
C61 B.n33 VSUBS 0.005959f
C62 B.n34 VSUBS 0.005959f
C63 B.n35 VSUBS 0.005959f
C64 B.n36 VSUBS 0.005609f
C65 B.n37 VSUBS 0.005959f
C66 B.t5 VSUBS 0.347668f
C67 B.t4 VSUBS 0.366098f
C68 B.t3 VSUBS 1.32225f
C69 B.n38 VSUBS 0.195127f
C70 B.n39 VSUBS 0.0616f
C71 B.n40 VSUBS 0.013807f
C72 B.n41 VSUBS 0.005959f
C73 B.n42 VSUBS 0.005959f
C74 B.n43 VSUBS 0.005959f
C75 B.n44 VSUBS 0.005959f
C76 B.t2 VSUBS 0.347661f
C77 B.t1 VSUBS 0.366092f
C78 B.t0 VSUBS 1.32225f
C79 B.n45 VSUBS 0.195133f
C80 B.n46 VSUBS 0.061607f
C81 B.n47 VSUBS 0.005959f
C82 B.n48 VSUBS 0.005959f
C83 B.n49 VSUBS 0.005959f
C84 B.n50 VSUBS 0.005959f
C85 B.n51 VSUBS 0.005959f
C86 B.n52 VSUBS 0.005959f
C87 B.n53 VSUBS 0.005959f
C88 B.n54 VSUBS 0.005959f
C89 B.n55 VSUBS 0.005959f
C90 B.n56 VSUBS 0.005959f
C91 B.n57 VSUBS 0.005959f
C92 B.n58 VSUBS 0.005959f
C93 B.n59 VSUBS 0.005959f
C94 B.n60 VSUBS 0.005959f
C95 B.n61 VSUBS 0.005959f
C96 B.n62 VSUBS 0.005959f
C97 B.n63 VSUBS 0.005959f
C98 B.n64 VSUBS 0.005959f
C99 B.n65 VSUBS 0.005959f
C100 B.n66 VSUBS 0.005959f
C101 B.n67 VSUBS 0.005959f
C102 B.n68 VSUBS 0.013149f
C103 B.n69 VSUBS 0.005959f
C104 B.n70 VSUBS 0.005959f
C105 B.n71 VSUBS 0.005959f
C106 B.n72 VSUBS 0.005959f
C107 B.n73 VSUBS 0.005959f
C108 B.n74 VSUBS 0.005959f
C109 B.n75 VSUBS 0.005959f
C110 B.n76 VSUBS 0.005959f
C111 B.n77 VSUBS 0.005959f
C112 B.n78 VSUBS 0.005959f
C113 B.n79 VSUBS 0.005959f
C114 B.n80 VSUBS 0.005959f
C115 B.n81 VSUBS 0.005959f
C116 B.n82 VSUBS 0.005959f
C117 B.n83 VSUBS 0.005959f
C118 B.n84 VSUBS 0.005959f
C119 B.n85 VSUBS 0.005959f
C120 B.n86 VSUBS 0.005959f
C121 B.n87 VSUBS 0.005959f
C122 B.n88 VSUBS 0.005959f
C123 B.n89 VSUBS 0.005959f
C124 B.n90 VSUBS 0.005959f
C125 B.n91 VSUBS 0.005959f
C126 B.n92 VSUBS 0.005959f
C127 B.n93 VSUBS 0.005959f
C128 B.n94 VSUBS 0.013149f
C129 B.n95 VSUBS 0.005959f
C130 B.n96 VSUBS 0.005959f
C131 B.n97 VSUBS 0.005959f
C132 B.n98 VSUBS 0.005959f
C133 B.n99 VSUBS 0.005959f
C134 B.n100 VSUBS 0.005959f
C135 B.n101 VSUBS 0.005959f
C136 B.n102 VSUBS 0.005959f
C137 B.n103 VSUBS 0.005959f
C138 B.n104 VSUBS 0.005959f
C139 B.n105 VSUBS 0.005959f
C140 B.n106 VSUBS 0.005959f
C141 B.n107 VSUBS 0.005959f
C142 B.n108 VSUBS 0.005959f
C143 B.n109 VSUBS 0.005959f
C144 B.n110 VSUBS 0.005959f
C145 B.n111 VSUBS 0.005959f
C146 B.n112 VSUBS 0.005959f
C147 B.n113 VSUBS 0.005959f
C148 B.n114 VSUBS 0.005959f
C149 B.n115 VSUBS 0.005959f
C150 B.n116 VSUBS 0.005959f
C151 B.t7 VSUBS 0.347661f
C152 B.t8 VSUBS 0.366092f
C153 B.t6 VSUBS 1.32225f
C154 B.n117 VSUBS 0.195133f
C155 B.n118 VSUBS 0.061607f
C156 B.n119 VSUBS 0.005959f
C157 B.n120 VSUBS 0.005959f
C158 B.n121 VSUBS 0.005959f
C159 B.n122 VSUBS 0.005959f
C160 B.t10 VSUBS 0.347668f
C161 B.t11 VSUBS 0.366098f
C162 B.t9 VSUBS 1.32225f
C163 B.n123 VSUBS 0.195127f
C164 B.n124 VSUBS 0.0616f
C165 B.n125 VSUBS 0.013807f
C166 B.n126 VSUBS 0.005959f
C167 B.n127 VSUBS 0.005959f
C168 B.n128 VSUBS 0.005959f
C169 B.n129 VSUBS 0.005959f
C170 B.n130 VSUBS 0.005959f
C171 B.n131 VSUBS 0.005959f
C172 B.n132 VSUBS 0.005959f
C173 B.n133 VSUBS 0.005959f
C174 B.n134 VSUBS 0.005959f
C175 B.n135 VSUBS 0.005959f
C176 B.n136 VSUBS 0.005959f
C177 B.n137 VSUBS 0.005959f
C178 B.n138 VSUBS 0.005959f
C179 B.n139 VSUBS 0.005959f
C180 B.n140 VSUBS 0.005959f
C181 B.n141 VSUBS 0.005959f
C182 B.n142 VSUBS 0.005959f
C183 B.n143 VSUBS 0.005959f
C184 B.n144 VSUBS 0.005959f
C185 B.n145 VSUBS 0.005959f
C186 B.n146 VSUBS 0.005959f
C187 B.n147 VSUBS 0.013149f
C188 B.n148 VSUBS 0.005959f
C189 B.n149 VSUBS 0.005959f
C190 B.n150 VSUBS 0.005959f
C191 B.n151 VSUBS 0.005959f
C192 B.n152 VSUBS 0.005959f
C193 B.n153 VSUBS 0.005959f
C194 B.n154 VSUBS 0.005959f
C195 B.n155 VSUBS 0.005959f
C196 B.n156 VSUBS 0.005959f
C197 B.n157 VSUBS 0.005959f
C198 B.n158 VSUBS 0.005959f
C199 B.n159 VSUBS 0.005959f
C200 B.n160 VSUBS 0.005959f
C201 B.n161 VSUBS 0.005959f
C202 B.n162 VSUBS 0.005959f
C203 B.n163 VSUBS 0.005959f
C204 B.n164 VSUBS 0.005959f
C205 B.n165 VSUBS 0.005959f
C206 B.n166 VSUBS 0.005959f
C207 B.n167 VSUBS 0.005959f
C208 B.n168 VSUBS 0.005959f
C209 B.n169 VSUBS 0.005959f
C210 B.n170 VSUBS 0.005959f
C211 B.n171 VSUBS 0.005959f
C212 B.n172 VSUBS 0.005959f
C213 B.n173 VSUBS 0.005959f
C214 B.n174 VSUBS 0.005959f
C215 B.n175 VSUBS 0.005959f
C216 B.n176 VSUBS 0.005959f
C217 B.n177 VSUBS 0.005959f
C218 B.n178 VSUBS 0.005959f
C219 B.n179 VSUBS 0.005959f
C220 B.n180 VSUBS 0.005959f
C221 B.n181 VSUBS 0.005959f
C222 B.n182 VSUBS 0.005959f
C223 B.n183 VSUBS 0.005959f
C224 B.n184 VSUBS 0.005959f
C225 B.n185 VSUBS 0.005959f
C226 B.n186 VSUBS 0.005959f
C227 B.n187 VSUBS 0.005959f
C228 B.n188 VSUBS 0.005959f
C229 B.n189 VSUBS 0.005959f
C230 B.n190 VSUBS 0.005959f
C231 B.n191 VSUBS 0.005959f
C232 B.n192 VSUBS 0.005959f
C233 B.n193 VSUBS 0.005959f
C234 B.n194 VSUBS 0.005959f
C235 B.n195 VSUBS 0.005959f
C236 B.n196 VSUBS 0.013149f
C237 B.n197 VSUBS 0.014193f
C238 B.n198 VSUBS 0.014193f
C239 B.n199 VSUBS 0.005959f
C240 B.n200 VSUBS 0.005959f
C241 B.n201 VSUBS 0.005959f
C242 B.n202 VSUBS 0.005959f
C243 B.n203 VSUBS 0.005959f
C244 B.n204 VSUBS 0.005959f
C245 B.n205 VSUBS 0.005959f
C246 B.n206 VSUBS 0.005959f
C247 B.n207 VSUBS 0.005959f
C248 B.n208 VSUBS 0.005959f
C249 B.n209 VSUBS 0.005959f
C250 B.n210 VSUBS 0.005959f
C251 B.n211 VSUBS 0.005959f
C252 B.n212 VSUBS 0.005959f
C253 B.n213 VSUBS 0.005959f
C254 B.n214 VSUBS 0.005959f
C255 B.n215 VSUBS 0.005959f
C256 B.n216 VSUBS 0.005959f
C257 B.n217 VSUBS 0.005959f
C258 B.n218 VSUBS 0.005959f
C259 B.n219 VSUBS 0.005959f
C260 B.n220 VSUBS 0.005959f
C261 B.n221 VSUBS 0.005959f
C262 B.n222 VSUBS 0.005959f
C263 B.n223 VSUBS 0.005959f
C264 B.n224 VSUBS 0.005959f
C265 B.n225 VSUBS 0.005959f
C266 B.n226 VSUBS 0.005959f
C267 B.n227 VSUBS 0.005959f
C268 B.n228 VSUBS 0.005959f
C269 B.n229 VSUBS 0.005959f
C270 B.n230 VSUBS 0.005959f
C271 B.n231 VSUBS 0.005959f
C272 B.n232 VSUBS 0.005959f
C273 B.n233 VSUBS 0.005959f
C274 B.n234 VSUBS 0.005959f
C275 B.n235 VSUBS 0.005959f
C276 B.n236 VSUBS 0.005959f
C277 B.n237 VSUBS 0.005959f
C278 B.n238 VSUBS 0.005959f
C279 B.n239 VSUBS 0.005959f
C280 B.n240 VSUBS 0.005959f
C281 B.n241 VSUBS 0.005959f
C282 B.n242 VSUBS 0.005959f
C283 B.n243 VSUBS 0.005959f
C284 B.n244 VSUBS 0.005959f
C285 B.n245 VSUBS 0.005959f
C286 B.n246 VSUBS 0.005959f
C287 B.n247 VSUBS 0.005959f
C288 B.n248 VSUBS 0.005959f
C289 B.n249 VSUBS 0.005959f
C290 B.n250 VSUBS 0.005959f
C291 B.n251 VSUBS 0.005959f
C292 B.n252 VSUBS 0.005959f
C293 B.n253 VSUBS 0.005959f
C294 B.n254 VSUBS 0.005959f
C295 B.n255 VSUBS 0.005959f
C296 B.n256 VSUBS 0.005959f
C297 B.n257 VSUBS 0.005959f
C298 B.n258 VSUBS 0.005959f
C299 B.n259 VSUBS 0.005959f
C300 B.n260 VSUBS 0.005609f
C301 B.n261 VSUBS 0.005959f
C302 B.n262 VSUBS 0.005959f
C303 B.n263 VSUBS 0.00333f
C304 B.n264 VSUBS 0.005959f
C305 B.n265 VSUBS 0.005959f
C306 B.n266 VSUBS 0.005959f
C307 B.n267 VSUBS 0.005959f
C308 B.n268 VSUBS 0.005959f
C309 B.n269 VSUBS 0.005959f
C310 B.n270 VSUBS 0.005959f
C311 B.n271 VSUBS 0.005959f
C312 B.n272 VSUBS 0.005959f
C313 B.n273 VSUBS 0.005959f
C314 B.n274 VSUBS 0.005959f
C315 B.n275 VSUBS 0.005959f
C316 B.n276 VSUBS 0.00333f
C317 B.n277 VSUBS 0.013807f
C318 B.n278 VSUBS 0.005609f
C319 B.n279 VSUBS 0.005959f
C320 B.n280 VSUBS 0.005959f
C321 B.n281 VSUBS 0.005959f
C322 B.n282 VSUBS 0.005959f
C323 B.n283 VSUBS 0.005959f
C324 B.n284 VSUBS 0.005959f
C325 B.n285 VSUBS 0.005959f
C326 B.n286 VSUBS 0.005959f
C327 B.n287 VSUBS 0.005959f
C328 B.n288 VSUBS 0.005959f
C329 B.n289 VSUBS 0.005959f
C330 B.n290 VSUBS 0.005959f
C331 B.n291 VSUBS 0.005959f
C332 B.n292 VSUBS 0.005959f
C333 B.n293 VSUBS 0.005959f
C334 B.n294 VSUBS 0.005959f
C335 B.n295 VSUBS 0.005959f
C336 B.n296 VSUBS 0.005959f
C337 B.n297 VSUBS 0.005959f
C338 B.n298 VSUBS 0.005959f
C339 B.n299 VSUBS 0.005959f
C340 B.n300 VSUBS 0.005959f
C341 B.n301 VSUBS 0.005959f
C342 B.n302 VSUBS 0.005959f
C343 B.n303 VSUBS 0.005959f
C344 B.n304 VSUBS 0.005959f
C345 B.n305 VSUBS 0.005959f
C346 B.n306 VSUBS 0.005959f
C347 B.n307 VSUBS 0.005959f
C348 B.n308 VSUBS 0.005959f
C349 B.n309 VSUBS 0.005959f
C350 B.n310 VSUBS 0.005959f
C351 B.n311 VSUBS 0.005959f
C352 B.n312 VSUBS 0.005959f
C353 B.n313 VSUBS 0.005959f
C354 B.n314 VSUBS 0.005959f
C355 B.n315 VSUBS 0.005959f
C356 B.n316 VSUBS 0.005959f
C357 B.n317 VSUBS 0.005959f
C358 B.n318 VSUBS 0.005959f
C359 B.n319 VSUBS 0.005959f
C360 B.n320 VSUBS 0.005959f
C361 B.n321 VSUBS 0.005959f
C362 B.n322 VSUBS 0.005959f
C363 B.n323 VSUBS 0.005959f
C364 B.n324 VSUBS 0.005959f
C365 B.n325 VSUBS 0.005959f
C366 B.n326 VSUBS 0.005959f
C367 B.n327 VSUBS 0.005959f
C368 B.n328 VSUBS 0.005959f
C369 B.n329 VSUBS 0.005959f
C370 B.n330 VSUBS 0.005959f
C371 B.n331 VSUBS 0.005959f
C372 B.n332 VSUBS 0.005959f
C373 B.n333 VSUBS 0.005959f
C374 B.n334 VSUBS 0.005959f
C375 B.n335 VSUBS 0.005959f
C376 B.n336 VSUBS 0.005959f
C377 B.n337 VSUBS 0.005959f
C378 B.n338 VSUBS 0.005959f
C379 B.n339 VSUBS 0.005959f
C380 B.n340 VSUBS 0.005959f
C381 B.n341 VSUBS 0.014193f
C382 B.n342 VSUBS 0.014193f
C383 B.n343 VSUBS 0.013149f
C384 B.n344 VSUBS 0.005959f
C385 B.n345 VSUBS 0.005959f
C386 B.n346 VSUBS 0.005959f
C387 B.n347 VSUBS 0.005959f
C388 B.n348 VSUBS 0.005959f
C389 B.n349 VSUBS 0.005959f
C390 B.n350 VSUBS 0.005959f
C391 B.n351 VSUBS 0.005959f
C392 B.n352 VSUBS 0.005959f
C393 B.n353 VSUBS 0.005959f
C394 B.n354 VSUBS 0.005959f
C395 B.n355 VSUBS 0.005959f
C396 B.n356 VSUBS 0.005959f
C397 B.n357 VSUBS 0.005959f
C398 B.n358 VSUBS 0.005959f
C399 B.n359 VSUBS 0.005959f
C400 B.n360 VSUBS 0.005959f
C401 B.n361 VSUBS 0.005959f
C402 B.n362 VSUBS 0.005959f
C403 B.n363 VSUBS 0.005959f
C404 B.n364 VSUBS 0.005959f
C405 B.n365 VSUBS 0.005959f
C406 B.n366 VSUBS 0.005959f
C407 B.n367 VSUBS 0.005959f
C408 B.n368 VSUBS 0.005959f
C409 B.n369 VSUBS 0.005959f
C410 B.n370 VSUBS 0.005959f
C411 B.n371 VSUBS 0.005959f
C412 B.n372 VSUBS 0.005959f
C413 B.n373 VSUBS 0.005959f
C414 B.n374 VSUBS 0.005959f
C415 B.n375 VSUBS 0.005959f
C416 B.n376 VSUBS 0.005959f
C417 B.n377 VSUBS 0.005959f
C418 B.n378 VSUBS 0.005959f
C419 B.n379 VSUBS 0.005959f
C420 B.n380 VSUBS 0.005959f
C421 B.n381 VSUBS 0.005959f
C422 B.n382 VSUBS 0.005959f
C423 B.n383 VSUBS 0.005959f
C424 B.n384 VSUBS 0.005959f
C425 B.n385 VSUBS 0.005959f
C426 B.n386 VSUBS 0.005959f
C427 B.n387 VSUBS 0.005959f
C428 B.n388 VSUBS 0.005959f
C429 B.n389 VSUBS 0.005959f
C430 B.n390 VSUBS 0.005959f
C431 B.n391 VSUBS 0.005959f
C432 B.n392 VSUBS 0.005959f
C433 B.n393 VSUBS 0.005959f
C434 B.n394 VSUBS 0.005959f
C435 B.n395 VSUBS 0.005959f
C436 B.n396 VSUBS 0.005959f
C437 B.n397 VSUBS 0.005959f
C438 B.n398 VSUBS 0.005959f
C439 B.n399 VSUBS 0.005959f
C440 B.n400 VSUBS 0.005959f
C441 B.n401 VSUBS 0.005959f
C442 B.n402 VSUBS 0.005959f
C443 B.n403 VSUBS 0.005959f
C444 B.n404 VSUBS 0.005959f
C445 B.n405 VSUBS 0.005959f
C446 B.n406 VSUBS 0.005959f
C447 B.n407 VSUBS 0.005959f
C448 B.n408 VSUBS 0.005959f
C449 B.n409 VSUBS 0.005959f
C450 B.n410 VSUBS 0.005959f
C451 B.n411 VSUBS 0.005959f
C452 B.n412 VSUBS 0.005959f
C453 B.n413 VSUBS 0.005959f
C454 B.n414 VSUBS 0.005959f
C455 B.n415 VSUBS 0.005959f
C456 B.n416 VSUBS 0.005959f
C457 B.n417 VSUBS 0.005959f
C458 B.n418 VSUBS 0.005959f
C459 B.n419 VSUBS 0.005959f
C460 B.n420 VSUBS 0.005959f
C461 B.n421 VSUBS 0.013875f
C462 B.n422 VSUBS 0.013467f
C463 B.n423 VSUBS 0.014193f
C464 B.n424 VSUBS 0.005959f
C465 B.n425 VSUBS 0.005959f
C466 B.n426 VSUBS 0.005959f
C467 B.n427 VSUBS 0.005959f
C468 B.n428 VSUBS 0.005959f
C469 B.n429 VSUBS 0.005959f
C470 B.n430 VSUBS 0.005959f
C471 B.n431 VSUBS 0.005959f
C472 B.n432 VSUBS 0.005959f
C473 B.n433 VSUBS 0.005959f
C474 B.n434 VSUBS 0.005959f
C475 B.n435 VSUBS 0.005959f
C476 B.n436 VSUBS 0.005959f
C477 B.n437 VSUBS 0.005959f
C478 B.n438 VSUBS 0.005959f
C479 B.n439 VSUBS 0.005959f
C480 B.n440 VSUBS 0.005959f
C481 B.n441 VSUBS 0.005959f
C482 B.n442 VSUBS 0.005959f
C483 B.n443 VSUBS 0.005959f
C484 B.n444 VSUBS 0.005959f
C485 B.n445 VSUBS 0.005959f
C486 B.n446 VSUBS 0.005959f
C487 B.n447 VSUBS 0.005959f
C488 B.n448 VSUBS 0.005959f
C489 B.n449 VSUBS 0.005959f
C490 B.n450 VSUBS 0.005959f
C491 B.n451 VSUBS 0.005959f
C492 B.n452 VSUBS 0.005959f
C493 B.n453 VSUBS 0.005959f
C494 B.n454 VSUBS 0.005959f
C495 B.n455 VSUBS 0.005959f
C496 B.n456 VSUBS 0.005959f
C497 B.n457 VSUBS 0.005959f
C498 B.n458 VSUBS 0.005959f
C499 B.n459 VSUBS 0.005959f
C500 B.n460 VSUBS 0.005959f
C501 B.n461 VSUBS 0.005959f
C502 B.n462 VSUBS 0.005959f
C503 B.n463 VSUBS 0.005959f
C504 B.n464 VSUBS 0.005959f
C505 B.n465 VSUBS 0.005959f
C506 B.n466 VSUBS 0.005959f
C507 B.n467 VSUBS 0.005959f
C508 B.n468 VSUBS 0.005959f
C509 B.n469 VSUBS 0.005959f
C510 B.n470 VSUBS 0.005959f
C511 B.n471 VSUBS 0.005959f
C512 B.n472 VSUBS 0.005959f
C513 B.n473 VSUBS 0.005959f
C514 B.n474 VSUBS 0.005959f
C515 B.n475 VSUBS 0.005959f
C516 B.n476 VSUBS 0.005959f
C517 B.n477 VSUBS 0.005959f
C518 B.n478 VSUBS 0.005959f
C519 B.n479 VSUBS 0.005959f
C520 B.n480 VSUBS 0.005959f
C521 B.n481 VSUBS 0.005959f
C522 B.n482 VSUBS 0.005959f
C523 B.n483 VSUBS 0.005959f
C524 B.n484 VSUBS 0.005959f
C525 B.n485 VSUBS 0.005959f
C526 B.n486 VSUBS 0.005609f
C527 B.n487 VSUBS 0.013807f
C528 B.n488 VSUBS 0.00333f
C529 B.n489 VSUBS 0.005959f
C530 B.n490 VSUBS 0.005959f
C531 B.n491 VSUBS 0.005959f
C532 B.n492 VSUBS 0.005959f
C533 B.n493 VSUBS 0.005959f
C534 B.n494 VSUBS 0.005959f
C535 B.n495 VSUBS 0.005959f
C536 B.n496 VSUBS 0.005959f
C537 B.n497 VSUBS 0.005959f
C538 B.n498 VSUBS 0.005959f
C539 B.n499 VSUBS 0.005959f
C540 B.n500 VSUBS 0.005959f
C541 B.n501 VSUBS 0.00333f
C542 B.n502 VSUBS 0.005959f
C543 B.n503 VSUBS 0.005959f
C544 B.n504 VSUBS 0.005959f
C545 B.n505 VSUBS 0.005959f
C546 B.n506 VSUBS 0.005959f
C547 B.n507 VSUBS 0.005959f
C548 B.n508 VSUBS 0.005959f
C549 B.n509 VSUBS 0.005959f
C550 B.n510 VSUBS 0.005959f
C551 B.n511 VSUBS 0.005959f
C552 B.n512 VSUBS 0.005959f
C553 B.n513 VSUBS 0.005959f
C554 B.n514 VSUBS 0.005959f
C555 B.n515 VSUBS 0.005959f
C556 B.n516 VSUBS 0.005959f
C557 B.n517 VSUBS 0.005959f
C558 B.n518 VSUBS 0.005959f
C559 B.n519 VSUBS 0.005959f
C560 B.n520 VSUBS 0.005959f
C561 B.n521 VSUBS 0.005959f
C562 B.n522 VSUBS 0.005959f
C563 B.n523 VSUBS 0.005959f
C564 B.n524 VSUBS 0.005959f
C565 B.n525 VSUBS 0.005959f
C566 B.n526 VSUBS 0.005959f
C567 B.n527 VSUBS 0.005959f
C568 B.n528 VSUBS 0.005959f
C569 B.n529 VSUBS 0.005959f
C570 B.n530 VSUBS 0.005959f
C571 B.n531 VSUBS 0.005959f
C572 B.n532 VSUBS 0.005959f
C573 B.n533 VSUBS 0.005959f
C574 B.n534 VSUBS 0.005959f
C575 B.n535 VSUBS 0.005959f
C576 B.n536 VSUBS 0.005959f
C577 B.n537 VSUBS 0.005959f
C578 B.n538 VSUBS 0.005959f
C579 B.n539 VSUBS 0.005959f
C580 B.n540 VSUBS 0.005959f
C581 B.n541 VSUBS 0.005959f
C582 B.n542 VSUBS 0.005959f
C583 B.n543 VSUBS 0.005959f
C584 B.n544 VSUBS 0.005959f
C585 B.n545 VSUBS 0.005959f
C586 B.n546 VSUBS 0.005959f
C587 B.n547 VSUBS 0.005959f
C588 B.n548 VSUBS 0.005959f
C589 B.n549 VSUBS 0.005959f
C590 B.n550 VSUBS 0.005959f
C591 B.n551 VSUBS 0.005959f
C592 B.n552 VSUBS 0.005959f
C593 B.n553 VSUBS 0.005959f
C594 B.n554 VSUBS 0.005959f
C595 B.n555 VSUBS 0.005959f
C596 B.n556 VSUBS 0.005959f
C597 B.n557 VSUBS 0.005959f
C598 B.n558 VSUBS 0.005959f
C599 B.n559 VSUBS 0.005959f
C600 B.n560 VSUBS 0.005959f
C601 B.n561 VSUBS 0.005959f
C602 B.n562 VSUBS 0.005959f
C603 B.n563 VSUBS 0.005959f
C604 B.n564 VSUBS 0.005959f
C605 B.n565 VSUBS 0.005959f
C606 B.n566 VSUBS 0.014193f
C607 B.n567 VSUBS 0.013149f
C608 B.n568 VSUBS 0.013149f
C609 B.n569 VSUBS 0.005959f
C610 B.n570 VSUBS 0.005959f
C611 B.n571 VSUBS 0.005959f
C612 B.n572 VSUBS 0.005959f
C613 B.n573 VSUBS 0.005959f
C614 B.n574 VSUBS 0.005959f
C615 B.n575 VSUBS 0.005959f
C616 B.n576 VSUBS 0.005959f
C617 B.n577 VSUBS 0.005959f
C618 B.n578 VSUBS 0.005959f
C619 B.n579 VSUBS 0.005959f
C620 B.n580 VSUBS 0.005959f
C621 B.n581 VSUBS 0.005959f
C622 B.n582 VSUBS 0.005959f
C623 B.n583 VSUBS 0.005959f
C624 B.n584 VSUBS 0.005959f
C625 B.n585 VSUBS 0.005959f
C626 B.n586 VSUBS 0.005959f
C627 B.n587 VSUBS 0.005959f
C628 B.n588 VSUBS 0.005959f
C629 B.n589 VSUBS 0.005959f
C630 B.n590 VSUBS 0.005959f
C631 B.n591 VSUBS 0.005959f
C632 B.n592 VSUBS 0.005959f
C633 B.n593 VSUBS 0.005959f
C634 B.n594 VSUBS 0.005959f
C635 B.n595 VSUBS 0.005959f
C636 B.n596 VSUBS 0.005959f
C637 B.n597 VSUBS 0.005959f
C638 B.n598 VSUBS 0.005959f
C639 B.n599 VSUBS 0.005959f
C640 B.n600 VSUBS 0.005959f
C641 B.n601 VSUBS 0.005959f
C642 B.n602 VSUBS 0.005959f
C643 B.n603 VSUBS 0.005959f
C644 B.n604 VSUBS 0.005959f
C645 B.n605 VSUBS 0.005959f
C646 B.n606 VSUBS 0.005959f
C647 B.n607 VSUBS 0.013494f
C648 VDD2.t1 VSUBS 2.63782f
C649 VDD2.t0 VSUBS 2.05508f
C650 VDD2.n0 VSUBS 3.37314f
C651 VN.t0 VSUBS 3.96781f
C652 VN.t1 VSUBS 4.68026f
C653 VDD1.t0 VSUBS 2.06602f
C654 VDD1.t1 VSUBS 2.68163f
C655 VTAIL.t2 VSUBS 2.80464f
C656 VTAIL.n0 VSUBS 2.83869f
C657 VTAIL.t1 VSUBS 2.80466f
C658 VTAIL.n1 VSUBS 2.89591f
C659 VTAIL.t3 VSUBS 2.80464f
C660 VTAIL.n2 VSUBS 2.64479f
C661 VTAIL.t0 VSUBS 2.80464f
C662 VTAIL.n3 VSUBS 2.53173f
C663 VP.t0 VSUBS 4.09127f
C664 VP.t1 VSUBS 4.82813f
C665 VP.n0 VSUBS 5.57418f
.ends

