* NGSPICE file created from diff_pair_sample_0123.ext - technology: sky130A

.subckt diff_pair_sample_0123 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9491 pd=26.16 as=4.9491 ps=26.16 w=12.69 l=0.74
X1 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.9491 pd=26.16 as=4.9491 ps=26.16 w=12.69 l=0.74
X2 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=4.9491 pd=26.16 as=0 ps=0 w=12.69 l=0.74
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=4.9491 pd=26.16 as=0 ps=0 w=12.69 l=0.74
X4 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.9491 pd=26.16 as=4.9491 ps=26.16 w=12.69 l=0.74
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=4.9491 pd=26.16 as=0 ps=0 w=12.69 l=0.74
X6 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.9491 pd=26.16 as=4.9491 ps=26.16 w=12.69 l=0.74
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.9491 pd=26.16 as=0 ps=0 w=12.69 l=0.74
R0 VP.n0 VP.t0 668.255
R1 VP.n0 VP.t1 627.994
R2 VP VP.n0 0.0516364
R3 VTAIL.n278 VTAIL.n277 289.615
R4 VTAIL.n68 VTAIL.n67 289.615
R5 VTAIL.n208 VTAIL.n207 289.615
R6 VTAIL.n138 VTAIL.n137 289.615
R7 VTAIL.n232 VTAIL.n231 185
R8 VTAIL.n237 VTAIL.n236 185
R9 VTAIL.n239 VTAIL.n238 185
R10 VTAIL.n228 VTAIL.n227 185
R11 VTAIL.n245 VTAIL.n244 185
R12 VTAIL.n247 VTAIL.n246 185
R13 VTAIL.n224 VTAIL.n223 185
R14 VTAIL.n253 VTAIL.n252 185
R15 VTAIL.n255 VTAIL.n254 185
R16 VTAIL.n220 VTAIL.n219 185
R17 VTAIL.n261 VTAIL.n260 185
R18 VTAIL.n263 VTAIL.n262 185
R19 VTAIL.n216 VTAIL.n215 185
R20 VTAIL.n269 VTAIL.n268 185
R21 VTAIL.n271 VTAIL.n270 185
R22 VTAIL.n212 VTAIL.n211 185
R23 VTAIL.n277 VTAIL.n276 185
R24 VTAIL.n22 VTAIL.n21 185
R25 VTAIL.n27 VTAIL.n26 185
R26 VTAIL.n29 VTAIL.n28 185
R27 VTAIL.n18 VTAIL.n17 185
R28 VTAIL.n35 VTAIL.n34 185
R29 VTAIL.n37 VTAIL.n36 185
R30 VTAIL.n14 VTAIL.n13 185
R31 VTAIL.n43 VTAIL.n42 185
R32 VTAIL.n45 VTAIL.n44 185
R33 VTAIL.n10 VTAIL.n9 185
R34 VTAIL.n51 VTAIL.n50 185
R35 VTAIL.n53 VTAIL.n52 185
R36 VTAIL.n6 VTAIL.n5 185
R37 VTAIL.n59 VTAIL.n58 185
R38 VTAIL.n61 VTAIL.n60 185
R39 VTAIL.n2 VTAIL.n1 185
R40 VTAIL.n67 VTAIL.n66 185
R41 VTAIL.n207 VTAIL.n206 185
R42 VTAIL.n142 VTAIL.n141 185
R43 VTAIL.n201 VTAIL.n200 185
R44 VTAIL.n199 VTAIL.n198 185
R45 VTAIL.n146 VTAIL.n145 185
R46 VTAIL.n193 VTAIL.n192 185
R47 VTAIL.n191 VTAIL.n190 185
R48 VTAIL.n150 VTAIL.n149 185
R49 VTAIL.n185 VTAIL.n184 185
R50 VTAIL.n183 VTAIL.n182 185
R51 VTAIL.n154 VTAIL.n153 185
R52 VTAIL.n177 VTAIL.n176 185
R53 VTAIL.n175 VTAIL.n174 185
R54 VTAIL.n158 VTAIL.n157 185
R55 VTAIL.n169 VTAIL.n168 185
R56 VTAIL.n167 VTAIL.n166 185
R57 VTAIL.n162 VTAIL.n161 185
R58 VTAIL.n137 VTAIL.n136 185
R59 VTAIL.n72 VTAIL.n71 185
R60 VTAIL.n131 VTAIL.n130 185
R61 VTAIL.n129 VTAIL.n128 185
R62 VTAIL.n76 VTAIL.n75 185
R63 VTAIL.n123 VTAIL.n122 185
R64 VTAIL.n121 VTAIL.n120 185
R65 VTAIL.n80 VTAIL.n79 185
R66 VTAIL.n115 VTAIL.n114 185
R67 VTAIL.n113 VTAIL.n112 185
R68 VTAIL.n84 VTAIL.n83 185
R69 VTAIL.n107 VTAIL.n106 185
R70 VTAIL.n105 VTAIL.n104 185
R71 VTAIL.n88 VTAIL.n87 185
R72 VTAIL.n99 VTAIL.n98 185
R73 VTAIL.n97 VTAIL.n96 185
R74 VTAIL.n92 VTAIL.n91 185
R75 VTAIL.n233 VTAIL.t1 147.659
R76 VTAIL.n23 VTAIL.t2 147.659
R77 VTAIL.n163 VTAIL.t3 147.659
R78 VTAIL.n93 VTAIL.t0 147.659
R79 VTAIL.n237 VTAIL.n231 104.615
R80 VTAIL.n238 VTAIL.n237 104.615
R81 VTAIL.n238 VTAIL.n227 104.615
R82 VTAIL.n245 VTAIL.n227 104.615
R83 VTAIL.n246 VTAIL.n245 104.615
R84 VTAIL.n246 VTAIL.n223 104.615
R85 VTAIL.n253 VTAIL.n223 104.615
R86 VTAIL.n254 VTAIL.n253 104.615
R87 VTAIL.n254 VTAIL.n219 104.615
R88 VTAIL.n261 VTAIL.n219 104.615
R89 VTAIL.n262 VTAIL.n261 104.615
R90 VTAIL.n262 VTAIL.n215 104.615
R91 VTAIL.n269 VTAIL.n215 104.615
R92 VTAIL.n270 VTAIL.n269 104.615
R93 VTAIL.n270 VTAIL.n211 104.615
R94 VTAIL.n277 VTAIL.n211 104.615
R95 VTAIL.n27 VTAIL.n21 104.615
R96 VTAIL.n28 VTAIL.n27 104.615
R97 VTAIL.n28 VTAIL.n17 104.615
R98 VTAIL.n35 VTAIL.n17 104.615
R99 VTAIL.n36 VTAIL.n35 104.615
R100 VTAIL.n36 VTAIL.n13 104.615
R101 VTAIL.n43 VTAIL.n13 104.615
R102 VTAIL.n44 VTAIL.n43 104.615
R103 VTAIL.n44 VTAIL.n9 104.615
R104 VTAIL.n51 VTAIL.n9 104.615
R105 VTAIL.n52 VTAIL.n51 104.615
R106 VTAIL.n52 VTAIL.n5 104.615
R107 VTAIL.n59 VTAIL.n5 104.615
R108 VTAIL.n60 VTAIL.n59 104.615
R109 VTAIL.n60 VTAIL.n1 104.615
R110 VTAIL.n67 VTAIL.n1 104.615
R111 VTAIL.n207 VTAIL.n141 104.615
R112 VTAIL.n200 VTAIL.n141 104.615
R113 VTAIL.n200 VTAIL.n199 104.615
R114 VTAIL.n199 VTAIL.n145 104.615
R115 VTAIL.n192 VTAIL.n145 104.615
R116 VTAIL.n192 VTAIL.n191 104.615
R117 VTAIL.n191 VTAIL.n149 104.615
R118 VTAIL.n184 VTAIL.n149 104.615
R119 VTAIL.n184 VTAIL.n183 104.615
R120 VTAIL.n183 VTAIL.n153 104.615
R121 VTAIL.n176 VTAIL.n153 104.615
R122 VTAIL.n176 VTAIL.n175 104.615
R123 VTAIL.n175 VTAIL.n157 104.615
R124 VTAIL.n168 VTAIL.n157 104.615
R125 VTAIL.n168 VTAIL.n167 104.615
R126 VTAIL.n167 VTAIL.n161 104.615
R127 VTAIL.n137 VTAIL.n71 104.615
R128 VTAIL.n130 VTAIL.n71 104.615
R129 VTAIL.n130 VTAIL.n129 104.615
R130 VTAIL.n129 VTAIL.n75 104.615
R131 VTAIL.n122 VTAIL.n75 104.615
R132 VTAIL.n122 VTAIL.n121 104.615
R133 VTAIL.n121 VTAIL.n79 104.615
R134 VTAIL.n114 VTAIL.n79 104.615
R135 VTAIL.n114 VTAIL.n113 104.615
R136 VTAIL.n113 VTAIL.n83 104.615
R137 VTAIL.n106 VTAIL.n83 104.615
R138 VTAIL.n106 VTAIL.n105 104.615
R139 VTAIL.n105 VTAIL.n87 104.615
R140 VTAIL.n98 VTAIL.n87 104.615
R141 VTAIL.n98 VTAIL.n97 104.615
R142 VTAIL.n97 VTAIL.n91 104.615
R143 VTAIL.t1 VTAIL.n231 52.3082
R144 VTAIL.t2 VTAIL.n21 52.3082
R145 VTAIL.t3 VTAIL.n161 52.3082
R146 VTAIL.t0 VTAIL.n91 52.3082
R147 VTAIL.n279 VTAIL.n278 35.8702
R148 VTAIL.n69 VTAIL.n68 35.8702
R149 VTAIL.n209 VTAIL.n208 35.8702
R150 VTAIL.n139 VTAIL.n138 35.8702
R151 VTAIL.n139 VTAIL.n69 25.1686
R152 VTAIL.n279 VTAIL.n209 24.2462
R153 VTAIL.n233 VTAIL.n232 15.6677
R154 VTAIL.n23 VTAIL.n22 15.6677
R155 VTAIL.n163 VTAIL.n162 15.6677
R156 VTAIL.n93 VTAIL.n92 15.6677
R157 VTAIL.n236 VTAIL.n235 12.8005
R158 VTAIL.n276 VTAIL.n210 12.8005
R159 VTAIL.n26 VTAIL.n25 12.8005
R160 VTAIL.n66 VTAIL.n0 12.8005
R161 VTAIL.n206 VTAIL.n140 12.8005
R162 VTAIL.n166 VTAIL.n165 12.8005
R163 VTAIL.n136 VTAIL.n70 12.8005
R164 VTAIL.n96 VTAIL.n95 12.8005
R165 VTAIL.n239 VTAIL.n230 12.0247
R166 VTAIL.n275 VTAIL.n212 12.0247
R167 VTAIL.n29 VTAIL.n20 12.0247
R168 VTAIL.n65 VTAIL.n2 12.0247
R169 VTAIL.n205 VTAIL.n142 12.0247
R170 VTAIL.n169 VTAIL.n160 12.0247
R171 VTAIL.n135 VTAIL.n72 12.0247
R172 VTAIL.n99 VTAIL.n90 12.0247
R173 VTAIL.n240 VTAIL.n228 11.249
R174 VTAIL.n272 VTAIL.n271 11.249
R175 VTAIL.n30 VTAIL.n18 11.249
R176 VTAIL.n62 VTAIL.n61 11.249
R177 VTAIL.n202 VTAIL.n201 11.249
R178 VTAIL.n170 VTAIL.n158 11.249
R179 VTAIL.n132 VTAIL.n131 11.249
R180 VTAIL.n100 VTAIL.n88 11.249
R181 VTAIL.n244 VTAIL.n243 10.4732
R182 VTAIL.n268 VTAIL.n214 10.4732
R183 VTAIL.n34 VTAIL.n33 10.4732
R184 VTAIL.n58 VTAIL.n4 10.4732
R185 VTAIL.n198 VTAIL.n144 10.4732
R186 VTAIL.n174 VTAIL.n173 10.4732
R187 VTAIL.n128 VTAIL.n74 10.4732
R188 VTAIL.n104 VTAIL.n103 10.4732
R189 VTAIL.n247 VTAIL.n226 9.69747
R190 VTAIL.n267 VTAIL.n216 9.69747
R191 VTAIL.n37 VTAIL.n16 9.69747
R192 VTAIL.n57 VTAIL.n6 9.69747
R193 VTAIL.n197 VTAIL.n146 9.69747
R194 VTAIL.n177 VTAIL.n156 9.69747
R195 VTAIL.n127 VTAIL.n76 9.69747
R196 VTAIL.n107 VTAIL.n86 9.69747
R197 VTAIL.n274 VTAIL.n210 9.45567
R198 VTAIL.n64 VTAIL.n0 9.45567
R199 VTAIL.n204 VTAIL.n140 9.45567
R200 VTAIL.n134 VTAIL.n70 9.45567
R201 VTAIL.n257 VTAIL.n256 9.3005
R202 VTAIL.n259 VTAIL.n258 9.3005
R203 VTAIL.n218 VTAIL.n217 9.3005
R204 VTAIL.n265 VTAIL.n264 9.3005
R205 VTAIL.n267 VTAIL.n266 9.3005
R206 VTAIL.n214 VTAIL.n213 9.3005
R207 VTAIL.n273 VTAIL.n272 9.3005
R208 VTAIL.n275 VTAIL.n274 9.3005
R209 VTAIL.n251 VTAIL.n250 9.3005
R210 VTAIL.n249 VTAIL.n248 9.3005
R211 VTAIL.n226 VTAIL.n225 9.3005
R212 VTAIL.n243 VTAIL.n242 9.3005
R213 VTAIL.n241 VTAIL.n240 9.3005
R214 VTAIL.n230 VTAIL.n229 9.3005
R215 VTAIL.n235 VTAIL.n234 9.3005
R216 VTAIL.n222 VTAIL.n221 9.3005
R217 VTAIL.n47 VTAIL.n46 9.3005
R218 VTAIL.n49 VTAIL.n48 9.3005
R219 VTAIL.n8 VTAIL.n7 9.3005
R220 VTAIL.n55 VTAIL.n54 9.3005
R221 VTAIL.n57 VTAIL.n56 9.3005
R222 VTAIL.n4 VTAIL.n3 9.3005
R223 VTAIL.n63 VTAIL.n62 9.3005
R224 VTAIL.n65 VTAIL.n64 9.3005
R225 VTAIL.n41 VTAIL.n40 9.3005
R226 VTAIL.n39 VTAIL.n38 9.3005
R227 VTAIL.n16 VTAIL.n15 9.3005
R228 VTAIL.n33 VTAIL.n32 9.3005
R229 VTAIL.n31 VTAIL.n30 9.3005
R230 VTAIL.n20 VTAIL.n19 9.3005
R231 VTAIL.n25 VTAIL.n24 9.3005
R232 VTAIL.n12 VTAIL.n11 9.3005
R233 VTAIL.n205 VTAIL.n204 9.3005
R234 VTAIL.n203 VTAIL.n202 9.3005
R235 VTAIL.n144 VTAIL.n143 9.3005
R236 VTAIL.n197 VTAIL.n196 9.3005
R237 VTAIL.n195 VTAIL.n194 9.3005
R238 VTAIL.n148 VTAIL.n147 9.3005
R239 VTAIL.n189 VTAIL.n188 9.3005
R240 VTAIL.n187 VTAIL.n186 9.3005
R241 VTAIL.n152 VTAIL.n151 9.3005
R242 VTAIL.n181 VTAIL.n180 9.3005
R243 VTAIL.n179 VTAIL.n178 9.3005
R244 VTAIL.n156 VTAIL.n155 9.3005
R245 VTAIL.n173 VTAIL.n172 9.3005
R246 VTAIL.n171 VTAIL.n170 9.3005
R247 VTAIL.n160 VTAIL.n159 9.3005
R248 VTAIL.n165 VTAIL.n164 9.3005
R249 VTAIL.n119 VTAIL.n118 9.3005
R250 VTAIL.n78 VTAIL.n77 9.3005
R251 VTAIL.n125 VTAIL.n124 9.3005
R252 VTAIL.n127 VTAIL.n126 9.3005
R253 VTAIL.n74 VTAIL.n73 9.3005
R254 VTAIL.n133 VTAIL.n132 9.3005
R255 VTAIL.n135 VTAIL.n134 9.3005
R256 VTAIL.n117 VTAIL.n116 9.3005
R257 VTAIL.n82 VTAIL.n81 9.3005
R258 VTAIL.n111 VTAIL.n110 9.3005
R259 VTAIL.n109 VTAIL.n108 9.3005
R260 VTAIL.n86 VTAIL.n85 9.3005
R261 VTAIL.n103 VTAIL.n102 9.3005
R262 VTAIL.n101 VTAIL.n100 9.3005
R263 VTAIL.n90 VTAIL.n89 9.3005
R264 VTAIL.n95 VTAIL.n94 9.3005
R265 VTAIL.n248 VTAIL.n224 8.92171
R266 VTAIL.n264 VTAIL.n263 8.92171
R267 VTAIL.n38 VTAIL.n14 8.92171
R268 VTAIL.n54 VTAIL.n53 8.92171
R269 VTAIL.n194 VTAIL.n193 8.92171
R270 VTAIL.n178 VTAIL.n154 8.92171
R271 VTAIL.n124 VTAIL.n123 8.92171
R272 VTAIL.n108 VTAIL.n84 8.92171
R273 VTAIL.n252 VTAIL.n251 8.14595
R274 VTAIL.n260 VTAIL.n218 8.14595
R275 VTAIL.n42 VTAIL.n41 8.14595
R276 VTAIL.n50 VTAIL.n8 8.14595
R277 VTAIL.n190 VTAIL.n148 8.14595
R278 VTAIL.n182 VTAIL.n181 8.14595
R279 VTAIL.n120 VTAIL.n78 8.14595
R280 VTAIL.n112 VTAIL.n111 8.14595
R281 VTAIL.n255 VTAIL.n222 7.3702
R282 VTAIL.n259 VTAIL.n220 7.3702
R283 VTAIL.n45 VTAIL.n12 7.3702
R284 VTAIL.n49 VTAIL.n10 7.3702
R285 VTAIL.n189 VTAIL.n150 7.3702
R286 VTAIL.n185 VTAIL.n152 7.3702
R287 VTAIL.n119 VTAIL.n80 7.3702
R288 VTAIL.n115 VTAIL.n82 7.3702
R289 VTAIL.n256 VTAIL.n255 6.59444
R290 VTAIL.n256 VTAIL.n220 6.59444
R291 VTAIL.n46 VTAIL.n45 6.59444
R292 VTAIL.n46 VTAIL.n10 6.59444
R293 VTAIL.n186 VTAIL.n150 6.59444
R294 VTAIL.n186 VTAIL.n185 6.59444
R295 VTAIL.n116 VTAIL.n80 6.59444
R296 VTAIL.n116 VTAIL.n115 6.59444
R297 VTAIL.n252 VTAIL.n222 5.81868
R298 VTAIL.n260 VTAIL.n259 5.81868
R299 VTAIL.n42 VTAIL.n12 5.81868
R300 VTAIL.n50 VTAIL.n49 5.81868
R301 VTAIL.n190 VTAIL.n189 5.81868
R302 VTAIL.n182 VTAIL.n152 5.81868
R303 VTAIL.n120 VTAIL.n119 5.81868
R304 VTAIL.n112 VTAIL.n82 5.81868
R305 VTAIL.n251 VTAIL.n224 5.04292
R306 VTAIL.n263 VTAIL.n218 5.04292
R307 VTAIL.n41 VTAIL.n14 5.04292
R308 VTAIL.n53 VTAIL.n8 5.04292
R309 VTAIL.n193 VTAIL.n148 5.04292
R310 VTAIL.n181 VTAIL.n154 5.04292
R311 VTAIL.n123 VTAIL.n78 5.04292
R312 VTAIL.n111 VTAIL.n84 5.04292
R313 VTAIL.n234 VTAIL.n233 4.38563
R314 VTAIL.n24 VTAIL.n23 4.38563
R315 VTAIL.n164 VTAIL.n163 4.38563
R316 VTAIL.n94 VTAIL.n93 4.38563
R317 VTAIL.n248 VTAIL.n247 4.26717
R318 VTAIL.n264 VTAIL.n216 4.26717
R319 VTAIL.n38 VTAIL.n37 4.26717
R320 VTAIL.n54 VTAIL.n6 4.26717
R321 VTAIL.n194 VTAIL.n146 4.26717
R322 VTAIL.n178 VTAIL.n177 4.26717
R323 VTAIL.n124 VTAIL.n76 4.26717
R324 VTAIL.n108 VTAIL.n107 4.26717
R325 VTAIL.n244 VTAIL.n226 3.49141
R326 VTAIL.n268 VTAIL.n267 3.49141
R327 VTAIL.n34 VTAIL.n16 3.49141
R328 VTAIL.n58 VTAIL.n57 3.49141
R329 VTAIL.n198 VTAIL.n197 3.49141
R330 VTAIL.n174 VTAIL.n156 3.49141
R331 VTAIL.n128 VTAIL.n127 3.49141
R332 VTAIL.n104 VTAIL.n86 3.49141
R333 VTAIL.n243 VTAIL.n228 2.71565
R334 VTAIL.n271 VTAIL.n214 2.71565
R335 VTAIL.n33 VTAIL.n18 2.71565
R336 VTAIL.n61 VTAIL.n4 2.71565
R337 VTAIL.n201 VTAIL.n144 2.71565
R338 VTAIL.n173 VTAIL.n158 2.71565
R339 VTAIL.n131 VTAIL.n74 2.71565
R340 VTAIL.n103 VTAIL.n88 2.71565
R341 VTAIL.n240 VTAIL.n239 1.93989
R342 VTAIL.n272 VTAIL.n212 1.93989
R343 VTAIL.n30 VTAIL.n29 1.93989
R344 VTAIL.n62 VTAIL.n2 1.93989
R345 VTAIL.n202 VTAIL.n142 1.93989
R346 VTAIL.n170 VTAIL.n169 1.93989
R347 VTAIL.n132 VTAIL.n72 1.93989
R348 VTAIL.n100 VTAIL.n99 1.93989
R349 VTAIL.n236 VTAIL.n230 1.16414
R350 VTAIL.n276 VTAIL.n275 1.16414
R351 VTAIL.n26 VTAIL.n20 1.16414
R352 VTAIL.n66 VTAIL.n65 1.16414
R353 VTAIL.n206 VTAIL.n205 1.16414
R354 VTAIL.n166 VTAIL.n160 1.16414
R355 VTAIL.n136 VTAIL.n135 1.16414
R356 VTAIL.n96 VTAIL.n90 1.16414
R357 VTAIL.n209 VTAIL.n139 0.931535
R358 VTAIL VTAIL.n69 0.759121
R359 VTAIL.n235 VTAIL.n232 0.388379
R360 VTAIL.n278 VTAIL.n210 0.388379
R361 VTAIL.n25 VTAIL.n22 0.388379
R362 VTAIL.n68 VTAIL.n0 0.388379
R363 VTAIL.n208 VTAIL.n140 0.388379
R364 VTAIL.n165 VTAIL.n162 0.388379
R365 VTAIL.n138 VTAIL.n70 0.388379
R366 VTAIL.n95 VTAIL.n92 0.388379
R367 VTAIL VTAIL.n279 0.172914
R368 VTAIL.n234 VTAIL.n229 0.155672
R369 VTAIL.n241 VTAIL.n229 0.155672
R370 VTAIL.n242 VTAIL.n241 0.155672
R371 VTAIL.n242 VTAIL.n225 0.155672
R372 VTAIL.n249 VTAIL.n225 0.155672
R373 VTAIL.n250 VTAIL.n249 0.155672
R374 VTAIL.n250 VTAIL.n221 0.155672
R375 VTAIL.n257 VTAIL.n221 0.155672
R376 VTAIL.n258 VTAIL.n257 0.155672
R377 VTAIL.n258 VTAIL.n217 0.155672
R378 VTAIL.n265 VTAIL.n217 0.155672
R379 VTAIL.n266 VTAIL.n265 0.155672
R380 VTAIL.n266 VTAIL.n213 0.155672
R381 VTAIL.n273 VTAIL.n213 0.155672
R382 VTAIL.n274 VTAIL.n273 0.155672
R383 VTAIL.n24 VTAIL.n19 0.155672
R384 VTAIL.n31 VTAIL.n19 0.155672
R385 VTAIL.n32 VTAIL.n31 0.155672
R386 VTAIL.n32 VTAIL.n15 0.155672
R387 VTAIL.n39 VTAIL.n15 0.155672
R388 VTAIL.n40 VTAIL.n39 0.155672
R389 VTAIL.n40 VTAIL.n11 0.155672
R390 VTAIL.n47 VTAIL.n11 0.155672
R391 VTAIL.n48 VTAIL.n47 0.155672
R392 VTAIL.n48 VTAIL.n7 0.155672
R393 VTAIL.n55 VTAIL.n7 0.155672
R394 VTAIL.n56 VTAIL.n55 0.155672
R395 VTAIL.n56 VTAIL.n3 0.155672
R396 VTAIL.n63 VTAIL.n3 0.155672
R397 VTAIL.n64 VTAIL.n63 0.155672
R398 VTAIL.n204 VTAIL.n203 0.155672
R399 VTAIL.n203 VTAIL.n143 0.155672
R400 VTAIL.n196 VTAIL.n143 0.155672
R401 VTAIL.n196 VTAIL.n195 0.155672
R402 VTAIL.n195 VTAIL.n147 0.155672
R403 VTAIL.n188 VTAIL.n147 0.155672
R404 VTAIL.n188 VTAIL.n187 0.155672
R405 VTAIL.n187 VTAIL.n151 0.155672
R406 VTAIL.n180 VTAIL.n151 0.155672
R407 VTAIL.n180 VTAIL.n179 0.155672
R408 VTAIL.n179 VTAIL.n155 0.155672
R409 VTAIL.n172 VTAIL.n155 0.155672
R410 VTAIL.n172 VTAIL.n171 0.155672
R411 VTAIL.n171 VTAIL.n159 0.155672
R412 VTAIL.n164 VTAIL.n159 0.155672
R413 VTAIL.n134 VTAIL.n133 0.155672
R414 VTAIL.n133 VTAIL.n73 0.155672
R415 VTAIL.n126 VTAIL.n73 0.155672
R416 VTAIL.n126 VTAIL.n125 0.155672
R417 VTAIL.n125 VTAIL.n77 0.155672
R418 VTAIL.n118 VTAIL.n77 0.155672
R419 VTAIL.n118 VTAIL.n117 0.155672
R420 VTAIL.n117 VTAIL.n81 0.155672
R421 VTAIL.n110 VTAIL.n81 0.155672
R422 VTAIL.n110 VTAIL.n109 0.155672
R423 VTAIL.n109 VTAIL.n85 0.155672
R424 VTAIL.n102 VTAIL.n85 0.155672
R425 VTAIL.n102 VTAIL.n101 0.155672
R426 VTAIL.n101 VTAIL.n89 0.155672
R427 VTAIL.n94 VTAIL.n89 0.155672
R428 VDD1.n68 VDD1.n67 289.615
R429 VDD1.n137 VDD1.n136 289.615
R430 VDD1.n67 VDD1.n66 185
R431 VDD1.n2 VDD1.n1 185
R432 VDD1.n61 VDD1.n60 185
R433 VDD1.n59 VDD1.n58 185
R434 VDD1.n6 VDD1.n5 185
R435 VDD1.n53 VDD1.n52 185
R436 VDD1.n51 VDD1.n50 185
R437 VDD1.n10 VDD1.n9 185
R438 VDD1.n45 VDD1.n44 185
R439 VDD1.n43 VDD1.n42 185
R440 VDD1.n14 VDD1.n13 185
R441 VDD1.n37 VDD1.n36 185
R442 VDD1.n35 VDD1.n34 185
R443 VDD1.n18 VDD1.n17 185
R444 VDD1.n29 VDD1.n28 185
R445 VDD1.n27 VDD1.n26 185
R446 VDD1.n22 VDD1.n21 185
R447 VDD1.n91 VDD1.n90 185
R448 VDD1.n96 VDD1.n95 185
R449 VDD1.n98 VDD1.n97 185
R450 VDD1.n87 VDD1.n86 185
R451 VDD1.n104 VDD1.n103 185
R452 VDD1.n106 VDD1.n105 185
R453 VDD1.n83 VDD1.n82 185
R454 VDD1.n112 VDD1.n111 185
R455 VDD1.n114 VDD1.n113 185
R456 VDD1.n79 VDD1.n78 185
R457 VDD1.n120 VDD1.n119 185
R458 VDD1.n122 VDD1.n121 185
R459 VDD1.n75 VDD1.n74 185
R460 VDD1.n128 VDD1.n127 185
R461 VDD1.n130 VDD1.n129 185
R462 VDD1.n71 VDD1.n70 185
R463 VDD1.n136 VDD1.n135 185
R464 VDD1.n92 VDD1.t0 147.659
R465 VDD1.n23 VDD1.t1 147.659
R466 VDD1.n67 VDD1.n1 104.615
R467 VDD1.n60 VDD1.n1 104.615
R468 VDD1.n60 VDD1.n59 104.615
R469 VDD1.n59 VDD1.n5 104.615
R470 VDD1.n52 VDD1.n5 104.615
R471 VDD1.n52 VDD1.n51 104.615
R472 VDD1.n51 VDD1.n9 104.615
R473 VDD1.n44 VDD1.n9 104.615
R474 VDD1.n44 VDD1.n43 104.615
R475 VDD1.n43 VDD1.n13 104.615
R476 VDD1.n36 VDD1.n13 104.615
R477 VDD1.n36 VDD1.n35 104.615
R478 VDD1.n35 VDD1.n17 104.615
R479 VDD1.n28 VDD1.n17 104.615
R480 VDD1.n28 VDD1.n27 104.615
R481 VDD1.n27 VDD1.n21 104.615
R482 VDD1.n96 VDD1.n90 104.615
R483 VDD1.n97 VDD1.n96 104.615
R484 VDD1.n97 VDD1.n86 104.615
R485 VDD1.n104 VDD1.n86 104.615
R486 VDD1.n105 VDD1.n104 104.615
R487 VDD1.n105 VDD1.n82 104.615
R488 VDD1.n112 VDD1.n82 104.615
R489 VDD1.n113 VDD1.n112 104.615
R490 VDD1.n113 VDD1.n78 104.615
R491 VDD1.n120 VDD1.n78 104.615
R492 VDD1.n121 VDD1.n120 104.615
R493 VDD1.n121 VDD1.n74 104.615
R494 VDD1.n128 VDD1.n74 104.615
R495 VDD1.n129 VDD1.n128 104.615
R496 VDD1.n129 VDD1.n70 104.615
R497 VDD1.n136 VDD1.n70 104.615
R498 VDD1 VDD1.n137 89.7656
R499 VDD1 VDD1.n68 52.8378
R500 VDD1.t1 VDD1.n21 52.3082
R501 VDD1.t0 VDD1.n90 52.3082
R502 VDD1.n23 VDD1.n22 15.6677
R503 VDD1.n92 VDD1.n91 15.6677
R504 VDD1.n66 VDD1.n0 12.8005
R505 VDD1.n26 VDD1.n25 12.8005
R506 VDD1.n95 VDD1.n94 12.8005
R507 VDD1.n135 VDD1.n69 12.8005
R508 VDD1.n65 VDD1.n2 12.0247
R509 VDD1.n29 VDD1.n20 12.0247
R510 VDD1.n98 VDD1.n89 12.0247
R511 VDD1.n134 VDD1.n71 12.0247
R512 VDD1.n62 VDD1.n61 11.249
R513 VDD1.n30 VDD1.n18 11.249
R514 VDD1.n99 VDD1.n87 11.249
R515 VDD1.n131 VDD1.n130 11.249
R516 VDD1.n58 VDD1.n4 10.4732
R517 VDD1.n34 VDD1.n33 10.4732
R518 VDD1.n103 VDD1.n102 10.4732
R519 VDD1.n127 VDD1.n73 10.4732
R520 VDD1.n57 VDD1.n6 9.69747
R521 VDD1.n37 VDD1.n16 9.69747
R522 VDD1.n106 VDD1.n85 9.69747
R523 VDD1.n126 VDD1.n75 9.69747
R524 VDD1.n64 VDD1.n0 9.45567
R525 VDD1.n133 VDD1.n69 9.45567
R526 VDD1.n65 VDD1.n64 9.3005
R527 VDD1.n63 VDD1.n62 9.3005
R528 VDD1.n4 VDD1.n3 9.3005
R529 VDD1.n57 VDD1.n56 9.3005
R530 VDD1.n55 VDD1.n54 9.3005
R531 VDD1.n8 VDD1.n7 9.3005
R532 VDD1.n49 VDD1.n48 9.3005
R533 VDD1.n47 VDD1.n46 9.3005
R534 VDD1.n12 VDD1.n11 9.3005
R535 VDD1.n41 VDD1.n40 9.3005
R536 VDD1.n39 VDD1.n38 9.3005
R537 VDD1.n16 VDD1.n15 9.3005
R538 VDD1.n33 VDD1.n32 9.3005
R539 VDD1.n31 VDD1.n30 9.3005
R540 VDD1.n20 VDD1.n19 9.3005
R541 VDD1.n25 VDD1.n24 9.3005
R542 VDD1.n116 VDD1.n115 9.3005
R543 VDD1.n118 VDD1.n117 9.3005
R544 VDD1.n77 VDD1.n76 9.3005
R545 VDD1.n124 VDD1.n123 9.3005
R546 VDD1.n126 VDD1.n125 9.3005
R547 VDD1.n73 VDD1.n72 9.3005
R548 VDD1.n132 VDD1.n131 9.3005
R549 VDD1.n134 VDD1.n133 9.3005
R550 VDD1.n110 VDD1.n109 9.3005
R551 VDD1.n108 VDD1.n107 9.3005
R552 VDD1.n85 VDD1.n84 9.3005
R553 VDD1.n102 VDD1.n101 9.3005
R554 VDD1.n100 VDD1.n99 9.3005
R555 VDD1.n89 VDD1.n88 9.3005
R556 VDD1.n94 VDD1.n93 9.3005
R557 VDD1.n81 VDD1.n80 9.3005
R558 VDD1.n54 VDD1.n53 8.92171
R559 VDD1.n38 VDD1.n14 8.92171
R560 VDD1.n107 VDD1.n83 8.92171
R561 VDD1.n123 VDD1.n122 8.92171
R562 VDD1.n50 VDD1.n8 8.14595
R563 VDD1.n42 VDD1.n41 8.14595
R564 VDD1.n111 VDD1.n110 8.14595
R565 VDD1.n119 VDD1.n77 8.14595
R566 VDD1.n49 VDD1.n10 7.3702
R567 VDD1.n45 VDD1.n12 7.3702
R568 VDD1.n114 VDD1.n81 7.3702
R569 VDD1.n118 VDD1.n79 7.3702
R570 VDD1.n46 VDD1.n10 6.59444
R571 VDD1.n46 VDD1.n45 6.59444
R572 VDD1.n115 VDD1.n114 6.59444
R573 VDD1.n115 VDD1.n79 6.59444
R574 VDD1.n50 VDD1.n49 5.81868
R575 VDD1.n42 VDD1.n12 5.81868
R576 VDD1.n111 VDD1.n81 5.81868
R577 VDD1.n119 VDD1.n118 5.81868
R578 VDD1.n53 VDD1.n8 5.04292
R579 VDD1.n41 VDD1.n14 5.04292
R580 VDD1.n110 VDD1.n83 5.04292
R581 VDD1.n122 VDD1.n77 5.04292
R582 VDD1.n93 VDD1.n92 4.38563
R583 VDD1.n24 VDD1.n23 4.38563
R584 VDD1.n54 VDD1.n6 4.26717
R585 VDD1.n38 VDD1.n37 4.26717
R586 VDD1.n107 VDD1.n106 4.26717
R587 VDD1.n123 VDD1.n75 4.26717
R588 VDD1.n58 VDD1.n57 3.49141
R589 VDD1.n34 VDD1.n16 3.49141
R590 VDD1.n103 VDD1.n85 3.49141
R591 VDD1.n127 VDD1.n126 3.49141
R592 VDD1.n61 VDD1.n4 2.71565
R593 VDD1.n33 VDD1.n18 2.71565
R594 VDD1.n102 VDD1.n87 2.71565
R595 VDD1.n130 VDD1.n73 2.71565
R596 VDD1.n62 VDD1.n2 1.93989
R597 VDD1.n30 VDD1.n29 1.93989
R598 VDD1.n99 VDD1.n98 1.93989
R599 VDD1.n131 VDD1.n71 1.93989
R600 VDD1.n66 VDD1.n65 1.16414
R601 VDD1.n26 VDD1.n20 1.16414
R602 VDD1.n95 VDD1.n89 1.16414
R603 VDD1.n135 VDD1.n134 1.16414
R604 VDD1.n68 VDD1.n0 0.388379
R605 VDD1.n25 VDD1.n22 0.388379
R606 VDD1.n94 VDD1.n91 0.388379
R607 VDD1.n137 VDD1.n69 0.388379
R608 VDD1.n64 VDD1.n63 0.155672
R609 VDD1.n63 VDD1.n3 0.155672
R610 VDD1.n56 VDD1.n3 0.155672
R611 VDD1.n56 VDD1.n55 0.155672
R612 VDD1.n55 VDD1.n7 0.155672
R613 VDD1.n48 VDD1.n7 0.155672
R614 VDD1.n48 VDD1.n47 0.155672
R615 VDD1.n47 VDD1.n11 0.155672
R616 VDD1.n40 VDD1.n11 0.155672
R617 VDD1.n40 VDD1.n39 0.155672
R618 VDD1.n39 VDD1.n15 0.155672
R619 VDD1.n32 VDD1.n15 0.155672
R620 VDD1.n32 VDD1.n31 0.155672
R621 VDD1.n31 VDD1.n19 0.155672
R622 VDD1.n24 VDD1.n19 0.155672
R623 VDD1.n93 VDD1.n88 0.155672
R624 VDD1.n100 VDD1.n88 0.155672
R625 VDD1.n101 VDD1.n100 0.155672
R626 VDD1.n101 VDD1.n84 0.155672
R627 VDD1.n108 VDD1.n84 0.155672
R628 VDD1.n109 VDD1.n108 0.155672
R629 VDD1.n109 VDD1.n80 0.155672
R630 VDD1.n116 VDD1.n80 0.155672
R631 VDD1.n117 VDD1.n116 0.155672
R632 VDD1.n117 VDD1.n76 0.155672
R633 VDD1.n124 VDD1.n76 0.155672
R634 VDD1.n125 VDD1.n124 0.155672
R635 VDD1.n125 VDD1.n72 0.155672
R636 VDD1.n132 VDD1.n72 0.155672
R637 VDD1.n133 VDD1.n132 0.155672
R638 B.n54 B.t6 615.783
R639 B.n60 B.t2 615.783
R640 B.n139 B.t13 615.783
R641 B.n133 B.t9 615.783
R642 B.n420 B.n83 585
R643 B.n83 B.n30 585
R644 B.n422 B.n421 585
R645 B.n424 B.n82 585
R646 B.n427 B.n426 585
R647 B.n428 B.n81 585
R648 B.n430 B.n429 585
R649 B.n432 B.n80 585
R650 B.n435 B.n434 585
R651 B.n436 B.n79 585
R652 B.n438 B.n437 585
R653 B.n440 B.n78 585
R654 B.n443 B.n442 585
R655 B.n444 B.n77 585
R656 B.n446 B.n445 585
R657 B.n448 B.n76 585
R658 B.n451 B.n450 585
R659 B.n452 B.n75 585
R660 B.n454 B.n453 585
R661 B.n456 B.n74 585
R662 B.n459 B.n458 585
R663 B.n460 B.n73 585
R664 B.n462 B.n461 585
R665 B.n464 B.n72 585
R666 B.n467 B.n466 585
R667 B.n468 B.n71 585
R668 B.n470 B.n469 585
R669 B.n472 B.n70 585
R670 B.n475 B.n474 585
R671 B.n476 B.n69 585
R672 B.n478 B.n477 585
R673 B.n480 B.n68 585
R674 B.n483 B.n482 585
R675 B.n484 B.n67 585
R676 B.n486 B.n485 585
R677 B.n488 B.n66 585
R678 B.n491 B.n490 585
R679 B.n492 B.n65 585
R680 B.n494 B.n493 585
R681 B.n496 B.n64 585
R682 B.n499 B.n498 585
R683 B.n500 B.n63 585
R684 B.n502 B.n501 585
R685 B.n504 B.n62 585
R686 B.n507 B.n506 585
R687 B.n509 B.n59 585
R688 B.n511 B.n510 585
R689 B.n513 B.n58 585
R690 B.n516 B.n515 585
R691 B.n517 B.n57 585
R692 B.n519 B.n518 585
R693 B.n521 B.n56 585
R694 B.n524 B.n523 585
R695 B.n525 B.n53 585
R696 B.n528 B.n527 585
R697 B.n530 B.n52 585
R698 B.n533 B.n532 585
R699 B.n534 B.n51 585
R700 B.n536 B.n535 585
R701 B.n538 B.n50 585
R702 B.n541 B.n540 585
R703 B.n542 B.n49 585
R704 B.n544 B.n543 585
R705 B.n546 B.n48 585
R706 B.n549 B.n548 585
R707 B.n550 B.n47 585
R708 B.n552 B.n551 585
R709 B.n554 B.n46 585
R710 B.n557 B.n556 585
R711 B.n558 B.n45 585
R712 B.n560 B.n559 585
R713 B.n562 B.n44 585
R714 B.n565 B.n564 585
R715 B.n566 B.n43 585
R716 B.n568 B.n567 585
R717 B.n570 B.n42 585
R718 B.n573 B.n572 585
R719 B.n574 B.n41 585
R720 B.n576 B.n575 585
R721 B.n578 B.n40 585
R722 B.n581 B.n580 585
R723 B.n582 B.n39 585
R724 B.n584 B.n583 585
R725 B.n586 B.n38 585
R726 B.n589 B.n588 585
R727 B.n590 B.n37 585
R728 B.n592 B.n591 585
R729 B.n594 B.n36 585
R730 B.n597 B.n596 585
R731 B.n598 B.n35 585
R732 B.n600 B.n599 585
R733 B.n602 B.n34 585
R734 B.n605 B.n604 585
R735 B.n606 B.n33 585
R736 B.n608 B.n607 585
R737 B.n610 B.n32 585
R738 B.n613 B.n612 585
R739 B.n614 B.n31 585
R740 B.n419 B.n29 585
R741 B.n617 B.n29 585
R742 B.n418 B.n28 585
R743 B.n618 B.n28 585
R744 B.n417 B.n27 585
R745 B.n619 B.n27 585
R746 B.n416 B.n415 585
R747 B.n415 B.n23 585
R748 B.n414 B.n22 585
R749 B.n625 B.n22 585
R750 B.n413 B.n21 585
R751 B.n626 B.n21 585
R752 B.n412 B.n20 585
R753 B.n627 B.n20 585
R754 B.n411 B.n410 585
R755 B.n410 B.n16 585
R756 B.n409 B.n15 585
R757 B.n633 B.n15 585
R758 B.n408 B.n14 585
R759 B.n634 B.n14 585
R760 B.n407 B.n13 585
R761 B.n635 B.n13 585
R762 B.n406 B.n405 585
R763 B.n405 B.n12 585
R764 B.n404 B.n403 585
R765 B.n404 B.n8 585
R766 B.n402 B.n7 585
R767 B.n642 B.n7 585
R768 B.n401 B.n6 585
R769 B.n643 B.n6 585
R770 B.n400 B.n5 585
R771 B.n644 B.n5 585
R772 B.n399 B.n398 585
R773 B.n398 B.n4 585
R774 B.n397 B.n84 585
R775 B.n397 B.n396 585
R776 B.n386 B.n85 585
R777 B.n389 B.n85 585
R778 B.n388 B.n387 585
R779 B.n390 B.n388 585
R780 B.n385 B.n90 585
R781 B.n90 B.n89 585
R782 B.n384 B.n383 585
R783 B.n383 B.n382 585
R784 B.n92 B.n91 585
R785 B.n93 B.n92 585
R786 B.n375 B.n374 585
R787 B.n376 B.n375 585
R788 B.n373 B.n98 585
R789 B.n98 B.n97 585
R790 B.n372 B.n371 585
R791 B.n371 B.n370 585
R792 B.n100 B.n99 585
R793 B.n101 B.n100 585
R794 B.n363 B.n362 585
R795 B.n364 B.n363 585
R796 B.n361 B.n106 585
R797 B.n106 B.n105 585
R798 B.n360 B.n359 585
R799 B.n359 B.n358 585
R800 B.n355 B.n110 585
R801 B.n354 B.n353 585
R802 B.n351 B.n111 585
R803 B.n351 B.n109 585
R804 B.n350 B.n349 585
R805 B.n348 B.n347 585
R806 B.n346 B.n113 585
R807 B.n344 B.n343 585
R808 B.n342 B.n114 585
R809 B.n341 B.n340 585
R810 B.n338 B.n115 585
R811 B.n336 B.n335 585
R812 B.n334 B.n116 585
R813 B.n333 B.n332 585
R814 B.n330 B.n117 585
R815 B.n328 B.n327 585
R816 B.n326 B.n118 585
R817 B.n325 B.n324 585
R818 B.n322 B.n119 585
R819 B.n320 B.n319 585
R820 B.n318 B.n120 585
R821 B.n317 B.n316 585
R822 B.n314 B.n121 585
R823 B.n312 B.n311 585
R824 B.n310 B.n122 585
R825 B.n309 B.n308 585
R826 B.n306 B.n123 585
R827 B.n304 B.n303 585
R828 B.n302 B.n124 585
R829 B.n301 B.n300 585
R830 B.n298 B.n125 585
R831 B.n296 B.n295 585
R832 B.n294 B.n126 585
R833 B.n293 B.n292 585
R834 B.n290 B.n127 585
R835 B.n288 B.n287 585
R836 B.n286 B.n128 585
R837 B.n285 B.n284 585
R838 B.n282 B.n129 585
R839 B.n280 B.n279 585
R840 B.n278 B.n130 585
R841 B.n277 B.n276 585
R842 B.n274 B.n131 585
R843 B.n272 B.n271 585
R844 B.n270 B.n132 585
R845 B.n268 B.n267 585
R846 B.n265 B.n135 585
R847 B.n263 B.n262 585
R848 B.n261 B.n136 585
R849 B.n260 B.n259 585
R850 B.n257 B.n137 585
R851 B.n255 B.n254 585
R852 B.n253 B.n138 585
R853 B.n252 B.n251 585
R854 B.n249 B.n248 585
R855 B.n247 B.n246 585
R856 B.n245 B.n143 585
R857 B.n243 B.n242 585
R858 B.n241 B.n144 585
R859 B.n240 B.n239 585
R860 B.n237 B.n145 585
R861 B.n235 B.n234 585
R862 B.n233 B.n146 585
R863 B.n232 B.n231 585
R864 B.n229 B.n147 585
R865 B.n227 B.n226 585
R866 B.n225 B.n148 585
R867 B.n224 B.n223 585
R868 B.n221 B.n149 585
R869 B.n219 B.n218 585
R870 B.n217 B.n150 585
R871 B.n216 B.n215 585
R872 B.n213 B.n151 585
R873 B.n211 B.n210 585
R874 B.n209 B.n152 585
R875 B.n208 B.n207 585
R876 B.n205 B.n153 585
R877 B.n203 B.n202 585
R878 B.n201 B.n154 585
R879 B.n200 B.n199 585
R880 B.n197 B.n155 585
R881 B.n195 B.n194 585
R882 B.n193 B.n156 585
R883 B.n192 B.n191 585
R884 B.n189 B.n157 585
R885 B.n187 B.n186 585
R886 B.n185 B.n158 585
R887 B.n184 B.n183 585
R888 B.n181 B.n159 585
R889 B.n179 B.n178 585
R890 B.n177 B.n160 585
R891 B.n176 B.n175 585
R892 B.n173 B.n161 585
R893 B.n171 B.n170 585
R894 B.n169 B.n162 585
R895 B.n168 B.n167 585
R896 B.n165 B.n163 585
R897 B.n108 B.n107 585
R898 B.n357 B.n356 585
R899 B.n358 B.n357 585
R900 B.n104 B.n103 585
R901 B.n105 B.n104 585
R902 B.n366 B.n365 585
R903 B.n365 B.n364 585
R904 B.n367 B.n102 585
R905 B.n102 B.n101 585
R906 B.n369 B.n368 585
R907 B.n370 B.n369 585
R908 B.n96 B.n95 585
R909 B.n97 B.n96 585
R910 B.n378 B.n377 585
R911 B.n377 B.n376 585
R912 B.n379 B.n94 585
R913 B.n94 B.n93 585
R914 B.n381 B.n380 585
R915 B.n382 B.n381 585
R916 B.n88 B.n87 585
R917 B.n89 B.n88 585
R918 B.n392 B.n391 585
R919 B.n391 B.n390 585
R920 B.n393 B.n86 585
R921 B.n389 B.n86 585
R922 B.n395 B.n394 585
R923 B.n396 B.n395 585
R924 B.n3 B.n0 585
R925 B.n4 B.n3 585
R926 B.n641 B.n1 585
R927 B.n642 B.n641 585
R928 B.n640 B.n639 585
R929 B.n640 B.n8 585
R930 B.n638 B.n9 585
R931 B.n12 B.n9 585
R932 B.n637 B.n636 585
R933 B.n636 B.n635 585
R934 B.n11 B.n10 585
R935 B.n634 B.n11 585
R936 B.n632 B.n631 585
R937 B.n633 B.n632 585
R938 B.n630 B.n17 585
R939 B.n17 B.n16 585
R940 B.n629 B.n628 585
R941 B.n628 B.n627 585
R942 B.n19 B.n18 585
R943 B.n626 B.n19 585
R944 B.n624 B.n623 585
R945 B.n625 B.n624 585
R946 B.n622 B.n24 585
R947 B.n24 B.n23 585
R948 B.n621 B.n620 585
R949 B.n620 B.n619 585
R950 B.n26 B.n25 585
R951 B.n618 B.n26 585
R952 B.n616 B.n615 585
R953 B.n617 B.n616 585
R954 B.n645 B.n644 585
R955 B.n643 B.n2 585
R956 B.n616 B.n31 482.89
R957 B.n83 B.n29 482.89
R958 B.n359 B.n108 482.89
R959 B.n357 B.n110 482.89
R960 B.n60 B.t4 314.666
R961 B.n139 B.t15 314.666
R962 B.n54 B.t7 314.666
R963 B.n133 B.t12 314.666
R964 B.n61 B.t5 293.914
R965 B.n140 B.t14 293.914
R966 B.n55 B.t8 293.914
R967 B.n134 B.t11 293.914
R968 B.n423 B.n30 256.663
R969 B.n425 B.n30 256.663
R970 B.n431 B.n30 256.663
R971 B.n433 B.n30 256.663
R972 B.n439 B.n30 256.663
R973 B.n441 B.n30 256.663
R974 B.n447 B.n30 256.663
R975 B.n449 B.n30 256.663
R976 B.n455 B.n30 256.663
R977 B.n457 B.n30 256.663
R978 B.n463 B.n30 256.663
R979 B.n465 B.n30 256.663
R980 B.n471 B.n30 256.663
R981 B.n473 B.n30 256.663
R982 B.n479 B.n30 256.663
R983 B.n481 B.n30 256.663
R984 B.n487 B.n30 256.663
R985 B.n489 B.n30 256.663
R986 B.n495 B.n30 256.663
R987 B.n497 B.n30 256.663
R988 B.n503 B.n30 256.663
R989 B.n505 B.n30 256.663
R990 B.n512 B.n30 256.663
R991 B.n514 B.n30 256.663
R992 B.n520 B.n30 256.663
R993 B.n522 B.n30 256.663
R994 B.n529 B.n30 256.663
R995 B.n531 B.n30 256.663
R996 B.n537 B.n30 256.663
R997 B.n539 B.n30 256.663
R998 B.n545 B.n30 256.663
R999 B.n547 B.n30 256.663
R1000 B.n553 B.n30 256.663
R1001 B.n555 B.n30 256.663
R1002 B.n561 B.n30 256.663
R1003 B.n563 B.n30 256.663
R1004 B.n569 B.n30 256.663
R1005 B.n571 B.n30 256.663
R1006 B.n577 B.n30 256.663
R1007 B.n579 B.n30 256.663
R1008 B.n585 B.n30 256.663
R1009 B.n587 B.n30 256.663
R1010 B.n593 B.n30 256.663
R1011 B.n595 B.n30 256.663
R1012 B.n601 B.n30 256.663
R1013 B.n603 B.n30 256.663
R1014 B.n609 B.n30 256.663
R1015 B.n611 B.n30 256.663
R1016 B.n352 B.n109 256.663
R1017 B.n112 B.n109 256.663
R1018 B.n345 B.n109 256.663
R1019 B.n339 B.n109 256.663
R1020 B.n337 B.n109 256.663
R1021 B.n331 B.n109 256.663
R1022 B.n329 B.n109 256.663
R1023 B.n323 B.n109 256.663
R1024 B.n321 B.n109 256.663
R1025 B.n315 B.n109 256.663
R1026 B.n313 B.n109 256.663
R1027 B.n307 B.n109 256.663
R1028 B.n305 B.n109 256.663
R1029 B.n299 B.n109 256.663
R1030 B.n297 B.n109 256.663
R1031 B.n291 B.n109 256.663
R1032 B.n289 B.n109 256.663
R1033 B.n283 B.n109 256.663
R1034 B.n281 B.n109 256.663
R1035 B.n275 B.n109 256.663
R1036 B.n273 B.n109 256.663
R1037 B.n266 B.n109 256.663
R1038 B.n264 B.n109 256.663
R1039 B.n258 B.n109 256.663
R1040 B.n256 B.n109 256.663
R1041 B.n250 B.n109 256.663
R1042 B.n142 B.n109 256.663
R1043 B.n244 B.n109 256.663
R1044 B.n238 B.n109 256.663
R1045 B.n236 B.n109 256.663
R1046 B.n230 B.n109 256.663
R1047 B.n228 B.n109 256.663
R1048 B.n222 B.n109 256.663
R1049 B.n220 B.n109 256.663
R1050 B.n214 B.n109 256.663
R1051 B.n212 B.n109 256.663
R1052 B.n206 B.n109 256.663
R1053 B.n204 B.n109 256.663
R1054 B.n198 B.n109 256.663
R1055 B.n196 B.n109 256.663
R1056 B.n190 B.n109 256.663
R1057 B.n188 B.n109 256.663
R1058 B.n182 B.n109 256.663
R1059 B.n180 B.n109 256.663
R1060 B.n174 B.n109 256.663
R1061 B.n172 B.n109 256.663
R1062 B.n166 B.n109 256.663
R1063 B.n164 B.n109 256.663
R1064 B.n647 B.n646 256.663
R1065 B.n612 B.n610 163.367
R1066 B.n608 B.n33 163.367
R1067 B.n604 B.n602 163.367
R1068 B.n600 B.n35 163.367
R1069 B.n596 B.n594 163.367
R1070 B.n592 B.n37 163.367
R1071 B.n588 B.n586 163.367
R1072 B.n584 B.n39 163.367
R1073 B.n580 B.n578 163.367
R1074 B.n576 B.n41 163.367
R1075 B.n572 B.n570 163.367
R1076 B.n568 B.n43 163.367
R1077 B.n564 B.n562 163.367
R1078 B.n560 B.n45 163.367
R1079 B.n556 B.n554 163.367
R1080 B.n552 B.n47 163.367
R1081 B.n548 B.n546 163.367
R1082 B.n544 B.n49 163.367
R1083 B.n540 B.n538 163.367
R1084 B.n536 B.n51 163.367
R1085 B.n532 B.n530 163.367
R1086 B.n528 B.n53 163.367
R1087 B.n523 B.n521 163.367
R1088 B.n519 B.n57 163.367
R1089 B.n515 B.n513 163.367
R1090 B.n511 B.n59 163.367
R1091 B.n506 B.n504 163.367
R1092 B.n502 B.n63 163.367
R1093 B.n498 B.n496 163.367
R1094 B.n494 B.n65 163.367
R1095 B.n490 B.n488 163.367
R1096 B.n486 B.n67 163.367
R1097 B.n482 B.n480 163.367
R1098 B.n478 B.n69 163.367
R1099 B.n474 B.n472 163.367
R1100 B.n470 B.n71 163.367
R1101 B.n466 B.n464 163.367
R1102 B.n462 B.n73 163.367
R1103 B.n458 B.n456 163.367
R1104 B.n454 B.n75 163.367
R1105 B.n450 B.n448 163.367
R1106 B.n446 B.n77 163.367
R1107 B.n442 B.n440 163.367
R1108 B.n438 B.n79 163.367
R1109 B.n434 B.n432 163.367
R1110 B.n430 B.n81 163.367
R1111 B.n426 B.n424 163.367
R1112 B.n422 B.n83 163.367
R1113 B.n359 B.n106 163.367
R1114 B.n363 B.n106 163.367
R1115 B.n363 B.n100 163.367
R1116 B.n371 B.n100 163.367
R1117 B.n371 B.n98 163.367
R1118 B.n375 B.n98 163.367
R1119 B.n375 B.n92 163.367
R1120 B.n383 B.n92 163.367
R1121 B.n383 B.n90 163.367
R1122 B.n388 B.n90 163.367
R1123 B.n388 B.n85 163.367
R1124 B.n397 B.n85 163.367
R1125 B.n398 B.n397 163.367
R1126 B.n398 B.n5 163.367
R1127 B.n6 B.n5 163.367
R1128 B.n7 B.n6 163.367
R1129 B.n404 B.n7 163.367
R1130 B.n405 B.n404 163.367
R1131 B.n405 B.n13 163.367
R1132 B.n14 B.n13 163.367
R1133 B.n15 B.n14 163.367
R1134 B.n410 B.n15 163.367
R1135 B.n410 B.n20 163.367
R1136 B.n21 B.n20 163.367
R1137 B.n22 B.n21 163.367
R1138 B.n415 B.n22 163.367
R1139 B.n415 B.n27 163.367
R1140 B.n28 B.n27 163.367
R1141 B.n29 B.n28 163.367
R1142 B.n353 B.n351 163.367
R1143 B.n351 B.n350 163.367
R1144 B.n347 B.n346 163.367
R1145 B.n344 B.n114 163.367
R1146 B.n340 B.n338 163.367
R1147 B.n336 B.n116 163.367
R1148 B.n332 B.n330 163.367
R1149 B.n328 B.n118 163.367
R1150 B.n324 B.n322 163.367
R1151 B.n320 B.n120 163.367
R1152 B.n316 B.n314 163.367
R1153 B.n312 B.n122 163.367
R1154 B.n308 B.n306 163.367
R1155 B.n304 B.n124 163.367
R1156 B.n300 B.n298 163.367
R1157 B.n296 B.n126 163.367
R1158 B.n292 B.n290 163.367
R1159 B.n288 B.n128 163.367
R1160 B.n284 B.n282 163.367
R1161 B.n280 B.n130 163.367
R1162 B.n276 B.n274 163.367
R1163 B.n272 B.n132 163.367
R1164 B.n267 B.n265 163.367
R1165 B.n263 B.n136 163.367
R1166 B.n259 B.n257 163.367
R1167 B.n255 B.n138 163.367
R1168 B.n251 B.n249 163.367
R1169 B.n246 B.n245 163.367
R1170 B.n243 B.n144 163.367
R1171 B.n239 B.n237 163.367
R1172 B.n235 B.n146 163.367
R1173 B.n231 B.n229 163.367
R1174 B.n227 B.n148 163.367
R1175 B.n223 B.n221 163.367
R1176 B.n219 B.n150 163.367
R1177 B.n215 B.n213 163.367
R1178 B.n211 B.n152 163.367
R1179 B.n207 B.n205 163.367
R1180 B.n203 B.n154 163.367
R1181 B.n199 B.n197 163.367
R1182 B.n195 B.n156 163.367
R1183 B.n191 B.n189 163.367
R1184 B.n187 B.n158 163.367
R1185 B.n183 B.n181 163.367
R1186 B.n179 B.n160 163.367
R1187 B.n175 B.n173 163.367
R1188 B.n171 B.n162 163.367
R1189 B.n167 B.n165 163.367
R1190 B.n357 B.n104 163.367
R1191 B.n365 B.n104 163.367
R1192 B.n365 B.n102 163.367
R1193 B.n369 B.n102 163.367
R1194 B.n369 B.n96 163.367
R1195 B.n377 B.n96 163.367
R1196 B.n377 B.n94 163.367
R1197 B.n381 B.n94 163.367
R1198 B.n381 B.n88 163.367
R1199 B.n391 B.n88 163.367
R1200 B.n391 B.n86 163.367
R1201 B.n395 B.n86 163.367
R1202 B.n395 B.n3 163.367
R1203 B.n645 B.n3 163.367
R1204 B.n641 B.n2 163.367
R1205 B.n641 B.n640 163.367
R1206 B.n640 B.n9 163.367
R1207 B.n636 B.n9 163.367
R1208 B.n636 B.n11 163.367
R1209 B.n632 B.n11 163.367
R1210 B.n632 B.n17 163.367
R1211 B.n628 B.n17 163.367
R1212 B.n628 B.n19 163.367
R1213 B.n624 B.n19 163.367
R1214 B.n624 B.n24 163.367
R1215 B.n620 B.n24 163.367
R1216 B.n620 B.n26 163.367
R1217 B.n616 B.n26 163.367
R1218 B.n611 B.n31 71.676
R1219 B.n610 B.n609 71.676
R1220 B.n603 B.n33 71.676
R1221 B.n602 B.n601 71.676
R1222 B.n595 B.n35 71.676
R1223 B.n594 B.n593 71.676
R1224 B.n587 B.n37 71.676
R1225 B.n586 B.n585 71.676
R1226 B.n579 B.n39 71.676
R1227 B.n578 B.n577 71.676
R1228 B.n571 B.n41 71.676
R1229 B.n570 B.n569 71.676
R1230 B.n563 B.n43 71.676
R1231 B.n562 B.n561 71.676
R1232 B.n555 B.n45 71.676
R1233 B.n554 B.n553 71.676
R1234 B.n547 B.n47 71.676
R1235 B.n546 B.n545 71.676
R1236 B.n539 B.n49 71.676
R1237 B.n538 B.n537 71.676
R1238 B.n531 B.n51 71.676
R1239 B.n530 B.n529 71.676
R1240 B.n522 B.n53 71.676
R1241 B.n521 B.n520 71.676
R1242 B.n514 B.n57 71.676
R1243 B.n513 B.n512 71.676
R1244 B.n505 B.n59 71.676
R1245 B.n504 B.n503 71.676
R1246 B.n497 B.n63 71.676
R1247 B.n496 B.n495 71.676
R1248 B.n489 B.n65 71.676
R1249 B.n488 B.n487 71.676
R1250 B.n481 B.n67 71.676
R1251 B.n480 B.n479 71.676
R1252 B.n473 B.n69 71.676
R1253 B.n472 B.n471 71.676
R1254 B.n465 B.n71 71.676
R1255 B.n464 B.n463 71.676
R1256 B.n457 B.n73 71.676
R1257 B.n456 B.n455 71.676
R1258 B.n449 B.n75 71.676
R1259 B.n448 B.n447 71.676
R1260 B.n441 B.n77 71.676
R1261 B.n440 B.n439 71.676
R1262 B.n433 B.n79 71.676
R1263 B.n432 B.n431 71.676
R1264 B.n425 B.n81 71.676
R1265 B.n424 B.n423 71.676
R1266 B.n423 B.n422 71.676
R1267 B.n426 B.n425 71.676
R1268 B.n431 B.n430 71.676
R1269 B.n434 B.n433 71.676
R1270 B.n439 B.n438 71.676
R1271 B.n442 B.n441 71.676
R1272 B.n447 B.n446 71.676
R1273 B.n450 B.n449 71.676
R1274 B.n455 B.n454 71.676
R1275 B.n458 B.n457 71.676
R1276 B.n463 B.n462 71.676
R1277 B.n466 B.n465 71.676
R1278 B.n471 B.n470 71.676
R1279 B.n474 B.n473 71.676
R1280 B.n479 B.n478 71.676
R1281 B.n482 B.n481 71.676
R1282 B.n487 B.n486 71.676
R1283 B.n490 B.n489 71.676
R1284 B.n495 B.n494 71.676
R1285 B.n498 B.n497 71.676
R1286 B.n503 B.n502 71.676
R1287 B.n506 B.n505 71.676
R1288 B.n512 B.n511 71.676
R1289 B.n515 B.n514 71.676
R1290 B.n520 B.n519 71.676
R1291 B.n523 B.n522 71.676
R1292 B.n529 B.n528 71.676
R1293 B.n532 B.n531 71.676
R1294 B.n537 B.n536 71.676
R1295 B.n540 B.n539 71.676
R1296 B.n545 B.n544 71.676
R1297 B.n548 B.n547 71.676
R1298 B.n553 B.n552 71.676
R1299 B.n556 B.n555 71.676
R1300 B.n561 B.n560 71.676
R1301 B.n564 B.n563 71.676
R1302 B.n569 B.n568 71.676
R1303 B.n572 B.n571 71.676
R1304 B.n577 B.n576 71.676
R1305 B.n580 B.n579 71.676
R1306 B.n585 B.n584 71.676
R1307 B.n588 B.n587 71.676
R1308 B.n593 B.n592 71.676
R1309 B.n596 B.n595 71.676
R1310 B.n601 B.n600 71.676
R1311 B.n604 B.n603 71.676
R1312 B.n609 B.n608 71.676
R1313 B.n612 B.n611 71.676
R1314 B.n352 B.n110 71.676
R1315 B.n350 B.n112 71.676
R1316 B.n346 B.n345 71.676
R1317 B.n339 B.n114 71.676
R1318 B.n338 B.n337 71.676
R1319 B.n331 B.n116 71.676
R1320 B.n330 B.n329 71.676
R1321 B.n323 B.n118 71.676
R1322 B.n322 B.n321 71.676
R1323 B.n315 B.n120 71.676
R1324 B.n314 B.n313 71.676
R1325 B.n307 B.n122 71.676
R1326 B.n306 B.n305 71.676
R1327 B.n299 B.n124 71.676
R1328 B.n298 B.n297 71.676
R1329 B.n291 B.n126 71.676
R1330 B.n290 B.n289 71.676
R1331 B.n283 B.n128 71.676
R1332 B.n282 B.n281 71.676
R1333 B.n275 B.n130 71.676
R1334 B.n274 B.n273 71.676
R1335 B.n266 B.n132 71.676
R1336 B.n265 B.n264 71.676
R1337 B.n258 B.n136 71.676
R1338 B.n257 B.n256 71.676
R1339 B.n250 B.n138 71.676
R1340 B.n249 B.n142 71.676
R1341 B.n245 B.n244 71.676
R1342 B.n238 B.n144 71.676
R1343 B.n237 B.n236 71.676
R1344 B.n230 B.n146 71.676
R1345 B.n229 B.n228 71.676
R1346 B.n222 B.n148 71.676
R1347 B.n221 B.n220 71.676
R1348 B.n214 B.n150 71.676
R1349 B.n213 B.n212 71.676
R1350 B.n206 B.n152 71.676
R1351 B.n205 B.n204 71.676
R1352 B.n198 B.n154 71.676
R1353 B.n197 B.n196 71.676
R1354 B.n190 B.n156 71.676
R1355 B.n189 B.n188 71.676
R1356 B.n182 B.n158 71.676
R1357 B.n181 B.n180 71.676
R1358 B.n174 B.n160 71.676
R1359 B.n173 B.n172 71.676
R1360 B.n166 B.n162 71.676
R1361 B.n165 B.n164 71.676
R1362 B.n353 B.n352 71.676
R1363 B.n347 B.n112 71.676
R1364 B.n345 B.n344 71.676
R1365 B.n340 B.n339 71.676
R1366 B.n337 B.n336 71.676
R1367 B.n332 B.n331 71.676
R1368 B.n329 B.n328 71.676
R1369 B.n324 B.n323 71.676
R1370 B.n321 B.n320 71.676
R1371 B.n316 B.n315 71.676
R1372 B.n313 B.n312 71.676
R1373 B.n308 B.n307 71.676
R1374 B.n305 B.n304 71.676
R1375 B.n300 B.n299 71.676
R1376 B.n297 B.n296 71.676
R1377 B.n292 B.n291 71.676
R1378 B.n289 B.n288 71.676
R1379 B.n284 B.n283 71.676
R1380 B.n281 B.n280 71.676
R1381 B.n276 B.n275 71.676
R1382 B.n273 B.n272 71.676
R1383 B.n267 B.n266 71.676
R1384 B.n264 B.n263 71.676
R1385 B.n259 B.n258 71.676
R1386 B.n256 B.n255 71.676
R1387 B.n251 B.n250 71.676
R1388 B.n246 B.n142 71.676
R1389 B.n244 B.n243 71.676
R1390 B.n239 B.n238 71.676
R1391 B.n236 B.n235 71.676
R1392 B.n231 B.n230 71.676
R1393 B.n228 B.n227 71.676
R1394 B.n223 B.n222 71.676
R1395 B.n220 B.n219 71.676
R1396 B.n215 B.n214 71.676
R1397 B.n212 B.n211 71.676
R1398 B.n207 B.n206 71.676
R1399 B.n204 B.n203 71.676
R1400 B.n199 B.n198 71.676
R1401 B.n196 B.n195 71.676
R1402 B.n191 B.n190 71.676
R1403 B.n188 B.n187 71.676
R1404 B.n183 B.n182 71.676
R1405 B.n180 B.n179 71.676
R1406 B.n175 B.n174 71.676
R1407 B.n172 B.n171 71.676
R1408 B.n167 B.n166 71.676
R1409 B.n164 B.n108 71.676
R1410 B.n646 B.n645 71.676
R1411 B.n646 B.n2 71.676
R1412 B.n358 B.n109 71.5601
R1413 B.n617 B.n30 71.5601
R1414 B.n526 B.n55 59.5399
R1415 B.n508 B.n61 59.5399
R1416 B.n141 B.n140 59.5399
R1417 B.n269 B.n134 59.5399
R1418 B.n358 B.n105 41.5907
R1419 B.n364 B.n105 41.5907
R1420 B.n364 B.n101 41.5907
R1421 B.n370 B.n101 41.5907
R1422 B.n376 B.n97 41.5907
R1423 B.n376 B.n93 41.5907
R1424 B.n382 B.n93 41.5907
R1425 B.n382 B.n89 41.5907
R1426 B.n390 B.n89 41.5907
R1427 B.n390 B.n389 41.5907
R1428 B.n396 B.n4 41.5907
R1429 B.n644 B.n4 41.5907
R1430 B.n644 B.n643 41.5907
R1431 B.n643 B.n642 41.5907
R1432 B.n642 B.n8 41.5907
R1433 B.n635 B.n12 41.5907
R1434 B.n635 B.n634 41.5907
R1435 B.n634 B.n633 41.5907
R1436 B.n633 B.n16 41.5907
R1437 B.n627 B.n16 41.5907
R1438 B.n627 B.n626 41.5907
R1439 B.n625 B.n23 41.5907
R1440 B.n619 B.n23 41.5907
R1441 B.n619 B.n618 41.5907
R1442 B.n618 B.n617 41.5907
R1443 B.n370 B.t10 40.3675
R1444 B.t3 B.n625 40.3675
R1445 B.n356 B.n355 31.3761
R1446 B.n360 B.n107 31.3761
R1447 B.n420 B.n419 31.3761
R1448 B.n615 B.n614 31.3761
R1449 B.n396 B.t0 28.1351
R1450 B.t1 B.n8 28.1351
R1451 B.n55 B.n54 20.752
R1452 B.n61 B.n60 20.752
R1453 B.n140 B.n139 20.752
R1454 B.n134 B.n133 20.752
R1455 B B.n647 18.0485
R1456 B.n389 B.t0 13.4562
R1457 B.n12 B.t1 13.4562
R1458 B.n356 B.n103 10.6151
R1459 B.n366 B.n103 10.6151
R1460 B.n367 B.n366 10.6151
R1461 B.n368 B.n367 10.6151
R1462 B.n368 B.n95 10.6151
R1463 B.n378 B.n95 10.6151
R1464 B.n379 B.n378 10.6151
R1465 B.n380 B.n379 10.6151
R1466 B.n380 B.n87 10.6151
R1467 B.n392 B.n87 10.6151
R1468 B.n393 B.n392 10.6151
R1469 B.n394 B.n393 10.6151
R1470 B.n394 B.n0 10.6151
R1471 B.n355 B.n354 10.6151
R1472 B.n354 B.n111 10.6151
R1473 B.n349 B.n111 10.6151
R1474 B.n349 B.n348 10.6151
R1475 B.n348 B.n113 10.6151
R1476 B.n343 B.n113 10.6151
R1477 B.n343 B.n342 10.6151
R1478 B.n342 B.n341 10.6151
R1479 B.n341 B.n115 10.6151
R1480 B.n335 B.n115 10.6151
R1481 B.n335 B.n334 10.6151
R1482 B.n334 B.n333 10.6151
R1483 B.n333 B.n117 10.6151
R1484 B.n327 B.n117 10.6151
R1485 B.n327 B.n326 10.6151
R1486 B.n326 B.n325 10.6151
R1487 B.n325 B.n119 10.6151
R1488 B.n319 B.n119 10.6151
R1489 B.n319 B.n318 10.6151
R1490 B.n318 B.n317 10.6151
R1491 B.n317 B.n121 10.6151
R1492 B.n311 B.n121 10.6151
R1493 B.n311 B.n310 10.6151
R1494 B.n310 B.n309 10.6151
R1495 B.n309 B.n123 10.6151
R1496 B.n303 B.n123 10.6151
R1497 B.n303 B.n302 10.6151
R1498 B.n302 B.n301 10.6151
R1499 B.n301 B.n125 10.6151
R1500 B.n295 B.n125 10.6151
R1501 B.n295 B.n294 10.6151
R1502 B.n294 B.n293 10.6151
R1503 B.n293 B.n127 10.6151
R1504 B.n287 B.n127 10.6151
R1505 B.n287 B.n286 10.6151
R1506 B.n286 B.n285 10.6151
R1507 B.n285 B.n129 10.6151
R1508 B.n279 B.n129 10.6151
R1509 B.n279 B.n278 10.6151
R1510 B.n278 B.n277 10.6151
R1511 B.n277 B.n131 10.6151
R1512 B.n271 B.n131 10.6151
R1513 B.n271 B.n270 10.6151
R1514 B.n268 B.n135 10.6151
R1515 B.n262 B.n135 10.6151
R1516 B.n262 B.n261 10.6151
R1517 B.n261 B.n260 10.6151
R1518 B.n260 B.n137 10.6151
R1519 B.n254 B.n137 10.6151
R1520 B.n254 B.n253 10.6151
R1521 B.n253 B.n252 10.6151
R1522 B.n248 B.n247 10.6151
R1523 B.n247 B.n143 10.6151
R1524 B.n242 B.n143 10.6151
R1525 B.n242 B.n241 10.6151
R1526 B.n241 B.n240 10.6151
R1527 B.n240 B.n145 10.6151
R1528 B.n234 B.n145 10.6151
R1529 B.n234 B.n233 10.6151
R1530 B.n233 B.n232 10.6151
R1531 B.n232 B.n147 10.6151
R1532 B.n226 B.n147 10.6151
R1533 B.n226 B.n225 10.6151
R1534 B.n225 B.n224 10.6151
R1535 B.n224 B.n149 10.6151
R1536 B.n218 B.n149 10.6151
R1537 B.n218 B.n217 10.6151
R1538 B.n217 B.n216 10.6151
R1539 B.n216 B.n151 10.6151
R1540 B.n210 B.n151 10.6151
R1541 B.n210 B.n209 10.6151
R1542 B.n209 B.n208 10.6151
R1543 B.n208 B.n153 10.6151
R1544 B.n202 B.n153 10.6151
R1545 B.n202 B.n201 10.6151
R1546 B.n201 B.n200 10.6151
R1547 B.n200 B.n155 10.6151
R1548 B.n194 B.n155 10.6151
R1549 B.n194 B.n193 10.6151
R1550 B.n193 B.n192 10.6151
R1551 B.n192 B.n157 10.6151
R1552 B.n186 B.n157 10.6151
R1553 B.n186 B.n185 10.6151
R1554 B.n185 B.n184 10.6151
R1555 B.n184 B.n159 10.6151
R1556 B.n178 B.n159 10.6151
R1557 B.n178 B.n177 10.6151
R1558 B.n177 B.n176 10.6151
R1559 B.n176 B.n161 10.6151
R1560 B.n170 B.n161 10.6151
R1561 B.n170 B.n169 10.6151
R1562 B.n169 B.n168 10.6151
R1563 B.n168 B.n163 10.6151
R1564 B.n163 B.n107 10.6151
R1565 B.n361 B.n360 10.6151
R1566 B.n362 B.n361 10.6151
R1567 B.n362 B.n99 10.6151
R1568 B.n372 B.n99 10.6151
R1569 B.n373 B.n372 10.6151
R1570 B.n374 B.n373 10.6151
R1571 B.n374 B.n91 10.6151
R1572 B.n384 B.n91 10.6151
R1573 B.n385 B.n384 10.6151
R1574 B.n387 B.n385 10.6151
R1575 B.n387 B.n386 10.6151
R1576 B.n386 B.n84 10.6151
R1577 B.n399 B.n84 10.6151
R1578 B.n400 B.n399 10.6151
R1579 B.n401 B.n400 10.6151
R1580 B.n402 B.n401 10.6151
R1581 B.n403 B.n402 10.6151
R1582 B.n406 B.n403 10.6151
R1583 B.n407 B.n406 10.6151
R1584 B.n408 B.n407 10.6151
R1585 B.n409 B.n408 10.6151
R1586 B.n411 B.n409 10.6151
R1587 B.n412 B.n411 10.6151
R1588 B.n413 B.n412 10.6151
R1589 B.n414 B.n413 10.6151
R1590 B.n416 B.n414 10.6151
R1591 B.n417 B.n416 10.6151
R1592 B.n418 B.n417 10.6151
R1593 B.n419 B.n418 10.6151
R1594 B.n639 B.n1 10.6151
R1595 B.n639 B.n638 10.6151
R1596 B.n638 B.n637 10.6151
R1597 B.n637 B.n10 10.6151
R1598 B.n631 B.n10 10.6151
R1599 B.n631 B.n630 10.6151
R1600 B.n630 B.n629 10.6151
R1601 B.n629 B.n18 10.6151
R1602 B.n623 B.n18 10.6151
R1603 B.n623 B.n622 10.6151
R1604 B.n622 B.n621 10.6151
R1605 B.n621 B.n25 10.6151
R1606 B.n615 B.n25 10.6151
R1607 B.n614 B.n613 10.6151
R1608 B.n613 B.n32 10.6151
R1609 B.n607 B.n32 10.6151
R1610 B.n607 B.n606 10.6151
R1611 B.n606 B.n605 10.6151
R1612 B.n605 B.n34 10.6151
R1613 B.n599 B.n34 10.6151
R1614 B.n599 B.n598 10.6151
R1615 B.n598 B.n597 10.6151
R1616 B.n597 B.n36 10.6151
R1617 B.n591 B.n36 10.6151
R1618 B.n591 B.n590 10.6151
R1619 B.n590 B.n589 10.6151
R1620 B.n589 B.n38 10.6151
R1621 B.n583 B.n38 10.6151
R1622 B.n583 B.n582 10.6151
R1623 B.n582 B.n581 10.6151
R1624 B.n581 B.n40 10.6151
R1625 B.n575 B.n40 10.6151
R1626 B.n575 B.n574 10.6151
R1627 B.n574 B.n573 10.6151
R1628 B.n573 B.n42 10.6151
R1629 B.n567 B.n42 10.6151
R1630 B.n567 B.n566 10.6151
R1631 B.n566 B.n565 10.6151
R1632 B.n565 B.n44 10.6151
R1633 B.n559 B.n44 10.6151
R1634 B.n559 B.n558 10.6151
R1635 B.n558 B.n557 10.6151
R1636 B.n557 B.n46 10.6151
R1637 B.n551 B.n46 10.6151
R1638 B.n551 B.n550 10.6151
R1639 B.n550 B.n549 10.6151
R1640 B.n549 B.n48 10.6151
R1641 B.n543 B.n48 10.6151
R1642 B.n543 B.n542 10.6151
R1643 B.n542 B.n541 10.6151
R1644 B.n541 B.n50 10.6151
R1645 B.n535 B.n50 10.6151
R1646 B.n535 B.n534 10.6151
R1647 B.n534 B.n533 10.6151
R1648 B.n533 B.n52 10.6151
R1649 B.n527 B.n52 10.6151
R1650 B.n525 B.n524 10.6151
R1651 B.n524 B.n56 10.6151
R1652 B.n518 B.n56 10.6151
R1653 B.n518 B.n517 10.6151
R1654 B.n517 B.n516 10.6151
R1655 B.n516 B.n58 10.6151
R1656 B.n510 B.n58 10.6151
R1657 B.n510 B.n509 10.6151
R1658 B.n507 B.n62 10.6151
R1659 B.n501 B.n62 10.6151
R1660 B.n501 B.n500 10.6151
R1661 B.n500 B.n499 10.6151
R1662 B.n499 B.n64 10.6151
R1663 B.n493 B.n64 10.6151
R1664 B.n493 B.n492 10.6151
R1665 B.n492 B.n491 10.6151
R1666 B.n491 B.n66 10.6151
R1667 B.n485 B.n66 10.6151
R1668 B.n485 B.n484 10.6151
R1669 B.n484 B.n483 10.6151
R1670 B.n483 B.n68 10.6151
R1671 B.n477 B.n68 10.6151
R1672 B.n477 B.n476 10.6151
R1673 B.n476 B.n475 10.6151
R1674 B.n475 B.n70 10.6151
R1675 B.n469 B.n70 10.6151
R1676 B.n469 B.n468 10.6151
R1677 B.n468 B.n467 10.6151
R1678 B.n467 B.n72 10.6151
R1679 B.n461 B.n72 10.6151
R1680 B.n461 B.n460 10.6151
R1681 B.n460 B.n459 10.6151
R1682 B.n459 B.n74 10.6151
R1683 B.n453 B.n74 10.6151
R1684 B.n453 B.n452 10.6151
R1685 B.n452 B.n451 10.6151
R1686 B.n451 B.n76 10.6151
R1687 B.n445 B.n76 10.6151
R1688 B.n445 B.n444 10.6151
R1689 B.n444 B.n443 10.6151
R1690 B.n443 B.n78 10.6151
R1691 B.n437 B.n78 10.6151
R1692 B.n437 B.n436 10.6151
R1693 B.n436 B.n435 10.6151
R1694 B.n435 B.n80 10.6151
R1695 B.n429 B.n80 10.6151
R1696 B.n429 B.n428 10.6151
R1697 B.n428 B.n427 10.6151
R1698 B.n427 B.n82 10.6151
R1699 B.n421 B.n82 10.6151
R1700 B.n421 B.n420 10.6151
R1701 B.n647 B.n0 8.11757
R1702 B.n647 B.n1 8.11757
R1703 B.n269 B.n268 7.18099
R1704 B.n252 B.n141 7.18099
R1705 B.n526 B.n525 7.18099
R1706 B.n509 B.n508 7.18099
R1707 B.n270 B.n269 3.43465
R1708 B.n248 B.n141 3.43465
R1709 B.n527 B.n526 3.43465
R1710 B.n508 B.n507 3.43465
R1711 B.t10 B.n97 1.22374
R1712 B.n626 B.t3 1.22374
R1713 VN VN.t0 668.635
R1714 VN VN.t1 628.044
R1715 VDD2.n137 VDD2.n136 289.615
R1716 VDD2.n68 VDD2.n67 289.615
R1717 VDD2.n136 VDD2.n135 185
R1718 VDD2.n71 VDD2.n70 185
R1719 VDD2.n130 VDD2.n129 185
R1720 VDD2.n128 VDD2.n127 185
R1721 VDD2.n75 VDD2.n74 185
R1722 VDD2.n122 VDD2.n121 185
R1723 VDD2.n120 VDD2.n119 185
R1724 VDD2.n79 VDD2.n78 185
R1725 VDD2.n114 VDD2.n113 185
R1726 VDD2.n112 VDD2.n111 185
R1727 VDD2.n83 VDD2.n82 185
R1728 VDD2.n106 VDD2.n105 185
R1729 VDD2.n104 VDD2.n103 185
R1730 VDD2.n87 VDD2.n86 185
R1731 VDD2.n98 VDD2.n97 185
R1732 VDD2.n96 VDD2.n95 185
R1733 VDD2.n91 VDD2.n90 185
R1734 VDD2.n22 VDD2.n21 185
R1735 VDD2.n27 VDD2.n26 185
R1736 VDD2.n29 VDD2.n28 185
R1737 VDD2.n18 VDD2.n17 185
R1738 VDD2.n35 VDD2.n34 185
R1739 VDD2.n37 VDD2.n36 185
R1740 VDD2.n14 VDD2.n13 185
R1741 VDD2.n43 VDD2.n42 185
R1742 VDD2.n45 VDD2.n44 185
R1743 VDD2.n10 VDD2.n9 185
R1744 VDD2.n51 VDD2.n50 185
R1745 VDD2.n53 VDD2.n52 185
R1746 VDD2.n6 VDD2.n5 185
R1747 VDD2.n59 VDD2.n58 185
R1748 VDD2.n61 VDD2.n60 185
R1749 VDD2.n2 VDD2.n1 185
R1750 VDD2.n67 VDD2.n66 185
R1751 VDD2.n23 VDD2.t0 147.659
R1752 VDD2.n92 VDD2.t1 147.659
R1753 VDD2.n136 VDD2.n70 104.615
R1754 VDD2.n129 VDD2.n70 104.615
R1755 VDD2.n129 VDD2.n128 104.615
R1756 VDD2.n128 VDD2.n74 104.615
R1757 VDD2.n121 VDD2.n74 104.615
R1758 VDD2.n121 VDD2.n120 104.615
R1759 VDD2.n120 VDD2.n78 104.615
R1760 VDD2.n113 VDD2.n78 104.615
R1761 VDD2.n113 VDD2.n112 104.615
R1762 VDD2.n112 VDD2.n82 104.615
R1763 VDD2.n105 VDD2.n82 104.615
R1764 VDD2.n105 VDD2.n104 104.615
R1765 VDD2.n104 VDD2.n86 104.615
R1766 VDD2.n97 VDD2.n86 104.615
R1767 VDD2.n97 VDD2.n96 104.615
R1768 VDD2.n96 VDD2.n90 104.615
R1769 VDD2.n27 VDD2.n21 104.615
R1770 VDD2.n28 VDD2.n27 104.615
R1771 VDD2.n28 VDD2.n17 104.615
R1772 VDD2.n35 VDD2.n17 104.615
R1773 VDD2.n36 VDD2.n35 104.615
R1774 VDD2.n36 VDD2.n13 104.615
R1775 VDD2.n43 VDD2.n13 104.615
R1776 VDD2.n44 VDD2.n43 104.615
R1777 VDD2.n44 VDD2.n9 104.615
R1778 VDD2.n51 VDD2.n9 104.615
R1779 VDD2.n52 VDD2.n51 104.615
R1780 VDD2.n52 VDD2.n5 104.615
R1781 VDD2.n59 VDD2.n5 104.615
R1782 VDD2.n60 VDD2.n59 104.615
R1783 VDD2.n60 VDD2.n1 104.615
R1784 VDD2.n67 VDD2.n1 104.615
R1785 VDD2.n138 VDD2.n68 89.0102
R1786 VDD2.n138 VDD2.n137 52.549
R1787 VDD2.t1 VDD2.n90 52.3082
R1788 VDD2.t0 VDD2.n21 52.3082
R1789 VDD2.n92 VDD2.n91 15.6677
R1790 VDD2.n23 VDD2.n22 15.6677
R1791 VDD2.n135 VDD2.n69 12.8005
R1792 VDD2.n95 VDD2.n94 12.8005
R1793 VDD2.n26 VDD2.n25 12.8005
R1794 VDD2.n66 VDD2.n0 12.8005
R1795 VDD2.n134 VDD2.n71 12.0247
R1796 VDD2.n98 VDD2.n89 12.0247
R1797 VDD2.n29 VDD2.n20 12.0247
R1798 VDD2.n65 VDD2.n2 12.0247
R1799 VDD2.n131 VDD2.n130 11.249
R1800 VDD2.n99 VDD2.n87 11.249
R1801 VDD2.n30 VDD2.n18 11.249
R1802 VDD2.n62 VDD2.n61 11.249
R1803 VDD2.n127 VDD2.n73 10.4732
R1804 VDD2.n103 VDD2.n102 10.4732
R1805 VDD2.n34 VDD2.n33 10.4732
R1806 VDD2.n58 VDD2.n4 10.4732
R1807 VDD2.n126 VDD2.n75 9.69747
R1808 VDD2.n106 VDD2.n85 9.69747
R1809 VDD2.n37 VDD2.n16 9.69747
R1810 VDD2.n57 VDD2.n6 9.69747
R1811 VDD2.n133 VDD2.n69 9.45567
R1812 VDD2.n64 VDD2.n0 9.45567
R1813 VDD2.n134 VDD2.n133 9.3005
R1814 VDD2.n132 VDD2.n131 9.3005
R1815 VDD2.n73 VDD2.n72 9.3005
R1816 VDD2.n126 VDD2.n125 9.3005
R1817 VDD2.n124 VDD2.n123 9.3005
R1818 VDD2.n77 VDD2.n76 9.3005
R1819 VDD2.n118 VDD2.n117 9.3005
R1820 VDD2.n116 VDD2.n115 9.3005
R1821 VDD2.n81 VDD2.n80 9.3005
R1822 VDD2.n110 VDD2.n109 9.3005
R1823 VDD2.n108 VDD2.n107 9.3005
R1824 VDD2.n85 VDD2.n84 9.3005
R1825 VDD2.n102 VDD2.n101 9.3005
R1826 VDD2.n100 VDD2.n99 9.3005
R1827 VDD2.n89 VDD2.n88 9.3005
R1828 VDD2.n94 VDD2.n93 9.3005
R1829 VDD2.n47 VDD2.n46 9.3005
R1830 VDD2.n49 VDD2.n48 9.3005
R1831 VDD2.n8 VDD2.n7 9.3005
R1832 VDD2.n55 VDD2.n54 9.3005
R1833 VDD2.n57 VDD2.n56 9.3005
R1834 VDD2.n4 VDD2.n3 9.3005
R1835 VDD2.n63 VDD2.n62 9.3005
R1836 VDD2.n65 VDD2.n64 9.3005
R1837 VDD2.n41 VDD2.n40 9.3005
R1838 VDD2.n39 VDD2.n38 9.3005
R1839 VDD2.n16 VDD2.n15 9.3005
R1840 VDD2.n33 VDD2.n32 9.3005
R1841 VDD2.n31 VDD2.n30 9.3005
R1842 VDD2.n20 VDD2.n19 9.3005
R1843 VDD2.n25 VDD2.n24 9.3005
R1844 VDD2.n12 VDD2.n11 9.3005
R1845 VDD2.n123 VDD2.n122 8.92171
R1846 VDD2.n107 VDD2.n83 8.92171
R1847 VDD2.n38 VDD2.n14 8.92171
R1848 VDD2.n54 VDD2.n53 8.92171
R1849 VDD2.n119 VDD2.n77 8.14595
R1850 VDD2.n111 VDD2.n110 8.14595
R1851 VDD2.n42 VDD2.n41 8.14595
R1852 VDD2.n50 VDD2.n8 8.14595
R1853 VDD2.n118 VDD2.n79 7.3702
R1854 VDD2.n114 VDD2.n81 7.3702
R1855 VDD2.n45 VDD2.n12 7.3702
R1856 VDD2.n49 VDD2.n10 7.3702
R1857 VDD2.n115 VDD2.n79 6.59444
R1858 VDD2.n115 VDD2.n114 6.59444
R1859 VDD2.n46 VDD2.n45 6.59444
R1860 VDD2.n46 VDD2.n10 6.59444
R1861 VDD2.n119 VDD2.n118 5.81868
R1862 VDD2.n111 VDD2.n81 5.81868
R1863 VDD2.n42 VDD2.n12 5.81868
R1864 VDD2.n50 VDD2.n49 5.81868
R1865 VDD2.n122 VDD2.n77 5.04292
R1866 VDD2.n110 VDD2.n83 5.04292
R1867 VDD2.n41 VDD2.n14 5.04292
R1868 VDD2.n53 VDD2.n8 5.04292
R1869 VDD2.n24 VDD2.n23 4.38563
R1870 VDD2.n93 VDD2.n92 4.38563
R1871 VDD2.n123 VDD2.n75 4.26717
R1872 VDD2.n107 VDD2.n106 4.26717
R1873 VDD2.n38 VDD2.n37 4.26717
R1874 VDD2.n54 VDD2.n6 4.26717
R1875 VDD2.n127 VDD2.n126 3.49141
R1876 VDD2.n103 VDD2.n85 3.49141
R1877 VDD2.n34 VDD2.n16 3.49141
R1878 VDD2.n58 VDD2.n57 3.49141
R1879 VDD2.n130 VDD2.n73 2.71565
R1880 VDD2.n102 VDD2.n87 2.71565
R1881 VDD2.n33 VDD2.n18 2.71565
R1882 VDD2.n61 VDD2.n4 2.71565
R1883 VDD2.n131 VDD2.n71 1.93989
R1884 VDD2.n99 VDD2.n98 1.93989
R1885 VDD2.n30 VDD2.n29 1.93989
R1886 VDD2.n62 VDD2.n2 1.93989
R1887 VDD2.n135 VDD2.n134 1.16414
R1888 VDD2.n95 VDD2.n89 1.16414
R1889 VDD2.n26 VDD2.n20 1.16414
R1890 VDD2.n66 VDD2.n65 1.16414
R1891 VDD2.n137 VDD2.n69 0.388379
R1892 VDD2.n94 VDD2.n91 0.388379
R1893 VDD2.n25 VDD2.n22 0.388379
R1894 VDD2.n68 VDD2.n0 0.388379
R1895 VDD2 VDD2.n138 0.289293
R1896 VDD2.n133 VDD2.n132 0.155672
R1897 VDD2.n132 VDD2.n72 0.155672
R1898 VDD2.n125 VDD2.n72 0.155672
R1899 VDD2.n125 VDD2.n124 0.155672
R1900 VDD2.n124 VDD2.n76 0.155672
R1901 VDD2.n117 VDD2.n76 0.155672
R1902 VDD2.n117 VDD2.n116 0.155672
R1903 VDD2.n116 VDD2.n80 0.155672
R1904 VDD2.n109 VDD2.n80 0.155672
R1905 VDD2.n109 VDD2.n108 0.155672
R1906 VDD2.n108 VDD2.n84 0.155672
R1907 VDD2.n101 VDD2.n84 0.155672
R1908 VDD2.n101 VDD2.n100 0.155672
R1909 VDD2.n100 VDD2.n88 0.155672
R1910 VDD2.n93 VDD2.n88 0.155672
R1911 VDD2.n24 VDD2.n19 0.155672
R1912 VDD2.n31 VDD2.n19 0.155672
R1913 VDD2.n32 VDD2.n31 0.155672
R1914 VDD2.n32 VDD2.n15 0.155672
R1915 VDD2.n39 VDD2.n15 0.155672
R1916 VDD2.n40 VDD2.n39 0.155672
R1917 VDD2.n40 VDD2.n11 0.155672
R1918 VDD2.n47 VDD2.n11 0.155672
R1919 VDD2.n48 VDD2.n47 0.155672
R1920 VDD2.n48 VDD2.n7 0.155672
R1921 VDD2.n55 VDD2.n7 0.155672
R1922 VDD2.n56 VDD2.n55 0.155672
R1923 VDD2.n56 VDD2.n3 0.155672
R1924 VDD2.n63 VDD2.n3 0.155672
R1925 VDD2.n64 VDD2.n63 0.155672
C0 VP VN 4.70762f
C1 VN VDD1 0.148607f
C2 VN VDD2 2.12749f
C3 VP VDD1 2.23112f
C4 VP VDD2 0.256763f
C5 VN VTAIL 1.5967f
C6 VDD1 VDD2 0.466174f
C7 VP VTAIL 1.61132f
C8 VTAIL VDD1 5.84165f
C9 VTAIL VDD2 5.87554f
C10 VDD2 B 3.894832f
C11 VDD1 B 6.381f
C12 VTAIL B 6.664948f
C13 VN B 8.27609f
C14 VP B 4.124895f
C15 VDD2.n0 B 0.011754f
C16 VDD2.n1 B 0.026469f
C17 VDD2.n2 B 0.011857f
C18 VDD2.n3 B 0.02084f
C19 VDD2.n4 B 0.011198f
C20 VDD2.n5 B 0.026469f
C21 VDD2.n6 B 0.011857f
C22 VDD2.n7 B 0.02084f
C23 VDD2.n8 B 0.011198f
C24 VDD2.n9 B 0.026469f
C25 VDD2.n10 B 0.011857f
C26 VDD2.n11 B 0.02084f
C27 VDD2.n12 B 0.011198f
C28 VDD2.n13 B 0.026469f
C29 VDD2.n14 B 0.011857f
C30 VDD2.n15 B 0.02084f
C31 VDD2.n16 B 0.011198f
C32 VDD2.n17 B 0.026469f
C33 VDD2.n18 B 0.011857f
C34 VDD2.n19 B 0.02084f
C35 VDD2.n20 B 0.011198f
C36 VDD2.n21 B 0.019852f
C37 VDD2.n22 B 0.015636f
C38 VDD2.t0 B 0.043479f
C39 VDD2.n23 B 0.123853f
C40 VDD2.n24 B 1.13525f
C41 VDD2.n25 B 0.011198f
C42 VDD2.n26 B 0.011857f
C43 VDD2.n27 B 0.026469f
C44 VDD2.n28 B 0.026469f
C45 VDD2.n29 B 0.011857f
C46 VDD2.n30 B 0.011198f
C47 VDD2.n31 B 0.02084f
C48 VDD2.n32 B 0.02084f
C49 VDD2.n33 B 0.011198f
C50 VDD2.n34 B 0.011857f
C51 VDD2.n35 B 0.026469f
C52 VDD2.n36 B 0.026469f
C53 VDD2.n37 B 0.011857f
C54 VDD2.n38 B 0.011198f
C55 VDD2.n39 B 0.02084f
C56 VDD2.n40 B 0.02084f
C57 VDD2.n41 B 0.011198f
C58 VDD2.n42 B 0.011857f
C59 VDD2.n43 B 0.026469f
C60 VDD2.n44 B 0.026469f
C61 VDD2.n45 B 0.011857f
C62 VDD2.n46 B 0.011198f
C63 VDD2.n47 B 0.02084f
C64 VDD2.n48 B 0.02084f
C65 VDD2.n49 B 0.011198f
C66 VDD2.n50 B 0.011857f
C67 VDD2.n51 B 0.026469f
C68 VDD2.n52 B 0.026469f
C69 VDD2.n53 B 0.011857f
C70 VDD2.n54 B 0.011198f
C71 VDD2.n55 B 0.02084f
C72 VDD2.n56 B 0.02084f
C73 VDD2.n57 B 0.011198f
C74 VDD2.n58 B 0.011857f
C75 VDD2.n59 B 0.026469f
C76 VDD2.n60 B 0.026469f
C77 VDD2.n61 B 0.011857f
C78 VDD2.n62 B 0.011198f
C79 VDD2.n63 B 0.02084f
C80 VDD2.n64 B 0.054149f
C81 VDD2.n65 B 0.011198f
C82 VDD2.n66 B 0.011857f
C83 VDD2.n67 B 0.054566f
C84 VDD2.n68 B 0.528626f
C85 VDD2.n69 B 0.011754f
C86 VDD2.n70 B 0.026469f
C87 VDD2.n71 B 0.011857f
C88 VDD2.n72 B 0.02084f
C89 VDD2.n73 B 0.011198f
C90 VDD2.n74 B 0.026469f
C91 VDD2.n75 B 0.011857f
C92 VDD2.n76 B 0.02084f
C93 VDD2.n77 B 0.011198f
C94 VDD2.n78 B 0.026469f
C95 VDD2.n79 B 0.011857f
C96 VDD2.n80 B 0.02084f
C97 VDD2.n81 B 0.011198f
C98 VDD2.n82 B 0.026469f
C99 VDD2.n83 B 0.011857f
C100 VDD2.n84 B 0.02084f
C101 VDD2.n85 B 0.011198f
C102 VDD2.n86 B 0.026469f
C103 VDD2.n87 B 0.011857f
C104 VDD2.n88 B 0.02084f
C105 VDD2.n89 B 0.011198f
C106 VDD2.n90 B 0.019852f
C107 VDD2.n91 B 0.015636f
C108 VDD2.t1 B 0.043479f
C109 VDD2.n92 B 0.123853f
C110 VDD2.n93 B 1.13525f
C111 VDD2.n94 B 0.011198f
C112 VDD2.n95 B 0.011857f
C113 VDD2.n96 B 0.026469f
C114 VDD2.n97 B 0.026469f
C115 VDD2.n98 B 0.011857f
C116 VDD2.n99 B 0.011198f
C117 VDD2.n100 B 0.02084f
C118 VDD2.n101 B 0.02084f
C119 VDD2.n102 B 0.011198f
C120 VDD2.n103 B 0.011857f
C121 VDD2.n104 B 0.026469f
C122 VDD2.n105 B 0.026469f
C123 VDD2.n106 B 0.011857f
C124 VDD2.n107 B 0.011198f
C125 VDD2.n108 B 0.02084f
C126 VDD2.n109 B 0.02084f
C127 VDD2.n110 B 0.011198f
C128 VDD2.n111 B 0.011857f
C129 VDD2.n112 B 0.026469f
C130 VDD2.n113 B 0.026469f
C131 VDD2.n114 B 0.011857f
C132 VDD2.n115 B 0.011198f
C133 VDD2.n116 B 0.02084f
C134 VDD2.n117 B 0.02084f
C135 VDD2.n118 B 0.011198f
C136 VDD2.n119 B 0.011857f
C137 VDD2.n120 B 0.026469f
C138 VDD2.n121 B 0.026469f
C139 VDD2.n122 B 0.011857f
C140 VDD2.n123 B 0.011198f
C141 VDD2.n124 B 0.02084f
C142 VDD2.n125 B 0.02084f
C143 VDD2.n126 B 0.011198f
C144 VDD2.n127 B 0.011857f
C145 VDD2.n128 B 0.026469f
C146 VDD2.n129 B 0.026469f
C147 VDD2.n130 B 0.011857f
C148 VDD2.n131 B 0.011198f
C149 VDD2.n132 B 0.02084f
C150 VDD2.n133 B 0.054149f
C151 VDD2.n134 B 0.011198f
C152 VDD2.n135 B 0.011857f
C153 VDD2.n136 B 0.054566f
C154 VDD2.n137 B 0.060433f
C155 VDD2.n138 B 2.32755f
C156 VN.t1 B 1.30157f
C157 VN.t0 B 1.42776f
C158 VDD1.n0 B 0.011642f
C159 VDD1.n1 B 0.026217f
C160 VDD1.n2 B 0.011744f
C161 VDD1.n3 B 0.020641f
C162 VDD1.n4 B 0.011092f
C163 VDD1.n5 B 0.026217f
C164 VDD1.n6 B 0.011744f
C165 VDD1.n7 B 0.020641f
C166 VDD1.n8 B 0.011092f
C167 VDD1.n9 B 0.026217f
C168 VDD1.n10 B 0.011744f
C169 VDD1.n11 B 0.020641f
C170 VDD1.n12 B 0.011092f
C171 VDD1.n13 B 0.026217f
C172 VDD1.n14 B 0.011744f
C173 VDD1.n15 B 0.020641f
C174 VDD1.n16 B 0.011092f
C175 VDD1.n17 B 0.026217f
C176 VDD1.n18 B 0.011744f
C177 VDD1.n19 B 0.020641f
C178 VDD1.n20 B 0.011092f
C179 VDD1.n21 B 0.019663f
C180 VDD1.n22 B 0.015487f
C181 VDD1.t1 B 0.043065f
C182 VDD1.n23 B 0.122673f
C183 VDD1.n24 B 1.12443f
C184 VDD1.n25 B 0.011092f
C185 VDD1.n26 B 0.011744f
C186 VDD1.n27 B 0.026217f
C187 VDD1.n28 B 0.026217f
C188 VDD1.n29 B 0.011744f
C189 VDD1.n30 B 0.011092f
C190 VDD1.n31 B 0.020641f
C191 VDD1.n32 B 0.020641f
C192 VDD1.n33 B 0.011092f
C193 VDD1.n34 B 0.011744f
C194 VDD1.n35 B 0.026217f
C195 VDD1.n36 B 0.026217f
C196 VDD1.n37 B 0.011744f
C197 VDD1.n38 B 0.011092f
C198 VDD1.n39 B 0.020641f
C199 VDD1.n40 B 0.020641f
C200 VDD1.n41 B 0.011092f
C201 VDD1.n42 B 0.011744f
C202 VDD1.n43 B 0.026217f
C203 VDD1.n44 B 0.026217f
C204 VDD1.n45 B 0.011744f
C205 VDD1.n46 B 0.011092f
C206 VDD1.n47 B 0.020641f
C207 VDD1.n48 B 0.020641f
C208 VDD1.n49 B 0.011092f
C209 VDD1.n50 B 0.011744f
C210 VDD1.n51 B 0.026217f
C211 VDD1.n52 B 0.026217f
C212 VDD1.n53 B 0.011744f
C213 VDD1.n54 B 0.011092f
C214 VDD1.n55 B 0.020641f
C215 VDD1.n56 B 0.020641f
C216 VDD1.n57 B 0.011092f
C217 VDD1.n58 B 0.011744f
C218 VDD1.n59 B 0.026217f
C219 VDD1.n60 B 0.026217f
C220 VDD1.n61 B 0.011744f
C221 VDD1.n62 B 0.011092f
C222 VDD1.n63 B 0.020641f
C223 VDD1.n64 B 0.053633f
C224 VDD1.n65 B 0.011092f
C225 VDD1.n66 B 0.011744f
C226 VDD1.n67 B 0.054046f
C227 VDD1.n68 B 0.060196f
C228 VDD1.n69 B 0.011642f
C229 VDD1.n70 B 0.026217f
C230 VDD1.n71 B 0.011744f
C231 VDD1.n72 B 0.020641f
C232 VDD1.n73 B 0.011092f
C233 VDD1.n74 B 0.026217f
C234 VDD1.n75 B 0.011744f
C235 VDD1.n76 B 0.020641f
C236 VDD1.n77 B 0.011092f
C237 VDD1.n78 B 0.026217f
C238 VDD1.n79 B 0.011744f
C239 VDD1.n80 B 0.020641f
C240 VDD1.n81 B 0.011092f
C241 VDD1.n82 B 0.026217f
C242 VDD1.n83 B 0.011744f
C243 VDD1.n84 B 0.020641f
C244 VDD1.n85 B 0.011092f
C245 VDD1.n86 B 0.026217f
C246 VDD1.n87 B 0.011744f
C247 VDD1.n88 B 0.020641f
C248 VDD1.n89 B 0.011092f
C249 VDD1.n90 B 0.019663f
C250 VDD1.n91 B 0.015487f
C251 VDD1.t0 B 0.043065f
C252 VDD1.n92 B 0.122673f
C253 VDD1.n93 B 1.12443f
C254 VDD1.n94 B 0.011092f
C255 VDD1.n95 B 0.011744f
C256 VDD1.n96 B 0.026217f
C257 VDD1.n97 B 0.026217f
C258 VDD1.n98 B 0.011744f
C259 VDD1.n99 B 0.011092f
C260 VDD1.n100 B 0.020641f
C261 VDD1.n101 B 0.020641f
C262 VDD1.n102 B 0.011092f
C263 VDD1.n103 B 0.011744f
C264 VDD1.n104 B 0.026217f
C265 VDD1.n105 B 0.026217f
C266 VDD1.n106 B 0.011744f
C267 VDD1.n107 B 0.011092f
C268 VDD1.n108 B 0.020641f
C269 VDD1.n109 B 0.020641f
C270 VDD1.n110 B 0.011092f
C271 VDD1.n111 B 0.011744f
C272 VDD1.n112 B 0.026217f
C273 VDD1.n113 B 0.026217f
C274 VDD1.n114 B 0.011744f
C275 VDD1.n115 B 0.011092f
C276 VDD1.n116 B 0.020641f
C277 VDD1.n117 B 0.020641f
C278 VDD1.n118 B 0.011092f
C279 VDD1.n119 B 0.011744f
C280 VDD1.n120 B 0.026217f
C281 VDD1.n121 B 0.026217f
C282 VDD1.n122 B 0.011744f
C283 VDD1.n123 B 0.011092f
C284 VDD1.n124 B 0.020641f
C285 VDD1.n125 B 0.020641f
C286 VDD1.n126 B 0.011092f
C287 VDD1.n127 B 0.011744f
C288 VDD1.n128 B 0.026217f
C289 VDD1.n129 B 0.026217f
C290 VDD1.n130 B 0.011744f
C291 VDD1.n131 B 0.011092f
C292 VDD1.n132 B 0.020641f
C293 VDD1.n133 B 0.053633f
C294 VDD1.n134 B 0.011092f
C295 VDD1.n135 B 0.011744f
C296 VDD1.n136 B 0.054046f
C297 VDD1.n137 B 0.55073f
C298 VTAIL.n0 B 0.00915f
C299 VTAIL.n1 B 0.020605f
C300 VTAIL.n2 B 0.00923f
C301 VTAIL.n3 B 0.016223f
C302 VTAIL.n4 B 0.008717f
C303 VTAIL.n5 B 0.020605f
C304 VTAIL.n6 B 0.00923f
C305 VTAIL.n7 B 0.016223f
C306 VTAIL.n8 B 0.008717f
C307 VTAIL.n9 B 0.020605f
C308 VTAIL.n10 B 0.00923f
C309 VTAIL.n11 B 0.016223f
C310 VTAIL.n12 B 0.008717f
C311 VTAIL.n13 B 0.020605f
C312 VTAIL.n14 B 0.00923f
C313 VTAIL.n15 B 0.016223f
C314 VTAIL.n16 B 0.008717f
C315 VTAIL.n17 B 0.020605f
C316 VTAIL.n18 B 0.00923f
C317 VTAIL.n19 B 0.016223f
C318 VTAIL.n20 B 0.008717f
C319 VTAIL.n21 B 0.015454f
C320 VTAIL.n22 B 0.012172f
C321 VTAIL.t2 B 0.033847f
C322 VTAIL.n23 B 0.096414f
C323 VTAIL.n24 B 0.883738f
C324 VTAIL.n25 B 0.008717f
C325 VTAIL.n26 B 0.00923f
C326 VTAIL.n27 B 0.020605f
C327 VTAIL.n28 B 0.020605f
C328 VTAIL.n29 B 0.00923f
C329 VTAIL.n30 B 0.008717f
C330 VTAIL.n31 B 0.016223f
C331 VTAIL.n32 B 0.016223f
C332 VTAIL.n33 B 0.008717f
C333 VTAIL.n34 B 0.00923f
C334 VTAIL.n35 B 0.020605f
C335 VTAIL.n36 B 0.020605f
C336 VTAIL.n37 B 0.00923f
C337 VTAIL.n38 B 0.008717f
C338 VTAIL.n39 B 0.016223f
C339 VTAIL.n40 B 0.016223f
C340 VTAIL.n41 B 0.008717f
C341 VTAIL.n42 B 0.00923f
C342 VTAIL.n43 B 0.020605f
C343 VTAIL.n44 B 0.020605f
C344 VTAIL.n45 B 0.00923f
C345 VTAIL.n46 B 0.008717f
C346 VTAIL.n47 B 0.016223f
C347 VTAIL.n48 B 0.016223f
C348 VTAIL.n49 B 0.008717f
C349 VTAIL.n50 B 0.00923f
C350 VTAIL.n51 B 0.020605f
C351 VTAIL.n52 B 0.020605f
C352 VTAIL.n53 B 0.00923f
C353 VTAIL.n54 B 0.008717f
C354 VTAIL.n55 B 0.016223f
C355 VTAIL.n56 B 0.016223f
C356 VTAIL.n57 B 0.008717f
C357 VTAIL.n58 B 0.00923f
C358 VTAIL.n59 B 0.020605f
C359 VTAIL.n60 B 0.020605f
C360 VTAIL.n61 B 0.00923f
C361 VTAIL.n62 B 0.008717f
C362 VTAIL.n63 B 0.016223f
C363 VTAIL.n64 B 0.042153f
C364 VTAIL.n65 B 0.008717f
C365 VTAIL.n66 B 0.00923f
C366 VTAIL.n67 B 0.042477f
C367 VTAIL.n68 B 0.035872f
C368 VTAIL.n69 B 0.94546f
C369 VTAIL.n70 B 0.00915f
C370 VTAIL.n71 B 0.020605f
C371 VTAIL.n72 B 0.00923f
C372 VTAIL.n73 B 0.016223f
C373 VTAIL.n74 B 0.008717f
C374 VTAIL.n75 B 0.020605f
C375 VTAIL.n76 B 0.00923f
C376 VTAIL.n77 B 0.016223f
C377 VTAIL.n78 B 0.008717f
C378 VTAIL.n79 B 0.020605f
C379 VTAIL.n80 B 0.00923f
C380 VTAIL.n81 B 0.016223f
C381 VTAIL.n82 B 0.008717f
C382 VTAIL.n83 B 0.020605f
C383 VTAIL.n84 B 0.00923f
C384 VTAIL.n85 B 0.016223f
C385 VTAIL.n86 B 0.008717f
C386 VTAIL.n87 B 0.020605f
C387 VTAIL.n88 B 0.00923f
C388 VTAIL.n89 B 0.016223f
C389 VTAIL.n90 B 0.008717f
C390 VTAIL.n91 B 0.015454f
C391 VTAIL.n92 B 0.012172f
C392 VTAIL.t0 B 0.033847f
C393 VTAIL.n93 B 0.096414f
C394 VTAIL.n94 B 0.883738f
C395 VTAIL.n95 B 0.008717f
C396 VTAIL.n96 B 0.00923f
C397 VTAIL.n97 B 0.020605f
C398 VTAIL.n98 B 0.020605f
C399 VTAIL.n99 B 0.00923f
C400 VTAIL.n100 B 0.008717f
C401 VTAIL.n101 B 0.016223f
C402 VTAIL.n102 B 0.016223f
C403 VTAIL.n103 B 0.008717f
C404 VTAIL.n104 B 0.00923f
C405 VTAIL.n105 B 0.020605f
C406 VTAIL.n106 B 0.020605f
C407 VTAIL.n107 B 0.00923f
C408 VTAIL.n108 B 0.008717f
C409 VTAIL.n109 B 0.016223f
C410 VTAIL.n110 B 0.016223f
C411 VTAIL.n111 B 0.008717f
C412 VTAIL.n112 B 0.00923f
C413 VTAIL.n113 B 0.020605f
C414 VTAIL.n114 B 0.020605f
C415 VTAIL.n115 B 0.00923f
C416 VTAIL.n116 B 0.008717f
C417 VTAIL.n117 B 0.016223f
C418 VTAIL.n118 B 0.016223f
C419 VTAIL.n119 B 0.008717f
C420 VTAIL.n120 B 0.00923f
C421 VTAIL.n121 B 0.020605f
C422 VTAIL.n122 B 0.020605f
C423 VTAIL.n123 B 0.00923f
C424 VTAIL.n124 B 0.008717f
C425 VTAIL.n125 B 0.016223f
C426 VTAIL.n126 B 0.016223f
C427 VTAIL.n127 B 0.008717f
C428 VTAIL.n128 B 0.00923f
C429 VTAIL.n129 B 0.020605f
C430 VTAIL.n130 B 0.020605f
C431 VTAIL.n131 B 0.00923f
C432 VTAIL.n132 B 0.008717f
C433 VTAIL.n133 B 0.016223f
C434 VTAIL.n134 B 0.042153f
C435 VTAIL.n135 B 0.008717f
C436 VTAIL.n136 B 0.00923f
C437 VTAIL.n137 B 0.042477f
C438 VTAIL.n138 B 0.035872f
C439 VTAIL.n139 B 0.954472f
C440 VTAIL.n140 B 0.00915f
C441 VTAIL.n141 B 0.020605f
C442 VTAIL.n142 B 0.00923f
C443 VTAIL.n143 B 0.016223f
C444 VTAIL.n144 B 0.008717f
C445 VTAIL.n145 B 0.020605f
C446 VTAIL.n146 B 0.00923f
C447 VTAIL.n147 B 0.016223f
C448 VTAIL.n148 B 0.008717f
C449 VTAIL.n149 B 0.020605f
C450 VTAIL.n150 B 0.00923f
C451 VTAIL.n151 B 0.016223f
C452 VTAIL.n152 B 0.008717f
C453 VTAIL.n153 B 0.020605f
C454 VTAIL.n154 B 0.00923f
C455 VTAIL.n155 B 0.016223f
C456 VTAIL.n156 B 0.008717f
C457 VTAIL.n157 B 0.020605f
C458 VTAIL.n158 B 0.00923f
C459 VTAIL.n159 B 0.016223f
C460 VTAIL.n160 B 0.008717f
C461 VTAIL.n161 B 0.015454f
C462 VTAIL.n162 B 0.012172f
C463 VTAIL.t3 B 0.033847f
C464 VTAIL.n163 B 0.096414f
C465 VTAIL.n164 B 0.883738f
C466 VTAIL.n165 B 0.008717f
C467 VTAIL.n166 B 0.00923f
C468 VTAIL.n167 B 0.020605f
C469 VTAIL.n168 B 0.020605f
C470 VTAIL.n169 B 0.00923f
C471 VTAIL.n170 B 0.008717f
C472 VTAIL.n171 B 0.016223f
C473 VTAIL.n172 B 0.016223f
C474 VTAIL.n173 B 0.008717f
C475 VTAIL.n174 B 0.00923f
C476 VTAIL.n175 B 0.020605f
C477 VTAIL.n176 B 0.020605f
C478 VTAIL.n177 B 0.00923f
C479 VTAIL.n178 B 0.008717f
C480 VTAIL.n179 B 0.016223f
C481 VTAIL.n180 B 0.016223f
C482 VTAIL.n181 B 0.008717f
C483 VTAIL.n182 B 0.00923f
C484 VTAIL.n183 B 0.020605f
C485 VTAIL.n184 B 0.020605f
C486 VTAIL.n185 B 0.00923f
C487 VTAIL.n186 B 0.008717f
C488 VTAIL.n187 B 0.016223f
C489 VTAIL.n188 B 0.016223f
C490 VTAIL.n189 B 0.008717f
C491 VTAIL.n190 B 0.00923f
C492 VTAIL.n191 B 0.020605f
C493 VTAIL.n192 B 0.020605f
C494 VTAIL.n193 B 0.00923f
C495 VTAIL.n194 B 0.008717f
C496 VTAIL.n195 B 0.016223f
C497 VTAIL.n196 B 0.016223f
C498 VTAIL.n197 B 0.008717f
C499 VTAIL.n198 B 0.00923f
C500 VTAIL.n199 B 0.020605f
C501 VTAIL.n200 B 0.020605f
C502 VTAIL.n201 B 0.00923f
C503 VTAIL.n202 B 0.008717f
C504 VTAIL.n203 B 0.016223f
C505 VTAIL.n204 B 0.042153f
C506 VTAIL.n205 B 0.008717f
C507 VTAIL.n206 B 0.00923f
C508 VTAIL.n207 B 0.042477f
C509 VTAIL.n208 B 0.035872f
C510 VTAIL.n209 B 0.906254f
C511 VTAIL.n210 B 0.00915f
C512 VTAIL.n211 B 0.020605f
C513 VTAIL.n212 B 0.00923f
C514 VTAIL.n213 B 0.016223f
C515 VTAIL.n214 B 0.008717f
C516 VTAIL.n215 B 0.020605f
C517 VTAIL.n216 B 0.00923f
C518 VTAIL.n217 B 0.016223f
C519 VTAIL.n218 B 0.008717f
C520 VTAIL.n219 B 0.020605f
C521 VTAIL.n220 B 0.00923f
C522 VTAIL.n221 B 0.016223f
C523 VTAIL.n222 B 0.008717f
C524 VTAIL.n223 B 0.020605f
C525 VTAIL.n224 B 0.00923f
C526 VTAIL.n225 B 0.016223f
C527 VTAIL.n226 B 0.008717f
C528 VTAIL.n227 B 0.020605f
C529 VTAIL.n228 B 0.00923f
C530 VTAIL.n229 B 0.016223f
C531 VTAIL.n230 B 0.008717f
C532 VTAIL.n231 B 0.015454f
C533 VTAIL.n232 B 0.012172f
C534 VTAIL.t1 B 0.033847f
C535 VTAIL.n233 B 0.096414f
C536 VTAIL.n234 B 0.883738f
C537 VTAIL.n235 B 0.008717f
C538 VTAIL.n236 B 0.00923f
C539 VTAIL.n237 B 0.020605f
C540 VTAIL.n238 B 0.020605f
C541 VTAIL.n239 B 0.00923f
C542 VTAIL.n240 B 0.008717f
C543 VTAIL.n241 B 0.016223f
C544 VTAIL.n242 B 0.016223f
C545 VTAIL.n243 B 0.008717f
C546 VTAIL.n244 B 0.00923f
C547 VTAIL.n245 B 0.020605f
C548 VTAIL.n246 B 0.020605f
C549 VTAIL.n247 B 0.00923f
C550 VTAIL.n248 B 0.008717f
C551 VTAIL.n249 B 0.016223f
C552 VTAIL.n250 B 0.016223f
C553 VTAIL.n251 B 0.008717f
C554 VTAIL.n252 B 0.00923f
C555 VTAIL.n253 B 0.020605f
C556 VTAIL.n254 B 0.020605f
C557 VTAIL.n255 B 0.00923f
C558 VTAIL.n256 B 0.008717f
C559 VTAIL.n257 B 0.016223f
C560 VTAIL.n258 B 0.016223f
C561 VTAIL.n259 B 0.008717f
C562 VTAIL.n260 B 0.00923f
C563 VTAIL.n261 B 0.020605f
C564 VTAIL.n262 B 0.020605f
C565 VTAIL.n263 B 0.00923f
C566 VTAIL.n264 B 0.008717f
C567 VTAIL.n265 B 0.016223f
C568 VTAIL.n266 B 0.016223f
C569 VTAIL.n267 B 0.008717f
C570 VTAIL.n268 B 0.00923f
C571 VTAIL.n269 B 0.020605f
C572 VTAIL.n270 B 0.020605f
C573 VTAIL.n271 B 0.00923f
C574 VTAIL.n272 B 0.008717f
C575 VTAIL.n273 B 0.016223f
C576 VTAIL.n274 B 0.042153f
C577 VTAIL.n275 B 0.008717f
C578 VTAIL.n276 B 0.00923f
C579 VTAIL.n277 B 0.042477f
C580 VTAIL.n278 B 0.035872f
C581 VTAIL.n279 B 0.866598f
C582 VP.t0 B 1.45919f
C583 VP.t1 B 1.33287f
C584 VP.n0 B 4.09105f
.ends

