* NGSPICE file created from diff_pair_sample_0874.ext - technology: sky130A

.subckt diff_pair_sample_0874 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=2.36775 ps=14.68 w=14.35 l=1.34
X1 VDD1.t0 VP.t1 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=2.36775 ps=14.68 w=14.35 l=1.34
X2 VTAIL.t13 VP.t2 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=5.5965 pd=29.48 as=2.36775 ps=14.68 w=14.35 l=1.34
X3 VTAIL.t2 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=5.5965 pd=29.48 as=2.36775 ps=14.68 w=14.35 l=1.34
X4 VDD2.t6 VN.t1 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=5.5965 ps=29.48 w=14.35 l=1.34
X5 VTAIL.t12 VP.t3 VDD1.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=2.36775 ps=14.68 w=14.35 l=1.34
X6 VTAIL.t3 VN.t2 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=2.36775 ps=14.68 w=14.35 l=1.34
X7 VDD1.t2 VP.t4 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=5.5965 ps=29.48 w=14.35 l=1.34
X8 VDD1.t3 VP.t5 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=5.5965 ps=29.48 w=14.35 l=1.34
X9 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=5.5965 pd=29.48 as=0 ps=0 w=14.35 l=1.34
X10 VDD2.t4 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=2.36775 ps=14.68 w=14.35 l=1.34
X11 VTAIL.t9 VP.t6 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=5.5965 pd=29.48 as=2.36775 ps=14.68 w=14.35 l=1.34
X12 VDD2.t3 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=5.5965 ps=29.48 w=14.35 l=1.34
X13 VTAIL.t5 VN.t5 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=2.36775 ps=14.68 w=14.35 l=1.34
X14 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=5.5965 pd=29.48 as=0 ps=0 w=14.35 l=1.34
X15 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.5965 pd=29.48 as=0 ps=0 w=14.35 l=1.34
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.5965 pd=29.48 as=0 ps=0 w=14.35 l=1.34
X17 VTAIL.t0 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=5.5965 pd=29.48 as=2.36775 ps=14.68 w=14.35 l=1.34
X18 VDD2.t0 VN.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=2.36775 ps=14.68 w=14.35 l=1.34
X19 VDD1.t1 VP.t7 VTAIL.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.36775 pd=14.68 as=2.36775 ps=14.68 w=14.35 l=1.34
R0 VP.n11 VP.t2 287.204
R1 VP.n5 VP.t6 258.087
R2 VP.n29 VP.t7 258.087
R3 VP.n36 VP.t3 258.087
R4 VP.n43 VP.t4 258.087
R5 VP.n23 VP.t5 258.087
R6 VP.n16 VP.t0 258.087
R7 VP.n10 VP.t1 258.087
R8 VP.n25 VP.n5 173.29
R9 VP.n44 VP.n43 173.29
R10 VP.n24 VP.n23 173.29
R11 VP.n12 VP.n9 161.3
R12 VP.n14 VP.n13 161.3
R13 VP.n15 VP.n8 161.3
R14 VP.n18 VP.n17 161.3
R15 VP.n19 VP.n7 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n6 161.3
R18 VP.n42 VP.n0 161.3
R19 VP.n41 VP.n40 161.3
R20 VP.n39 VP.n1 161.3
R21 VP.n38 VP.n37 161.3
R22 VP.n35 VP.n2 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n32 VP.n3 161.3
R25 VP.n31 VP.n30 161.3
R26 VP.n28 VP.n4 161.3
R27 VP.n27 VP.n26 161.3
R28 VP.n11 VP.n10 61.1116
R29 VP.n35 VP.n34 56.5193
R30 VP.n15 VP.n14 56.5193
R31 VP.n30 VP.n28 48.2635
R32 VP.n41 VP.n1 48.2635
R33 VP.n21 VP.n7 48.2635
R34 VP.n25 VP.n24 46.705
R35 VP.n28 VP.n27 32.7233
R36 VP.n42 VP.n41 32.7233
R37 VP.n22 VP.n21 32.7233
R38 VP.n12 VP.n11 27.209
R39 VP.n34 VP.n3 24.4675
R40 VP.n37 VP.n35 24.4675
R41 VP.n17 VP.n15 24.4675
R42 VP.n14 VP.n9 24.4675
R43 VP.n30 VP.n29 20.3081
R44 VP.n36 VP.n1 20.3081
R45 VP.n16 VP.n7 20.3081
R46 VP.n27 VP.n5 12.4787
R47 VP.n43 VP.n42 12.4787
R48 VP.n23 VP.n22 12.4787
R49 VP.n29 VP.n3 4.15989
R50 VP.n37 VP.n36 4.15989
R51 VP.n17 VP.n16 4.15989
R52 VP.n10 VP.n9 4.15989
R53 VP.n13 VP.n12 0.189894
R54 VP.n13 VP.n8 0.189894
R55 VP.n18 VP.n8 0.189894
R56 VP.n19 VP.n18 0.189894
R57 VP.n20 VP.n19 0.189894
R58 VP.n20 VP.n6 0.189894
R59 VP.n24 VP.n6 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n4 0.189894
R62 VP.n31 VP.n4 0.189894
R63 VP.n32 VP.n31 0.189894
R64 VP.n33 VP.n32 0.189894
R65 VP.n33 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP.n44 VP.n0 0.189894
R71 VP VP.n44 0.0516364
R72 VDD1 VDD1.n0 63.1015
R73 VDD1.n3 VDD1.n2 62.9877
R74 VDD1.n3 VDD1.n1 62.9877
R75 VDD1.n5 VDD1.n4 62.3233
R76 VDD1.n5 VDD1.n3 43.1474
R77 VDD1.n4 VDD1.t7 1.38029
R78 VDD1.n4 VDD1.t3 1.38029
R79 VDD1.n0 VDD1.t4 1.38029
R80 VDD1.n0 VDD1.t0 1.38029
R81 VDD1.n2 VDD1.t6 1.38029
R82 VDD1.n2 VDD1.t2 1.38029
R83 VDD1.n1 VDD1.t5 1.38029
R84 VDD1.n1 VDD1.t1 1.38029
R85 VDD1 VDD1.n5 0.662138
R86 VTAIL.n11 VTAIL.t13 47.0244
R87 VTAIL.n10 VTAIL.t4 47.0244
R88 VTAIL.n7 VTAIL.t2 47.0244
R89 VTAIL.n15 VTAIL.t6 47.0243
R90 VTAIL.n2 VTAIL.t0 47.0243
R91 VTAIL.n3 VTAIL.t11 47.0243
R92 VTAIL.n6 VTAIL.t9 47.0243
R93 VTAIL.n14 VTAIL.t10 47.0243
R94 VTAIL.n13 VTAIL.n12 45.6447
R95 VTAIL.n9 VTAIL.n8 45.6447
R96 VTAIL.n1 VTAIL.n0 45.6444
R97 VTAIL.n5 VTAIL.n4 45.6444
R98 VTAIL.n15 VTAIL.n14 26.1772
R99 VTAIL.n7 VTAIL.n6 26.1772
R100 VTAIL.n9 VTAIL.n7 1.44016
R101 VTAIL.n10 VTAIL.n9 1.44016
R102 VTAIL.n13 VTAIL.n11 1.44016
R103 VTAIL.n14 VTAIL.n13 1.44016
R104 VTAIL.n6 VTAIL.n5 1.44016
R105 VTAIL.n5 VTAIL.n3 1.44016
R106 VTAIL.n2 VTAIL.n1 1.44016
R107 VTAIL VTAIL.n15 1.38197
R108 VTAIL.n0 VTAIL.t1 1.38029
R109 VTAIL.n0 VTAIL.t3 1.38029
R110 VTAIL.n4 VTAIL.t8 1.38029
R111 VTAIL.n4 VTAIL.t12 1.38029
R112 VTAIL.n12 VTAIL.t14 1.38029
R113 VTAIL.n12 VTAIL.t15 1.38029
R114 VTAIL.n8 VTAIL.t7 1.38029
R115 VTAIL.n8 VTAIL.t5 1.38029
R116 VTAIL.n11 VTAIL.n10 0.470328
R117 VTAIL.n3 VTAIL.n2 0.470328
R118 VTAIL VTAIL.n1 0.0586897
R119 B.n807 B.n806 585
R120 B.n808 B.n807 585
R121 B.n330 B.n115 585
R122 B.n329 B.n328 585
R123 B.n327 B.n326 585
R124 B.n325 B.n324 585
R125 B.n323 B.n322 585
R126 B.n321 B.n320 585
R127 B.n319 B.n318 585
R128 B.n317 B.n316 585
R129 B.n315 B.n314 585
R130 B.n313 B.n312 585
R131 B.n311 B.n310 585
R132 B.n309 B.n308 585
R133 B.n307 B.n306 585
R134 B.n305 B.n304 585
R135 B.n303 B.n302 585
R136 B.n301 B.n300 585
R137 B.n299 B.n298 585
R138 B.n297 B.n296 585
R139 B.n295 B.n294 585
R140 B.n293 B.n292 585
R141 B.n291 B.n290 585
R142 B.n289 B.n288 585
R143 B.n287 B.n286 585
R144 B.n285 B.n284 585
R145 B.n283 B.n282 585
R146 B.n281 B.n280 585
R147 B.n279 B.n278 585
R148 B.n277 B.n276 585
R149 B.n275 B.n274 585
R150 B.n273 B.n272 585
R151 B.n271 B.n270 585
R152 B.n269 B.n268 585
R153 B.n267 B.n266 585
R154 B.n265 B.n264 585
R155 B.n263 B.n262 585
R156 B.n261 B.n260 585
R157 B.n259 B.n258 585
R158 B.n257 B.n256 585
R159 B.n255 B.n254 585
R160 B.n253 B.n252 585
R161 B.n251 B.n250 585
R162 B.n249 B.n248 585
R163 B.n247 B.n246 585
R164 B.n245 B.n244 585
R165 B.n243 B.n242 585
R166 B.n241 B.n240 585
R167 B.n239 B.n238 585
R168 B.n237 B.n236 585
R169 B.n235 B.n234 585
R170 B.n233 B.n232 585
R171 B.n231 B.n230 585
R172 B.n229 B.n228 585
R173 B.n227 B.n226 585
R174 B.n225 B.n224 585
R175 B.n223 B.n222 585
R176 B.n221 B.n220 585
R177 B.n219 B.n218 585
R178 B.n216 B.n215 585
R179 B.n214 B.n213 585
R180 B.n212 B.n211 585
R181 B.n210 B.n209 585
R182 B.n208 B.n207 585
R183 B.n206 B.n205 585
R184 B.n204 B.n203 585
R185 B.n202 B.n201 585
R186 B.n200 B.n199 585
R187 B.n198 B.n197 585
R188 B.n196 B.n195 585
R189 B.n194 B.n193 585
R190 B.n192 B.n191 585
R191 B.n190 B.n189 585
R192 B.n188 B.n187 585
R193 B.n186 B.n185 585
R194 B.n184 B.n183 585
R195 B.n182 B.n181 585
R196 B.n180 B.n179 585
R197 B.n178 B.n177 585
R198 B.n176 B.n175 585
R199 B.n174 B.n173 585
R200 B.n172 B.n171 585
R201 B.n170 B.n169 585
R202 B.n168 B.n167 585
R203 B.n166 B.n165 585
R204 B.n164 B.n163 585
R205 B.n162 B.n161 585
R206 B.n160 B.n159 585
R207 B.n158 B.n157 585
R208 B.n156 B.n155 585
R209 B.n154 B.n153 585
R210 B.n152 B.n151 585
R211 B.n150 B.n149 585
R212 B.n148 B.n147 585
R213 B.n146 B.n145 585
R214 B.n144 B.n143 585
R215 B.n142 B.n141 585
R216 B.n140 B.n139 585
R217 B.n138 B.n137 585
R218 B.n136 B.n135 585
R219 B.n134 B.n133 585
R220 B.n132 B.n131 585
R221 B.n130 B.n129 585
R222 B.n128 B.n127 585
R223 B.n126 B.n125 585
R224 B.n124 B.n123 585
R225 B.n122 B.n121 585
R226 B.n60 B.n59 585
R227 B.n805 B.n61 585
R228 B.n809 B.n61 585
R229 B.n804 B.n803 585
R230 B.n803 B.n57 585
R231 B.n802 B.n56 585
R232 B.n815 B.n56 585
R233 B.n801 B.n55 585
R234 B.n816 B.n55 585
R235 B.n800 B.n54 585
R236 B.n817 B.n54 585
R237 B.n799 B.n798 585
R238 B.n798 B.n53 585
R239 B.n797 B.n49 585
R240 B.n823 B.n49 585
R241 B.n796 B.n48 585
R242 B.n824 B.n48 585
R243 B.n795 B.n47 585
R244 B.n825 B.n47 585
R245 B.n794 B.n793 585
R246 B.n793 B.n43 585
R247 B.n792 B.n42 585
R248 B.n831 B.n42 585
R249 B.n791 B.n41 585
R250 B.n832 B.n41 585
R251 B.n790 B.n40 585
R252 B.n833 B.n40 585
R253 B.n789 B.n788 585
R254 B.n788 B.n39 585
R255 B.n787 B.n35 585
R256 B.n839 B.n35 585
R257 B.n786 B.n34 585
R258 B.n840 B.n34 585
R259 B.n785 B.n33 585
R260 B.n841 B.n33 585
R261 B.n784 B.n783 585
R262 B.n783 B.n29 585
R263 B.n782 B.n28 585
R264 B.n847 B.n28 585
R265 B.n781 B.n27 585
R266 B.n848 B.n27 585
R267 B.n780 B.n26 585
R268 B.n849 B.n26 585
R269 B.n779 B.n778 585
R270 B.n778 B.n22 585
R271 B.n777 B.n21 585
R272 B.n855 B.n21 585
R273 B.n776 B.n20 585
R274 B.n856 B.n20 585
R275 B.n775 B.n19 585
R276 B.n857 B.n19 585
R277 B.n774 B.n773 585
R278 B.n773 B.n15 585
R279 B.n772 B.n14 585
R280 B.n863 B.n14 585
R281 B.n771 B.n13 585
R282 B.n864 B.n13 585
R283 B.n770 B.n12 585
R284 B.n865 B.n12 585
R285 B.n769 B.n768 585
R286 B.n768 B.n767 585
R287 B.n766 B.n765 585
R288 B.n766 B.n8 585
R289 B.n764 B.n7 585
R290 B.n872 B.n7 585
R291 B.n763 B.n6 585
R292 B.n873 B.n6 585
R293 B.n762 B.n5 585
R294 B.n874 B.n5 585
R295 B.n761 B.n760 585
R296 B.n760 B.n4 585
R297 B.n759 B.n331 585
R298 B.n759 B.n758 585
R299 B.n749 B.n332 585
R300 B.n333 B.n332 585
R301 B.n751 B.n750 585
R302 B.n752 B.n751 585
R303 B.n748 B.n338 585
R304 B.n338 B.n337 585
R305 B.n747 B.n746 585
R306 B.n746 B.n745 585
R307 B.n340 B.n339 585
R308 B.n341 B.n340 585
R309 B.n738 B.n737 585
R310 B.n739 B.n738 585
R311 B.n736 B.n345 585
R312 B.n349 B.n345 585
R313 B.n735 B.n734 585
R314 B.n734 B.n733 585
R315 B.n347 B.n346 585
R316 B.n348 B.n347 585
R317 B.n726 B.n725 585
R318 B.n727 B.n726 585
R319 B.n724 B.n354 585
R320 B.n354 B.n353 585
R321 B.n723 B.n722 585
R322 B.n722 B.n721 585
R323 B.n356 B.n355 585
R324 B.n357 B.n356 585
R325 B.n714 B.n713 585
R326 B.n715 B.n714 585
R327 B.n712 B.n362 585
R328 B.n362 B.n361 585
R329 B.n711 B.n710 585
R330 B.n710 B.n709 585
R331 B.n364 B.n363 585
R332 B.n702 B.n364 585
R333 B.n701 B.n700 585
R334 B.n703 B.n701 585
R335 B.n699 B.n369 585
R336 B.n369 B.n368 585
R337 B.n698 B.n697 585
R338 B.n697 B.n696 585
R339 B.n371 B.n370 585
R340 B.n372 B.n371 585
R341 B.n689 B.n688 585
R342 B.n690 B.n689 585
R343 B.n687 B.n377 585
R344 B.n377 B.n376 585
R345 B.n686 B.n685 585
R346 B.n685 B.n684 585
R347 B.n379 B.n378 585
R348 B.n677 B.n379 585
R349 B.n676 B.n675 585
R350 B.n678 B.n676 585
R351 B.n674 B.n384 585
R352 B.n384 B.n383 585
R353 B.n673 B.n672 585
R354 B.n672 B.n671 585
R355 B.n386 B.n385 585
R356 B.n387 B.n386 585
R357 B.n664 B.n663 585
R358 B.n665 B.n664 585
R359 B.n390 B.n389 585
R360 B.n452 B.n451 585
R361 B.n453 B.n449 585
R362 B.n449 B.n391 585
R363 B.n455 B.n454 585
R364 B.n457 B.n448 585
R365 B.n460 B.n459 585
R366 B.n461 B.n447 585
R367 B.n463 B.n462 585
R368 B.n465 B.n446 585
R369 B.n468 B.n467 585
R370 B.n469 B.n445 585
R371 B.n471 B.n470 585
R372 B.n473 B.n444 585
R373 B.n476 B.n475 585
R374 B.n477 B.n443 585
R375 B.n479 B.n478 585
R376 B.n481 B.n442 585
R377 B.n484 B.n483 585
R378 B.n485 B.n441 585
R379 B.n487 B.n486 585
R380 B.n489 B.n440 585
R381 B.n492 B.n491 585
R382 B.n493 B.n439 585
R383 B.n495 B.n494 585
R384 B.n497 B.n438 585
R385 B.n500 B.n499 585
R386 B.n501 B.n437 585
R387 B.n503 B.n502 585
R388 B.n505 B.n436 585
R389 B.n508 B.n507 585
R390 B.n509 B.n435 585
R391 B.n511 B.n510 585
R392 B.n513 B.n434 585
R393 B.n516 B.n515 585
R394 B.n517 B.n433 585
R395 B.n519 B.n518 585
R396 B.n521 B.n432 585
R397 B.n524 B.n523 585
R398 B.n525 B.n431 585
R399 B.n527 B.n526 585
R400 B.n529 B.n430 585
R401 B.n532 B.n531 585
R402 B.n533 B.n429 585
R403 B.n535 B.n534 585
R404 B.n537 B.n428 585
R405 B.n540 B.n539 585
R406 B.n541 B.n427 585
R407 B.n543 B.n542 585
R408 B.n545 B.n426 585
R409 B.n548 B.n547 585
R410 B.n549 B.n422 585
R411 B.n551 B.n550 585
R412 B.n553 B.n421 585
R413 B.n556 B.n555 585
R414 B.n557 B.n420 585
R415 B.n559 B.n558 585
R416 B.n561 B.n419 585
R417 B.n564 B.n563 585
R418 B.n566 B.n416 585
R419 B.n568 B.n567 585
R420 B.n570 B.n415 585
R421 B.n573 B.n572 585
R422 B.n574 B.n414 585
R423 B.n576 B.n575 585
R424 B.n578 B.n413 585
R425 B.n581 B.n580 585
R426 B.n582 B.n412 585
R427 B.n584 B.n583 585
R428 B.n586 B.n411 585
R429 B.n589 B.n588 585
R430 B.n590 B.n410 585
R431 B.n592 B.n591 585
R432 B.n594 B.n409 585
R433 B.n597 B.n596 585
R434 B.n598 B.n408 585
R435 B.n600 B.n599 585
R436 B.n602 B.n407 585
R437 B.n605 B.n604 585
R438 B.n606 B.n406 585
R439 B.n608 B.n607 585
R440 B.n610 B.n405 585
R441 B.n613 B.n612 585
R442 B.n614 B.n404 585
R443 B.n616 B.n615 585
R444 B.n618 B.n403 585
R445 B.n621 B.n620 585
R446 B.n622 B.n402 585
R447 B.n624 B.n623 585
R448 B.n626 B.n401 585
R449 B.n629 B.n628 585
R450 B.n630 B.n400 585
R451 B.n632 B.n631 585
R452 B.n634 B.n399 585
R453 B.n637 B.n636 585
R454 B.n638 B.n398 585
R455 B.n640 B.n639 585
R456 B.n642 B.n397 585
R457 B.n645 B.n644 585
R458 B.n646 B.n396 585
R459 B.n648 B.n647 585
R460 B.n650 B.n395 585
R461 B.n653 B.n652 585
R462 B.n654 B.n394 585
R463 B.n656 B.n655 585
R464 B.n658 B.n393 585
R465 B.n661 B.n660 585
R466 B.n662 B.n392 585
R467 B.n667 B.n666 585
R468 B.n666 B.n665 585
R469 B.n668 B.n388 585
R470 B.n388 B.n387 585
R471 B.n670 B.n669 585
R472 B.n671 B.n670 585
R473 B.n382 B.n381 585
R474 B.n383 B.n382 585
R475 B.n680 B.n679 585
R476 B.n679 B.n678 585
R477 B.n681 B.n380 585
R478 B.n677 B.n380 585
R479 B.n683 B.n682 585
R480 B.n684 B.n683 585
R481 B.n375 B.n374 585
R482 B.n376 B.n375 585
R483 B.n692 B.n691 585
R484 B.n691 B.n690 585
R485 B.n693 B.n373 585
R486 B.n373 B.n372 585
R487 B.n695 B.n694 585
R488 B.n696 B.n695 585
R489 B.n367 B.n366 585
R490 B.n368 B.n367 585
R491 B.n705 B.n704 585
R492 B.n704 B.n703 585
R493 B.n706 B.n365 585
R494 B.n702 B.n365 585
R495 B.n708 B.n707 585
R496 B.n709 B.n708 585
R497 B.n360 B.n359 585
R498 B.n361 B.n360 585
R499 B.n717 B.n716 585
R500 B.n716 B.n715 585
R501 B.n718 B.n358 585
R502 B.n358 B.n357 585
R503 B.n720 B.n719 585
R504 B.n721 B.n720 585
R505 B.n352 B.n351 585
R506 B.n353 B.n352 585
R507 B.n729 B.n728 585
R508 B.n728 B.n727 585
R509 B.n730 B.n350 585
R510 B.n350 B.n348 585
R511 B.n732 B.n731 585
R512 B.n733 B.n732 585
R513 B.n344 B.n343 585
R514 B.n349 B.n344 585
R515 B.n741 B.n740 585
R516 B.n740 B.n739 585
R517 B.n742 B.n342 585
R518 B.n342 B.n341 585
R519 B.n744 B.n743 585
R520 B.n745 B.n744 585
R521 B.n336 B.n335 585
R522 B.n337 B.n336 585
R523 B.n754 B.n753 585
R524 B.n753 B.n752 585
R525 B.n755 B.n334 585
R526 B.n334 B.n333 585
R527 B.n757 B.n756 585
R528 B.n758 B.n757 585
R529 B.n3 B.n0 585
R530 B.n4 B.n3 585
R531 B.n871 B.n1 585
R532 B.n872 B.n871 585
R533 B.n870 B.n869 585
R534 B.n870 B.n8 585
R535 B.n868 B.n9 585
R536 B.n767 B.n9 585
R537 B.n867 B.n866 585
R538 B.n866 B.n865 585
R539 B.n11 B.n10 585
R540 B.n864 B.n11 585
R541 B.n862 B.n861 585
R542 B.n863 B.n862 585
R543 B.n860 B.n16 585
R544 B.n16 B.n15 585
R545 B.n859 B.n858 585
R546 B.n858 B.n857 585
R547 B.n18 B.n17 585
R548 B.n856 B.n18 585
R549 B.n854 B.n853 585
R550 B.n855 B.n854 585
R551 B.n852 B.n23 585
R552 B.n23 B.n22 585
R553 B.n851 B.n850 585
R554 B.n850 B.n849 585
R555 B.n25 B.n24 585
R556 B.n848 B.n25 585
R557 B.n846 B.n845 585
R558 B.n847 B.n846 585
R559 B.n844 B.n30 585
R560 B.n30 B.n29 585
R561 B.n843 B.n842 585
R562 B.n842 B.n841 585
R563 B.n32 B.n31 585
R564 B.n840 B.n32 585
R565 B.n838 B.n837 585
R566 B.n839 B.n838 585
R567 B.n836 B.n36 585
R568 B.n39 B.n36 585
R569 B.n835 B.n834 585
R570 B.n834 B.n833 585
R571 B.n38 B.n37 585
R572 B.n832 B.n38 585
R573 B.n830 B.n829 585
R574 B.n831 B.n830 585
R575 B.n828 B.n44 585
R576 B.n44 B.n43 585
R577 B.n827 B.n826 585
R578 B.n826 B.n825 585
R579 B.n46 B.n45 585
R580 B.n824 B.n46 585
R581 B.n822 B.n821 585
R582 B.n823 B.n822 585
R583 B.n820 B.n50 585
R584 B.n53 B.n50 585
R585 B.n819 B.n818 585
R586 B.n818 B.n817 585
R587 B.n52 B.n51 585
R588 B.n816 B.n52 585
R589 B.n814 B.n813 585
R590 B.n815 B.n814 585
R591 B.n812 B.n58 585
R592 B.n58 B.n57 585
R593 B.n811 B.n810 585
R594 B.n810 B.n809 585
R595 B.n875 B.n874 585
R596 B.n873 B.n2 585
R597 B.n810 B.n60 497.305
R598 B.n807 B.n61 497.305
R599 B.n664 B.n392 497.305
R600 B.n666 B.n390 497.305
R601 B.n119 B.t8 462.875
R602 B.n116 B.t12 462.875
R603 B.n417 B.t19 462.875
R604 B.n423 B.t15 462.875
R605 B.n808 B.n114 256.663
R606 B.n808 B.n113 256.663
R607 B.n808 B.n112 256.663
R608 B.n808 B.n111 256.663
R609 B.n808 B.n110 256.663
R610 B.n808 B.n109 256.663
R611 B.n808 B.n108 256.663
R612 B.n808 B.n107 256.663
R613 B.n808 B.n106 256.663
R614 B.n808 B.n105 256.663
R615 B.n808 B.n104 256.663
R616 B.n808 B.n103 256.663
R617 B.n808 B.n102 256.663
R618 B.n808 B.n101 256.663
R619 B.n808 B.n100 256.663
R620 B.n808 B.n99 256.663
R621 B.n808 B.n98 256.663
R622 B.n808 B.n97 256.663
R623 B.n808 B.n96 256.663
R624 B.n808 B.n95 256.663
R625 B.n808 B.n94 256.663
R626 B.n808 B.n93 256.663
R627 B.n808 B.n92 256.663
R628 B.n808 B.n91 256.663
R629 B.n808 B.n90 256.663
R630 B.n808 B.n89 256.663
R631 B.n808 B.n88 256.663
R632 B.n808 B.n87 256.663
R633 B.n808 B.n86 256.663
R634 B.n808 B.n85 256.663
R635 B.n808 B.n84 256.663
R636 B.n808 B.n83 256.663
R637 B.n808 B.n82 256.663
R638 B.n808 B.n81 256.663
R639 B.n808 B.n80 256.663
R640 B.n808 B.n79 256.663
R641 B.n808 B.n78 256.663
R642 B.n808 B.n77 256.663
R643 B.n808 B.n76 256.663
R644 B.n808 B.n75 256.663
R645 B.n808 B.n74 256.663
R646 B.n808 B.n73 256.663
R647 B.n808 B.n72 256.663
R648 B.n808 B.n71 256.663
R649 B.n808 B.n70 256.663
R650 B.n808 B.n69 256.663
R651 B.n808 B.n68 256.663
R652 B.n808 B.n67 256.663
R653 B.n808 B.n66 256.663
R654 B.n808 B.n65 256.663
R655 B.n808 B.n64 256.663
R656 B.n808 B.n63 256.663
R657 B.n808 B.n62 256.663
R658 B.n450 B.n391 256.663
R659 B.n456 B.n391 256.663
R660 B.n458 B.n391 256.663
R661 B.n464 B.n391 256.663
R662 B.n466 B.n391 256.663
R663 B.n472 B.n391 256.663
R664 B.n474 B.n391 256.663
R665 B.n480 B.n391 256.663
R666 B.n482 B.n391 256.663
R667 B.n488 B.n391 256.663
R668 B.n490 B.n391 256.663
R669 B.n496 B.n391 256.663
R670 B.n498 B.n391 256.663
R671 B.n504 B.n391 256.663
R672 B.n506 B.n391 256.663
R673 B.n512 B.n391 256.663
R674 B.n514 B.n391 256.663
R675 B.n520 B.n391 256.663
R676 B.n522 B.n391 256.663
R677 B.n528 B.n391 256.663
R678 B.n530 B.n391 256.663
R679 B.n536 B.n391 256.663
R680 B.n538 B.n391 256.663
R681 B.n544 B.n391 256.663
R682 B.n546 B.n391 256.663
R683 B.n552 B.n391 256.663
R684 B.n554 B.n391 256.663
R685 B.n560 B.n391 256.663
R686 B.n562 B.n391 256.663
R687 B.n569 B.n391 256.663
R688 B.n571 B.n391 256.663
R689 B.n577 B.n391 256.663
R690 B.n579 B.n391 256.663
R691 B.n585 B.n391 256.663
R692 B.n587 B.n391 256.663
R693 B.n593 B.n391 256.663
R694 B.n595 B.n391 256.663
R695 B.n601 B.n391 256.663
R696 B.n603 B.n391 256.663
R697 B.n609 B.n391 256.663
R698 B.n611 B.n391 256.663
R699 B.n617 B.n391 256.663
R700 B.n619 B.n391 256.663
R701 B.n625 B.n391 256.663
R702 B.n627 B.n391 256.663
R703 B.n633 B.n391 256.663
R704 B.n635 B.n391 256.663
R705 B.n641 B.n391 256.663
R706 B.n643 B.n391 256.663
R707 B.n649 B.n391 256.663
R708 B.n651 B.n391 256.663
R709 B.n657 B.n391 256.663
R710 B.n659 B.n391 256.663
R711 B.n877 B.n876 256.663
R712 B.n123 B.n122 163.367
R713 B.n127 B.n126 163.367
R714 B.n131 B.n130 163.367
R715 B.n135 B.n134 163.367
R716 B.n139 B.n138 163.367
R717 B.n143 B.n142 163.367
R718 B.n147 B.n146 163.367
R719 B.n151 B.n150 163.367
R720 B.n155 B.n154 163.367
R721 B.n159 B.n158 163.367
R722 B.n163 B.n162 163.367
R723 B.n167 B.n166 163.367
R724 B.n171 B.n170 163.367
R725 B.n175 B.n174 163.367
R726 B.n179 B.n178 163.367
R727 B.n183 B.n182 163.367
R728 B.n187 B.n186 163.367
R729 B.n191 B.n190 163.367
R730 B.n195 B.n194 163.367
R731 B.n199 B.n198 163.367
R732 B.n203 B.n202 163.367
R733 B.n207 B.n206 163.367
R734 B.n211 B.n210 163.367
R735 B.n215 B.n214 163.367
R736 B.n220 B.n219 163.367
R737 B.n224 B.n223 163.367
R738 B.n228 B.n227 163.367
R739 B.n232 B.n231 163.367
R740 B.n236 B.n235 163.367
R741 B.n240 B.n239 163.367
R742 B.n244 B.n243 163.367
R743 B.n248 B.n247 163.367
R744 B.n252 B.n251 163.367
R745 B.n256 B.n255 163.367
R746 B.n260 B.n259 163.367
R747 B.n264 B.n263 163.367
R748 B.n268 B.n267 163.367
R749 B.n272 B.n271 163.367
R750 B.n276 B.n275 163.367
R751 B.n280 B.n279 163.367
R752 B.n284 B.n283 163.367
R753 B.n288 B.n287 163.367
R754 B.n292 B.n291 163.367
R755 B.n296 B.n295 163.367
R756 B.n300 B.n299 163.367
R757 B.n304 B.n303 163.367
R758 B.n308 B.n307 163.367
R759 B.n312 B.n311 163.367
R760 B.n316 B.n315 163.367
R761 B.n320 B.n319 163.367
R762 B.n324 B.n323 163.367
R763 B.n328 B.n327 163.367
R764 B.n807 B.n115 163.367
R765 B.n664 B.n386 163.367
R766 B.n672 B.n386 163.367
R767 B.n672 B.n384 163.367
R768 B.n676 B.n384 163.367
R769 B.n676 B.n379 163.367
R770 B.n685 B.n379 163.367
R771 B.n685 B.n377 163.367
R772 B.n689 B.n377 163.367
R773 B.n689 B.n371 163.367
R774 B.n697 B.n371 163.367
R775 B.n697 B.n369 163.367
R776 B.n701 B.n369 163.367
R777 B.n701 B.n364 163.367
R778 B.n710 B.n364 163.367
R779 B.n710 B.n362 163.367
R780 B.n714 B.n362 163.367
R781 B.n714 B.n356 163.367
R782 B.n722 B.n356 163.367
R783 B.n722 B.n354 163.367
R784 B.n726 B.n354 163.367
R785 B.n726 B.n347 163.367
R786 B.n734 B.n347 163.367
R787 B.n734 B.n345 163.367
R788 B.n738 B.n345 163.367
R789 B.n738 B.n340 163.367
R790 B.n746 B.n340 163.367
R791 B.n746 B.n338 163.367
R792 B.n751 B.n338 163.367
R793 B.n751 B.n332 163.367
R794 B.n759 B.n332 163.367
R795 B.n760 B.n759 163.367
R796 B.n760 B.n5 163.367
R797 B.n6 B.n5 163.367
R798 B.n7 B.n6 163.367
R799 B.n766 B.n7 163.367
R800 B.n768 B.n766 163.367
R801 B.n768 B.n12 163.367
R802 B.n13 B.n12 163.367
R803 B.n14 B.n13 163.367
R804 B.n773 B.n14 163.367
R805 B.n773 B.n19 163.367
R806 B.n20 B.n19 163.367
R807 B.n21 B.n20 163.367
R808 B.n778 B.n21 163.367
R809 B.n778 B.n26 163.367
R810 B.n27 B.n26 163.367
R811 B.n28 B.n27 163.367
R812 B.n783 B.n28 163.367
R813 B.n783 B.n33 163.367
R814 B.n34 B.n33 163.367
R815 B.n35 B.n34 163.367
R816 B.n788 B.n35 163.367
R817 B.n788 B.n40 163.367
R818 B.n41 B.n40 163.367
R819 B.n42 B.n41 163.367
R820 B.n793 B.n42 163.367
R821 B.n793 B.n47 163.367
R822 B.n48 B.n47 163.367
R823 B.n49 B.n48 163.367
R824 B.n798 B.n49 163.367
R825 B.n798 B.n54 163.367
R826 B.n55 B.n54 163.367
R827 B.n56 B.n55 163.367
R828 B.n803 B.n56 163.367
R829 B.n803 B.n61 163.367
R830 B.n451 B.n449 163.367
R831 B.n455 B.n449 163.367
R832 B.n459 B.n457 163.367
R833 B.n463 B.n447 163.367
R834 B.n467 B.n465 163.367
R835 B.n471 B.n445 163.367
R836 B.n475 B.n473 163.367
R837 B.n479 B.n443 163.367
R838 B.n483 B.n481 163.367
R839 B.n487 B.n441 163.367
R840 B.n491 B.n489 163.367
R841 B.n495 B.n439 163.367
R842 B.n499 B.n497 163.367
R843 B.n503 B.n437 163.367
R844 B.n507 B.n505 163.367
R845 B.n511 B.n435 163.367
R846 B.n515 B.n513 163.367
R847 B.n519 B.n433 163.367
R848 B.n523 B.n521 163.367
R849 B.n527 B.n431 163.367
R850 B.n531 B.n529 163.367
R851 B.n535 B.n429 163.367
R852 B.n539 B.n537 163.367
R853 B.n543 B.n427 163.367
R854 B.n547 B.n545 163.367
R855 B.n551 B.n422 163.367
R856 B.n555 B.n553 163.367
R857 B.n559 B.n420 163.367
R858 B.n563 B.n561 163.367
R859 B.n568 B.n416 163.367
R860 B.n572 B.n570 163.367
R861 B.n576 B.n414 163.367
R862 B.n580 B.n578 163.367
R863 B.n584 B.n412 163.367
R864 B.n588 B.n586 163.367
R865 B.n592 B.n410 163.367
R866 B.n596 B.n594 163.367
R867 B.n600 B.n408 163.367
R868 B.n604 B.n602 163.367
R869 B.n608 B.n406 163.367
R870 B.n612 B.n610 163.367
R871 B.n616 B.n404 163.367
R872 B.n620 B.n618 163.367
R873 B.n624 B.n402 163.367
R874 B.n628 B.n626 163.367
R875 B.n632 B.n400 163.367
R876 B.n636 B.n634 163.367
R877 B.n640 B.n398 163.367
R878 B.n644 B.n642 163.367
R879 B.n648 B.n396 163.367
R880 B.n652 B.n650 163.367
R881 B.n656 B.n394 163.367
R882 B.n660 B.n658 163.367
R883 B.n666 B.n388 163.367
R884 B.n670 B.n388 163.367
R885 B.n670 B.n382 163.367
R886 B.n679 B.n382 163.367
R887 B.n679 B.n380 163.367
R888 B.n683 B.n380 163.367
R889 B.n683 B.n375 163.367
R890 B.n691 B.n375 163.367
R891 B.n691 B.n373 163.367
R892 B.n695 B.n373 163.367
R893 B.n695 B.n367 163.367
R894 B.n704 B.n367 163.367
R895 B.n704 B.n365 163.367
R896 B.n708 B.n365 163.367
R897 B.n708 B.n360 163.367
R898 B.n716 B.n360 163.367
R899 B.n716 B.n358 163.367
R900 B.n720 B.n358 163.367
R901 B.n720 B.n352 163.367
R902 B.n728 B.n352 163.367
R903 B.n728 B.n350 163.367
R904 B.n732 B.n350 163.367
R905 B.n732 B.n344 163.367
R906 B.n740 B.n344 163.367
R907 B.n740 B.n342 163.367
R908 B.n744 B.n342 163.367
R909 B.n744 B.n336 163.367
R910 B.n753 B.n336 163.367
R911 B.n753 B.n334 163.367
R912 B.n757 B.n334 163.367
R913 B.n757 B.n3 163.367
R914 B.n875 B.n3 163.367
R915 B.n871 B.n2 163.367
R916 B.n871 B.n870 163.367
R917 B.n870 B.n9 163.367
R918 B.n866 B.n9 163.367
R919 B.n866 B.n11 163.367
R920 B.n862 B.n11 163.367
R921 B.n862 B.n16 163.367
R922 B.n858 B.n16 163.367
R923 B.n858 B.n18 163.367
R924 B.n854 B.n18 163.367
R925 B.n854 B.n23 163.367
R926 B.n850 B.n23 163.367
R927 B.n850 B.n25 163.367
R928 B.n846 B.n25 163.367
R929 B.n846 B.n30 163.367
R930 B.n842 B.n30 163.367
R931 B.n842 B.n32 163.367
R932 B.n838 B.n32 163.367
R933 B.n838 B.n36 163.367
R934 B.n834 B.n36 163.367
R935 B.n834 B.n38 163.367
R936 B.n830 B.n38 163.367
R937 B.n830 B.n44 163.367
R938 B.n826 B.n44 163.367
R939 B.n826 B.n46 163.367
R940 B.n822 B.n46 163.367
R941 B.n822 B.n50 163.367
R942 B.n818 B.n50 163.367
R943 B.n818 B.n52 163.367
R944 B.n814 B.n52 163.367
R945 B.n814 B.n58 163.367
R946 B.n810 B.n58 163.367
R947 B.n116 B.t13 101.269
R948 B.n417 B.t21 101.269
R949 B.n119 B.t10 101.249
R950 B.n423 B.t18 101.249
R951 B.n665 B.n391 75.6693
R952 B.n809 B.n808 75.6693
R953 B.n62 B.n60 71.676
R954 B.n123 B.n63 71.676
R955 B.n127 B.n64 71.676
R956 B.n131 B.n65 71.676
R957 B.n135 B.n66 71.676
R958 B.n139 B.n67 71.676
R959 B.n143 B.n68 71.676
R960 B.n147 B.n69 71.676
R961 B.n151 B.n70 71.676
R962 B.n155 B.n71 71.676
R963 B.n159 B.n72 71.676
R964 B.n163 B.n73 71.676
R965 B.n167 B.n74 71.676
R966 B.n171 B.n75 71.676
R967 B.n175 B.n76 71.676
R968 B.n179 B.n77 71.676
R969 B.n183 B.n78 71.676
R970 B.n187 B.n79 71.676
R971 B.n191 B.n80 71.676
R972 B.n195 B.n81 71.676
R973 B.n199 B.n82 71.676
R974 B.n203 B.n83 71.676
R975 B.n207 B.n84 71.676
R976 B.n211 B.n85 71.676
R977 B.n215 B.n86 71.676
R978 B.n220 B.n87 71.676
R979 B.n224 B.n88 71.676
R980 B.n228 B.n89 71.676
R981 B.n232 B.n90 71.676
R982 B.n236 B.n91 71.676
R983 B.n240 B.n92 71.676
R984 B.n244 B.n93 71.676
R985 B.n248 B.n94 71.676
R986 B.n252 B.n95 71.676
R987 B.n256 B.n96 71.676
R988 B.n260 B.n97 71.676
R989 B.n264 B.n98 71.676
R990 B.n268 B.n99 71.676
R991 B.n272 B.n100 71.676
R992 B.n276 B.n101 71.676
R993 B.n280 B.n102 71.676
R994 B.n284 B.n103 71.676
R995 B.n288 B.n104 71.676
R996 B.n292 B.n105 71.676
R997 B.n296 B.n106 71.676
R998 B.n300 B.n107 71.676
R999 B.n304 B.n108 71.676
R1000 B.n308 B.n109 71.676
R1001 B.n312 B.n110 71.676
R1002 B.n316 B.n111 71.676
R1003 B.n320 B.n112 71.676
R1004 B.n324 B.n113 71.676
R1005 B.n328 B.n114 71.676
R1006 B.n115 B.n114 71.676
R1007 B.n327 B.n113 71.676
R1008 B.n323 B.n112 71.676
R1009 B.n319 B.n111 71.676
R1010 B.n315 B.n110 71.676
R1011 B.n311 B.n109 71.676
R1012 B.n307 B.n108 71.676
R1013 B.n303 B.n107 71.676
R1014 B.n299 B.n106 71.676
R1015 B.n295 B.n105 71.676
R1016 B.n291 B.n104 71.676
R1017 B.n287 B.n103 71.676
R1018 B.n283 B.n102 71.676
R1019 B.n279 B.n101 71.676
R1020 B.n275 B.n100 71.676
R1021 B.n271 B.n99 71.676
R1022 B.n267 B.n98 71.676
R1023 B.n263 B.n97 71.676
R1024 B.n259 B.n96 71.676
R1025 B.n255 B.n95 71.676
R1026 B.n251 B.n94 71.676
R1027 B.n247 B.n93 71.676
R1028 B.n243 B.n92 71.676
R1029 B.n239 B.n91 71.676
R1030 B.n235 B.n90 71.676
R1031 B.n231 B.n89 71.676
R1032 B.n227 B.n88 71.676
R1033 B.n223 B.n87 71.676
R1034 B.n219 B.n86 71.676
R1035 B.n214 B.n85 71.676
R1036 B.n210 B.n84 71.676
R1037 B.n206 B.n83 71.676
R1038 B.n202 B.n82 71.676
R1039 B.n198 B.n81 71.676
R1040 B.n194 B.n80 71.676
R1041 B.n190 B.n79 71.676
R1042 B.n186 B.n78 71.676
R1043 B.n182 B.n77 71.676
R1044 B.n178 B.n76 71.676
R1045 B.n174 B.n75 71.676
R1046 B.n170 B.n74 71.676
R1047 B.n166 B.n73 71.676
R1048 B.n162 B.n72 71.676
R1049 B.n158 B.n71 71.676
R1050 B.n154 B.n70 71.676
R1051 B.n150 B.n69 71.676
R1052 B.n146 B.n68 71.676
R1053 B.n142 B.n67 71.676
R1054 B.n138 B.n66 71.676
R1055 B.n134 B.n65 71.676
R1056 B.n130 B.n64 71.676
R1057 B.n126 B.n63 71.676
R1058 B.n122 B.n62 71.676
R1059 B.n450 B.n390 71.676
R1060 B.n456 B.n455 71.676
R1061 B.n459 B.n458 71.676
R1062 B.n464 B.n463 71.676
R1063 B.n467 B.n466 71.676
R1064 B.n472 B.n471 71.676
R1065 B.n475 B.n474 71.676
R1066 B.n480 B.n479 71.676
R1067 B.n483 B.n482 71.676
R1068 B.n488 B.n487 71.676
R1069 B.n491 B.n490 71.676
R1070 B.n496 B.n495 71.676
R1071 B.n499 B.n498 71.676
R1072 B.n504 B.n503 71.676
R1073 B.n507 B.n506 71.676
R1074 B.n512 B.n511 71.676
R1075 B.n515 B.n514 71.676
R1076 B.n520 B.n519 71.676
R1077 B.n523 B.n522 71.676
R1078 B.n528 B.n527 71.676
R1079 B.n531 B.n530 71.676
R1080 B.n536 B.n535 71.676
R1081 B.n539 B.n538 71.676
R1082 B.n544 B.n543 71.676
R1083 B.n547 B.n546 71.676
R1084 B.n552 B.n551 71.676
R1085 B.n555 B.n554 71.676
R1086 B.n560 B.n559 71.676
R1087 B.n563 B.n562 71.676
R1088 B.n569 B.n568 71.676
R1089 B.n572 B.n571 71.676
R1090 B.n577 B.n576 71.676
R1091 B.n580 B.n579 71.676
R1092 B.n585 B.n584 71.676
R1093 B.n588 B.n587 71.676
R1094 B.n593 B.n592 71.676
R1095 B.n596 B.n595 71.676
R1096 B.n601 B.n600 71.676
R1097 B.n604 B.n603 71.676
R1098 B.n609 B.n608 71.676
R1099 B.n612 B.n611 71.676
R1100 B.n617 B.n616 71.676
R1101 B.n620 B.n619 71.676
R1102 B.n625 B.n624 71.676
R1103 B.n628 B.n627 71.676
R1104 B.n633 B.n632 71.676
R1105 B.n636 B.n635 71.676
R1106 B.n641 B.n640 71.676
R1107 B.n644 B.n643 71.676
R1108 B.n649 B.n648 71.676
R1109 B.n652 B.n651 71.676
R1110 B.n657 B.n656 71.676
R1111 B.n660 B.n659 71.676
R1112 B.n451 B.n450 71.676
R1113 B.n457 B.n456 71.676
R1114 B.n458 B.n447 71.676
R1115 B.n465 B.n464 71.676
R1116 B.n466 B.n445 71.676
R1117 B.n473 B.n472 71.676
R1118 B.n474 B.n443 71.676
R1119 B.n481 B.n480 71.676
R1120 B.n482 B.n441 71.676
R1121 B.n489 B.n488 71.676
R1122 B.n490 B.n439 71.676
R1123 B.n497 B.n496 71.676
R1124 B.n498 B.n437 71.676
R1125 B.n505 B.n504 71.676
R1126 B.n506 B.n435 71.676
R1127 B.n513 B.n512 71.676
R1128 B.n514 B.n433 71.676
R1129 B.n521 B.n520 71.676
R1130 B.n522 B.n431 71.676
R1131 B.n529 B.n528 71.676
R1132 B.n530 B.n429 71.676
R1133 B.n537 B.n536 71.676
R1134 B.n538 B.n427 71.676
R1135 B.n545 B.n544 71.676
R1136 B.n546 B.n422 71.676
R1137 B.n553 B.n552 71.676
R1138 B.n554 B.n420 71.676
R1139 B.n561 B.n560 71.676
R1140 B.n562 B.n416 71.676
R1141 B.n570 B.n569 71.676
R1142 B.n571 B.n414 71.676
R1143 B.n578 B.n577 71.676
R1144 B.n579 B.n412 71.676
R1145 B.n586 B.n585 71.676
R1146 B.n587 B.n410 71.676
R1147 B.n594 B.n593 71.676
R1148 B.n595 B.n408 71.676
R1149 B.n602 B.n601 71.676
R1150 B.n603 B.n406 71.676
R1151 B.n610 B.n609 71.676
R1152 B.n611 B.n404 71.676
R1153 B.n618 B.n617 71.676
R1154 B.n619 B.n402 71.676
R1155 B.n626 B.n625 71.676
R1156 B.n627 B.n400 71.676
R1157 B.n634 B.n633 71.676
R1158 B.n635 B.n398 71.676
R1159 B.n642 B.n641 71.676
R1160 B.n643 B.n396 71.676
R1161 B.n650 B.n649 71.676
R1162 B.n651 B.n394 71.676
R1163 B.n658 B.n657 71.676
R1164 B.n659 B.n392 71.676
R1165 B.n876 B.n875 71.676
R1166 B.n876 B.n2 71.676
R1167 B.n117 B.t14 68.8808
R1168 B.n418 B.t20 68.8808
R1169 B.n120 B.t11 68.862
R1170 B.n424 B.t17 68.862
R1171 B.n217 B.n120 59.5399
R1172 B.n118 B.n117 59.5399
R1173 B.n565 B.n418 59.5399
R1174 B.n425 B.n424 59.5399
R1175 B.n665 B.n387 38.1151
R1176 B.n671 B.n387 38.1151
R1177 B.n671 B.n383 38.1151
R1178 B.n678 B.n383 38.1151
R1179 B.n678 B.n677 38.1151
R1180 B.n684 B.n376 38.1151
R1181 B.n690 B.n376 38.1151
R1182 B.n690 B.n372 38.1151
R1183 B.n696 B.n372 38.1151
R1184 B.n696 B.n368 38.1151
R1185 B.n703 B.n368 38.1151
R1186 B.n703 B.n702 38.1151
R1187 B.n709 B.n361 38.1151
R1188 B.n715 B.n361 38.1151
R1189 B.n715 B.n357 38.1151
R1190 B.n721 B.n357 38.1151
R1191 B.n727 B.n353 38.1151
R1192 B.n727 B.n348 38.1151
R1193 B.n733 B.n348 38.1151
R1194 B.n733 B.n349 38.1151
R1195 B.n739 B.n341 38.1151
R1196 B.n745 B.n341 38.1151
R1197 B.n745 B.n337 38.1151
R1198 B.n752 B.n337 38.1151
R1199 B.n758 B.n333 38.1151
R1200 B.n758 B.n4 38.1151
R1201 B.n874 B.n4 38.1151
R1202 B.n874 B.n873 38.1151
R1203 B.n873 B.n872 38.1151
R1204 B.n872 B.n8 38.1151
R1205 B.n767 B.n8 38.1151
R1206 B.n865 B.n864 38.1151
R1207 B.n864 B.n863 38.1151
R1208 B.n863 B.n15 38.1151
R1209 B.n857 B.n15 38.1151
R1210 B.n856 B.n855 38.1151
R1211 B.n855 B.n22 38.1151
R1212 B.n849 B.n22 38.1151
R1213 B.n849 B.n848 38.1151
R1214 B.n847 B.n29 38.1151
R1215 B.n841 B.n29 38.1151
R1216 B.n841 B.n840 38.1151
R1217 B.n840 B.n839 38.1151
R1218 B.n833 B.n39 38.1151
R1219 B.n833 B.n832 38.1151
R1220 B.n832 B.n831 38.1151
R1221 B.n831 B.n43 38.1151
R1222 B.n825 B.n43 38.1151
R1223 B.n825 B.n824 38.1151
R1224 B.n824 B.n823 38.1151
R1225 B.n817 B.n53 38.1151
R1226 B.n817 B.n816 38.1151
R1227 B.n816 B.n815 38.1151
R1228 B.n815 B.n57 38.1151
R1229 B.n809 B.n57 38.1151
R1230 B.n120 B.n119 32.3884
R1231 B.n117 B.n116 32.3884
R1232 B.n418 B.n417 32.3884
R1233 B.n424 B.n423 32.3884
R1234 B.n667 B.n389 32.3127
R1235 B.n663 B.n662 32.3127
R1236 B.n806 B.n805 32.3127
R1237 B.n811 B.n59 32.3127
R1238 B.n702 B.t2 26.905
R1239 B.n39 B.t6 26.905
R1240 B.n721 B.t7 23.5419
R1241 B.t3 B.n847 23.5419
R1242 B.n677 B.t16 22.4209
R1243 B.n53 B.t9 22.4209
R1244 B.t4 B.n333 21.2999
R1245 B.n767 B.t0 21.2999
R1246 B.n349 B.t5 20.1788
R1247 B.t1 B.n856 20.1788
R1248 B B.n877 18.0485
R1249 B.n739 B.t5 17.9368
R1250 B.n857 B.t1 17.9368
R1251 B.n752 B.t4 16.8158
R1252 B.n865 B.t0 16.8158
R1253 B.n684 B.t16 15.6948
R1254 B.n823 B.t9 15.6948
R1255 B.t7 B.n353 14.5737
R1256 B.n848 B.t3 14.5737
R1257 B.n709 B.t2 11.2107
R1258 B.n839 B.t6 11.2107
R1259 B.n668 B.n667 10.6151
R1260 B.n669 B.n668 10.6151
R1261 B.n669 B.n381 10.6151
R1262 B.n680 B.n381 10.6151
R1263 B.n681 B.n680 10.6151
R1264 B.n682 B.n681 10.6151
R1265 B.n682 B.n374 10.6151
R1266 B.n692 B.n374 10.6151
R1267 B.n693 B.n692 10.6151
R1268 B.n694 B.n693 10.6151
R1269 B.n694 B.n366 10.6151
R1270 B.n705 B.n366 10.6151
R1271 B.n706 B.n705 10.6151
R1272 B.n707 B.n706 10.6151
R1273 B.n707 B.n359 10.6151
R1274 B.n717 B.n359 10.6151
R1275 B.n718 B.n717 10.6151
R1276 B.n719 B.n718 10.6151
R1277 B.n719 B.n351 10.6151
R1278 B.n729 B.n351 10.6151
R1279 B.n730 B.n729 10.6151
R1280 B.n731 B.n730 10.6151
R1281 B.n731 B.n343 10.6151
R1282 B.n741 B.n343 10.6151
R1283 B.n742 B.n741 10.6151
R1284 B.n743 B.n742 10.6151
R1285 B.n743 B.n335 10.6151
R1286 B.n754 B.n335 10.6151
R1287 B.n755 B.n754 10.6151
R1288 B.n756 B.n755 10.6151
R1289 B.n756 B.n0 10.6151
R1290 B.n452 B.n389 10.6151
R1291 B.n453 B.n452 10.6151
R1292 B.n454 B.n453 10.6151
R1293 B.n454 B.n448 10.6151
R1294 B.n460 B.n448 10.6151
R1295 B.n461 B.n460 10.6151
R1296 B.n462 B.n461 10.6151
R1297 B.n462 B.n446 10.6151
R1298 B.n468 B.n446 10.6151
R1299 B.n469 B.n468 10.6151
R1300 B.n470 B.n469 10.6151
R1301 B.n470 B.n444 10.6151
R1302 B.n476 B.n444 10.6151
R1303 B.n477 B.n476 10.6151
R1304 B.n478 B.n477 10.6151
R1305 B.n478 B.n442 10.6151
R1306 B.n484 B.n442 10.6151
R1307 B.n485 B.n484 10.6151
R1308 B.n486 B.n485 10.6151
R1309 B.n486 B.n440 10.6151
R1310 B.n492 B.n440 10.6151
R1311 B.n493 B.n492 10.6151
R1312 B.n494 B.n493 10.6151
R1313 B.n494 B.n438 10.6151
R1314 B.n500 B.n438 10.6151
R1315 B.n501 B.n500 10.6151
R1316 B.n502 B.n501 10.6151
R1317 B.n502 B.n436 10.6151
R1318 B.n508 B.n436 10.6151
R1319 B.n509 B.n508 10.6151
R1320 B.n510 B.n509 10.6151
R1321 B.n510 B.n434 10.6151
R1322 B.n516 B.n434 10.6151
R1323 B.n517 B.n516 10.6151
R1324 B.n518 B.n517 10.6151
R1325 B.n518 B.n432 10.6151
R1326 B.n524 B.n432 10.6151
R1327 B.n525 B.n524 10.6151
R1328 B.n526 B.n525 10.6151
R1329 B.n526 B.n430 10.6151
R1330 B.n532 B.n430 10.6151
R1331 B.n533 B.n532 10.6151
R1332 B.n534 B.n533 10.6151
R1333 B.n534 B.n428 10.6151
R1334 B.n540 B.n428 10.6151
R1335 B.n541 B.n540 10.6151
R1336 B.n542 B.n541 10.6151
R1337 B.n542 B.n426 10.6151
R1338 B.n549 B.n548 10.6151
R1339 B.n550 B.n549 10.6151
R1340 B.n550 B.n421 10.6151
R1341 B.n556 B.n421 10.6151
R1342 B.n557 B.n556 10.6151
R1343 B.n558 B.n557 10.6151
R1344 B.n558 B.n419 10.6151
R1345 B.n564 B.n419 10.6151
R1346 B.n567 B.n566 10.6151
R1347 B.n567 B.n415 10.6151
R1348 B.n573 B.n415 10.6151
R1349 B.n574 B.n573 10.6151
R1350 B.n575 B.n574 10.6151
R1351 B.n575 B.n413 10.6151
R1352 B.n581 B.n413 10.6151
R1353 B.n582 B.n581 10.6151
R1354 B.n583 B.n582 10.6151
R1355 B.n583 B.n411 10.6151
R1356 B.n589 B.n411 10.6151
R1357 B.n590 B.n589 10.6151
R1358 B.n591 B.n590 10.6151
R1359 B.n591 B.n409 10.6151
R1360 B.n597 B.n409 10.6151
R1361 B.n598 B.n597 10.6151
R1362 B.n599 B.n598 10.6151
R1363 B.n599 B.n407 10.6151
R1364 B.n605 B.n407 10.6151
R1365 B.n606 B.n605 10.6151
R1366 B.n607 B.n606 10.6151
R1367 B.n607 B.n405 10.6151
R1368 B.n613 B.n405 10.6151
R1369 B.n614 B.n613 10.6151
R1370 B.n615 B.n614 10.6151
R1371 B.n615 B.n403 10.6151
R1372 B.n621 B.n403 10.6151
R1373 B.n622 B.n621 10.6151
R1374 B.n623 B.n622 10.6151
R1375 B.n623 B.n401 10.6151
R1376 B.n629 B.n401 10.6151
R1377 B.n630 B.n629 10.6151
R1378 B.n631 B.n630 10.6151
R1379 B.n631 B.n399 10.6151
R1380 B.n637 B.n399 10.6151
R1381 B.n638 B.n637 10.6151
R1382 B.n639 B.n638 10.6151
R1383 B.n639 B.n397 10.6151
R1384 B.n645 B.n397 10.6151
R1385 B.n646 B.n645 10.6151
R1386 B.n647 B.n646 10.6151
R1387 B.n647 B.n395 10.6151
R1388 B.n653 B.n395 10.6151
R1389 B.n654 B.n653 10.6151
R1390 B.n655 B.n654 10.6151
R1391 B.n655 B.n393 10.6151
R1392 B.n661 B.n393 10.6151
R1393 B.n662 B.n661 10.6151
R1394 B.n663 B.n385 10.6151
R1395 B.n673 B.n385 10.6151
R1396 B.n674 B.n673 10.6151
R1397 B.n675 B.n674 10.6151
R1398 B.n675 B.n378 10.6151
R1399 B.n686 B.n378 10.6151
R1400 B.n687 B.n686 10.6151
R1401 B.n688 B.n687 10.6151
R1402 B.n688 B.n370 10.6151
R1403 B.n698 B.n370 10.6151
R1404 B.n699 B.n698 10.6151
R1405 B.n700 B.n699 10.6151
R1406 B.n700 B.n363 10.6151
R1407 B.n711 B.n363 10.6151
R1408 B.n712 B.n711 10.6151
R1409 B.n713 B.n712 10.6151
R1410 B.n713 B.n355 10.6151
R1411 B.n723 B.n355 10.6151
R1412 B.n724 B.n723 10.6151
R1413 B.n725 B.n724 10.6151
R1414 B.n725 B.n346 10.6151
R1415 B.n735 B.n346 10.6151
R1416 B.n736 B.n735 10.6151
R1417 B.n737 B.n736 10.6151
R1418 B.n737 B.n339 10.6151
R1419 B.n747 B.n339 10.6151
R1420 B.n748 B.n747 10.6151
R1421 B.n750 B.n748 10.6151
R1422 B.n750 B.n749 10.6151
R1423 B.n749 B.n331 10.6151
R1424 B.n761 B.n331 10.6151
R1425 B.n762 B.n761 10.6151
R1426 B.n763 B.n762 10.6151
R1427 B.n764 B.n763 10.6151
R1428 B.n765 B.n764 10.6151
R1429 B.n769 B.n765 10.6151
R1430 B.n770 B.n769 10.6151
R1431 B.n771 B.n770 10.6151
R1432 B.n772 B.n771 10.6151
R1433 B.n774 B.n772 10.6151
R1434 B.n775 B.n774 10.6151
R1435 B.n776 B.n775 10.6151
R1436 B.n777 B.n776 10.6151
R1437 B.n779 B.n777 10.6151
R1438 B.n780 B.n779 10.6151
R1439 B.n781 B.n780 10.6151
R1440 B.n782 B.n781 10.6151
R1441 B.n784 B.n782 10.6151
R1442 B.n785 B.n784 10.6151
R1443 B.n786 B.n785 10.6151
R1444 B.n787 B.n786 10.6151
R1445 B.n789 B.n787 10.6151
R1446 B.n790 B.n789 10.6151
R1447 B.n791 B.n790 10.6151
R1448 B.n792 B.n791 10.6151
R1449 B.n794 B.n792 10.6151
R1450 B.n795 B.n794 10.6151
R1451 B.n796 B.n795 10.6151
R1452 B.n797 B.n796 10.6151
R1453 B.n799 B.n797 10.6151
R1454 B.n800 B.n799 10.6151
R1455 B.n801 B.n800 10.6151
R1456 B.n802 B.n801 10.6151
R1457 B.n804 B.n802 10.6151
R1458 B.n805 B.n804 10.6151
R1459 B.n869 B.n1 10.6151
R1460 B.n869 B.n868 10.6151
R1461 B.n868 B.n867 10.6151
R1462 B.n867 B.n10 10.6151
R1463 B.n861 B.n10 10.6151
R1464 B.n861 B.n860 10.6151
R1465 B.n860 B.n859 10.6151
R1466 B.n859 B.n17 10.6151
R1467 B.n853 B.n17 10.6151
R1468 B.n853 B.n852 10.6151
R1469 B.n852 B.n851 10.6151
R1470 B.n851 B.n24 10.6151
R1471 B.n845 B.n24 10.6151
R1472 B.n845 B.n844 10.6151
R1473 B.n844 B.n843 10.6151
R1474 B.n843 B.n31 10.6151
R1475 B.n837 B.n31 10.6151
R1476 B.n837 B.n836 10.6151
R1477 B.n836 B.n835 10.6151
R1478 B.n835 B.n37 10.6151
R1479 B.n829 B.n37 10.6151
R1480 B.n829 B.n828 10.6151
R1481 B.n828 B.n827 10.6151
R1482 B.n827 B.n45 10.6151
R1483 B.n821 B.n45 10.6151
R1484 B.n821 B.n820 10.6151
R1485 B.n820 B.n819 10.6151
R1486 B.n819 B.n51 10.6151
R1487 B.n813 B.n51 10.6151
R1488 B.n813 B.n812 10.6151
R1489 B.n812 B.n811 10.6151
R1490 B.n121 B.n59 10.6151
R1491 B.n124 B.n121 10.6151
R1492 B.n125 B.n124 10.6151
R1493 B.n128 B.n125 10.6151
R1494 B.n129 B.n128 10.6151
R1495 B.n132 B.n129 10.6151
R1496 B.n133 B.n132 10.6151
R1497 B.n136 B.n133 10.6151
R1498 B.n137 B.n136 10.6151
R1499 B.n140 B.n137 10.6151
R1500 B.n141 B.n140 10.6151
R1501 B.n144 B.n141 10.6151
R1502 B.n145 B.n144 10.6151
R1503 B.n148 B.n145 10.6151
R1504 B.n149 B.n148 10.6151
R1505 B.n152 B.n149 10.6151
R1506 B.n153 B.n152 10.6151
R1507 B.n156 B.n153 10.6151
R1508 B.n157 B.n156 10.6151
R1509 B.n160 B.n157 10.6151
R1510 B.n161 B.n160 10.6151
R1511 B.n164 B.n161 10.6151
R1512 B.n165 B.n164 10.6151
R1513 B.n168 B.n165 10.6151
R1514 B.n169 B.n168 10.6151
R1515 B.n172 B.n169 10.6151
R1516 B.n173 B.n172 10.6151
R1517 B.n176 B.n173 10.6151
R1518 B.n177 B.n176 10.6151
R1519 B.n180 B.n177 10.6151
R1520 B.n181 B.n180 10.6151
R1521 B.n184 B.n181 10.6151
R1522 B.n185 B.n184 10.6151
R1523 B.n188 B.n185 10.6151
R1524 B.n189 B.n188 10.6151
R1525 B.n192 B.n189 10.6151
R1526 B.n193 B.n192 10.6151
R1527 B.n196 B.n193 10.6151
R1528 B.n197 B.n196 10.6151
R1529 B.n200 B.n197 10.6151
R1530 B.n201 B.n200 10.6151
R1531 B.n204 B.n201 10.6151
R1532 B.n205 B.n204 10.6151
R1533 B.n208 B.n205 10.6151
R1534 B.n209 B.n208 10.6151
R1535 B.n212 B.n209 10.6151
R1536 B.n213 B.n212 10.6151
R1537 B.n216 B.n213 10.6151
R1538 B.n221 B.n218 10.6151
R1539 B.n222 B.n221 10.6151
R1540 B.n225 B.n222 10.6151
R1541 B.n226 B.n225 10.6151
R1542 B.n229 B.n226 10.6151
R1543 B.n230 B.n229 10.6151
R1544 B.n233 B.n230 10.6151
R1545 B.n234 B.n233 10.6151
R1546 B.n238 B.n237 10.6151
R1547 B.n241 B.n238 10.6151
R1548 B.n242 B.n241 10.6151
R1549 B.n245 B.n242 10.6151
R1550 B.n246 B.n245 10.6151
R1551 B.n249 B.n246 10.6151
R1552 B.n250 B.n249 10.6151
R1553 B.n253 B.n250 10.6151
R1554 B.n254 B.n253 10.6151
R1555 B.n257 B.n254 10.6151
R1556 B.n258 B.n257 10.6151
R1557 B.n261 B.n258 10.6151
R1558 B.n262 B.n261 10.6151
R1559 B.n265 B.n262 10.6151
R1560 B.n266 B.n265 10.6151
R1561 B.n269 B.n266 10.6151
R1562 B.n270 B.n269 10.6151
R1563 B.n273 B.n270 10.6151
R1564 B.n274 B.n273 10.6151
R1565 B.n277 B.n274 10.6151
R1566 B.n278 B.n277 10.6151
R1567 B.n281 B.n278 10.6151
R1568 B.n282 B.n281 10.6151
R1569 B.n285 B.n282 10.6151
R1570 B.n286 B.n285 10.6151
R1571 B.n289 B.n286 10.6151
R1572 B.n290 B.n289 10.6151
R1573 B.n293 B.n290 10.6151
R1574 B.n294 B.n293 10.6151
R1575 B.n297 B.n294 10.6151
R1576 B.n298 B.n297 10.6151
R1577 B.n301 B.n298 10.6151
R1578 B.n302 B.n301 10.6151
R1579 B.n305 B.n302 10.6151
R1580 B.n306 B.n305 10.6151
R1581 B.n309 B.n306 10.6151
R1582 B.n310 B.n309 10.6151
R1583 B.n313 B.n310 10.6151
R1584 B.n314 B.n313 10.6151
R1585 B.n317 B.n314 10.6151
R1586 B.n318 B.n317 10.6151
R1587 B.n321 B.n318 10.6151
R1588 B.n322 B.n321 10.6151
R1589 B.n325 B.n322 10.6151
R1590 B.n326 B.n325 10.6151
R1591 B.n329 B.n326 10.6151
R1592 B.n330 B.n329 10.6151
R1593 B.n806 B.n330 10.6151
R1594 B.n877 B.n0 8.11757
R1595 B.n877 B.n1 8.11757
R1596 B.n548 B.n425 6.5566
R1597 B.n565 B.n564 6.5566
R1598 B.n218 B.n217 6.5566
R1599 B.n234 B.n118 6.5566
R1600 B.n426 B.n425 4.05904
R1601 B.n566 B.n565 4.05904
R1602 B.n217 B.n216 4.05904
R1603 B.n237 B.n118 4.05904
R1604 VN.n5 VN.t6 287.204
R1605 VN.n25 VN.t4 287.204
R1606 VN.n4 VN.t3 258.087
R1607 VN.n10 VN.t2 258.087
R1608 VN.n17 VN.t1 258.087
R1609 VN.n24 VN.t5 258.087
R1610 VN.n22 VN.t7 258.087
R1611 VN.n36 VN.t0 258.087
R1612 VN.n18 VN.n17 173.29
R1613 VN.n37 VN.n36 173.29
R1614 VN.n35 VN.n19 161.3
R1615 VN.n34 VN.n33 161.3
R1616 VN.n32 VN.n20 161.3
R1617 VN.n31 VN.n30 161.3
R1618 VN.n29 VN.n21 161.3
R1619 VN.n28 VN.n27 161.3
R1620 VN.n26 VN.n23 161.3
R1621 VN.n16 VN.n0 161.3
R1622 VN.n15 VN.n14 161.3
R1623 VN.n13 VN.n1 161.3
R1624 VN.n12 VN.n11 161.3
R1625 VN.n9 VN.n2 161.3
R1626 VN.n8 VN.n7 161.3
R1627 VN.n6 VN.n3 161.3
R1628 VN.n5 VN.n4 61.1116
R1629 VN.n25 VN.n24 61.1116
R1630 VN.n9 VN.n8 56.5193
R1631 VN.n29 VN.n28 56.5193
R1632 VN.n15 VN.n1 48.2635
R1633 VN.n34 VN.n20 48.2635
R1634 VN VN.n37 47.0857
R1635 VN.n16 VN.n15 32.7233
R1636 VN.n35 VN.n34 32.7233
R1637 VN.n26 VN.n25 27.209
R1638 VN.n6 VN.n5 27.209
R1639 VN.n8 VN.n3 24.4675
R1640 VN.n11 VN.n9 24.4675
R1641 VN.n28 VN.n23 24.4675
R1642 VN.n30 VN.n29 24.4675
R1643 VN.n10 VN.n1 20.3081
R1644 VN.n22 VN.n20 20.3081
R1645 VN.n17 VN.n16 12.4787
R1646 VN.n36 VN.n35 12.4787
R1647 VN.n4 VN.n3 4.15989
R1648 VN.n11 VN.n10 4.15989
R1649 VN.n24 VN.n23 4.15989
R1650 VN.n30 VN.n22 4.15989
R1651 VN.n37 VN.n19 0.189894
R1652 VN.n33 VN.n19 0.189894
R1653 VN.n33 VN.n32 0.189894
R1654 VN.n32 VN.n31 0.189894
R1655 VN.n31 VN.n21 0.189894
R1656 VN.n27 VN.n21 0.189894
R1657 VN.n27 VN.n26 0.189894
R1658 VN.n7 VN.n6 0.189894
R1659 VN.n7 VN.n2 0.189894
R1660 VN.n12 VN.n2 0.189894
R1661 VN.n13 VN.n12 0.189894
R1662 VN.n14 VN.n13 0.189894
R1663 VN.n14 VN.n0 0.189894
R1664 VN.n18 VN.n0 0.189894
R1665 VN VN.n18 0.0516364
R1666 VDD2.n2 VDD2.n1 62.9877
R1667 VDD2.n2 VDD2.n0 62.9877
R1668 VDD2 VDD2.n5 62.9849
R1669 VDD2.n4 VDD2.n3 62.3235
R1670 VDD2.n4 VDD2.n2 42.5644
R1671 VDD2.n5 VDD2.t2 1.38029
R1672 VDD2.n5 VDD2.t3 1.38029
R1673 VDD2.n3 VDD2.t7 1.38029
R1674 VDD2.n3 VDD2.t0 1.38029
R1675 VDD2.n1 VDD2.t5 1.38029
R1676 VDD2.n1 VDD2.t6 1.38029
R1677 VDD2.n0 VDD2.t1 1.38029
R1678 VDD2.n0 VDD2.t4 1.38029
R1679 VDD2 VDD2.n4 0.778517
C0 VP VDD1 8.87287f
C1 VTAIL VDD1 9.8747f
C2 VDD1 VDD2 1.14581f
C3 VN VDD1 0.149195f
C4 VTAIL VP 8.54457f
C5 VP VDD2 0.385338f
C6 VTAIL VDD2 9.920671f
C7 VP VN 6.55739f
C8 VN VDD2 8.63749f
C9 VTAIL VN 8.53046f
C10 VDD2 B 4.281921f
C11 VDD1 B 4.586419f
C12 VTAIL B 10.882407f
C13 VN B 11.034531f
C14 VP B 9.297294f
C15 VDD2.t1 B 0.285299f
C16 VDD2.t4 B 0.285299f
C17 VDD2.n0 B 2.57899f
C18 VDD2.t5 B 0.285299f
C19 VDD2.t6 B 0.285299f
C20 VDD2.n1 B 2.57899f
C21 VDD2.n2 B 2.70194f
C22 VDD2.t7 B 0.285299f
C23 VDD2.t0 B 0.285299f
C24 VDD2.n3 B 2.57493f
C25 VDD2.n4 B 2.70688f
C26 VDD2.t2 B 0.285299f
C27 VDD2.t3 B 0.285299f
C28 VDD2.n5 B 2.57896f
C29 VN.n0 B 0.032474f
C30 VN.t1 B 1.70932f
C31 VN.n1 B 0.055734f
C32 VN.n2 B 0.032474f
C33 VN.n3 B 0.035721f
C34 VN.t6 B 1.78224f
C35 VN.t3 B 1.70932f
C36 VN.n4 B 0.658115f
C37 VN.n5 B 0.694239f
C38 VN.n6 B 0.172307f
C39 VN.n7 B 0.032474f
C40 VN.n8 B 0.047406f
C41 VN.n9 B 0.047406f
C42 VN.t2 B 1.70932f
C43 VN.n10 B 0.6132f
C44 VN.n11 B 0.035721f
C45 VN.n12 B 0.032474f
C46 VN.n13 B 0.032474f
C47 VN.n14 B 0.032474f
C48 VN.n15 B 0.029023f
C49 VN.n16 B 0.050853f
C50 VN.n17 B 0.674819f
C51 VN.n18 B 0.029746f
C52 VN.n19 B 0.032474f
C53 VN.t0 B 1.70932f
C54 VN.n20 B 0.055734f
C55 VN.n21 B 0.032474f
C56 VN.t7 B 1.70932f
C57 VN.n22 B 0.6132f
C58 VN.n23 B 0.035721f
C59 VN.t4 B 1.78224f
C60 VN.t5 B 1.70932f
C61 VN.n24 B 0.658115f
C62 VN.n25 B 0.694239f
C63 VN.n26 B 0.172307f
C64 VN.n27 B 0.032474f
C65 VN.n28 B 0.047406f
C66 VN.n29 B 0.047406f
C67 VN.n30 B 0.035721f
C68 VN.n31 B 0.032474f
C69 VN.n32 B 0.032474f
C70 VN.n33 B 0.032474f
C71 VN.n34 B 0.029023f
C72 VN.n35 B 0.050853f
C73 VN.n36 B 0.674819f
C74 VN.n37 B 1.61628f
C75 VTAIL.t1 B 0.212936f
C76 VTAIL.t3 B 0.212936f
C77 VTAIL.n0 B 1.86756f
C78 VTAIL.n1 B 0.271447f
C79 VTAIL.t0 B 2.38269f
C80 VTAIL.n2 B 0.361951f
C81 VTAIL.t11 B 2.38269f
C82 VTAIL.n3 B 0.361951f
C83 VTAIL.t8 B 0.212936f
C84 VTAIL.t12 B 0.212936f
C85 VTAIL.n4 B 1.86756f
C86 VTAIL.n5 B 0.355033f
C87 VTAIL.t9 B 2.38269f
C88 VTAIL.n6 B 1.42421f
C89 VTAIL.t2 B 2.38271f
C90 VTAIL.n7 B 1.42419f
C91 VTAIL.t7 B 0.212936f
C92 VTAIL.t5 B 0.212936f
C93 VTAIL.n8 B 1.86756f
C94 VTAIL.n9 B 0.355031f
C95 VTAIL.t4 B 2.38271f
C96 VTAIL.n10 B 0.361934f
C97 VTAIL.t13 B 2.38271f
C98 VTAIL.n11 B 0.361934f
C99 VTAIL.t14 B 0.212936f
C100 VTAIL.t15 B 0.212936f
C101 VTAIL.n12 B 1.86756f
C102 VTAIL.n13 B 0.355031f
C103 VTAIL.t10 B 2.38269f
C104 VTAIL.n14 B 1.42421f
C105 VTAIL.t6 B 2.38269f
C106 VTAIL.n15 B 1.42068f
C107 VDD1.t4 B 0.288477f
C108 VDD1.t0 B 0.288477f
C109 VDD1.n0 B 2.60851f
C110 VDD1.t5 B 0.288477f
C111 VDD1.t1 B 0.288477f
C112 VDD1.n1 B 2.60772f
C113 VDD1.t6 B 0.288477f
C114 VDD1.t2 B 0.288477f
C115 VDD1.n2 B 2.60772f
C116 VDD1.n3 B 2.78571f
C117 VDD1.t7 B 0.288477f
C118 VDD1.t3 B 0.288477f
C119 VDD1.n4 B 2.6036f
C120 VDD1.n5 B 2.76778f
C121 VP.n0 B 0.032948f
C122 VP.t4 B 1.7343f
C123 VP.n1 B 0.056548f
C124 VP.n2 B 0.032948f
C125 VP.n3 B 0.036243f
C126 VP.n4 B 0.032948f
C127 VP.t6 B 1.7343f
C128 VP.n5 B 0.68468f
C129 VP.n6 B 0.032948f
C130 VP.t5 B 1.7343f
C131 VP.n7 B 0.056548f
C132 VP.n8 B 0.032948f
C133 VP.n9 B 0.036243f
C134 VP.t2 B 1.80829f
C135 VP.t1 B 1.7343f
C136 VP.n10 B 0.667732f
C137 VP.n11 B 0.704383f
C138 VP.n12 B 0.174825f
C139 VP.n13 B 0.032948f
C140 VP.n14 B 0.048099f
C141 VP.n15 B 0.048099f
C142 VP.t0 B 1.7343f
C143 VP.n16 B 0.622161f
C144 VP.n17 B 0.036243f
C145 VP.n18 B 0.032948f
C146 VP.n19 B 0.032948f
C147 VP.n20 B 0.032948f
C148 VP.n21 B 0.029447f
C149 VP.n22 B 0.051596f
C150 VP.n23 B 0.68468f
C151 VP.n24 B 1.6184f
C152 VP.n25 B 1.64376f
C153 VP.n26 B 0.032948f
C154 VP.n27 B 0.051596f
C155 VP.n28 B 0.029447f
C156 VP.t7 B 1.7343f
C157 VP.n29 B 0.622161f
C158 VP.n30 B 0.056548f
C159 VP.n31 B 0.032948f
C160 VP.n32 B 0.032948f
C161 VP.n33 B 0.032948f
C162 VP.n34 B 0.048099f
C163 VP.n35 B 0.048099f
C164 VP.t3 B 1.7343f
C165 VP.n36 B 0.622161f
C166 VP.n37 B 0.036243f
C167 VP.n38 B 0.032948f
C168 VP.n39 B 0.032948f
C169 VP.n40 B 0.032948f
C170 VP.n41 B 0.029447f
C171 VP.n42 B 0.051596f
C172 VP.n43 B 0.68468f
C173 VP.n44 B 0.03018f
.ends

