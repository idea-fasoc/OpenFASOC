* NGSPICE file created from diff_pair_sample_0020.ext - technology: sky130A

.subckt diff_pair_sample_0020 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.858 pd=5.18 as=0 ps=0 w=2.2 l=2.59
X1 B.t8 B.t6 B.t7 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.858 pd=5.18 as=0 ps=0 w=2.2 l=2.59
X2 VDD1.t3 VP.t0 VTAIL.t5 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.363 pd=2.53 as=0.858 ps=5.18 w=2.2 l=2.59
X3 VDD2.t3 VN.t0 VTAIL.t1 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.363 pd=2.53 as=0.858 ps=5.18 w=2.2 l=2.59
X4 VDD1.t2 VP.t1 VTAIL.t4 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.363 pd=2.53 as=0.858 ps=5.18 w=2.2 l=2.59
X5 VTAIL.t7 VP.t2 VDD1.t1 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.858 pd=5.18 as=0.363 ps=2.53 w=2.2 l=2.59
X6 VDD2.t2 VN.t1 VTAIL.t2 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.363 pd=2.53 as=0.858 ps=5.18 w=2.2 l=2.59
X7 VTAIL.t0 VN.t2 VDD2.t1 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.858 pd=5.18 as=0.363 ps=2.53 w=2.2 l=2.59
X8 VTAIL.t3 VN.t3 VDD2.t0 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.858 pd=5.18 as=0.363 ps=2.53 w=2.2 l=2.59
X9 B.t5 B.t3 B.t4 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.858 pd=5.18 as=0 ps=0 w=2.2 l=2.59
X10 B.t2 B.t0 B.t1 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.858 pd=5.18 as=0 ps=0 w=2.2 l=2.59
X11 VTAIL.t6 VP.t3 VDD1.t0 w_n2722_n1408# sky130_fd_pr__pfet_01v8 ad=0.858 pd=5.18 as=0.363 ps=2.53 w=2.2 l=2.59
R0 B.n322 B.n321 585
R1 B.n323 B.n40 585
R2 B.n325 B.n324 585
R3 B.n326 B.n39 585
R4 B.n328 B.n327 585
R5 B.n329 B.n38 585
R6 B.n331 B.n330 585
R7 B.n332 B.n37 585
R8 B.n334 B.n333 585
R9 B.n335 B.n36 585
R10 B.n337 B.n336 585
R11 B.n338 B.n35 585
R12 B.n340 B.n339 585
R13 B.n342 B.n341 585
R14 B.n343 B.n31 585
R15 B.n345 B.n344 585
R16 B.n346 B.n30 585
R17 B.n348 B.n347 585
R18 B.n349 B.n29 585
R19 B.n351 B.n350 585
R20 B.n352 B.n28 585
R21 B.n354 B.n353 585
R22 B.n356 B.n25 585
R23 B.n358 B.n357 585
R24 B.n359 B.n24 585
R25 B.n361 B.n360 585
R26 B.n362 B.n23 585
R27 B.n364 B.n363 585
R28 B.n365 B.n22 585
R29 B.n367 B.n366 585
R30 B.n368 B.n21 585
R31 B.n370 B.n369 585
R32 B.n371 B.n20 585
R33 B.n373 B.n372 585
R34 B.n374 B.n19 585
R35 B.n320 B.n41 585
R36 B.n319 B.n318 585
R37 B.n317 B.n42 585
R38 B.n316 B.n315 585
R39 B.n314 B.n43 585
R40 B.n313 B.n312 585
R41 B.n311 B.n44 585
R42 B.n310 B.n309 585
R43 B.n308 B.n45 585
R44 B.n307 B.n306 585
R45 B.n305 B.n46 585
R46 B.n304 B.n303 585
R47 B.n302 B.n47 585
R48 B.n301 B.n300 585
R49 B.n299 B.n48 585
R50 B.n298 B.n297 585
R51 B.n296 B.n49 585
R52 B.n295 B.n294 585
R53 B.n293 B.n50 585
R54 B.n292 B.n291 585
R55 B.n290 B.n51 585
R56 B.n289 B.n288 585
R57 B.n287 B.n52 585
R58 B.n286 B.n285 585
R59 B.n284 B.n53 585
R60 B.n283 B.n282 585
R61 B.n281 B.n54 585
R62 B.n280 B.n279 585
R63 B.n278 B.n55 585
R64 B.n277 B.n276 585
R65 B.n275 B.n56 585
R66 B.n274 B.n273 585
R67 B.n272 B.n57 585
R68 B.n271 B.n270 585
R69 B.n269 B.n58 585
R70 B.n268 B.n267 585
R71 B.n266 B.n59 585
R72 B.n265 B.n264 585
R73 B.n263 B.n60 585
R74 B.n262 B.n261 585
R75 B.n260 B.n61 585
R76 B.n259 B.n258 585
R77 B.n257 B.n62 585
R78 B.n256 B.n255 585
R79 B.n254 B.n63 585
R80 B.n253 B.n252 585
R81 B.n251 B.n64 585
R82 B.n250 B.n249 585
R83 B.n248 B.n65 585
R84 B.n247 B.n246 585
R85 B.n245 B.n66 585
R86 B.n244 B.n243 585
R87 B.n242 B.n67 585
R88 B.n241 B.n240 585
R89 B.n239 B.n68 585
R90 B.n238 B.n237 585
R91 B.n236 B.n69 585
R92 B.n235 B.n234 585
R93 B.n233 B.n70 585
R94 B.n232 B.n231 585
R95 B.n230 B.n71 585
R96 B.n229 B.n228 585
R97 B.n227 B.n72 585
R98 B.n226 B.n225 585
R99 B.n224 B.n73 585
R100 B.n223 B.n222 585
R101 B.n221 B.n74 585
R102 B.n220 B.n219 585
R103 B.n218 B.n75 585
R104 B.n164 B.n97 585
R105 B.n166 B.n165 585
R106 B.n167 B.n96 585
R107 B.n169 B.n168 585
R108 B.n170 B.n95 585
R109 B.n172 B.n171 585
R110 B.n173 B.n94 585
R111 B.n175 B.n174 585
R112 B.n176 B.n93 585
R113 B.n178 B.n177 585
R114 B.n179 B.n92 585
R115 B.n181 B.n180 585
R116 B.n182 B.n89 585
R117 B.n185 B.n184 585
R118 B.n186 B.n88 585
R119 B.n188 B.n187 585
R120 B.n189 B.n87 585
R121 B.n191 B.n190 585
R122 B.n192 B.n86 585
R123 B.n194 B.n193 585
R124 B.n195 B.n85 585
R125 B.n197 B.n196 585
R126 B.n199 B.n198 585
R127 B.n200 B.n81 585
R128 B.n202 B.n201 585
R129 B.n203 B.n80 585
R130 B.n205 B.n204 585
R131 B.n206 B.n79 585
R132 B.n208 B.n207 585
R133 B.n209 B.n78 585
R134 B.n211 B.n210 585
R135 B.n212 B.n77 585
R136 B.n214 B.n213 585
R137 B.n215 B.n76 585
R138 B.n217 B.n216 585
R139 B.n163 B.n162 585
R140 B.n161 B.n98 585
R141 B.n160 B.n159 585
R142 B.n158 B.n99 585
R143 B.n157 B.n156 585
R144 B.n155 B.n100 585
R145 B.n154 B.n153 585
R146 B.n152 B.n101 585
R147 B.n151 B.n150 585
R148 B.n149 B.n102 585
R149 B.n148 B.n147 585
R150 B.n146 B.n103 585
R151 B.n145 B.n144 585
R152 B.n143 B.n104 585
R153 B.n142 B.n141 585
R154 B.n140 B.n105 585
R155 B.n139 B.n138 585
R156 B.n137 B.n106 585
R157 B.n136 B.n135 585
R158 B.n134 B.n107 585
R159 B.n133 B.n132 585
R160 B.n131 B.n108 585
R161 B.n130 B.n129 585
R162 B.n128 B.n109 585
R163 B.n127 B.n126 585
R164 B.n125 B.n110 585
R165 B.n124 B.n123 585
R166 B.n122 B.n111 585
R167 B.n121 B.n120 585
R168 B.n119 B.n112 585
R169 B.n118 B.n117 585
R170 B.n116 B.n113 585
R171 B.n115 B.n114 585
R172 B.n2 B.n0 585
R173 B.n425 B.n1 585
R174 B.n424 B.n423 585
R175 B.n422 B.n3 585
R176 B.n421 B.n420 585
R177 B.n419 B.n4 585
R178 B.n418 B.n417 585
R179 B.n416 B.n5 585
R180 B.n415 B.n414 585
R181 B.n413 B.n6 585
R182 B.n412 B.n411 585
R183 B.n410 B.n7 585
R184 B.n409 B.n408 585
R185 B.n407 B.n8 585
R186 B.n406 B.n405 585
R187 B.n404 B.n9 585
R188 B.n403 B.n402 585
R189 B.n401 B.n10 585
R190 B.n400 B.n399 585
R191 B.n398 B.n11 585
R192 B.n397 B.n396 585
R193 B.n395 B.n12 585
R194 B.n394 B.n393 585
R195 B.n392 B.n13 585
R196 B.n391 B.n390 585
R197 B.n389 B.n14 585
R198 B.n388 B.n387 585
R199 B.n386 B.n15 585
R200 B.n385 B.n384 585
R201 B.n383 B.n16 585
R202 B.n382 B.n381 585
R203 B.n380 B.n17 585
R204 B.n379 B.n378 585
R205 B.n377 B.n18 585
R206 B.n376 B.n375 585
R207 B.n427 B.n426 585
R208 B.n162 B.n97 492.5
R209 B.n376 B.n19 492.5
R210 B.n216 B.n75 492.5
R211 B.n322 B.n41 492.5
R212 B.n82 B.t5 229.478
R213 B.n32 B.t7 229.478
R214 B.n90 B.t2 229.478
R215 B.n26 B.t10 229.478
R216 B.n82 B.t3 228.504
R217 B.n90 B.t0 228.504
R218 B.n26 B.t9 228.504
R219 B.n32 B.t6 228.504
R220 B.n83 B.t4 172.849
R221 B.n33 B.t8 172.849
R222 B.n91 B.t1 172.847
R223 B.n27 B.t11 172.847
R224 B.n162 B.n161 163.367
R225 B.n161 B.n160 163.367
R226 B.n160 B.n99 163.367
R227 B.n156 B.n99 163.367
R228 B.n156 B.n155 163.367
R229 B.n155 B.n154 163.367
R230 B.n154 B.n101 163.367
R231 B.n150 B.n101 163.367
R232 B.n150 B.n149 163.367
R233 B.n149 B.n148 163.367
R234 B.n148 B.n103 163.367
R235 B.n144 B.n103 163.367
R236 B.n144 B.n143 163.367
R237 B.n143 B.n142 163.367
R238 B.n142 B.n105 163.367
R239 B.n138 B.n105 163.367
R240 B.n138 B.n137 163.367
R241 B.n137 B.n136 163.367
R242 B.n136 B.n107 163.367
R243 B.n132 B.n107 163.367
R244 B.n132 B.n131 163.367
R245 B.n131 B.n130 163.367
R246 B.n130 B.n109 163.367
R247 B.n126 B.n109 163.367
R248 B.n126 B.n125 163.367
R249 B.n125 B.n124 163.367
R250 B.n124 B.n111 163.367
R251 B.n120 B.n111 163.367
R252 B.n120 B.n119 163.367
R253 B.n119 B.n118 163.367
R254 B.n118 B.n113 163.367
R255 B.n114 B.n113 163.367
R256 B.n114 B.n2 163.367
R257 B.n426 B.n2 163.367
R258 B.n426 B.n425 163.367
R259 B.n425 B.n424 163.367
R260 B.n424 B.n3 163.367
R261 B.n420 B.n3 163.367
R262 B.n420 B.n419 163.367
R263 B.n419 B.n418 163.367
R264 B.n418 B.n5 163.367
R265 B.n414 B.n5 163.367
R266 B.n414 B.n413 163.367
R267 B.n413 B.n412 163.367
R268 B.n412 B.n7 163.367
R269 B.n408 B.n7 163.367
R270 B.n408 B.n407 163.367
R271 B.n407 B.n406 163.367
R272 B.n406 B.n9 163.367
R273 B.n402 B.n9 163.367
R274 B.n402 B.n401 163.367
R275 B.n401 B.n400 163.367
R276 B.n400 B.n11 163.367
R277 B.n396 B.n11 163.367
R278 B.n396 B.n395 163.367
R279 B.n395 B.n394 163.367
R280 B.n394 B.n13 163.367
R281 B.n390 B.n13 163.367
R282 B.n390 B.n389 163.367
R283 B.n389 B.n388 163.367
R284 B.n388 B.n15 163.367
R285 B.n384 B.n15 163.367
R286 B.n384 B.n383 163.367
R287 B.n383 B.n382 163.367
R288 B.n382 B.n17 163.367
R289 B.n378 B.n17 163.367
R290 B.n378 B.n377 163.367
R291 B.n377 B.n376 163.367
R292 B.n166 B.n97 163.367
R293 B.n167 B.n166 163.367
R294 B.n168 B.n167 163.367
R295 B.n168 B.n95 163.367
R296 B.n172 B.n95 163.367
R297 B.n173 B.n172 163.367
R298 B.n174 B.n173 163.367
R299 B.n174 B.n93 163.367
R300 B.n178 B.n93 163.367
R301 B.n179 B.n178 163.367
R302 B.n180 B.n179 163.367
R303 B.n180 B.n89 163.367
R304 B.n185 B.n89 163.367
R305 B.n186 B.n185 163.367
R306 B.n187 B.n186 163.367
R307 B.n187 B.n87 163.367
R308 B.n191 B.n87 163.367
R309 B.n192 B.n191 163.367
R310 B.n193 B.n192 163.367
R311 B.n193 B.n85 163.367
R312 B.n197 B.n85 163.367
R313 B.n198 B.n197 163.367
R314 B.n198 B.n81 163.367
R315 B.n202 B.n81 163.367
R316 B.n203 B.n202 163.367
R317 B.n204 B.n203 163.367
R318 B.n204 B.n79 163.367
R319 B.n208 B.n79 163.367
R320 B.n209 B.n208 163.367
R321 B.n210 B.n209 163.367
R322 B.n210 B.n77 163.367
R323 B.n214 B.n77 163.367
R324 B.n215 B.n214 163.367
R325 B.n216 B.n215 163.367
R326 B.n220 B.n75 163.367
R327 B.n221 B.n220 163.367
R328 B.n222 B.n221 163.367
R329 B.n222 B.n73 163.367
R330 B.n226 B.n73 163.367
R331 B.n227 B.n226 163.367
R332 B.n228 B.n227 163.367
R333 B.n228 B.n71 163.367
R334 B.n232 B.n71 163.367
R335 B.n233 B.n232 163.367
R336 B.n234 B.n233 163.367
R337 B.n234 B.n69 163.367
R338 B.n238 B.n69 163.367
R339 B.n239 B.n238 163.367
R340 B.n240 B.n239 163.367
R341 B.n240 B.n67 163.367
R342 B.n244 B.n67 163.367
R343 B.n245 B.n244 163.367
R344 B.n246 B.n245 163.367
R345 B.n246 B.n65 163.367
R346 B.n250 B.n65 163.367
R347 B.n251 B.n250 163.367
R348 B.n252 B.n251 163.367
R349 B.n252 B.n63 163.367
R350 B.n256 B.n63 163.367
R351 B.n257 B.n256 163.367
R352 B.n258 B.n257 163.367
R353 B.n258 B.n61 163.367
R354 B.n262 B.n61 163.367
R355 B.n263 B.n262 163.367
R356 B.n264 B.n263 163.367
R357 B.n264 B.n59 163.367
R358 B.n268 B.n59 163.367
R359 B.n269 B.n268 163.367
R360 B.n270 B.n269 163.367
R361 B.n270 B.n57 163.367
R362 B.n274 B.n57 163.367
R363 B.n275 B.n274 163.367
R364 B.n276 B.n275 163.367
R365 B.n276 B.n55 163.367
R366 B.n280 B.n55 163.367
R367 B.n281 B.n280 163.367
R368 B.n282 B.n281 163.367
R369 B.n282 B.n53 163.367
R370 B.n286 B.n53 163.367
R371 B.n287 B.n286 163.367
R372 B.n288 B.n287 163.367
R373 B.n288 B.n51 163.367
R374 B.n292 B.n51 163.367
R375 B.n293 B.n292 163.367
R376 B.n294 B.n293 163.367
R377 B.n294 B.n49 163.367
R378 B.n298 B.n49 163.367
R379 B.n299 B.n298 163.367
R380 B.n300 B.n299 163.367
R381 B.n300 B.n47 163.367
R382 B.n304 B.n47 163.367
R383 B.n305 B.n304 163.367
R384 B.n306 B.n305 163.367
R385 B.n306 B.n45 163.367
R386 B.n310 B.n45 163.367
R387 B.n311 B.n310 163.367
R388 B.n312 B.n311 163.367
R389 B.n312 B.n43 163.367
R390 B.n316 B.n43 163.367
R391 B.n317 B.n316 163.367
R392 B.n318 B.n317 163.367
R393 B.n318 B.n41 163.367
R394 B.n372 B.n19 163.367
R395 B.n372 B.n371 163.367
R396 B.n371 B.n370 163.367
R397 B.n370 B.n21 163.367
R398 B.n366 B.n21 163.367
R399 B.n366 B.n365 163.367
R400 B.n365 B.n364 163.367
R401 B.n364 B.n23 163.367
R402 B.n360 B.n23 163.367
R403 B.n360 B.n359 163.367
R404 B.n359 B.n358 163.367
R405 B.n358 B.n25 163.367
R406 B.n353 B.n25 163.367
R407 B.n353 B.n352 163.367
R408 B.n352 B.n351 163.367
R409 B.n351 B.n29 163.367
R410 B.n347 B.n29 163.367
R411 B.n347 B.n346 163.367
R412 B.n346 B.n345 163.367
R413 B.n345 B.n31 163.367
R414 B.n341 B.n31 163.367
R415 B.n341 B.n340 163.367
R416 B.n340 B.n35 163.367
R417 B.n336 B.n35 163.367
R418 B.n336 B.n335 163.367
R419 B.n335 B.n334 163.367
R420 B.n334 B.n37 163.367
R421 B.n330 B.n37 163.367
R422 B.n330 B.n329 163.367
R423 B.n329 B.n328 163.367
R424 B.n328 B.n39 163.367
R425 B.n324 B.n39 163.367
R426 B.n324 B.n323 163.367
R427 B.n323 B.n322 163.367
R428 B.n84 B.n83 59.5399
R429 B.n183 B.n91 59.5399
R430 B.n355 B.n27 59.5399
R431 B.n34 B.n33 59.5399
R432 B.n83 B.n82 56.6308
R433 B.n91 B.n90 56.6308
R434 B.n27 B.n26 56.6308
R435 B.n33 B.n32 56.6308
R436 B.n375 B.n374 32.0005
R437 B.n321 B.n320 32.0005
R438 B.n218 B.n217 32.0005
R439 B.n164 B.n163 32.0005
R440 B B.n427 18.0485
R441 B.n374 B.n373 10.6151
R442 B.n373 B.n20 10.6151
R443 B.n369 B.n20 10.6151
R444 B.n369 B.n368 10.6151
R445 B.n368 B.n367 10.6151
R446 B.n367 B.n22 10.6151
R447 B.n363 B.n22 10.6151
R448 B.n363 B.n362 10.6151
R449 B.n362 B.n361 10.6151
R450 B.n361 B.n24 10.6151
R451 B.n357 B.n24 10.6151
R452 B.n357 B.n356 10.6151
R453 B.n354 B.n28 10.6151
R454 B.n350 B.n28 10.6151
R455 B.n350 B.n349 10.6151
R456 B.n349 B.n348 10.6151
R457 B.n348 B.n30 10.6151
R458 B.n344 B.n30 10.6151
R459 B.n344 B.n343 10.6151
R460 B.n343 B.n342 10.6151
R461 B.n339 B.n338 10.6151
R462 B.n338 B.n337 10.6151
R463 B.n337 B.n36 10.6151
R464 B.n333 B.n36 10.6151
R465 B.n333 B.n332 10.6151
R466 B.n332 B.n331 10.6151
R467 B.n331 B.n38 10.6151
R468 B.n327 B.n38 10.6151
R469 B.n327 B.n326 10.6151
R470 B.n326 B.n325 10.6151
R471 B.n325 B.n40 10.6151
R472 B.n321 B.n40 10.6151
R473 B.n219 B.n218 10.6151
R474 B.n219 B.n74 10.6151
R475 B.n223 B.n74 10.6151
R476 B.n224 B.n223 10.6151
R477 B.n225 B.n224 10.6151
R478 B.n225 B.n72 10.6151
R479 B.n229 B.n72 10.6151
R480 B.n230 B.n229 10.6151
R481 B.n231 B.n230 10.6151
R482 B.n231 B.n70 10.6151
R483 B.n235 B.n70 10.6151
R484 B.n236 B.n235 10.6151
R485 B.n237 B.n236 10.6151
R486 B.n237 B.n68 10.6151
R487 B.n241 B.n68 10.6151
R488 B.n242 B.n241 10.6151
R489 B.n243 B.n242 10.6151
R490 B.n243 B.n66 10.6151
R491 B.n247 B.n66 10.6151
R492 B.n248 B.n247 10.6151
R493 B.n249 B.n248 10.6151
R494 B.n249 B.n64 10.6151
R495 B.n253 B.n64 10.6151
R496 B.n254 B.n253 10.6151
R497 B.n255 B.n254 10.6151
R498 B.n255 B.n62 10.6151
R499 B.n259 B.n62 10.6151
R500 B.n260 B.n259 10.6151
R501 B.n261 B.n260 10.6151
R502 B.n261 B.n60 10.6151
R503 B.n265 B.n60 10.6151
R504 B.n266 B.n265 10.6151
R505 B.n267 B.n266 10.6151
R506 B.n267 B.n58 10.6151
R507 B.n271 B.n58 10.6151
R508 B.n272 B.n271 10.6151
R509 B.n273 B.n272 10.6151
R510 B.n273 B.n56 10.6151
R511 B.n277 B.n56 10.6151
R512 B.n278 B.n277 10.6151
R513 B.n279 B.n278 10.6151
R514 B.n279 B.n54 10.6151
R515 B.n283 B.n54 10.6151
R516 B.n284 B.n283 10.6151
R517 B.n285 B.n284 10.6151
R518 B.n285 B.n52 10.6151
R519 B.n289 B.n52 10.6151
R520 B.n290 B.n289 10.6151
R521 B.n291 B.n290 10.6151
R522 B.n291 B.n50 10.6151
R523 B.n295 B.n50 10.6151
R524 B.n296 B.n295 10.6151
R525 B.n297 B.n296 10.6151
R526 B.n297 B.n48 10.6151
R527 B.n301 B.n48 10.6151
R528 B.n302 B.n301 10.6151
R529 B.n303 B.n302 10.6151
R530 B.n303 B.n46 10.6151
R531 B.n307 B.n46 10.6151
R532 B.n308 B.n307 10.6151
R533 B.n309 B.n308 10.6151
R534 B.n309 B.n44 10.6151
R535 B.n313 B.n44 10.6151
R536 B.n314 B.n313 10.6151
R537 B.n315 B.n314 10.6151
R538 B.n315 B.n42 10.6151
R539 B.n319 B.n42 10.6151
R540 B.n320 B.n319 10.6151
R541 B.n165 B.n164 10.6151
R542 B.n165 B.n96 10.6151
R543 B.n169 B.n96 10.6151
R544 B.n170 B.n169 10.6151
R545 B.n171 B.n170 10.6151
R546 B.n171 B.n94 10.6151
R547 B.n175 B.n94 10.6151
R548 B.n176 B.n175 10.6151
R549 B.n177 B.n176 10.6151
R550 B.n177 B.n92 10.6151
R551 B.n181 B.n92 10.6151
R552 B.n182 B.n181 10.6151
R553 B.n184 B.n88 10.6151
R554 B.n188 B.n88 10.6151
R555 B.n189 B.n188 10.6151
R556 B.n190 B.n189 10.6151
R557 B.n190 B.n86 10.6151
R558 B.n194 B.n86 10.6151
R559 B.n195 B.n194 10.6151
R560 B.n196 B.n195 10.6151
R561 B.n200 B.n199 10.6151
R562 B.n201 B.n200 10.6151
R563 B.n201 B.n80 10.6151
R564 B.n205 B.n80 10.6151
R565 B.n206 B.n205 10.6151
R566 B.n207 B.n206 10.6151
R567 B.n207 B.n78 10.6151
R568 B.n211 B.n78 10.6151
R569 B.n212 B.n211 10.6151
R570 B.n213 B.n212 10.6151
R571 B.n213 B.n76 10.6151
R572 B.n217 B.n76 10.6151
R573 B.n163 B.n98 10.6151
R574 B.n159 B.n98 10.6151
R575 B.n159 B.n158 10.6151
R576 B.n158 B.n157 10.6151
R577 B.n157 B.n100 10.6151
R578 B.n153 B.n100 10.6151
R579 B.n153 B.n152 10.6151
R580 B.n152 B.n151 10.6151
R581 B.n151 B.n102 10.6151
R582 B.n147 B.n102 10.6151
R583 B.n147 B.n146 10.6151
R584 B.n146 B.n145 10.6151
R585 B.n145 B.n104 10.6151
R586 B.n141 B.n104 10.6151
R587 B.n141 B.n140 10.6151
R588 B.n140 B.n139 10.6151
R589 B.n139 B.n106 10.6151
R590 B.n135 B.n106 10.6151
R591 B.n135 B.n134 10.6151
R592 B.n134 B.n133 10.6151
R593 B.n133 B.n108 10.6151
R594 B.n129 B.n108 10.6151
R595 B.n129 B.n128 10.6151
R596 B.n128 B.n127 10.6151
R597 B.n127 B.n110 10.6151
R598 B.n123 B.n110 10.6151
R599 B.n123 B.n122 10.6151
R600 B.n122 B.n121 10.6151
R601 B.n121 B.n112 10.6151
R602 B.n117 B.n112 10.6151
R603 B.n117 B.n116 10.6151
R604 B.n116 B.n115 10.6151
R605 B.n115 B.n0 10.6151
R606 B.n423 B.n1 10.6151
R607 B.n423 B.n422 10.6151
R608 B.n422 B.n421 10.6151
R609 B.n421 B.n4 10.6151
R610 B.n417 B.n4 10.6151
R611 B.n417 B.n416 10.6151
R612 B.n416 B.n415 10.6151
R613 B.n415 B.n6 10.6151
R614 B.n411 B.n6 10.6151
R615 B.n411 B.n410 10.6151
R616 B.n410 B.n409 10.6151
R617 B.n409 B.n8 10.6151
R618 B.n405 B.n8 10.6151
R619 B.n405 B.n404 10.6151
R620 B.n404 B.n403 10.6151
R621 B.n403 B.n10 10.6151
R622 B.n399 B.n10 10.6151
R623 B.n399 B.n398 10.6151
R624 B.n398 B.n397 10.6151
R625 B.n397 B.n12 10.6151
R626 B.n393 B.n12 10.6151
R627 B.n393 B.n392 10.6151
R628 B.n392 B.n391 10.6151
R629 B.n391 B.n14 10.6151
R630 B.n387 B.n14 10.6151
R631 B.n387 B.n386 10.6151
R632 B.n386 B.n385 10.6151
R633 B.n385 B.n16 10.6151
R634 B.n381 B.n16 10.6151
R635 B.n381 B.n380 10.6151
R636 B.n380 B.n379 10.6151
R637 B.n379 B.n18 10.6151
R638 B.n375 B.n18 10.6151
R639 B.n355 B.n354 6.5566
R640 B.n342 B.n34 6.5566
R641 B.n184 B.n183 6.5566
R642 B.n196 B.n84 6.5566
R643 B.n356 B.n355 4.05904
R644 B.n339 B.n34 4.05904
R645 B.n183 B.n182 4.05904
R646 B.n199 B.n84 4.05904
R647 B.n427 B.n0 2.81026
R648 B.n427 B.n1 2.81026
R649 VP.n14 VP.n0 161.3
R650 VP.n13 VP.n12 161.3
R651 VP.n11 VP.n1 161.3
R652 VP.n10 VP.n9 161.3
R653 VP.n8 VP.n2 161.3
R654 VP.n7 VP.n6 161.3
R655 VP.n5 VP.n3 100.579
R656 VP.n16 VP.n15 100.579
R657 VP.n4 VP.t3 56.6708
R658 VP.n9 VP.n1 56.5617
R659 VP.n4 VP.t1 55.8963
R660 VP.n5 VP.n4 43.2062
R661 VP.n8 VP.n7 24.5923
R662 VP.n9 VP.n8 24.5923
R663 VP.n13 VP.n1 24.5923
R664 VP.n14 VP.n13 24.5923
R665 VP.n3 VP.t2 20.4715
R666 VP.n15 VP.t0 20.4715
R667 VP.n7 VP.n3 10.3291
R668 VP.n15 VP.n14 10.3291
R669 VP.n6 VP.n5 0.278335
R670 VP.n16 VP.n0 0.278335
R671 VP.n6 VP.n2 0.189894
R672 VP.n10 VP.n2 0.189894
R673 VP.n11 VP.n10 0.189894
R674 VP.n12 VP.n11 0.189894
R675 VP.n12 VP.n0 0.189894
R676 VP VP.n16 0.153485
R677 VTAIL.n7 VTAIL.t1 172.038
R678 VTAIL.n0 VTAIL.t3 172.038
R679 VTAIL.n1 VTAIL.t5 172.038
R680 VTAIL.n2 VTAIL.t7 172.038
R681 VTAIL.n6 VTAIL.t4 172.038
R682 VTAIL.n5 VTAIL.t6 172.038
R683 VTAIL.n4 VTAIL.t2 172.038
R684 VTAIL.n3 VTAIL.t0 172.038
R685 VTAIL.n7 VTAIL.n6 16.7807
R686 VTAIL.n3 VTAIL.n2 16.7807
R687 VTAIL.n4 VTAIL.n3 2.51774
R688 VTAIL.n6 VTAIL.n5 2.51774
R689 VTAIL.n2 VTAIL.n1 2.51774
R690 VTAIL VTAIL.n0 1.31731
R691 VTAIL VTAIL.n7 1.20093
R692 VTAIL.n5 VTAIL.n4 0.470328
R693 VTAIL.n1 VTAIL.n0 0.470328
R694 VDD1 VDD1.n1 207.631
R695 VDD1 VDD1.n0 174
R696 VDD1.n0 VDD1.t0 14.7755
R697 VDD1.n0 VDD1.t2 14.7755
R698 VDD1.n1 VDD1.t1 14.7755
R699 VDD1.n1 VDD1.t3 14.7755
R700 VN.n0 VN.t3 56.6708
R701 VN.n1 VN.t1 56.6708
R702 VN.n0 VN.t0 55.8963
R703 VN.n1 VN.t2 55.8963
R704 VN VN.n1 43.4851
R705 VN VN.n0 4.33734
R706 VDD2.n2 VDD2.n0 207.106
R707 VDD2.n2 VDD2.n1 173.942
R708 VDD2.n1 VDD2.t1 14.7755
R709 VDD2.n1 VDD2.t2 14.7755
R710 VDD2.n0 VDD2.t0 14.7755
R711 VDD2.n0 VDD2.t3 14.7755
R712 VDD2 VDD2.n2 0.0586897
C0 VTAIL B 1.63826f
C1 VTAIL VDD2 3.12526f
C2 VN w_n2722_n1408# 4.4011f
C3 w_n2722_n1408# VP 4.74707f
C4 VN VDD1 0.155023f
C5 w_n2722_n1408# B 6.51749f
C6 VDD1 VP 1.37563f
C7 VDD2 w_n2722_n1408# 1.24177f
C8 VDD1 B 0.99411f
C9 VDD2 VDD1 1.01803f
C10 VN VP 4.37078f
C11 VTAIL w_n2722_n1408# 1.72766f
C12 VN B 0.974517f
C13 VTAIL VDD1 3.07112f
C14 VDD2 VN 1.13181f
C15 B VP 1.55444f
C16 VDD2 VP 0.400527f
C17 VDD2 B 1.04641f
C18 VTAIL VN 1.67477f
C19 VDD1 w_n2722_n1408# 1.18657f
C20 VTAIL VP 1.68888f
C21 VDD2 VSUBS 0.66324f
C22 VDD1 VSUBS 3.355631f
C23 VTAIL VSUBS 0.428256f
C24 VN VSUBS 4.99758f
C25 VP VSUBS 1.743651f
C26 B VSUBS 3.249855f
C27 w_n2722_n1408# VSUBS 48.8327f
C28 VDD2.t0 VSUBS 0.036523f
C29 VDD2.t3 VSUBS 0.036523f
C30 VDD2.n0 VSUBS 0.307193f
C31 VDD2.t1 VSUBS 0.036523f
C32 VDD2.t2 VSUBS 0.036523f
C33 VDD2.n1 VSUBS 0.167904f
C34 VDD2.n2 VSUBS 2.30389f
C35 VN.t3 VSUBS 0.916773f
C36 VN.t0 VSUBS 0.909555f
C37 VN.n0 VSUBS 0.570062f
C38 VN.t1 VSUBS 0.916773f
C39 VN.t2 VSUBS 0.909555f
C40 VN.n1 VSUBS 2.35629f
C41 VDD1.t0 VSUBS 0.035631f
C42 VDD1.t2 VSUBS 0.035631f
C43 VDD1.n0 VSUBS 0.163939f
C44 VDD1.t1 VSUBS 0.035631f
C45 VDD1.t3 VSUBS 0.035631f
C46 VDD1.n1 VSUBS 0.308233f
C47 VTAIL.t3 VSUBS 0.183854f
C48 VTAIL.n0 VSUBS 0.299679f
C49 VTAIL.t5 VSUBS 0.183854f
C50 VTAIL.n1 VSUBS 0.365942f
C51 VTAIL.t7 VSUBS 0.183854f
C52 VTAIL.n2 VSUBS 0.81635f
C53 VTAIL.t0 VSUBS 0.183855f
C54 VTAIL.n3 VSUBS 0.816349f
C55 VTAIL.t2 VSUBS 0.183855f
C56 VTAIL.n4 VSUBS 0.365942f
C57 VTAIL.t6 VSUBS 0.183855f
C58 VTAIL.n5 VSUBS 0.365942f
C59 VTAIL.t4 VSUBS 0.183854f
C60 VTAIL.n6 VSUBS 0.81635f
C61 VTAIL.t1 VSUBS 0.183854f
C62 VTAIL.n7 VSUBS 0.743663f
C63 VP.n0 VSUBS 0.058127f
C64 VP.t0 VSUBS 0.597393f
C65 VP.n1 VSUBS 0.064094f
C66 VP.n2 VSUBS 0.044091f
C67 VP.t2 VSUBS 0.597393f
C68 VP.n3 VSUBS 0.422219f
C69 VP.t1 VSUBS 0.946969f
C70 VP.t3 VSUBS 0.954484f
C71 VP.n4 VSUBS 2.42958f
C72 VP.n5 VSUBS 1.90012f
C73 VP.n6 VSUBS 0.058127f
C74 VP.n7 VSUBS 0.058352f
C75 VP.n8 VSUBS 0.081763f
C76 VP.n9 VSUBS 0.064094f
C77 VP.n10 VSUBS 0.044091f
C78 VP.n11 VSUBS 0.044091f
C79 VP.n12 VSUBS 0.044091f
C80 VP.n13 VSUBS 0.081763f
C81 VP.n14 VSUBS 0.058352f
C82 VP.n15 VSUBS 0.422219f
C83 VP.n16 VSUBS 0.071231f
C84 B.n0 VSUBS 0.005519f
C85 B.n1 VSUBS 0.005519f
C86 B.n2 VSUBS 0.008728f
C87 B.n3 VSUBS 0.008728f
C88 B.n4 VSUBS 0.008728f
C89 B.n5 VSUBS 0.008728f
C90 B.n6 VSUBS 0.008728f
C91 B.n7 VSUBS 0.008728f
C92 B.n8 VSUBS 0.008728f
C93 B.n9 VSUBS 0.008728f
C94 B.n10 VSUBS 0.008728f
C95 B.n11 VSUBS 0.008728f
C96 B.n12 VSUBS 0.008728f
C97 B.n13 VSUBS 0.008728f
C98 B.n14 VSUBS 0.008728f
C99 B.n15 VSUBS 0.008728f
C100 B.n16 VSUBS 0.008728f
C101 B.n17 VSUBS 0.008728f
C102 B.n18 VSUBS 0.008728f
C103 B.n19 VSUBS 0.020472f
C104 B.n20 VSUBS 0.008728f
C105 B.n21 VSUBS 0.008728f
C106 B.n22 VSUBS 0.008728f
C107 B.n23 VSUBS 0.008728f
C108 B.n24 VSUBS 0.008728f
C109 B.n25 VSUBS 0.008728f
C110 B.t11 VSUBS 0.06048f
C111 B.t10 VSUBS 0.075867f
C112 B.t9 VSUBS 0.34898f
C113 B.n26 VSUBS 0.091719f
C114 B.n27 VSUBS 0.074799f
C115 B.n28 VSUBS 0.008728f
C116 B.n29 VSUBS 0.008728f
C117 B.n30 VSUBS 0.008728f
C118 B.n31 VSUBS 0.008728f
C119 B.t8 VSUBS 0.06048f
C120 B.t7 VSUBS 0.075867f
C121 B.t6 VSUBS 0.34898f
C122 B.n32 VSUBS 0.091719f
C123 B.n33 VSUBS 0.074799f
C124 B.n34 VSUBS 0.020221f
C125 B.n35 VSUBS 0.008728f
C126 B.n36 VSUBS 0.008728f
C127 B.n37 VSUBS 0.008728f
C128 B.n38 VSUBS 0.008728f
C129 B.n39 VSUBS 0.008728f
C130 B.n40 VSUBS 0.008728f
C131 B.n41 VSUBS 0.01983f
C132 B.n42 VSUBS 0.008728f
C133 B.n43 VSUBS 0.008728f
C134 B.n44 VSUBS 0.008728f
C135 B.n45 VSUBS 0.008728f
C136 B.n46 VSUBS 0.008728f
C137 B.n47 VSUBS 0.008728f
C138 B.n48 VSUBS 0.008728f
C139 B.n49 VSUBS 0.008728f
C140 B.n50 VSUBS 0.008728f
C141 B.n51 VSUBS 0.008728f
C142 B.n52 VSUBS 0.008728f
C143 B.n53 VSUBS 0.008728f
C144 B.n54 VSUBS 0.008728f
C145 B.n55 VSUBS 0.008728f
C146 B.n56 VSUBS 0.008728f
C147 B.n57 VSUBS 0.008728f
C148 B.n58 VSUBS 0.008728f
C149 B.n59 VSUBS 0.008728f
C150 B.n60 VSUBS 0.008728f
C151 B.n61 VSUBS 0.008728f
C152 B.n62 VSUBS 0.008728f
C153 B.n63 VSUBS 0.008728f
C154 B.n64 VSUBS 0.008728f
C155 B.n65 VSUBS 0.008728f
C156 B.n66 VSUBS 0.008728f
C157 B.n67 VSUBS 0.008728f
C158 B.n68 VSUBS 0.008728f
C159 B.n69 VSUBS 0.008728f
C160 B.n70 VSUBS 0.008728f
C161 B.n71 VSUBS 0.008728f
C162 B.n72 VSUBS 0.008728f
C163 B.n73 VSUBS 0.008728f
C164 B.n74 VSUBS 0.008728f
C165 B.n75 VSUBS 0.01983f
C166 B.n76 VSUBS 0.008728f
C167 B.n77 VSUBS 0.008728f
C168 B.n78 VSUBS 0.008728f
C169 B.n79 VSUBS 0.008728f
C170 B.n80 VSUBS 0.008728f
C171 B.n81 VSUBS 0.008728f
C172 B.t4 VSUBS 0.06048f
C173 B.t5 VSUBS 0.075867f
C174 B.t3 VSUBS 0.34898f
C175 B.n82 VSUBS 0.091719f
C176 B.n83 VSUBS 0.074799f
C177 B.n84 VSUBS 0.020221f
C178 B.n85 VSUBS 0.008728f
C179 B.n86 VSUBS 0.008728f
C180 B.n87 VSUBS 0.008728f
C181 B.n88 VSUBS 0.008728f
C182 B.n89 VSUBS 0.008728f
C183 B.t1 VSUBS 0.06048f
C184 B.t2 VSUBS 0.075867f
C185 B.t0 VSUBS 0.34898f
C186 B.n90 VSUBS 0.091719f
C187 B.n91 VSUBS 0.074799f
C188 B.n92 VSUBS 0.008728f
C189 B.n93 VSUBS 0.008728f
C190 B.n94 VSUBS 0.008728f
C191 B.n95 VSUBS 0.008728f
C192 B.n96 VSUBS 0.008728f
C193 B.n97 VSUBS 0.020472f
C194 B.n98 VSUBS 0.008728f
C195 B.n99 VSUBS 0.008728f
C196 B.n100 VSUBS 0.008728f
C197 B.n101 VSUBS 0.008728f
C198 B.n102 VSUBS 0.008728f
C199 B.n103 VSUBS 0.008728f
C200 B.n104 VSUBS 0.008728f
C201 B.n105 VSUBS 0.008728f
C202 B.n106 VSUBS 0.008728f
C203 B.n107 VSUBS 0.008728f
C204 B.n108 VSUBS 0.008728f
C205 B.n109 VSUBS 0.008728f
C206 B.n110 VSUBS 0.008728f
C207 B.n111 VSUBS 0.008728f
C208 B.n112 VSUBS 0.008728f
C209 B.n113 VSUBS 0.008728f
C210 B.n114 VSUBS 0.008728f
C211 B.n115 VSUBS 0.008728f
C212 B.n116 VSUBS 0.008728f
C213 B.n117 VSUBS 0.008728f
C214 B.n118 VSUBS 0.008728f
C215 B.n119 VSUBS 0.008728f
C216 B.n120 VSUBS 0.008728f
C217 B.n121 VSUBS 0.008728f
C218 B.n122 VSUBS 0.008728f
C219 B.n123 VSUBS 0.008728f
C220 B.n124 VSUBS 0.008728f
C221 B.n125 VSUBS 0.008728f
C222 B.n126 VSUBS 0.008728f
C223 B.n127 VSUBS 0.008728f
C224 B.n128 VSUBS 0.008728f
C225 B.n129 VSUBS 0.008728f
C226 B.n130 VSUBS 0.008728f
C227 B.n131 VSUBS 0.008728f
C228 B.n132 VSUBS 0.008728f
C229 B.n133 VSUBS 0.008728f
C230 B.n134 VSUBS 0.008728f
C231 B.n135 VSUBS 0.008728f
C232 B.n136 VSUBS 0.008728f
C233 B.n137 VSUBS 0.008728f
C234 B.n138 VSUBS 0.008728f
C235 B.n139 VSUBS 0.008728f
C236 B.n140 VSUBS 0.008728f
C237 B.n141 VSUBS 0.008728f
C238 B.n142 VSUBS 0.008728f
C239 B.n143 VSUBS 0.008728f
C240 B.n144 VSUBS 0.008728f
C241 B.n145 VSUBS 0.008728f
C242 B.n146 VSUBS 0.008728f
C243 B.n147 VSUBS 0.008728f
C244 B.n148 VSUBS 0.008728f
C245 B.n149 VSUBS 0.008728f
C246 B.n150 VSUBS 0.008728f
C247 B.n151 VSUBS 0.008728f
C248 B.n152 VSUBS 0.008728f
C249 B.n153 VSUBS 0.008728f
C250 B.n154 VSUBS 0.008728f
C251 B.n155 VSUBS 0.008728f
C252 B.n156 VSUBS 0.008728f
C253 B.n157 VSUBS 0.008728f
C254 B.n158 VSUBS 0.008728f
C255 B.n159 VSUBS 0.008728f
C256 B.n160 VSUBS 0.008728f
C257 B.n161 VSUBS 0.008728f
C258 B.n162 VSUBS 0.01983f
C259 B.n163 VSUBS 0.01983f
C260 B.n164 VSUBS 0.020472f
C261 B.n165 VSUBS 0.008728f
C262 B.n166 VSUBS 0.008728f
C263 B.n167 VSUBS 0.008728f
C264 B.n168 VSUBS 0.008728f
C265 B.n169 VSUBS 0.008728f
C266 B.n170 VSUBS 0.008728f
C267 B.n171 VSUBS 0.008728f
C268 B.n172 VSUBS 0.008728f
C269 B.n173 VSUBS 0.008728f
C270 B.n174 VSUBS 0.008728f
C271 B.n175 VSUBS 0.008728f
C272 B.n176 VSUBS 0.008728f
C273 B.n177 VSUBS 0.008728f
C274 B.n178 VSUBS 0.008728f
C275 B.n179 VSUBS 0.008728f
C276 B.n180 VSUBS 0.008728f
C277 B.n181 VSUBS 0.008728f
C278 B.n182 VSUBS 0.006032f
C279 B.n183 VSUBS 0.020221f
C280 B.n184 VSUBS 0.007059f
C281 B.n185 VSUBS 0.008728f
C282 B.n186 VSUBS 0.008728f
C283 B.n187 VSUBS 0.008728f
C284 B.n188 VSUBS 0.008728f
C285 B.n189 VSUBS 0.008728f
C286 B.n190 VSUBS 0.008728f
C287 B.n191 VSUBS 0.008728f
C288 B.n192 VSUBS 0.008728f
C289 B.n193 VSUBS 0.008728f
C290 B.n194 VSUBS 0.008728f
C291 B.n195 VSUBS 0.008728f
C292 B.n196 VSUBS 0.007059f
C293 B.n197 VSUBS 0.008728f
C294 B.n198 VSUBS 0.008728f
C295 B.n199 VSUBS 0.006032f
C296 B.n200 VSUBS 0.008728f
C297 B.n201 VSUBS 0.008728f
C298 B.n202 VSUBS 0.008728f
C299 B.n203 VSUBS 0.008728f
C300 B.n204 VSUBS 0.008728f
C301 B.n205 VSUBS 0.008728f
C302 B.n206 VSUBS 0.008728f
C303 B.n207 VSUBS 0.008728f
C304 B.n208 VSUBS 0.008728f
C305 B.n209 VSUBS 0.008728f
C306 B.n210 VSUBS 0.008728f
C307 B.n211 VSUBS 0.008728f
C308 B.n212 VSUBS 0.008728f
C309 B.n213 VSUBS 0.008728f
C310 B.n214 VSUBS 0.008728f
C311 B.n215 VSUBS 0.008728f
C312 B.n216 VSUBS 0.020472f
C313 B.n217 VSUBS 0.020472f
C314 B.n218 VSUBS 0.01983f
C315 B.n219 VSUBS 0.008728f
C316 B.n220 VSUBS 0.008728f
C317 B.n221 VSUBS 0.008728f
C318 B.n222 VSUBS 0.008728f
C319 B.n223 VSUBS 0.008728f
C320 B.n224 VSUBS 0.008728f
C321 B.n225 VSUBS 0.008728f
C322 B.n226 VSUBS 0.008728f
C323 B.n227 VSUBS 0.008728f
C324 B.n228 VSUBS 0.008728f
C325 B.n229 VSUBS 0.008728f
C326 B.n230 VSUBS 0.008728f
C327 B.n231 VSUBS 0.008728f
C328 B.n232 VSUBS 0.008728f
C329 B.n233 VSUBS 0.008728f
C330 B.n234 VSUBS 0.008728f
C331 B.n235 VSUBS 0.008728f
C332 B.n236 VSUBS 0.008728f
C333 B.n237 VSUBS 0.008728f
C334 B.n238 VSUBS 0.008728f
C335 B.n239 VSUBS 0.008728f
C336 B.n240 VSUBS 0.008728f
C337 B.n241 VSUBS 0.008728f
C338 B.n242 VSUBS 0.008728f
C339 B.n243 VSUBS 0.008728f
C340 B.n244 VSUBS 0.008728f
C341 B.n245 VSUBS 0.008728f
C342 B.n246 VSUBS 0.008728f
C343 B.n247 VSUBS 0.008728f
C344 B.n248 VSUBS 0.008728f
C345 B.n249 VSUBS 0.008728f
C346 B.n250 VSUBS 0.008728f
C347 B.n251 VSUBS 0.008728f
C348 B.n252 VSUBS 0.008728f
C349 B.n253 VSUBS 0.008728f
C350 B.n254 VSUBS 0.008728f
C351 B.n255 VSUBS 0.008728f
C352 B.n256 VSUBS 0.008728f
C353 B.n257 VSUBS 0.008728f
C354 B.n258 VSUBS 0.008728f
C355 B.n259 VSUBS 0.008728f
C356 B.n260 VSUBS 0.008728f
C357 B.n261 VSUBS 0.008728f
C358 B.n262 VSUBS 0.008728f
C359 B.n263 VSUBS 0.008728f
C360 B.n264 VSUBS 0.008728f
C361 B.n265 VSUBS 0.008728f
C362 B.n266 VSUBS 0.008728f
C363 B.n267 VSUBS 0.008728f
C364 B.n268 VSUBS 0.008728f
C365 B.n269 VSUBS 0.008728f
C366 B.n270 VSUBS 0.008728f
C367 B.n271 VSUBS 0.008728f
C368 B.n272 VSUBS 0.008728f
C369 B.n273 VSUBS 0.008728f
C370 B.n274 VSUBS 0.008728f
C371 B.n275 VSUBS 0.008728f
C372 B.n276 VSUBS 0.008728f
C373 B.n277 VSUBS 0.008728f
C374 B.n278 VSUBS 0.008728f
C375 B.n279 VSUBS 0.008728f
C376 B.n280 VSUBS 0.008728f
C377 B.n281 VSUBS 0.008728f
C378 B.n282 VSUBS 0.008728f
C379 B.n283 VSUBS 0.008728f
C380 B.n284 VSUBS 0.008728f
C381 B.n285 VSUBS 0.008728f
C382 B.n286 VSUBS 0.008728f
C383 B.n287 VSUBS 0.008728f
C384 B.n288 VSUBS 0.008728f
C385 B.n289 VSUBS 0.008728f
C386 B.n290 VSUBS 0.008728f
C387 B.n291 VSUBS 0.008728f
C388 B.n292 VSUBS 0.008728f
C389 B.n293 VSUBS 0.008728f
C390 B.n294 VSUBS 0.008728f
C391 B.n295 VSUBS 0.008728f
C392 B.n296 VSUBS 0.008728f
C393 B.n297 VSUBS 0.008728f
C394 B.n298 VSUBS 0.008728f
C395 B.n299 VSUBS 0.008728f
C396 B.n300 VSUBS 0.008728f
C397 B.n301 VSUBS 0.008728f
C398 B.n302 VSUBS 0.008728f
C399 B.n303 VSUBS 0.008728f
C400 B.n304 VSUBS 0.008728f
C401 B.n305 VSUBS 0.008728f
C402 B.n306 VSUBS 0.008728f
C403 B.n307 VSUBS 0.008728f
C404 B.n308 VSUBS 0.008728f
C405 B.n309 VSUBS 0.008728f
C406 B.n310 VSUBS 0.008728f
C407 B.n311 VSUBS 0.008728f
C408 B.n312 VSUBS 0.008728f
C409 B.n313 VSUBS 0.008728f
C410 B.n314 VSUBS 0.008728f
C411 B.n315 VSUBS 0.008728f
C412 B.n316 VSUBS 0.008728f
C413 B.n317 VSUBS 0.008728f
C414 B.n318 VSUBS 0.008728f
C415 B.n319 VSUBS 0.008728f
C416 B.n320 VSUBS 0.020883f
C417 B.n321 VSUBS 0.019419f
C418 B.n322 VSUBS 0.020472f
C419 B.n323 VSUBS 0.008728f
C420 B.n324 VSUBS 0.008728f
C421 B.n325 VSUBS 0.008728f
C422 B.n326 VSUBS 0.008728f
C423 B.n327 VSUBS 0.008728f
C424 B.n328 VSUBS 0.008728f
C425 B.n329 VSUBS 0.008728f
C426 B.n330 VSUBS 0.008728f
C427 B.n331 VSUBS 0.008728f
C428 B.n332 VSUBS 0.008728f
C429 B.n333 VSUBS 0.008728f
C430 B.n334 VSUBS 0.008728f
C431 B.n335 VSUBS 0.008728f
C432 B.n336 VSUBS 0.008728f
C433 B.n337 VSUBS 0.008728f
C434 B.n338 VSUBS 0.008728f
C435 B.n339 VSUBS 0.006032f
C436 B.n340 VSUBS 0.008728f
C437 B.n341 VSUBS 0.008728f
C438 B.n342 VSUBS 0.007059f
C439 B.n343 VSUBS 0.008728f
C440 B.n344 VSUBS 0.008728f
C441 B.n345 VSUBS 0.008728f
C442 B.n346 VSUBS 0.008728f
C443 B.n347 VSUBS 0.008728f
C444 B.n348 VSUBS 0.008728f
C445 B.n349 VSUBS 0.008728f
C446 B.n350 VSUBS 0.008728f
C447 B.n351 VSUBS 0.008728f
C448 B.n352 VSUBS 0.008728f
C449 B.n353 VSUBS 0.008728f
C450 B.n354 VSUBS 0.007059f
C451 B.n355 VSUBS 0.020221f
C452 B.n356 VSUBS 0.006032f
C453 B.n357 VSUBS 0.008728f
C454 B.n358 VSUBS 0.008728f
C455 B.n359 VSUBS 0.008728f
C456 B.n360 VSUBS 0.008728f
C457 B.n361 VSUBS 0.008728f
C458 B.n362 VSUBS 0.008728f
C459 B.n363 VSUBS 0.008728f
C460 B.n364 VSUBS 0.008728f
C461 B.n365 VSUBS 0.008728f
C462 B.n366 VSUBS 0.008728f
C463 B.n367 VSUBS 0.008728f
C464 B.n368 VSUBS 0.008728f
C465 B.n369 VSUBS 0.008728f
C466 B.n370 VSUBS 0.008728f
C467 B.n371 VSUBS 0.008728f
C468 B.n372 VSUBS 0.008728f
C469 B.n373 VSUBS 0.008728f
C470 B.n374 VSUBS 0.020472f
C471 B.n375 VSUBS 0.01983f
C472 B.n376 VSUBS 0.01983f
C473 B.n377 VSUBS 0.008728f
C474 B.n378 VSUBS 0.008728f
C475 B.n379 VSUBS 0.008728f
C476 B.n380 VSUBS 0.008728f
C477 B.n381 VSUBS 0.008728f
C478 B.n382 VSUBS 0.008728f
C479 B.n383 VSUBS 0.008728f
C480 B.n384 VSUBS 0.008728f
C481 B.n385 VSUBS 0.008728f
C482 B.n386 VSUBS 0.008728f
C483 B.n387 VSUBS 0.008728f
C484 B.n388 VSUBS 0.008728f
C485 B.n389 VSUBS 0.008728f
C486 B.n390 VSUBS 0.008728f
C487 B.n391 VSUBS 0.008728f
C488 B.n392 VSUBS 0.008728f
C489 B.n393 VSUBS 0.008728f
C490 B.n394 VSUBS 0.008728f
C491 B.n395 VSUBS 0.008728f
C492 B.n396 VSUBS 0.008728f
C493 B.n397 VSUBS 0.008728f
C494 B.n398 VSUBS 0.008728f
C495 B.n399 VSUBS 0.008728f
C496 B.n400 VSUBS 0.008728f
C497 B.n401 VSUBS 0.008728f
C498 B.n402 VSUBS 0.008728f
C499 B.n403 VSUBS 0.008728f
C500 B.n404 VSUBS 0.008728f
C501 B.n405 VSUBS 0.008728f
C502 B.n406 VSUBS 0.008728f
C503 B.n407 VSUBS 0.008728f
C504 B.n408 VSUBS 0.008728f
C505 B.n409 VSUBS 0.008728f
C506 B.n410 VSUBS 0.008728f
C507 B.n411 VSUBS 0.008728f
C508 B.n412 VSUBS 0.008728f
C509 B.n413 VSUBS 0.008728f
C510 B.n414 VSUBS 0.008728f
C511 B.n415 VSUBS 0.008728f
C512 B.n416 VSUBS 0.008728f
C513 B.n417 VSUBS 0.008728f
C514 B.n418 VSUBS 0.008728f
C515 B.n419 VSUBS 0.008728f
C516 B.n420 VSUBS 0.008728f
C517 B.n421 VSUBS 0.008728f
C518 B.n422 VSUBS 0.008728f
C519 B.n423 VSUBS 0.008728f
C520 B.n424 VSUBS 0.008728f
C521 B.n425 VSUBS 0.008728f
C522 B.n426 VSUBS 0.008728f
C523 B.n427 VSUBS 0.019763f
.ends

