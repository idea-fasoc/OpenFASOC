* NGSPICE file created from diff_pair_sample_1016.ext - technology: sky130A

.subckt diff_pair_sample_1016 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.7176 pd=4.46 as=0.3036 ps=2.17 w=1.84 l=1.82
X1 VTAIL.t14 VP.t1 VDD1.t5 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.3036 ps=2.17 w=1.84 l=1.82
X2 B.t11 B.t9 B.t10 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.7176 pd=4.46 as=0 ps=0 w=1.84 l=1.82
X3 VTAIL.t3 VN.t0 VDD2.t7 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.7176 pd=4.46 as=0.3036 ps=2.17 w=1.84 l=1.82
X4 VDD2.t6 VN.t1 VTAIL.t1 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.7176 ps=4.46 w=1.84 l=1.82
X5 B.t8 B.t6 B.t7 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.7176 pd=4.46 as=0 ps=0 w=1.84 l=1.82
X6 VDD2.t5 VN.t2 VTAIL.t2 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.3036 ps=2.17 w=1.84 l=1.82
X7 B.t5 B.t3 B.t4 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.7176 pd=4.46 as=0 ps=0 w=1.84 l=1.82
X8 VTAIL.t5 VN.t3 VDD2.t4 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.3036 ps=2.17 w=1.84 l=1.82
X9 VTAIL.t6 VN.t4 VDD2.t3 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.3036 ps=2.17 w=1.84 l=1.82
X10 VDD2.t2 VN.t5 VTAIL.t7 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.7176 ps=4.46 w=1.84 l=1.82
X11 VTAIL.t13 VP.t2 VDD1.t2 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.3036 ps=2.17 w=1.84 l=1.82
X12 VTAIL.t12 VP.t3 VDD1.t0 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.7176 pd=4.46 as=0.3036 ps=2.17 w=1.84 l=1.82
X13 VDD2.t1 VN.t6 VTAIL.t0 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.3036 ps=2.17 w=1.84 l=1.82
X14 VDD1.t1 VP.t4 VTAIL.t11 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.7176 ps=4.46 w=1.84 l=1.82
X15 VDD1.t3 VP.t5 VTAIL.t10 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.3036 ps=2.17 w=1.84 l=1.82
X16 VTAIL.t4 VN.t7 VDD2.t0 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.7176 pd=4.46 as=0.3036 ps=2.17 w=1.84 l=1.82
X17 VDD1.t4 VP.t6 VTAIL.t9 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.7176 ps=4.46 w=1.84 l=1.82
X18 VDD1.t6 VP.t7 VTAIL.t8 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.3036 pd=2.17 as=0.3036 ps=2.17 w=1.84 l=1.82
X19 B.t2 B.t0 B.t1 w_n3120_n1336# sky130_fd_pr__pfet_01v8 ad=0.7176 pd=4.46 as=0 ps=0 w=1.84 l=1.82
R0 VP.n13 VP.n12 161.3
R1 VP.n14 VP.n9 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n17 VP.n8 161.3
R4 VP.n20 VP.n19 161.3
R5 VP.n21 VP.n7 161.3
R6 VP.n23 VP.n22 161.3
R7 VP.n24 VP.n6 161.3
R8 VP.n48 VP.n0 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n45 VP.n1 161.3
R11 VP.n44 VP.n43 161.3
R12 VP.n41 VP.n2 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n3 161.3
R15 VP.n37 VP.n36 161.3
R16 VP.n34 VP.n4 161.3
R17 VP.n33 VP.n32 161.3
R18 VP.n31 VP.n5 161.3
R19 VP.n30 VP.n29 161.3
R20 VP.n28 VP.n27 87.546
R21 VP.n50 VP.n49 87.546
R22 VP.n26 VP.n25 87.546
R23 VP.n40 VP.n3 56.5617
R24 VP.n16 VP.n9 56.5617
R25 VP.n10 VP.t3 55.8733
R26 VP.n11 VP.n10 54.0319
R27 VP.n33 VP.n5 50.2647
R28 VP.n47 VP.n1 50.2647
R29 VP.n23 VP.n7 50.2647
R30 VP.n27 VP.n26 39.583
R31 VP.n29 VP.n5 30.8893
R32 VP.n48 VP.n47 30.8893
R33 VP.n24 VP.n23 30.8893
R34 VP.n34 VP.n33 24.5923
R35 VP.n36 VP.n3 24.5923
R36 VP.n41 VP.n40 24.5923
R37 VP.n43 VP.n1 24.5923
R38 VP.n17 VP.n16 24.5923
R39 VP.n19 VP.n7 24.5923
R40 VP.n12 VP.n9 24.5923
R41 VP.n28 VP.t0 24.3653
R42 VP.n35 VP.t7 24.3653
R43 VP.n42 VP.t1 24.3653
R44 VP.n49 VP.t6 24.3653
R45 VP.n25 VP.t4 24.3653
R46 VP.n18 VP.t2 24.3653
R47 VP.n11 VP.t5 24.3653
R48 VP.n29 VP.n28 23.3627
R49 VP.n49 VP.n48 23.3627
R50 VP.n25 VP.n24 23.3627
R51 VP.n36 VP.n35 15.9852
R52 VP.n42 VP.n41 15.9852
R53 VP.n18 VP.n17 15.9852
R54 VP.n12 VP.n11 15.9852
R55 VP.n13 VP.n10 12.7521
R56 VP.n35 VP.n34 8.60764
R57 VP.n43 VP.n42 8.60764
R58 VP.n19 VP.n18 8.60764
R59 VP.n26 VP.n6 0.278335
R60 VP.n30 VP.n27 0.278335
R61 VP.n50 VP.n0 0.278335
R62 VP.n14 VP.n13 0.189894
R63 VP.n15 VP.n14 0.189894
R64 VP.n15 VP.n8 0.189894
R65 VP.n20 VP.n8 0.189894
R66 VP.n21 VP.n20 0.189894
R67 VP.n22 VP.n21 0.189894
R68 VP.n22 VP.n6 0.189894
R69 VP.n31 VP.n30 0.189894
R70 VP.n32 VP.n31 0.189894
R71 VP.n32 VP.n4 0.189894
R72 VP.n37 VP.n4 0.189894
R73 VP.n38 VP.n37 0.189894
R74 VP.n39 VP.n38 0.189894
R75 VP.n39 VP.n2 0.189894
R76 VP.n44 VP.n2 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n46 VP.n45 0.189894
R79 VP.n46 VP.n0 0.189894
R80 VP VP.n50 0.153485
R81 VDD1 VDD1.n0 203.647
R82 VDD1.n3 VDD1.n2 203.534
R83 VDD1.n3 VDD1.n1 203.534
R84 VDD1.n5 VDD1.n4 202.661
R85 VDD1.n5 VDD1.n3 34.225
R86 VDD1.n4 VDD1.t2 17.6663
R87 VDD1.n4 VDD1.t1 17.6663
R88 VDD1.n0 VDD1.t0 17.6663
R89 VDD1.n0 VDD1.t3 17.6663
R90 VDD1.n2 VDD1.t5 17.6663
R91 VDD1.n2 VDD1.t4 17.6663
R92 VDD1.n1 VDD1.t7 17.6663
R93 VDD1.n1 VDD1.t6 17.6663
R94 VDD1 VDD1.n5 0.869035
R95 VTAIL.n66 VTAIL.n64 756.745
R96 VTAIL.n4 VTAIL.n2 756.745
R97 VTAIL.n12 VTAIL.n10 756.745
R98 VTAIL.n22 VTAIL.n20 756.745
R99 VTAIL.n58 VTAIL.n56 756.745
R100 VTAIL.n48 VTAIL.n46 756.745
R101 VTAIL.n40 VTAIL.n38 756.745
R102 VTAIL.n30 VTAIL.n28 756.745
R103 VTAIL.n67 VTAIL.n66 585
R104 VTAIL.n5 VTAIL.n4 585
R105 VTAIL.n13 VTAIL.n12 585
R106 VTAIL.n23 VTAIL.n22 585
R107 VTAIL.n59 VTAIL.n58 585
R108 VTAIL.n49 VTAIL.n48 585
R109 VTAIL.n41 VTAIL.n40 585
R110 VTAIL.n31 VTAIL.n30 585
R111 VTAIL.t7 VTAIL.n65 415.613
R112 VTAIL.t3 VTAIL.n3 415.613
R113 VTAIL.t9 VTAIL.n11 415.613
R114 VTAIL.t15 VTAIL.n21 415.613
R115 VTAIL.t11 VTAIL.n57 415.613
R116 VTAIL.t12 VTAIL.n47 415.613
R117 VTAIL.t1 VTAIL.n39 415.613
R118 VTAIL.t4 VTAIL.n29 415.613
R119 VTAIL.n55 VTAIL.n54 185.982
R120 VTAIL.n37 VTAIL.n36 185.982
R121 VTAIL.n1 VTAIL.n0 185.982
R122 VTAIL.n19 VTAIL.n18 185.982
R123 VTAIL.n66 VTAIL.t7 85.8723
R124 VTAIL.n4 VTAIL.t3 85.8723
R125 VTAIL.n12 VTAIL.t9 85.8723
R126 VTAIL.n22 VTAIL.t15 85.8723
R127 VTAIL.n58 VTAIL.t11 85.8723
R128 VTAIL.n48 VTAIL.t12 85.8723
R129 VTAIL.n40 VTAIL.t1 85.8723
R130 VTAIL.n30 VTAIL.t4 85.8723
R131 VTAIL.n71 VTAIL.n70 35.2884
R132 VTAIL.n9 VTAIL.n8 35.2884
R133 VTAIL.n17 VTAIL.n16 35.2884
R134 VTAIL.n27 VTAIL.n26 35.2884
R135 VTAIL.n63 VTAIL.n62 35.2884
R136 VTAIL.n53 VTAIL.n52 35.2884
R137 VTAIL.n45 VTAIL.n44 35.2884
R138 VTAIL.n35 VTAIL.n34 35.2884
R139 VTAIL.n0 VTAIL.t2 17.6663
R140 VTAIL.n0 VTAIL.t6 17.6663
R141 VTAIL.n18 VTAIL.t8 17.6663
R142 VTAIL.n18 VTAIL.t14 17.6663
R143 VTAIL.n54 VTAIL.t10 17.6663
R144 VTAIL.n54 VTAIL.t13 17.6663
R145 VTAIL.n36 VTAIL.t0 17.6663
R146 VTAIL.n36 VTAIL.t5 17.6663
R147 VTAIL.n71 VTAIL.n63 15.8065
R148 VTAIL.n35 VTAIL.n27 15.8065
R149 VTAIL.n67 VTAIL.n65 14.9339
R150 VTAIL.n5 VTAIL.n3 14.9339
R151 VTAIL.n13 VTAIL.n11 14.9339
R152 VTAIL.n23 VTAIL.n21 14.9339
R153 VTAIL.n59 VTAIL.n57 14.9339
R154 VTAIL.n49 VTAIL.n47 14.9339
R155 VTAIL.n41 VTAIL.n39 14.9339
R156 VTAIL.n31 VTAIL.n29 14.9339
R157 VTAIL.n68 VTAIL.n64 12.8005
R158 VTAIL.n6 VTAIL.n2 12.8005
R159 VTAIL.n14 VTAIL.n10 12.8005
R160 VTAIL.n24 VTAIL.n20 12.8005
R161 VTAIL.n60 VTAIL.n56 12.8005
R162 VTAIL.n50 VTAIL.n46 12.8005
R163 VTAIL.n42 VTAIL.n38 12.8005
R164 VTAIL.n32 VTAIL.n28 12.8005
R165 VTAIL.n70 VTAIL.n69 9.45567
R166 VTAIL.n8 VTAIL.n7 9.45567
R167 VTAIL.n16 VTAIL.n15 9.45567
R168 VTAIL.n26 VTAIL.n25 9.45567
R169 VTAIL.n62 VTAIL.n61 9.45567
R170 VTAIL.n52 VTAIL.n51 9.45567
R171 VTAIL.n44 VTAIL.n43 9.45567
R172 VTAIL.n34 VTAIL.n33 9.45567
R173 VTAIL.n69 VTAIL.n68 9.3005
R174 VTAIL.n7 VTAIL.n6 9.3005
R175 VTAIL.n15 VTAIL.n14 9.3005
R176 VTAIL.n25 VTAIL.n24 9.3005
R177 VTAIL.n61 VTAIL.n60 9.3005
R178 VTAIL.n51 VTAIL.n50 9.3005
R179 VTAIL.n43 VTAIL.n42 9.3005
R180 VTAIL.n33 VTAIL.n32 9.3005
R181 VTAIL.n69 VTAIL.n65 5.44463
R182 VTAIL.n7 VTAIL.n3 5.44463
R183 VTAIL.n15 VTAIL.n11 5.44463
R184 VTAIL.n25 VTAIL.n21 5.44463
R185 VTAIL.n61 VTAIL.n57 5.44463
R186 VTAIL.n51 VTAIL.n47 5.44463
R187 VTAIL.n43 VTAIL.n39 5.44463
R188 VTAIL.n33 VTAIL.n29 5.44463
R189 VTAIL.n37 VTAIL.n35 1.85395
R190 VTAIL.n45 VTAIL.n37 1.85395
R191 VTAIL.n55 VTAIL.n53 1.85395
R192 VTAIL.n63 VTAIL.n55 1.85395
R193 VTAIL.n27 VTAIL.n19 1.85395
R194 VTAIL.n19 VTAIL.n17 1.85395
R195 VTAIL.n9 VTAIL.n1 1.85395
R196 VTAIL VTAIL.n71 1.79576
R197 VTAIL.n70 VTAIL.n64 1.16414
R198 VTAIL.n8 VTAIL.n2 1.16414
R199 VTAIL.n16 VTAIL.n10 1.16414
R200 VTAIL.n26 VTAIL.n20 1.16414
R201 VTAIL.n62 VTAIL.n56 1.16414
R202 VTAIL.n52 VTAIL.n46 1.16414
R203 VTAIL.n44 VTAIL.n38 1.16414
R204 VTAIL.n34 VTAIL.n28 1.16414
R205 VTAIL.n53 VTAIL.n45 0.470328
R206 VTAIL.n17 VTAIL.n9 0.470328
R207 VTAIL.n68 VTAIL.n67 0.388379
R208 VTAIL.n6 VTAIL.n5 0.388379
R209 VTAIL.n14 VTAIL.n13 0.388379
R210 VTAIL.n24 VTAIL.n23 0.388379
R211 VTAIL.n60 VTAIL.n59 0.388379
R212 VTAIL.n50 VTAIL.n49 0.388379
R213 VTAIL.n42 VTAIL.n41 0.388379
R214 VTAIL.n32 VTAIL.n31 0.388379
R215 VTAIL VTAIL.n1 0.0586897
R216 B.n230 B.n229 585
R217 B.n228 B.n83 585
R218 B.n227 B.n226 585
R219 B.n225 B.n84 585
R220 B.n224 B.n223 585
R221 B.n222 B.n85 585
R222 B.n221 B.n220 585
R223 B.n219 B.n86 585
R224 B.n218 B.n217 585
R225 B.n216 B.n87 585
R226 B.n215 B.n214 585
R227 B.n213 B.n88 585
R228 B.n212 B.n211 585
R229 B.n207 B.n89 585
R230 B.n206 B.n205 585
R231 B.n204 B.n90 585
R232 B.n203 B.n202 585
R233 B.n201 B.n91 585
R234 B.n200 B.n199 585
R235 B.n198 B.n92 585
R236 B.n197 B.n196 585
R237 B.n194 B.n93 585
R238 B.n193 B.n192 585
R239 B.n191 B.n96 585
R240 B.n190 B.n189 585
R241 B.n188 B.n97 585
R242 B.n187 B.n186 585
R243 B.n185 B.n98 585
R244 B.n184 B.n183 585
R245 B.n182 B.n99 585
R246 B.n181 B.n180 585
R247 B.n179 B.n100 585
R248 B.n178 B.n177 585
R249 B.n231 B.n82 585
R250 B.n233 B.n232 585
R251 B.n234 B.n81 585
R252 B.n236 B.n235 585
R253 B.n237 B.n80 585
R254 B.n239 B.n238 585
R255 B.n240 B.n79 585
R256 B.n242 B.n241 585
R257 B.n243 B.n78 585
R258 B.n245 B.n244 585
R259 B.n246 B.n77 585
R260 B.n248 B.n247 585
R261 B.n249 B.n76 585
R262 B.n251 B.n250 585
R263 B.n252 B.n75 585
R264 B.n254 B.n253 585
R265 B.n255 B.n74 585
R266 B.n257 B.n256 585
R267 B.n258 B.n73 585
R268 B.n260 B.n259 585
R269 B.n261 B.n72 585
R270 B.n263 B.n262 585
R271 B.n264 B.n71 585
R272 B.n266 B.n265 585
R273 B.n267 B.n70 585
R274 B.n269 B.n268 585
R275 B.n270 B.n69 585
R276 B.n272 B.n271 585
R277 B.n273 B.n68 585
R278 B.n275 B.n274 585
R279 B.n276 B.n67 585
R280 B.n278 B.n277 585
R281 B.n279 B.n66 585
R282 B.n281 B.n280 585
R283 B.n282 B.n65 585
R284 B.n284 B.n283 585
R285 B.n285 B.n64 585
R286 B.n287 B.n286 585
R287 B.n288 B.n63 585
R288 B.n290 B.n289 585
R289 B.n291 B.n62 585
R290 B.n293 B.n292 585
R291 B.n294 B.n61 585
R292 B.n296 B.n295 585
R293 B.n297 B.n60 585
R294 B.n299 B.n298 585
R295 B.n300 B.n59 585
R296 B.n302 B.n301 585
R297 B.n303 B.n58 585
R298 B.n305 B.n304 585
R299 B.n306 B.n57 585
R300 B.n308 B.n307 585
R301 B.n309 B.n56 585
R302 B.n311 B.n310 585
R303 B.n312 B.n55 585
R304 B.n314 B.n313 585
R305 B.n315 B.n54 585
R306 B.n317 B.n316 585
R307 B.n318 B.n53 585
R308 B.n320 B.n319 585
R309 B.n321 B.n52 585
R310 B.n323 B.n322 585
R311 B.n324 B.n51 585
R312 B.n326 B.n325 585
R313 B.n327 B.n50 585
R314 B.n329 B.n328 585
R315 B.n330 B.n49 585
R316 B.n332 B.n331 585
R317 B.n333 B.n48 585
R318 B.n335 B.n334 585
R319 B.n336 B.n47 585
R320 B.n338 B.n337 585
R321 B.n339 B.n46 585
R322 B.n341 B.n340 585
R323 B.n342 B.n45 585
R324 B.n344 B.n343 585
R325 B.n345 B.n44 585
R326 B.n347 B.n346 585
R327 B.n348 B.n43 585
R328 B.n350 B.n349 585
R329 B.n401 B.n400 585
R330 B.n399 B.n22 585
R331 B.n398 B.n397 585
R332 B.n396 B.n23 585
R333 B.n395 B.n394 585
R334 B.n393 B.n24 585
R335 B.n392 B.n391 585
R336 B.n390 B.n25 585
R337 B.n389 B.n388 585
R338 B.n387 B.n26 585
R339 B.n386 B.n385 585
R340 B.n384 B.n27 585
R341 B.n382 B.n381 585
R342 B.n380 B.n30 585
R343 B.n379 B.n378 585
R344 B.n377 B.n31 585
R345 B.n376 B.n375 585
R346 B.n374 B.n32 585
R347 B.n373 B.n372 585
R348 B.n371 B.n33 585
R349 B.n370 B.n369 585
R350 B.n368 B.n367 585
R351 B.n366 B.n37 585
R352 B.n365 B.n364 585
R353 B.n363 B.n38 585
R354 B.n362 B.n361 585
R355 B.n360 B.n39 585
R356 B.n359 B.n358 585
R357 B.n357 B.n40 585
R358 B.n356 B.n355 585
R359 B.n354 B.n41 585
R360 B.n353 B.n352 585
R361 B.n351 B.n42 585
R362 B.n402 B.n21 585
R363 B.n404 B.n403 585
R364 B.n405 B.n20 585
R365 B.n407 B.n406 585
R366 B.n408 B.n19 585
R367 B.n410 B.n409 585
R368 B.n411 B.n18 585
R369 B.n413 B.n412 585
R370 B.n414 B.n17 585
R371 B.n416 B.n415 585
R372 B.n417 B.n16 585
R373 B.n419 B.n418 585
R374 B.n420 B.n15 585
R375 B.n422 B.n421 585
R376 B.n423 B.n14 585
R377 B.n425 B.n424 585
R378 B.n426 B.n13 585
R379 B.n428 B.n427 585
R380 B.n429 B.n12 585
R381 B.n431 B.n430 585
R382 B.n432 B.n11 585
R383 B.n434 B.n433 585
R384 B.n435 B.n10 585
R385 B.n437 B.n436 585
R386 B.n438 B.n9 585
R387 B.n440 B.n439 585
R388 B.n441 B.n8 585
R389 B.n443 B.n442 585
R390 B.n444 B.n7 585
R391 B.n446 B.n445 585
R392 B.n447 B.n6 585
R393 B.n449 B.n448 585
R394 B.n450 B.n5 585
R395 B.n452 B.n451 585
R396 B.n453 B.n4 585
R397 B.n455 B.n454 585
R398 B.n456 B.n3 585
R399 B.n458 B.n457 585
R400 B.n459 B.n0 585
R401 B.n2 B.n1 585
R402 B.n121 B.n120 585
R403 B.n122 B.n119 585
R404 B.n124 B.n123 585
R405 B.n125 B.n118 585
R406 B.n127 B.n126 585
R407 B.n128 B.n117 585
R408 B.n130 B.n129 585
R409 B.n131 B.n116 585
R410 B.n133 B.n132 585
R411 B.n134 B.n115 585
R412 B.n136 B.n135 585
R413 B.n137 B.n114 585
R414 B.n139 B.n138 585
R415 B.n140 B.n113 585
R416 B.n142 B.n141 585
R417 B.n143 B.n112 585
R418 B.n145 B.n144 585
R419 B.n146 B.n111 585
R420 B.n148 B.n147 585
R421 B.n149 B.n110 585
R422 B.n151 B.n150 585
R423 B.n152 B.n109 585
R424 B.n154 B.n153 585
R425 B.n155 B.n108 585
R426 B.n157 B.n156 585
R427 B.n158 B.n107 585
R428 B.n160 B.n159 585
R429 B.n161 B.n106 585
R430 B.n163 B.n162 585
R431 B.n164 B.n105 585
R432 B.n166 B.n165 585
R433 B.n167 B.n104 585
R434 B.n169 B.n168 585
R435 B.n170 B.n103 585
R436 B.n172 B.n171 585
R437 B.n173 B.n102 585
R438 B.n175 B.n174 585
R439 B.n176 B.n101 585
R440 B.n178 B.n101 540.549
R441 B.n231 B.n230 540.549
R442 B.n351 B.n350 540.549
R443 B.n400 B.n21 540.549
R444 B.n208 B.t7 286.932
R445 B.n34 B.t2 286.932
R446 B.n94 B.t4 286.932
R447 B.n28 B.t11 286.932
R448 B.n461 B.n460 256.663
R449 B.n209 B.t8 245.234
R450 B.n35 B.t1 245.234
R451 B.n95 B.t5 245.234
R452 B.n29 B.t10 245.234
R453 B.n460 B.n459 235.042
R454 B.n460 B.n2 235.042
R455 B.n94 B.t3 230.827
R456 B.n208 B.t6 230.827
R457 B.n34 B.t0 230.827
R458 B.n28 B.t9 230.827
R459 B.n179 B.n178 163.367
R460 B.n180 B.n179 163.367
R461 B.n180 B.n99 163.367
R462 B.n184 B.n99 163.367
R463 B.n185 B.n184 163.367
R464 B.n186 B.n185 163.367
R465 B.n186 B.n97 163.367
R466 B.n190 B.n97 163.367
R467 B.n191 B.n190 163.367
R468 B.n192 B.n191 163.367
R469 B.n192 B.n93 163.367
R470 B.n197 B.n93 163.367
R471 B.n198 B.n197 163.367
R472 B.n199 B.n198 163.367
R473 B.n199 B.n91 163.367
R474 B.n203 B.n91 163.367
R475 B.n204 B.n203 163.367
R476 B.n205 B.n204 163.367
R477 B.n205 B.n89 163.367
R478 B.n212 B.n89 163.367
R479 B.n213 B.n212 163.367
R480 B.n214 B.n213 163.367
R481 B.n214 B.n87 163.367
R482 B.n218 B.n87 163.367
R483 B.n219 B.n218 163.367
R484 B.n220 B.n219 163.367
R485 B.n220 B.n85 163.367
R486 B.n224 B.n85 163.367
R487 B.n225 B.n224 163.367
R488 B.n226 B.n225 163.367
R489 B.n226 B.n83 163.367
R490 B.n230 B.n83 163.367
R491 B.n350 B.n43 163.367
R492 B.n346 B.n43 163.367
R493 B.n346 B.n345 163.367
R494 B.n345 B.n344 163.367
R495 B.n344 B.n45 163.367
R496 B.n340 B.n45 163.367
R497 B.n340 B.n339 163.367
R498 B.n339 B.n338 163.367
R499 B.n338 B.n47 163.367
R500 B.n334 B.n47 163.367
R501 B.n334 B.n333 163.367
R502 B.n333 B.n332 163.367
R503 B.n332 B.n49 163.367
R504 B.n328 B.n49 163.367
R505 B.n328 B.n327 163.367
R506 B.n327 B.n326 163.367
R507 B.n326 B.n51 163.367
R508 B.n322 B.n51 163.367
R509 B.n322 B.n321 163.367
R510 B.n321 B.n320 163.367
R511 B.n320 B.n53 163.367
R512 B.n316 B.n53 163.367
R513 B.n316 B.n315 163.367
R514 B.n315 B.n314 163.367
R515 B.n314 B.n55 163.367
R516 B.n310 B.n55 163.367
R517 B.n310 B.n309 163.367
R518 B.n309 B.n308 163.367
R519 B.n308 B.n57 163.367
R520 B.n304 B.n57 163.367
R521 B.n304 B.n303 163.367
R522 B.n303 B.n302 163.367
R523 B.n302 B.n59 163.367
R524 B.n298 B.n59 163.367
R525 B.n298 B.n297 163.367
R526 B.n297 B.n296 163.367
R527 B.n296 B.n61 163.367
R528 B.n292 B.n61 163.367
R529 B.n292 B.n291 163.367
R530 B.n291 B.n290 163.367
R531 B.n290 B.n63 163.367
R532 B.n286 B.n63 163.367
R533 B.n286 B.n285 163.367
R534 B.n285 B.n284 163.367
R535 B.n284 B.n65 163.367
R536 B.n280 B.n65 163.367
R537 B.n280 B.n279 163.367
R538 B.n279 B.n278 163.367
R539 B.n278 B.n67 163.367
R540 B.n274 B.n67 163.367
R541 B.n274 B.n273 163.367
R542 B.n273 B.n272 163.367
R543 B.n272 B.n69 163.367
R544 B.n268 B.n69 163.367
R545 B.n268 B.n267 163.367
R546 B.n267 B.n266 163.367
R547 B.n266 B.n71 163.367
R548 B.n262 B.n71 163.367
R549 B.n262 B.n261 163.367
R550 B.n261 B.n260 163.367
R551 B.n260 B.n73 163.367
R552 B.n256 B.n73 163.367
R553 B.n256 B.n255 163.367
R554 B.n255 B.n254 163.367
R555 B.n254 B.n75 163.367
R556 B.n250 B.n75 163.367
R557 B.n250 B.n249 163.367
R558 B.n249 B.n248 163.367
R559 B.n248 B.n77 163.367
R560 B.n244 B.n77 163.367
R561 B.n244 B.n243 163.367
R562 B.n243 B.n242 163.367
R563 B.n242 B.n79 163.367
R564 B.n238 B.n79 163.367
R565 B.n238 B.n237 163.367
R566 B.n237 B.n236 163.367
R567 B.n236 B.n81 163.367
R568 B.n232 B.n81 163.367
R569 B.n232 B.n231 163.367
R570 B.n400 B.n399 163.367
R571 B.n399 B.n398 163.367
R572 B.n398 B.n23 163.367
R573 B.n394 B.n23 163.367
R574 B.n394 B.n393 163.367
R575 B.n393 B.n392 163.367
R576 B.n392 B.n25 163.367
R577 B.n388 B.n25 163.367
R578 B.n388 B.n387 163.367
R579 B.n387 B.n386 163.367
R580 B.n386 B.n27 163.367
R581 B.n381 B.n27 163.367
R582 B.n381 B.n380 163.367
R583 B.n380 B.n379 163.367
R584 B.n379 B.n31 163.367
R585 B.n375 B.n31 163.367
R586 B.n375 B.n374 163.367
R587 B.n374 B.n373 163.367
R588 B.n373 B.n33 163.367
R589 B.n369 B.n33 163.367
R590 B.n369 B.n368 163.367
R591 B.n368 B.n37 163.367
R592 B.n364 B.n37 163.367
R593 B.n364 B.n363 163.367
R594 B.n363 B.n362 163.367
R595 B.n362 B.n39 163.367
R596 B.n358 B.n39 163.367
R597 B.n358 B.n357 163.367
R598 B.n357 B.n356 163.367
R599 B.n356 B.n41 163.367
R600 B.n352 B.n41 163.367
R601 B.n352 B.n351 163.367
R602 B.n404 B.n21 163.367
R603 B.n405 B.n404 163.367
R604 B.n406 B.n405 163.367
R605 B.n406 B.n19 163.367
R606 B.n410 B.n19 163.367
R607 B.n411 B.n410 163.367
R608 B.n412 B.n411 163.367
R609 B.n412 B.n17 163.367
R610 B.n416 B.n17 163.367
R611 B.n417 B.n416 163.367
R612 B.n418 B.n417 163.367
R613 B.n418 B.n15 163.367
R614 B.n422 B.n15 163.367
R615 B.n423 B.n422 163.367
R616 B.n424 B.n423 163.367
R617 B.n424 B.n13 163.367
R618 B.n428 B.n13 163.367
R619 B.n429 B.n428 163.367
R620 B.n430 B.n429 163.367
R621 B.n430 B.n11 163.367
R622 B.n434 B.n11 163.367
R623 B.n435 B.n434 163.367
R624 B.n436 B.n435 163.367
R625 B.n436 B.n9 163.367
R626 B.n440 B.n9 163.367
R627 B.n441 B.n440 163.367
R628 B.n442 B.n441 163.367
R629 B.n442 B.n7 163.367
R630 B.n446 B.n7 163.367
R631 B.n447 B.n446 163.367
R632 B.n448 B.n447 163.367
R633 B.n448 B.n5 163.367
R634 B.n452 B.n5 163.367
R635 B.n453 B.n452 163.367
R636 B.n454 B.n453 163.367
R637 B.n454 B.n3 163.367
R638 B.n458 B.n3 163.367
R639 B.n459 B.n458 163.367
R640 B.n120 B.n2 163.367
R641 B.n120 B.n119 163.367
R642 B.n124 B.n119 163.367
R643 B.n125 B.n124 163.367
R644 B.n126 B.n125 163.367
R645 B.n126 B.n117 163.367
R646 B.n130 B.n117 163.367
R647 B.n131 B.n130 163.367
R648 B.n132 B.n131 163.367
R649 B.n132 B.n115 163.367
R650 B.n136 B.n115 163.367
R651 B.n137 B.n136 163.367
R652 B.n138 B.n137 163.367
R653 B.n138 B.n113 163.367
R654 B.n142 B.n113 163.367
R655 B.n143 B.n142 163.367
R656 B.n144 B.n143 163.367
R657 B.n144 B.n111 163.367
R658 B.n148 B.n111 163.367
R659 B.n149 B.n148 163.367
R660 B.n150 B.n149 163.367
R661 B.n150 B.n109 163.367
R662 B.n154 B.n109 163.367
R663 B.n155 B.n154 163.367
R664 B.n156 B.n155 163.367
R665 B.n156 B.n107 163.367
R666 B.n160 B.n107 163.367
R667 B.n161 B.n160 163.367
R668 B.n162 B.n161 163.367
R669 B.n162 B.n105 163.367
R670 B.n166 B.n105 163.367
R671 B.n167 B.n166 163.367
R672 B.n168 B.n167 163.367
R673 B.n168 B.n103 163.367
R674 B.n172 B.n103 163.367
R675 B.n173 B.n172 163.367
R676 B.n174 B.n173 163.367
R677 B.n174 B.n101 163.367
R678 B.n195 B.n95 59.5399
R679 B.n210 B.n209 59.5399
R680 B.n36 B.n35 59.5399
R681 B.n383 B.n29 59.5399
R682 B.n95 B.n94 41.6975
R683 B.n209 B.n208 41.6975
R684 B.n35 B.n34 41.6975
R685 B.n29 B.n28 41.6975
R686 B.n402 B.n401 35.1225
R687 B.n349 B.n42 35.1225
R688 B.n229 B.n82 35.1225
R689 B.n177 B.n176 35.1225
R690 B B.n461 18.0485
R691 B.n403 B.n402 10.6151
R692 B.n403 B.n20 10.6151
R693 B.n407 B.n20 10.6151
R694 B.n408 B.n407 10.6151
R695 B.n409 B.n408 10.6151
R696 B.n409 B.n18 10.6151
R697 B.n413 B.n18 10.6151
R698 B.n414 B.n413 10.6151
R699 B.n415 B.n414 10.6151
R700 B.n415 B.n16 10.6151
R701 B.n419 B.n16 10.6151
R702 B.n420 B.n419 10.6151
R703 B.n421 B.n420 10.6151
R704 B.n421 B.n14 10.6151
R705 B.n425 B.n14 10.6151
R706 B.n426 B.n425 10.6151
R707 B.n427 B.n426 10.6151
R708 B.n427 B.n12 10.6151
R709 B.n431 B.n12 10.6151
R710 B.n432 B.n431 10.6151
R711 B.n433 B.n432 10.6151
R712 B.n433 B.n10 10.6151
R713 B.n437 B.n10 10.6151
R714 B.n438 B.n437 10.6151
R715 B.n439 B.n438 10.6151
R716 B.n439 B.n8 10.6151
R717 B.n443 B.n8 10.6151
R718 B.n444 B.n443 10.6151
R719 B.n445 B.n444 10.6151
R720 B.n445 B.n6 10.6151
R721 B.n449 B.n6 10.6151
R722 B.n450 B.n449 10.6151
R723 B.n451 B.n450 10.6151
R724 B.n451 B.n4 10.6151
R725 B.n455 B.n4 10.6151
R726 B.n456 B.n455 10.6151
R727 B.n457 B.n456 10.6151
R728 B.n457 B.n0 10.6151
R729 B.n401 B.n22 10.6151
R730 B.n397 B.n22 10.6151
R731 B.n397 B.n396 10.6151
R732 B.n396 B.n395 10.6151
R733 B.n395 B.n24 10.6151
R734 B.n391 B.n24 10.6151
R735 B.n391 B.n390 10.6151
R736 B.n390 B.n389 10.6151
R737 B.n389 B.n26 10.6151
R738 B.n385 B.n26 10.6151
R739 B.n385 B.n384 10.6151
R740 B.n382 B.n30 10.6151
R741 B.n378 B.n30 10.6151
R742 B.n378 B.n377 10.6151
R743 B.n377 B.n376 10.6151
R744 B.n376 B.n32 10.6151
R745 B.n372 B.n32 10.6151
R746 B.n372 B.n371 10.6151
R747 B.n371 B.n370 10.6151
R748 B.n367 B.n366 10.6151
R749 B.n366 B.n365 10.6151
R750 B.n365 B.n38 10.6151
R751 B.n361 B.n38 10.6151
R752 B.n361 B.n360 10.6151
R753 B.n360 B.n359 10.6151
R754 B.n359 B.n40 10.6151
R755 B.n355 B.n40 10.6151
R756 B.n355 B.n354 10.6151
R757 B.n354 B.n353 10.6151
R758 B.n353 B.n42 10.6151
R759 B.n349 B.n348 10.6151
R760 B.n348 B.n347 10.6151
R761 B.n347 B.n44 10.6151
R762 B.n343 B.n44 10.6151
R763 B.n343 B.n342 10.6151
R764 B.n342 B.n341 10.6151
R765 B.n341 B.n46 10.6151
R766 B.n337 B.n46 10.6151
R767 B.n337 B.n336 10.6151
R768 B.n336 B.n335 10.6151
R769 B.n335 B.n48 10.6151
R770 B.n331 B.n48 10.6151
R771 B.n331 B.n330 10.6151
R772 B.n330 B.n329 10.6151
R773 B.n329 B.n50 10.6151
R774 B.n325 B.n50 10.6151
R775 B.n325 B.n324 10.6151
R776 B.n324 B.n323 10.6151
R777 B.n323 B.n52 10.6151
R778 B.n319 B.n52 10.6151
R779 B.n319 B.n318 10.6151
R780 B.n318 B.n317 10.6151
R781 B.n317 B.n54 10.6151
R782 B.n313 B.n54 10.6151
R783 B.n313 B.n312 10.6151
R784 B.n312 B.n311 10.6151
R785 B.n311 B.n56 10.6151
R786 B.n307 B.n56 10.6151
R787 B.n307 B.n306 10.6151
R788 B.n306 B.n305 10.6151
R789 B.n305 B.n58 10.6151
R790 B.n301 B.n58 10.6151
R791 B.n301 B.n300 10.6151
R792 B.n300 B.n299 10.6151
R793 B.n299 B.n60 10.6151
R794 B.n295 B.n60 10.6151
R795 B.n295 B.n294 10.6151
R796 B.n294 B.n293 10.6151
R797 B.n293 B.n62 10.6151
R798 B.n289 B.n62 10.6151
R799 B.n289 B.n288 10.6151
R800 B.n288 B.n287 10.6151
R801 B.n287 B.n64 10.6151
R802 B.n283 B.n64 10.6151
R803 B.n283 B.n282 10.6151
R804 B.n282 B.n281 10.6151
R805 B.n281 B.n66 10.6151
R806 B.n277 B.n66 10.6151
R807 B.n277 B.n276 10.6151
R808 B.n276 B.n275 10.6151
R809 B.n275 B.n68 10.6151
R810 B.n271 B.n68 10.6151
R811 B.n271 B.n270 10.6151
R812 B.n270 B.n269 10.6151
R813 B.n269 B.n70 10.6151
R814 B.n265 B.n70 10.6151
R815 B.n265 B.n264 10.6151
R816 B.n264 B.n263 10.6151
R817 B.n263 B.n72 10.6151
R818 B.n259 B.n72 10.6151
R819 B.n259 B.n258 10.6151
R820 B.n258 B.n257 10.6151
R821 B.n257 B.n74 10.6151
R822 B.n253 B.n74 10.6151
R823 B.n253 B.n252 10.6151
R824 B.n252 B.n251 10.6151
R825 B.n251 B.n76 10.6151
R826 B.n247 B.n76 10.6151
R827 B.n247 B.n246 10.6151
R828 B.n246 B.n245 10.6151
R829 B.n245 B.n78 10.6151
R830 B.n241 B.n78 10.6151
R831 B.n241 B.n240 10.6151
R832 B.n240 B.n239 10.6151
R833 B.n239 B.n80 10.6151
R834 B.n235 B.n80 10.6151
R835 B.n235 B.n234 10.6151
R836 B.n234 B.n233 10.6151
R837 B.n233 B.n82 10.6151
R838 B.n121 B.n1 10.6151
R839 B.n122 B.n121 10.6151
R840 B.n123 B.n122 10.6151
R841 B.n123 B.n118 10.6151
R842 B.n127 B.n118 10.6151
R843 B.n128 B.n127 10.6151
R844 B.n129 B.n128 10.6151
R845 B.n129 B.n116 10.6151
R846 B.n133 B.n116 10.6151
R847 B.n134 B.n133 10.6151
R848 B.n135 B.n134 10.6151
R849 B.n135 B.n114 10.6151
R850 B.n139 B.n114 10.6151
R851 B.n140 B.n139 10.6151
R852 B.n141 B.n140 10.6151
R853 B.n141 B.n112 10.6151
R854 B.n145 B.n112 10.6151
R855 B.n146 B.n145 10.6151
R856 B.n147 B.n146 10.6151
R857 B.n147 B.n110 10.6151
R858 B.n151 B.n110 10.6151
R859 B.n152 B.n151 10.6151
R860 B.n153 B.n152 10.6151
R861 B.n153 B.n108 10.6151
R862 B.n157 B.n108 10.6151
R863 B.n158 B.n157 10.6151
R864 B.n159 B.n158 10.6151
R865 B.n159 B.n106 10.6151
R866 B.n163 B.n106 10.6151
R867 B.n164 B.n163 10.6151
R868 B.n165 B.n164 10.6151
R869 B.n165 B.n104 10.6151
R870 B.n169 B.n104 10.6151
R871 B.n170 B.n169 10.6151
R872 B.n171 B.n170 10.6151
R873 B.n171 B.n102 10.6151
R874 B.n175 B.n102 10.6151
R875 B.n176 B.n175 10.6151
R876 B.n177 B.n100 10.6151
R877 B.n181 B.n100 10.6151
R878 B.n182 B.n181 10.6151
R879 B.n183 B.n182 10.6151
R880 B.n183 B.n98 10.6151
R881 B.n187 B.n98 10.6151
R882 B.n188 B.n187 10.6151
R883 B.n189 B.n188 10.6151
R884 B.n189 B.n96 10.6151
R885 B.n193 B.n96 10.6151
R886 B.n194 B.n193 10.6151
R887 B.n196 B.n92 10.6151
R888 B.n200 B.n92 10.6151
R889 B.n201 B.n200 10.6151
R890 B.n202 B.n201 10.6151
R891 B.n202 B.n90 10.6151
R892 B.n206 B.n90 10.6151
R893 B.n207 B.n206 10.6151
R894 B.n211 B.n207 10.6151
R895 B.n215 B.n88 10.6151
R896 B.n216 B.n215 10.6151
R897 B.n217 B.n216 10.6151
R898 B.n217 B.n86 10.6151
R899 B.n221 B.n86 10.6151
R900 B.n222 B.n221 10.6151
R901 B.n223 B.n222 10.6151
R902 B.n223 B.n84 10.6151
R903 B.n227 B.n84 10.6151
R904 B.n228 B.n227 10.6151
R905 B.n229 B.n228 10.6151
R906 B.n461 B.n0 8.11757
R907 B.n461 B.n1 8.11757
R908 B.n383 B.n382 6.5566
R909 B.n370 B.n36 6.5566
R910 B.n196 B.n195 6.5566
R911 B.n211 B.n210 6.5566
R912 B.n384 B.n383 4.05904
R913 B.n367 B.n36 4.05904
R914 B.n195 B.n194 4.05904
R915 B.n210 B.n88 4.05904
R916 VN.n39 VN.n21 161.3
R917 VN.n38 VN.n37 161.3
R918 VN.n36 VN.n22 161.3
R919 VN.n35 VN.n34 161.3
R920 VN.n32 VN.n23 161.3
R921 VN.n31 VN.n30 161.3
R922 VN.n29 VN.n24 161.3
R923 VN.n28 VN.n27 161.3
R924 VN.n18 VN.n0 161.3
R925 VN.n17 VN.n16 161.3
R926 VN.n15 VN.n1 161.3
R927 VN.n14 VN.n13 161.3
R928 VN.n11 VN.n2 161.3
R929 VN.n10 VN.n9 161.3
R930 VN.n8 VN.n3 161.3
R931 VN.n7 VN.n6 161.3
R932 VN.n20 VN.n19 87.546
R933 VN.n41 VN.n40 87.546
R934 VN.n10 VN.n3 56.5617
R935 VN.n31 VN.n24 56.5617
R936 VN.n4 VN.t0 55.8733
R937 VN.n25 VN.t1 55.8733
R938 VN.n5 VN.n4 54.0319
R939 VN.n26 VN.n25 54.0319
R940 VN.n17 VN.n1 50.2647
R941 VN.n38 VN.n22 50.2647
R942 VN VN.n41 39.8618
R943 VN.n18 VN.n17 30.8893
R944 VN.n39 VN.n38 30.8893
R945 VN.n6 VN.n3 24.5923
R946 VN.n11 VN.n10 24.5923
R947 VN.n13 VN.n1 24.5923
R948 VN.n27 VN.n24 24.5923
R949 VN.n34 VN.n22 24.5923
R950 VN.n32 VN.n31 24.5923
R951 VN.n5 VN.t2 24.3653
R952 VN.n12 VN.t4 24.3653
R953 VN.n19 VN.t5 24.3653
R954 VN.n26 VN.t3 24.3653
R955 VN.n33 VN.t6 24.3653
R956 VN.n40 VN.t7 24.3653
R957 VN.n19 VN.n18 23.3627
R958 VN.n40 VN.n39 23.3627
R959 VN.n6 VN.n5 15.9852
R960 VN.n12 VN.n11 15.9852
R961 VN.n27 VN.n26 15.9852
R962 VN.n33 VN.n32 15.9852
R963 VN.n28 VN.n25 12.7521
R964 VN.n7 VN.n4 12.7521
R965 VN.n13 VN.n12 8.60764
R966 VN.n34 VN.n33 8.60764
R967 VN.n41 VN.n21 0.278335
R968 VN.n20 VN.n0 0.278335
R969 VN.n37 VN.n21 0.189894
R970 VN.n37 VN.n36 0.189894
R971 VN.n36 VN.n35 0.189894
R972 VN.n35 VN.n23 0.189894
R973 VN.n30 VN.n23 0.189894
R974 VN.n30 VN.n29 0.189894
R975 VN.n29 VN.n28 0.189894
R976 VN.n8 VN.n7 0.189894
R977 VN.n9 VN.n8 0.189894
R978 VN.n9 VN.n2 0.189894
R979 VN.n14 VN.n2 0.189894
R980 VN.n15 VN.n14 0.189894
R981 VN.n16 VN.n15 0.189894
R982 VN.n16 VN.n0 0.189894
R983 VN VN.n20 0.153485
R984 VDD2.n2 VDD2.n1 203.534
R985 VDD2.n2 VDD2.n0 203.534
R986 VDD2 VDD2.n5 203.53
R987 VDD2.n4 VDD2.n3 202.661
R988 VDD2.n4 VDD2.n2 33.642
R989 VDD2.n5 VDD2.t4 17.6663
R990 VDD2.n5 VDD2.t6 17.6663
R991 VDD2.n3 VDD2.t0 17.6663
R992 VDD2.n3 VDD2.t1 17.6663
R993 VDD2.n1 VDD2.t3 17.6663
R994 VDD2.n1 VDD2.t2 17.6663
R995 VDD2.n0 VDD2.t7 17.6663
R996 VDD2.n0 VDD2.t5 17.6663
R997 VDD2 VDD2.n4 0.985414
C0 VDD1 w_n3120_n1336# 1.41905f
C1 VN VDD1 0.156486f
C2 VDD1 B 1.13738f
C3 VP w_n3120_n1336# 6.33309f
C4 VN VP 4.83243f
C5 VDD2 VDD1 1.3704f
C6 VN w_n3120_n1336# 5.93549f
C7 B VP 1.5914f
C8 B w_n3120_n1336# 6.09719f
C9 VN B 0.921238f
C10 VTAIL VDD1 3.99863f
C11 VDD2 VP 0.443932f
C12 VDD2 w_n3120_n1336# 1.50027f
C13 VDD2 VN 1.59774f
C14 VTAIL VP 2.39892f
C15 VDD2 B 1.20916f
C16 VTAIL w_n3120_n1336# 1.76021f
C17 VTAIL VN 2.38481f
C18 VTAIL B 1.35684f
C19 VDD1 VP 1.88288f
C20 VDD2 VTAIL 4.04782f
C21 VDD2 VSUBS 0.954869f
C22 VDD1 VSUBS 1.44742f
C23 VTAIL VSUBS 0.44555f
C24 VN VSUBS 5.44241f
C25 VP VSUBS 2.226272f
C26 B VSUBS 3.081581f
C27 w_n3120_n1336# VSUBS 53.277103f
C28 VDD2.t7 VSUBS 0.02509f
C29 VDD2.t5 VSUBS 0.02509f
C30 VDD2.n0 VSUBS 0.10773f
C31 VDD2.t3 VSUBS 0.02509f
C32 VDD2.t2 VSUBS 0.02509f
C33 VDD2.n1 VSUBS 0.10773f
C34 VDD2.n2 VSUBS 1.60254f
C35 VDD2.t0 VSUBS 0.02509f
C36 VDD2.t1 VSUBS 0.02509f
C37 VDD2.n3 VSUBS 0.106295f
C38 VDD2.n4 VSUBS 1.33098f
C39 VDD2.t4 VSUBS 0.02509f
C40 VDD2.t6 VSUBS 0.02509f
C41 VDD2.n5 VSUBS 0.107723f
C42 VN.n0 VSUBS 0.069182f
C43 VN.t5 VSUBS 0.403276f
C44 VN.n1 VSUBS 0.095842f
C45 VN.n2 VSUBS 0.052477f
C46 VN.t4 VSUBS 0.403276f
C47 VN.n3 VSUBS 0.076284f
C48 VN.t0 VSUBS 0.660769f
C49 VN.n4 VSUBS 0.310759f
C50 VN.t2 VSUBS 0.403276f
C51 VN.n5 VSUBS 0.336307f
C52 VN.n6 VSUBS 0.0805f
C53 VN.n7 VSUBS 0.384435f
C54 VN.n8 VSUBS 0.052477f
C55 VN.n9 VSUBS 0.052477f
C56 VN.n10 VSUBS 0.076284f
C57 VN.n11 VSUBS 0.0805f
C58 VN.n12 VSUBS 0.212207f
C59 VN.n13 VSUBS 0.066087f
C60 VN.n14 VSUBS 0.052477f
C61 VN.n15 VSUBS 0.052477f
C62 VN.n16 VSUBS 0.052477f
C63 VN.n17 VSUBS 0.049479f
C64 VN.n18 VSUBS 0.10216f
C65 VN.n19 VSUBS 0.368606f
C66 VN.n20 VSUBS 0.057044f
C67 VN.n21 VSUBS 0.069182f
C68 VN.t7 VSUBS 0.403276f
C69 VN.n22 VSUBS 0.095842f
C70 VN.n23 VSUBS 0.052477f
C71 VN.t6 VSUBS 0.403276f
C72 VN.n24 VSUBS 0.076284f
C73 VN.t1 VSUBS 0.660769f
C74 VN.n25 VSUBS 0.310759f
C75 VN.t3 VSUBS 0.403276f
C76 VN.n26 VSUBS 0.336307f
C77 VN.n27 VSUBS 0.0805f
C78 VN.n28 VSUBS 0.384435f
C79 VN.n29 VSUBS 0.052477f
C80 VN.n30 VSUBS 0.052477f
C81 VN.n31 VSUBS 0.076284f
C82 VN.n32 VSUBS 0.0805f
C83 VN.n33 VSUBS 0.212207f
C84 VN.n34 VSUBS 0.066087f
C85 VN.n35 VSUBS 0.052477f
C86 VN.n36 VSUBS 0.052477f
C87 VN.n37 VSUBS 0.052477f
C88 VN.n38 VSUBS 0.049479f
C89 VN.n39 VSUBS 0.10216f
C90 VN.n40 VSUBS 0.368606f
C91 VN.n41 VSUBS 2.0245f
C92 B.n0 VSUBS 0.007761f
C93 B.n1 VSUBS 0.007761f
C94 B.n2 VSUBS 0.011478f
C95 B.n3 VSUBS 0.008796f
C96 B.n4 VSUBS 0.008796f
C97 B.n5 VSUBS 0.008796f
C98 B.n6 VSUBS 0.008796f
C99 B.n7 VSUBS 0.008796f
C100 B.n8 VSUBS 0.008796f
C101 B.n9 VSUBS 0.008796f
C102 B.n10 VSUBS 0.008796f
C103 B.n11 VSUBS 0.008796f
C104 B.n12 VSUBS 0.008796f
C105 B.n13 VSUBS 0.008796f
C106 B.n14 VSUBS 0.008796f
C107 B.n15 VSUBS 0.008796f
C108 B.n16 VSUBS 0.008796f
C109 B.n17 VSUBS 0.008796f
C110 B.n18 VSUBS 0.008796f
C111 B.n19 VSUBS 0.008796f
C112 B.n20 VSUBS 0.008796f
C113 B.n21 VSUBS 0.020976f
C114 B.n22 VSUBS 0.008796f
C115 B.n23 VSUBS 0.008796f
C116 B.n24 VSUBS 0.008796f
C117 B.n25 VSUBS 0.008796f
C118 B.n26 VSUBS 0.008796f
C119 B.n27 VSUBS 0.008796f
C120 B.t10 VSUBS 0.039216f
C121 B.t11 VSUBS 0.048547f
C122 B.t9 VSUBS 0.20678f
C123 B.n28 VSUBS 0.088649f
C124 B.n29 VSUBS 0.076752f
C125 B.n30 VSUBS 0.008796f
C126 B.n31 VSUBS 0.008796f
C127 B.n32 VSUBS 0.008796f
C128 B.n33 VSUBS 0.008796f
C129 B.t1 VSUBS 0.039216f
C130 B.t2 VSUBS 0.048547f
C131 B.t0 VSUBS 0.20678f
C132 B.n34 VSUBS 0.088649f
C133 B.n35 VSUBS 0.076752f
C134 B.n36 VSUBS 0.020379f
C135 B.n37 VSUBS 0.008796f
C136 B.n38 VSUBS 0.008796f
C137 B.n39 VSUBS 0.008796f
C138 B.n40 VSUBS 0.008796f
C139 B.n41 VSUBS 0.008796f
C140 B.n42 VSUBS 0.022226f
C141 B.n43 VSUBS 0.008796f
C142 B.n44 VSUBS 0.008796f
C143 B.n45 VSUBS 0.008796f
C144 B.n46 VSUBS 0.008796f
C145 B.n47 VSUBS 0.008796f
C146 B.n48 VSUBS 0.008796f
C147 B.n49 VSUBS 0.008796f
C148 B.n50 VSUBS 0.008796f
C149 B.n51 VSUBS 0.008796f
C150 B.n52 VSUBS 0.008796f
C151 B.n53 VSUBS 0.008796f
C152 B.n54 VSUBS 0.008796f
C153 B.n55 VSUBS 0.008796f
C154 B.n56 VSUBS 0.008796f
C155 B.n57 VSUBS 0.008796f
C156 B.n58 VSUBS 0.008796f
C157 B.n59 VSUBS 0.008796f
C158 B.n60 VSUBS 0.008796f
C159 B.n61 VSUBS 0.008796f
C160 B.n62 VSUBS 0.008796f
C161 B.n63 VSUBS 0.008796f
C162 B.n64 VSUBS 0.008796f
C163 B.n65 VSUBS 0.008796f
C164 B.n66 VSUBS 0.008796f
C165 B.n67 VSUBS 0.008796f
C166 B.n68 VSUBS 0.008796f
C167 B.n69 VSUBS 0.008796f
C168 B.n70 VSUBS 0.008796f
C169 B.n71 VSUBS 0.008796f
C170 B.n72 VSUBS 0.008796f
C171 B.n73 VSUBS 0.008796f
C172 B.n74 VSUBS 0.008796f
C173 B.n75 VSUBS 0.008796f
C174 B.n76 VSUBS 0.008796f
C175 B.n77 VSUBS 0.008796f
C176 B.n78 VSUBS 0.008796f
C177 B.n79 VSUBS 0.008796f
C178 B.n80 VSUBS 0.008796f
C179 B.n81 VSUBS 0.008796f
C180 B.n82 VSUBS 0.021943f
C181 B.n83 VSUBS 0.008796f
C182 B.n84 VSUBS 0.008796f
C183 B.n85 VSUBS 0.008796f
C184 B.n86 VSUBS 0.008796f
C185 B.n87 VSUBS 0.008796f
C186 B.n88 VSUBS 0.006079f
C187 B.n89 VSUBS 0.008796f
C188 B.n90 VSUBS 0.008796f
C189 B.n91 VSUBS 0.008796f
C190 B.n92 VSUBS 0.008796f
C191 B.n93 VSUBS 0.008796f
C192 B.t5 VSUBS 0.039216f
C193 B.t4 VSUBS 0.048547f
C194 B.t3 VSUBS 0.20678f
C195 B.n94 VSUBS 0.088649f
C196 B.n95 VSUBS 0.076752f
C197 B.n96 VSUBS 0.008796f
C198 B.n97 VSUBS 0.008796f
C199 B.n98 VSUBS 0.008796f
C200 B.n99 VSUBS 0.008796f
C201 B.n100 VSUBS 0.008796f
C202 B.n101 VSUBS 0.020976f
C203 B.n102 VSUBS 0.008796f
C204 B.n103 VSUBS 0.008796f
C205 B.n104 VSUBS 0.008796f
C206 B.n105 VSUBS 0.008796f
C207 B.n106 VSUBS 0.008796f
C208 B.n107 VSUBS 0.008796f
C209 B.n108 VSUBS 0.008796f
C210 B.n109 VSUBS 0.008796f
C211 B.n110 VSUBS 0.008796f
C212 B.n111 VSUBS 0.008796f
C213 B.n112 VSUBS 0.008796f
C214 B.n113 VSUBS 0.008796f
C215 B.n114 VSUBS 0.008796f
C216 B.n115 VSUBS 0.008796f
C217 B.n116 VSUBS 0.008796f
C218 B.n117 VSUBS 0.008796f
C219 B.n118 VSUBS 0.008796f
C220 B.n119 VSUBS 0.008796f
C221 B.n120 VSUBS 0.008796f
C222 B.n121 VSUBS 0.008796f
C223 B.n122 VSUBS 0.008796f
C224 B.n123 VSUBS 0.008796f
C225 B.n124 VSUBS 0.008796f
C226 B.n125 VSUBS 0.008796f
C227 B.n126 VSUBS 0.008796f
C228 B.n127 VSUBS 0.008796f
C229 B.n128 VSUBS 0.008796f
C230 B.n129 VSUBS 0.008796f
C231 B.n130 VSUBS 0.008796f
C232 B.n131 VSUBS 0.008796f
C233 B.n132 VSUBS 0.008796f
C234 B.n133 VSUBS 0.008796f
C235 B.n134 VSUBS 0.008796f
C236 B.n135 VSUBS 0.008796f
C237 B.n136 VSUBS 0.008796f
C238 B.n137 VSUBS 0.008796f
C239 B.n138 VSUBS 0.008796f
C240 B.n139 VSUBS 0.008796f
C241 B.n140 VSUBS 0.008796f
C242 B.n141 VSUBS 0.008796f
C243 B.n142 VSUBS 0.008796f
C244 B.n143 VSUBS 0.008796f
C245 B.n144 VSUBS 0.008796f
C246 B.n145 VSUBS 0.008796f
C247 B.n146 VSUBS 0.008796f
C248 B.n147 VSUBS 0.008796f
C249 B.n148 VSUBS 0.008796f
C250 B.n149 VSUBS 0.008796f
C251 B.n150 VSUBS 0.008796f
C252 B.n151 VSUBS 0.008796f
C253 B.n152 VSUBS 0.008796f
C254 B.n153 VSUBS 0.008796f
C255 B.n154 VSUBS 0.008796f
C256 B.n155 VSUBS 0.008796f
C257 B.n156 VSUBS 0.008796f
C258 B.n157 VSUBS 0.008796f
C259 B.n158 VSUBS 0.008796f
C260 B.n159 VSUBS 0.008796f
C261 B.n160 VSUBS 0.008796f
C262 B.n161 VSUBS 0.008796f
C263 B.n162 VSUBS 0.008796f
C264 B.n163 VSUBS 0.008796f
C265 B.n164 VSUBS 0.008796f
C266 B.n165 VSUBS 0.008796f
C267 B.n166 VSUBS 0.008796f
C268 B.n167 VSUBS 0.008796f
C269 B.n168 VSUBS 0.008796f
C270 B.n169 VSUBS 0.008796f
C271 B.n170 VSUBS 0.008796f
C272 B.n171 VSUBS 0.008796f
C273 B.n172 VSUBS 0.008796f
C274 B.n173 VSUBS 0.008796f
C275 B.n174 VSUBS 0.008796f
C276 B.n175 VSUBS 0.008796f
C277 B.n176 VSUBS 0.020976f
C278 B.n177 VSUBS 0.022226f
C279 B.n178 VSUBS 0.022226f
C280 B.n179 VSUBS 0.008796f
C281 B.n180 VSUBS 0.008796f
C282 B.n181 VSUBS 0.008796f
C283 B.n182 VSUBS 0.008796f
C284 B.n183 VSUBS 0.008796f
C285 B.n184 VSUBS 0.008796f
C286 B.n185 VSUBS 0.008796f
C287 B.n186 VSUBS 0.008796f
C288 B.n187 VSUBS 0.008796f
C289 B.n188 VSUBS 0.008796f
C290 B.n189 VSUBS 0.008796f
C291 B.n190 VSUBS 0.008796f
C292 B.n191 VSUBS 0.008796f
C293 B.n192 VSUBS 0.008796f
C294 B.n193 VSUBS 0.008796f
C295 B.n194 VSUBS 0.006079f
C296 B.n195 VSUBS 0.020379f
C297 B.n196 VSUBS 0.007114f
C298 B.n197 VSUBS 0.008796f
C299 B.n198 VSUBS 0.008796f
C300 B.n199 VSUBS 0.008796f
C301 B.n200 VSUBS 0.008796f
C302 B.n201 VSUBS 0.008796f
C303 B.n202 VSUBS 0.008796f
C304 B.n203 VSUBS 0.008796f
C305 B.n204 VSUBS 0.008796f
C306 B.n205 VSUBS 0.008796f
C307 B.n206 VSUBS 0.008796f
C308 B.n207 VSUBS 0.008796f
C309 B.t8 VSUBS 0.039216f
C310 B.t7 VSUBS 0.048547f
C311 B.t6 VSUBS 0.20678f
C312 B.n208 VSUBS 0.088649f
C313 B.n209 VSUBS 0.076752f
C314 B.n210 VSUBS 0.020379f
C315 B.n211 VSUBS 0.007114f
C316 B.n212 VSUBS 0.008796f
C317 B.n213 VSUBS 0.008796f
C318 B.n214 VSUBS 0.008796f
C319 B.n215 VSUBS 0.008796f
C320 B.n216 VSUBS 0.008796f
C321 B.n217 VSUBS 0.008796f
C322 B.n218 VSUBS 0.008796f
C323 B.n219 VSUBS 0.008796f
C324 B.n220 VSUBS 0.008796f
C325 B.n221 VSUBS 0.008796f
C326 B.n222 VSUBS 0.008796f
C327 B.n223 VSUBS 0.008796f
C328 B.n224 VSUBS 0.008796f
C329 B.n225 VSUBS 0.008796f
C330 B.n226 VSUBS 0.008796f
C331 B.n227 VSUBS 0.008796f
C332 B.n228 VSUBS 0.008796f
C333 B.n229 VSUBS 0.021259f
C334 B.n230 VSUBS 0.022226f
C335 B.n231 VSUBS 0.020976f
C336 B.n232 VSUBS 0.008796f
C337 B.n233 VSUBS 0.008796f
C338 B.n234 VSUBS 0.008796f
C339 B.n235 VSUBS 0.008796f
C340 B.n236 VSUBS 0.008796f
C341 B.n237 VSUBS 0.008796f
C342 B.n238 VSUBS 0.008796f
C343 B.n239 VSUBS 0.008796f
C344 B.n240 VSUBS 0.008796f
C345 B.n241 VSUBS 0.008796f
C346 B.n242 VSUBS 0.008796f
C347 B.n243 VSUBS 0.008796f
C348 B.n244 VSUBS 0.008796f
C349 B.n245 VSUBS 0.008796f
C350 B.n246 VSUBS 0.008796f
C351 B.n247 VSUBS 0.008796f
C352 B.n248 VSUBS 0.008796f
C353 B.n249 VSUBS 0.008796f
C354 B.n250 VSUBS 0.008796f
C355 B.n251 VSUBS 0.008796f
C356 B.n252 VSUBS 0.008796f
C357 B.n253 VSUBS 0.008796f
C358 B.n254 VSUBS 0.008796f
C359 B.n255 VSUBS 0.008796f
C360 B.n256 VSUBS 0.008796f
C361 B.n257 VSUBS 0.008796f
C362 B.n258 VSUBS 0.008796f
C363 B.n259 VSUBS 0.008796f
C364 B.n260 VSUBS 0.008796f
C365 B.n261 VSUBS 0.008796f
C366 B.n262 VSUBS 0.008796f
C367 B.n263 VSUBS 0.008796f
C368 B.n264 VSUBS 0.008796f
C369 B.n265 VSUBS 0.008796f
C370 B.n266 VSUBS 0.008796f
C371 B.n267 VSUBS 0.008796f
C372 B.n268 VSUBS 0.008796f
C373 B.n269 VSUBS 0.008796f
C374 B.n270 VSUBS 0.008796f
C375 B.n271 VSUBS 0.008796f
C376 B.n272 VSUBS 0.008796f
C377 B.n273 VSUBS 0.008796f
C378 B.n274 VSUBS 0.008796f
C379 B.n275 VSUBS 0.008796f
C380 B.n276 VSUBS 0.008796f
C381 B.n277 VSUBS 0.008796f
C382 B.n278 VSUBS 0.008796f
C383 B.n279 VSUBS 0.008796f
C384 B.n280 VSUBS 0.008796f
C385 B.n281 VSUBS 0.008796f
C386 B.n282 VSUBS 0.008796f
C387 B.n283 VSUBS 0.008796f
C388 B.n284 VSUBS 0.008796f
C389 B.n285 VSUBS 0.008796f
C390 B.n286 VSUBS 0.008796f
C391 B.n287 VSUBS 0.008796f
C392 B.n288 VSUBS 0.008796f
C393 B.n289 VSUBS 0.008796f
C394 B.n290 VSUBS 0.008796f
C395 B.n291 VSUBS 0.008796f
C396 B.n292 VSUBS 0.008796f
C397 B.n293 VSUBS 0.008796f
C398 B.n294 VSUBS 0.008796f
C399 B.n295 VSUBS 0.008796f
C400 B.n296 VSUBS 0.008796f
C401 B.n297 VSUBS 0.008796f
C402 B.n298 VSUBS 0.008796f
C403 B.n299 VSUBS 0.008796f
C404 B.n300 VSUBS 0.008796f
C405 B.n301 VSUBS 0.008796f
C406 B.n302 VSUBS 0.008796f
C407 B.n303 VSUBS 0.008796f
C408 B.n304 VSUBS 0.008796f
C409 B.n305 VSUBS 0.008796f
C410 B.n306 VSUBS 0.008796f
C411 B.n307 VSUBS 0.008796f
C412 B.n308 VSUBS 0.008796f
C413 B.n309 VSUBS 0.008796f
C414 B.n310 VSUBS 0.008796f
C415 B.n311 VSUBS 0.008796f
C416 B.n312 VSUBS 0.008796f
C417 B.n313 VSUBS 0.008796f
C418 B.n314 VSUBS 0.008796f
C419 B.n315 VSUBS 0.008796f
C420 B.n316 VSUBS 0.008796f
C421 B.n317 VSUBS 0.008796f
C422 B.n318 VSUBS 0.008796f
C423 B.n319 VSUBS 0.008796f
C424 B.n320 VSUBS 0.008796f
C425 B.n321 VSUBS 0.008796f
C426 B.n322 VSUBS 0.008796f
C427 B.n323 VSUBS 0.008796f
C428 B.n324 VSUBS 0.008796f
C429 B.n325 VSUBS 0.008796f
C430 B.n326 VSUBS 0.008796f
C431 B.n327 VSUBS 0.008796f
C432 B.n328 VSUBS 0.008796f
C433 B.n329 VSUBS 0.008796f
C434 B.n330 VSUBS 0.008796f
C435 B.n331 VSUBS 0.008796f
C436 B.n332 VSUBS 0.008796f
C437 B.n333 VSUBS 0.008796f
C438 B.n334 VSUBS 0.008796f
C439 B.n335 VSUBS 0.008796f
C440 B.n336 VSUBS 0.008796f
C441 B.n337 VSUBS 0.008796f
C442 B.n338 VSUBS 0.008796f
C443 B.n339 VSUBS 0.008796f
C444 B.n340 VSUBS 0.008796f
C445 B.n341 VSUBS 0.008796f
C446 B.n342 VSUBS 0.008796f
C447 B.n343 VSUBS 0.008796f
C448 B.n344 VSUBS 0.008796f
C449 B.n345 VSUBS 0.008796f
C450 B.n346 VSUBS 0.008796f
C451 B.n347 VSUBS 0.008796f
C452 B.n348 VSUBS 0.008796f
C453 B.n349 VSUBS 0.020976f
C454 B.n350 VSUBS 0.020976f
C455 B.n351 VSUBS 0.022226f
C456 B.n352 VSUBS 0.008796f
C457 B.n353 VSUBS 0.008796f
C458 B.n354 VSUBS 0.008796f
C459 B.n355 VSUBS 0.008796f
C460 B.n356 VSUBS 0.008796f
C461 B.n357 VSUBS 0.008796f
C462 B.n358 VSUBS 0.008796f
C463 B.n359 VSUBS 0.008796f
C464 B.n360 VSUBS 0.008796f
C465 B.n361 VSUBS 0.008796f
C466 B.n362 VSUBS 0.008796f
C467 B.n363 VSUBS 0.008796f
C468 B.n364 VSUBS 0.008796f
C469 B.n365 VSUBS 0.008796f
C470 B.n366 VSUBS 0.008796f
C471 B.n367 VSUBS 0.006079f
C472 B.n368 VSUBS 0.008796f
C473 B.n369 VSUBS 0.008796f
C474 B.n370 VSUBS 0.007114f
C475 B.n371 VSUBS 0.008796f
C476 B.n372 VSUBS 0.008796f
C477 B.n373 VSUBS 0.008796f
C478 B.n374 VSUBS 0.008796f
C479 B.n375 VSUBS 0.008796f
C480 B.n376 VSUBS 0.008796f
C481 B.n377 VSUBS 0.008796f
C482 B.n378 VSUBS 0.008796f
C483 B.n379 VSUBS 0.008796f
C484 B.n380 VSUBS 0.008796f
C485 B.n381 VSUBS 0.008796f
C486 B.n382 VSUBS 0.007114f
C487 B.n383 VSUBS 0.020379f
C488 B.n384 VSUBS 0.006079f
C489 B.n385 VSUBS 0.008796f
C490 B.n386 VSUBS 0.008796f
C491 B.n387 VSUBS 0.008796f
C492 B.n388 VSUBS 0.008796f
C493 B.n389 VSUBS 0.008796f
C494 B.n390 VSUBS 0.008796f
C495 B.n391 VSUBS 0.008796f
C496 B.n392 VSUBS 0.008796f
C497 B.n393 VSUBS 0.008796f
C498 B.n394 VSUBS 0.008796f
C499 B.n395 VSUBS 0.008796f
C500 B.n396 VSUBS 0.008796f
C501 B.n397 VSUBS 0.008796f
C502 B.n398 VSUBS 0.008796f
C503 B.n399 VSUBS 0.008796f
C504 B.n400 VSUBS 0.022226f
C505 B.n401 VSUBS 0.022226f
C506 B.n402 VSUBS 0.020976f
C507 B.n403 VSUBS 0.008796f
C508 B.n404 VSUBS 0.008796f
C509 B.n405 VSUBS 0.008796f
C510 B.n406 VSUBS 0.008796f
C511 B.n407 VSUBS 0.008796f
C512 B.n408 VSUBS 0.008796f
C513 B.n409 VSUBS 0.008796f
C514 B.n410 VSUBS 0.008796f
C515 B.n411 VSUBS 0.008796f
C516 B.n412 VSUBS 0.008796f
C517 B.n413 VSUBS 0.008796f
C518 B.n414 VSUBS 0.008796f
C519 B.n415 VSUBS 0.008796f
C520 B.n416 VSUBS 0.008796f
C521 B.n417 VSUBS 0.008796f
C522 B.n418 VSUBS 0.008796f
C523 B.n419 VSUBS 0.008796f
C524 B.n420 VSUBS 0.008796f
C525 B.n421 VSUBS 0.008796f
C526 B.n422 VSUBS 0.008796f
C527 B.n423 VSUBS 0.008796f
C528 B.n424 VSUBS 0.008796f
C529 B.n425 VSUBS 0.008796f
C530 B.n426 VSUBS 0.008796f
C531 B.n427 VSUBS 0.008796f
C532 B.n428 VSUBS 0.008796f
C533 B.n429 VSUBS 0.008796f
C534 B.n430 VSUBS 0.008796f
C535 B.n431 VSUBS 0.008796f
C536 B.n432 VSUBS 0.008796f
C537 B.n433 VSUBS 0.008796f
C538 B.n434 VSUBS 0.008796f
C539 B.n435 VSUBS 0.008796f
C540 B.n436 VSUBS 0.008796f
C541 B.n437 VSUBS 0.008796f
C542 B.n438 VSUBS 0.008796f
C543 B.n439 VSUBS 0.008796f
C544 B.n440 VSUBS 0.008796f
C545 B.n441 VSUBS 0.008796f
C546 B.n442 VSUBS 0.008796f
C547 B.n443 VSUBS 0.008796f
C548 B.n444 VSUBS 0.008796f
C549 B.n445 VSUBS 0.008796f
C550 B.n446 VSUBS 0.008796f
C551 B.n447 VSUBS 0.008796f
C552 B.n448 VSUBS 0.008796f
C553 B.n449 VSUBS 0.008796f
C554 B.n450 VSUBS 0.008796f
C555 B.n451 VSUBS 0.008796f
C556 B.n452 VSUBS 0.008796f
C557 B.n453 VSUBS 0.008796f
C558 B.n454 VSUBS 0.008796f
C559 B.n455 VSUBS 0.008796f
C560 B.n456 VSUBS 0.008796f
C561 B.n457 VSUBS 0.008796f
C562 B.n458 VSUBS 0.008796f
C563 B.n459 VSUBS 0.011478f
C564 B.n460 VSUBS 0.012227f
C565 B.n461 VSUBS 0.024314f
C566 VTAIL.t2 VSUBS 0.043907f
C567 VTAIL.t6 VSUBS 0.043907f
C568 VTAIL.n0 VSUBS 0.158854f
C569 VTAIL.n1 VSUBS 0.480728f
C570 VTAIL.n2 VSUBS 0.03203f
C571 VTAIL.n3 VSUBS 0.085813f
C572 VTAIL.t3 VSUBS 0.082414f
C573 VTAIL.n4 VSUBS 0.079343f
C574 VTAIL.n5 VSUBS 0.02037f
C575 VTAIL.n6 VSUBS 0.016227f
C576 VTAIL.n7 VSUBS 0.182859f
C577 VTAIL.n8 VSUBS 0.044744f
C578 VTAIL.n9 VSUBS 0.255582f
C579 VTAIL.n10 VSUBS 0.03203f
C580 VTAIL.n11 VSUBS 0.085813f
C581 VTAIL.t9 VSUBS 0.082414f
C582 VTAIL.n12 VSUBS 0.079343f
C583 VTAIL.n13 VSUBS 0.02037f
C584 VTAIL.n14 VSUBS 0.016227f
C585 VTAIL.n15 VSUBS 0.182859f
C586 VTAIL.n16 VSUBS 0.044744f
C587 VTAIL.n17 VSUBS 0.255582f
C588 VTAIL.t8 VSUBS 0.043907f
C589 VTAIL.t14 VSUBS 0.043907f
C590 VTAIL.n18 VSUBS 0.158854f
C591 VTAIL.n19 VSUBS 0.65541f
C592 VTAIL.n20 VSUBS 0.03203f
C593 VTAIL.n21 VSUBS 0.085813f
C594 VTAIL.t15 VSUBS 0.082414f
C595 VTAIL.n22 VSUBS 0.079343f
C596 VTAIL.n23 VSUBS 0.02037f
C597 VTAIL.n24 VSUBS 0.016227f
C598 VTAIL.n25 VSUBS 0.182859f
C599 VTAIL.n26 VSUBS 0.044744f
C600 VTAIL.n27 VSUBS 0.954741f
C601 VTAIL.n28 VSUBS 0.03203f
C602 VTAIL.n29 VSUBS 0.085813f
C603 VTAIL.t4 VSUBS 0.082414f
C604 VTAIL.n30 VSUBS 0.079343f
C605 VTAIL.n31 VSUBS 0.02037f
C606 VTAIL.n32 VSUBS 0.016227f
C607 VTAIL.n33 VSUBS 0.182859f
C608 VTAIL.n34 VSUBS 0.044744f
C609 VTAIL.n35 VSUBS 0.954741f
C610 VTAIL.t0 VSUBS 0.043907f
C611 VTAIL.t5 VSUBS 0.043907f
C612 VTAIL.n36 VSUBS 0.158855f
C613 VTAIL.n37 VSUBS 0.655409f
C614 VTAIL.n38 VSUBS 0.03203f
C615 VTAIL.n39 VSUBS 0.085813f
C616 VTAIL.t1 VSUBS 0.082414f
C617 VTAIL.n40 VSUBS 0.079343f
C618 VTAIL.n41 VSUBS 0.02037f
C619 VTAIL.n42 VSUBS 0.016227f
C620 VTAIL.n43 VSUBS 0.182859f
C621 VTAIL.n44 VSUBS 0.044744f
C622 VTAIL.n45 VSUBS 0.255582f
C623 VTAIL.n46 VSUBS 0.03203f
C624 VTAIL.n47 VSUBS 0.085813f
C625 VTAIL.t12 VSUBS 0.082414f
C626 VTAIL.n48 VSUBS 0.079343f
C627 VTAIL.n49 VSUBS 0.02037f
C628 VTAIL.n50 VSUBS 0.016227f
C629 VTAIL.n51 VSUBS 0.182859f
C630 VTAIL.n52 VSUBS 0.044744f
C631 VTAIL.n53 VSUBS 0.255582f
C632 VTAIL.t10 VSUBS 0.043907f
C633 VTAIL.t13 VSUBS 0.043907f
C634 VTAIL.n54 VSUBS 0.158855f
C635 VTAIL.n55 VSUBS 0.655409f
C636 VTAIL.n56 VSUBS 0.03203f
C637 VTAIL.n57 VSUBS 0.085813f
C638 VTAIL.t11 VSUBS 0.082414f
C639 VTAIL.n58 VSUBS 0.079343f
C640 VTAIL.n59 VSUBS 0.02037f
C641 VTAIL.n60 VSUBS 0.016227f
C642 VTAIL.n61 VSUBS 0.182859f
C643 VTAIL.n62 VSUBS 0.044744f
C644 VTAIL.n63 VSUBS 0.954741f
C645 VTAIL.n64 VSUBS 0.03203f
C646 VTAIL.n65 VSUBS 0.085813f
C647 VTAIL.t7 VSUBS 0.082414f
C648 VTAIL.n66 VSUBS 0.079343f
C649 VTAIL.n67 VSUBS 0.02037f
C650 VTAIL.n68 VSUBS 0.016227f
C651 VTAIL.n69 VSUBS 0.182859f
C652 VTAIL.n70 VSUBS 0.044744f
C653 VTAIL.n71 VSUBS 0.949079f
C654 VDD1.t0 VSUBS 0.024697f
C655 VDD1.t3 VSUBS 0.024697f
C656 VDD1.n0 VSUBS 0.106252f
C657 VDD1.t7 VSUBS 0.024697f
C658 VDD1.t6 VSUBS 0.024697f
C659 VDD1.n1 VSUBS 0.106041f
C660 VDD1.t5 VSUBS 0.024697f
C661 VDD1.t4 VSUBS 0.024697f
C662 VDD1.n2 VSUBS 0.106041f
C663 VDD1.n3 VSUBS 1.61326f
C664 VDD1.t2 VSUBS 0.024697f
C665 VDD1.t1 VSUBS 0.024697f
C666 VDD1.n4 VSUBS 0.104628f
C667 VDD1.n5 VSUBS 1.33063f
C668 VP.n0 VSUBS 0.071699f
C669 VP.t6 VSUBS 0.417943f
C670 VP.n1 VSUBS 0.099328f
C671 VP.n2 VSUBS 0.054386f
C672 VP.t1 VSUBS 0.417943f
C673 VP.n3 VSUBS 0.079059f
C674 VP.n4 VSUBS 0.054386f
C675 VP.t7 VSUBS 0.417943f
C676 VP.n5 VSUBS 0.051278f
C677 VP.n6 VSUBS 0.071699f
C678 VP.t4 VSUBS 0.417943f
C679 VP.n7 VSUBS 0.099328f
C680 VP.n8 VSUBS 0.054386f
C681 VP.t2 VSUBS 0.417943f
C682 VP.n9 VSUBS 0.079059f
C683 VP.t3 VSUBS 0.684801f
C684 VP.n10 VSUBS 0.322061f
C685 VP.t5 VSUBS 0.417943f
C686 VP.n11 VSUBS 0.348539f
C687 VP.n12 VSUBS 0.083428f
C688 VP.n13 VSUBS 0.398417f
C689 VP.n14 VSUBS 0.054386f
C690 VP.n15 VSUBS 0.054386f
C691 VP.n16 VSUBS 0.079059f
C692 VP.n17 VSUBS 0.083428f
C693 VP.n18 VSUBS 0.219925f
C694 VP.n19 VSUBS 0.068491f
C695 VP.n20 VSUBS 0.054386f
C696 VP.n21 VSUBS 0.054386f
C697 VP.n22 VSUBS 0.054386f
C698 VP.n23 VSUBS 0.051278f
C699 VP.n24 VSUBS 0.105876f
C700 VP.n25 VSUBS 0.382012f
C701 VP.n26 VSUBS 2.06769f
C702 VP.n27 VSUBS 2.11722f
C703 VP.t0 VSUBS 0.417943f
C704 VP.n28 VSUBS 0.382012f
C705 VP.n29 VSUBS 0.105876f
C706 VP.n30 VSUBS 0.071699f
C707 VP.n31 VSUBS 0.054386f
C708 VP.n32 VSUBS 0.054386f
C709 VP.n33 VSUBS 0.099328f
C710 VP.n34 VSUBS 0.068491f
C711 VP.n35 VSUBS 0.219925f
C712 VP.n36 VSUBS 0.083428f
C713 VP.n37 VSUBS 0.054386f
C714 VP.n38 VSUBS 0.054386f
C715 VP.n39 VSUBS 0.054386f
C716 VP.n40 VSUBS 0.079059f
C717 VP.n41 VSUBS 0.083428f
C718 VP.n42 VSUBS 0.219925f
C719 VP.n43 VSUBS 0.068491f
C720 VP.n44 VSUBS 0.054386f
C721 VP.n45 VSUBS 0.054386f
C722 VP.n46 VSUBS 0.054386f
C723 VP.n47 VSUBS 0.051278f
C724 VP.n48 VSUBS 0.105876f
C725 VP.n49 VSUBS 0.382012f
C726 VP.n50 VSUBS 0.059119f
.ends

