* NGSPICE file created from diff_pair_sample_0944.ext - technology: sky130A

.subckt diff_pair_sample_0944 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=1.6071 pd=10.07 as=3.7986 ps=20.26 w=9.74 l=1.7
X1 VTAIL.t3 VN.t0 VDD2.t3 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=3.7986 pd=20.26 as=1.6071 ps=10.07 w=9.74 l=1.7
X2 VTAIL.t6 VP.t1 VDD1.t2 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=3.7986 pd=20.26 as=1.6071 ps=10.07 w=9.74 l=1.7
X3 VDD2.t2 VN.t1 VTAIL.t0 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=1.6071 pd=10.07 as=3.7986 ps=20.26 w=9.74 l=1.7
X4 B.t11 B.t9 B.t10 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=3.7986 pd=20.26 as=0 ps=0 w=9.74 l=1.7
X5 VTAIL.t7 VP.t2 VDD1.t1 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=3.7986 pd=20.26 as=1.6071 ps=10.07 w=9.74 l=1.7
X6 VDD2.t1 VN.t2 VTAIL.t1 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=1.6071 pd=10.07 as=3.7986 ps=20.26 w=9.74 l=1.7
X7 B.t8 B.t6 B.t7 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=3.7986 pd=20.26 as=0 ps=0 w=9.74 l=1.7
X8 VDD1.t0 VP.t3 VTAIL.t4 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=1.6071 pd=10.07 as=3.7986 ps=20.26 w=9.74 l=1.7
X9 VTAIL.t2 VN.t3 VDD2.t0 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=3.7986 pd=20.26 as=1.6071 ps=10.07 w=9.74 l=1.7
X10 B.t5 B.t3 B.t4 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=3.7986 pd=20.26 as=0 ps=0 w=9.74 l=1.7
X11 B.t2 B.t0 B.t1 w_n2188_n2916# sky130_fd_pr__pfet_01v8 ad=3.7986 pd=20.26 as=0 ps=0 w=9.74 l=1.7
R0 VP.n5 VP.n4 184.913
R1 VP.n14 VP.n13 184.913
R2 VP.n3 VP.t1 173.042
R3 VP.n3 VP.t0 172.623
R4 VP.n12 VP.n0 161.3
R5 VP.n11 VP.n10 161.3
R6 VP.n9 VP.n1 161.3
R7 VP.n8 VP.n7 161.3
R8 VP.n6 VP.n2 161.3
R9 VP.n5 VP.t2 138.079
R10 VP.n13 VP.t3 138.079
R11 VP.n4 VP.n3 51.2586
R12 VP.n7 VP.n1 40.4106
R13 VP.n11 VP.n1 40.4106
R14 VP.n7 VP.n6 24.3439
R15 VP.n12 VP.n11 24.3439
R16 VP.n6 VP.n5 0.730803
R17 VP.n13 VP.n12 0.730803
R18 VP.n4 VP.n2 0.189894
R19 VP.n8 VP.n2 0.189894
R20 VP.n9 VP.n8 0.189894
R21 VP.n10 VP.n9 0.189894
R22 VP.n10 VP.n0 0.189894
R23 VP.n14 VP.n0 0.189894
R24 VP VP.n14 0.0516364
R25 VTAIL.n5 VTAIL.t6 67.194
R26 VTAIL.n4 VTAIL.t0 67.194
R27 VTAIL.n3 VTAIL.t3 67.194
R28 VTAIL.n7 VTAIL.t1 67.1938
R29 VTAIL.n0 VTAIL.t2 67.1938
R30 VTAIL.n1 VTAIL.t4 67.1938
R31 VTAIL.n2 VTAIL.t7 67.1938
R32 VTAIL.n6 VTAIL.t5 67.1938
R33 VTAIL.n7 VTAIL.n6 22.5134
R34 VTAIL.n3 VTAIL.n2 22.5134
R35 VTAIL.n4 VTAIL.n3 1.7505
R36 VTAIL.n6 VTAIL.n5 1.7505
R37 VTAIL.n2 VTAIL.n1 1.7505
R38 VTAIL VTAIL.n0 0.93369
R39 VTAIL VTAIL.n7 0.81731
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 VDD1 VDD1.n1 118.421
R43 VDD1 VDD1.n0 80.5935
R44 VDD1.n0 VDD1.t2 3.33777
R45 VDD1.n0 VDD1.t3 3.33777
R46 VDD1.n1 VDD1.t1 3.33777
R47 VDD1.n1 VDD1.t0 3.33777
R48 VN.n0 VN.t3 173.042
R49 VN.n1 VN.t1 173.042
R50 VN.n0 VN.t2 172.623
R51 VN.n1 VN.t0 172.623
R52 VN VN.n1 51.6393
R53 VN VN.n0 9.58248
R54 VDD2.n2 VDD2.n0 117.897
R55 VDD2.n2 VDD2.n1 80.5354
R56 VDD2.n1 VDD2.t3 3.33777
R57 VDD2.n1 VDD2.t2 3.33777
R58 VDD2.n0 VDD2.t0 3.33777
R59 VDD2.n0 VDD2.t1 3.33777
R60 VDD2 VDD2.n2 0.0586897
R61 B.n380 B.n59 585
R62 B.n382 B.n381 585
R63 B.n383 B.n58 585
R64 B.n385 B.n384 585
R65 B.n386 B.n57 585
R66 B.n388 B.n387 585
R67 B.n389 B.n56 585
R68 B.n391 B.n390 585
R69 B.n392 B.n55 585
R70 B.n394 B.n393 585
R71 B.n395 B.n54 585
R72 B.n397 B.n396 585
R73 B.n398 B.n53 585
R74 B.n400 B.n399 585
R75 B.n401 B.n52 585
R76 B.n403 B.n402 585
R77 B.n404 B.n51 585
R78 B.n406 B.n405 585
R79 B.n407 B.n50 585
R80 B.n409 B.n408 585
R81 B.n410 B.n49 585
R82 B.n412 B.n411 585
R83 B.n413 B.n48 585
R84 B.n415 B.n414 585
R85 B.n416 B.n47 585
R86 B.n418 B.n417 585
R87 B.n419 B.n46 585
R88 B.n421 B.n420 585
R89 B.n422 B.n45 585
R90 B.n424 B.n423 585
R91 B.n425 B.n44 585
R92 B.n427 B.n426 585
R93 B.n428 B.n43 585
R94 B.n430 B.n429 585
R95 B.n431 B.n40 585
R96 B.n434 B.n433 585
R97 B.n435 B.n39 585
R98 B.n437 B.n436 585
R99 B.n438 B.n38 585
R100 B.n440 B.n439 585
R101 B.n441 B.n37 585
R102 B.n443 B.n442 585
R103 B.n444 B.n33 585
R104 B.n446 B.n445 585
R105 B.n447 B.n32 585
R106 B.n449 B.n448 585
R107 B.n450 B.n31 585
R108 B.n452 B.n451 585
R109 B.n453 B.n30 585
R110 B.n455 B.n454 585
R111 B.n456 B.n29 585
R112 B.n458 B.n457 585
R113 B.n459 B.n28 585
R114 B.n461 B.n460 585
R115 B.n462 B.n27 585
R116 B.n464 B.n463 585
R117 B.n465 B.n26 585
R118 B.n467 B.n466 585
R119 B.n468 B.n25 585
R120 B.n470 B.n469 585
R121 B.n471 B.n24 585
R122 B.n473 B.n472 585
R123 B.n474 B.n23 585
R124 B.n476 B.n475 585
R125 B.n477 B.n22 585
R126 B.n479 B.n478 585
R127 B.n480 B.n21 585
R128 B.n482 B.n481 585
R129 B.n483 B.n20 585
R130 B.n485 B.n484 585
R131 B.n486 B.n19 585
R132 B.n488 B.n487 585
R133 B.n489 B.n18 585
R134 B.n491 B.n490 585
R135 B.n492 B.n17 585
R136 B.n494 B.n493 585
R137 B.n495 B.n16 585
R138 B.n497 B.n496 585
R139 B.n498 B.n15 585
R140 B.n379 B.n378 585
R141 B.n377 B.n60 585
R142 B.n376 B.n375 585
R143 B.n374 B.n61 585
R144 B.n373 B.n372 585
R145 B.n371 B.n62 585
R146 B.n370 B.n369 585
R147 B.n368 B.n63 585
R148 B.n367 B.n366 585
R149 B.n365 B.n64 585
R150 B.n364 B.n363 585
R151 B.n362 B.n65 585
R152 B.n361 B.n360 585
R153 B.n359 B.n66 585
R154 B.n358 B.n357 585
R155 B.n356 B.n67 585
R156 B.n355 B.n354 585
R157 B.n353 B.n68 585
R158 B.n352 B.n351 585
R159 B.n350 B.n69 585
R160 B.n349 B.n348 585
R161 B.n347 B.n70 585
R162 B.n346 B.n345 585
R163 B.n344 B.n71 585
R164 B.n343 B.n342 585
R165 B.n341 B.n72 585
R166 B.n340 B.n339 585
R167 B.n338 B.n73 585
R168 B.n337 B.n336 585
R169 B.n335 B.n74 585
R170 B.n334 B.n333 585
R171 B.n332 B.n75 585
R172 B.n331 B.n330 585
R173 B.n329 B.n76 585
R174 B.n328 B.n327 585
R175 B.n326 B.n77 585
R176 B.n325 B.n324 585
R177 B.n323 B.n78 585
R178 B.n322 B.n321 585
R179 B.n320 B.n79 585
R180 B.n319 B.n318 585
R181 B.n317 B.n80 585
R182 B.n316 B.n315 585
R183 B.n314 B.n81 585
R184 B.n313 B.n312 585
R185 B.n311 B.n82 585
R186 B.n310 B.n309 585
R187 B.n308 B.n83 585
R188 B.n307 B.n306 585
R189 B.n305 B.n84 585
R190 B.n304 B.n303 585
R191 B.n302 B.n85 585
R192 B.n301 B.n300 585
R193 B.n178 B.n127 585
R194 B.n180 B.n179 585
R195 B.n181 B.n126 585
R196 B.n183 B.n182 585
R197 B.n184 B.n125 585
R198 B.n186 B.n185 585
R199 B.n187 B.n124 585
R200 B.n189 B.n188 585
R201 B.n190 B.n123 585
R202 B.n192 B.n191 585
R203 B.n193 B.n122 585
R204 B.n195 B.n194 585
R205 B.n196 B.n121 585
R206 B.n198 B.n197 585
R207 B.n199 B.n120 585
R208 B.n201 B.n200 585
R209 B.n202 B.n119 585
R210 B.n204 B.n203 585
R211 B.n205 B.n118 585
R212 B.n207 B.n206 585
R213 B.n208 B.n117 585
R214 B.n210 B.n209 585
R215 B.n211 B.n116 585
R216 B.n213 B.n212 585
R217 B.n214 B.n115 585
R218 B.n216 B.n215 585
R219 B.n217 B.n114 585
R220 B.n219 B.n218 585
R221 B.n220 B.n113 585
R222 B.n222 B.n221 585
R223 B.n223 B.n112 585
R224 B.n225 B.n224 585
R225 B.n226 B.n111 585
R226 B.n228 B.n227 585
R227 B.n229 B.n108 585
R228 B.n232 B.n231 585
R229 B.n233 B.n107 585
R230 B.n235 B.n234 585
R231 B.n236 B.n106 585
R232 B.n238 B.n237 585
R233 B.n239 B.n105 585
R234 B.n241 B.n240 585
R235 B.n242 B.n104 585
R236 B.n247 B.n246 585
R237 B.n248 B.n103 585
R238 B.n250 B.n249 585
R239 B.n251 B.n102 585
R240 B.n253 B.n252 585
R241 B.n254 B.n101 585
R242 B.n256 B.n255 585
R243 B.n257 B.n100 585
R244 B.n259 B.n258 585
R245 B.n260 B.n99 585
R246 B.n262 B.n261 585
R247 B.n263 B.n98 585
R248 B.n265 B.n264 585
R249 B.n266 B.n97 585
R250 B.n268 B.n267 585
R251 B.n269 B.n96 585
R252 B.n271 B.n270 585
R253 B.n272 B.n95 585
R254 B.n274 B.n273 585
R255 B.n275 B.n94 585
R256 B.n277 B.n276 585
R257 B.n278 B.n93 585
R258 B.n280 B.n279 585
R259 B.n281 B.n92 585
R260 B.n283 B.n282 585
R261 B.n284 B.n91 585
R262 B.n286 B.n285 585
R263 B.n287 B.n90 585
R264 B.n289 B.n288 585
R265 B.n290 B.n89 585
R266 B.n292 B.n291 585
R267 B.n293 B.n88 585
R268 B.n295 B.n294 585
R269 B.n296 B.n87 585
R270 B.n298 B.n297 585
R271 B.n299 B.n86 585
R272 B.n177 B.n176 585
R273 B.n175 B.n128 585
R274 B.n174 B.n173 585
R275 B.n172 B.n129 585
R276 B.n171 B.n170 585
R277 B.n169 B.n130 585
R278 B.n168 B.n167 585
R279 B.n166 B.n131 585
R280 B.n165 B.n164 585
R281 B.n163 B.n132 585
R282 B.n162 B.n161 585
R283 B.n160 B.n133 585
R284 B.n159 B.n158 585
R285 B.n157 B.n134 585
R286 B.n156 B.n155 585
R287 B.n154 B.n135 585
R288 B.n153 B.n152 585
R289 B.n151 B.n136 585
R290 B.n150 B.n149 585
R291 B.n148 B.n137 585
R292 B.n147 B.n146 585
R293 B.n145 B.n138 585
R294 B.n144 B.n143 585
R295 B.n142 B.n139 585
R296 B.n141 B.n140 585
R297 B.n2 B.n0 585
R298 B.n537 B.n1 585
R299 B.n536 B.n535 585
R300 B.n534 B.n3 585
R301 B.n533 B.n532 585
R302 B.n531 B.n4 585
R303 B.n530 B.n529 585
R304 B.n528 B.n5 585
R305 B.n527 B.n526 585
R306 B.n525 B.n6 585
R307 B.n524 B.n523 585
R308 B.n522 B.n7 585
R309 B.n521 B.n520 585
R310 B.n519 B.n8 585
R311 B.n518 B.n517 585
R312 B.n516 B.n9 585
R313 B.n515 B.n514 585
R314 B.n513 B.n10 585
R315 B.n512 B.n511 585
R316 B.n510 B.n11 585
R317 B.n509 B.n508 585
R318 B.n507 B.n12 585
R319 B.n506 B.n505 585
R320 B.n504 B.n13 585
R321 B.n503 B.n502 585
R322 B.n501 B.n14 585
R323 B.n500 B.n499 585
R324 B.n539 B.n538 585
R325 B.n178 B.n177 545.355
R326 B.n500 B.n15 545.355
R327 B.n301 B.n86 545.355
R328 B.n380 B.n379 545.355
R329 B.n243 B.t0 344.193
R330 B.n109 B.t6 344.193
R331 B.n34 B.t3 344.193
R332 B.n41 B.t9 344.193
R333 B.n177 B.n128 163.367
R334 B.n173 B.n128 163.367
R335 B.n173 B.n172 163.367
R336 B.n172 B.n171 163.367
R337 B.n171 B.n130 163.367
R338 B.n167 B.n130 163.367
R339 B.n167 B.n166 163.367
R340 B.n166 B.n165 163.367
R341 B.n165 B.n132 163.367
R342 B.n161 B.n132 163.367
R343 B.n161 B.n160 163.367
R344 B.n160 B.n159 163.367
R345 B.n159 B.n134 163.367
R346 B.n155 B.n134 163.367
R347 B.n155 B.n154 163.367
R348 B.n154 B.n153 163.367
R349 B.n153 B.n136 163.367
R350 B.n149 B.n136 163.367
R351 B.n149 B.n148 163.367
R352 B.n148 B.n147 163.367
R353 B.n147 B.n138 163.367
R354 B.n143 B.n138 163.367
R355 B.n143 B.n142 163.367
R356 B.n142 B.n141 163.367
R357 B.n141 B.n2 163.367
R358 B.n538 B.n2 163.367
R359 B.n538 B.n537 163.367
R360 B.n537 B.n536 163.367
R361 B.n536 B.n3 163.367
R362 B.n532 B.n3 163.367
R363 B.n532 B.n531 163.367
R364 B.n531 B.n530 163.367
R365 B.n530 B.n5 163.367
R366 B.n526 B.n5 163.367
R367 B.n526 B.n525 163.367
R368 B.n525 B.n524 163.367
R369 B.n524 B.n7 163.367
R370 B.n520 B.n7 163.367
R371 B.n520 B.n519 163.367
R372 B.n519 B.n518 163.367
R373 B.n518 B.n9 163.367
R374 B.n514 B.n9 163.367
R375 B.n514 B.n513 163.367
R376 B.n513 B.n512 163.367
R377 B.n512 B.n11 163.367
R378 B.n508 B.n11 163.367
R379 B.n508 B.n507 163.367
R380 B.n507 B.n506 163.367
R381 B.n506 B.n13 163.367
R382 B.n502 B.n13 163.367
R383 B.n502 B.n501 163.367
R384 B.n501 B.n500 163.367
R385 B.n179 B.n178 163.367
R386 B.n179 B.n126 163.367
R387 B.n183 B.n126 163.367
R388 B.n184 B.n183 163.367
R389 B.n185 B.n184 163.367
R390 B.n185 B.n124 163.367
R391 B.n189 B.n124 163.367
R392 B.n190 B.n189 163.367
R393 B.n191 B.n190 163.367
R394 B.n191 B.n122 163.367
R395 B.n195 B.n122 163.367
R396 B.n196 B.n195 163.367
R397 B.n197 B.n196 163.367
R398 B.n197 B.n120 163.367
R399 B.n201 B.n120 163.367
R400 B.n202 B.n201 163.367
R401 B.n203 B.n202 163.367
R402 B.n203 B.n118 163.367
R403 B.n207 B.n118 163.367
R404 B.n208 B.n207 163.367
R405 B.n209 B.n208 163.367
R406 B.n209 B.n116 163.367
R407 B.n213 B.n116 163.367
R408 B.n214 B.n213 163.367
R409 B.n215 B.n214 163.367
R410 B.n215 B.n114 163.367
R411 B.n219 B.n114 163.367
R412 B.n220 B.n219 163.367
R413 B.n221 B.n220 163.367
R414 B.n221 B.n112 163.367
R415 B.n225 B.n112 163.367
R416 B.n226 B.n225 163.367
R417 B.n227 B.n226 163.367
R418 B.n227 B.n108 163.367
R419 B.n232 B.n108 163.367
R420 B.n233 B.n232 163.367
R421 B.n234 B.n233 163.367
R422 B.n234 B.n106 163.367
R423 B.n238 B.n106 163.367
R424 B.n239 B.n238 163.367
R425 B.n240 B.n239 163.367
R426 B.n240 B.n104 163.367
R427 B.n247 B.n104 163.367
R428 B.n248 B.n247 163.367
R429 B.n249 B.n248 163.367
R430 B.n249 B.n102 163.367
R431 B.n253 B.n102 163.367
R432 B.n254 B.n253 163.367
R433 B.n255 B.n254 163.367
R434 B.n255 B.n100 163.367
R435 B.n259 B.n100 163.367
R436 B.n260 B.n259 163.367
R437 B.n261 B.n260 163.367
R438 B.n261 B.n98 163.367
R439 B.n265 B.n98 163.367
R440 B.n266 B.n265 163.367
R441 B.n267 B.n266 163.367
R442 B.n267 B.n96 163.367
R443 B.n271 B.n96 163.367
R444 B.n272 B.n271 163.367
R445 B.n273 B.n272 163.367
R446 B.n273 B.n94 163.367
R447 B.n277 B.n94 163.367
R448 B.n278 B.n277 163.367
R449 B.n279 B.n278 163.367
R450 B.n279 B.n92 163.367
R451 B.n283 B.n92 163.367
R452 B.n284 B.n283 163.367
R453 B.n285 B.n284 163.367
R454 B.n285 B.n90 163.367
R455 B.n289 B.n90 163.367
R456 B.n290 B.n289 163.367
R457 B.n291 B.n290 163.367
R458 B.n291 B.n88 163.367
R459 B.n295 B.n88 163.367
R460 B.n296 B.n295 163.367
R461 B.n297 B.n296 163.367
R462 B.n297 B.n86 163.367
R463 B.n302 B.n301 163.367
R464 B.n303 B.n302 163.367
R465 B.n303 B.n84 163.367
R466 B.n307 B.n84 163.367
R467 B.n308 B.n307 163.367
R468 B.n309 B.n308 163.367
R469 B.n309 B.n82 163.367
R470 B.n313 B.n82 163.367
R471 B.n314 B.n313 163.367
R472 B.n315 B.n314 163.367
R473 B.n315 B.n80 163.367
R474 B.n319 B.n80 163.367
R475 B.n320 B.n319 163.367
R476 B.n321 B.n320 163.367
R477 B.n321 B.n78 163.367
R478 B.n325 B.n78 163.367
R479 B.n326 B.n325 163.367
R480 B.n327 B.n326 163.367
R481 B.n327 B.n76 163.367
R482 B.n331 B.n76 163.367
R483 B.n332 B.n331 163.367
R484 B.n333 B.n332 163.367
R485 B.n333 B.n74 163.367
R486 B.n337 B.n74 163.367
R487 B.n338 B.n337 163.367
R488 B.n339 B.n338 163.367
R489 B.n339 B.n72 163.367
R490 B.n343 B.n72 163.367
R491 B.n344 B.n343 163.367
R492 B.n345 B.n344 163.367
R493 B.n345 B.n70 163.367
R494 B.n349 B.n70 163.367
R495 B.n350 B.n349 163.367
R496 B.n351 B.n350 163.367
R497 B.n351 B.n68 163.367
R498 B.n355 B.n68 163.367
R499 B.n356 B.n355 163.367
R500 B.n357 B.n356 163.367
R501 B.n357 B.n66 163.367
R502 B.n361 B.n66 163.367
R503 B.n362 B.n361 163.367
R504 B.n363 B.n362 163.367
R505 B.n363 B.n64 163.367
R506 B.n367 B.n64 163.367
R507 B.n368 B.n367 163.367
R508 B.n369 B.n368 163.367
R509 B.n369 B.n62 163.367
R510 B.n373 B.n62 163.367
R511 B.n374 B.n373 163.367
R512 B.n375 B.n374 163.367
R513 B.n375 B.n60 163.367
R514 B.n379 B.n60 163.367
R515 B.n496 B.n15 163.367
R516 B.n496 B.n495 163.367
R517 B.n495 B.n494 163.367
R518 B.n494 B.n17 163.367
R519 B.n490 B.n17 163.367
R520 B.n490 B.n489 163.367
R521 B.n489 B.n488 163.367
R522 B.n488 B.n19 163.367
R523 B.n484 B.n19 163.367
R524 B.n484 B.n483 163.367
R525 B.n483 B.n482 163.367
R526 B.n482 B.n21 163.367
R527 B.n478 B.n21 163.367
R528 B.n478 B.n477 163.367
R529 B.n477 B.n476 163.367
R530 B.n476 B.n23 163.367
R531 B.n472 B.n23 163.367
R532 B.n472 B.n471 163.367
R533 B.n471 B.n470 163.367
R534 B.n470 B.n25 163.367
R535 B.n466 B.n25 163.367
R536 B.n466 B.n465 163.367
R537 B.n465 B.n464 163.367
R538 B.n464 B.n27 163.367
R539 B.n460 B.n27 163.367
R540 B.n460 B.n459 163.367
R541 B.n459 B.n458 163.367
R542 B.n458 B.n29 163.367
R543 B.n454 B.n29 163.367
R544 B.n454 B.n453 163.367
R545 B.n453 B.n452 163.367
R546 B.n452 B.n31 163.367
R547 B.n448 B.n31 163.367
R548 B.n448 B.n447 163.367
R549 B.n447 B.n446 163.367
R550 B.n446 B.n33 163.367
R551 B.n442 B.n33 163.367
R552 B.n442 B.n441 163.367
R553 B.n441 B.n440 163.367
R554 B.n440 B.n38 163.367
R555 B.n436 B.n38 163.367
R556 B.n436 B.n435 163.367
R557 B.n435 B.n434 163.367
R558 B.n434 B.n40 163.367
R559 B.n429 B.n40 163.367
R560 B.n429 B.n428 163.367
R561 B.n428 B.n427 163.367
R562 B.n427 B.n44 163.367
R563 B.n423 B.n44 163.367
R564 B.n423 B.n422 163.367
R565 B.n422 B.n421 163.367
R566 B.n421 B.n46 163.367
R567 B.n417 B.n46 163.367
R568 B.n417 B.n416 163.367
R569 B.n416 B.n415 163.367
R570 B.n415 B.n48 163.367
R571 B.n411 B.n48 163.367
R572 B.n411 B.n410 163.367
R573 B.n410 B.n409 163.367
R574 B.n409 B.n50 163.367
R575 B.n405 B.n50 163.367
R576 B.n405 B.n404 163.367
R577 B.n404 B.n403 163.367
R578 B.n403 B.n52 163.367
R579 B.n399 B.n52 163.367
R580 B.n399 B.n398 163.367
R581 B.n398 B.n397 163.367
R582 B.n397 B.n54 163.367
R583 B.n393 B.n54 163.367
R584 B.n393 B.n392 163.367
R585 B.n392 B.n391 163.367
R586 B.n391 B.n56 163.367
R587 B.n387 B.n56 163.367
R588 B.n387 B.n386 163.367
R589 B.n386 B.n385 163.367
R590 B.n385 B.n58 163.367
R591 B.n381 B.n58 163.367
R592 B.n381 B.n380 163.367
R593 B.n243 B.t2 151.413
R594 B.n41 B.t10 151.413
R595 B.n109 B.t8 151.403
R596 B.n34 B.t4 151.403
R597 B.n244 B.t1 112.043
R598 B.n42 B.t11 112.043
R599 B.n110 B.t7 112.032
R600 B.n35 B.t5 112.032
R601 B.n245 B.n244 59.5399
R602 B.n230 B.n110 59.5399
R603 B.n36 B.n35 59.5399
R604 B.n432 B.n42 59.5399
R605 B.n244 B.n243 39.3702
R606 B.n110 B.n109 39.3702
R607 B.n35 B.n34 39.3702
R608 B.n42 B.n41 39.3702
R609 B.n499 B.n498 35.4346
R610 B.n378 B.n59 35.4346
R611 B.n300 B.n299 35.4346
R612 B.n176 B.n127 35.4346
R613 B B.n539 18.0485
R614 B.n498 B.n497 10.6151
R615 B.n497 B.n16 10.6151
R616 B.n493 B.n16 10.6151
R617 B.n493 B.n492 10.6151
R618 B.n492 B.n491 10.6151
R619 B.n491 B.n18 10.6151
R620 B.n487 B.n18 10.6151
R621 B.n487 B.n486 10.6151
R622 B.n486 B.n485 10.6151
R623 B.n485 B.n20 10.6151
R624 B.n481 B.n20 10.6151
R625 B.n481 B.n480 10.6151
R626 B.n480 B.n479 10.6151
R627 B.n479 B.n22 10.6151
R628 B.n475 B.n22 10.6151
R629 B.n475 B.n474 10.6151
R630 B.n474 B.n473 10.6151
R631 B.n473 B.n24 10.6151
R632 B.n469 B.n24 10.6151
R633 B.n469 B.n468 10.6151
R634 B.n468 B.n467 10.6151
R635 B.n467 B.n26 10.6151
R636 B.n463 B.n26 10.6151
R637 B.n463 B.n462 10.6151
R638 B.n462 B.n461 10.6151
R639 B.n461 B.n28 10.6151
R640 B.n457 B.n28 10.6151
R641 B.n457 B.n456 10.6151
R642 B.n456 B.n455 10.6151
R643 B.n455 B.n30 10.6151
R644 B.n451 B.n30 10.6151
R645 B.n451 B.n450 10.6151
R646 B.n450 B.n449 10.6151
R647 B.n449 B.n32 10.6151
R648 B.n445 B.n444 10.6151
R649 B.n444 B.n443 10.6151
R650 B.n443 B.n37 10.6151
R651 B.n439 B.n37 10.6151
R652 B.n439 B.n438 10.6151
R653 B.n438 B.n437 10.6151
R654 B.n437 B.n39 10.6151
R655 B.n433 B.n39 10.6151
R656 B.n431 B.n430 10.6151
R657 B.n430 B.n43 10.6151
R658 B.n426 B.n43 10.6151
R659 B.n426 B.n425 10.6151
R660 B.n425 B.n424 10.6151
R661 B.n424 B.n45 10.6151
R662 B.n420 B.n45 10.6151
R663 B.n420 B.n419 10.6151
R664 B.n419 B.n418 10.6151
R665 B.n418 B.n47 10.6151
R666 B.n414 B.n47 10.6151
R667 B.n414 B.n413 10.6151
R668 B.n413 B.n412 10.6151
R669 B.n412 B.n49 10.6151
R670 B.n408 B.n49 10.6151
R671 B.n408 B.n407 10.6151
R672 B.n407 B.n406 10.6151
R673 B.n406 B.n51 10.6151
R674 B.n402 B.n51 10.6151
R675 B.n402 B.n401 10.6151
R676 B.n401 B.n400 10.6151
R677 B.n400 B.n53 10.6151
R678 B.n396 B.n53 10.6151
R679 B.n396 B.n395 10.6151
R680 B.n395 B.n394 10.6151
R681 B.n394 B.n55 10.6151
R682 B.n390 B.n55 10.6151
R683 B.n390 B.n389 10.6151
R684 B.n389 B.n388 10.6151
R685 B.n388 B.n57 10.6151
R686 B.n384 B.n57 10.6151
R687 B.n384 B.n383 10.6151
R688 B.n383 B.n382 10.6151
R689 B.n382 B.n59 10.6151
R690 B.n300 B.n85 10.6151
R691 B.n304 B.n85 10.6151
R692 B.n305 B.n304 10.6151
R693 B.n306 B.n305 10.6151
R694 B.n306 B.n83 10.6151
R695 B.n310 B.n83 10.6151
R696 B.n311 B.n310 10.6151
R697 B.n312 B.n311 10.6151
R698 B.n312 B.n81 10.6151
R699 B.n316 B.n81 10.6151
R700 B.n317 B.n316 10.6151
R701 B.n318 B.n317 10.6151
R702 B.n318 B.n79 10.6151
R703 B.n322 B.n79 10.6151
R704 B.n323 B.n322 10.6151
R705 B.n324 B.n323 10.6151
R706 B.n324 B.n77 10.6151
R707 B.n328 B.n77 10.6151
R708 B.n329 B.n328 10.6151
R709 B.n330 B.n329 10.6151
R710 B.n330 B.n75 10.6151
R711 B.n334 B.n75 10.6151
R712 B.n335 B.n334 10.6151
R713 B.n336 B.n335 10.6151
R714 B.n336 B.n73 10.6151
R715 B.n340 B.n73 10.6151
R716 B.n341 B.n340 10.6151
R717 B.n342 B.n341 10.6151
R718 B.n342 B.n71 10.6151
R719 B.n346 B.n71 10.6151
R720 B.n347 B.n346 10.6151
R721 B.n348 B.n347 10.6151
R722 B.n348 B.n69 10.6151
R723 B.n352 B.n69 10.6151
R724 B.n353 B.n352 10.6151
R725 B.n354 B.n353 10.6151
R726 B.n354 B.n67 10.6151
R727 B.n358 B.n67 10.6151
R728 B.n359 B.n358 10.6151
R729 B.n360 B.n359 10.6151
R730 B.n360 B.n65 10.6151
R731 B.n364 B.n65 10.6151
R732 B.n365 B.n364 10.6151
R733 B.n366 B.n365 10.6151
R734 B.n366 B.n63 10.6151
R735 B.n370 B.n63 10.6151
R736 B.n371 B.n370 10.6151
R737 B.n372 B.n371 10.6151
R738 B.n372 B.n61 10.6151
R739 B.n376 B.n61 10.6151
R740 B.n377 B.n376 10.6151
R741 B.n378 B.n377 10.6151
R742 B.n180 B.n127 10.6151
R743 B.n181 B.n180 10.6151
R744 B.n182 B.n181 10.6151
R745 B.n182 B.n125 10.6151
R746 B.n186 B.n125 10.6151
R747 B.n187 B.n186 10.6151
R748 B.n188 B.n187 10.6151
R749 B.n188 B.n123 10.6151
R750 B.n192 B.n123 10.6151
R751 B.n193 B.n192 10.6151
R752 B.n194 B.n193 10.6151
R753 B.n194 B.n121 10.6151
R754 B.n198 B.n121 10.6151
R755 B.n199 B.n198 10.6151
R756 B.n200 B.n199 10.6151
R757 B.n200 B.n119 10.6151
R758 B.n204 B.n119 10.6151
R759 B.n205 B.n204 10.6151
R760 B.n206 B.n205 10.6151
R761 B.n206 B.n117 10.6151
R762 B.n210 B.n117 10.6151
R763 B.n211 B.n210 10.6151
R764 B.n212 B.n211 10.6151
R765 B.n212 B.n115 10.6151
R766 B.n216 B.n115 10.6151
R767 B.n217 B.n216 10.6151
R768 B.n218 B.n217 10.6151
R769 B.n218 B.n113 10.6151
R770 B.n222 B.n113 10.6151
R771 B.n223 B.n222 10.6151
R772 B.n224 B.n223 10.6151
R773 B.n224 B.n111 10.6151
R774 B.n228 B.n111 10.6151
R775 B.n229 B.n228 10.6151
R776 B.n231 B.n107 10.6151
R777 B.n235 B.n107 10.6151
R778 B.n236 B.n235 10.6151
R779 B.n237 B.n236 10.6151
R780 B.n237 B.n105 10.6151
R781 B.n241 B.n105 10.6151
R782 B.n242 B.n241 10.6151
R783 B.n246 B.n242 10.6151
R784 B.n250 B.n103 10.6151
R785 B.n251 B.n250 10.6151
R786 B.n252 B.n251 10.6151
R787 B.n252 B.n101 10.6151
R788 B.n256 B.n101 10.6151
R789 B.n257 B.n256 10.6151
R790 B.n258 B.n257 10.6151
R791 B.n258 B.n99 10.6151
R792 B.n262 B.n99 10.6151
R793 B.n263 B.n262 10.6151
R794 B.n264 B.n263 10.6151
R795 B.n264 B.n97 10.6151
R796 B.n268 B.n97 10.6151
R797 B.n269 B.n268 10.6151
R798 B.n270 B.n269 10.6151
R799 B.n270 B.n95 10.6151
R800 B.n274 B.n95 10.6151
R801 B.n275 B.n274 10.6151
R802 B.n276 B.n275 10.6151
R803 B.n276 B.n93 10.6151
R804 B.n280 B.n93 10.6151
R805 B.n281 B.n280 10.6151
R806 B.n282 B.n281 10.6151
R807 B.n282 B.n91 10.6151
R808 B.n286 B.n91 10.6151
R809 B.n287 B.n286 10.6151
R810 B.n288 B.n287 10.6151
R811 B.n288 B.n89 10.6151
R812 B.n292 B.n89 10.6151
R813 B.n293 B.n292 10.6151
R814 B.n294 B.n293 10.6151
R815 B.n294 B.n87 10.6151
R816 B.n298 B.n87 10.6151
R817 B.n299 B.n298 10.6151
R818 B.n176 B.n175 10.6151
R819 B.n175 B.n174 10.6151
R820 B.n174 B.n129 10.6151
R821 B.n170 B.n129 10.6151
R822 B.n170 B.n169 10.6151
R823 B.n169 B.n168 10.6151
R824 B.n168 B.n131 10.6151
R825 B.n164 B.n131 10.6151
R826 B.n164 B.n163 10.6151
R827 B.n163 B.n162 10.6151
R828 B.n162 B.n133 10.6151
R829 B.n158 B.n133 10.6151
R830 B.n158 B.n157 10.6151
R831 B.n157 B.n156 10.6151
R832 B.n156 B.n135 10.6151
R833 B.n152 B.n135 10.6151
R834 B.n152 B.n151 10.6151
R835 B.n151 B.n150 10.6151
R836 B.n150 B.n137 10.6151
R837 B.n146 B.n137 10.6151
R838 B.n146 B.n145 10.6151
R839 B.n145 B.n144 10.6151
R840 B.n144 B.n139 10.6151
R841 B.n140 B.n139 10.6151
R842 B.n140 B.n0 10.6151
R843 B.n535 B.n1 10.6151
R844 B.n535 B.n534 10.6151
R845 B.n534 B.n533 10.6151
R846 B.n533 B.n4 10.6151
R847 B.n529 B.n4 10.6151
R848 B.n529 B.n528 10.6151
R849 B.n528 B.n527 10.6151
R850 B.n527 B.n6 10.6151
R851 B.n523 B.n6 10.6151
R852 B.n523 B.n522 10.6151
R853 B.n522 B.n521 10.6151
R854 B.n521 B.n8 10.6151
R855 B.n517 B.n8 10.6151
R856 B.n517 B.n516 10.6151
R857 B.n516 B.n515 10.6151
R858 B.n515 B.n10 10.6151
R859 B.n511 B.n10 10.6151
R860 B.n511 B.n510 10.6151
R861 B.n510 B.n509 10.6151
R862 B.n509 B.n12 10.6151
R863 B.n505 B.n12 10.6151
R864 B.n505 B.n504 10.6151
R865 B.n504 B.n503 10.6151
R866 B.n503 B.n14 10.6151
R867 B.n499 B.n14 10.6151
R868 B.n445 B.n36 6.5566
R869 B.n433 B.n432 6.5566
R870 B.n231 B.n230 6.5566
R871 B.n246 B.n245 6.5566
R872 B.n36 B.n32 4.05904
R873 B.n432 B.n431 4.05904
R874 B.n230 B.n229 4.05904
R875 B.n245 B.n103 4.05904
R876 B.n539 B.n0 2.81026
R877 B.n539 B.n1 2.81026
C0 VDD1 w_n2188_n2916# 1.2129f
C1 VTAIL VDD2 4.85031f
C2 VDD1 B 1.04271f
C3 VDD2 VN 3.57594f
C4 VDD2 VP 0.336523f
C5 VTAIL VN 3.44807f
C6 VDD2 w_n2188_n2916# 1.24888f
C7 VTAIL VP 3.46217f
C8 VTAIL w_n2188_n2916# 3.45317f
C9 B VDD2 1.08015f
C10 VP VN 5.12994f
C11 VTAIL B 3.79834f
C12 w_n2188_n2916# VN 3.51049f
C13 VDD1 VDD2 0.806964f
C14 w_n2188_n2916# VP 3.78949f
C15 VDD1 VTAIL 4.80214f
C16 B VN 0.908376f
C17 B VP 1.36718f
C18 B w_n2188_n2916# 7.5045f
C19 VDD1 VN 0.147673f
C20 VDD1 VP 3.76428f
C21 VDD2 VSUBS 0.753813f
C22 VDD1 VSUBS 4.948347f
C23 VTAIL VSUBS 0.969721f
C24 VN VSUBS 5.0335f
C25 VP VSUBS 1.710596f
C26 B VSUBS 3.306152f
C27 w_n2188_n2916# VSUBS 78.846794f
C28 B.n0 VSUBS 0.004847f
C29 B.n1 VSUBS 0.004847f
C30 B.n2 VSUBS 0.007666f
C31 B.n3 VSUBS 0.007666f
C32 B.n4 VSUBS 0.007666f
C33 B.n5 VSUBS 0.007666f
C34 B.n6 VSUBS 0.007666f
C35 B.n7 VSUBS 0.007666f
C36 B.n8 VSUBS 0.007666f
C37 B.n9 VSUBS 0.007666f
C38 B.n10 VSUBS 0.007666f
C39 B.n11 VSUBS 0.007666f
C40 B.n12 VSUBS 0.007666f
C41 B.n13 VSUBS 0.007666f
C42 B.n14 VSUBS 0.007666f
C43 B.n15 VSUBS 0.019173f
C44 B.n16 VSUBS 0.007666f
C45 B.n17 VSUBS 0.007666f
C46 B.n18 VSUBS 0.007666f
C47 B.n19 VSUBS 0.007666f
C48 B.n20 VSUBS 0.007666f
C49 B.n21 VSUBS 0.007666f
C50 B.n22 VSUBS 0.007666f
C51 B.n23 VSUBS 0.007666f
C52 B.n24 VSUBS 0.007666f
C53 B.n25 VSUBS 0.007666f
C54 B.n26 VSUBS 0.007666f
C55 B.n27 VSUBS 0.007666f
C56 B.n28 VSUBS 0.007666f
C57 B.n29 VSUBS 0.007666f
C58 B.n30 VSUBS 0.007666f
C59 B.n31 VSUBS 0.007666f
C60 B.n32 VSUBS 0.005298f
C61 B.n33 VSUBS 0.007666f
C62 B.t5 VSUBS 0.338976f
C63 B.t4 VSUBS 0.355465f
C64 B.t3 VSUBS 0.812263f
C65 B.n34 VSUBS 0.169612f
C66 B.n35 VSUBS 0.074342f
C67 B.n36 VSUBS 0.017761f
C68 B.n37 VSUBS 0.007666f
C69 B.n38 VSUBS 0.007666f
C70 B.n39 VSUBS 0.007666f
C71 B.n40 VSUBS 0.007666f
C72 B.t11 VSUBS 0.338972f
C73 B.t10 VSUBS 0.35546f
C74 B.t9 VSUBS 0.812263f
C75 B.n41 VSUBS 0.169616f
C76 B.n42 VSUBS 0.074346f
C77 B.n43 VSUBS 0.007666f
C78 B.n44 VSUBS 0.007666f
C79 B.n45 VSUBS 0.007666f
C80 B.n46 VSUBS 0.007666f
C81 B.n47 VSUBS 0.007666f
C82 B.n48 VSUBS 0.007666f
C83 B.n49 VSUBS 0.007666f
C84 B.n50 VSUBS 0.007666f
C85 B.n51 VSUBS 0.007666f
C86 B.n52 VSUBS 0.007666f
C87 B.n53 VSUBS 0.007666f
C88 B.n54 VSUBS 0.007666f
C89 B.n55 VSUBS 0.007666f
C90 B.n56 VSUBS 0.007666f
C91 B.n57 VSUBS 0.007666f
C92 B.n58 VSUBS 0.007666f
C93 B.n59 VSUBS 0.018338f
C94 B.n60 VSUBS 0.007666f
C95 B.n61 VSUBS 0.007666f
C96 B.n62 VSUBS 0.007666f
C97 B.n63 VSUBS 0.007666f
C98 B.n64 VSUBS 0.007666f
C99 B.n65 VSUBS 0.007666f
C100 B.n66 VSUBS 0.007666f
C101 B.n67 VSUBS 0.007666f
C102 B.n68 VSUBS 0.007666f
C103 B.n69 VSUBS 0.007666f
C104 B.n70 VSUBS 0.007666f
C105 B.n71 VSUBS 0.007666f
C106 B.n72 VSUBS 0.007666f
C107 B.n73 VSUBS 0.007666f
C108 B.n74 VSUBS 0.007666f
C109 B.n75 VSUBS 0.007666f
C110 B.n76 VSUBS 0.007666f
C111 B.n77 VSUBS 0.007666f
C112 B.n78 VSUBS 0.007666f
C113 B.n79 VSUBS 0.007666f
C114 B.n80 VSUBS 0.007666f
C115 B.n81 VSUBS 0.007666f
C116 B.n82 VSUBS 0.007666f
C117 B.n83 VSUBS 0.007666f
C118 B.n84 VSUBS 0.007666f
C119 B.n85 VSUBS 0.007666f
C120 B.n86 VSUBS 0.019173f
C121 B.n87 VSUBS 0.007666f
C122 B.n88 VSUBS 0.007666f
C123 B.n89 VSUBS 0.007666f
C124 B.n90 VSUBS 0.007666f
C125 B.n91 VSUBS 0.007666f
C126 B.n92 VSUBS 0.007666f
C127 B.n93 VSUBS 0.007666f
C128 B.n94 VSUBS 0.007666f
C129 B.n95 VSUBS 0.007666f
C130 B.n96 VSUBS 0.007666f
C131 B.n97 VSUBS 0.007666f
C132 B.n98 VSUBS 0.007666f
C133 B.n99 VSUBS 0.007666f
C134 B.n100 VSUBS 0.007666f
C135 B.n101 VSUBS 0.007666f
C136 B.n102 VSUBS 0.007666f
C137 B.n103 VSUBS 0.005298f
C138 B.n104 VSUBS 0.007666f
C139 B.n105 VSUBS 0.007666f
C140 B.n106 VSUBS 0.007666f
C141 B.n107 VSUBS 0.007666f
C142 B.n108 VSUBS 0.007666f
C143 B.t7 VSUBS 0.338976f
C144 B.t8 VSUBS 0.355465f
C145 B.t6 VSUBS 0.812263f
C146 B.n109 VSUBS 0.169612f
C147 B.n110 VSUBS 0.074342f
C148 B.n111 VSUBS 0.007666f
C149 B.n112 VSUBS 0.007666f
C150 B.n113 VSUBS 0.007666f
C151 B.n114 VSUBS 0.007666f
C152 B.n115 VSUBS 0.007666f
C153 B.n116 VSUBS 0.007666f
C154 B.n117 VSUBS 0.007666f
C155 B.n118 VSUBS 0.007666f
C156 B.n119 VSUBS 0.007666f
C157 B.n120 VSUBS 0.007666f
C158 B.n121 VSUBS 0.007666f
C159 B.n122 VSUBS 0.007666f
C160 B.n123 VSUBS 0.007666f
C161 B.n124 VSUBS 0.007666f
C162 B.n125 VSUBS 0.007666f
C163 B.n126 VSUBS 0.007666f
C164 B.n127 VSUBS 0.019173f
C165 B.n128 VSUBS 0.007666f
C166 B.n129 VSUBS 0.007666f
C167 B.n130 VSUBS 0.007666f
C168 B.n131 VSUBS 0.007666f
C169 B.n132 VSUBS 0.007666f
C170 B.n133 VSUBS 0.007666f
C171 B.n134 VSUBS 0.007666f
C172 B.n135 VSUBS 0.007666f
C173 B.n136 VSUBS 0.007666f
C174 B.n137 VSUBS 0.007666f
C175 B.n138 VSUBS 0.007666f
C176 B.n139 VSUBS 0.007666f
C177 B.n140 VSUBS 0.007666f
C178 B.n141 VSUBS 0.007666f
C179 B.n142 VSUBS 0.007666f
C180 B.n143 VSUBS 0.007666f
C181 B.n144 VSUBS 0.007666f
C182 B.n145 VSUBS 0.007666f
C183 B.n146 VSUBS 0.007666f
C184 B.n147 VSUBS 0.007666f
C185 B.n148 VSUBS 0.007666f
C186 B.n149 VSUBS 0.007666f
C187 B.n150 VSUBS 0.007666f
C188 B.n151 VSUBS 0.007666f
C189 B.n152 VSUBS 0.007666f
C190 B.n153 VSUBS 0.007666f
C191 B.n154 VSUBS 0.007666f
C192 B.n155 VSUBS 0.007666f
C193 B.n156 VSUBS 0.007666f
C194 B.n157 VSUBS 0.007666f
C195 B.n158 VSUBS 0.007666f
C196 B.n159 VSUBS 0.007666f
C197 B.n160 VSUBS 0.007666f
C198 B.n161 VSUBS 0.007666f
C199 B.n162 VSUBS 0.007666f
C200 B.n163 VSUBS 0.007666f
C201 B.n164 VSUBS 0.007666f
C202 B.n165 VSUBS 0.007666f
C203 B.n166 VSUBS 0.007666f
C204 B.n167 VSUBS 0.007666f
C205 B.n168 VSUBS 0.007666f
C206 B.n169 VSUBS 0.007666f
C207 B.n170 VSUBS 0.007666f
C208 B.n171 VSUBS 0.007666f
C209 B.n172 VSUBS 0.007666f
C210 B.n173 VSUBS 0.007666f
C211 B.n174 VSUBS 0.007666f
C212 B.n175 VSUBS 0.007666f
C213 B.n176 VSUBS 0.018705f
C214 B.n177 VSUBS 0.018705f
C215 B.n178 VSUBS 0.019173f
C216 B.n179 VSUBS 0.007666f
C217 B.n180 VSUBS 0.007666f
C218 B.n181 VSUBS 0.007666f
C219 B.n182 VSUBS 0.007666f
C220 B.n183 VSUBS 0.007666f
C221 B.n184 VSUBS 0.007666f
C222 B.n185 VSUBS 0.007666f
C223 B.n186 VSUBS 0.007666f
C224 B.n187 VSUBS 0.007666f
C225 B.n188 VSUBS 0.007666f
C226 B.n189 VSUBS 0.007666f
C227 B.n190 VSUBS 0.007666f
C228 B.n191 VSUBS 0.007666f
C229 B.n192 VSUBS 0.007666f
C230 B.n193 VSUBS 0.007666f
C231 B.n194 VSUBS 0.007666f
C232 B.n195 VSUBS 0.007666f
C233 B.n196 VSUBS 0.007666f
C234 B.n197 VSUBS 0.007666f
C235 B.n198 VSUBS 0.007666f
C236 B.n199 VSUBS 0.007666f
C237 B.n200 VSUBS 0.007666f
C238 B.n201 VSUBS 0.007666f
C239 B.n202 VSUBS 0.007666f
C240 B.n203 VSUBS 0.007666f
C241 B.n204 VSUBS 0.007666f
C242 B.n205 VSUBS 0.007666f
C243 B.n206 VSUBS 0.007666f
C244 B.n207 VSUBS 0.007666f
C245 B.n208 VSUBS 0.007666f
C246 B.n209 VSUBS 0.007666f
C247 B.n210 VSUBS 0.007666f
C248 B.n211 VSUBS 0.007666f
C249 B.n212 VSUBS 0.007666f
C250 B.n213 VSUBS 0.007666f
C251 B.n214 VSUBS 0.007666f
C252 B.n215 VSUBS 0.007666f
C253 B.n216 VSUBS 0.007666f
C254 B.n217 VSUBS 0.007666f
C255 B.n218 VSUBS 0.007666f
C256 B.n219 VSUBS 0.007666f
C257 B.n220 VSUBS 0.007666f
C258 B.n221 VSUBS 0.007666f
C259 B.n222 VSUBS 0.007666f
C260 B.n223 VSUBS 0.007666f
C261 B.n224 VSUBS 0.007666f
C262 B.n225 VSUBS 0.007666f
C263 B.n226 VSUBS 0.007666f
C264 B.n227 VSUBS 0.007666f
C265 B.n228 VSUBS 0.007666f
C266 B.n229 VSUBS 0.005298f
C267 B.n230 VSUBS 0.017761f
C268 B.n231 VSUBS 0.0062f
C269 B.n232 VSUBS 0.007666f
C270 B.n233 VSUBS 0.007666f
C271 B.n234 VSUBS 0.007666f
C272 B.n235 VSUBS 0.007666f
C273 B.n236 VSUBS 0.007666f
C274 B.n237 VSUBS 0.007666f
C275 B.n238 VSUBS 0.007666f
C276 B.n239 VSUBS 0.007666f
C277 B.n240 VSUBS 0.007666f
C278 B.n241 VSUBS 0.007666f
C279 B.n242 VSUBS 0.007666f
C280 B.t1 VSUBS 0.338972f
C281 B.t2 VSUBS 0.35546f
C282 B.t0 VSUBS 0.812263f
C283 B.n243 VSUBS 0.169616f
C284 B.n244 VSUBS 0.074346f
C285 B.n245 VSUBS 0.017761f
C286 B.n246 VSUBS 0.0062f
C287 B.n247 VSUBS 0.007666f
C288 B.n248 VSUBS 0.007666f
C289 B.n249 VSUBS 0.007666f
C290 B.n250 VSUBS 0.007666f
C291 B.n251 VSUBS 0.007666f
C292 B.n252 VSUBS 0.007666f
C293 B.n253 VSUBS 0.007666f
C294 B.n254 VSUBS 0.007666f
C295 B.n255 VSUBS 0.007666f
C296 B.n256 VSUBS 0.007666f
C297 B.n257 VSUBS 0.007666f
C298 B.n258 VSUBS 0.007666f
C299 B.n259 VSUBS 0.007666f
C300 B.n260 VSUBS 0.007666f
C301 B.n261 VSUBS 0.007666f
C302 B.n262 VSUBS 0.007666f
C303 B.n263 VSUBS 0.007666f
C304 B.n264 VSUBS 0.007666f
C305 B.n265 VSUBS 0.007666f
C306 B.n266 VSUBS 0.007666f
C307 B.n267 VSUBS 0.007666f
C308 B.n268 VSUBS 0.007666f
C309 B.n269 VSUBS 0.007666f
C310 B.n270 VSUBS 0.007666f
C311 B.n271 VSUBS 0.007666f
C312 B.n272 VSUBS 0.007666f
C313 B.n273 VSUBS 0.007666f
C314 B.n274 VSUBS 0.007666f
C315 B.n275 VSUBS 0.007666f
C316 B.n276 VSUBS 0.007666f
C317 B.n277 VSUBS 0.007666f
C318 B.n278 VSUBS 0.007666f
C319 B.n279 VSUBS 0.007666f
C320 B.n280 VSUBS 0.007666f
C321 B.n281 VSUBS 0.007666f
C322 B.n282 VSUBS 0.007666f
C323 B.n283 VSUBS 0.007666f
C324 B.n284 VSUBS 0.007666f
C325 B.n285 VSUBS 0.007666f
C326 B.n286 VSUBS 0.007666f
C327 B.n287 VSUBS 0.007666f
C328 B.n288 VSUBS 0.007666f
C329 B.n289 VSUBS 0.007666f
C330 B.n290 VSUBS 0.007666f
C331 B.n291 VSUBS 0.007666f
C332 B.n292 VSUBS 0.007666f
C333 B.n293 VSUBS 0.007666f
C334 B.n294 VSUBS 0.007666f
C335 B.n295 VSUBS 0.007666f
C336 B.n296 VSUBS 0.007666f
C337 B.n297 VSUBS 0.007666f
C338 B.n298 VSUBS 0.007666f
C339 B.n299 VSUBS 0.019173f
C340 B.n300 VSUBS 0.018705f
C341 B.n301 VSUBS 0.018705f
C342 B.n302 VSUBS 0.007666f
C343 B.n303 VSUBS 0.007666f
C344 B.n304 VSUBS 0.007666f
C345 B.n305 VSUBS 0.007666f
C346 B.n306 VSUBS 0.007666f
C347 B.n307 VSUBS 0.007666f
C348 B.n308 VSUBS 0.007666f
C349 B.n309 VSUBS 0.007666f
C350 B.n310 VSUBS 0.007666f
C351 B.n311 VSUBS 0.007666f
C352 B.n312 VSUBS 0.007666f
C353 B.n313 VSUBS 0.007666f
C354 B.n314 VSUBS 0.007666f
C355 B.n315 VSUBS 0.007666f
C356 B.n316 VSUBS 0.007666f
C357 B.n317 VSUBS 0.007666f
C358 B.n318 VSUBS 0.007666f
C359 B.n319 VSUBS 0.007666f
C360 B.n320 VSUBS 0.007666f
C361 B.n321 VSUBS 0.007666f
C362 B.n322 VSUBS 0.007666f
C363 B.n323 VSUBS 0.007666f
C364 B.n324 VSUBS 0.007666f
C365 B.n325 VSUBS 0.007666f
C366 B.n326 VSUBS 0.007666f
C367 B.n327 VSUBS 0.007666f
C368 B.n328 VSUBS 0.007666f
C369 B.n329 VSUBS 0.007666f
C370 B.n330 VSUBS 0.007666f
C371 B.n331 VSUBS 0.007666f
C372 B.n332 VSUBS 0.007666f
C373 B.n333 VSUBS 0.007666f
C374 B.n334 VSUBS 0.007666f
C375 B.n335 VSUBS 0.007666f
C376 B.n336 VSUBS 0.007666f
C377 B.n337 VSUBS 0.007666f
C378 B.n338 VSUBS 0.007666f
C379 B.n339 VSUBS 0.007666f
C380 B.n340 VSUBS 0.007666f
C381 B.n341 VSUBS 0.007666f
C382 B.n342 VSUBS 0.007666f
C383 B.n343 VSUBS 0.007666f
C384 B.n344 VSUBS 0.007666f
C385 B.n345 VSUBS 0.007666f
C386 B.n346 VSUBS 0.007666f
C387 B.n347 VSUBS 0.007666f
C388 B.n348 VSUBS 0.007666f
C389 B.n349 VSUBS 0.007666f
C390 B.n350 VSUBS 0.007666f
C391 B.n351 VSUBS 0.007666f
C392 B.n352 VSUBS 0.007666f
C393 B.n353 VSUBS 0.007666f
C394 B.n354 VSUBS 0.007666f
C395 B.n355 VSUBS 0.007666f
C396 B.n356 VSUBS 0.007666f
C397 B.n357 VSUBS 0.007666f
C398 B.n358 VSUBS 0.007666f
C399 B.n359 VSUBS 0.007666f
C400 B.n360 VSUBS 0.007666f
C401 B.n361 VSUBS 0.007666f
C402 B.n362 VSUBS 0.007666f
C403 B.n363 VSUBS 0.007666f
C404 B.n364 VSUBS 0.007666f
C405 B.n365 VSUBS 0.007666f
C406 B.n366 VSUBS 0.007666f
C407 B.n367 VSUBS 0.007666f
C408 B.n368 VSUBS 0.007666f
C409 B.n369 VSUBS 0.007666f
C410 B.n370 VSUBS 0.007666f
C411 B.n371 VSUBS 0.007666f
C412 B.n372 VSUBS 0.007666f
C413 B.n373 VSUBS 0.007666f
C414 B.n374 VSUBS 0.007666f
C415 B.n375 VSUBS 0.007666f
C416 B.n376 VSUBS 0.007666f
C417 B.n377 VSUBS 0.007666f
C418 B.n378 VSUBS 0.01954f
C419 B.n379 VSUBS 0.018705f
C420 B.n380 VSUBS 0.019173f
C421 B.n381 VSUBS 0.007666f
C422 B.n382 VSUBS 0.007666f
C423 B.n383 VSUBS 0.007666f
C424 B.n384 VSUBS 0.007666f
C425 B.n385 VSUBS 0.007666f
C426 B.n386 VSUBS 0.007666f
C427 B.n387 VSUBS 0.007666f
C428 B.n388 VSUBS 0.007666f
C429 B.n389 VSUBS 0.007666f
C430 B.n390 VSUBS 0.007666f
C431 B.n391 VSUBS 0.007666f
C432 B.n392 VSUBS 0.007666f
C433 B.n393 VSUBS 0.007666f
C434 B.n394 VSUBS 0.007666f
C435 B.n395 VSUBS 0.007666f
C436 B.n396 VSUBS 0.007666f
C437 B.n397 VSUBS 0.007666f
C438 B.n398 VSUBS 0.007666f
C439 B.n399 VSUBS 0.007666f
C440 B.n400 VSUBS 0.007666f
C441 B.n401 VSUBS 0.007666f
C442 B.n402 VSUBS 0.007666f
C443 B.n403 VSUBS 0.007666f
C444 B.n404 VSUBS 0.007666f
C445 B.n405 VSUBS 0.007666f
C446 B.n406 VSUBS 0.007666f
C447 B.n407 VSUBS 0.007666f
C448 B.n408 VSUBS 0.007666f
C449 B.n409 VSUBS 0.007666f
C450 B.n410 VSUBS 0.007666f
C451 B.n411 VSUBS 0.007666f
C452 B.n412 VSUBS 0.007666f
C453 B.n413 VSUBS 0.007666f
C454 B.n414 VSUBS 0.007666f
C455 B.n415 VSUBS 0.007666f
C456 B.n416 VSUBS 0.007666f
C457 B.n417 VSUBS 0.007666f
C458 B.n418 VSUBS 0.007666f
C459 B.n419 VSUBS 0.007666f
C460 B.n420 VSUBS 0.007666f
C461 B.n421 VSUBS 0.007666f
C462 B.n422 VSUBS 0.007666f
C463 B.n423 VSUBS 0.007666f
C464 B.n424 VSUBS 0.007666f
C465 B.n425 VSUBS 0.007666f
C466 B.n426 VSUBS 0.007666f
C467 B.n427 VSUBS 0.007666f
C468 B.n428 VSUBS 0.007666f
C469 B.n429 VSUBS 0.007666f
C470 B.n430 VSUBS 0.007666f
C471 B.n431 VSUBS 0.005298f
C472 B.n432 VSUBS 0.017761f
C473 B.n433 VSUBS 0.0062f
C474 B.n434 VSUBS 0.007666f
C475 B.n435 VSUBS 0.007666f
C476 B.n436 VSUBS 0.007666f
C477 B.n437 VSUBS 0.007666f
C478 B.n438 VSUBS 0.007666f
C479 B.n439 VSUBS 0.007666f
C480 B.n440 VSUBS 0.007666f
C481 B.n441 VSUBS 0.007666f
C482 B.n442 VSUBS 0.007666f
C483 B.n443 VSUBS 0.007666f
C484 B.n444 VSUBS 0.007666f
C485 B.n445 VSUBS 0.0062f
C486 B.n446 VSUBS 0.007666f
C487 B.n447 VSUBS 0.007666f
C488 B.n448 VSUBS 0.007666f
C489 B.n449 VSUBS 0.007666f
C490 B.n450 VSUBS 0.007666f
C491 B.n451 VSUBS 0.007666f
C492 B.n452 VSUBS 0.007666f
C493 B.n453 VSUBS 0.007666f
C494 B.n454 VSUBS 0.007666f
C495 B.n455 VSUBS 0.007666f
C496 B.n456 VSUBS 0.007666f
C497 B.n457 VSUBS 0.007666f
C498 B.n458 VSUBS 0.007666f
C499 B.n459 VSUBS 0.007666f
C500 B.n460 VSUBS 0.007666f
C501 B.n461 VSUBS 0.007666f
C502 B.n462 VSUBS 0.007666f
C503 B.n463 VSUBS 0.007666f
C504 B.n464 VSUBS 0.007666f
C505 B.n465 VSUBS 0.007666f
C506 B.n466 VSUBS 0.007666f
C507 B.n467 VSUBS 0.007666f
C508 B.n468 VSUBS 0.007666f
C509 B.n469 VSUBS 0.007666f
C510 B.n470 VSUBS 0.007666f
C511 B.n471 VSUBS 0.007666f
C512 B.n472 VSUBS 0.007666f
C513 B.n473 VSUBS 0.007666f
C514 B.n474 VSUBS 0.007666f
C515 B.n475 VSUBS 0.007666f
C516 B.n476 VSUBS 0.007666f
C517 B.n477 VSUBS 0.007666f
C518 B.n478 VSUBS 0.007666f
C519 B.n479 VSUBS 0.007666f
C520 B.n480 VSUBS 0.007666f
C521 B.n481 VSUBS 0.007666f
C522 B.n482 VSUBS 0.007666f
C523 B.n483 VSUBS 0.007666f
C524 B.n484 VSUBS 0.007666f
C525 B.n485 VSUBS 0.007666f
C526 B.n486 VSUBS 0.007666f
C527 B.n487 VSUBS 0.007666f
C528 B.n488 VSUBS 0.007666f
C529 B.n489 VSUBS 0.007666f
C530 B.n490 VSUBS 0.007666f
C531 B.n491 VSUBS 0.007666f
C532 B.n492 VSUBS 0.007666f
C533 B.n493 VSUBS 0.007666f
C534 B.n494 VSUBS 0.007666f
C535 B.n495 VSUBS 0.007666f
C536 B.n496 VSUBS 0.007666f
C537 B.n497 VSUBS 0.007666f
C538 B.n498 VSUBS 0.019173f
C539 B.n499 VSUBS 0.018705f
C540 B.n500 VSUBS 0.018705f
C541 B.n501 VSUBS 0.007666f
C542 B.n502 VSUBS 0.007666f
C543 B.n503 VSUBS 0.007666f
C544 B.n504 VSUBS 0.007666f
C545 B.n505 VSUBS 0.007666f
C546 B.n506 VSUBS 0.007666f
C547 B.n507 VSUBS 0.007666f
C548 B.n508 VSUBS 0.007666f
C549 B.n509 VSUBS 0.007666f
C550 B.n510 VSUBS 0.007666f
C551 B.n511 VSUBS 0.007666f
C552 B.n512 VSUBS 0.007666f
C553 B.n513 VSUBS 0.007666f
C554 B.n514 VSUBS 0.007666f
C555 B.n515 VSUBS 0.007666f
C556 B.n516 VSUBS 0.007666f
C557 B.n517 VSUBS 0.007666f
C558 B.n518 VSUBS 0.007666f
C559 B.n519 VSUBS 0.007666f
C560 B.n520 VSUBS 0.007666f
C561 B.n521 VSUBS 0.007666f
C562 B.n522 VSUBS 0.007666f
C563 B.n523 VSUBS 0.007666f
C564 B.n524 VSUBS 0.007666f
C565 B.n525 VSUBS 0.007666f
C566 B.n526 VSUBS 0.007666f
C567 B.n527 VSUBS 0.007666f
C568 B.n528 VSUBS 0.007666f
C569 B.n529 VSUBS 0.007666f
C570 B.n530 VSUBS 0.007666f
C571 B.n531 VSUBS 0.007666f
C572 B.n532 VSUBS 0.007666f
C573 B.n533 VSUBS 0.007666f
C574 B.n534 VSUBS 0.007666f
C575 B.n535 VSUBS 0.007666f
C576 B.n536 VSUBS 0.007666f
C577 B.n537 VSUBS 0.007666f
C578 B.n538 VSUBS 0.007666f
C579 B.n539 VSUBS 0.017358f
C580 VDD2.t0 VSUBS 0.208147f
C581 VDD2.t1 VSUBS 0.208147f
C582 VDD2.n0 VSUBS 2.12008f
C583 VDD2.t3 VSUBS 0.208147f
C584 VDD2.t2 VSUBS 0.208147f
C585 VDD2.n1 VSUBS 1.57156f
C586 VDD2.n2 VSUBS 3.81745f
C587 VN.t3 VSUBS 2.10498f
C588 VN.t2 VSUBS 2.10274f
C589 VN.n0 VSUBS 1.51373f
C590 VN.t1 VSUBS 2.10498f
C591 VN.t0 VSUBS 2.10274f
C592 VN.n1 VSUBS 3.1917f
C593 VDD1.t2 VSUBS 0.20815f
C594 VDD1.t3 VSUBS 0.20815f
C595 VDD1.n0 VSUBS 1.57205f
C596 VDD1.t1 VSUBS 0.20815f
C597 VDD1.t0 VSUBS 0.20815f
C598 VDD1.n1 VSUBS 2.14279f
C599 VTAIL.t2 VSUBS 1.70285f
C600 VTAIL.n0 VSUBS 0.686562f
C601 VTAIL.t4 VSUBS 1.70285f
C602 VTAIL.n1 VSUBS 0.749492f
C603 VTAIL.t7 VSUBS 1.70285f
C604 VTAIL.n2 VSUBS 1.8198f
C605 VTAIL.t3 VSUBS 1.70286f
C606 VTAIL.n3 VSUBS 1.81979f
C607 VTAIL.t0 VSUBS 1.70286f
C608 VTAIL.n4 VSUBS 0.74948f
C609 VTAIL.t6 VSUBS 1.70286f
C610 VTAIL.n5 VSUBS 0.74948f
C611 VTAIL.t5 VSUBS 1.70285f
C612 VTAIL.n6 VSUBS 1.8198f
C613 VTAIL.t1 VSUBS 1.70285f
C614 VTAIL.n7 VSUBS 1.74791f
C615 VP.n0 VSUBS 0.044722f
C616 VP.t3 VSUBS 2.00423f
C617 VP.n1 VSUBS 0.03619f
C618 VP.n2 VSUBS 0.044722f
C619 VP.t2 VSUBS 2.00423f
C620 VP.t1 VSUBS 2.19442f
C621 VP.t0 VSUBS 2.19209f
C622 VP.n3 VSUBS 3.30047f
C623 VP.n4 VSUBS 2.2713f
C624 VP.n5 VSUBS 0.821697f
C625 VP.n6 VSUBS 0.04365f
C626 VP.n7 VSUBS 0.08936f
C627 VP.n8 VSUBS 0.044722f
C628 VP.n9 VSUBS 0.044722f
C629 VP.n10 VSUBS 0.044722f
C630 VP.n11 VSUBS 0.08936f
C631 VP.n12 VSUBS 0.04365f
C632 VP.n13 VSUBS 0.821697f
C633 VP.n14 VSUBS 0.047626f
.ends

