* NGSPICE file created from diff_pair_sample_0610.ext - technology: sky130A

.subckt diff_pair_sample_0610 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=0 ps=0 w=18.21 l=1.53
X1 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=0 ps=0 w=18.21 l=1.53
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=0 ps=0 w=18.21 l=1.53
X3 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=0 ps=0 w=18.21 l=1.53
X4 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=7.1019 ps=37.2 w=18.21 l=1.53
X5 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=7.1019 ps=37.2 w=18.21 l=1.53
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=7.1019 ps=37.2 w=18.21 l=1.53
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.1019 pd=37.2 as=7.1019 ps=37.2 w=18.21 l=1.53
R0 B.n808 B.n807 585
R1 B.n809 B.n808 585
R2 B.n361 B.n103 585
R3 B.n360 B.n359 585
R4 B.n358 B.n357 585
R5 B.n356 B.n355 585
R6 B.n354 B.n353 585
R7 B.n352 B.n351 585
R8 B.n350 B.n349 585
R9 B.n348 B.n347 585
R10 B.n346 B.n345 585
R11 B.n344 B.n343 585
R12 B.n342 B.n341 585
R13 B.n340 B.n339 585
R14 B.n338 B.n337 585
R15 B.n336 B.n335 585
R16 B.n334 B.n333 585
R17 B.n332 B.n331 585
R18 B.n330 B.n329 585
R19 B.n328 B.n327 585
R20 B.n326 B.n325 585
R21 B.n324 B.n323 585
R22 B.n322 B.n321 585
R23 B.n320 B.n319 585
R24 B.n318 B.n317 585
R25 B.n316 B.n315 585
R26 B.n314 B.n313 585
R27 B.n312 B.n311 585
R28 B.n310 B.n309 585
R29 B.n308 B.n307 585
R30 B.n306 B.n305 585
R31 B.n304 B.n303 585
R32 B.n302 B.n301 585
R33 B.n300 B.n299 585
R34 B.n298 B.n297 585
R35 B.n296 B.n295 585
R36 B.n294 B.n293 585
R37 B.n292 B.n291 585
R38 B.n290 B.n289 585
R39 B.n288 B.n287 585
R40 B.n286 B.n285 585
R41 B.n284 B.n283 585
R42 B.n282 B.n281 585
R43 B.n280 B.n279 585
R44 B.n278 B.n277 585
R45 B.n276 B.n275 585
R46 B.n274 B.n273 585
R47 B.n272 B.n271 585
R48 B.n270 B.n269 585
R49 B.n268 B.n267 585
R50 B.n266 B.n265 585
R51 B.n264 B.n263 585
R52 B.n262 B.n261 585
R53 B.n260 B.n259 585
R54 B.n258 B.n257 585
R55 B.n256 B.n255 585
R56 B.n254 B.n253 585
R57 B.n252 B.n251 585
R58 B.n250 B.n249 585
R59 B.n248 B.n247 585
R60 B.n246 B.n245 585
R61 B.n243 B.n242 585
R62 B.n241 B.n240 585
R63 B.n239 B.n238 585
R64 B.n237 B.n236 585
R65 B.n235 B.n234 585
R66 B.n233 B.n232 585
R67 B.n231 B.n230 585
R68 B.n229 B.n228 585
R69 B.n227 B.n226 585
R70 B.n225 B.n224 585
R71 B.n223 B.n222 585
R72 B.n221 B.n220 585
R73 B.n219 B.n218 585
R74 B.n217 B.n216 585
R75 B.n215 B.n214 585
R76 B.n213 B.n212 585
R77 B.n211 B.n210 585
R78 B.n209 B.n208 585
R79 B.n207 B.n206 585
R80 B.n205 B.n204 585
R81 B.n203 B.n202 585
R82 B.n201 B.n200 585
R83 B.n199 B.n198 585
R84 B.n197 B.n196 585
R85 B.n195 B.n194 585
R86 B.n193 B.n192 585
R87 B.n191 B.n190 585
R88 B.n189 B.n188 585
R89 B.n187 B.n186 585
R90 B.n185 B.n184 585
R91 B.n183 B.n182 585
R92 B.n181 B.n180 585
R93 B.n179 B.n178 585
R94 B.n177 B.n176 585
R95 B.n175 B.n174 585
R96 B.n173 B.n172 585
R97 B.n171 B.n170 585
R98 B.n169 B.n168 585
R99 B.n167 B.n166 585
R100 B.n165 B.n164 585
R101 B.n163 B.n162 585
R102 B.n161 B.n160 585
R103 B.n159 B.n158 585
R104 B.n157 B.n156 585
R105 B.n155 B.n154 585
R106 B.n153 B.n152 585
R107 B.n151 B.n150 585
R108 B.n149 B.n148 585
R109 B.n147 B.n146 585
R110 B.n145 B.n144 585
R111 B.n143 B.n142 585
R112 B.n141 B.n140 585
R113 B.n139 B.n138 585
R114 B.n137 B.n136 585
R115 B.n135 B.n134 585
R116 B.n133 B.n132 585
R117 B.n131 B.n130 585
R118 B.n129 B.n128 585
R119 B.n127 B.n126 585
R120 B.n125 B.n124 585
R121 B.n123 B.n122 585
R122 B.n121 B.n120 585
R123 B.n119 B.n118 585
R124 B.n117 B.n116 585
R125 B.n115 B.n114 585
R126 B.n113 B.n112 585
R127 B.n111 B.n110 585
R128 B.n39 B.n38 585
R129 B.n812 B.n811 585
R130 B.n806 B.n104 585
R131 B.n104 B.n36 585
R132 B.n805 B.n35 585
R133 B.n816 B.n35 585
R134 B.n804 B.n34 585
R135 B.n817 B.n34 585
R136 B.n803 B.n33 585
R137 B.n818 B.n33 585
R138 B.n802 B.n801 585
R139 B.n801 B.n29 585
R140 B.n800 B.n28 585
R141 B.n824 B.n28 585
R142 B.n799 B.n27 585
R143 B.n825 B.n27 585
R144 B.n798 B.n26 585
R145 B.n826 B.n26 585
R146 B.n797 B.n796 585
R147 B.n796 B.n22 585
R148 B.n795 B.n21 585
R149 B.n832 B.n21 585
R150 B.n794 B.n20 585
R151 B.n833 B.n20 585
R152 B.n793 B.n19 585
R153 B.n834 B.n19 585
R154 B.n792 B.n791 585
R155 B.n791 B.n15 585
R156 B.n790 B.n14 585
R157 B.n840 B.n14 585
R158 B.n789 B.n13 585
R159 B.n841 B.n13 585
R160 B.n788 B.n12 585
R161 B.n842 B.n12 585
R162 B.n787 B.n786 585
R163 B.n786 B.n8 585
R164 B.n785 B.n7 585
R165 B.n848 B.n7 585
R166 B.n784 B.n6 585
R167 B.n849 B.n6 585
R168 B.n783 B.n5 585
R169 B.n850 B.n5 585
R170 B.n782 B.n781 585
R171 B.n781 B.n4 585
R172 B.n780 B.n362 585
R173 B.n780 B.n779 585
R174 B.n770 B.n363 585
R175 B.n364 B.n363 585
R176 B.n772 B.n771 585
R177 B.n773 B.n772 585
R178 B.n769 B.n368 585
R179 B.n372 B.n368 585
R180 B.n768 B.n767 585
R181 B.n767 B.n766 585
R182 B.n370 B.n369 585
R183 B.n371 B.n370 585
R184 B.n759 B.n758 585
R185 B.n760 B.n759 585
R186 B.n757 B.n377 585
R187 B.n377 B.n376 585
R188 B.n756 B.n755 585
R189 B.n755 B.n754 585
R190 B.n379 B.n378 585
R191 B.n380 B.n379 585
R192 B.n747 B.n746 585
R193 B.n748 B.n747 585
R194 B.n745 B.n385 585
R195 B.n385 B.n384 585
R196 B.n744 B.n743 585
R197 B.n743 B.n742 585
R198 B.n387 B.n386 585
R199 B.n388 B.n387 585
R200 B.n735 B.n734 585
R201 B.n736 B.n735 585
R202 B.n733 B.n393 585
R203 B.n393 B.n392 585
R204 B.n732 B.n731 585
R205 B.n731 B.n730 585
R206 B.n395 B.n394 585
R207 B.n396 B.n395 585
R208 B.n726 B.n725 585
R209 B.n399 B.n398 585
R210 B.n722 B.n721 585
R211 B.n723 B.n722 585
R212 B.n720 B.n463 585
R213 B.n719 B.n718 585
R214 B.n717 B.n716 585
R215 B.n715 B.n714 585
R216 B.n713 B.n712 585
R217 B.n711 B.n710 585
R218 B.n709 B.n708 585
R219 B.n707 B.n706 585
R220 B.n705 B.n704 585
R221 B.n703 B.n702 585
R222 B.n701 B.n700 585
R223 B.n699 B.n698 585
R224 B.n697 B.n696 585
R225 B.n695 B.n694 585
R226 B.n693 B.n692 585
R227 B.n691 B.n690 585
R228 B.n689 B.n688 585
R229 B.n687 B.n686 585
R230 B.n685 B.n684 585
R231 B.n683 B.n682 585
R232 B.n681 B.n680 585
R233 B.n679 B.n678 585
R234 B.n677 B.n676 585
R235 B.n675 B.n674 585
R236 B.n673 B.n672 585
R237 B.n671 B.n670 585
R238 B.n669 B.n668 585
R239 B.n667 B.n666 585
R240 B.n665 B.n664 585
R241 B.n663 B.n662 585
R242 B.n661 B.n660 585
R243 B.n659 B.n658 585
R244 B.n657 B.n656 585
R245 B.n655 B.n654 585
R246 B.n653 B.n652 585
R247 B.n651 B.n650 585
R248 B.n649 B.n648 585
R249 B.n647 B.n646 585
R250 B.n645 B.n644 585
R251 B.n643 B.n642 585
R252 B.n641 B.n640 585
R253 B.n639 B.n638 585
R254 B.n637 B.n636 585
R255 B.n635 B.n634 585
R256 B.n633 B.n632 585
R257 B.n631 B.n630 585
R258 B.n629 B.n628 585
R259 B.n627 B.n626 585
R260 B.n625 B.n624 585
R261 B.n623 B.n622 585
R262 B.n621 B.n620 585
R263 B.n619 B.n618 585
R264 B.n617 B.n616 585
R265 B.n615 B.n614 585
R266 B.n613 B.n612 585
R267 B.n611 B.n610 585
R268 B.n609 B.n608 585
R269 B.n606 B.n605 585
R270 B.n604 B.n603 585
R271 B.n602 B.n601 585
R272 B.n600 B.n599 585
R273 B.n598 B.n597 585
R274 B.n596 B.n595 585
R275 B.n594 B.n593 585
R276 B.n592 B.n591 585
R277 B.n590 B.n589 585
R278 B.n588 B.n587 585
R279 B.n586 B.n585 585
R280 B.n584 B.n583 585
R281 B.n582 B.n581 585
R282 B.n580 B.n579 585
R283 B.n578 B.n577 585
R284 B.n576 B.n575 585
R285 B.n574 B.n573 585
R286 B.n572 B.n571 585
R287 B.n570 B.n569 585
R288 B.n568 B.n567 585
R289 B.n566 B.n565 585
R290 B.n564 B.n563 585
R291 B.n562 B.n561 585
R292 B.n560 B.n559 585
R293 B.n558 B.n557 585
R294 B.n556 B.n555 585
R295 B.n554 B.n553 585
R296 B.n552 B.n551 585
R297 B.n550 B.n549 585
R298 B.n548 B.n547 585
R299 B.n546 B.n545 585
R300 B.n544 B.n543 585
R301 B.n542 B.n541 585
R302 B.n540 B.n539 585
R303 B.n538 B.n537 585
R304 B.n536 B.n535 585
R305 B.n534 B.n533 585
R306 B.n532 B.n531 585
R307 B.n530 B.n529 585
R308 B.n528 B.n527 585
R309 B.n526 B.n525 585
R310 B.n524 B.n523 585
R311 B.n522 B.n521 585
R312 B.n520 B.n519 585
R313 B.n518 B.n517 585
R314 B.n516 B.n515 585
R315 B.n514 B.n513 585
R316 B.n512 B.n511 585
R317 B.n510 B.n509 585
R318 B.n508 B.n507 585
R319 B.n506 B.n505 585
R320 B.n504 B.n503 585
R321 B.n502 B.n501 585
R322 B.n500 B.n499 585
R323 B.n498 B.n497 585
R324 B.n496 B.n495 585
R325 B.n494 B.n493 585
R326 B.n492 B.n491 585
R327 B.n490 B.n489 585
R328 B.n488 B.n487 585
R329 B.n486 B.n485 585
R330 B.n484 B.n483 585
R331 B.n482 B.n481 585
R332 B.n480 B.n479 585
R333 B.n478 B.n477 585
R334 B.n476 B.n475 585
R335 B.n474 B.n473 585
R336 B.n472 B.n471 585
R337 B.n470 B.n469 585
R338 B.n727 B.n397 585
R339 B.n397 B.n396 585
R340 B.n729 B.n728 585
R341 B.n730 B.n729 585
R342 B.n391 B.n390 585
R343 B.n392 B.n391 585
R344 B.n738 B.n737 585
R345 B.n737 B.n736 585
R346 B.n739 B.n389 585
R347 B.n389 B.n388 585
R348 B.n741 B.n740 585
R349 B.n742 B.n741 585
R350 B.n383 B.n382 585
R351 B.n384 B.n383 585
R352 B.n750 B.n749 585
R353 B.n749 B.n748 585
R354 B.n751 B.n381 585
R355 B.n381 B.n380 585
R356 B.n753 B.n752 585
R357 B.n754 B.n753 585
R358 B.n375 B.n374 585
R359 B.n376 B.n375 585
R360 B.n762 B.n761 585
R361 B.n761 B.n760 585
R362 B.n763 B.n373 585
R363 B.n373 B.n371 585
R364 B.n765 B.n764 585
R365 B.n766 B.n765 585
R366 B.n367 B.n366 585
R367 B.n372 B.n367 585
R368 B.n775 B.n774 585
R369 B.n774 B.n773 585
R370 B.n776 B.n365 585
R371 B.n365 B.n364 585
R372 B.n778 B.n777 585
R373 B.n779 B.n778 585
R374 B.n2 B.n0 585
R375 B.n4 B.n2 585
R376 B.n3 B.n1 585
R377 B.n849 B.n3 585
R378 B.n847 B.n846 585
R379 B.n848 B.n847 585
R380 B.n845 B.n9 585
R381 B.n9 B.n8 585
R382 B.n844 B.n843 585
R383 B.n843 B.n842 585
R384 B.n11 B.n10 585
R385 B.n841 B.n11 585
R386 B.n839 B.n838 585
R387 B.n840 B.n839 585
R388 B.n837 B.n16 585
R389 B.n16 B.n15 585
R390 B.n836 B.n835 585
R391 B.n835 B.n834 585
R392 B.n18 B.n17 585
R393 B.n833 B.n18 585
R394 B.n831 B.n830 585
R395 B.n832 B.n831 585
R396 B.n829 B.n23 585
R397 B.n23 B.n22 585
R398 B.n828 B.n827 585
R399 B.n827 B.n826 585
R400 B.n25 B.n24 585
R401 B.n825 B.n25 585
R402 B.n823 B.n822 585
R403 B.n824 B.n823 585
R404 B.n821 B.n30 585
R405 B.n30 B.n29 585
R406 B.n820 B.n819 585
R407 B.n819 B.n818 585
R408 B.n32 B.n31 585
R409 B.n817 B.n32 585
R410 B.n815 B.n814 585
R411 B.n816 B.n815 585
R412 B.n813 B.n37 585
R413 B.n37 B.n36 585
R414 B.n852 B.n851 585
R415 B.n851 B.n850 585
R416 B.n725 B.n397 535.745
R417 B.n811 B.n37 535.745
R418 B.n469 B.n395 535.745
R419 B.n808 B.n104 535.745
R420 B.n466 B.t6 492.387
R421 B.n464 B.t10 492.387
R422 B.n107 B.t13 492.387
R423 B.n105 B.t2 492.387
R424 B.n466 B.t9 425.238
R425 B.n464 B.t12 425.238
R426 B.n107 B.t14 425.238
R427 B.n105 B.t4 425.238
R428 B.n467 B.t8 389.166
R429 B.n106 B.t5 389.166
R430 B.n465 B.t11 389.166
R431 B.n108 B.t15 389.166
R432 B.n809 B.n102 256.663
R433 B.n809 B.n101 256.663
R434 B.n809 B.n100 256.663
R435 B.n809 B.n99 256.663
R436 B.n809 B.n98 256.663
R437 B.n809 B.n97 256.663
R438 B.n809 B.n96 256.663
R439 B.n809 B.n95 256.663
R440 B.n809 B.n94 256.663
R441 B.n809 B.n93 256.663
R442 B.n809 B.n92 256.663
R443 B.n809 B.n91 256.663
R444 B.n809 B.n90 256.663
R445 B.n809 B.n89 256.663
R446 B.n809 B.n88 256.663
R447 B.n809 B.n87 256.663
R448 B.n809 B.n86 256.663
R449 B.n809 B.n85 256.663
R450 B.n809 B.n84 256.663
R451 B.n809 B.n83 256.663
R452 B.n809 B.n82 256.663
R453 B.n809 B.n81 256.663
R454 B.n809 B.n80 256.663
R455 B.n809 B.n79 256.663
R456 B.n809 B.n78 256.663
R457 B.n809 B.n77 256.663
R458 B.n809 B.n76 256.663
R459 B.n809 B.n75 256.663
R460 B.n809 B.n74 256.663
R461 B.n809 B.n73 256.663
R462 B.n809 B.n72 256.663
R463 B.n809 B.n71 256.663
R464 B.n809 B.n70 256.663
R465 B.n809 B.n69 256.663
R466 B.n809 B.n68 256.663
R467 B.n809 B.n67 256.663
R468 B.n809 B.n66 256.663
R469 B.n809 B.n65 256.663
R470 B.n809 B.n64 256.663
R471 B.n809 B.n63 256.663
R472 B.n809 B.n62 256.663
R473 B.n809 B.n61 256.663
R474 B.n809 B.n60 256.663
R475 B.n809 B.n59 256.663
R476 B.n809 B.n58 256.663
R477 B.n809 B.n57 256.663
R478 B.n809 B.n56 256.663
R479 B.n809 B.n55 256.663
R480 B.n809 B.n54 256.663
R481 B.n809 B.n53 256.663
R482 B.n809 B.n52 256.663
R483 B.n809 B.n51 256.663
R484 B.n809 B.n50 256.663
R485 B.n809 B.n49 256.663
R486 B.n809 B.n48 256.663
R487 B.n809 B.n47 256.663
R488 B.n809 B.n46 256.663
R489 B.n809 B.n45 256.663
R490 B.n809 B.n44 256.663
R491 B.n809 B.n43 256.663
R492 B.n809 B.n42 256.663
R493 B.n809 B.n41 256.663
R494 B.n809 B.n40 256.663
R495 B.n810 B.n809 256.663
R496 B.n724 B.n723 256.663
R497 B.n723 B.n400 256.663
R498 B.n723 B.n401 256.663
R499 B.n723 B.n402 256.663
R500 B.n723 B.n403 256.663
R501 B.n723 B.n404 256.663
R502 B.n723 B.n405 256.663
R503 B.n723 B.n406 256.663
R504 B.n723 B.n407 256.663
R505 B.n723 B.n408 256.663
R506 B.n723 B.n409 256.663
R507 B.n723 B.n410 256.663
R508 B.n723 B.n411 256.663
R509 B.n723 B.n412 256.663
R510 B.n723 B.n413 256.663
R511 B.n723 B.n414 256.663
R512 B.n723 B.n415 256.663
R513 B.n723 B.n416 256.663
R514 B.n723 B.n417 256.663
R515 B.n723 B.n418 256.663
R516 B.n723 B.n419 256.663
R517 B.n723 B.n420 256.663
R518 B.n723 B.n421 256.663
R519 B.n723 B.n422 256.663
R520 B.n723 B.n423 256.663
R521 B.n723 B.n424 256.663
R522 B.n723 B.n425 256.663
R523 B.n723 B.n426 256.663
R524 B.n723 B.n427 256.663
R525 B.n723 B.n428 256.663
R526 B.n723 B.n429 256.663
R527 B.n723 B.n430 256.663
R528 B.n723 B.n431 256.663
R529 B.n723 B.n432 256.663
R530 B.n723 B.n433 256.663
R531 B.n723 B.n434 256.663
R532 B.n723 B.n435 256.663
R533 B.n723 B.n436 256.663
R534 B.n723 B.n437 256.663
R535 B.n723 B.n438 256.663
R536 B.n723 B.n439 256.663
R537 B.n723 B.n440 256.663
R538 B.n723 B.n441 256.663
R539 B.n723 B.n442 256.663
R540 B.n723 B.n443 256.663
R541 B.n723 B.n444 256.663
R542 B.n723 B.n445 256.663
R543 B.n723 B.n446 256.663
R544 B.n723 B.n447 256.663
R545 B.n723 B.n448 256.663
R546 B.n723 B.n449 256.663
R547 B.n723 B.n450 256.663
R548 B.n723 B.n451 256.663
R549 B.n723 B.n452 256.663
R550 B.n723 B.n453 256.663
R551 B.n723 B.n454 256.663
R552 B.n723 B.n455 256.663
R553 B.n723 B.n456 256.663
R554 B.n723 B.n457 256.663
R555 B.n723 B.n458 256.663
R556 B.n723 B.n459 256.663
R557 B.n723 B.n460 256.663
R558 B.n723 B.n461 256.663
R559 B.n723 B.n462 256.663
R560 B.n729 B.n397 163.367
R561 B.n729 B.n391 163.367
R562 B.n737 B.n391 163.367
R563 B.n737 B.n389 163.367
R564 B.n741 B.n389 163.367
R565 B.n741 B.n383 163.367
R566 B.n749 B.n383 163.367
R567 B.n749 B.n381 163.367
R568 B.n753 B.n381 163.367
R569 B.n753 B.n375 163.367
R570 B.n761 B.n375 163.367
R571 B.n761 B.n373 163.367
R572 B.n765 B.n373 163.367
R573 B.n765 B.n367 163.367
R574 B.n774 B.n367 163.367
R575 B.n774 B.n365 163.367
R576 B.n778 B.n365 163.367
R577 B.n778 B.n2 163.367
R578 B.n851 B.n2 163.367
R579 B.n851 B.n3 163.367
R580 B.n847 B.n3 163.367
R581 B.n847 B.n9 163.367
R582 B.n843 B.n9 163.367
R583 B.n843 B.n11 163.367
R584 B.n839 B.n11 163.367
R585 B.n839 B.n16 163.367
R586 B.n835 B.n16 163.367
R587 B.n835 B.n18 163.367
R588 B.n831 B.n18 163.367
R589 B.n831 B.n23 163.367
R590 B.n827 B.n23 163.367
R591 B.n827 B.n25 163.367
R592 B.n823 B.n25 163.367
R593 B.n823 B.n30 163.367
R594 B.n819 B.n30 163.367
R595 B.n819 B.n32 163.367
R596 B.n815 B.n32 163.367
R597 B.n815 B.n37 163.367
R598 B.n722 B.n399 163.367
R599 B.n722 B.n463 163.367
R600 B.n718 B.n717 163.367
R601 B.n714 B.n713 163.367
R602 B.n710 B.n709 163.367
R603 B.n706 B.n705 163.367
R604 B.n702 B.n701 163.367
R605 B.n698 B.n697 163.367
R606 B.n694 B.n693 163.367
R607 B.n690 B.n689 163.367
R608 B.n686 B.n685 163.367
R609 B.n682 B.n681 163.367
R610 B.n678 B.n677 163.367
R611 B.n674 B.n673 163.367
R612 B.n670 B.n669 163.367
R613 B.n666 B.n665 163.367
R614 B.n662 B.n661 163.367
R615 B.n658 B.n657 163.367
R616 B.n654 B.n653 163.367
R617 B.n650 B.n649 163.367
R618 B.n646 B.n645 163.367
R619 B.n642 B.n641 163.367
R620 B.n638 B.n637 163.367
R621 B.n634 B.n633 163.367
R622 B.n630 B.n629 163.367
R623 B.n626 B.n625 163.367
R624 B.n622 B.n621 163.367
R625 B.n618 B.n617 163.367
R626 B.n614 B.n613 163.367
R627 B.n610 B.n609 163.367
R628 B.n605 B.n604 163.367
R629 B.n601 B.n600 163.367
R630 B.n597 B.n596 163.367
R631 B.n593 B.n592 163.367
R632 B.n589 B.n588 163.367
R633 B.n585 B.n584 163.367
R634 B.n581 B.n580 163.367
R635 B.n577 B.n576 163.367
R636 B.n573 B.n572 163.367
R637 B.n569 B.n568 163.367
R638 B.n565 B.n564 163.367
R639 B.n561 B.n560 163.367
R640 B.n557 B.n556 163.367
R641 B.n553 B.n552 163.367
R642 B.n549 B.n548 163.367
R643 B.n545 B.n544 163.367
R644 B.n541 B.n540 163.367
R645 B.n537 B.n536 163.367
R646 B.n533 B.n532 163.367
R647 B.n529 B.n528 163.367
R648 B.n525 B.n524 163.367
R649 B.n521 B.n520 163.367
R650 B.n517 B.n516 163.367
R651 B.n513 B.n512 163.367
R652 B.n509 B.n508 163.367
R653 B.n505 B.n504 163.367
R654 B.n501 B.n500 163.367
R655 B.n497 B.n496 163.367
R656 B.n493 B.n492 163.367
R657 B.n489 B.n488 163.367
R658 B.n485 B.n484 163.367
R659 B.n481 B.n480 163.367
R660 B.n477 B.n476 163.367
R661 B.n473 B.n472 163.367
R662 B.n731 B.n395 163.367
R663 B.n731 B.n393 163.367
R664 B.n735 B.n393 163.367
R665 B.n735 B.n387 163.367
R666 B.n743 B.n387 163.367
R667 B.n743 B.n385 163.367
R668 B.n747 B.n385 163.367
R669 B.n747 B.n379 163.367
R670 B.n755 B.n379 163.367
R671 B.n755 B.n377 163.367
R672 B.n759 B.n377 163.367
R673 B.n759 B.n370 163.367
R674 B.n767 B.n370 163.367
R675 B.n767 B.n368 163.367
R676 B.n772 B.n368 163.367
R677 B.n772 B.n363 163.367
R678 B.n780 B.n363 163.367
R679 B.n781 B.n780 163.367
R680 B.n781 B.n5 163.367
R681 B.n6 B.n5 163.367
R682 B.n7 B.n6 163.367
R683 B.n786 B.n7 163.367
R684 B.n786 B.n12 163.367
R685 B.n13 B.n12 163.367
R686 B.n14 B.n13 163.367
R687 B.n791 B.n14 163.367
R688 B.n791 B.n19 163.367
R689 B.n20 B.n19 163.367
R690 B.n21 B.n20 163.367
R691 B.n796 B.n21 163.367
R692 B.n796 B.n26 163.367
R693 B.n27 B.n26 163.367
R694 B.n28 B.n27 163.367
R695 B.n801 B.n28 163.367
R696 B.n801 B.n33 163.367
R697 B.n34 B.n33 163.367
R698 B.n35 B.n34 163.367
R699 B.n104 B.n35 163.367
R700 B.n110 B.n39 163.367
R701 B.n114 B.n113 163.367
R702 B.n118 B.n117 163.367
R703 B.n122 B.n121 163.367
R704 B.n126 B.n125 163.367
R705 B.n130 B.n129 163.367
R706 B.n134 B.n133 163.367
R707 B.n138 B.n137 163.367
R708 B.n142 B.n141 163.367
R709 B.n146 B.n145 163.367
R710 B.n150 B.n149 163.367
R711 B.n154 B.n153 163.367
R712 B.n158 B.n157 163.367
R713 B.n162 B.n161 163.367
R714 B.n166 B.n165 163.367
R715 B.n170 B.n169 163.367
R716 B.n174 B.n173 163.367
R717 B.n178 B.n177 163.367
R718 B.n182 B.n181 163.367
R719 B.n186 B.n185 163.367
R720 B.n190 B.n189 163.367
R721 B.n194 B.n193 163.367
R722 B.n198 B.n197 163.367
R723 B.n202 B.n201 163.367
R724 B.n206 B.n205 163.367
R725 B.n210 B.n209 163.367
R726 B.n214 B.n213 163.367
R727 B.n218 B.n217 163.367
R728 B.n222 B.n221 163.367
R729 B.n226 B.n225 163.367
R730 B.n230 B.n229 163.367
R731 B.n234 B.n233 163.367
R732 B.n238 B.n237 163.367
R733 B.n242 B.n241 163.367
R734 B.n247 B.n246 163.367
R735 B.n251 B.n250 163.367
R736 B.n255 B.n254 163.367
R737 B.n259 B.n258 163.367
R738 B.n263 B.n262 163.367
R739 B.n267 B.n266 163.367
R740 B.n271 B.n270 163.367
R741 B.n275 B.n274 163.367
R742 B.n279 B.n278 163.367
R743 B.n283 B.n282 163.367
R744 B.n287 B.n286 163.367
R745 B.n291 B.n290 163.367
R746 B.n295 B.n294 163.367
R747 B.n299 B.n298 163.367
R748 B.n303 B.n302 163.367
R749 B.n307 B.n306 163.367
R750 B.n311 B.n310 163.367
R751 B.n315 B.n314 163.367
R752 B.n319 B.n318 163.367
R753 B.n323 B.n322 163.367
R754 B.n327 B.n326 163.367
R755 B.n331 B.n330 163.367
R756 B.n335 B.n334 163.367
R757 B.n339 B.n338 163.367
R758 B.n343 B.n342 163.367
R759 B.n347 B.n346 163.367
R760 B.n351 B.n350 163.367
R761 B.n355 B.n354 163.367
R762 B.n359 B.n358 163.367
R763 B.n808 B.n103 163.367
R764 B.n725 B.n724 71.676
R765 B.n463 B.n400 71.676
R766 B.n717 B.n401 71.676
R767 B.n713 B.n402 71.676
R768 B.n709 B.n403 71.676
R769 B.n705 B.n404 71.676
R770 B.n701 B.n405 71.676
R771 B.n697 B.n406 71.676
R772 B.n693 B.n407 71.676
R773 B.n689 B.n408 71.676
R774 B.n685 B.n409 71.676
R775 B.n681 B.n410 71.676
R776 B.n677 B.n411 71.676
R777 B.n673 B.n412 71.676
R778 B.n669 B.n413 71.676
R779 B.n665 B.n414 71.676
R780 B.n661 B.n415 71.676
R781 B.n657 B.n416 71.676
R782 B.n653 B.n417 71.676
R783 B.n649 B.n418 71.676
R784 B.n645 B.n419 71.676
R785 B.n641 B.n420 71.676
R786 B.n637 B.n421 71.676
R787 B.n633 B.n422 71.676
R788 B.n629 B.n423 71.676
R789 B.n625 B.n424 71.676
R790 B.n621 B.n425 71.676
R791 B.n617 B.n426 71.676
R792 B.n613 B.n427 71.676
R793 B.n609 B.n428 71.676
R794 B.n604 B.n429 71.676
R795 B.n600 B.n430 71.676
R796 B.n596 B.n431 71.676
R797 B.n592 B.n432 71.676
R798 B.n588 B.n433 71.676
R799 B.n584 B.n434 71.676
R800 B.n580 B.n435 71.676
R801 B.n576 B.n436 71.676
R802 B.n572 B.n437 71.676
R803 B.n568 B.n438 71.676
R804 B.n564 B.n439 71.676
R805 B.n560 B.n440 71.676
R806 B.n556 B.n441 71.676
R807 B.n552 B.n442 71.676
R808 B.n548 B.n443 71.676
R809 B.n544 B.n444 71.676
R810 B.n540 B.n445 71.676
R811 B.n536 B.n446 71.676
R812 B.n532 B.n447 71.676
R813 B.n528 B.n448 71.676
R814 B.n524 B.n449 71.676
R815 B.n520 B.n450 71.676
R816 B.n516 B.n451 71.676
R817 B.n512 B.n452 71.676
R818 B.n508 B.n453 71.676
R819 B.n504 B.n454 71.676
R820 B.n500 B.n455 71.676
R821 B.n496 B.n456 71.676
R822 B.n492 B.n457 71.676
R823 B.n488 B.n458 71.676
R824 B.n484 B.n459 71.676
R825 B.n480 B.n460 71.676
R826 B.n476 B.n461 71.676
R827 B.n472 B.n462 71.676
R828 B.n811 B.n810 71.676
R829 B.n110 B.n40 71.676
R830 B.n114 B.n41 71.676
R831 B.n118 B.n42 71.676
R832 B.n122 B.n43 71.676
R833 B.n126 B.n44 71.676
R834 B.n130 B.n45 71.676
R835 B.n134 B.n46 71.676
R836 B.n138 B.n47 71.676
R837 B.n142 B.n48 71.676
R838 B.n146 B.n49 71.676
R839 B.n150 B.n50 71.676
R840 B.n154 B.n51 71.676
R841 B.n158 B.n52 71.676
R842 B.n162 B.n53 71.676
R843 B.n166 B.n54 71.676
R844 B.n170 B.n55 71.676
R845 B.n174 B.n56 71.676
R846 B.n178 B.n57 71.676
R847 B.n182 B.n58 71.676
R848 B.n186 B.n59 71.676
R849 B.n190 B.n60 71.676
R850 B.n194 B.n61 71.676
R851 B.n198 B.n62 71.676
R852 B.n202 B.n63 71.676
R853 B.n206 B.n64 71.676
R854 B.n210 B.n65 71.676
R855 B.n214 B.n66 71.676
R856 B.n218 B.n67 71.676
R857 B.n222 B.n68 71.676
R858 B.n226 B.n69 71.676
R859 B.n230 B.n70 71.676
R860 B.n234 B.n71 71.676
R861 B.n238 B.n72 71.676
R862 B.n242 B.n73 71.676
R863 B.n247 B.n74 71.676
R864 B.n251 B.n75 71.676
R865 B.n255 B.n76 71.676
R866 B.n259 B.n77 71.676
R867 B.n263 B.n78 71.676
R868 B.n267 B.n79 71.676
R869 B.n271 B.n80 71.676
R870 B.n275 B.n81 71.676
R871 B.n279 B.n82 71.676
R872 B.n283 B.n83 71.676
R873 B.n287 B.n84 71.676
R874 B.n291 B.n85 71.676
R875 B.n295 B.n86 71.676
R876 B.n299 B.n87 71.676
R877 B.n303 B.n88 71.676
R878 B.n307 B.n89 71.676
R879 B.n311 B.n90 71.676
R880 B.n315 B.n91 71.676
R881 B.n319 B.n92 71.676
R882 B.n323 B.n93 71.676
R883 B.n327 B.n94 71.676
R884 B.n331 B.n95 71.676
R885 B.n335 B.n96 71.676
R886 B.n339 B.n97 71.676
R887 B.n343 B.n98 71.676
R888 B.n347 B.n99 71.676
R889 B.n351 B.n100 71.676
R890 B.n355 B.n101 71.676
R891 B.n359 B.n102 71.676
R892 B.n103 B.n102 71.676
R893 B.n358 B.n101 71.676
R894 B.n354 B.n100 71.676
R895 B.n350 B.n99 71.676
R896 B.n346 B.n98 71.676
R897 B.n342 B.n97 71.676
R898 B.n338 B.n96 71.676
R899 B.n334 B.n95 71.676
R900 B.n330 B.n94 71.676
R901 B.n326 B.n93 71.676
R902 B.n322 B.n92 71.676
R903 B.n318 B.n91 71.676
R904 B.n314 B.n90 71.676
R905 B.n310 B.n89 71.676
R906 B.n306 B.n88 71.676
R907 B.n302 B.n87 71.676
R908 B.n298 B.n86 71.676
R909 B.n294 B.n85 71.676
R910 B.n290 B.n84 71.676
R911 B.n286 B.n83 71.676
R912 B.n282 B.n82 71.676
R913 B.n278 B.n81 71.676
R914 B.n274 B.n80 71.676
R915 B.n270 B.n79 71.676
R916 B.n266 B.n78 71.676
R917 B.n262 B.n77 71.676
R918 B.n258 B.n76 71.676
R919 B.n254 B.n75 71.676
R920 B.n250 B.n74 71.676
R921 B.n246 B.n73 71.676
R922 B.n241 B.n72 71.676
R923 B.n237 B.n71 71.676
R924 B.n233 B.n70 71.676
R925 B.n229 B.n69 71.676
R926 B.n225 B.n68 71.676
R927 B.n221 B.n67 71.676
R928 B.n217 B.n66 71.676
R929 B.n213 B.n65 71.676
R930 B.n209 B.n64 71.676
R931 B.n205 B.n63 71.676
R932 B.n201 B.n62 71.676
R933 B.n197 B.n61 71.676
R934 B.n193 B.n60 71.676
R935 B.n189 B.n59 71.676
R936 B.n185 B.n58 71.676
R937 B.n181 B.n57 71.676
R938 B.n177 B.n56 71.676
R939 B.n173 B.n55 71.676
R940 B.n169 B.n54 71.676
R941 B.n165 B.n53 71.676
R942 B.n161 B.n52 71.676
R943 B.n157 B.n51 71.676
R944 B.n153 B.n50 71.676
R945 B.n149 B.n49 71.676
R946 B.n145 B.n48 71.676
R947 B.n141 B.n47 71.676
R948 B.n137 B.n46 71.676
R949 B.n133 B.n45 71.676
R950 B.n129 B.n44 71.676
R951 B.n125 B.n43 71.676
R952 B.n121 B.n42 71.676
R953 B.n117 B.n41 71.676
R954 B.n113 B.n40 71.676
R955 B.n810 B.n39 71.676
R956 B.n724 B.n399 71.676
R957 B.n718 B.n400 71.676
R958 B.n714 B.n401 71.676
R959 B.n710 B.n402 71.676
R960 B.n706 B.n403 71.676
R961 B.n702 B.n404 71.676
R962 B.n698 B.n405 71.676
R963 B.n694 B.n406 71.676
R964 B.n690 B.n407 71.676
R965 B.n686 B.n408 71.676
R966 B.n682 B.n409 71.676
R967 B.n678 B.n410 71.676
R968 B.n674 B.n411 71.676
R969 B.n670 B.n412 71.676
R970 B.n666 B.n413 71.676
R971 B.n662 B.n414 71.676
R972 B.n658 B.n415 71.676
R973 B.n654 B.n416 71.676
R974 B.n650 B.n417 71.676
R975 B.n646 B.n418 71.676
R976 B.n642 B.n419 71.676
R977 B.n638 B.n420 71.676
R978 B.n634 B.n421 71.676
R979 B.n630 B.n422 71.676
R980 B.n626 B.n423 71.676
R981 B.n622 B.n424 71.676
R982 B.n618 B.n425 71.676
R983 B.n614 B.n426 71.676
R984 B.n610 B.n427 71.676
R985 B.n605 B.n428 71.676
R986 B.n601 B.n429 71.676
R987 B.n597 B.n430 71.676
R988 B.n593 B.n431 71.676
R989 B.n589 B.n432 71.676
R990 B.n585 B.n433 71.676
R991 B.n581 B.n434 71.676
R992 B.n577 B.n435 71.676
R993 B.n573 B.n436 71.676
R994 B.n569 B.n437 71.676
R995 B.n565 B.n438 71.676
R996 B.n561 B.n439 71.676
R997 B.n557 B.n440 71.676
R998 B.n553 B.n441 71.676
R999 B.n549 B.n442 71.676
R1000 B.n545 B.n443 71.676
R1001 B.n541 B.n444 71.676
R1002 B.n537 B.n445 71.676
R1003 B.n533 B.n446 71.676
R1004 B.n529 B.n447 71.676
R1005 B.n525 B.n448 71.676
R1006 B.n521 B.n449 71.676
R1007 B.n517 B.n450 71.676
R1008 B.n513 B.n451 71.676
R1009 B.n509 B.n452 71.676
R1010 B.n505 B.n453 71.676
R1011 B.n501 B.n454 71.676
R1012 B.n497 B.n455 71.676
R1013 B.n493 B.n456 71.676
R1014 B.n489 B.n457 71.676
R1015 B.n485 B.n458 71.676
R1016 B.n481 B.n459 71.676
R1017 B.n477 B.n460 71.676
R1018 B.n473 B.n461 71.676
R1019 B.n469 B.n462 71.676
R1020 B.n468 B.n467 59.5399
R1021 B.n607 B.n465 59.5399
R1022 B.n109 B.n108 59.5399
R1023 B.n244 B.n106 59.5399
R1024 B.n723 B.n396 59.4853
R1025 B.n809 B.n36 59.4853
R1026 B.n467 B.n466 36.0732
R1027 B.n465 B.n464 36.0732
R1028 B.n108 B.n107 36.0732
R1029 B.n106 B.n105 36.0732
R1030 B.n813 B.n812 34.8103
R1031 B.n807 B.n806 34.8103
R1032 B.n470 B.n394 34.8103
R1033 B.n727 B.n726 34.8103
R1034 B.n730 B.n396 31.8506
R1035 B.n730 B.n392 31.8506
R1036 B.n736 B.n392 31.8506
R1037 B.n736 B.n388 31.8506
R1038 B.n742 B.n388 31.8506
R1039 B.n748 B.n384 31.8506
R1040 B.n748 B.n380 31.8506
R1041 B.n754 B.n380 31.8506
R1042 B.n754 B.n376 31.8506
R1043 B.n760 B.n376 31.8506
R1044 B.n760 B.n371 31.8506
R1045 B.n766 B.n371 31.8506
R1046 B.n766 B.n372 31.8506
R1047 B.n773 B.n364 31.8506
R1048 B.n779 B.n364 31.8506
R1049 B.n779 B.n4 31.8506
R1050 B.n850 B.n4 31.8506
R1051 B.n850 B.n849 31.8506
R1052 B.n849 B.n848 31.8506
R1053 B.n848 B.n8 31.8506
R1054 B.n842 B.n8 31.8506
R1055 B.n841 B.n840 31.8506
R1056 B.n840 B.n15 31.8506
R1057 B.n834 B.n15 31.8506
R1058 B.n834 B.n833 31.8506
R1059 B.n833 B.n832 31.8506
R1060 B.n832 B.n22 31.8506
R1061 B.n826 B.n22 31.8506
R1062 B.n826 B.n825 31.8506
R1063 B.n824 B.n29 31.8506
R1064 B.n818 B.n29 31.8506
R1065 B.n818 B.n817 31.8506
R1066 B.n817 B.n816 31.8506
R1067 B.n816 B.n36 31.8506
R1068 B.n742 B.t7 31.3822
R1069 B.t3 B.n824 31.3822
R1070 B.n372 B.t1 21.0778
R1071 B.t0 B.n841 21.0778
R1072 B B.n852 18.0485
R1073 B.n773 B.t1 10.7733
R1074 B.n842 B.t0 10.7733
R1075 B.n812 B.n38 10.6151
R1076 B.n111 B.n38 10.6151
R1077 B.n112 B.n111 10.6151
R1078 B.n115 B.n112 10.6151
R1079 B.n116 B.n115 10.6151
R1080 B.n119 B.n116 10.6151
R1081 B.n120 B.n119 10.6151
R1082 B.n123 B.n120 10.6151
R1083 B.n124 B.n123 10.6151
R1084 B.n127 B.n124 10.6151
R1085 B.n128 B.n127 10.6151
R1086 B.n131 B.n128 10.6151
R1087 B.n132 B.n131 10.6151
R1088 B.n135 B.n132 10.6151
R1089 B.n136 B.n135 10.6151
R1090 B.n139 B.n136 10.6151
R1091 B.n140 B.n139 10.6151
R1092 B.n143 B.n140 10.6151
R1093 B.n144 B.n143 10.6151
R1094 B.n147 B.n144 10.6151
R1095 B.n148 B.n147 10.6151
R1096 B.n151 B.n148 10.6151
R1097 B.n152 B.n151 10.6151
R1098 B.n155 B.n152 10.6151
R1099 B.n156 B.n155 10.6151
R1100 B.n159 B.n156 10.6151
R1101 B.n160 B.n159 10.6151
R1102 B.n163 B.n160 10.6151
R1103 B.n164 B.n163 10.6151
R1104 B.n167 B.n164 10.6151
R1105 B.n168 B.n167 10.6151
R1106 B.n171 B.n168 10.6151
R1107 B.n172 B.n171 10.6151
R1108 B.n175 B.n172 10.6151
R1109 B.n176 B.n175 10.6151
R1110 B.n179 B.n176 10.6151
R1111 B.n180 B.n179 10.6151
R1112 B.n183 B.n180 10.6151
R1113 B.n184 B.n183 10.6151
R1114 B.n187 B.n184 10.6151
R1115 B.n188 B.n187 10.6151
R1116 B.n191 B.n188 10.6151
R1117 B.n192 B.n191 10.6151
R1118 B.n195 B.n192 10.6151
R1119 B.n196 B.n195 10.6151
R1120 B.n199 B.n196 10.6151
R1121 B.n200 B.n199 10.6151
R1122 B.n203 B.n200 10.6151
R1123 B.n204 B.n203 10.6151
R1124 B.n207 B.n204 10.6151
R1125 B.n208 B.n207 10.6151
R1126 B.n211 B.n208 10.6151
R1127 B.n212 B.n211 10.6151
R1128 B.n215 B.n212 10.6151
R1129 B.n216 B.n215 10.6151
R1130 B.n219 B.n216 10.6151
R1131 B.n220 B.n219 10.6151
R1132 B.n223 B.n220 10.6151
R1133 B.n224 B.n223 10.6151
R1134 B.n228 B.n227 10.6151
R1135 B.n231 B.n228 10.6151
R1136 B.n232 B.n231 10.6151
R1137 B.n235 B.n232 10.6151
R1138 B.n236 B.n235 10.6151
R1139 B.n239 B.n236 10.6151
R1140 B.n240 B.n239 10.6151
R1141 B.n243 B.n240 10.6151
R1142 B.n248 B.n245 10.6151
R1143 B.n249 B.n248 10.6151
R1144 B.n252 B.n249 10.6151
R1145 B.n253 B.n252 10.6151
R1146 B.n256 B.n253 10.6151
R1147 B.n257 B.n256 10.6151
R1148 B.n260 B.n257 10.6151
R1149 B.n261 B.n260 10.6151
R1150 B.n264 B.n261 10.6151
R1151 B.n265 B.n264 10.6151
R1152 B.n268 B.n265 10.6151
R1153 B.n269 B.n268 10.6151
R1154 B.n272 B.n269 10.6151
R1155 B.n273 B.n272 10.6151
R1156 B.n276 B.n273 10.6151
R1157 B.n277 B.n276 10.6151
R1158 B.n280 B.n277 10.6151
R1159 B.n281 B.n280 10.6151
R1160 B.n284 B.n281 10.6151
R1161 B.n285 B.n284 10.6151
R1162 B.n288 B.n285 10.6151
R1163 B.n289 B.n288 10.6151
R1164 B.n292 B.n289 10.6151
R1165 B.n293 B.n292 10.6151
R1166 B.n296 B.n293 10.6151
R1167 B.n297 B.n296 10.6151
R1168 B.n300 B.n297 10.6151
R1169 B.n301 B.n300 10.6151
R1170 B.n304 B.n301 10.6151
R1171 B.n305 B.n304 10.6151
R1172 B.n308 B.n305 10.6151
R1173 B.n309 B.n308 10.6151
R1174 B.n312 B.n309 10.6151
R1175 B.n313 B.n312 10.6151
R1176 B.n316 B.n313 10.6151
R1177 B.n317 B.n316 10.6151
R1178 B.n320 B.n317 10.6151
R1179 B.n321 B.n320 10.6151
R1180 B.n324 B.n321 10.6151
R1181 B.n325 B.n324 10.6151
R1182 B.n328 B.n325 10.6151
R1183 B.n329 B.n328 10.6151
R1184 B.n332 B.n329 10.6151
R1185 B.n333 B.n332 10.6151
R1186 B.n336 B.n333 10.6151
R1187 B.n337 B.n336 10.6151
R1188 B.n340 B.n337 10.6151
R1189 B.n341 B.n340 10.6151
R1190 B.n344 B.n341 10.6151
R1191 B.n345 B.n344 10.6151
R1192 B.n348 B.n345 10.6151
R1193 B.n349 B.n348 10.6151
R1194 B.n352 B.n349 10.6151
R1195 B.n353 B.n352 10.6151
R1196 B.n356 B.n353 10.6151
R1197 B.n357 B.n356 10.6151
R1198 B.n360 B.n357 10.6151
R1199 B.n361 B.n360 10.6151
R1200 B.n807 B.n361 10.6151
R1201 B.n732 B.n394 10.6151
R1202 B.n733 B.n732 10.6151
R1203 B.n734 B.n733 10.6151
R1204 B.n734 B.n386 10.6151
R1205 B.n744 B.n386 10.6151
R1206 B.n745 B.n744 10.6151
R1207 B.n746 B.n745 10.6151
R1208 B.n746 B.n378 10.6151
R1209 B.n756 B.n378 10.6151
R1210 B.n757 B.n756 10.6151
R1211 B.n758 B.n757 10.6151
R1212 B.n758 B.n369 10.6151
R1213 B.n768 B.n369 10.6151
R1214 B.n769 B.n768 10.6151
R1215 B.n771 B.n769 10.6151
R1216 B.n771 B.n770 10.6151
R1217 B.n770 B.n362 10.6151
R1218 B.n782 B.n362 10.6151
R1219 B.n783 B.n782 10.6151
R1220 B.n784 B.n783 10.6151
R1221 B.n785 B.n784 10.6151
R1222 B.n787 B.n785 10.6151
R1223 B.n788 B.n787 10.6151
R1224 B.n789 B.n788 10.6151
R1225 B.n790 B.n789 10.6151
R1226 B.n792 B.n790 10.6151
R1227 B.n793 B.n792 10.6151
R1228 B.n794 B.n793 10.6151
R1229 B.n795 B.n794 10.6151
R1230 B.n797 B.n795 10.6151
R1231 B.n798 B.n797 10.6151
R1232 B.n799 B.n798 10.6151
R1233 B.n800 B.n799 10.6151
R1234 B.n802 B.n800 10.6151
R1235 B.n803 B.n802 10.6151
R1236 B.n804 B.n803 10.6151
R1237 B.n805 B.n804 10.6151
R1238 B.n806 B.n805 10.6151
R1239 B.n726 B.n398 10.6151
R1240 B.n721 B.n398 10.6151
R1241 B.n721 B.n720 10.6151
R1242 B.n720 B.n719 10.6151
R1243 B.n719 B.n716 10.6151
R1244 B.n716 B.n715 10.6151
R1245 B.n715 B.n712 10.6151
R1246 B.n712 B.n711 10.6151
R1247 B.n711 B.n708 10.6151
R1248 B.n708 B.n707 10.6151
R1249 B.n707 B.n704 10.6151
R1250 B.n704 B.n703 10.6151
R1251 B.n703 B.n700 10.6151
R1252 B.n700 B.n699 10.6151
R1253 B.n699 B.n696 10.6151
R1254 B.n696 B.n695 10.6151
R1255 B.n695 B.n692 10.6151
R1256 B.n692 B.n691 10.6151
R1257 B.n691 B.n688 10.6151
R1258 B.n688 B.n687 10.6151
R1259 B.n687 B.n684 10.6151
R1260 B.n684 B.n683 10.6151
R1261 B.n683 B.n680 10.6151
R1262 B.n680 B.n679 10.6151
R1263 B.n679 B.n676 10.6151
R1264 B.n676 B.n675 10.6151
R1265 B.n675 B.n672 10.6151
R1266 B.n672 B.n671 10.6151
R1267 B.n671 B.n668 10.6151
R1268 B.n668 B.n667 10.6151
R1269 B.n667 B.n664 10.6151
R1270 B.n664 B.n663 10.6151
R1271 B.n663 B.n660 10.6151
R1272 B.n660 B.n659 10.6151
R1273 B.n659 B.n656 10.6151
R1274 B.n656 B.n655 10.6151
R1275 B.n655 B.n652 10.6151
R1276 B.n652 B.n651 10.6151
R1277 B.n651 B.n648 10.6151
R1278 B.n648 B.n647 10.6151
R1279 B.n647 B.n644 10.6151
R1280 B.n644 B.n643 10.6151
R1281 B.n643 B.n640 10.6151
R1282 B.n640 B.n639 10.6151
R1283 B.n639 B.n636 10.6151
R1284 B.n636 B.n635 10.6151
R1285 B.n635 B.n632 10.6151
R1286 B.n632 B.n631 10.6151
R1287 B.n631 B.n628 10.6151
R1288 B.n628 B.n627 10.6151
R1289 B.n627 B.n624 10.6151
R1290 B.n624 B.n623 10.6151
R1291 B.n623 B.n620 10.6151
R1292 B.n620 B.n619 10.6151
R1293 B.n619 B.n616 10.6151
R1294 B.n616 B.n615 10.6151
R1295 B.n615 B.n612 10.6151
R1296 B.n612 B.n611 10.6151
R1297 B.n611 B.n608 10.6151
R1298 B.n606 B.n603 10.6151
R1299 B.n603 B.n602 10.6151
R1300 B.n602 B.n599 10.6151
R1301 B.n599 B.n598 10.6151
R1302 B.n598 B.n595 10.6151
R1303 B.n595 B.n594 10.6151
R1304 B.n594 B.n591 10.6151
R1305 B.n591 B.n590 10.6151
R1306 B.n587 B.n586 10.6151
R1307 B.n586 B.n583 10.6151
R1308 B.n583 B.n582 10.6151
R1309 B.n582 B.n579 10.6151
R1310 B.n579 B.n578 10.6151
R1311 B.n578 B.n575 10.6151
R1312 B.n575 B.n574 10.6151
R1313 B.n574 B.n571 10.6151
R1314 B.n571 B.n570 10.6151
R1315 B.n570 B.n567 10.6151
R1316 B.n567 B.n566 10.6151
R1317 B.n566 B.n563 10.6151
R1318 B.n563 B.n562 10.6151
R1319 B.n562 B.n559 10.6151
R1320 B.n559 B.n558 10.6151
R1321 B.n558 B.n555 10.6151
R1322 B.n555 B.n554 10.6151
R1323 B.n554 B.n551 10.6151
R1324 B.n551 B.n550 10.6151
R1325 B.n550 B.n547 10.6151
R1326 B.n547 B.n546 10.6151
R1327 B.n546 B.n543 10.6151
R1328 B.n543 B.n542 10.6151
R1329 B.n542 B.n539 10.6151
R1330 B.n539 B.n538 10.6151
R1331 B.n538 B.n535 10.6151
R1332 B.n535 B.n534 10.6151
R1333 B.n534 B.n531 10.6151
R1334 B.n531 B.n530 10.6151
R1335 B.n530 B.n527 10.6151
R1336 B.n527 B.n526 10.6151
R1337 B.n526 B.n523 10.6151
R1338 B.n523 B.n522 10.6151
R1339 B.n522 B.n519 10.6151
R1340 B.n519 B.n518 10.6151
R1341 B.n518 B.n515 10.6151
R1342 B.n515 B.n514 10.6151
R1343 B.n514 B.n511 10.6151
R1344 B.n511 B.n510 10.6151
R1345 B.n510 B.n507 10.6151
R1346 B.n507 B.n506 10.6151
R1347 B.n506 B.n503 10.6151
R1348 B.n503 B.n502 10.6151
R1349 B.n502 B.n499 10.6151
R1350 B.n499 B.n498 10.6151
R1351 B.n498 B.n495 10.6151
R1352 B.n495 B.n494 10.6151
R1353 B.n494 B.n491 10.6151
R1354 B.n491 B.n490 10.6151
R1355 B.n490 B.n487 10.6151
R1356 B.n487 B.n486 10.6151
R1357 B.n486 B.n483 10.6151
R1358 B.n483 B.n482 10.6151
R1359 B.n482 B.n479 10.6151
R1360 B.n479 B.n478 10.6151
R1361 B.n478 B.n475 10.6151
R1362 B.n475 B.n474 10.6151
R1363 B.n474 B.n471 10.6151
R1364 B.n471 B.n470 10.6151
R1365 B.n728 B.n727 10.6151
R1366 B.n728 B.n390 10.6151
R1367 B.n738 B.n390 10.6151
R1368 B.n739 B.n738 10.6151
R1369 B.n740 B.n739 10.6151
R1370 B.n740 B.n382 10.6151
R1371 B.n750 B.n382 10.6151
R1372 B.n751 B.n750 10.6151
R1373 B.n752 B.n751 10.6151
R1374 B.n752 B.n374 10.6151
R1375 B.n762 B.n374 10.6151
R1376 B.n763 B.n762 10.6151
R1377 B.n764 B.n763 10.6151
R1378 B.n764 B.n366 10.6151
R1379 B.n775 B.n366 10.6151
R1380 B.n776 B.n775 10.6151
R1381 B.n777 B.n776 10.6151
R1382 B.n777 B.n0 10.6151
R1383 B.n846 B.n1 10.6151
R1384 B.n846 B.n845 10.6151
R1385 B.n845 B.n844 10.6151
R1386 B.n844 B.n10 10.6151
R1387 B.n838 B.n10 10.6151
R1388 B.n838 B.n837 10.6151
R1389 B.n837 B.n836 10.6151
R1390 B.n836 B.n17 10.6151
R1391 B.n830 B.n17 10.6151
R1392 B.n830 B.n829 10.6151
R1393 B.n829 B.n828 10.6151
R1394 B.n828 B.n24 10.6151
R1395 B.n822 B.n24 10.6151
R1396 B.n822 B.n821 10.6151
R1397 B.n821 B.n820 10.6151
R1398 B.n820 B.n31 10.6151
R1399 B.n814 B.n31 10.6151
R1400 B.n814 B.n813 10.6151
R1401 B.n227 B.n109 6.5566
R1402 B.n244 B.n243 6.5566
R1403 B.n607 B.n606 6.5566
R1404 B.n590 B.n468 6.5566
R1405 B.n224 B.n109 4.05904
R1406 B.n245 B.n244 4.05904
R1407 B.n608 B.n607 4.05904
R1408 B.n587 B.n468 4.05904
R1409 B.n852 B.n0 2.81026
R1410 B.n852 B.n1 2.81026
R1411 B.t7 B.n384 0.468884
R1412 B.n825 B.t3 0.468884
R1413 VP.n0 VP.t1 439.798
R1414 VP.n0 VP.t0 393.274
R1415 VP VP.n0 0.146778
R1416 VTAIL.n402 VTAIL.n306 289.615
R1417 VTAIL.n96 VTAIL.n0 289.615
R1418 VTAIL.n300 VTAIL.n204 289.615
R1419 VTAIL.n198 VTAIL.n102 289.615
R1420 VTAIL.n338 VTAIL.n337 185
R1421 VTAIL.n343 VTAIL.n342 185
R1422 VTAIL.n345 VTAIL.n344 185
R1423 VTAIL.n334 VTAIL.n333 185
R1424 VTAIL.n351 VTAIL.n350 185
R1425 VTAIL.n353 VTAIL.n352 185
R1426 VTAIL.n330 VTAIL.n329 185
R1427 VTAIL.n359 VTAIL.n358 185
R1428 VTAIL.n361 VTAIL.n360 185
R1429 VTAIL.n326 VTAIL.n325 185
R1430 VTAIL.n367 VTAIL.n366 185
R1431 VTAIL.n369 VTAIL.n368 185
R1432 VTAIL.n322 VTAIL.n321 185
R1433 VTAIL.n375 VTAIL.n374 185
R1434 VTAIL.n377 VTAIL.n376 185
R1435 VTAIL.n318 VTAIL.n317 185
R1436 VTAIL.n384 VTAIL.n383 185
R1437 VTAIL.n385 VTAIL.n316 185
R1438 VTAIL.n387 VTAIL.n386 185
R1439 VTAIL.n314 VTAIL.n313 185
R1440 VTAIL.n393 VTAIL.n392 185
R1441 VTAIL.n395 VTAIL.n394 185
R1442 VTAIL.n310 VTAIL.n309 185
R1443 VTAIL.n401 VTAIL.n400 185
R1444 VTAIL.n403 VTAIL.n402 185
R1445 VTAIL.n32 VTAIL.n31 185
R1446 VTAIL.n37 VTAIL.n36 185
R1447 VTAIL.n39 VTAIL.n38 185
R1448 VTAIL.n28 VTAIL.n27 185
R1449 VTAIL.n45 VTAIL.n44 185
R1450 VTAIL.n47 VTAIL.n46 185
R1451 VTAIL.n24 VTAIL.n23 185
R1452 VTAIL.n53 VTAIL.n52 185
R1453 VTAIL.n55 VTAIL.n54 185
R1454 VTAIL.n20 VTAIL.n19 185
R1455 VTAIL.n61 VTAIL.n60 185
R1456 VTAIL.n63 VTAIL.n62 185
R1457 VTAIL.n16 VTAIL.n15 185
R1458 VTAIL.n69 VTAIL.n68 185
R1459 VTAIL.n71 VTAIL.n70 185
R1460 VTAIL.n12 VTAIL.n11 185
R1461 VTAIL.n78 VTAIL.n77 185
R1462 VTAIL.n79 VTAIL.n10 185
R1463 VTAIL.n81 VTAIL.n80 185
R1464 VTAIL.n8 VTAIL.n7 185
R1465 VTAIL.n87 VTAIL.n86 185
R1466 VTAIL.n89 VTAIL.n88 185
R1467 VTAIL.n4 VTAIL.n3 185
R1468 VTAIL.n95 VTAIL.n94 185
R1469 VTAIL.n97 VTAIL.n96 185
R1470 VTAIL.n301 VTAIL.n300 185
R1471 VTAIL.n299 VTAIL.n298 185
R1472 VTAIL.n208 VTAIL.n207 185
R1473 VTAIL.n293 VTAIL.n292 185
R1474 VTAIL.n291 VTAIL.n290 185
R1475 VTAIL.n212 VTAIL.n211 185
R1476 VTAIL.n285 VTAIL.n284 185
R1477 VTAIL.n283 VTAIL.n214 185
R1478 VTAIL.n282 VTAIL.n281 185
R1479 VTAIL.n217 VTAIL.n215 185
R1480 VTAIL.n276 VTAIL.n275 185
R1481 VTAIL.n274 VTAIL.n273 185
R1482 VTAIL.n221 VTAIL.n220 185
R1483 VTAIL.n268 VTAIL.n267 185
R1484 VTAIL.n266 VTAIL.n265 185
R1485 VTAIL.n225 VTAIL.n224 185
R1486 VTAIL.n260 VTAIL.n259 185
R1487 VTAIL.n258 VTAIL.n257 185
R1488 VTAIL.n229 VTAIL.n228 185
R1489 VTAIL.n252 VTAIL.n251 185
R1490 VTAIL.n250 VTAIL.n249 185
R1491 VTAIL.n233 VTAIL.n232 185
R1492 VTAIL.n244 VTAIL.n243 185
R1493 VTAIL.n242 VTAIL.n241 185
R1494 VTAIL.n237 VTAIL.n236 185
R1495 VTAIL.n199 VTAIL.n198 185
R1496 VTAIL.n197 VTAIL.n196 185
R1497 VTAIL.n106 VTAIL.n105 185
R1498 VTAIL.n191 VTAIL.n190 185
R1499 VTAIL.n189 VTAIL.n188 185
R1500 VTAIL.n110 VTAIL.n109 185
R1501 VTAIL.n183 VTAIL.n182 185
R1502 VTAIL.n181 VTAIL.n112 185
R1503 VTAIL.n180 VTAIL.n179 185
R1504 VTAIL.n115 VTAIL.n113 185
R1505 VTAIL.n174 VTAIL.n173 185
R1506 VTAIL.n172 VTAIL.n171 185
R1507 VTAIL.n119 VTAIL.n118 185
R1508 VTAIL.n166 VTAIL.n165 185
R1509 VTAIL.n164 VTAIL.n163 185
R1510 VTAIL.n123 VTAIL.n122 185
R1511 VTAIL.n158 VTAIL.n157 185
R1512 VTAIL.n156 VTAIL.n155 185
R1513 VTAIL.n127 VTAIL.n126 185
R1514 VTAIL.n150 VTAIL.n149 185
R1515 VTAIL.n148 VTAIL.n147 185
R1516 VTAIL.n131 VTAIL.n130 185
R1517 VTAIL.n142 VTAIL.n141 185
R1518 VTAIL.n140 VTAIL.n139 185
R1519 VTAIL.n135 VTAIL.n134 185
R1520 VTAIL.n339 VTAIL.t0 147.659
R1521 VTAIL.n33 VTAIL.t2 147.659
R1522 VTAIL.n238 VTAIL.t3 147.659
R1523 VTAIL.n136 VTAIL.t1 147.659
R1524 VTAIL.n343 VTAIL.n337 104.615
R1525 VTAIL.n344 VTAIL.n343 104.615
R1526 VTAIL.n344 VTAIL.n333 104.615
R1527 VTAIL.n351 VTAIL.n333 104.615
R1528 VTAIL.n352 VTAIL.n351 104.615
R1529 VTAIL.n352 VTAIL.n329 104.615
R1530 VTAIL.n359 VTAIL.n329 104.615
R1531 VTAIL.n360 VTAIL.n359 104.615
R1532 VTAIL.n360 VTAIL.n325 104.615
R1533 VTAIL.n367 VTAIL.n325 104.615
R1534 VTAIL.n368 VTAIL.n367 104.615
R1535 VTAIL.n368 VTAIL.n321 104.615
R1536 VTAIL.n375 VTAIL.n321 104.615
R1537 VTAIL.n376 VTAIL.n375 104.615
R1538 VTAIL.n376 VTAIL.n317 104.615
R1539 VTAIL.n384 VTAIL.n317 104.615
R1540 VTAIL.n385 VTAIL.n384 104.615
R1541 VTAIL.n386 VTAIL.n385 104.615
R1542 VTAIL.n386 VTAIL.n313 104.615
R1543 VTAIL.n393 VTAIL.n313 104.615
R1544 VTAIL.n394 VTAIL.n393 104.615
R1545 VTAIL.n394 VTAIL.n309 104.615
R1546 VTAIL.n401 VTAIL.n309 104.615
R1547 VTAIL.n402 VTAIL.n401 104.615
R1548 VTAIL.n37 VTAIL.n31 104.615
R1549 VTAIL.n38 VTAIL.n37 104.615
R1550 VTAIL.n38 VTAIL.n27 104.615
R1551 VTAIL.n45 VTAIL.n27 104.615
R1552 VTAIL.n46 VTAIL.n45 104.615
R1553 VTAIL.n46 VTAIL.n23 104.615
R1554 VTAIL.n53 VTAIL.n23 104.615
R1555 VTAIL.n54 VTAIL.n53 104.615
R1556 VTAIL.n54 VTAIL.n19 104.615
R1557 VTAIL.n61 VTAIL.n19 104.615
R1558 VTAIL.n62 VTAIL.n61 104.615
R1559 VTAIL.n62 VTAIL.n15 104.615
R1560 VTAIL.n69 VTAIL.n15 104.615
R1561 VTAIL.n70 VTAIL.n69 104.615
R1562 VTAIL.n70 VTAIL.n11 104.615
R1563 VTAIL.n78 VTAIL.n11 104.615
R1564 VTAIL.n79 VTAIL.n78 104.615
R1565 VTAIL.n80 VTAIL.n79 104.615
R1566 VTAIL.n80 VTAIL.n7 104.615
R1567 VTAIL.n87 VTAIL.n7 104.615
R1568 VTAIL.n88 VTAIL.n87 104.615
R1569 VTAIL.n88 VTAIL.n3 104.615
R1570 VTAIL.n95 VTAIL.n3 104.615
R1571 VTAIL.n96 VTAIL.n95 104.615
R1572 VTAIL.n300 VTAIL.n299 104.615
R1573 VTAIL.n299 VTAIL.n207 104.615
R1574 VTAIL.n292 VTAIL.n207 104.615
R1575 VTAIL.n292 VTAIL.n291 104.615
R1576 VTAIL.n291 VTAIL.n211 104.615
R1577 VTAIL.n284 VTAIL.n211 104.615
R1578 VTAIL.n284 VTAIL.n283 104.615
R1579 VTAIL.n283 VTAIL.n282 104.615
R1580 VTAIL.n282 VTAIL.n215 104.615
R1581 VTAIL.n275 VTAIL.n215 104.615
R1582 VTAIL.n275 VTAIL.n274 104.615
R1583 VTAIL.n274 VTAIL.n220 104.615
R1584 VTAIL.n267 VTAIL.n220 104.615
R1585 VTAIL.n267 VTAIL.n266 104.615
R1586 VTAIL.n266 VTAIL.n224 104.615
R1587 VTAIL.n259 VTAIL.n224 104.615
R1588 VTAIL.n259 VTAIL.n258 104.615
R1589 VTAIL.n258 VTAIL.n228 104.615
R1590 VTAIL.n251 VTAIL.n228 104.615
R1591 VTAIL.n251 VTAIL.n250 104.615
R1592 VTAIL.n250 VTAIL.n232 104.615
R1593 VTAIL.n243 VTAIL.n232 104.615
R1594 VTAIL.n243 VTAIL.n242 104.615
R1595 VTAIL.n242 VTAIL.n236 104.615
R1596 VTAIL.n198 VTAIL.n197 104.615
R1597 VTAIL.n197 VTAIL.n105 104.615
R1598 VTAIL.n190 VTAIL.n105 104.615
R1599 VTAIL.n190 VTAIL.n189 104.615
R1600 VTAIL.n189 VTAIL.n109 104.615
R1601 VTAIL.n182 VTAIL.n109 104.615
R1602 VTAIL.n182 VTAIL.n181 104.615
R1603 VTAIL.n181 VTAIL.n180 104.615
R1604 VTAIL.n180 VTAIL.n113 104.615
R1605 VTAIL.n173 VTAIL.n113 104.615
R1606 VTAIL.n173 VTAIL.n172 104.615
R1607 VTAIL.n172 VTAIL.n118 104.615
R1608 VTAIL.n165 VTAIL.n118 104.615
R1609 VTAIL.n165 VTAIL.n164 104.615
R1610 VTAIL.n164 VTAIL.n122 104.615
R1611 VTAIL.n157 VTAIL.n122 104.615
R1612 VTAIL.n157 VTAIL.n156 104.615
R1613 VTAIL.n156 VTAIL.n126 104.615
R1614 VTAIL.n149 VTAIL.n126 104.615
R1615 VTAIL.n149 VTAIL.n148 104.615
R1616 VTAIL.n148 VTAIL.n130 104.615
R1617 VTAIL.n141 VTAIL.n130 104.615
R1618 VTAIL.n141 VTAIL.n140 104.615
R1619 VTAIL.n140 VTAIL.n134 104.615
R1620 VTAIL.t0 VTAIL.n337 52.3082
R1621 VTAIL.t2 VTAIL.n31 52.3082
R1622 VTAIL.t3 VTAIL.n236 52.3082
R1623 VTAIL.t1 VTAIL.n134 52.3082
R1624 VTAIL.n407 VTAIL.n406 31.6035
R1625 VTAIL.n101 VTAIL.n100 31.6035
R1626 VTAIL.n305 VTAIL.n304 31.6035
R1627 VTAIL.n203 VTAIL.n202 31.6035
R1628 VTAIL.n203 VTAIL.n101 31.2721
R1629 VTAIL.n407 VTAIL.n305 29.6686
R1630 VTAIL.n339 VTAIL.n338 15.6677
R1631 VTAIL.n33 VTAIL.n32 15.6677
R1632 VTAIL.n238 VTAIL.n237 15.6677
R1633 VTAIL.n136 VTAIL.n135 15.6677
R1634 VTAIL.n387 VTAIL.n316 13.1884
R1635 VTAIL.n81 VTAIL.n10 13.1884
R1636 VTAIL.n285 VTAIL.n214 13.1884
R1637 VTAIL.n183 VTAIL.n112 13.1884
R1638 VTAIL.n342 VTAIL.n341 12.8005
R1639 VTAIL.n383 VTAIL.n382 12.8005
R1640 VTAIL.n388 VTAIL.n314 12.8005
R1641 VTAIL.n36 VTAIL.n35 12.8005
R1642 VTAIL.n77 VTAIL.n76 12.8005
R1643 VTAIL.n82 VTAIL.n8 12.8005
R1644 VTAIL.n286 VTAIL.n212 12.8005
R1645 VTAIL.n281 VTAIL.n216 12.8005
R1646 VTAIL.n241 VTAIL.n240 12.8005
R1647 VTAIL.n184 VTAIL.n110 12.8005
R1648 VTAIL.n179 VTAIL.n114 12.8005
R1649 VTAIL.n139 VTAIL.n138 12.8005
R1650 VTAIL.n345 VTAIL.n336 12.0247
R1651 VTAIL.n381 VTAIL.n318 12.0247
R1652 VTAIL.n392 VTAIL.n391 12.0247
R1653 VTAIL.n39 VTAIL.n30 12.0247
R1654 VTAIL.n75 VTAIL.n12 12.0247
R1655 VTAIL.n86 VTAIL.n85 12.0247
R1656 VTAIL.n290 VTAIL.n289 12.0247
R1657 VTAIL.n280 VTAIL.n217 12.0247
R1658 VTAIL.n244 VTAIL.n235 12.0247
R1659 VTAIL.n188 VTAIL.n187 12.0247
R1660 VTAIL.n178 VTAIL.n115 12.0247
R1661 VTAIL.n142 VTAIL.n133 12.0247
R1662 VTAIL.n346 VTAIL.n334 11.249
R1663 VTAIL.n378 VTAIL.n377 11.249
R1664 VTAIL.n395 VTAIL.n312 11.249
R1665 VTAIL.n40 VTAIL.n28 11.249
R1666 VTAIL.n72 VTAIL.n71 11.249
R1667 VTAIL.n89 VTAIL.n6 11.249
R1668 VTAIL.n293 VTAIL.n210 11.249
R1669 VTAIL.n277 VTAIL.n276 11.249
R1670 VTAIL.n245 VTAIL.n233 11.249
R1671 VTAIL.n191 VTAIL.n108 11.249
R1672 VTAIL.n175 VTAIL.n174 11.249
R1673 VTAIL.n143 VTAIL.n131 11.249
R1674 VTAIL.n350 VTAIL.n349 10.4732
R1675 VTAIL.n374 VTAIL.n320 10.4732
R1676 VTAIL.n396 VTAIL.n310 10.4732
R1677 VTAIL.n44 VTAIL.n43 10.4732
R1678 VTAIL.n68 VTAIL.n14 10.4732
R1679 VTAIL.n90 VTAIL.n4 10.4732
R1680 VTAIL.n294 VTAIL.n208 10.4732
R1681 VTAIL.n273 VTAIL.n219 10.4732
R1682 VTAIL.n249 VTAIL.n248 10.4732
R1683 VTAIL.n192 VTAIL.n106 10.4732
R1684 VTAIL.n171 VTAIL.n117 10.4732
R1685 VTAIL.n147 VTAIL.n146 10.4732
R1686 VTAIL.n353 VTAIL.n332 9.69747
R1687 VTAIL.n373 VTAIL.n322 9.69747
R1688 VTAIL.n400 VTAIL.n399 9.69747
R1689 VTAIL.n47 VTAIL.n26 9.69747
R1690 VTAIL.n67 VTAIL.n16 9.69747
R1691 VTAIL.n94 VTAIL.n93 9.69747
R1692 VTAIL.n298 VTAIL.n297 9.69747
R1693 VTAIL.n272 VTAIL.n221 9.69747
R1694 VTAIL.n252 VTAIL.n231 9.69747
R1695 VTAIL.n196 VTAIL.n195 9.69747
R1696 VTAIL.n170 VTAIL.n119 9.69747
R1697 VTAIL.n150 VTAIL.n129 9.69747
R1698 VTAIL.n406 VTAIL.n405 9.45567
R1699 VTAIL.n100 VTAIL.n99 9.45567
R1700 VTAIL.n304 VTAIL.n303 9.45567
R1701 VTAIL.n202 VTAIL.n201 9.45567
R1702 VTAIL.n405 VTAIL.n404 9.3005
R1703 VTAIL.n308 VTAIL.n307 9.3005
R1704 VTAIL.n399 VTAIL.n398 9.3005
R1705 VTAIL.n397 VTAIL.n396 9.3005
R1706 VTAIL.n312 VTAIL.n311 9.3005
R1707 VTAIL.n391 VTAIL.n390 9.3005
R1708 VTAIL.n389 VTAIL.n388 9.3005
R1709 VTAIL.n328 VTAIL.n327 9.3005
R1710 VTAIL.n357 VTAIL.n356 9.3005
R1711 VTAIL.n355 VTAIL.n354 9.3005
R1712 VTAIL.n332 VTAIL.n331 9.3005
R1713 VTAIL.n349 VTAIL.n348 9.3005
R1714 VTAIL.n347 VTAIL.n346 9.3005
R1715 VTAIL.n336 VTAIL.n335 9.3005
R1716 VTAIL.n341 VTAIL.n340 9.3005
R1717 VTAIL.n363 VTAIL.n362 9.3005
R1718 VTAIL.n365 VTAIL.n364 9.3005
R1719 VTAIL.n324 VTAIL.n323 9.3005
R1720 VTAIL.n371 VTAIL.n370 9.3005
R1721 VTAIL.n373 VTAIL.n372 9.3005
R1722 VTAIL.n320 VTAIL.n319 9.3005
R1723 VTAIL.n379 VTAIL.n378 9.3005
R1724 VTAIL.n381 VTAIL.n380 9.3005
R1725 VTAIL.n382 VTAIL.n315 9.3005
R1726 VTAIL.n99 VTAIL.n98 9.3005
R1727 VTAIL.n2 VTAIL.n1 9.3005
R1728 VTAIL.n93 VTAIL.n92 9.3005
R1729 VTAIL.n91 VTAIL.n90 9.3005
R1730 VTAIL.n6 VTAIL.n5 9.3005
R1731 VTAIL.n85 VTAIL.n84 9.3005
R1732 VTAIL.n83 VTAIL.n82 9.3005
R1733 VTAIL.n22 VTAIL.n21 9.3005
R1734 VTAIL.n51 VTAIL.n50 9.3005
R1735 VTAIL.n49 VTAIL.n48 9.3005
R1736 VTAIL.n26 VTAIL.n25 9.3005
R1737 VTAIL.n43 VTAIL.n42 9.3005
R1738 VTAIL.n41 VTAIL.n40 9.3005
R1739 VTAIL.n30 VTAIL.n29 9.3005
R1740 VTAIL.n35 VTAIL.n34 9.3005
R1741 VTAIL.n57 VTAIL.n56 9.3005
R1742 VTAIL.n59 VTAIL.n58 9.3005
R1743 VTAIL.n18 VTAIL.n17 9.3005
R1744 VTAIL.n65 VTAIL.n64 9.3005
R1745 VTAIL.n67 VTAIL.n66 9.3005
R1746 VTAIL.n14 VTAIL.n13 9.3005
R1747 VTAIL.n73 VTAIL.n72 9.3005
R1748 VTAIL.n75 VTAIL.n74 9.3005
R1749 VTAIL.n76 VTAIL.n9 9.3005
R1750 VTAIL.n264 VTAIL.n263 9.3005
R1751 VTAIL.n223 VTAIL.n222 9.3005
R1752 VTAIL.n270 VTAIL.n269 9.3005
R1753 VTAIL.n272 VTAIL.n271 9.3005
R1754 VTAIL.n219 VTAIL.n218 9.3005
R1755 VTAIL.n278 VTAIL.n277 9.3005
R1756 VTAIL.n280 VTAIL.n279 9.3005
R1757 VTAIL.n216 VTAIL.n213 9.3005
R1758 VTAIL.n303 VTAIL.n302 9.3005
R1759 VTAIL.n206 VTAIL.n205 9.3005
R1760 VTAIL.n297 VTAIL.n296 9.3005
R1761 VTAIL.n295 VTAIL.n294 9.3005
R1762 VTAIL.n210 VTAIL.n209 9.3005
R1763 VTAIL.n289 VTAIL.n288 9.3005
R1764 VTAIL.n287 VTAIL.n286 9.3005
R1765 VTAIL.n262 VTAIL.n261 9.3005
R1766 VTAIL.n227 VTAIL.n226 9.3005
R1767 VTAIL.n256 VTAIL.n255 9.3005
R1768 VTAIL.n254 VTAIL.n253 9.3005
R1769 VTAIL.n231 VTAIL.n230 9.3005
R1770 VTAIL.n248 VTAIL.n247 9.3005
R1771 VTAIL.n246 VTAIL.n245 9.3005
R1772 VTAIL.n235 VTAIL.n234 9.3005
R1773 VTAIL.n240 VTAIL.n239 9.3005
R1774 VTAIL.n162 VTAIL.n161 9.3005
R1775 VTAIL.n121 VTAIL.n120 9.3005
R1776 VTAIL.n168 VTAIL.n167 9.3005
R1777 VTAIL.n170 VTAIL.n169 9.3005
R1778 VTAIL.n117 VTAIL.n116 9.3005
R1779 VTAIL.n176 VTAIL.n175 9.3005
R1780 VTAIL.n178 VTAIL.n177 9.3005
R1781 VTAIL.n114 VTAIL.n111 9.3005
R1782 VTAIL.n201 VTAIL.n200 9.3005
R1783 VTAIL.n104 VTAIL.n103 9.3005
R1784 VTAIL.n195 VTAIL.n194 9.3005
R1785 VTAIL.n193 VTAIL.n192 9.3005
R1786 VTAIL.n108 VTAIL.n107 9.3005
R1787 VTAIL.n187 VTAIL.n186 9.3005
R1788 VTAIL.n185 VTAIL.n184 9.3005
R1789 VTAIL.n160 VTAIL.n159 9.3005
R1790 VTAIL.n125 VTAIL.n124 9.3005
R1791 VTAIL.n154 VTAIL.n153 9.3005
R1792 VTAIL.n152 VTAIL.n151 9.3005
R1793 VTAIL.n129 VTAIL.n128 9.3005
R1794 VTAIL.n146 VTAIL.n145 9.3005
R1795 VTAIL.n144 VTAIL.n143 9.3005
R1796 VTAIL.n133 VTAIL.n132 9.3005
R1797 VTAIL.n138 VTAIL.n137 9.3005
R1798 VTAIL.n354 VTAIL.n330 8.92171
R1799 VTAIL.n370 VTAIL.n369 8.92171
R1800 VTAIL.n403 VTAIL.n308 8.92171
R1801 VTAIL.n48 VTAIL.n24 8.92171
R1802 VTAIL.n64 VTAIL.n63 8.92171
R1803 VTAIL.n97 VTAIL.n2 8.92171
R1804 VTAIL.n301 VTAIL.n206 8.92171
R1805 VTAIL.n269 VTAIL.n268 8.92171
R1806 VTAIL.n253 VTAIL.n229 8.92171
R1807 VTAIL.n199 VTAIL.n104 8.92171
R1808 VTAIL.n167 VTAIL.n166 8.92171
R1809 VTAIL.n151 VTAIL.n127 8.92171
R1810 VTAIL.n358 VTAIL.n357 8.14595
R1811 VTAIL.n366 VTAIL.n324 8.14595
R1812 VTAIL.n404 VTAIL.n306 8.14595
R1813 VTAIL.n52 VTAIL.n51 8.14595
R1814 VTAIL.n60 VTAIL.n18 8.14595
R1815 VTAIL.n98 VTAIL.n0 8.14595
R1816 VTAIL.n302 VTAIL.n204 8.14595
R1817 VTAIL.n265 VTAIL.n223 8.14595
R1818 VTAIL.n257 VTAIL.n256 8.14595
R1819 VTAIL.n200 VTAIL.n102 8.14595
R1820 VTAIL.n163 VTAIL.n121 8.14595
R1821 VTAIL.n155 VTAIL.n154 8.14595
R1822 VTAIL.n361 VTAIL.n328 7.3702
R1823 VTAIL.n365 VTAIL.n326 7.3702
R1824 VTAIL.n55 VTAIL.n22 7.3702
R1825 VTAIL.n59 VTAIL.n20 7.3702
R1826 VTAIL.n264 VTAIL.n225 7.3702
R1827 VTAIL.n260 VTAIL.n227 7.3702
R1828 VTAIL.n162 VTAIL.n123 7.3702
R1829 VTAIL.n158 VTAIL.n125 7.3702
R1830 VTAIL.n362 VTAIL.n361 6.59444
R1831 VTAIL.n362 VTAIL.n326 6.59444
R1832 VTAIL.n56 VTAIL.n55 6.59444
R1833 VTAIL.n56 VTAIL.n20 6.59444
R1834 VTAIL.n261 VTAIL.n225 6.59444
R1835 VTAIL.n261 VTAIL.n260 6.59444
R1836 VTAIL.n159 VTAIL.n123 6.59444
R1837 VTAIL.n159 VTAIL.n158 6.59444
R1838 VTAIL.n358 VTAIL.n328 5.81868
R1839 VTAIL.n366 VTAIL.n365 5.81868
R1840 VTAIL.n406 VTAIL.n306 5.81868
R1841 VTAIL.n52 VTAIL.n22 5.81868
R1842 VTAIL.n60 VTAIL.n59 5.81868
R1843 VTAIL.n100 VTAIL.n0 5.81868
R1844 VTAIL.n304 VTAIL.n204 5.81868
R1845 VTAIL.n265 VTAIL.n264 5.81868
R1846 VTAIL.n257 VTAIL.n227 5.81868
R1847 VTAIL.n202 VTAIL.n102 5.81868
R1848 VTAIL.n163 VTAIL.n162 5.81868
R1849 VTAIL.n155 VTAIL.n125 5.81868
R1850 VTAIL.n357 VTAIL.n330 5.04292
R1851 VTAIL.n369 VTAIL.n324 5.04292
R1852 VTAIL.n404 VTAIL.n403 5.04292
R1853 VTAIL.n51 VTAIL.n24 5.04292
R1854 VTAIL.n63 VTAIL.n18 5.04292
R1855 VTAIL.n98 VTAIL.n97 5.04292
R1856 VTAIL.n302 VTAIL.n301 5.04292
R1857 VTAIL.n268 VTAIL.n223 5.04292
R1858 VTAIL.n256 VTAIL.n229 5.04292
R1859 VTAIL.n200 VTAIL.n199 5.04292
R1860 VTAIL.n166 VTAIL.n121 5.04292
R1861 VTAIL.n154 VTAIL.n127 5.04292
R1862 VTAIL.n340 VTAIL.n339 4.38563
R1863 VTAIL.n34 VTAIL.n33 4.38563
R1864 VTAIL.n239 VTAIL.n238 4.38563
R1865 VTAIL.n137 VTAIL.n136 4.38563
R1866 VTAIL.n354 VTAIL.n353 4.26717
R1867 VTAIL.n370 VTAIL.n322 4.26717
R1868 VTAIL.n400 VTAIL.n308 4.26717
R1869 VTAIL.n48 VTAIL.n47 4.26717
R1870 VTAIL.n64 VTAIL.n16 4.26717
R1871 VTAIL.n94 VTAIL.n2 4.26717
R1872 VTAIL.n298 VTAIL.n206 4.26717
R1873 VTAIL.n269 VTAIL.n221 4.26717
R1874 VTAIL.n253 VTAIL.n252 4.26717
R1875 VTAIL.n196 VTAIL.n104 4.26717
R1876 VTAIL.n167 VTAIL.n119 4.26717
R1877 VTAIL.n151 VTAIL.n150 4.26717
R1878 VTAIL.n350 VTAIL.n332 3.49141
R1879 VTAIL.n374 VTAIL.n373 3.49141
R1880 VTAIL.n399 VTAIL.n310 3.49141
R1881 VTAIL.n44 VTAIL.n26 3.49141
R1882 VTAIL.n68 VTAIL.n67 3.49141
R1883 VTAIL.n93 VTAIL.n4 3.49141
R1884 VTAIL.n297 VTAIL.n208 3.49141
R1885 VTAIL.n273 VTAIL.n272 3.49141
R1886 VTAIL.n249 VTAIL.n231 3.49141
R1887 VTAIL.n195 VTAIL.n106 3.49141
R1888 VTAIL.n171 VTAIL.n170 3.49141
R1889 VTAIL.n147 VTAIL.n129 3.49141
R1890 VTAIL.n349 VTAIL.n334 2.71565
R1891 VTAIL.n377 VTAIL.n320 2.71565
R1892 VTAIL.n396 VTAIL.n395 2.71565
R1893 VTAIL.n43 VTAIL.n28 2.71565
R1894 VTAIL.n71 VTAIL.n14 2.71565
R1895 VTAIL.n90 VTAIL.n89 2.71565
R1896 VTAIL.n294 VTAIL.n293 2.71565
R1897 VTAIL.n276 VTAIL.n219 2.71565
R1898 VTAIL.n248 VTAIL.n233 2.71565
R1899 VTAIL.n192 VTAIL.n191 2.71565
R1900 VTAIL.n174 VTAIL.n117 2.71565
R1901 VTAIL.n146 VTAIL.n131 2.71565
R1902 VTAIL.n346 VTAIL.n345 1.93989
R1903 VTAIL.n378 VTAIL.n318 1.93989
R1904 VTAIL.n392 VTAIL.n312 1.93989
R1905 VTAIL.n40 VTAIL.n39 1.93989
R1906 VTAIL.n72 VTAIL.n12 1.93989
R1907 VTAIL.n86 VTAIL.n6 1.93989
R1908 VTAIL.n290 VTAIL.n210 1.93989
R1909 VTAIL.n277 VTAIL.n217 1.93989
R1910 VTAIL.n245 VTAIL.n244 1.93989
R1911 VTAIL.n188 VTAIL.n108 1.93989
R1912 VTAIL.n175 VTAIL.n115 1.93989
R1913 VTAIL.n143 VTAIL.n142 1.93989
R1914 VTAIL.n305 VTAIL.n203 1.27205
R1915 VTAIL.n342 VTAIL.n336 1.16414
R1916 VTAIL.n383 VTAIL.n381 1.16414
R1917 VTAIL.n391 VTAIL.n314 1.16414
R1918 VTAIL.n36 VTAIL.n30 1.16414
R1919 VTAIL.n77 VTAIL.n75 1.16414
R1920 VTAIL.n85 VTAIL.n8 1.16414
R1921 VTAIL.n289 VTAIL.n212 1.16414
R1922 VTAIL.n281 VTAIL.n280 1.16414
R1923 VTAIL.n241 VTAIL.n235 1.16414
R1924 VTAIL.n187 VTAIL.n110 1.16414
R1925 VTAIL.n179 VTAIL.n178 1.16414
R1926 VTAIL.n139 VTAIL.n133 1.16414
R1927 VTAIL VTAIL.n101 0.929379
R1928 VTAIL.n341 VTAIL.n338 0.388379
R1929 VTAIL.n382 VTAIL.n316 0.388379
R1930 VTAIL.n388 VTAIL.n387 0.388379
R1931 VTAIL.n35 VTAIL.n32 0.388379
R1932 VTAIL.n76 VTAIL.n10 0.388379
R1933 VTAIL.n82 VTAIL.n81 0.388379
R1934 VTAIL.n286 VTAIL.n285 0.388379
R1935 VTAIL.n216 VTAIL.n214 0.388379
R1936 VTAIL.n240 VTAIL.n237 0.388379
R1937 VTAIL.n184 VTAIL.n183 0.388379
R1938 VTAIL.n114 VTAIL.n112 0.388379
R1939 VTAIL.n138 VTAIL.n135 0.388379
R1940 VTAIL VTAIL.n407 0.343172
R1941 VTAIL.n340 VTAIL.n335 0.155672
R1942 VTAIL.n347 VTAIL.n335 0.155672
R1943 VTAIL.n348 VTAIL.n347 0.155672
R1944 VTAIL.n348 VTAIL.n331 0.155672
R1945 VTAIL.n355 VTAIL.n331 0.155672
R1946 VTAIL.n356 VTAIL.n355 0.155672
R1947 VTAIL.n356 VTAIL.n327 0.155672
R1948 VTAIL.n363 VTAIL.n327 0.155672
R1949 VTAIL.n364 VTAIL.n363 0.155672
R1950 VTAIL.n364 VTAIL.n323 0.155672
R1951 VTAIL.n371 VTAIL.n323 0.155672
R1952 VTAIL.n372 VTAIL.n371 0.155672
R1953 VTAIL.n372 VTAIL.n319 0.155672
R1954 VTAIL.n379 VTAIL.n319 0.155672
R1955 VTAIL.n380 VTAIL.n379 0.155672
R1956 VTAIL.n380 VTAIL.n315 0.155672
R1957 VTAIL.n389 VTAIL.n315 0.155672
R1958 VTAIL.n390 VTAIL.n389 0.155672
R1959 VTAIL.n390 VTAIL.n311 0.155672
R1960 VTAIL.n397 VTAIL.n311 0.155672
R1961 VTAIL.n398 VTAIL.n397 0.155672
R1962 VTAIL.n398 VTAIL.n307 0.155672
R1963 VTAIL.n405 VTAIL.n307 0.155672
R1964 VTAIL.n34 VTAIL.n29 0.155672
R1965 VTAIL.n41 VTAIL.n29 0.155672
R1966 VTAIL.n42 VTAIL.n41 0.155672
R1967 VTAIL.n42 VTAIL.n25 0.155672
R1968 VTAIL.n49 VTAIL.n25 0.155672
R1969 VTAIL.n50 VTAIL.n49 0.155672
R1970 VTAIL.n50 VTAIL.n21 0.155672
R1971 VTAIL.n57 VTAIL.n21 0.155672
R1972 VTAIL.n58 VTAIL.n57 0.155672
R1973 VTAIL.n58 VTAIL.n17 0.155672
R1974 VTAIL.n65 VTAIL.n17 0.155672
R1975 VTAIL.n66 VTAIL.n65 0.155672
R1976 VTAIL.n66 VTAIL.n13 0.155672
R1977 VTAIL.n73 VTAIL.n13 0.155672
R1978 VTAIL.n74 VTAIL.n73 0.155672
R1979 VTAIL.n74 VTAIL.n9 0.155672
R1980 VTAIL.n83 VTAIL.n9 0.155672
R1981 VTAIL.n84 VTAIL.n83 0.155672
R1982 VTAIL.n84 VTAIL.n5 0.155672
R1983 VTAIL.n91 VTAIL.n5 0.155672
R1984 VTAIL.n92 VTAIL.n91 0.155672
R1985 VTAIL.n92 VTAIL.n1 0.155672
R1986 VTAIL.n99 VTAIL.n1 0.155672
R1987 VTAIL.n303 VTAIL.n205 0.155672
R1988 VTAIL.n296 VTAIL.n205 0.155672
R1989 VTAIL.n296 VTAIL.n295 0.155672
R1990 VTAIL.n295 VTAIL.n209 0.155672
R1991 VTAIL.n288 VTAIL.n209 0.155672
R1992 VTAIL.n288 VTAIL.n287 0.155672
R1993 VTAIL.n287 VTAIL.n213 0.155672
R1994 VTAIL.n279 VTAIL.n213 0.155672
R1995 VTAIL.n279 VTAIL.n278 0.155672
R1996 VTAIL.n278 VTAIL.n218 0.155672
R1997 VTAIL.n271 VTAIL.n218 0.155672
R1998 VTAIL.n271 VTAIL.n270 0.155672
R1999 VTAIL.n270 VTAIL.n222 0.155672
R2000 VTAIL.n263 VTAIL.n222 0.155672
R2001 VTAIL.n263 VTAIL.n262 0.155672
R2002 VTAIL.n262 VTAIL.n226 0.155672
R2003 VTAIL.n255 VTAIL.n226 0.155672
R2004 VTAIL.n255 VTAIL.n254 0.155672
R2005 VTAIL.n254 VTAIL.n230 0.155672
R2006 VTAIL.n247 VTAIL.n230 0.155672
R2007 VTAIL.n247 VTAIL.n246 0.155672
R2008 VTAIL.n246 VTAIL.n234 0.155672
R2009 VTAIL.n239 VTAIL.n234 0.155672
R2010 VTAIL.n201 VTAIL.n103 0.155672
R2011 VTAIL.n194 VTAIL.n103 0.155672
R2012 VTAIL.n194 VTAIL.n193 0.155672
R2013 VTAIL.n193 VTAIL.n107 0.155672
R2014 VTAIL.n186 VTAIL.n107 0.155672
R2015 VTAIL.n186 VTAIL.n185 0.155672
R2016 VTAIL.n185 VTAIL.n111 0.155672
R2017 VTAIL.n177 VTAIL.n111 0.155672
R2018 VTAIL.n177 VTAIL.n176 0.155672
R2019 VTAIL.n176 VTAIL.n116 0.155672
R2020 VTAIL.n169 VTAIL.n116 0.155672
R2021 VTAIL.n169 VTAIL.n168 0.155672
R2022 VTAIL.n168 VTAIL.n120 0.155672
R2023 VTAIL.n161 VTAIL.n120 0.155672
R2024 VTAIL.n161 VTAIL.n160 0.155672
R2025 VTAIL.n160 VTAIL.n124 0.155672
R2026 VTAIL.n153 VTAIL.n124 0.155672
R2027 VTAIL.n153 VTAIL.n152 0.155672
R2028 VTAIL.n152 VTAIL.n128 0.155672
R2029 VTAIL.n145 VTAIL.n128 0.155672
R2030 VTAIL.n145 VTAIL.n144 0.155672
R2031 VTAIL.n144 VTAIL.n132 0.155672
R2032 VTAIL.n137 VTAIL.n132 0.155672
R2033 VDD1.n96 VDD1.n0 289.615
R2034 VDD1.n197 VDD1.n101 289.615
R2035 VDD1.n97 VDD1.n96 185
R2036 VDD1.n95 VDD1.n94 185
R2037 VDD1.n4 VDD1.n3 185
R2038 VDD1.n89 VDD1.n88 185
R2039 VDD1.n87 VDD1.n86 185
R2040 VDD1.n8 VDD1.n7 185
R2041 VDD1.n81 VDD1.n80 185
R2042 VDD1.n79 VDD1.n10 185
R2043 VDD1.n78 VDD1.n77 185
R2044 VDD1.n13 VDD1.n11 185
R2045 VDD1.n72 VDD1.n71 185
R2046 VDD1.n70 VDD1.n69 185
R2047 VDD1.n17 VDD1.n16 185
R2048 VDD1.n64 VDD1.n63 185
R2049 VDD1.n62 VDD1.n61 185
R2050 VDD1.n21 VDD1.n20 185
R2051 VDD1.n56 VDD1.n55 185
R2052 VDD1.n54 VDD1.n53 185
R2053 VDD1.n25 VDD1.n24 185
R2054 VDD1.n48 VDD1.n47 185
R2055 VDD1.n46 VDD1.n45 185
R2056 VDD1.n29 VDD1.n28 185
R2057 VDD1.n40 VDD1.n39 185
R2058 VDD1.n38 VDD1.n37 185
R2059 VDD1.n33 VDD1.n32 185
R2060 VDD1.n133 VDD1.n132 185
R2061 VDD1.n138 VDD1.n137 185
R2062 VDD1.n140 VDD1.n139 185
R2063 VDD1.n129 VDD1.n128 185
R2064 VDD1.n146 VDD1.n145 185
R2065 VDD1.n148 VDD1.n147 185
R2066 VDD1.n125 VDD1.n124 185
R2067 VDD1.n154 VDD1.n153 185
R2068 VDD1.n156 VDD1.n155 185
R2069 VDD1.n121 VDD1.n120 185
R2070 VDD1.n162 VDD1.n161 185
R2071 VDD1.n164 VDD1.n163 185
R2072 VDD1.n117 VDD1.n116 185
R2073 VDD1.n170 VDD1.n169 185
R2074 VDD1.n172 VDD1.n171 185
R2075 VDD1.n113 VDD1.n112 185
R2076 VDD1.n179 VDD1.n178 185
R2077 VDD1.n180 VDD1.n111 185
R2078 VDD1.n182 VDD1.n181 185
R2079 VDD1.n109 VDD1.n108 185
R2080 VDD1.n188 VDD1.n187 185
R2081 VDD1.n190 VDD1.n189 185
R2082 VDD1.n105 VDD1.n104 185
R2083 VDD1.n196 VDD1.n195 185
R2084 VDD1.n198 VDD1.n197 185
R2085 VDD1.n34 VDD1.t0 147.659
R2086 VDD1.n134 VDD1.t1 147.659
R2087 VDD1.n96 VDD1.n95 104.615
R2088 VDD1.n95 VDD1.n3 104.615
R2089 VDD1.n88 VDD1.n3 104.615
R2090 VDD1.n88 VDD1.n87 104.615
R2091 VDD1.n87 VDD1.n7 104.615
R2092 VDD1.n80 VDD1.n7 104.615
R2093 VDD1.n80 VDD1.n79 104.615
R2094 VDD1.n79 VDD1.n78 104.615
R2095 VDD1.n78 VDD1.n11 104.615
R2096 VDD1.n71 VDD1.n11 104.615
R2097 VDD1.n71 VDD1.n70 104.615
R2098 VDD1.n70 VDD1.n16 104.615
R2099 VDD1.n63 VDD1.n16 104.615
R2100 VDD1.n63 VDD1.n62 104.615
R2101 VDD1.n62 VDD1.n20 104.615
R2102 VDD1.n55 VDD1.n20 104.615
R2103 VDD1.n55 VDD1.n54 104.615
R2104 VDD1.n54 VDD1.n24 104.615
R2105 VDD1.n47 VDD1.n24 104.615
R2106 VDD1.n47 VDD1.n46 104.615
R2107 VDD1.n46 VDD1.n28 104.615
R2108 VDD1.n39 VDD1.n28 104.615
R2109 VDD1.n39 VDD1.n38 104.615
R2110 VDD1.n38 VDD1.n32 104.615
R2111 VDD1.n138 VDD1.n132 104.615
R2112 VDD1.n139 VDD1.n138 104.615
R2113 VDD1.n139 VDD1.n128 104.615
R2114 VDD1.n146 VDD1.n128 104.615
R2115 VDD1.n147 VDD1.n146 104.615
R2116 VDD1.n147 VDD1.n124 104.615
R2117 VDD1.n154 VDD1.n124 104.615
R2118 VDD1.n155 VDD1.n154 104.615
R2119 VDD1.n155 VDD1.n120 104.615
R2120 VDD1.n162 VDD1.n120 104.615
R2121 VDD1.n163 VDD1.n162 104.615
R2122 VDD1.n163 VDD1.n116 104.615
R2123 VDD1.n170 VDD1.n116 104.615
R2124 VDD1.n171 VDD1.n170 104.615
R2125 VDD1.n171 VDD1.n112 104.615
R2126 VDD1.n179 VDD1.n112 104.615
R2127 VDD1.n180 VDD1.n179 104.615
R2128 VDD1.n181 VDD1.n180 104.615
R2129 VDD1.n181 VDD1.n108 104.615
R2130 VDD1.n188 VDD1.n108 104.615
R2131 VDD1.n189 VDD1.n188 104.615
R2132 VDD1.n189 VDD1.n104 104.615
R2133 VDD1.n196 VDD1.n104 104.615
R2134 VDD1.n197 VDD1.n196 104.615
R2135 VDD1 VDD1.n201 91.7726
R2136 VDD1.t0 VDD1.n32 52.3082
R2137 VDD1.t1 VDD1.n132 52.3082
R2138 VDD1 VDD1.n100 48.7414
R2139 VDD1.n34 VDD1.n33 15.6677
R2140 VDD1.n134 VDD1.n133 15.6677
R2141 VDD1.n81 VDD1.n10 13.1884
R2142 VDD1.n182 VDD1.n111 13.1884
R2143 VDD1.n82 VDD1.n8 12.8005
R2144 VDD1.n77 VDD1.n12 12.8005
R2145 VDD1.n37 VDD1.n36 12.8005
R2146 VDD1.n137 VDD1.n136 12.8005
R2147 VDD1.n178 VDD1.n177 12.8005
R2148 VDD1.n183 VDD1.n109 12.8005
R2149 VDD1.n86 VDD1.n85 12.0247
R2150 VDD1.n76 VDD1.n13 12.0247
R2151 VDD1.n40 VDD1.n31 12.0247
R2152 VDD1.n140 VDD1.n131 12.0247
R2153 VDD1.n176 VDD1.n113 12.0247
R2154 VDD1.n187 VDD1.n186 12.0247
R2155 VDD1.n89 VDD1.n6 11.249
R2156 VDD1.n73 VDD1.n72 11.249
R2157 VDD1.n41 VDD1.n29 11.249
R2158 VDD1.n141 VDD1.n129 11.249
R2159 VDD1.n173 VDD1.n172 11.249
R2160 VDD1.n190 VDD1.n107 11.249
R2161 VDD1.n90 VDD1.n4 10.4732
R2162 VDD1.n69 VDD1.n15 10.4732
R2163 VDD1.n45 VDD1.n44 10.4732
R2164 VDD1.n145 VDD1.n144 10.4732
R2165 VDD1.n169 VDD1.n115 10.4732
R2166 VDD1.n191 VDD1.n105 10.4732
R2167 VDD1.n94 VDD1.n93 9.69747
R2168 VDD1.n68 VDD1.n17 9.69747
R2169 VDD1.n48 VDD1.n27 9.69747
R2170 VDD1.n148 VDD1.n127 9.69747
R2171 VDD1.n168 VDD1.n117 9.69747
R2172 VDD1.n195 VDD1.n194 9.69747
R2173 VDD1.n100 VDD1.n99 9.45567
R2174 VDD1.n201 VDD1.n200 9.45567
R2175 VDD1.n60 VDD1.n59 9.3005
R2176 VDD1.n19 VDD1.n18 9.3005
R2177 VDD1.n66 VDD1.n65 9.3005
R2178 VDD1.n68 VDD1.n67 9.3005
R2179 VDD1.n15 VDD1.n14 9.3005
R2180 VDD1.n74 VDD1.n73 9.3005
R2181 VDD1.n76 VDD1.n75 9.3005
R2182 VDD1.n12 VDD1.n9 9.3005
R2183 VDD1.n99 VDD1.n98 9.3005
R2184 VDD1.n2 VDD1.n1 9.3005
R2185 VDD1.n93 VDD1.n92 9.3005
R2186 VDD1.n91 VDD1.n90 9.3005
R2187 VDD1.n6 VDD1.n5 9.3005
R2188 VDD1.n85 VDD1.n84 9.3005
R2189 VDD1.n83 VDD1.n82 9.3005
R2190 VDD1.n58 VDD1.n57 9.3005
R2191 VDD1.n23 VDD1.n22 9.3005
R2192 VDD1.n52 VDD1.n51 9.3005
R2193 VDD1.n50 VDD1.n49 9.3005
R2194 VDD1.n27 VDD1.n26 9.3005
R2195 VDD1.n44 VDD1.n43 9.3005
R2196 VDD1.n42 VDD1.n41 9.3005
R2197 VDD1.n31 VDD1.n30 9.3005
R2198 VDD1.n36 VDD1.n35 9.3005
R2199 VDD1.n200 VDD1.n199 9.3005
R2200 VDD1.n103 VDD1.n102 9.3005
R2201 VDD1.n194 VDD1.n193 9.3005
R2202 VDD1.n192 VDD1.n191 9.3005
R2203 VDD1.n107 VDD1.n106 9.3005
R2204 VDD1.n186 VDD1.n185 9.3005
R2205 VDD1.n184 VDD1.n183 9.3005
R2206 VDD1.n123 VDD1.n122 9.3005
R2207 VDD1.n152 VDD1.n151 9.3005
R2208 VDD1.n150 VDD1.n149 9.3005
R2209 VDD1.n127 VDD1.n126 9.3005
R2210 VDD1.n144 VDD1.n143 9.3005
R2211 VDD1.n142 VDD1.n141 9.3005
R2212 VDD1.n131 VDD1.n130 9.3005
R2213 VDD1.n136 VDD1.n135 9.3005
R2214 VDD1.n158 VDD1.n157 9.3005
R2215 VDD1.n160 VDD1.n159 9.3005
R2216 VDD1.n119 VDD1.n118 9.3005
R2217 VDD1.n166 VDD1.n165 9.3005
R2218 VDD1.n168 VDD1.n167 9.3005
R2219 VDD1.n115 VDD1.n114 9.3005
R2220 VDD1.n174 VDD1.n173 9.3005
R2221 VDD1.n176 VDD1.n175 9.3005
R2222 VDD1.n177 VDD1.n110 9.3005
R2223 VDD1.n97 VDD1.n2 8.92171
R2224 VDD1.n65 VDD1.n64 8.92171
R2225 VDD1.n49 VDD1.n25 8.92171
R2226 VDD1.n149 VDD1.n125 8.92171
R2227 VDD1.n165 VDD1.n164 8.92171
R2228 VDD1.n198 VDD1.n103 8.92171
R2229 VDD1.n98 VDD1.n0 8.14595
R2230 VDD1.n61 VDD1.n19 8.14595
R2231 VDD1.n53 VDD1.n52 8.14595
R2232 VDD1.n153 VDD1.n152 8.14595
R2233 VDD1.n161 VDD1.n119 8.14595
R2234 VDD1.n199 VDD1.n101 8.14595
R2235 VDD1.n60 VDD1.n21 7.3702
R2236 VDD1.n56 VDD1.n23 7.3702
R2237 VDD1.n156 VDD1.n123 7.3702
R2238 VDD1.n160 VDD1.n121 7.3702
R2239 VDD1.n57 VDD1.n21 6.59444
R2240 VDD1.n57 VDD1.n56 6.59444
R2241 VDD1.n157 VDD1.n156 6.59444
R2242 VDD1.n157 VDD1.n121 6.59444
R2243 VDD1.n100 VDD1.n0 5.81868
R2244 VDD1.n61 VDD1.n60 5.81868
R2245 VDD1.n53 VDD1.n23 5.81868
R2246 VDD1.n153 VDD1.n123 5.81868
R2247 VDD1.n161 VDD1.n160 5.81868
R2248 VDD1.n201 VDD1.n101 5.81868
R2249 VDD1.n98 VDD1.n97 5.04292
R2250 VDD1.n64 VDD1.n19 5.04292
R2251 VDD1.n52 VDD1.n25 5.04292
R2252 VDD1.n152 VDD1.n125 5.04292
R2253 VDD1.n164 VDD1.n119 5.04292
R2254 VDD1.n199 VDD1.n198 5.04292
R2255 VDD1.n35 VDD1.n34 4.38563
R2256 VDD1.n135 VDD1.n134 4.38563
R2257 VDD1.n94 VDD1.n2 4.26717
R2258 VDD1.n65 VDD1.n17 4.26717
R2259 VDD1.n49 VDD1.n48 4.26717
R2260 VDD1.n149 VDD1.n148 4.26717
R2261 VDD1.n165 VDD1.n117 4.26717
R2262 VDD1.n195 VDD1.n103 4.26717
R2263 VDD1.n93 VDD1.n4 3.49141
R2264 VDD1.n69 VDD1.n68 3.49141
R2265 VDD1.n45 VDD1.n27 3.49141
R2266 VDD1.n145 VDD1.n127 3.49141
R2267 VDD1.n169 VDD1.n168 3.49141
R2268 VDD1.n194 VDD1.n105 3.49141
R2269 VDD1.n90 VDD1.n89 2.71565
R2270 VDD1.n72 VDD1.n15 2.71565
R2271 VDD1.n44 VDD1.n29 2.71565
R2272 VDD1.n144 VDD1.n129 2.71565
R2273 VDD1.n172 VDD1.n115 2.71565
R2274 VDD1.n191 VDD1.n190 2.71565
R2275 VDD1.n86 VDD1.n6 1.93989
R2276 VDD1.n73 VDD1.n13 1.93989
R2277 VDD1.n41 VDD1.n40 1.93989
R2278 VDD1.n141 VDD1.n140 1.93989
R2279 VDD1.n173 VDD1.n113 1.93989
R2280 VDD1.n187 VDD1.n107 1.93989
R2281 VDD1.n85 VDD1.n8 1.16414
R2282 VDD1.n77 VDD1.n76 1.16414
R2283 VDD1.n37 VDD1.n31 1.16414
R2284 VDD1.n137 VDD1.n131 1.16414
R2285 VDD1.n178 VDD1.n176 1.16414
R2286 VDD1.n186 VDD1.n109 1.16414
R2287 VDD1.n82 VDD1.n81 0.388379
R2288 VDD1.n12 VDD1.n10 0.388379
R2289 VDD1.n36 VDD1.n33 0.388379
R2290 VDD1.n136 VDD1.n133 0.388379
R2291 VDD1.n177 VDD1.n111 0.388379
R2292 VDD1.n183 VDD1.n182 0.388379
R2293 VDD1.n99 VDD1.n1 0.155672
R2294 VDD1.n92 VDD1.n1 0.155672
R2295 VDD1.n92 VDD1.n91 0.155672
R2296 VDD1.n91 VDD1.n5 0.155672
R2297 VDD1.n84 VDD1.n5 0.155672
R2298 VDD1.n84 VDD1.n83 0.155672
R2299 VDD1.n83 VDD1.n9 0.155672
R2300 VDD1.n75 VDD1.n9 0.155672
R2301 VDD1.n75 VDD1.n74 0.155672
R2302 VDD1.n74 VDD1.n14 0.155672
R2303 VDD1.n67 VDD1.n14 0.155672
R2304 VDD1.n67 VDD1.n66 0.155672
R2305 VDD1.n66 VDD1.n18 0.155672
R2306 VDD1.n59 VDD1.n18 0.155672
R2307 VDD1.n59 VDD1.n58 0.155672
R2308 VDD1.n58 VDD1.n22 0.155672
R2309 VDD1.n51 VDD1.n22 0.155672
R2310 VDD1.n51 VDD1.n50 0.155672
R2311 VDD1.n50 VDD1.n26 0.155672
R2312 VDD1.n43 VDD1.n26 0.155672
R2313 VDD1.n43 VDD1.n42 0.155672
R2314 VDD1.n42 VDD1.n30 0.155672
R2315 VDD1.n35 VDD1.n30 0.155672
R2316 VDD1.n135 VDD1.n130 0.155672
R2317 VDD1.n142 VDD1.n130 0.155672
R2318 VDD1.n143 VDD1.n142 0.155672
R2319 VDD1.n143 VDD1.n126 0.155672
R2320 VDD1.n150 VDD1.n126 0.155672
R2321 VDD1.n151 VDD1.n150 0.155672
R2322 VDD1.n151 VDD1.n122 0.155672
R2323 VDD1.n158 VDD1.n122 0.155672
R2324 VDD1.n159 VDD1.n158 0.155672
R2325 VDD1.n159 VDD1.n118 0.155672
R2326 VDD1.n166 VDD1.n118 0.155672
R2327 VDD1.n167 VDD1.n166 0.155672
R2328 VDD1.n167 VDD1.n114 0.155672
R2329 VDD1.n174 VDD1.n114 0.155672
R2330 VDD1.n175 VDD1.n174 0.155672
R2331 VDD1.n175 VDD1.n110 0.155672
R2332 VDD1.n184 VDD1.n110 0.155672
R2333 VDD1.n185 VDD1.n184 0.155672
R2334 VDD1.n185 VDD1.n106 0.155672
R2335 VDD1.n192 VDD1.n106 0.155672
R2336 VDD1.n193 VDD1.n192 0.155672
R2337 VDD1.n193 VDD1.n102 0.155672
R2338 VDD1.n200 VDD1.n102 0.155672
R2339 VN VN.t0 440.082
R2340 VN VN.t1 393.42
R2341 VDD2.n197 VDD2.n101 289.615
R2342 VDD2.n96 VDD2.n0 289.615
R2343 VDD2.n198 VDD2.n197 185
R2344 VDD2.n196 VDD2.n195 185
R2345 VDD2.n105 VDD2.n104 185
R2346 VDD2.n190 VDD2.n189 185
R2347 VDD2.n188 VDD2.n187 185
R2348 VDD2.n109 VDD2.n108 185
R2349 VDD2.n182 VDD2.n181 185
R2350 VDD2.n180 VDD2.n111 185
R2351 VDD2.n179 VDD2.n178 185
R2352 VDD2.n114 VDD2.n112 185
R2353 VDD2.n173 VDD2.n172 185
R2354 VDD2.n171 VDD2.n170 185
R2355 VDD2.n118 VDD2.n117 185
R2356 VDD2.n165 VDD2.n164 185
R2357 VDD2.n163 VDD2.n162 185
R2358 VDD2.n122 VDD2.n121 185
R2359 VDD2.n157 VDD2.n156 185
R2360 VDD2.n155 VDD2.n154 185
R2361 VDD2.n126 VDD2.n125 185
R2362 VDD2.n149 VDD2.n148 185
R2363 VDD2.n147 VDD2.n146 185
R2364 VDD2.n130 VDD2.n129 185
R2365 VDD2.n141 VDD2.n140 185
R2366 VDD2.n139 VDD2.n138 185
R2367 VDD2.n134 VDD2.n133 185
R2368 VDD2.n32 VDD2.n31 185
R2369 VDD2.n37 VDD2.n36 185
R2370 VDD2.n39 VDD2.n38 185
R2371 VDD2.n28 VDD2.n27 185
R2372 VDD2.n45 VDD2.n44 185
R2373 VDD2.n47 VDD2.n46 185
R2374 VDD2.n24 VDD2.n23 185
R2375 VDD2.n53 VDD2.n52 185
R2376 VDD2.n55 VDD2.n54 185
R2377 VDD2.n20 VDD2.n19 185
R2378 VDD2.n61 VDD2.n60 185
R2379 VDD2.n63 VDD2.n62 185
R2380 VDD2.n16 VDD2.n15 185
R2381 VDD2.n69 VDD2.n68 185
R2382 VDD2.n71 VDD2.n70 185
R2383 VDD2.n12 VDD2.n11 185
R2384 VDD2.n78 VDD2.n77 185
R2385 VDD2.n79 VDD2.n10 185
R2386 VDD2.n81 VDD2.n80 185
R2387 VDD2.n8 VDD2.n7 185
R2388 VDD2.n87 VDD2.n86 185
R2389 VDD2.n89 VDD2.n88 185
R2390 VDD2.n4 VDD2.n3 185
R2391 VDD2.n95 VDD2.n94 185
R2392 VDD2.n97 VDD2.n96 185
R2393 VDD2.n135 VDD2.t1 147.659
R2394 VDD2.n33 VDD2.t0 147.659
R2395 VDD2.n197 VDD2.n196 104.615
R2396 VDD2.n196 VDD2.n104 104.615
R2397 VDD2.n189 VDD2.n104 104.615
R2398 VDD2.n189 VDD2.n188 104.615
R2399 VDD2.n188 VDD2.n108 104.615
R2400 VDD2.n181 VDD2.n108 104.615
R2401 VDD2.n181 VDD2.n180 104.615
R2402 VDD2.n180 VDD2.n179 104.615
R2403 VDD2.n179 VDD2.n112 104.615
R2404 VDD2.n172 VDD2.n112 104.615
R2405 VDD2.n172 VDD2.n171 104.615
R2406 VDD2.n171 VDD2.n117 104.615
R2407 VDD2.n164 VDD2.n117 104.615
R2408 VDD2.n164 VDD2.n163 104.615
R2409 VDD2.n163 VDD2.n121 104.615
R2410 VDD2.n156 VDD2.n121 104.615
R2411 VDD2.n156 VDD2.n155 104.615
R2412 VDD2.n155 VDD2.n125 104.615
R2413 VDD2.n148 VDD2.n125 104.615
R2414 VDD2.n148 VDD2.n147 104.615
R2415 VDD2.n147 VDD2.n129 104.615
R2416 VDD2.n140 VDD2.n129 104.615
R2417 VDD2.n140 VDD2.n139 104.615
R2418 VDD2.n139 VDD2.n133 104.615
R2419 VDD2.n37 VDD2.n31 104.615
R2420 VDD2.n38 VDD2.n37 104.615
R2421 VDD2.n38 VDD2.n27 104.615
R2422 VDD2.n45 VDD2.n27 104.615
R2423 VDD2.n46 VDD2.n45 104.615
R2424 VDD2.n46 VDD2.n23 104.615
R2425 VDD2.n53 VDD2.n23 104.615
R2426 VDD2.n54 VDD2.n53 104.615
R2427 VDD2.n54 VDD2.n19 104.615
R2428 VDD2.n61 VDD2.n19 104.615
R2429 VDD2.n62 VDD2.n61 104.615
R2430 VDD2.n62 VDD2.n15 104.615
R2431 VDD2.n69 VDD2.n15 104.615
R2432 VDD2.n70 VDD2.n69 104.615
R2433 VDD2.n70 VDD2.n11 104.615
R2434 VDD2.n78 VDD2.n11 104.615
R2435 VDD2.n79 VDD2.n78 104.615
R2436 VDD2.n80 VDD2.n79 104.615
R2437 VDD2.n80 VDD2.n7 104.615
R2438 VDD2.n87 VDD2.n7 104.615
R2439 VDD2.n88 VDD2.n87 104.615
R2440 VDD2.n88 VDD2.n3 104.615
R2441 VDD2.n95 VDD2.n3 104.615
R2442 VDD2.n96 VDD2.n95 104.615
R2443 VDD2.n202 VDD2.n100 90.8469
R2444 VDD2.t1 VDD2.n133 52.3082
R2445 VDD2.t0 VDD2.n31 52.3082
R2446 VDD2.n202 VDD2.n201 48.2823
R2447 VDD2.n135 VDD2.n134 15.6677
R2448 VDD2.n33 VDD2.n32 15.6677
R2449 VDD2.n182 VDD2.n111 13.1884
R2450 VDD2.n81 VDD2.n10 13.1884
R2451 VDD2.n183 VDD2.n109 12.8005
R2452 VDD2.n178 VDD2.n113 12.8005
R2453 VDD2.n138 VDD2.n137 12.8005
R2454 VDD2.n36 VDD2.n35 12.8005
R2455 VDD2.n77 VDD2.n76 12.8005
R2456 VDD2.n82 VDD2.n8 12.8005
R2457 VDD2.n187 VDD2.n186 12.0247
R2458 VDD2.n177 VDD2.n114 12.0247
R2459 VDD2.n141 VDD2.n132 12.0247
R2460 VDD2.n39 VDD2.n30 12.0247
R2461 VDD2.n75 VDD2.n12 12.0247
R2462 VDD2.n86 VDD2.n85 12.0247
R2463 VDD2.n190 VDD2.n107 11.249
R2464 VDD2.n174 VDD2.n173 11.249
R2465 VDD2.n142 VDD2.n130 11.249
R2466 VDD2.n40 VDD2.n28 11.249
R2467 VDD2.n72 VDD2.n71 11.249
R2468 VDD2.n89 VDD2.n6 11.249
R2469 VDD2.n191 VDD2.n105 10.4732
R2470 VDD2.n170 VDD2.n116 10.4732
R2471 VDD2.n146 VDD2.n145 10.4732
R2472 VDD2.n44 VDD2.n43 10.4732
R2473 VDD2.n68 VDD2.n14 10.4732
R2474 VDD2.n90 VDD2.n4 10.4732
R2475 VDD2.n195 VDD2.n194 9.69747
R2476 VDD2.n169 VDD2.n118 9.69747
R2477 VDD2.n149 VDD2.n128 9.69747
R2478 VDD2.n47 VDD2.n26 9.69747
R2479 VDD2.n67 VDD2.n16 9.69747
R2480 VDD2.n94 VDD2.n93 9.69747
R2481 VDD2.n201 VDD2.n200 9.45567
R2482 VDD2.n100 VDD2.n99 9.45567
R2483 VDD2.n161 VDD2.n160 9.3005
R2484 VDD2.n120 VDD2.n119 9.3005
R2485 VDD2.n167 VDD2.n166 9.3005
R2486 VDD2.n169 VDD2.n168 9.3005
R2487 VDD2.n116 VDD2.n115 9.3005
R2488 VDD2.n175 VDD2.n174 9.3005
R2489 VDD2.n177 VDD2.n176 9.3005
R2490 VDD2.n113 VDD2.n110 9.3005
R2491 VDD2.n200 VDD2.n199 9.3005
R2492 VDD2.n103 VDD2.n102 9.3005
R2493 VDD2.n194 VDD2.n193 9.3005
R2494 VDD2.n192 VDD2.n191 9.3005
R2495 VDD2.n107 VDD2.n106 9.3005
R2496 VDD2.n186 VDD2.n185 9.3005
R2497 VDD2.n184 VDD2.n183 9.3005
R2498 VDD2.n159 VDD2.n158 9.3005
R2499 VDD2.n124 VDD2.n123 9.3005
R2500 VDD2.n153 VDD2.n152 9.3005
R2501 VDD2.n151 VDD2.n150 9.3005
R2502 VDD2.n128 VDD2.n127 9.3005
R2503 VDD2.n145 VDD2.n144 9.3005
R2504 VDD2.n143 VDD2.n142 9.3005
R2505 VDD2.n132 VDD2.n131 9.3005
R2506 VDD2.n137 VDD2.n136 9.3005
R2507 VDD2.n99 VDD2.n98 9.3005
R2508 VDD2.n2 VDD2.n1 9.3005
R2509 VDD2.n93 VDD2.n92 9.3005
R2510 VDD2.n91 VDD2.n90 9.3005
R2511 VDD2.n6 VDD2.n5 9.3005
R2512 VDD2.n85 VDD2.n84 9.3005
R2513 VDD2.n83 VDD2.n82 9.3005
R2514 VDD2.n22 VDD2.n21 9.3005
R2515 VDD2.n51 VDD2.n50 9.3005
R2516 VDD2.n49 VDD2.n48 9.3005
R2517 VDD2.n26 VDD2.n25 9.3005
R2518 VDD2.n43 VDD2.n42 9.3005
R2519 VDD2.n41 VDD2.n40 9.3005
R2520 VDD2.n30 VDD2.n29 9.3005
R2521 VDD2.n35 VDD2.n34 9.3005
R2522 VDD2.n57 VDD2.n56 9.3005
R2523 VDD2.n59 VDD2.n58 9.3005
R2524 VDD2.n18 VDD2.n17 9.3005
R2525 VDD2.n65 VDD2.n64 9.3005
R2526 VDD2.n67 VDD2.n66 9.3005
R2527 VDD2.n14 VDD2.n13 9.3005
R2528 VDD2.n73 VDD2.n72 9.3005
R2529 VDD2.n75 VDD2.n74 9.3005
R2530 VDD2.n76 VDD2.n9 9.3005
R2531 VDD2.n198 VDD2.n103 8.92171
R2532 VDD2.n166 VDD2.n165 8.92171
R2533 VDD2.n150 VDD2.n126 8.92171
R2534 VDD2.n48 VDD2.n24 8.92171
R2535 VDD2.n64 VDD2.n63 8.92171
R2536 VDD2.n97 VDD2.n2 8.92171
R2537 VDD2.n199 VDD2.n101 8.14595
R2538 VDD2.n162 VDD2.n120 8.14595
R2539 VDD2.n154 VDD2.n153 8.14595
R2540 VDD2.n52 VDD2.n51 8.14595
R2541 VDD2.n60 VDD2.n18 8.14595
R2542 VDD2.n98 VDD2.n0 8.14595
R2543 VDD2.n161 VDD2.n122 7.3702
R2544 VDD2.n157 VDD2.n124 7.3702
R2545 VDD2.n55 VDD2.n22 7.3702
R2546 VDD2.n59 VDD2.n20 7.3702
R2547 VDD2.n158 VDD2.n122 6.59444
R2548 VDD2.n158 VDD2.n157 6.59444
R2549 VDD2.n56 VDD2.n55 6.59444
R2550 VDD2.n56 VDD2.n20 6.59444
R2551 VDD2.n201 VDD2.n101 5.81868
R2552 VDD2.n162 VDD2.n161 5.81868
R2553 VDD2.n154 VDD2.n124 5.81868
R2554 VDD2.n52 VDD2.n22 5.81868
R2555 VDD2.n60 VDD2.n59 5.81868
R2556 VDD2.n100 VDD2.n0 5.81868
R2557 VDD2.n199 VDD2.n198 5.04292
R2558 VDD2.n165 VDD2.n120 5.04292
R2559 VDD2.n153 VDD2.n126 5.04292
R2560 VDD2.n51 VDD2.n24 5.04292
R2561 VDD2.n63 VDD2.n18 5.04292
R2562 VDD2.n98 VDD2.n97 5.04292
R2563 VDD2.n136 VDD2.n135 4.38563
R2564 VDD2.n34 VDD2.n33 4.38563
R2565 VDD2.n195 VDD2.n103 4.26717
R2566 VDD2.n166 VDD2.n118 4.26717
R2567 VDD2.n150 VDD2.n149 4.26717
R2568 VDD2.n48 VDD2.n47 4.26717
R2569 VDD2.n64 VDD2.n16 4.26717
R2570 VDD2.n94 VDD2.n2 4.26717
R2571 VDD2.n194 VDD2.n105 3.49141
R2572 VDD2.n170 VDD2.n169 3.49141
R2573 VDD2.n146 VDD2.n128 3.49141
R2574 VDD2.n44 VDD2.n26 3.49141
R2575 VDD2.n68 VDD2.n67 3.49141
R2576 VDD2.n93 VDD2.n4 3.49141
R2577 VDD2.n191 VDD2.n190 2.71565
R2578 VDD2.n173 VDD2.n116 2.71565
R2579 VDD2.n145 VDD2.n130 2.71565
R2580 VDD2.n43 VDD2.n28 2.71565
R2581 VDD2.n71 VDD2.n14 2.71565
R2582 VDD2.n90 VDD2.n89 2.71565
R2583 VDD2.n187 VDD2.n107 1.93989
R2584 VDD2.n174 VDD2.n114 1.93989
R2585 VDD2.n142 VDD2.n141 1.93989
R2586 VDD2.n40 VDD2.n39 1.93989
R2587 VDD2.n72 VDD2.n12 1.93989
R2588 VDD2.n86 VDD2.n6 1.93989
R2589 VDD2.n186 VDD2.n109 1.16414
R2590 VDD2.n178 VDD2.n177 1.16414
R2591 VDD2.n138 VDD2.n132 1.16414
R2592 VDD2.n36 VDD2.n30 1.16414
R2593 VDD2.n77 VDD2.n75 1.16414
R2594 VDD2.n85 VDD2.n8 1.16414
R2595 VDD2 VDD2.n202 0.459552
R2596 VDD2.n183 VDD2.n182 0.388379
R2597 VDD2.n113 VDD2.n111 0.388379
R2598 VDD2.n137 VDD2.n134 0.388379
R2599 VDD2.n35 VDD2.n32 0.388379
R2600 VDD2.n76 VDD2.n10 0.388379
R2601 VDD2.n82 VDD2.n81 0.388379
R2602 VDD2.n200 VDD2.n102 0.155672
R2603 VDD2.n193 VDD2.n102 0.155672
R2604 VDD2.n193 VDD2.n192 0.155672
R2605 VDD2.n192 VDD2.n106 0.155672
R2606 VDD2.n185 VDD2.n106 0.155672
R2607 VDD2.n185 VDD2.n184 0.155672
R2608 VDD2.n184 VDD2.n110 0.155672
R2609 VDD2.n176 VDD2.n110 0.155672
R2610 VDD2.n176 VDD2.n175 0.155672
R2611 VDD2.n175 VDD2.n115 0.155672
R2612 VDD2.n168 VDD2.n115 0.155672
R2613 VDD2.n168 VDD2.n167 0.155672
R2614 VDD2.n167 VDD2.n119 0.155672
R2615 VDD2.n160 VDD2.n119 0.155672
R2616 VDD2.n160 VDD2.n159 0.155672
R2617 VDD2.n159 VDD2.n123 0.155672
R2618 VDD2.n152 VDD2.n123 0.155672
R2619 VDD2.n152 VDD2.n151 0.155672
R2620 VDD2.n151 VDD2.n127 0.155672
R2621 VDD2.n144 VDD2.n127 0.155672
R2622 VDD2.n144 VDD2.n143 0.155672
R2623 VDD2.n143 VDD2.n131 0.155672
R2624 VDD2.n136 VDD2.n131 0.155672
R2625 VDD2.n34 VDD2.n29 0.155672
R2626 VDD2.n41 VDD2.n29 0.155672
R2627 VDD2.n42 VDD2.n41 0.155672
R2628 VDD2.n42 VDD2.n25 0.155672
R2629 VDD2.n49 VDD2.n25 0.155672
R2630 VDD2.n50 VDD2.n49 0.155672
R2631 VDD2.n50 VDD2.n21 0.155672
R2632 VDD2.n57 VDD2.n21 0.155672
R2633 VDD2.n58 VDD2.n57 0.155672
R2634 VDD2.n58 VDD2.n17 0.155672
R2635 VDD2.n65 VDD2.n17 0.155672
R2636 VDD2.n66 VDD2.n65 0.155672
R2637 VDD2.n66 VDD2.n13 0.155672
R2638 VDD2.n73 VDD2.n13 0.155672
R2639 VDD2.n74 VDD2.n73 0.155672
R2640 VDD2.n74 VDD2.n9 0.155672
R2641 VDD2.n83 VDD2.n9 0.155672
R2642 VDD2.n84 VDD2.n83 0.155672
R2643 VDD2.n84 VDD2.n5 0.155672
R2644 VDD2.n91 VDD2.n5 0.155672
R2645 VDD2.n92 VDD2.n91 0.155672
R2646 VDD2.n92 VDD2.n1 0.155672
R2647 VDD2.n99 VDD2.n1 0.155672
C0 VP VDD2 0.288939f
C1 VDD2 VN 3.68435f
C2 VDD2 VTAIL 6.93191f
C3 VP VDD1 3.82082f
C4 VDD1 VN 0.147632f
C5 VDD1 VTAIL 6.89234f
C6 VP VN 6.10054f
C7 VP VTAIL 3.02949f
C8 VN VTAIL 3.01492f
C9 VDD1 VDD2 0.550674f
C10 VDD2 B 5.171494f
C11 VDD1 B 8.146781f
C12 VTAIL B 9.244756f
C13 VN B 11.183779f
C14 VP B 5.472183f
C15 VDD2.n0 B 0.027649f
C16 VDD2.n1 B 0.019958f
C17 VDD2.n2 B 0.010725f
C18 VDD2.n3 B 0.025349f
C19 VDD2.n4 B 0.011355f
C20 VDD2.n5 B 0.019958f
C21 VDD2.n6 B 0.010725f
C22 VDD2.n7 B 0.025349f
C23 VDD2.n8 B 0.011355f
C24 VDD2.n9 B 0.019958f
C25 VDD2.n10 B 0.01104f
C26 VDD2.n11 B 0.025349f
C27 VDD2.n12 B 0.011355f
C28 VDD2.n13 B 0.019958f
C29 VDD2.n14 B 0.010725f
C30 VDD2.n15 B 0.025349f
C31 VDD2.n16 B 0.011355f
C32 VDD2.n17 B 0.019958f
C33 VDD2.n18 B 0.010725f
C34 VDD2.n19 B 0.025349f
C35 VDD2.n20 B 0.011355f
C36 VDD2.n21 B 0.019958f
C37 VDD2.n22 B 0.010725f
C38 VDD2.n23 B 0.025349f
C39 VDD2.n24 B 0.011355f
C40 VDD2.n25 B 0.019958f
C41 VDD2.n26 B 0.010725f
C42 VDD2.n27 B 0.025349f
C43 VDD2.n28 B 0.011355f
C44 VDD2.n29 B 0.019958f
C45 VDD2.n30 B 0.010725f
C46 VDD2.n31 B 0.019012f
C47 VDD2.n32 B 0.014975f
C48 VDD2.t0 B 0.042017f
C49 VDD2.n33 B 0.146234f
C50 VDD2.n34 B 1.59211f
C51 VDD2.n35 B 0.010725f
C52 VDD2.n36 B 0.011355f
C53 VDD2.n37 B 0.025349f
C54 VDD2.n38 B 0.025349f
C55 VDD2.n39 B 0.011355f
C56 VDD2.n40 B 0.010725f
C57 VDD2.n41 B 0.019958f
C58 VDD2.n42 B 0.019958f
C59 VDD2.n43 B 0.010725f
C60 VDD2.n44 B 0.011355f
C61 VDD2.n45 B 0.025349f
C62 VDD2.n46 B 0.025349f
C63 VDD2.n47 B 0.011355f
C64 VDD2.n48 B 0.010725f
C65 VDD2.n49 B 0.019958f
C66 VDD2.n50 B 0.019958f
C67 VDD2.n51 B 0.010725f
C68 VDD2.n52 B 0.011355f
C69 VDD2.n53 B 0.025349f
C70 VDD2.n54 B 0.025349f
C71 VDD2.n55 B 0.011355f
C72 VDD2.n56 B 0.010725f
C73 VDD2.n57 B 0.019958f
C74 VDD2.n58 B 0.019958f
C75 VDD2.n59 B 0.010725f
C76 VDD2.n60 B 0.011355f
C77 VDD2.n61 B 0.025349f
C78 VDD2.n62 B 0.025349f
C79 VDD2.n63 B 0.011355f
C80 VDD2.n64 B 0.010725f
C81 VDD2.n65 B 0.019958f
C82 VDD2.n66 B 0.019958f
C83 VDD2.n67 B 0.010725f
C84 VDD2.n68 B 0.011355f
C85 VDD2.n69 B 0.025349f
C86 VDD2.n70 B 0.025349f
C87 VDD2.n71 B 0.011355f
C88 VDD2.n72 B 0.010725f
C89 VDD2.n73 B 0.019958f
C90 VDD2.n74 B 0.019958f
C91 VDD2.n75 B 0.010725f
C92 VDD2.n76 B 0.010725f
C93 VDD2.n77 B 0.011355f
C94 VDD2.n78 B 0.025349f
C95 VDD2.n79 B 0.025349f
C96 VDD2.n80 B 0.025349f
C97 VDD2.n81 B 0.01104f
C98 VDD2.n82 B 0.010725f
C99 VDD2.n83 B 0.019958f
C100 VDD2.n84 B 0.019958f
C101 VDD2.n85 B 0.010725f
C102 VDD2.n86 B 0.011355f
C103 VDD2.n87 B 0.025349f
C104 VDD2.n88 B 0.025349f
C105 VDD2.n89 B 0.011355f
C106 VDD2.n90 B 0.010725f
C107 VDD2.n91 B 0.019958f
C108 VDD2.n92 B 0.019958f
C109 VDD2.n93 B 0.010725f
C110 VDD2.n94 B 0.011355f
C111 VDD2.n95 B 0.025349f
C112 VDD2.n96 B 0.054162f
C113 VDD2.n97 B 0.011355f
C114 VDD2.n98 B 0.010725f
C115 VDD2.n99 B 0.045314f
C116 VDD2.n100 B 0.715412f
C117 VDD2.n101 B 0.027649f
C118 VDD2.n102 B 0.019958f
C119 VDD2.n103 B 0.010725f
C120 VDD2.n104 B 0.025349f
C121 VDD2.n105 B 0.011355f
C122 VDD2.n106 B 0.019958f
C123 VDD2.n107 B 0.010725f
C124 VDD2.n108 B 0.025349f
C125 VDD2.n109 B 0.011355f
C126 VDD2.n110 B 0.019958f
C127 VDD2.n111 B 0.01104f
C128 VDD2.n112 B 0.025349f
C129 VDD2.n113 B 0.010725f
C130 VDD2.n114 B 0.011355f
C131 VDD2.n115 B 0.019958f
C132 VDD2.n116 B 0.010725f
C133 VDD2.n117 B 0.025349f
C134 VDD2.n118 B 0.011355f
C135 VDD2.n119 B 0.019958f
C136 VDD2.n120 B 0.010725f
C137 VDD2.n121 B 0.025349f
C138 VDD2.n122 B 0.011355f
C139 VDD2.n123 B 0.019958f
C140 VDD2.n124 B 0.010725f
C141 VDD2.n125 B 0.025349f
C142 VDD2.n126 B 0.011355f
C143 VDD2.n127 B 0.019958f
C144 VDD2.n128 B 0.010725f
C145 VDD2.n129 B 0.025349f
C146 VDD2.n130 B 0.011355f
C147 VDD2.n131 B 0.019958f
C148 VDD2.n132 B 0.010725f
C149 VDD2.n133 B 0.019012f
C150 VDD2.n134 B 0.014975f
C151 VDD2.t1 B 0.042017f
C152 VDD2.n135 B 0.146234f
C153 VDD2.n136 B 1.59211f
C154 VDD2.n137 B 0.010725f
C155 VDD2.n138 B 0.011355f
C156 VDD2.n139 B 0.025349f
C157 VDD2.n140 B 0.025349f
C158 VDD2.n141 B 0.011355f
C159 VDD2.n142 B 0.010725f
C160 VDD2.n143 B 0.019958f
C161 VDD2.n144 B 0.019958f
C162 VDD2.n145 B 0.010725f
C163 VDD2.n146 B 0.011355f
C164 VDD2.n147 B 0.025349f
C165 VDD2.n148 B 0.025349f
C166 VDD2.n149 B 0.011355f
C167 VDD2.n150 B 0.010725f
C168 VDD2.n151 B 0.019958f
C169 VDD2.n152 B 0.019958f
C170 VDD2.n153 B 0.010725f
C171 VDD2.n154 B 0.011355f
C172 VDD2.n155 B 0.025349f
C173 VDD2.n156 B 0.025349f
C174 VDD2.n157 B 0.011355f
C175 VDD2.n158 B 0.010725f
C176 VDD2.n159 B 0.019958f
C177 VDD2.n160 B 0.019958f
C178 VDD2.n161 B 0.010725f
C179 VDD2.n162 B 0.011355f
C180 VDD2.n163 B 0.025349f
C181 VDD2.n164 B 0.025349f
C182 VDD2.n165 B 0.011355f
C183 VDD2.n166 B 0.010725f
C184 VDD2.n167 B 0.019958f
C185 VDD2.n168 B 0.019958f
C186 VDD2.n169 B 0.010725f
C187 VDD2.n170 B 0.011355f
C188 VDD2.n171 B 0.025349f
C189 VDD2.n172 B 0.025349f
C190 VDD2.n173 B 0.011355f
C191 VDD2.n174 B 0.010725f
C192 VDD2.n175 B 0.019958f
C193 VDD2.n176 B 0.019958f
C194 VDD2.n177 B 0.010725f
C195 VDD2.n178 B 0.011355f
C196 VDD2.n179 B 0.025349f
C197 VDD2.n180 B 0.025349f
C198 VDD2.n181 B 0.025349f
C199 VDD2.n182 B 0.01104f
C200 VDD2.n183 B 0.010725f
C201 VDD2.n184 B 0.019958f
C202 VDD2.n185 B 0.019958f
C203 VDD2.n186 B 0.010725f
C204 VDD2.n187 B 0.011355f
C205 VDD2.n188 B 0.025349f
C206 VDD2.n189 B 0.025349f
C207 VDD2.n190 B 0.011355f
C208 VDD2.n191 B 0.010725f
C209 VDD2.n192 B 0.019958f
C210 VDD2.n193 B 0.019958f
C211 VDD2.n194 B 0.010725f
C212 VDD2.n195 B 0.011355f
C213 VDD2.n196 B 0.025349f
C214 VDD2.n197 B 0.054162f
C215 VDD2.n198 B 0.011355f
C216 VDD2.n199 B 0.010725f
C217 VDD2.n200 B 0.045314f
C218 VDD2.n201 B 0.043994f
C219 VDD2.n202 B 2.77321f
C220 VN.t1 B 3.41916f
C221 VN.t0 B 3.73358f
C222 VDD1.n0 B 0.027717f
C223 VDD1.n1 B 0.020007f
C224 VDD1.n2 B 0.010751f
C225 VDD1.n3 B 0.025412f
C226 VDD1.n4 B 0.011383f
C227 VDD1.n5 B 0.020007f
C228 VDD1.n6 B 0.010751f
C229 VDD1.n7 B 0.025412f
C230 VDD1.n8 B 0.011383f
C231 VDD1.n9 B 0.020007f
C232 VDD1.n10 B 0.011067f
C233 VDD1.n11 B 0.025412f
C234 VDD1.n12 B 0.010751f
C235 VDD1.n13 B 0.011383f
C236 VDD1.n14 B 0.020007f
C237 VDD1.n15 B 0.010751f
C238 VDD1.n16 B 0.025412f
C239 VDD1.n17 B 0.011383f
C240 VDD1.n18 B 0.020007f
C241 VDD1.n19 B 0.010751f
C242 VDD1.n20 B 0.025412f
C243 VDD1.n21 B 0.011383f
C244 VDD1.n22 B 0.020007f
C245 VDD1.n23 B 0.010751f
C246 VDD1.n24 B 0.025412f
C247 VDD1.n25 B 0.011383f
C248 VDD1.n26 B 0.020007f
C249 VDD1.n27 B 0.010751f
C250 VDD1.n28 B 0.025412f
C251 VDD1.n29 B 0.011383f
C252 VDD1.n30 B 0.020007f
C253 VDD1.n31 B 0.010751f
C254 VDD1.n32 B 0.019059f
C255 VDD1.n33 B 0.015011f
C256 VDD1.t0 B 0.042121f
C257 VDD1.n34 B 0.146594f
C258 VDD1.n35 B 1.59603f
C259 VDD1.n36 B 0.010751f
C260 VDD1.n37 B 0.011383f
C261 VDD1.n38 B 0.025412f
C262 VDD1.n39 B 0.025412f
C263 VDD1.n40 B 0.011383f
C264 VDD1.n41 B 0.010751f
C265 VDD1.n42 B 0.020007f
C266 VDD1.n43 B 0.020007f
C267 VDD1.n44 B 0.010751f
C268 VDD1.n45 B 0.011383f
C269 VDD1.n46 B 0.025412f
C270 VDD1.n47 B 0.025412f
C271 VDD1.n48 B 0.011383f
C272 VDD1.n49 B 0.010751f
C273 VDD1.n50 B 0.020007f
C274 VDD1.n51 B 0.020007f
C275 VDD1.n52 B 0.010751f
C276 VDD1.n53 B 0.011383f
C277 VDD1.n54 B 0.025412f
C278 VDD1.n55 B 0.025412f
C279 VDD1.n56 B 0.011383f
C280 VDD1.n57 B 0.010751f
C281 VDD1.n58 B 0.020007f
C282 VDD1.n59 B 0.020007f
C283 VDD1.n60 B 0.010751f
C284 VDD1.n61 B 0.011383f
C285 VDD1.n62 B 0.025412f
C286 VDD1.n63 B 0.025412f
C287 VDD1.n64 B 0.011383f
C288 VDD1.n65 B 0.010751f
C289 VDD1.n66 B 0.020007f
C290 VDD1.n67 B 0.020007f
C291 VDD1.n68 B 0.010751f
C292 VDD1.n69 B 0.011383f
C293 VDD1.n70 B 0.025412f
C294 VDD1.n71 B 0.025412f
C295 VDD1.n72 B 0.011383f
C296 VDD1.n73 B 0.010751f
C297 VDD1.n74 B 0.020007f
C298 VDD1.n75 B 0.020007f
C299 VDD1.n76 B 0.010751f
C300 VDD1.n77 B 0.011383f
C301 VDD1.n78 B 0.025412f
C302 VDD1.n79 B 0.025412f
C303 VDD1.n80 B 0.025412f
C304 VDD1.n81 B 0.011067f
C305 VDD1.n82 B 0.010751f
C306 VDD1.n83 B 0.020007f
C307 VDD1.n84 B 0.020007f
C308 VDD1.n85 B 0.010751f
C309 VDD1.n86 B 0.011383f
C310 VDD1.n87 B 0.025412f
C311 VDD1.n88 B 0.025412f
C312 VDD1.n89 B 0.011383f
C313 VDD1.n90 B 0.010751f
C314 VDD1.n91 B 0.020007f
C315 VDD1.n92 B 0.020007f
C316 VDD1.n93 B 0.010751f
C317 VDD1.n94 B 0.011383f
C318 VDD1.n95 B 0.025412f
C319 VDD1.n96 B 0.054295f
C320 VDD1.n97 B 0.011383f
C321 VDD1.n98 B 0.010751f
C322 VDD1.n99 B 0.045426f
C323 VDD1.n100 B 0.04474f
C324 VDD1.n101 B 0.027717f
C325 VDD1.n102 B 0.020007f
C326 VDD1.n103 B 0.010751f
C327 VDD1.n104 B 0.025412f
C328 VDD1.n105 B 0.011383f
C329 VDD1.n106 B 0.020007f
C330 VDD1.n107 B 0.010751f
C331 VDD1.n108 B 0.025412f
C332 VDD1.n109 B 0.011383f
C333 VDD1.n110 B 0.020007f
C334 VDD1.n111 B 0.011067f
C335 VDD1.n112 B 0.025412f
C336 VDD1.n113 B 0.011383f
C337 VDD1.n114 B 0.020007f
C338 VDD1.n115 B 0.010751f
C339 VDD1.n116 B 0.025412f
C340 VDD1.n117 B 0.011383f
C341 VDD1.n118 B 0.020007f
C342 VDD1.n119 B 0.010751f
C343 VDD1.n120 B 0.025412f
C344 VDD1.n121 B 0.011383f
C345 VDD1.n122 B 0.020007f
C346 VDD1.n123 B 0.010751f
C347 VDD1.n124 B 0.025412f
C348 VDD1.n125 B 0.011383f
C349 VDD1.n126 B 0.020007f
C350 VDD1.n127 B 0.010751f
C351 VDD1.n128 B 0.025412f
C352 VDD1.n129 B 0.011383f
C353 VDD1.n130 B 0.020007f
C354 VDD1.n131 B 0.010751f
C355 VDD1.n132 B 0.019059f
C356 VDD1.n133 B 0.015011f
C357 VDD1.t1 B 0.042121f
C358 VDD1.n134 B 0.146594f
C359 VDD1.n135 B 1.59603f
C360 VDD1.n136 B 0.010751f
C361 VDD1.n137 B 0.011383f
C362 VDD1.n138 B 0.025412f
C363 VDD1.n139 B 0.025412f
C364 VDD1.n140 B 0.011383f
C365 VDD1.n141 B 0.010751f
C366 VDD1.n142 B 0.020007f
C367 VDD1.n143 B 0.020007f
C368 VDD1.n144 B 0.010751f
C369 VDD1.n145 B 0.011383f
C370 VDD1.n146 B 0.025412f
C371 VDD1.n147 B 0.025412f
C372 VDD1.n148 B 0.011383f
C373 VDD1.n149 B 0.010751f
C374 VDD1.n150 B 0.020007f
C375 VDD1.n151 B 0.020007f
C376 VDD1.n152 B 0.010751f
C377 VDD1.n153 B 0.011383f
C378 VDD1.n154 B 0.025412f
C379 VDD1.n155 B 0.025412f
C380 VDD1.n156 B 0.011383f
C381 VDD1.n157 B 0.010751f
C382 VDD1.n158 B 0.020007f
C383 VDD1.n159 B 0.020007f
C384 VDD1.n160 B 0.010751f
C385 VDD1.n161 B 0.011383f
C386 VDD1.n162 B 0.025412f
C387 VDD1.n163 B 0.025412f
C388 VDD1.n164 B 0.011383f
C389 VDD1.n165 B 0.010751f
C390 VDD1.n166 B 0.020007f
C391 VDD1.n167 B 0.020007f
C392 VDD1.n168 B 0.010751f
C393 VDD1.n169 B 0.011383f
C394 VDD1.n170 B 0.025412f
C395 VDD1.n171 B 0.025412f
C396 VDD1.n172 B 0.011383f
C397 VDD1.n173 B 0.010751f
C398 VDD1.n174 B 0.020007f
C399 VDD1.n175 B 0.020007f
C400 VDD1.n176 B 0.010751f
C401 VDD1.n177 B 0.010751f
C402 VDD1.n178 B 0.011383f
C403 VDD1.n179 B 0.025412f
C404 VDD1.n180 B 0.025412f
C405 VDD1.n181 B 0.025412f
C406 VDD1.n182 B 0.011067f
C407 VDD1.n183 B 0.010751f
C408 VDD1.n184 B 0.020007f
C409 VDD1.n185 B 0.020007f
C410 VDD1.n186 B 0.010751f
C411 VDD1.n187 B 0.011383f
C412 VDD1.n188 B 0.025412f
C413 VDD1.n189 B 0.025412f
C414 VDD1.n190 B 0.011383f
C415 VDD1.n191 B 0.010751f
C416 VDD1.n192 B 0.020007f
C417 VDD1.n193 B 0.020007f
C418 VDD1.n194 B 0.010751f
C419 VDD1.n195 B 0.011383f
C420 VDD1.n196 B 0.025412f
C421 VDD1.n197 B 0.054295f
C422 VDD1.n198 B 0.011383f
C423 VDD1.n199 B 0.010751f
C424 VDD1.n200 B 0.045426f
C425 VDD1.n201 B 0.752498f
C426 VTAIL.n0 B 0.027065f
C427 VTAIL.n1 B 0.019537f
C428 VTAIL.n2 B 0.010498f
C429 VTAIL.n3 B 0.024814f
C430 VTAIL.n4 B 0.011116f
C431 VTAIL.n5 B 0.019537f
C432 VTAIL.n6 B 0.010498f
C433 VTAIL.n7 B 0.024814f
C434 VTAIL.n8 B 0.011116f
C435 VTAIL.n9 B 0.019537f
C436 VTAIL.n10 B 0.010807f
C437 VTAIL.n11 B 0.024814f
C438 VTAIL.n12 B 0.011116f
C439 VTAIL.n13 B 0.019537f
C440 VTAIL.n14 B 0.010498f
C441 VTAIL.n15 B 0.024814f
C442 VTAIL.n16 B 0.011116f
C443 VTAIL.n17 B 0.019537f
C444 VTAIL.n18 B 0.010498f
C445 VTAIL.n19 B 0.024814f
C446 VTAIL.n20 B 0.011116f
C447 VTAIL.n21 B 0.019537f
C448 VTAIL.n22 B 0.010498f
C449 VTAIL.n23 B 0.024814f
C450 VTAIL.n24 B 0.011116f
C451 VTAIL.n25 B 0.019537f
C452 VTAIL.n26 B 0.010498f
C453 VTAIL.n27 B 0.024814f
C454 VTAIL.n28 B 0.011116f
C455 VTAIL.n29 B 0.019537f
C456 VTAIL.n30 B 0.010498f
C457 VTAIL.n31 B 0.01861f
C458 VTAIL.n32 B 0.014658f
C459 VTAIL.t2 B 0.04113f
C460 VTAIL.n33 B 0.143146f
C461 VTAIL.n34 B 1.5585f
C462 VTAIL.n35 B 0.010498f
C463 VTAIL.n36 B 0.011116f
C464 VTAIL.n37 B 0.024814f
C465 VTAIL.n38 B 0.024814f
C466 VTAIL.n39 B 0.011116f
C467 VTAIL.n40 B 0.010498f
C468 VTAIL.n41 B 0.019537f
C469 VTAIL.n42 B 0.019537f
C470 VTAIL.n43 B 0.010498f
C471 VTAIL.n44 B 0.011116f
C472 VTAIL.n45 B 0.024814f
C473 VTAIL.n46 B 0.024814f
C474 VTAIL.n47 B 0.011116f
C475 VTAIL.n48 B 0.010498f
C476 VTAIL.n49 B 0.019537f
C477 VTAIL.n50 B 0.019537f
C478 VTAIL.n51 B 0.010498f
C479 VTAIL.n52 B 0.011116f
C480 VTAIL.n53 B 0.024814f
C481 VTAIL.n54 B 0.024814f
C482 VTAIL.n55 B 0.011116f
C483 VTAIL.n56 B 0.010498f
C484 VTAIL.n57 B 0.019537f
C485 VTAIL.n58 B 0.019537f
C486 VTAIL.n59 B 0.010498f
C487 VTAIL.n60 B 0.011116f
C488 VTAIL.n61 B 0.024814f
C489 VTAIL.n62 B 0.024814f
C490 VTAIL.n63 B 0.011116f
C491 VTAIL.n64 B 0.010498f
C492 VTAIL.n65 B 0.019537f
C493 VTAIL.n66 B 0.019537f
C494 VTAIL.n67 B 0.010498f
C495 VTAIL.n68 B 0.011116f
C496 VTAIL.n69 B 0.024814f
C497 VTAIL.n70 B 0.024814f
C498 VTAIL.n71 B 0.011116f
C499 VTAIL.n72 B 0.010498f
C500 VTAIL.n73 B 0.019537f
C501 VTAIL.n74 B 0.019537f
C502 VTAIL.n75 B 0.010498f
C503 VTAIL.n76 B 0.010498f
C504 VTAIL.n77 B 0.011116f
C505 VTAIL.n78 B 0.024814f
C506 VTAIL.n79 B 0.024814f
C507 VTAIL.n80 B 0.024814f
C508 VTAIL.n81 B 0.010807f
C509 VTAIL.n82 B 0.010498f
C510 VTAIL.n83 B 0.019537f
C511 VTAIL.n84 B 0.019537f
C512 VTAIL.n85 B 0.010498f
C513 VTAIL.n86 B 0.011116f
C514 VTAIL.n87 B 0.024814f
C515 VTAIL.n88 B 0.024814f
C516 VTAIL.n89 B 0.011116f
C517 VTAIL.n90 B 0.010498f
C518 VTAIL.n91 B 0.019537f
C519 VTAIL.n92 B 0.019537f
C520 VTAIL.n93 B 0.010498f
C521 VTAIL.n94 B 0.011116f
C522 VTAIL.n95 B 0.024814f
C523 VTAIL.n96 B 0.053019f
C524 VTAIL.n97 B 0.011116f
C525 VTAIL.n98 B 0.010498f
C526 VTAIL.n99 B 0.044357f
C527 VTAIL.n100 B 0.029569f
C528 VTAIL.n101 B 1.5302f
C529 VTAIL.n102 B 0.027065f
C530 VTAIL.n103 B 0.019537f
C531 VTAIL.n104 B 0.010498f
C532 VTAIL.n105 B 0.024814f
C533 VTAIL.n106 B 0.011116f
C534 VTAIL.n107 B 0.019537f
C535 VTAIL.n108 B 0.010498f
C536 VTAIL.n109 B 0.024814f
C537 VTAIL.n110 B 0.011116f
C538 VTAIL.n111 B 0.019537f
C539 VTAIL.n112 B 0.010807f
C540 VTAIL.n113 B 0.024814f
C541 VTAIL.n114 B 0.010498f
C542 VTAIL.n115 B 0.011116f
C543 VTAIL.n116 B 0.019537f
C544 VTAIL.n117 B 0.010498f
C545 VTAIL.n118 B 0.024814f
C546 VTAIL.n119 B 0.011116f
C547 VTAIL.n120 B 0.019537f
C548 VTAIL.n121 B 0.010498f
C549 VTAIL.n122 B 0.024814f
C550 VTAIL.n123 B 0.011116f
C551 VTAIL.n124 B 0.019537f
C552 VTAIL.n125 B 0.010498f
C553 VTAIL.n126 B 0.024814f
C554 VTAIL.n127 B 0.011116f
C555 VTAIL.n128 B 0.019537f
C556 VTAIL.n129 B 0.010498f
C557 VTAIL.n130 B 0.024814f
C558 VTAIL.n131 B 0.011116f
C559 VTAIL.n132 B 0.019537f
C560 VTAIL.n133 B 0.010498f
C561 VTAIL.n134 B 0.01861f
C562 VTAIL.n135 B 0.014658f
C563 VTAIL.t1 B 0.04113f
C564 VTAIL.n136 B 0.143146f
C565 VTAIL.n137 B 1.5585f
C566 VTAIL.n138 B 0.010498f
C567 VTAIL.n139 B 0.011116f
C568 VTAIL.n140 B 0.024814f
C569 VTAIL.n141 B 0.024814f
C570 VTAIL.n142 B 0.011116f
C571 VTAIL.n143 B 0.010498f
C572 VTAIL.n144 B 0.019537f
C573 VTAIL.n145 B 0.019537f
C574 VTAIL.n146 B 0.010498f
C575 VTAIL.n147 B 0.011116f
C576 VTAIL.n148 B 0.024814f
C577 VTAIL.n149 B 0.024814f
C578 VTAIL.n150 B 0.011116f
C579 VTAIL.n151 B 0.010498f
C580 VTAIL.n152 B 0.019537f
C581 VTAIL.n153 B 0.019537f
C582 VTAIL.n154 B 0.010498f
C583 VTAIL.n155 B 0.011116f
C584 VTAIL.n156 B 0.024814f
C585 VTAIL.n157 B 0.024814f
C586 VTAIL.n158 B 0.011116f
C587 VTAIL.n159 B 0.010498f
C588 VTAIL.n160 B 0.019537f
C589 VTAIL.n161 B 0.019537f
C590 VTAIL.n162 B 0.010498f
C591 VTAIL.n163 B 0.011116f
C592 VTAIL.n164 B 0.024814f
C593 VTAIL.n165 B 0.024814f
C594 VTAIL.n166 B 0.011116f
C595 VTAIL.n167 B 0.010498f
C596 VTAIL.n168 B 0.019537f
C597 VTAIL.n169 B 0.019537f
C598 VTAIL.n170 B 0.010498f
C599 VTAIL.n171 B 0.011116f
C600 VTAIL.n172 B 0.024814f
C601 VTAIL.n173 B 0.024814f
C602 VTAIL.n174 B 0.011116f
C603 VTAIL.n175 B 0.010498f
C604 VTAIL.n176 B 0.019537f
C605 VTAIL.n177 B 0.019537f
C606 VTAIL.n178 B 0.010498f
C607 VTAIL.n179 B 0.011116f
C608 VTAIL.n180 B 0.024814f
C609 VTAIL.n181 B 0.024814f
C610 VTAIL.n182 B 0.024814f
C611 VTAIL.n183 B 0.010807f
C612 VTAIL.n184 B 0.010498f
C613 VTAIL.n185 B 0.019537f
C614 VTAIL.n186 B 0.019537f
C615 VTAIL.n187 B 0.010498f
C616 VTAIL.n188 B 0.011116f
C617 VTAIL.n189 B 0.024814f
C618 VTAIL.n190 B 0.024814f
C619 VTAIL.n191 B 0.011116f
C620 VTAIL.n192 B 0.010498f
C621 VTAIL.n193 B 0.019537f
C622 VTAIL.n194 B 0.019537f
C623 VTAIL.n195 B 0.010498f
C624 VTAIL.n196 B 0.011116f
C625 VTAIL.n197 B 0.024814f
C626 VTAIL.n198 B 0.053019f
C627 VTAIL.n199 B 0.011116f
C628 VTAIL.n200 B 0.010498f
C629 VTAIL.n201 B 0.044357f
C630 VTAIL.n202 B 0.029569f
C631 VTAIL.n203 B 1.55177f
C632 VTAIL.n204 B 0.027065f
C633 VTAIL.n205 B 0.019537f
C634 VTAIL.n206 B 0.010498f
C635 VTAIL.n207 B 0.024814f
C636 VTAIL.n208 B 0.011116f
C637 VTAIL.n209 B 0.019537f
C638 VTAIL.n210 B 0.010498f
C639 VTAIL.n211 B 0.024814f
C640 VTAIL.n212 B 0.011116f
C641 VTAIL.n213 B 0.019537f
C642 VTAIL.n214 B 0.010807f
C643 VTAIL.n215 B 0.024814f
C644 VTAIL.n216 B 0.010498f
C645 VTAIL.n217 B 0.011116f
C646 VTAIL.n218 B 0.019537f
C647 VTAIL.n219 B 0.010498f
C648 VTAIL.n220 B 0.024814f
C649 VTAIL.n221 B 0.011116f
C650 VTAIL.n222 B 0.019537f
C651 VTAIL.n223 B 0.010498f
C652 VTAIL.n224 B 0.024814f
C653 VTAIL.n225 B 0.011116f
C654 VTAIL.n226 B 0.019537f
C655 VTAIL.n227 B 0.010498f
C656 VTAIL.n228 B 0.024814f
C657 VTAIL.n229 B 0.011116f
C658 VTAIL.n230 B 0.019537f
C659 VTAIL.n231 B 0.010498f
C660 VTAIL.n232 B 0.024814f
C661 VTAIL.n233 B 0.011116f
C662 VTAIL.n234 B 0.019537f
C663 VTAIL.n235 B 0.010498f
C664 VTAIL.n236 B 0.01861f
C665 VTAIL.n237 B 0.014658f
C666 VTAIL.t3 B 0.04113f
C667 VTAIL.n238 B 0.143146f
C668 VTAIL.n239 B 1.5585f
C669 VTAIL.n240 B 0.010498f
C670 VTAIL.n241 B 0.011116f
C671 VTAIL.n242 B 0.024814f
C672 VTAIL.n243 B 0.024814f
C673 VTAIL.n244 B 0.011116f
C674 VTAIL.n245 B 0.010498f
C675 VTAIL.n246 B 0.019537f
C676 VTAIL.n247 B 0.019537f
C677 VTAIL.n248 B 0.010498f
C678 VTAIL.n249 B 0.011116f
C679 VTAIL.n250 B 0.024814f
C680 VTAIL.n251 B 0.024814f
C681 VTAIL.n252 B 0.011116f
C682 VTAIL.n253 B 0.010498f
C683 VTAIL.n254 B 0.019537f
C684 VTAIL.n255 B 0.019537f
C685 VTAIL.n256 B 0.010498f
C686 VTAIL.n257 B 0.011116f
C687 VTAIL.n258 B 0.024814f
C688 VTAIL.n259 B 0.024814f
C689 VTAIL.n260 B 0.011116f
C690 VTAIL.n261 B 0.010498f
C691 VTAIL.n262 B 0.019537f
C692 VTAIL.n263 B 0.019537f
C693 VTAIL.n264 B 0.010498f
C694 VTAIL.n265 B 0.011116f
C695 VTAIL.n266 B 0.024814f
C696 VTAIL.n267 B 0.024814f
C697 VTAIL.n268 B 0.011116f
C698 VTAIL.n269 B 0.010498f
C699 VTAIL.n270 B 0.019537f
C700 VTAIL.n271 B 0.019537f
C701 VTAIL.n272 B 0.010498f
C702 VTAIL.n273 B 0.011116f
C703 VTAIL.n274 B 0.024814f
C704 VTAIL.n275 B 0.024814f
C705 VTAIL.n276 B 0.011116f
C706 VTAIL.n277 B 0.010498f
C707 VTAIL.n278 B 0.019537f
C708 VTAIL.n279 B 0.019537f
C709 VTAIL.n280 B 0.010498f
C710 VTAIL.n281 B 0.011116f
C711 VTAIL.n282 B 0.024814f
C712 VTAIL.n283 B 0.024814f
C713 VTAIL.n284 B 0.024814f
C714 VTAIL.n285 B 0.010807f
C715 VTAIL.n286 B 0.010498f
C716 VTAIL.n287 B 0.019537f
C717 VTAIL.n288 B 0.019537f
C718 VTAIL.n289 B 0.010498f
C719 VTAIL.n290 B 0.011116f
C720 VTAIL.n291 B 0.024814f
C721 VTAIL.n292 B 0.024814f
C722 VTAIL.n293 B 0.011116f
C723 VTAIL.n294 B 0.010498f
C724 VTAIL.n295 B 0.019537f
C725 VTAIL.n296 B 0.019537f
C726 VTAIL.n297 B 0.010498f
C727 VTAIL.n298 B 0.011116f
C728 VTAIL.n299 B 0.024814f
C729 VTAIL.n300 B 0.053019f
C730 VTAIL.n301 B 0.011116f
C731 VTAIL.n302 B 0.010498f
C732 VTAIL.n303 B 0.044357f
C733 VTAIL.n304 B 0.029569f
C734 VTAIL.n305 B 1.45083f
C735 VTAIL.n306 B 0.027065f
C736 VTAIL.n307 B 0.019537f
C737 VTAIL.n308 B 0.010498f
C738 VTAIL.n309 B 0.024814f
C739 VTAIL.n310 B 0.011116f
C740 VTAIL.n311 B 0.019537f
C741 VTAIL.n312 B 0.010498f
C742 VTAIL.n313 B 0.024814f
C743 VTAIL.n314 B 0.011116f
C744 VTAIL.n315 B 0.019537f
C745 VTAIL.n316 B 0.010807f
C746 VTAIL.n317 B 0.024814f
C747 VTAIL.n318 B 0.011116f
C748 VTAIL.n319 B 0.019537f
C749 VTAIL.n320 B 0.010498f
C750 VTAIL.n321 B 0.024814f
C751 VTAIL.n322 B 0.011116f
C752 VTAIL.n323 B 0.019537f
C753 VTAIL.n324 B 0.010498f
C754 VTAIL.n325 B 0.024814f
C755 VTAIL.n326 B 0.011116f
C756 VTAIL.n327 B 0.019537f
C757 VTAIL.n328 B 0.010498f
C758 VTAIL.n329 B 0.024814f
C759 VTAIL.n330 B 0.011116f
C760 VTAIL.n331 B 0.019537f
C761 VTAIL.n332 B 0.010498f
C762 VTAIL.n333 B 0.024814f
C763 VTAIL.n334 B 0.011116f
C764 VTAIL.n335 B 0.019537f
C765 VTAIL.n336 B 0.010498f
C766 VTAIL.n337 B 0.01861f
C767 VTAIL.n338 B 0.014658f
C768 VTAIL.t0 B 0.04113f
C769 VTAIL.n339 B 0.143146f
C770 VTAIL.n340 B 1.5585f
C771 VTAIL.n341 B 0.010498f
C772 VTAIL.n342 B 0.011116f
C773 VTAIL.n343 B 0.024814f
C774 VTAIL.n344 B 0.024814f
C775 VTAIL.n345 B 0.011116f
C776 VTAIL.n346 B 0.010498f
C777 VTAIL.n347 B 0.019537f
C778 VTAIL.n348 B 0.019537f
C779 VTAIL.n349 B 0.010498f
C780 VTAIL.n350 B 0.011116f
C781 VTAIL.n351 B 0.024814f
C782 VTAIL.n352 B 0.024814f
C783 VTAIL.n353 B 0.011116f
C784 VTAIL.n354 B 0.010498f
C785 VTAIL.n355 B 0.019537f
C786 VTAIL.n356 B 0.019537f
C787 VTAIL.n357 B 0.010498f
C788 VTAIL.n358 B 0.011116f
C789 VTAIL.n359 B 0.024814f
C790 VTAIL.n360 B 0.024814f
C791 VTAIL.n361 B 0.011116f
C792 VTAIL.n362 B 0.010498f
C793 VTAIL.n363 B 0.019537f
C794 VTAIL.n364 B 0.019537f
C795 VTAIL.n365 B 0.010498f
C796 VTAIL.n366 B 0.011116f
C797 VTAIL.n367 B 0.024814f
C798 VTAIL.n368 B 0.024814f
C799 VTAIL.n369 B 0.011116f
C800 VTAIL.n370 B 0.010498f
C801 VTAIL.n371 B 0.019537f
C802 VTAIL.n372 B 0.019537f
C803 VTAIL.n373 B 0.010498f
C804 VTAIL.n374 B 0.011116f
C805 VTAIL.n375 B 0.024814f
C806 VTAIL.n376 B 0.024814f
C807 VTAIL.n377 B 0.011116f
C808 VTAIL.n378 B 0.010498f
C809 VTAIL.n379 B 0.019537f
C810 VTAIL.n380 B 0.019537f
C811 VTAIL.n381 B 0.010498f
C812 VTAIL.n382 B 0.010498f
C813 VTAIL.n383 B 0.011116f
C814 VTAIL.n384 B 0.024814f
C815 VTAIL.n385 B 0.024814f
C816 VTAIL.n386 B 0.024814f
C817 VTAIL.n387 B 0.010807f
C818 VTAIL.n388 B 0.010498f
C819 VTAIL.n389 B 0.019537f
C820 VTAIL.n390 B 0.019537f
C821 VTAIL.n391 B 0.010498f
C822 VTAIL.n392 B 0.011116f
C823 VTAIL.n393 B 0.024814f
C824 VTAIL.n394 B 0.024814f
C825 VTAIL.n395 B 0.011116f
C826 VTAIL.n396 B 0.010498f
C827 VTAIL.n397 B 0.019537f
C828 VTAIL.n398 B 0.019537f
C829 VTAIL.n399 B 0.010498f
C830 VTAIL.n400 B 0.011116f
C831 VTAIL.n401 B 0.024814f
C832 VTAIL.n402 B 0.053019f
C833 VTAIL.n403 B 0.011116f
C834 VTAIL.n404 B 0.010498f
C835 VTAIL.n405 B 0.044357f
C836 VTAIL.n406 B 0.029569f
C837 VTAIL.n407 B 1.39236f
C838 VP.t1 B 3.77533f
C839 VP.t0 B 3.46078f
C840 VP.n0 B 5.6209f
.ends

