* NGSPICE file created from diff_pair_sample_0754.ext - technology: sky130A

.subckt diff_pair_sample_0754 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=0.26565 pd=1.94 as=0.6279 ps=4 w=1.61 l=0.49
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=0.6279 pd=4 as=0 ps=0 w=1.61 l=0.49
X2 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=0.6279 pd=4 as=0 ps=0 w=1.61 l=0.49
X3 VDD2.t3 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.26565 pd=1.94 as=0.6279 ps=4 w=1.61 l=0.49
X4 VTAIL.t1 VN.t1 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6279 pd=4 as=0.26565 ps=1.94 w=1.61 l=0.49
X5 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6279 pd=4 as=0 ps=0 w=1.61 l=0.49
X6 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.6279 pd=4 as=0 ps=0 w=1.61 l=0.49
X7 VDD2.t1 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.26565 pd=1.94 as=0.6279 ps=4 w=1.61 l=0.49
X8 VTAIL.t5 VP.t1 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6279 pd=4 as=0.26565 ps=1.94 w=1.61 l=0.49
X9 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6279 pd=4 as=0.26565 ps=1.94 w=1.61 l=0.49
X10 VTAIL.t6 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6279 pd=4 as=0.26565 ps=1.94 w=1.61 l=0.49
X11 VDD1.t0 VP.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.26565 pd=1.94 as=0.6279 ps=4 w=1.61 l=0.49
R0 VP.n0 VP.t2 180.829
R1 VP.n0 VP.t3 180.804
R2 VP.n4 VP.n3 161.3
R3 VP.n2 VP.n1 161.3
R4 VP.n2 VP.t1 159.847
R5 VP.n3 VP.t0 159.847
R6 VP.n1 VP.n0 102.145
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.189894
R9 VP VP.n4 0.0516364
R10 VTAIL.n7 VTAIL.t2 111.013
R11 VTAIL.n0 VTAIL.t1 111.013
R12 VTAIL.n1 VTAIL.t7 111.013
R13 VTAIL.n2 VTAIL.t5 111.013
R14 VTAIL.n6 VTAIL.t4 111.013
R15 VTAIL.n5 VTAIL.t6 111.013
R16 VTAIL.n4 VTAIL.t0 111.013
R17 VTAIL.n3 VTAIL.t3 111.013
R18 VTAIL.n7 VTAIL.n6 14.4617
R19 VTAIL.n3 VTAIL.n2 14.4617
R20 VTAIL.n4 VTAIL.n3 0.707397
R21 VTAIL.n6 VTAIL.n5 0.707397
R22 VTAIL.n2 VTAIL.n1 0.707397
R23 VTAIL.n5 VTAIL.n4 0.470328
R24 VTAIL.n1 VTAIL.n0 0.470328
R25 VTAIL VTAIL.n0 0.412138
R26 VTAIL VTAIL.n7 0.295759
R27 VDD1 VDD1.n1 143.143
R28 VDD1 VDD1.n0 115.453
R29 VDD1.n0 VDD1.t1 12.2986
R30 VDD1.n0 VDD1.t0 12.2986
R31 VDD1.n1 VDD1.t2 12.2986
R32 VDD1.n1 VDD1.t3 12.2986
R33 B.n293 B.n292 585
R34 B.n112 B.n48 585
R35 B.n111 B.n110 585
R36 B.n109 B.n108 585
R37 B.n107 B.n106 585
R38 B.n105 B.n104 585
R39 B.n103 B.n102 585
R40 B.n101 B.n100 585
R41 B.n99 B.n98 585
R42 B.n97 B.n96 585
R43 B.n95 B.n94 585
R44 B.n92 B.n91 585
R45 B.n90 B.n89 585
R46 B.n88 B.n87 585
R47 B.n86 B.n85 585
R48 B.n84 B.n83 585
R49 B.n82 B.n81 585
R50 B.n80 B.n79 585
R51 B.n78 B.n77 585
R52 B.n76 B.n75 585
R53 B.n74 B.n73 585
R54 B.n71 B.n70 585
R55 B.n69 B.n68 585
R56 B.n67 B.n66 585
R57 B.n65 B.n64 585
R58 B.n63 B.n62 585
R59 B.n61 B.n60 585
R60 B.n59 B.n58 585
R61 B.n57 B.n56 585
R62 B.n55 B.n54 585
R63 B.n33 B.n32 585
R64 B.n298 B.n297 585
R65 B.n291 B.n49 585
R66 B.n49 B.n30 585
R67 B.n290 B.n29 585
R68 B.n302 B.n29 585
R69 B.n289 B.n28 585
R70 B.n303 B.n28 585
R71 B.n288 B.n27 585
R72 B.n304 B.n27 585
R73 B.n287 B.n286 585
R74 B.n286 B.n26 585
R75 B.n285 B.n22 585
R76 B.n310 B.n22 585
R77 B.n284 B.n21 585
R78 B.n311 B.n21 585
R79 B.n283 B.n20 585
R80 B.n312 B.n20 585
R81 B.n282 B.n281 585
R82 B.n281 B.n16 585
R83 B.n280 B.n15 585
R84 B.n318 B.n15 585
R85 B.n279 B.n14 585
R86 B.n319 B.n14 585
R87 B.n278 B.n13 585
R88 B.n320 B.n13 585
R89 B.n277 B.n276 585
R90 B.n276 B.n12 585
R91 B.n275 B.n274 585
R92 B.n275 B.n8 585
R93 B.n273 B.n7 585
R94 B.n327 B.n7 585
R95 B.n272 B.n6 585
R96 B.n328 B.n6 585
R97 B.n271 B.n5 585
R98 B.n329 B.n5 585
R99 B.n270 B.n269 585
R100 B.n269 B.n4 585
R101 B.n268 B.n113 585
R102 B.n268 B.n267 585
R103 B.n257 B.n114 585
R104 B.n260 B.n114 585
R105 B.n259 B.n258 585
R106 B.n261 B.n259 585
R107 B.n256 B.n118 585
R108 B.n122 B.n118 585
R109 B.n255 B.n254 585
R110 B.n254 B.n253 585
R111 B.n120 B.n119 585
R112 B.n121 B.n120 585
R113 B.n246 B.n245 585
R114 B.n247 B.n246 585
R115 B.n244 B.n127 585
R116 B.n127 B.n126 585
R117 B.n243 B.n242 585
R118 B.n242 B.n241 585
R119 B.n129 B.n128 585
R120 B.n234 B.n129 585
R121 B.n233 B.n232 585
R122 B.n235 B.n233 585
R123 B.n231 B.n134 585
R124 B.n134 B.n133 585
R125 B.n230 B.n229 585
R126 B.n229 B.n228 585
R127 B.n136 B.n135 585
R128 B.n137 B.n136 585
R129 B.n224 B.n223 585
R130 B.n140 B.n139 585
R131 B.n220 B.n219 585
R132 B.n221 B.n220 585
R133 B.n218 B.n156 585
R134 B.n217 B.n216 585
R135 B.n215 B.n214 585
R136 B.n213 B.n212 585
R137 B.n211 B.n210 585
R138 B.n209 B.n208 585
R139 B.n207 B.n206 585
R140 B.n205 B.n204 585
R141 B.n203 B.n202 585
R142 B.n201 B.n200 585
R143 B.n199 B.n198 585
R144 B.n197 B.n196 585
R145 B.n195 B.n194 585
R146 B.n193 B.n192 585
R147 B.n191 B.n190 585
R148 B.n189 B.n188 585
R149 B.n187 B.n186 585
R150 B.n185 B.n184 585
R151 B.n183 B.n182 585
R152 B.n181 B.n180 585
R153 B.n179 B.n178 585
R154 B.n177 B.n176 585
R155 B.n175 B.n174 585
R156 B.n173 B.n172 585
R157 B.n171 B.n170 585
R158 B.n169 B.n168 585
R159 B.n167 B.n166 585
R160 B.n165 B.n164 585
R161 B.n163 B.n155 585
R162 B.n221 B.n155 585
R163 B.n225 B.n138 585
R164 B.n138 B.n137 585
R165 B.n227 B.n226 585
R166 B.n228 B.n227 585
R167 B.n132 B.n131 585
R168 B.n133 B.n132 585
R169 B.n237 B.n236 585
R170 B.n236 B.n235 585
R171 B.n238 B.n130 585
R172 B.n234 B.n130 585
R173 B.n240 B.n239 585
R174 B.n241 B.n240 585
R175 B.n125 B.n124 585
R176 B.n126 B.n125 585
R177 B.n249 B.n248 585
R178 B.n248 B.n247 585
R179 B.n250 B.n123 585
R180 B.n123 B.n121 585
R181 B.n252 B.n251 585
R182 B.n253 B.n252 585
R183 B.n117 B.n116 585
R184 B.n122 B.n117 585
R185 B.n263 B.n262 585
R186 B.n262 B.n261 585
R187 B.n264 B.n115 585
R188 B.n260 B.n115 585
R189 B.n266 B.n265 585
R190 B.n267 B.n266 585
R191 B.n3 B.n0 585
R192 B.n4 B.n3 585
R193 B.n326 B.n1 585
R194 B.n327 B.n326 585
R195 B.n325 B.n324 585
R196 B.n325 B.n8 585
R197 B.n323 B.n9 585
R198 B.n12 B.n9 585
R199 B.n322 B.n321 585
R200 B.n321 B.n320 585
R201 B.n11 B.n10 585
R202 B.n319 B.n11 585
R203 B.n317 B.n316 585
R204 B.n318 B.n317 585
R205 B.n315 B.n17 585
R206 B.n17 B.n16 585
R207 B.n314 B.n313 585
R208 B.n313 B.n312 585
R209 B.n19 B.n18 585
R210 B.n311 B.n19 585
R211 B.n309 B.n308 585
R212 B.n310 B.n309 585
R213 B.n307 B.n23 585
R214 B.n26 B.n23 585
R215 B.n306 B.n305 585
R216 B.n305 B.n304 585
R217 B.n25 B.n24 585
R218 B.n303 B.n25 585
R219 B.n301 B.n300 585
R220 B.n302 B.n301 585
R221 B.n299 B.n31 585
R222 B.n31 B.n30 585
R223 B.n330 B.n329 585
R224 B.n328 B.n2 585
R225 B.n297 B.n31 449.257
R226 B.n293 B.n49 449.257
R227 B.n155 B.n136 449.257
R228 B.n223 B.n138 449.257
R229 B.n50 B.t4 286.57
R230 B.n160 B.t15 286.57
R231 B.n52 B.t8 286.332
R232 B.n157 B.t11 286.332
R233 B.n295 B.n294 256.663
R234 B.n295 B.n47 256.663
R235 B.n295 B.n46 256.663
R236 B.n295 B.n45 256.663
R237 B.n295 B.n44 256.663
R238 B.n295 B.n43 256.663
R239 B.n295 B.n42 256.663
R240 B.n295 B.n41 256.663
R241 B.n295 B.n40 256.663
R242 B.n295 B.n39 256.663
R243 B.n295 B.n38 256.663
R244 B.n295 B.n37 256.663
R245 B.n295 B.n36 256.663
R246 B.n295 B.n35 256.663
R247 B.n295 B.n34 256.663
R248 B.n296 B.n295 256.663
R249 B.n222 B.n221 256.663
R250 B.n221 B.n141 256.663
R251 B.n221 B.n142 256.663
R252 B.n221 B.n143 256.663
R253 B.n221 B.n144 256.663
R254 B.n221 B.n145 256.663
R255 B.n221 B.n146 256.663
R256 B.n221 B.n147 256.663
R257 B.n221 B.n148 256.663
R258 B.n221 B.n149 256.663
R259 B.n221 B.n150 256.663
R260 B.n221 B.n151 256.663
R261 B.n221 B.n152 256.663
R262 B.n221 B.n153 256.663
R263 B.n221 B.n154 256.663
R264 B.n332 B.n331 256.663
R265 B.n221 B.n137 180.537
R266 B.n295 B.n30 180.537
R267 B.n54 B.n33 163.367
R268 B.n58 B.n57 163.367
R269 B.n62 B.n61 163.367
R270 B.n66 B.n65 163.367
R271 B.n70 B.n69 163.367
R272 B.n75 B.n74 163.367
R273 B.n79 B.n78 163.367
R274 B.n83 B.n82 163.367
R275 B.n87 B.n86 163.367
R276 B.n91 B.n90 163.367
R277 B.n96 B.n95 163.367
R278 B.n100 B.n99 163.367
R279 B.n104 B.n103 163.367
R280 B.n108 B.n107 163.367
R281 B.n110 B.n48 163.367
R282 B.n229 B.n136 163.367
R283 B.n229 B.n134 163.367
R284 B.n233 B.n134 163.367
R285 B.n233 B.n129 163.367
R286 B.n242 B.n129 163.367
R287 B.n242 B.n127 163.367
R288 B.n246 B.n127 163.367
R289 B.n246 B.n120 163.367
R290 B.n254 B.n120 163.367
R291 B.n254 B.n118 163.367
R292 B.n259 B.n118 163.367
R293 B.n259 B.n114 163.367
R294 B.n268 B.n114 163.367
R295 B.n269 B.n268 163.367
R296 B.n269 B.n5 163.367
R297 B.n6 B.n5 163.367
R298 B.n7 B.n6 163.367
R299 B.n275 B.n7 163.367
R300 B.n276 B.n275 163.367
R301 B.n276 B.n13 163.367
R302 B.n14 B.n13 163.367
R303 B.n15 B.n14 163.367
R304 B.n281 B.n15 163.367
R305 B.n281 B.n20 163.367
R306 B.n21 B.n20 163.367
R307 B.n22 B.n21 163.367
R308 B.n286 B.n22 163.367
R309 B.n286 B.n27 163.367
R310 B.n28 B.n27 163.367
R311 B.n29 B.n28 163.367
R312 B.n49 B.n29 163.367
R313 B.n220 B.n140 163.367
R314 B.n220 B.n156 163.367
R315 B.n216 B.n215 163.367
R316 B.n212 B.n211 163.367
R317 B.n208 B.n207 163.367
R318 B.n204 B.n203 163.367
R319 B.n200 B.n199 163.367
R320 B.n196 B.n195 163.367
R321 B.n192 B.n191 163.367
R322 B.n188 B.n187 163.367
R323 B.n184 B.n183 163.367
R324 B.n180 B.n179 163.367
R325 B.n176 B.n175 163.367
R326 B.n172 B.n171 163.367
R327 B.n168 B.n167 163.367
R328 B.n164 B.n155 163.367
R329 B.n227 B.n138 163.367
R330 B.n227 B.n132 163.367
R331 B.n236 B.n132 163.367
R332 B.n236 B.n130 163.367
R333 B.n240 B.n130 163.367
R334 B.n240 B.n125 163.367
R335 B.n248 B.n125 163.367
R336 B.n248 B.n123 163.367
R337 B.n252 B.n123 163.367
R338 B.n252 B.n117 163.367
R339 B.n262 B.n117 163.367
R340 B.n262 B.n115 163.367
R341 B.n266 B.n115 163.367
R342 B.n266 B.n3 163.367
R343 B.n330 B.n3 163.367
R344 B.n326 B.n2 163.367
R345 B.n326 B.n325 163.367
R346 B.n325 B.n9 163.367
R347 B.n321 B.n9 163.367
R348 B.n321 B.n11 163.367
R349 B.n317 B.n11 163.367
R350 B.n317 B.n17 163.367
R351 B.n313 B.n17 163.367
R352 B.n313 B.n19 163.367
R353 B.n309 B.n19 163.367
R354 B.n309 B.n23 163.367
R355 B.n305 B.n23 163.367
R356 B.n305 B.n25 163.367
R357 B.n301 B.n25 163.367
R358 B.n301 B.n31 163.367
R359 B.n50 B.t6 124.668
R360 B.n160 B.t17 124.668
R361 B.n52 B.t9 124.668
R362 B.n157 B.t14 124.668
R363 B.n51 B.t7 108.764
R364 B.n161 B.t16 108.764
R365 B.n53 B.t10 108.764
R366 B.n158 B.t13 108.764
R367 B.n228 B.n137 108.642
R368 B.n228 B.n133 108.642
R369 B.n235 B.n133 108.642
R370 B.n235 B.n234 108.642
R371 B.n241 B.n126 108.642
R372 B.n247 B.n126 108.642
R373 B.n247 B.n121 108.642
R374 B.n253 B.n121 108.642
R375 B.n253 B.n122 108.642
R376 B.n261 B.n260 108.642
R377 B.n267 B.n4 108.642
R378 B.n329 B.n4 108.642
R379 B.n329 B.n328 108.642
R380 B.n328 B.n327 108.642
R381 B.n327 B.n8 108.642
R382 B.n320 B.n12 108.642
R383 B.n319 B.n318 108.642
R384 B.n318 B.n16 108.642
R385 B.n312 B.n16 108.642
R386 B.n312 B.n311 108.642
R387 B.n311 B.n310 108.642
R388 B.n304 B.n26 108.642
R389 B.n304 B.n303 108.642
R390 B.n303 B.n302 108.642
R391 B.n302 B.n30 108.642
R392 B.n261 B.t3 78.2866
R393 B.n320 B.t2 78.2866
R394 B.n260 B.t0 75.0913
R395 B.n12 B.t1 75.0913
R396 B.n234 B.t12 71.8959
R397 B.n26 B.t5 71.8959
R398 B.n297 B.n296 71.676
R399 B.n54 B.n34 71.676
R400 B.n58 B.n35 71.676
R401 B.n62 B.n36 71.676
R402 B.n66 B.n37 71.676
R403 B.n70 B.n38 71.676
R404 B.n75 B.n39 71.676
R405 B.n79 B.n40 71.676
R406 B.n83 B.n41 71.676
R407 B.n87 B.n42 71.676
R408 B.n91 B.n43 71.676
R409 B.n96 B.n44 71.676
R410 B.n100 B.n45 71.676
R411 B.n104 B.n46 71.676
R412 B.n108 B.n47 71.676
R413 B.n294 B.n48 71.676
R414 B.n294 B.n293 71.676
R415 B.n110 B.n47 71.676
R416 B.n107 B.n46 71.676
R417 B.n103 B.n45 71.676
R418 B.n99 B.n44 71.676
R419 B.n95 B.n43 71.676
R420 B.n90 B.n42 71.676
R421 B.n86 B.n41 71.676
R422 B.n82 B.n40 71.676
R423 B.n78 B.n39 71.676
R424 B.n74 B.n38 71.676
R425 B.n69 B.n37 71.676
R426 B.n65 B.n36 71.676
R427 B.n61 B.n35 71.676
R428 B.n57 B.n34 71.676
R429 B.n296 B.n33 71.676
R430 B.n223 B.n222 71.676
R431 B.n156 B.n141 71.676
R432 B.n215 B.n142 71.676
R433 B.n211 B.n143 71.676
R434 B.n207 B.n144 71.676
R435 B.n203 B.n145 71.676
R436 B.n199 B.n146 71.676
R437 B.n195 B.n147 71.676
R438 B.n191 B.n148 71.676
R439 B.n187 B.n149 71.676
R440 B.n183 B.n150 71.676
R441 B.n179 B.n151 71.676
R442 B.n175 B.n152 71.676
R443 B.n171 B.n153 71.676
R444 B.n167 B.n154 71.676
R445 B.n222 B.n140 71.676
R446 B.n216 B.n141 71.676
R447 B.n212 B.n142 71.676
R448 B.n208 B.n143 71.676
R449 B.n204 B.n144 71.676
R450 B.n200 B.n145 71.676
R451 B.n196 B.n146 71.676
R452 B.n192 B.n147 71.676
R453 B.n188 B.n148 71.676
R454 B.n184 B.n149 71.676
R455 B.n180 B.n150 71.676
R456 B.n176 B.n151 71.676
R457 B.n172 B.n152 71.676
R458 B.n168 B.n153 71.676
R459 B.n164 B.n154 71.676
R460 B.n331 B.n330 71.676
R461 B.n331 B.n2 71.676
R462 B.n72 B.n53 59.5399
R463 B.n93 B.n51 59.5399
R464 B.n162 B.n161 59.5399
R465 B.n159 B.n158 59.5399
R466 B.n241 B.t12 36.7471
R467 B.n310 B.t5 36.7471
R468 B.n267 B.t0 33.5517
R469 B.t1 B.n8 33.5517
R470 B.n122 B.t3 30.3563
R471 B.t2 B.n319 30.3563
R472 B.n225 B.n224 29.1907
R473 B.n163 B.n135 29.1907
R474 B.n292 B.n291 29.1907
R475 B.n299 B.n298 29.1907
R476 B B.n332 18.0485
R477 B.n53 B.n52 15.9035
R478 B.n51 B.n50 15.9035
R479 B.n161 B.n160 15.9035
R480 B.n158 B.n157 15.9035
R481 B.n226 B.n225 10.6151
R482 B.n226 B.n131 10.6151
R483 B.n237 B.n131 10.6151
R484 B.n238 B.n237 10.6151
R485 B.n239 B.n238 10.6151
R486 B.n239 B.n124 10.6151
R487 B.n249 B.n124 10.6151
R488 B.n250 B.n249 10.6151
R489 B.n251 B.n250 10.6151
R490 B.n251 B.n116 10.6151
R491 B.n263 B.n116 10.6151
R492 B.n264 B.n263 10.6151
R493 B.n265 B.n264 10.6151
R494 B.n265 B.n0 10.6151
R495 B.n224 B.n139 10.6151
R496 B.n219 B.n139 10.6151
R497 B.n219 B.n218 10.6151
R498 B.n218 B.n217 10.6151
R499 B.n217 B.n214 10.6151
R500 B.n214 B.n213 10.6151
R501 B.n213 B.n210 10.6151
R502 B.n210 B.n209 10.6151
R503 B.n209 B.n206 10.6151
R504 B.n206 B.n205 10.6151
R505 B.n202 B.n201 10.6151
R506 B.n201 B.n198 10.6151
R507 B.n198 B.n197 10.6151
R508 B.n197 B.n194 10.6151
R509 B.n194 B.n193 10.6151
R510 B.n193 B.n190 10.6151
R511 B.n190 B.n189 10.6151
R512 B.n189 B.n186 10.6151
R513 B.n186 B.n185 10.6151
R514 B.n182 B.n181 10.6151
R515 B.n181 B.n178 10.6151
R516 B.n178 B.n177 10.6151
R517 B.n177 B.n174 10.6151
R518 B.n174 B.n173 10.6151
R519 B.n173 B.n170 10.6151
R520 B.n170 B.n169 10.6151
R521 B.n169 B.n166 10.6151
R522 B.n166 B.n165 10.6151
R523 B.n165 B.n163 10.6151
R524 B.n230 B.n135 10.6151
R525 B.n231 B.n230 10.6151
R526 B.n232 B.n231 10.6151
R527 B.n232 B.n128 10.6151
R528 B.n243 B.n128 10.6151
R529 B.n244 B.n243 10.6151
R530 B.n245 B.n244 10.6151
R531 B.n245 B.n119 10.6151
R532 B.n255 B.n119 10.6151
R533 B.n256 B.n255 10.6151
R534 B.n258 B.n256 10.6151
R535 B.n258 B.n257 10.6151
R536 B.n257 B.n113 10.6151
R537 B.n270 B.n113 10.6151
R538 B.n271 B.n270 10.6151
R539 B.n272 B.n271 10.6151
R540 B.n273 B.n272 10.6151
R541 B.n274 B.n273 10.6151
R542 B.n277 B.n274 10.6151
R543 B.n278 B.n277 10.6151
R544 B.n279 B.n278 10.6151
R545 B.n280 B.n279 10.6151
R546 B.n282 B.n280 10.6151
R547 B.n283 B.n282 10.6151
R548 B.n284 B.n283 10.6151
R549 B.n285 B.n284 10.6151
R550 B.n287 B.n285 10.6151
R551 B.n288 B.n287 10.6151
R552 B.n289 B.n288 10.6151
R553 B.n290 B.n289 10.6151
R554 B.n291 B.n290 10.6151
R555 B.n324 B.n1 10.6151
R556 B.n324 B.n323 10.6151
R557 B.n323 B.n322 10.6151
R558 B.n322 B.n10 10.6151
R559 B.n316 B.n10 10.6151
R560 B.n316 B.n315 10.6151
R561 B.n315 B.n314 10.6151
R562 B.n314 B.n18 10.6151
R563 B.n308 B.n18 10.6151
R564 B.n308 B.n307 10.6151
R565 B.n307 B.n306 10.6151
R566 B.n306 B.n24 10.6151
R567 B.n300 B.n24 10.6151
R568 B.n300 B.n299 10.6151
R569 B.n298 B.n32 10.6151
R570 B.n55 B.n32 10.6151
R571 B.n56 B.n55 10.6151
R572 B.n59 B.n56 10.6151
R573 B.n60 B.n59 10.6151
R574 B.n63 B.n60 10.6151
R575 B.n64 B.n63 10.6151
R576 B.n67 B.n64 10.6151
R577 B.n68 B.n67 10.6151
R578 B.n71 B.n68 10.6151
R579 B.n76 B.n73 10.6151
R580 B.n77 B.n76 10.6151
R581 B.n80 B.n77 10.6151
R582 B.n81 B.n80 10.6151
R583 B.n84 B.n81 10.6151
R584 B.n85 B.n84 10.6151
R585 B.n88 B.n85 10.6151
R586 B.n89 B.n88 10.6151
R587 B.n92 B.n89 10.6151
R588 B.n97 B.n94 10.6151
R589 B.n98 B.n97 10.6151
R590 B.n101 B.n98 10.6151
R591 B.n102 B.n101 10.6151
R592 B.n105 B.n102 10.6151
R593 B.n106 B.n105 10.6151
R594 B.n109 B.n106 10.6151
R595 B.n111 B.n109 10.6151
R596 B.n112 B.n111 10.6151
R597 B.n292 B.n112 10.6151
R598 B.n205 B.n159 9.52245
R599 B.n182 B.n162 9.52245
R600 B.n72 B.n71 9.52245
R601 B.n94 B.n93 9.52245
R602 B.n332 B.n0 8.11757
R603 B.n332 B.n1 8.11757
R604 B.n202 B.n159 1.09318
R605 B.n185 B.n162 1.09318
R606 B.n73 B.n72 1.09318
R607 B.n93 B.n92 1.09318
R608 VN.n0 VN.t1 180.829
R609 VN.n1 VN.t2 180.829
R610 VN.n0 VN.t0 180.804
R611 VN.n1 VN.t3 180.804
R612 VN VN.n1 102.526
R613 VN VN.n0 70.265
R614 VDD2.n2 VDD2.n0 142.618
R615 VDD2.n2 VDD2.n1 115.394
R616 VDD2.n1 VDD2.t0 12.2986
R617 VDD2.n1 VDD2.t1 12.2986
R618 VDD2.n0 VDD2.t2 12.2986
R619 VDD2.n0 VDD2.t3 12.2986
R620 VDD2 VDD2.n2 0.0586897
C0 VP VDD1 0.711978f
C1 VTAIL VDD2 2.25665f
C2 VTAIL VN 0.682286f
C3 VDD2 VN 0.599259f
C4 VTAIL VP 0.696393f
C5 VTAIL VDD1 2.21659f
C6 VP VDD2 0.267117f
C7 VDD2 VDD1 0.521669f
C8 VP VN 2.75529f
C9 VDD1 VN 0.153381f
C10 VDD2 B 1.745034f
C11 VDD1 B 3.5001f
C12 VTAIL B 2.597132f
C13 VN B 5.47779f
C14 VP B 3.597478f
C15 VDD2.t2 B 0.028034f
C16 VDD2.t3 B 0.028034f
C17 VDD2.n0 B 0.2962f
C18 VDD2.t0 B 0.028034f
C19 VDD2.t1 B 0.028034f
C20 VDD2.n1 B 0.161003f
C21 VDD2.n2 B 1.67573f
C22 VN.t1 B 0.105434f
C23 VN.t0 B 0.105418f
C24 VN.n0 B 0.137867f
C25 VN.t2 B 0.105434f
C26 VN.t3 B 0.105418f
C27 VN.n1 B 0.461896f
C28 VDD1.t1 B 0.025899f
C29 VDD1.t0 B 0.025899f
C30 VDD1.n0 B 0.148845f
C31 VDD1.t2 B 0.025899f
C32 VDD1.t3 B 0.025899f
C33 VDD1.n1 B 0.283768f
C34 VTAIL.t1 B 0.16237f
C35 VTAIL.n0 B 0.205612f
C36 VTAIL.t7 B 0.16237f
C37 VTAIL.n1 B 0.223473f
C38 VTAIL.t5 B 0.16237f
C39 VTAIL.n2 B 0.576786f
C40 VTAIL.t3 B 0.162371f
C41 VTAIL.n3 B 0.576786f
C42 VTAIL.t0 B 0.162371f
C43 VTAIL.n4 B 0.223472f
C44 VTAIL.t6 B 0.162371f
C45 VTAIL.n5 B 0.223472f
C46 VTAIL.t4 B 0.162371f
C47 VTAIL.n6 B 0.576786f
C48 VTAIL.t2 B 0.16237f
C49 VTAIL.n7 B 0.551885f
C50 VP.t3 B 0.107503f
C51 VP.t2 B 0.107519f
C52 VP.n0 B 0.460109f
C53 VP.n1 B 1.72243f
C54 VP.t1 B 0.098293f
C55 VP.n2 B 0.07946f
C56 VP.t0 B 0.098293f
C57 VP.n3 B 0.07946f
C58 VP.n4 B 0.030535f
.ends

