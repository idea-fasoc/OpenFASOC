* NGSPICE file created from diff_pair_sample_1313.ext - technology: sky130A

.subckt diff_pair_sample_1313 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5171 pd=8.56 as=0.64185 ps=4.22 w=3.89 l=1.85
X1 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5171 pd=8.56 as=0.64185 ps=4.22 w=3.89 l=1.85
X2 VDD1.t4 VP.t1 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.64185 pd=4.22 as=1.5171 ps=8.56 w=3.89 l=1.85
X3 VTAIL.t10 VP.t2 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.64185 pd=4.22 as=0.64185 ps=4.22 w=3.89 l=1.85
X4 VDD2.t4 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.64185 pd=4.22 as=1.5171 ps=8.56 w=3.89 l=1.85
X5 VDD2.t3 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5171 pd=8.56 as=0.64185 ps=4.22 w=3.89 l=1.85
X6 VTAIL.t1 VN.t3 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.64185 pd=4.22 as=0.64185 ps=4.22 w=3.89 l=1.85
X7 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5171 pd=8.56 as=0 ps=0 w=3.89 l=1.85
X8 VDD2.t1 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.64185 pd=4.22 as=1.5171 ps=8.56 w=3.89 l=1.85
X9 VDD1.t2 VP.t3 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=0.64185 pd=4.22 as=1.5171 ps=8.56 w=3.89 l=1.85
X10 VTAIL.t2 VN.t5 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.64185 pd=4.22 as=0.64185 ps=4.22 w=3.89 l=1.85
X11 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5171 pd=8.56 as=0 ps=0 w=3.89 l=1.85
X12 VTAIL.t8 VP.t4 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.64185 pd=4.22 as=0.64185 ps=4.22 w=3.89 l=1.85
X13 VDD1.t0 VP.t5 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5171 pd=8.56 as=0.64185 ps=4.22 w=3.89 l=1.85
X14 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.5171 pd=8.56 as=0 ps=0 w=3.89 l=1.85
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5171 pd=8.56 as=0 ps=0 w=3.89 l=1.85
R0 VP.n9 VP.n8 161.3
R1 VP.n10 VP.n5 161.3
R2 VP.n12 VP.n11 161.3
R3 VP.n13 VP.n4 161.3
R4 VP.n30 VP.n0 161.3
R5 VP.n29 VP.n28 161.3
R6 VP.n27 VP.n1 161.3
R7 VP.n26 VP.n25 161.3
R8 VP.n23 VP.n2 161.3
R9 VP.n22 VP.n21 161.3
R10 VP.n20 VP.n3 161.3
R11 VP.n19 VP.n18 161.3
R12 VP.n17 VP.n16 89.7148
R13 VP.n32 VP.n31 89.7148
R14 VP.n15 VP.n14 89.7148
R15 VP.n6 VP.t0 81.2706
R16 VP.n7 VP.n6 57.6865
R17 VP.n22 VP.n3 56.0336
R18 VP.n29 VP.n1 56.0336
R19 VP.n12 VP.n5 56.0336
R20 VP.n17 VP.t5 50.6756
R21 VP.n24 VP.t4 50.6756
R22 VP.n31 VP.t3 50.6756
R23 VP.n14 VP.t1 50.6756
R24 VP.n7 VP.t2 50.6756
R25 VP.n16 VP.n15 39.5981
R26 VP.n18 VP.n3 24.9531
R27 VP.n30 VP.n29 24.9531
R28 VP.n13 VP.n12 24.9531
R29 VP.n23 VP.n22 24.4675
R30 VP.n25 VP.n1 24.4675
R31 VP.n8 VP.n5 24.4675
R32 VP.n18 VP.n17 21.0421
R33 VP.n31 VP.n30 21.0421
R34 VP.n14 VP.n13 21.0421
R35 VP.n9 VP.n6 13.151
R36 VP.n24 VP.n23 12.234
R37 VP.n25 VP.n24 12.234
R38 VP.n8 VP.n7 12.234
R39 VP.n15 VP.n4 0.278367
R40 VP.n19 VP.n16 0.278367
R41 VP.n32 VP.n0 0.278367
R42 VP.n10 VP.n9 0.189894
R43 VP.n11 VP.n10 0.189894
R44 VP.n11 VP.n4 0.189894
R45 VP.n20 VP.n19 0.189894
R46 VP.n21 VP.n20 0.189894
R47 VP.n21 VP.n2 0.189894
R48 VP.n26 VP.n2 0.189894
R49 VP.n27 VP.n26 0.189894
R50 VP.n28 VP.n27 0.189894
R51 VP.n28 VP.n0 0.189894
R52 VP VP.n32 0.153454
R53 VTAIL.n82 VTAIL.n68 289.615
R54 VTAIL.n16 VTAIL.n2 289.615
R55 VTAIL.n62 VTAIL.n48 289.615
R56 VTAIL.n40 VTAIL.n26 289.615
R57 VTAIL.n75 VTAIL.n74 185
R58 VTAIL.n72 VTAIL.n71 185
R59 VTAIL.n81 VTAIL.n80 185
R60 VTAIL.n83 VTAIL.n82 185
R61 VTAIL.n9 VTAIL.n8 185
R62 VTAIL.n6 VTAIL.n5 185
R63 VTAIL.n15 VTAIL.n14 185
R64 VTAIL.n17 VTAIL.n16 185
R65 VTAIL.n63 VTAIL.n62 185
R66 VTAIL.n61 VTAIL.n60 185
R67 VTAIL.n52 VTAIL.n51 185
R68 VTAIL.n55 VTAIL.n54 185
R69 VTAIL.n41 VTAIL.n40 185
R70 VTAIL.n39 VTAIL.n38 185
R71 VTAIL.n30 VTAIL.n29 185
R72 VTAIL.n33 VTAIL.n32 185
R73 VTAIL.t5 VTAIL.n73 147.888
R74 VTAIL.t9 VTAIL.n7 147.888
R75 VTAIL.t6 VTAIL.n53 147.888
R76 VTAIL.t4 VTAIL.n31 147.888
R77 VTAIL.n74 VTAIL.n71 104.615
R78 VTAIL.n81 VTAIL.n71 104.615
R79 VTAIL.n82 VTAIL.n81 104.615
R80 VTAIL.n8 VTAIL.n5 104.615
R81 VTAIL.n15 VTAIL.n5 104.615
R82 VTAIL.n16 VTAIL.n15 104.615
R83 VTAIL.n62 VTAIL.n61 104.615
R84 VTAIL.n61 VTAIL.n51 104.615
R85 VTAIL.n54 VTAIL.n51 104.615
R86 VTAIL.n40 VTAIL.n39 104.615
R87 VTAIL.n39 VTAIL.n29 104.615
R88 VTAIL.n32 VTAIL.n29 104.615
R89 VTAIL.n47 VTAIL.n46 57.755
R90 VTAIL.n25 VTAIL.n24 57.755
R91 VTAIL.n1 VTAIL.n0 57.7549
R92 VTAIL.n23 VTAIL.n22 57.7549
R93 VTAIL.n74 VTAIL.t5 52.3082
R94 VTAIL.n8 VTAIL.t9 52.3082
R95 VTAIL.n54 VTAIL.t6 52.3082
R96 VTAIL.n32 VTAIL.t4 52.3082
R97 VTAIL.n87 VTAIL.n86 33.155
R98 VTAIL.n21 VTAIL.n20 33.155
R99 VTAIL.n67 VTAIL.n66 33.155
R100 VTAIL.n45 VTAIL.n44 33.155
R101 VTAIL.n25 VTAIL.n23 19.4789
R102 VTAIL.n87 VTAIL.n67 17.5996
R103 VTAIL.n75 VTAIL.n73 15.6496
R104 VTAIL.n9 VTAIL.n7 15.6496
R105 VTAIL.n55 VTAIL.n53 15.6496
R106 VTAIL.n33 VTAIL.n31 15.6496
R107 VTAIL.n76 VTAIL.n72 12.8005
R108 VTAIL.n10 VTAIL.n6 12.8005
R109 VTAIL.n56 VTAIL.n52 12.8005
R110 VTAIL.n34 VTAIL.n30 12.8005
R111 VTAIL.n80 VTAIL.n79 12.0247
R112 VTAIL.n14 VTAIL.n13 12.0247
R113 VTAIL.n60 VTAIL.n59 12.0247
R114 VTAIL.n38 VTAIL.n37 12.0247
R115 VTAIL.n83 VTAIL.n70 11.249
R116 VTAIL.n17 VTAIL.n4 11.249
R117 VTAIL.n63 VTAIL.n50 11.249
R118 VTAIL.n41 VTAIL.n28 11.249
R119 VTAIL.n84 VTAIL.n68 10.4732
R120 VTAIL.n18 VTAIL.n2 10.4732
R121 VTAIL.n64 VTAIL.n48 10.4732
R122 VTAIL.n42 VTAIL.n26 10.4732
R123 VTAIL.n86 VTAIL.n85 9.45567
R124 VTAIL.n20 VTAIL.n19 9.45567
R125 VTAIL.n66 VTAIL.n65 9.45567
R126 VTAIL.n44 VTAIL.n43 9.45567
R127 VTAIL.n85 VTAIL.n84 9.3005
R128 VTAIL.n70 VTAIL.n69 9.3005
R129 VTAIL.n79 VTAIL.n78 9.3005
R130 VTAIL.n77 VTAIL.n76 9.3005
R131 VTAIL.n19 VTAIL.n18 9.3005
R132 VTAIL.n4 VTAIL.n3 9.3005
R133 VTAIL.n13 VTAIL.n12 9.3005
R134 VTAIL.n11 VTAIL.n10 9.3005
R135 VTAIL.n65 VTAIL.n64 9.3005
R136 VTAIL.n50 VTAIL.n49 9.3005
R137 VTAIL.n59 VTAIL.n58 9.3005
R138 VTAIL.n57 VTAIL.n56 9.3005
R139 VTAIL.n43 VTAIL.n42 9.3005
R140 VTAIL.n28 VTAIL.n27 9.3005
R141 VTAIL.n37 VTAIL.n36 9.3005
R142 VTAIL.n35 VTAIL.n34 9.3005
R143 VTAIL.n0 VTAIL.t0 5.09047
R144 VTAIL.n0 VTAIL.t1 5.09047
R145 VTAIL.n22 VTAIL.t7 5.09047
R146 VTAIL.n22 VTAIL.t8 5.09047
R147 VTAIL.n46 VTAIL.t11 5.09047
R148 VTAIL.n46 VTAIL.t10 5.09047
R149 VTAIL.n24 VTAIL.t3 5.09047
R150 VTAIL.n24 VTAIL.t2 5.09047
R151 VTAIL.n77 VTAIL.n73 4.40546
R152 VTAIL.n11 VTAIL.n7 4.40546
R153 VTAIL.n57 VTAIL.n53 4.40546
R154 VTAIL.n35 VTAIL.n31 4.40546
R155 VTAIL.n86 VTAIL.n68 3.49141
R156 VTAIL.n20 VTAIL.n2 3.49141
R157 VTAIL.n66 VTAIL.n48 3.49141
R158 VTAIL.n44 VTAIL.n26 3.49141
R159 VTAIL.n84 VTAIL.n83 2.71565
R160 VTAIL.n18 VTAIL.n17 2.71565
R161 VTAIL.n64 VTAIL.n63 2.71565
R162 VTAIL.n42 VTAIL.n41 2.71565
R163 VTAIL.n80 VTAIL.n70 1.93989
R164 VTAIL.n14 VTAIL.n4 1.93989
R165 VTAIL.n60 VTAIL.n50 1.93989
R166 VTAIL.n38 VTAIL.n28 1.93989
R167 VTAIL.n45 VTAIL.n25 1.87981
R168 VTAIL.n67 VTAIL.n47 1.87981
R169 VTAIL.n23 VTAIL.n21 1.87981
R170 VTAIL.n47 VTAIL.n45 1.40998
R171 VTAIL.n21 VTAIL.n1 1.40998
R172 VTAIL VTAIL.n87 1.35179
R173 VTAIL.n79 VTAIL.n72 1.16414
R174 VTAIL.n13 VTAIL.n6 1.16414
R175 VTAIL.n59 VTAIL.n52 1.16414
R176 VTAIL.n37 VTAIL.n30 1.16414
R177 VTAIL VTAIL.n1 0.528517
R178 VTAIL.n76 VTAIL.n75 0.388379
R179 VTAIL.n10 VTAIL.n9 0.388379
R180 VTAIL.n56 VTAIL.n55 0.388379
R181 VTAIL.n34 VTAIL.n33 0.388379
R182 VTAIL.n78 VTAIL.n77 0.155672
R183 VTAIL.n78 VTAIL.n69 0.155672
R184 VTAIL.n85 VTAIL.n69 0.155672
R185 VTAIL.n12 VTAIL.n11 0.155672
R186 VTAIL.n12 VTAIL.n3 0.155672
R187 VTAIL.n19 VTAIL.n3 0.155672
R188 VTAIL.n65 VTAIL.n49 0.155672
R189 VTAIL.n58 VTAIL.n49 0.155672
R190 VTAIL.n58 VTAIL.n57 0.155672
R191 VTAIL.n43 VTAIL.n27 0.155672
R192 VTAIL.n36 VTAIL.n27 0.155672
R193 VTAIL.n36 VTAIL.n35 0.155672
R194 VDD1.n14 VDD1.n0 289.615
R195 VDD1.n33 VDD1.n19 289.615
R196 VDD1.n15 VDD1.n14 185
R197 VDD1.n13 VDD1.n12 185
R198 VDD1.n4 VDD1.n3 185
R199 VDD1.n7 VDD1.n6 185
R200 VDD1.n26 VDD1.n25 185
R201 VDD1.n23 VDD1.n22 185
R202 VDD1.n32 VDD1.n31 185
R203 VDD1.n34 VDD1.n33 185
R204 VDD1.t5 VDD1.n5 147.888
R205 VDD1.t0 VDD1.n24 147.888
R206 VDD1.n14 VDD1.n13 104.615
R207 VDD1.n13 VDD1.n3 104.615
R208 VDD1.n6 VDD1.n3 104.615
R209 VDD1.n25 VDD1.n22 104.615
R210 VDD1.n32 VDD1.n22 104.615
R211 VDD1.n33 VDD1.n32 104.615
R212 VDD1.n39 VDD1.n38 74.8481
R213 VDD1.n41 VDD1.n40 74.4337
R214 VDD1.n6 VDD1.t5 52.3082
R215 VDD1.n25 VDD1.t0 52.3082
R216 VDD1 VDD1.n18 51.3015
R217 VDD1.n39 VDD1.n37 51.188
R218 VDD1.n41 VDD1.n39 34.6992
R219 VDD1.n7 VDD1.n5 15.6496
R220 VDD1.n26 VDD1.n24 15.6496
R221 VDD1.n8 VDD1.n4 12.8005
R222 VDD1.n27 VDD1.n23 12.8005
R223 VDD1.n12 VDD1.n11 12.0247
R224 VDD1.n31 VDD1.n30 12.0247
R225 VDD1.n15 VDD1.n2 11.249
R226 VDD1.n34 VDD1.n21 11.249
R227 VDD1.n16 VDD1.n0 10.4732
R228 VDD1.n35 VDD1.n19 10.4732
R229 VDD1.n18 VDD1.n17 9.45567
R230 VDD1.n37 VDD1.n36 9.45567
R231 VDD1.n17 VDD1.n16 9.3005
R232 VDD1.n2 VDD1.n1 9.3005
R233 VDD1.n11 VDD1.n10 9.3005
R234 VDD1.n9 VDD1.n8 9.3005
R235 VDD1.n36 VDD1.n35 9.3005
R236 VDD1.n21 VDD1.n20 9.3005
R237 VDD1.n30 VDD1.n29 9.3005
R238 VDD1.n28 VDD1.n27 9.3005
R239 VDD1.n40 VDD1.t3 5.09047
R240 VDD1.n40 VDD1.t4 5.09047
R241 VDD1.n38 VDD1.t1 5.09047
R242 VDD1.n38 VDD1.t2 5.09047
R243 VDD1.n9 VDD1.n5 4.40546
R244 VDD1.n28 VDD1.n24 4.40546
R245 VDD1.n18 VDD1.n0 3.49141
R246 VDD1.n37 VDD1.n19 3.49141
R247 VDD1.n16 VDD1.n15 2.71565
R248 VDD1.n35 VDD1.n34 2.71565
R249 VDD1.n12 VDD1.n2 1.93989
R250 VDD1.n31 VDD1.n21 1.93989
R251 VDD1.n11 VDD1.n4 1.16414
R252 VDD1.n30 VDD1.n23 1.16414
R253 VDD1 VDD1.n41 0.412138
R254 VDD1.n8 VDD1.n7 0.388379
R255 VDD1.n27 VDD1.n26 0.388379
R256 VDD1.n17 VDD1.n1 0.155672
R257 VDD1.n10 VDD1.n1 0.155672
R258 VDD1.n10 VDD1.n9 0.155672
R259 VDD1.n29 VDD1.n28 0.155672
R260 VDD1.n29 VDD1.n20 0.155672
R261 VDD1.n36 VDD1.n20 0.155672
R262 B.n506 B.n505 585
R263 B.n507 B.n506 585
R264 B.n179 B.n86 585
R265 B.n178 B.n177 585
R266 B.n176 B.n175 585
R267 B.n174 B.n173 585
R268 B.n172 B.n171 585
R269 B.n170 B.n169 585
R270 B.n168 B.n167 585
R271 B.n166 B.n165 585
R272 B.n164 B.n163 585
R273 B.n162 B.n161 585
R274 B.n160 B.n159 585
R275 B.n158 B.n157 585
R276 B.n156 B.n155 585
R277 B.n154 B.n153 585
R278 B.n152 B.n151 585
R279 B.n150 B.n149 585
R280 B.n148 B.n147 585
R281 B.n145 B.n144 585
R282 B.n143 B.n142 585
R283 B.n141 B.n140 585
R284 B.n139 B.n138 585
R285 B.n137 B.n136 585
R286 B.n135 B.n134 585
R287 B.n133 B.n132 585
R288 B.n131 B.n130 585
R289 B.n129 B.n128 585
R290 B.n127 B.n126 585
R291 B.n125 B.n124 585
R292 B.n123 B.n122 585
R293 B.n121 B.n120 585
R294 B.n119 B.n118 585
R295 B.n117 B.n116 585
R296 B.n115 B.n114 585
R297 B.n113 B.n112 585
R298 B.n111 B.n110 585
R299 B.n109 B.n108 585
R300 B.n107 B.n106 585
R301 B.n105 B.n104 585
R302 B.n103 B.n102 585
R303 B.n101 B.n100 585
R304 B.n99 B.n98 585
R305 B.n97 B.n96 585
R306 B.n95 B.n94 585
R307 B.n93 B.n92 585
R308 B.n504 B.n63 585
R309 B.n508 B.n63 585
R310 B.n503 B.n62 585
R311 B.n509 B.n62 585
R312 B.n502 B.n501 585
R313 B.n501 B.n58 585
R314 B.n500 B.n57 585
R315 B.n515 B.n57 585
R316 B.n499 B.n56 585
R317 B.n516 B.n56 585
R318 B.n498 B.n55 585
R319 B.n517 B.n55 585
R320 B.n497 B.n496 585
R321 B.n496 B.n54 585
R322 B.n495 B.n50 585
R323 B.n523 B.n50 585
R324 B.n494 B.n49 585
R325 B.n524 B.n49 585
R326 B.n493 B.n48 585
R327 B.n525 B.n48 585
R328 B.n492 B.n491 585
R329 B.n491 B.n44 585
R330 B.n490 B.n43 585
R331 B.n531 B.n43 585
R332 B.n489 B.n42 585
R333 B.n532 B.n42 585
R334 B.n488 B.n41 585
R335 B.n533 B.n41 585
R336 B.n487 B.n486 585
R337 B.n486 B.n37 585
R338 B.n485 B.n36 585
R339 B.n539 B.n36 585
R340 B.n484 B.n35 585
R341 B.n540 B.n35 585
R342 B.n483 B.n34 585
R343 B.n541 B.n34 585
R344 B.n482 B.n481 585
R345 B.n481 B.n30 585
R346 B.n480 B.n29 585
R347 B.n547 B.n29 585
R348 B.n479 B.n28 585
R349 B.n548 B.n28 585
R350 B.n478 B.n27 585
R351 B.n549 B.n27 585
R352 B.n477 B.n476 585
R353 B.n476 B.n26 585
R354 B.n475 B.n22 585
R355 B.n555 B.n22 585
R356 B.n474 B.n21 585
R357 B.n556 B.n21 585
R358 B.n473 B.n20 585
R359 B.n557 B.n20 585
R360 B.n472 B.n471 585
R361 B.n471 B.n16 585
R362 B.n470 B.n15 585
R363 B.n563 B.n15 585
R364 B.n469 B.n14 585
R365 B.n564 B.n14 585
R366 B.n468 B.n13 585
R367 B.n565 B.n13 585
R368 B.n467 B.n466 585
R369 B.n466 B.n12 585
R370 B.n465 B.n464 585
R371 B.n465 B.n8 585
R372 B.n463 B.n7 585
R373 B.n572 B.n7 585
R374 B.n462 B.n6 585
R375 B.n573 B.n6 585
R376 B.n461 B.n5 585
R377 B.n574 B.n5 585
R378 B.n460 B.n459 585
R379 B.n459 B.n4 585
R380 B.n458 B.n180 585
R381 B.n458 B.n457 585
R382 B.n448 B.n181 585
R383 B.n182 B.n181 585
R384 B.n450 B.n449 585
R385 B.n451 B.n450 585
R386 B.n447 B.n186 585
R387 B.n190 B.n186 585
R388 B.n446 B.n445 585
R389 B.n445 B.n444 585
R390 B.n188 B.n187 585
R391 B.n189 B.n188 585
R392 B.n437 B.n436 585
R393 B.n438 B.n437 585
R394 B.n435 B.n195 585
R395 B.n195 B.n194 585
R396 B.n434 B.n433 585
R397 B.n433 B.n432 585
R398 B.n197 B.n196 585
R399 B.n425 B.n197 585
R400 B.n424 B.n423 585
R401 B.n426 B.n424 585
R402 B.n422 B.n202 585
R403 B.n202 B.n201 585
R404 B.n421 B.n420 585
R405 B.n420 B.n419 585
R406 B.n204 B.n203 585
R407 B.n205 B.n204 585
R408 B.n412 B.n411 585
R409 B.n413 B.n412 585
R410 B.n410 B.n210 585
R411 B.n210 B.n209 585
R412 B.n409 B.n408 585
R413 B.n408 B.n407 585
R414 B.n212 B.n211 585
R415 B.n213 B.n212 585
R416 B.n400 B.n399 585
R417 B.n401 B.n400 585
R418 B.n398 B.n218 585
R419 B.n218 B.n217 585
R420 B.n397 B.n396 585
R421 B.n396 B.n395 585
R422 B.n220 B.n219 585
R423 B.n221 B.n220 585
R424 B.n388 B.n387 585
R425 B.n389 B.n388 585
R426 B.n386 B.n226 585
R427 B.n226 B.n225 585
R428 B.n385 B.n384 585
R429 B.n384 B.n383 585
R430 B.n228 B.n227 585
R431 B.n376 B.n228 585
R432 B.n375 B.n374 585
R433 B.n377 B.n375 585
R434 B.n373 B.n233 585
R435 B.n233 B.n232 585
R436 B.n372 B.n371 585
R437 B.n371 B.n370 585
R438 B.n235 B.n234 585
R439 B.n236 B.n235 585
R440 B.n363 B.n362 585
R441 B.n364 B.n363 585
R442 B.n361 B.n241 585
R443 B.n241 B.n240 585
R444 B.n355 B.n354 585
R445 B.n353 B.n265 585
R446 B.n352 B.n264 585
R447 B.n357 B.n264 585
R448 B.n351 B.n350 585
R449 B.n349 B.n348 585
R450 B.n347 B.n346 585
R451 B.n345 B.n344 585
R452 B.n343 B.n342 585
R453 B.n341 B.n340 585
R454 B.n339 B.n338 585
R455 B.n337 B.n336 585
R456 B.n335 B.n334 585
R457 B.n333 B.n332 585
R458 B.n331 B.n330 585
R459 B.n329 B.n328 585
R460 B.n327 B.n326 585
R461 B.n325 B.n324 585
R462 B.n323 B.n322 585
R463 B.n320 B.n319 585
R464 B.n318 B.n317 585
R465 B.n316 B.n315 585
R466 B.n314 B.n313 585
R467 B.n312 B.n311 585
R468 B.n310 B.n309 585
R469 B.n308 B.n307 585
R470 B.n306 B.n305 585
R471 B.n304 B.n303 585
R472 B.n302 B.n301 585
R473 B.n300 B.n299 585
R474 B.n298 B.n297 585
R475 B.n296 B.n295 585
R476 B.n294 B.n293 585
R477 B.n292 B.n291 585
R478 B.n290 B.n289 585
R479 B.n288 B.n287 585
R480 B.n286 B.n285 585
R481 B.n284 B.n283 585
R482 B.n282 B.n281 585
R483 B.n280 B.n279 585
R484 B.n278 B.n277 585
R485 B.n276 B.n275 585
R486 B.n274 B.n273 585
R487 B.n272 B.n271 585
R488 B.n243 B.n242 585
R489 B.n360 B.n359 585
R490 B.n239 B.n238 585
R491 B.n240 B.n239 585
R492 B.n366 B.n365 585
R493 B.n365 B.n364 585
R494 B.n367 B.n237 585
R495 B.n237 B.n236 585
R496 B.n369 B.n368 585
R497 B.n370 B.n369 585
R498 B.n231 B.n230 585
R499 B.n232 B.n231 585
R500 B.n379 B.n378 585
R501 B.n378 B.n377 585
R502 B.n380 B.n229 585
R503 B.n376 B.n229 585
R504 B.n382 B.n381 585
R505 B.n383 B.n382 585
R506 B.n224 B.n223 585
R507 B.n225 B.n224 585
R508 B.n391 B.n390 585
R509 B.n390 B.n389 585
R510 B.n392 B.n222 585
R511 B.n222 B.n221 585
R512 B.n394 B.n393 585
R513 B.n395 B.n394 585
R514 B.n216 B.n215 585
R515 B.n217 B.n216 585
R516 B.n403 B.n402 585
R517 B.n402 B.n401 585
R518 B.n404 B.n214 585
R519 B.n214 B.n213 585
R520 B.n406 B.n405 585
R521 B.n407 B.n406 585
R522 B.n208 B.n207 585
R523 B.n209 B.n208 585
R524 B.n415 B.n414 585
R525 B.n414 B.n413 585
R526 B.n416 B.n206 585
R527 B.n206 B.n205 585
R528 B.n418 B.n417 585
R529 B.n419 B.n418 585
R530 B.n200 B.n199 585
R531 B.n201 B.n200 585
R532 B.n428 B.n427 585
R533 B.n427 B.n426 585
R534 B.n429 B.n198 585
R535 B.n425 B.n198 585
R536 B.n431 B.n430 585
R537 B.n432 B.n431 585
R538 B.n193 B.n192 585
R539 B.n194 B.n193 585
R540 B.n440 B.n439 585
R541 B.n439 B.n438 585
R542 B.n441 B.n191 585
R543 B.n191 B.n189 585
R544 B.n443 B.n442 585
R545 B.n444 B.n443 585
R546 B.n185 B.n184 585
R547 B.n190 B.n185 585
R548 B.n453 B.n452 585
R549 B.n452 B.n451 585
R550 B.n454 B.n183 585
R551 B.n183 B.n182 585
R552 B.n456 B.n455 585
R553 B.n457 B.n456 585
R554 B.n3 B.n0 585
R555 B.n4 B.n3 585
R556 B.n571 B.n1 585
R557 B.n572 B.n571 585
R558 B.n570 B.n569 585
R559 B.n570 B.n8 585
R560 B.n568 B.n9 585
R561 B.n12 B.n9 585
R562 B.n567 B.n566 585
R563 B.n566 B.n565 585
R564 B.n11 B.n10 585
R565 B.n564 B.n11 585
R566 B.n562 B.n561 585
R567 B.n563 B.n562 585
R568 B.n560 B.n17 585
R569 B.n17 B.n16 585
R570 B.n559 B.n558 585
R571 B.n558 B.n557 585
R572 B.n19 B.n18 585
R573 B.n556 B.n19 585
R574 B.n554 B.n553 585
R575 B.n555 B.n554 585
R576 B.n552 B.n23 585
R577 B.n26 B.n23 585
R578 B.n551 B.n550 585
R579 B.n550 B.n549 585
R580 B.n25 B.n24 585
R581 B.n548 B.n25 585
R582 B.n546 B.n545 585
R583 B.n547 B.n546 585
R584 B.n544 B.n31 585
R585 B.n31 B.n30 585
R586 B.n543 B.n542 585
R587 B.n542 B.n541 585
R588 B.n33 B.n32 585
R589 B.n540 B.n33 585
R590 B.n538 B.n537 585
R591 B.n539 B.n538 585
R592 B.n536 B.n38 585
R593 B.n38 B.n37 585
R594 B.n535 B.n534 585
R595 B.n534 B.n533 585
R596 B.n40 B.n39 585
R597 B.n532 B.n40 585
R598 B.n530 B.n529 585
R599 B.n531 B.n530 585
R600 B.n528 B.n45 585
R601 B.n45 B.n44 585
R602 B.n527 B.n526 585
R603 B.n526 B.n525 585
R604 B.n47 B.n46 585
R605 B.n524 B.n47 585
R606 B.n522 B.n521 585
R607 B.n523 B.n522 585
R608 B.n520 B.n51 585
R609 B.n54 B.n51 585
R610 B.n519 B.n518 585
R611 B.n518 B.n517 585
R612 B.n53 B.n52 585
R613 B.n516 B.n53 585
R614 B.n514 B.n513 585
R615 B.n515 B.n514 585
R616 B.n512 B.n59 585
R617 B.n59 B.n58 585
R618 B.n511 B.n510 585
R619 B.n510 B.n509 585
R620 B.n61 B.n60 585
R621 B.n508 B.n61 585
R622 B.n575 B.n574 585
R623 B.n573 B.n2 585
R624 B.n92 B.n61 550.159
R625 B.n506 B.n63 550.159
R626 B.n359 B.n241 550.159
R627 B.n355 B.n239 550.159
R628 B.n87 B.t17 257.868
R629 B.n268 B.t6 257.868
R630 B.n89 B.t10 257.454
R631 B.n266 B.t14 257.454
R632 B.n507 B.n85 256.663
R633 B.n507 B.n84 256.663
R634 B.n507 B.n83 256.663
R635 B.n507 B.n82 256.663
R636 B.n507 B.n81 256.663
R637 B.n507 B.n80 256.663
R638 B.n507 B.n79 256.663
R639 B.n507 B.n78 256.663
R640 B.n507 B.n77 256.663
R641 B.n507 B.n76 256.663
R642 B.n507 B.n75 256.663
R643 B.n507 B.n74 256.663
R644 B.n507 B.n73 256.663
R645 B.n507 B.n72 256.663
R646 B.n507 B.n71 256.663
R647 B.n507 B.n70 256.663
R648 B.n507 B.n69 256.663
R649 B.n507 B.n68 256.663
R650 B.n507 B.n67 256.663
R651 B.n507 B.n66 256.663
R652 B.n507 B.n65 256.663
R653 B.n507 B.n64 256.663
R654 B.n357 B.n356 256.663
R655 B.n357 B.n244 256.663
R656 B.n357 B.n245 256.663
R657 B.n357 B.n246 256.663
R658 B.n357 B.n247 256.663
R659 B.n357 B.n248 256.663
R660 B.n357 B.n249 256.663
R661 B.n357 B.n250 256.663
R662 B.n357 B.n251 256.663
R663 B.n357 B.n252 256.663
R664 B.n357 B.n253 256.663
R665 B.n357 B.n254 256.663
R666 B.n357 B.n255 256.663
R667 B.n357 B.n256 256.663
R668 B.n357 B.n257 256.663
R669 B.n357 B.n258 256.663
R670 B.n357 B.n259 256.663
R671 B.n357 B.n260 256.663
R672 B.n357 B.n261 256.663
R673 B.n357 B.n262 256.663
R674 B.n357 B.n263 256.663
R675 B.n358 B.n357 256.663
R676 B.n577 B.n576 256.663
R677 B.n87 B.t18 185.6
R678 B.n268 B.t9 185.6
R679 B.n89 B.t12 185.6
R680 B.n266 B.t16 185.6
R681 B.n357 B.n240 169.232
R682 B.n508 B.n507 169.232
R683 B.n96 B.n95 163.367
R684 B.n100 B.n99 163.367
R685 B.n104 B.n103 163.367
R686 B.n108 B.n107 163.367
R687 B.n112 B.n111 163.367
R688 B.n116 B.n115 163.367
R689 B.n120 B.n119 163.367
R690 B.n124 B.n123 163.367
R691 B.n128 B.n127 163.367
R692 B.n132 B.n131 163.367
R693 B.n136 B.n135 163.367
R694 B.n140 B.n139 163.367
R695 B.n144 B.n143 163.367
R696 B.n149 B.n148 163.367
R697 B.n153 B.n152 163.367
R698 B.n157 B.n156 163.367
R699 B.n161 B.n160 163.367
R700 B.n165 B.n164 163.367
R701 B.n169 B.n168 163.367
R702 B.n173 B.n172 163.367
R703 B.n177 B.n176 163.367
R704 B.n506 B.n86 163.367
R705 B.n363 B.n241 163.367
R706 B.n363 B.n235 163.367
R707 B.n371 B.n235 163.367
R708 B.n371 B.n233 163.367
R709 B.n375 B.n233 163.367
R710 B.n375 B.n228 163.367
R711 B.n384 B.n228 163.367
R712 B.n384 B.n226 163.367
R713 B.n388 B.n226 163.367
R714 B.n388 B.n220 163.367
R715 B.n396 B.n220 163.367
R716 B.n396 B.n218 163.367
R717 B.n400 B.n218 163.367
R718 B.n400 B.n212 163.367
R719 B.n408 B.n212 163.367
R720 B.n408 B.n210 163.367
R721 B.n412 B.n210 163.367
R722 B.n412 B.n204 163.367
R723 B.n420 B.n204 163.367
R724 B.n420 B.n202 163.367
R725 B.n424 B.n202 163.367
R726 B.n424 B.n197 163.367
R727 B.n433 B.n197 163.367
R728 B.n433 B.n195 163.367
R729 B.n437 B.n195 163.367
R730 B.n437 B.n188 163.367
R731 B.n445 B.n188 163.367
R732 B.n445 B.n186 163.367
R733 B.n450 B.n186 163.367
R734 B.n450 B.n181 163.367
R735 B.n458 B.n181 163.367
R736 B.n459 B.n458 163.367
R737 B.n459 B.n5 163.367
R738 B.n6 B.n5 163.367
R739 B.n7 B.n6 163.367
R740 B.n465 B.n7 163.367
R741 B.n466 B.n465 163.367
R742 B.n466 B.n13 163.367
R743 B.n14 B.n13 163.367
R744 B.n15 B.n14 163.367
R745 B.n471 B.n15 163.367
R746 B.n471 B.n20 163.367
R747 B.n21 B.n20 163.367
R748 B.n22 B.n21 163.367
R749 B.n476 B.n22 163.367
R750 B.n476 B.n27 163.367
R751 B.n28 B.n27 163.367
R752 B.n29 B.n28 163.367
R753 B.n481 B.n29 163.367
R754 B.n481 B.n34 163.367
R755 B.n35 B.n34 163.367
R756 B.n36 B.n35 163.367
R757 B.n486 B.n36 163.367
R758 B.n486 B.n41 163.367
R759 B.n42 B.n41 163.367
R760 B.n43 B.n42 163.367
R761 B.n491 B.n43 163.367
R762 B.n491 B.n48 163.367
R763 B.n49 B.n48 163.367
R764 B.n50 B.n49 163.367
R765 B.n496 B.n50 163.367
R766 B.n496 B.n55 163.367
R767 B.n56 B.n55 163.367
R768 B.n57 B.n56 163.367
R769 B.n501 B.n57 163.367
R770 B.n501 B.n62 163.367
R771 B.n63 B.n62 163.367
R772 B.n265 B.n264 163.367
R773 B.n350 B.n264 163.367
R774 B.n348 B.n347 163.367
R775 B.n344 B.n343 163.367
R776 B.n340 B.n339 163.367
R777 B.n336 B.n335 163.367
R778 B.n332 B.n331 163.367
R779 B.n328 B.n327 163.367
R780 B.n324 B.n323 163.367
R781 B.n319 B.n318 163.367
R782 B.n315 B.n314 163.367
R783 B.n311 B.n310 163.367
R784 B.n307 B.n306 163.367
R785 B.n303 B.n302 163.367
R786 B.n299 B.n298 163.367
R787 B.n295 B.n294 163.367
R788 B.n291 B.n290 163.367
R789 B.n287 B.n286 163.367
R790 B.n283 B.n282 163.367
R791 B.n279 B.n278 163.367
R792 B.n275 B.n274 163.367
R793 B.n271 B.n243 163.367
R794 B.n365 B.n239 163.367
R795 B.n365 B.n237 163.367
R796 B.n369 B.n237 163.367
R797 B.n369 B.n231 163.367
R798 B.n378 B.n231 163.367
R799 B.n378 B.n229 163.367
R800 B.n382 B.n229 163.367
R801 B.n382 B.n224 163.367
R802 B.n390 B.n224 163.367
R803 B.n390 B.n222 163.367
R804 B.n394 B.n222 163.367
R805 B.n394 B.n216 163.367
R806 B.n402 B.n216 163.367
R807 B.n402 B.n214 163.367
R808 B.n406 B.n214 163.367
R809 B.n406 B.n208 163.367
R810 B.n414 B.n208 163.367
R811 B.n414 B.n206 163.367
R812 B.n418 B.n206 163.367
R813 B.n418 B.n200 163.367
R814 B.n427 B.n200 163.367
R815 B.n427 B.n198 163.367
R816 B.n431 B.n198 163.367
R817 B.n431 B.n193 163.367
R818 B.n439 B.n193 163.367
R819 B.n439 B.n191 163.367
R820 B.n443 B.n191 163.367
R821 B.n443 B.n185 163.367
R822 B.n452 B.n185 163.367
R823 B.n452 B.n183 163.367
R824 B.n456 B.n183 163.367
R825 B.n456 B.n3 163.367
R826 B.n575 B.n3 163.367
R827 B.n571 B.n2 163.367
R828 B.n571 B.n570 163.367
R829 B.n570 B.n9 163.367
R830 B.n566 B.n9 163.367
R831 B.n566 B.n11 163.367
R832 B.n562 B.n11 163.367
R833 B.n562 B.n17 163.367
R834 B.n558 B.n17 163.367
R835 B.n558 B.n19 163.367
R836 B.n554 B.n19 163.367
R837 B.n554 B.n23 163.367
R838 B.n550 B.n23 163.367
R839 B.n550 B.n25 163.367
R840 B.n546 B.n25 163.367
R841 B.n546 B.n31 163.367
R842 B.n542 B.n31 163.367
R843 B.n542 B.n33 163.367
R844 B.n538 B.n33 163.367
R845 B.n538 B.n38 163.367
R846 B.n534 B.n38 163.367
R847 B.n534 B.n40 163.367
R848 B.n530 B.n40 163.367
R849 B.n530 B.n45 163.367
R850 B.n526 B.n45 163.367
R851 B.n526 B.n47 163.367
R852 B.n522 B.n47 163.367
R853 B.n522 B.n51 163.367
R854 B.n518 B.n51 163.367
R855 B.n518 B.n53 163.367
R856 B.n514 B.n53 163.367
R857 B.n514 B.n59 163.367
R858 B.n510 B.n59 163.367
R859 B.n510 B.n61 163.367
R860 B.n88 B.t19 143.321
R861 B.n269 B.t8 143.321
R862 B.n90 B.t13 143.321
R863 B.n267 B.t15 143.321
R864 B.n364 B.n240 81.6153
R865 B.n364 B.n236 81.6153
R866 B.n370 B.n236 81.6153
R867 B.n370 B.n232 81.6153
R868 B.n377 B.n232 81.6153
R869 B.n377 B.n376 81.6153
R870 B.n383 B.n225 81.6153
R871 B.n389 B.n225 81.6153
R872 B.n389 B.n221 81.6153
R873 B.n395 B.n221 81.6153
R874 B.n395 B.n217 81.6153
R875 B.n401 B.n217 81.6153
R876 B.n401 B.n213 81.6153
R877 B.n407 B.n213 81.6153
R878 B.n413 B.n209 81.6153
R879 B.n413 B.n205 81.6153
R880 B.n419 B.n205 81.6153
R881 B.n419 B.n201 81.6153
R882 B.n426 B.n201 81.6153
R883 B.n426 B.n425 81.6153
R884 B.n432 B.n194 81.6153
R885 B.n438 B.n194 81.6153
R886 B.n438 B.n189 81.6153
R887 B.n444 B.n189 81.6153
R888 B.n444 B.n190 81.6153
R889 B.n451 B.n182 81.6153
R890 B.n457 B.n182 81.6153
R891 B.n457 B.n4 81.6153
R892 B.n574 B.n4 81.6153
R893 B.n574 B.n573 81.6153
R894 B.n573 B.n572 81.6153
R895 B.n572 B.n8 81.6153
R896 B.n12 B.n8 81.6153
R897 B.n565 B.n12 81.6153
R898 B.n564 B.n563 81.6153
R899 B.n563 B.n16 81.6153
R900 B.n557 B.n16 81.6153
R901 B.n557 B.n556 81.6153
R902 B.n556 B.n555 81.6153
R903 B.n549 B.n26 81.6153
R904 B.n549 B.n548 81.6153
R905 B.n548 B.n547 81.6153
R906 B.n547 B.n30 81.6153
R907 B.n541 B.n30 81.6153
R908 B.n541 B.n540 81.6153
R909 B.n539 B.n37 81.6153
R910 B.n533 B.n37 81.6153
R911 B.n533 B.n532 81.6153
R912 B.n532 B.n531 81.6153
R913 B.n531 B.n44 81.6153
R914 B.n525 B.n44 81.6153
R915 B.n525 B.n524 81.6153
R916 B.n524 B.n523 81.6153
R917 B.n517 B.n54 81.6153
R918 B.n517 B.n516 81.6153
R919 B.n516 B.n515 81.6153
R920 B.n515 B.n58 81.6153
R921 B.n509 B.n58 81.6153
R922 B.n509 B.n508 81.6153
R923 B.n92 B.n64 71.676
R924 B.n96 B.n65 71.676
R925 B.n100 B.n66 71.676
R926 B.n104 B.n67 71.676
R927 B.n108 B.n68 71.676
R928 B.n112 B.n69 71.676
R929 B.n116 B.n70 71.676
R930 B.n120 B.n71 71.676
R931 B.n124 B.n72 71.676
R932 B.n128 B.n73 71.676
R933 B.n132 B.n74 71.676
R934 B.n136 B.n75 71.676
R935 B.n140 B.n76 71.676
R936 B.n144 B.n77 71.676
R937 B.n149 B.n78 71.676
R938 B.n153 B.n79 71.676
R939 B.n157 B.n80 71.676
R940 B.n161 B.n81 71.676
R941 B.n165 B.n82 71.676
R942 B.n169 B.n83 71.676
R943 B.n173 B.n84 71.676
R944 B.n177 B.n85 71.676
R945 B.n86 B.n85 71.676
R946 B.n176 B.n84 71.676
R947 B.n172 B.n83 71.676
R948 B.n168 B.n82 71.676
R949 B.n164 B.n81 71.676
R950 B.n160 B.n80 71.676
R951 B.n156 B.n79 71.676
R952 B.n152 B.n78 71.676
R953 B.n148 B.n77 71.676
R954 B.n143 B.n76 71.676
R955 B.n139 B.n75 71.676
R956 B.n135 B.n74 71.676
R957 B.n131 B.n73 71.676
R958 B.n127 B.n72 71.676
R959 B.n123 B.n71 71.676
R960 B.n119 B.n70 71.676
R961 B.n115 B.n69 71.676
R962 B.n111 B.n68 71.676
R963 B.n107 B.n67 71.676
R964 B.n103 B.n66 71.676
R965 B.n99 B.n65 71.676
R966 B.n95 B.n64 71.676
R967 B.n356 B.n355 71.676
R968 B.n350 B.n244 71.676
R969 B.n347 B.n245 71.676
R970 B.n343 B.n246 71.676
R971 B.n339 B.n247 71.676
R972 B.n335 B.n248 71.676
R973 B.n331 B.n249 71.676
R974 B.n327 B.n250 71.676
R975 B.n323 B.n251 71.676
R976 B.n318 B.n252 71.676
R977 B.n314 B.n253 71.676
R978 B.n310 B.n254 71.676
R979 B.n306 B.n255 71.676
R980 B.n302 B.n256 71.676
R981 B.n298 B.n257 71.676
R982 B.n294 B.n258 71.676
R983 B.n290 B.n259 71.676
R984 B.n286 B.n260 71.676
R985 B.n282 B.n261 71.676
R986 B.n278 B.n262 71.676
R987 B.n274 B.n263 71.676
R988 B.n358 B.n243 71.676
R989 B.n356 B.n265 71.676
R990 B.n348 B.n244 71.676
R991 B.n344 B.n245 71.676
R992 B.n340 B.n246 71.676
R993 B.n336 B.n247 71.676
R994 B.n332 B.n248 71.676
R995 B.n328 B.n249 71.676
R996 B.n324 B.n250 71.676
R997 B.n319 B.n251 71.676
R998 B.n315 B.n252 71.676
R999 B.n311 B.n253 71.676
R1000 B.n307 B.n254 71.676
R1001 B.n303 B.n255 71.676
R1002 B.n299 B.n256 71.676
R1003 B.n295 B.n257 71.676
R1004 B.n291 B.n258 71.676
R1005 B.n287 B.n259 71.676
R1006 B.n283 B.n260 71.676
R1007 B.n279 B.n261 71.676
R1008 B.n275 B.n262 71.676
R1009 B.n271 B.n263 71.676
R1010 B.n359 B.n358 71.676
R1011 B.n576 B.n575 71.676
R1012 B.n576 B.n2 71.676
R1013 B.n407 B.t3 70.8134
R1014 B.t5 B.n539 70.8134
R1015 B.n383 B.t7 61.2116
R1016 B.n523 B.t11 61.2116
R1017 B.n91 B.n90 59.5399
R1018 B.n146 B.n88 59.5399
R1019 B.n270 B.n269 59.5399
R1020 B.n321 B.n267 59.5399
R1021 B.n432 B.t2 58.8112
R1022 B.n555 B.t1 58.8112
R1023 B.n190 B.t4 56.4108
R1024 B.t0 B.n564 56.4108
R1025 B.n90 B.n89 42.2793
R1026 B.n88 B.n87 42.2793
R1027 B.n269 B.n268 42.2793
R1028 B.n267 B.n266 42.2793
R1029 B.n505 B.n504 35.7468
R1030 B.n354 B.n238 35.7468
R1031 B.n361 B.n360 35.7468
R1032 B.n93 B.n60 35.7468
R1033 B.n451 B.t4 25.2051
R1034 B.n565 B.t0 25.2051
R1035 B.n425 B.t2 22.8046
R1036 B.n26 B.t1 22.8046
R1037 B.n376 B.t7 20.4042
R1038 B.n54 B.t11 20.4042
R1039 B B.n577 18.0485
R1040 B.t3 B.n209 10.8025
R1041 B.n540 B.t5 10.8025
R1042 B.n366 B.n238 10.6151
R1043 B.n367 B.n366 10.6151
R1044 B.n368 B.n367 10.6151
R1045 B.n368 B.n230 10.6151
R1046 B.n379 B.n230 10.6151
R1047 B.n380 B.n379 10.6151
R1048 B.n381 B.n380 10.6151
R1049 B.n381 B.n223 10.6151
R1050 B.n391 B.n223 10.6151
R1051 B.n392 B.n391 10.6151
R1052 B.n393 B.n392 10.6151
R1053 B.n393 B.n215 10.6151
R1054 B.n403 B.n215 10.6151
R1055 B.n404 B.n403 10.6151
R1056 B.n405 B.n404 10.6151
R1057 B.n405 B.n207 10.6151
R1058 B.n415 B.n207 10.6151
R1059 B.n416 B.n415 10.6151
R1060 B.n417 B.n416 10.6151
R1061 B.n417 B.n199 10.6151
R1062 B.n428 B.n199 10.6151
R1063 B.n429 B.n428 10.6151
R1064 B.n430 B.n429 10.6151
R1065 B.n430 B.n192 10.6151
R1066 B.n440 B.n192 10.6151
R1067 B.n441 B.n440 10.6151
R1068 B.n442 B.n441 10.6151
R1069 B.n442 B.n184 10.6151
R1070 B.n453 B.n184 10.6151
R1071 B.n454 B.n453 10.6151
R1072 B.n455 B.n454 10.6151
R1073 B.n455 B.n0 10.6151
R1074 B.n354 B.n353 10.6151
R1075 B.n353 B.n352 10.6151
R1076 B.n352 B.n351 10.6151
R1077 B.n351 B.n349 10.6151
R1078 B.n349 B.n346 10.6151
R1079 B.n346 B.n345 10.6151
R1080 B.n345 B.n342 10.6151
R1081 B.n342 B.n341 10.6151
R1082 B.n341 B.n338 10.6151
R1083 B.n338 B.n337 10.6151
R1084 B.n337 B.n334 10.6151
R1085 B.n334 B.n333 10.6151
R1086 B.n333 B.n330 10.6151
R1087 B.n330 B.n329 10.6151
R1088 B.n329 B.n326 10.6151
R1089 B.n326 B.n325 10.6151
R1090 B.n325 B.n322 10.6151
R1091 B.n320 B.n317 10.6151
R1092 B.n317 B.n316 10.6151
R1093 B.n316 B.n313 10.6151
R1094 B.n313 B.n312 10.6151
R1095 B.n312 B.n309 10.6151
R1096 B.n309 B.n308 10.6151
R1097 B.n308 B.n305 10.6151
R1098 B.n305 B.n304 10.6151
R1099 B.n301 B.n300 10.6151
R1100 B.n300 B.n297 10.6151
R1101 B.n297 B.n296 10.6151
R1102 B.n296 B.n293 10.6151
R1103 B.n293 B.n292 10.6151
R1104 B.n292 B.n289 10.6151
R1105 B.n289 B.n288 10.6151
R1106 B.n288 B.n285 10.6151
R1107 B.n285 B.n284 10.6151
R1108 B.n284 B.n281 10.6151
R1109 B.n281 B.n280 10.6151
R1110 B.n280 B.n277 10.6151
R1111 B.n277 B.n276 10.6151
R1112 B.n276 B.n273 10.6151
R1113 B.n273 B.n272 10.6151
R1114 B.n272 B.n242 10.6151
R1115 B.n360 B.n242 10.6151
R1116 B.n362 B.n361 10.6151
R1117 B.n362 B.n234 10.6151
R1118 B.n372 B.n234 10.6151
R1119 B.n373 B.n372 10.6151
R1120 B.n374 B.n373 10.6151
R1121 B.n374 B.n227 10.6151
R1122 B.n385 B.n227 10.6151
R1123 B.n386 B.n385 10.6151
R1124 B.n387 B.n386 10.6151
R1125 B.n387 B.n219 10.6151
R1126 B.n397 B.n219 10.6151
R1127 B.n398 B.n397 10.6151
R1128 B.n399 B.n398 10.6151
R1129 B.n399 B.n211 10.6151
R1130 B.n409 B.n211 10.6151
R1131 B.n410 B.n409 10.6151
R1132 B.n411 B.n410 10.6151
R1133 B.n411 B.n203 10.6151
R1134 B.n421 B.n203 10.6151
R1135 B.n422 B.n421 10.6151
R1136 B.n423 B.n422 10.6151
R1137 B.n423 B.n196 10.6151
R1138 B.n434 B.n196 10.6151
R1139 B.n435 B.n434 10.6151
R1140 B.n436 B.n435 10.6151
R1141 B.n436 B.n187 10.6151
R1142 B.n446 B.n187 10.6151
R1143 B.n447 B.n446 10.6151
R1144 B.n449 B.n447 10.6151
R1145 B.n449 B.n448 10.6151
R1146 B.n448 B.n180 10.6151
R1147 B.n460 B.n180 10.6151
R1148 B.n461 B.n460 10.6151
R1149 B.n462 B.n461 10.6151
R1150 B.n463 B.n462 10.6151
R1151 B.n464 B.n463 10.6151
R1152 B.n467 B.n464 10.6151
R1153 B.n468 B.n467 10.6151
R1154 B.n469 B.n468 10.6151
R1155 B.n470 B.n469 10.6151
R1156 B.n472 B.n470 10.6151
R1157 B.n473 B.n472 10.6151
R1158 B.n474 B.n473 10.6151
R1159 B.n475 B.n474 10.6151
R1160 B.n477 B.n475 10.6151
R1161 B.n478 B.n477 10.6151
R1162 B.n479 B.n478 10.6151
R1163 B.n480 B.n479 10.6151
R1164 B.n482 B.n480 10.6151
R1165 B.n483 B.n482 10.6151
R1166 B.n484 B.n483 10.6151
R1167 B.n485 B.n484 10.6151
R1168 B.n487 B.n485 10.6151
R1169 B.n488 B.n487 10.6151
R1170 B.n489 B.n488 10.6151
R1171 B.n490 B.n489 10.6151
R1172 B.n492 B.n490 10.6151
R1173 B.n493 B.n492 10.6151
R1174 B.n494 B.n493 10.6151
R1175 B.n495 B.n494 10.6151
R1176 B.n497 B.n495 10.6151
R1177 B.n498 B.n497 10.6151
R1178 B.n499 B.n498 10.6151
R1179 B.n500 B.n499 10.6151
R1180 B.n502 B.n500 10.6151
R1181 B.n503 B.n502 10.6151
R1182 B.n504 B.n503 10.6151
R1183 B.n569 B.n1 10.6151
R1184 B.n569 B.n568 10.6151
R1185 B.n568 B.n567 10.6151
R1186 B.n567 B.n10 10.6151
R1187 B.n561 B.n10 10.6151
R1188 B.n561 B.n560 10.6151
R1189 B.n560 B.n559 10.6151
R1190 B.n559 B.n18 10.6151
R1191 B.n553 B.n18 10.6151
R1192 B.n553 B.n552 10.6151
R1193 B.n552 B.n551 10.6151
R1194 B.n551 B.n24 10.6151
R1195 B.n545 B.n24 10.6151
R1196 B.n545 B.n544 10.6151
R1197 B.n544 B.n543 10.6151
R1198 B.n543 B.n32 10.6151
R1199 B.n537 B.n32 10.6151
R1200 B.n537 B.n536 10.6151
R1201 B.n536 B.n535 10.6151
R1202 B.n535 B.n39 10.6151
R1203 B.n529 B.n39 10.6151
R1204 B.n529 B.n528 10.6151
R1205 B.n528 B.n527 10.6151
R1206 B.n527 B.n46 10.6151
R1207 B.n521 B.n46 10.6151
R1208 B.n521 B.n520 10.6151
R1209 B.n520 B.n519 10.6151
R1210 B.n519 B.n52 10.6151
R1211 B.n513 B.n52 10.6151
R1212 B.n513 B.n512 10.6151
R1213 B.n512 B.n511 10.6151
R1214 B.n511 B.n60 10.6151
R1215 B.n94 B.n93 10.6151
R1216 B.n97 B.n94 10.6151
R1217 B.n98 B.n97 10.6151
R1218 B.n101 B.n98 10.6151
R1219 B.n102 B.n101 10.6151
R1220 B.n105 B.n102 10.6151
R1221 B.n106 B.n105 10.6151
R1222 B.n109 B.n106 10.6151
R1223 B.n110 B.n109 10.6151
R1224 B.n113 B.n110 10.6151
R1225 B.n114 B.n113 10.6151
R1226 B.n117 B.n114 10.6151
R1227 B.n118 B.n117 10.6151
R1228 B.n121 B.n118 10.6151
R1229 B.n122 B.n121 10.6151
R1230 B.n125 B.n122 10.6151
R1231 B.n126 B.n125 10.6151
R1232 B.n130 B.n129 10.6151
R1233 B.n133 B.n130 10.6151
R1234 B.n134 B.n133 10.6151
R1235 B.n137 B.n134 10.6151
R1236 B.n138 B.n137 10.6151
R1237 B.n141 B.n138 10.6151
R1238 B.n142 B.n141 10.6151
R1239 B.n145 B.n142 10.6151
R1240 B.n150 B.n147 10.6151
R1241 B.n151 B.n150 10.6151
R1242 B.n154 B.n151 10.6151
R1243 B.n155 B.n154 10.6151
R1244 B.n158 B.n155 10.6151
R1245 B.n159 B.n158 10.6151
R1246 B.n162 B.n159 10.6151
R1247 B.n163 B.n162 10.6151
R1248 B.n166 B.n163 10.6151
R1249 B.n167 B.n166 10.6151
R1250 B.n170 B.n167 10.6151
R1251 B.n171 B.n170 10.6151
R1252 B.n174 B.n171 10.6151
R1253 B.n175 B.n174 10.6151
R1254 B.n178 B.n175 10.6151
R1255 B.n179 B.n178 10.6151
R1256 B.n505 B.n179 10.6151
R1257 B.n577 B.n0 8.11757
R1258 B.n577 B.n1 8.11757
R1259 B.n321 B.n320 6.4005
R1260 B.n304 B.n270 6.4005
R1261 B.n129 B.n91 6.4005
R1262 B.n146 B.n145 6.4005
R1263 B.n322 B.n321 4.21513
R1264 B.n301 B.n270 4.21513
R1265 B.n126 B.n91 4.21513
R1266 B.n147 B.n146 4.21513
R1267 VN.n21 VN.n12 161.3
R1268 VN.n20 VN.n19 161.3
R1269 VN.n18 VN.n13 161.3
R1270 VN.n17 VN.n16 161.3
R1271 VN.n9 VN.n0 161.3
R1272 VN.n8 VN.n7 161.3
R1273 VN.n6 VN.n1 161.3
R1274 VN.n5 VN.n4 161.3
R1275 VN.n11 VN.n10 89.7148
R1276 VN.n23 VN.n22 89.7148
R1277 VN.n2 VN.t2 81.2706
R1278 VN.n14 VN.t4 81.2706
R1279 VN.n3 VN.n2 57.6865
R1280 VN.n15 VN.n14 57.6865
R1281 VN.n8 VN.n1 56.0336
R1282 VN.n20 VN.n13 56.0336
R1283 VN.n3 VN.t3 50.6756
R1284 VN.n10 VN.t1 50.6756
R1285 VN.n15 VN.t5 50.6756
R1286 VN.n22 VN.t0 50.6756
R1287 VN VN.n23 39.8769
R1288 VN.n9 VN.n8 24.9531
R1289 VN.n21 VN.n20 24.9531
R1290 VN.n4 VN.n1 24.4675
R1291 VN.n16 VN.n13 24.4675
R1292 VN.n10 VN.n9 21.0421
R1293 VN.n22 VN.n21 21.0421
R1294 VN.n17 VN.n14 13.151
R1295 VN.n5 VN.n2 13.151
R1296 VN.n4 VN.n3 12.234
R1297 VN.n16 VN.n15 12.234
R1298 VN.n23 VN.n12 0.278367
R1299 VN.n11 VN.n0 0.278367
R1300 VN.n19 VN.n12 0.189894
R1301 VN.n19 VN.n18 0.189894
R1302 VN.n18 VN.n17 0.189894
R1303 VN.n6 VN.n5 0.189894
R1304 VN.n7 VN.n6 0.189894
R1305 VN.n7 VN.n0 0.189894
R1306 VN VN.n11 0.153454
R1307 VDD2.n35 VDD2.n21 289.615
R1308 VDD2.n14 VDD2.n0 289.615
R1309 VDD2.n36 VDD2.n35 185
R1310 VDD2.n34 VDD2.n33 185
R1311 VDD2.n25 VDD2.n24 185
R1312 VDD2.n28 VDD2.n27 185
R1313 VDD2.n7 VDD2.n6 185
R1314 VDD2.n4 VDD2.n3 185
R1315 VDD2.n13 VDD2.n12 185
R1316 VDD2.n15 VDD2.n14 185
R1317 VDD2.t5 VDD2.n26 147.888
R1318 VDD2.t3 VDD2.n5 147.888
R1319 VDD2.n35 VDD2.n34 104.615
R1320 VDD2.n34 VDD2.n24 104.615
R1321 VDD2.n27 VDD2.n24 104.615
R1322 VDD2.n6 VDD2.n3 104.615
R1323 VDD2.n13 VDD2.n3 104.615
R1324 VDD2.n14 VDD2.n13 104.615
R1325 VDD2.n20 VDD2.n19 74.8481
R1326 VDD2 VDD2.n41 74.8453
R1327 VDD2.n27 VDD2.t5 52.3082
R1328 VDD2.n6 VDD2.t3 52.3082
R1329 VDD2.n20 VDD2.n18 51.188
R1330 VDD2.n40 VDD2.n39 49.8338
R1331 VDD2.n40 VDD2.n20 33.1765
R1332 VDD2.n28 VDD2.n26 15.6496
R1333 VDD2.n7 VDD2.n5 15.6496
R1334 VDD2.n29 VDD2.n25 12.8005
R1335 VDD2.n8 VDD2.n4 12.8005
R1336 VDD2.n33 VDD2.n32 12.0247
R1337 VDD2.n12 VDD2.n11 12.0247
R1338 VDD2.n36 VDD2.n23 11.249
R1339 VDD2.n15 VDD2.n2 11.249
R1340 VDD2.n37 VDD2.n21 10.4732
R1341 VDD2.n16 VDD2.n0 10.4732
R1342 VDD2.n39 VDD2.n38 9.45567
R1343 VDD2.n18 VDD2.n17 9.45567
R1344 VDD2.n38 VDD2.n37 9.3005
R1345 VDD2.n23 VDD2.n22 9.3005
R1346 VDD2.n32 VDD2.n31 9.3005
R1347 VDD2.n30 VDD2.n29 9.3005
R1348 VDD2.n17 VDD2.n16 9.3005
R1349 VDD2.n2 VDD2.n1 9.3005
R1350 VDD2.n11 VDD2.n10 9.3005
R1351 VDD2.n9 VDD2.n8 9.3005
R1352 VDD2.n41 VDD2.t0 5.09047
R1353 VDD2.n41 VDD2.t1 5.09047
R1354 VDD2.n19 VDD2.t2 5.09047
R1355 VDD2.n19 VDD2.t4 5.09047
R1356 VDD2.n30 VDD2.n26 4.40546
R1357 VDD2.n9 VDD2.n5 4.40546
R1358 VDD2.n39 VDD2.n21 3.49141
R1359 VDD2.n18 VDD2.n0 3.49141
R1360 VDD2.n37 VDD2.n36 2.71565
R1361 VDD2.n16 VDD2.n15 2.71565
R1362 VDD2.n33 VDD2.n23 1.93989
R1363 VDD2.n12 VDD2.n2 1.93989
R1364 VDD2 VDD2.n40 1.46817
R1365 VDD2.n32 VDD2.n25 1.16414
R1366 VDD2.n11 VDD2.n4 1.16414
R1367 VDD2.n29 VDD2.n28 0.388379
R1368 VDD2.n8 VDD2.n7 0.388379
R1369 VDD2.n38 VDD2.n22 0.155672
R1370 VDD2.n31 VDD2.n22 0.155672
R1371 VDD2.n31 VDD2.n30 0.155672
R1372 VDD2.n10 VDD2.n9 0.155672
R1373 VDD2.n10 VDD2.n1 0.155672
R1374 VDD2.n17 VDD2.n1 0.155672
C0 VDD2 VTAIL 4.44355f
C1 VN VP 4.70509f
C2 VDD1 VTAIL 4.39621f
C3 VDD2 VP 0.398886f
C4 VDD1 VP 2.51473f
C5 VTAIL VP 2.74917f
C6 VDD2 VN 2.27223f
C7 VDD1 VN 0.154133f
C8 VTAIL VN 2.73498f
C9 VDD2 VDD1 1.1388f
C10 VDD2 B 3.925388f
C11 VDD1 B 4.021509f
C12 VTAIL B 3.859866f
C13 VN B 9.95096f
C14 VP B 8.551014f
C15 VDD2.n0 B 0.030093f
C16 VDD2.n1 B 0.022154f
C17 VDD2.n2 B 0.011905f
C18 VDD2.n3 B 0.028139f
C19 VDD2.n4 B 0.012605f
C20 VDD2.n5 B 0.084587f
C21 VDD2.t3 B 0.046582f
C22 VDD2.n6 B 0.021104f
C23 VDD2.n7 B 0.016561f
C24 VDD2.n8 B 0.011905f
C25 VDD2.n9 B 0.310581f
C26 VDD2.n10 B 0.022154f
C27 VDD2.n11 B 0.011905f
C28 VDD2.n12 B 0.012605f
C29 VDD2.n13 B 0.028139f
C30 VDD2.n14 B 0.059065f
C31 VDD2.n15 B 0.012605f
C32 VDD2.n16 B 0.011905f
C33 VDD2.n17 B 0.052722f
C34 VDD2.n18 B 0.051909f
C35 VDD2.t2 B 0.068102f
C36 VDD2.t4 B 0.068102f
C37 VDD2.n19 B 0.53469f
C38 VDD2.n20 B 1.64753f
C39 VDD2.n21 B 0.030093f
C40 VDD2.n22 B 0.022154f
C41 VDD2.n23 B 0.011905f
C42 VDD2.n24 B 0.028139f
C43 VDD2.n25 B 0.012605f
C44 VDD2.n26 B 0.084587f
C45 VDD2.t5 B 0.046582f
C46 VDD2.n27 B 0.021104f
C47 VDD2.n28 B 0.016561f
C48 VDD2.n29 B 0.011905f
C49 VDD2.n30 B 0.310581f
C50 VDD2.n31 B 0.022154f
C51 VDD2.n32 B 0.011905f
C52 VDD2.n33 B 0.012605f
C53 VDD2.n34 B 0.028139f
C54 VDD2.n35 B 0.059065f
C55 VDD2.n36 B 0.012605f
C56 VDD2.n37 B 0.011905f
C57 VDD2.n38 B 0.052722f
C58 VDD2.n39 B 0.04819f
C59 VDD2.n40 B 1.51965f
C60 VDD2.t0 B 0.068102f
C61 VDD2.t1 B 0.068102f
C62 VDD2.n41 B 0.534669f
C63 VN.n0 B 0.043736f
C64 VN.t1 B 0.610561f
C65 VN.n1 B 0.056665f
C66 VN.t2 B 0.763906f
C67 VN.n2 B 0.328832f
C68 VN.t3 B 0.610561f
C69 VN.n3 B 0.328675f
C70 VN.n4 B 0.046565f
C71 VN.n5 B 0.243925f
C72 VN.n6 B 0.033173f
C73 VN.n7 B 0.033173f
C74 VN.n8 B 0.039608f
C75 VN.n9 B 0.058134f
C76 VN.n10 B 0.350095f
C77 VN.n11 B 0.038326f
C78 VN.n12 B 0.043736f
C79 VN.t0 B 0.610561f
C80 VN.n13 B 0.056665f
C81 VN.t4 B 0.763906f
C82 VN.n14 B 0.328832f
C83 VN.t5 B 0.610561f
C84 VN.n15 B 0.328675f
C85 VN.n16 B 0.046565f
C86 VN.n17 B 0.243925f
C87 VN.n18 B 0.033173f
C88 VN.n19 B 0.033173f
C89 VN.n20 B 0.039608f
C90 VN.n21 B 0.058134f
C91 VN.n22 B 0.350095f
C92 VN.n23 B 1.28259f
C93 VDD1.n0 B 0.030618f
C94 VDD1.n1 B 0.02254f
C95 VDD1.n2 B 0.012112f
C96 VDD1.n3 B 0.028629f
C97 VDD1.n4 B 0.012825f
C98 VDD1.n5 B 0.086061f
C99 VDD1.t5 B 0.047393f
C100 VDD1.n6 B 0.021472f
C101 VDD1.n7 B 0.01685f
C102 VDD1.n8 B 0.012112f
C103 VDD1.n9 B 0.315993f
C104 VDD1.n10 B 0.02254f
C105 VDD1.n11 B 0.012112f
C106 VDD1.n12 B 0.012825f
C107 VDD1.n13 B 0.028629f
C108 VDD1.n14 B 0.060094f
C109 VDD1.n15 B 0.012825f
C110 VDD1.n16 B 0.012112f
C111 VDD1.n17 B 0.05364f
C112 VDD1.n18 B 0.053346f
C113 VDD1.n19 B 0.030618f
C114 VDD1.n20 B 0.02254f
C115 VDD1.n21 B 0.012112f
C116 VDD1.n22 B 0.028629f
C117 VDD1.n23 B 0.012825f
C118 VDD1.n24 B 0.086061f
C119 VDD1.t0 B 0.047393f
C120 VDD1.n25 B 0.021472f
C121 VDD1.n26 B 0.01685f
C122 VDD1.n27 B 0.012112f
C123 VDD1.n28 B 0.315993f
C124 VDD1.n29 B 0.02254f
C125 VDD1.n30 B 0.012112f
C126 VDD1.n31 B 0.012825f
C127 VDD1.n32 B 0.028629f
C128 VDD1.n33 B 0.060094f
C129 VDD1.n34 B 0.012825f
C130 VDD1.n35 B 0.012112f
C131 VDD1.n36 B 0.05364f
C132 VDD1.n37 B 0.052813f
C133 VDD1.t1 B 0.069289f
C134 VDD1.t2 B 0.069289f
C135 VDD1.n38 B 0.544007f
C136 VDD1.n39 B 1.76476f
C137 VDD1.t3 B 0.069289f
C138 VDD1.t4 B 0.069289f
C139 VDD1.n40 B 0.54206f
C140 VDD1.n41 B 1.74003f
C141 VTAIL.t0 B 0.086935f
C142 VTAIL.t1 B 0.086935f
C143 VTAIL.n0 B 0.618404f
C144 VTAIL.n1 B 0.418877f
C145 VTAIL.n2 B 0.038416f
C146 VTAIL.n3 B 0.028281f
C147 VTAIL.n4 B 0.015197f
C148 VTAIL.n5 B 0.03592f
C149 VTAIL.n6 B 0.016091f
C150 VTAIL.n7 B 0.107979f
C151 VTAIL.t9 B 0.059463f
C152 VTAIL.n8 B 0.02694f
C153 VTAIL.n9 B 0.021141f
C154 VTAIL.n10 B 0.015197f
C155 VTAIL.n11 B 0.396469f
C156 VTAIL.n12 B 0.028281f
C157 VTAIL.n13 B 0.015197f
C158 VTAIL.n14 B 0.016091f
C159 VTAIL.n15 B 0.03592f
C160 VTAIL.n16 B 0.075398f
C161 VTAIL.n17 B 0.016091f
C162 VTAIL.n18 B 0.015197f
C163 VTAIL.n19 B 0.067301f
C164 VTAIL.n20 B 0.042004f
C165 VTAIL.n21 B 0.324943f
C166 VTAIL.t7 B 0.086935f
C167 VTAIL.t8 B 0.086935f
C168 VTAIL.n22 B 0.618404f
C169 VTAIL.n23 B 1.44584f
C170 VTAIL.t3 B 0.086935f
C171 VTAIL.t2 B 0.086935f
C172 VTAIL.n24 B 0.618409f
C173 VTAIL.n25 B 1.44583f
C174 VTAIL.n26 B 0.038416f
C175 VTAIL.n27 B 0.028281f
C176 VTAIL.n28 B 0.015197f
C177 VTAIL.n29 B 0.03592f
C178 VTAIL.n30 B 0.016091f
C179 VTAIL.n31 B 0.107979f
C180 VTAIL.t4 B 0.059463f
C181 VTAIL.n32 B 0.02694f
C182 VTAIL.n33 B 0.021141f
C183 VTAIL.n34 B 0.015197f
C184 VTAIL.n35 B 0.396469f
C185 VTAIL.n36 B 0.028281f
C186 VTAIL.n37 B 0.015197f
C187 VTAIL.n38 B 0.016091f
C188 VTAIL.n39 B 0.03592f
C189 VTAIL.n40 B 0.075398f
C190 VTAIL.n41 B 0.016091f
C191 VTAIL.n42 B 0.015197f
C192 VTAIL.n43 B 0.067301f
C193 VTAIL.n44 B 0.042004f
C194 VTAIL.n45 B 0.324943f
C195 VTAIL.t11 B 0.086935f
C196 VTAIL.t10 B 0.086935f
C197 VTAIL.n46 B 0.618409f
C198 VTAIL.n47 B 0.542012f
C199 VTAIL.n48 B 0.038416f
C200 VTAIL.n49 B 0.028281f
C201 VTAIL.n50 B 0.015197f
C202 VTAIL.n51 B 0.03592f
C203 VTAIL.n52 B 0.016091f
C204 VTAIL.n53 B 0.107979f
C205 VTAIL.t6 B 0.059463f
C206 VTAIL.n54 B 0.02694f
C207 VTAIL.n55 B 0.021141f
C208 VTAIL.n56 B 0.015197f
C209 VTAIL.n57 B 0.396469f
C210 VTAIL.n58 B 0.028281f
C211 VTAIL.n59 B 0.015197f
C212 VTAIL.n60 B 0.016091f
C213 VTAIL.n61 B 0.03592f
C214 VTAIL.n62 B 0.075398f
C215 VTAIL.n63 B 0.016091f
C216 VTAIL.n64 B 0.015197f
C217 VTAIL.n65 B 0.067301f
C218 VTAIL.n66 B 0.042004f
C219 VTAIL.n67 B 1.05751f
C220 VTAIL.n68 B 0.038416f
C221 VTAIL.n69 B 0.028281f
C222 VTAIL.n70 B 0.015197f
C223 VTAIL.n71 B 0.03592f
C224 VTAIL.n72 B 0.016091f
C225 VTAIL.n73 B 0.107979f
C226 VTAIL.t5 B 0.059463f
C227 VTAIL.n74 B 0.02694f
C228 VTAIL.n75 B 0.021141f
C229 VTAIL.n76 B 0.015197f
C230 VTAIL.n77 B 0.396469f
C231 VTAIL.n78 B 0.028281f
C232 VTAIL.n79 B 0.015197f
C233 VTAIL.n80 B 0.016091f
C234 VTAIL.n81 B 0.03592f
C235 VTAIL.n82 B 0.075398f
C236 VTAIL.n83 B 0.016091f
C237 VTAIL.n84 B 0.015197f
C238 VTAIL.n85 B 0.067301f
C239 VTAIL.n86 B 0.042004f
C240 VTAIL.n87 B 1.00939f
C241 VP.n0 B 0.044853f
C242 VP.t3 B 0.626161f
C243 VP.n1 B 0.058113f
C244 VP.n2 B 0.034021f
C245 VP.t4 B 0.626161f
C246 VP.n3 B 0.04062f
C247 VP.n4 B 0.044853f
C248 VP.t1 B 0.626161f
C249 VP.n5 B 0.058113f
C250 VP.t0 B 0.783423f
C251 VP.n6 B 0.337234f
C252 VP.t2 B 0.626161f
C253 VP.n7 B 0.337072f
C254 VP.n8 B 0.047754f
C255 VP.n9 B 0.250157f
C256 VP.n10 B 0.034021f
C257 VP.n11 B 0.034021f
C258 VP.n12 B 0.04062f
C259 VP.n13 B 0.059619f
C260 VP.n14 B 0.359039f
C261 VP.n15 B 1.29631f
C262 VP.n16 B 1.3272f
C263 VP.t5 B 0.626161f
C264 VP.n17 B 0.359039f
C265 VP.n18 B 0.059619f
C266 VP.n19 B 0.044853f
C267 VP.n20 B 0.034021f
C268 VP.n21 B 0.034021f
C269 VP.n22 B 0.058113f
C270 VP.n23 B 0.047754f
C271 VP.n24 B 0.260014f
C272 VP.n25 B 0.047754f
C273 VP.n26 B 0.034021f
C274 VP.n27 B 0.034021f
C275 VP.n28 B 0.034021f
C276 VP.n29 B 0.04062f
C277 VP.n30 B 0.059619f
C278 VP.n31 B 0.359039f
C279 VP.n32 B 0.039305f
.ends

