* NGSPICE file created from diff_pair_sample_0403.ext - technology: sky130A

.subckt diff_pair_sample_0403 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VN.t0 VDD2.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=0.97845 ps=6.26 w=5.93 l=1.6
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=2.3127 pd=12.64 as=0 ps=0 w=5.93 l=1.6
X2 VTAIL.t15 VP.t0 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3127 pd=12.64 as=0.97845 ps=6.26 w=5.93 l=1.6
X3 VDD1.t6 VP.t1 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=2.3127 ps=12.64 w=5.93 l=1.6
X4 VDD2.t0 VN.t1 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=0.97845 ps=6.26 w=5.93 l=1.6
X5 VDD2.t1 VN.t2 VTAIL.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=0.97845 ps=6.26 w=5.93 l=1.6
X6 VTAIL.t6 VN.t3 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=0.97845 ps=6.26 w=5.93 l=1.6
X7 VDD1.t5 VP.t2 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=2.3127 ps=12.64 w=5.93 l=1.6
X8 VDD1.t4 VP.t3 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=0.97845 ps=6.26 w=5.93 l=1.6
X9 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.3127 pd=12.64 as=0 ps=0 w=5.93 l=1.6
X10 VDD2.t4 VN.t4 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=2.3127 ps=12.64 w=5.93 l=1.6
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=2.3127 pd=12.64 as=0 ps=0 w=5.93 l=1.6
X12 VDD2.t7 VN.t5 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=2.3127 ps=12.64 w=5.93 l=1.6
X13 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.3127 pd=12.64 as=0 ps=0 w=5.93 l=1.6
X14 VTAIL.t0 VP.t4 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=0.97845 ps=6.26 w=5.93 l=1.6
X15 VTAIL.t1 VP.t5 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3127 pd=12.64 as=0.97845 ps=6.26 w=5.93 l=1.6
X16 VTAIL.t3 VN.t6 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.3127 pd=12.64 as=0.97845 ps=6.26 w=5.93 l=1.6
X17 VTAIL.t11 VP.t6 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=0.97845 ps=6.26 w=5.93 l=1.6
X18 VDD1.t0 VP.t7 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.97845 pd=6.26 as=0.97845 ps=6.26 w=5.93 l=1.6
X19 VTAIL.t2 VN.t7 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3127 pd=12.64 as=0.97845 ps=6.26 w=5.93 l=1.6
R0 VN.n20 VN.n19 178.673
R1 VN.n41 VN.n40 178.673
R2 VN.n39 VN.n21 161.3
R3 VN.n38 VN.n37 161.3
R4 VN.n36 VN.n22 161.3
R5 VN.n35 VN.n34 161.3
R6 VN.n32 VN.n23 161.3
R7 VN.n31 VN.n30 161.3
R8 VN.n29 VN.n24 161.3
R9 VN.n28 VN.n27 161.3
R10 VN.n18 VN.n0 161.3
R11 VN.n17 VN.n16 161.3
R12 VN.n15 VN.n1 161.3
R13 VN.n14 VN.n13 161.3
R14 VN.n11 VN.n2 161.3
R15 VN.n10 VN.n9 161.3
R16 VN.n8 VN.n3 161.3
R17 VN.n7 VN.n6 161.3
R18 VN.n4 VN.t7 121.507
R19 VN.n25 VN.t4 121.507
R20 VN.n5 VN.t1 89.3211
R21 VN.n12 VN.t3 89.3211
R22 VN.n19 VN.t5 89.3211
R23 VN.n26 VN.t0 89.3211
R24 VN.n33 VN.t2 89.3211
R25 VN.n40 VN.t6 89.3211
R26 VN.n17 VN.n1 56.5193
R27 VN.n38 VN.n22 56.5193
R28 VN.n10 VN.n3 56.5193
R29 VN.n31 VN.n24 56.5193
R30 VN.n5 VN.n4 55.5644
R31 VN.n26 VN.n25 55.5644
R32 VN VN.n41 41.9039
R33 VN.n6 VN.n3 24.4675
R34 VN.n11 VN.n10 24.4675
R35 VN.n13 VN.n1 24.4675
R36 VN.n18 VN.n17 24.4675
R37 VN.n27 VN.n24 24.4675
R38 VN.n34 VN.n22 24.4675
R39 VN.n32 VN.n31 24.4675
R40 VN.n39 VN.n38 24.4675
R41 VN.n28 VN.n25 18.0716
R42 VN.n7 VN.n4 18.0716
R43 VN.n13 VN.n12 13.9467
R44 VN.n34 VN.n33 13.9467
R45 VN.n6 VN.n5 10.5213
R46 VN.n12 VN.n11 10.5213
R47 VN.n27 VN.n26 10.5213
R48 VN.n33 VN.n32 10.5213
R49 VN.n19 VN.n18 7.09593
R50 VN.n40 VN.n39 7.09593
R51 VN.n41 VN.n21 0.189894
R52 VN.n37 VN.n21 0.189894
R53 VN.n37 VN.n36 0.189894
R54 VN.n36 VN.n35 0.189894
R55 VN.n35 VN.n23 0.189894
R56 VN.n30 VN.n23 0.189894
R57 VN.n30 VN.n29 0.189894
R58 VN.n29 VN.n28 0.189894
R59 VN.n8 VN.n7 0.189894
R60 VN.n9 VN.n8 0.189894
R61 VN.n9 VN.n2 0.189894
R62 VN.n14 VN.n2 0.189894
R63 VN.n15 VN.n14 0.189894
R64 VN.n16 VN.n15 0.189894
R65 VN.n16 VN.n0 0.189894
R66 VN.n20 VN.n0 0.189894
R67 VN VN.n20 0.0516364
R68 VDD2.n2 VDD2.n1 66.6096
R69 VDD2.n2 VDD2.n0 66.6096
R70 VDD2 VDD2.n5 66.6068
R71 VDD2.n4 VDD2.n3 65.8332
R72 VDD2.n4 VDD2.n2 36.3144
R73 VDD2.n5 VDD2.t5 3.33945
R74 VDD2.n5 VDD2.t4 3.33945
R75 VDD2.n3 VDD2.t2 3.33945
R76 VDD2.n3 VDD2.t1 3.33945
R77 VDD2.n1 VDD2.t6 3.33945
R78 VDD2.n1 VDD2.t7 3.33945
R79 VDD2.n0 VDD2.t3 3.33945
R80 VDD2.n0 VDD2.t0 3.33945
R81 VDD2 VDD2.n4 0.890586
R82 VTAIL.n258 VTAIL.n232 289.615
R83 VTAIL.n28 VTAIL.n2 289.615
R84 VTAIL.n60 VTAIL.n34 289.615
R85 VTAIL.n94 VTAIL.n68 289.615
R86 VTAIL.n226 VTAIL.n200 289.615
R87 VTAIL.n192 VTAIL.n166 289.615
R88 VTAIL.n160 VTAIL.n134 289.615
R89 VTAIL.n126 VTAIL.n100 289.615
R90 VTAIL.n243 VTAIL.n242 185
R91 VTAIL.n240 VTAIL.n239 185
R92 VTAIL.n249 VTAIL.n248 185
R93 VTAIL.n251 VTAIL.n250 185
R94 VTAIL.n236 VTAIL.n235 185
R95 VTAIL.n257 VTAIL.n256 185
R96 VTAIL.n259 VTAIL.n258 185
R97 VTAIL.n13 VTAIL.n12 185
R98 VTAIL.n10 VTAIL.n9 185
R99 VTAIL.n19 VTAIL.n18 185
R100 VTAIL.n21 VTAIL.n20 185
R101 VTAIL.n6 VTAIL.n5 185
R102 VTAIL.n27 VTAIL.n26 185
R103 VTAIL.n29 VTAIL.n28 185
R104 VTAIL.n45 VTAIL.n44 185
R105 VTAIL.n42 VTAIL.n41 185
R106 VTAIL.n51 VTAIL.n50 185
R107 VTAIL.n53 VTAIL.n52 185
R108 VTAIL.n38 VTAIL.n37 185
R109 VTAIL.n59 VTAIL.n58 185
R110 VTAIL.n61 VTAIL.n60 185
R111 VTAIL.n79 VTAIL.n78 185
R112 VTAIL.n76 VTAIL.n75 185
R113 VTAIL.n85 VTAIL.n84 185
R114 VTAIL.n87 VTAIL.n86 185
R115 VTAIL.n72 VTAIL.n71 185
R116 VTAIL.n93 VTAIL.n92 185
R117 VTAIL.n95 VTAIL.n94 185
R118 VTAIL.n227 VTAIL.n226 185
R119 VTAIL.n225 VTAIL.n224 185
R120 VTAIL.n204 VTAIL.n203 185
R121 VTAIL.n219 VTAIL.n218 185
R122 VTAIL.n217 VTAIL.n216 185
R123 VTAIL.n208 VTAIL.n207 185
R124 VTAIL.n211 VTAIL.n210 185
R125 VTAIL.n193 VTAIL.n192 185
R126 VTAIL.n191 VTAIL.n190 185
R127 VTAIL.n170 VTAIL.n169 185
R128 VTAIL.n185 VTAIL.n184 185
R129 VTAIL.n183 VTAIL.n182 185
R130 VTAIL.n174 VTAIL.n173 185
R131 VTAIL.n177 VTAIL.n176 185
R132 VTAIL.n161 VTAIL.n160 185
R133 VTAIL.n159 VTAIL.n158 185
R134 VTAIL.n138 VTAIL.n137 185
R135 VTAIL.n153 VTAIL.n152 185
R136 VTAIL.n151 VTAIL.n150 185
R137 VTAIL.n142 VTAIL.n141 185
R138 VTAIL.n145 VTAIL.n144 185
R139 VTAIL.n127 VTAIL.n126 185
R140 VTAIL.n125 VTAIL.n124 185
R141 VTAIL.n104 VTAIL.n103 185
R142 VTAIL.n119 VTAIL.n118 185
R143 VTAIL.n117 VTAIL.n116 185
R144 VTAIL.n108 VTAIL.n107 185
R145 VTAIL.n111 VTAIL.n110 185
R146 VTAIL.t4 VTAIL.n241 147.661
R147 VTAIL.t2 VTAIL.n11 147.661
R148 VTAIL.t12 VTAIL.n43 147.661
R149 VTAIL.t1 VTAIL.n77 147.661
R150 VTAIL.t14 VTAIL.n209 147.661
R151 VTAIL.t15 VTAIL.n175 147.661
R152 VTAIL.t5 VTAIL.n143 147.661
R153 VTAIL.t3 VTAIL.n109 147.661
R154 VTAIL.n242 VTAIL.n239 104.615
R155 VTAIL.n249 VTAIL.n239 104.615
R156 VTAIL.n250 VTAIL.n249 104.615
R157 VTAIL.n250 VTAIL.n235 104.615
R158 VTAIL.n257 VTAIL.n235 104.615
R159 VTAIL.n258 VTAIL.n257 104.615
R160 VTAIL.n12 VTAIL.n9 104.615
R161 VTAIL.n19 VTAIL.n9 104.615
R162 VTAIL.n20 VTAIL.n19 104.615
R163 VTAIL.n20 VTAIL.n5 104.615
R164 VTAIL.n27 VTAIL.n5 104.615
R165 VTAIL.n28 VTAIL.n27 104.615
R166 VTAIL.n44 VTAIL.n41 104.615
R167 VTAIL.n51 VTAIL.n41 104.615
R168 VTAIL.n52 VTAIL.n51 104.615
R169 VTAIL.n52 VTAIL.n37 104.615
R170 VTAIL.n59 VTAIL.n37 104.615
R171 VTAIL.n60 VTAIL.n59 104.615
R172 VTAIL.n78 VTAIL.n75 104.615
R173 VTAIL.n85 VTAIL.n75 104.615
R174 VTAIL.n86 VTAIL.n85 104.615
R175 VTAIL.n86 VTAIL.n71 104.615
R176 VTAIL.n93 VTAIL.n71 104.615
R177 VTAIL.n94 VTAIL.n93 104.615
R178 VTAIL.n226 VTAIL.n225 104.615
R179 VTAIL.n225 VTAIL.n203 104.615
R180 VTAIL.n218 VTAIL.n203 104.615
R181 VTAIL.n218 VTAIL.n217 104.615
R182 VTAIL.n217 VTAIL.n207 104.615
R183 VTAIL.n210 VTAIL.n207 104.615
R184 VTAIL.n192 VTAIL.n191 104.615
R185 VTAIL.n191 VTAIL.n169 104.615
R186 VTAIL.n184 VTAIL.n169 104.615
R187 VTAIL.n184 VTAIL.n183 104.615
R188 VTAIL.n183 VTAIL.n173 104.615
R189 VTAIL.n176 VTAIL.n173 104.615
R190 VTAIL.n160 VTAIL.n159 104.615
R191 VTAIL.n159 VTAIL.n137 104.615
R192 VTAIL.n152 VTAIL.n137 104.615
R193 VTAIL.n152 VTAIL.n151 104.615
R194 VTAIL.n151 VTAIL.n141 104.615
R195 VTAIL.n144 VTAIL.n141 104.615
R196 VTAIL.n126 VTAIL.n125 104.615
R197 VTAIL.n125 VTAIL.n103 104.615
R198 VTAIL.n118 VTAIL.n103 104.615
R199 VTAIL.n118 VTAIL.n117 104.615
R200 VTAIL.n117 VTAIL.n107 104.615
R201 VTAIL.n110 VTAIL.n107 104.615
R202 VTAIL.n242 VTAIL.t4 52.3082
R203 VTAIL.n12 VTAIL.t2 52.3082
R204 VTAIL.n44 VTAIL.t12 52.3082
R205 VTAIL.n78 VTAIL.t1 52.3082
R206 VTAIL.n210 VTAIL.t14 52.3082
R207 VTAIL.n176 VTAIL.t15 52.3082
R208 VTAIL.n144 VTAIL.t5 52.3082
R209 VTAIL.n110 VTAIL.t3 52.3082
R210 VTAIL.n199 VTAIL.n198 49.1545
R211 VTAIL.n133 VTAIL.n132 49.1545
R212 VTAIL.n1 VTAIL.n0 49.1543
R213 VTAIL.n67 VTAIL.n66 49.1543
R214 VTAIL.n263 VTAIL.n262 30.8278
R215 VTAIL.n33 VTAIL.n32 30.8278
R216 VTAIL.n65 VTAIL.n64 30.8278
R217 VTAIL.n99 VTAIL.n98 30.8278
R218 VTAIL.n231 VTAIL.n230 30.8278
R219 VTAIL.n197 VTAIL.n196 30.8278
R220 VTAIL.n165 VTAIL.n164 30.8278
R221 VTAIL.n131 VTAIL.n130 30.8278
R222 VTAIL.n263 VTAIL.n231 19.1427
R223 VTAIL.n131 VTAIL.n99 19.1427
R224 VTAIL.n243 VTAIL.n241 15.6674
R225 VTAIL.n13 VTAIL.n11 15.6674
R226 VTAIL.n45 VTAIL.n43 15.6674
R227 VTAIL.n79 VTAIL.n77 15.6674
R228 VTAIL.n211 VTAIL.n209 15.6674
R229 VTAIL.n177 VTAIL.n175 15.6674
R230 VTAIL.n145 VTAIL.n143 15.6674
R231 VTAIL.n111 VTAIL.n109 15.6674
R232 VTAIL.n244 VTAIL.n240 12.8005
R233 VTAIL.n14 VTAIL.n10 12.8005
R234 VTAIL.n46 VTAIL.n42 12.8005
R235 VTAIL.n80 VTAIL.n76 12.8005
R236 VTAIL.n212 VTAIL.n208 12.8005
R237 VTAIL.n178 VTAIL.n174 12.8005
R238 VTAIL.n146 VTAIL.n142 12.8005
R239 VTAIL.n112 VTAIL.n108 12.8005
R240 VTAIL.n248 VTAIL.n247 12.0247
R241 VTAIL.n18 VTAIL.n17 12.0247
R242 VTAIL.n50 VTAIL.n49 12.0247
R243 VTAIL.n84 VTAIL.n83 12.0247
R244 VTAIL.n216 VTAIL.n215 12.0247
R245 VTAIL.n182 VTAIL.n181 12.0247
R246 VTAIL.n150 VTAIL.n149 12.0247
R247 VTAIL.n116 VTAIL.n115 12.0247
R248 VTAIL.n251 VTAIL.n238 11.249
R249 VTAIL.n21 VTAIL.n8 11.249
R250 VTAIL.n53 VTAIL.n40 11.249
R251 VTAIL.n87 VTAIL.n74 11.249
R252 VTAIL.n219 VTAIL.n206 11.249
R253 VTAIL.n185 VTAIL.n172 11.249
R254 VTAIL.n153 VTAIL.n140 11.249
R255 VTAIL.n119 VTAIL.n106 11.249
R256 VTAIL.n252 VTAIL.n236 10.4732
R257 VTAIL.n22 VTAIL.n6 10.4732
R258 VTAIL.n54 VTAIL.n38 10.4732
R259 VTAIL.n88 VTAIL.n72 10.4732
R260 VTAIL.n220 VTAIL.n204 10.4732
R261 VTAIL.n186 VTAIL.n170 10.4732
R262 VTAIL.n154 VTAIL.n138 10.4732
R263 VTAIL.n120 VTAIL.n104 10.4732
R264 VTAIL.n256 VTAIL.n255 9.69747
R265 VTAIL.n26 VTAIL.n25 9.69747
R266 VTAIL.n58 VTAIL.n57 9.69747
R267 VTAIL.n92 VTAIL.n91 9.69747
R268 VTAIL.n224 VTAIL.n223 9.69747
R269 VTAIL.n190 VTAIL.n189 9.69747
R270 VTAIL.n158 VTAIL.n157 9.69747
R271 VTAIL.n124 VTAIL.n123 9.69747
R272 VTAIL.n262 VTAIL.n261 9.45567
R273 VTAIL.n32 VTAIL.n31 9.45567
R274 VTAIL.n64 VTAIL.n63 9.45567
R275 VTAIL.n98 VTAIL.n97 9.45567
R276 VTAIL.n230 VTAIL.n229 9.45567
R277 VTAIL.n196 VTAIL.n195 9.45567
R278 VTAIL.n164 VTAIL.n163 9.45567
R279 VTAIL.n130 VTAIL.n129 9.45567
R280 VTAIL.n261 VTAIL.n260 9.3005
R281 VTAIL.n234 VTAIL.n233 9.3005
R282 VTAIL.n255 VTAIL.n254 9.3005
R283 VTAIL.n253 VTAIL.n252 9.3005
R284 VTAIL.n238 VTAIL.n237 9.3005
R285 VTAIL.n247 VTAIL.n246 9.3005
R286 VTAIL.n245 VTAIL.n244 9.3005
R287 VTAIL.n31 VTAIL.n30 9.3005
R288 VTAIL.n4 VTAIL.n3 9.3005
R289 VTAIL.n25 VTAIL.n24 9.3005
R290 VTAIL.n23 VTAIL.n22 9.3005
R291 VTAIL.n8 VTAIL.n7 9.3005
R292 VTAIL.n17 VTAIL.n16 9.3005
R293 VTAIL.n15 VTAIL.n14 9.3005
R294 VTAIL.n63 VTAIL.n62 9.3005
R295 VTAIL.n36 VTAIL.n35 9.3005
R296 VTAIL.n57 VTAIL.n56 9.3005
R297 VTAIL.n55 VTAIL.n54 9.3005
R298 VTAIL.n40 VTAIL.n39 9.3005
R299 VTAIL.n49 VTAIL.n48 9.3005
R300 VTAIL.n47 VTAIL.n46 9.3005
R301 VTAIL.n97 VTAIL.n96 9.3005
R302 VTAIL.n70 VTAIL.n69 9.3005
R303 VTAIL.n91 VTAIL.n90 9.3005
R304 VTAIL.n89 VTAIL.n88 9.3005
R305 VTAIL.n74 VTAIL.n73 9.3005
R306 VTAIL.n83 VTAIL.n82 9.3005
R307 VTAIL.n81 VTAIL.n80 9.3005
R308 VTAIL.n229 VTAIL.n228 9.3005
R309 VTAIL.n202 VTAIL.n201 9.3005
R310 VTAIL.n223 VTAIL.n222 9.3005
R311 VTAIL.n221 VTAIL.n220 9.3005
R312 VTAIL.n206 VTAIL.n205 9.3005
R313 VTAIL.n215 VTAIL.n214 9.3005
R314 VTAIL.n213 VTAIL.n212 9.3005
R315 VTAIL.n195 VTAIL.n194 9.3005
R316 VTAIL.n168 VTAIL.n167 9.3005
R317 VTAIL.n189 VTAIL.n188 9.3005
R318 VTAIL.n187 VTAIL.n186 9.3005
R319 VTAIL.n172 VTAIL.n171 9.3005
R320 VTAIL.n181 VTAIL.n180 9.3005
R321 VTAIL.n179 VTAIL.n178 9.3005
R322 VTAIL.n163 VTAIL.n162 9.3005
R323 VTAIL.n136 VTAIL.n135 9.3005
R324 VTAIL.n157 VTAIL.n156 9.3005
R325 VTAIL.n155 VTAIL.n154 9.3005
R326 VTAIL.n140 VTAIL.n139 9.3005
R327 VTAIL.n149 VTAIL.n148 9.3005
R328 VTAIL.n147 VTAIL.n146 9.3005
R329 VTAIL.n129 VTAIL.n128 9.3005
R330 VTAIL.n102 VTAIL.n101 9.3005
R331 VTAIL.n123 VTAIL.n122 9.3005
R332 VTAIL.n121 VTAIL.n120 9.3005
R333 VTAIL.n106 VTAIL.n105 9.3005
R334 VTAIL.n115 VTAIL.n114 9.3005
R335 VTAIL.n113 VTAIL.n112 9.3005
R336 VTAIL.n259 VTAIL.n234 8.92171
R337 VTAIL.n29 VTAIL.n4 8.92171
R338 VTAIL.n61 VTAIL.n36 8.92171
R339 VTAIL.n95 VTAIL.n70 8.92171
R340 VTAIL.n227 VTAIL.n202 8.92171
R341 VTAIL.n193 VTAIL.n168 8.92171
R342 VTAIL.n161 VTAIL.n136 8.92171
R343 VTAIL.n127 VTAIL.n102 8.92171
R344 VTAIL.n260 VTAIL.n232 8.14595
R345 VTAIL.n30 VTAIL.n2 8.14595
R346 VTAIL.n62 VTAIL.n34 8.14595
R347 VTAIL.n96 VTAIL.n68 8.14595
R348 VTAIL.n228 VTAIL.n200 8.14595
R349 VTAIL.n194 VTAIL.n166 8.14595
R350 VTAIL.n162 VTAIL.n134 8.14595
R351 VTAIL.n128 VTAIL.n100 8.14595
R352 VTAIL.n262 VTAIL.n232 5.81868
R353 VTAIL.n32 VTAIL.n2 5.81868
R354 VTAIL.n64 VTAIL.n34 5.81868
R355 VTAIL.n98 VTAIL.n68 5.81868
R356 VTAIL.n230 VTAIL.n200 5.81868
R357 VTAIL.n196 VTAIL.n166 5.81868
R358 VTAIL.n164 VTAIL.n134 5.81868
R359 VTAIL.n130 VTAIL.n100 5.81868
R360 VTAIL.n260 VTAIL.n259 5.04292
R361 VTAIL.n30 VTAIL.n29 5.04292
R362 VTAIL.n62 VTAIL.n61 5.04292
R363 VTAIL.n96 VTAIL.n95 5.04292
R364 VTAIL.n228 VTAIL.n227 5.04292
R365 VTAIL.n194 VTAIL.n193 5.04292
R366 VTAIL.n162 VTAIL.n161 5.04292
R367 VTAIL.n128 VTAIL.n127 5.04292
R368 VTAIL.n245 VTAIL.n241 4.38594
R369 VTAIL.n15 VTAIL.n11 4.38594
R370 VTAIL.n47 VTAIL.n43 4.38594
R371 VTAIL.n81 VTAIL.n77 4.38594
R372 VTAIL.n213 VTAIL.n209 4.38594
R373 VTAIL.n179 VTAIL.n175 4.38594
R374 VTAIL.n147 VTAIL.n143 4.38594
R375 VTAIL.n113 VTAIL.n109 4.38594
R376 VTAIL.n256 VTAIL.n234 4.26717
R377 VTAIL.n26 VTAIL.n4 4.26717
R378 VTAIL.n58 VTAIL.n36 4.26717
R379 VTAIL.n92 VTAIL.n70 4.26717
R380 VTAIL.n224 VTAIL.n202 4.26717
R381 VTAIL.n190 VTAIL.n168 4.26717
R382 VTAIL.n158 VTAIL.n136 4.26717
R383 VTAIL.n124 VTAIL.n102 4.26717
R384 VTAIL.n255 VTAIL.n236 3.49141
R385 VTAIL.n25 VTAIL.n6 3.49141
R386 VTAIL.n57 VTAIL.n38 3.49141
R387 VTAIL.n91 VTAIL.n72 3.49141
R388 VTAIL.n223 VTAIL.n204 3.49141
R389 VTAIL.n189 VTAIL.n170 3.49141
R390 VTAIL.n157 VTAIL.n138 3.49141
R391 VTAIL.n123 VTAIL.n104 3.49141
R392 VTAIL.n0 VTAIL.t8 3.33945
R393 VTAIL.n0 VTAIL.t6 3.33945
R394 VTAIL.n66 VTAIL.t10 3.33945
R395 VTAIL.n66 VTAIL.t11 3.33945
R396 VTAIL.n198 VTAIL.t13 3.33945
R397 VTAIL.n198 VTAIL.t0 3.33945
R398 VTAIL.n132 VTAIL.t7 3.33945
R399 VTAIL.n132 VTAIL.t9 3.33945
R400 VTAIL.n252 VTAIL.n251 2.71565
R401 VTAIL.n22 VTAIL.n21 2.71565
R402 VTAIL.n54 VTAIL.n53 2.71565
R403 VTAIL.n88 VTAIL.n87 2.71565
R404 VTAIL.n220 VTAIL.n219 2.71565
R405 VTAIL.n186 VTAIL.n185 2.71565
R406 VTAIL.n154 VTAIL.n153 2.71565
R407 VTAIL.n120 VTAIL.n119 2.71565
R408 VTAIL.n248 VTAIL.n238 1.93989
R409 VTAIL.n18 VTAIL.n8 1.93989
R410 VTAIL.n50 VTAIL.n40 1.93989
R411 VTAIL.n84 VTAIL.n74 1.93989
R412 VTAIL.n216 VTAIL.n206 1.93989
R413 VTAIL.n182 VTAIL.n172 1.93989
R414 VTAIL.n150 VTAIL.n140 1.93989
R415 VTAIL.n116 VTAIL.n106 1.93989
R416 VTAIL.n133 VTAIL.n131 1.66429
R417 VTAIL.n165 VTAIL.n133 1.66429
R418 VTAIL.n199 VTAIL.n197 1.66429
R419 VTAIL.n231 VTAIL.n199 1.66429
R420 VTAIL.n99 VTAIL.n67 1.66429
R421 VTAIL.n67 VTAIL.n65 1.66429
R422 VTAIL.n33 VTAIL.n1 1.66429
R423 VTAIL VTAIL.n263 1.6061
R424 VTAIL.n247 VTAIL.n240 1.16414
R425 VTAIL.n17 VTAIL.n10 1.16414
R426 VTAIL.n49 VTAIL.n42 1.16414
R427 VTAIL.n83 VTAIL.n76 1.16414
R428 VTAIL.n215 VTAIL.n208 1.16414
R429 VTAIL.n181 VTAIL.n174 1.16414
R430 VTAIL.n149 VTAIL.n142 1.16414
R431 VTAIL.n115 VTAIL.n108 1.16414
R432 VTAIL.n197 VTAIL.n165 0.470328
R433 VTAIL.n65 VTAIL.n33 0.470328
R434 VTAIL.n244 VTAIL.n243 0.388379
R435 VTAIL.n14 VTAIL.n13 0.388379
R436 VTAIL.n46 VTAIL.n45 0.388379
R437 VTAIL.n80 VTAIL.n79 0.388379
R438 VTAIL.n212 VTAIL.n211 0.388379
R439 VTAIL.n178 VTAIL.n177 0.388379
R440 VTAIL.n146 VTAIL.n145 0.388379
R441 VTAIL.n112 VTAIL.n111 0.388379
R442 VTAIL.n246 VTAIL.n245 0.155672
R443 VTAIL.n246 VTAIL.n237 0.155672
R444 VTAIL.n253 VTAIL.n237 0.155672
R445 VTAIL.n254 VTAIL.n253 0.155672
R446 VTAIL.n254 VTAIL.n233 0.155672
R447 VTAIL.n261 VTAIL.n233 0.155672
R448 VTAIL.n16 VTAIL.n15 0.155672
R449 VTAIL.n16 VTAIL.n7 0.155672
R450 VTAIL.n23 VTAIL.n7 0.155672
R451 VTAIL.n24 VTAIL.n23 0.155672
R452 VTAIL.n24 VTAIL.n3 0.155672
R453 VTAIL.n31 VTAIL.n3 0.155672
R454 VTAIL.n48 VTAIL.n47 0.155672
R455 VTAIL.n48 VTAIL.n39 0.155672
R456 VTAIL.n55 VTAIL.n39 0.155672
R457 VTAIL.n56 VTAIL.n55 0.155672
R458 VTAIL.n56 VTAIL.n35 0.155672
R459 VTAIL.n63 VTAIL.n35 0.155672
R460 VTAIL.n82 VTAIL.n81 0.155672
R461 VTAIL.n82 VTAIL.n73 0.155672
R462 VTAIL.n89 VTAIL.n73 0.155672
R463 VTAIL.n90 VTAIL.n89 0.155672
R464 VTAIL.n90 VTAIL.n69 0.155672
R465 VTAIL.n97 VTAIL.n69 0.155672
R466 VTAIL.n229 VTAIL.n201 0.155672
R467 VTAIL.n222 VTAIL.n201 0.155672
R468 VTAIL.n222 VTAIL.n221 0.155672
R469 VTAIL.n221 VTAIL.n205 0.155672
R470 VTAIL.n214 VTAIL.n205 0.155672
R471 VTAIL.n214 VTAIL.n213 0.155672
R472 VTAIL.n195 VTAIL.n167 0.155672
R473 VTAIL.n188 VTAIL.n167 0.155672
R474 VTAIL.n188 VTAIL.n187 0.155672
R475 VTAIL.n187 VTAIL.n171 0.155672
R476 VTAIL.n180 VTAIL.n171 0.155672
R477 VTAIL.n180 VTAIL.n179 0.155672
R478 VTAIL.n163 VTAIL.n135 0.155672
R479 VTAIL.n156 VTAIL.n135 0.155672
R480 VTAIL.n156 VTAIL.n155 0.155672
R481 VTAIL.n155 VTAIL.n139 0.155672
R482 VTAIL.n148 VTAIL.n139 0.155672
R483 VTAIL.n148 VTAIL.n147 0.155672
R484 VTAIL.n129 VTAIL.n101 0.155672
R485 VTAIL.n122 VTAIL.n101 0.155672
R486 VTAIL.n122 VTAIL.n121 0.155672
R487 VTAIL.n121 VTAIL.n105 0.155672
R488 VTAIL.n114 VTAIL.n105 0.155672
R489 VTAIL.n114 VTAIL.n113 0.155672
R490 VTAIL VTAIL.n1 0.0586897
R491 B.n589 B.n588 585
R492 B.n590 B.n589 585
R493 B.n212 B.n97 585
R494 B.n211 B.n210 585
R495 B.n209 B.n208 585
R496 B.n207 B.n206 585
R497 B.n205 B.n204 585
R498 B.n203 B.n202 585
R499 B.n201 B.n200 585
R500 B.n199 B.n198 585
R501 B.n197 B.n196 585
R502 B.n195 B.n194 585
R503 B.n193 B.n192 585
R504 B.n191 B.n190 585
R505 B.n189 B.n188 585
R506 B.n187 B.n186 585
R507 B.n185 B.n184 585
R508 B.n183 B.n182 585
R509 B.n181 B.n180 585
R510 B.n179 B.n178 585
R511 B.n177 B.n176 585
R512 B.n175 B.n174 585
R513 B.n173 B.n172 585
R514 B.n171 B.n170 585
R515 B.n169 B.n168 585
R516 B.n166 B.n165 585
R517 B.n164 B.n163 585
R518 B.n162 B.n161 585
R519 B.n160 B.n159 585
R520 B.n158 B.n157 585
R521 B.n156 B.n155 585
R522 B.n154 B.n153 585
R523 B.n152 B.n151 585
R524 B.n150 B.n149 585
R525 B.n148 B.n147 585
R526 B.n146 B.n145 585
R527 B.n144 B.n143 585
R528 B.n142 B.n141 585
R529 B.n140 B.n139 585
R530 B.n138 B.n137 585
R531 B.n136 B.n135 585
R532 B.n134 B.n133 585
R533 B.n132 B.n131 585
R534 B.n130 B.n129 585
R535 B.n128 B.n127 585
R536 B.n126 B.n125 585
R537 B.n124 B.n123 585
R538 B.n122 B.n121 585
R539 B.n120 B.n119 585
R540 B.n118 B.n117 585
R541 B.n116 B.n115 585
R542 B.n114 B.n113 585
R543 B.n112 B.n111 585
R544 B.n110 B.n109 585
R545 B.n108 B.n107 585
R546 B.n106 B.n105 585
R547 B.n104 B.n103 585
R548 B.n67 B.n66 585
R549 B.n587 B.n68 585
R550 B.n591 B.n68 585
R551 B.n586 B.n585 585
R552 B.n585 B.n64 585
R553 B.n584 B.n63 585
R554 B.n597 B.n63 585
R555 B.n583 B.n62 585
R556 B.n598 B.n62 585
R557 B.n582 B.n61 585
R558 B.n599 B.n61 585
R559 B.n581 B.n580 585
R560 B.n580 B.n57 585
R561 B.n579 B.n56 585
R562 B.n605 B.n56 585
R563 B.n578 B.n55 585
R564 B.n606 B.n55 585
R565 B.n577 B.n54 585
R566 B.n607 B.n54 585
R567 B.n576 B.n575 585
R568 B.n575 B.n50 585
R569 B.n574 B.n49 585
R570 B.n613 B.n49 585
R571 B.n573 B.n48 585
R572 B.n614 B.n48 585
R573 B.n572 B.n47 585
R574 B.n615 B.n47 585
R575 B.n571 B.n570 585
R576 B.n570 B.n43 585
R577 B.n569 B.n42 585
R578 B.n621 B.n42 585
R579 B.n568 B.n41 585
R580 B.n622 B.n41 585
R581 B.n567 B.n40 585
R582 B.n623 B.n40 585
R583 B.n566 B.n565 585
R584 B.n565 B.n36 585
R585 B.n564 B.n35 585
R586 B.n629 B.n35 585
R587 B.n563 B.n34 585
R588 B.n630 B.n34 585
R589 B.n562 B.n33 585
R590 B.n631 B.n33 585
R591 B.n561 B.n560 585
R592 B.n560 B.n29 585
R593 B.n559 B.n28 585
R594 B.n637 B.n28 585
R595 B.n558 B.n27 585
R596 B.n638 B.n27 585
R597 B.n557 B.n26 585
R598 B.n639 B.n26 585
R599 B.n556 B.n555 585
R600 B.n555 B.n22 585
R601 B.n554 B.n21 585
R602 B.n645 B.n21 585
R603 B.n553 B.n20 585
R604 B.n646 B.n20 585
R605 B.n552 B.n19 585
R606 B.n647 B.n19 585
R607 B.n551 B.n550 585
R608 B.n550 B.n15 585
R609 B.n549 B.n14 585
R610 B.n653 B.n14 585
R611 B.n548 B.n13 585
R612 B.n654 B.n13 585
R613 B.n547 B.n12 585
R614 B.n655 B.n12 585
R615 B.n546 B.n545 585
R616 B.n545 B.n544 585
R617 B.n543 B.n542 585
R618 B.n543 B.n8 585
R619 B.n541 B.n7 585
R620 B.n662 B.n7 585
R621 B.n540 B.n6 585
R622 B.n663 B.n6 585
R623 B.n539 B.n5 585
R624 B.n664 B.n5 585
R625 B.n538 B.n537 585
R626 B.n537 B.n4 585
R627 B.n536 B.n213 585
R628 B.n536 B.n535 585
R629 B.n526 B.n214 585
R630 B.n215 B.n214 585
R631 B.n528 B.n527 585
R632 B.n529 B.n528 585
R633 B.n525 B.n220 585
R634 B.n220 B.n219 585
R635 B.n524 B.n523 585
R636 B.n523 B.n522 585
R637 B.n222 B.n221 585
R638 B.n223 B.n222 585
R639 B.n515 B.n514 585
R640 B.n516 B.n515 585
R641 B.n513 B.n228 585
R642 B.n228 B.n227 585
R643 B.n512 B.n511 585
R644 B.n511 B.n510 585
R645 B.n230 B.n229 585
R646 B.n231 B.n230 585
R647 B.n503 B.n502 585
R648 B.n504 B.n503 585
R649 B.n501 B.n236 585
R650 B.n236 B.n235 585
R651 B.n500 B.n499 585
R652 B.n499 B.n498 585
R653 B.n238 B.n237 585
R654 B.n239 B.n238 585
R655 B.n491 B.n490 585
R656 B.n492 B.n491 585
R657 B.n489 B.n244 585
R658 B.n244 B.n243 585
R659 B.n488 B.n487 585
R660 B.n487 B.n486 585
R661 B.n246 B.n245 585
R662 B.n247 B.n246 585
R663 B.n479 B.n478 585
R664 B.n480 B.n479 585
R665 B.n477 B.n251 585
R666 B.n255 B.n251 585
R667 B.n476 B.n475 585
R668 B.n475 B.n474 585
R669 B.n253 B.n252 585
R670 B.n254 B.n253 585
R671 B.n467 B.n466 585
R672 B.n468 B.n467 585
R673 B.n465 B.n260 585
R674 B.n260 B.n259 585
R675 B.n464 B.n463 585
R676 B.n463 B.n462 585
R677 B.n262 B.n261 585
R678 B.n263 B.n262 585
R679 B.n455 B.n454 585
R680 B.n456 B.n455 585
R681 B.n453 B.n268 585
R682 B.n268 B.n267 585
R683 B.n452 B.n451 585
R684 B.n451 B.n450 585
R685 B.n270 B.n269 585
R686 B.n271 B.n270 585
R687 B.n443 B.n442 585
R688 B.n444 B.n443 585
R689 B.n441 B.n276 585
R690 B.n276 B.n275 585
R691 B.n440 B.n439 585
R692 B.n439 B.n438 585
R693 B.n278 B.n277 585
R694 B.n279 B.n278 585
R695 B.n431 B.n430 585
R696 B.n432 B.n431 585
R697 B.n282 B.n281 585
R698 B.n318 B.n316 585
R699 B.n319 B.n315 585
R700 B.n319 B.n283 585
R701 B.n322 B.n321 585
R702 B.n323 B.n314 585
R703 B.n325 B.n324 585
R704 B.n327 B.n313 585
R705 B.n330 B.n329 585
R706 B.n331 B.n312 585
R707 B.n333 B.n332 585
R708 B.n335 B.n311 585
R709 B.n338 B.n337 585
R710 B.n339 B.n310 585
R711 B.n341 B.n340 585
R712 B.n343 B.n309 585
R713 B.n346 B.n345 585
R714 B.n347 B.n308 585
R715 B.n349 B.n348 585
R716 B.n351 B.n307 585
R717 B.n354 B.n353 585
R718 B.n355 B.n306 585
R719 B.n357 B.n356 585
R720 B.n359 B.n305 585
R721 B.n362 B.n361 585
R722 B.n364 B.n302 585
R723 B.n366 B.n365 585
R724 B.n368 B.n301 585
R725 B.n371 B.n370 585
R726 B.n372 B.n300 585
R727 B.n374 B.n373 585
R728 B.n376 B.n299 585
R729 B.n379 B.n378 585
R730 B.n380 B.n296 585
R731 B.n383 B.n382 585
R732 B.n385 B.n295 585
R733 B.n388 B.n387 585
R734 B.n389 B.n294 585
R735 B.n391 B.n390 585
R736 B.n393 B.n293 585
R737 B.n396 B.n395 585
R738 B.n397 B.n292 585
R739 B.n399 B.n398 585
R740 B.n401 B.n291 585
R741 B.n404 B.n403 585
R742 B.n405 B.n290 585
R743 B.n407 B.n406 585
R744 B.n409 B.n289 585
R745 B.n412 B.n411 585
R746 B.n413 B.n288 585
R747 B.n415 B.n414 585
R748 B.n417 B.n287 585
R749 B.n420 B.n419 585
R750 B.n421 B.n286 585
R751 B.n423 B.n422 585
R752 B.n425 B.n285 585
R753 B.n428 B.n427 585
R754 B.n429 B.n284 585
R755 B.n434 B.n433 585
R756 B.n433 B.n432 585
R757 B.n435 B.n280 585
R758 B.n280 B.n279 585
R759 B.n437 B.n436 585
R760 B.n438 B.n437 585
R761 B.n274 B.n273 585
R762 B.n275 B.n274 585
R763 B.n446 B.n445 585
R764 B.n445 B.n444 585
R765 B.n447 B.n272 585
R766 B.n272 B.n271 585
R767 B.n449 B.n448 585
R768 B.n450 B.n449 585
R769 B.n266 B.n265 585
R770 B.n267 B.n266 585
R771 B.n458 B.n457 585
R772 B.n457 B.n456 585
R773 B.n459 B.n264 585
R774 B.n264 B.n263 585
R775 B.n461 B.n460 585
R776 B.n462 B.n461 585
R777 B.n258 B.n257 585
R778 B.n259 B.n258 585
R779 B.n470 B.n469 585
R780 B.n469 B.n468 585
R781 B.n471 B.n256 585
R782 B.n256 B.n254 585
R783 B.n473 B.n472 585
R784 B.n474 B.n473 585
R785 B.n250 B.n249 585
R786 B.n255 B.n250 585
R787 B.n482 B.n481 585
R788 B.n481 B.n480 585
R789 B.n483 B.n248 585
R790 B.n248 B.n247 585
R791 B.n485 B.n484 585
R792 B.n486 B.n485 585
R793 B.n242 B.n241 585
R794 B.n243 B.n242 585
R795 B.n494 B.n493 585
R796 B.n493 B.n492 585
R797 B.n495 B.n240 585
R798 B.n240 B.n239 585
R799 B.n497 B.n496 585
R800 B.n498 B.n497 585
R801 B.n234 B.n233 585
R802 B.n235 B.n234 585
R803 B.n506 B.n505 585
R804 B.n505 B.n504 585
R805 B.n507 B.n232 585
R806 B.n232 B.n231 585
R807 B.n509 B.n508 585
R808 B.n510 B.n509 585
R809 B.n226 B.n225 585
R810 B.n227 B.n226 585
R811 B.n518 B.n517 585
R812 B.n517 B.n516 585
R813 B.n519 B.n224 585
R814 B.n224 B.n223 585
R815 B.n521 B.n520 585
R816 B.n522 B.n521 585
R817 B.n218 B.n217 585
R818 B.n219 B.n218 585
R819 B.n531 B.n530 585
R820 B.n530 B.n529 585
R821 B.n532 B.n216 585
R822 B.n216 B.n215 585
R823 B.n534 B.n533 585
R824 B.n535 B.n534 585
R825 B.n3 B.n0 585
R826 B.n4 B.n3 585
R827 B.n661 B.n1 585
R828 B.n662 B.n661 585
R829 B.n660 B.n659 585
R830 B.n660 B.n8 585
R831 B.n658 B.n9 585
R832 B.n544 B.n9 585
R833 B.n657 B.n656 585
R834 B.n656 B.n655 585
R835 B.n11 B.n10 585
R836 B.n654 B.n11 585
R837 B.n652 B.n651 585
R838 B.n653 B.n652 585
R839 B.n650 B.n16 585
R840 B.n16 B.n15 585
R841 B.n649 B.n648 585
R842 B.n648 B.n647 585
R843 B.n18 B.n17 585
R844 B.n646 B.n18 585
R845 B.n644 B.n643 585
R846 B.n645 B.n644 585
R847 B.n642 B.n23 585
R848 B.n23 B.n22 585
R849 B.n641 B.n640 585
R850 B.n640 B.n639 585
R851 B.n25 B.n24 585
R852 B.n638 B.n25 585
R853 B.n636 B.n635 585
R854 B.n637 B.n636 585
R855 B.n634 B.n30 585
R856 B.n30 B.n29 585
R857 B.n633 B.n632 585
R858 B.n632 B.n631 585
R859 B.n32 B.n31 585
R860 B.n630 B.n32 585
R861 B.n628 B.n627 585
R862 B.n629 B.n628 585
R863 B.n626 B.n37 585
R864 B.n37 B.n36 585
R865 B.n625 B.n624 585
R866 B.n624 B.n623 585
R867 B.n39 B.n38 585
R868 B.n622 B.n39 585
R869 B.n620 B.n619 585
R870 B.n621 B.n620 585
R871 B.n618 B.n44 585
R872 B.n44 B.n43 585
R873 B.n617 B.n616 585
R874 B.n616 B.n615 585
R875 B.n46 B.n45 585
R876 B.n614 B.n46 585
R877 B.n612 B.n611 585
R878 B.n613 B.n612 585
R879 B.n610 B.n51 585
R880 B.n51 B.n50 585
R881 B.n609 B.n608 585
R882 B.n608 B.n607 585
R883 B.n53 B.n52 585
R884 B.n606 B.n53 585
R885 B.n604 B.n603 585
R886 B.n605 B.n604 585
R887 B.n602 B.n58 585
R888 B.n58 B.n57 585
R889 B.n601 B.n600 585
R890 B.n600 B.n599 585
R891 B.n60 B.n59 585
R892 B.n598 B.n60 585
R893 B.n596 B.n595 585
R894 B.n597 B.n596 585
R895 B.n594 B.n65 585
R896 B.n65 B.n64 585
R897 B.n593 B.n592 585
R898 B.n592 B.n591 585
R899 B.n665 B.n664 585
R900 B.n663 B.n2 585
R901 B.n592 B.n67 506.916
R902 B.n589 B.n68 506.916
R903 B.n431 B.n284 506.916
R904 B.n433 B.n282 506.916
R905 B.n100 B.t8 295.115
R906 B.n98 B.t16 295.115
R907 B.n297 B.t19 295.115
R908 B.n303 B.t12 295.115
R909 B.n590 B.n96 256.663
R910 B.n590 B.n95 256.663
R911 B.n590 B.n94 256.663
R912 B.n590 B.n93 256.663
R913 B.n590 B.n92 256.663
R914 B.n590 B.n91 256.663
R915 B.n590 B.n90 256.663
R916 B.n590 B.n89 256.663
R917 B.n590 B.n88 256.663
R918 B.n590 B.n87 256.663
R919 B.n590 B.n86 256.663
R920 B.n590 B.n85 256.663
R921 B.n590 B.n84 256.663
R922 B.n590 B.n83 256.663
R923 B.n590 B.n82 256.663
R924 B.n590 B.n81 256.663
R925 B.n590 B.n80 256.663
R926 B.n590 B.n79 256.663
R927 B.n590 B.n78 256.663
R928 B.n590 B.n77 256.663
R929 B.n590 B.n76 256.663
R930 B.n590 B.n75 256.663
R931 B.n590 B.n74 256.663
R932 B.n590 B.n73 256.663
R933 B.n590 B.n72 256.663
R934 B.n590 B.n71 256.663
R935 B.n590 B.n70 256.663
R936 B.n590 B.n69 256.663
R937 B.n317 B.n283 256.663
R938 B.n320 B.n283 256.663
R939 B.n326 B.n283 256.663
R940 B.n328 B.n283 256.663
R941 B.n334 B.n283 256.663
R942 B.n336 B.n283 256.663
R943 B.n342 B.n283 256.663
R944 B.n344 B.n283 256.663
R945 B.n350 B.n283 256.663
R946 B.n352 B.n283 256.663
R947 B.n358 B.n283 256.663
R948 B.n360 B.n283 256.663
R949 B.n367 B.n283 256.663
R950 B.n369 B.n283 256.663
R951 B.n375 B.n283 256.663
R952 B.n377 B.n283 256.663
R953 B.n384 B.n283 256.663
R954 B.n386 B.n283 256.663
R955 B.n392 B.n283 256.663
R956 B.n394 B.n283 256.663
R957 B.n400 B.n283 256.663
R958 B.n402 B.n283 256.663
R959 B.n408 B.n283 256.663
R960 B.n410 B.n283 256.663
R961 B.n416 B.n283 256.663
R962 B.n418 B.n283 256.663
R963 B.n424 B.n283 256.663
R964 B.n426 B.n283 256.663
R965 B.n667 B.n666 256.663
R966 B.n98 B.t17 215.06
R967 B.n297 B.t21 215.06
R968 B.n100 B.t10 215.06
R969 B.n303 B.t15 215.06
R970 B.n99 B.t18 177.63
R971 B.n298 B.t20 177.63
R972 B.n101 B.t11 177.629
R973 B.n304 B.t14 177.629
R974 B.n105 B.n104 163.367
R975 B.n109 B.n108 163.367
R976 B.n113 B.n112 163.367
R977 B.n117 B.n116 163.367
R978 B.n121 B.n120 163.367
R979 B.n125 B.n124 163.367
R980 B.n129 B.n128 163.367
R981 B.n133 B.n132 163.367
R982 B.n137 B.n136 163.367
R983 B.n141 B.n140 163.367
R984 B.n145 B.n144 163.367
R985 B.n149 B.n148 163.367
R986 B.n153 B.n152 163.367
R987 B.n157 B.n156 163.367
R988 B.n161 B.n160 163.367
R989 B.n165 B.n164 163.367
R990 B.n170 B.n169 163.367
R991 B.n174 B.n173 163.367
R992 B.n178 B.n177 163.367
R993 B.n182 B.n181 163.367
R994 B.n186 B.n185 163.367
R995 B.n190 B.n189 163.367
R996 B.n194 B.n193 163.367
R997 B.n198 B.n197 163.367
R998 B.n202 B.n201 163.367
R999 B.n206 B.n205 163.367
R1000 B.n210 B.n209 163.367
R1001 B.n589 B.n97 163.367
R1002 B.n431 B.n278 163.367
R1003 B.n439 B.n278 163.367
R1004 B.n439 B.n276 163.367
R1005 B.n443 B.n276 163.367
R1006 B.n443 B.n270 163.367
R1007 B.n451 B.n270 163.367
R1008 B.n451 B.n268 163.367
R1009 B.n455 B.n268 163.367
R1010 B.n455 B.n262 163.367
R1011 B.n463 B.n262 163.367
R1012 B.n463 B.n260 163.367
R1013 B.n467 B.n260 163.367
R1014 B.n467 B.n253 163.367
R1015 B.n475 B.n253 163.367
R1016 B.n475 B.n251 163.367
R1017 B.n479 B.n251 163.367
R1018 B.n479 B.n246 163.367
R1019 B.n487 B.n246 163.367
R1020 B.n487 B.n244 163.367
R1021 B.n491 B.n244 163.367
R1022 B.n491 B.n238 163.367
R1023 B.n499 B.n238 163.367
R1024 B.n499 B.n236 163.367
R1025 B.n503 B.n236 163.367
R1026 B.n503 B.n230 163.367
R1027 B.n511 B.n230 163.367
R1028 B.n511 B.n228 163.367
R1029 B.n515 B.n228 163.367
R1030 B.n515 B.n222 163.367
R1031 B.n523 B.n222 163.367
R1032 B.n523 B.n220 163.367
R1033 B.n528 B.n220 163.367
R1034 B.n528 B.n214 163.367
R1035 B.n536 B.n214 163.367
R1036 B.n537 B.n536 163.367
R1037 B.n537 B.n5 163.367
R1038 B.n6 B.n5 163.367
R1039 B.n7 B.n6 163.367
R1040 B.n543 B.n7 163.367
R1041 B.n545 B.n543 163.367
R1042 B.n545 B.n12 163.367
R1043 B.n13 B.n12 163.367
R1044 B.n14 B.n13 163.367
R1045 B.n550 B.n14 163.367
R1046 B.n550 B.n19 163.367
R1047 B.n20 B.n19 163.367
R1048 B.n21 B.n20 163.367
R1049 B.n555 B.n21 163.367
R1050 B.n555 B.n26 163.367
R1051 B.n27 B.n26 163.367
R1052 B.n28 B.n27 163.367
R1053 B.n560 B.n28 163.367
R1054 B.n560 B.n33 163.367
R1055 B.n34 B.n33 163.367
R1056 B.n35 B.n34 163.367
R1057 B.n565 B.n35 163.367
R1058 B.n565 B.n40 163.367
R1059 B.n41 B.n40 163.367
R1060 B.n42 B.n41 163.367
R1061 B.n570 B.n42 163.367
R1062 B.n570 B.n47 163.367
R1063 B.n48 B.n47 163.367
R1064 B.n49 B.n48 163.367
R1065 B.n575 B.n49 163.367
R1066 B.n575 B.n54 163.367
R1067 B.n55 B.n54 163.367
R1068 B.n56 B.n55 163.367
R1069 B.n580 B.n56 163.367
R1070 B.n580 B.n61 163.367
R1071 B.n62 B.n61 163.367
R1072 B.n63 B.n62 163.367
R1073 B.n585 B.n63 163.367
R1074 B.n585 B.n68 163.367
R1075 B.n319 B.n318 163.367
R1076 B.n321 B.n319 163.367
R1077 B.n325 B.n314 163.367
R1078 B.n329 B.n327 163.367
R1079 B.n333 B.n312 163.367
R1080 B.n337 B.n335 163.367
R1081 B.n341 B.n310 163.367
R1082 B.n345 B.n343 163.367
R1083 B.n349 B.n308 163.367
R1084 B.n353 B.n351 163.367
R1085 B.n357 B.n306 163.367
R1086 B.n361 B.n359 163.367
R1087 B.n366 B.n302 163.367
R1088 B.n370 B.n368 163.367
R1089 B.n374 B.n300 163.367
R1090 B.n378 B.n376 163.367
R1091 B.n383 B.n296 163.367
R1092 B.n387 B.n385 163.367
R1093 B.n391 B.n294 163.367
R1094 B.n395 B.n393 163.367
R1095 B.n399 B.n292 163.367
R1096 B.n403 B.n401 163.367
R1097 B.n407 B.n290 163.367
R1098 B.n411 B.n409 163.367
R1099 B.n415 B.n288 163.367
R1100 B.n419 B.n417 163.367
R1101 B.n423 B.n286 163.367
R1102 B.n427 B.n425 163.367
R1103 B.n433 B.n280 163.367
R1104 B.n437 B.n280 163.367
R1105 B.n437 B.n274 163.367
R1106 B.n445 B.n274 163.367
R1107 B.n445 B.n272 163.367
R1108 B.n449 B.n272 163.367
R1109 B.n449 B.n266 163.367
R1110 B.n457 B.n266 163.367
R1111 B.n457 B.n264 163.367
R1112 B.n461 B.n264 163.367
R1113 B.n461 B.n258 163.367
R1114 B.n469 B.n258 163.367
R1115 B.n469 B.n256 163.367
R1116 B.n473 B.n256 163.367
R1117 B.n473 B.n250 163.367
R1118 B.n481 B.n250 163.367
R1119 B.n481 B.n248 163.367
R1120 B.n485 B.n248 163.367
R1121 B.n485 B.n242 163.367
R1122 B.n493 B.n242 163.367
R1123 B.n493 B.n240 163.367
R1124 B.n497 B.n240 163.367
R1125 B.n497 B.n234 163.367
R1126 B.n505 B.n234 163.367
R1127 B.n505 B.n232 163.367
R1128 B.n509 B.n232 163.367
R1129 B.n509 B.n226 163.367
R1130 B.n517 B.n226 163.367
R1131 B.n517 B.n224 163.367
R1132 B.n521 B.n224 163.367
R1133 B.n521 B.n218 163.367
R1134 B.n530 B.n218 163.367
R1135 B.n530 B.n216 163.367
R1136 B.n534 B.n216 163.367
R1137 B.n534 B.n3 163.367
R1138 B.n665 B.n3 163.367
R1139 B.n661 B.n2 163.367
R1140 B.n661 B.n660 163.367
R1141 B.n660 B.n9 163.367
R1142 B.n656 B.n9 163.367
R1143 B.n656 B.n11 163.367
R1144 B.n652 B.n11 163.367
R1145 B.n652 B.n16 163.367
R1146 B.n648 B.n16 163.367
R1147 B.n648 B.n18 163.367
R1148 B.n644 B.n18 163.367
R1149 B.n644 B.n23 163.367
R1150 B.n640 B.n23 163.367
R1151 B.n640 B.n25 163.367
R1152 B.n636 B.n25 163.367
R1153 B.n636 B.n30 163.367
R1154 B.n632 B.n30 163.367
R1155 B.n632 B.n32 163.367
R1156 B.n628 B.n32 163.367
R1157 B.n628 B.n37 163.367
R1158 B.n624 B.n37 163.367
R1159 B.n624 B.n39 163.367
R1160 B.n620 B.n39 163.367
R1161 B.n620 B.n44 163.367
R1162 B.n616 B.n44 163.367
R1163 B.n616 B.n46 163.367
R1164 B.n612 B.n46 163.367
R1165 B.n612 B.n51 163.367
R1166 B.n608 B.n51 163.367
R1167 B.n608 B.n53 163.367
R1168 B.n604 B.n53 163.367
R1169 B.n604 B.n58 163.367
R1170 B.n600 B.n58 163.367
R1171 B.n600 B.n60 163.367
R1172 B.n596 B.n60 163.367
R1173 B.n596 B.n65 163.367
R1174 B.n592 B.n65 163.367
R1175 B.n432 B.n283 120.751
R1176 B.n591 B.n590 120.751
R1177 B.n69 B.n67 71.676
R1178 B.n105 B.n70 71.676
R1179 B.n109 B.n71 71.676
R1180 B.n113 B.n72 71.676
R1181 B.n117 B.n73 71.676
R1182 B.n121 B.n74 71.676
R1183 B.n125 B.n75 71.676
R1184 B.n129 B.n76 71.676
R1185 B.n133 B.n77 71.676
R1186 B.n137 B.n78 71.676
R1187 B.n141 B.n79 71.676
R1188 B.n145 B.n80 71.676
R1189 B.n149 B.n81 71.676
R1190 B.n153 B.n82 71.676
R1191 B.n157 B.n83 71.676
R1192 B.n161 B.n84 71.676
R1193 B.n165 B.n85 71.676
R1194 B.n170 B.n86 71.676
R1195 B.n174 B.n87 71.676
R1196 B.n178 B.n88 71.676
R1197 B.n182 B.n89 71.676
R1198 B.n186 B.n90 71.676
R1199 B.n190 B.n91 71.676
R1200 B.n194 B.n92 71.676
R1201 B.n198 B.n93 71.676
R1202 B.n202 B.n94 71.676
R1203 B.n206 B.n95 71.676
R1204 B.n210 B.n96 71.676
R1205 B.n97 B.n96 71.676
R1206 B.n209 B.n95 71.676
R1207 B.n205 B.n94 71.676
R1208 B.n201 B.n93 71.676
R1209 B.n197 B.n92 71.676
R1210 B.n193 B.n91 71.676
R1211 B.n189 B.n90 71.676
R1212 B.n185 B.n89 71.676
R1213 B.n181 B.n88 71.676
R1214 B.n177 B.n87 71.676
R1215 B.n173 B.n86 71.676
R1216 B.n169 B.n85 71.676
R1217 B.n164 B.n84 71.676
R1218 B.n160 B.n83 71.676
R1219 B.n156 B.n82 71.676
R1220 B.n152 B.n81 71.676
R1221 B.n148 B.n80 71.676
R1222 B.n144 B.n79 71.676
R1223 B.n140 B.n78 71.676
R1224 B.n136 B.n77 71.676
R1225 B.n132 B.n76 71.676
R1226 B.n128 B.n75 71.676
R1227 B.n124 B.n74 71.676
R1228 B.n120 B.n73 71.676
R1229 B.n116 B.n72 71.676
R1230 B.n112 B.n71 71.676
R1231 B.n108 B.n70 71.676
R1232 B.n104 B.n69 71.676
R1233 B.n317 B.n282 71.676
R1234 B.n321 B.n320 71.676
R1235 B.n326 B.n325 71.676
R1236 B.n329 B.n328 71.676
R1237 B.n334 B.n333 71.676
R1238 B.n337 B.n336 71.676
R1239 B.n342 B.n341 71.676
R1240 B.n345 B.n344 71.676
R1241 B.n350 B.n349 71.676
R1242 B.n353 B.n352 71.676
R1243 B.n358 B.n357 71.676
R1244 B.n361 B.n360 71.676
R1245 B.n367 B.n366 71.676
R1246 B.n370 B.n369 71.676
R1247 B.n375 B.n374 71.676
R1248 B.n378 B.n377 71.676
R1249 B.n384 B.n383 71.676
R1250 B.n387 B.n386 71.676
R1251 B.n392 B.n391 71.676
R1252 B.n395 B.n394 71.676
R1253 B.n400 B.n399 71.676
R1254 B.n403 B.n402 71.676
R1255 B.n408 B.n407 71.676
R1256 B.n411 B.n410 71.676
R1257 B.n416 B.n415 71.676
R1258 B.n419 B.n418 71.676
R1259 B.n424 B.n423 71.676
R1260 B.n427 B.n426 71.676
R1261 B.n318 B.n317 71.676
R1262 B.n320 B.n314 71.676
R1263 B.n327 B.n326 71.676
R1264 B.n328 B.n312 71.676
R1265 B.n335 B.n334 71.676
R1266 B.n336 B.n310 71.676
R1267 B.n343 B.n342 71.676
R1268 B.n344 B.n308 71.676
R1269 B.n351 B.n350 71.676
R1270 B.n352 B.n306 71.676
R1271 B.n359 B.n358 71.676
R1272 B.n360 B.n302 71.676
R1273 B.n368 B.n367 71.676
R1274 B.n369 B.n300 71.676
R1275 B.n376 B.n375 71.676
R1276 B.n377 B.n296 71.676
R1277 B.n385 B.n384 71.676
R1278 B.n386 B.n294 71.676
R1279 B.n393 B.n392 71.676
R1280 B.n394 B.n292 71.676
R1281 B.n401 B.n400 71.676
R1282 B.n402 B.n290 71.676
R1283 B.n409 B.n408 71.676
R1284 B.n410 B.n288 71.676
R1285 B.n417 B.n416 71.676
R1286 B.n418 B.n286 71.676
R1287 B.n425 B.n424 71.676
R1288 B.n426 B.n284 71.676
R1289 B.n666 B.n665 71.676
R1290 B.n666 B.n2 71.676
R1291 B.n432 B.n279 66.7564
R1292 B.n438 B.n279 66.7564
R1293 B.n438 B.n275 66.7564
R1294 B.n444 B.n275 66.7564
R1295 B.n444 B.n271 66.7564
R1296 B.n450 B.n271 66.7564
R1297 B.n456 B.n267 66.7564
R1298 B.n456 B.n263 66.7564
R1299 B.n462 B.n263 66.7564
R1300 B.n462 B.n259 66.7564
R1301 B.n468 B.n259 66.7564
R1302 B.n468 B.n254 66.7564
R1303 B.n474 B.n254 66.7564
R1304 B.n474 B.n255 66.7564
R1305 B.n480 B.n247 66.7564
R1306 B.n486 B.n247 66.7564
R1307 B.n486 B.n243 66.7564
R1308 B.n492 B.n243 66.7564
R1309 B.n498 B.n239 66.7564
R1310 B.n498 B.n235 66.7564
R1311 B.n504 B.n235 66.7564
R1312 B.n504 B.n231 66.7564
R1313 B.n510 B.n231 66.7564
R1314 B.n516 B.n227 66.7564
R1315 B.n516 B.n223 66.7564
R1316 B.n522 B.n223 66.7564
R1317 B.n522 B.n219 66.7564
R1318 B.n529 B.n219 66.7564
R1319 B.n535 B.n215 66.7564
R1320 B.n535 B.n4 66.7564
R1321 B.n664 B.n4 66.7564
R1322 B.n664 B.n663 66.7564
R1323 B.n663 B.n662 66.7564
R1324 B.n662 B.n8 66.7564
R1325 B.n544 B.n8 66.7564
R1326 B.n655 B.n654 66.7564
R1327 B.n654 B.n653 66.7564
R1328 B.n653 B.n15 66.7564
R1329 B.n647 B.n15 66.7564
R1330 B.n647 B.n646 66.7564
R1331 B.n645 B.n22 66.7564
R1332 B.n639 B.n22 66.7564
R1333 B.n639 B.n638 66.7564
R1334 B.n638 B.n637 66.7564
R1335 B.n637 B.n29 66.7564
R1336 B.n631 B.n630 66.7564
R1337 B.n630 B.n629 66.7564
R1338 B.n629 B.n36 66.7564
R1339 B.n623 B.n36 66.7564
R1340 B.n622 B.n621 66.7564
R1341 B.n621 B.n43 66.7564
R1342 B.n615 B.n43 66.7564
R1343 B.n615 B.n614 66.7564
R1344 B.n614 B.n613 66.7564
R1345 B.n613 B.n50 66.7564
R1346 B.n607 B.n50 66.7564
R1347 B.n607 B.n606 66.7564
R1348 B.n605 B.n57 66.7564
R1349 B.n599 B.n57 66.7564
R1350 B.n599 B.n598 66.7564
R1351 B.n598 B.n597 66.7564
R1352 B.n597 B.n64 66.7564
R1353 B.n591 B.n64 66.7564
R1354 B.n480 B.t1 64.793
R1355 B.n623 B.t3 64.793
R1356 B.t4 B.n215 62.8296
R1357 B.n544 B.t2 62.8296
R1358 B.n102 B.n101 59.5399
R1359 B.n167 B.n99 59.5399
R1360 B.n381 B.n298 59.5399
R1361 B.n363 B.n304 59.5399
R1362 B.t13 B.n267 56.9394
R1363 B.n606 B.t9 56.9394
R1364 B.n492 B.t5 47.1223
R1365 B.n631 B.t0 47.1223
R1366 B.t7 B.n227 41.2321
R1367 B.n646 B.t6 41.2321
R1368 B.n101 B.n100 37.4308
R1369 B.n99 B.n98 37.4308
R1370 B.n298 B.n297 37.4308
R1371 B.n304 B.n303 37.4308
R1372 B.n434 B.n281 32.9371
R1373 B.n430 B.n429 32.9371
R1374 B.n588 B.n587 32.9371
R1375 B.n593 B.n66 32.9371
R1376 B.n510 B.t7 25.5248
R1377 B.t6 B.n645 25.5248
R1378 B.t5 B.n239 19.6346
R1379 B.t0 B.n29 19.6346
R1380 B B.n667 18.0485
R1381 B.n435 B.n434 10.6151
R1382 B.n436 B.n435 10.6151
R1383 B.n436 B.n273 10.6151
R1384 B.n446 B.n273 10.6151
R1385 B.n447 B.n446 10.6151
R1386 B.n448 B.n447 10.6151
R1387 B.n448 B.n265 10.6151
R1388 B.n458 B.n265 10.6151
R1389 B.n459 B.n458 10.6151
R1390 B.n460 B.n459 10.6151
R1391 B.n460 B.n257 10.6151
R1392 B.n470 B.n257 10.6151
R1393 B.n471 B.n470 10.6151
R1394 B.n472 B.n471 10.6151
R1395 B.n472 B.n249 10.6151
R1396 B.n482 B.n249 10.6151
R1397 B.n483 B.n482 10.6151
R1398 B.n484 B.n483 10.6151
R1399 B.n484 B.n241 10.6151
R1400 B.n494 B.n241 10.6151
R1401 B.n495 B.n494 10.6151
R1402 B.n496 B.n495 10.6151
R1403 B.n496 B.n233 10.6151
R1404 B.n506 B.n233 10.6151
R1405 B.n507 B.n506 10.6151
R1406 B.n508 B.n507 10.6151
R1407 B.n508 B.n225 10.6151
R1408 B.n518 B.n225 10.6151
R1409 B.n519 B.n518 10.6151
R1410 B.n520 B.n519 10.6151
R1411 B.n520 B.n217 10.6151
R1412 B.n531 B.n217 10.6151
R1413 B.n532 B.n531 10.6151
R1414 B.n533 B.n532 10.6151
R1415 B.n533 B.n0 10.6151
R1416 B.n316 B.n281 10.6151
R1417 B.n316 B.n315 10.6151
R1418 B.n322 B.n315 10.6151
R1419 B.n323 B.n322 10.6151
R1420 B.n324 B.n323 10.6151
R1421 B.n324 B.n313 10.6151
R1422 B.n330 B.n313 10.6151
R1423 B.n331 B.n330 10.6151
R1424 B.n332 B.n331 10.6151
R1425 B.n332 B.n311 10.6151
R1426 B.n338 B.n311 10.6151
R1427 B.n339 B.n338 10.6151
R1428 B.n340 B.n339 10.6151
R1429 B.n340 B.n309 10.6151
R1430 B.n346 B.n309 10.6151
R1431 B.n347 B.n346 10.6151
R1432 B.n348 B.n347 10.6151
R1433 B.n348 B.n307 10.6151
R1434 B.n354 B.n307 10.6151
R1435 B.n355 B.n354 10.6151
R1436 B.n356 B.n355 10.6151
R1437 B.n356 B.n305 10.6151
R1438 B.n362 B.n305 10.6151
R1439 B.n365 B.n364 10.6151
R1440 B.n365 B.n301 10.6151
R1441 B.n371 B.n301 10.6151
R1442 B.n372 B.n371 10.6151
R1443 B.n373 B.n372 10.6151
R1444 B.n373 B.n299 10.6151
R1445 B.n379 B.n299 10.6151
R1446 B.n380 B.n379 10.6151
R1447 B.n382 B.n295 10.6151
R1448 B.n388 B.n295 10.6151
R1449 B.n389 B.n388 10.6151
R1450 B.n390 B.n389 10.6151
R1451 B.n390 B.n293 10.6151
R1452 B.n396 B.n293 10.6151
R1453 B.n397 B.n396 10.6151
R1454 B.n398 B.n397 10.6151
R1455 B.n398 B.n291 10.6151
R1456 B.n404 B.n291 10.6151
R1457 B.n405 B.n404 10.6151
R1458 B.n406 B.n405 10.6151
R1459 B.n406 B.n289 10.6151
R1460 B.n412 B.n289 10.6151
R1461 B.n413 B.n412 10.6151
R1462 B.n414 B.n413 10.6151
R1463 B.n414 B.n287 10.6151
R1464 B.n420 B.n287 10.6151
R1465 B.n421 B.n420 10.6151
R1466 B.n422 B.n421 10.6151
R1467 B.n422 B.n285 10.6151
R1468 B.n428 B.n285 10.6151
R1469 B.n429 B.n428 10.6151
R1470 B.n430 B.n277 10.6151
R1471 B.n440 B.n277 10.6151
R1472 B.n441 B.n440 10.6151
R1473 B.n442 B.n441 10.6151
R1474 B.n442 B.n269 10.6151
R1475 B.n452 B.n269 10.6151
R1476 B.n453 B.n452 10.6151
R1477 B.n454 B.n453 10.6151
R1478 B.n454 B.n261 10.6151
R1479 B.n464 B.n261 10.6151
R1480 B.n465 B.n464 10.6151
R1481 B.n466 B.n465 10.6151
R1482 B.n466 B.n252 10.6151
R1483 B.n476 B.n252 10.6151
R1484 B.n477 B.n476 10.6151
R1485 B.n478 B.n477 10.6151
R1486 B.n478 B.n245 10.6151
R1487 B.n488 B.n245 10.6151
R1488 B.n489 B.n488 10.6151
R1489 B.n490 B.n489 10.6151
R1490 B.n490 B.n237 10.6151
R1491 B.n500 B.n237 10.6151
R1492 B.n501 B.n500 10.6151
R1493 B.n502 B.n501 10.6151
R1494 B.n502 B.n229 10.6151
R1495 B.n512 B.n229 10.6151
R1496 B.n513 B.n512 10.6151
R1497 B.n514 B.n513 10.6151
R1498 B.n514 B.n221 10.6151
R1499 B.n524 B.n221 10.6151
R1500 B.n525 B.n524 10.6151
R1501 B.n527 B.n525 10.6151
R1502 B.n527 B.n526 10.6151
R1503 B.n526 B.n213 10.6151
R1504 B.n538 B.n213 10.6151
R1505 B.n539 B.n538 10.6151
R1506 B.n540 B.n539 10.6151
R1507 B.n541 B.n540 10.6151
R1508 B.n542 B.n541 10.6151
R1509 B.n546 B.n542 10.6151
R1510 B.n547 B.n546 10.6151
R1511 B.n548 B.n547 10.6151
R1512 B.n549 B.n548 10.6151
R1513 B.n551 B.n549 10.6151
R1514 B.n552 B.n551 10.6151
R1515 B.n553 B.n552 10.6151
R1516 B.n554 B.n553 10.6151
R1517 B.n556 B.n554 10.6151
R1518 B.n557 B.n556 10.6151
R1519 B.n558 B.n557 10.6151
R1520 B.n559 B.n558 10.6151
R1521 B.n561 B.n559 10.6151
R1522 B.n562 B.n561 10.6151
R1523 B.n563 B.n562 10.6151
R1524 B.n564 B.n563 10.6151
R1525 B.n566 B.n564 10.6151
R1526 B.n567 B.n566 10.6151
R1527 B.n568 B.n567 10.6151
R1528 B.n569 B.n568 10.6151
R1529 B.n571 B.n569 10.6151
R1530 B.n572 B.n571 10.6151
R1531 B.n573 B.n572 10.6151
R1532 B.n574 B.n573 10.6151
R1533 B.n576 B.n574 10.6151
R1534 B.n577 B.n576 10.6151
R1535 B.n578 B.n577 10.6151
R1536 B.n579 B.n578 10.6151
R1537 B.n581 B.n579 10.6151
R1538 B.n582 B.n581 10.6151
R1539 B.n583 B.n582 10.6151
R1540 B.n584 B.n583 10.6151
R1541 B.n586 B.n584 10.6151
R1542 B.n587 B.n586 10.6151
R1543 B.n659 B.n1 10.6151
R1544 B.n659 B.n658 10.6151
R1545 B.n658 B.n657 10.6151
R1546 B.n657 B.n10 10.6151
R1547 B.n651 B.n10 10.6151
R1548 B.n651 B.n650 10.6151
R1549 B.n650 B.n649 10.6151
R1550 B.n649 B.n17 10.6151
R1551 B.n643 B.n17 10.6151
R1552 B.n643 B.n642 10.6151
R1553 B.n642 B.n641 10.6151
R1554 B.n641 B.n24 10.6151
R1555 B.n635 B.n24 10.6151
R1556 B.n635 B.n634 10.6151
R1557 B.n634 B.n633 10.6151
R1558 B.n633 B.n31 10.6151
R1559 B.n627 B.n31 10.6151
R1560 B.n627 B.n626 10.6151
R1561 B.n626 B.n625 10.6151
R1562 B.n625 B.n38 10.6151
R1563 B.n619 B.n38 10.6151
R1564 B.n619 B.n618 10.6151
R1565 B.n618 B.n617 10.6151
R1566 B.n617 B.n45 10.6151
R1567 B.n611 B.n45 10.6151
R1568 B.n611 B.n610 10.6151
R1569 B.n610 B.n609 10.6151
R1570 B.n609 B.n52 10.6151
R1571 B.n603 B.n52 10.6151
R1572 B.n603 B.n602 10.6151
R1573 B.n602 B.n601 10.6151
R1574 B.n601 B.n59 10.6151
R1575 B.n595 B.n59 10.6151
R1576 B.n595 B.n594 10.6151
R1577 B.n594 B.n593 10.6151
R1578 B.n103 B.n66 10.6151
R1579 B.n106 B.n103 10.6151
R1580 B.n107 B.n106 10.6151
R1581 B.n110 B.n107 10.6151
R1582 B.n111 B.n110 10.6151
R1583 B.n114 B.n111 10.6151
R1584 B.n115 B.n114 10.6151
R1585 B.n118 B.n115 10.6151
R1586 B.n119 B.n118 10.6151
R1587 B.n122 B.n119 10.6151
R1588 B.n123 B.n122 10.6151
R1589 B.n126 B.n123 10.6151
R1590 B.n127 B.n126 10.6151
R1591 B.n130 B.n127 10.6151
R1592 B.n131 B.n130 10.6151
R1593 B.n134 B.n131 10.6151
R1594 B.n135 B.n134 10.6151
R1595 B.n138 B.n135 10.6151
R1596 B.n139 B.n138 10.6151
R1597 B.n142 B.n139 10.6151
R1598 B.n143 B.n142 10.6151
R1599 B.n146 B.n143 10.6151
R1600 B.n147 B.n146 10.6151
R1601 B.n151 B.n150 10.6151
R1602 B.n154 B.n151 10.6151
R1603 B.n155 B.n154 10.6151
R1604 B.n158 B.n155 10.6151
R1605 B.n159 B.n158 10.6151
R1606 B.n162 B.n159 10.6151
R1607 B.n163 B.n162 10.6151
R1608 B.n166 B.n163 10.6151
R1609 B.n171 B.n168 10.6151
R1610 B.n172 B.n171 10.6151
R1611 B.n175 B.n172 10.6151
R1612 B.n176 B.n175 10.6151
R1613 B.n179 B.n176 10.6151
R1614 B.n180 B.n179 10.6151
R1615 B.n183 B.n180 10.6151
R1616 B.n184 B.n183 10.6151
R1617 B.n187 B.n184 10.6151
R1618 B.n188 B.n187 10.6151
R1619 B.n191 B.n188 10.6151
R1620 B.n192 B.n191 10.6151
R1621 B.n195 B.n192 10.6151
R1622 B.n196 B.n195 10.6151
R1623 B.n199 B.n196 10.6151
R1624 B.n200 B.n199 10.6151
R1625 B.n203 B.n200 10.6151
R1626 B.n204 B.n203 10.6151
R1627 B.n207 B.n204 10.6151
R1628 B.n208 B.n207 10.6151
R1629 B.n211 B.n208 10.6151
R1630 B.n212 B.n211 10.6151
R1631 B.n588 B.n212 10.6151
R1632 B.n450 B.t13 9.81755
R1633 B.t9 B.n605 9.81755
R1634 B.n667 B.n0 8.11757
R1635 B.n667 B.n1 8.11757
R1636 B.n364 B.n363 6.5566
R1637 B.n381 B.n380 6.5566
R1638 B.n150 B.n102 6.5566
R1639 B.n167 B.n166 6.5566
R1640 B.n363 B.n362 4.05904
R1641 B.n382 B.n381 4.05904
R1642 B.n147 B.n102 4.05904
R1643 B.n168 B.n167 4.05904
R1644 B.n529 B.t4 3.92732
R1645 B.n655 B.t2 3.92732
R1646 B.n255 B.t1 1.96391
R1647 B.t3 B.n622 1.96391
R1648 VP.n28 VP.n27 178.673
R1649 VP.n50 VP.n49 178.673
R1650 VP.n26 VP.n25 178.673
R1651 VP.n13 VP.n12 161.3
R1652 VP.n14 VP.n9 161.3
R1653 VP.n16 VP.n15 161.3
R1654 VP.n17 VP.n8 161.3
R1655 VP.n20 VP.n19 161.3
R1656 VP.n21 VP.n7 161.3
R1657 VP.n23 VP.n22 161.3
R1658 VP.n24 VP.n6 161.3
R1659 VP.n48 VP.n0 161.3
R1660 VP.n47 VP.n46 161.3
R1661 VP.n45 VP.n1 161.3
R1662 VP.n44 VP.n43 161.3
R1663 VP.n41 VP.n2 161.3
R1664 VP.n40 VP.n39 161.3
R1665 VP.n38 VP.n3 161.3
R1666 VP.n37 VP.n36 161.3
R1667 VP.n34 VP.n4 161.3
R1668 VP.n33 VP.n32 161.3
R1669 VP.n31 VP.n5 161.3
R1670 VP.n30 VP.n29 161.3
R1671 VP.n10 VP.t0 121.507
R1672 VP.n28 VP.t5 89.3211
R1673 VP.n35 VP.t7 89.3211
R1674 VP.n42 VP.t6 89.3211
R1675 VP.n49 VP.t2 89.3211
R1676 VP.n25 VP.t1 89.3211
R1677 VP.n18 VP.t4 89.3211
R1678 VP.n11 VP.t3 89.3211
R1679 VP.n47 VP.n1 56.5193
R1680 VP.n33 VP.n5 56.5193
R1681 VP.n40 VP.n3 56.5193
R1682 VP.n23 VP.n7 56.5193
R1683 VP.n16 VP.n9 56.5193
R1684 VP.n11 VP.n10 55.5644
R1685 VP.n27 VP.n26 41.5232
R1686 VP.n29 VP.n5 24.4675
R1687 VP.n34 VP.n33 24.4675
R1688 VP.n36 VP.n3 24.4675
R1689 VP.n41 VP.n40 24.4675
R1690 VP.n43 VP.n1 24.4675
R1691 VP.n48 VP.n47 24.4675
R1692 VP.n24 VP.n23 24.4675
R1693 VP.n17 VP.n16 24.4675
R1694 VP.n19 VP.n7 24.4675
R1695 VP.n12 VP.n9 24.4675
R1696 VP.n13 VP.n10 18.0716
R1697 VP.n35 VP.n34 13.9467
R1698 VP.n43 VP.n42 13.9467
R1699 VP.n19 VP.n18 13.9467
R1700 VP.n36 VP.n35 10.5213
R1701 VP.n42 VP.n41 10.5213
R1702 VP.n18 VP.n17 10.5213
R1703 VP.n12 VP.n11 10.5213
R1704 VP.n29 VP.n28 7.09593
R1705 VP.n49 VP.n48 7.09593
R1706 VP.n25 VP.n24 7.09593
R1707 VP.n14 VP.n13 0.189894
R1708 VP.n15 VP.n14 0.189894
R1709 VP.n15 VP.n8 0.189894
R1710 VP.n20 VP.n8 0.189894
R1711 VP.n21 VP.n20 0.189894
R1712 VP.n22 VP.n21 0.189894
R1713 VP.n22 VP.n6 0.189894
R1714 VP.n26 VP.n6 0.189894
R1715 VP.n30 VP.n27 0.189894
R1716 VP.n31 VP.n30 0.189894
R1717 VP.n32 VP.n31 0.189894
R1718 VP.n32 VP.n4 0.189894
R1719 VP.n37 VP.n4 0.189894
R1720 VP.n38 VP.n37 0.189894
R1721 VP.n39 VP.n38 0.189894
R1722 VP.n39 VP.n2 0.189894
R1723 VP.n44 VP.n2 0.189894
R1724 VP.n45 VP.n44 0.189894
R1725 VP.n46 VP.n45 0.189894
R1726 VP.n46 VP.n0 0.189894
R1727 VP.n50 VP.n0 0.189894
R1728 VP VP.n50 0.0516364
R1729 VDD1 VDD1.n0 66.7233
R1730 VDD1.n3 VDD1.n2 66.6096
R1731 VDD1.n3 VDD1.n1 66.6096
R1732 VDD1.n5 VDD1.n4 65.8331
R1733 VDD1.n5 VDD1.n3 36.8974
R1734 VDD1.n4 VDD1.t3 3.33945
R1735 VDD1.n4 VDD1.t6 3.33945
R1736 VDD1.n0 VDD1.t7 3.33945
R1737 VDD1.n0 VDD1.t4 3.33945
R1738 VDD1.n2 VDD1.t1 3.33945
R1739 VDD1.n2 VDD1.t5 3.33945
R1740 VDD1.n1 VDD1.t2 3.33945
R1741 VDD1.n1 VDD1.t0 3.33945
R1742 VDD1 VDD1.n5 0.774207
C0 VN VDD2 4.02374f
C1 VP VDD1 4.28619f
C2 VTAIL VDD1 5.65737f
C3 VTAIL VP 4.4747f
C4 VDD1 VDD2 1.26037f
C5 VP VDD2 0.413332f
C6 VTAIL VDD2 5.70508f
C7 VDD1 VN 0.149992f
C8 VP VN 5.31562f
C9 VTAIL VN 4.46059f
C10 VDD2 B 3.909242f
C11 VDD1 B 4.246265f
C12 VTAIL B 5.926992f
C13 VN B 11.061761f
C14 VP B 9.610196f
C15 VDD1.t7 B 0.117943f
C16 VDD1.t4 B 0.117943f
C17 VDD1.n0 B 0.987351f
C18 VDD1.t2 B 0.117943f
C19 VDD1.t0 B 0.117943f
C20 VDD1.n1 B 0.986539f
C21 VDD1.t1 B 0.117943f
C22 VDD1.t5 B 0.117943f
C23 VDD1.n2 B 0.986539f
C24 VDD1.n3 B 2.39245f
C25 VDD1.t3 B 0.117943f
C26 VDD1.t6 B 0.117943f
C27 VDD1.n4 B 0.98172f
C28 VDD1.n5 B 2.17073f
C29 VP.n0 B 0.032774f
C30 VP.t2 B 0.82248f
C31 VP.n1 B 0.041452f
C32 VP.n2 B 0.032774f
C33 VP.t6 B 0.82248f
C34 VP.n3 B 0.047845f
C35 VP.n4 B 0.032774f
C36 VP.t7 B 0.82248f
C37 VP.n5 B 0.054238f
C38 VP.n6 B 0.032774f
C39 VP.t1 B 0.82248f
C40 VP.n7 B 0.041452f
C41 VP.n8 B 0.032774f
C42 VP.t4 B 0.82248f
C43 VP.n9 B 0.047845f
C44 VP.t0 B 0.942704f
C45 VP.n10 B 0.394054f
C46 VP.t3 B 0.82248f
C47 VP.n11 B 0.382467f
C48 VP.n12 B 0.043892f
C49 VP.n13 B 0.208401f
C50 VP.n14 B 0.032774f
C51 VP.n15 B 0.032774f
C52 VP.n16 B 0.047845f
C53 VP.n17 B 0.043892f
C54 VP.n18 B 0.320643f
C55 VP.n19 B 0.048114f
C56 VP.n20 B 0.032774f
C57 VP.n21 B 0.032774f
C58 VP.n22 B 0.032774f
C59 VP.n23 B 0.054238f
C60 VP.n24 B 0.03967f
C61 VP.n25 B 0.389126f
C62 VP.n26 B 1.33461f
C63 VP.n27 B 1.36298f
C64 VP.t5 B 0.82248f
C65 VP.n28 B 0.389126f
C66 VP.n29 B 0.03967f
C67 VP.n30 B 0.032774f
C68 VP.n31 B 0.032774f
C69 VP.n32 B 0.032774f
C70 VP.n33 B 0.041452f
C71 VP.n34 B 0.048114f
C72 VP.n35 B 0.320643f
C73 VP.n36 B 0.043892f
C74 VP.n37 B 0.032774f
C75 VP.n38 B 0.032774f
C76 VP.n39 B 0.032774f
C77 VP.n40 B 0.047845f
C78 VP.n41 B 0.043892f
C79 VP.n42 B 0.320643f
C80 VP.n43 B 0.048114f
C81 VP.n44 B 0.032774f
C82 VP.n45 B 0.032774f
C83 VP.n46 B 0.032774f
C84 VP.n47 B 0.054238f
C85 VP.n48 B 0.03967f
C86 VP.n49 B 0.389126f
C87 VP.n50 B 0.032774f
C88 VTAIL.t8 B 0.103625f
C89 VTAIL.t6 B 0.103625f
C90 VTAIL.n0 B 0.80298f
C91 VTAIL.n1 B 0.331934f
C92 VTAIL.n2 B 0.030038f
C93 VTAIL.n3 B 0.022113f
C94 VTAIL.n4 B 0.011883f
C95 VTAIL.n5 B 0.028087f
C96 VTAIL.n6 B 0.012582f
C97 VTAIL.n7 B 0.022113f
C98 VTAIL.n8 B 0.011883f
C99 VTAIL.n9 B 0.028087f
C100 VTAIL.n10 B 0.012582f
C101 VTAIL.n11 B 0.0942f
C102 VTAIL.t2 B 0.045752f
C103 VTAIL.n12 B 0.021065f
C104 VTAIL.n13 B 0.01659f
C105 VTAIL.n14 B 0.011883f
C106 VTAIL.n15 B 0.519133f
C107 VTAIL.n16 B 0.022113f
C108 VTAIL.n17 B 0.011883f
C109 VTAIL.n18 B 0.012582f
C110 VTAIL.n19 B 0.028087f
C111 VTAIL.n20 B 0.028087f
C112 VTAIL.n21 B 0.012582f
C113 VTAIL.n22 B 0.011883f
C114 VTAIL.n23 B 0.022113f
C115 VTAIL.n24 B 0.022113f
C116 VTAIL.n25 B 0.011883f
C117 VTAIL.n26 B 0.012582f
C118 VTAIL.n27 B 0.028087f
C119 VTAIL.n28 B 0.058956f
C120 VTAIL.n29 B 0.012582f
C121 VTAIL.n30 B 0.011883f
C122 VTAIL.n31 B 0.048999f
C123 VTAIL.n32 B 0.032732f
C124 VTAIL.n33 B 0.169724f
C125 VTAIL.n34 B 0.030038f
C126 VTAIL.n35 B 0.022113f
C127 VTAIL.n36 B 0.011883f
C128 VTAIL.n37 B 0.028087f
C129 VTAIL.n38 B 0.012582f
C130 VTAIL.n39 B 0.022113f
C131 VTAIL.n40 B 0.011883f
C132 VTAIL.n41 B 0.028087f
C133 VTAIL.n42 B 0.012582f
C134 VTAIL.n43 B 0.0942f
C135 VTAIL.t12 B 0.045752f
C136 VTAIL.n44 B 0.021065f
C137 VTAIL.n45 B 0.01659f
C138 VTAIL.n46 B 0.011883f
C139 VTAIL.n47 B 0.519133f
C140 VTAIL.n48 B 0.022113f
C141 VTAIL.n49 B 0.011883f
C142 VTAIL.n50 B 0.012582f
C143 VTAIL.n51 B 0.028087f
C144 VTAIL.n52 B 0.028087f
C145 VTAIL.n53 B 0.012582f
C146 VTAIL.n54 B 0.011883f
C147 VTAIL.n55 B 0.022113f
C148 VTAIL.n56 B 0.022113f
C149 VTAIL.n57 B 0.011883f
C150 VTAIL.n58 B 0.012582f
C151 VTAIL.n59 B 0.028087f
C152 VTAIL.n60 B 0.058956f
C153 VTAIL.n61 B 0.012582f
C154 VTAIL.n62 B 0.011883f
C155 VTAIL.n63 B 0.048999f
C156 VTAIL.n64 B 0.032732f
C157 VTAIL.n65 B 0.169724f
C158 VTAIL.t10 B 0.103625f
C159 VTAIL.t11 B 0.103625f
C160 VTAIL.n66 B 0.80298f
C161 VTAIL.n67 B 0.44634f
C162 VTAIL.n68 B 0.030038f
C163 VTAIL.n69 B 0.022113f
C164 VTAIL.n70 B 0.011883f
C165 VTAIL.n71 B 0.028087f
C166 VTAIL.n72 B 0.012582f
C167 VTAIL.n73 B 0.022113f
C168 VTAIL.n74 B 0.011883f
C169 VTAIL.n75 B 0.028087f
C170 VTAIL.n76 B 0.012582f
C171 VTAIL.n77 B 0.0942f
C172 VTAIL.t1 B 0.045752f
C173 VTAIL.n78 B 0.021065f
C174 VTAIL.n79 B 0.01659f
C175 VTAIL.n80 B 0.011883f
C176 VTAIL.n81 B 0.519133f
C177 VTAIL.n82 B 0.022113f
C178 VTAIL.n83 B 0.011883f
C179 VTAIL.n84 B 0.012582f
C180 VTAIL.n85 B 0.028087f
C181 VTAIL.n86 B 0.028087f
C182 VTAIL.n87 B 0.012582f
C183 VTAIL.n88 B 0.011883f
C184 VTAIL.n89 B 0.022113f
C185 VTAIL.n90 B 0.022113f
C186 VTAIL.n91 B 0.011883f
C187 VTAIL.n92 B 0.012582f
C188 VTAIL.n93 B 0.028087f
C189 VTAIL.n94 B 0.058956f
C190 VTAIL.n95 B 0.012582f
C191 VTAIL.n96 B 0.011883f
C192 VTAIL.n97 B 0.048999f
C193 VTAIL.n98 B 0.032732f
C194 VTAIL.n99 B 0.919439f
C195 VTAIL.n100 B 0.030038f
C196 VTAIL.n101 B 0.022113f
C197 VTAIL.n102 B 0.011883f
C198 VTAIL.n103 B 0.028087f
C199 VTAIL.n104 B 0.012582f
C200 VTAIL.n105 B 0.022113f
C201 VTAIL.n106 B 0.011883f
C202 VTAIL.n107 B 0.028087f
C203 VTAIL.n108 B 0.012582f
C204 VTAIL.n109 B 0.0942f
C205 VTAIL.t3 B 0.045752f
C206 VTAIL.n110 B 0.021065f
C207 VTAIL.n111 B 0.01659f
C208 VTAIL.n112 B 0.011883f
C209 VTAIL.n113 B 0.519133f
C210 VTAIL.n114 B 0.022113f
C211 VTAIL.n115 B 0.011883f
C212 VTAIL.n116 B 0.012582f
C213 VTAIL.n117 B 0.028087f
C214 VTAIL.n118 B 0.028087f
C215 VTAIL.n119 B 0.012582f
C216 VTAIL.n120 B 0.011883f
C217 VTAIL.n121 B 0.022113f
C218 VTAIL.n122 B 0.022113f
C219 VTAIL.n123 B 0.011883f
C220 VTAIL.n124 B 0.012582f
C221 VTAIL.n125 B 0.028087f
C222 VTAIL.n126 B 0.058956f
C223 VTAIL.n127 B 0.012582f
C224 VTAIL.n128 B 0.011883f
C225 VTAIL.n129 B 0.048999f
C226 VTAIL.n130 B 0.032732f
C227 VTAIL.n131 B 0.919439f
C228 VTAIL.t7 B 0.103625f
C229 VTAIL.t9 B 0.103625f
C230 VTAIL.n132 B 0.802986f
C231 VTAIL.n133 B 0.446335f
C232 VTAIL.n134 B 0.030038f
C233 VTAIL.n135 B 0.022113f
C234 VTAIL.n136 B 0.011883f
C235 VTAIL.n137 B 0.028087f
C236 VTAIL.n138 B 0.012582f
C237 VTAIL.n139 B 0.022113f
C238 VTAIL.n140 B 0.011883f
C239 VTAIL.n141 B 0.028087f
C240 VTAIL.n142 B 0.012582f
C241 VTAIL.n143 B 0.0942f
C242 VTAIL.t5 B 0.045752f
C243 VTAIL.n144 B 0.021065f
C244 VTAIL.n145 B 0.01659f
C245 VTAIL.n146 B 0.011883f
C246 VTAIL.n147 B 0.519133f
C247 VTAIL.n148 B 0.022113f
C248 VTAIL.n149 B 0.011883f
C249 VTAIL.n150 B 0.012582f
C250 VTAIL.n151 B 0.028087f
C251 VTAIL.n152 B 0.028087f
C252 VTAIL.n153 B 0.012582f
C253 VTAIL.n154 B 0.011883f
C254 VTAIL.n155 B 0.022113f
C255 VTAIL.n156 B 0.022113f
C256 VTAIL.n157 B 0.011883f
C257 VTAIL.n158 B 0.012582f
C258 VTAIL.n159 B 0.028087f
C259 VTAIL.n160 B 0.058956f
C260 VTAIL.n161 B 0.012582f
C261 VTAIL.n162 B 0.011883f
C262 VTAIL.n163 B 0.048999f
C263 VTAIL.n164 B 0.032732f
C264 VTAIL.n165 B 0.169724f
C265 VTAIL.n166 B 0.030038f
C266 VTAIL.n167 B 0.022113f
C267 VTAIL.n168 B 0.011883f
C268 VTAIL.n169 B 0.028087f
C269 VTAIL.n170 B 0.012582f
C270 VTAIL.n171 B 0.022113f
C271 VTAIL.n172 B 0.011883f
C272 VTAIL.n173 B 0.028087f
C273 VTAIL.n174 B 0.012582f
C274 VTAIL.n175 B 0.0942f
C275 VTAIL.t15 B 0.045752f
C276 VTAIL.n176 B 0.021065f
C277 VTAIL.n177 B 0.01659f
C278 VTAIL.n178 B 0.011883f
C279 VTAIL.n179 B 0.519133f
C280 VTAIL.n180 B 0.022113f
C281 VTAIL.n181 B 0.011883f
C282 VTAIL.n182 B 0.012582f
C283 VTAIL.n183 B 0.028087f
C284 VTAIL.n184 B 0.028087f
C285 VTAIL.n185 B 0.012582f
C286 VTAIL.n186 B 0.011883f
C287 VTAIL.n187 B 0.022113f
C288 VTAIL.n188 B 0.022113f
C289 VTAIL.n189 B 0.011883f
C290 VTAIL.n190 B 0.012582f
C291 VTAIL.n191 B 0.028087f
C292 VTAIL.n192 B 0.058956f
C293 VTAIL.n193 B 0.012582f
C294 VTAIL.n194 B 0.011883f
C295 VTAIL.n195 B 0.048999f
C296 VTAIL.n196 B 0.032732f
C297 VTAIL.n197 B 0.169724f
C298 VTAIL.t13 B 0.103625f
C299 VTAIL.t0 B 0.103625f
C300 VTAIL.n198 B 0.802986f
C301 VTAIL.n199 B 0.446335f
C302 VTAIL.n200 B 0.030038f
C303 VTAIL.n201 B 0.022113f
C304 VTAIL.n202 B 0.011883f
C305 VTAIL.n203 B 0.028087f
C306 VTAIL.n204 B 0.012582f
C307 VTAIL.n205 B 0.022113f
C308 VTAIL.n206 B 0.011883f
C309 VTAIL.n207 B 0.028087f
C310 VTAIL.n208 B 0.012582f
C311 VTAIL.n209 B 0.0942f
C312 VTAIL.t14 B 0.045752f
C313 VTAIL.n210 B 0.021065f
C314 VTAIL.n211 B 0.01659f
C315 VTAIL.n212 B 0.011883f
C316 VTAIL.n213 B 0.519133f
C317 VTAIL.n214 B 0.022113f
C318 VTAIL.n215 B 0.011883f
C319 VTAIL.n216 B 0.012582f
C320 VTAIL.n217 B 0.028087f
C321 VTAIL.n218 B 0.028087f
C322 VTAIL.n219 B 0.012582f
C323 VTAIL.n220 B 0.011883f
C324 VTAIL.n221 B 0.022113f
C325 VTAIL.n222 B 0.022113f
C326 VTAIL.n223 B 0.011883f
C327 VTAIL.n224 B 0.012582f
C328 VTAIL.n225 B 0.028087f
C329 VTAIL.n226 B 0.058956f
C330 VTAIL.n227 B 0.012582f
C331 VTAIL.n228 B 0.011883f
C332 VTAIL.n229 B 0.048999f
C333 VTAIL.n230 B 0.032732f
C334 VTAIL.n231 B 0.919438f
C335 VTAIL.n232 B 0.030038f
C336 VTAIL.n233 B 0.022113f
C337 VTAIL.n234 B 0.011883f
C338 VTAIL.n235 B 0.028087f
C339 VTAIL.n236 B 0.012582f
C340 VTAIL.n237 B 0.022113f
C341 VTAIL.n238 B 0.011883f
C342 VTAIL.n239 B 0.028087f
C343 VTAIL.n240 B 0.012582f
C344 VTAIL.n241 B 0.0942f
C345 VTAIL.t4 B 0.045752f
C346 VTAIL.n242 B 0.021065f
C347 VTAIL.n243 B 0.01659f
C348 VTAIL.n244 B 0.011883f
C349 VTAIL.n245 B 0.519133f
C350 VTAIL.n246 B 0.022113f
C351 VTAIL.n247 B 0.011883f
C352 VTAIL.n248 B 0.012582f
C353 VTAIL.n249 B 0.028087f
C354 VTAIL.n250 B 0.028087f
C355 VTAIL.n251 B 0.012582f
C356 VTAIL.n252 B 0.011883f
C357 VTAIL.n253 B 0.022113f
C358 VTAIL.n254 B 0.022113f
C359 VTAIL.n255 B 0.011883f
C360 VTAIL.n256 B 0.012582f
C361 VTAIL.n257 B 0.028087f
C362 VTAIL.n258 B 0.058956f
C363 VTAIL.n259 B 0.012582f
C364 VTAIL.n260 B 0.011883f
C365 VTAIL.n261 B 0.048999f
C366 VTAIL.n262 B 0.032732f
C367 VTAIL.n263 B 0.915292f
C368 VDD2.t3 B 0.115478f
C369 VDD2.t0 B 0.115478f
C370 VDD2.n0 B 0.965922f
C371 VDD2.t6 B 0.115478f
C372 VDD2.t7 B 0.115478f
C373 VDD2.n1 B 0.965922f
C374 VDD2.n2 B 2.29032f
C375 VDD2.t2 B 0.115478f
C376 VDD2.t1 B 0.115478f
C377 VDD2.n3 B 0.961208f
C378 VDD2.n4 B 2.09572f
C379 VDD2.t5 B 0.115478f
C380 VDD2.t4 B 0.115478f
C381 VDD2.n5 B 0.965894f
C382 VN.n0 B 0.031973f
C383 VN.t5 B 0.802359f
C384 VN.n1 B 0.040438f
C385 VN.n2 B 0.031973f
C386 VN.t3 B 0.802359f
C387 VN.n3 B 0.046674f
C388 VN.t7 B 0.919642f
C389 VN.n4 B 0.384414f
C390 VN.t1 B 0.802359f
C391 VN.n5 B 0.37311f
C392 VN.n6 B 0.042818f
C393 VN.n7 B 0.203302f
C394 VN.n8 B 0.031973f
C395 VN.n9 B 0.031973f
C396 VN.n10 B 0.046674f
C397 VN.n11 B 0.042818f
C398 VN.n12 B 0.312799f
C399 VN.n13 B 0.046937f
C400 VN.n14 B 0.031973f
C401 VN.n15 B 0.031973f
C402 VN.n16 B 0.031973f
C403 VN.n17 B 0.052911f
C404 VN.n18 B 0.0387f
C405 VN.n19 B 0.379607f
C406 VN.n20 B 0.031973f
C407 VN.n21 B 0.031973f
C408 VN.t6 B 0.802359f
C409 VN.n22 B 0.040438f
C410 VN.n23 B 0.031973f
C411 VN.t2 B 0.802359f
C412 VN.n24 B 0.046674f
C413 VN.t4 B 0.919642f
C414 VN.n25 B 0.384414f
C415 VN.t0 B 0.802359f
C416 VN.n26 B 0.37311f
C417 VN.n27 B 0.042818f
C418 VN.n28 B 0.203302f
C419 VN.n29 B 0.031973f
C420 VN.n30 B 0.031973f
C421 VN.n31 B 0.046674f
C422 VN.n32 B 0.042818f
C423 VN.n33 B 0.312799f
C424 VN.n34 B 0.046937f
C425 VN.n35 B 0.031973f
C426 VN.n36 B 0.031973f
C427 VN.n37 B 0.031973f
C428 VN.n38 B 0.052911f
C429 VN.n39 B 0.0387f
C430 VN.n40 B 0.379607f
C431 VN.n41 B 1.32296f
.ends

