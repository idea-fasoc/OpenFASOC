* NGSPICE file created from diff_pair_sample_0917.ext - technology: sky130A

.subckt diff_pair_sample_0917 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VN.t0 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=2.53275 ps=15.68 w=15.35 l=3.95
X1 VTAIL.t1 VP.t0 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=2.53275 ps=15.68 w=15.35 l=3.95
X2 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=5.9865 pd=31.48 as=0 ps=0 w=15.35 l=3.95
X3 VTAIL.t13 VN.t1 VDD2.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=5.9865 pd=31.48 as=2.53275 ps=15.68 w=15.35 l=3.95
X4 VDD2.t5 VN.t2 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=5.9865 ps=31.48 w=15.35 l=3.95
X5 VDD1.t6 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=2.53275 ps=15.68 w=15.35 l=3.95
X6 VDD1.t5 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=5.9865 ps=31.48 w=15.35 l=3.95
X7 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.9865 pd=31.48 as=0 ps=0 w=15.35 l=3.95
X8 VTAIL.t6 VP.t3 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=5.9865 pd=31.48 as=2.53275 ps=15.68 w=15.35 l=3.95
X9 VTAIL.t4 VP.t4 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=5.9865 pd=31.48 as=2.53275 ps=15.68 w=15.35 l=3.95
X10 B.t13 B.t11 B.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=5.9865 pd=31.48 as=0 ps=0 w=15.35 l=3.95
X11 VTAIL.t11 VN.t3 VDD2.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=5.9865 pd=31.48 as=2.53275 ps=15.68 w=15.35 l=3.95
X12 VDD2.t0 VN.t4 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=5.9865 ps=31.48 w=15.35 l=3.95
X13 VDD1.t2 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=5.9865 ps=31.48 w=15.35 l=3.95
X14 VDD1.t1 VP.t6 VTAIL.t15 B.t21 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=2.53275 ps=15.68 w=15.35 l=3.95
X15 VDD2.t3 VN.t5 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=2.53275 ps=15.68 w=15.35 l=3.95
X16 VDD2.t2 VN.t6 VTAIL.t8 B.t21 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=2.53275 ps=15.68 w=15.35 l=3.95
X17 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=5.9865 pd=31.48 as=0 ps=0 w=15.35 l=3.95
X18 VTAIL.t7 VN.t7 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=2.53275 ps=15.68 w=15.35 l=3.95
X19 VTAIL.t2 VP.t7 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=2.53275 pd=15.68 as=2.53275 ps=15.68 w=15.35 l=3.95
R0 VN.n75 VN.n39 161.3
R1 VN.n74 VN.n73 161.3
R2 VN.n72 VN.n40 161.3
R3 VN.n71 VN.n70 161.3
R4 VN.n69 VN.n41 161.3
R5 VN.n68 VN.n67 161.3
R6 VN.n66 VN.n42 161.3
R7 VN.n65 VN.n64 161.3
R8 VN.n62 VN.n43 161.3
R9 VN.n61 VN.n60 161.3
R10 VN.n59 VN.n44 161.3
R11 VN.n58 VN.n57 161.3
R12 VN.n56 VN.n45 161.3
R13 VN.n55 VN.n54 161.3
R14 VN.n53 VN.n46 161.3
R15 VN.n52 VN.n51 161.3
R16 VN.n50 VN.n47 161.3
R17 VN.n36 VN.n0 161.3
R18 VN.n35 VN.n34 161.3
R19 VN.n33 VN.n1 161.3
R20 VN.n32 VN.n31 161.3
R21 VN.n30 VN.n2 161.3
R22 VN.n29 VN.n28 161.3
R23 VN.n27 VN.n3 161.3
R24 VN.n26 VN.n25 161.3
R25 VN.n23 VN.n4 161.3
R26 VN.n22 VN.n21 161.3
R27 VN.n20 VN.n5 161.3
R28 VN.n19 VN.n18 161.3
R29 VN.n17 VN.n6 161.3
R30 VN.n16 VN.n15 161.3
R31 VN.n14 VN.n7 161.3
R32 VN.n13 VN.n12 161.3
R33 VN.n11 VN.n8 161.3
R34 VN.n9 VN.t3 125.903
R35 VN.n48 VN.t4 125.903
R36 VN.n10 VN.t6 93.6549
R37 VN.n24 VN.t7 93.6549
R38 VN.n37 VN.t2 93.6549
R39 VN.n49 VN.t0 93.6549
R40 VN.n63 VN.t5 93.6549
R41 VN.n76 VN.t1 93.6549
R42 VN.n10 VN.n9 68.2271
R43 VN.n49 VN.n48 68.2271
R44 VN.n38 VN.n37 61.6295
R45 VN.n77 VN.n76 61.6295
R46 VN VN.n77 60.0269
R47 VN.n31 VN.n30 56.5193
R48 VN.n70 VN.n69 56.5193
R49 VN.n17 VN.n16 40.4934
R50 VN.n18 VN.n17 40.4934
R51 VN.n56 VN.n55 40.4934
R52 VN.n57 VN.n56 40.4934
R53 VN.n12 VN.n11 24.4675
R54 VN.n12 VN.n7 24.4675
R55 VN.n16 VN.n7 24.4675
R56 VN.n18 VN.n5 24.4675
R57 VN.n22 VN.n5 24.4675
R58 VN.n23 VN.n22 24.4675
R59 VN.n25 VN.n3 24.4675
R60 VN.n29 VN.n3 24.4675
R61 VN.n30 VN.n29 24.4675
R62 VN.n31 VN.n1 24.4675
R63 VN.n35 VN.n1 24.4675
R64 VN.n36 VN.n35 24.4675
R65 VN.n55 VN.n46 24.4675
R66 VN.n51 VN.n46 24.4675
R67 VN.n51 VN.n50 24.4675
R68 VN.n69 VN.n68 24.4675
R69 VN.n68 VN.n42 24.4675
R70 VN.n64 VN.n42 24.4675
R71 VN.n62 VN.n61 24.4675
R72 VN.n61 VN.n44 24.4675
R73 VN.n57 VN.n44 24.4675
R74 VN.n75 VN.n74 24.4675
R75 VN.n74 VN.n40 24.4675
R76 VN.n70 VN.n40 24.4675
R77 VN.n37 VN.n36 20.5528
R78 VN.n76 VN.n75 20.5528
R79 VN.n25 VN.n24 17.6167
R80 VN.n64 VN.n63 17.6167
R81 VN.n11 VN.n10 6.85126
R82 VN.n24 VN.n23 6.85126
R83 VN.n50 VN.n49 6.85126
R84 VN.n63 VN.n62 6.85126
R85 VN.n48 VN.n47 2.67497
R86 VN.n9 VN.n8 2.67497
R87 VN.n77 VN.n39 0.417535
R88 VN.n38 VN.n0 0.417535
R89 VN VN.n38 0.394291
R90 VN.n73 VN.n39 0.189894
R91 VN.n73 VN.n72 0.189894
R92 VN.n72 VN.n71 0.189894
R93 VN.n71 VN.n41 0.189894
R94 VN.n67 VN.n41 0.189894
R95 VN.n67 VN.n66 0.189894
R96 VN.n66 VN.n65 0.189894
R97 VN.n65 VN.n43 0.189894
R98 VN.n60 VN.n43 0.189894
R99 VN.n60 VN.n59 0.189894
R100 VN.n59 VN.n58 0.189894
R101 VN.n58 VN.n45 0.189894
R102 VN.n54 VN.n45 0.189894
R103 VN.n54 VN.n53 0.189894
R104 VN.n53 VN.n52 0.189894
R105 VN.n52 VN.n47 0.189894
R106 VN.n13 VN.n8 0.189894
R107 VN.n14 VN.n13 0.189894
R108 VN.n15 VN.n14 0.189894
R109 VN.n15 VN.n6 0.189894
R110 VN.n19 VN.n6 0.189894
R111 VN.n20 VN.n19 0.189894
R112 VN.n21 VN.n20 0.189894
R113 VN.n21 VN.n4 0.189894
R114 VN.n26 VN.n4 0.189894
R115 VN.n27 VN.n26 0.189894
R116 VN.n28 VN.n27 0.189894
R117 VN.n28 VN.n2 0.189894
R118 VN.n32 VN.n2 0.189894
R119 VN.n33 VN.n32 0.189894
R120 VN.n34 VN.n33 0.189894
R121 VN.n34 VN.n0 0.189894
R122 VDD2.n2 VDD2.n1 62.4379
R123 VDD2.n2 VDD2.n0 62.4379
R124 VDD2 VDD2.n5 62.4351
R125 VDD2.n4 VDD2.n3 60.6486
R126 VDD2.n4 VDD2.n2 53.5515
R127 VDD2 VDD2.n4 1.90352
R128 VDD2.n5 VDD2.t7 1.2904
R129 VDD2.n5 VDD2.t0 1.2904
R130 VDD2.n3 VDD2.t6 1.2904
R131 VDD2.n3 VDD2.t3 1.2904
R132 VDD2.n1 VDD2.t4 1.2904
R133 VDD2.n1 VDD2.t5 1.2904
R134 VDD2.n0 VDD2.t1 1.2904
R135 VDD2.n0 VDD2.t2 1.2904
R136 VTAIL.n690 VTAIL.n610 289.615
R137 VTAIL.n82 VTAIL.n2 289.615
R138 VTAIL.n168 VTAIL.n88 289.615
R139 VTAIL.n256 VTAIL.n176 289.615
R140 VTAIL.n604 VTAIL.n524 289.615
R141 VTAIL.n516 VTAIL.n436 289.615
R142 VTAIL.n430 VTAIL.n350 289.615
R143 VTAIL.n342 VTAIL.n262 289.615
R144 VTAIL.n639 VTAIL.n638 185
R145 VTAIL.n641 VTAIL.n640 185
R146 VTAIL.n634 VTAIL.n633 185
R147 VTAIL.n647 VTAIL.n646 185
R148 VTAIL.n649 VTAIL.n648 185
R149 VTAIL.n630 VTAIL.n629 185
R150 VTAIL.n655 VTAIL.n654 185
R151 VTAIL.n657 VTAIL.n656 185
R152 VTAIL.n626 VTAIL.n625 185
R153 VTAIL.n663 VTAIL.n662 185
R154 VTAIL.n665 VTAIL.n664 185
R155 VTAIL.n622 VTAIL.n621 185
R156 VTAIL.n671 VTAIL.n670 185
R157 VTAIL.n673 VTAIL.n672 185
R158 VTAIL.n618 VTAIL.n617 185
R159 VTAIL.n680 VTAIL.n679 185
R160 VTAIL.n681 VTAIL.n616 185
R161 VTAIL.n683 VTAIL.n682 185
R162 VTAIL.n614 VTAIL.n613 185
R163 VTAIL.n689 VTAIL.n688 185
R164 VTAIL.n691 VTAIL.n690 185
R165 VTAIL.n31 VTAIL.n30 185
R166 VTAIL.n33 VTAIL.n32 185
R167 VTAIL.n26 VTAIL.n25 185
R168 VTAIL.n39 VTAIL.n38 185
R169 VTAIL.n41 VTAIL.n40 185
R170 VTAIL.n22 VTAIL.n21 185
R171 VTAIL.n47 VTAIL.n46 185
R172 VTAIL.n49 VTAIL.n48 185
R173 VTAIL.n18 VTAIL.n17 185
R174 VTAIL.n55 VTAIL.n54 185
R175 VTAIL.n57 VTAIL.n56 185
R176 VTAIL.n14 VTAIL.n13 185
R177 VTAIL.n63 VTAIL.n62 185
R178 VTAIL.n65 VTAIL.n64 185
R179 VTAIL.n10 VTAIL.n9 185
R180 VTAIL.n72 VTAIL.n71 185
R181 VTAIL.n73 VTAIL.n8 185
R182 VTAIL.n75 VTAIL.n74 185
R183 VTAIL.n6 VTAIL.n5 185
R184 VTAIL.n81 VTAIL.n80 185
R185 VTAIL.n83 VTAIL.n82 185
R186 VTAIL.n117 VTAIL.n116 185
R187 VTAIL.n119 VTAIL.n118 185
R188 VTAIL.n112 VTAIL.n111 185
R189 VTAIL.n125 VTAIL.n124 185
R190 VTAIL.n127 VTAIL.n126 185
R191 VTAIL.n108 VTAIL.n107 185
R192 VTAIL.n133 VTAIL.n132 185
R193 VTAIL.n135 VTAIL.n134 185
R194 VTAIL.n104 VTAIL.n103 185
R195 VTAIL.n141 VTAIL.n140 185
R196 VTAIL.n143 VTAIL.n142 185
R197 VTAIL.n100 VTAIL.n99 185
R198 VTAIL.n149 VTAIL.n148 185
R199 VTAIL.n151 VTAIL.n150 185
R200 VTAIL.n96 VTAIL.n95 185
R201 VTAIL.n158 VTAIL.n157 185
R202 VTAIL.n159 VTAIL.n94 185
R203 VTAIL.n161 VTAIL.n160 185
R204 VTAIL.n92 VTAIL.n91 185
R205 VTAIL.n167 VTAIL.n166 185
R206 VTAIL.n169 VTAIL.n168 185
R207 VTAIL.n205 VTAIL.n204 185
R208 VTAIL.n207 VTAIL.n206 185
R209 VTAIL.n200 VTAIL.n199 185
R210 VTAIL.n213 VTAIL.n212 185
R211 VTAIL.n215 VTAIL.n214 185
R212 VTAIL.n196 VTAIL.n195 185
R213 VTAIL.n221 VTAIL.n220 185
R214 VTAIL.n223 VTAIL.n222 185
R215 VTAIL.n192 VTAIL.n191 185
R216 VTAIL.n229 VTAIL.n228 185
R217 VTAIL.n231 VTAIL.n230 185
R218 VTAIL.n188 VTAIL.n187 185
R219 VTAIL.n237 VTAIL.n236 185
R220 VTAIL.n239 VTAIL.n238 185
R221 VTAIL.n184 VTAIL.n183 185
R222 VTAIL.n246 VTAIL.n245 185
R223 VTAIL.n247 VTAIL.n182 185
R224 VTAIL.n249 VTAIL.n248 185
R225 VTAIL.n180 VTAIL.n179 185
R226 VTAIL.n255 VTAIL.n254 185
R227 VTAIL.n257 VTAIL.n256 185
R228 VTAIL.n605 VTAIL.n604 185
R229 VTAIL.n603 VTAIL.n602 185
R230 VTAIL.n528 VTAIL.n527 185
R231 VTAIL.n532 VTAIL.n530 185
R232 VTAIL.n597 VTAIL.n596 185
R233 VTAIL.n595 VTAIL.n594 185
R234 VTAIL.n534 VTAIL.n533 185
R235 VTAIL.n589 VTAIL.n588 185
R236 VTAIL.n587 VTAIL.n586 185
R237 VTAIL.n538 VTAIL.n537 185
R238 VTAIL.n581 VTAIL.n580 185
R239 VTAIL.n579 VTAIL.n578 185
R240 VTAIL.n542 VTAIL.n541 185
R241 VTAIL.n573 VTAIL.n572 185
R242 VTAIL.n571 VTAIL.n570 185
R243 VTAIL.n546 VTAIL.n545 185
R244 VTAIL.n565 VTAIL.n564 185
R245 VTAIL.n563 VTAIL.n562 185
R246 VTAIL.n550 VTAIL.n549 185
R247 VTAIL.n557 VTAIL.n556 185
R248 VTAIL.n555 VTAIL.n554 185
R249 VTAIL.n517 VTAIL.n516 185
R250 VTAIL.n515 VTAIL.n514 185
R251 VTAIL.n440 VTAIL.n439 185
R252 VTAIL.n444 VTAIL.n442 185
R253 VTAIL.n509 VTAIL.n508 185
R254 VTAIL.n507 VTAIL.n506 185
R255 VTAIL.n446 VTAIL.n445 185
R256 VTAIL.n501 VTAIL.n500 185
R257 VTAIL.n499 VTAIL.n498 185
R258 VTAIL.n450 VTAIL.n449 185
R259 VTAIL.n493 VTAIL.n492 185
R260 VTAIL.n491 VTAIL.n490 185
R261 VTAIL.n454 VTAIL.n453 185
R262 VTAIL.n485 VTAIL.n484 185
R263 VTAIL.n483 VTAIL.n482 185
R264 VTAIL.n458 VTAIL.n457 185
R265 VTAIL.n477 VTAIL.n476 185
R266 VTAIL.n475 VTAIL.n474 185
R267 VTAIL.n462 VTAIL.n461 185
R268 VTAIL.n469 VTAIL.n468 185
R269 VTAIL.n467 VTAIL.n466 185
R270 VTAIL.n431 VTAIL.n430 185
R271 VTAIL.n429 VTAIL.n428 185
R272 VTAIL.n354 VTAIL.n353 185
R273 VTAIL.n358 VTAIL.n356 185
R274 VTAIL.n423 VTAIL.n422 185
R275 VTAIL.n421 VTAIL.n420 185
R276 VTAIL.n360 VTAIL.n359 185
R277 VTAIL.n415 VTAIL.n414 185
R278 VTAIL.n413 VTAIL.n412 185
R279 VTAIL.n364 VTAIL.n363 185
R280 VTAIL.n407 VTAIL.n406 185
R281 VTAIL.n405 VTAIL.n404 185
R282 VTAIL.n368 VTAIL.n367 185
R283 VTAIL.n399 VTAIL.n398 185
R284 VTAIL.n397 VTAIL.n396 185
R285 VTAIL.n372 VTAIL.n371 185
R286 VTAIL.n391 VTAIL.n390 185
R287 VTAIL.n389 VTAIL.n388 185
R288 VTAIL.n376 VTAIL.n375 185
R289 VTAIL.n383 VTAIL.n382 185
R290 VTAIL.n381 VTAIL.n380 185
R291 VTAIL.n343 VTAIL.n342 185
R292 VTAIL.n341 VTAIL.n340 185
R293 VTAIL.n266 VTAIL.n265 185
R294 VTAIL.n270 VTAIL.n268 185
R295 VTAIL.n335 VTAIL.n334 185
R296 VTAIL.n333 VTAIL.n332 185
R297 VTAIL.n272 VTAIL.n271 185
R298 VTAIL.n327 VTAIL.n326 185
R299 VTAIL.n325 VTAIL.n324 185
R300 VTAIL.n276 VTAIL.n275 185
R301 VTAIL.n319 VTAIL.n318 185
R302 VTAIL.n317 VTAIL.n316 185
R303 VTAIL.n280 VTAIL.n279 185
R304 VTAIL.n311 VTAIL.n310 185
R305 VTAIL.n309 VTAIL.n308 185
R306 VTAIL.n284 VTAIL.n283 185
R307 VTAIL.n303 VTAIL.n302 185
R308 VTAIL.n301 VTAIL.n300 185
R309 VTAIL.n288 VTAIL.n287 185
R310 VTAIL.n295 VTAIL.n294 185
R311 VTAIL.n293 VTAIL.n292 185
R312 VTAIL.n637 VTAIL.t12 147.659
R313 VTAIL.n29 VTAIL.t11 147.659
R314 VTAIL.n115 VTAIL.t3 147.659
R315 VTAIL.n203 VTAIL.t6 147.659
R316 VTAIL.n553 VTAIL.t0 147.659
R317 VTAIL.n465 VTAIL.t4 147.659
R318 VTAIL.n379 VTAIL.t10 147.659
R319 VTAIL.n291 VTAIL.t13 147.659
R320 VTAIL.n640 VTAIL.n639 104.615
R321 VTAIL.n640 VTAIL.n633 104.615
R322 VTAIL.n647 VTAIL.n633 104.615
R323 VTAIL.n648 VTAIL.n647 104.615
R324 VTAIL.n648 VTAIL.n629 104.615
R325 VTAIL.n655 VTAIL.n629 104.615
R326 VTAIL.n656 VTAIL.n655 104.615
R327 VTAIL.n656 VTAIL.n625 104.615
R328 VTAIL.n663 VTAIL.n625 104.615
R329 VTAIL.n664 VTAIL.n663 104.615
R330 VTAIL.n664 VTAIL.n621 104.615
R331 VTAIL.n671 VTAIL.n621 104.615
R332 VTAIL.n672 VTAIL.n671 104.615
R333 VTAIL.n672 VTAIL.n617 104.615
R334 VTAIL.n680 VTAIL.n617 104.615
R335 VTAIL.n681 VTAIL.n680 104.615
R336 VTAIL.n682 VTAIL.n681 104.615
R337 VTAIL.n682 VTAIL.n613 104.615
R338 VTAIL.n689 VTAIL.n613 104.615
R339 VTAIL.n690 VTAIL.n689 104.615
R340 VTAIL.n32 VTAIL.n31 104.615
R341 VTAIL.n32 VTAIL.n25 104.615
R342 VTAIL.n39 VTAIL.n25 104.615
R343 VTAIL.n40 VTAIL.n39 104.615
R344 VTAIL.n40 VTAIL.n21 104.615
R345 VTAIL.n47 VTAIL.n21 104.615
R346 VTAIL.n48 VTAIL.n47 104.615
R347 VTAIL.n48 VTAIL.n17 104.615
R348 VTAIL.n55 VTAIL.n17 104.615
R349 VTAIL.n56 VTAIL.n55 104.615
R350 VTAIL.n56 VTAIL.n13 104.615
R351 VTAIL.n63 VTAIL.n13 104.615
R352 VTAIL.n64 VTAIL.n63 104.615
R353 VTAIL.n64 VTAIL.n9 104.615
R354 VTAIL.n72 VTAIL.n9 104.615
R355 VTAIL.n73 VTAIL.n72 104.615
R356 VTAIL.n74 VTAIL.n73 104.615
R357 VTAIL.n74 VTAIL.n5 104.615
R358 VTAIL.n81 VTAIL.n5 104.615
R359 VTAIL.n82 VTAIL.n81 104.615
R360 VTAIL.n118 VTAIL.n117 104.615
R361 VTAIL.n118 VTAIL.n111 104.615
R362 VTAIL.n125 VTAIL.n111 104.615
R363 VTAIL.n126 VTAIL.n125 104.615
R364 VTAIL.n126 VTAIL.n107 104.615
R365 VTAIL.n133 VTAIL.n107 104.615
R366 VTAIL.n134 VTAIL.n133 104.615
R367 VTAIL.n134 VTAIL.n103 104.615
R368 VTAIL.n141 VTAIL.n103 104.615
R369 VTAIL.n142 VTAIL.n141 104.615
R370 VTAIL.n142 VTAIL.n99 104.615
R371 VTAIL.n149 VTAIL.n99 104.615
R372 VTAIL.n150 VTAIL.n149 104.615
R373 VTAIL.n150 VTAIL.n95 104.615
R374 VTAIL.n158 VTAIL.n95 104.615
R375 VTAIL.n159 VTAIL.n158 104.615
R376 VTAIL.n160 VTAIL.n159 104.615
R377 VTAIL.n160 VTAIL.n91 104.615
R378 VTAIL.n167 VTAIL.n91 104.615
R379 VTAIL.n168 VTAIL.n167 104.615
R380 VTAIL.n206 VTAIL.n205 104.615
R381 VTAIL.n206 VTAIL.n199 104.615
R382 VTAIL.n213 VTAIL.n199 104.615
R383 VTAIL.n214 VTAIL.n213 104.615
R384 VTAIL.n214 VTAIL.n195 104.615
R385 VTAIL.n221 VTAIL.n195 104.615
R386 VTAIL.n222 VTAIL.n221 104.615
R387 VTAIL.n222 VTAIL.n191 104.615
R388 VTAIL.n229 VTAIL.n191 104.615
R389 VTAIL.n230 VTAIL.n229 104.615
R390 VTAIL.n230 VTAIL.n187 104.615
R391 VTAIL.n237 VTAIL.n187 104.615
R392 VTAIL.n238 VTAIL.n237 104.615
R393 VTAIL.n238 VTAIL.n183 104.615
R394 VTAIL.n246 VTAIL.n183 104.615
R395 VTAIL.n247 VTAIL.n246 104.615
R396 VTAIL.n248 VTAIL.n247 104.615
R397 VTAIL.n248 VTAIL.n179 104.615
R398 VTAIL.n255 VTAIL.n179 104.615
R399 VTAIL.n256 VTAIL.n255 104.615
R400 VTAIL.n604 VTAIL.n603 104.615
R401 VTAIL.n603 VTAIL.n527 104.615
R402 VTAIL.n532 VTAIL.n527 104.615
R403 VTAIL.n596 VTAIL.n532 104.615
R404 VTAIL.n596 VTAIL.n595 104.615
R405 VTAIL.n595 VTAIL.n533 104.615
R406 VTAIL.n588 VTAIL.n533 104.615
R407 VTAIL.n588 VTAIL.n587 104.615
R408 VTAIL.n587 VTAIL.n537 104.615
R409 VTAIL.n580 VTAIL.n537 104.615
R410 VTAIL.n580 VTAIL.n579 104.615
R411 VTAIL.n579 VTAIL.n541 104.615
R412 VTAIL.n572 VTAIL.n541 104.615
R413 VTAIL.n572 VTAIL.n571 104.615
R414 VTAIL.n571 VTAIL.n545 104.615
R415 VTAIL.n564 VTAIL.n545 104.615
R416 VTAIL.n564 VTAIL.n563 104.615
R417 VTAIL.n563 VTAIL.n549 104.615
R418 VTAIL.n556 VTAIL.n549 104.615
R419 VTAIL.n556 VTAIL.n555 104.615
R420 VTAIL.n516 VTAIL.n515 104.615
R421 VTAIL.n515 VTAIL.n439 104.615
R422 VTAIL.n444 VTAIL.n439 104.615
R423 VTAIL.n508 VTAIL.n444 104.615
R424 VTAIL.n508 VTAIL.n507 104.615
R425 VTAIL.n507 VTAIL.n445 104.615
R426 VTAIL.n500 VTAIL.n445 104.615
R427 VTAIL.n500 VTAIL.n499 104.615
R428 VTAIL.n499 VTAIL.n449 104.615
R429 VTAIL.n492 VTAIL.n449 104.615
R430 VTAIL.n492 VTAIL.n491 104.615
R431 VTAIL.n491 VTAIL.n453 104.615
R432 VTAIL.n484 VTAIL.n453 104.615
R433 VTAIL.n484 VTAIL.n483 104.615
R434 VTAIL.n483 VTAIL.n457 104.615
R435 VTAIL.n476 VTAIL.n457 104.615
R436 VTAIL.n476 VTAIL.n475 104.615
R437 VTAIL.n475 VTAIL.n461 104.615
R438 VTAIL.n468 VTAIL.n461 104.615
R439 VTAIL.n468 VTAIL.n467 104.615
R440 VTAIL.n430 VTAIL.n429 104.615
R441 VTAIL.n429 VTAIL.n353 104.615
R442 VTAIL.n358 VTAIL.n353 104.615
R443 VTAIL.n422 VTAIL.n358 104.615
R444 VTAIL.n422 VTAIL.n421 104.615
R445 VTAIL.n421 VTAIL.n359 104.615
R446 VTAIL.n414 VTAIL.n359 104.615
R447 VTAIL.n414 VTAIL.n413 104.615
R448 VTAIL.n413 VTAIL.n363 104.615
R449 VTAIL.n406 VTAIL.n363 104.615
R450 VTAIL.n406 VTAIL.n405 104.615
R451 VTAIL.n405 VTAIL.n367 104.615
R452 VTAIL.n398 VTAIL.n367 104.615
R453 VTAIL.n398 VTAIL.n397 104.615
R454 VTAIL.n397 VTAIL.n371 104.615
R455 VTAIL.n390 VTAIL.n371 104.615
R456 VTAIL.n390 VTAIL.n389 104.615
R457 VTAIL.n389 VTAIL.n375 104.615
R458 VTAIL.n382 VTAIL.n375 104.615
R459 VTAIL.n382 VTAIL.n381 104.615
R460 VTAIL.n342 VTAIL.n341 104.615
R461 VTAIL.n341 VTAIL.n265 104.615
R462 VTAIL.n270 VTAIL.n265 104.615
R463 VTAIL.n334 VTAIL.n270 104.615
R464 VTAIL.n334 VTAIL.n333 104.615
R465 VTAIL.n333 VTAIL.n271 104.615
R466 VTAIL.n326 VTAIL.n271 104.615
R467 VTAIL.n326 VTAIL.n325 104.615
R468 VTAIL.n325 VTAIL.n275 104.615
R469 VTAIL.n318 VTAIL.n275 104.615
R470 VTAIL.n318 VTAIL.n317 104.615
R471 VTAIL.n317 VTAIL.n279 104.615
R472 VTAIL.n310 VTAIL.n279 104.615
R473 VTAIL.n310 VTAIL.n309 104.615
R474 VTAIL.n309 VTAIL.n283 104.615
R475 VTAIL.n302 VTAIL.n283 104.615
R476 VTAIL.n302 VTAIL.n301 104.615
R477 VTAIL.n301 VTAIL.n287 104.615
R478 VTAIL.n294 VTAIL.n287 104.615
R479 VTAIL.n294 VTAIL.n293 104.615
R480 VTAIL.n639 VTAIL.t12 52.3082
R481 VTAIL.n31 VTAIL.t11 52.3082
R482 VTAIL.n117 VTAIL.t3 52.3082
R483 VTAIL.n205 VTAIL.t6 52.3082
R484 VTAIL.n555 VTAIL.t0 52.3082
R485 VTAIL.n467 VTAIL.t4 52.3082
R486 VTAIL.n381 VTAIL.t10 52.3082
R487 VTAIL.n293 VTAIL.t13 52.3082
R488 VTAIL.n523 VTAIL.n522 43.9698
R489 VTAIL.n349 VTAIL.n348 43.9698
R490 VTAIL.n1 VTAIL.n0 43.9697
R491 VTAIL.n175 VTAIL.n174 43.9697
R492 VTAIL.n695 VTAIL.n694 31.9914
R493 VTAIL.n87 VTAIL.n86 31.9914
R494 VTAIL.n173 VTAIL.n172 31.9914
R495 VTAIL.n261 VTAIL.n260 31.9914
R496 VTAIL.n609 VTAIL.n608 31.9914
R497 VTAIL.n521 VTAIL.n520 31.9914
R498 VTAIL.n435 VTAIL.n434 31.9914
R499 VTAIL.n347 VTAIL.n346 31.9914
R500 VTAIL.n695 VTAIL.n609 29.2893
R501 VTAIL.n347 VTAIL.n261 29.2893
R502 VTAIL.n638 VTAIL.n637 15.6677
R503 VTAIL.n30 VTAIL.n29 15.6677
R504 VTAIL.n116 VTAIL.n115 15.6677
R505 VTAIL.n204 VTAIL.n203 15.6677
R506 VTAIL.n554 VTAIL.n553 15.6677
R507 VTAIL.n466 VTAIL.n465 15.6677
R508 VTAIL.n380 VTAIL.n379 15.6677
R509 VTAIL.n292 VTAIL.n291 15.6677
R510 VTAIL.n683 VTAIL.n614 13.1884
R511 VTAIL.n75 VTAIL.n6 13.1884
R512 VTAIL.n161 VTAIL.n92 13.1884
R513 VTAIL.n249 VTAIL.n180 13.1884
R514 VTAIL.n530 VTAIL.n528 13.1884
R515 VTAIL.n442 VTAIL.n440 13.1884
R516 VTAIL.n356 VTAIL.n354 13.1884
R517 VTAIL.n268 VTAIL.n266 13.1884
R518 VTAIL.n641 VTAIL.n636 12.8005
R519 VTAIL.n684 VTAIL.n616 12.8005
R520 VTAIL.n688 VTAIL.n687 12.8005
R521 VTAIL.n33 VTAIL.n28 12.8005
R522 VTAIL.n76 VTAIL.n8 12.8005
R523 VTAIL.n80 VTAIL.n79 12.8005
R524 VTAIL.n119 VTAIL.n114 12.8005
R525 VTAIL.n162 VTAIL.n94 12.8005
R526 VTAIL.n166 VTAIL.n165 12.8005
R527 VTAIL.n207 VTAIL.n202 12.8005
R528 VTAIL.n250 VTAIL.n182 12.8005
R529 VTAIL.n254 VTAIL.n253 12.8005
R530 VTAIL.n602 VTAIL.n601 12.8005
R531 VTAIL.n598 VTAIL.n597 12.8005
R532 VTAIL.n557 VTAIL.n552 12.8005
R533 VTAIL.n514 VTAIL.n513 12.8005
R534 VTAIL.n510 VTAIL.n509 12.8005
R535 VTAIL.n469 VTAIL.n464 12.8005
R536 VTAIL.n428 VTAIL.n427 12.8005
R537 VTAIL.n424 VTAIL.n423 12.8005
R538 VTAIL.n383 VTAIL.n378 12.8005
R539 VTAIL.n340 VTAIL.n339 12.8005
R540 VTAIL.n336 VTAIL.n335 12.8005
R541 VTAIL.n295 VTAIL.n290 12.8005
R542 VTAIL.n642 VTAIL.n634 12.0247
R543 VTAIL.n679 VTAIL.n678 12.0247
R544 VTAIL.n691 VTAIL.n612 12.0247
R545 VTAIL.n34 VTAIL.n26 12.0247
R546 VTAIL.n71 VTAIL.n70 12.0247
R547 VTAIL.n83 VTAIL.n4 12.0247
R548 VTAIL.n120 VTAIL.n112 12.0247
R549 VTAIL.n157 VTAIL.n156 12.0247
R550 VTAIL.n169 VTAIL.n90 12.0247
R551 VTAIL.n208 VTAIL.n200 12.0247
R552 VTAIL.n245 VTAIL.n244 12.0247
R553 VTAIL.n257 VTAIL.n178 12.0247
R554 VTAIL.n605 VTAIL.n526 12.0247
R555 VTAIL.n594 VTAIL.n531 12.0247
R556 VTAIL.n558 VTAIL.n550 12.0247
R557 VTAIL.n517 VTAIL.n438 12.0247
R558 VTAIL.n506 VTAIL.n443 12.0247
R559 VTAIL.n470 VTAIL.n462 12.0247
R560 VTAIL.n431 VTAIL.n352 12.0247
R561 VTAIL.n420 VTAIL.n357 12.0247
R562 VTAIL.n384 VTAIL.n376 12.0247
R563 VTAIL.n343 VTAIL.n264 12.0247
R564 VTAIL.n332 VTAIL.n269 12.0247
R565 VTAIL.n296 VTAIL.n288 12.0247
R566 VTAIL.n646 VTAIL.n645 11.249
R567 VTAIL.n677 VTAIL.n618 11.249
R568 VTAIL.n692 VTAIL.n610 11.249
R569 VTAIL.n38 VTAIL.n37 11.249
R570 VTAIL.n69 VTAIL.n10 11.249
R571 VTAIL.n84 VTAIL.n2 11.249
R572 VTAIL.n124 VTAIL.n123 11.249
R573 VTAIL.n155 VTAIL.n96 11.249
R574 VTAIL.n170 VTAIL.n88 11.249
R575 VTAIL.n212 VTAIL.n211 11.249
R576 VTAIL.n243 VTAIL.n184 11.249
R577 VTAIL.n258 VTAIL.n176 11.249
R578 VTAIL.n606 VTAIL.n524 11.249
R579 VTAIL.n593 VTAIL.n534 11.249
R580 VTAIL.n562 VTAIL.n561 11.249
R581 VTAIL.n518 VTAIL.n436 11.249
R582 VTAIL.n505 VTAIL.n446 11.249
R583 VTAIL.n474 VTAIL.n473 11.249
R584 VTAIL.n432 VTAIL.n350 11.249
R585 VTAIL.n419 VTAIL.n360 11.249
R586 VTAIL.n388 VTAIL.n387 11.249
R587 VTAIL.n344 VTAIL.n262 11.249
R588 VTAIL.n331 VTAIL.n272 11.249
R589 VTAIL.n300 VTAIL.n299 11.249
R590 VTAIL.n649 VTAIL.n632 10.4732
R591 VTAIL.n674 VTAIL.n673 10.4732
R592 VTAIL.n41 VTAIL.n24 10.4732
R593 VTAIL.n66 VTAIL.n65 10.4732
R594 VTAIL.n127 VTAIL.n110 10.4732
R595 VTAIL.n152 VTAIL.n151 10.4732
R596 VTAIL.n215 VTAIL.n198 10.4732
R597 VTAIL.n240 VTAIL.n239 10.4732
R598 VTAIL.n590 VTAIL.n589 10.4732
R599 VTAIL.n565 VTAIL.n548 10.4732
R600 VTAIL.n502 VTAIL.n501 10.4732
R601 VTAIL.n477 VTAIL.n460 10.4732
R602 VTAIL.n416 VTAIL.n415 10.4732
R603 VTAIL.n391 VTAIL.n374 10.4732
R604 VTAIL.n328 VTAIL.n327 10.4732
R605 VTAIL.n303 VTAIL.n286 10.4732
R606 VTAIL.n650 VTAIL.n630 9.69747
R607 VTAIL.n670 VTAIL.n620 9.69747
R608 VTAIL.n42 VTAIL.n22 9.69747
R609 VTAIL.n62 VTAIL.n12 9.69747
R610 VTAIL.n128 VTAIL.n108 9.69747
R611 VTAIL.n148 VTAIL.n98 9.69747
R612 VTAIL.n216 VTAIL.n196 9.69747
R613 VTAIL.n236 VTAIL.n186 9.69747
R614 VTAIL.n586 VTAIL.n536 9.69747
R615 VTAIL.n566 VTAIL.n546 9.69747
R616 VTAIL.n498 VTAIL.n448 9.69747
R617 VTAIL.n478 VTAIL.n458 9.69747
R618 VTAIL.n412 VTAIL.n362 9.69747
R619 VTAIL.n392 VTAIL.n372 9.69747
R620 VTAIL.n324 VTAIL.n274 9.69747
R621 VTAIL.n304 VTAIL.n284 9.69747
R622 VTAIL.n694 VTAIL.n693 9.45567
R623 VTAIL.n86 VTAIL.n85 9.45567
R624 VTAIL.n172 VTAIL.n171 9.45567
R625 VTAIL.n260 VTAIL.n259 9.45567
R626 VTAIL.n608 VTAIL.n607 9.45567
R627 VTAIL.n520 VTAIL.n519 9.45567
R628 VTAIL.n434 VTAIL.n433 9.45567
R629 VTAIL.n346 VTAIL.n345 9.45567
R630 VTAIL.n693 VTAIL.n692 9.3005
R631 VTAIL.n612 VTAIL.n611 9.3005
R632 VTAIL.n687 VTAIL.n686 9.3005
R633 VTAIL.n659 VTAIL.n658 9.3005
R634 VTAIL.n628 VTAIL.n627 9.3005
R635 VTAIL.n653 VTAIL.n652 9.3005
R636 VTAIL.n651 VTAIL.n650 9.3005
R637 VTAIL.n632 VTAIL.n631 9.3005
R638 VTAIL.n645 VTAIL.n644 9.3005
R639 VTAIL.n643 VTAIL.n642 9.3005
R640 VTAIL.n636 VTAIL.n635 9.3005
R641 VTAIL.n661 VTAIL.n660 9.3005
R642 VTAIL.n624 VTAIL.n623 9.3005
R643 VTAIL.n667 VTAIL.n666 9.3005
R644 VTAIL.n669 VTAIL.n668 9.3005
R645 VTAIL.n620 VTAIL.n619 9.3005
R646 VTAIL.n675 VTAIL.n674 9.3005
R647 VTAIL.n677 VTAIL.n676 9.3005
R648 VTAIL.n678 VTAIL.n615 9.3005
R649 VTAIL.n685 VTAIL.n684 9.3005
R650 VTAIL.n85 VTAIL.n84 9.3005
R651 VTAIL.n4 VTAIL.n3 9.3005
R652 VTAIL.n79 VTAIL.n78 9.3005
R653 VTAIL.n51 VTAIL.n50 9.3005
R654 VTAIL.n20 VTAIL.n19 9.3005
R655 VTAIL.n45 VTAIL.n44 9.3005
R656 VTAIL.n43 VTAIL.n42 9.3005
R657 VTAIL.n24 VTAIL.n23 9.3005
R658 VTAIL.n37 VTAIL.n36 9.3005
R659 VTAIL.n35 VTAIL.n34 9.3005
R660 VTAIL.n28 VTAIL.n27 9.3005
R661 VTAIL.n53 VTAIL.n52 9.3005
R662 VTAIL.n16 VTAIL.n15 9.3005
R663 VTAIL.n59 VTAIL.n58 9.3005
R664 VTAIL.n61 VTAIL.n60 9.3005
R665 VTAIL.n12 VTAIL.n11 9.3005
R666 VTAIL.n67 VTAIL.n66 9.3005
R667 VTAIL.n69 VTAIL.n68 9.3005
R668 VTAIL.n70 VTAIL.n7 9.3005
R669 VTAIL.n77 VTAIL.n76 9.3005
R670 VTAIL.n171 VTAIL.n170 9.3005
R671 VTAIL.n90 VTAIL.n89 9.3005
R672 VTAIL.n165 VTAIL.n164 9.3005
R673 VTAIL.n137 VTAIL.n136 9.3005
R674 VTAIL.n106 VTAIL.n105 9.3005
R675 VTAIL.n131 VTAIL.n130 9.3005
R676 VTAIL.n129 VTAIL.n128 9.3005
R677 VTAIL.n110 VTAIL.n109 9.3005
R678 VTAIL.n123 VTAIL.n122 9.3005
R679 VTAIL.n121 VTAIL.n120 9.3005
R680 VTAIL.n114 VTAIL.n113 9.3005
R681 VTAIL.n139 VTAIL.n138 9.3005
R682 VTAIL.n102 VTAIL.n101 9.3005
R683 VTAIL.n145 VTAIL.n144 9.3005
R684 VTAIL.n147 VTAIL.n146 9.3005
R685 VTAIL.n98 VTAIL.n97 9.3005
R686 VTAIL.n153 VTAIL.n152 9.3005
R687 VTAIL.n155 VTAIL.n154 9.3005
R688 VTAIL.n156 VTAIL.n93 9.3005
R689 VTAIL.n163 VTAIL.n162 9.3005
R690 VTAIL.n259 VTAIL.n258 9.3005
R691 VTAIL.n178 VTAIL.n177 9.3005
R692 VTAIL.n253 VTAIL.n252 9.3005
R693 VTAIL.n225 VTAIL.n224 9.3005
R694 VTAIL.n194 VTAIL.n193 9.3005
R695 VTAIL.n219 VTAIL.n218 9.3005
R696 VTAIL.n217 VTAIL.n216 9.3005
R697 VTAIL.n198 VTAIL.n197 9.3005
R698 VTAIL.n211 VTAIL.n210 9.3005
R699 VTAIL.n209 VTAIL.n208 9.3005
R700 VTAIL.n202 VTAIL.n201 9.3005
R701 VTAIL.n227 VTAIL.n226 9.3005
R702 VTAIL.n190 VTAIL.n189 9.3005
R703 VTAIL.n233 VTAIL.n232 9.3005
R704 VTAIL.n235 VTAIL.n234 9.3005
R705 VTAIL.n186 VTAIL.n185 9.3005
R706 VTAIL.n241 VTAIL.n240 9.3005
R707 VTAIL.n243 VTAIL.n242 9.3005
R708 VTAIL.n244 VTAIL.n181 9.3005
R709 VTAIL.n251 VTAIL.n250 9.3005
R710 VTAIL.n540 VTAIL.n539 9.3005
R711 VTAIL.n583 VTAIL.n582 9.3005
R712 VTAIL.n585 VTAIL.n584 9.3005
R713 VTAIL.n536 VTAIL.n535 9.3005
R714 VTAIL.n591 VTAIL.n590 9.3005
R715 VTAIL.n593 VTAIL.n592 9.3005
R716 VTAIL.n531 VTAIL.n529 9.3005
R717 VTAIL.n599 VTAIL.n598 9.3005
R718 VTAIL.n607 VTAIL.n606 9.3005
R719 VTAIL.n526 VTAIL.n525 9.3005
R720 VTAIL.n601 VTAIL.n600 9.3005
R721 VTAIL.n577 VTAIL.n576 9.3005
R722 VTAIL.n575 VTAIL.n574 9.3005
R723 VTAIL.n544 VTAIL.n543 9.3005
R724 VTAIL.n569 VTAIL.n568 9.3005
R725 VTAIL.n567 VTAIL.n566 9.3005
R726 VTAIL.n548 VTAIL.n547 9.3005
R727 VTAIL.n561 VTAIL.n560 9.3005
R728 VTAIL.n559 VTAIL.n558 9.3005
R729 VTAIL.n552 VTAIL.n551 9.3005
R730 VTAIL.n452 VTAIL.n451 9.3005
R731 VTAIL.n495 VTAIL.n494 9.3005
R732 VTAIL.n497 VTAIL.n496 9.3005
R733 VTAIL.n448 VTAIL.n447 9.3005
R734 VTAIL.n503 VTAIL.n502 9.3005
R735 VTAIL.n505 VTAIL.n504 9.3005
R736 VTAIL.n443 VTAIL.n441 9.3005
R737 VTAIL.n511 VTAIL.n510 9.3005
R738 VTAIL.n519 VTAIL.n518 9.3005
R739 VTAIL.n438 VTAIL.n437 9.3005
R740 VTAIL.n513 VTAIL.n512 9.3005
R741 VTAIL.n489 VTAIL.n488 9.3005
R742 VTAIL.n487 VTAIL.n486 9.3005
R743 VTAIL.n456 VTAIL.n455 9.3005
R744 VTAIL.n481 VTAIL.n480 9.3005
R745 VTAIL.n479 VTAIL.n478 9.3005
R746 VTAIL.n460 VTAIL.n459 9.3005
R747 VTAIL.n473 VTAIL.n472 9.3005
R748 VTAIL.n471 VTAIL.n470 9.3005
R749 VTAIL.n464 VTAIL.n463 9.3005
R750 VTAIL.n366 VTAIL.n365 9.3005
R751 VTAIL.n409 VTAIL.n408 9.3005
R752 VTAIL.n411 VTAIL.n410 9.3005
R753 VTAIL.n362 VTAIL.n361 9.3005
R754 VTAIL.n417 VTAIL.n416 9.3005
R755 VTAIL.n419 VTAIL.n418 9.3005
R756 VTAIL.n357 VTAIL.n355 9.3005
R757 VTAIL.n425 VTAIL.n424 9.3005
R758 VTAIL.n433 VTAIL.n432 9.3005
R759 VTAIL.n352 VTAIL.n351 9.3005
R760 VTAIL.n427 VTAIL.n426 9.3005
R761 VTAIL.n403 VTAIL.n402 9.3005
R762 VTAIL.n401 VTAIL.n400 9.3005
R763 VTAIL.n370 VTAIL.n369 9.3005
R764 VTAIL.n395 VTAIL.n394 9.3005
R765 VTAIL.n393 VTAIL.n392 9.3005
R766 VTAIL.n374 VTAIL.n373 9.3005
R767 VTAIL.n387 VTAIL.n386 9.3005
R768 VTAIL.n385 VTAIL.n384 9.3005
R769 VTAIL.n378 VTAIL.n377 9.3005
R770 VTAIL.n278 VTAIL.n277 9.3005
R771 VTAIL.n321 VTAIL.n320 9.3005
R772 VTAIL.n323 VTAIL.n322 9.3005
R773 VTAIL.n274 VTAIL.n273 9.3005
R774 VTAIL.n329 VTAIL.n328 9.3005
R775 VTAIL.n331 VTAIL.n330 9.3005
R776 VTAIL.n269 VTAIL.n267 9.3005
R777 VTAIL.n337 VTAIL.n336 9.3005
R778 VTAIL.n345 VTAIL.n344 9.3005
R779 VTAIL.n264 VTAIL.n263 9.3005
R780 VTAIL.n339 VTAIL.n338 9.3005
R781 VTAIL.n315 VTAIL.n314 9.3005
R782 VTAIL.n313 VTAIL.n312 9.3005
R783 VTAIL.n282 VTAIL.n281 9.3005
R784 VTAIL.n307 VTAIL.n306 9.3005
R785 VTAIL.n305 VTAIL.n304 9.3005
R786 VTAIL.n286 VTAIL.n285 9.3005
R787 VTAIL.n299 VTAIL.n298 9.3005
R788 VTAIL.n297 VTAIL.n296 9.3005
R789 VTAIL.n290 VTAIL.n289 9.3005
R790 VTAIL.n654 VTAIL.n653 8.92171
R791 VTAIL.n669 VTAIL.n622 8.92171
R792 VTAIL.n46 VTAIL.n45 8.92171
R793 VTAIL.n61 VTAIL.n14 8.92171
R794 VTAIL.n132 VTAIL.n131 8.92171
R795 VTAIL.n147 VTAIL.n100 8.92171
R796 VTAIL.n220 VTAIL.n219 8.92171
R797 VTAIL.n235 VTAIL.n188 8.92171
R798 VTAIL.n585 VTAIL.n538 8.92171
R799 VTAIL.n570 VTAIL.n569 8.92171
R800 VTAIL.n497 VTAIL.n450 8.92171
R801 VTAIL.n482 VTAIL.n481 8.92171
R802 VTAIL.n411 VTAIL.n364 8.92171
R803 VTAIL.n396 VTAIL.n395 8.92171
R804 VTAIL.n323 VTAIL.n276 8.92171
R805 VTAIL.n308 VTAIL.n307 8.92171
R806 VTAIL.n657 VTAIL.n628 8.14595
R807 VTAIL.n666 VTAIL.n665 8.14595
R808 VTAIL.n49 VTAIL.n20 8.14595
R809 VTAIL.n58 VTAIL.n57 8.14595
R810 VTAIL.n135 VTAIL.n106 8.14595
R811 VTAIL.n144 VTAIL.n143 8.14595
R812 VTAIL.n223 VTAIL.n194 8.14595
R813 VTAIL.n232 VTAIL.n231 8.14595
R814 VTAIL.n582 VTAIL.n581 8.14595
R815 VTAIL.n573 VTAIL.n544 8.14595
R816 VTAIL.n494 VTAIL.n493 8.14595
R817 VTAIL.n485 VTAIL.n456 8.14595
R818 VTAIL.n408 VTAIL.n407 8.14595
R819 VTAIL.n399 VTAIL.n370 8.14595
R820 VTAIL.n320 VTAIL.n319 8.14595
R821 VTAIL.n311 VTAIL.n282 8.14595
R822 VTAIL.n658 VTAIL.n626 7.3702
R823 VTAIL.n662 VTAIL.n624 7.3702
R824 VTAIL.n50 VTAIL.n18 7.3702
R825 VTAIL.n54 VTAIL.n16 7.3702
R826 VTAIL.n136 VTAIL.n104 7.3702
R827 VTAIL.n140 VTAIL.n102 7.3702
R828 VTAIL.n224 VTAIL.n192 7.3702
R829 VTAIL.n228 VTAIL.n190 7.3702
R830 VTAIL.n578 VTAIL.n540 7.3702
R831 VTAIL.n574 VTAIL.n542 7.3702
R832 VTAIL.n490 VTAIL.n452 7.3702
R833 VTAIL.n486 VTAIL.n454 7.3702
R834 VTAIL.n404 VTAIL.n366 7.3702
R835 VTAIL.n400 VTAIL.n368 7.3702
R836 VTAIL.n316 VTAIL.n278 7.3702
R837 VTAIL.n312 VTAIL.n280 7.3702
R838 VTAIL.n661 VTAIL.n626 6.59444
R839 VTAIL.n662 VTAIL.n661 6.59444
R840 VTAIL.n53 VTAIL.n18 6.59444
R841 VTAIL.n54 VTAIL.n53 6.59444
R842 VTAIL.n139 VTAIL.n104 6.59444
R843 VTAIL.n140 VTAIL.n139 6.59444
R844 VTAIL.n227 VTAIL.n192 6.59444
R845 VTAIL.n228 VTAIL.n227 6.59444
R846 VTAIL.n578 VTAIL.n577 6.59444
R847 VTAIL.n577 VTAIL.n542 6.59444
R848 VTAIL.n490 VTAIL.n489 6.59444
R849 VTAIL.n489 VTAIL.n454 6.59444
R850 VTAIL.n404 VTAIL.n403 6.59444
R851 VTAIL.n403 VTAIL.n368 6.59444
R852 VTAIL.n316 VTAIL.n315 6.59444
R853 VTAIL.n315 VTAIL.n280 6.59444
R854 VTAIL.n658 VTAIL.n657 5.81868
R855 VTAIL.n665 VTAIL.n624 5.81868
R856 VTAIL.n50 VTAIL.n49 5.81868
R857 VTAIL.n57 VTAIL.n16 5.81868
R858 VTAIL.n136 VTAIL.n135 5.81868
R859 VTAIL.n143 VTAIL.n102 5.81868
R860 VTAIL.n224 VTAIL.n223 5.81868
R861 VTAIL.n231 VTAIL.n190 5.81868
R862 VTAIL.n581 VTAIL.n540 5.81868
R863 VTAIL.n574 VTAIL.n573 5.81868
R864 VTAIL.n493 VTAIL.n452 5.81868
R865 VTAIL.n486 VTAIL.n485 5.81868
R866 VTAIL.n407 VTAIL.n366 5.81868
R867 VTAIL.n400 VTAIL.n399 5.81868
R868 VTAIL.n319 VTAIL.n278 5.81868
R869 VTAIL.n312 VTAIL.n311 5.81868
R870 VTAIL.n654 VTAIL.n628 5.04292
R871 VTAIL.n666 VTAIL.n622 5.04292
R872 VTAIL.n46 VTAIL.n20 5.04292
R873 VTAIL.n58 VTAIL.n14 5.04292
R874 VTAIL.n132 VTAIL.n106 5.04292
R875 VTAIL.n144 VTAIL.n100 5.04292
R876 VTAIL.n220 VTAIL.n194 5.04292
R877 VTAIL.n232 VTAIL.n188 5.04292
R878 VTAIL.n582 VTAIL.n538 5.04292
R879 VTAIL.n570 VTAIL.n544 5.04292
R880 VTAIL.n494 VTAIL.n450 5.04292
R881 VTAIL.n482 VTAIL.n456 5.04292
R882 VTAIL.n408 VTAIL.n364 5.04292
R883 VTAIL.n396 VTAIL.n370 5.04292
R884 VTAIL.n320 VTAIL.n276 5.04292
R885 VTAIL.n308 VTAIL.n282 5.04292
R886 VTAIL.n637 VTAIL.n635 4.38563
R887 VTAIL.n29 VTAIL.n27 4.38563
R888 VTAIL.n115 VTAIL.n113 4.38563
R889 VTAIL.n203 VTAIL.n201 4.38563
R890 VTAIL.n553 VTAIL.n551 4.38563
R891 VTAIL.n465 VTAIL.n463 4.38563
R892 VTAIL.n379 VTAIL.n377 4.38563
R893 VTAIL.n291 VTAIL.n289 4.38563
R894 VTAIL.n653 VTAIL.n630 4.26717
R895 VTAIL.n670 VTAIL.n669 4.26717
R896 VTAIL.n45 VTAIL.n22 4.26717
R897 VTAIL.n62 VTAIL.n61 4.26717
R898 VTAIL.n131 VTAIL.n108 4.26717
R899 VTAIL.n148 VTAIL.n147 4.26717
R900 VTAIL.n219 VTAIL.n196 4.26717
R901 VTAIL.n236 VTAIL.n235 4.26717
R902 VTAIL.n586 VTAIL.n585 4.26717
R903 VTAIL.n569 VTAIL.n546 4.26717
R904 VTAIL.n498 VTAIL.n497 4.26717
R905 VTAIL.n481 VTAIL.n458 4.26717
R906 VTAIL.n412 VTAIL.n411 4.26717
R907 VTAIL.n395 VTAIL.n372 4.26717
R908 VTAIL.n324 VTAIL.n323 4.26717
R909 VTAIL.n307 VTAIL.n284 4.26717
R910 VTAIL.n349 VTAIL.n347 3.69016
R911 VTAIL.n435 VTAIL.n349 3.69016
R912 VTAIL.n523 VTAIL.n521 3.69016
R913 VTAIL.n609 VTAIL.n523 3.69016
R914 VTAIL.n261 VTAIL.n175 3.69016
R915 VTAIL.n175 VTAIL.n173 3.69016
R916 VTAIL.n87 VTAIL.n1 3.69016
R917 VTAIL VTAIL.n695 3.63197
R918 VTAIL.n650 VTAIL.n649 3.49141
R919 VTAIL.n673 VTAIL.n620 3.49141
R920 VTAIL.n42 VTAIL.n41 3.49141
R921 VTAIL.n65 VTAIL.n12 3.49141
R922 VTAIL.n128 VTAIL.n127 3.49141
R923 VTAIL.n151 VTAIL.n98 3.49141
R924 VTAIL.n216 VTAIL.n215 3.49141
R925 VTAIL.n239 VTAIL.n186 3.49141
R926 VTAIL.n589 VTAIL.n536 3.49141
R927 VTAIL.n566 VTAIL.n565 3.49141
R928 VTAIL.n501 VTAIL.n448 3.49141
R929 VTAIL.n478 VTAIL.n477 3.49141
R930 VTAIL.n415 VTAIL.n362 3.49141
R931 VTAIL.n392 VTAIL.n391 3.49141
R932 VTAIL.n327 VTAIL.n274 3.49141
R933 VTAIL.n304 VTAIL.n303 3.49141
R934 VTAIL.n646 VTAIL.n632 2.71565
R935 VTAIL.n674 VTAIL.n618 2.71565
R936 VTAIL.n694 VTAIL.n610 2.71565
R937 VTAIL.n38 VTAIL.n24 2.71565
R938 VTAIL.n66 VTAIL.n10 2.71565
R939 VTAIL.n86 VTAIL.n2 2.71565
R940 VTAIL.n124 VTAIL.n110 2.71565
R941 VTAIL.n152 VTAIL.n96 2.71565
R942 VTAIL.n172 VTAIL.n88 2.71565
R943 VTAIL.n212 VTAIL.n198 2.71565
R944 VTAIL.n240 VTAIL.n184 2.71565
R945 VTAIL.n260 VTAIL.n176 2.71565
R946 VTAIL.n608 VTAIL.n524 2.71565
R947 VTAIL.n590 VTAIL.n534 2.71565
R948 VTAIL.n562 VTAIL.n548 2.71565
R949 VTAIL.n520 VTAIL.n436 2.71565
R950 VTAIL.n502 VTAIL.n446 2.71565
R951 VTAIL.n474 VTAIL.n460 2.71565
R952 VTAIL.n434 VTAIL.n350 2.71565
R953 VTAIL.n416 VTAIL.n360 2.71565
R954 VTAIL.n388 VTAIL.n374 2.71565
R955 VTAIL.n346 VTAIL.n262 2.71565
R956 VTAIL.n328 VTAIL.n272 2.71565
R957 VTAIL.n300 VTAIL.n286 2.71565
R958 VTAIL.n645 VTAIL.n634 1.93989
R959 VTAIL.n679 VTAIL.n677 1.93989
R960 VTAIL.n692 VTAIL.n691 1.93989
R961 VTAIL.n37 VTAIL.n26 1.93989
R962 VTAIL.n71 VTAIL.n69 1.93989
R963 VTAIL.n84 VTAIL.n83 1.93989
R964 VTAIL.n123 VTAIL.n112 1.93989
R965 VTAIL.n157 VTAIL.n155 1.93989
R966 VTAIL.n170 VTAIL.n169 1.93989
R967 VTAIL.n211 VTAIL.n200 1.93989
R968 VTAIL.n245 VTAIL.n243 1.93989
R969 VTAIL.n258 VTAIL.n257 1.93989
R970 VTAIL.n606 VTAIL.n605 1.93989
R971 VTAIL.n594 VTAIL.n593 1.93989
R972 VTAIL.n561 VTAIL.n550 1.93989
R973 VTAIL.n518 VTAIL.n517 1.93989
R974 VTAIL.n506 VTAIL.n505 1.93989
R975 VTAIL.n473 VTAIL.n462 1.93989
R976 VTAIL.n432 VTAIL.n431 1.93989
R977 VTAIL.n420 VTAIL.n419 1.93989
R978 VTAIL.n387 VTAIL.n376 1.93989
R979 VTAIL.n344 VTAIL.n343 1.93989
R980 VTAIL.n332 VTAIL.n331 1.93989
R981 VTAIL.n299 VTAIL.n288 1.93989
R982 VTAIL.n0 VTAIL.t8 1.2904
R983 VTAIL.n0 VTAIL.t7 1.2904
R984 VTAIL.n174 VTAIL.t5 1.2904
R985 VTAIL.n174 VTAIL.t2 1.2904
R986 VTAIL.n522 VTAIL.t15 1.2904
R987 VTAIL.n522 VTAIL.t1 1.2904
R988 VTAIL.n348 VTAIL.t9 1.2904
R989 VTAIL.n348 VTAIL.t14 1.2904
R990 VTAIL.n642 VTAIL.n641 1.16414
R991 VTAIL.n678 VTAIL.n616 1.16414
R992 VTAIL.n688 VTAIL.n612 1.16414
R993 VTAIL.n34 VTAIL.n33 1.16414
R994 VTAIL.n70 VTAIL.n8 1.16414
R995 VTAIL.n80 VTAIL.n4 1.16414
R996 VTAIL.n120 VTAIL.n119 1.16414
R997 VTAIL.n156 VTAIL.n94 1.16414
R998 VTAIL.n166 VTAIL.n90 1.16414
R999 VTAIL.n208 VTAIL.n207 1.16414
R1000 VTAIL.n244 VTAIL.n182 1.16414
R1001 VTAIL.n254 VTAIL.n178 1.16414
R1002 VTAIL.n602 VTAIL.n526 1.16414
R1003 VTAIL.n597 VTAIL.n531 1.16414
R1004 VTAIL.n558 VTAIL.n557 1.16414
R1005 VTAIL.n514 VTAIL.n438 1.16414
R1006 VTAIL.n509 VTAIL.n443 1.16414
R1007 VTAIL.n470 VTAIL.n469 1.16414
R1008 VTAIL.n428 VTAIL.n352 1.16414
R1009 VTAIL.n423 VTAIL.n357 1.16414
R1010 VTAIL.n384 VTAIL.n383 1.16414
R1011 VTAIL.n340 VTAIL.n264 1.16414
R1012 VTAIL.n335 VTAIL.n269 1.16414
R1013 VTAIL.n296 VTAIL.n295 1.16414
R1014 VTAIL.n521 VTAIL.n435 0.470328
R1015 VTAIL.n173 VTAIL.n87 0.470328
R1016 VTAIL.n638 VTAIL.n636 0.388379
R1017 VTAIL.n684 VTAIL.n683 0.388379
R1018 VTAIL.n687 VTAIL.n614 0.388379
R1019 VTAIL.n30 VTAIL.n28 0.388379
R1020 VTAIL.n76 VTAIL.n75 0.388379
R1021 VTAIL.n79 VTAIL.n6 0.388379
R1022 VTAIL.n116 VTAIL.n114 0.388379
R1023 VTAIL.n162 VTAIL.n161 0.388379
R1024 VTAIL.n165 VTAIL.n92 0.388379
R1025 VTAIL.n204 VTAIL.n202 0.388379
R1026 VTAIL.n250 VTAIL.n249 0.388379
R1027 VTAIL.n253 VTAIL.n180 0.388379
R1028 VTAIL.n601 VTAIL.n528 0.388379
R1029 VTAIL.n598 VTAIL.n530 0.388379
R1030 VTAIL.n554 VTAIL.n552 0.388379
R1031 VTAIL.n513 VTAIL.n440 0.388379
R1032 VTAIL.n510 VTAIL.n442 0.388379
R1033 VTAIL.n466 VTAIL.n464 0.388379
R1034 VTAIL.n427 VTAIL.n354 0.388379
R1035 VTAIL.n424 VTAIL.n356 0.388379
R1036 VTAIL.n380 VTAIL.n378 0.388379
R1037 VTAIL.n339 VTAIL.n266 0.388379
R1038 VTAIL.n336 VTAIL.n268 0.388379
R1039 VTAIL.n292 VTAIL.n290 0.388379
R1040 VTAIL.n643 VTAIL.n635 0.155672
R1041 VTAIL.n644 VTAIL.n643 0.155672
R1042 VTAIL.n644 VTAIL.n631 0.155672
R1043 VTAIL.n651 VTAIL.n631 0.155672
R1044 VTAIL.n652 VTAIL.n651 0.155672
R1045 VTAIL.n652 VTAIL.n627 0.155672
R1046 VTAIL.n659 VTAIL.n627 0.155672
R1047 VTAIL.n660 VTAIL.n659 0.155672
R1048 VTAIL.n660 VTAIL.n623 0.155672
R1049 VTAIL.n667 VTAIL.n623 0.155672
R1050 VTAIL.n668 VTAIL.n667 0.155672
R1051 VTAIL.n668 VTAIL.n619 0.155672
R1052 VTAIL.n675 VTAIL.n619 0.155672
R1053 VTAIL.n676 VTAIL.n675 0.155672
R1054 VTAIL.n676 VTAIL.n615 0.155672
R1055 VTAIL.n685 VTAIL.n615 0.155672
R1056 VTAIL.n686 VTAIL.n685 0.155672
R1057 VTAIL.n686 VTAIL.n611 0.155672
R1058 VTAIL.n693 VTAIL.n611 0.155672
R1059 VTAIL.n35 VTAIL.n27 0.155672
R1060 VTAIL.n36 VTAIL.n35 0.155672
R1061 VTAIL.n36 VTAIL.n23 0.155672
R1062 VTAIL.n43 VTAIL.n23 0.155672
R1063 VTAIL.n44 VTAIL.n43 0.155672
R1064 VTAIL.n44 VTAIL.n19 0.155672
R1065 VTAIL.n51 VTAIL.n19 0.155672
R1066 VTAIL.n52 VTAIL.n51 0.155672
R1067 VTAIL.n52 VTAIL.n15 0.155672
R1068 VTAIL.n59 VTAIL.n15 0.155672
R1069 VTAIL.n60 VTAIL.n59 0.155672
R1070 VTAIL.n60 VTAIL.n11 0.155672
R1071 VTAIL.n67 VTAIL.n11 0.155672
R1072 VTAIL.n68 VTAIL.n67 0.155672
R1073 VTAIL.n68 VTAIL.n7 0.155672
R1074 VTAIL.n77 VTAIL.n7 0.155672
R1075 VTAIL.n78 VTAIL.n77 0.155672
R1076 VTAIL.n78 VTAIL.n3 0.155672
R1077 VTAIL.n85 VTAIL.n3 0.155672
R1078 VTAIL.n121 VTAIL.n113 0.155672
R1079 VTAIL.n122 VTAIL.n121 0.155672
R1080 VTAIL.n122 VTAIL.n109 0.155672
R1081 VTAIL.n129 VTAIL.n109 0.155672
R1082 VTAIL.n130 VTAIL.n129 0.155672
R1083 VTAIL.n130 VTAIL.n105 0.155672
R1084 VTAIL.n137 VTAIL.n105 0.155672
R1085 VTAIL.n138 VTAIL.n137 0.155672
R1086 VTAIL.n138 VTAIL.n101 0.155672
R1087 VTAIL.n145 VTAIL.n101 0.155672
R1088 VTAIL.n146 VTAIL.n145 0.155672
R1089 VTAIL.n146 VTAIL.n97 0.155672
R1090 VTAIL.n153 VTAIL.n97 0.155672
R1091 VTAIL.n154 VTAIL.n153 0.155672
R1092 VTAIL.n154 VTAIL.n93 0.155672
R1093 VTAIL.n163 VTAIL.n93 0.155672
R1094 VTAIL.n164 VTAIL.n163 0.155672
R1095 VTAIL.n164 VTAIL.n89 0.155672
R1096 VTAIL.n171 VTAIL.n89 0.155672
R1097 VTAIL.n209 VTAIL.n201 0.155672
R1098 VTAIL.n210 VTAIL.n209 0.155672
R1099 VTAIL.n210 VTAIL.n197 0.155672
R1100 VTAIL.n217 VTAIL.n197 0.155672
R1101 VTAIL.n218 VTAIL.n217 0.155672
R1102 VTAIL.n218 VTAIL.n193 0.155672
R1103 VTAIL.n225 VTAIL.n193 0.155672
R1104 VTAIL.n226 VTAIL.n225 0.155672
R1105 VTAIL.n226 VTAIL.n189 0.155672
R1106 VTAIL.n233 VTAIL.n189 0.155672
R1107 VTAIL.n234 VTAIL.n233 0.155672
R1108 VTAIL.n234 VTAIL.n185 0.155672
R1109 VTAIL.n241 VTAIL.n185 0.155672
R1110 VTAIL.n242 VTAIL.n241 0.155672
R1111 VTAIL.n242 VTAIL.n181 0.155672
R1112 VTAIL.n251 VTAIL.n181 0.155672
R1113 VTAIL.n252 VTAIL.n251 0.155672
R1114 VTAIL.n252 VTAIL.n177 0.155672
R1115 VTAIL.n259 VTAIL.n177 0.155672
R1116 VTAIL.n607 VTAIL.n525 0.155672
R1117 VTAIL.n600 VTAIL.n525 0.155672
R1118 VTAIL.n600 VTAIL.n599 0.155672
R1119 VTAIL.n599 VTAIL.n529 0.155672
R1120 VTAIL.n592 VTAIL.n529 0.155672
R1121 VTAIL.n592 VTAIL.n591 0.155672
R1122 VTAIL.n591 VTAIL.n535 0.155672
R1123 VTAIL.n584 VTAIL.n535 0.155672
R1124 VTAIL.n584 VTAIL.n583 0.155672
R1125 VTAIL.n583 VTAIL.n539 0.155672
R1126 VTAIL.n576 VTAIL.n539 0.155672
R1127 VTAIL.n576 VTAIL.n575 0.155672
R1128 VTAIL.n575 VTAIL.n543 0.155672
R1129 VTAIL.n568 VTAIL.n543 0.155672
R1130 VTAIL.n568 VTAIL.n567 0.155672
R1131 VTAIL.n567 VTAIL.n547 0.155672
R1132 VTAIL.n560 VTAIL.n547 0.155672
R1133 VTAIL.n560 VTAIL.n559 0.155672
R1134 VTAIL.n559 VTAIL.n551 0.155672
R1135 VTAIL.n519 VTAIL.n437 0.155672
R1136 VTAIL.n512 VTAIL.n437 0.155672
R1137 VTAIL.n512 VTAIL.n511 0.155672
R1138 VTAIL.n511 VTAIL.n441 0.155672
R1139 VTAIL.n504 VTAIL.n441 0.155672
R1140 VTAIL.n504 VTAIL.n503 0.155672
R1141 VTAIL.n503 VTAIL.n447 0.155672
R1142 VTAIL.n496 VTAIL.n447 0.155672
R1143 VTAIL.n496 VTAIL.n495 0.155672
R1144 VTAIL.n495 VTAIL.n451 0.155672
R1145 VTAIL.n488 VTAIL.n451 0.155672
R1146 VTAIL.n488 VTAIL.n487 0.155672
R1147 VTAIL.n487 VTAIL.n455 0.155672
R1148 VTAIL.n480 VTAIL.n455 0.155672
R1149 VTAIL.n480 VTAIL.n479 0.155672
R1150 VTAIL.n479 VTAIL.n459 0.155672
R1151 VTAIL.n472 VTAIL.n459 0.155672
R1152 VTAIL.n472 VTAIL.n471 0.155672
R1153 VTAIL.n471 VTAIL.n463 0.155672
R1154 VTAIL.n433 VTAIL.n351 0.155672
R1155 VTAIL.n426 VTAIL.n351 0.155672
R1156 VTAIL.n426 VTAIL.n425 0.155672
R1157 VTAIL.n425 VTAIL.n355 0.155672
R1158 VTAIL.n418 VTAIL.n355 0.155672
R1159 VTAIL.n418 VTAIL.n417 0.155672
R1160 VTAIL.n417 VTAIL.n361 0.155672
R1161 VTAIL.n410 VTAIL.n361 0.155672
R1162 VTAIL.n410 VTAIL.n409 0.155672
R1163 VTAIL.n409 VTAIL.n365 0.155672
R1164 VTAIL.n402 VTAIL.n365 0.155672
R1165 VTAIL.n402 VTAIL.n401 0.155672
R1166 VTAIL.n401 VTAIL.n369 0.155672
R1167 VTAIL.n394 VTAIL.n369 0.155672
R1168 VTAIL.n394 VTAIL.n393 0.155672
R1169 VTAIL.n393 VTAIL.n373 0.155672
R1170 VTAIL.n386 VTAIL.n373 0.155672
R1171 VTAIL.n386 VTAIL.n385 0.155672
R1172 VTAIL.n385 VTAIL.n377 0.155672
R1173 VTAIL.n345 VTAIL.n263 0.155672
R1174 VTAIL.n338 VTAIL.n263 0.155672
R1175 VTAIL.n338 VTAIL.n337 0.155672
R1176 VTAIL.n337 VTAIL.n267 0.155672
R1177 VTAIL.n330 VTAIL.n267 0.155672
R1178 VTAIL.n330 VTAIL.n329 0.155672
R1179 VTAIL.n329 VTAIL.n273 0.155672
R1180 VTAIL.n322 VTAIL.n273 0.155672
R1181 VTAIL.n322 VTAIL.n321 0.155672
R1182 VTAIL.n321 VTAIL.n277 0.155672
R1183 VTAIL.n314 VTAIL.n277 0.155672
R1184 VTAIL.n314 VTAIL.n313 0.155672
R1185 VTAIL.n313 VTAIL.n281 0.155672
R1186 VTAIL.n306 VTAIL.n281 0.155672
R1187 VTAIL.n306 VTAIL.n305 0.155672
R1188 VTAIL.n305 VTAIL.n285 0.155672
R1189 VTAIL.n298 VTAIL.n285 0.155672
R1190 VTAIL.n298 VTAIL.n297 0.155672
R1191 VTAIL.n297 VTAIL.n289 0.155672
R1192 VTAIL VTAIL.n1 0.0586897
R1193 B.n1138 B.n1137 585
R1194 B.n409 B.n185 585
R1195 B.n408 B.n407 585
R1196 B.n406 B.n405 585
R1197 B.n404 B.n403 585
R1198 B.n402 B.n401 585
R1199 B.n400 B.n399 585
R1200 B.n398 B.n397 585
R1201 B.n396 B.n395 585
R1202 B.n394 B.n393 585
R1203 B.n392 B.n391 585
R1204 B.n390 B.n389 585
R1205 B.n388 B.n387 585
R1206 B.n386 B.n385 585
R1207 B.n384 B.n383 585
R1208 B.n382 B.n381 585
R1209 B.n380 B.n379 585
R1210 B.n378 B.n377 585
R1211 B.n376 B.n375 585
R1212 B.n374 B.n373 585
R1213 B.n372 B.n371 585
R1214 B.n370 B.n369 585
R1215 B.n368 B.n367 585
R1216 B.n366 B.n365 585
R1217 B.n364 B.n363 585
R1218 B.n362 B.n361 585
R1219 B.n360 B.n359 585
R1220 B.n358 B.n357 585
R1221 B.n356 B.n355 585
R1222 B.n354 B.n353 585
R1223 B.n352 B.n351 585
R1224 B.n350 B.n349 585
R1225 B.n348 B.n347 585
R1226 B.n346 B.n345 585
R1227 B.n344 B.n343 585
R1228 B.n342 B.n341 585
R1229 B.n340 B.n339 585
R1230 B.n338 B.n337 585
R1231 B.n336 B.n335 585
R1232 B.n334 B.n333 585
R1233 B.n332 B.n331 585
R1234 B.n330 B.n329 585
R1235 B.n328 B.n327 585
R1236 B.n326 B.n325 585
R1237 B.n324 B.n323 585
R1238 B.n322 B.n321 585
R1239 B.n320 B.n319 585
R1240 B.n318 B.n317 585
R1241 B.n316 B.n315 585
R1242 B.n314 B.n313 585
R1243 B.n312 B.n311 585
R1244 B.n309 B.n308 585
R1245 B.n307 B.n306 585
R1246 B.n305 B.n304 585
R1247 B.n303 B.n302 585
R1248 B.n301 B.n300 585
R1249 B.n299 B.n298 585
R1250 B.n297 B.n296 585
R1251 B.n295 B.n294 585
R1252 B.n293 B.n292 585
R1253 B.n291 B.n290 585
R1254 B.n288 B.n287 585
R1255 B.n286 B.n285 585
R1256 B.n284 B.n283 585
R1257 B.n282 B.n281 585
R1258 B.n280 B.n279 585
R1259 B.n278 B.n277 585
R1260 B.n276 B.n275 585
R1261 B.n274 B.n273 585
R1262 B.n272 B.n271 585
R1263 B.n270 B.n269 585
R1264 B.n268 B.n267 585
R1265 B.n266 B.n265 585
R1266 B.n264 B.n263 585
R1267 B.n262 B.n261 585
R1268 B.n260 B.n259 585
R1269 B.n258 B.n257 585
R1270 B.n256 B.n255 585
R1271 B.n254 B.n253 585
R1272 B.n252 B.n251 585
R1273 B.n250 B.n249 585
R1274 B.n248 B.n247 585
R1275 B.n246 B.n245 585
R1276 B.n244 B.n243 585
R1277 B.n242 B.n241 585
R1278 B.n240 B.n239 585
R1279 B.n238 B.n237 585
R1280 B.n236 B.n235 585
R1281 B.n234 B.n233 585
R1282 B.n232 B.n231 585
R1283 B.n230 B.n229 585
R1284 B.n228 B.n227 585
R1285 B.n226 B.n225 585
R1286 B.n224 B.n223 585
R1287 B.n222 B.n221 585
R1288 B.n220 B.n219 585
R1289 B.n218 B.n217 585
R1290 B.n216 B.n215 585
R1291 B.n214 B.n213 585
R1292 B.n212 B.n211 585
R1293 B.n210 B.n209 585
R1294 B.n208 B.n207 585
R1295 B.n206 B.n205 585
R1296 B.n204 B.n203 585
R1297 B.n202 B.n201 585
R1298 B.n200 B.n199 585
R1299 B.n198 B.n197 585
R1300 B.n196 B.n195 585
R1301 B.n194 B.n193 585
R1302 B.n192 B.n191 585
R1303 B.n130 B.n129 585
R1304 B.n1143 B.n1142 585
R1305 B.n1136 B.n186 585
R1306 B.n186 B.n127 585
R1307 B.n1135 B.n126 585
R1308 B.n1147 B.n126 585
R1309 B.n1134 B.n125 585
R1310 B.n1148 B.n125 585
R1311 B.n1133 B.n124 585
R1312 B.n1149 B.n124 585
R1313 B.n1132 B.n1131 585
R1314 B.n1131 B.n120 585
R1315 B.n1130 B.n119 585
R1316 B.n1155 B.n119 585
R1317 B.n1129 B.n118 585
R1318 B.n1156 B.n118 585
R1319 B.n1128 B.n117 585
R1320 B.n1157 B.n117 585
R1321 B.n1127 B.n1126 585
R1322 B.n1126 B.n113 585
R1323 B.n1125 B.n112 585
R1324 B.n1163 B.n112 585
R1325 B.n1124 B.n111 585
R1326 B.n1164 B.n111 585
R1327 B.n1123 B.n110 585
R1328 B.n1165 B.n110 585
R1329 B.n1122 B.n1121 585
R1330 B.n1121 B.n106 585
R1331 B.n1120 B.n105 585
R1332 B.n1171 B.n105 585
R1333 B.n1119 B.n104 585
R1334 B.n1172 B.n104 585
R1335 B.n1118 B.n103 585
R1336 B.n1173 B.n103 585
R1337 B.n1117 B.n1116 585
R1338 B.n1116 B.n99 585
R1339 B.n1115 B.n98 585
R1340 B.n1179 B.n98 585
R1341 B.n1114 B.n97 585
R1342 B.n1180 B.n97 585
R1343 B.n1113 B.n96 585
R1344 B.n1181 B.n96 585
R1345 B.n1112 B.n1111 585
R1346 B.n1111 B.n92 585
R1347 B.n1110 B.n91 585
R1348 B.n1187 B.n91 585
R1349 B.n1109 B.n90 585
R1350 B.n1188 B.n90 585
R1351 B.n1108 B.n89 585
R1352 B.n1189 B.n89 585
R1353 B.n1107 B.n1106 585
R1354 B.n1106 B.n85 585
R1355 B.n1105 B.n84 585
R1356 B.n1195 B.n84 585
R1357 B.n1104 B.n83 585
R1358 B.n1196 B.n83 585
R1359 B.n1103 B.n82 585
R1360 B.n1197 B.n82 585
R1361 B.n1102 B.n1101 585
R1362 B.n1101 B.n78 585
R1363 B.n1100 B.n77 585
R1364 B.n1203 B.n77 585
R1365 B.n1099 B.n76 585
R1366 B.n1204 B.n76 585
R1367 B.n1098 B.n75 585
R1368 B.n1205 B.n75 585
R1369 B.n1097 B.n1096 585
R1370 B.n1096 B.n71 585
R1371 B.n1095 B.n70 585
R1372 B.n1211 B.n70 585
R1373 B.n1094 B.n69 585
R1374 B.n1212 B.n69 585
R1375 B.n1093 B.n68 585
R1376 B.n1213 B.n68 585
R1377 B.n1092 B.n1091 585
R1378 B.n1091 B.n64 585
R1379 B.n1090 B.n63 585
R1380 B.n1219 B.n63 585
R1381 B.n1089 B.n62 585
R1382 B.n1220 B.n62 585
R1383 B.n1088 B.n61 585
R1384 B.n1221 B.n61 585
R1385 B.n1087 B.n1086 585
R1386 B.n1086 B.n57 585
R1387 B.n1085 B.n56 585
R1388 B.n1227 B.n56 585
R1389 B.n1084 B.n55 585
R1390 B.n1228 B.n55 585
R1391 B.n1083 B.n54 585
R1392 B.n1229 B.n54 585
R1393 B.n1082 B.n1081 585
R1394 B.n1081 B.n50 585
R1395 B.n1080 B.n49 585
R1396 B.n1235 B.n49 585
R1397 B.n1079 B.n48 585
R1398 B.n1236 B.n48 585
R1399 B.n1078 B.n47 585
R1400 B.n1237 B.n47 585
R1401 B.n1077 B.n1076 585
R1402 B.n1076 B.n43 585
R1403 B.n1075 B.n42 585
R1404 B.n1243 B.n42 585
R1405 B.n1074 B.n41 585
R1406 B.n1244 B.n41 585
R1407 B.n1073 B.n40 585
R1408 B.n1245 B.n40 585
R1409 B.n1072 B.n1071 585
R1410 B.n1071 B.n36 585
R1411 B.n1070 B.n35 585
R1412 B.n1251 B.n35 585
R1413 B.n1069 B.n34 585
R1414 B.n1252 B.n34 585
R1415 B.n1068 B.n33 585
R1416 B.n1253 B.n33 585
R1417 B.n1067 B.n1066 585
R1418 B.n1066 B.n29 585
R1419 B.n1065 B.n28 585
R1420 B.n1259 B.n28 585
R1421 B.n1064 B.n27 585
R1422 B.n1260 B.n27 585
R1423 B.n1063 B.n26 585
R1424 B.n1261 B.n26 585
R1425 B.n1062 B.n1061 585
R1426 B.n1061 B.n22 585
R1427 B.n1060 B.n21 585
R1428 B.n1267 B.n21 585
R1429 B.n1059 B.n20 585
R1430 B.n1268 B.n20 585
R1431 B.n1058 B.n19 585
R1432 B.n1269 B.n19 585
R1433 B.n1057 B.n1056 585
R1434 B.n1056 B.n15 585
R1435 B.n1055 B.n14 585
R1436 B.n1275 B.n14 585
R1437 B.n1054 B.n13 585
R1438 B.n1276 B.n13 585
R1439 B.n1053 B.n12 585
R1440 B.n1277 B.n12 585
R1441 B.n1052 B.n1051 585
R1442 B.n1051 B.n8 585
R1443 B.n1050 B.n7 585
R1444 B.n1283 B.n7 585
R1445 B.n1049 B.n6 585
R1446 B.n1284 B.n6 585
R1447 B.n1048 B.n5 585
R1448 B.n1285 B.n5 585
R1449 B.n1047 B.n1046 585
R1450 B.n1046 B.n4 585
R1451 B.n1045 B.n410 585
R1452 B.n1045 B.n1044 585
R1453 B.n1035 B.n411 585
R1454 B.n412 B.n411 585
R1455 B.n1037 B.n1036 585
R1456 B.n1038 B.n1037 585
R1457 B.n1034 B.n417 585
R1458 B.n417 B.n416 585
R1459 B.n1033 B.n1032 585
R1460 B.n1032 B.n1031 585
R1461 B.n419 B.n418 585
R1462 B.n420 B.n419 585
R1463 B.n1024 B.n1023 585
R1464 B.n1025 B.n1024 585
R1465 B.n1022 B.n425 585
R1466 B.n425 B.n424 585
R1467 B.n1021 B.n1020 585
R1468 B.n1020 B.n1019 585
R1469 B.n427 B.n426 585
R1470 B.n428 B.n427 585
R1471 B.n1012 B.n1011 585
R1472 B.n1013 B.n1012 585
R1473 B.n1010 B.n433 585
R1474 B.n433 B.n432 585
R1475 B.n1009 B.n1008 585
R1476 B.n1008 B.n1007 585
R1477 B.n435 B.n434 585
R1478 B.n436 B.n435 585
R1479 B.n1000 B.n999 585
R1480 B.n1001 B.n1000 585
R1481 B.n998 B.n441 585
R1482 B.n441 B.n440 585
R1483 B.n997 B.n996 585
R1484 B.n996 B.n995 585
R1485 B.n443 B.n442 585
R1486 B.n444 B.n443 585
R1487 B.n988 B.n987 585
R1488 B.n989 B.n988 585
R1489 B.n986 B.n448 585
R1490 B.n452 B.n448 585
R1491 B.n985 B.n984 585
R1492 B.n984 B.n983 585
R1493 B.n450 B.n449 585
R1494 B.n451 B.n450 585
R1495 B.n976 B.n975 585
R1496 B.n977 B.n976 585
R1497 B.n974 B.n457 585
R1498 B.n457 B.n456 585
R1499 B.n973 B.n972 585
R1500 B.n972 B.n971 585
R1501 B.n459 B.n458 585
R1502 B.n460 B.n459 585
R1503 B.n964 B.n963 585
R1504 B.n965 B.n964 585
R1505 B.n962 B.n465 585
R1506 B.n465 B.n464 585
R1507 B.n961 B.n960 585
R1508 B.n960 B.n959 585
R1509 B.n467 B.n466 585
R1510 B.n468 B.n467 585
R1511 B.n952 B.n951 585
R1512 B.n953 B.n952 585
R1513 B.n950 B.n473 585
R1514 B.n473 B.n472 585
R1515 B.n949 B.n948 585
R1516 B.n948 B.n947 585
R1517 B.n475 B.n474 585
R1518 B.n476 B.n475 585
R1519 B.n940 B.n939 585
R1520 B.n941 B.n940 585
R1521 B.n938 B.n481 585
R1522 B.n481 B.n480 585
R1523 B.n937 B.n936 585
R1524 B.n936 B.n935 585
R1525 B.n483 B.n482 585
R1526 B.n484 B.n483 585
R1527 B.n928 B.n927 585
R1528 B.n929 B.n928 585
R1529 B.n926 B.n489 585
R1530 B.n489 B.n488 585
R1531 B.n925 B.n924 585
R1532 B.n924 B.n923 585
R1533 B.n491 B.n490 585
R1534 B.n492 B.n491 585
R1535 B.n916 B.n915 585
R1536 B.n917 B.n916 585
R1537 B.n914 B.n497 585
R1538 B.n497 B.n496 585
R1539 B.n913 B.n912 585
R1540 B.n912 B.n911 585
R1541 B.n499 B.n498 585
R1542 B.n500 B.n499 585
R1543 B.n904 B.n903 585
R1544 B.n905 B.n904 585
R1545 B.n902 B.n505 585
R1546 B.n505 B.n504 585
R1547 B.n901 B.n900 585
R1548 B.n900 B.n899 585
R1549 B.n507 B.n506 585
R1550 B.n508 B.n507 585
R1551 B.n892 B.n891 585
R1552 B.n893 B.n892 585
R1553 B.n890 B.n513 585
R1554 B.n513 B.n512 585
R1555 B.n889 B.n888 585
R1556 B.n888 B.n887 585
R1557 B.n515 B.n514 585
R1558 B.n516 B.n515 585
R1559 B.n880 B.n879 585
R1560 B.n881 B.n880 585
R1561 B.n878 B.n521 585
R1562 B.n521 B.n520 585
R1563 B.n877 B.n876 585
R1564 B.n876 B.n875 585
R1565 B.n523 B.n522 585
R1566 B.n524 B.n523 585
R1567 B.n868 B.n867 585
R1568 B.n869 B.n868 585
R1569 B.n866 B.n529 585
R1570 B.n529 B.n528 585
R1571 B.n865 B.n864 585
R1572 B.n864 B.n863 585
R1573 B.n531 B.n530 585
R1574 B.n532 B.n531 585
R1575 B.n856 B.n855 585
R1576 B.n857 B.n856 585
R1577 B.n854 B.n537 585
R1578 B.n537 B.n536 585
R1579 B.n853 B.n852 585
R1580 B.n852 B.n851 585
R1581 B.n539 B.n538 585
R1582 B.n540 B.n539 585
R1583 B.n844 B.n843 585
R1584 B.n845 B.n844 585
R1585 B.n842 B.n545 585
R1586 B.n545 B.n544 585
R1587 B.n841 B.n840 585
R1588 B.n840 B.n839 585
R1589 B.n547 B.n546 585
R1590 B.n548 B.n547 585
R1591 B.n835 B.n834 585
R1592 B.n551 B.n550 585
R1593 B.n831 B.n830 585
R1594 B.n832 B.n831 585
R1595 B.n829 B.n607 585
R1596 B.n828 B.n827 585
R1597 B.n826 B.n825 585
R1598 B.n824 B.n823 585
R1599 B.n822 B.n821 585
R1600 B.n820 B.n819 585
R1601 B.n818 B.n817 585
R1602 B.n816 B.n815 585
R1603 B.n814 B.n813 585
R1604 B.n812 B.n811 585
R1605 B.n810 B.n809 585
R1606 B.n808 B.n807 585
R1607 B.n806 B.n805 585
R1608 B.n804 B.n803 585
R1609 B.n802 B.n801 585
R1610 B.n800 B.n799 585
R1611 B.n798 B.n797 585
R1612 B.n796 B.n795 585
R1613 B.n794 B.n793 585
R1614 B.n792 B.n791 585
R1615 B.n790 B.n789 585
R1616 B.n788 B.n787 585
R1617 B.n786 B.n785 585
R1618 B.n784 B.n783 585
R1619 B.n782 B.n781 585
R1620 B.n780 B.n779 585
R1621 B.n778 B.n777 585
R1622 B.n776 B.n775 585
R1623 B.n774 B.n773 585
R1624 B.n772 B.n771 585
R1625 B.n770 B.n769 585
R1626 B.n768 B.n767 585
R1627 B.n766 B.n765 585
R1628 B.n764 B.n763 585
R1629 B.n762 B.n761 585
R1630 B.n760 B.n759 585
R1631 B.n758 B.n757 585
R1632 B.n756 B.n755 585
R1633 B.n754 B.n753 585
R1634 B.n752 B.n751 585
R1635 B.n750 B.n749 585
R1636 B.n748 B.n747 585
R1637 B.n746 B.n745 585
R1638 B.n744 B.n743 585
R1639 B.n742 B.n741 585
R1640 B.n740 B.n739 585
R1641 B.n738 B.n737 585
R1642 B.n736 B.n735 585
R1643 B.n734 B.n733 585
R1644 B.n732 B.n731 585
R1645 B.n730 B.n729 585
R1646 B.n728 B.n727 585
R1647 B.n726 B.n725 585
R1648 B.n724 B.n723 585
R1649 B.n722 B.n721 585
R1650 B.n720 B.n719 585
R1651 B.n718 B.n717 585
R1652 B.n716 B.n715 585
R1653 B.n714 B.n713 585
R1654 B.n712 B.n711 585
R1655 B.n710 B.n709 585
R1656 B.n708 B.n707 585
R1657 B.n706 B.n705 585
R1658 B.n704 B.n703 585
R1659 B.n702 B.n701 585
R1660 B.n700 B.n699 585
R1661 B.n698 B.n697 585
R1662 B.n696 B.n695 585
R1663 B.n694 B.n693 585
R1664 B.n692 B.n691 585
R1665 B.n690 B.n689 585
R1666 B.n688 B.n687 585
R1667 B.n686 B.n685 585
R1668 B.n684 B.n683 585
R1669 B.n682 B.n681 585
R1670 B.n680 B.n679 585
R1671 B.n678 B.n677 585
R1672 B.n676 B.n675 585
R1673 B.n674 B.n673 585
R1674 B.n672 B.n671 585
R1675 B.n670 B.n669 585
R1676 B.n668 B.n667 585
R1677 B.n666 B.n665 585
R1678 B.n664 B.n663 585
R1679 B.n662 B.n661 585
R1680 B.n660 B.n659 585
R1681 B.n658 B.n657 585
R1682 B.n656 B.n655 585
R1683 B.n654 B.n653 585
R1684 B.n652 B.n651 585
R1685 B.n650 B.n649 585
R1686 B.n648 B.n647 585
R1687 B.n646 B.n645 585
R1688 B.n644 B.n643 585
R1689 B.n642 B.n641 585
R1690 B.n640 B.n639 585
R1691 B.n638 B.n637 585
R1692 B.n636 B.n635 585
R1693 B.n634 B.n633 585
R1694 B.n632 B.n631 585
R1695 B.n630 B.n629 585
R1696 B.n628 B.n627 585
R1697 B.n626 B.n625 585
R1698 B.n624 B.n623 585
R1699 B.n622 B.n621 585
R1700 B.n620 B.n619 585
R1701 B.n618 B.n617 585
R1702 B.n616 B.n615 585
R1703 B.n614 B.n606 585
R1704 B.n832 B.n606 585
R1705 B.n836 B.n549 585
R1706 B.n549 B.n548 585
R1707 B.n838 B.n837 585
R1708 B.n839 B.n838 585
R1709 B.n543 B.n542 585
R1710 B.n544 B.n543 585
R1711 B.n847 B.n846 585
R1712 B.n846 B.n845 585
R1713 B.n848 B.n541 585
R1714 B.n541 B.n540 585
R1715 B.n850 B.n849 585
R1716 B.n851 B.n850 585
R1717 B.n535 B.n534 585
R1718 B.n536 B.n535 585
R1719 B.n859 B.n858 585
R1720 B.n858 B.n857 585
R1721 B.n860 B.n533 585
R1722 B.n533 B.n532 585
R1723 B.n862 B.n861 585
R1724 B.n863 B.n862 585
R1725 B.n527 B.n526 585
R1726 B.n528 B.n527 585
R1727 B.n871 B.n870 585
R1728 B.n870 B.n869 585
R1729 B.n872 B.n525 585
R1730 B.n525 B.n524 585
R1731 B.n874 B.n873 585
R1732 B.n875 B.n874 585
R1733 B.n519 B.n518 585
R1734 B.n520 B.n519 585
R1735 B.n883 B.n882 585
R1736 B.n882 B.n881 585
R1737 B.n884 B.n517 585
R1738 B.n517 B.n516 585
R1739 B.n886 B.n885 585
R1740 B.n887 B.n886 585
R1741 B.n511 B.n510 585
R1742 B.n512 B.n511 585
R1743 B.n895 B.n894 585
R1744 B.n894 B.n893 585
R1745 B.n896 B.n509 585
R1746 B.n509 B.n508 585
R1747 B.n898 B.n897 585
R1748 B.n899 B.n898 585
R1749 B.n503 B.n502 585
R1750 B.n504 B.n503 585
R1751 B.n907 B.n906 585
R1752 B.n906 B.n905 585
R1753 B.n908 B.n501 585
R1754 B.n501 B.n500 585
R1755 B.n910 B.n909 585
R1756 B.n911 B.n910 585
R1757 B.n495 B.n494 585
R1758 B.n496 B.n495 585
R1759 B.n919 B.n918 585
R1760 B.n918 B.n917 585
R1761 B.n920 B.n493 585
R1762 B.n493 B.n492 585
R1763 B.n922 B.n921 585
R1764 B.n923 B.n922 585
R1765 B.n487 B.n486 585
R1766 B.n488 B.n487 585
R1767 B.n931 B.n930 585
R1768 B.n930 B.n929 585
R1769 B.n932 B.n485 585
R1770 B.n485 B.n484 585
R1771 B.n934 B.n933 585
R1772 B.n935 B.n934 585
R1773 B.n479 B.n478 585
R1774 B.n480 B.n479 585
R1775 B.n943 B.n942 585
R1776 B.n942 B.n941 585
R1777 B.n944 B.n477 585
R1778 B.n477 B.n476 585
R1779 B.n946 B.n945 585
R1780 B.n947 B.n946 585
R1781 B.n471 B.n470 585
R1782 B.n472 B.n471 585
R1783 B.n955 B.n954 585
R1784 B.n954 B.n953 585
R1785 B.n956 B.n469 585
R1786 B.n469 B.n468 585
R1787 B.n958 B.n957 585
R1788 B.n959 B.n958 585
R1789 B.n463 B.n462 585
R1790 B.n464 B.n463 585
R1791 B.n967 B.n966 585
R1792 B.n966 B.n965 585
R1793 B.n968 B.n461 585
R1794 B.n461 B.n460 585
R1795 B.n970 B.n969 585
R1796 B.n971 B.n970 585
R1797 B.n455 B.n454 585
R1798 B.n456 B.n455 585
R1799 B.n979 B.n978 585
R1800 B.n978 B.n977 585
R1801 B.n980 B.n453 585
R1802 B.n453 B.n451 585
R1803 B.n982 B.n981 585
R1804 B.n983 B.n982 585
R1805 B.n447 B.n446 585
R1806 B.n452 B.n447 585
R1807 B.n991 B.n990 585
R1808 B.n990 B.n989 585
R1809 B.n992 B.n445 585
R1810 B.n445 B.n444 585
R1811 B.n994 B.n993 585
R1812 B.n995 B.n994 585
R1813 B.n439 B.n438 585
R1814 B.n440 B.n439 585
R1815 B.n1003 B.n1002 585
R1816 B.n1002 B.n1001 585
R1817 B.n1004 B.n437 585
R1818 B.n437 B.n436 585
R1819 B.n1006 B.n1005 585
R1820 B.n1007 B.n1006 585
R1821 B.n431 B.n430 585
R1822 B.n432 B.n431 585
R1823 B.n1015 B.n1014 585
R1824 B.n1014 B.n1013 585
R1825 B.n1016 B.n429 585
R1826 B.n429 B.n428 585
R1827 B.n1018 B.n1017 585
R1828 B.n1019 B.n1018 585
R1829 B.n423 B.n422 585
R1830 B.n424 B.n423 585
R1831 B.n1027 B.n1026 585
R1832 B.n1026 B.n1025 585
R1833 B.n1028 B.n421 585
R1834 B.n421 B.n420 585
R1835 B.n1030 B.n1029 585
R1836 B.n1031 B.n1030 585
R1837 B.n415 B.n414 585
R1838 B.n416 B.n415 585
R1839 B.n1040 B.n1039 585
R1840 B.n1039 B.n1038 585
R1841 B.n1041 B.n413 585
R1842 B.n413 B.n412 585
R1843 B.n1043 B.n1042 585
R1844 B.n1044 B.n1043 585
R1845 B.n2 B.n0 585
R1846 B.n4 B.n2 585
R1847 B.n3 B.n1 585
R1848 B.n1284 B.n3 585
R1849 B.n1282 B.n1281 585
R1850 B.n1283 B.n1282 585
R1851 B.n1280 B.n9 585
R1852 B.n9 B.n8 585
R1853 B.n1279 B.n1278 585
R1854 B.n1278 B.n1277 585
R1855 B.n11 B.n10 585
R1856 B.n1276 B.n11 585
R1857 B.n1274 B.n1273 585
R1858 B.n1275 B.n1274 585
R1859 B.n1272 B.n16 585
R1860 B.n16 B.n15 585
R1861 B.n1271 B.n1270 585
R1862 B.n1270 B.n1269 585
R1863 B.n18 B.n17 585
R1864 B.n1268 B.n18 585
R1865 B.n1266 B.n1265 585
R1866 B.n1267 B.n1266 585
R1867 B.n1264 B.n23 585
R1868 B.n23 B.n22 585
R1869 B.n1263 B.n1262 585
R1870 B.n1262 B.n1261 585
R1871 B.n25 B.n24 585
R1872 B.n1260 B.n25 585
R1873 B.n1258 B.n1257 585
R1874 B.n1259 B.n1258 585
R1875 B.n1256 B.n30 585
R1876 B.n30 B.n29 585
R1877 B.n1255 B.n1254 585
R1878 B.n1254 B.n1253 585
R1879 B.n32 B.n31 585
R1880 B.n1252 B.n32 585
R1881 B.n1250 B.n1249 585
R1882 B.n1251 B.n1250 585
R1883 B.n1248 B.n37 585
R1884 B.n37 B.n36 585
R1885 B.n1247 B.n1246 585
R1886 B.n1246 B.n1245 585
R1887 B.n39 B.n38 585
R1888 B.n1244 B.n39 585
R1889 B.n1242 B.n1241 585
R1890 B.n1243 B.n1242 585
R1891 B.n1240 B.n44 585
R1892 B.n44 B.n43 585
R1893 B.n1239 B.n1238 585
R1894 B.n1238 B.n1237 585
R1895 B.n46 B.n45 585
R1896 B.n1236 B.n46 585
R1897 B.n1234 B.n1233 585
R1898 B.n1235 B.n1234 585
R1899 B.n1232 B.n51 585
R1900 B.n51 B.n50 585
R1901 B.n1231 B.n1230 585
R1902 B.n1230 B.n1229 585
R1903 B.n53 B.n52 585
R1904 B.n1228 B.n53 585
R1905 B.n1226 B.n1225 585
R1906 B.n1227 B.n1226 585
R1907 B.n1224 B.n58 585
R1908 B.n58 B.n57 585
R1909 B.n1223 B.n1222 585
R1910 B.n1222 B.n1221 585
R1911 B.n60 B.n59 585
R1912 B.n1220 B.n60 585
R1913 B.n1218 B.n1217 585
R1914 B.n1219 B.n1218 585
R1915 B.n1216 B.n65 585
R1916 B.n65 B.n64 585
R1917 B.n1215 B.n1214 585
R1918 B.n1214 B.n1213 585
R1919 B.n67 B.n66 585
R1920 B.n1212 B.n67 585
R1921 B.n1210 B.n1209 585
R1922 B.n1211 B.n1210 585
R1923 B.n1208 B.n72 585
R1924 B.n72 B.n71 585
R1925 B.n1207 B.n1206 585
R1926 B.n1206 B.n1205 585
R1927 B.n74 B.n73 585
R1928 B.n1204 B.n74 585
R1929 B.n1202 B.n1201 585
R1930 B.n1203 B.n1202 585
R1931 B.n1200 B.n79 585
R1932 B.n79 B.n78 585
R1933 B.n1199 B.n1198 585
R1934 B.n1198 B.n1197 585
R1935 B.n81 B.n80 585
R1936 B.n1196 B.n81 585
R1937 B.n1194 B.n1193 585
R1938 B.n1195 B.n1194 585
R1939 B.n1192 B.n86 585
R1940 B.n86 B.n85 585
R1941 B.n1191 B.n1190 585
R1942 B.n1190 B.n1189 585
R1943 B.n88 B.n87 585
R1944 B.n1188 B.n88 585
R1945 B.n1186 B.n1185 585
R1946 B.n1187 B.n1186 585
R1947 B.n1184 B.n93 585
R1948 B.n93 B.n92 585
R1949 B.n1183 B.n1182 585
R1950 B.n1182 B.n1181 585
R1951 B.n95 B.n94 585
R1952 B.n1180 B.n95 585
R1953 B.n1178 B.n1177 585
R1954 B.n1179 B.n1178 585
R1955 B.n1176 B.n100 585
R1956 B.n100 B.n99 585
R1957 B.n1175 B.n1174 585
R1958 B.n1174 B.n1173 585
R1959 B.n102 B.n101 585
R1960 B.n1172 B.n102 585
R1961 B.n1170 B.n1169 585
R1962 B.n1171 B.n1170 585
R1963 B.n1168 B.n107 585
R1964 B.n107 B.n106 585
R1965 B.n1167 B.n1166 585
R1966 B.n1166 B.n1165 585
R1967 B.n109 B.n108 585
R1968 B.n1164 B.n109 585
R1969 B.n1162 B.n1161 585
R1970 B.n1163 B.n1162 585
R1971 B.n1160 B.n114 585
R1972 B.n114 B.n113 585
R1973 B.n1159 B.n1158 585
R1974 B.n1158 B.n1157 585
R1975 B.n116 B.n115 585
R1976 B.n1156 B.n116 585
R1977 B.n1154 B.n1153 585
R1978 B.n1155 B.n1154 585
R1979 B.n1152 B.n121 585
R1980 B.n121 B.n120 585
R1981 B.n1151 B.n1150 585
R1982 B.n1150 B.n1149 585
R1983 B.n123 B.n122 585
R1984 B.n1148 B.n123 585
R1985 B.n1146 B.n1145 585
R1986 B.n1147 B.n1146 585
R1987 B.n1144 B.n128 585
R1988 B.n128 B.n127 585
R1989 B.n1287 B.n1286 585
R1990 B.n1286 B.n1285 585
R1991 B.n834 B.n549 550.159
R1992 B.n1142 B.n128 550.159
R1993 B.n606 B.n547 550.159
R1994 B.n1138 B.n186 550.159
R1995 B.n611 B.t13 422.606
R1996 B.n608 B.t10 422.606
R1997 B.n189 B.t19 422.606
R1998 B.n187 B.t16 422.606
R1999 B.n612 B.t12 339.601
R2000 B.n188 B.t17 339.601
R2001 B.n609 B.t9 339.601
R2002 B.n190 B.t20 339.601
R2003 B.n611 B.t11 303.111
R2004 B.n608 B.t7 303.111
R2005 B.n189 B.t18 303.111
R2006 B.n187 B.t14 303.111
R2007 B.n1140 B.n1139 256.663
R2008 B.n1140 B.n184 256.663
R2009 B.n1140 B.n183 256.663
R2010 B.n1140 B.n182 256.663
R2011 B.n1140 B.n181 256.663
R2012 B.n1140 B.n180 256.663
R2013 B.n1140 B.n179 256.663
R2014 B.n1140 B.n178 256.663
R2015 B.n1140 B.n177 256.663
R2016 B.n1140 B.n176 256.663
R2017 B.n1140 B.n175 256.663
R2018 B.n1140 B.n174 256.663
R2019 B.n1140 B.n173 256.663
R2020 B.n1140 B.n172 256.663
R2021 B.n1140 B.n171 256.663
R2022 B.n1140 B.n170 256.663
R2023 B.n1140 B.n169 256.663
R2024 B.n1140 B.n168 256.663
R2025 B.n1140 B.n167 256.663
R2026 B.n1140 B.n166 256.663
R2027 B.n1140 B.n165 256.663
R2028 B.n1140 B.n164 256.663
R2029 B.n1140 B.n163 256.663
R2030 B.n1140 B.n162 256.663
R2031 B.n1140 B.n161 256.663
R2032 B.n1140 B.n160 256.663
R2033 B.n1140 B.n159 256.663
R2034 B.n1140 B.n158 256.663
R2035 B.n1140 B.n157 256.663
R2036 B.n1140 B.n156 256.663
R2037 B.n1140 B.n155 256.663
R2038 B.n1140 B.n154 256.663
R2039 B.n1140 B.n153 256.663
R2040 B.n1140 B.n152 256.663
R2041 B.n1140 B.n151 256.663
R2042 B.n1140 B.n150 256.663
R2043 B.n1140 B.n149 256.663
R2044 B.n1140 B.n148 256.663
R2045 B.n1140 B.n147 256.663
R2046 B.n1140 B.n146 256.663
R2047 B.n1140 B.n145 256.663
R2048 B.n1140 B.n144 256.663
R2049 B.n1140 B.n143 256.663
R2050 B.n1140 B.n142 256.663
R2051 B.n1140 B.n141 256.663
R2052 B.n1140 B.n140 256.663
R2053 B.n1140 B.n139 256.663
R2054 B.n1140 B.n138 256.663
R2055 B.n1140 B.n137 256.663
R2056 B.n1140 B.n136 256.663
R2057 B.n1140 B.n135 256.663
R2058 B.n1140 B.n134 256.663
R2059 B.n1140 B.n133 256.663
R2060 B.n1140 B.n132 256.663
R2061 B.n1140 B.n131 256.663
R2062 B.n1141 B.n1140 256.663
R2063 B.n833 B.n832 256.663
R2064 B.n832 B.n552 256.663
R2065 B.n832 B.n553 256.663
R2066 B.n832 B.n554 256.663
R2067 B.n832 B.n555 256.663
R2068 B.n832 B.n556 256.663
R2069 B.n832 B.n557 256.663
R2070 B.n832 B.n558 256.663
R2071 B.n832 B.n559 256.663
R2072 B.n832 B.n560 256.663
R2073 B.n832 B.n561 256.663
R2074 B.n832 B.n562 256.663
R2075 B.n832 B.n563 256.663
R2076 B.n832 B.n564 256.663
R2077 B.n832 B.n565 256.663
R2078 B.n832 B.n566 256.663
R2079 B.n832 B.n567 256.663
R2080 B.n832 B.n568 256.663
R2081 B.n832 B.n569 256.663
R2082 B.n832 B.n570 256.663
R2083 B.n832 B.n571 256.663
R2084 B.n832 B.n572 256.663
R2085 B.n832 B.n573 256.663
R2086 B.n832 B.n574 256.663
R2087 B.n832 B.n575 256.663
R2088 B.n832 B.n576 256.663
R2089 B.n832 B.n577 256.663
R2090 B.n832 B.n578 256.663
R2091 B.n832 B.n579 256.663
R2092 B.n832 B.n580 256.663
R2093 B.n832 B.n581 256.663
R2094 B.n832 B.n582 256.663
R2095 B.n832 B.n583 256.663
R2096 B.n832 B.n584 256.663
R2097 B.n832 B.n585 256.663
R2098 B.n832 B.n586 256.663
R2099 B.n832 B.n587 256.663
R2100 B.n832 B.n588 256.663
R2101 B.n832 B.n589 256.663
R2102 B.n832 B.n590 256.663
R2103 B.n832 B.n591 256.663
R2104 B.n832 B.n592 256.663
R2105 B.n832 B.n593 256.663
R2106 B.n832 B.n594 256.663
R2107 B.n832 B.n595 256.663
R2108 B.n832 B.n596 256.663
R2109 B.n832 B.n597 256.663
R2110 B.n832 B.n598 256.663
R2111 B.n832 B.n599 256.663
R2112 B.n832 B.n600 256.663
R2113 B.n832 B.n601 256.663
R2114 B.n832 B.n602 256.663
R2115 B.n832 B.n603 256.663
R2116 B.n832 B.n604 256.663
R2117 B.n832 B.n605 256.663
R2118 B.n838 B.n549 163.367
R2119 B.n838 B.n543 163.367
R2120 B.n846 B.n543 163.367
R2121 B.n846 B.n541 163.367
R2122 B.n850 B.n541 163.367
R2123 B.n850 B.n535 163.367
R2124 B.n858 B.n535 163.367
R2125 B.n858 B.n533 163.367
R2126 B.n862 B.n533 163.367
R2127 B.n862 B.n527 163.367
R2128 B.n870 B.n527 163.367
R2129 B.n870 B.n525 163.367
R2130 B.n874 B.n525 163.367
R2131 B.n874 B.n519 163.367
R2132 B.n882 B.n519 163.367
R2133 B.n882 B.n517 163.367
R2134 B.n886 B.n517 163.367
R2135 B.n886 B.n511 163.367
R2136 B.n894 B.n511 163.367
R2137 B.n894 B.n509 163.367
R2138 B.n898 B.n509 163.367
R2139 B.n898 B.n503 163.367
R2140 B.n906 B.n503 163.367
R2141 B.n906 B.n501 163.367
R2142 B.n910 B.n501 163.367
R2143 B.n910 B.n495 163.367
R2144 B.n918 B.n495 163.367
R2145 B.n918 B.n493 163.367
R2146 B.n922 B.n493 163.367
R2147 B.n922 B.n487 163.367
R2148 B.n930 B.n487 163.367
R2149 B.n930 B.n485 163.367
R2150 B.n934 B.n485 163.367
R2151 B.n934 B.n479 163.367
R2152 B.n942 B.n479 163.367
R2153 B.n942 B.n477 163.367
R2154 B.n946 B.n477 163.367
R2155 B.n946 B.n471 163.367
R2156 B.n954 B.n471 163.367
R2157 B.n954 B.n469 163.367
R2158 B.n958 B.n469 163.367
R2159 B.n958 B.n463 163.367
R2160 B.n966 B.n463 163.367
R2161 B.n966 B.n461 163.367
R2162 B.n970 B.n461 163.367
R2163 B.n970 B.n455 163.367
R2164 B.n978 B.n455 163.367
R2165 B.n978 B.n453 163.367
R2166 B.n982 B.n453 163.367
R2167 B.n982 B.n447 163.367
R2168 B.n990 B.n447 163.367
R2169 B.n990 B.n445 163.367
R2170 B.n994 B.n445 163.367
R2171 B.n994 B.n439 163.367
R2172 B.n1002 B.n439 163.367
R2173 B.n1002 B.n437 163.367
R2174 B.n1006 B.n437 163.367
R2175 B.n1006 B.n431 163.367
R2176 B.n1014 B.n431 163.367
R2177 B.n1014 B.n429 163.367
R2178 B.n1018 B.n429 163.367
R2179 B.n1018 B.n423 163.367
R2180 B.n1026 B.n423 163.367
R2181 B.n1026 B.n421 163.367
R2182 B.n1030 B.n421 163.367
R2183 B.n1030 B.n415 163.367
R2184 B.n1039 B.n415 163.367
R2185 B.n1039 B.n413 163.367
R2186 B.n1043 B.n413 163.367
R2187 B.n1043 B.n2 163.367
R2188 B.n1286 B.n2 163.367
R2189 B.n1286 B.n3 163.367
R2190 B.n1282 B.n3 163.367
R2191 B.n1282 B.n9 163.367
R2192 B.n1278 B.n9 163.367
R2193 B.n1278 B.n11 163.367
R2194 B.n1274 B.n11 163.367
R2195 B.n1274 B.n16 163.367
R2196 B.n1270 B.n16 163.367
R2197 B.n1270 B.n18 163.367
R2198 B.n1266 B.n18 163.367
R2199 B.n1266 B.n23 163.367
R2200 B.n1262 B.n23 163.367
R2201 B.n1262 B.n25 163.367
R2202 B.n1258 B.n25 163.367
R2203 B.n1258 B.n30 163.367
R2204 B.n1254 B.n30 163.367
R2205 B.n1254 B.n32 163.367
R2206 B.n1250 B.n32 163.367
R2207 B.n1250 B.n37 163.367
R2208 B.n1246 B.n37 163.367
R2209 B.n1246 B.n39 163.367
R2210 B.n1242 B.n39 163.367
R2211 B.n1242 B.n44 163.367
R2212 B.n1238 B.n44 163.367
R2213 B.n1238 B.n46 163.367
R2214 B.n1234 B.n46 163.367
R2215 B.n1234 B.n51 163.367
R2216 B.n1230 B.n51 163.367
R2217 B.n1230 B.n53 163.367
R2218 B.n1226 B.n53 163.367
R2219 B.n1226 B.n58 163.367
R2220 B.n1222 B.n58 163.367
R2221 B.n1222 B.n60 163.367
R2222 B.n1218 B.n60 163.367
R2223 B.n1218 B.n65 163.367
R2224 B.n1214 B.n65 163.367
R2225 B.n1214 B.n67 163.367
R2226 B.n1210 B.n67 163.367
R2227 B.n1210 B.n72 163.367
R2228 B.n1206 B.n72 163.367
R2229 B.n1206 B.n74 163.367
R2230 B.n1202 B.n74 163.367
R2231 B.n1202 B.n79 163.367
R2232 B.n1198 B.n79 163.367
R2233 B.n1198 B.n81 163.367
R2234 B.n1194 B.n81 163.367
R2235 B.n1194 B.n86 163.367
R2236 B.n1190 B.n86 163.367
R2237 B.n1190 B.n88 163.367
R2238 B.n1186 B.n88 163.367
R2239 B.n1186 B.n93 163.367
R2240 B.n1182 B.n93 163.367
R2241 B.n1182 B.n95 163.367
R2242 B.n1178 B.n95 163.367
R2243 B.n1178 B.n100 163.367
R2244 B.n1174 B.n100 163.367
R2245 B.n1174 B.n102 163.367
R2246 B.n1170 B.n102 163.367
R2247 B.n1170 B.n107 163.367
R2248 B.n1166 B.n107 163.367
R2249 B.n1166 B.n109 163.367
R2250 B.n1162 B.n109 163.367
R2251 B.n1162 B.n114 163.367
R2252 B.n1158 B.n114 163.367
R2253 B.n1158 B.n116 163.367
R2254 B.n1154 B.n116 163.367
R2255 B.n1154 B.n121 163.367
R2256 B.n1150 B.n121 163.367
R2257 B.n1150 B.n123 163.367
R2258 B.n1146 B.n123 163.367
R2259 B.n1146 B.n128 163.367
R2260 B.n831 B.n551 163.367
R2261 B.n831 B.n607 163.367
R2262 B.n827 B.n826 163.367
R2263 B.n823 B.n822 163.367
R2264 B.n819 B.n818 163.367
R2265 B.n815 B.n814 163.367
R2266 B.n811 B.n810 163.367
R2267 B.n807 B.n806 163.367
R2268 B.n803 B.n802 163.367
R2269 B.n799 B.n798 163.367
R2270 B.n795 B.n794 163.367
R2271 B.n791 B.n790 163.367
R2272 B.n787 B.n786 163.367
R2273 B.n783 B.n782 163.367
R2274 B.n779 B.n778 163.367
R2275 B.n775 B.n774 163.367
R2276 B.n771 B.n770 163.367
R2277 B.n767 B.n766 163.367
R2278 B.n763 B.n762 163.367
R2279 B.n759 B.n758 163.367
R2280 B.n755 B.n754 163.367
R2281 B.n751 B.n750 163.367
R2282 B.n747 B.n746 163.367
R2283 B.n743 B.n742 163.367
R2284 B.n739 B.n738 163.367
R2285 B.n735 B.n734 163.367
R2286 B.n731 B.n730 163.367
R2287 B.n727 B.n726 163.367
R2288 B.n723 B.n722 163.367
R2289 B.n719 B.n718 163.367
R2290 B.n715 B.n714 163.367
R2291 B.n711 B.n710 163.367
R2292 B.n707 B.n706 163.367
R2293 B.n703 B.n702 163.367
R2294 B.n699 B.n698 163.367
R2295 B.n695 B.n694 163.367
R2296 B.n691 B.n690 163.367
R2297 B.n687 B.n686 163.367
R2298 B.n683 B.n682 163.367
R2299 B.n679 B.n678 163.367
R2300 B.n675 B.n674 163.367
R2301 B.n671 B.n670 163.367
R2302 B.n667 B.n666 163.367
R2303 B.n663 B.n662 163.367
R2304 B.n659 B.n658 163.367
R2305 B.n655 B.n654 163.367
R2306 B.n651 B.n650 163.367
R2307 B.n647 B.n646 163.367
R2308 B.n643 B.n642 163.367
R2309 B.n639 B.n638 163.367
R2310 B.n635 B.n634 163.367
R2311 B.n631 B.n630 163.367
R2312 B.n627 B.n626 163.367
R2313 B.n623 B.n622 163.367
R2314 B.n619 B.n618 163.367
R2315 B.n615 B.n606 163.367
R2316 B.n840 B.n547 163.367
R2317 B.n840 B.n545 163.367
R2318 B.n844 B.n545 163.367
R2319 B.n844 B.n539 163.367
R2320 B.n852 B.n539 163.367
R2321 B.n852 B.n537 163.367
R2322 B.n856 B.n537 163.367
R2323 B.n856 B.n531 163.367
R2324 B.n864 B.n531 163.367
R2325 B.n864 B.n529 163.367
R2326 B.n868 B.n529 163.367
R2327 B.n868 B.n523 163.367
R2328 B.n876 B.n523 163.367
R2329 B.n876 B.n521 163.367
R2330 B.n880 B.n521 163.367
R2331 B.n880 B.n515 163.367
R2332 B.n888 B.n515 163.367
R2333 B.n888 B.n513 163.367
R2334 B.n892 B.n513 163.367
R2335 B.n892 B.n507 163.367
R2336 B.n900 B.n507 163.367
R2337 B.n900 B.n505 163.367
R2338 B.n904 B.n505 163.367
R2339 B.n904 B.n499 163.367
R2340 B.n912 B.n499 163.367
R2341 B.n912 B.n497 163.367
R2342 B.n916 B.n497 163.367
R2343 B.n916 B.n491 163.367
R2344 B.n924 B.n491 163.367
R2345 B.n924 B.n489 163.367
R2346 B.n928 B.n489 163.367
R2347 B.n928 B.n483 163.367
R2348 B.n936 B.n483 163.367
R2349 B.n936 B.n481 163.367
R2350 B.n940 B.n481 163.367
R2351 B.n940 B.n475 163.367
R2352 B.n948 B.n475 163.367
R2353 B.n948 B.n473 163.367
R2354 B.n952 B.n473 163.367
R2355 B.n952 B.n467 163.367
R2356 B.n960 B.n467 163.367
R2357 B.n960 B.n465 163.367
R2358 B.n964 B.n465 163.367
R2359 B.n964 B.n459 163.367
R2360 B.n972 B.n459 163.367
R2361 B.n972 B.n457 163.367
R2362 B.n976 B.n457 163.367
R2363 B.n976 B.n450 163.367
R2364 B.n984 B.n450 163.367
R2365 B.n984 B.n448 163.367
R2366 B.n988 B.n448 163.367
R2367 B.n988 B.n443 163.367
R2368 B.n996 B.n443 163.367
R2369 B.n996 B.n441 163.367
R2370 B.n1000 B.n441 163.367
R2371 B.n1000 B.n435 163.367
R2372 B.n1008 B.n435 163.367
R2373 B.n1008 B.n433 163.367
R2374 B.n1012 B.n433 163.367
R2375 B.n1012 B.n427 163.367
R2376 B.n1020 B.n427 163.367
R2377 B.n1020 B.n425 163.367
R2378 B.n1024 B.n425 163.367
R2379 B.n1024 B.n419 163.367
R2380 B.n1032 B.n419 163.367
R2381 B.n1032 B.n417 163.367
R2382 B.n1037 B.n417 163.367
R2383 B.n1037 B.n411 163.367
R2384 B.n1045 B.n411 163.367
R2385 B.n1046 B.n1045 163.367
R2386 B.n1046 B.n5 163.367
R2387 B.n6 B.n5 163.367
R2388 B.n7 B.n6 163.367
R2389 B.n1051 B.n7 163.367
R2390 B.n1051 B.n12 163.367
R2391 B.n13 B.n12 163.367
R2392 B.n14 B.n13 163.367
R2393 B.n1056 B.n14 163.367
R2394 B.n1056 B.n19 163.367
R2395 B.n20 B.n19 163.367
R2396 B.n21 B.n20 163.367
R2397 B.n1061 B.n21 163.367
R2398 B.n1061 B.n26 163.367
R2399 B.n27 B.n26 163.367
R2400 B.n28 B.n27 163.367
R2401 B.n1066 B.n28 163.367
R2402 B.n1066 B.n33 163.367
R2403 B.n34 B.n33 163.367
R2404 B.n35 B.n34 163.367
R2405 B.n1071 B.n35 163.367
R2406 B.n1071 B.n40 163.367
R2407 B.n41 B.n40 163.367
R2408 B.n42 B.n41 163.367
R2409 B.n1076 B.n42 163.367
R2410 B.n1076 B.n47 163.367
R2411 B.n48 B.n47 163.367
R2412 B.n49 B.n48 163.367
R2413 B.n1081 B.n49 163.367
R2414 B.n1081 B.n54 163.367
R2415 B.n55 B.n54 163.367
R2416 B.n56 B.n55 163.367
R2417 B.n1086 B.n56 163.367
R2418 B.n1086 B.n61 163.367
R2419 B.n62 B.n61 163.367
R2420 B.n63 B.n62 163.367
R2421 B.n1091 B.n63 163.367
R2422 B.n1091 B.n68 163.367
R2423 B.n69 B.n68 163.367
R2424 B.n70 B.n69 163.367
R2425 B.n1096 B.n70 163.367
R2426 B.n1096 B.n75 163.367
R2427 B.n76 B.n75 163.367
R2428 B.n77 B.n76 163.367
R2429 B.n1101 B.n77 163.367
R2430 B.n1101 B.n82 163.367
R2431 B.n83 B.n82 163.367
R2432 B.n84 B.n83 163.367
R2433 B.n1106 B.n84 163.367
R2434 B.n1106 B.n89 163.367
R2435 B.n90 B.n89 163.367
R2436 B.n91 B.n90 163.367
R2437 B.n1111 B.n91 163.367
R2438 B.n1111 B.n96 163.367
R2439 B.n97 B.n96 163.367
R2440 B.n98 B.n97 163.367
R2441 B.n1116 B.n98 163.367
R2442 B.n1116 B.n103 163.367
R2443 B.n104 B.n103 163.367
R2444 B.n105 B.n104 163.367
R2445 B.n1121 B.n105 163.367
R2446 B.n1121 B.n110 163.367
R2447 B.n111 B.n110 163.367
R2448 B.n112 B.n111 163.367
R2449 B.n1126 B.n112 163.367
R2450 B.n1126 B.n117 163.367
R2451 B.n118 B.n117 163.367
R2452 B.n119 B.n118 163.367
R2453 B.n1131 B.n119 163.367
R2454 B.n1131 B.n124 163.367
R2455 B.n125 B.n124 163.367
R2456 B.n126 B.n125 163.367
R2457 B.n186 B.n126 163.367
R2458 B.n191 B.n130 163.367
R2459 B.n195 B.n194 163.367
R2460 B.n199 B.n198 163.367
R2461 B.n203 B.n202 163.367
R2462 B.n207 B.n206 163.367
R2463 B.n211 B.n210 163.367
R2464 B.n215 B.n214 163.367
R2465 B.n219 B.n218 163.367
R2466 B.n223 B.n222 163.367
R2467 B.n227 B.n226 163.367
R2468 B.n231 B.n230 163.367
R2469 B.n235 B.n234 163.367
R2470 B.n239 B.n238 163.367
R2471 B.n243 B.n242 163.367
R2472 B.n247 B.n246 163.367
R2473 B.n251 B.n250 163.367
R2474 B.n255 B.n254 163.367
R2475 B.n259 B.n258 163.367
R2476 B.n263 B.n262 163.367
R2477 B.n267 B.n266 163.367
R2478 B.n271 B.n270 163.367
R2479 B.n275 B.n274 163.367
R2480 B.n279 B.n278 163.367
R2481 B.n283 B.n282 163.367
R2482 B.n287 B.n286 163.367
R2483 B.n292 B.n291 163.367
R2484 B.n296 B.n295 163.367
R2485 B.n300 B.n299 163.367
R2486 B.n304 B.n303 163.367
R2487 B.n308 B.n307 163.367
R2488 B.n313 B.n312 163.367
R2489 B.n317 B.n316 163.367
R2490 B.n321 B.n320 163.367
R2491 B.n325 B.n324 163.367
R2492 B.n329 B.n328 163.367
R2493 B.n333 B.n332 163.367
R2494 B.n337 B.n336 163.367
R2495 B.n341 B.n340 163.367
R2496 B.n345 B.n344 163.367
R2497 B.n349 B.n348 163.367
R2498 B.n353 B.n352 163.367
R2499 B.n357 B.n356 163.367
R2500 B.n361 B.n360 163.367
R2501 B.n365 B.n364 163.367
R2502 B.n369 B.n368 163.367
R2503 B.n373 B.n372 163.367
R2504 B.n377 B.n376 163.367
R2505 B.n381 B.n380 163.367
R2506 B.n385 B.n384 163.367
R2507 B.n389 B.n388 163.367
R2508 B.n393 B.n392 163.367
R2509 B.n397 B.n396 163.367
R2510 B.n401 B.n400 163.367
R2511 B.n405 B.n404 163.367
R2512 B.n407 B.n185 163.367
R2513 B.n612 B.n611 83.0066
R2514 B.n609 B.n608 83.0066
R2515 B.n190 B.n189 83.0066
R2516 B.n188 B.n187 83.0066
R2517 B.n834 B.n833 71.676
R2518 B.n607 B.n552 71.676
R2519 B.n826 B.n553 71.676
R2520 B.n822 B.n554 71.676
R2521 B.n818 B.n555 71.676
R2522 B.n814 B.n556 71.676
R2523 B.n810 B.n557 71.676
R2524 B.n806 B.n558 71.676
R2525 B.n802 B.n559 71.676
R2526 B.n798 B.n560 71.676
R2527 B.n794 B.n561 71.676
R2528 B.n790 B.n562 71.676
R2529 B.n786 B.n563 71.676
R2530 B.n782 B.n564 71.676
R2531 B.n778 B.n565 71.676
R2532 B.n774 B.n566 71.676
R2533 B.n770 B.n567 71.676
R2534 B.n766 B.n568 71.676
R2535 B.n762 B.n569 71.676
R2536 B.n758 B.n570 71.676
R2537 B.n754 B.n571 71.676
R2538 B.n750 B.n572 71.676
R2539 B.n746 B.n573 71.676
R2540 B.n742 B.n574 71.676
R2541 B.n738 B.n575 71.676
R2542 B.n734 B.n576 71.676
R2543 B.n730 B.n577 71.676
R2544 B.n726 B.n578 71.676
R2545 B.n722 B.n579 71.676
R2546 B.n718 B.n580 71.676
R2547 B.n714 B.n581 71.676
R2548 B.n710 B.n582 71.676
R2549 B.n706 B.n583 71.676
R2550 B.n702 B.n584 71.676
R2551 B.n698 B.n585 71.676
R2552 B.n694 B.n586 71.676
R2553 B.n690 B.n587 71.676
R2554 B.n686 B.n588 71.676
R2555 B.n682 B.n589 71.676
R2556 B.n678 B.n590 71.676
R2557 B.n674 B.n591 71.676
R2558 B.n670 B.n592 71.676
R2559 B.n666 B.n593 71.676
R2560 B.n662 B.n594 71.676
R2561 B.n658 B.n595 71.676
R2562 B.n654 B.n596 71.676
R2563 B.n650 B.n597 71.676
R2564 B.n646 B.n598 71.676
R2565 B.n642 B.n599 71.676
R2566 B.n638 B.n600 71.676
R2567 B.n634 B.n601 71.676
R2568 B.n630 B.n602 71.676
R2569 B.n626 B.n603 71.676
R2570 B.n622 B.n604 71.676
R2571 B.n618 B.n605 71.676
R2572 B.n1142 B.n1141 71.676
R2573 B.n191 B.n131 71.676
R2574 B.n195 B.n132 71.676
R2575 B.n199 B.n133 71.676
R2576 B.n203 B.n134 71.676
R2577 B.n207 B.n135 71.676
R2578 B.n211 B.n136 71.676
R2579 B.n215 B.n137 71.676
R2580 B.n219 B.n138 71.676
R2581 B.n223 B.n139 71.676
R2582 B.n227 B.n140 71.676
R2583 B.n231 B.n141 71.676
R2584 B.n235 B.n142 71.676
R2585 B.n239 B.n143 71.676
R2586 B.n243 B.n144 71.676
R2587 B.n247 B.n145 71.676
R2588 B.n251 B.n146 71.676
R2589 B.n255 B.n147 71.676
R2590 B.n259 B.n148 71.676
R2591 B.n263 B.n149 71.676
R2592 B.n267 B.n150 71.676
R2593 B.n271 B.n151 71.676
R2594 B.n275 B.n152 71.676
R2595 B.n279 B.n153 71.676
R2596 B.n283 B.n154 71.676
R2597 B.n287 B.n155 71.676
R2598 B.n292 B.n156 71.676
R2599 B.n296 B.n157 71.676
R2600 B.n300 B.n158 71.676
R2601 B.n304 B.n159 71.676
R2602 B.n308 B.n160 71.676
R2603 B.n313 B.n161 71.676
R2604 B.n317 B.n162 71.676
R2605 B.n321 B.n163 71.676
R2606 B.n325 B.n164 71.676
R2607 B.n329 B.n165 71.676
R2608 B.n333 B.n166 71.676
R2609 B.n337 B.n167 71.676
R2610 B.n341 B.n168 71.676
R2611 B.n345 B.n169 71.676
R2612 B.n349 B.n170 71.676
R2613 B.n353 B.n171 71.676
R2614 B.n357 B.n172 71.676
R2615 B.n361 B.n173 71.676
R2616 B.n365 B.n174 71.676
R2617 B.n369 B.n175 71.676
R2618 B.n373 B.n176 71.676
R2619 B.n377 B.n177 71.676
R2620 B.n381 B.n178 71.676
R2621 B.n385 B.n179 71.676
R2622 B.n389 B.n180 71.676
R2623 B.n393 B.n181 71.676
R2624 B.n397 B.n182 71.676
R2625 B.n401 B.n183 71.676
R2626 B.n405 B.n184 71.676
R2627 B.n1139 B.n185 71.676
R2628 B.n1139 B.n1138 71.676
R2629 B.n407 B.n184 71.676
R2630 B.n404 B.n183 71.676
R2631 B.n400 B.n182 71.676
R2632 B.n396 B.n181 71.676
R2633 B.n392 B.n180 71.676
R2634 B.n388 B.n179 71.676
R2635 B.n384 B.n178 71.676
R2636 B.n380 B.n177 71.676
R2637 B.n376 B.n176 71.676
R2638 B.n372 B.n175 71.676
R2639 B.n368 B.n174 71.676
R2640 B.n364 B.n173 71.676
R2641 B.n360 B.n172 71.676
R2642 B.n356 B.n171 71.676
R2643 B.n352 B.n170 71.676
R2644 B.n348 B.n169 71.676
R2645 B.n344 B.n168 71.676
R2646 B.n340 B.n167 71.676
R2647 B.n336 B.n166 71.676
R2648 B.n332 B.n165 71.676
R2649 B.n328 B.n164 71.676
R2650 B.n324 B.n163 71.676
R2651 B.n320 B.n162 71.676
R2652 B.n316 B.n161 71.676
R2653 B.n312 B.n160 71.676
R2654 B.n307 B.n159 71.676
R2655 B.n303 B.n158 71.676
R2656 B.n299 B.n157 71.676
R2657 B.n295 B.n156 71.676
R2658 B.n291 B.n155 71.676
R2659 B.n286 B.n154 71.676
R2660 B.n282 B.n153 71.676
R2661 B.n278 B.n152 71.676
R2662 B.n274 B.n151 71.676
R2663 B.n270 B.n150 71.676
R2664 B.n266 B.n149 71.676
R2665 B.n262 B.n148 71.676
R2666 B.n258 B.n147 71.676
R2667 B.n254 B.n146 71.676
R2668 B.n250 B.n145 71.676
R2669 B.n246 B.n144 71.676
R2670 B.n242 B.n143 71.676
R2671 B.n238 B.n142 71.676
R2672 B.n234 B.n141 71.676
R2673 B.n230 B.n140 71.676
R2674 B.n226 B.n139 71.676
R2675 B.n222 B.n138 71.676
R2676 B.n218 B.n137 71.676
R2677 B.n214 B.n136 71.676
R2678 B.n210 B.n135 71.676
R2679 B.n206 B.n134 71.676
R2680 B.n202 B.n133 71.676
R2681 B.n198 B.n132 71.676
R2682 B.n194 B.n131 71.676
R2683 B.n1141 B.n130 71.676
R2684 B.n833 B.n551 71.676
R2685 B.n827 B.n552 71.676
R2686 B.n823 B.n553 71.676
R2687 B.n819 B.n554 71.676
R2688 B.n815 B.n555 71.676
R2689 B.n811 B.n556 71.676
R2690 B.n807 B.n557 71.676
R2691 B.n803 B.n558 71.676
R2692 B.n799 B.n559 71.676
R2693 B.n795 B.n560 71.676
R2694 B.n791 B.n561 71.676
R2695 B.n787 B.n562 71.676
R2696 B.n783 B.n563 71.676
R2697 B.n779 B.n564 71.676
R2698 B.n775 B.n565 71.676
R2699 B.n771 B.n566 71.676
R2700 B.n767 B.n567 71.676
R2701 B.n763 B.n568 71.676
R2702 B.n759 B.n569 71.676
R2703 B.n755 B.n570 71.676
R2704 B.n751 B.n571 71.676
R2705 B.n747 B.n572 71.676
R2706 B.n743 B.n573 71.676
R2707 B.n739 B.n574 71.676
R2708 B.n735 B.n575 71.676
R2709 B.n731 B.n576 71.676
R2710 B.n727 B.n577 71.676
R2711 B.n723 B.n578 71.676
R2712 B.n719 B.n579 71.676
R2713 B.n715 B.n580 71.676
R2714 B.n711 B.n581 71.676
R2715 B.n707 B.n582 71.676
R2716 B.n703 B.n583 71.676
R2717 B.n699 B.n584 71.676
R2718 B.n695 B.n585 71.676
R2719 B.n691 B.n586 71.676
R2720 B.n687 B.n587 71.676
R2721 B.n683 B.n588 71.676
R2722 B.n679 B.n589 71.676
R2723 B.n675 B.n590 71.676
R2724 B.n671 B.n591 71.676
R2725 B.n667 B.n592 71.676
R2726 B.n663 B.n593 71.676
R2727 B.n659 B.n594 71.676
R2728 B.n655 B.n595 71.676
R2729 B.n651 B.n596 71.676
R2730 B.n647 B.n597 71.676
R2731 B.n643 B.n598 71.676
R2732 B.n639 B.n599 71.676
R2733 B.n635 B.n600 71.676
R2734 B.n631 B.n601 71.676
R2735 B.n627 B.n602 71.676
R2736 B.n623 B.n603 71.676
R2737 B.n619 B.n604 71.676
R2738 B.n615 B.n605 71.676
R2739 B.n832 B.n548 67.7338
R2740 B.n1140 B.n127 67.7338
R2741 B.n613 B.n612 59.5399
R2742 B.n610 B.n609 59.5399
R2743 B.n289 B.n190 59.5399
R2744 B.n310 B.n188 59.5399
R2745 B.n839 B.n548 36.2672
R2746 B.n839 B.n544 36.2672
R2747 B.n845 B.n544 36.2672
R2748 B.n845 B.n540 36.2672
R2749 B.n851 B.n540 36.2672
R2750 B.n851 B.n536 36.2672
R2751 B.n857 B.n536 36.2672
R2752 B.n857 B.n532 36.2672
R2753 B.n863 B.n532 36.2672
R2754 B.n869 B.n528 36.2672
R2755 B.n869 B.n524 36.2672
R2756 B.n875 B.n524 36.2672
R2757 B.n875 B.n520 36.2672
R2758 B.n881 B.n520 36.2672
R2759 B.n881 B.n516 36.2672
R2760 B.n887 B.n516 36.2672
R2761 B.n887 B.n512 36.2672
R2762 B.n893 B.n512 36.2672
R2763 B.n893 B.n508 36.2672
R2764 B.n899 B.n508 36.2672
R2765 B.n899 B.n504 36.2672
R2766 B.n905 B.n504 36.2672
R2767 B.n905 B.n500 36.2672
R2768 B.n911 B.n500 36.2672
R2769 B.n917 B.n496 36.2672
R2770 B.n917 B.n492 36.2672
R2771 B.n923 B.n492 36.2672
R2772 B.n923 B.n488 36.2672
R2773 B.n929 B.n488 36.2672
R2774 B.n929 B.n484 36.2672
R2775 B.n935 B.n484 36.2672
R2776 B.n935 B.n480 36.2672
R2777 B.n941 B.n480 36.2672
R2778 B.n941 B.n476 36.2672
R2779 B.n947 B.n476 36.2672
R2780 B.n953 B.n472 36.2672
R2781 B.n953 B.n468 36.2672
R2782 B.n959 B.n468 36.2672
R2783 B.n959 B.n464 36.2672
R2784 B.n965 B.n464 36.2672
R2785 B.n965 B.n460 36.2672
R2786 B.n971 B.n460 36.2672
R2787 B.n971 B.n456 36.2672
R2788 B.n977 B.n456 36.2672
R2789 B.n977 B.n451 36.2672
R2790 B.n983 B.n451 36.2672
R2791 B.n983 B.n452 36.2672
R2792 B.n989 B.n444 36.2672
R2793 B.n995 B.n444 36.2672
R2794 B.n995 B.n440 36.2672
R2795 B.n1001 B.n440 36.2672
R2796 B.n1001 B.n436 36.2672
R2797 B.n1007 B.n436 36.2672
R2798 B.n1007 B.n432 36.2672
R2799 B.n1013 B.n432 36.2672
R2800 B.n1013 B.n428 36.2672
R2801 B.n1019 B.n428 36.2672
R2802 B.n1019 B.n424 36.2672
R2803 B.n1025 B.n424 36.2672
R2804 B.n1031 B.n420 36.2672
R2805 B.n1031 B.n416 36.2672
R2806 B.n1038 B.n416 36.2672
R2807 B.n1038 B.n412 36.2672
R2808 B.n1044 B.n412 36.2672
R2809 B.n1044 B.n4 36.2672
R2810 B.n1285 B.n4 36.2672
R2811 B.n1285 B.n1284 36.2672
R2812 B.n1284 B.n1283 36.2672
R2813 B.n1283 B.n8 36.2672
R2814 B.n1277 B.n8 36.2672
R2815 B.n1277 B.n1276 36.2672
R2816 B.n1276 B.n1275 36.2672
R2817 B.n1275 B.n15 36.2672
R2818 B.n1269 B.n1268 36.2672
R2819 B.n1268 B.n1267 36.2672
R2820 B.n1267 B.n22 36.2672
R2821 B.n1261 B.n22 36.2672
R2822 B.n1261 B.n1260 36.2672
R2823 B.n1260 B.n1259 36.2672
R2824 B.n1259 B.n29 36.2672
R2825 B.n1253 B.n29 36.2672
R2826 B.n1253 B.n1252 36.2672
R2827 B.n1252 B.n1251 36.2672
R2828 B.n1251 B.n36 36.2672
R2829 B.n1245 B.n36 36.2672
R2830 B.n1244 B.n1243 36.2672
R2831 B.n1243 B.n43 36.2672
R2832 B.n1237 B.n43 36.2672
R2833 B.n1237 B.n1236 36.2672
R2834 B.n1236 B.n1235 36.2672
R2835 B.n1235 B.n50 36.2672
R2836 B.n1229 B.n50 36.2672
R2837 B.n1229 B.n1228 36.2672
R2838 B.n1228 B.n1227 36.2672
R2839 B.n1227 B.n57 36.2672
R2840 B.n1221 B.n57 36.2672
R2841 B.n1221 B.n1220 36.2672
R2842 B.n1219 B.n64 36.2672
R2843 B.n1213 B.n64 36.2672
R2844 B.n1213 B.n1212 36.2672
R2845 B.n1212 B.n1211 36.2672
R2846 B.n1211 B.n71 36.2672
R2847 B.n1205 B.n71 36.2672
R2848 B.n1205 B.n1204 36.2672
R2849 B.n1204 B.n1203 36.2672
R2850 B.n1203 B.n78 36.2672
R2851 B.n1197 B.n78 36.2672
R2852 B.n1197 B.n1196 36.2672
R2853 B.n1195 B.n85 36.2672
R2854 B.n1189 B.n85 36.2672
R2855 B.n1189 B.n1188 36.2672
R2856 B.n1188 B.n1187 36.2672
R2857 B.n1187 B.n92 36.2672
R2858 B.n1181 B.n92 36.2672
R2859 B.n1181 B.n1180 36.2672
R2860 B.n1180 B.n1179 36.2672
R2861 B.n1179 B.n99 36.2672
R2862 B.n1173 B.n99 36.2672
R2863 B.n1173 B.n1172 36.2672
R2864 B.n1172 B.n1171 36.2672
R2865 B.n1171 B.n106 36.2672
R2866 B.n1165 B.n106 36.2672
R2867 B.n1165 B.n1164 36.2672
R2868 B.n1163 B.n113 36.2672
R2869 B.n1157 B.n113 36.2672
R2870 B.n1157 B.n1156 36.2672
R2871 B.n1156 B.n1155 36.2672
R2872 B.n1155 B.n120 36.2672
R2873 B.n1149 B.n120 36.2672
R2874 B.n1149 B.n1148 36.2672
R2875 B.n1148 B.n1147 36.2672
R2876 B.n1147 B.n127 36.2672
R2877 B.n1144 B.n1143 35.7468
R2878 B.n1137 B.n1136 35.7468
R2879 B.n614 B.n546 35.7468
R2880 B.n836 B.n835 35.7468
R2881 B.n947 B.t5 33.6005
R2882 B.t1 B.n1219 33.6005
R2883 B.t3 B.n420 32.5338
R2884 B.t4 B.n15 32.5338
R2885 B.t6 B.n496 24.0005
R2886 B.n1196 B.t0 24.0005
R2887 B.n863 B.t8 19.7338
R2888 B.t15 B.n1163 19.7338
R2889 B.n452 B.t2 18.6672
R2890 B.t21 B.n1244 18.6672
R2891 B B.n1287 18.0485
R2892 B.n989 B.t2 17.6005
R2893 B.n1245 B.t21 17.6005
R2894 B.t8 B.n528 16.5338
R2895 B.n1164 B.t15 16.5338
R2896 B.n911 B.t6 12.2672
R2897 B.t0 B.n1195 12.2672
R2898 B.n1143 B.n129 10.6151
R2899 B.n192 B.n129 10.6151
R2900 B.n193 B.n192 10.6151
R2901 B.n196 B.n193 10.6151
R2902 B.n197 B.n196 10.6151
R2903 B.n200 B.n197 10.6151
R2904 B.n201 B.n200 10.6151
R2905 B.n204 B.n201 10.6151
R2906 B.n205 B.n204 10.6151
R2907 B.n208 B.n205 10.6151
R2908 B.n209 B.n208 10.6151
R2909 B.n212 B.n209 10.6151
R2910 B.n213 B.n212 10.6151
R2911 B.n216 B.n213 10.6151
R2912 B.n217 B.n216 10.6151
R2913 B.n220 B.n217 10.6151
R2914 B.n221 B.n220 10.6151
R2915 B.n224 B.n221 10.6151
R2916 B.n225 B.n224 10.6151
R2917 B.n228 B.n225 10.6151
R2918 B.n229 B.n228 10.6151
R2919 B.n232 B.n229 10.6151
R2920 B.n233 B.n232 10.6151
R2921 B.n236 B.n233 10.6151
R2922 B.n237 B.n236 10.6151
R2923 B.n240 B.n237 10.6151
R2924 B.n241 B.n240 10.6151
R2925 B.n244 B.n241 10.6151
R2926 B.n245 B.n244 10.6151
R2927 B.n248 B.n245 10.6151
R2928 B.n249 B.n248 10.6151
R2929 B.n252 B.n249 10.6151
R2930 B.n253 B.n252 10.6151
R2931 B.n256 B.n253 10.6151
R2932 B.n257 B.n256 10.6151
R2933 B.n260 B.n257 10.6151
R2934 B.n261 B.n260 10.6151
R2935 B.n264 B.n261 10.6151
R2936 B.n265 B.n264 10.6151
R2937 B.n268 B.n265 10.6151
R2938 B.n269 B.n268 10.6151
R2939 B.n272 B.n269 10.6151
R2940 B.n273 B.n272 10.6151
R2941 B.n276 B.n273 10.6151
R2942 B.n277 B.n276 10.6151
R2943 B.n280 B.n277 10.6151
R2944 B.n281 B.n280 10.6151
R2945 B.n284 B.n281 10.6151
R2946 B.n285 B.n284 10.6151
R2947 B.n288 B.n285 10.6151
R2948 B.n293 B.n290 10.6151
R2949 B.n294 B.n293 10.6151
R2950 B.n297 B.n294 10.6151
R2951 B.n298 B.n297 10.6151
R2952 B.n301 B.n298 10.6151
R2953 B.n302 B.n301 10.6151
R2954 B.n305 B.n302 10.6151
R2955 B.n306 B.n305 10.6151
R2956 B.n309 B.n306 10.6151
R2957 B.n314 B.n311 10.6151
R2958 B.n315 B.n314 10.6151
R2959 B.n318 B.n315 10.6151
R2960 B.n319 B.n318 10.6151
R2961 B.n322 B.n319 10.6151
R2962 B.n323 B.n322 10.6151
R2963 B.n326 B.n323 10.6151
R2964 B.n327 B.n326 10.6151
R2965 B.n330 B.n327 10.6151
R2966 B.n331 B.n330 10.6151
R2967 B.n334 B.n331 10.6151
R2968 B.n335 B.n334 10.6151
R2969 B.n338 B.n335 10.6151
R2970 B.n339 B.n338 10.6151
R2971 B.n342 B.n339 10.6151
R2972 B.n343 B.n342 10.6151
R2973 B.n346 B.n343 10.6151
R2974 B.n347 B.n346 10.6151
R2975 B.n350 B.n347 10.6151
R2976 B.n351 B.n350 10.6151
R2977 B.n354 B.n351 10.6151
R2978 B.n355 B.n354 10.6151
R2979 B.n358 B.n355 10.6151
R2980 B.n359 B.n358 10.6151
R2981 B.n362 B.n359 10.6151
R2982 B.n363 B.n362 10.6151
R2983 B.n366 B.n363 10.6151
R2984 B.n367 B.n366 10.6151
R2985 B.n370 B.n367 10.6151
R2986 B.n371 B.n370 10.6151
R2987 B.n374 B.n371 10.6151
R2988 B.n375 B.n374 10.6151
R2989 B.n378 B.n375 10.6151
R2990 B.n379 B.n378 10.6151
R2991 B.n382 B.n379 10.6151
R2992 B.n383 B.n382 10.6151
R2993 B.n386 B.n383 10.6151
R2994 B.n387 B.n386 10.6151
R2995 B.n390 B.n387 10.6151
R2996 B.n391 B.n390 10.6151
R2997 B.n394 B.n391 10.6151
R2998 B.n395 B.n394 10.6151
R2999 B.n398 B.n395 10.6151
R3000 B.n399 B.n398 10.6151
R3001 B.n402 B.n399 10.6151
R3002 B.n403 B.n402 10.6151
R3003 B.n406 B.n403 10.6151
R3004 B.n408 B.n406 10.6151
R3005 B.n409 B.n408 10.6151
R3006 B.n1137 B.n409 10.6151
R3007 B.n841 B.n546 10.6151
R3008 B.n842 B.n841 10.6151
R3009 B.n843 B.n842 10.6151
R3010 B.n843 B.n538 10.6151
R3011 B.n853 B.n538 10.6151
R3012 B.n854 B.n853 10.6151
R3013 B.n855 B.n854 10.6151
R3014 B.n855 B.n530 10.6151
R3015 B.n865 B.n530 10.6151
R3016 B.n866 B.n865 10.6151
R3017 B.n867 B.n866 10.6151
R3018 B.n867 B.n522 10.6151
R3019 B.n877 B.n522 10.6151
R3020 B.n878 B.n877 10.6151
R3021 B.n879 B.n878 10.6151
R3022 B.n879 B.n514 10.6151
R3023 B.n889 B.n514 10.6151
R3024 B.n890 B.n889 10.6151
R3025 B.n891 B.n890 10.6151
R3026 B.n891 B.n506 10.6151
R3027 B.n901 B.n506 10.6151
R3028 B.n902 B.n901 10.6151
R3029 B.n903 B.n902 10.6151
R3030 B.n903 B.n498 10.6151
R3031 B.n913 B.n498 10.6151
R3032 B.n914 B.n913 10.6151
R3033 B.n915 B.n914 10.6151
R3034 B.n915 B.n490 10.6151
R3035 B.n925 B.n490 10.6151
R3036 B.n926 B.n925 10.6151
R3037 B.n927 B.n926 10.6151
R3038 B.n927 B.n482 10.6151
R3039 B.n937 B.n482 10.6151
R3040 B.n938 B.n937 10.6151
R3041 B.n939 B.n938 10.6151
R3042 B.n939 B.n474 10.6151
R3043 B.n949 B.n474 10.6151
R3044 B.n950 B.n949 10.6151
R3045 B.n951 B.n950 10.6151
R3046 B.n951 B.n466 10.6151
R3047 B.n961 B.n466 10.6151
R3048 B.n962 B.n961 10.6151
R3049 B.n963 B.n962 10.6151
R3050 B.n963 B.n458 10.6151
R3051 B.n973 B.n458 10.6151
R3052 B.n974 B.n973 10.6151
R3053 B.n975 B.n974 10.6151
R3054 B.n975 B.n449 10.6151
R3055 B.n985 B.n449 10.6151
R3056 B.n986 B.n985 10.6151
R3057 B.n987 B.n986 10.6151
R3058 B.n987 B.n442 10.6151
R3059 B.n997 B.n442 10.6151
R3060 B.n998 B.n997 10.6151
R3061 B.n999 B.n998 10.6151
R3062 B.n999 B.n434 10.6151
R3063 B.n1009 B.n434 10.6151
R3064 B.n1010 B.n1009 10.6151
R3065 B.n1011 B.n1010 10.6151
R3066 B.n1011 B.n426 10.6151
R3067 B.n1021 B.n426 10.6151
R3068 B.n1022 B.n1021 10.6151
R3069 B.n1023 B.n1022 10.6151
R3070 B.n1023 B.n418 10.6151
R3071 B.n1033 B.n418 10.6151
R3072 B.n1034 B.n1033 10.6151
R3073 B.n1036 B.n1034 10.6151
R3074 B.n1036 B.n1035 10.6151
R3075 B.n1035 B.n410 10.6151
R3076 B.n1047 B.n410 10.6151
R3077 B.n1048 B.n1047 10.6151
R3078 B.n1049 B.n1048 10.6151
R3079 B.n1050 B.n1049 10.6151
R3080 B.n1052 B.n1050 10.6151
R3081 B.n1053 B.n1052 10.6151
R3082 B.n1054 B.n1053 10.6151
R3083 B.n1055 B.n1054 10.6151
R3084 B.n1057 B.n1055 10.6151
R3085 B.n1058 B.n1057 10.6151
R3086 B.n1059 B.n1058 10.6151
R3087 B.n1060 B.n1059 10.6151
R3088 B.n1062 B.n1060 10.6151
R3089 B.n1063 B.n1062 10.6151
R3090 B.n1064 B.n1063 10.6151
R3091 B.n1065 B.n1064 10.6151
R3092 B.n1067 B.n1065 10.6151
R3093 B.n1068 B.n1067 10.6151
R3094 B.n1069 B.n1068 10.6151
R3095 B.n1070 B.n1069 10.6151
R3096 B.n1072 B.n1070 10.6151
R3097 B.n1073 B.n1072 10.6151
R3098 B.n1074 B.n1073 10.6151
R3099 B.n1075 B.n1074 10.6151
R3100 B.n1077 B.n1075 10.6151
R3101 B.n1078 B.n1077 10.6151
R3102 B.n1079 B.n1078 10.6151
R3103 B.n1080 B.n1079 10.6151
R3104 B.n1082 B.n1080 10.6151
R3105 B.n1083 B.n1082 10.6151
R3106 B.n1084 B.n1083 10.6151
R3107 B.n1085 B.n1084 10.6151
R3108 B.n1087 B.n1085 10.6151
R3109 B.n1088 B.n1087 10.6151
R3110 B.n1089 B.n1088 10.6151
R3111 B.n1090 B.n1089 10.6151
R3112 B.n1092 B.n1090 10.6151
R3113 B.n1093 B.n1092 10.6151
R3114 B.n1094 B.n1093 10.6151
R3115 B.n1095 B.n1094 10.6151
R3116 B.n1097 B.n1095 10.6151
R3117 B.n1098 B.n1097 10.6151
R3118 B.n1099 B.n1098 10.6151
R3119 B.n1100 B.n1099 10.6151
R3120 B.n1102 B.n1100 10.6151
R3121 B.n1103 B.n1102 10.6151
R3122 B.n1104 B.n1103 10.6151
R3123 B.n1105 B.n1104 10.6151
R3124 B.n1107 B.n1105 10.6151
R3125 B.n1108 B.n1107 10.6151
R3126 B.n1109 B.n1108 10.6151
R3127 B.n1110 B.n1109 10.6151
R3128 B.n1112 B.n1110 10.6151
R3129 B.n1113 B.n1112 10.6151
R3130 B.n1114 B.n1113 10.6151
R3131 B.n1115 B.n1114 10.6151
R3132 B.n1117 B.n1115 10.6151
R3133 B.n1118 B.n1117 10.6151
R3134 B.n1119 B.n1118 10.6151
R3135 B.n1120 B.n1119 10.6151
R3136 B.n1122 B.n1120 10.6151
R3137 B.n1123 B.n1122 10.6151
R3138 B.n1124 B.n1123 10.6151
R3139 B.n1125 B.n1124 10.6151
R3140 B.n1127 B.n1125 10.6151
R3141 B.n1128 B.n1127 10.6151
R3142 B.n1129 B.n1128 10.6151
R3143 B.n1130 B.n1129 10.6151
R3144 B.n1132 B.n1130 10.6151
R3145 B.n1133 B.n1132 10.6151
R3146 B.n1134 B.n1133 10.6151
R3147 B.n1135 B.n1134 10.6151
R3148 B.n1136 B.n1135 10.6151
R3149 B.n835 B.n550 10.6151
R3150 B.n830 B.n550 10.6151
R3151 B.n830 B.n829 10.6151
R3152 B.n829 B.n828 10.6151
R3153 B.n828 B.n825 10.6151
R3154 B.n825 B.n824 10.6151
R3155 B.n824 B.n821 10.6151
R3156 B.n821 B.n820 10.6151
R3157 B.n820 B.n817 10.6151
R3158 B.n817 B.n816 10.6151
R3159 B.n816 B.n813 10.6151
R3160 B.n813 B.n812 10.6151
R3161 B.n812 B.n809 10.6151
R3162 B.n809 B.n808 10.6151
R3163 B.n808 B.n805 10.6151
R3164 B.n805 B.n804 10.6151
R3165 B.n804 B.n801 10.6151
R3166 B.n801 B.n800 10.6151
R3167 B.n800 B.n797 10.6151
R3168 B.n797 B.n796 10.6151
R3169 B.n796 B.n793 10.6151
R3170 B.n793 B.n792 10.6151
R3171 B.n792 B.n789 10.6151
R3172 B.n789 B.n788 10.6151
R3173 B.n788 B.n785 10.6151
R3174 B.n785 B.n784 10.6151
R3175 B.n784 B.n781 10.6151
R3176 B.n781 B.n780 10.6151
R3177 B.n780 B.n777 10.6151
R3178 B.n777 B.n776 10.6151
R3179 B.n776 B.n773 10.6151
R3180 B.n773 B.n772 10.6151
R3181 B.n772 B.n769 10.6151
R3182 B.n769 B.n768 10.6151
R3183 B.n768 B.n765 10.6151
R3184 B.n765 B.n764 10.6151
R3185 B.n764 B.n761 10.6151
R3186 B.n761 B.n760 10.6151
R3187 B.n760 B.n757 10.6151
R3188 B.n757 B.n756 10.6151
R3189 B.n756 B.n753 10.6151
R3190 B.n753 B.n752 10.6151
R3191 B.n752 B.n749 10.6151
R3192 B.n749 B.n748 10.6151
R3193 B.n748 B.n745 10.6151
R3194 B.n745 B.n744 10.6151
R3195 B.n744 B.n741 10.6151
R3196 B.n741 B.n740 10.6151
R3197 B.n740 B.n737 10.6151
R3198 B.n737 B.n736 10.6151
R3199 B.n733 B.n732 10.6151
R3200 B.n732 B.n729 10.6151
R3201 B.n729 B.n728 10.6151
R3202 B.n728 B.n725 10.6151
R3203 B.n725 B.n724 10.6151
R3204 B.n724 B.n721 10.6151
R3205 B.n721 B.n720 10.6151
R3206 B.n720 B.n717 10.6151
R3207 B.n717 B.n716 10.6151
R3208 B.n713 B.n712 10.6151
R3209 B.n712 B.n709 10.6151
R3210 B.n709 B.n708 10.6151
R3211 B.n708 B.n705 10.6151
R3212 B.n705 B.n704 10.6151
R3213 B.n704 B.n701 10.6151
R3214 B.n701 B.n700 10.6151
R3215 B.n700 B.n697 10.6151
R3216 B.n697 B.n696 10.6151
R3217 B.n696 B.n693 10.6151
R3218 B.n693 B.n692 10.6151
R3219 B.n692 B.n689 10.6151
R3220 B.n689 B.n688 10.6151
R3221 B.n688 B.n685 10.6151
R3222 B.n685 B.n684 10.6151
R3223 B.n684 B.n681 10.6151
R3224 B.n681 B.n680 10.6151
R3225 B.n680 B.n677 10.6151
R3226 B.n677 B.n676 10.6151
R3227 B.n676 B.n673 10.6151
R3228 B.n673 B.n672 10.6151
R3229 B.n672 B.n669 10.6151
R3230 B.n669 B.n668 10.6151
R3231 B.n668 B.n665 10.6151
R3232 B.n665 B.n664 10.6151
R3233 B.n664 B.n661 10.6151
R3234 B.n661 B.n660 10.6151
R3235 B.n660 B.n657 10.6151
R3236 B.n657 B.n656 10.6151
R3237 B.n656 B.n653 10.6151
R3238 B.n653 B.n652 10.6151
R3239 B.n652 B.n649 10.6151
R3240 B.n649 B.n648 10.6151
R3241 B.n648 B.n645 10.6151
R3242 B.n645 B.n644 10.6151
R3243 B.n644 B.n641 10.6151
R3244 B.n641 B.n640 10.6151
R3245 B.n640 B.n637 10.6151
R3246 B.n637 B.n636 10.6151
R3247 B.n636 B.n633 10.6151
R3248 B.n633 B.n632 10.6151
R3249 B.n632 B.n629 10.6151
R3250 B.n629 B.n628 10.6151
R3251 B.n628 B.n625 10.6151
R3252 B.n625 B.n624 10.6151
R3253 B.n624 B.n621 10.6151
R3254 B.n621 B.n620 10.6151
R3255 B.n620 B.n617 10.6151
R3256 B.n617 B.n616 10.6151
R3257 B.n616 B.n614 10.6151
R3258 B.n837 B.n836 10.6151
R3259 B.n837 B.n542 10.6151
R3260 B.n847 B.n542 10.6151
R3261 B.n848 B.n847 10.6151
R3262 B.n849 B.n848 10.6151
R3263 B.n849 B.n534 10.6151
R3264 B.n859 B.n534 10.6151
R3265 B.n860 B.n859 10.6151
R3266 B.n861 B.n860 10.6151
R3267 B.n861 B.n526 10.6151
R3268 B.n871 B.n526 10.6151
R3269 B.n872 B.n871 10.6151
R3270 B.n873 B.n872 10.6151
R3271 B.n873 B.n518 10.6151
R3272 B.n883 B.n518 10.6151
R3273 B.n884 B.n883 10.6151
R3274 B.n885 B.n884 10.6151
R3275 B.n885 B.n510 10.6151
R3276 B.n895 B.n510 10.6151
R3277 B.n896 B.n895 10.6151
R3278 B.n897 B.n896 10.6151
R3279 B.n897 B.n502 10.6151
R3280 B.n907 B.n502 10.6151
R3281 B.n908 B.n907 10.6151
R3282 B.n909 B.n908 10.6151
R3283 B.n909 B.n494 10.6151
R3284 B.n919 B.n494 10.6151
R3285 B.n920 B.n919 10.6151
R3286 B.n921 B.n920 10.6151
R3287 B.n921 B.n486 10.6151
R3288 B.n931 B.n486 10.6151
R3289 B.n932 B.n931 10.6151
R3290 B.n933 B.n932 10.6151
R3291 B.n933 B.n478 10.6151
R3292 B.n943 B.n478 10.6151
R3293 B.n944 B.n943 10.6151
R3294 B.n945 B.n944 10.6151
R3295 B.n945 B.n470 10.6151
R3296 B.n955 B.n470 10.6151
R3297 B.n956 B.n955 10.6151
R3298 B.n957 B.n956 10.6151
R3299 B.n957 B.n462 10.6151
R3300 B.n967 B.n462 10.6151
R3301 B.n968 B.n967 10.6151
R3302 B.n969 B.n968 10.6151
R3303 B.n969 B.n454 10.6151
R3304 B.n979 B.n454 10.6151
R3305 B.n980 B.n979 10.6151
R3306 B.n981 B.n980 10.6151
R3307 B.n981 B.n446 10.6151
R3308 B.n991 B.n446 10.6151
R3309 B.n992 B.n991 10.6151
R3310 B.n993 B.n992 10.6151
R3311 B.n993 B.n438 10.6151
R3312 B.n1003 B.n438 10.6151
R3313 B.n1004 B.n1003 10.6151
R3314 B.n1005 B.n1004 10.6151
R3315 B.n1005 B.n430 10.6151
R3316 B.n1015 B.n430 10.6151
R3317 B.n1016 B.n1015 10.6151
R3318 B.n1017 B.n1016 10.6151
R3319 B.n1017 B.n422 10.6151
R3320 B.n1027 B.n422 10.6151
R3321 B.n1028 B.n1027 10.6151
R3322 B.n1029 B.n1028 10.6151
R3323 B.n1029 B.n414 10.6151
R3324 B.n1040 B.n414 10.6151
R3325 B.n1041 B.n1040 10.6151
R3326 B.n1042 B.n1041 10.6151
R3327 B.n1042 B.n0 10.6151
R3328 B.n1281 B.n1 10.6151
R3329 B.n1281 B.n1280 10.6151
R3330 B.n1280 B.n1279 10.6151
R3331 B.n1279 B.n10 10.6151
R3332 B.n1273 B.n10 10.6151
R3333 B.n1273 B.n1272 10.6151
R3334 B.n1272 B.n1271 10.6151
R3335 B.n1271 B.n17 10.6151
R3336 B.n1265 B.n17 10.6151
R3337 B.n1265 B.n1264 10.6151
R3338 B.n1264 B.n1263 10.6151
R3339 B.n1263 B.n24 10.6151
R3340 B.n1257 B.n24 10.6151
R3341 B.n1257 B.n1256 10.6151
R3342 B.n1256 B.n1255 10.6151
R3343 B.n1255 B.n31 10.6151
R3344 B.n1249 B.n31 10.6151
R3345 B.n1249 B.n1248 10.6151
R3346 B.n1248 B.n1247 10.6151
R3347 B.n1247 B.n38 10.6151
R3348 B.n1241 B.n38 10.6151
R3349 B.n1241 B.n1240 10.6151
R3350 B.n1240 B.n1239 10.6151
R3351 B.n1239 B.n45 10.6151
R3352 B.n1233 B.n45 10.6151
R3353 B.n1233 B.n1232 10.6151
R3354 B.n1232 B.n1231 10.6151
R3355 B.n1231 B.n52 10.6151
R3356 B.n1225 B.n52 10.6151
R3357 B.n1225 B.n1224 10.6151
R3358 B.n1224 B.n1223 10.6151
R3359 B.n1223 B.n59 10.6151
R3360 B.n1217 B.n59 10.6151
R3361 B.n1217 B.n1216 10.6151
R3362 B.n1216 B.n1215 10.6151
R3363 B.n1215 B.n66 10.6151
R3364 B.n1209 B.n66 10.6151
R3365 B.n1209 B.n1208 10.6151
R3366 B.n1208 B.n1207 10.6151
R3367 B.n1207 B.n73 10.6151
R3368 B.n1201 B.n73 10.6151
R3369 B.n1201 B.n1200 10.6151
R3370 B.n1200 B.n1199 10.6151
R3371 B.n1199 B.n80 10.6151
R3372 B.n1193 B.n80 10.6151
R3373 B.n1193 B.n1192 10.6151
R3374 B.n1192 B.n1191 10.6151
R3375 B.n1191 B.n87 10.6151
R3376 B.n1185 B.n87 10.6151
R3377 B.n1185 B.n1184 10.6151
R3378 B.n1184 B.n1183 10.6151
R3379 B.n1183 B.n94 10.6151
R3380 B.n1177 B.n94 10.6151
R3381 B.n1177 B.n1176 10.6151
R3382 B.n1176 B.n1175 10.6151
R3383 B.n1175 B.n101 10.6151
R3384 B.n1169 B.n101 10.6151
R3385 B.n1169 B.n1168 10.6151
R3386 B.n1168 B.n1167 10.6151
R3387 B.n1167 B.n108 10.6151
R3388 B.n1161 B.n108 10.6151
R3389 B.n1161 B.n1160 10.6151
R3390 B.n1160 B.n1159 10.6151
R3391 B.n1159 B.n115 10.6151
R3392 B.n1153 B.n115 10.6151
R3393 B.n1153 B.n1152 10.6151
R3394 B.n1152 B.n1151 10.6151
R3395 B.n1151 B.n122 10.6151
R3396 B.n1145 B.n122 10.6151
R3397 B.n1145 B.n1144 10.6151
R3398 B.n289 B.n288 9.36635
R3399 B.n311 B.n310 9.36635
R3400 B.n736 B.n610 9.36635
R3401 B.n713 B.n613 9.36635
R3402 B.n1025 B.t3 3.73383
R3403 B.n1269 B.t4 3.73383
R3404 B.n1287 B.n0 2.81026
R3405 B.n1287 B.n1 2.81026
R3406 B.t5 B.n472 2.66717
R3407 B.n1220 B.t1 2.66717
R3408 B.n290 B.n289 1.24928
R3409 B.n310 B.n309 1.24928
R3410 B.n733 B.n610 1.24928
R3411 B.n716 B.n613 1.24928
R3412 VP.n24 VP.n21 161.3
R3413 VP.n26 VP.n25 161.3
R3414 VP.n27 VP.n20 161.3
R3415 VP.n29 VP.n28 161.3
R3416 VP.n30 VP.n19 161.3
R3417 VP.n32 VP.n31 161.3
R3418 VP.n33 VP.n18 161.3
R3419 VP.n35 VP.n34 161.3
R3420 VP.n36 VP.n17 161.3
R3421 VP.n39 VP.n38 161.3
R3422 VP.n40 VP.n16 161.3
R3423 VP.n42 VP.n41 161.3
R3424 VP.n43 VP.n15 161.3
R3425 VP.n45 VP.n44 161.3
R3426 VP.n46 VP.n14 161.3
R3427 VP.n48 VP.n47 161.3
R3428 VP.n49 VP.n13 161.3
R3429 VP.n92 VP.n0 161.3
R3430 VP.n91 VP.n90 161.3
R3431 VP.n89 VP.n1 161.3
R3432 VP.n88 VP.n87 161.3
R3433 VP.n86 VP.n2 161.3
R3434 VP.n85 VP.n84 161.3
R3435 VP.n83 VP.n3 161.3
R3436 VP.n82 VP.n81 161.3
R3437 VP.n79 VP.n4 161.3
R3438 VP.n78 VP.n77 161.3
R3439 VP.n76 VP.n5 161.3
R3440 VP.n75 VP.n74 161.3
R3441 VP.n73 VP.n6 161.3
R3442 VP.n72 VP.n71 161.3
R3443 VP.n70 VP.n7 161.3
R3444 VP.n69 VP.n68 161.3
R3445 VP.n67 VP.n8 161.3
R3446 VP.n65 VP.n64 161.3
R3447 VP.n63 VP.n9 161.3
R3448 VP.n62 VP.n61 161.3
R3449 VP.n60 VP.n10 161.3
R3450 VP.n59 VP.n58 161.3
R3451 VP.n57 VP.n11 161.3
R3452 VP.n56 VP.n55 161.3
R3453 VP.n54 VP.n12 161.3
R3454 VP.n22 VP.t4 125.903
R3455 VP.n53 VP.t3 93.6549
R3456 VP.n66 VP.t1 93.6549
R3457 VP.n80 VP.t7 93.6549
R3458 VP.n93 VP.t5 93.6549
R3459 VP.n50 VP.t2 93.6549
R3460 VP.n37 VP.t0 93.6549
R3461 VP.n23 VP.t6 93.6549
R3462 VP.n23 VP.n22 68.2271
R3463 VP.n53 VP.n52 61.6295
R3464 VP.n94 VP.n93 61.6295
R3465 VP.n51 VP.n50 61.6295
R3466 VP.n52 VP.n51 59.9888
R3467 VP.n60 VP.n59 56.5193
R3468 VP.n87 VP.n86 56.5193
R3469 VP.n44 VP.n43 56.5193
R3470 VP.n73 VP.n72 40.4934
R3471 VP.n74 VP.n73 40.4934
R3472 VP.n31 VP.n30 40.4934
R3473 VP.n30 VP.n29 40.4934
R3474 VP.n55 VP.n54 24.4675
R3475 VP.n55 VP.n11 24.4675
R3476 VP.n59 VP.n11 24.4675
R3477 VP.n61 VP.n60 24.4675
R3478 VP.n61 VP.n9 24.4675
R3479 VP.n65 VP.n9 24.4675
R3480 VP.n68 VP.n67 24.4675
R3481 VP.n68 VP.n7 24.4675
R3482 VP.n72 VP.n7 24.4675
R3483 VP.n74 VP.n5 24.4675
R3484 VP.n78 VP.n5 24.4675
R3485 VP.n79 VP.n78 24.4675
R3486 VP.n81 VP.n3 24.4675
R3487 VP.n85 VP.n3 24.4675
R3488 VP.n86 VP.n85 24.4675
R3489 VP.n87 VP.n1 24.4675
R3490 VP.n91 VP.n1 24.4675
R3491 VP.n92 VP.n91 24.4675
R3492 VP.n44 VP.n14 24.4675
R3493 VP.n48 VP.n14 24.4675
R3494 VP.n49 VP.n48 24.4675
R3495 VP.n31 VP.n18 24.4675
R3496 VP.n35 VP.n18 24.4675
R3497 VP.n36 VP.n35 24.4675
R3498 VP.n38 VP.n16 24.4675
R3499 VP.n42 VP.n16 24.4675
R3500 VP.n43 VP.n42 24.4675
R3501 VP.n25 VP.n24 24.4675
R3502 VP.n25 VP.n20 24.4675
R3503 VP.n29 VP.n20 24.4675
R3504 VP.n54 VP.n53 20.5528
R3505 VP.n93 VP.n92 20.5528
R3506 VP.n50 VP.n49 20.5528
R3507 VP.n66 VP.n65 17.6167
R3508 VP.n81 VP.n80 17.6167
R3509 VP.n38 VP.n37 17.6167
R3510 VP.n67 VP.n66 6.85126
R3511 VP.n80 VP.n79 6.85126
R3512 VP.n37 VP.n36 6.85126
R3513 VP.n24 VP.n23 6.85126
R3514 VP.n22 VP.n21 2.67494
R3515 VP.n51 VP.n13 0.417535
R3516 VP.n52 VP.n12 0.417535
R3517 VP.n94 VP.n0 0.417535
R3518 VP VP.n94 0.394291
R3519 VP.n26 VP.n21 0.189894
R3520 VP.n27 VP.n26 0.189894
R3521 VP.n28 VP.n27 0.189894
R3522 VP.n28 VP.n19 0.189894
R3523 VP.n32 VP.n19 0.189894
R3524 VP.n33 VP.n32 0.189894
R3525 VP.n34 VP.n33 0.189894
R3526 VP.n34 VP.n17 0.189894
R3527 VP.n39 VP.n17 0.189894
R3528 VP.n40 VP.n39 0.189894
R3529 VP.n41 VP.n40 0.189894
R3530 VP.n41 VP.n15 0.189894
R3531 VP.n45 VP.n15 0.189894
R3532 VP.n46 VP.n45 0.189894
R3533 VP.n47 VP.n46 0.189894
R3534 VP.n47 VP.n13 0.189894
R3535 VP.n56 VP.n12 0.189894
R3536 VP.n57 VP.n56 0.189894
R3537 VP.n58 VP.n57 0.189894
R3538 VP.n58 VP.n10 0.189894
R3539 VP.n62 VP.n10 0.189894
R3540 VP.n63 VP.n62 0.189894
R3541 VP.n64 VP.n63 0.189894
R3542 VP.n64 VP.n8 0.189894
R3543 VP.n69 VP.n8 0.189894
R3544 VP.n70 VP.n69 0.189894
R3545 VP.n71 VP.n70 0.189894
R3546 VP.n71 VP.n6 0.189894
R3547 VP.n75 VP.n6 0.189894
R3548 VP.n76 VP.n75 0.189894
R3549 VP.n77 VP.n76 0.189894
R3550 VP.n77 VP.n4 0.189894
R3551 VP.n82 VP.n4 0.189894
R3552 VP.n83 VP.n82 0.189894
R3553 VP.n84 VP.n83 0.189894
R3554 VP.n84 VP.n2 0.189894
R3555 VP.n88 VP.n2 0.189894
R3556 VP.n89 VP.n88 0.189894
R3557 VP.n90 VP.n89 0.189894
R3558 VP.n90 VP.n0 0.189894
R3559 VDD1 VDD1.n0 62.5516
R3560 VDD1.n3 VDD1.n2 62.4379
R3561 VDD1.n3 VDD1.n1 62.4379
R3562 VDD1.n5 VDD1.n4 60.6485
R3563 VDD1.n5 VDD1.n3 54.1345
R3564 VDD1 VDD1.n5 1.78714
R3565 VDD1.n4 VDD1.t7 1.2904
R3566 VDD1.n4 VDD1.t5 1.2904
R3567 VDD1.n0 VDD1.t3 1.2904
R3568 VDD1.n0 VDD1.t1 1.2904
R3569 VDD1.n2 VDD1.t0 1.2904
R3570 VDD1.n2 VDD1.t2 1.2904
R3571 VDD1.n1 VDD1.t4 1.2904
R3572 VDD1.n1 VDD1.t6 1.2904
C0 VN VDD1 0.154322f
C1 VP VDD2 0.663478f
C2 VTAIL VDD1 9.611821f
C3 VN VDD2 11.767f
C4 VP VN 9.937309f
C5 VDD2 VTAIL 9.675281f
C6 VP VTAIL 12.4769f
C7 VDD2 VDD1 2.47962f
C8 VP VDD1 12.274f
C9 VN VTAIL 12.4628f
C10 VDD2 B 7.00494f
C11 VDD1 B 7.585299f
C12 VTAIL B 13.413213f
C13 VN B 20.993052f
C14 VP B 19.63601f
C15 VDD1.t3 B 0.32997f
C16 VDD1.t1 B 0.32997f
C17 VDD1.n0 B 3.00748f
C18 VDD1.t4 B 0.32997f
C19 VDD1.t6 B 0.32997f
C20 VDD1.n1 B 3.00591f
C21 VDD1.t0 B 0.32997f
C22 VDD1.t2 B 0.32997f
C23 VDD1.n2 B 3.00591f
C24 VDD1.n3 B 4.70082f
C25 VDD1.t7 B 0.32997f
C26 VDD1.t5 B 0.32997f
C27 VDD1.n4 B 2.98542f
C28 VDD1.n5 B 4.02866f
C29 VP.n0 B 0.030973f
C30 VP.t5 B 2.73717f
C31 VP.n1 B 0.030689f
C32 VP.n2 B 0.016466f
C33 VP.n3 B 0.030689f
C34 VP.n4 B 0.016466f
C35 VP.t7 B 2.73717f
C36 VP.n5 B 0.030689f
C37 VP.n6 B 0.016466f
C38 VP.n7 B 0.030689f
C39 VP.n8 B 0.016466f
C40 VP.t1 B 2.73717f
C41 VP.n9 B 0.030689f
C42 VP.n10 B 0.016466f
C43 VP.n11 B 0.030689f
C44 VP.n12 B 0.030973f
C45 VP.t3 B 2.73717f
C46 VP.n13 B 0.030973f
C47 VP.t2 B 2.73717f
C48 VP.n14 B 0.030689f
C49 VP.n15 B 0.016466f
C50 VP.n16 B 0.030689f
C51 VP.n17 B 0.016466f
C52 VP.t0 B 2.73717f
C53 VP.n18 B 0.030689f
C54 VP.n19 B 0.016466f
C55 VP.n20 B 0.030689f
C56 VP.n21 B 0.218971f
C57 VP.t6 B 2.73717f
C58 VP.t4 B 3.0132f
C59 VP.n22 B 0.957414f
C60 VP.n23 B 1.00454f
C61 VP.n24 B 0.01978f
C62 VP.n25 B 0.030689f
C63 VP.n26 B 0.016466f
C64 VP.n27 B 0.016466f
C65 VP.n28 B 0.016466f
C66 VP.n29 B 0.032726f
C67 VP.n30 B 0.013311f
C68 VP.n31 B 0.032726f
C69 VP.n32 B 0.016466f
C70 VP.n33 B 0.016466f
C71 VP.n34 B 0.016466f
C72 VP.n35 B 0.030689f
C73 VP.n36 B 0.01978f
C74 VP.n37 B 0.947795f
C75 VP.n38 B 0.026446f
C76 VP.n39 B 0.016466f
C77 VP.n40 B 0.016466f
C78 VP.n41 B 0.016466f
C79 VP.n42 B 0.030689f
C80 VP.n43 B 0.025414f
C81 VP.n44 B 0.022661f
C82 VP.n45 B 0.016466f
C83 VP.n46 B 0.016466f
C84 VP.n47 B 0.016466f
C85 VP.n48 B 0.030689f
C86 VP.n49 B 0.028265f
C87 VP.n50 B 1.02007f
C88 VP.n51 B 1.22697f
C89 VP.n52 B 1.23684f
C90 VP.n53 B 1.02007f
C91 VP.n54 B 0.028265f
C92 VP.n55 B 0.030689f
C93 VP.n56 B 0.016466f
C94 VP.n57 B 0.016466f
C95 VP.n58 B 0.016466f
C96 VP.n59 B 0.022661f
C97 VP.n60 B 0.025414f
C98 VP.n61 B 0.030689f
C99 VP.n62 B 0.016466f
C100 VP.n63 B 0.016466f
C101 VP.n64 B 0.016466f
C102 VP.n65 B 0.026446f
C103 VP.n66 B 0.947795f
C104 VP.n67 B 0.01978f
C105 VP.n68 B 0.030689f
C106 VP.n69 B 0.016466f
C107 VP.n70 B 0.016466f
C108 VP.n71 B 0.016466f
C109 VP.n72 B 0.032726f
C110 VP.n73 B 0.013311f
C111 VP.n74 B 0.032726f
C112 VP.n75 B 0.016466f
C113 VP.n76 B 0.016466f
C114 VP.n77 B 0.016466f
C115 VP.n78 B 0.030689f
C116 VP.n79 B 0.01978f
C117 VP.n80 B 0.947795f
C118 VP.n81 B 0.026446f
C119 VP.n82 B 0.016466f
C120 VP.n83 B 0.016466f
C121 VP.n84 B 0.016466f
C122 VP.n85 B 0.030689f
C123 VP.n86 B 0.025414f
C124 VP.n87 B 0.022661f
C125 VP.n88 B 0.016466f
C126 VP.n89 B 0.016466f
C127 VP.n90 B 0.016466f
C128 VP.n91 B 0.030689f
C129 VP.n92 B 0.028265f
C130 VP.n93 B 1.02007f
C131 VP.n94 B 0.052031f
C132 VTAIL.t8 B 0.241004f
C133 VTAIL.t7 B 0.241004f
C134 VTAIL.n0 B 2.12f
C135 VTAIL.n1 B 0.436679f
C136 VTAIL.n2 B 0.025648f
C137 VTAIL.n3 B 0.019868f
C138 VTAIL.n4 B 0.010676f
C139 VTAIL.n5 B 0.025235f
C140 VTAIL.n6 B 0.01099f
C141 VTAIL.n7 B 0.019868f
C142 VTAIL.n8 B 0.011304f
C143 VTAIL.n9 B 0.025235f
C144 VTAIL.n10 B 0.011304f
C145 VTAIL.n11 B 0.019868f
C146 VTAIL.n12 B 0.010676f
C147 VTAIL.n13 B 0.025235f
C148 VTAIL.n14 B 0.011304f
C149 VTAIL.n15 B 0.019868f
C150 VTAIL.n16 B 0.010676f
C151 VTAIL.n17 B 0.025235f
C152 VTAIL.n18 B 0.011304f
C153 VTAIL.n19 B 0.019868f
C154 VTAIL.n20 B 0.010676f
C155 VTAIL.n21 B 0.025235f
C156 VTAIL.n22 B 0.011304f
C157 VTAIL.n23 B 0.019868f
C158 VTAIL.n24 B 0.010676f
C159 VTAIL.n25 B 0.025235f
C160 VTAIL.n26 B 0.011304f
C161 VTAIL.n27 B 1.32454f
C162 VTAIL.n28 B 0.010676f
C163 VTAIL.t11 B 0.041634f
C164 VTAIL.n29 B 0.131329f
C165 VTAIL.n30 B 0.014907f
C166 VTAIL.n31 B 0.018926f
C167 VTAIL.n32 B 0.025235f
C168 VTAIL.n33 B 0.011304f
C169 VTAIL.n34 B 0.010676f
C170 VTAIL.n35 B 0.019868f
C171 VTAIL.n36 B 0.019868f
C172 VTAIL.n37 B 0.010676f
C173 VTAIL.n38 B 0.011304f
C174 VTAIL.n39 B 0.025235f
C175 VTAIL.n40 B 0.025235f
C176 VTAIL.n41 B 0.011304f
C177 VTAIL.n42 B 0.010676f
C178 VTAIL.n43 B 0.019868f
C179 VTAIL.n44 B 0.019868f
C180 VTAIL.n45 B 0.010676f
C181 VTAIL.n46 B 0.011304f
C182 VTAIL.n47 B 0.025235f
C183 VTAIL.n48 B 0.025235f
C184 VTAIL.n49 B 0.011304f
C185 VTAIL.n50 B 0.010676f
C186 VTAIL.n51 B 0.019868f
C187 VTAIL.n52 B 0.019868f
C188 VTAIL.n53 B 0.010676f
C189 VTAIL.n54 B 0.011304f
C190 VTAIL.n55 B 0.025235f
C191 VTAIL.n56 B 0.025235f
C192 VTAIL.n57 B 0.011304f
C193 VTAIL.n58 B 0.010676f
C194 VTAIL.n59 B 0.019868f
C195 VTAIL.n60 B 0.019868f
C196 VTAIL.n61 B 0.010676f
C197 VTAIL.n62 B 0.011304f
C198 VTAIL.n63 B 0.025235f
C199 VTAIL.n64 B 0.025235f
C200 VTAIL.n65 B 0.011304f
C201 VTAIL.n66 B 0.010676f
C202 VTAIL.n67 B 0.019868f
C203 VTAIL.n68 B 0.019868f
C204 VTAIL.n69 B 0.010676f
C205 VTAIL.n70 B 0.010676f
C206 VTAIL.n71 B 0.011304f
C207 VTAIL.n72 B 0.025235f
C208 VTAIL.n73 B 0.025235f
C209 VTAIL.n74 B 0.025235f
C210 VTAIL.n75 B 0.01099f
C211 VTAIL.n76 B 0.010676f
C212 VTAIL.n77 B 0.019868f
C213 VTAIL.n78 B 0.019868f
C214 VTAIL.n79 B 0.010676f
C215 VTAIL.n80 B 0.011304f
C216 VTAIL.n81 B 0.025235f
C217 VTAIL.n82 B 0.0506f
C218 VTAIL.n83 B 0.011304f
C219 VTAIL.n84 B 0.010676f
C220 VTAIL.n85 B 0.045653f
C221 VTAIL.n86 B 0.02789f
C222 VTAIL.n87 B 0.283108f
C223 VTAIL.n88 B 0.025648f
C224 VTAIL.n89 B 0.019868f
C225 VTAIL.n90 B 0.010676f
C226 VTAIL.n91 B 0.025235f
C227 VTAIL.n92 B 0.01099f
C228 VTAIL.n93 B 0.019868f
C229 VTAIL.n94 B 0.011304f
C230 VTAIL.n95 B 0.025235f
C231 VTAIL.n96 B 0.011304f
C232 VTAIL.n97 B 0.019868f
C233 VTAIL.n98 B 0.010676f
C234 VTAIL.n99 B 0.025235f
C235 VTAIL.n100 B 0.011304f
C236 VTAIL.n101 B 0.019868f
C237 VTAIL.n102 B 0.010676f
C238 VTAIL.n103 B 0.025235f
C239 VTAIL.n104 B 0.011304f
C240 VTAIL.n105 B 0.019868f
C241 VTAIL.n106 B 0.010676f
C242 VTAIL.n107 B 0.025235f
C243 VTAIL.n108 B 0.011304f
C244 VTAIL.n109 B 0.019868f
C245 VTAIL.n110 B 0.010676f
C246 VTAIL.n111 B 0.025235f
C247 VTAIL.n112 B 0.011304f
C248 VTAIL.n113 B 1.32454f
C249 VTAIL.n114 B 0.010676f
C250 VTAIL.t3 B 0.041634f
C251 VTAIL.n115 B 0.131329f
C252 VTAIL.n116 B 0.014907f
C253 VTAIL.n117 B 0.018926f
C254 VTAIL.n118 B 0.025235f
C255 VTAIL.n119 B 0.011304f
C256 VTAIL.n120 B 0.010676f
C257 VTAIL.n121 B 0.019868f
C258 VTAIL.n122 B 0.019868f
C259 VTAIL.n123 B 0.010676f
C260 VTAIL.n124 B 0.011304f
C261 VTAIL.n125 B 0.025235f
C262 VTAIL.n126 B 0.025235f
C263 VTAIL.n127 B 0.011304f
C264 VTAIL.n128 B 0.010676f
C265 VTAIL.n129 B 0.019868f
C266 VTAIL.n130 B 0.019868f
C267 VTAIL.n131 B 0.010676f
C268 VTAIL.n132 B 0.011304f
C269 VTAIL.n133 B 0.025235f
C270 VTAIL.n134 B 0.025235f
C271 VTAIL.n135 B 0.011304f
C272 VTAIL.n136 B 0.010676f
C273 VTAIL.n137 B 0.019868f
C274 VTAIL.n138 B 0.019868f
C275 VTAIL.n139 B 0.010676f
C276 VTAIL.n140 B 0.011304f
C277 VTAIL.n141 B 0.025235f
C278 VTAIL.n142 B 0.025235f
C279 VTAIL.n143 B 0.011304f
C280 VTAIL.n144 B 0.010676f
C281 VTAIL.n145 B 0.019868f
C282 VTAIL.n146 B 0.019868f
C283 VTAIL.n147 B 0.010676f
C284 VTAIL.n148 B 0.011304f
C285 VTAIL.n149 B 0.025235f
C286 VTAIL.n150 B 0.025235f
C287 VTAIL.n151 B 0.011304f
C288 VTAIL.n152 B 0.010676f
C289 VTAIL.n153 B 0.019868f
C290 VTAIL.n154 B 0.019868f
C291 VTAIL.n155 B 0.010676f
C292 VTAIL.n156 B 0.010676f
C293 VTAIL.n157 B 0.011304f
C294 VTAIL.n158 B 0.025235f
C295 VTAIL.n159 B 0.025235f
C296 VTAIL.n160 B 0.025235f
C297 VTAIL.n161 B 0.01099f
C298 VTAIL.n162 B 0.010676f
C299 VTAIL.n163 B 0.019868f
C300 VTAIL.n164 B 0.019868f
C301 VTAIL.n165 B 0.010676f
C302 VTAIL.n166 B 0.011304f
C303 VTAIL.n167 B 0.025235f
C304 VTAIL.n168 B 0.0506f
C305 VTAIL.n169 B 0.011304f
C306 VTAIL.n170 B 0.010676f
C307 VTAIL.n171 B 0.045653f
C308 VTAIL.n172 B 0.02789f
C309 VTAIL.n173 B 0.283108f
C310 VTAIL.t5 B 0.241004f
C311 VTAIL.t2 B 0.241004f
C312 VTAIL.n174 B 2.12f
C313 VTAIL.n175 B 0.669167f
C314 VTAIL.n176 B 0.025648f
C315 VTAIL.n177 B 0.019868f
C316 VTAIL.n178 B 0.010676f
C317 VTAIL.n179 B 0.025235f
C318 VTAIL.n180 B 0.01099f
C319 VTAIL.n181 B 0.019868f
C320 VTAIL.n182 B 0.011304f
C321 VTAIL.n183 B 0.025235f
C322 VTAIL.n184 B 0.011304f
C323 VTAIL.n185 B 0.019868f
C324 VTAIL.n186 B 0.010676f
C325 VTAIL.n187 B 0.025235f
C326 VTAIL.n188 B 0.011304f
C327 VTAIL.n189 B 0.019868f
C328 VTAIL.n190 B 0.010676f
C329 VTAIL.n191 B 0.025235f
C330 VTAIL.n192 B 0.011304f
C331 VTAIL.n193 B 0.019868f
C332 VTAIL.n194 B 0.010676f
C333 VTAIL.n195 B 0.025235f
C334 VTAIL.n196 B 0.011304f
C335 VTAIL.n197 B 0.019868f
C336 VTAIL.n198 B 0.010676f
C337 VTAIL.n199 B 0.025235f
C338 VTAIL.n200 B 0.011304f
C339 VTAIL.n201 B 1.32454f
C340 VTAIL.n202 B 0.010676f
C341 VTAIL.t6 B 0.041634f
C342 VTAIL.n203 B 0.131329f
C343 VTAIL.n204 B 0.014907f
C344 VTAIL.n205 B 0.018926f
C345 VTAIL.n206 B 0.025235f
C346 VTAIL.n207 B 0.011304f
C347 VTAIL.n208 B 0.010676f
C348 VTAIL.n209 B 0.019868f
C349 VTAIL.n210 B 0.019868f
C350 VTAIL.n211 B 0.010676f
C351 VTAIL.n212 B 0.011304f
C352 VTAIL.n213 B 0.025235f
C353 VTAIL.n214 B 0.025235f
C354 VTAIL.n215 B 0.011304f
C355 VTAIL.n216 B 0.010676f
C356 VTAIL.n217 B 0.019868f
C357 VTAIL.n218 B 0.019868f
C358 VTAIL.n219 B 0.010676f
C359 VTAIL.n220 B 0.011304f
C360 VTAIL.n221 B 0.025235f
C361 VTAIL.n222 B 0.025235f
C362 VTAIL.n223 B 0.011304f
C363 VTAIL.n224 B 0.010676f
C364 VTAIL.n225 B 0.019868f
C365 VTAIL.n226 B 0.019868f
C366 VTAIL.n227 B 0.010676f
C367 VTAIL.n228 B 0.011304f
C368 VTAIL.n229 B 0.025235f
C369 VTAIL.n230 B 0.025235f
C370 VTAIL.n231 B 0.011304f
C371 VTAIL.n232 B 0.010676f
C372 VTAIL.n233 B 0.019868f
C373 VTAIL.n234 B 0.019868f
C374 VTAIL.n235 B 0.010676f
C375 VTAIL.n236 B 0.011304f
C376 VTAIL.n237 B 0.025235f
C377 VTAIL.n238 B 0.025235f
C378 VTAIL.n239 B 0.011304f
C379 VTAIL.n240 B 0.010676f
C380 VTAIL.n241 B 0.019868f
C381 VTAIL.n242 B 0.019868f
C382 VTAIL.n243 B 0.010676f
C383 VTAIL.n244 B 0.010676f
C384 VTAIL.n245 B 0.011304f
C385 VTAIL.n246 B 0.025235f
C386 VTAIL.n247 B 0.025235f
C387 VTAIL.n248 B 0.025235f
C388 VTAIL.n249 B 0.01099f
C389 VTAIL.n250 B 0.010676f
C390 VTAIL.n251 B 0.019868f
C391 VTAIL.n252 B 0.019868f
C392 VTAIL.n253 B 0.010676f
C393 VTAIL.n254 B 0.011304f
C394 VTAIL.n255 B 0.025235f
C395 VTAIL.n256 B 0.0506f
C396 VTAIL.n257 B 0.011304f
C397 VTAIL.n258 B 0.010676f
C398 VTAIL.n259 B 0.045653f
C399 VTAIL.n260 B 0.02789f
C400 VTAIL.n261 B 1.6063f
C401 VTAIL.n262 B 0.025648f
C402 VTAIL.n263 B 0.019868f
C403 VTAIL.n264 B 0.010676f
C404 VTAIL.n265 B 0.025235f
C405 VTAIL.n266 B 0.01099f
C406 VTAIL.n267 B 0.019868f
C407 VTAIL.n268 B 0.01099f
C408 VTAIL.n269 B 0.010676f
C409 VTAIL.n270 B 0.025235f
C410 VTAIL.n271 B 0.025235f
C411 VTAIL.n272 B 0.011304f
C412 VTAIL.n273 B 0.019868f
C413 VTAIL.n274 B 0.010676f
C414 VTAIL.n275 B 0.025235f
C415 VTAIL.n276 B 0.011304f
C416 VTAIL.n277 B 0.019868f
C417 VTAIL.n278 B 0.010676f
C418 VTAIL.n279 B 0.025235f
C419 VTAIL.n280 B 0.011304f
C420 VTAIL.n281 B 0.019868f
C421 VTAIL.n282 B 0.010676f
C422 VTAIL.n283 B 0.025235f
C423 VTAIL.n284 B 0.011304f
C424 VTAIL.n285 B 0.019868f
C425 VTAIL.n286 B 0.010676f
C426 VTAIL.n287 B 0.025235f
C427 VTAIL.n288 B 0.011304f
C428 VTAIL.n289 B 1.32454f
C429 VTAIL.n290 B 0.010676f
C430 VTAIL.t13 B 0.041634f
C431 VTAIL.n291 B 0.131329f
C432 VTAIL.n292 B 0.014907f
C433 VTAIL.n293 B 0.018926f
C434 VTAIL.n294 B 0.025235f
C435 VTAIL.n295 B 0.011304f
C436 VTAIL.n296 B 0.010676f
C437 VTAIL.n297 B 0.019868f
C438 VTAIL.n298 B 0.019868f
C439 VTAIL.n299 B 0.010676f
C440 VTAIL.n300 B 0.011304f
C441 VTAIL.n301 B 0.025235f
C442 VTAIL.n302 B 0.025235f
C443 VTAIL.n303 B 0.011304f
C444 VTAIL.n304 B 0.010676f
C445 VTAIL.n305 B 0.019868f
C446 VTAIL.n306 B 0.019868f
C447 VTAIL.n307 B 0.010676f
C448 VTAIL.n308 B 0.011304f
C449 VTAIL.n309 B 0.025235f
C450 VTAIL.n310 B 0.025235f
C451 VTAIL.n311 B 0.011304f
C452 VTAIL.n312 B 0.010676f
C453 VTAIL.n313 B 0.019868f
C454 VTAIL.n314 B 0.019868f
C455 VTAIL.n315 B 0.010676f
C456 VTAIL.n316 B 0.011304f
C457 VTAIL.n317 B 0.025235f
C458 VTAIL.n318 B 0.025235f
C459 VTAIL.n319 B 0.011304f
C460 VTAIL.n320 B 0.010676f
C461 VTAIL.n321 B 0.019868f
C462 VTAIL.n322 B 0.019868f
C463 VTAIL.n323 B 0.010676f
C464 VTAIL.n324 B 0.011304f
C465 VTAIL.n325 B 0.025235f
C466 VTAIL.n326 B 0.025235f
C467 VTAIL.n327 B 0.011304f
C468 VTAIL.n328 B 0.010676f
C469 VTAIL.n329 B 0.019868f
C470 VTAIL.n330 B 0.019868f
C471 VTAIL.n331 B 0.010676f
C472 VTAIL.n332 B 0.011304f
C473 VTAIL.n333 B 0.025235f
C474 VTAIL.n334 B 0.025235f
C475 VTAIL.n335 B 0.011304f
C476 VTAIL.n336 B 0.010676f
C477 VTAIL.n337 B 0.019868f
C478 VTAIL.n338 B 0.019868f
C479 VTAIL.n339 B 0.010676f
C480 VTAIL.n340 B 0.011304f
C481 VTAIL.n341 B 0.025235f
C482 VTAIL.n342 B 0.0506f
C483 VTAIL.n343 B 0.011304f
C484 VTAIL.n344 B 0.010676f
C485 VTAIL.n345 B 0.045653f
C486 VTAIL.n346 B 0.02789f
C487 VTAIL.n347 B 1.6063f
C488 VTAIL.t9 B 0.241004f
C489 VTAIL.t14 B 0.241004f
C490 VTAIL.n348 B 2.12001f
C491 VTAIL.n349 B 0.669157f
C492 VTAIL.n350 B 0.025648f
C493 VTAIL.n351 B 0.019868f
C494 VTAIL.n352 B 0.010676f
C495 VTAIL.n353 B 0.025235f
C496 VTAIL.n354 B 0.01099f
C497 VTAIL.n355 B 0.019868f
C498 VTAIL.n356 B 0.01099f
C499 VTAIL.n357 B 0.010676f
C500 VTAIL.n358 B 0.025235f
C501 VTAIL.n359 B 0.025235f
C502 VTAIL.n360 B 0.011304f
C503 VTAIL.n361 B 0.019868f
C504 VTAIL.n362 B 0.010676f
C505 VTAIL.n363 B 0.025235f
C506 VTAIL.n364 B 0.011304f
C507 VTAIL.n365 B 0.019868f
C508 VTAIL.n366 B 0.010676f
C509 VTAIL.n367 B 0.025235f
C510 VTAIL.n368 B 0.011304f
C511 VTAIL.n369 B 0.019868f
C512 VTAIL.n370 B 0.010676f
C513 VTAIL.n371 B 0.025235f
C514 VTAIL.n372 B 0.011304f
C515 VTAIL.n373 B 0.019868f
C516 VTAIL.n374 B 0.010676f
C517 VTAIL.n375 B 0.025235f
C518 VTAIL.n376 B 0.011304f
C519 VTAIL.n377 B 1.32454f
C520 VTAIL.n378 B 0.010676f
C521 VTAIL.t10 B 0.041634f
C522 VTAIL.n379 B 0.131329f
C523 VTAIL.n380 B 0.014907f
C524 VTAIL.n381 B 0.018926f
C525 VTAIL.n382 B 0.025235f
C526 VTAIL.n383 B 0.011304f
C527 VTAIL.n384 B 0.010676f
C528 VTAIL.n385 B 0.019868f
C529 VTAIL.n386 B 0.019868f
C530 VTAIL.n387 B 0.010676f
C531 VTAIL.n388 B 0.011304f
C532 VTAIL.n389 B 0.025235f
C533 VTAIL.n390 B 0.025235f
C534 VTAIL.n391 B 0.011304f
C535 VTAIL.n392 B 0.010676f
C536 VTAIL.n393 B 0.019868f
C537 VTAIL.n394 B 0.019868f
C538 VTAIL.n395 B 0.010676f
C539 VTAIL.n396 B 0.011304f
C540 VTAIL.n397 B 0.025235f
C541 VTAIL.n398 B 0.025235f
C542 VTAIL.n399 B 0.011304f
C543 VTAIL.n400 B 0.010676f
C544 VTAIL.n401 B 0.019868f
C545 VTAIL.n402 B 0.019868f
C546 VTAIL.n403 B 0.010676f
C547 VTAIL.n404 B 0.011304f
C548 VTAIL.n405 B 0.025235f
C549 VTAIL.n406 B 0.025235f
C550 VTAIL.n407 B 0.011304f
C551 VTAIL.n408 B 0.010676f
C552 VTAIL.n409 B 0.019868f
C553 VTAIL.n410 B 0.019868f
C554 VTAIL.n411 B 0.010676f
C555 VTAIL.n412 B 0.011304f
C556 VTAIL.n413 B 0.025235f
C557 VTAIL.n414 B 0.025235f
C558 VTAIL.n415 B 0.011304f
C559 VTAIL.n416 B 0.010676f
C560 VTAIL.n417 B 0.019868f
C561 VTAIL.n418 B 0.019868f
C562 VTAIL.n419 B 0.010676f
C563 VTAIL.n420 B 0.011304f
C564 VTAIL.n421 B 0.025235f
C565 VTAIL.n422 B 0.025235f
C566 VTAIL.n423 B 0.011304f
C567 VTAIL.n424 B 0.010676f
C568 VTAIL.n425 B 0.019868f
C569 VTAIL.n426 B 0.019868f
C570 VTAIL.n427 B 0.010676f
C571 VTAIL.n428 B 0.011304f
C572 VTAIL.n429 B 0.025235f
C573 VTAIL.n430 B 0.0506f
C574 VTAIL.n431 B 0.011304f
C575 VTAIL.n432 B 0.010676f
C576 VTAIL.n433 B 0.045653f
C577 VTAIL.n434 B 0.02789f
C578 VTAIL.n435 B 0.283108f
C579 VTAIL.n436 B 0.025648f
C580 VTAIL.n437 B 0.019868f
C581 VTAIL.n438 B 0.010676f
C582 VTAIL.n439 B 0.025235f
C583 VTAIL.n440 B 0.01099f
C584 VTAIL.n441 B 0.019868f
C585 VTAIL.n442 B 0.01099f
C586 VTAIL.n443 B 0.010676f
C587 VTAIL.n444 B 0.025235f
C588 VTAIL.n445 B 0.025235f
C589 VTAIL.n446 B 0.011304f
C590 VTAIL.n447 B 0.019868f
C591 VTAIL.n448 B 0.010676f
C592 VTAIL.n449 B 0.025235f
C593 VTAIL.n450 B 0.011304f
C594 VTAIL.n451 B 0.019868f
C595 VTAIL.n452 B 0.010676f
C596 VTAIL.n453 B 0.025235f
C597 VTAIL.n454 B 0.011304f
C598 VTAIL.n455 B 0.019868f
C599 VTAIL.n456 B 0.010676f
C600 VTAIL.n457 B 0.025235f
C601 VTAIL.n458 B 0.011304f
C602 VTAIL.n459 B 0.019868f
C603 VTAIL.n460 B 0.010676f
C604 VTAIL.n461 B 0.025235f
C605 VTAIL.n462 B 0.011304f
C606 VTAIL.n463 B 1.32454f
C607 VTAIL.n464 B 0.010676f
C608 VTAIL.t4 B 0.041634f
C609 VTAIL.n465 B 0.131329f
C610 VTAIL.n466 B 0.014907f
C611 VTAIL.n467 B 0.018926f
C612 VTAIL.n468 B 0.025235f
C613 VTAIL.n469 B 0.011304f
C614 VTAIL.n470 B 0.010676f
C615 VTAIL.n471 B 0.019868f
C616 VTAIL.n472 B 0.019868f
C617 VTAIL.n473 B 0.010676f
C618 VTAIL.n474 B 0.011304f
C619 VTAIL.n475 B 0.025235f
C620 VTAIL.n476 B 0.025235f
C621 VTAIL.n477 B 0.011304f
C622 VTAIL.n478 B 0.010676f
C623 VTAIL.n479 B 0.019868f
C624 VTAIL.n480 B 0.019868f
C625 VTAIL.n481 B 0.010676f
C626 VTAIL.n482 B 0.011304f
C627 VTAIL.n483 B 0.025235f
C628 VTAIL.n484 B 0.025235f
C629 VTAIL.n485 B 0.011304f
C630 VTAIL.n486 B 0.010676f
C631 VTAIL.n487 B 0.019868f
C632 VTAIL.n488 B 0.019868f
C633 VTAIL.n489 B 0.010676f
C634 VTAIL.n490 B 0.011304f
C635 VTAIL.n491 B 0.025235f
C636 VTAIL.n492 B 0.025235f
C637 VTAIL.n493 B 0.011304f
C638 VTAIL.n494 B 0.010676f
C639 VTAIL.n495 B 0.019868f
C640 VTAIL.n496 B 0.019868f
C641 VTAIL.n497 B 0.010676f
C642 VTAIL.n498 B 0.011304f
C643 VTAIL.n499 B 0.025235f
C644 VTAIL.n500 B 0.025235f
C645 VTAIL.n501 B 0.011304f
C646 VTAIL.n502 B 0.010676f
C647 VTAIL.n503 B 0.019868f
C648 VTAIL.n504 B 0.019868f
C649 VTAIL.n505 B 0.010676f
C650 VTAIL.n506 B 0.011304f
C651 VTAIL.n507 B 0.025235f
C652 VTAIL.n508 B 0.025235f
C653 VTAIL.n509 B 0.011304f
C654 VTAIL.n510 B 0.010676f
C655 VTAIL.n511 B 0.019868f
C656 VTAIL.n512 B 0.019868f
C657 VTAIL.n513 B 0.010676f
C658 VTAIL.n514 B 0.011304f
C659 VTAIL.n515 B 0.025235f
C660 VTAIL.n516 B 0.0506f
C661 VTAIL.n517 B 0.011304f
C662 VTAIL.n518 B 0.010676f
C663 VTAIL.n519 B 0.045653f
C664 VTAIL.n520 B 0.02789f
C665 VTAIL.n521 B 0.283108f
C666 VTAIL.t15 B 0.241004f
C667 VTAIL.t1 B 0.241004f
C668 VTAIL.n522 B 2.12001f
C669 VTAIL.n523 B 0.669157f
C670 VTAIL.n524 B 0.025648f
C671 VTAIL.n525 B 0.019868f
C672 VTAIL.n526 B 0.010676f
C673 VTAIL.n527 B 0.025235f
C674 VTAIL.n528 B 0.01099f
C675 VTAIL.n529 B 0.019868f
C676 VTAIL.n530 B 0.01099f
C677 VTAIL.n531 B 0.010676f
C678 VTAIL.n532 B 0.025235f
C679 VTAIL.n533 B 0.025235f
C680 VTAIL.n534 B 0.011304f
C681 VTAIL.n535 B 0.019868f
C682 VTAIL.n536 B 0.010676f
C683 VTAIL.n537 B 0.025235f
C684 VTAIL.n538 B 0.011304f
C685 VTAIL.n539 B 0.019868f
C686 VTAIL.n540 B 0.010676f
C687 VTAIL.n541 B 0.025235f
C688 VTAIL.n542 B 0.011304f
C689 VTAIL.n543 B 0.019868f
C690 VTAIL.n544 B 0.010676f
C691 VTAIL.n545 B 0.025235f
C692 VTAIL.n546 B 0.011304f
C693 VTAIL.n547 B 0.019868f
C694 VTAIL.n548 B 0.010676f
C695 VTAIL.n549 B 0.025235f
C696 VTAIL.n550 B 0.011304f
C697 VTAIL.n551 B 1.32454f
C698 VTAIL.n552 B 0.010676f
C699 VTAIL.t0 B 0.041634f
C700 VTAIL.n553 B 0.131329f
C701 VTAIL.n554 B 0.014907f
C702 VTAIL.n555 B 0.018926f
C703 VTAIL.n556 B 0.025235f
C704 VTAIL.n557 B 0.011304f
C705 VTAIL.n558 B 0.010676f
C706 VTAIL.n559 B 0.019868f
C707 VTAIL.n560 B 0.019868f
C708 VTAIL.n561 B 0.010676f
C709 VTAIL.n562 B 0.011304f
C710 VTAIL.n563 B 0.025235f
C711 VTAIL.n564 B 0.025235f
C712 VTAIL.n565 B 0.011304f
C713 VTAIL.n566 B 0.010676f
C714 VTAIL.n567 B 0.019868f
C715 VTAIL.n568 B 0.019868f
C716 VTAIL.n569 B 0.010676f
C717 VTAIL.n570 B 0.011304f
C718 VTAIL.n571 B 0.025235f
C719 VTAIL.n572 B 0.025235f
C720 VTAIL.n573 B 0.011304f
C721 VTAIL.n574 B 0.010676f
C722 VTAIL.n575 B 0.019868f
C723 VTAIL.n576 B 0.019868f
C724 VTAIL.n577 B 0.010676f
C725 VTAIL.n578 B 0.011304f
C726 VTAIL.n579 B 0.025235f
C727 VTAIL.n580 B 0.025235f
C728 VTAIL.n581 B 0.011304f
C729 VTAIL.n582 B 0.010676f
C730 VTAIL.n583 B 0.019868f
C731 VTAIL.n584 B 0.019868f
C732 VTAIL.n585 B 0.010676f
C733 VTAIL.n586 B 0.011304f
C734 VTAIL.n587 B 0.025235f
C735 VTAIL.n588 B 0.025235f
C736 VTAIL.n589 B 0.011304f
C737 VTAIL.n590 B 0.010676f
C738 VTAIL.n591 B 0.019868f
C739 VTAIL.n592 B 0.019868f
C740 VTAIL.n593 B 0.010676f
C741 VTAIL.n594 B 0.011304f
C742 VTAIL.n595 B 0.025235f
C743 VTAIL.n596 B 0.025235f
C744 VTAIL.n597 B 0.011304f
C745 VTAIL.n598 B 0.010676f
C746 VTAIL.n599 B 0.019868f
C747 VTAIL.n600 B 0.019868f
C748 VTAIL.n601 B 0.010676f
C749 VTAIL.n602 B 0.011304f
C750 VTAIL.n603 B 0.025235f
C751 VTAIL.n604 B 0.0506f
C752 VTAIL.n605 B 0.011304f
C753 VTAIL.n606 B 0.010676f
C754 VTAIL.n607 B 0.045653f
C755 VTAIL.n608 B 0.02789f
C756 VTAIL.n609 B 1.6063f
C757 VTAIL.n610 B 0.025648f
C758 VTAIL.n611 B 0.019868f
C759 VTAIL.n612 B 0.010676f
C760 VTAIL.n613 B 0.025235f
C761 VTAIL.n614 B 0.01099f
C762 VTAIL.n615 B 0.019868f
C763 VTAIL.n616 B 0.011304f
C764 VTAIL.n617 B 0.025235f
C765 VTAIL.n618 B 0.011304f
C766 VTAIL.n619 B 0.019868f
C767 VTAIL.n620 B 0.010676f
C768 VTAIL.n621 B 0.025235f
C769 VTAIL.n622 B 0.011304f
C770 VTAIL.n623 B 0.019868f
C771 VTAIL.n624 B 0.010676f
C772 VTAIL.n625 B 0.025235f
C773 VTAIL.n626 B 0.011304f
C774 VTAIL.n627 B 0.019868f
C775 VTAIL.n628 B 0.010676f
C776 VTAIL.n629 B 0.025235f
C777 VTAIL.n630 B 0.011304f
C778 VTAIL.n631 B 0.019868f
C779 VTAIL.n632 B 0.010676f
C780 VTAIL.n633 B 0.025235f
C781 VTAIL.n634 B 0.011304f
C782 VTAIL.n635 B 1.32454f
C783 VTAIL.n636 B 0.010676f
C784 VTAIL.t12 B 0.041634f
C785 VTAIL.n637 B 0.131329f
C786 VTAIL.n638 B 0.014907f
C787 VTAIL.n639 B 0.018926f
C788 VTAIL.n640 B 0.025235f
C789 VTAIL.n641 B 0.011304f
C790 VTAIL.n642 B 0.010676f
C791 VTAIL.n643 B 0.019868f
C792 VTAIL.n644 B 0.019868f
C793 VTAIL.n645 B 0.010676f
C794 VTAIL.n646 B 0.011304f
C795 VTAIL.n647 B 0.025235f
C796 VTAIL.n648 B 0.025235f
C797 VTAIL.n649 B 0.011304f
C798 VTAIL.n650 B 0.010676f
C799 VTAIL.n651 B 0.019868f
C800 VTAIL.n652 B 0.019868f
C801 VTAIL.n653 B 0.010676f
C802 VTAIL.n654 B 0.011304f
C803 VTAIL.n655 B 0.025235f
C804 VTAIL.n656 B 0.025235f
C805 VTAIL.n657 B 0.011304f
C806 VTAIL.n658 B 0.010676f
C807 VTAIL.n659 B 0.019868f
C808 VTAIL.n660 B 0.019868f
C809 VTAIL.n661 B 0.010676f
C810 VTAIL.n662 B 0.011304f
C811 VTAIL.n663 B 0.025235f
C812 VTAIL.n664 B 0.025235f
C813 VTAIL.n665 B 0.011304f
C814 VTAIL.n666 B 0.010676f
C815 VTAIL.n667 B 0.019868f
C816 VTAIL.n668 B 0.019868f
C817 VTAIL.n669 B 0.010676f
C818 VTAIL.n670 B 0.011304f
C819 VTAIL.n671 B 0.025235f
C820 VTAIL.n672 B 0.025235f
C821 VTAIL.n673 B 0.011304f
C822 VTAIL.n674 B 0.010676f
C823 VTAIL.n675 B 0.019868f
C824 VTAIL.n676 B 0.019868f
C825 VTAIL.n677 B 0.010676f
C826 VTAIL.n678 B 0.010676f
C827 VTAIL.n679 B 0.011304f
C828 VTAIL.n680 B 0.025235f
C829 VTAIL.n681 B 0.025235f
C830 VTAIL.n682 B 0.025235f
C831 VTAIL.n683 B 0.01099f
C832 VTAIL.n684 B 0.010676f
C833 VTAIL.n685 B 0.019868f
C834 VTAIL.n686 B 0.019868f
C835 VTAIL.n687 B 0.010676f
C836 VTAIL.n688 B 0.011304f
C837 VTAIL.n689 B 0.025235f
C838 VTAIL.n690 B 0.0506f
C839 VTAIL.n691 B 0.011304f
C840 VTAIL.n692 B 0.010676f
C841 VTAIL.n693 B 0.045653f
C842 VTAIL.n694 B 0.02789f
C843 VTAIL.n695 B 1.60257f
C844 VDD2.t1 B 0.325903f
C845 VDD2.t2 B 0.325903f
C846 VDD2.n0 B 2.96886f
C847 VDD2.t4 B 0.325903f
C848 VDD2.t5 B 0.325903f
C849 VDD2.n1 B 2.96886f
C850 VDD2.n2 B 4.587759f
C851 VDD2.t6 B 0.325903f
C852 VDD2.t3 B 0.325903f
C853 VDD2.n3 B 2.94863f
C854 VDD2.n4 B 3.94494f
C855 VDD2.t7 B 0.325903f
C856 VDD2.t0 B 0.325903f
C857 VDD2.n5 B 2.96881f
C858 VN.n0 B 0.030506f
C859 VN.t2 B 2.69593f
C860 VN.n1 B 0.030226f
C861 VN.n2 B 0.016218f
C862 VN.n3 B 0.030226f
C863 VN.n4 B 0.016218f
C864 VN.t7 B 2.69593f
C865 VN.n5 B 0.030226f
C866 VN.n6 B 0.016218f
C867 VN.n7 B 0.030226f
C868 VN.n8 B 0.215671f
C869 VN.t6 B 2.69593f
C870 VN.t3 B 2.9678f
C871 VN.n9 B 0.942988f
C872 VN.n10 B 0.989404f
C873 VN.n11 B 0.019482f
C874 VN.n12 B 0.030226f
C875 VN.n13 B 0.016218f
C876 VN.n14 B 0.016218f
C877 VN.n15 B 0.016218f
C878 VN.n16 B 0.032233f
C879 VN.n17 B 0.013111f
C880 VN.n18 B 0.032233f
C881 VN.n19 B 0.016218f
C882 VN.n20 B 0.016218f
C883 VN.n21 B 0.016218f
C884 VN.n22 B 0.030226f
C885 VN.n23 B 0.019482f
C886 VN.n24 B 0.933515f
C887 VN.n25 B 0.026048f
C888 VN.n26 B 0.016218f
C889 VN.n27 B 0.016218f
C890 VN.n28 B 0.016218f
C891 VN.n29 B 0.030226f
C892 VN.n30 B 0.025031f
C893 VN.n31 B 0.02232f
C894 VN.n32 B 0.016218f
C895 VN.n33 B 0.016218f
C896 VN.n34 B 0.016218f
C897 VN.n35 B 0.030226f
C898 VN.n36 B 0.027839f
C899 VN.n37 B 1.0047f
C900 VN.n38 B 0.051247f
C901 VN.n39 B 0.030506f
C902 VN.t1 B 2.69593f
C903 VN.n40 B 0.030226f
C904 VN.n41 B 0.016218f
C905 VN.n42 B 0.030226f
C906 VN.n43 B 0.016218f
C907 VN.t5 B 2.69593f
C908 VN.n44 B 0.030226f
C909 VN.n45 B 0.016218f
C910 VN.n46 B 0.030226f
C911 VN.n47 B 0.215671f
C912 VN.t0 B 2.69593f
C913 VN.t4 B 2.9678f
C914 VN.n48 B 0.942988f
C915 VN.n49 B 0.989404f
C916 VN.n50 B 0.019482f
C917 VN.n51 B 0.030226f
C918 VN.n52 B 0.016218f
C919 VN.n53 B 0.016218f
C920 VN.n54 B 0.016218f
C921 VN.n55 B 0.032233f
C922 VN.n56 B 0.013111f
C923 VN.n57 B 0.032233f
C924 VN.n58 B 0.016218f
C925 VN.n59 B 0.016218f
C926 VN.n60 B 0.016218f
C927 VN.n61 B 0.030226f
C928 VN.n62 B 0.019482f
C929 VN.n63 B 0.933515f
C930 VN.n64 B 0.026048f
C931 VN.n65 B 0.016218f
C932 VN.n66 B 0.016218f
C933 VN.n67 B 0.016218f
C934 VN.n68 B 0.030226f
C935 VN.n69 B 0.025031f
C936 VN.n70 B 0.02232f
C937 VN.n71 B 0.016218f
C938 VN.n72 B 0.016218f
C939 VN.n73 B 0.016218f
C940 VN.n74 B 0.030226f
C941 VN.n75 B 0.027839f
C942 VN.n76 B 1.0047f
C943 VN.n77 B 1.21219f
.ends

