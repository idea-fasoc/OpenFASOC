* NGSPICE file created from diff_pair_sample_1523.ext - technology: sky130A

.subckt diff_pair_sample_1523 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VP.t0 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X1 VTAIL.t8 VN.t0 VDD2.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X2 VDD2.t8 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.1175 pd=37.28 as=3.01125 ps=18.58 w=18.25 l=1.41
X3 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1175 pd=37.28 as=0 ps=0 w=18.25 l=1.41
X4 VDD2.t7 VN.t2 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X5 VTAIL.t18 VP.t1 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X6 VTAIL.t7 VN.t3 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X7 VDD1.t7 VP.t2 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X8 VDD2.t5 VN.t4 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.1175 pd=37.28 as=3.01125 ps=18.58 w=18.25 l=1.41
X9 VTAIL.t3 VN.t5 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X10 VDD1.t6 VP.t3 VTAIL.t16 B.t2 sky130_fd_pr__nfet_01v8 ad=7.1175 pd=37.28 as=3.01125 ps=18.58 w=18.25 l=1.41
X11 VDD1.t9 VP.t4 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=7.1175 ps=37.28 w=18.25 l=1.41
X12 VTAIL.t1 VN.t6 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X13 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=7.1175 pd=37.28 as=0 ps=0 w=18.25 l=1.41
X14 VTAIL.t14 VP.t5 VDD1.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X15 VDD1.t5 VP.t6 VTAIL.t13 B.t6 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X16 VDD2.t2 VN.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=7.1175 ps=37.28 w=18.25 l=1.41
X17 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.1175 pd=37.28 as=0 ps=0 w=18.25 l=1.41
X18 VDD1.t4 VP.t7 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=7.1175 pd=37.28 as=3.01125 ps=18.58 w=18.25 l=1.41
X19 VDD2.t1 VN.t8 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=7.1175 ps=37.28 w=18.25 l=1.41
X20 VDD1.t3 VP.t8 VTAIL.t11 B.t9 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=7.1175 ps=37.28 w=18.25 l=1.41
X21 VDD2.t0 VN.t9 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X22 VTAIL.t10 VP.t9 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.01125 pd=18.58 as=3.01125 ps=18.58 w=18.25 l=1.41
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.1175 pd=37.28 as=0 ps=0 w=18.25 l=1.41
R0 VP.n14 VP.t3 346.658
R1 VP.n34 VP.t7 311.933
R2 VP.n5 VP.t1 311.933
R3 VP.n45 VP.t2 311.933
R4 VP.n52 VP.t5 311.933
R5 VP.n59 VP.t4 311.933
R6 VP.n32 VP.t8 311.933
R7 VP.n25 VP.t0 311.933
R8 VP.n18 VP.t6 311.933
R9 VP.n13 VP.t9 311.933
R10 VP.n35 VP.n34 174.512
R11 VP.n60 VP.n59 174.512
R12 VP.n33 VP.n32 174.512
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n12 161.3
R15 VP.n20 VP.n19 161.3
R16 VP.n21 VP.n11 161.3
R17 VP.n23 VP.n22 161.3
R18 VP.n24 VP.n10 161.3
R19 VP.n27 VP.n26 161.3
R20 VP.n28 VP.n9 161.3
R21 VP.n30 VP.n29 161.3
R22 VP.n31 VP.n8 161.3
R23 VP.n58 VP.n0 161.3
R24 VP.n57 VP.n56 161.3
R25 VP.n55 VP.n1 161.3
R26 VP.n54 VP.n53 161.3
R27 VP.n51 VP.n2 161.3
R28 VP.n50 VP.n49 161.3
R29 VP.n48 VP.n3 161.3
R30 VP.n47 VP.n46 161.3
R31 VP.n44 VP.n4 161.3
R32 VP.n43 VP.n42 161.3
R33 VP.n41 VP.n40 161.3
R34 VP.n39 VP.n6 161.3
R35 VP.n38 VP.n37 161.3
R36 VP.n36 VP.n7 161.3
R37 VP.n39 VP.n38 54.0911
R38 VP.n57 VP.n1 54.0911
R39 VP.n30 VP.n9 54.0911
R40 VP.n44 VP.n43 52.1486
R41 VP.n51 VP.n50 52.1486
R42 VP.n24 VP.n23 52.1486
R43 VP.n17 VP.n16 52.1486
R44 VP.n35 VP.n33 51.3035
R45 VP.n14 VP.n13 42.3338
R46 VP.n46 VP.n44 28.8382
R47 VP.n50 VP.n3 28.8382
R48 VP.n23 VP.n11 28.8382
R49 VP.n19 VP.n17 28.8382
R50 VP.n38 VP.n7 26.8957
R51 VP.n58 VP.n57 26.8957
R52 VP.n31 VP.n30 26.8957
R53 VP.n40 VP.n39 24.4675
R54 VP.n53 VP.n1 24.4675
R55 VP.n26 VP.n9 24.4675
R56 VP.n43 VP.n5 23.9782
R57 VP.n52 VP.n51 23.9782
R58 VP.n25 VP.n24 23.9782
R59 VP.n16 VP.n13 23.9782
R60 VP.n15 VP.n14 17.64
R61 VP.n46 VP.n45 12.234
R62 VP.n45 VP.n3 12.234
R63 VP.n19 VP.n18 12.234
R64 VP.n18 VP.n11 12.234
R65 VP.n34 VP.n7 11.2553
R66 VP.n59 VP.n58 11.2553
R67 VP.n32 VP.n31 11.2553
R68 VP.n40 VP.n5 0.48984
R69 VP.n53 VP.n52 0.48984
R70 VP.n26 VP.n25 0.48984
R71 VP.n15 VP.n12 0.189894
R72 VP.n20 VP.n12 0.189894
R73 VP.n21 VP.n20 0.189894
R74 VP.n22 VP.n21 0.189894
R75 VP.n22 VP.n10 0.189894
R76 VP.n27 VP.n10 0.189894
R77 VP.n28 VP.n27 0.189894
R78 VP.n29 VP.n28 0.189894
R79 VP.n29 VP.n8 0.189894
R80 VP.n33 VP.n8 0.189894
R81 VP.n36 VP.n35 0.189894
R82 VP.n37 VP.n36 0.189894
R83 VP.n37 VP.n6 0.189894
R84 VP.n41 VP.n6 0.189894
R85 VP.n42 VP.n41 0.189894
R86 VP.n42 VP.n4 0.189894
R87 VP.n47 VP.n4 0.189894
R88 VP.n48 VP.n47 0.189894
R89 VP.n49 VP.n48 0.189894
R90 VP.n49 VP.n2 0.189894
R91 VP.n54 VP.n2 0.189894
R92 VP.n55 VP.n54 0.189894
R93 VP.n56 VP.n55 0.189894
R94 VP.n56 VP.n0 0.189894
R95 VP.n60 VP.n0 0.189894
R96 VP VP.n60 0.0516364
R97 VDD1.n96 VDD1.n0 289.615
R98 VDD1.n199 VDD1.n103 289.615
R99 VDD1.n97 VDD1.n96 185
R100 VDD1.n95 VDD1.n94 185
R101 VDD1.n4 VDD1.n3 185
R102 VDD1.n89 VDD1.n88 185
R103 VDD1.n87 VDD1.n86 185
R104 VDD1.n8 VDD1.n7 185
R105 VDD1.n81 VDD1.n80 185
R106 VDD1.n79 VDD1.n10 185
R107 VDD1.n78 VDD1.n77 185
R108 VDD1.n13 VDD1.n11 185
R109 VDD1.n72 VDD1.n71 185
R110 VDD1.n70 VDD1.n69 185
R111 VDD1.n17 VDD1.n16 185
R112 VDD1.n64 VDD1.n63 185
R113 VDD1.n62 VDD1.n61 185
R114 VDD1.n21 VDD1.n20 185
R115 VDD1.n56 VDD1.n55 185
R116 VDD1.n54 VDD1.n53 185
R117 VDD1.n25 VDD1.n24 185
R118 VDD1.n48 VDD1.n47 185
R119 VDD1.n46 VDD1.n45 185
R120 VDD1.n29 VDD1.n28 185
R121 VDD1.n40 VDD1.n39 185
R122 VDD1.n38 VDD1.n37 185
R123 VDD1.n33 VDD1.n32 185
R124 VDD1.n135 VDD1.n134 185
R125 VDD1.n140 VDD1.n139 185
R126 VDD1.n142 VDD1.n141 185
R127 VDD1.n131 VDD1.n130 185
R128 VDD1.n148 VDD1.n147 185
R129 VDD1.n150 VDD1.n149 185
R130 VDD1.n127 VDD1.n126 185
R131 VDD1.n156 VDD1.n155 185
R132 VDD1.n158 VDD1.n157 185
R133 VDD1.n123 VDD1.n122 185
R134 VDD1.n164 VDD1.n163 185
R135 VDD1.n166 VDD1.n165 185
R136 VDD1.n119 VDD1.n118 185
R137 VDD1.n172 VDD1.n171 185
R138 VDD1.n174 VDD1.n173 185
R139 VDD1.n115 VDD1.n114 185
R140 VDD1.n181 VDD1.n180 185
R141 VDD1.n182 VDD1.n113 185
R142 VDD1.n184 VDD1.n183 185
R143 VDD1.n111 VDD1.n110 185
R144 VDD1.n190 VDD1.n189 185
R145 VDD1.n192 VDD1.n191 185
R146 VDD1.n107 VDD1.n106 185
R147 VDD1.n198 VDD1.n197 185
R148 VDD1.n200 VDD1.n199 185
R149 VDD1.n34 VDD1.t6 147.659
R150 VDD1.n136 VDD1.t4 147.659
R151 VDD1.n96 VDD1.n95 104.615
R152 VDD1.n95 VDD1.n3 104.615
R153 VDD1.n88 VDD1.n3 104.615
R154 VDD1.n88 VDD1.n87 104.615
R155 VDD1.n87 VDD1.n7 104.615
R156 VDD1.n80 VDD1.n7 104.615
R157 VDD1.n80 VDD1.n79 104.615
R158 VDD1.n79 VDD1.n78 104.615
R159 VDD1.n78 VDD1.n11 104.615
R160 VDD1.n71 VDD1.n11 104.615
R161 VDD1.n71 VDD1.n70 104.615
R162 VDD1.n70 VDD1.n16 104.615
R163 VDD1.n63 VDD1.n16 104.615
R164 VDD1.n63 VDD1.n62 104.615
R165 VDD1.n62 VDD1.n20 104.615
R166 VDD1.n55 VDD1.n20 104.615
R167 VDD1.n55 VDD1.n54 104.615
R168 VDD1.n54 VDD1.n24 104.615
R169 VDD1.n47 VDD1.n24 104.615
R170 VDD1.n47 VDD1.n46 104.615
R171 VDD1.n46 VDD1.n28 104.615
R172 VDD1.n39 VDD1.n28 104.615
R173 VDD1.n39 VDD1.n38 104.615
R174 VDD1.n38 VDD1.n32 104.615
R175 VDD1.n140 VDD1.n134 104.615
R176 VDD1.n141 VDD1.n140 104.615
R177 VDD1.n141 VDD1.n130 104.615
R178 VDD1.n148 VDD1.n130 104.615
R179 VDD1.n149 VDD1.n148 104.615
R180 VDD1.n149 VDD1.n126 104.615
R181 VDD1.n156 VDD1.n126 104.615
R182 VDD1.n157 VDD1.n156 104.615
R183 VDD1.n157 VDD1.n122 104.615
R184 VDD1.n164 VDD1.n122 104.615
R185 VDD1.n165 VDD1.n164 104.615
R186 VDD1.n165 VDD1.n118 104.615
R187 VDD1.n172 VDD1.n118 104.615
R188 VDD1.n173 VDD1.n172 104.615
R189 VDD1.n173 VDD1.n114 104.615
R190 VDD1.n181 VDD1.n114 104.615
R191 VDD1.n182 VDD1.n181 104.615
R192 VDD1.n183 VDD1.n182 104.615
R193 VDD1.n183 VDD1.n110 104.615
R194 VDD1.n190 VDD1.n110 104.615
R195 VDD1.n191 VDD1.n190 104.615
R196 VDD1.n191 VDD1.n106 104.615
R197 VDD1.n198 VDD1.n106 104.615
R198 VDD1.n199 VDD1.n198 104.615
R199 VDD1.n207 VDD1.n206 61.9117
R200 VDD1.n102 VDD1.n101 60.8422
R201 VDD1.n209 VDD1.n208 60.842
R202 VDD1.n205 VDD1.n204 60.842
R203 VDD1.t6 VDD1.n32 52.3082
R204 VDD1.t4 VDD1.n134 52.3082
R205 VDD1.n102 VDD1.n100 50.5581
R206 VDD1.n205 VDD1.n203 50.5581
R207 VDD1.n209 VDD1.n207 47.9061
R208 VDD1.n34 VDD1.n33 15.6677
R209 VDD1.n136 VDD1.n135 15.6677
R210 VDD1.n81 VDD1.n10 13.1884
R211 VDD1.n184 VDD1.n113 13.1884
R212 VDD1.n82 VDD1.n8 12.8005
R213 VDD1.n77 VDD1.n12 12.8005
R214 VDD1.n37 VDD1.n36 12.8005
R215 VDD1.n139 VDD1.n138 12.8005
R216 VDD1.n180 VDD1.n179 12.8005
R217 VDD1.n185 VDD1.n111 12.8005
R218 VDD1.n86 VDD1.n85 12.0247
R219 VDD1.n76 VDD1.n13 12.0247
R220 VDD1.n40 VDD1.n31 12.0247
R221 VDD1.n142 VDD1.n133 12.0247
R222 VDD1.n178 VDD1.n115 12.0247
R223 VDD1.n189 VDD1.n188 12.0247
R224 VDD1.n89 VDD1.n6 11.249
R225 VDD1.n73 VDD1.n72 11.249
R226 VDD1.n41 VDD1.n29 11.249
R227 VDD1.n143 VDD1.n131 11.249
R228 VDD1.n175 VDD1.n174 11.249
R229 VDD1.n192 VDD1.n109 11.249
R230 VDD1.n90 VDD1.n4 10.4732
R231 VDD1.n69 VDD1.n15 10.4732
R232 VDD1.n45 VDD1.n44 10.4732
R233 VDD1.n147 VDD1.n146 10.4732
R234 VDD1.n171 VDD1.n117 10.4732
R235 VDD1.n193 VDD1.n107 10.4732
R236 VDD1.n94 VDD1.n93 9.69747
R237 VDD1.n68 VDD1.n17 9.69747
R238 VDD1.n48 VDD1.n27 9.69747
R239 VDD1.n150 VDD1.n129 9.69747
R240 VDD1.n170 VDD1.n119 9.69747
R241 VDD1.n197 VDD1.n196 9.69747
R242 VDD1.n100 VDD1.n99 9.45567
R243 VDD1.n203 VDD1.n202 9.45567
R244 VDD1.n60 VDD1.n59 9.3005
R245 VDD1.n19 VDD1.n18 9.3005
R246 VDD1.n66 VDD1.n65 9.3005
R247 VDD1.n68 VDD1.n67 9.3005
R248 VDD1.n15 VDD1.n14 9.3005
R249 VDD1.n74 VDD1.n73 9.3005
R250 VDD1.n76 VDD1.n75 9.3005
R251 VDD1.n12 VDD1.n9 9.3005
R252 VDD1.n99 VDD1.n98 9.3005
R253 VDD1.n2 VDD1.n1 9.3005
R254 VDD1.n93 VDD1.n92 9.3005
R255 VDD1.n91 VDD1.n90 9.3005
R256 VDD1.n6 VDD1.n5 9.3005
R257 VDD1.n85 VDD1.n84 9.3005
R258 VDD1.n83 VDD1.n82 9.3005
R259 VDD1.n58 VDD1.n57 9.3005
R260 VDD1.n23 VDD1.n22 9.3005
R261 VDD1.n52 VDD1.n51 9.3005
R262 VDD1.n50 VDD1.n49 9.3005
R263 VDD1.n27 VDD1.n26 9.3005
R264 VDD1.n44 VDD1.n43 9.3005
R265 VDD1.n42 VDD1.n41 9.3005
R266 VDD1.n31 VDD1.n30 9.3005
R267 VDD1.n36 VDD1.n35 9.3005
R268 VDD1.n202 VDD1.n201 9.3005
R269 VDD1.n105 VDD1.n104 9.3005
R270 VDD1.n196 VDD1.n195 9.3005
R271 VDD1.n194 VDD1.n193 9.3005
R272 VDD1.n109 VDD1.n108 9.3005
R273 VDD1.n188 VDD1.n187 9.3005
R274 VDD1.n186 VDD1.n185 9.3005
R275 VDD1.n125 VDD1.n124 9.3005
R276 VDD1.n154 VDD1.n153 9.3005
R277 VDD1.n152 VDD1.n151 9.3005
R278 VDD1.n129 VDD1.n128 9.3005
R279 VDD1.n146 VDD1.n145 9.3005
R280 VDD1.n144 VDD1.n143 9.3005
R281 VDD1.n133 VDD1.n132 9.3005
R282 VDD1.n138 VDD1.n137 9.3005
R283 VDD1.n160 VDD1.n159 9.3005
R284 VDD1.n162 VDD1.n161 9.3005
R285 VDD1.n121 VDD1.n120 9.3005
R286 VDD1.n168 VDD1.n167 9.3005
R287 VDD1.n170 VDD1.n169 9.3005
R288 VDD1.n117 VDD1.n116 9.3005
R289 VDD1.n176 VDD1.n175 9.3005
R290 VDD1.n178 VDD1.n177 9.3005
R291 VDD1.n179 VDD1.n112 9.3005
R292 VDD1.n97 VDD1.n2 8.92171
R293 VDD1.n65 VDD1.n64 8.92171
R294 VDD1.n49 VDD1.n25 8.92171
R295 VDD1.n151 VDD1.n127 8.92171
R296 VDD1.n167 VDD1.n166 8.92171
R297 VDD1.n200 VDD1.n105 8.92171
R298 VDD1.n98 VDD1.n0 8.14595
R299 VDD1.n61 VDD1.n19 8.14595
R300 VDD1.n53 VDD1.n52 8.14595
R301 VDD1.n155 VDD1.n154 8.14595
R302 VDD1.n163 VDD1.n121 8.14595
R303 VDD1.n201 VDD1.n103 8.14595
R304 VDD1.n60 VDD1.n21 7.3702
R305 VDD1.n56 VDD1.n23 7.3702
R306 VDD1.n158 VDD1.n125 7.3702
R307 VDD1.n162 VDD1.n123 7.3702
R308 VDD1.n57 VDD1.n21 6.59444
R309 VDD1.n57 VDD1.n56 6.59444
R310 VDD1.n159 VDD1.n158 6.59444
R311 VDD1.n159 VDD1.n123 6.59444
R312 VDD1.n100 VDD1.n0 5.81868
R313 VDD1.n61 VDD1.n60 5.81868
R314 VDD1.n53 VDD1.n23 5.81868
R315 VDD1.n155 VDD1.n125 5.81868
R316 VDD1.n163 VDD1.n162 5.81868
R317 VDD1.n203 VDD1.n103 5.81868
R318 VDD1.n98 VDD1.n97 5.04292
R319 VDD1.n64 VDD1.n19 5.04292
R320 VDD1.n52 VDD1.n25 5.04292
R321 VDD1.n154 VDD1.n127 5.04292
R322 VDD1.n166 VDD1.n121 5.04292
R323 VDD1.n201 VDD1.n200 5.04292
R324 VDD1.n35 VDD1.n34 4.38563
R325 VDD1.n137 VDD1.n136 4.38563
R326 VDD1.n94 VDD1.n2 4.26717
R327 VDD1.n65 VDD1.n17 4.26717
R328 VDD1.n49 VDD1.n48 4.26717
R329 VDD1.n151 VDD1.n150 4.26717
R330 VDD1.n167 VDD1.n119 4.26717
R331 VDD1.n197 VDD1.n105 4.26717
R332 VDD1.n93 VDD1.n4 3.49141
R333 VDD1.n69 VDD1.n68 3.49141
R334 VDD1.n45 VDD1.n27 3.49141
R335 VDD1.n147 VDD1.n129 3.49141
R336 VDD1.n171 VDD1.n170 3.49141
R337 VDD1.n196 VDD1.n107 3.49141
R338 VDD1.n90 VDD1.n89 2.71565
R339 VDD1.n72 VDD1.n15 2.71565
R340 VDD1.n44 VDD1.n29 2.71565
R341 VDD1.n146 VDD1.n131 2.71565
R342 VDD1.n174 VDD1.n117 2.71565
R343 VDD1.n193 VDD1.n192 2.71565
R344 VDD1.n86 VDD1.n6 1.93989
R345 VDD1.n73 VDD1.n13 1.93989
R346 VDD1.n41 VDD1.n40 1.93989
R347 VDD1.n143 VDD1.n142 1.93989
R348 VDD1.n175 VDD1.n115 1.93989
R349 VDD1.n189 VDD1.n109 1.93989
R350 VDD1.n85 VDD1.n8 1.16414
R351 VDD1.n77 VDD1.n76 1.16414
R352 VDD1.n37 VDD1.n31 1.16414
R353 VDD1.n139 VDD1.n133 1.16414
R354 VDD1.n180 VDD1.n178 1.16414
R355 VDD1.n188 VDD1.n111 1.16414
R356 VDD1.n208 VDD1.t1 1.08543
R357 VDD1.n208 VDD1.t3 1.08543
R358 VDD1.n101 VDD1.t2 1.08543
R359 VDD1.n101 VDD1.t5 1.08543
R360 VDD1.n206 VDD1.t8 1.08543
R361 VDD1.n206 VDD1.t9 1.08543
R362 VDD1.n204 VDD1.t0 1.08543
R363 VDD1.n204 VDD1.t7 1.08543
R364 VDD1 VDD1.n209 1.06731
R365 VDD1 VDD1.n102 0.43369
R366 VDD1.n82 VDD1.n81 0.388379
R367 VDD1.n12 VDD1.n10 0.388379
R368 VDD1.n36 VDD1.n33 0.388379
R369 VDD1.n138 VDD1.n135 0.388379
R370 VDD1.n179 VDD1.n113 0.388379
R371 VDD1.n185 VDD1.n184 0.388379
R372 VDD1.n207 VDD1.n205 0.320154
R373 VDD1.n99 VDD1.n1 0.155672
R374 VDD1.n92 VDD1.n1 0.155672
R375 VDD1.n92 VDD1.n91 0.155672
R376 VDD1.n91 VDD1.n5 0.155672
R377 VDD1.n84 VDD1.n5 0.155672
R378 VDD1.n84 VDD1.n83 0.155672
R379 VDD1.n83 VDD1.n9 0.155672
R380 VDD1.n75 VDD1.n9 0.155672
R381 VDD1.n75 VDD1.n74 0.155672
R382 VDD1.n74 VDD1.n14 0.155672
R383 VDD1.n67 VDD1.n14 0.155672
R384 VDD1.n67 VDD1.n66 0.155672
R385 VDD1.n66 VDD1.n18 0.155672
R386 VDD1.n59 VDD1.n18 0.155672
R387 VDD1.n59 VDD1.n58 0.155672
R388 VDD1.n58 VDD1.n22 0.155672
R389 VDD1.n51 VDD1.n22 0.155672
R390 VDD1.n51 VDD1.n50 0.155672
R391 VDD1.n50 VDD1.n26 0.155672
R392 VDD1.n43 VDD1.n26 0.155672
R393 VDD1.n43 VDD1.n42 0.155672
R394 VDD1.n42 VDD1.n30 0.155672
R395 VDD1.n35 VDD1.n30 0.155672
R396 VDD1.n137 VDD1.n132 0.155672
R397 VDD1.n144 VDD1.n132 0.155672
R398 VDD1.n145 VDD1.n144 0.155672
R399 VDD1.n145 VDD1.n128 0.155672
R400 VDD1.n152 VDD1.n128 0.155672
R401 VDD1.n153 VDD1.n152 0.155672
R402 VDD1.n153 VDD1.n124 0.155672
R403 VDD1.n160 VDD1.n124 0.155672
R404 VDD1.n161 VDD1.n160 0.155672
R405 VDD1.n161 VDD1.n120 0.155672
R406 VDD1.n168 VDD1.n120 0.155672
R407 VDD1.n169 VDD1.n168 0.155672
R408 VDD1.n169 VDD1.n116 0.155672
R409 VDD1.n176 VDD1.n116 0.155672
R410 VDD1.n177 VDD1.n176 0.155672
R411 VDD1.n177 VDD1.n112 0.155672
R412 VDD1.n186 VDD1.n112 0.155672
R413 VDD1.n187 VDD1.n186 0.155672
R414 VDD1.n187 VDD1.n108 0.155672
R415 VDD1.n194 VDD1.n108 0.155672
R416 VDD1.n195 VDD1.n194 0.155672
R417 VDD1.n195 VDD1.n104 0.155672
R418 VDD1.n202 VDD1.n104 0.155672
R419 VTAIL.n416 VTAIL.n320 289.615
R420 VTAIL.n98 VTAIL.n2 289.615
R421 VTAIL.n314 VTAIL.n218 289.615
R422 VTAIL.n208 VTAIL.n112 289.615
R423 VTAIL.n352 VTAIL.n351 185
R424 VTAIL.n357 VTAIL.n356 185
R425 VTAIL.n359 VTAIL.n358 185
R426 VTAIL.n348 VTAIL.n347 185
R427 VTAIL.n365 VTAIL.n364 185
R428 VTAIL.n367 VTAIL.n366 185
R429 VTAIL.n344 VTAIL.n343 185
R430 VTAIL.n373 VTAIL.n372 185
R431 VTAIL.n375 VTAIL.n374 185
R432 VTAIL.n340 VTAIL.n339 185
R433 VTAIL.n381 VTAIL.n380 185
R434 VTAIL.n383 VTAIL.n382 185
R435 VTAIL.n336 VTAIL.n335 185
R436 VTAIL.n389 VTAIL.n388 185
R437 VTAIL.n391 VTAIL.n390 185
R438 VTAIL.n332 VTAIL.n331 185
R439 VTAIL.n398 VTAIL.n397 185
R440 VTAIL.n399 VTAIL.n330 185
R441 VTAIL.n401 VTAIL.n400 185
R442 VTAIL.n328 VTAIL.n327 185
R443 VTAIL.n407 VTAIL.n406 185
R444 VTAIL.n409 VTAIL.n408 185
R445 VTAIL.n324 VTAIL.n323 185
R446 VTAIL.n415 VTAIL.n414 185
R447 VTAIL.n417 VTAIL.n416 185
R448 VTAIL.n34 VTAIL.n33 185
R449 VTAIL.n39 VTAIL.n38 185
R450 VTAIL.n41 VTAIL.n40 185
R451 VTAIL.n30 VTAIL.n29 185
R452 VTAIL.n47 VTAIL.n46 185
R453 VTAIL.n49 VTAIL.n48 185
R454 VTAIL.n26 VTAIL.n25 185
R455 VTAIL.n55 VTAIL.n54 185
R456 VTAIL.n57 VTAIL.n56 185
R457 VTAIL.n22 VTAIL.n21 185
R458 VTAIL.n63 VTAIL.n62 185
R459 VTAIL.n65 VTAIL.n64 185
R460 VTAIL.n18 VTAIL.n17 185
R461 VTAIL.n71 VTAIL.n70 185
R462 VTAIL.n73 VTAIL.n72 185
R463 VTAIL.n14 VTAIL.n13 185
R464 VTAIL.n80 VTAIL.n79 185
R465 VTAIL.n81 VTAIL.n12 185
R466 VTAIL.n83 VTAIL.n82 185
R467 VTAIL.n10 VTAIL.n9 185
R468 VTAIL.n89 VTAIL.n88 185
R469 VTAIL.n91 VTAIL.n90 185
R470 VTAIL.n6 VTAIL.n5 185
R471 VTAIL.n97 VTAIL.n96 185
R472 VTAIL.n99 VTAIL.n98 185
R473 VTAIL.n315 VTAIL.n314 185
R474 VTAIL.n313 VTAIL.n312 185
R475 VTAIL.n222 VTAIL.n221 185
R476 VTAIL.n307 VTAIL.n306 185
R477 VTAIL.n305 VTAIL.n304 185
R478 VTAIL.n226 VTAIL.n225 185
R479 VTAIL.n299 VTAIL.n298 185
R480 VTAIL.n297 VTAIL.n228 185
R481 VTAIL.n296 VTAIL.n295 185
R482 VTAIL.n231 VTAIL.n229 185
R483 VTAIL.n290 VTAIL.n289 185
R484 VTAIL.n288 VTAIL.n287 185
R485 VTAIL.n235 VTAIL.n234 185
R486 VTAIL.n282 VTAIL.n281 185
R487 VTAIL.n280 VTAIL.n279 185
R488 VTAIL.n239 VTAIL.n238 185
R489 VTAIL.n274 VTAIL.n273 185
R490 VTAIL.n272 VTAIL.n271 185
R491 VTAIL.n243 VTAIL.n242 185
R492 VTAIL.n266 VTAIL.n265 185
R493 VTAIL.n264 VTAIL.n263 185
R494 VTAIL.n247 VTAIL.n246 185
R495 VTAIL.n258 VTAIL.n257 185
R496 VTAIL.n256 VTAIL.n255 185
R497 VTAIL.n251 VTAIL.n250 185
R498 VTAIL.n209 VTAIL.n208 185
R499 VTAIL.n207 VTAIL.n206 185
R500 VTAIL.n116 VTAIL.n115 185
R501 VTAIL.n201 VTAIL.n200 185
R502 VTAIL.n199 VTAIL.n198 185
R503 VTAIL.n120 VTAIL.n119 185
R504 VTAIL.n193 VTAIL.n192 185
R505 VTAIL.n191 VTAIL.n122 185
R506 VTAIL.n190 VTAIL.n189 185
R507 VTAIL.n125 VTAIL.n123 185
R508 VTAIL.n184 VTAIL.n183 185
R509 VTAIL.n182 VTAIL.n181 185
R510 VTAIL.n129 VTAIL.n128 185
R511 VTAIL.n176 VTAIL.n175 185
R512 VTAIL.n174 VTAIL.n173 185
R513 VTAIL.n133 VTAIL.n132 185
R514 VTAIL.n168 VTAIL.n167 185
R515 VTAIL.n166 VTAIL.n165 185
R516 VTAIL.n137 VTAIL.n136 185
R517 VTAIL.n160 VTAIL.n159 185
R518 VTAIL.n158 VTAIL.n157 185
R519 VTAIL.n141 VTAIL.n140 185
R520 VTAIL.n152 VTAIL.n151 185
R521 VTAIL.n150 VTAIL.n149 185
R522 VTAIL.n145 VTAIL.n144 185
R523 VTAIL.n353 VTAIL.t9 147.659
R524 VTAIL.n35 VTAIL.t15 147.659
R525 VTAIL.n252 VTAIL.t11 147.659
R526 VTAIL.n146 VTAIL.t5 147.659
R527 VTAIL.n357 VTAIL.n351 104.615
R528 VTAIL.n358 VTAIL.n357 104.615
R529 VTAIL.n358 VTAIL.n347 104.615
R530 VTAIL.n365 VTAIL.n347 104.615
R531 VTAIL.n366 VTAIL.n365 104.615
R532 VTAIL.n366 VTAIL.n343 104.615
R533 VTAIL.n373 VTAIL.n343 104.615
R534 VTAIL.n374 VTAIL.n373 104.615
R535 VTAIL.n374 VTAIL.n339 104.615
R536 VTAIL.n381 VTAIL.n339 104.615
R537 VTAIL.n382 VTAIL.n381 104.615
R538 VTAIL.n382 VTAIL.n335 104.615
R539 VTAIL.n389 VTAIL.n335 104.615
R540 VTAIL.n390 VTAIL.n389 104.615
R541 VTAIL.n390 VTAIL.n331 104.615
R542 VTAIL.n398 VTAIL.n331 104.615
R543 VTAIL.n399 VTAIL.n398 104.615
R544 VTAIL.n400 VTAIL.n399 104.615
R545 VTAIL.n400 VTAIL.n327 104.615
R546 VTAIL.n407 VTAIL.n327 104.615
R547 VTAIL.n408 VTAIL.n407 104.615
R548 VTAIL.n408 VTAIL.n323 104.615
R549 VTAIL.n415 VTAIL.n323 104.615
R550 VTAIL.n416 VTAIL.n415 104.615
R551 VTAIL.n39 VTAIL.n33 104.615
R552 VTAIL.n40 VTAIL.n39 104.615
R553 VTAIL.n40 VTAIL.n29 104.615
R554 VTAIL.n47 VTAIL.n29 104.615
R555 VTAIL.n48 VTAIL.n47 104.615
R556 VTAIL.n48 VTAIL.n25 104.615
R557 VTAIL.n55 VTAIL.n25 104.615
R558 VTAIL.n56 VTAIL.n55 104.615
R559 VTAIL.n56 VTAIL.n21 104.615
R560 VTAIL.n63 VTAIL.n21 104.615
R561 VTAIL.n64 VTAIL.n63 104.615
R562 VTAIL.n64 VTAIL.n17 104.615
R563 VTAIL.n71 VTAIL.n17 104.615
R564 VTAIL.n72 VTAIL.n71 104.615
R565 VTAIL.n72 VTAIL.n13 104.615
R566 VTAIL.n80 VTAIL.n13 104.615
R567 VTAIL.n81 VTAIL.n80 104.615
R568 VTAIL.n82 VTAIL.n81 104.615
R569 VTAIL.n82 VTAIL.n9 104.615
R570 VTAIL.n89 VTAIL.n9 104.615
R571 VTAIL.n90 VTAIL.n89 104.615
R572 VTAIL.n90 VTAIL.n5 104.615
R573 VTAIL.n97 VTAIL.n5 104.615
R574 VTAIL.n98 VTAIL.n97 104.615
R575 VTAIL.n314 VTAIL.n313 104.615
R576 VTAIL.n313 VTAIL.n221 104.615
R577 VTAIL.n306 VTAIL.n221 104.615
R578 VTAIL.n306 VTAIL.n305 104.615
R579 VTAIL.n305 VTAIL.n225 104.615
R580 VTAIL.n298 VTAIL.n225 104.615
R581 VTAIL.n298 VTAIL.n297 104.615
R582 VTAIL.n297 VTAIL.n296 104.615
R583 VTAIL.n296 VTAIL.n229 104.615
R584 VTAIL.n289 VTAIL.n229 104.615
R585 VTAIL.n289 VTAIL.n288 104.615
R586 VTAIL.n288 VTAIL.n234 104.615
R587 VTAIL.n281 VTAIL.n234 104.615
R588 VTAIL.n281 VTAIL.n280 104.615
R589 VTAIL.n280 VTAIL.n238 104.615
R590 VTAIL.n273 VTAIL.n238 104.615
R591 VTAIL.n273 VTAIL.n272 104.615
R592 VTAIL.n272 VTAIL.n242 104.615
R593 VTAIL.n265 VTAIL.n242 104.615
R594 VTAIL.n265 VTAIL.n264 104.615
R595 VTAIL.n264 VTAIL.n246 104.615
R596 VTAIL.n257 VTAIL.n246 104.615
R597 VTAIL.n257 VTAIL.n256 104.615
R598 VTAIL.n256 VTAIL.n250 104.615
R599 VTAIL.n208 VTAIL.n207 104.615
R600 VTAIL.n207 VTAIL.n115 104.615
R601 VTAIL.n200 VTAIL.n115 104.615
R602 VTAIL.n200 VTAIL.n199 104.615
R603 VTAIL.n199 VTAIL.n119 104.615
R604 VTAIL.n192 VTAIL.n119 104.615
R605 VTAIL.n192 VTAIL.n191 104.615
R606 VTAIL.n191 VTAIL.n190 104.615
R607 VTAIL.n190 VTAIL.n123 104.615
R608 VTAIL.n183 VTAIL.n123 104.615
R609 VTAIL.n183 VTAIL.n182 104.615
R610 VTAIL.n182 VTAIL.n128 104.615
R611 VTAIL.n175 VTAIL.n128 104.615
R612 VTAIL.n175 VTAIL.n174 104.615
R613 VTAIL.n174 VTAIL.n132 104.615
R614 VTAIL.n167 VTAIL.n132 104.615
R615 VTAIL.n167 VTAIL.n166 104.615
R616 VTAIL.n166 VTAIL.n136 104.615
R617 VTAIL.n159 VTAIL.n136 104.615
R618 VTAIL.n159 VTAIL.n158 104.615
R619 VTAIL.n158 VTAIL.n140 104.615
R620 VTAIL.n151 VTAIL.n140 104.615
R621 VTAIL.n151 VTAIL.n150 104.615
R622 VTAIL.n150 VTAIL.n144 104.615
R623 VTAIL.t9 VTAIL.n351 52.3082
R624 VTAIL.t15 VTAIL.n33 52.3082
R625 VTAIL.t11 VTAIL.n250 52.3082
R626 VTAIL.t5 VTAIL.n144 52.3082
R627 VTAIL.n217 VTAIL.n216 44.1634
R628 VTAIL.n215 VTAIL.n214 44.1634
R629 VTAIL.n111 VTAIL.n110 44.1634
R630 VTAIL.n109 VTAIL.n108 44.1634
R631 VTAIL.n423 VTAIL.n422 44.1633
R632 VTAIL.n1 VTAIL.n0 44.1633
R633 VTAIL.n105 VTAIL.n104 44.1633
R634 VTAIL.n107 VTAIL.n106 44.1633
R635 VTAIL.n421 VTAIL.n420 32.3793
R636 VTAIL.n103 VTAIL.n102 32.3793
R637 VTAIL.n319 VTAIL.n318 32.3793
R638 VTAIL.n213 VTAIL.n212 32.3793
R639 VTAIL.n109 VTAIL.n107 31.0996
R640 VTAIL.n421 VTAIL.n319 29.5996
R641 VTAIL.n353 VTAIL.n352 15.6677
R642 VTAIL.n35 VTAIL.n34 15.6677
R643 VTAIL.n252 VTAIL.n251 15.6677
R644 VTAIL.n146 VTAIL.n145 15.6677
R645 VTAIL.n401 VTAIL.n330 13.1884
R646 VTAIL.n83 VTAIL.n12 13.1884
R647 VTAIL.n299 VTAIL.n228 13.1884
R648 VTAIL.n193 VTAIL.n122 13.1884
R649 VTAIL.n356 VTAIL.n355 12.8005
R650 VTAIL.n397 VTAIL.n396 12.8005
R651 VTAIL.n402 VTAIL.n328 12.8005
R652 VTAIL.n38 VTAIL.n37 12.8005
R653 VTAIL.n79 VTAIL.n78 12.8005
R654 VTAIL.n84 VTAIL.n10 12.8005
R655 VTAIL.n300 VTAIL.n226 12.8005
R656 VTAIL.n295 VTAIL.n230 12.8005
R657 VTAIL.n255 VTAIL.n254 12.8005
R658 VTAIL.n194 VTAIL.n120 12.8005
R659 VTAIL.n189 VTAIL.n124 12.8005
R660 VTAIL.n149 VTAIL.n148 12.8005
R661 VTAIL.n359 VTAIL.n350 12.0247
R662 VTAIL.n395 VTAIL.n332 12.0247
R663 VTAIL.n406 VTAIL.n405 12.0247
R664 VTAIL.n41 VTAIL.n32 12.0247
R665 VTAIL.n77 VTAIL.n14 12.0247
R666 VTAIL.n88 VTAIL.n87 12.0247
R667 VTAIL.n304 VTAIL.n303 12.0247
R668 VTAIL.n294 VTAIL.n231 12.0247
R669 VTAIL.n258 VTAIL.n249 12.0247
R670 VTAIL.n198 VTAIL.n197 12.0247
R671 VTAIL.n188 VTAIL.n125 12.0247
R672 VTAIL.n152 VTAIL.n143 12.0247
R673 VTAIL.n360 VTAIL.n348 11.249
R674 VTAIL.n392 VTAIL.n391 11.249
R675 VTAIL.n409 VTAIL.n326 11.249
R676 VTAIL.n42 VTAIL.n30 11.249
R677 VTAIL.n74 VTAIL.n73 11.249
R678 VTAIL.n91 VTAIL.n8 11.249
R679 VTAIL.n307 VTAIL.n224 11.249
R680 VTAIL.n291 VTAIL.n290 11.249
R681 VTAIL.n259 VTAIL.n247 11.249
R682 VTAIL.n201 VTAIL.n118 11.249
R683 VTAIL.n185 VTAIL.n184 11.249
R684 VTAIL.n153 VTAIL.n141 11.249
R685 VTAIL.n364 VTAIL.n363 10.4732
R686 VTAIL.n388 VTAIL.n334 10.4732
R687 VTAIL.n410 VTAIL.n324 10.4732
R688 VTAIL.n46 VTAIL.n45 10.4732
R689 VTAIL.n70 VTAIL.n16 10.4732
R690 VTAIL.n92 VTAIL.n6 10.4732
R691 VTAIL.n308 VTAIL.n222 10.4732
R692 VTAIL.n287 VTAIL.n233 10.4732
R693 VTAIL.n263 VTAIL.n262 10.4732
R694 VTAIL.n202 VTAIL.n116 10.4732
R695 VTAIL.n181 VTAIL.n127 10.4732
R696 VTAIL.n157 VTAIL.n156 10.4732
R697 VTAIL.n367 VTAIL.n346 9.69747
R698 VTAIL.n387 VTAIL.n336 9.69747
R699 VTAIL.n414 VTAIL.n413 9.69747
R700 VTAIL.n49 VTAIL.n28 9.69747
R701 VTAIL.n69 VTAIL.n18 9.69747
R702 VTAIL.n96 VTAIL.n95 9.69747
R703 VTAIL.n312 VTAIL.n311 9.69747
R704 VTAIL.n286 VTAIL.n235 9.69747
R705 VTAIL.n266 VTAIL.n245 9.69747
R706 VTAIL.n206 VTAIL.n205 9.69747
R707 VTAIL.n180 VTAIL.n129 9.69747
R708 VTAIL.n160 VTAIL.n139 9.69747
R709 VTAIL.n420 VTAIL.n419 9.45567
R710 VTAIL.n102 VTAIL.n101 9.45567
R711 VTAIL.n318 VTAIL.n317 9.45567
R712 VTAIL.n212 VTAIL.n211 9.45567
R713 VTAIL.n419 VTAIL.n418 9.3005
R714 VTAIL.n322 VTAIL.n321 9.3005
R715 VTAIL.n413 VTAIL.n412 9.3005
R716 VTAIL.n411 VTAIL.n410 9.3005
R717 VTAIL.n326 VTAIL.n325 9.3005
R718 VTAIL.n405 VTAIL.n404 9.3005
R719 VTAIL.n403 VTAIL.n402 9.3005
R720 VTAIL.n342 VTAIL.n341 9.3005
R721 VTAIL.n371 VTAIL.n370 9.3005
R722 VTAIL.n369 VTAIL.n368 9.3005
R723 VTAIL.n346 VTAIL.n345 9.3005
R724 VTAIL.n363 VTAIL.n362 9.3005
R725 VTAIL.n361 VTAIL.n360 9.3005
R726 VTAIL.n350 VTAIL.n349 9.3005
R727 VTAIL.n355 VTAIL.n354 9.3005
R728 VTAIL.n377 VTAIL.n376 9.3005
R729 VTAIL.n379 VTAIL.n378 9.3005
R730 VTAIL.n338 VTAIL.n337 9.3005
R731 VTAIL.n385 VTAIL.n384 9.3005
R732 VTAIL.n387 VTAIL.n386 9.3005
R733 VTAIL.n334 VTAIL.n333 9.3005
R734 VTAIL.n393 VTAIL.n392 9.3005
R735 VTAIL.n395 VTAIL.n394 9.3005
R736 VTAIL.n396 VTAIL.n329 9.3005
R737 VTAIL.n101 VTAIL.n100 9.3005
R738 VTAIL.n4 VTAIL.n3 9.3005
R739 VTAIL.n95 VTAIL.n94 9.3005
R740 VTAIL.n93 VTAIL.n92 9.3005
R741 VTAIL.n8 VTAIL.n7 9.3005
R742 VTAIL.n87 VTAIL.n86 9.3005
R743 VTAIL.n85 VTAIL.n84 9.3005
R744 VTAIL.n24 VTAIL.n23 9.3005
R745 VTAIL.n53 VTAIL.n52 9.3005
R746 VTAIL.n51 VTAIL.n50 9.3005
R747 VTAIL.n28 VTAIL.n27 9.3005
R748 VTAIL.n45 VTAIL.n44 9.3005
R749 VTAIL.n43 VTAIL.n42 9.3005
R750 VTAIL.n32 VTAIL.n31 9.3005
R751 VTAIL.n37 VTAIL.n36 9.3005
R752 VTAIL.n59 VTAIL.n58 9.3005
R753 VTAIL.n61 VTAIL.n60 9.3005
R754 VTAIL.n20 VTAIL.n19 9.3005
R755 VTAIL.n67 VTAIL.n66 9.3005
R756 VTAIL.n69 VTAIL.n68 9.3005
R757 VTAIL.n16 VTAIL.n15 9.3005
R758 VTAIL.n75 VTAIL.n74 9.3005
R759 VTAIL.n77 VTAIL.n76 9.3005
R760 VTAIL.n78 VTAIL.n11 9.3005
R761 VTAIL.n278 VTAIL.n277 9.3005
R762 VTAIL.n237 VTAIL.n236 9.3005
R763 VTAIL.n284 VTAIL.n283 9.3005
R764 VTAIL.n286 VTAIL.n285 9.3005
R765 VTAIL.n233 VTAIL.n232 9.3005
R766 VTAIL.n292 VTAIL.n291 9.3005
R767 VTAIL.n294 VTAIL.n293 9.3005
R768 VTAIL.n230 VTAIL.n227 9.3005
R769 VTAIL.n317 VTAIL.n316 9.3005
R770 VTAIL.n220 VTAIL.n219 9.3005
R771 VTAIL.n311 VTAIL.n310 9.3005
R772 VTAIL.n309 VTAIL.n308 9.3005
R773 VTAIL.n224 VTAIL.n223 9.3005
R774 VTAIL.n303 VTAIL.n302 9.3005
R775 VTAIL.n301 VTAIL.n300 9.3005
R776 VTAIL.n276 VTAIL.n275 9.3005
R777 VTAIL.n241 VTAIL.n240 9.3005
R778 VTAIL.n270 VTAIL.n269 9.3005
R779 VTAIL.n268 VTAIL.n267 9.3005
R780 VTAIL.n245 VTAIL.n244 9.3005
R781 VTAIL.n262 VTAIL.n261 9.3005
R782 VTAIL.n260 VTAIL.n259 9.3005
R783 VTAIL.n249 VTAIL.n248 9.3005
R784 VTAIL.n254 VTAIL.n253 9.3005
R785 VTAIL.n172 VTAIL.n171 9.3005
R786 VTAIL.n131 VTAIL.n130 9.3005
R787 VTAIL.n178 VTAIL.n177 9.3005
R788 VTAIL.n180 VTAIL.n179 9.3005
R789 VTAIL.n127 VTAIL.n126 9.3005
R790 VTAIL.n186 VTAIL.n185 9.3005
R791 VTAIL.n188 VTAIL.n187 9.3005
R792 VTAIL.n124 VTAIL.n121 9.3005
R793 VTAIL.n211 VTAIL.n210 9.3005
R794 VTAIL.n114 VTAIL.n113 9.3005
R795 VTAIL.n205 VTAIL.n204 9.3005
R796 VTAIL.n203 VTAIL.n202 9.3005
R797 VTAIL.n118 VTAIL.n117 9.3005
R798 VTAIL.n197 VTAIL.n196 9.3005
R799 VTAIL.n195 VTAIL.n194 9.3005
R800 VTAIL.n170 VTAIL.n169 9.3005
R801 VTAIL.n135 VTAIL.n134 9.3005
R802 VTAIL.n164 VTAIL.n163 9.3005
R803 VTAIL.n162 VTAIL.n161 9.3005
R804 VTAIL.n139 VTAIL.n138 9.3005
R805 VTAIL.n156 VTAIL.n155 9.3005
R806 VTAIL.n154 VTAIL.n153 9.3005
R807 VTAIL.n143 VTAIL.n142 9.3005
R808 VTAIL.n148 VTAIL.n147 9.3005
R809 VTAIL.n368 VTAIL.n344 8.92171
R810 VTAIL.n384 VTAIL.n383 8.92171
R811 VTAIL.n417 VTAIL.n322 8.92171
R812 VTAIL.n50 VTAIL.n26 8.92171
R813 VTAIL.n66 VTAIL.n65 8.92171
R814 VTAIL.n99 VTAIL.n4 8.92171
R815 VTAIL.n315 VTAIL.n220 8.92171
R816 VTAIL.n283 VTAIL.n282 8.92171
R817 VTAIL.n267 VTAIL.n243 8.92171
R818 VTAIL.n209 VTAIL.n114 8.92171
R819 VTAIL.n177 VTAIL.n176 8.92171
R820 VTAIL.n161 VTAIL.n137 8.92171
R821 VTAIL.n372 VTAIL.n371 8.14595
R822 VTAIL.n380 VTAIL.n338 8.14595
R823 VTAIL.n418 VTAIL.n320 8.14595
R824 VTAIL.n54 VTAIL.n53 8.14595
R825 VTAIL.n62 VTAIL.n20 8.14595
R826 VTAIL.n100 VTAIL.n2 8.14595
R827 VTAIL.n316 VTAIL.n218 8.14595
R828 VTAIL.n279 VTAIL.n237 8.14595
R829 VTAIL.n271 VTAIL.n270 8.14595
R830 VTAIL.n210 VTAIL.n112 8.14595
R831 VTAIL.n173 VTAIL.n131 8.14595
R832 VTAIL.n165 VTAIL.n164 8.14595
R833 VTAIL.n375 VTAIL.n342 7.3702
R834 VTAIL.n379 VTAIL.n340 7.3702
R835 VTAIL.n57 VTAIL.n24 7.3702
R836 VTAIL.n61 VTAIL.n22 7.3702
R837 VTAIL.n278 VTAIL.n239 7.3702
R838 VTAIL.n274 VTAIL.n241 7.3702
R839 VTAIL.n172 VTAIL.n133 7.3702
R840 VTAIL.n168 VTAIL.n135 7.3702
R841 VTAIL.n376 VTAIL.n375 6.59444
R842 VTAIL.n376 VTAIL.n340 6.59444
R843 VTAIL.n58 VTAIL.n57 6.59444
R844 VTAIL.n58 VTAIL.n22 6.59444
R845 VTAIL.n275 VTAIL.n239 6.59444
R846 VTAIL.n275 VTAIL.n274 6.59444
R847 VTAIL.n169 VTAIL.n133 6.59444
R848 VTAIL.n169 VTAIL.n168 6.59444
R849 VTAIL.n372 VTAIL.n342 5.81868
R850 VTAIL.n380 VTAIL.n379 5.81868
R851 VTAIL.n420 VTAIL.n320 5.81868
R852 VTAIL.n54 VTAIL.n24 5.81868
R853 VTAIL.n62 VTAIL.n61 5.81868
R854 VTAIL.n102 VTAIL.n2 5.81868
R855 VTAIL.n318 VTAIL.n218 5.81868
R856 VTAIL.n279 VTAIL.n278 5.81868
R857 VTAIL.n271 VTAIL.n241 5.81868
R858 VTAIL.n212 VTAIL.n112 5.81868
R859 VTAIL.n173 VTAIL.n172 5.81868
R860 VTAIL.n165 VTAIL.n135 5.81868
R861 VTAIL.n371 VTAIL.n344 5.04292
R862 VTAIL.n383 VTAIL.n338 5.04292
R863 VTAIL.n418 VTAIL.n417 5.04292
R864 VTAIL.n53 VTAIL.n26 5.04292
R865 VTAIL.n65 VTAIL.n20 5.04292
R866 VTAIL.n100 VTAIL.n99 5.04292
R867 VTAIL.n316 VTAIL.n315 5.04292
R868 VTAIL.n282 VTAIL.n237 5.04292
R869 VTAIL.n270 VTAIL.n243 5.04292
R870 VTAIL.n210 VTAIL.n209 5.04292
R871 VTAIL.n176 VTAIL.n131 5.04292
R872 VTAIL.n164 VTAIL.n137 5.04292
R873 VTAIL.n354 VTAIL.n353 4.38563
R874 VTAIL.n36 VTAIL.n35 4.38563
R875 VTAIL.n253 VTAIL.n252 4.38563
R876 VTAIL.n147 VTAIL.n146 4.38563
R877 VTAIL.n368 VTAIL.n367 4.26717
R878 VTAIL.n384 VTAIL.n336 4.26717
R879 VTAIL.n414 VTAIL.n322 4.26717
R880 VTAIL.n50 VTAIL.n49 4.26717
R881 VTAIL.n66 VTAIL.n18 4.26717
R882 VTAIL.n96 VTAIL.n4 4.26717
R883 VTAIL.n312 VTAIL.n220 4.26717
R884 VTAIL.n283 VTAIL.n235 4.26717
R885 VTAIL.n267 VTAIL.n266 4.26717
R886 VTAIL.n206 VTAIL.n114 4.26717
R887 VTAIL.n177 VTAIL.n129 4.26717
R888 VTAIL.n161 VTAIL.n160 4.26717
R889 VTAIL.n364 VTAIL.n346 3.49141
R890 VTAIL.n388 VTAIL.n387 3.49141
R891 VTAIL.n413 VTAIL.n324 3.49141
R892 VTAIL.n46 VTAIL.n28 3.49141
R893 VTAIL.n70 VTAIL.n69 3.49141
R894 VTAIL.n95 VTAIL.n6 3.49141
R895 VTAIL.n311 VTAIL.n222 3.49141
R896 VTAIL.n287 VTAIL.n286 3.49141
R897 VTAIL.n263 VTAIL.n245 3.49141
R898 VTAIL.n205 VTAIL.n116 3.49141
R899 VTAIL.n181 VTAIL.n180 3.49141
R900 VTAIL.n157 VTAIL.n139 3.49141
R901 VTAIL.n363 VTAIL.n348 2.71565
R902 VTAIL.n391 VTAIL.n334 2.71565
R903 VTAIL.n410 VTAIL.n409 2.71565
R904 VTAIL.n45 VTAIL.n30 2.71565
R905 VTAIL.n73 VTAIL.n16 2.71565
R906 VTAIL.n92 VTAIL.n91 2.71565
R907 VTAIL.n308 VTAIL.n307 2.71565
R908 VTAIL.n290 VTAIL.n233 2.71565
R909 VTAIL.n262 VTAIL.n247 2.71565
R910 VTAIL.n202 VTAIL.n201 2.71565
R911 VTAIL.n184 VTAIL.n127 2.71565
R912 VTAIL.n156 VTAIL.n141 2.71565
R913 VTAIL.n360 VTAIL.n359 1.93989
R914 VTAIL.n392 VTAIL.n332 1.93989
R915 VTAIL.n406 VTAIL.n326 1.93989
R916 VTAIL.n42 VTAIL.n41 1.93989
R917 VTAIL.n74 VTAIL.n14 1.93989
R918 VTAIL.n88 VTAIL.n8 1.93989
R919 VTAIL.n304 VTAIL.n224 1.93989
R920 VTAIL.n291 VTAIL.n231 1.93989
R921 VTAIL.n259 VTAIL.n258 1.93989
R922 VTAIL.n198 VTAIL.n118 1.93989
R923 VTAIL.n185 VTAIL.n125 1.93989
R924 VTAIL.n153 VTAIL.n152 1.93989
R925 VTAIL.n111 VTAIL.n109 1.5005
R926 VTAIL.n213 VTAIL.n111 1.5005
R927 VTAIL.n217 VTAIL.n215 1.5005
R928 VTAIL.n319 VTAIL.n217 1.5005
R929 VTAIL.n107 VTAIL.n105 1.5005
R930 VTAIL.n105 VTAIL.n103 1.5005
R931 VTAIL.n423 VTAIL.n421 1.5005
R932 VTAIL.n215 VTAIL.n213 1.22033
R933 VTAIL.n103 VTAIL.n1 1.22033
R934 VTAIL VTAIL.n1 1.18369
R935 VTAIL.n356 VTAIL.n350 1.16414
R936 VTAIL.n397 VTAIL.n395 1.16414
R937 VTAIL.n405 VTAIL.n328 1.16414
R938 VTAIL.n38 VTAIL.n32 1.16414
R939 VTAIL.n79 VTAIL.n77 1.16414
R940 VTAIL.n87 VTAIL.n10 1.16414
R941 VTAIL.n303 VTAIL.n226 1.16414
R942 VTAIL.n295 VTAIL.n294 1.16414
R943 VTAIL.n255 VTAIL.n249 1.16414
R944 VTAIL.n197 VTAIL.n120 1.16414
R945 VTAIL.n189 VTAIL.n188 1.16414
R946 VTAIL.n149 VTAIL.n143 1.16414
R947 VTAIL.n422 VTAIL.t6 1.08543
R948 VTAIL.n422 VTAIL.t7 1.08543
R949 VTAIL.n0 VTAIL.t2 1.08543
R950 VTAIL.n0 VTAIL.t1 1.08543
R951 VTAIL.n104 VTAIL.t17 1.08543
R952 VTAIL.n104 VTAIL.t14 1.08543
R953 VTAIL.n106 VTAIL.t12 1.08543
R954 VTAIL.n106 VTAIL.t18 1.08543
R955 VTAIL.n216 VTAIL.t13 1.08543
R956 VTAIL.n216 VTAIL.t19 1.08543
R957 VTAIL.n214 VTAIL.t16 1.08543
R958 VTAIL.n214 VTAIL.t10 1.08543
R959 VTAIL.n110 VTAIL.t4 1.08543
R960 VTAIL.n110 VTAIL.t8 1.08543
R961 VTAIL.n108 VTAIL.t0 1.08543
R962 VTAIL.n108 VTAIL.t3 1.08543
R963 VTAIL.n355 VTAIL.n352 0.388379
R964 VTAIL.n396 VTAIL.n330 0.388379
R965 VTAIL.n402 VTAIL.n401 0.388379
R966 VTAIL.n37 VTAIL.n34 0.388379
R967 VTAIL.n78 VTAIL.n12 0.388379
R968 VTAIL.n84 VTAIL.n83 0.388379
R969 VTAIL.n300 VTAIL.n299 0.388379
R970 VTAIL.n230 VTAIL.n228 0.388379
R971 VTAIL.n254 VTAIL.n251 0.388379
R972 VTAIL.n194 VTAIL.n193 0.388379
R973 VTAIL.n124 VTAIL.n122 0.388379
R974 VTAIL.n148 VTAIL.n145 0.388379
R975 VTAIL VTAIL.n423 0.31731
R976 VTAIL.n354 VTAIL.n349 0.155672
R977 VTAIL.n361 VTAIL.n349 0.155672
R978 VTAIL.n362 VTAIL.n361 0.155672
R979 VTAIL.n362 VTAIL.n345 0.155672
R980 VTAIL.n369 VTAIL.n345 0.155672
R981 VTAIL.n370 VTAIL.n369 0.155672
R982 VTAIL.n370 VTAIL.n341 0.155672
R983 VTAIL.n377 VTAIL.n341 0.155672
R984 VTAIL.n378 VTAIL.n377 0.155672
R985 VTAIL.n378 VTAIL.n337 0.155672
R986 VTAIL.n385 VTAIL.n337 0.155672
R987 VTAIL.n386 VTAIL.n385 0.155672
R988 VTAIL.n386 VTAIL.n333 0.155672
R989 VTAIL.n393 VTAIL.n333 0.155672
R990 VTAIL.n394 VTAIL.n393 0.155672
R991 VTAIL.n394 VTAIL.n329 0.155672
R992 VTAIL.n403 VTAIL.n329 0.155672
R993 VTAIL.n404 VTAIL.n403 0.155672
R994 VTAIL.n404 VTAIL.n325 0.155672
R995 VTAIL.n411 VTAIL.n325 0.155672
R996 VTAIL.n412 VTAIL.n411 0.155672
R997 VTAIL.n412 VTAIL.n321 0.155672
R998 VTAIL.n419 VTAIL.n321 0.155672
R999 VTAIL.n36 VTAIL.n31 0.155672
R1000 VTAIL.n43 VTAIL.n31 0.155672
R1001 VTAIL.n44 VTAIL.n43 0.155672
R1002 VTAIL.n44 VTAIL.n27 0.155672
R1003 VTAIL.n51 VTAIL.n27 0.155672
R1004 VTAIL.n52 VTAIL.n51 0.155672
R1005 VTAIL.n52 VTAIL.n23 0.155672
R1006 VTAIL.n59 VTAIL.n23 0.155672
R1007 VTAIL.n60 VTAIL.n59 0.155672
R1008 VTAIL.n60 VTAIL.n19 0.155672
R1009 VTAIL.n67 VTAIL.n19 0.155672
R1010 VTAIL.n68 VTAIL.n67 0.155672
R1011 VTAIL.n68 VTAIL.n15 0.155672
R1012 VTAIL.n75 VTAIL.n15 0.155672
R1013 VTAIL.n76 VTAIL.n75 0.155672
R1014 VTAIL.n76 VTAIL.n11 0.155672
R1015 VTAIL.n85 VTAIL.n11 0.155672
R1016 VTAIL.n86 VTAIL.n85 0.155672
R1017 VTAIL.n86 VTAIL.n7 0.155672
R1018 VTAIL.n93 VTAIL.n7 0.155672
R1019 VTAIL.n94 VTAIL.n93 0.155672
R1020 VTAIL.n94 VTAIL.n3 0.155672
R1021 VTAIL.n101 VTAIL.n3 0.155672
R1022 VTAIL.n317 VTAIL.n219 0.155672
R1023 VTAIL.n310 VTAIL.n219 0.155672
R1024 VTAIL.n310 VTAIL.n309 0.155672
R1025 VTAIL.n309 VTAIL.n223 0.155672
R1026 VTAIL.n302 VTAIL.n223 0.155672
R1027 VTAIL.n302 VTAIL.n301 0.155672
R1028 VTAIL.n301 VTAIL.n227 0.155672
R1029 VTAIL.n293 VTAIL.n227 0.155672
R1030 VTAIL.n293 VTAIL.n292 0.155672
R1031 VTAIL.n292 VTAIL.n232 0.155672
R1032 VTAIL.n285 VTAIL.n232 0.155672
R1033 VTAIL.n285 VTAIL.n284 0.155672
R1034 VTAIL.n284 VTAIL.n236 0.155672
R1035 VTAIL.n277 VTAIL.n236 0.155672
R1036 VTAIL.n277 VTAIL.n276 0.155672
R1037 VTAIL.n276 VTAIL.n240 0.155672
R1038 VTAIL.n269 VTAIL.n240 0.155672
R1039 VTAIL.n269 VTAIL.n268 0.155672
R1040 VTAIL.n268 VTAIL.n244 0.155672
R1041 VTAIL.n261 VTAIL.n244 0.155672
R1042 VTAIL.n261 VTAIL.n260 0.155672
R1043 VTAIL.n260 VTAIL.n248 0.155672
R1044 VTAIL.n253 VTAIL.n248 0.155672
R1045 VTAIL.n211 VTAIL.n113 0.155672
R1046 VTAIL.n204 VTAIL.n113 0.155672
R1047 VTAIL.n204 VTAIL.n203 0.155672
R1048 VTAIL.n203 VTAIL.n117 0.155672
R1049 VTAIL.n196 VTAIL.n117 0.155672
R1050 VTAIL.n196 VTAIL.n195 0.155672
R1051 VTAIL.n195 VTAIL.n121 0.155672
R1052 VTAIL.n187 VTAIL.n121 0.155672
R1053 VTAIL.n187 VTAIL.n186 0.155672
R1054 VTAIL.n186 VTAIL.n126 0.155672
R1055 VTAIL.n179 VTAIL.n126 0.155672
R1056 VTAIL.n179 VTAIL.n178 0.155672
R1057 VTAIL.n178 VTAIL.n130 0.155672
R1058 VTAIL.n171 VTAIL.n130 0.155672
R1059 VTAIL.n171 VTAIL.n170 0.155672
R1060 VTAIL.n170 VTAIL.n134 0.155672
R1061 VTAIL.n163 VTAIL.n134 0.155672
R1062 VTAIL.n163 VTAIL.n162 0.155672
R1063 VTAIL.n162 VTAIL.n138 0.155672
R1064 VTAIL.n155 VTAIL.n138 0.155672
R1065 VTAIL.n155 VTAIL.n154 0.155672
R1066 VTAIL.n154 VTAIL.n142 0.155672
R1067 VTAIL.n147 VTAIL.n142 0.155672
R1068 B.n972 B.n971 585
R1069 B.n398 B.n138 585
R1070 B.n397 B.n396 585
R1071 B.n395 B.n394 585
R1072 B.n393 B.n392 585
R1073 B.n391 B.n390 585
R1074 B.n389 B.n388 585
R1075 B.n387 B.n386 585
R1076 B.n385 B.n384 585
R1077 B.n383 B.n382 585
R1078 B.n381 B.n380 585
R1079 B.n379 B.n378 585
R1080 B.n377 B.n376 585
R1081 B.n375 B.n374 585
R1082 B.n373 B.n372 585
R1083 B.n371 B.n370 585
R1084 B.n369 B.n368 585
R1085 B.n367 B.n366 585
R1086 B.n365 B.n364 585
R1087 B.n363 B.n362 585
R1088 B.n361 B.n360 585
R1089 B.n359 B.n358 585
R1090 B.n357 B.n356 585
R1091 B.n355 B.n354 585
R1092 B.n353 B.n352 585
R1093 B.n351 B.n350 585
R1094 B.n349 B.n348 585
R1095 B.n347 B.n346 585
R1096 B.n345 B.n344 585
R1097 B.n343 B.n342 585
R1098 B.n341 B.n340 585
R1099 B.n339 B.n338 585
R1100 B.n337 B.n336 585
R1101 B.n335 B.n334 585
R1102 B.n333 B.n332 585
R1103 B.n331 B.n330 585
R1104 B.n329 B.n328 585
R1105 B.n327 B.n326 585
R1106 B.n325 B.n324 585
R1107 B.n323 B.n322 585
R1108 B.n321 B.n320 585
R1109 B.n319 B.n318 585
R1110 B.n317 B.n316 585
R1111 B.n315 B.n314 585
R1112 B.n313 B.n312 585
R1113 B.n311 B.n310 585
R1114 B.n309 B.n308 585
R1115 B.n307 B.n306 585
R1116 B.n305 B.n304 585
R1117 B.n303 B.n302 585
R1118 B.n301 B.n300 585
R1119 B.n299 B.n298 585
R1120 B.n297 B.n296 585
R1121 B.n295 B.n294 585
R1122 B.n293 B.n292 585
R1123 B.n291 B.n290 585
R1124 B.n289 B.n288 585
R1125 B.n287 B.n286 585
R1126 B.n285 B.n284 585
R1127 B.n283 B.n282 585
R1128 B.n281 B.n280 585
R1129 B.n279 B.n278 585
R1130 B.n277 B.n276 585
R1131 B.n275 B.n274 585
R1132 B.n273 B.n272 585
R1133 B.n271 B.n270 585
R1134 B.n269 B.n268 585
R1135 B.n267 B.n266 585
R1136 B.n265 B.n264 585
R1137 B.n263 B.n262 585
R1138 B.n261 B.n260 585
R1139 B.n259 B.n258 585
R1140 B.n257 B.n256 585
R1141 B.n255 B.n254 585
R1142 B.n253 B.n252 585
R1143 B.n251 B.n250 585
R1144 B.n249 B.n248 585
R1145 B.n247 B.n246 585
R1146 B.n245 B.n244 585
R1147 B.n243 B.n242 585
R1148 B.n241 B.n240 585
R1149 B.n239 B.n238 585
R1150 B.n237 B.n236 585
R1151 B.n235 B.n234 585
R1152 B.n233 B.n232 585
R1153 B.n231 B.n230 585
R1154 B.n229 B.n228 585
R1155 B.n227 B.n226 585
R1156 B.n225 B.n224 585
R1157 B.n223 B.n222 585
R1158 B.n221 B.n220 585
R1159 B.n219 B.n218 585
R1160 B.n217 B.n216 585
R1161 B.n215 B.n214 585
R1162 B.n213 B.n212 585
R1163 B.n211 B.n210 585
R1164 B.n209 B.n208 585
R1165 B.n207 B.n206 585
R1166 B.n205 B.n204 585
R1167 B.n203 B.n202 585
R1168 B.n201 B.n200 585
R1169 B.n199 B.n198 585
R1170 B.n197 B.n196 585
R1171 B.n195 B.n194 585
R1172 B.n193 B.n192 585
R1173 B.n191 B.n190 585
R1174 B.n189 B.n188 585
R1175 B.n187 B.n186 585
R1176 B.n185 B.n184 585
R1177 B.n183 B.n182 585
R1178 B.n181 B.n180 585
R1179 B.n179 B.n178 585
R1180 B.n177 B.n176 585
R1181 B.n175 B.n174 585
R1182 B.n173 B.n172 585
R1183 B.n171 B.n170 585
R1184 B.n169 B.n168 585
R1185 B.n167 B.n166 585
R1186 B.n165 B.n164 585
R1187 B.n163 B.n162 585
R1188 B.n161 B.n160 585
R1189 B.n159 B.n158 585
R1190 B.n157 B.n156 585
R1191 B.n155 B.n154 585
R1192 B.n153 B.n152 585
R1193 B.n151 B.n150 585
R1194 B.n149 B.n148 585
R1195 B.n147 B.n146 585
R1196 B.n74 B.n73 585
R1197 B.n977 B.n976 585
R1198 B.n970 B.n139 585
R1199 B.n139 B.n71 585
R1200 B.n969 B.n70 585
R1201 B.n981 B.n70 585
R1202 B.n968 B.n69 585
R1203 B.n982 B.n69 585
R1204 B.n967 B.n68 585
R1205 B.n983 B.n68 585
R1206 B.n966 B.n965 585
R1207 B.n965 B.n64 585
R1208 B.n964 B.n63 585
R1209 B.n989 B.n63 585
R1210 B.n963 B.n62 585
R1211 B.n990 B.n62 585
R1212 B.n962 B.n61 585
R1213 B.n991 B.n61 585
R1214 B.n961 B.n960 585
R1215 B.n960 B.n57 585
R1216 B.n959 B.n56 585
R1217 B.n997 B.n56 585
R1218 B.n958 B.n55 585
R1219 B.n998 B.n55 585
R1220 B.n957 B.n54 585
R1221 B.n999 B.n54 585
R1222 B.n956 B.n955 585
R1223 B.n955 B.n50 585
R1224 B.n954 B.n49 585
R1225 B.n1005 B.n49 585
R1226 B.n953 B.n48 585
R1227 B.n1006 B.n48 585
R1228 B.n952 B.n47 585
R1229 B.n1007 B.n47 585
R1230 B.n951 B.n950 585
R1231 B.n950 B.n43 585
R1232 B.n949 B.n42 585
R1233 B.n1013 B.n42 585
R1234 B.n948 B.n41 585
R1235 B.n1014 B.n41 585
R1236 B.n947 B.n40 585
R1237 B.n1015 B.n40 585
R1238 B.n946 B.n945 585
R1239 B.n945 B.n36 585
R1240 B.n944 B.n35 585
R1241 B.n1021 B.n35 585
R1242 B.n943 B.n34 585
R1243 B.n1022 B.n34 585
R1244 B.n942 B.n33 585
R1245 B.n1023 B.n33 585
R1246 B.n941 B.n940 585
R1247 B.n940 B.n32 585
R1248 B.n939 B.n28 585
R1249 B.n1029 B.n28 585
R1250 B.n938 B.n27 585
R1251 B.n1030 B.n27 585
R1252 B.n937 B.n26 585
R1253 B.n1031 B.n26 585
R1254 B.n936 B.n935 585
R1255 B.n935 B.n22 585
R1256 B.n934 B.n21 585
R1257 B.n1037 B.n21 585
R1258 B.n933 B.n20 585
R1259 B.n1038 B.n20 585
R1260 B.n932 B.n19 585
R1261 B.n1039 B.n19 585
R1262 B.n931 B.n930 585
R1263 B.n930 B.n15 585
R1264 B.n929 B.n14 585
R1265 B.n1045 B.n14 585
R1266 B.n928 B.n13 585
R1267 B.n1046 B.n13 585
R1268 B.n927 B.n12 585
R1269 B.n1047 B.n12 585
R1270 B.n926 B.n925 585
R1271 B.n925 B.n8 585
R1272 B.n924 B.n7 585
R1273 B.n1053 B.n7 585
R1274 B.n923 B.n6 585
R1275 B.n1054 B.n6 585
R1276 B.n922 B.n5 585
R1277 B.n1055 B.n5 585
R1278 B.n921 B.n920 585
R1279 B.n920 B.n4 585
R1280 B.n919 B.n399 585
R1281 B.n919 B.n918 585
R1282 B.n909 B.n400 585
R1283 B.n401 B.n400 585
R1284 B.n911 B.n910 585
R1285 B.n912 B.n911 585
R1286 B.n908 B.n405 585
R1287 B.n409 B.n405 585
R1288 B.n907 B.n906 585
R1289 B.n906 B.n905 585
R1290 B.n407 B.n406 585
R1291 B.n408 B.n407 585
R1292 B.n898 B.n897 585
R1293 B.n899 B.n898 585
R1294 B.n896 B.n414 585
R1295 B.n414 B.n413 585
R1296 B.n895 B.n894 585
R1297 B.n894 B.n893 585
R1298 B.n416 B.n415 585
R1299 B.n417 B.n416 585
R1300 B.n886 B.n885 585
R1301 B.n887 B.n886 585
R1302 B.n884 B.n422 585
R1303 B.n422 B.n421 585
R1304 B.n883 B.n882 585
R1305 B.n882 B.n881 585
R1306 B.n424 B.n423 585
R1307 B.n874 B.n424 585
R1308 B.n873 B.n872 585
R1309 B.n875 B.n873 585
R1310 B.n871 B.n429 585
R1311 B.n429 B.n428 585
R1312 B.n870 B.n869 585
R1313 B.n869 B.n868 585
R1314 B.n431 B.n430 585
R1315 B.n432 B.n431 585
R1316 B.n861 B.n860 585
R1317 B.n862 B.n861 585
R1318 B.n859 B.n437 585
R1319 B.n437 B.n436 585
R1320 B.n858 B.n857 585
R1321 B.n857 B.n856 585
R1322 B.n439 B.n438 585
R1323 B.n440 B.n439 585
R1324 B.n849 B.n848 585
R1325 B.n850 B.n849 585
R1326 B.n847 B.n444 585
R1327 B.n448 B.n444 585
R1328 B.n846 B.n845 585
R1329 B.n845 B.n844 585
R1330 B.n446 B.n445 585
R1331 B.n447 B.n446 585
R1332 B.n837 B.n836 585
R1333 B.n838 B.n837 585
R1334 B.n835 B.n453 585
R1335 B.n453 B.n452 585
R1336 B.n834 B.n833 585
R1337 B.n833 B.n832 585
R1338 B.n455 B.n454 585
R1339 B.n456 B.n455 585
R1340 B.n825 B.n824 585
R1341 B.n826 B.n825 585
R1342 B.n823 B.n460 585
R1343 B.n464 B.n460 585
R1344 B.n822 B.n821 585
R1345 B.n821 B.n820 585
R1346 B.n462 B.n461 585
R1347 B.n463 B.n462 585
R1348 B.n813 B.n812 585
R1349 B.n814 B.n813 585
R1350 B.n811 B.n469 585
R1351 B.n469 B.n468 585
R1352 B.n810 B.n809 585
R1353 B.n809 B.n808 585
R1354 B.n471 B.n470 585
R1355 B.n472 B.n471 585
R1356 B.n804 B.n803 585
R1357 B.n475 B.n474 585
R1358 B.n800 B.n799 585
R1359 B.n801 B.n800 585
R1360 B.n798 B.n540 585
R1361 B.n797 B.n796 585
R1362 B.n795 B.n794 585
R1363 B.n793 B.n792 585
R1364 B.n791 B.n790 585
R1365 B.n789 B.n788 585
R1366 B.n787 B.n786 585
R1367 B.n785 B.n784 585
R1368 B.n783 B.n782 585
R1369 B.n781 B.n780 585
R1370 B.n779 B.n778 585
R1371 B.n777 B.n776 585
R1372 B.n775 B.n774 585
R1373 B.n773 B.n772 585
R1374 B.n771 B.n770 585
R1375 B.n769 B.n768 585
R1376 B.n767 B.n766 585
R1377 B.n765 B.n764 585
R1378 B.n763 B.n762 585
R1379 B.n761 B.n760 585
R1380 B.n759 B.n758 585
R1381 B.n757 B.n756 585
R1382 B.n755 B.n754 585
R1383 B.n753 B.n752 585
R1384 B.n751 B.n750 585
R1385 B.n749 B.n748 585
R1386 B.n747 B.n746 585
R1387 B.n745 B.n744 585
R1388 B.n743 B.n742 585
R1389 B.n741 B.n740 585
R1390 B.n739 B.n738 585
R1391 B.n737 B.n736 585
R1392 B.n735 B.n734 585
R1393 B.n733 B.n732 585
R1394 B.n731 B.n730 585
R1395 B.n729 B.n728 585
R1396 B.n727 B.n726 585
R1397 B.n725 B.n724 585
R1398 B.n723 B.n722 585
R1399 B.n721 B.n720 585
R1400 B.n719 B.n718 585
R1401 B.n717 B.n716 585
R1402 B.n715 B.n714 585
R1403 B.n713 B.n712 585
R1404 B.n711 B.n710 585
R1405 B.n709 B.n708 585
R1406 B.n707 B.n706 585
R1407 B.n705 B.n704 585
R1408 B.n703 B.n702 585
R1409 B.n701 B.n700 585
R1410 B.n699 B.n698 585
R1411 B.n697 B.n696 585
R1412 B.n695 B.n694 585
R1413 B.n693 B.n692 585
R1414 B.n691 B.n690 585
R1415 B.n689 B.n688 585
R1416 B.n687 B.n686 585
R1417 B.n684 B.n683 585
R1418 B.n682 B.n681 585
R1419 B.n680 B.n679 585
R1420 B.n678 B.n677 585
R1421 B.n676 B.n675 585
R1422 B.n674 B.n673 585
R1423 B.n672 B.n671 585
R1424 B.n670 B.n669 585
R1425 B.n668 B.n667 585
R1426 B.n666 B.n665 585
R1427 B.n663 B.n662 585
R1428 B.n661 B.n660 585
R1429 B.n659 B.n658 585
R1430 B.n657 B.n656 585
R1431 B.n655 B.n654 585
R1432 B.n653 B.n652 585
R1433 B.n651 B.n650 585
R1434 B.n649 B.n648 585
R1435 B.n647 B.n646 585
R1436 B.n645 B.n644 585
R1437 B.n643 B.n642 585
R1438 B.n641 B.n640 585
R1439 B.n639 B.n638 585
R1440 B.n637 B.n636 585
R1441 B.n635 B.n634 585
R1442 B.n633 B.n632 585
R1443 B.n631 B.n630 585
R1444 B.n629 B.n628 585
R1445 B.n627 B.n626 585
R1446 B.n625 B.n624 585
R1447 B.n623 B.n622 585
R1448 B.n621 B.n620 585
R1449 B.n619 B.n618 585
R1450 B.n617 B.n616 585
R1451 B.n615 B.n614 585
R1452 B.n613 B.n612 585
R1453 B.n611 B.n610 585
R1454 B.n609 B.n608 585
R1455 B.n607 B.n606 585
R1456 B.n605 B.n604 585
R1457 B.n603 B.n602 585
R1458 B.n601 B.n600 585
R1459 B.n599 B.n598 585
R1460 B.n597 B.n596 585
R1461 B.n595 B.n594 585
R1462 B.n593 B.n592 585
R1463 B.n591 B.n590 585
R1464 B.n589 B.n588 585
R1465 B.n587 B.n586 585
R1466 B.n585 B.n584 585
R1467 B.n583 B.n582 585
R1468 B.n581 B.n580 585
R1469 B.n579 B.n578 585
R1470 B.n577 B.n576 585
R1471 B.n575 B.n574 585
R1472 B.n573 B.n572 585
R1473 B.n571 B.n570 585
R1474 B.n569 B.n568 585
R1475 B.n567 B.n566 585
R1476 B.n565 B.n564 585
R1477 B.n563 B.n562 585
R1478 B.n561 B.n560 585
R1479 B.n559 B.n558 585
R1480 B.n557 B.n556 585
R1481 B.n555 B.n554 585
R1482 B.n553 B.n552 585
R1483 B.n551 B.n550 585
R1484 B.n549 B.n548 585
R1485 B.n547 B.n546 585
R1486 B.n545 B.n539 585
R1487 B.n801 B.n539 585
R1488 B.n805 B.n473 585
R1489 B.n473 B.n472 585
R1490 B.n807 B.n806 585
R1491 B.n808 B.n807 585
R1492 B.n467 B.n466 585
R1493 B.n468 B.n467 585
R1494 B.n816 B.n815 585
R1495 B.n815 B.n814 585
R1496 B.n817 B.n465 585
R1497 B.n465 B.n463 585
R1498 B.n819 B.n818 585
R1499 B.n820 B.n819 585
R1500 B.n459 B.n458 585
R1501 B.n464 B.n459 585
R1502 B.n828 B.n827 585
R1503 B.n827 B.n826 585
R1504 B.n829 B.n457 585
R1505 B.n457 B.n456 585
R1506 B.n831 B.n830 585
R1507 B.n832 B.n831 585
R1508 B.n451 B.n450 585
R1509 B.n452 B.n451 585
R1510 B.n840 B.n839 585
R1511 B.n839 B.n838 585
R1512 B.n841 B.n449 585
R1513 B.n449 B.n447 585
R1514 B.n843 B.n842 585
R1515 B.n844 B.n843 585
R1516 B.n443 B.n442 585
R1517 B.n448 B.n443 585
R1518 B.n852 B.n851 585
R1519 B.n851 B.n850 585
R1520 B.n853 B.n441 585
R1521 B.n441 B.n440 585
R1522 B.n855 B.n854 585
R1523 B.n856 B.n855 585
R1524 B.n435 B.n434 585
R1525 B.n436 B.n435 585
R1526 B.n864 B.n863 585
R1527 B.n863 B.n862 585
R1528 B.n865 B.n433 585
R1529 B.n433 B.n432 585
R1530 B.n867 B.n866 585
R1531 B.n868 B.n867 585
R1532 B.n427 B.n426 585
R1533 B.n428 B.n427 585
R1534 B.n877 B.n876 585
R1535 B.n876 B.n875 585
R1536 B.n878 B.n425 585
R1537 B.n874 B.n425 585
R1538 B.n880 B.n879 585
R1539 B.n881 B.n880 585
R1540 B.n420 B.n419 585
R1541 B.n421 B.n420 585
R1542 B.n889 B.n888 585
R1543 B.n888 B.n887 585
R1544 B.n890 B.n418 585
R1545 B.n418 B.n417 585
R1546 B.n892 B.n891 585
R1547 B.n893 B.n892 585
R1548 B.n412 B.n411 585
R1549 B.n413 B.n412 585
R1550 B.n901 B.n900 585
R1551 B.n900 B.n899 585
R1552 B.n902 B.n410 585
R1553 B.n410 B.n408 585
R1554 B.n904 B.n903 585
R1555 B.n905 B.n904 585
R1556 B.n404 B.n403 585
R1557 B.n409 B.n404 585
R1558 B.n914 B.n913 585
R1559 B.n913 B.n912 585
R1560 B.n915 B.n402 585
R1561 B.n402 B.n401 585
R1562 B.n917 B.n916 585
R1563 B.n918 B.n917 585
R1564 B.n2 B.n0 585
R1565 B.n4 B.n2 585
R1566 B.n3 B.n1 585
R1567 B.n1054 B.n3 585
R1568 B.n1052 B.n1051 585
R1569 B.n1053 B.n1052 585
R1570 B.n1050 B.n9 585
R1571 B.n9 B.n8 585
R1572 B.n1049 B.n1048 585
R1573 B.n1048 B.n1047 585
R1574 B.n11 B.n10 585
R1575 B.n1046 B.n11 585
R1576 B.n1044 B.n1043 585
R1577 B.n1045 B.n1044 585
R1578 B.n1042 B.n16 585
R1579 B.n16 B.n15 585
R1580 B.n1041 B.n1040 585
R1581 B.n1040 B.n1039 585
R1582 B.n18 B.n17 585
R1583 B.n1038 B.n18 585
R1584 B.n1036 B.n1035 585
R1585 B.n1037 B.n1036 585
R1586 B.n1034 B.n23 585
R1587 B.n23 B.n22 585
R1588 B.n1033 B.n1032 585
R1589 B.n1032 B.n1031 585
R1590 B.n25 B.n24 585
R1591 B.n1030 B.n25 585
R1592 B.n1028 B.n1027 585
R1593 B.n1029 B.n1028 585
R1594 B.n1026 B.n29 585
R1595 B.n32 B.n29 585
R1596 B.n1025 B.n1024 585
R1597 B.n1024 B.n1023 585
R1598 B.n31 B.n30 585
R1599 B.n1022 B.n31 585
R1600 B.n1020 B.n1019 585
R1601 B.n1021 B.n1020 585
R1602 B.n1018 B.n37 585
R1603 B.n37 B.n36 585
R1604 B.n1017 B.n1016 585
R1605 B.n1016 B.n1015 585
R1606 B.n39 B.n38 585
R1607 B.n1014 B.n39 585
R1608 B.n1012 B.n1011 585
R1609 B.n1013 B.n1012 585
R1610 B.n1010 B.n44 585
R1611 B.n44 B.n43 585
R1612 B.n1009 B.n1008 585
R1613 B.n1008 B.n1007 585
R1614 B.n46 B.n45 585
R1615 B.n1006 B.n46 585
R1616 B.n1004 B.n1003 585
R1617 B.n1005 B.n1004 585
R1618 B.n1002 B.n51 585
R1619 B.n51 B.n50 585
R1620 B.n1001 B.n1000 585
R1621 B.n1000 B.n999 585
R1622 B.n53 B.n52 585
R1623 B.n998 B.n53 585
R1624 B.n996 B.n995 585
R1625 B.n997 B.n996 585
R1626 B.n994 B.n58 585
R1627 B.n58 B.n57 585
R1628 B.n993 B.n992 585
R1629 B.n992 B.n991 585
R1630 B.n60 B.n59 585
R1631 B.n990 B.n60 585
R1632 B.n988 B.n987 585
R1633 B.n989 B.n988 585
R1634 B.n986 B.n65 585
R1635 B.n65 B.n64 585
R1636 B.n985 B.n984 585
R1637 B.n984 B.n983 585
R1638 B.n67 B.n66 585
R1639 B.n982 B.n67 585
R1640 B.n980 B.n979 585
R1641 B.n981 B.n980 585
R1642 B.n978 B.n72 585
R1643 B.n72 B.n71 585
R1644 B.n1057 B.n1056 585
R1645 B.n1056 B.n1055 585
R1646 B.n543 B.t10 517.021
R1647 B.n541 B.t21 517.021
R1648 B.n143 B.t18 517.021
R1649 B.n140 B.t14 517.021
R1650 B.n803 B.n473 434.841
R1651 B.n976 B.n72 434.841
R1652 B.n539 B.n471 434.841
R1653 B.n972 B.n139 434.841
R1654 B.n543 B.t13 423.687
R1655 B.n541 B.t23 423.687
R1656 B.n143 B.t19 423.687
R1657 B.n140 B.t16 423.687
R1658 B.n544 B.t12 389.942
R1659 B.n141 B.t17 389.942
R1660 B.n542 B.t22 389.94
R1661 B.n144 B.t20 389.94
R1662 B.n974 B.n973 256.663
R1663 B.n974 B.n137 256.663
R1664 B.n974 B.n136 256.663
R1665 B.n974 B.n135 256.663
R1666 B.n974 B.n134 256.663
R1667 B.n974 B.n133 256.663
R1668 B.n974 B.n132 256.663
R1669 B.n974 B.n131 256.663
R1670 B.n974 B.n130 256.663
R1671 B.n974 B.n129 256.663
R1672 B.n974 B.n128 256.663
R1673 B.n974 B.n127 256.663
R1674 B.n974 B.n126 256.663
R1675 B.n974 B.n125 256.663
R1676 B.n974 B.n124 256.663
R1677 B.n974 B.n123 256.663
R1678 B.n974 B.n122 256.663
R1679 B.n974 B.n121 256.663
R1680 B.n974 B.n120 256.663
R1681 B.n974 B.n119 256.663
R1682 B.n974 B.n118 256.663
R1683 B.n974 B.n117 256.663
R1684 B.n974 B.n116 256.663
R1685 B.n974 B.n115 256.663
R1686 B.n974 B.n114 256.663
R1687 B.n974 B.n113 256.663
R1688 B.n974 B.n112 256.663
R1689 B.n974 B.n111 256.663
R1690 B.n974 B.n110 256.663
R1691 B.n974 B.n109 256.663
R1692 B.n974 B.n108 256.663
R1693 B.n974 B.n107 256.663
R1694 B.n974 B.n106 256.663
R1695 B.n974 B.n105 256.663
R1696 B.n974 B.n104 256.663
R1697 B.n974 B.n103 256.663
R1698 B.n974 B.n102 256.663
R1699 B.n974 B.n101 256.663
R1700 B.n974 B.n100 256.663
R1701 B.n974 B.n99 256.663
R1702 B.n974 B.n98 256.663
R1703 B.n974 B.n97 256.663
R1704 B.n974 B.n96 256.663
R1705 B.n974 B.n95 256.663
R1706 B.n974 B.n94 256.663
R1707 B.n974 B.n93 256.663
R1708 B.n974 B.n92 256.663
R1709 B.n974 B.n91 256.663
R1710 B.n974 B.n90 256.663
R1711 B.n974 B.n89 256.663
R1712 B.n974 B.n88 256.663
R1713 B.n974 B.n87 256.663
R1714 B.n974 B.n86 256.663
R1715 B.n974 B.n85 256.663
R1716 B.n974 B.n84 256.663
R1717 B.n974 B.n83 256.663
R1718 B.n974 B.n82 256.663
R1719 B.n974 B.n81 256.663
R1720 B.n974 B.n80 256.663
R1721 B.n974 B.n79 256.663
R1722 B.n974 B.n78 256.663
R1723 B.n974 B.n77 256.663
R1724 B.n974 B.n76 256.663
R1725 B.n974 B.n75 256.663
R1726 B.n975 B.n974 256.663
R1727 B.n802 B.n801 256.663
R1728 B.n801 B.n476 256.663
R1729 B.n801 B.n477 256.663
R1730 B.n801 B.n478 256.663
R1731 B.n801 B.n479 256.663
R1732 B.n801 B.n480 256.663
R1733 B.n801 B.n481 256.663
R1734 B.n801 B.n482 256.663
R1735 B.n801 B.n483 256.663
R1736 B.n801 B.n484 256.663
R1737 B.n801 B.n485 256.663
R1738 B.n801 B.n486 256.663
R1739 B.n801 B.n487 256.663
R1740 B.n801 B.n488 256.663
R1741 B.n801 B.n489 256.663
R1742 B.n801 B.n490 256.663
R1743 B.n801 B.n491 256.663
R1744 B.n801 B.n492 256.663
R1745 B.n801 B.n493 256.663
R1746 B.n801 B.n494 256.663
R1747 B.n801 B.n495 256.663
R1748 B.n801 B.n496 256.663
R1749 B.n801 B.n497 256.663
R1750 B.n801 B.n498 256.663
R1751 B.n801 B.n499 256.663
R1752 B.n801 B.n500 256.663
R1753 B.n801 B.n501 256.663
R1754 B.n801 B.n502 256.663
R1755 B.n801 B.n503 256.663
R1756 B.n801 B.n504 256.663
R1757 B.n801 B.n505 256.663
R1758 B.n801 B.n506 256.663
R1759 B.n801 B.n507 256.663
R1760 B.n801 B.n508 256.663
R1761 B.n801 B.n509 256.663
R1762 B.n801 B.n510 256.663
R1763 B.n801 B.n511 256.663
R1764 B.n801 B.n512 256.663
R1765 B.n801 B.n513 256.663
R1766 B.n801 B.n514 256.663
R1767 B.n801 B.n515 256.663
R1768 B.n801 B.n516 256.663
R1769 B.n801 B.n517 256.663
R1770 B.n801 B.n518 256.663
R1771 B.n801 B.n519 256.663
R1772 B.n801 B.n520 256.663
R1773 B.n801 B.n521 256.663
R1774 B.n801 B.n522 256.663
R1775 B.n801 B.n523 256.663
R1776 B.n801 B.n524 256.663
R1777 B.n801 B.n525 256.663
R1778 B.n801 B.n526 256.663
R1779 B.n801 B.n527 256.663
R1780 B.n801 B.n528 256.663
R1781 B.n801 B.n529 256.663
R1782 B.n801 B.n530 256.663
R1783 B.n801 B.n531 256.663
R1784 B.n801 B.n532 256.663
R1785 B.n801 B.n533 256.663
R1786 B.n801 B.n534 256.663
R1787 B.n801 B.n535 256.663
R1788 B.n801 B.n536 256.663
R1789 B.n801 B.n537 256.663
R1790 B.n801 B.n538 256.663
R1791 B.n807 B.n473 163.367
R1792 B.n807 B.n467 163.367
R1793 B.n815 B.n467 163.367
R1794 B.n815 B.n465 163.367
R1795 B.n819 B.n465 163.367
R1796 B.n819 B.n459 163.367
R1797 B.n827 B.n459 163.367
R1798 B.n827 B.n457 163.367
R1799 B.n831 B.n457 163.367
R1800 B.n831 B.n451 163.367
R1801 B.n839 B.n451 163.367
R1802 B.n839 B.n449 163.367
R1803 B.n843 B.n449 163.367
R1804 B.n843 B.n443 163.367
R1805 B.n851 B.n443 163.367
R1806 B.n851 B.n441 163.367
R1807 B.n855 B.n441 163.367
R1808 B.n855 B.n435 163.367
R1809 B.n863 B.n435 163.367
R1810 B.n863 B.n433 163.367
R1811 B.n867 B.n433 163.367
R1812 B.n867 B.n427 163.367
R1813 B.n876 B.n427 163.367
R1814 B.n876 B.n425 163.367
R1815 B.n880 B.n425 163.367
R1816 B.n880 B.n420 163.367
R1817 B.n888 B.n420 163.367
R1818 B.n888 B.n418 163.367
R1819 B.n892 B.n418 163.367
R1820 B.n892 B.n412 163.367
R1821 B.n900 B.n412 163.367
R1822 B.n900 B.n410 163.367
R1823 B.n904 B.n410 163.367
R1824 B.n904 B.n404 163.367
R1825 B.n913 B.n404 163.367
R1826 B.n913 B.n402 163.367
R1827 B.n917 B.n402 163.367
R1828 B.n917 B.n2 163.367
R1829 B.n1056 B.n2 163.367
R1830 B.n1056 B.n3 163.367
R1831 B.n1052 B.n3 163.367
R1832 B.n1052 B.n9 163.367
R1833 B.n1048 B.n9 163.367
R1834 B.n1048 B.n11 163.367
R1835 B.n1044 B.n11 163.367
R1836 B.n1044 B.n16 163.367
R1837 B.n1040 B.n16 163.367
R1838 B.n1040 B.n18 163.367
R1839 B.n1036 B.n18 163.367
R1840 B.n1036 B.n23 163.367
R1841 B.n1032 B.n23 163.367
R1842 B.n1032 B.n25 163.367
R1843 B.n1028 B.n25 163.367
R1844 B.n1028 B.n29 163.367
R1845 B.n1024 B.n29 163.367
R1846 B.n1024 B.n31 163.367
R1847 B.n1020 B.n31 163.367
R1848 B.n1020 B.n37 163.367
R1849 B.n1016 B.n37 163.367
R1850 B.n1016 B.n39 163.367
R1851 B.n1012 B.n39 163.367
R1852 B.n1012 B.n44 163.367
R1853 B.n1008 B.n44 163.367
R1854 B.n1008 B.n46 163.367
R1855 B.n1004 B.n46 163.367
R1856 B.n1004 B.n51 163.367
R1857 B.n1000 B.n51 163.367
R1858 B.n1000 B.n53 163.367
R1859 B.n996 B.n53 163.367
R1860 B.n996 B.n58 163.367
R1861 B.n992 B.n58 163.367
R1862 B.n992 B.n60 163.367
R1863 B.n988 B.n60 163.367
R1864 B.n988 B.n65 163.367
R1865 B.n984 B.n65 163.367
R1866 B.n984 B.n67 163.367
R1867 B.n980 B.n67 163.367
R1868 B.n980 B.n72 163.367
R1869 B.n800 B.n475 163.367
R1870 B.n800 B.n540 163.367
R1871 B.n796 B.n795 163.367
R1872 B.n792 B.n791 163.367
R1873 B.n788 B.n787 163.367
R1874 B.n784 B.n783 163.367
R1875 B.n780 B.n779 163.367
R1876 B.n776 B.n775 163.367
R1877 B.n772 B.n771 163.367
R1878 B.n768 B.n767 163.367
R1879 B.n764 B.n763 163.367
R1880 B.n760 B.n759 163.367
R1881 B.n756 B.n755 163.367
R1882 B.n752 B.n751 163.367
R1883 B.n748 B.n747 163.367
R1884 B.n744 B.n743 163.367
R1885 B.n740 B.n739 163.367
R1886 B.n736 B.n735 163.367
R1887 B.n732 B.n731 163.367
R1888 B.n728 B.n727 163.367
R1889 B.n724 B.n723 163.367
R1890 B.n720 B.n719 163.367
R1891 B.n716 B.n715 163.367
R1892 B.n712 B.n711 163.367
R1893 B.n708 B.n707 163.367
R1894 B.n704 B.n703 163.367
R1895 B.n700 B.n699 163.367
R1896 B.n696 B.n695 163.367
R1897 B.n692 B.n691 163.367
R1898 B.n688 B.n687 163.367
R1899 B.n683 B.n682 163.367
R1900 B.n679 B.n678 163.367
R1901 B.n675 B.n674 163.367
R1902 B.n671 B.n670 163.367
R1903 B.n667 B.n666 163.367
R1904 B.n662 B.n661 163.367
R1905 B.n658 B.n657 163.367
R1906 B.n654 B.n653 163.367
R1907 B.n650 B.n649 163.367
R1908 B.n646 B.n645 163.367
R1909 B.n642 B.n641 163.367
R1910 B.n638 B.n637 163.367
R1911 B.n634 B.n633 163.367
R1912 B.n630 B.n629 163.367
R1913 B.n626 B.n625 163.367
R1914 B.n622 B.n621 163.367
R1915 B.n618 B.n617 163.367
R1916 B.n614 B.n613 163.367
R1917 B.n610 B.n609 163.367
R1918 B.n606 B.n605 163.367
R1919 B.n602 B.n601 163.367
R1920 B.n598 B.n597 163.367
R1921 B.n594 B.n593 163.367
R1922 B.n590 B.n589 163.367
R1923 B.n586 B.n585 163.367
R1924 B.n582 B.n581 163.367
R1925 B.n578 B.n577 163.367
R1926 B.n574 B.n573 163.367
R1927 B.n570 B.n569 163.367
R1928 B.n566 B.n565 163.367
R1929 B.n562 B.n561 163.367
R1930 B.n558 B.n557 163.367
R1931 B.n554 B.n553 163.367
R1932 B.n550 B.n549 163.367
R1933 B.n546 B.n539 163.367
R1934 B.n809 B.n471 163.367
R1935 B.n809 B.n469 163.367
R1936 B.n813 B.n469 163.367
R1937 B.n813 B.n462 163.367
R1938 B.n821 B.n462 163.367
R1939 B.n821 B.n460 163.367
R1940 B.n825 B.n460 163.367
R1941 B.n825 B.n455 163.367
R1942 B.n833 B.n455 163.367
R1943 B.n833 B.n453 163.367
R1944 B.n837 B.n453 163.367
R1945 B.n837 B.n446 163.367
R1946 B.n845 B.n446 163.367
R1947 B.n845 B.n444 163.367
R1948 B.n849 B.n444 163.367
R1949 B.n849 B.n439 163.367
R1950 B.n857 B.n439 163.367
R1951 B.n857 B.n437 163.367
R1952 B.n861 B.n437 163.367
R1953 B.n861 B.n431 163.367
R1954 B.n869 B.n431 163.367
R1955 B.n869 B.n429 163.367
R1956 B.n873 B.n429 163.367
R1957 B.n873 B.n424 163.367
R1958 B.n882 B.n424 163.367
R1959 B.n882 B.n422 163.367
R1960 B.n886 B.n422 163.367
R1961 B.n886 B.n416 163.367
R1962 B.n894 B.n416 163.367
R1963 B.n894 B.n414 163.367
R1964 B.n898 B.n414 163.367
R1965 B.n898 B.n407 163.367
R1966 B.n906 B.n407 163.367
R1967 B.n906 B.n405 163.367
R1968 B.n911 B.n405 163.367
R1969 B.n911 B.n400 163.367
R1970 B.n919 B.n400 163.367
R1971 B.n920 B.n919 163.367
R1972 B.n920 B.n5 163.367
R1973 B.n6 B.n5 163.367
R1974 B.n7 B.n6 163.367
R1975 B.n925 B.n7 163.367
R1976 B.n925 B.n12 163.367
R1977 B.n13 B.n12 163.367
R1978 B.n14 B.n13 163.367
R1979 B.n930 B.n14 163.367
R1980 B.n930 B.n19 163.367
R1981 B.n20 B.n19 163.367
R1982 B.n21 B.n20 163.367
R1983 B.n935 B.n21 163.367
R1984 B.n935 B.n26 163.367
R1985 B.n27 B.n26 163.367
R1986 B.n28 B.n27 163.367
R1987 B.n940 B.n28 163.367
R1988 B.n940 B.n33 163.367
R1989 B.n34 B.n33 163.367
R1990 B.n35 B.n34 163.367
R1991 B.n945 B.n35 163.367
R1992 B.n945 B.n40 163.367
R1993 B.n41 B.n40 163.367
R1994 B.n42 B.n41 163.367
R1995 B.n950 B.n42 163.367
R1996 B.n950 B.n47 163.367
R1997 B.n48 B.n47 163.367
R1998 B.n49 B.n48 163.367
R1999 B.n955 B.n49 163.367
R2000 B.n955 B.n54 163.367
R2001 B.n55 B.n54 163.367
R2002 B.n56 B.n55 163.367
R2003 B.n960 B.n56 163.367
R2004 B.n960 B.n61 163.367
R2005 B.n62 B.n61 163.367
R2006 B.n63 B.n62 163.367
R2007 B.n965 B.n63 163.367
R2008 B.n965 B.n68 163.367
R2009 B.n69 B.n68 163.367
R2010 B.n70 B.n69 163.367
R2011 B.n139 B.n70 163.367
R2012 B.n146 B.n74 163.367
R2013 B.n150 B.n149 163.367
R2014 B.n154 B.n153 163.367
R2015 B.n158 B.n157 163.367
R2016 B.n162 B.n161 163.367
R2017 B.n166 B.n165 163.367
R2018 B.n170 B.n169 163.367
R2019 B.n174 B.n173 163.367
R2020 B.n178 B.n177 163.367
R2021 B.n182 B.n181 163.367
R2022 B.n186 B.n185 163.367
R2023 B.n190 B.n189 163.367
R2024 B.n194 B.n193 163.367
R2025 B.n198 B.n197 163.367
R2026 B.n202 B.n201 163.367
R2027 B.n206 B.n205 163.367
R2028 B.n210 B.n209 163.367
R2029 B.n214 B.n213 163.367
R2030 B.n218 B.n217 163.367
R2031 B.n222 B.n221 163.367
R2032 B.n226 B.n225 163.367
R2033 B.n230 B.n229 163.367
R2034 B.n234 B.n233 163.367
R2035 B.n238 B.n237 163.367
R2036 B.n242 B.n241 163.367
R2037 B.n246 B.n245 163.367
R2038 B.n250 B.n249 163.367
R2039 B.n254 B.n253 163.367
R2040 B.n258 B.n257 163.367
R2041 B.n262 B.n261 163.367
R2042 B.n266 B.n265 163.367
R2043 B.n270 B.n269 163.367
R2044 B.n274 B.n273 163.367
R2045 B.n278 B.n277 163.367
R2046 B.n282 B.n281 163.367
R2047 B.n286 B.n285 163.367
R2048 B.n290 B.n289 163.367
R2049 B.n294 B.n293 163.367
R2050 B.n298 B.n297 163.367
R2051 B.n302 B.n301 163.367
R2052 B.n306 B.n305 163.367
R2053 B.n310 B.n309 163.367
R2054 B.n314 B.n313 163.367
R2055 B.n318 B.n317 163.367
R2056 B.n322 B.n321 163.367
R2057 B.n326 B.n325 163.367
R2058 B.n330 B.n329 163.367
R2059 B.n334 B.n333 163.367
R2060 B.n338 B.n337 163.367
R2061 B.n342 B.n341 163.367
R2062 B.n346 B.n345 163.367
R2063 B.n350 B.n349 163.367
R2064 B.n354 B.n353 163.367
R2065 B.n358 B.n357 163.367
R2066 B.n362 B.n361 163.367
R2067 B.n366 B.n365 163.367
R2068 B.n370 B.n369 163.367
R2069 B.n374 B.n373 163.367
R2070 B.n378 B.n377 163.367
R2071 B.n382 B.n381 163.367
R2072 B.n386 B.n385 163.367
R2073 B.n390 B.n389 163.367
R2074 B.n394 B.n393 163.367
R2075 B.n396 B.n138 163.367
R2076 B.n803 B.n802 71.676
R2077 B.n540 B.n476 71.676
R2078 B.n795 B.n477 71.676
R2079 B.n791 B.n478 71.676
R2080 B.n787 B.n479 71.676
R2081 B.n783 B.n480 71.676
R2082 B.n779 B.n481 71.676
R2083 B.n775 B.n482 71.676
R2084 B.n771 B.n483 71.676
R2085 B.n767 B.n484 71.676
R2086 B.n763 B.n485 71.676
R2087 B.n759 B.n486 71.676
R2088 B.n755 B.n487 71.676
R2089 B.n751 B.n488 71.676
R2090 B.n747 B.n489 71.676
R2091 B.n743 B.n490 71.676
R2092 B.n739 B.n491 71.676
R2093 B.n735 B.n492 71.676
R2094 B.n731 B.n493 71.676
R2095 B.n727 B.n494 71.676
R2096 B.n723 B.n495 71.676
R2097 B.n719 B.n496 71.676
R2098 B.n715 B.n497 71.676
R2099 B.n711 B.n498 71.676
R2100 B.n707 B.n499 71.676
R2101 B.n703 B.n500 71.676
R2102 B.n699 B.n501 71.676
R2103 B.n695 B.n502 71.676
R2104 B.n691 B.n503 71.676
R2105 B.n687 B.n504 71.676
R2106 B.n682 B.n505 71.676
R2107 B.n678 B.n506 71.676
R2108 B.n674 B.n507 71.676
R2109 B.n670 B.n508 71.676
R2110 B.n666 B.n509 71.676
R2111 B.n661 B.n510 71.676
R2112 B.n657 B.n511 71.676
R2113 B.n653 B.n512 71.676
R2114 B.n649 B.n513 71.676
R2115 B.n645 B.n514 71.676
R2116 B.n641 B.n515 71.676
R2117 B.n637 B.n516 71.676
R2118 B.n633 B.n517 71.676
R2119 B.n629 B.n518 71.676
R2120 B.n625 B.n519 71.676
R2121 B.n621 B.n520 71.676
R2122 B.n617 B.n521 71.676
R2123 B.n613 B.n522 71.676
R2124 B.n609 B.n523 71.676
R2125 B.n605 B.n524 71.676
R2126 B.n601 B.n525 71.676
R2127 B.n597 B.n526 71.676
R2128 B.n593 B.n527 71.676
R2129 B.n589 B.n528 71.676
R2130 B.n585 B.n529 71.676
R2131 B.n581 B.n530 71.676
R2132 B.n577 B.n531 71.676
R2133 B.n573 B.n532 71.676
R2134 B.n569 B.n533 71.676
R2135 B.n565 B.n534 71.676
R2136 B.n561 B.n535 71.676
R2137 B.n557 B.n536 71.676
R2138 B.n553 B.n537 71.676
R2139 B.n549 B.n538 71.676
R2140 B.n976 B.n975 71.676
R2141 B.n146 B.n75 71.676
R2142 B.n150 B.n76 71.676
R2143 B.n154 B.n77 71.676
R2144 B.n158 B.n78 71.676
R2145 B.n162 B.n79 71.676
R2146 B.n166 B.n80 71.676
R2147 B.n170 B.n81 71.676
R2148 B.n174 B.n82 71.676
R2149 B.n178 B.n83 71.676
R2150 B.n182 B.n84 71.676
R2151 B.n186 B.n85 71.676
R2152 B.n190 B.n86 71.676
R2153 B.n194 B.n87 71.676
R2154 B.n198 B.n88 71.676
R2155 B.n202 B.n89 71.676
R2156 B.n206 B.n90 71.676
R2157 B.n210 B.n91 71.676
R2158 B.n214 B.n92 71.676
R2159 B.n218 B.n93 71.676
R2160 B.n222 B.n94 71.676
R2161 B.n226 B.n95 71.676
R2162 B.n230 B.n96 71.676
R2163 B.n234 B.n97 71.676
R2164 B.n238 B.n98 71.676
R2165 B.n242 B.n99 71.676
R2166 B.n246 B.n100 71.676
R2167 B.n250 B.n101 71.676
R2168 B.n254 B.n102 71.676
R2169 B.n258 B.n103 71.676
R2170 B.n262 B.n104 71.676
R2171 B.n266 B.n105 71.676
R2172 B.n270 B.n106 71.676
R2173 B.n274 B.n107 71.676
R2174 B.n278 B.n108 71.676
R2175 B.n282 B.n109 71.676
R2176 B.n286 B.n110 71.676
R2177 B.n290 B.n111 71.676
R2178 B.n294 B.n112 71.676
R2179 B.n298 B.n113 71.676
R2180 B.n302 B.n114 71.676
R2181 B.n306 B.n115 71.676
R2182 B.n310 B.n116 71.676
R2183 B.n314 B.n117 71.676
R2184 B.n318 B.n118 71.676
R2185 B.n322 B.n119 71.676
R2186 B.n326 B.n120 71.676
R2187 B.n330 B.n121 71.676
R2188 B.n334 B.n122 71.676
R2189 B.n338 B.n123 71.676
R2190 B.n342 B.n124 71.676
R2191 B.n346 B.n125 71.676
R2192 B.n350 B.n126 71.676
R2193 B.n354 B.n127 71.676
R2194 B.n358 B.n128 71.676
R2195 B.n362 B.n129 71.676
R2196 B.n366 B.n130 71.676
R2197 B.n370 B.n131 71.676
R2198 B.n374 B.n132 71.676
R2199 B.n378 B.n133 71.676
R2200 B.n382 B.n134 71.676
R2201 B.n386 B.n135 71.676
R2202 B.n390 B.n136 71.676
R2203 B.n394 B.n137 71.676
R2204 B.n973 B.n138 71.676
R2205 B.n973 B.n972 71.676
R2206 B.n396 B.n137 71.676
R2207 B.n393 B.n136 71.676
R2208 B.n389 B.n135 71.676
R2209 B.n385 B.n134 71.676
R2210 B.n381 B.n133 71.676
R2211 B.n377 B.n132 71.676
R2212 B.n373 B.n131 71.676
R2213 B.n369 B.n130 71.676
R2214 B.n365 B.n129 71.676
R2215 B.n361 B.n128 71.676
R2216 B.n357 B.n127 71.676
R2217 B.n353 B.n126 71.676
R2218 B.n349 B.n125 71.676
R2219 B.n345 B.n124 71.676
R2220 B.n341 B.n123 71.676
R2221 B.n337 B.n122 71.676
R2222 B.n333 B.n121 71.676
R2223 B.n329 B.n120 71.676
R2224 B.n325 B.n119 71.676
R2225 B.n321 B.n118 71.676
R2226 B.n317 B.n117 71.676
R2227 B.n313 B.n116 71.676
R2228 B.n309 B.n115 71.676
R2229 B.n305 B.n114 71.676
R2230 B.n301 B.n113 71.676
R2231 B.n297 B.n112 71.676
R2232 B.n293 B.n111 71.676
R2233 B.n289 B.n110 71.676
R2234 B.n285 B.n109 71.676
R2235 B.n281 B.n108 71.676
R2236 B.n277 B.n107 71.676
R2237 B.n273 B.n106 71.676
R2238 B.n269 B.n105 71.676
R2239 B.n265 B.n104 71.676
R2240 B.n261 B.n103 71.676
R2241 B.n257 B.n102 71.676
R2242 B.n253 B.n101 71.676
R2243 B.n249 B.n100 71.676
R2244 B.n245 B.n99 71.676
R2245 B.n241 B.n98 71.676
R2246 B.n237 B.n97 71.676
R2247 B.n233 B.n96 71.676
R2248 B.n229 B.n95 71.676
R2249 B.n225 B.n94 71.676
R2250 B.n221 B.n93 71.676
R2251 B.n217 B.n92 71.676
R2252 B.n213 B.n91 71.676
R2253 B.n209 B.n90 71.676
R2254 B.n205 B.n89 71.676
R2255 B.n201 B.n88 71.676
R2256 B.n197 B.n87 71.676
R2257 B.n193 B.n86 71.676
R2258 B.n189 B.n85 71.676
R2259 B.n185 B.n84 71.676
R2260 B.n181 B.n83 71.676
R2261 B.n177 B.n82 71.676
R2262 B.n173 B.n81 71.676
R2263 B.n169 B.n80 71.676
R2264 B.n165 B.n79 71.676
R2265 B.n161 B.n78 71.676
R2266 B.n157 B.n77 71.676
R2267 B.n153 B.n76 71.676
R2268 B.n149 B.n75 71.676
R2269 B.n975 B.n74 71.676
R2270 B.n802 B.n475 71.676
R2271 B.n796 B.n476 71.676
R2272 B.n792 B.n477 71.676
R2273 B.n788 B.n478 71.676
R2274 B.n784 B.n479 71.676
R2275 B.n780 B.n480 71.676
R2276 B.n776 B.n481 71.676
R2277 B.n772 B.n482 71.676
R2278 B.n768 B.n483 71.676
R2279 B.n764 B.n484 71.676
R2280 B.n760 B.n485 71.676
R2281 B.n756 B.n486 71.676
R2282 B.n752 B.n487 71.676
R2283 B.n748 B.n488 71.676
R2284 B.n744 B.n489 71.676
R2285 B.n740 B.n490 71.676
R2286 B.n736 B.n491 71.676
R2287 B.n732 B.n492 71.676
R2288 B.n728 B.n493 71.676
R2289 B.n724 B.n494 71.676
R2290 B.n720 B.n495 71.676
R2291 B.n716 B.n496 71.676
R2292 B.n712 B.n497 71.676
R2293 B.n708 B.n498 71.676
R2294 B.n704 B.n499 71.676
R2295 B.n700 B.n500 71.676
R2296 B.n696 B.n501 71.676
R2297 B.n692 B.n502 71.676
R2298 B.n688 B.n503 71.676
R2299 B.n683 B.n504 71.676
R2300 B.n679 B.n505 71.676
R2301 B.n675 B.n506 71.676
R2302 B.n671 B.n507 71.676
R2303 B.n667 B.n508 71.676
R2304 B.n662 B.n509 71.676
R2305 B.n658 B.n510 71.676
R2306 B.n654 B.n511 71.676
R2307 B.n650 B.n512 71.676
R2308 B.n646 B.n513 71.676
R2309 B.n642 B.n514 71.676
R2310 B.n638 B.n515 71.676
R2311 B.n634 B.n516 71.676
R2312 B.n630 B.n517 71.676
R2313 B.n626 B.n518 71.676
R2314 B.n622 B.n519 71.676
R2315 B.n618 B.n520 71.676
R2316 B.n614 B.n521 71.676
R2317 B.n610 B.n522 71.676
R2318 B.n606 B.n523 71.676
R2319 B.n602 B.n524 71.676
R2320 B.n598 B.n525 71.676
R2321 B.n594 B.n526 71.676
R2322 B.n590 B.n527 71.676
R2323 B.n586 B.n528 71.676
R2324 B.n582 B.n529 71.676
R2325 B.n578 B.n530 71.676
R2326 B.n574 B.n531 71.676
R2327 B.n570 B.n532 71.676
R2328 B.n566 B.n533 71.676
R2329 B.n562 B.n534 71.676
R2330 B.n558 B.n535 71.676
R2331 B.n554 B.n536 71.676
R2332 B.n550 B.n537 71.676
R2333 B.n546 B.n538 71.676
R2334 B.n664 B.n544 59.5399
R2335 B.n685 B.n542 59.5399
R2336 B.n145 B.n144 59.5399
R2337 B.n142 B.n141 59.5399
R2338 B.n801 B.n472 51.9027
R2339 B.n974 B.n71 51.9027
R2340 B.n544 B.n543 33.746
R2341 B.n542 B.n541 33.746
R2342 B.n144 B.n143 33.746
R2343 B.n141 B.n140 33.746
R2344 B.n808 B.n472 31.7965
R2345 B.n808 B.n468 31.7965
R2346 B.n814 B.n468 31.7965
R2347 B.n814 B.n463 31.7965
R2348 B.n820 B.n463 31.7965
R2349 B.n820 B.n464 31.7965
R2350 B.n826 B.n456 31.7965
R2351 B.n832 B.n456 31.7965
R2352 B.n832 B.n452 31.7965
R2353 B.n838 B.n452 31.7965
R2354 B.n838 B.n447 31.7965
R2355 B.n844 B.n447 31.7965
R2356 B.n844 B.n448 31.7965
R2357 B.n850 B.n440 31.7965
R2358 B.n856 B.n440 31.7965
R2359 B.n856 B.n436 31.7965
R2360 B.n862 B.n436 31.7965
R2361 B.n868 B.n432 31.7965
R2362 B.n868 B.n428 31.7965
R2363 B.n875 B.n428 31.7965
R2364 B.n875 B.n874 31.7965
R2365 B.n881 B.n421 31.7965
R2366 B.n887 B.n421 31.7965
R2367 B.n887 B.n417 31.7965
R2368 B.n893 B.n417 31.7965
R2369 B.n899 B.n413 31.7965
R2370 B.n899 B.n408 31.7965
R2371 B.n905 B.n408 31.7965
R2372 B.n905 B.n409 31.7965
R2373 B.n912 B.n401 31.7965
R2374 B.n918 B.n401 31.7965
R2375 B.n918 B.n4 31.7965
R2376 B.n1055 B.n4 31.7965
R2377 B.n1055 B.n1054 31.7965
R2378 B.n1054 B.n1053 31.7965
R2379 B.n1053 B.n8 31.7965
R2380 B.n1047 B.n8 31.7965
R2381 B.n1046 B.n1045 31.7965
R2382 B.n1045 B.n15 31.7965
R2383 B.n1039 B.n15 31.7965
R2384 B.n1039 B.n1038 31.7965
R2385 B.n1037 B.n22 31.7965
R2386 B.n1031 B.n22 31.7965
R2387 B.n1031 B.n1030 31.7965
R2388 B.n1030 B.n1029 31.7965
R2389 B.n1023 B.n32 31.7965
R2390 B.n1023 B.n1022 31.7965
R2391 B.n1022 B.n1021 31.7965
R2392 B.n1021 B.n36 31.7965
R2393 B.n1015 B.n1014 31.7965
R2394 B.n1014 B.n1013 31.7965
R2395 B.n1013 B.n43 31.7965
R2396 B.n1007 B.n43 31.7965
R2397 B.n1006 B.n1005 31.7965
R2398 B.n1005 B.n50 31.7965
R2399 B.n999 B.n50 31.7965
R2400 B.n999 B.n998 31.7965
R2401 B.n998 B.n997 31.7965
R2402 B.n997 B.n57 31.7965
R2403 B.n991 B.n57 31.7965
R2404 B.n990 B.n989 31.7965
R2405 B.n989 B.n64 31.7965
R2406 B.n983 B.n64 31.7965
R2407 B.n983 B.n982 31.7965
R2408 B.n982 B.n981 31.7965
R2409 B.n981 B.n71 31.7965
R2410 B.n826 B.t11 30.3937
R2411 B.n991 B.t15 30.3937
R2412 B.n978 B.n977 28.2542
R2413 B.n971 B.n970 28.2542
R2414 B.n545 B.n470 28.2542
R2415 B.n805 B.n804 28.2542
R2416 B.n409 B.t5 26.653
R2417 B.t2 B.n1046 26.653
R2418 B.n893 B.t8 22.9123
R2419 B.t1 B.n1037 22.9123
R2420 B.n850 B.t0 20.1068
R2421 B.n1007 B.t9 20.1068
R2422 B.n874 B.t4 19.1716
R2423 B.n32 B.t6 19.1716
R2424 B B.n1057 18.0485
R2425 B.t3 B.n432 16.3661
R2426 B.t7 B.n36 16.3661
R2427 B.n862 B.t3 15.4309
R2428 B.n1015 B.t7 15.4309
R2429 B.n881 B.t4 12.6254
R2430 B.n1029 B.t6 12.6254
R2431 B.n448 B.t0 11.6902
R2432 B.t9 B.n1006 11.6902
R2433 B.n977 B.n73 10.6151
R2434 B.n147 B.n73 10.6151
R2435 B.n148 B.n147 10.6151
R2436 B.n151 B.n148 10.6151
R2437 B.n152 B.n151 10.6151
R2438 B.n155 B.n152 10.6151
R2439 B.n156 B.n155 10.6151
R2440 B.n159 B.n156 10.6151
R2441 B.n160 B.n159 10.6151
R2442 B.n163 B.n160 10.6151
R2443 B.n164 B.n163 10.6151
R2444 B.n167 B.n164 10.6151
R2445 B.n168 B.n167 10.6151
R2446 B.n171 B.n168 10.6151
R2447 B.n172 B.n171 10.6151
R2448 B.n175 B.n172 10.6151
R2449 B.n176 B.n175 10.6151
R2450 B.n179 B.n176 10.6151
R2451 B.n180 B.n179 10.6151
R2452 B.n183 B.n180 10.6151
R2453 B.n184 B.n183 10.6151
R2454 B.n187 B.n184 10.6151
R2455 B.n188 B.n187 10.6151
R2456 B.n191 B.n188 10.6151
R2457 B.n192 B.n191 10.6151
R2458 B.n195 B.n192 10.6151
R2459 B.n196 B.n195 10.6151
R2460 B.n199 B.n196 10.6151
R2461 B.n200 B.n199 10.6151
R2462 B.n203 B.n200 10.6151
R2463 B.n204 B.n203 10.6151
R2464 B.n207 B.n204 10.6151
R2465 B.n208 B.n207 10.6151
R2466 B.n211 B.n208 10.6151
R2467 B.n212 B.n211 10.6151
R2468 B.n215 B.n212 10.6151
R2469 B.n216 B.n215 10.6151
R2470 B.n219 B.n216 10.6151
R2471 B.n220 B.n219 10.6151
R2472 B.n223 B.n220 10.6151
R2473 B.n224 B.n223 10.6151
R2474 B.n227 B.n224 10.6151
R2475 B.n228 B.n227 10.6151
R2476 B.n231 B.n228 10.6151
R2477 B.n232 B.n231 10.6151
R2478 B.n235 B.n232 10.6151
R2479 B.n236 B.n235 10.6151
R2480 B.n239 B.n236 10.6151
R2481 B.n240 B.n239 10.6151
R2482 B.n243 B.n240 10.6151
R2483 B.n244 B.n243 10.6151
R2484 B.n247 B.n244 10.6151
R2485 B.n248 B.n247 10.6151
R2486 B.n251 B.n248 10.6151
R2487 B.n252 B.n251 10.6151
R2488 B.n255 B.n252 10.6151
R2489 B.n256 B.n255 10.6151
R2490 B.n259 B.n256 10.6151
R2491 B.n260 B.n259 10.6151
R2492 B.n264 B.n263 10.6151
R2493 B.n267 B.n264 10.6151
R2494 B.n268 B.n267 10.6151
R2495 B.n271 B.n268 10.6151
R2496 B.n272 B.n271 10.6151
R2497 B.n275 B.n272 10.6151
R2498 B.n276 B.n275 10.6151
R2499 B.n279 B.n276 10.6151
R2500 B.n280 B.n279 10.6151
R2501 B.n284 B.n283 10.6151
R2502 B.n287 B.n284 10.6151
R2503 B.n288 B.n287 10.6151
R2504 B.n291 B.n288 10.6151
R2505 B.n292 B.n291 10.6151
R2506 B.n295 B.n292 10.6151
R2507 B.n296 B.n295 10.6151
R2508 B.n299 B.n296 10.6151
R2509 B.n300 B.n299 10.6151
R2510 B.n303 B.n300 10.6151
R2511 B.n304 B.n303 10.6151
R2512 B.n307 B.n304 10.6151
R2513 B.n308 B.n307 10.6151
R2514 B.n311 B.n308 10.6151
R2515 B.n312 B.n311 10.6151
R2516 B.n315 B.n312 10.6151
R2517 B.n316 B.n315 10.6151
R2518 B.n319 B.n316 10.6151
R2519 B.n320 B.n319 10.6151
R2520 B.n323 B.n320 10.6151
R2521 B.n324 B.n323 10.6151
R2522 B.n327 B.n324 10.6151
R2523 B.n328 B.n327 10.6151
R2524 B.n331 B.n328 10.6151
R2525 B.n332 B.n331 10.6151
R2526 B.n335 B.n332 10.6151
R2527 B.n336 B.n335 10.6151
R2528 B.n339 B.n336 10.6151
R2529 B.n340 B.n339 10.6151
R2530 B.n343 B.n340 10.6151
R2531 B.n344 B.n343 10.6151
R2532 B.n347 B.n344 10.6151
R2533 B.n348 B.n347 10.6151
R2534 B.n351 B.n348 10.6151
R2535 B.n352 B.n351 10.6151
R2536 B.n355 B.n352 10.6151
R2537 B.n356 B.n355 10.6151
R2538 B.n359 B.n356 10.6151
R2539 B.n360 B.n359 10.6151
R2540 B.n363 B.n360 10.6151
R2541 B.n364 B.n363 10.6151
R2542 B.n367 B.n364 10.6151
R2543 B.n368 B.n367 10.6151
R2544 B.n371 B.n368 10.6151
R2545 B.n372 B.n371 10.6151
R2546 B.n375 B.n372 10.6151
R2547 B.n376 B.n375 10.6151
R2548 B.n379 B.n376 10.6151
R2549 B.n380 B.n379 10.6151
R2550 B.n383 B.n380 10.6151
R2551 B.n384 B.n383 10.6151
R2552 B.n387 B.n384 10.6151
R2553 B.n388 B.n387 10.6151
R2554 B.n391 B.n388 10.6151
R2555 B.n392 B.n391 10.6151
R2556 B.n395 B.n392 10.6151
R2557 B.n397 B.n395 10.6151
R2558 B.n398 B.n397 10.6151
R2559 B.n971 B.n398 10.6151
R2560 B.n810 B.n470 10.6151
R2561 B.n811 B.n810 10.6151
R2562 B.n812 B.n811 10.6151
R2563 B.n812 B.n461 10.6151
R2564 B.n822 B.n461 10.6151
R2565 B.n823 B.n822 10.6151
R2566 B.n824 B.n823 10.6151
R2567 B.n824 B.n454 10.6151
R2568 B.n834 B.n454 10.6151
R2569 B.n835 B.n834 10.6151
R2570 B.n836 B.n835 10.6151
R2571 B.n836 B.n445 10.6151
R2572 B.n846 B.n445 10.6151
R2573 B.n847 B.n846 10.6151
R2574 B.n848 B.n847 10.6151
R2575 B.n848 B.n438 10.6151
R2576 B.n858 B.n438 10.6151
R2577 B.n859 B.n858 10.6151
R2578 B.n860 B.n859 10.6151
R2579 B.n860 B.n430 10.6151
R2580 B.n870 B.n430 10.6151
R2581 B.n871 B.n870 10.6151
R2582 B.n872 B.n871 10.6151
R2583 B.n872 B.n423 10.6151
R2584 B.n883 B.n423 10.6151
R2585 B.n884 B.n883 10.6151
R2586 B.n885 B.n884 10.6151
R2587 B.n885 B.n415 10.6151
R2588 B.n895 B.n415 10.6151
R2589 B.n896 B.n895 10.6151
R2590 B.n897 B.n896 10.6151
R2591 B.n897 B.n406 10.6151
R2592 B.n907 B.n406 10.6151
R2593 B.n908 B.n907 10.6151
R2594 B.n910 B.n908 10.6151
R2595 B.n910 B.n909 10.6151
R2596 B.n909 B.n399 10.6151
R2597 B.n921 B.n399 10.6151
R2598 B.n922 B.n921 10.6151
R2599 B.n923 B.n922 10.6151
R2600 B.n924 B.n923 10.6151
R2601 B.n926 B.n924 10.6151
R2602 B.n927 B.n926 10.6151
R2603 B.n928 B.n927 10.6151
R2604 B.n929 B.n928 10.6151
R2605 B.n931 B.n929 10.6151
R2606 B.n932 B.n931 10.6151
R2607 B.n933 B.n932 10.6151
R2608 B.n934 B.n933 10.6151
R2609 B.n936 B.n934 10.6151
R2610 B.n937 B.n936 10.6151
R2611 B.n938 B.n937 10.6151
R2612 B.n939 B.n938 10.6151
R2613 B.n941 B.n939 10.6151
R2614 B.n942 B.n941 10.6151
R2615 B.n943 B.n942 10.6151
R2616 B.n944 B.n943 10.6151
R2617 B.n946 B.n944 10.6151
R2618 B.n947 B.n946 10.6151
R2619 B.n948 B.n947 10.6151
R2620 B.n949 B.n948 10.6151
R2621 B.n951 B.n949 10.6151
R2622 B.n952 B.n951 10.6151
R2623 B.n953 B.n952 10.6151
R2624 B.n954 B.n953 10.6151
R2625 B.n956 B.n954 10.6151
R2626 B.n957 B.n956 10.6151
R2627 B.n958 B.n957 10.6151
R2628 B.n959 B.n958 10.6151
R2629 B.n961 B.n959 10.6151
R2630 B.n962 B.n961 10.6151
R2631 B.n963 B.n962 10.6151
R2632 B.n964 B.n963 10.6151
R2633 B.n966 B.n964 10.6151
R2634 B.n967 B.n966 10.6151
R2635 B.n968 B.n967 10.6151
R2636 B.n969 B.n968 10.6151
R2637 B.n970 B.n969 10.6151
R2638 B.n804 B.n474 10.6151
R2639 B.n799 B.n474 10.6151
R2640 B.n799 B.n798 10.6151
R2641 B.n798 B.n797 10.6151
R2642 B.n797 B.n794 10.6151
R2643 B.n794 B.n793 10.6151
R2644 B.n793 B.n790 10.6151
R2645 B.n790 B.n789 10.6151
R2646 B.n789 B.n786 10.6151
R2647 B.n786 B.n785 10.6151
R2648 B.n785 B.n782 10.6151
R2649 B.n782 B.n781 10.6151
R2650 B.n781 B.n778 10.6151
R2651 B.n778 B.n777 10.6151
R2652 B.n777 B.n774 10.6151
R2653 B.n774 B.n773 10.6151
R2654 B.n773 B.n770 10.6151
R2655 B.n770 B.n769 10.6151
R2656 B.n769 B.n766 10.6151
R2657 B.n766 B.n765 10.6151
R2658 B.n765 B.n762 10.6151
R2659 B.n762 B.n761 10.6151
R2660 B.n761 B.n758 10.6151
R2661 B.n758 B.n757 10.6151
R2662 B.n757 B.n754 10.6151
R2663 B.n754 B.n753 10.6151
R2664 B.n753 B.n750 10.6151
R2665 B.n750 B.n749 10.6151
R2666 B.n749 B.n746 10.6151
R2667 B.n746 B.n745 10.6151
R2668 B.n745 B.n742 10.6151
R2669 B.n742 B.n741 10.6151
R2670 B.n741 B.n738 10.6151
R2671 B.n738 B.n737 10.6151
R2672 B.n737 B.n734 10.6151
R2673 B.n734 B.n733 10.6151
R2674 B.n733 B.n730 10.6151
R2675 B.n730 B.n729 10.6151
R2676 B.n729 B.n726 10.6151
R2677 B.n726 B.n725 10.6151
R2678 B.n725 B.n722 10.6151
R2679 B.n722 B.n721 10.6151
R2680 B.n721 B.n718 10.6151
R2681 B.n718 B.n717 10.6151
R2682 B.n717 B.n714 10.6151
R2683 B.n714 B.n713 10.6151
R2684 B.n713 B.n710 10.6151
R2685 B.n710 B.n709 10.6151
R2686 B.n709 B.n706 10.6151
R2687 B.n706 B.n705 10.6151
R2688 B.n705 B.n702 10.6151
R2689 B.n702 B.n701 10.6151
R2690 B.n701 B.n698 10.6151
R2691 B.n698 B.n697 10.6151
R2692 B.n697 B.n694 10.6151
R2693 B.n694 B.n693 10.6151
R2694 B.n693 B.n690 10.6151
R2695 B.n690 B.n689 10.6151
R2696 B.n689 B.n686 10.6151
R2697 B.n684 B.n681 10.6151
R2698 B.n681 B.n680 10.6151
R2699 B.n680 B.n677 10.6151
R2700 B.n677 B.n676 10.6151
R2701 B.n676 B.n673 10.6151
R2702 B.n673 B.n672 10.6151
R2703 B.n672 B.n669 10.6151
R2704 B.n669 B.n668 10.6151
R2705 B.n668 B.n665 10.6151
R2706 B.n663 B.n660 10.6151
R2707 B.n660 B.n659 10.6151
R2708 B.n659 B.n656 10.6151
R2709 B.n656 B.n655 10.6151
R2710 B.n655 B.n652 10.6151
R2711 B.n652 B.n651 10.6151
R2712 B.n651 B.n648 10.6151
R2713 B.n648 B.n647 10.6151
R2714 B.n647 B.n644 10.6151
R2715 B.n644 B.n643 10.6151
R2716 B.n643 B.n640 10.6151
R2717 B.n640 B.n639 10.6151
R2718 B.n639 B.n636 10.6151
R2719 B.n636 B.n635 10.6151
R2720 B.n635 B.n632 10.6151
R2721 B.n632 B.n631 10.6151
R2722 B.n631 B.n628 10.6151
R2723 B.n628 B.n627 10.6151
R2724 B.n627 B.n624 10.6151
R2725 B.n624 B.n623 10.6151
R2726 B.n623 B.n620 10.6151
R2727 B.n620 B.n619 10.6151
R2728 B.n619 B.n616 10.6151
R2729 B.n616 B.n615 10.6151
R2730 B.n615 B.n612 10.6151
R2731 B.n612 B.n611 10.6151
R2732 B.n611 B.n608 10.6151
R2733 B.n608 B.n607 10.6151
R2734 B.n607 B.n604 10.6151
R2735 B.n604 B.n603 10.6151
R2736 B.n603 B.n600 10.6151
R2737 B.n600 B.n599 10.6151
R2738 B.n599 B.n596 10.6151
R2739 B.n596 B.n595 10.6151
R2740 B.n595 B.n592 10.6151
R2741 B.n592 B.n591 10.6151
R2742 B.n591 B.n588 10.6151
R2743 B.n588 B.n587 10.6151
R2744 B.n587 B.n584 10.6151
R2745 B.n584 B.n583 10.6151
R2746 B.n583 B.n580 10.6151
R2747 B.n580 B.n579 10.6151
R2748 B.n579 B.n576 10.6151
R2749 B.n576 B.n575 10.6151
R2750 B.n575 B.n572 10.6151
R2751 B.n572 B.n571 10.6151
R2752 B.n571 B.n568 10.6151
R2753 B.n568 B.n567 10.6151
R2754 B.n567 B.n564 10.6151
R2755 B.n564 B.n563 10.6151
R2756 B.n563 B.n560 10.6151
R2757 B.n560 B.n559 10.6151
R2758 B.n559 B.n556 10.6151
R2759 B.n556 B.n555 10.6151
R2760 B.n555 B.n552 10.6151
R2761 B.n552 B.n551 10.6151
R2762 B.n551 B.n548 10.6151
R2763 B.n548 B.n547 10.6151
R2764 B.n547 B.n545 10.6151
R2765 B.n806 B.n805 10.6151
R2766 B.n806 B.n466 10.6151
R2767 B.n816 B.n466 10.6151
R2768 B.n817 B.n816 10.6151
R2769 B.n818 B.n817 10.6151
R2770 B.n818 B.n458 10.6151
R2771 B.n828 B.n458 10.6151
R2772 B.n829 B.n828 10.6151
R2773 B.n830 B.n829 10.6151
R2774 B.n830 B.n450 10.6151
R2775 B.n840 B.n450 10.6151
R2776 B.n841 B.n840 10.6151
R2777 B.n842 B.n841 10.6151
R2778 B.n842 B.n442 10.6151
R2779 B.n852 B.n442 10.6151
R2780 B.n853 B.n852 10.6151
R2781 B.n854 B.n853 10.6151
R2782 B.n854 B.n434 10.6151
R2783 B.n864 B.n434 10.6151
R2784 B.n865 B.n864 10.6151
R2785 B.n866 B.n865 10.6151
R2786 B.n866 B.n426 10.6151
R2787 B.n877 B.n426 10.6151
R2788 B.n878 B.n877 10.6151
R2789 B.n879 B.n878 10.6151
R2790 B.n879 B.n419 10.6151
R2791 B.n889 B.n419 10.6151
R2792 B.n890 B.n889 10.6151
R2793 B.n891 B.n890 10.6151
R2794 B.n891 B.n411 10.6151
R2795 B.n901 B.n411 10.6151
R2796 B.n902 B.n901 10.6151
R2797 B.n903 B.n902 10.6151
R2798 B.n903 B.n403 10.6151
R2799 B.n914 B.n403 10.6151
R2800 B.n915 B.n914 10.6151
R2801 B.n916 B.n915 10.6151
R2802 B.n916 B.n0 10.6151
R2803 B.n1051 B.n1 10.6151
R2804 B.n1051 B.n1050 10.6151
R2805 B.n1050 B.n1049 10.6151
R2806 B.n1049 B.n10 10.6151
R2807 B.n1043 B.n10 10.6151
R2808 B.n1043 B.n1042 10.6151
R2809 B.n1042 B.n1041 10.6151
R2810 B.n1041 B.n17 10.6151
R2811 B.n1035 B.n17 10.6151
R2812 B.n1035 B.n1034 10.6151
R2813 B.n1034 B.n1033 10.6151
R2814 B.n1033 B.n24 10.6151
R2815 B.n1027 B.n24 10.6151
R2816 B.n1027 B.n1026 10.6151
R2817 B.n1026 B.n1025 10.6151
R2818 B.n1025 B.n30 10.6151
R2819 B.n1019 B.n30 10.6151
R2820 B.n1019 B.n1018 10.6151
R2821 B.n1018 B.n1017 10.6151
R2822 B.n1017 B.n38 10.6151
R2823 B.n1011 B.n38 10.6151
R2824 B.n1011 B.n1010 10.6151
R2825 B.n1010 B.n1009 10.6151
R2826 B.n1009 B.n45 10.6151
R2827 B.n1003 B.n45 10.6151
R2828 B.n1003 B.n1002 10.6151
R2829 B.n1002 B.n1001 10.6151
R2830 B.n1001 B.n52 10.6151
R2831 B.n995 B.n52 10.6151
R2832 B.n995 B.n994 10.6151
R2833 B.n994 B.n993 10.6151
R2834 B.n993 B.n59 10.6151
R2835 B.n987 B.n59 10.6151
R2836 B.n987 B.n986 10.6151
R2837 B.n986 B.n985 10.6151
R2838 B.n985 B.n66 10.6151
R2839 B.n979 B.n66 10.6151
R2840 B.n979 B.n978 10.6151
R2841 B.n260 B.n145 9.36635
R2842 B.n283 B.n142 9.36635
R2843 B.n686 B.n685 9.36635
R2844 B.n664 B.n663 9.36635
R2845 B.t8 B.n413 8.88467
R2846 B.n1038 B.t1 8.88467
R2847 B.n912 B.t5 5.14396
R2848 B.n1047 B.t2 5.14396
R2849 B.n1057 B.n0 2.81026
R2850 B.n1057 B.n1 2.81026
R2851 B.n464 B.t11 1.40326
R2852 B.t15 B.n990 1.40326
R2853 B.n263 B.n145 1.24928
R2854 B.n280 B.n142 1.24928
R2855 B.n685 B.n684 1.24928
R2856 B.n665 B.n664 1.24928
R2857 VN.n6 VN.t4 346.658
R2858 VN.n33 VN.t7 346.658
R2859 VN.n5 VN.t6 311.933
R2860 VN.n10 VN.t2 311.933
R2861 VN.n17 VN.t3 311.933
R2862 VN.n24 VN.t8 311.933
R2863 VN.n32 VN.t0 311.933
R2864 VN.n31 VN.t9 311.933
R2865 VN.n43 VN.t5 311.933
R2866 VN.n50 VN.t1 311.933
R2867 VN.n25 VN.n24 174.512
R2868 VN.n51 VN.n50 174.512
R2869 VN.n49 VN.n26 161.3
R2870 VN.n48 VN.n47 161.3
R2871 VN.n46 VN.n27 161.3
R2872 VN.n45 VN.n44 161.3
R2873 VN.n42 VN.n28 161.3
R2874 VN.n41 VN.n40 161.3
R2875 VN.n39 VN.n29 161.3
R2876 VN.n38 VN.n37 161.3
R2877 VN.n36 VN.n30 161.3
R2878 VN.n35 VN.n34 161.3
R2879 VN.n23 VN.n0 161.3
R2880 VN.n22 VN.n21 161.3
R2881 VN.n20 VN.n1 161.3
R2882 VN.n19 VN.n18 161.3
R2883 VN.n16 VN.n2 161.3
R2884 VN.n15 VN.n14 161.3
R2885 VN.n13 VN.n3 161.3
R2886 VN.n12 VN.n11 161.3
R2887 VN.n9 VN.n4 161.3
R2888 VN.n8 VN.n7 161.3
R2889 VN.n22 VN.n1 54.0911
R2890 VN.n48 VN.n27 54.0911
R2891 VN.n9 VN.n8 52.1486
R2892 VN.n16 VN.n15 52.1486
R2893 VN.n36 VN.n35 52.1486
R2894 VN.n42 VN.n41 52.1486
R2895 VN VN.n51 51.6842
R2896 VN.n6 VN.n5 42.3338
R2897 VN.n33 VN.n32 42.3338
R2898 VN.n11 VN.n9 28.8382
R2899 VN.n15 VN.n3 28.8382
R2900 VN.n37 VN.n36 28.8382
R2901 VN.n41 VN.n29 28.8382
R2902 VN.n23 VN.n22 26.8957
R2903 VN.n49 VN.n48 26.8957
R2904 VN.n18 VN.n1 24.4675
R2905 VN.n44 VN.n27 24.4675
R2906 VN.n8 VN.n5 23.9782
R2907 VN.n17 VN.n16 23.9782
R2908 VN.n35 VN.n32 23.9782
R2909 VN.n43 VN.n42 23.9782
R2910 VN.n34 VN.n33 17.64
R2911 VN.n7 VN.n6 17.64
R2912 VN.n11 VN.n10 12.234
R2913 VN.n10 VN.n3 12.234
R2914 VN.n31 VN.n29 12.234
R2915 VN.n37 VN.n31 12.234
R2916 VN.n24 VN.n23 11.2553
R2917 VN.n50 VN.n49 11.2553
R2918 VN.n18 VN.n17 0.48984
R2919 VN.n44 VN.n43 0.48984
R2920 VN.n51 VN.n26 0.189894
R2921 VN.n47 VN.n26 0.189894
R2922 VN.n47 VN.n46 0.189894
R2923 VN.n46 VN.n45 0.189894
R2924 VN.n45 VN.n28 0.189894
R2925 VN.n40 VN.n28 0.189894
R2926 VN.n40 VN.n39 0.189894
R2927 VN.n39 VN.n38 0.189894
R2928 VN.n38 VN.n30 0.189894
R2929 VN.n34 VN.n30 0.189894
R2930 VN.n7 VN.n4 0.189894
R2931 VN.n12 VN.n4 0.189894
R2932 VN.n13 VN.n12 0.189894
R2933 VN.n14 VN.n13 0.189894
R2934 VN.n14 VN.n2 0.189894
R2935 VN.n19 VN.n2 0.189894
R2936 VN.n20 VN.n19 0.189894
R2937 VN.n21 VN.n20 0.189894
R2938 VN.n21 VN.n0 0.189894
R2939 VN.n25 VN.n0 0.189894
R2940 VN VN.n25 0.0516364
R2941 VDD2.n201 VDD2.n105 289.615
R2942 VDD2.n96 VDD2.n0 289.615
R2943 VDD2.n202 VDD2.n201 185
R2944 VDD2.n200 VDD2.n199 185
R2945 VDD2.n109 VDD2.n108 185
R2946 VDD2.n194 VDD2.n193 185
R2947 VDD2.n192 VDD2.n191 185
R2948 VDD2.n113 VDD2.n112 185
R2949 VDD2.n186 VDD2.n185 185
R2950 VDD2.n184 VDD2.n115 185
R2951 VDD2.n183 VDD2.n182 185
R2952 VDD2.n118 VDD2.n116 185
R2953 VDD2.n177 VDD2.n176 185
R2954 VDD2.n175 VDD2.n174 185
R2955 VDD2.n122 VDD2.n121 185
R2956 VDD2.n169 VDD2.n168 185
R2957 VDD2.n167 VDD2.n166 185
R2958 VDD2.n126 VDD2.n125 185
R2959 VDD2.n161 VDD2.n160 185
R2960 VDD2.n159 VDD2.n158 185
R2961 VDD2.n130 VDD2.n129 185
R2962 VDD2.n153 VDD2.n152 185
R2963 VDD2.n151 VDD2.n150 185
R2964 VDD2.n134 VDD2.n133 185
R2965 VDD2.n145 VDD2.n144 185
R2966 VDD2.n143 VDD2.n142 185
R2967 VDD2.n138 VDD2.n137 185
R2968 VDD2.n32 VDD2.n31 185
R2969 VDD2.n37 VDD2.n36 185
R2970 VDD2.n39 VDD2.n38 185
R2971 VDD2.n28 VDD2.n27 185
R2972 VDD2.n45 VDD2.n44 185
R2973 VDD2.n47 VDD2.n46 185
R2974 VDD2.n24 VDD2.n23 185
R2975 VDD2.n53 VDD2.n52 185
R2976 VDD2.n55 VDD2.n54 185
R2977 VDD2.n20 VDD2.n19 185
R2978 VDD2.n61 VDD2.n60 185
R2979 VDD2.n63 VDD2.n62 185
R2980 VDD2.n16 VDD2.n15 185
R2981 VDD2.n69 VDD2.n68 185
R2982 VDD2.n71 VDD2.n70 185
R2983 VDD2.n12 VDD2.n11 185
R2984 VDD2.n78 VDD2.n77 185
R2985 VDD2.n79 VDD2.n10 185
R2986 VDD2.n81 VDD2.n80 185
R2987 VDD2.n8 VDD2.n7 185
R2988 VDD2.n87 VDD2.n86 185
R2989 VDD2.n89 VDD2.n88 185
R2990 VDD2.n4 VDD2.n3 185
R2991 VDD2.n95 VDD2.n94 185
R2992 VDD2.n97 VDD2.n96 185
R2993 VDD2.n139 VDD2.t8 147.659
R2994 VDD2.n33 VDD2.t5 147.659
R2995 VDD2.n201 VDD2.n200 104.615
R2996 VDD2.n200 VDD2.n108 104.615
R2997 VDD2.n193 VDD2.n108 104.615
R2998 VDD2.n193 VDD2.n192 104.615
R2999 VDD2.n192 VDD2.n112 104.615
R3000 VDD2.n185 VDD2.n112 104.615
R3001 VDD2.n185 VDD2.n184 104.615
R3002 VDD2.n184 VDD2.n183 104.615
R3003 VDD2.n183 VDD2.n116 104.615
R3004 VDD2.n176 VDD2.n116 104.615
R3005 VDD2.n176 VDD2.n175 104.615
R3006 VDD2.n175 VDD2.n121 104.615
R3007 VDD2.n168 VDD2.n121 104.615
R3008 VDD2.n168 VDD2.n167 104.615
R3009 VDD2.n167 VDD2.n125 104.615
R3010 VDD2.n160 VDD2.n125 104.615
R3011 VDD2.n160 VDD2.n159 104.615
R3012 VDD2.n159 VDD2.n129 104.615
R3013 VDD2.n152 VDD2.n129 104.615
R3014 VDD2.n152 VDD2.n151 104.615
R3015 VDD2.n151 VDD2.n133 104.615
R3016 VDD2.n144 VDD2.n133 104.615
R3017 VDD2.n144 VDD2.n143 104.615
R3018 VDD2.n143 VDD2.n137 104.615
R3019 VDD2.n37 VDD2.n31 104.615
R3020 VDD2.n38 VDD2.n37 104.615
R3021 VDD2.n38 VDD2.n27 104.615
R3022 VDD2.n45 VDD2.n27 104.615
R3023 VDD2.n46 VDD2.n45 104.615
R3024 VDD2.n46 VDD2.n23 104.615
R3025 VDD2.n53 VDD2.n23 104.615
R3026 VDD2.n54 VDD2.n53 104.615
R3027 VDD2.n54 VDD2.n19 104.615
R3028 VDD2.n61 VDD2.n19 104.615
R3029 VDD2.n62 VDD2.n61 104.615
R3030 VDD2.n62 VDD2.n15 104.615
R3031 VDD2.n69 VDD2.n15 104.615
R3032 VDD2.n70 VDD2.n69 104.615
R3033 VDD2.n70 VDD2.n11 104.615
R3034 VDD2.n78 VDD2.n11 104.615
R3035 VDD2.n79 VDD2.n78 104.615
R3036 VDD2.n80 VDD2.n79 104.615
R3037 VDD2.n80 VDD2.n7 104.615
R3038 VDD2.n87 VDD2.n7 104.615
R3039 VDD2.n88 VDD2.n87 104.615
R3040 VDD2.n88 VDD2.n3 104.615
R3041 VDD2.n95 VDD2.n3 104.615
R3042 VDD2.n96 VDD2.n95 104.615
R3043 VDD2.n104 VDD2.n103 61.9117
R3044 VDD2 VDD2.n209 61.9089
R3045 VDD2.n208 VDD2.n207 60.8422
R3046 VDD2.n102 VDD2.n101 60.842
R3047 VDD2.t8 VDD2.n137 52.3082
R3048 VDD2.t5 VDD2.n31 52.3082
R3049 VDD2.n102 VDD2.n100 50.5581
R3050 VDD2.n206 VDD2.n205 49.0581
R3051 VDD2.n206 VDD2.n104 46.5731
R3052 VDD2.n139 VDD2.n138 15.6677
R3053 VDD2.n33 VDD2.n32 15.6677
R3054 VDD2.n186 VDD2.n115 13.1884
R3055 VDD2.n81 VDD2.n10 13.1884
R3056 VDD2.n187 VDD2.n113 12.8005
R3057 VDD2.n182 VDD2.n117 12.8005
R3058 VDD2.n142 VDD2.n141 12.8005
R3059 VDD2.n36 VDD2.n35 12.8005
R3060 VDD2.n77 VDD2.n76 12.8005
R3061 VDD2.n82 VDD2.n8 12.8005
R3062 VDD2.n191 VDD2.n190 12.0247
R3063 VDD2.n181 VDD2.n118 12.0247
R3064 VDD2.n145 VDD2.n136 12.0247
R3065 VDD2.n39 VDD2.n30 12.0247
R3066 VDD2.n75 VDD2.n12 12.0247
R3067 VDD2.n86 VDD2.n85 12.0247
R3068 VDD2.n194 VDD2.n111 11.249
R3069 VDD2.n178 VDD2.n177 11.249
R3070 VDD2.n146 VDD2.n134 11.249
R3071 VDD2.n40 VDD2.n28 11.249
R3072 VDD2.n72 VDD2.n71 11.249
R3073 VDD2.n89 VDD2.n6 11.249
R3074 VDD2.n195 VDD2.n109 10.4732
R3075 VDD2.n174 VDD2.n120 10.4732
R3076 VDD2.n150 VDD2.n149 10.4732
R3077 VDD2.n44 VDD2.n43 10.4732
R3078 VDD2.n68 VDD2.n14 10.4732
R3079 VDD2.n90 VDD2.n4 10.4732
R3080 VDD2.n199 VDD2.n198 9.69747
R3081 VDD2.n173 VDD2.n122 9.69747
R3082 VDD2.n153 VDD2.n132 9.69747
R3083 VDD2.n47 VDD2.n26 9.69747
R3084 VDD2.n67 VDD2.n16 9.69747
R3085 VDD2.n94 VDD2.n93 9.69747
R3086 VDD2.n205 VDD2.n204 9.45567
R3087 VDD2.n100 VDD2.n99 9.45567
R3088 VDD2.n165 VDD2.n164 9.3005
R3089 VDD2.n124 VDD2.n123 9.3005
R3090 VDD2.n171 VDD2.n170 9.3005
R3091 VDD2.n173 VDD2.n172 9.3005
R3092 VDD2.n120 VDD2.n119 9.3005
R3093 VDD2.n179 VDD2.n178 9.3005
R3094 VDD2.n181 VDD2.n180 9.3005
R3095 VDD2.n117 VDD2.n114 9.3005
R3096 VDD2.n204 VDD2.n203 9.3005
R3097 VDD2.n107 VDD2.n106 9.3005
R3098 VDD2.n198 VDD2.n197 9.3005
R3099 VDD2.n196 VDD2.n195 9.3005
R3100 VDD2.n111 VDD2.n110 9.3005
R3101 VDD2.n190 VDD2.n189 9.3005
R3102 VDD2.n188 VDD2.n187 9.3005
R3103 VDD2.n163 VDD2.n162 9.3005
R3104 VDD2.n128 VDD2.n127 9.3005
R3105 VDD2.n157 VDD2.n156 9.3005
R3106 VDD2.n155 VDD2.n154 9.3005
R3107 VDD2.n132 VDD2.n131 9.3005
R3108 VDD2.n149 VDD2.n148 9.3005
R3109 VDD2.n147 VDD2.n146 9.3005
R3110 VDD2.n136 VDD2.n135 9.3005
R3111 VDD2.n141 VDD2.n140 9.3005
R3112 VDD2.n99 VDD2.n98 9.3005
R3113 VDD2.n2 VDD2.n1 9.3005
R3114 VDD2.n93 VDD2.n92 9.3005
R3115 VDD2.n91 VDD2.n90 9.3005
R3116 VDD2.n6 VDD2.n5 9.3005
R3117 VDD2.n85 VDD2.n84 9.3005
R3118 VDD2.n83 VDD2.n82 9.3005
R3119 VDD2.n22 VDD2.n21 9.3005
R3120 VDD2.n51 VDD2.n50 9.3005
R3121 VDD2.n49 VDD2.n48 9.3005
R3122 VDD2.n26 VDD2.n25 9.3005
R3123 VDD2.n43 VDD2.n42 9.3005
R3124 VDD2.n41 VDD2.n40 9.3005
R3125 VDD2.n30 VDD2.n29 9.3005
R3126 VDD2.n35 VDD2.n34 9.3005
R3127 VDD2.n57 VDD2.n56 9.3005
R3128 VDD2.n59 VDD2.n58 9.3005
R3129 VDD2.n18 VDD2.n17 9.3005
R3130 VDD2.n65 VDD2.n64 9.3005
R3131 VDD2.n67 VDD2.n66 9.3005
R3132 VDD2.n14 VDD2.n13 9.3005
R3133 VDD2.n73 VDD2.n72 9.3005
R3134 VDD2.n75 VDD2.n74 9.3005
R3135 VDD2.n76 VDD2.n9 9.3005
R3136 VDD2.n202 VDD2.n107 8.92171
R3137 VDD2.n170 VDD2.n169 8.92171
R3138 VDD2.n154 VDD2.n130 8.92171
R3139 VDD2.n48 VDD2.n24 8.92171
R3140 VDD2.n64 VDD2.n63 8.92171
R3141 VDD2.n97 VDD2.n2 8.92171
R3142 VDD2.n203 VDD2.n105 8.14595
R3143 VDD2.n166 VDD2.n124 8.14595
R3144 VDD2.n158 VDD2.n157 8.14595
R3145 VDD2.n52 VDD2.n51 8.14595
R3146 VDD2.n60 VDD2.n18 8.14595
R3147 VDD2.n98 VDD2.n0 8.14595
R3148 VDD2.n165 VDD2.n126 7.3702
R3149 VDD2.n161 VDD2.n128 7.3702
R3150 VDD2.n55 VDD2.n22 7.3702
R3151 VDD2.n59 VDD2.n20 7.3702
R3152 VDD2.n162 VDD2.n126 6.59444
R3153 VDD2.n162 VDD2.n161 6.59444
R3154 VDD2.n56 VDD2.n55 6.59444
R3155 VDD2.n56 VDD2.n20 6.59444
R3156 VDD2.n205 VDD2.n105 5.81868
R3157 VDD2.n166 VDD2.n165 5.81868
R3158 VDD2.n158 VDD2.n128 5.81868
R3159 VDD2.n52 VDD2.n22 5.81868
R3160 VDD2.n60 VDD2.n59 5.81868
R3161 VDD2.n100 VDD2.n0 5.81868
R3162 VDD2.n203 VDD2.n202 5.04292
R3163 VDD2.n169 VDD2.n124 5.04292
R3164 VDD2.n157 VDD2.n130 5.04292
R3165 VDD2.n51 VDD2.n24 5.04292
R3166 VDD2.n63 VDD2.n18 5.04292
R3167 VDD2.n98 VDD2.n97 5.04292
R3168 VDD2.n140 VDD2.n139 4.38563
R3169 VDD2.n34 VDD2.n33 4.38563
R3170 VDD2.n199 VDD2.n107 4.26717
R3171 VDD2.n170 VDD2.n122 4.26717
R3172 VDD2.n154 VDD2.n153 4.26717
R3173 VDD2.n48 VDD2.n47 4.26717
R3174 VDD2.n64 VDD2.n16 4.26717
R3175 VDD2.n94 VDD2.n2 4.26717
R3176 VDD2.n198 VDD2.n109 3.49141
R3177 VDD2.n174 VDD2.n173 3.49141
R3178 VDD2.n150 VDD2.n132 3.49141
R3179 VDD2.n44 VDD2.n26 3.49141
R3180 VDD2.n68 VDD2.n67 3.49141
R3181 VDD2.n93 VDD2.n4 3.49141
R3182 VDD2.n195 VDD2.n194 2.71565
R3183 VDD2.n177 VDD2.n120 2.71565
R3184 VDD2.n149 VDD2.n134 2.71565
R3185 VDD2.n43 VDD2.n28 2.71565
R3186 VDD2.n71 VDD2.n14 2.71565
R3187 VDD2.n90 VDD2.n89 2.71565
R3188 VDD2.n191 VDD2.n111 1.93989
R3189 VDD2.n178 VDD2.n118 1.93989
R3190 VDD2.n146 VDD2.n145 1.93989
R3191 VDD2.n40 VDD2.n39 1.93989
R3192 VDD2.n72 VDD2.n12 1.93989
R3193 VDD2.n86 VDD2.n6 1.93989
R3194 VDD2.n208 VDD2.n206 1.5005
R3195 VDD2.n190 VDD2.n113 1.16414
R3196 VDD2.n182 VDD2.n181 1.16414
R3197 VDD2.n142 VDD2.n136 1.16414
R3198 VDD2.n36 VDD2.n30 1.16414
R3199 VDD2.n77 VDD2.n75 1.16414
R3200 VDD2.n85 VDD2.n8 1.16414
R3201 VDD2.n209 VDD2.t9 1.08543
R3202 VDD2.n209 VDD2.t2 1.08543
R3203 VDD2.n207 VDD2.t4 1.08543
R3204 VDD2.n207 VDD2.t0 1.08543
R3205 VDD2.n103 VDD2.t6 1.08543
R3206 VDD2.n103 VDD2.t1 1.08543
R3207 VDD2.n101 VDD2.t3 1.08543
R3208 VDD2.n101 VDD2.t7 1.08543
R3209 VDD2 VDD2.n208 0.43369
R3210 VDD2.n187 VDD2.n186 0.388379
R3211 VDD2.n117 VDD2.n115 0.388379
R3212 VDD2.n141 VDD2.n138 0.388379
R3213 VDD2.n35 VDD2.n32 0.388379
R3214 VDD2.n76 VDD2.n10 0.388379
R3215 VDD2.n82 VDD2.n81 0.388379
R3216 VDD2.n104 VDD2.n102 0.320154
R3217 VDD2.n204 VDD2.n106 0.155672
R3218 VDD2.n197 VDD2.n106 0.155672
R3219 VDD2.n197 VDD2.n196 0.155672
R3220 VDD2.n196 VDD2.n110 0.155672
R3221 VDD2.n189 VDD2.n110 0.155672
R3222 VDD2.n189 VDD2.n188 0.155672
R3223 VDD2.n188 VDD2.n114 0.155672
R3224 VDD2.n180 VDD2.n114 0.155672
R3225 VDD2.n180 VDD2.n179 0.155672
R3226 VDD2.n179 VDD2.n119 0.155672
R3227 VDD2.n172 VDD2.n119 0.155672
R3228 VDD2.n172 VDD2.n171 0.155672
R3229 VDD2.n171 VDD2.n123 0.155672
R3230 VDD2.n164 VDD2.n123 0.155672
R3231 VDD2.n164 VDD2.n163 0.155672
R3232 VDD2.n163 VDD2.n127 0.155672
R3233 VDD2.n156 VDD2.n127 0.155672
R3234 VDD2.n156 VDD2.n155 0.155672
R3235 VDD2.n155 VDD2.n131 0.155672
R3236 VDD2.n148 VDD2.n131 0.155672
R3237 VDD2.n148 VDD2.n147 0.155672
R3238 VDD2.n147 VDD2.n135 0.155672
R3239 VDD2.n140 VDD2.n135 0.155672
R3240 VDD2.n34 VDD2.n29 0.155672
R3241 VDD2.n41 VDD2.n29 0.155672
R3242 VDD2.n42 VDD2.n41 0.155672
R3243 VDD2.n42 VDD2.n25 0.155672
R3244 VDD2.n49 VDD2.n25 0.155672
R3245 VDD2.n50 VDD2.n49 0.155672
R3246 VDD2.n50 VDD2.n21 0.155672
R3247 VDD2.n57 VDD2.n21 0.155672
R3248 VDD2.n58 VDD2.n57 0.155672
R3249 VDD2.n58 VDD2.n17 0.155672
R3250 VDD2.n65 VDD2.n17 0.155672
R3251 VDD2.n66 VDD2.n65 0.155672
R3252 VDD2.n66 VDD2.n13 0.155672
R3253 VDD2.n73 VDD2.n13 0.155672
R3254 VDD2.n74 VDD2.n73 0.155672
R3255 VDD2.n74 VDD2.n9 0.155672
R3256 VDD2.n83 VDD2.n9 0.155672
R3257 VDD2.n84 VDD2.n83 0.155672
R3258 VDD2.n84 VDD2.n5 0.155672
R3259 VDD2.n91 VDD2.n5 0.155672
R3260 VDD2.n92 VDD2.n91 0.155672
R3261 VDD2.n92 VDD2.n1 0.155672
R3262 VDD2.n99 VDD2.n1 0.155672
C0 VP VTAIL 13.458401f
C1 VDD1 VDD2 1.40204f
C2 VDD1 VP 13.8229f
C3 VN VTAIL 13.443799f
C4 VDD2 VP 0.432634f
C5 VDD1 VN 0.150637f
C6 VDD1 VTAIL 15.0946f
C7 VDD2 VN 13.546599f
C8 VP VN 7.80184f
C9 VDD2 VTAIL 15.133299f
C10 VDD2 B 6.929022f
C11 VDD1 B 6.897244f
C12 VTAIL B 9.60502f
C13 VN B 13.20382f
C14 VP B 11.34165f
C15 VDD2.n0 B 0.031627f
C16 VDD2.n1 B 0.022393f
C17 VDD2.n2 B 0.012033f
C18 VDD2.n3 B 0.028442f
C19 VDD2.n4 B 0.012741f
C20 VDD2.n5 B 0.022393f
C21 VDD2.n6 B 0.012033f
C22 VDD2.n7 B 0.028442f
C23 VDD2.n8 B 0.012741f
C24 VDD2.n9 B 0.022393f
C25 VDD2.n10 B 0.012387f
C26 VDD2.n11 B 0.028442f
C27 VDD2.n12 B 0.012741f
C28 VDD2.n13 B 0.022393f
C29 VDD2.n14 B 0.012033f
C30 VDD2.n15 B 0.028442f
C31 VDD2.n16 B 0.012741f
C32 VDD2.n17 B 0.022393f
C33 VDD2.n18 B 0.012033f
C34 VDD2.n19 B 0.028442f
C35 VDD2.n20 B 0.012741f
C36 VDD2.n21 B 0.022393f
C37 VDD2.n22 B 0.012033f
C38 VDD2.n23 B 0.028442f
C39 VDD2.n24 B 0.012741f
C40 VDD2.n25 B 0.022393f
C41 VDD2.n26 B 0.012033f
C42 VDD2.n27 B 0.028442f
C43 VDD2.n28 B 0.012741f
C44 VDD2.n29 B 0.022393f
C45 VDD2.n30 B 0.012033f
C46 VDD2.n31 B 0.021331f
C47 VDD2.n32 B 0.016802f
C48 VDD2.t5 B 0.047147f
C49 VDD2.n33 B 0.164301f
C50 VDD2.n34 B 1.79048f
C51 VDD2.n35 B 0.012033f
C52 VDD2.n36 B 0.012741f
C53 VDD2.n37 B 0.028442f
C54 VDD2.n38 B 0.028442f
C55 VDD2.n39 B 0.012741f
C56 VDD2.n40 B 0.012033f
C57 VDD2.n41 B 0.022393f
C58 VDD2.n42 B 0.022393f
C59 VDD2.n43 B 0.012033f
C60 VDD2.n44 B 0.012741f
C61 VDD2.n45 B 0.028442f
C62 VDD2.n46 B 0.028442f
C63 VDD2.n47 B 0.012741f
C64 VDD2.n48 B 0.012033f
C65 VDD2.n49 B 0.022393f
C66 VDD2.n50 B 0.022393f
C67 VDD2.n51 B 0.012033f
C68 VDD2.n52 B 0.012741f
C69 VDD2.n53 B 0.028442f
C70 VDD2.n54 B 0.028442f
C71 VDD2.n55 B 0.012741f
C72 VDD2.n56 B 0.012033f
C73 VDD2.n57 B 0.022393f
C74 VDD2.n58 B 0.022393f
C75 VDD2.n59 B 0.012033f
C76 VDD2.n60 B 0.012741f
C77 VDD2.n61 B 0.028442f
C78 VDD2.n62 B 0.028442f
C79 VDD2.n63 B 0.012741f
C80 VDD2.n64 B 0.012033f
C81 VDD2.n65 B 0.022393f
C82 VDD2.n66 B 0.022393f
C83 VDD2.n67 B 0.012033f
C84 VDD2.n68 B 0.012741f
C85 VDD2.n69 B 0.028442f
C86 VDD2.n70 B 0.028442f
C87 VDD2.n71 B 0.012741f
C88 VDD2.n72 B 0.012033f
C89 VDD2.n73 B 0.022393f
C90 VDD2.n74 B 0.022393f
C91 VDD2.n75 B 0.012033f
C92 VDD2.n76 B 0.012033f
C93 VDD2.n77 B 0.012741f
C94 VDD2.n78 B 0.028442f
C95 VDD2.n79 B 0.028442f
C96 VDD2.n80 B 0.028442f
C97 VDD2.n81 B 0.012387f
C98 VDD2.n82 B 0.012033f
C99 VDD2.n83 B 0.022393f
C100 VDD2.n84 B 0.022393f
C101 VDD2.n85 B 0.012033f
C102 VDD2.n86 B 0.012741f
C103 VDD2.n87 B 0.028442f
C104 VDD2.n88 B 0.028442f
C105 VDD2.n89 B 0.012741f
C106 VDD2.n90 B 0.012033f
C107 VDD2.n91 B 0.022393f
C108 VDD2.n92 B 0.022393f
C109 VDD2.n93 B 0.012033f
C110 VDD2.n94 B 0.012741f
C111 VDD2.n95 B 0.028442f
C112 VDD2.n96 B 0.061839f
C113 VDD2.n97 B 0.012741f
C114 VDD2.n98 B 0.012033f
C115 VDD2.n99 B 0.052067f
C116 VDD2.n100 B 0.054594f
C117 VDD2.t3 B 0.322949f
C118 VDD2.t7 B 0.322949f
C119 VDD2.n101 B 2.94357f
C120 VDD2.n102 B 0.466272f
C121 VDD2.t6 B 0.322949f
C122 VDD2.t1 B 0.322949f
C123 VDD2.n103 B 2.95016f
C124 VDD2.n104 B 2.39266f
C125 VDD2.n105 B 0.031627f
C126 VDD2.n106 B 0.022393f
C127 VDD2.n107 B 0.012033f
C128 VDD2.n108 B 0.028442f
C129 VDD2.n109 B 0.012741f
C130 VDD2.n110 B 0.022393f
C131 VDD2.n111 B 0.012033f
C132 VDD2.n112 B 0.028442f
C133 VDD2.n113 B 0.012741f
C134 VDD2.n114 B 0.022393f
C135 VDD2.n115 B 0.012387f
C136 VDD2.n116 B 0.028442f
C137 VDD2.n117 B 0.012033f
C138 VDD2.n118 B 0.012741f
C139 VDD2.n119 B 0.022393f
C140 VDD2.n120 B 0.012033f
C141 VDD2.n121 B 0.028442f
C142 VDD2.n122 B 0.012741f
C143 VDD2.n123 B 0.022393f
C144 VDD2.n124 B 0.012033f
C145 VDD2.n125 B 0.028442f
C146 VDD2.n126 B 0.012741f
C147 VDD2.n127 B 0.022393f
C148 VDD2.n128 B 0.012033f
C149 VDD2.n129 B 0.028442f
C150 VDD2.n130 B 0.012741f
C151 VDD2.n131 B 0.022393f
C152 VDD2.n132 B 0.012033f
C153 VDD2.n133 B 0.028442f
C154 VDD2.n134 B 0.012741f
C155 VDD2.n135 B 0.022393f
C156 VDD2.n136 B 0.012033f
C157 VDD2.n137 B 0.021331f
C158 VDD2.n138 B 0.016802f
C159 VDD2.t8 B 0.047147f
C160 VDD2.n139 B 0.164301f
C161 VDD2.n140 B 1.79048f
C162 VDD2.n141 B 0.012033f
C163 VDD2.n142 B 0.012741f
C164 VDD2.n143 B 0.028442f
C165 VDD2.n144 B 0.028442f
C166 VDD2.n145 B 0.012741f
C167 VDD2.n146 B 0.012033f
C168 VDD2.n147 B 0.022393f
C169 VDD2.n148 B 0.022393f
C170 VDD2.n149 B 0.012033f
C171 VDD2.n150 B 0.012741f
C172 VDD2.n151 B 0.028442f
C173 VDD2.n152 B 0.028442f
C174 VDD2.n153 B 0.012741f
C175 VDD2.n154 B 0.012033f
C176 VDD2.n155 B 0.022393f
C177 VDD2.n156 B 0.022393f
C178 VDD2.n157 B 0.012033f
C179 VDD2.n158 B 0.012741f
C180 VDD2.n159 B 0.028442f
C181 VDD2.n160 B 0.028442f
C182 VDD2.n161 B 0.012741f
C183 VDD2.n162 B 0.012033f
C184 VDD2.n163 B 0.022393f
C185 VDD2.n164 B 0.022393f
C186 VDD2.n165 B 0.012033f
C187 VDD2.n166 B 0.012741f
C188 VDD2.n167 B 0.028442f
C189 VDD2.n168 B 0.028442f
C190 VDD2.n169 B 0.012741f
C191 VDD2.n170 B 0.012033f
C192 VDD2.n171 B 0.022393f
C193 VDD2.n172 B 0.022393f
C194 VDD2.n173 B 0.012033f
C195 VDD2.n174 B 0.012741f
C196 VDD2.n175 B 0.028442f
C197 VDD2.n176 B 0.028442f
C198 VDD2.n177 B 0.012741f
C199 VDD2.n178 B 0.012033f
C200 VDD2.n179 B 0.022393f
C201 VDD2.n180 B 0.022393f
C202 VDD2.n181 B 0.012033f
C203 VDD2.n182 B 0.012741f
C204 VDD2.n183 B 0.028442f
C205 VDD2.n184 B 0.028442f
C206 VDD2.n185 B 0.028442f
C207 VDD2.n186 B 0.012387f
C208 VDD2.n187 B 0.012033f
C209 VDD2.n188 B 0.022393f
C210 VDD2.n189 B 0.022393f
C211 VDD2.n190 B 0.012033f
C212 VDD2.n191 B 0.012741f
C213 VDD2.n192 B 0.028442f
C214 VDD2.n193 B 0.028442f
C215 VDD2.n194 B 0.012741f
C216 VDD2.n195 B 0.012033f
C217 VDD2.n196 B 0.022393f
C218 VDD2.n197 B 0.022393f
C219 VDD2.n198 B 0.012033f
C220 VDD2.n199 B 0.012741f
C221 VDD2.n200 B 0.028442f
C222 VDD2.n201 B 0.061839f
C223 VDD2.n202 B 0.012741f
C224 VDD2.n203 B 0.012033f
C225 VDD2.n204 B 0.052067f
C226 VDD2.n205 B 0.050098f
C227 VDD2.n206 B 2.60477f
C228 VDD2.t4 B 0.322949f
C229 VDD2.t0 B 0.322949f
C230 VDD2.n207 B 2.94358f
C231 VDD2.n208 B 0.325798f
C232 VDD2.t9 B 0.322949f
C233 VDD2.t2 B 0.322949f
C234 VDD2.n209 B 2.95013f
C235 VN.n0 B 0.030179f
C236 VN.t8 B 2.13658f
C237 VN.n1 B 0.052897f
C238 VN.n2 B 0.030179f
C239 VN.t3 B 2.13658f
C240 VN.n3 B 0.045811f
C241 VN.n4 B 0.030179f
C242 VN.t6 B 2.13658f
C243 VN.n5 B 0.821308f
C244 VN.t4 B 2.22323f
C245 VN.n6 B 0.819287f
C246 VN.n7 B 0.189553f
C247 VN.n8 B 0.053624f
C248 VN.n9 B 0.030482f
C249 VN.t2 B 2.13658f
C250 VN.n10 B 0.753212f
C251 VN.n11 B 0.045811f
C252 VN.n12 B 0.030179f
C253 VN.n13 B 0.030179f
C254 VN.n14 B 0.030179f
C255 VN.n15 B 0.030482f
C256 VN.n16 B 0.053624f
C257 VN.n17 B 0.753212f
C258 VN.n18 B 0.029032f
C259 VN.n19 B 0.030179f
C260 VN.n20 B 0.030179f
C261 VN.n21 B 0.030179f
C262 VN.n22 B 0.032959f
C263 VN.n23 B 0.043505f
C264 VN.n24 B 0.812386f
C265 VN.n25 B 0.028234f
C266 VN.n26 B 0.030179f
C267 VN.t1 B 2.13658f
C268 VN.n27 B 0.052897f
C269 VN.n28 B 0.030179f
C270 VN.t5 B 2.13658f
C271 VN.n29 B 0.045811f
C272 VN.n30 B 0.030179f
C273 VN.t9 B 2.13658f
C274 VN.n31 B 0.753212f
C275 VN.t0 B 2.13658f
C276 VN.n32 B 0.821308f
C277 VN.t7 B 2.22323f
C278 VN.n33 B 0.819287f
C279 VN.n34 B 0.189553f
C280 VN.n35 B 0.053624f
C281 VN.n36 B 0.030482f
C282 VN.n37 B 0.045811f
C283 VN.n38 B 0.030179f
C284 VN.n39 B 0.030179f
C285 VN.n40 B 0.030179f
C286 VN.n41 B 0.030482f
C287 VN.n42 B 0.053624f
C288 VN.n43 B 0.753212f
C289 VN.n44 B 0.029032f
C290 VN.n45 B 0.030179f
C291 VN.n46 B 0.030179f
C292 VN.n47 B 0.030179f
C293 VN.n48 B 0.032959f
C294 VN.n49 B 0.043505f
C295 VN.n50 B 0.812386f
C296 VN.n51 B 1.72947f
C297 VTAIL.t2 B 0.339137f
C298 VTAIL.t1 B 0.339137f
C299 VTAIL.n0 B 3.01892f
C300 VTAIL.n1 B 0.417977f
C301 VTAIL.n2 B 0.033212f
C302 VTAIL.n3 B 0.023516f
C303 VTAIL.n4 B 0.012636f
C304 VTAIL.n5 B 0.029868f
C305 VTAIL.n6 B 0.01338f
C306 VTAIL.n7 B 0.023516f
C307 VTAIL.n8 B 0.012636f
C308 VTAIL.n9 B 0.029868f
C309 VTAIL.n10 B 0.01338f
C310 VTAIL.n11 B 0.023516f
C311 VTAIL.n12 B 0.013008f
C312 VTAIL.n13 B 0.029868f
C313 VTAIL.n14 B 0.01338f
C314 VTAIL.n15 B 0.023516f
C315 VTAIL.n16 B 0.012636f
C316 VTAIL.n17 B 0.029868f
C317 VTAIL.n18 B 0.01338f
C318 VTAIL.n19 B 0.023516f
C319 VTAIL.n20 B 0.012636f
C320 VTAIL.n21 B 0.029868f
C321 VTAIL.n22 B 0.01338f
C322 VTAIL.n23 B 0.023516f
C323 VTAIL.n24 B 0.012636f
C324 VTAIL.n25 B 0.029868f
C325 VTAIL.n26 B 0.01338f
C326 VTAIL.n27 B 0.023516f
C327 VTAIL.n28 B 0.012636f
C328 VTAIL.n29 B 0.029868f
C329 VTAIL.n30 B 0.01338f
C330 VTAIL.n31 B 0.023516f
C331 VTAIL.n32 B 0.012636f
C332 VTAIL.n33 B 0.022401f
C333 VTAIL.n34 B 0.017644f
C334 VTAIL.t15 B 0.04951f
C335 VTAIL.n35 B 0.172536f
C336 VTAIL.n36 B 1.88023f
C337 VTAIL.n37 B 0.012636f
C338 VTAIL.n38 B 0.01338f
C339 VTAIL.n39 B 0.029868f
C340 VTAIL.n40 B 0.029868f
C341 VTAIL.n41 B 0.01338f
C342 VTAIL.n42 B 0.012636f
C343 VTAIL.n43 B 0.023516f
C344 VTAIL.n44 B 0.023516f
C345 VTAIL.n45 B 0.012636f
C346 VTAIL.n46 B 0.01338f
C347 VTAIL.n47 B 0.029868f
C348 VTAIL.n48 B 0.029868f
C349 VTAIL.n49 B 0.01338f
C350 VTAIL.n50 B 0.012636f
C351 VTAIL.n51 B 0.023516f
C352 VTAIL.n52 B 0.023516f
C353 VTAIL.n53 B 0.012636f
C354 VTAIL.n54 B 0.01338f
C355 VTAIL.n55 B 0.029868f
C356 VTAIL.n56 B 0.029868f
C357 VTAIL.n57 B 0.01338f
C358 VTAIL.n58 B 0.012636f
C359 VTAIL.n59 B 0.023516f
C360 VTAIL.n60 B 0.023516f
C361 VTAIL.n61 B 0.012636f
C362 VTAIL.n62 B 0.01338f
C363 VTAIL.n63 B 0.029868f
C364 VTAIL.n64 B 0.029868f
C365 VTAIL.n65 B 0.01338f
C366 VTAIL.n66 B 0.012636f
C367 VTAIL.n67 B 0.023516f
C368 VTAIL.n68 B 0.023516f
C369 VTAIL.n69 B 0.012636f
C370 VTAIL.n70 B 0.01338f
C371 VTAIL.n71 B 0.029868f
C372 VTAIL.n72 B 0.029868f
C373 VTAIL.n73 B 0.01338f
C374 VTAIL.n74 B 0.012636f
C375 VTAIL.n75 B 0.023516f
C376 VTAIL.n76 B 0.023516f
C377 VTAIL.n77 B 0.012636f
C378 VTAIL.n78 B 0.012636f
C379 VTAIL.n79 B 0.01338f
C380 VTAIL.n80 B 0.029868f
C381 VTAIL.n81 B 0.029868f
C382 VTAIL.n82 B 0.029868f
C383 VTAIL.n83 B 0.013008f
C384 VTAIL.n84 B 0.012636f
C385 VTAIL.n85 B 0.023516f
C386 VTAIL.n86 B 0.023516f
C387 VTAIL.n87 B 0.012636f
C388 VTAIL.n88 B 0.01338f
C389 VTAIL.n89 B 0.029868f
C390 VTAIL.n90 B 0.029868f
C391 VTAIL.n91 B 0.01338f
C392 VTAIL.n92 B 0.012636f
C393 VTAIL.n93 B 0.023516f
C394 VTAIL.n94 B 0.023516f
C395 VTAIL.n95 B 0.012636f
C396 VTAIL.n96 B 0.01338f
C397 VTAIL.n97 B 0.029868f
C398 VTAIL.n98 B 0.064939f
C399 VTAIL.n99 B 0.01338f
C400 VTAIL.n100 B 0.012636f
C401 VTAIL.n101 B 0.054677f
C402 VTAIL.n102 B 0.036375f
C403 VTAIL.n103 B 0.226355f
C404 VTAIL.t17 B 0.339137f
C405 VTAIL.t14 B 0.339137f
C406 VTAIL.n104 B 3.01892f
C407 VTAIL.n105 B 0.463212f
C408 VTAIL.t12 B 0.339137f
C409 VTAIL.t18 B 0.339137f
C410 VTAIL.n106 B 3.01892f
C411 VTAIL.n107 B 2.08842f
C412 VTAIL.t0 B 0.339137f
C413 VTAIL.t3 B 0.339137f
C414 VTAIL.n108 B 3.01893f
C415 VTAIL.n109 B 2.08841f
C416 VTAIL.t4 B 0.339137f
C417 VTAIL.t8 B 0.339137f
C418 VTAIL.n110 B 3.01893f
C419 VTAIL.n111 B 0.463198f
C420 VTAIL.n112 B 0.033212f
C421 VTAIL.n113 B 0.023516f
C422 VTAIL.n114 B 0.012636f
C423 VTAIL.n115 B 0.029868f
C424 VTAIL.n116 B 0.01338f
C425 VTAIL.n117 B 0.023516f
C426 VTAIL.n118 B 0.012636f
C427 VTAIL.n119 B 0.029868f
C428 VTAIL.n120 B 0.01338f
C429 VTAIL.n121 B 0.023516f
C430 VTAIL.n122 B 0.013008f
C431 VTAIL.n123 B 0.029868f
C432 VTAIL.n124 B 0.012636f
C433 VTAIL.n125 B 0.01338f
C434 VTAIL.n126 B 0.023516f
C435 VTAIL.n127 B 0.012636f
C436 VTAIL.n128 B 0.029868f
C437 VTAIL.n129 B 0.01338f
C438 VTAIL.n130 B 0.023516f
C439 VTAIL.n131 B 0.012636f
C440 VTAIL.n132 B 0.029868f
C441 VTAIL.n133 B 0.01338f
C442 VTAIL.n134 B 0.023516f
C443 VTAIL.n135 B 0.012636f
C444 VTAIL.n136 B 0.029868f
C445 VTAIL.n137 B 0.01338f
C446 VTAIL.n138 B 0.023516f
C447 VTAIL.n139 B 0.012636f
C448 VTAIL.n140 B 0.029868f
C449 VTAIL.n141 B 0.01338f
C450 VTAIL.n142 B 0.023516f
C451 VTAIL.n143 B 0.012636f
C452 VTAIL.n144 B 0.022401f
C453 VTAIL.n145 B 0.017644f
C454 VTAIL.t5 B 0.04951f
C455 VTAIL.n146 B 0.172536f
C456 VTAIL.n147 B 1.88023f
C457 VTAIL.n148 B 0.012636f
C458 VTAIL.n149 B 0.01338f
C459 VTAIL.n150 B 0.029868f
C460 VTAIL.n151 B 0.029868f
C461 VTAIL.n152 B 0.01338f
C462 VTAIL.n153 B 0.012636f
C463 VTAIL.n154 B 0.023516f
C464 VTAIL.n155 B 0.023516f
C465 VTAIL.n156 B 0.012636f
C466 VTAIL.n157 B 0.01338f
C467 VTAIL.n158 B 0.029868f
C468 VTAIL.n159 B 0.029868f
C469 VTAIL.n160 B 0.01338f
C470 VTAIL.n161 B 0.012636f
C471 VTAIL.n162 B 0.023516f
C472 VTAIL.n163 B 0.023516f
C473 VTAIL.n164 B 0.012636f
C474 VTAIL.n165 B 0.01338f
C475 VTAIL.n166 B 0.029868f
C476 VTAIL.n167 B 0.029868f
C477 VTAIL.n168 B 0.01338f
C478 VTAIL.n169 B 0.012636f
C479 VTAIL.n170 B 0.023516f
C480 VTAIL.n171 B 0.023516f
C481 VTAIL.n172 B 0.012636f
C482 VTAIL.n173 B 0.01338f
C483 VTAIL.n174 B 0.029868f
C484 VTAIL.n175 B 0.029868f
C485 VTAIL.n176 B 0.01338f
C486 VTAIL.n177 B 0.012636f
C487 VTAIL.n178 B 0.023516f
C488 VTAIL.n179 B 0.023516f
C489 VTAIL.n180 B 0.012636f
C490 VTAIL.n181 B 0.01338f
C491 VTAIL.n182 B 0.029868f
C492 VTAIL.n183 B 0.029868f
C493 VTAIL.n184 B 0.01338f
C494 VTAIL.n185 B 0.012636f
C495 VTAIL.n186 B 0.023516f
C496 VTAIL.n187 B 0.023516f
C497 VTAIL.n188 B 0.012636f
C498 VTAIL.n189 B 0.01338f
C499 VTAIL.n190 B 0.029868f
C500 VTAIL.n191 B 0.029868f
C501 VTAIL.n192 B 0.029868f
C502 VTAIL.n193 B 0.013008f
C503 VTAIL.n194 B 0.012636f
C504 VTAIL.n195 B 0.023516f
C505 VTAIL.n196 B 0.023516f
C506 VTAIL.n197 B 0.012636f
C507 VTAIL.n198 B 0.01338f
C508 VTAIL.n199 B 0.029868f
C509 VTAIL.n200 B 0.029868f
C510 VTAIL.n201 B 0.01338f
C511 VTAIL.n202 B 0.012636f
C512 VTAIL.n203 B 0.023516f
C513 VTAIL.n204 B 0.023516f
C514 VTAIL.n205 B 0.012636f
C515 VTAIL.n206 B 0.01338f
C516 VTAIL.n207 B 0.029868f
C517 VTAIL.n208 B 0.064939f
C518 VTAIL.n209 B 0.01338f
C519 VTAIL.n210 B 0.012636f
C520 VTAIL.n211 B 0.054677f
C521 VTAIL.n212 B 0.036375f
C522 VTAIL.n213 B 0.226355f
C523 VTAIL.t16 B 0.339137f
C524 VTAIL.t10 B 0.339137f
C525 VTAIL.n214 B 3.01893f
C526 VTAIL.n215 B 0.441969f
C527 VTAIL.t13 B 0.339137f
C528 VTAIL.t19 B 0.339137f
C529 VTAIL.n216 B 3.01893f
C530 VTAIL.n217 B 0.463198f
C531 VTAIL.n218 B 0.033212f
C532 VTAIL.n219 B 0.023516f
C533 VTAIL.n220 B 0.012636f
C534 VTAIL.n221 B 0.029868f
C535 VTAIL.n222 B 0.01338f
C536 VTAIL.n223 B 0.023516f
C537 VTAIL.n224 B 0.012636f
C538 VTAIL.n225 B 0.029868f
C539 VTAIL.n226 B 0.01338f
C540 VTAIL.n227 B 0.023516f
C541 VTAIL.n228 B 0.013008f
C542 VTAIL.n229 B 0.029868f
C543 VTAIL.n230 B 0.012636f
C544 VTAIL.n231 B 0.01338f
C545 VTAIL.n232 B 0.023516f
C546 VTAIL.n233 B 0.012636f
C547 VTAIL.n234 B 0.029868f
C548 VTAIL.n235 B 0.01338f
C549 VTAIL.n236 B 0.023516f
C550 VTAIL.n237 B 0.012636f
C551 VTAIL.n238 B 0.029868f
C552 VTAIL.n239 B 0.01338f
C553 VTAIL.n240 B 0.023516f
C554 VTAIL.n241 B 0.012636f
C555 VTAIL.n242 B 0.029868f
C556 VTAIL.n243 B 0.01338f
C557 VTAIL.n244 B 0.023516f
C558 VTAIL.n245 B 0.012636f
C559 VTAIL.n246 B 0.029868f
C560 VTAIL.n247 B 0.01338f
C561 VTAIL.n248 B 0.023516f
C562 VTAIL.n249 B 0.012636f
C563 VTAIL.n250 B 0.022401f
C564 VTAIL.n251 B 0.017644f
C565 VTAIL.t11 B 0.04951f
C566 VTAIL.n252 B 0.172536f
C567 VTAIL.n253 B 1.88023f
C568 VTAIL.n254 B 0.012636f
C569 VTAIL.n255 B 0.01338f
C570 VTAIL.n256 B 0.029868f
C571 VTAIL.n257 B 0.029868f
C572 VTAIL.n258 B 0.01338f
C573 VTAIL.n259 B 0.012636f
C574 VTAIL.n260 B 0.023516f
C575 VTAIL.n261 B 0.023516f
C576 VTAIL.n262 B 0.012636f
C577 VTAIL.n263 B 0.01338f
C578 VTAIL.n264 B 0.029868f
C579 VTAIL.n265 B 0.029868f
C580 VTAIL.n266 B 0.01338f
C581 VTAIL.n267 B 0.012636f
C582 VTAIL.n268 B 0.023516f
C583 VTAIL.n269 B 0.023516f
C584 VTAIL.n270 B 0.012636f
C585 VTAIL.n271 B 0.01338f
C586 VTAIL.n272 B 0.029868f
C587 VTAIL.n273 B 0.029868f
C588 VTAIL.n274 B 0.01338f
C589 VTAIL.n275 B 0.012636f
C590 VTAIL.n276 B 0.023516f
C591 VTAIL.n277 B 0.023516f
C592 VTAIL.n278 B 0.012636f
C593 VTAIL.n279 B 0.01338f
C594 VTAIL.n280 B 0.029868f
C595 VTAIL.n281 B 0.029868f
C596 VTAIL.n282 B 0.01338f
C597 VTAIL.n283 B 0.012636f
C598 VTAIL.n284 B 0.023516f
C599 VTAIL.n285 B 0.023516f
C600 VTAIL.n286 B 0.012636f
C601 VTAIL.n287 B 0.01338f
C602 VTAIL.n288 B 0.029868f
C603 VTAIL.n289 B 0.029868f
C604 VTAIL.n290 B 0.01338f
C605 VTAIL.n291 B 0.012636f
C606 VTAIL.n292 B 0.023516f
C607 VTAIL.n293 B 0.023516f
C608 VTAIL.n294 B 0.012636f
C609 VTAIL.n295 B 0.01338f
C610 VTAIL.n296 B 0.029868f
C611 VTAIL.n297 B 0.029868f
C612 VTAIL.n298 B 0.029868f
C613 VTAIL.n299 B 0.013008f
C614 VTAIL.n300 B 0.012636f
C615 VTAIL.n301 B 0.023516f
C616 VTAIL.n302 B 0.023516f
C617 VTAIL.n303 B 0.012636f
C618 VTAIL.n304 B 0.01338f
C619 VTAIL.n305 B 0.029868f
C620 VTAIL.n306 B 0.029868f
C621 VTAIL.n307 B 0.01338f
C622 VTAIL.n308 B 0.012636f
C623 VTAIL.n309 B 0.023516f
C624 VTAIL.n310 B 0.023516f
C625 VTAIL.n311 B 0.012636f
C626 VTAIL.n312 B 0.01338f
C627 VTAIL.n313 B 0.029868f
C628 VTAIL.n314 B 0.064939f
C629 VTAIL.n315 B 0.01338f
C630 VTAIL.n316 B 0.012636f
C631 VTAIL.n317 B 0.054677f
C632 VTAIL.n318 B 0.036375f
C633 VTAIL.n319 B 1.75913f
C634 VTAIL.n320 B 0.033212f
C635 VTAIL.n321 B 0.023516f
C636 VTAIL.n322 B 0.012636f
C637 VTAIL.n323 B 0.029868f
C638 VTAIL.n324 B 0.01338f
C639 VTAIL.n325 B 0.023516f
C640 VTAIL.n326 B 0.012636f
C641 VTAIL.n327 B 0.029868f
C642 VTAIL.n328 B 0.01338f
C643 VTAIL.n329 B 0.023516f
C644 VTAIL.n330 B 0.013008f
C645 VTAIL.n331 B 0.029868f
C646 VTAIL.n332 B 0.01338f
C647 VTAIL.n333 B 0.023516f
C648 VTAIL.n334 B 0.012636f
C649 VTAIL.n335 B 0.029868f
C650 VTAIL.n336 B 0.01338f
C651 VTAIL.n337 B 0.023516f
C652 VTAIL.n338 B 0.012636f
C653 VTAIL.n339 B 0.029868f
C654 VTAIL.n340 B 0.01338f
C655 VTAIL.n341 B 0.023516f
C656 VTAIL.n342 B 0.012636f
C657 VTAIL.n343 B 0.029868f
C658 VTAIL.n344 B 0.01338f
C659 VTAIL.n345 B 0.023516f
C660 VTAIL.n346 B 0.012636f
C661 VTAIL.n347 B 0.029868f
C662 VTAIL.n348 B 0.01338f
C663 VTAIL.n349 B 0.023516f
C664 VTAIL.n350 B 0.012636f
C665 VTAIL.n351 B 0.022401f
C666 VTAIL.n352 B 0.017644f
C667 VTAIL.t9 B 0.04951f
C668 VTAIL.n353 B 0.172536f
C669 VTAIL.n354 B 1.88023f
C670 VTAIL.n355 B 0.012636f
C671 VTAIL.n356 B 0.01338f
C672 VTAIL.n357 B 0.029868f
C673 VTAIL.n358 B 0.029868f
C674 VTAIL.n359 B 0.01338f
C675 VTAIL.n360 B 0.012636f
C676 VTAIL.n361 B 0.023516f
C677 VTAIL.n362 B 0.023516f
C678 VTAIL.n363 B 0.012636f
C679 VTAIL.n364 B 0.01338f
C680 VTAIL.n365 B 0.029868f
C681 VTAIL.n366 B 0.029868f
C682 VTAIL.n367 B 0.01338f
C683 VTAIL.n368 B 0.012636f
C684 VTAIL.n369 B 0.023516f
C685 VTAIL.n370 B 0.023516f
C686 VTAIL.n371 B 0.012636f
C687 VTAIL.n372 B 0.01338f
C688 VTAIL.n373 B 0.029868f
C689 VTAIL.n374 B 0.029868f
C690 VTAIL.n375 B 0.01338f
C691 VTAIL.n376 B 0.012636f
C692 VTAIL.n377 B 0.023516f
C693 VTAIL.n378 B 0.023516f
C694 VTAIL.n379 B 0.012636f
C695 VTAIL.n380 B 0.01338f
C696 VTAIL.n381 B 0.029868f
C697 VTAIL.n382 B 0.029868f
C698 VTAIL.n383 B 0.01338f
C699 VTAIL.n384 B 0.012636f
C700 VTAIL.n385 B 0.023516f
C701 VTAIL.n386 B 0.023516f
C702 VTAIL.n387 B 0.012636f
C703 VTAIL.n388 B 0.01338f
C704 VTAIL.n389 B 0.029868f
C705 VTAIL.n390 B 0.029868f
C706 VTAIL.n391 B 0.01338f
C707 VTAIL.n392 B 0.012636f
C708 VTAIL.n393 B 0.023516f
C709 VTAIL.n394 B 0.023516f
C710 VTAIL.n395 B 0.012636f
C711 VTAIL.n396 B 0.012636f
C712 VTAIL.n397 B 0.01338f
C713 VTAIL.n398 B 0.029868f
C714 VTAIL.n399 B 0.029868f
C715 VTAIL.n400 B 0.029868f
C716 VTAIL.n401 B 0.013008f
C717 VTAIL.n402 B 0.012636f
C718 VTAIL.n403 B 0.023516f
C719 VTAIL.n404 B 0.023516f
C720 VTAIL.n405 B 0.012636f
C721 VTAIL.n406 B 0.01338f
C722 VTAIL.n407 B 0.029868f
C723 VTAIL.n408 B 0.029868f
C724 VTAIL.n409 B 0.01338f
C725 VTAIL.n410 B 0.012636f
C726 VTAIL.n411 B 0.023516f
C727 VTAIL.n412 B 0.023516f
C728 VTAIL.n413 B 0.012636f
C729 VTAIL.n414 B 0.01338f
C730 VTAIL.n415 B 0.029868f
C731 VTAIL.n416 B 0.064939f
C732 VTAIL.n417 B 0.01338f
C733 VTAIL.n418 B 0.012636f
C734 VTAIL.n419 B 0.054677f
C735 VTAIL.n420 B 0.036375f
C736 VTAIL.n421 B 1.75913f
C737 VTAIL.t6 B 0.339137f
C738 VTAIL.t7 B 0.339137f
C739 VTAIL.n422 B 3.01892f
C740 VTAIL.n423 B 0.373558f
C741 VDD1.n0 B 0.031866f
C742 VDD1.n1 B 0.022563f
C743 VDD1.n2 B 0.012124f
C744 VDD1.n3 B 0.028657f
C745 VDD1.n4 B 0.012837f
C746 VDD1.n5 B 0.022563f
C747 VDD1.n6 B 0.012124f
C748 VDD1.n7 B 0.028657f
C749 VDD1.n8 B 0.012837f
C750 VDD1.n9 B 0.022563f
C751 VDD1.n10 B 0.012481f
C752 VDD1.n11 B 0.028657f
C753 VDD1.n12 B 0.012124f
C754 VDD1.n13 B 0.012837f
C755 VDD1.n14 B 0.022563f
C756 VDD1.n15 B 0.012124f
C757 VDD1.n16 B 0.028657f
C758 VDD1.n17 B 0.012837f
C759 VDD1.n18 B 0.022563f
C760 VDD1.n19 B 0.012124f
C761 VDD1.n20 B 0.028657f
C762 VDD1.n21 B 0.012837f
C763 VDD1.n22 B 0.022563f
C764 VDD1.n23 B 0.012124f
C765 VDD1.n24 B 0.028657f
C766 VDD1.n25 B 0.012837f
C767 VDD1.n26 B 0.022563f
C768 VDD1.n27 B 0.012124f
C769 VDD1.n28 B 0.028657f
C770 VDD1.n29 B 0.012837f
C771 VDD1.n30 B 0.022563f
C772 VDD1.n31 B 0.012124f
C773 VDD1.n32 B 0.021493f
C774 VDD1.n33 B 0.016929f
C775 VDD1.t6 B 0.047504f
C776 VDD1.n34 B 0.165545f
C777 VDD1.n35 B 1.80404f
C778 VDD1.n36 B 0.012124f
C779 VDD1.n37 B 0.012837f
C780 VDD1.n38 B 0.028657f
C781 VDD1.n39 B 0.028657f
C782 VDD1.n40 B 0.012837f
C783 VDD1.n41 B 0.012124f
C784 VDD1.n42 B 0.022563f
C785 VDD1.n43 B 0.022563f
C786 VDD1.n44 B 0.012124f
C787 VDD1.n45 B 0.012837f
C788 VDD1.n46 B 0.028657f
C789 VDD1.n47 B 0.028657f
C790 VDD1.n48 B 0.012837f
C791 VDD1.n49 B 0.012124f
C792 VDD1.n50 B 0.022563f
C793 VDD1.n51 B 0.022563f
C794 VDD1.n52 B 0.012124f
C795 VDD1.n53 B 0.012837f
C796 VDD1.n54 B 0.028657f
C797 VDD1.n55 B 0.028657f
C798 VDD1.n56 B 0.012837f
C799 VDD1.n57 B 0.012124f
C800 VDD1.n58 B 0.022563f
C801 VDD1.n59 B 0.022563f
C802 VDD1.n60 B 0.012124f
C803 VDD1.n61 B 0.012837f
C804 VDD1.n62 B 0.028657f
C805 VDD1.n63 B 0.028657f
C806 VDD1.n64 B 0.012837f
C807 VDD1.n65 B 0.012124f
C808 VDD1.n66 B 0.022563f
C809 VDD1.n67 B 0.022563f
C810 VDD1.n68 B 0.012124f
C811 VDD1.n69 B 0.012837f
C812 VDD1.n70 B 0.028657f
C813 VDD1.n71 B 0.028657f
C814 VDD1.n72 B 0.012837f
C815 VDD1.n73 B 0.012124f
C816 VDD1.n74 B 0.022563f
C817 VDD1.n75 B 0.022563f
C818 VDD1.n76 B 0.012124f
C819 VDD1.n77 B 0.012837f
C820 VDD1.n78 B 0.028657f
C821 VDD1.n79 B 0.028657f
C822 VDD1.n80 B 0.028657f
C823 VDD1.n81 B 0.012481f
C824 VDD1.n82 B 0.012124f
C825 VDD1.n83 B 0.022563f
C826 VDD1.n84 B 0.022563f
C827 VDD1.n85 B 0.012124f
C828 VDD1.n86 B 0.012837f
C829 VDD1.n87 B 0.028657f
C830 VDD1.n88 B 0.028657f
C831 VDD1.n89 B 0.012837f
C832 VDD1.n90 B 0.012124f
C833 VDD1.n91 B 0.022563f
C834 VDD1.n92 B 0.022563f
C835 VDD1.n93 B 0.012124f
C836 VDD1.n94 B 0.012837f
C837 VDD1.n95 B 0.028657f
C838 VDD1.n96 B 0.062308f
C839 VDD1.n97 B 0.012837f
C840 VDD1.n98 B 0.012124f
C841 VDD1.n99 B 0.052461f
C842 VDD1.n100 B 0.055007f
C843 VDD1.t2 B 0.325395f
C844 VDD1.t5 B 0.325395f
C845 VDD1.n101 B 2.96588f
C846 VDD1.n102 B 0.476413f
C847 VDD1.n103 B 0.031866f
C848 VDD1.n104 B 0.022563f
C849 VDD1.n105 B 0.012124f
C850 VDD1.n106 B 0.028657f
C851 VDD1.n107 B 0.012837f
C852 VDD1.n108 B 0.022563f
C853 VDD1.n109 B 0.012124f
C854 VDD1.n110 B 0.028657f
C855 VDD1.n111 B 0.012837f
C856 VDD1.n112 B 0.022563f
C857 VDD1.n113 B 0.012481f
C858 VDD1.n114 B 0.028657f
C859 VDD1.n115 B 0.012837f
C860 VDD1.n116 B 0.022563f
C861 VDD1.n117 B 0.012124f
C862 VDD1.n118 B 0.028657f
C863 VDD1.n119 B 0.012837f
C864 VDD1.n120 B 0.022563f
C865 VDD1.n121 B 0.012124f
C866 VDD1.n122 B 0.028657f
C867 VDD1.n123 B 0.012837f
C868 VDD1.n124 B 0.022563f
C869 VDD1.n125 B 0.012124f
C870 VDD1.n126 B 0.028657f
C871 VDD1.n127 B 0.012837f
C872 VDD1.n128 B 0.022563f
C873 VDD1.n129 B 0.012124f
C874 VDD1.n130 B 0.028657f
C875 VDD1.n131 B 0.012837f
C876 VDD1.n132 B 0.022563f
C877 VDD1.n133 B 0.012124f
C878 VDD1.n134 B 0.021493f
C879 VDD1.n135 B 0.016929f
C880 VDD1.t4 B 0.047504f
C881 VDD1.n136 B 0.165545f
C882 VDD1.n137 B 1.80404f
C883 VDD1.n138 B 0.012124f
C884 VDD1.n139 B 0.012837f
C885 VDD1.n140 B 0.028657f
C886 VDD1.n141 B 0.028657f
C887 VDD1.n142 B 0.012837f
C888 VDD1.n143 B 0.012124f
C889 VDD1.n144 B 0.022563f
C890 VDD1.n145 B 0.022563f
C891 VDD1.n146 B 0.012124f
C892 VDD1.n147 B 0.012837f
C893 VDD1.n148 B 0.028657f
C894 VDD1.n149 B 0.028657f
C895 VDD1.n150 B 0.012837f
C896 VDD1.n151 B 0.012124f
C897 VDD1.n152 B 0.022563f
C898 VDD1.n153 B 0.022563f
C899 VDD1.n154 B 0.012124f
C900 VDD1.n155 B 0.012837f
C901 VDD1.n156 B 0.028657f
C902 VDD1.n157 B 0.028657f
C903 VDD1.n158 B 0.012837f
C904 VDD1.n159 B 0.012124f
C905 VDD1.n160 B 0.022563f
C906 VDD1.n161 B 0.022563f
C907 VDD1.n162 B 0.012124f
C908 VDD1.n163 B 0.012837f
C909 VDD1.n164 B 0.028657f
C910 VDD1.n165 B 0.028657f
C911 VDD1.n166 B 0.012837f
C912 VDD1.n167 B 0.012124f
C913 VDD1.n168 B 0.022563f
C914 VDD1.n169 B 0.022563f
C915 VDD1.n170 B 0.012124f
C916 VDD1.n171 B 0.012837f
C917 VDD1.n172 B 0.028657f
C918 VDD1.n173 B 0.028657f
C919 VDD1.n174 B 0.012837f
C920 VDD1.n175 B 0.012124f
C921 VDD1.n176 B 0.022563f
C922 VDD1.n177 B 0.022563f
C923 VDD1.n178 B 0.012124f
C924 VDD1.n179 B 0.012124f
C925 VDD1.n180 B 0.012837f
C926 VDD1.n181 B 0.028657f
C927 VDD1.n182 B 0.028657f
C928 VDD1.n183 B 0.028657f
C929 VDD1.n184 B 0.012481f
C930 VDD1.n185 B 0.012124f
C931 VDD1.n186 B 0.022563f
C932 VDD1.n187 B 0.022563f
C933 VDD1.n188 B 0.012124f
C934 VDD1.n189 B 0.012837f
C935 VDD1.n190 B 0.028657f
C936 VDD1.n191 B 0.028657f
C937 VDD1.n192 B 0.012837f
C938 VDD1.n193 B 0.012124f
C939 VDD1.n194 B 0.022563f
C940 VDD1.n195 B 0.022563f
C941 VDD1.n196 B 0.012124f
C942 VDD1.n197 B 0.012837f
C943 VDD1.n198 B 0.028657f
C944 VDD1.n199 B 0.062308f
C945 VDD1.n200 B 0.012837f
C946 VDD1.n201 B 0.012124f
C947 VDD1.n202 B 0.052461f
C948 VDD1.n203 B 0.055007f
C949 VDD1.t0 B 0.325395f
C950 VDD1.t7 B 0.325395f
C951 VDD1.n204 B 2.96587f
C952 VDD1.n205 B 0.469804f
C953 VDD1.t8 B 0.325395f
C954 VDD1.t9 B 0.325395f
C955 VDD1.n206 B 2.97251f
C956 VDD1.n207 B 2.4981f
C957 VDD1.t1 B 0.325395f
C958 VDD1.t3 B 0.325395f
C959 VDD1.n208 B 2.96587f
C960 VDD1.n209 B 2.85127f
C961 VP.n0 B 0.030564f
C962 VP.t4 B 2.16385f
C963 VP.n1 B 0.053573f
C964 VP.n2 B 0.030564f
C965 VP.t5 B 2.16385f
C966 VP.n3 B 0.046396f
C967 VP.n4 B 0.030564f
C968 VP.t1 B 2.16385f
C969 VP.n5 B 0.762827f
C970 VP.n6 B 0.030564f
C971 VP.n7 B 0.044061f
C972 VP.n8 B 0.030564f
C973 VP.t8 B 2.16385f
C974 VP.n9 B 0.053573f
C975 VP.n10 B 0.030564f
C976 VP.t0 B 2.16385f
C977 VP.n11 B 0.046396f
C978 VP.n12 B 0.030564f
C979 VP.t9 B 2.16385f
C980 VP.n13 B 0.831792f
C981 VP.t3 B 2.25161f
C982 VP.n14 B 0.829745f
C983 VP.n15 B 0.191973f
C984 VP.n16 B 0.054309f
C985 VP.n17 B 0.030871f
C986 VP.t6 B 2.16385f
C987 VP.n18 B 0.762827f
C988 VP.n19 B 0.046396f
C989 VP.n20 B 0.030564f
C990 VP.n21 B 0.030564f
C991 VP.n22 B 0.030564f
C992 VP.n23 B 0.030871f
C993 VP.n24 B 0.054309f
C994 VP.n25 B 0.762827f
C995 VP.n26 B 0.029403f
C996 VP.n27 B 0.030564f
C997 VP.n28 B 0.030564f
C998 VP.n29 B 0.030564f
C999 VP.n30 B 0.03338f
C1000 VP.n31 B 0.044061f
C1001 VP.n32 B 0.822757f
C1002 VP.n33 B 1.7317f
C1003 VP.t7 B 2.16385f
C1004 VP.n34 B 0.822757f
C1005 VP.n35 B 1.75312f
C1006 VP.n36 B 0.030564f
C1007 VP.n37 B 0.030564f
C1008 VP.n38 B 0.03338f
C1009 VP.n39 B 0.053573f
C1010 VP.n40 B 0.029403f
C1011 VP.n41 B 0.030564f
C1012 VP.n42 B 0.030564f
C1013 VP.n43 B 0.054309f
C1014 VP.n44 B 0.030871f
C1015 VP.t2 B 2.16385f
C1016 VP.n45 B 0.762827f
C1017 VP.n46 B 0.046396f
C1018 VP.n47 B 0.030564f
C1019 VP.n48 B 0.030564f
C1020 VP.n49 B 0.030564f
C1021 VP.n50 B 0.030871f
C1022 VP.n51 B 0.054309f
C1023 VP.n52 B 0.762827f
C1024 VP.n53 B 0.029403f
C1025 VP.n54 B 0.030564f
C1026 VP.n55 B 0.030564f
C1027 VP.n56 B 0.030564f
C1028 VP.n57 B 0.03338f
C1029 VP.n58 B 0.044061f
C1030 VP.n59 B 0.822756f
C1031 VP.n60 B 0.028595f
.ends

