* NGSPICE file created from diff_pair_sample_0820.ext - technology: sky130A

.subckt diff_pair_sample_0820 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=6.3921 pd=33.56 as=0 ps=0 w=16.39 l=2.28
X1 VTAIL.t19 VN.t0 VDD2.t7 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X2 VDD1.t9 VP.t0 VTAIL.t9 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=6.3921 ps=33.56 w=16.39 l=2.28
X3 B.t8 B.t6 B.t7 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=6.3921 pd=33.56 as=0 ps=0 w=16.39 l=2.28
X4 VDD2.t4 VN.t1 VTAIL.t18 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X5 VTAIL.t8 VP.t1 VDD1.t8 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X6 VDD2.t8 VN.t2 VTAIL.t17 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=6.3921 ps=33.56 w=16.39 l=2.28
X7 VTAIL.t7 VP.t2 VDD1.t7 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X8 VTAIL.t5 VP.t3 VDD1.t6 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X9 VDD1.t5 VP.t4 VTAIL.t6 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=6.3921 pd=33.56 as=2.70435 ps=16.72 w=16.39 l=2.28
X10 VDD2.t3 VN.t3 VTAIL.t16 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=6.3921 ps=33.56 w=16.39 l=2.28
X11 VTAIL.t15 VN.t4 VDD2.t5 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X12 VDD1.t4 VP.t5 VTAIL.t0 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X13 VDD1.t3 VP.t6 VTAIL.t2 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X14 B.t5 B.t3 B.t4 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=6.3921 pd=33.56 as=0 ps=0 w=16.39 l=2.28
X15 VTAIL.t14 VN.t5 VDD2.t2 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X16 VDD2.t1 VN.t6 VTAIL.t13 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X17 VDD2.t6 VN.t7 VTAIL.t12 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=6.3921 pd=33.56 as=2.70435 ps=16.72 w=16.39 l=2.28
X18 VTAIL.t11 VN.t8 VDD2.t0 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X19 VTAIL.t4 VP.t7 VDD1.t2 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=2.70435 ps=16.72 w=16.39 l=2.28
X20 VDD2.t9 VN.t9 VTAIL.t10 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=6.3921 pd=33.56 as=2.70435 ps=16.72 w=16.39 l=2.28
X21 VDD1.t1 VP.t8 VTAIL.t3 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=2.70435 pd=16.72 as=6.3921 ps=33.56 w=16.39 l=2.28
X22 B.t2 B.t0 B.t1 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=6.3921 pd=33.56 as=0 ps=0 w=16.39 l=2.28
X23 VDD1.t0 VP.t9 VTAIL.t1 w_n4102_n4246# sky130_fd_pr__pfet_01v8 ad=6.3921 pd=33.56 as=2.70435 ps=16.72 w=16.39 l=2.28
R0 B.n662 B.n93 585
R1 B.n664 B.n663 585
R2 B.n665 B.n92 585
R3 B.n667 B.n666 585
R4 B.n668 B.n91 585
R5 B.n670 B.n669 585
R6 B.n671 B.n90 585
R7 B.n673 B.n672 585
R8 B.n674 B.n89 585
R9 B.n676 B.n675 585
R10 B.n677 B.n88 585
R11 B.n679 B.n678 585
R12 B.n680 B.n87 585
R13 B.n682 B.n681 585
R14 B.n683 B.n86 585
R15 B.n685 B.n684 585
R16 B.n686 B.n85 585
R17 B.n688 B.n687 585
R18 B.n689 B.n84 585
R19 B.n691 B.n690 585
R20 B.n692 B.n83 585
R21 B.n694 B.n693 585
R22 B.n695 B.n82 585
R23 B.n697 B.n696 585
R24 B.n698 B.n81 585
R25 B.n700 B.n699 585
R26 B.n701 B.n80 585
R27 B.n703 B.n702 585
R28 B.n704 B.n79 585
R29 B.n706 B.n705 585
R30 B.n707 B.n78 585
R31 B.n709 B.n708 585
R32 B.n710 B.n77 585
R33 B.n712 B.n711 585
R34 B.n713 B.n76 585
R35 B.n715 B.n714 585
R36 B.n716 B.n75 585
R37 B.n718 B.n717 585
R38 B.n719 B.n74 585
R39 B.n721 B.n720 585
R40 B.n722 B.n73 585
R41 B.n724 B.n723 585
R42 B.n725 B.n72 585
R43 B.n727 B.n726 585
R44 B.n728 B.n71 585
R45 B.n730 B.n729 585
R46 B.n731 B.n70 585
R47 B.n733 B.n732 585
R48 B.n734 B.n69 585
R49 B.n736 B.n735 585
R50 B.n737 B.n68 585
R51 B.n739 B.n738 585
R52 B.n740 B.n67 585
R53 B.n742 B.n741 585
R54 B.n743 B.n64 585
R55 B.n746 B.n745 585
R56 B.n747 B.n63 585
R57 B.n749 B.n748 585
R58 B.n750 B.n62 585
R59 B.n752 B.n751 585
R60 B.n753 B.n61 585
R61 B.n755 B.n754 585
R62 B.n756 B.n57 585
R63 B.n758 B.n757 585
R64 B.n759 B.n56 585
R65 B.n761 B.n760 585
R66 B.n762 B.n55 585
R67 B.n764 B.n763 585
R68 B.n765 B.n54 585
R69 B.n767 B.n766 585
R70 B.n768 B.n53 585
R71 B.n770 B.n769 585
R72 B.n771 B.n52 585
R73 B.n773 B.n772 585
R74 B.n774 B.n51 585
R75 B.n776 B.n775 585
R76 B.n777 B.n50 585
R77 B.n779 B.n778 585
R78 B.n780 B.n49 585
R79 B.n782 B.n781 585
R80 B.n783 B.n48 585
R81 B.n785 B.n784 585
R82 B.n786 B.n47 585
R83 B.n788 B.n787 585
R84 B.n789 B.n46 585
R85 B.n791 B.n790 585
R86 B.n792 B.n45 585
R87 B.n794 B.n793 585
R88 B.n795 B.n44 585
R89 B.n797 B.n796 585
R90 B.n798 B.n43 585
R91 B.n800 B.n799 585
R92 B.n801 B.n42 585
R93 B.n803 B.n802 585
R94 B.n804 B.n41 585
R95 B.n806 B.n805 585
R96 B.n807 B.n40 585
R97 B.n809 B.n808 585
R98 B.n810 B.n39 585
R99 B.n812 B.n811 585
R100 B.n813 B.n38 585
R101 B.n815 B.n814 585
R102 B.n816 B.n37 585
R103 B.n818 B.n817 585
R104 B.n819 B.n36 585
R105 B.n821 B.n820 585
R106 B.n822 B.n35 585
R107 B.n824 B.n823 585
R108 B.n825 B.n34 585
R109 B.n827 B.n826 585
R110 B.n828 B.n33 585
R111 B.n830 B.n829 585
R112 B.n831 B.n32 585
R113 B.n833 B.n832 585
R114 B.n834 B.n31 585
R115 B.n836 B.n835 585
R116 B.n837 B.n30 585
R117 B.n839 B.n838 585
R118 B.n840 B.n29 585
R119 B.n661 B.n660 585
R120 B.n659 B.n94 585
R121 B.n658 B.n657 585
R122 B.n656 B.n95 585
R123 B.n655 B.n654 585
R124 B.n653 B.n96 585
R125 B.n652 B.n651 585
R126 B.n650 B.n97 585
R127 B.n649 B.n648 585
R128 B.n647 B.n98 585
R129 B.n646 B.n645 585
R130 B.n644 B.n99 585
R131 B.n643 B.n642 585
R132 B.n641 B.n100 585
R133 B.n640 B.n639 585
R134 B.n638 B.n101 585
R135 B.n637 B.n636 585
R136 B.n635 B.n102 585
R137 B.n634 B.n633 585
R138 B.n632 B.n103 585
R139 B.n631 B.n630 585
R140 B.n629 B.n104 585
R141 B.n628 B.n627 585
R142 B.n626 B.n105 585
R143 B.n625 B.n624 585
R144 B.n623 B.n106 585
R145 B.n622 B.n621 585
R146 B.n620 B.n107 585
R147 B.n619 B.n618 585
R148 B.n617 B.n108 585
R149 B.n616 B.n615 585
R150 B.n614 B.n109 585
R151 B.n613 B.n612 585
R152 B.n611 B.n110 585
R153 B.n610 B.n609 585
R154 B.n608 B.n111 585
R155 B.n607 B.n606 585
R156 B.n605 B.n112 585
R157 B.n604 B.n603 585
R158 B.n602 B.n113 585
R159 B.n601 B.n600 585
R160 B.n599 B.n114 585
R161 B.n598 B.n597 585
R162 B.n596 B.n115 585
R163 B.n595 B.n594 585
R164 B.n593 B.n116 585
R165 B.n592 B.n591 585
R166 B.n590 B.n117 585
R167 B.n589 B.n588 585
R168 B.n587 B.n118 585
R169 B.n586 B.n585 585
R170 B.n584 B.n119 585
R171 B.n583 B.n582 585
R172 B.n581 B.n120 585
R173 B.n580 B.n579 585
R174 B.n578 B.n121 585
R175 B.n577 B.n576 585
R176 B.n575 B.n122 585
R177 B.n574 B.n573 585
R178 B.n572 B.n123 585
R179 B.n571 B.n570 585
R180 B.n569 B.n124 585
R181 B.n568 B.n567 585
R182 B.n566 B.n125 585
R183 B.n565 B.n564 585
R184 B.n563 B.n126 585
R185 B.n562 B.n561 585
R186 B.n560 B.n127 585
R187 B.n559 B.n558 585
R188 B.n557 B.n128 585
R189 B.n556 B.n555 585
R190 B.n554 B.n129 585
R191 B.n553 B.n552 585
R192 B.n551 B.n130 585
R193 B.n550 B.n549 585
R194 B.n548 B.n131 585
R195 B.n547 B.n546 585
R196 B.n545 B.n132 585
R197 B.n544 B.n543 585
R198 B.n542 B.n133 585
R199 B.n541 B.n540 585
R200 B.n539 B.n134 585
R201 B.n538 B.n537 585
R202 B.n536 B.n135 585
R203 B.n535 B.n534 585
R204 B.n533 B.n136 585
R205 B.n532 B.n531 585
R206 B.n530 B.n137 585
R207 B.n529 B.n528 585
R208 B.n527 B.n138 585
R209 B.n526 B.n525 585
R210 B.n524 B.n139 585
R211 B.n523 B.n522 585
R212 B.n521 B.n140 585
R213 B.n520 B.n519 585
R214 B.n518 B.n141 585
R215 B.n517 B.n516 585
R216 B.n515 B.n142 585
R217 B.n514 B.n513 585
R218 B.n512 B.n143 585
R219 B.n511 B.n510 585
R220 B.n509 B.n144 585
R221 B.n508 B.n507 585
R222 B.n506 B.n145 585
R223 B.n505 B.n504 585
R224 B.n503 B.n146 585
R225 B.n502 B.n501 585
R226 B.n500 B.n147 585
R227 B.n499 B.n498 585
R228 B.n316 B.n209 585
R229 B.n318 B.n317 585
R230 B.n319 B.n208 585
R231 B.n321 B.n320 585
R232 B.n322 B.n207 585
R233 B.n324 B.n323 585
R234 B.n325 B.n206 585
R235 B.n327 B.n326 585
R236 B.n328 B.n205 585
R237 B.n330 B.n329 585
R238 B.n331 B.n204 585
R239 B.n333 B.n332 585
R240 B.n334 B.n203 585
R241 B.n336 B.n335 585
R242 B.n337 B.n202 585
R243 B.n339 B.n338 585
R244 B.n340 B.n201 585
R245 B.n342 B.n341 585
R246 B.n343 B.n200 585
R247 B.n345 B.n344 585
R248 B.n346 B.n199 585
R249 B.n348 B.n347 585
R250 B.n349 B.n198 585
R251 B.n351 B.n350 585
R252 B.n352 B.n197 585
R253 B.n354 B.n353 585
R254 B.n355 B.n196 585
R255 B.n357 B.n356 585
R256 B.n358 B.n195 585
R257 B.n360 B.n359 585
R258 B.n361 B.n194 585
R259 B.n363 B.n362 585
R260 B.n364 B.n193 585
R261 B.n366 B.n365 585
R262 B.n367 B.n192 585
R263 B.n369 B.n368 585
R264 B.n370 B.n191 585
R265 B.n372 B.n371 585
R266 B.n373 B.n190 585
R267 B.n375 B.n374 585
R268 B.n376 B.n189 585
R269 B.n378 B.n377 585
R270 B.n379 B.n188 585
R271 B.n381 B.n380 585
R272 B.n382 B.n187 585
R273 B.n384 B.n383 585
R274 B.n385 B.n186 585
R275 B.n387 B.n386 585
R276 B.n388 B.n185 585
R277 B.n390 B.n389 585
R278 B.n391 B.n184 585
R279 B.n393 B.n392 585
R280 B.n394 B.n183 585
R281 B.n396 B.n395 585
R282 B.n397 B.n180 585
R283 B.n400 B.n399 585
R284 B.n401 B.n179 585
R285 B.n403 B.n402 585
R286 B.n404 B.n178 585
R287 B.n406 B.n405 585
R288 B.n407 B.n177 585
R289 B.n409 B.n408 585
R290 B.n410 B.n176 585
R291 B.n415 B.n414 585
R292 B.n416 B.n175 585
R293 B.n418 B.n417 585
R294 B.n419 B.n174 585
R295 B.n421 B.n420 585
R296 B.n422 B.n173 585
R297 B.n424 B.n423 585
R298 B.n425 B.n172 585
R299 B.n427 B.n426 585
R300 B.n428 B.n171 585
R301 B.n430 B.n429 585
R302 B.n431 B.n170 585
R303 B.n433 B.n432 585
R304 B.n434 B.n169 585
R305 B.n436 B.n435 585
R306 B.n437 B.n168 585
R307 B.n439 B.n438 585
R308 B.n440 B.n167 585
R309 B.n442 B.n441 585
R310 B.n443 B.n166 585
R311 B.n445 B.n444 585
R312 B.n446 B.n165 585
R313 B.n448 B.n447 585
R314 B.n449 B.n164 585
R315 B.n451 B.n450 585
R316 B.n452 B.n163 585
R317 B.n454 B.n453 585
R318 B.n455 B.n162 585
R319 B.n457 B.n456 585
R320 B.n458 B.n161 585
R321 B.n460 B.n459 585
R322 B.n461 B.n160 585
R323 B.n463 B.n462 585
R324 B.n464 B.n159 585
R325 B.n466 B.n465 585
R326 B.n467 B.n158 585
R327 B.n469 B.n468 585
R328 B.n470 B.n157 585
R329 B.n472 B.n471 585
R330 B.n473 B.n156 585
R331 B.n475 B.n474 585
R332 B.n476 B.n155 585
R333 B.n478 B.n477 585
R334 B.n479 B.n154 585
R335 B.n481 B.n480 585
R336 B.n482 B.n153 585
R337 B.n484 B.n483 585
R338 B.n485 B.n152 585
R339 B.n487 B.n486 585
R340 B.n488 B.n151 585
R341 B.n490 B.n489 585
R342 B.n491 B.n150 585
R343 B.n493 B.n492 585
R344 B.n494 B.n149 585
R345 B.n496 B.n495 585
R346 B.n497 B.n148 585
R347 B.n315 B.n314 585
R348 B.n313 B.n210 585
R349 B.n312 B.n311 585
R350 B.n310 B.n211 585
R351 B.n309 B.n308 585
R352 B.n307 B.n212 585
R353 B.n306 B.n305 585
R354 B.n304 B.n213 585
R355 B.n303 B.n302 585
R356 B.n301 B.n214 585
R357 B.n300 B.n299 585
R358 B.n298 B.n215 585
R359 B.n297 B.n296 585
R360 B.n295 B.n216 585
R361 B.n294 B.n293 585
R362 B.n292 B.n217 585
R363 B.n291 B.n290 585
R364 B.n289 B.n218 585
R365 B.n288 B.n287 585
R366 B.n286 B.n219 585
R367 B.n285 B.n284 585
R368 B.n283 B.n220 585
R369 B.n282 B.n281 585
R370 B.n280 B.n221 585
R371 B.n279 B.n278 585
R372 B.n277 B.n222 585
R373 B.n276 B.n275 585
R374 B.n274 B.n223 585
R375 B.n273 B.n272 585
R376 B.n271 B.n224 585
R377 B.n270 B.n269 585
R378 B.n268 B.n225 585
R379 B.n267 B.n266 585
R380 B.n265 B.n226 585
R381 B.n264 B.n263 585
R382 B.n262 B.n227 585
R383 B.n261 B.n260 585
R384 B.n259 B.n228 585
R385 B.n258 B.n257 585
R386 B.n256 B.n229 585
R387 B.n255 B.n254 585
R388 B.n253 B.n230 585
R389 B.n252 B.n251 585
R390 B.n250 B.n231 585
R391 B.n249 B.n248 585
R392 B.n247 B.n232 585
R393 B.n246 B.n245 585
R394 B.n244 B.n233 585
R395 B.n243 B.n242 585
R396 B.n241 B.n234 585
R397 B.n240 B.n239 585
R398 B.n238 B.n235 585
R399 B.n237 B.n236 585
R400 B.n2 B.n0 585
R401 B.n921 B.n1 585
R402 B.n920 B.n919 585
R403 B.n918 B.n3 585
R404 B.n917 B.n916 585
R405 B.n915 B.n4 585
R406 B.n914 B.n913 585
R407 B.n912 B.n5 585
R408 B.n911 B.n910 585
R409 B.n909 B.n6 585
R410 B.n908 B.n907 585
R411 B.n906 B.n7 585
R412 B.n905 B.n904 585
R413 B.n903 B.n8 585
R414 B.n902 B.n901 585
R415 B.n900 B.n9 585
R416 B.n899 B.n898 585
R417 B.n897 B.n10 585
R418 B.n896 B.n895 585
R419 B.n894 B.n11 585
R420 B.n893 B.n892 585
R421 B.n891 B.n12 585
R422 B.n890 B.n889 585
R423 B.n888 B.n13 585
R424 B.n887 B.n886 585
R425 B.n885 B.n14 585
R426 B.n884 B.n883 585
R427 B.n882 B.n15 585
R428 B.n881 B.n880 585
R429 B.n879 B.n16 585
R430 B.n878 B.n877 585
R431 B.n876 B.n17 585
R432 B.n875 B.n874 585
R433 B.n873 B.n18 585
R434 B.n872 B.n871 585
R435 B.n870 B.n19 585
R436 B.n869 B.n868 585
R437 B.n867 B.n20 585
R438 B.n866 B.n865 585
R439 B.n864 B.n21 585
R440 B.n863 B.n862 585
R441 B.n861 B.n22 585
R442 B.n860 B.n859 585
R443 B.n858 B.n23 585
R444 B.n857 B.n856 585
R445 B.n855 B.n24 585
R446 B.n854 B.n853 585
R447 B.n852 B.n25 585
R448 B.n851 B.n850 585
R449 B.n849 B.n26 585
R450 B.n848 B.n847 585
R451 B.n846 B.n27 585
R452 B.n845 B.n844 585
R453 B.n843 B.n28 585
R454 B.n842 B.n841 585
R455 B.n923 B.n922 585
R456 B.n316 B.n315 497.305
R457 B.n842 B.n29 497.305
R458 B.n499 B.n148 497.305
R459 B.n662 B.n661 497.305
R460 B.n411 B.t0 380.752
R461 B.n181 B.t3 380.752
R462 B.n58 B.t9 380.752
R463 B.n65 B.t6 380.752
R464 B.n315 B.n210 163.367
R465 B.n311 B.n210 163.367
R466 B.n311 B.n310 163.367
R467 B.n310 B.n309 163.367
R468 B.n309 B.n212 163.367
R469 B.n305 B.n212 163.367
R470 B.n305 B.n304 163.367
R471 B.n304 B.n303 163.367
R472 B.n303 B.n214 163.367
R473 B.n299 B.n214 163.367
R474 B.n299 B.n298 163.367
R475 B.n298 B.n297 163.367
R476 B.n297 B.n216 163.367
R477 B.n293 B.n216 163.367
R478 B.n293 B.n292 163.367
R479 B.n292 B.n291 163.367
R480 B.n291 B.n218 163.367
R481 B.n287 B.n218 163.367
R482 B.n287 B.n286 163.367
R483 B.n286 B.n285 163.367
R484 B.n285 B.n220 163.367
R485 B.n281 B.n220 163.367
R486 B.n281 B.n280 163.367
R487 B.n280 B.n279 163.367
R488 B.n279 B.n222 163.367
R489 B.n275 B.n222 163.367
R490 B.n275 B.n274 163.367
R491 B.n274 B.n273 163.367
R492 B.n273 B.n224 163.367
R493 B.n269 B.n224 163.367
R494 B.n269 B.n268 163.367
R495 B.n268 B.n267 163.367
R496 B.n267 B.n226 163.367
R497 B.n263 B.n226 163.367
R498 B.n263 B.n262 163.367
R499 B.n262 B.n261 163.367
R500 B.n261 B.n228 163.367
R501 B.n257 B.n228 163.367
R502 B.n257 B.n256 163.367
R503 B.n256 B.n255 163.367
R504 B.n255 B.n230 163.367
R505 B.n251 B.n230 163.367
R506 B.n251 B.n250 163.367
R507 B.n250 B.n249 163.367
R508 B.n249 B.n232 163.367
R509 B.n245 B.n232 163.367
R510 B.n245 B.n244 163.367
R511 B.n244 B.n243 163.367
R512 B.n243 B.n234 163.367
R513 B.n239 B.n234 163.367
R514 B.n239 B.n238 163.367
R515 B.n238 B.n237 163.367
R516 B.n237 B.n2 163.367
R517 B.n922 B.n2 163.367
R518 B.n922 B.n921 163.367
R519 B.n921 B.n920 163.367
R520 B.n920 B.n3 163.367
R521 B.n916 B.n3 163.367
R522 B.n916 B.n915 163.367
R523 B.n915 B.n914 163.367
R524 B.n914 B.n5 163.367
R525 B.n910 B.n5 163.367
R526 B.n910 B.n909 163.367
R527 B.n909 B.n908 163.367
R528 B.n908 B.n7 163.367
R529 B.n904 B.n7 163.367
R530 B.n904 B.n903 163.367
R531 B.n903 B.n902 163.367
R532 B.n902 B.n9 163.367
R533 B.n898 B.n9 163.367
R534 B.n898 B.n897 163.367
R535 B.n897 B.n896 163.367
R536 B.n896 B.n11 163.367
R537 B.n892 B.n11 163.367
R538 B.n892 B.n891 163.367
R539 B.n891 B.n890 163.367
R540 B.n890 B.n13 163.367
R541 B.n886 B.n13 163.367
R542 B.n886 B.n885 163.367
R543 B.n885 B.n884 163.367
R544 B.n884 B.n15 163.367
R545 B.n880 B.n15 163.367
R546 B.n880 B.n879 163.367
R547 B.n879 B.n878 163.367
R548 B.n878 B.n17 163.367
R549 B.n874 B.n17 163.367
R550 B.n874 B.n873 163.367
R551 B.n873 B.n872 163.367
R552 B.n872 B.n19 163.367
R553 B.n868 B.n19 163.367
R554 B.n868 B.n867 163.367
R555 B.n867 B.n866 163.367
R556 B.n866 B.n21 163.367
R557 B.n862 B.n21 163.367
R558 B.n862 B.n861 163.367
R559 B.n861 B.n860 163.367
R560 B.n860 B.n23 163.367
R561 B.n856 B.n23 163.367
R562 B.n856 B.n855 163.367
R563 B.n855 B.n854 163.367
R564 B.n854 B.n25 163.367
R565 B.n850 B.n25 163.367
R566 B.n850 B.n849 163.367
R567 B.n849 B.n848 163.367
R568 B.n848 B.n27 163.367
R569 B.n844 B.n27 163.367
R570 B.n844 B.n843 163.367
R571 B.n843 B.n842 163.367
R572 B.n317 B.n316 163.367
R573 B.n317 B.n208 163.367
R574 B.n321 B.n208 163.367
R575 B.n322 B.n321 163.367
R576 B.n323 B.n322 163.367
R577 B.n323 B.n206 163.367
R578 B.n327 B.n206 163.367
R579 B.n328 B.n327 163.367
R580 B.n329 B.n328 163.367
R581 B.n329 B.n204 163.367
R582 B.n333 B.n204 163.367
R583 B.n334 B.n333 163.367
R584 B.n335 B.n334 163.367
R585 B.n335 B.n202 163.367
R586 B.n339 B.n202 163.367
R587 B.n340 B.n339 163.367
R588 B.n341 B.n340 163.367
R589 B.n341 B.n200 163.367
R590 B.n345 B.n200 163.367
R591 B.n346 B.n345 163.367
R592 B.n347 B.n346 163.367
R593 B.n347 B.n198 163.367
R594 B.n351 B.n198 163.367
R595 B.n352 B.n351 163.367
R596 B.n353 B.n352 163.367
R597 B.n353 B.n196 163.367
R598 B.n357 B.n196 163.367
R599 B.n358 B.n357 163.367
R600 B.n359 B.n358 163.367
R601 B.n359 B.n194 163.367
R602 B.n363 B.n194 163.367
R603 B.n364 B.n363 163.367
R604 B.n365 B.n364 163.367
R605 B.n365 B.n192 163.367
R606 B.n369 B.n192 163.367
R607 B.n370 B.n369 163.367
R608 B.n371 B.n370 163.367
R609 B.n371 B.n190 163.367
R610 B.n375 B.n190 163.367
R611 B.n376 B.n375 163.367
R612 B.n377 B.n376 163.367
R613 B.n377 B.n188 163.367
R614 B.n381 B.n188 163.367
R615 B.n382 B.n381 163.367
R616 B.n383 B.n382 163.367
R617 B.n383 B.n186 163.367
R618 B.n387 B.n186 163.367
R619 B.n388 B.n387 163.367
R620 B.n389 B.n388 163.367
R621 B.n389 B.n184 163.367
R622 B.n393 B.n184 163.367
R623 B.n394 B.n393 163.367
R624 B.n395 B.n394 163.367
R625 B.n395 B.n180 163.367
R626 B.n400 B.n180 163.367
R627 B.n401 B.n400 163.367
R628 B.n402 B.n401 163.367
R629 B.n402 B.n178 163.367
R630 B.n406 B.n178 163.367
R631 B.n407 B.n406 163.367
R632 B.n408 B.n407 163.367
R633 B.n408 B.n176 163.367
R634 B.n415 B.n176 163.367
R635 B.n416 B.n415 163.367
R636 B.n417 B.n416 163.367
R637 B.n417 B.n174 163.367
R638 B.n421 B.n174 163.367
R639 B.n422 B.n421 163.367
R640 B.n423 B.n422 163.367
R641 B.n423 B.n172 163.367
R642 B.n427 B.n172 163.367
R643 B.n428 B.n427 163.367
R644 B.n429 B.n428 163.367
R645 B.n429 B.n170 163.367
R646 B.n433 B.n170 163.367
R647 B.n434 B.n433 163.367
R648 B.n435 B.n434 163.367
R649 B.n435 B.n168 163.367
R650 B.n439 B.n168 163.367
R651 B.n440 B.n439 163.367
R652 B.n441 B.n440 163.367
R653 B.n441 B.n166 163.367
R654 B.n445 B.n166 163.367
R655 B.n446 B.n445 163.367
R656 B.n447 B.n446 163.367
R657 B.n447 B.n164 163.367
R658 B.n451 B.n164 163.367
R659 B.n452 B.n451 163.367
R660 B.n453 B.n452 163.367
R661 B.n453 B.n162 163.367
R662 B.n457 B.n162 163.367
R663 B.n458 B.n457 163.367
R664 B.n459 B.n458 163.367
R665 B.n459 B.n160 163.367
R666 B.n463 B.n160 163.367
R667 B.n464 B.n463 163.367
R668 B.n465 B.n464 163.367
R669 B.n465 B.n158 163.367
R670 B.n469 B.n158 163.367
R671 B.n470 B.n469 163.367
R672 B.n471 B.n470 163.367
R673 B.n471 B.n156 163.367
R674 B.n475 B.n156 163.367
R675 B.n476 B.n475 163.367
R676 B.n477 B.n476 163.367
R677 B.n477 B.n154 163.367
R678 B.n481 B.n154 163.367
R679 B.n482 B.n481 163.367
R680 B.n483 B.n482 163.367
R681 B.n483 B.n152 163.367
R682 B.n487 B.n152 163.367
R683 B.n488 B.n487 163.367
R684 B.n489 B.n488 163.367
R685 B.n489 B.n150 163.367
R686 B.n493 B.n150 163.367
R687 B.n494 B.n493 163.367
R688 B.n495 B.n494 163.367
R689 B.n495 B.n148 163.367
R690 B.n500 B.n499 163.367
R691 B.n501 B.n500 163.367
R692 B.n501 B.n146 163.367
R693 B.n505 B.n146 163.367
R694 B.n506 B.n505 163.367
R695 B.n507 B.n506 163.367
R696 B.n507 B.n144 163.367
R697 B.n511 B.n144 163.367
R698 B.n512 B.n511 163.367
R699 B.n513 B.n512 163.367
R700 B.n513 B.n142 163.367
R701 B.n517 B.n142 163.367
R702 B.n518 B.n517 163.367
R703 B.n519 B.n518 163.367
R704 B.n519 B.n140 163.367
R705 B.n523 B.n140 163.367
R706 B.n524 B.n523 163.367
R707 B.n525 B.n524 163.367
R708 B.n525 B.n138 163.367
R709 B.n529 B.n138 163.367
R710 B.n530 B.n529 163.367
R711 B.n531 B.n530 163.367
R712 B.n531 B.n136 163.367
R713 B.n535 B.n136 163.367
R714 B.n536 B.n535 163.367
R715 B.n537 B.n536 163.367
R716 B.n537 B.n134 163.367
R717 B.n541 B.n134 163.367
R718 B.n542 B.n541 163.367
R719 B.n543 B.n542 163.367
R720 B.n543 B.n132 163.367
R721 B.n547 B.n132 163.367
R722 B.n548 B.n547 163.367
R723 B.n549 B.n548 163.367
R724 B.n549 B.n130 163.367
R725 B.n553 B.n130 163.367
R726 B.n554 B.n553 163.367
R727 B.n555 B.n554 163.367
R728 B.n555 B.n128 163.367
R729 B.n559 B.n128 163.367
R730 B.n560 B.n559 163.367
R731 B.n561 B.n560 163.367
R732 B.n561 B.n126 163.367
R733 B.n565 B.n126 163.367
R734 B.n566 B.n565 163.367
R735 B.n567 B.n566 163.367
R736 B.n567 B.n124 163.367
R737 B.n571 B.n124 163.367
R738 B.n572 B.n571 163.367
R739 B.n573 B.n572 163.367
R740 B.n573 B.n122 163.367
R741 B.n577 B.n122 163.367
R742 B.n578 B.n577 163.367
R743 B.n579 B.n578 163.367
R744 B.n579 B.n120 163.367
R745 B.n583 B.n120 163.367
R746 B.n584 B.n583 163.367
R747 B.n585 B.n584 163.367
R748 B.n585 B.n118 163.367
R749 B.n589 B.n118 163.367
R750 B.n590 B.n589 163.367
R751 B.n591 B.n590 163.367
R752 B.n591 B.n116 163.367
R753 B.n595 B.n116 163.367
R754 B.n596 B.n595 163.367
R755 B.n597 B.n596 163.367
R756 B.n597 B.n114 163.367
R757 B.n601 B.n114 163.367
R758 B.n602 B.n601 163.367
R759 B.n603 B.n602 163.367
R760 B.n603 B.n112 163.367
R761 B.n607 B.n112 163.367
R762 B.n608 B.n607 163.367
R763 B.n609 B.n608 163.367
R764 B.n609 B.n110 163.367
R765 B.n613 B.n110 163.367
R766 B.n614 B.n613 163.367
R767 B.n615 B.n614 163.367
R768 B.n615 B.n108 163.367
R769 B.n619 B.n108 163.367
R770 B.n620 B.n619 163.367
R771 B.n621 B.n620 163.367
R772 B.n621 B.n106 163.367
R773 B.n625 B.n106 163.367
R774 B.n626 B.n625 163.367
R775 B.n627 B.n626 163.367
R776 B.n627 B.n104 163.367
R777 B.n631 B.n104 163.367
R778 B.n632 B.n631 163.367
R779 B.n633 B.n632 163.367
R780 B.n633 B.n102 163.367
R781 B.n637 B.n102 163.367
R782 B.n638 B.n637 163.367
R783 B.n639 B.n638 163.367
R784 B.n639 B.n100 163.367
R785 B.n643 B.n100 163.367
R786 B.n644 B.n643 163.367
R787 B.n645 B.n644 163.367
R788 B.n645 B.n98 163.367
R789 B.n649 B.n98 163.367
R790 B.n650 B.n649 163.367
R791 B.n651 B.n650 163.367
R792 B.n651 B.n96 163.367
R793 B.n655 B.n96 163.367
R794 B.n656 B.n655 163.367
R795 B.n657 B.n656 163.367
R796 B.n657 B.n94 163.367
R797 B.n661 B.n94 163.367
R798 B.n838 B.n29 163.367
R799 B.n838 B.n837 163.367
R800 B.n837 B.n836 163.367
R801 B.n836 B.n31 163.367
R802 B.n832 B.n31 163.367
R803 B.n832 B.n831 163.367
R804 B.n831 B.n830 163.367
R805 B.n830 B.n33 163.367
R806 B.n826 B.n33 163.367
R807 B.n826 B.n825 163.367
R808 B.n825 B.n824 163.367
R809 B.n824 B.n35 163.367
R810 B.n820 B.n35 163.367
R811 B.n820 B.n819 163.367
R812 B.n819 B.n818 163.367
R813 B.n818 B.n37 163.367
R814 B.n814 B.n37 163.367
R815 B.n814 B.n813 163.367
R816 B.n813 B.n812 163.367
R817 B.n812 B.n39 163.367
R818 B.n808 B.n39 163.367
R819 B.n808 B.n807 163.367
R820 B.n807 B.n806 163.367
R821 B.n806 B.n41 163.367
R822 B.n802 B.n41 163.367
R823 B.n802 B.n801 163.367
R824 B.n801 B.n800 163.367
R825 B.n800 B.n43 163.367
R826 B.n796 B.n43 163.367
R827 B.n796 B.n795 163.367
R828 B.n795 B.n794 163.367
R829 B.n794 B.n45 163.367
R830 B.n790 B.n45 163.367
R831 B.n790 B.n789 163.367
R832 B.n789 B.n788 163.367
R833 B.n788 B.n47 163.367
R834 B.n784 B.n47 163.367
R835 B.n784 B.n783 163.367
R836 B.n783 B.n782 163.367
R837 B.n782 B.n49 163.367
R838 B.n778 B.n49 163.367
R839 B.n778 B.n777 163.367
R840 B.n777 B.n776 163.367
R841 B.n776 B.n51 163.367
R842 B.n772 B.n51 163.367
R843 B.n772 B.n771 163.367
R844 B.n771 B.n770 163.367
R845 B.n770 B.n53 163.367
R846 B.n766 B.n53 163.367
R847 B.n766 B.n765 163.367
R848 B.n765 B.n764 163.367
R849 B.n764 B.n55 163.367
R850 B.n760 B.n55 163.367
R851 B.n760 B.n759 163.367
R852 B.n759 B.n758 163.367
R853 B.n758 B.n57 163.367
R854 B.n754 B.n57 163.367
R855 B.n754 B.n753 163.367
R856 B.n753 B.n752 163.367
R857 B.n752 B.n62 163.367
R858 B.n748 B.n62 163.367
R859 B.n748 B.n747 163.367
R860 B.n747 B.n746 163.367
R861 B.n746 B.n64 163.367
R862 B.n741 B.n64 163.367
R863 B.n741 B.n740 163.367
R864 B.n740 B.n739 163.367
R865 B.n739 B.n68 163.367
R866 B.n735 B.n68 163.367
R867 B.n735 B.n734 163.367
R868 B.n734 B.n733 163.367
R869 B.n733 B.n70 163.367
R870 B.n729 B.n70 163.367
R871 B.n729 B.n728 163.367
R872 B.n728 B.n727 163.367
R873 B.n727 B.n72 163.367
R874 B.n723 B.n72 163.367
R875 B.n723 B.n722 163.367
R876 B.n722 B.n721 163.367
R877 B.n721 B.n74 163.367
R878 B.n717 B.n74 163.367
R879 B.n717 B.n716 163.367
R880 B.n716 B.n715 163.367
R881 B.n715 B.n76 163.367
R882 B.n711 B.n76 163.367
R883 B.n711 B.n710 163.367
R884 B.n710 B.n709 163.367
R885 B.n709 B.n78 163.367
R886 B.n705 B.n78 163.367
R887 B.n705 B.n704 163.367
R888 B.n704 B.n703 163.367
R889 B.n703 B.n80 163.367
R890 B.n699 B.n80 163.367
R891 B.n699 B.n698 163.367
R892 B.n698 B.n697 163.367
R893 B.n697 B.n82 163.367
R894 B.n693 B.n82 163.367
R895 B.n693 B.n692 163.367
R896 B.n692 B.n691 163.367
R897 B.n691 B.n84 163.367
R898 B.n687 B.n84 163.367
R899 B.n687 B.n686 163.367
R900 B.n686 B.n685 163.367
R901 B.n685 B.n86 163.367
R902 B.n681 B.n86 163.367
R903 B.n681 B.n680 163.367
R904 B.n680 B.n679 163.367
R905 B.n679 B.n88 163.367
R906 B.n675 B.n88 163.367
R907 B.n675 B.n674 163.367
R908 B.n674 B.n673 163.367
R909 B.n673 B.n90 163.367
R910 B.n669 B.n90 163.367
R911 B.n669 B.n668 163.367
R912 B.n668 B.n667 163.367
R913 B.n667 B.n92 163.367
R914 B.n663 B.n92 163.367
R915 B.n663 B.n662 163.367
R916 B.n411 B.t2 158.356
R917 B.n65 B.t7 158.356
R918 B.n181 B.t5 158.334
R919 B.n58 B.t10 158.334
R920 B.n412 B.t1 107.737
R921 B.n66 B.t8 107.737
R922 B.n182 B.t4 107.716
R923 B.n59 B.t11 107.716
R924 B.n413 B.n412 59.5399
R925 B.n398 B.n182 59.5399
R926 B.n60 B.n59 59.5399
R927 B.n744 B.n66 59.5399
R928 B.n412 B.n411 50.6187
R929 B.n182 B.n181 50.6187
R930 B.n59 B.n58 50.6187
R931 B.n66 B.n65 50.6187
R932 B.n841 B.n840 32.3127
R933 B.n660 B.n93 32.3127
R934 B.n498 B.n497 32.3127
R935 B.n314 B.n209 32.3127
R936 B B.n923 18.0485
R937 B.n840 B.n839 10.6151
R938 B.n839 B.n30 10.6151
R939 B.n835 B.n30 10.6151
R940 B.n835 B.n834 10.6151
R941 B.n834 B.n833 10.6151
R942 B.n833 B.n32 10.6151
R943 B.n829 B.n32 10.6151
R944 B.n829 B.n828 10.6151
R945 B.n828 B.n827 10.6151
R946 B.n827 B.n34 10.6151
R947 B.n823 B.n34 10.6151
R948 B.n823 B.n822 10.6151
R949 B.n822 B.n821 10.6151
R950 B.n821 B.n36 10.6151
R951 B.n817 B.n36 10.6151
R952 B.n817 B.n816 10.6151
R953 B.n816 B.n815 10.6151
R954 B.n815 B.n38 10.6151
R955 B.n811 B.n38 10.6151
R956 B.n811 B.n810 10.6151
R957 B.n810 B.n809 10.6151
R958 B.n809 B.n40 10.6151
R959 B.n805 B.n40 10.6151
R960 B.n805 B.n804 10.6151
R961 B.n804 B.n803 10.6151
R962 B.n803 B.n42 10.6151
R963 B.n799 B.n42 10.6151
R964 B.n799 B.n798 10.6151
R965 B.n798 B.n797 10.6151
R966 B.n797 B.n44 10.6151
R967 B.n793 B.n44 10.6151
R968 B.n793 B.n792 10.6151
R969 B.n792 B.n791 10.6151
R970 B.n791 B.n46 10.6151
R971 B.n787 B.n46 10.6151
R972 B.n787 B.n786 10.6151
R973 B.n786 B.n785 10.6151
R974 B.n785 B.n48 10.6151
R975 B.n781 B.n48 10.6151
R976 B.n781 B.n780 10.6151
R977 B.n780 B.n779 10.6151
R978 B.n779 B.n50 10.6151
R979 B.n775 B.n50 10.6151
R980 B.n775 B.n774 10.6151
R981 B.n774 B.n773 10.6151
R982 B.n773 B.n52 10.6151
R983 B.n769 B.n52 10.6151
R984 B.n769 B.n768 10.6151
R985 B.n768 B.n767 10.6151
R986 B.n767 B.n54 10.6151
R987 B.n763 B.n54 10.6151
R988 B.n763 B.n762 10.6151
R989 B.n762 B.n761 10.6151
R990 B.n761 B.n56 10.6151
R991 B.n757 B.n756 10.6151
R992 B.n756 B.n755 10.6151
R993 B.n755 B.n61 10.6151
R994 B.n751 B.n61 10.6151
R995 B.n751 B.n750 10.6151
R996 B.n750 B.n749 10.6151
R997 B.n749 B.n63 10.6151
R998 B.n745 B.n63 10.6151
R999 B.n743 B.n742 10.6151
R1000 B.n742 B.n67 10.6151
R1001 B.n738 B.n67 10.6151
R1002 B.n738 B.n737 10.6151
R1003 B.n737 B.n736 10.6151
R1004 B.n736 B.n69 10.6151
R1005 B.n732 B.n69 10.6151
R1006 B.n732 B.n731 10.6151
R1007 B.n731 B.n730 10.6151
R1008 B.n730 B.n71 10.6151
R1009 B.n726 B.n71 10.6151
R1010 B.n726 B.n725 10.6151
R1011 B.n725 B.n724 10.6151
R1012 B.n724 B.n73 10.6151
R1013 B.n720 B.n73 10.6151
R1014 B.n720 B.n719 10.6151
R1015 B.n719 B.n718 10.6151
R1016 B.n718 B.n75 10.6151
R1017 B.n714 B.n75 10.6151
R1018 B.n714 B.n713 10.6151
R1019 B.n713 B.n712 10.6151
R1020 B.n712 B.n77 10.6151
R1021 B.n708 B.n77 10.6151
R1022 B.n708 B.n707 10.6151
R1023 B.n707 B.n706 10.6151
R1024 B.n706 B.n79 10.6151
R1025 B.n702 B.n79 10.6151
R1026 B.n702 B.n701 10.6151
R1027 B.n701 B.n700 10.6151
R1028 B.n700 B.n81 10.6151
R1029 B.n696 B.n81 10.6151
R1030 B.n696 B.n695 10.6151
R1031 B.n695 B.n694 10.6151
R1032 B.n694 B.n83 10.6151
R1033 B.n690 B.n83 10.6151
R1034 B.n690 B.n689 10.6151
R1035 B.n689 B.n688 10.6151
R1036 B.n688 B.n85 10.6151
R1037 B.n684 B.n85 10.6151
R1038 B.n684 B.n683 10.6151
R1039 B.n683 B.n682 10.6151
R1040 B.n682 B.n87 10.6151
R1041 B.n678 B.n87 10.6151
R1042 B.n678 B.n677 10.6151
R1043 B.n677 B.n676 10.6151
R1044 B.n676 B.n89 10.6151
R1045 B.n672 B.n89 10.6151
R1046 B.n672 B.n671 10.6151
R1047 B.n671 B.n670 10.6151
R1048 B.n670 B.n91 10.6151
R1049 B.n666 B.n91 10.6151
R1050 B.n666 B.n665 10.6151
R1051 B.n665 B.n664 10.6151
R1052 B.n664 B.n93 10.6151
R1053 B.n498 B.n147 10.6151
R1054 B.n502 B.n147 10.6151
R1055 B.n503 B.n502 10.6151
R1056 B.n504 B.n503 10.6151
R1057 B.n504 B.n145 10.6151
R1058 B.n508 B.n145 10.6151
R1059 B.n509 B.n508 10.6151
R1060 B.n510 B.n509 10.6151
R1061 B.n510 B.n143 10.6151
R1062 B.n514 B.n143 10.6151
R1063 B.n515 B.n514 10.6151
R1064 B.n516 B.n515 10.6151
R1065 B.n516 B.n141 10.6151
R1066 B.n520 B.n141 10.6151
R1067 B.n521 B.n520 10.6151
R1068 B.n522 B.n521 10.6151
R1069 B.n522 B.n139 10.6151
R1070 B.n526 B.n139 10.6151
R1071 B.n527 B.n526 10.6151
R1072 B.n528 B.n527 10.6151
R1073 B.n528 B.n137 10.6151
R1074 B.n532 B.n137 10.6151
R1075 B.n533 B.n532 10.6151
R1076 B.n534 B.n533 10.6151
R1077 B.n534 B.n135 10.6151
R1078 B.n538 B.n135 10.6151
R1079 B.n539 B.n538 10.6151
R1080 B.n540 B.n539 10.6151
R1081 B.n540 B.n133 10.6151
R1082 B.n544 B.n133 10.6151
R1083 B.n545 B.n544 10.6151
R1084 B.n546 B.n545 10.6151
R1085 B.n546 B.n131 10.6151
R1086 B.n550 B.n131 10.6151
R1087 B.n551 B.n550 10.6151
R1088 B.n552 B.n551 10.6151
R1089 B.n552 B.n129 10.6151
R1090 B.n556 B.n129 10.6151
R1091 B.n557 B.n556 10.6151
R1092 B.n558 B.n557 10.6151
R1093 B.n558 B.n127 10.6151
R1094 B.n562 B.n127 10.6151
R1095 B.n563 B.n562 10.6151
R1096 B.n564 B.n563 10.6151
R1097 B.n564 B.n125 10.6151
R1098 B.n568 B.n125 10.6151
R1099 B.n569 B.n568 10.6151
R1100 B.n570 B.n569 10.6151
R1101 B.n570 B.n123 10.6151
R1102 B.n574 B.n123 10.6151
R1103 B.n575 B.n574 10.6151
R1104 B.n576 B.n575 10.6151
R1105 B.n576 B.n121 10.6151
R1106 B.n580 B.n121 10.6151
R1107 B.n581 B.n580 10.6151
R1108 B.n582 B.n581 10.6151
R1109 B.n582 B.n119 10.6151
R1110 B.n586 B.n119 10.6151
R1111 B.n587 B.n586 10.6151
R1112 B.n588 B.n587 10.6151
R1113 B.n588 B.n117 10.6151
R1114 B.n592 B.n117 10.6151
R1115 B.n593 B.n592 10.6151
R1116 B.n594 B.n593 10.6151
R1117 B.n594 B.n115 10.6151
R1118 B.n598 B.n115 10.6151
R1119 B.n599 B.n598 10.6151
R1120 B.n600 B.n599 10.6151
R1121 B.n600 B.n113 10.6151
R1122 B.n604 B.n113 10.6151
R1123 B.n605 B.n604 10.6151
R1124 B.n606 B.n605 10.6151
R1125 B.n606 B.n111 10.6151
R1126 B.n610 B.n111 10.6151
R1127 B.n611 B.n610 10.6151
R1128 B.n612 B.n611 10.6151
R1129 B.n612 B.n109 10.6151
R1130 B.n616 B.n109 10.6151
R1131 B.n617 B.n616 10.6151
R1132 B.n618 B.n617 10.6151
R1133 B.n618 B.n107 10.6151
R1134 B.n622 B.n107 10.6151
R1135 B.n623 B.n622 10.6151
R1136 B.n624 B.n623 10.6151
R1137 B.n624 B.n105 10.6151
R1138 B.n628 B.n105 10.6151
R1139 B.n629 B.n628 10.6151
R1140 B.n630 B.n629 10.6151
R1141 B.n630 B.n103 10.6151
R1142 B.n634 B.n103 10.6151
R1143 B.n635 B.n634 10.6151
R1144 B.n636 B.n635 10.6151
R1145 B.n636 B.n101 10.6151
R1146 B.n640 B.n101 10.6151
R1147 B.n641 B.n640 10.6151
R1148 B.n642 B.n641 10.6151
R1149 B.n642 B.n99 10.6151
R1150 B.n646 B.n99 10.6151
R1151 B.n647 B.n646 10.6151
R1152 B.n648 B.n647 10.6151
R1153 B.n648 B.n97 10.6151
R1154 B.n652 B.n97 10.6151
R1155 B.n653 B.n652 10.6151
R1156 B.n654 B.n653 10.6151
R1157 B.n654 B.n95 10.6151
R1158 B.n658 B.n95 10.6151
R1159 B.n659 B.n658 10.6151
R1160 B.n660 B.n659 10.6151
R1161 B.n318 B.n209 10.6151
R1162 B.n319 B.n318 10.6151
R1163 B.n320 B.n319 10.6151
R1164 B.n320 B.n207 10.6151
R1165 B.n324 B.n207 10.6151
R1166 B.n325 B.n324 10.6151
R1167 B.n326 B.n325 10.6151
R1168 B.n326 B.n205 10.6151
R1169 B.n330 B.n205 10.6151
R1170 B.n331 B.n330 10.6151
R1171 B.n332 B.n331 10.6151
R1172 B.n332 B.n203 10.6151
R1173 B.n336 B.n203 10.6151
R1174 B.n337 B.n336 10.6151
R1175 B.n338 B.n337 10.6151
R1176 B.n338 B.n201 10.6151
R1177 B.n342 B.n201 10.6151
R1178 B.n343 B.n342 10.6151
R1179 B.n344 B.n343 10.6151
R1180 B.n344 B.n199 10.6151
R1181 B.n348 B.n199 10.6151
R1182 B.n349 B.n348 10.6151
R1183 B.n350 B.n349 10.6151
R1184 B.n350 B.n197 10.6151
R1185 B.n354 B.n197 10.6151
R1186 B.n355 B.n354 10.6151
R1187 B.n356 B.n355 10.6151
R1188 B.n356 B.n195 10.6151
R1189 B.n360 B.n195 10.6151
R1190 B.n361 B.n360 10.6151
R1191 B.n362 B.n361 10.6151
R1192 B.n362 B.n193 10.6151
R1193 B.n366 B.n193 10.6151
R1194 B.n367 B.n366 10.6151
R1195 B.n368 B.n367 10.6151
R1196 B.n368 B.n191 10.6151
R1197 B.n372 B.n191 10.6151
R1198 B.n373 B.n372 10.6151
R1199 B.n374 B.n373 10.6151
R1200 B.n374 B.n189 10.6151
R1201 B.n378 B.n189 10.6151
R1202 B.n379 B.n378 10.6151
R1203 B.n380 B.n379 10.6151
R1204 B.n380 B.n187 10.6151
R1205 B.n384 B.n187 10.6151
R1206 B.n385 B.n384 10.6151
R1207 B.n386 B.n385 10.6151
R1208 B.n386 B.n185 10.6151
R1209 B.n390 B.n185 10.6151
R1210 B.n391 B.n390 10.6151
R1211 B.n392 B.n391 10.6151
R1212 B.n392 B.n183 10.6151
R1213 B.n396 B.n183 10.6151
R1214 B.n397 B.n396 10.6151
R1215 B.n399 B.n179 10.6151
R1216 B.n403 B.n179 10.6151
R1217 B.n404 B.n403 10.6151
R1218 B.n405 B.n404 10.6151
R1219 B.n405 B.n177 10.6151
R1220 B.n409 B.n177 10.6151
R1221 B.n410 B.n409 10.6151
R1222 B.n414 B.n410 10.6151
R1223 B.n418 B.n175 10.6151
R1224 B.n419 B.n418 10.6151
R1225 B.n420 B.n419 10.6151
R1226 B.n420 B.n173 10.6151
R1227 B.n424 B.n173 10.6151
R1228 B.n425 B.n424 10.6151
R1229 B.n426 B.n425 10.6151
R1230 B.n426 B.n171 10.6151
R1231 B.n430 B.n171 10.6151
R1232 B.n431 B.n430 10.6151
R1233 B.n432 B.n431 10.6151
R1234 B.n432 B.n169 10.6151
R1235 B.n436 B.n169 10.6151
R1236 B.n437 B.n436 10.6151
R1237 B.n438 B.n437 10.6151
R1238 B.n438 B.n167 10.6151
R1239 B.n442 B.n167 10.6151
R1240 B.n443 B.n442 10.6151
R1241 B.n444 B.n443 10.6151
R1242 B.n444 B.n165 10.6151
R1243 B.n448 B.n165 10.6151
R1244 B.n449 B.n448 10.6151
R1245 B.n450 B.n449 10.6151
R1246 B.n450 B.n163 10.6151
R1247 B.n454 B.n163 10.6151
R1248 B.n455 B.n454 10.6151
R1249 B.n456 B.n455 10.6151
R1250 B.n456 B.n161 10.6151
R1251 B.n460 B.n161 10.6151
R1252 B.n461 B.n460 10.6151
R1253 B.n462 B.n461 10.6151
R1254 B.n462 B.n159 10.6151
R1255 B.n466 B.n159 10.6151
R1256 B.n467 B.n466 10.6151
R1257 B.n468 B.n467 10.6151
R1258 B.n468 B.n157 10.6151
R1259 B.n472 B.n157 10.6151
R1260 B.n473 B.n472 10.6151
R1261 B.n474 B.n473 10.6151
R1262 B.n474 B.n155 10.6151
R1263 B.n478 B.n155 10.6151
R1264 B.n479 B.n478 10.6151
R1265 B.n480 B.n479 10.6151
R1266 B.n480 B.n153 10.6151
R1267 B.n484 B.n153 10.6151
R1268 B.n485 B.n484 10.6151
R1269 B.n486 B.n485 10.6151
R1270 B.n486 B.n151 10.6151
R1271 B.n490 B.n151 10.6151
R1272 B.n491 B.n490 10.6151
R1273 B.n492 B.n491 10.6151
R1274 B.n492 B.n149 10.6151
R1275 B.n496 B.n149 10.6151
R1276 B.n497 B.n496 10.6151
R1277 B.n314 B.n313 10.6151
R1278 B.n313 B.n312 10.6151
R1279 B.n312 B.n211 10.6151
R1280 B.n308 B.n211 10.6151
R1281 B.n308 B.n307 10.6151
R1282 B.n307 B.n306 10.6151
R1283 B.n306 B.n213 10.6151
R1284 B.n302 B.n213 10.6151
R1285 B.n302 B.n301 10.6151
R1286 B.n301 B.n300 10.6151
R1287 B.n300 B.n215 10.6151
R1288 B.n296 B.n215 10.6151
R1289 B.n296 B.n295 10.6151
R1290 B.n295 B.n294 10.6151
R1291 B.n294 B.n217 10.6151
R1292 B.n290 B.n217 10.6151
R1293 B.n290 B.n289 10.6151
R1294 B.n289 B.n288 10.6151
R1295 B.n288 B.n219 10.6151
R1296 B.n284 B.n219 10.6151
R1297 B.n284 B.n283 10.6151
R1298 B.n283 B.n282 10.6151
R1299 B.n282 B.n221 10.6151
R1300 B.n278 B.n221 10.6151
R1301 B.n278 B.n277 10.6151
R1302 B.n277 B.n276 10.6151
R1303 B.n276 B.n223 10.6151
R1304 B.n272 B.n223 10.6151
R1305 B.n272 B.n271 10.6151
R1306 B.n271 B.n270 10.6151
R1307 B.n270 B.n225 10.6151
R1308 B.n266 B.n225 10.6151
R1309 B.n266 B.n265 10.6151
R1310 B.n265 B.n264 10.6151
R1311 B.n264 B.n227 10.6151
R1312 B.n260 B.n227 10.6151
R1313 B.n260 B.n259 10.6151
R1314 B.n259 B.n258 10.6151
R1315 B.n258 B.n229 10.6151
R1316 B.n254 B.n229 10.6151
R1317 B.n254 B.n253 10.6151
R1318 B.n253 B.n252 10.6151
R1319 B.n252 B.n231 10.6151
R1320 B.n248 B.n231 10.6151
R1321 B.n248 B.n247 10.6151
R1322 B.n247 B.n246 10.6151
R1323 B.n246 B.n233 10.6151
R1324 B.n242 B.n233 10.6151
R1325 B.n242 B.n241 10.6151
R1326 B.n241 B.n240 10.6151
R1327 B.n240 B.n235 10.6151
R1328 B.n236 B.n235 10.6151
R1329 B.n236 B.n0 10.6151
R1330 B.n919 B.n1 10.6151
R1331 B.n919 B.n918 10.6151
R1332 B.n918 B.n917 10.6151
R1333 B.n917 B.n4 10.6151
R1334 B.n913 B.n4 10.6151
R1335 B.n913 B.n912 10.6151
R1336 B.n912 B.n911 10.6151
R1337 B.n911 B.n6 10.6151
R1338 B.n907 B.n6 10.6151
R1339 B.n907 B.n906 10.6151
R1340 B.n906 B.n905 10.6151
R1341 B.n905 B.n8 10.6151
R1342 B.n901 B.n8 10.6151
R1343 B.n901 B.n900 10.6151
R1344 B.n900 B.n899 10.6151
R1345 B.n899 B.n10 10.6151
R1346 B.n895 B.n10 10.6151
R1347 B.n895 B.n894 10.6151
R1348 B.n894 B.n893 10.6151
R1349 B.n893 B.n12 10.6151
R1350 B.n889 B.n12 10.6151
R1351 B.n889 B.n888 10.6151
R1352 B.n888 B.n887 10.6151
R1353 B.n887 B.n14 10.6151
R1354 B.n883 B.n14 10.6151
R1355 B.n883 B.n882 10.6151
R1356 B.n882 B.n881 10.6151
R1357 B.n881 B.n16 10.6151
R1358 B.n877 B.n16 10.6151
R1359 B.n877 B.n876 10.6151
R1360 B.n876 B.n875 10.6151
R1361 B.n875 B.n18 10.6151
R1362 B.n871 B.n18 10.6151
R1363 B.n871 B.n870 10.6151
R1364 B.n870 B.n869 10.6151
R1365 B.n869 B.n20 10.6151
R1366 B.n865 B.n20 10.6151
R1367 B.n865 B.n864 10.6151
R1368 B.n864 B.n863 10.6151
R1369 B.n863 B.n22 10.6151
R1370 B.n859 B.n22 10.6151
R1371 B.n859 B.n858 10.6151
R1372 B.n858 B.n857 10.6151
R1373 B.n857 B.n24 10.6151
R1374 B.n853 B.n24 10.6151
R1375 B.n853 B.n852 10.6151
R1376 B.n852 B.n851 10.6151
R1377 B.n851 B.n26 10.6151
R1378 B.n847 B.n26 10.6151
R1379 B.n847 B.n846 10.6151
R1380 B.n846 B.n845 10.6151
R1381 B.n845 B.n28 10.6151
R1382 B.n841 B.n28 10.6151
R1383 B.n757 B.n60 6.5566
R1384 B.n745 B.n744 6.5566
R1385 B.n399 B.n398 6.5566
R1386 B.n414 B.n413 6.5566
R1387 B.n60 B.n56 4.05904
R1388 B.n744 B.n743 4.05904
R1389 B.n398 B.n397 4.05904
R1390 B.n413 B.n175 4.05904
R1391 B.n923 B.n0 2.81026
R1392 B.n923 B.n1 2.81026
R1393 VN.n8 VN.t7 204.478
R1394 VN.n45 VN.t2 204.478
R1395 VN.n5 VN.t6 173.245
R1396 VN.n9 VN.t4 173.245
R1397 VN.n27 VN.t0 173.245
R1398 VN.n35 VN.t3 173.245
R1399 VN.n42 VN.t1 173.245
R1400 VN.n46 VN.t5 173.245
R1401 VN.n64 VN.t8 173.245
R1402 VN.n72 VN.t9 173.245
R1403 VN.n71 VN.n37 161.3
R1404 VN.n70 VN.n69 161.3
R1405 VN.n68 VN.n38 161.3
R1406 VN.n67 VN.n66 161.3
R1407 VN.n65 VN.n39 161.3
R1408 VN.n63 VN.n62 161.3
R1409 VN.n61 VN.n40 161.3
R1410 VN.n60 VN.n59 161.3
R1411 VN.n58 VN.n41 161.3
R1412 VN.n57 VN.n56 161.3
R1413 VN.n55 VN.n42 161.3
R1414 VN.n54 VN.n53 161.3
R1415 VN.n52 VN.n43 161.3
R1416 VN.n51 VN.n50 161.3
R1417 VN.n49 VN.n44 161.3
R1418 VN.n48 VN.n47 161.3
R1419 VN.n34 VN.n0 161.3
R1420 VN.n33 VN.n32 161.3
R1421 VN.n31 VN.n1 161.3
R1422 VN.n30 VN.n29 161.3
R1423 VN.n28 VN.n2 161.3
R1424 VN.n26 VN.n25 161.3
R1425 VN.n24 VN.n3 161.3
R1426 VN.n23 VN.n22 161.3
R1427 VN.n21 VN.n4 161.3
R1428 VN.n20 VN.n19 161.3
R1429 VN.n18 VN.n5 161.3
R1430 VN.n17 VN.n16 161.3
R1431 VN.n15 VN.n6 161.3
R1432 VN.n14 VN.n13 161.3
R1433 VN.n12 VN.n7 161.3
R1434 VN.n11 VN.n10 161.3
R1435 VN.n36 VN.n35 99.991
R1436 VN.n73 VN.n72 99.991
R1437 VN.n9 VN.n8 66.6814
R1438 VN.n46 VN.n45 66.6814
R1439 VN.n15 VN.n14 56.5193
R1440 VN.n22 VN.n21 56.5193
R1441 VN.n52 VN.n51 56.5193
R1442 VN.n59 VN.n58 56.5193
R1443 VN VN.n73 54.9338
R1444 VN.n29 VN.n1 48.7492
R1445 VN.n66 VN.n38 48.7492
R1446 VN.n33 VN.n1 32.2376
R1447 VN.n70 VN.n38 32.2376
R1448 VN.n10 VN.n7 24.4675
R1449 VN.n14 VN.n7 24.4675
R1450 VN.n16 VN.n15 24.4675
R1451 VN.n16 VN.n5 24.4675
R1452 VN.n20 VN.n5 24.4675
R1453 VN.n21 VN.n20 24.4675
R1454 VN.n22 VN.n3 24.4675
R1455 VN.n26 VN.n3 24.4675
R1456 VN.n29 VN.n28 24.4675
R1457 VN.n34 VN.n33 24.4675
R1458 VN.n51 VN.n44 24.4675
R1459 VN.n47 VN.n44 24.4675
R1460 VN.n58 VN.n57 24.4675
R1461 VN.n57 VN.n42 24.4675
R1462 VN.n53 VN.n42 24.4675
R1463 VN.n53 VN.n52 24.4675
R1464 VN.n66 VN.n65 24.4675
R1465 VN.n63 VN.n40 24.4675
R1466 VN.n59 VN.n40 24.4675
R1467 VN.n71 VN.n70 24.4675
R1468 VN.n28 VN.n27 19.0848
R1469 VN.n65 VN.n64 19.0848
R1470 VN.n35 VN.n34 10.766
R1471 VN.n72 VN.n71 10.766
R1472 VN.n48 VN.n45 9.92074
R1473 VN.n11 VN.n8 9.92074
R1474 VN.n10 VN.n9 5.38324
R1475 VN.n27 VN.n26 5.38324
R1476 VN.n47 VN.n46 5.38324
R1477 VN.n64 VN.n63 5.38324
R1478 VN.n73 VN.n37 0.278367
R1479 VN.n36 VN.n0 0.278367
R1480 VN.n69 VN.n37 0.189894
R1481 VN.n69 VN.n68 0.189894
R1482 VN.n68 VN.n67 0.189894
R1483 VN.n67 VN.n39 0.189894
R1484 VN.n62 VN.n39 0.189894
R1485 VN.n62 VN.n61 0.189894
R1486 VN.n61 VN.n60 0.189894
R1487 VN.n60 VN.n41 0.189894
R1488 VN.n56 VN.n41 0.189894
R1489 VN.n56 VN.n55 0.189894
R1490 VN.n55 VN.n54 0.189894
R1491 VN.n54 VN.n43 0.189894
R1492 VN.n50 VN.n43 0.189894
R1493 VN.n50 VN.n49 0.189894
R1494 VN.n49 VN.n48 0.189894
R1495 VN.n12 VN.n11 0.189894
R1496 VN.n13 VN.n12 0.189894
R1497 VN.n13 VN.n6 0.189894
R1498 VN.n17 VN.n6 0.189894
R1499 VN.n18 VN.n17 0.189894
R1500 VN.n19 VN.n18 0.189894
R1501 VN.n19 VN.n4 0.189894
R1502 VN.n23 VN.n4 0.189894
R1503 VN.n24 VN.n23 0.189894
R1504 VN.n25 VN.n24 0.189894
R1505 VN.n25 VN.n2 0.189894
R1506 VN.n30 VN.n2 0.189894
R1507 VN.n31 VN.n30 0.189894
R1508 VN.n32 VN.n31 0.189894
R1509 VN.n32 VN.n0 0.189894
R1510 VN VN.n36 0.153454
R1511 VDD2.n1 VDD2.t6 72.8547
R1512 VDD2.n4 VDD2.t9 70.605
R1513 VDD2.n3 VDD2.n2 70.2537
R1514 VDD2 VDD2.n7 70.2509
R1515 VDD2.n6 VDD2.n5 68.6218
R1516 VDD2.n1 VDD2.n0 68.6215
R1517 VDD2.n4 VDD2.n3 48.5321
R1518 VDD2.n6 VDD2.n4 2.2505
R1519 VDD2.n7 VDD2.t2 1.98372
R1520 VDD2.n7 VDD2.t8 1.98372
R1521 VDD2.n5 VDD2.t0 1.98372
R1522 VDD2.n5 VDD2.t4 1.98372
R1523 VDD2.n2 VDD2.t7 1.98372
R1524 VDD2.n2 VDD2.t3 1.98372
R1525 VDD2.n0 VDD2.t5 1.98372
R1526 VDD2.n0 VDD2.t1 1.98372
R1527 VDD2 VDD2.n6 0.62119
R1528 VDD2.n3 VDD2.n1 0.507654
R1529 VTAIL.n11 VTAIL.t17 53.9262
R1530 VTAIL.n17 VTAIL.t16 53.926
R1531 VTAIL.n2 VTAIL.t3 53.926
R1532 VTAIL.n16 VTAIL.t9 53.926
R1533 VTAIL.n15 VTAIL.n14 51.943
R1534 VTAIL.n13 VTAIL.n12 51.943
R1535 VTAIL.n10 VTAIL.n9 51.943
R1536 VTAIL.n8 VTAIL.n7 51.943
R1537 VTAIL.n19 VTAIL.n18 51.9427
R1538 VTAIL.n1 VTAIL.n0 51.9427
R1539 VTAIL.n4 VTAIL.n3 51.9427
R1540 VTAIL.n6 VTAIL.n5 51.9427
R1541 VTAIL.n8 VTAIL.n6 30.9962
R1542 VTAIL.n17 VTAIL.n16 28.7462
R1543 VTAIL.n10 VTAIL.n8 2.2505
R1544 VTAIL.n11 VTAIL.n10 2.2505
R1545 VTAIL.n15 VTAIL.n13 2.2505
R1546 VTAIL.n16 VTAIL.n15 2.2505
R1547 VTAIL.n6 VTAIL.n4 2.2505
R1548 VTAIL.n4 VTAIL.n2 2.2505
R1549 VTAIL.n19 VTAIL.n17 2.2505
R1550 VTAIL.n18 VTAIL.t13 1.98372
R1551 VTAIL.n18 VTAIL.t19 1.98372
R1552 VTAIL.n0 VTAIL.t12 1.98372
R1553 VTAIL.n0 VTAIL.t15 1.98372
R1554 VTAIL.n3 VTAIL.t0 1.98372
R1555 VTAIL.n3 VTAIL.t8 1.98372
R1556 VTAIL.n5 VTAIL.t6 1.98372
R1557 VTAIL.n5 VTAIL.t7 1.98372
R1558 VTAIL.n14 VTAIL.t2 1.98372
R1559 VTAIL.n14 VTAIL.t4 1.98372
R1560 VTAIL.n12 VTAIL.t1 1.98372
R1561 VTAIL.n12 VTAIL.t5 1.98372
R1562 VTAIL.n9 VTAIL.t18 1.98372
R1563 VTAIL.n9 VTAIL.t14 1.98372
R1564 VTAIL.n7 VTAIL.t10 1.98372
R1565 VTAIL.n7 VTAIL.t11 1.98372
R1566 VTAIL VTAIL.n1 1.74619
R1567 VTAIL.n13 VTAIL.n11 1.59533
R1568 VTAIL.n2 VTAIL.n1 1.59533
R1569 VTAIL VTAIL.n19 0.50481
R1570 VP.n19 VP.t9 204.478
R1571 VP.n5 VP.t5 173.245
R1572 VP.n49 VP.t4 173.245
R1573 VP.n57 VP.t2 173.245
R1574 VP.n75 VP.t1 173.245
R1575 VP.n83 VP.t8 173.245
R1576 VP.n16 VP.t6 173.245
R1577 VP.n46 VP.t0 173.245
R1578 VP.n38 VP.t7 173.245
R1579 VP.n20 VP.t3 173.245
R1580 VP.n22 VP.n21 161.3
R1581 VP.n23 VP.n18 161.3
R1582 VP.n25 VP.n24 161.3
R1583 VP.n26 VP.n17 161.3
R1584 VP.n28 VP.n27 161.3
R1585 VP.n29 VP.n16 161.3
R1586 VP.n31 VP.n30 161.3
R1587 VP.n32 VP.n15 161.3
R1588 VP.n34 VP.n33 161.3
R1589 VP.n35 VP.n14 161.3
R1590 VP.n37 VP.n36 161.3
R1591 VP.n39 VP.n13 161.3
R1592 VP.n41 VP.n40 161.3
R1593 VP.n42 VP.n12 161.3
R1594 VP.n44 VP.n43 161.3
R1595 VP.n45 VP.n11 161.3
R1596 VP.n82 VP.n0 161.3
R1597 VP.n81 VP.n80 161.3
R1598 VP.n79 VP.n1 161.3
R1599 VP.n78 VP.n77 161.3
R1600 VP.n76 VP.n2 161.3
R1601 VP.n74 VP.n73 161.3
R1602 VP.n72 VP.n3 161.3
R1603 VP.n71 VP.n70 161.3
R1604 VP.n69 VP.n4 161.3
R1605 VP.n68 VP.n67 161.3
R1606 VP.n66 VP.n5 161.3
R1607 VP.n65 VP.n64 161.3
R1608 VP.n63 VP.n6 161.3
R1609 VP.n62 VP.n61 161.3
R1610 VP.n60 VP.n7 161.3
R1611 VP.n59 VP.n58 161.3
R1612 VP.n56 VP.n8 161.3
R1613 VP.n55 VP.n54 161.3
R1614 VP.n53 VP.n9 161.3
R1615 VP.n52 VP.n51 161.3
R1616 VP.n50 VP.n10 161.3
R1617 VP.n49 VP.n48 99.991
R1618 VP.n84 VP.n83 99.991
R1619 VP.n47 VP.n46 99.991
R1620 VP.n20 VP.n19 66.6814
R1621 VP.n63 VP.n62 56.5193
R1622 VP.n70 VP.n69 56.5193
R1623 VP.n33 VP.n32 56.5193
R1624 VP.n26 VP.n25 56.5193
R1625 VP.n48 VP.n47 54.6549
R1626 VP.n55 VP.n9 48.7492
R1627 VP.n77 VP.n1 48.7492
R1628 VP.n40 VP.n12 48.7492
R1629 VP.n51 VP.n9 32.2376
R1630 VP.n81 VP.n1 32.2376
R1631 VP.n44 VP.n12 32.2376
R1632 VP.n51 VP.n50 24.4675
R1633 VP.n56 VP.n55 24.4675
R1634 VP.n58 VP.n7 24.4675
R1635 VP.n62 VP.n7 24.4675
R1636 VP.n64 VP.n63 24.4675
R1637 VP.n64 VP.n5 24.4675
R1638 VP.n68 VP.n5 24.4675
R1639 VP.n69 VP.n68 24.4675
R1640 VP.n70 VP.n3 24.4675
R1641 VP.n74 VP.n3 24.4675
R1642 VP.n77 VP.n76 24.4675
R1643 VP.n82 VP.n81 24.4675
R1644 VP.n45 VP.n44 24.4675
R1645 VP.n33 VP.n14 24.4675
R1646 VP.n37 VP.n14 24.4675
R1647 VP.n40 VP.n39 24.4675
R1648 VP.n27 VP.n26 24.4675
R1649 VP.n27 VP.n16 24.4675
R1650 VP.n31 VP.n16 24.4675
R1651 VP.n32 VP.n31 24.4675
R1652 VP.n21 VP.n18 24.4675
R1653 VP.n25 VP.n18 24.4675
R1654 VP.n57 VP.n56 19.0848
R1655 VP.n76 VP.n75 19.0848
R1656 VP.n39 VP.n38 19.0848
R1657 VP.n50 VP.n49 10.766
R1658 VP.n83 VP.n82 10.766
R1659 VP.n46 VP.n45 10.766
R1660 VP.n22 VP.n19 9.92074
R1661 VP.n58 VP.n57 5.38324
R1662 VP.n75 VP.n74 5.38324
R1663 VP.n38 VP.n37 5.38324
R1664 VP.n21 VP.n20 5.38324
R1665 VP.n47 VP.n11 0.278367
R1666 VP.n48 VP.n10 0.278367
R1667 VP.n84 VP.n0 0.278367
R1668 VP.n23 VP.n22 0.189894
R1669 VP.n24 VP.n23 0.189894
R1670 VP.n24 VP.n17 0.189894
R1671 VP.n28 VP.n17 0.189894
R1672 VP.n29 VP.n28 0.189894
R1673 VP.n30 VP.n29 0.189894
R1674 VP.n30 VP.n15 0.189894
R1675 VP.n34 VP.n15 0.189894
R1676 VP.n35 VP.n34 0.189894
R1677 VP.n36 VP.n35 0.189894
R1678 VP.n36 VP.n13 0.189894
R1679 VP.n41 VP.n13 0.189894
R1680 VP.n42 VP.n41 0.189894
R1681 VP.n43 VP.n42 0.189894
R1682 VP.n43 VP.n11 0.189894
R1683 VP.n52 VP.n10 0.189894
R1684 VP.n53 VP.n52 0.189894
R1685 VP.n54 VP.n53 0.189894
R1686 VP.n54 VP.n8 0.189894
R1687 VP.n59 VP.n8 0.189894
R1688 VP.n60 VP.n59 0.189894
R1689 VP.n61 VP.n60 0.189894
R1690 VP.n61 VP.n6 0.189894
R1691 VP.n65 VP.n6 0.189894
R1692 VP.n66 VP.n65 0.189894
R1693 VP.n67 VP.n66 0.189894
R1694 VP.n67 VP.n4 0.189894
R1695 VP.n71 VP.n4 0.189894
R1696 VP.n72 VP.n71 0.189894
R1697 VP.n73 VP.n72 0.189894
R1698 VP.n73 VP.n2 0.189894
R1699 VP.n78 VP.n2 0.189894
R1700 VP.n79 VP.n78 0.189894
R1701 VP.n80 VP.n79 0.189894
R1702 VP.n80 VP.n0 0.189894
R1703 VP VP.n84 0.153454
R1704 VDD1.n1 VDD1.t0 72.855
R1705 VDD1.n3 VDD1.t5 72.8547
R1706 VDD1.n5 VDD1.n4 70.2537
R1707 VDD1.n1 VDD1.n0 68.6218
R1708 VDD1.n7 VDD1.n6 68.6216
R1709 VDD1.n3 VDD1.n2 68.6215
R1710 VDD1.n7 VDD1.n5 50.2401
R1711 VDD1.n6 VDD1.t2 1.98372
R1712 VDD1.n6 VDD1.t9 1.98372
R1713 VDD1.n0 VDD1.t6 1.98372
R1714 VDD1.n0 VDD1.t3 1.98372
R1715 VDD1.n4 VDD1.t8 1.98372
R1716 VDD1.n4 VDD1.t1 1.98372
R1717 VDD1.n2 VDD1.t7 1.98372
R1718 VDD1.n2 VDD1.t4 1.98372
R1719 VDD1 VDD1.n7 1.62981
R1720 VDD1 VDD1.n1 0.62119
R1721 VDD1.n5 VDD1.n3 0.507654
C0 VP VDD1 14.3703f
C1 VDD2 VDD1 1.96678f
C2 w_n4102_n4246# VN 8.765429f
C3 B VP 2.14813f
C4 B VDD2 2.80475f
C5 w_n4102_n4246# VDD1 2.97442f
C6 B w_n4102_n4246# 11.239599f
C7 VP VTAIL 14.3161f
C8 VTAIL VDD2 12.583599f
C9 VDD1 VN 0.152632f
C10 B VN 1.25351f
C11 w_n4102_n4246# VTAIL 3.78892f
C12 VP VDD2 0.543159f
C13 B VDD1 2.6993f
C14 w_n4102_n4246# VP 9.29851f
C15 w_n4102_n4246# VDD2 3.10143f
C16 VTAIL VN 14.301701f
C17 VTAIL VDD1 12.536301f
C18 VP VN 8.74304f
C19 VDD2 VN 13.9845f
C20 B VTAIL 4.55414f
C21 VDD2 VSUBS 2.10485f
C22 VDD1 VSUBS 1.936082f
C23 VTAIL VSUBS 1.374031f
C24 VN VSUBS 7.334899f
C25 VP VSUBS 3.989917f
C26 B VSUBS 5.339225f
C27 w_n4102_n4246# VSUBS 0.213288p
C28 VDD1.t0 VSUBS 3.72761f
C29 VDD1.t6 VSUBS 0.347811f
C30 VDD1.t3 VSUBS 0.347811f
C31 VDD1.n0 VSUBS 2.85034f
C32 VDD1.n1 VSUBS 1.58015f
C33 VDD1.t5 VSUBS 3.72761f
C34 VDD1.t7 VSUBS 0.347811f
C35 VDD1.t4 VSUBS 0.347811f
C36 VDD1.n2 VSUBS 2.85034f
C37 VDD1.n3 VSUBS 1.57156f
C38 VDD1.t8 VSUBS 0.347811f
C39 VDD1.t1 VSUBS 0.347811f
C40 VDD1.n4 VSUBS 2.87066f
C41 VDD1.n5 VSUBS 3.66338f
C42 VDD1.t2 VSUBS 0.347811f
C43 VDD1.t9 VSUBS 0.347811f
C44 VDD1.n6 VSUBS 2.85033f
C45 VDD1.n7 VSUBS 3.93085f
C46 VP.n0 VSUBS 0.039336f
C47 VP.t8 VSUBS 3.06106f
C48 VP.n1 VSUBS 0.02701f
C49 VP.n2 VSUBS 0.029836f
C50 VP.t1 VSUBS 3.06106f
C51 VP.n3 VSUBS 0.055607f
C52 VP.n4 VSUBS 0.029836f
C53 VP.t5 VSUBS 3.06106f
C54 VP.n5 VSUBS 1.09714f
C55 VP.n6 VSUBS 0.029836f
C56 VP.n7 VSUBS 0.055607f
C57 VP.n8 VSUBS 0.029836f
C58 VP.t2 VSUBS 3.06106f
C59 VP.n9 VSUBS 0.02701f
C60 VP.n10 VSUBS 0.039336f
C61 VP.t4 VSUBS 3.06106f
C62 VP.n11 VSUBS 0.039336f
C63 VP.t0 VSUBS 3.06106f
C64 VP.n12 VSUBS 0.02701f
C65 VP.n13 VSUBS 0.029836f
C66 VP.t7 VSUBS 3.06106f
C67 VP.n14 VSUBS 0.055607f
C68 VP.n15 VSUBS 0.029836f
C69 VP.t6 VSUBS 3.06106f
C70 VP.n16 VSUBS 1.09714f
C71 VP.n17 VSUBS 0.029836f
C72 VP.n18 VSUBS 0.055607f
C73 VP.t9 VSUBS 3.24892f
C74 VP.n19 VSUBS 1.13933f
C75 VP.t3 VSUBS 3.06106f
C76 VP.n20 VSUBS 1.14118f
C77 VP.n21 VSUBS 0.034193f
C78 VP.n22 VSUBS 0.256074f
C79 VP.n23 VSUBS 0.029836f
C80 VP.n24 VSUBS 0.029836f
C81 VP.n25 VSUBS 0.038985f
C82 VP.n26 VSUBS 0.048131f
C83 VP.n27 VSUBS 0.055607f
C84 VP.n28 VSUBS 0.029836f
C85 VP.n29 VSUBS 0.029836f
C86 VP.n30 VSUBS 0.029836f
C87 VP.n31 VSUBS 0.055607f
C88 VP.n32 VSUBS 0.048131f
C89 VP.n33 VSUBS 0.038985f
C90 VP.n34 VSUBS 0.029836f
C91 VP.n35 VSUBS 0.029836f
C92 VP.n36 VSUBS 0.029836f
C93 VP.n37 VSUBS 0.034193f
C94 VP.n38 VSUBS 1.06899f
C95 VP.n39 VSUBS 0.049567f
C96 VP.n40 VSUBS 0.055607f
C97 VP.n41 VSUBS 0.029836f
C98 VP.n42 VSUBS 0.029836f
C99 VP.n43 VSUBS 0.029836f
C100 VP.n44 VSUBS 0.060106f
C101 VP.n45 VSUBS 0.040233f
C102 VP.n46 VSUBS 1.15727f
C103 VP.n47 VSUBS 1.88244f
C104 VP.n48 VSUBS 1.90206f
C105 VP.n49 VSUBS 1.15727f
C106 VP.n50 VSUBS 0.040233f
C107 VP.n51 VSUBS 0.060106f
C108 VP.n52 VSUBS 0.029836f
C109 VP.n53 VSUBS 0.029836f
C110 VP.n54 VSUBS 0.029836f
C111 VP.n55 VSUBS 0.055607f
C112 VP.n56 VSUBS 0.049567f
C113 VP.n57 VSUBS 1.06899f
C114 VP.n58 VSUBS 0.034193f
C115 VP.n59 VSUBS 0.029836f
C116 VP.n60 VSUBS 0.029836f
C117 VP.n61 VSUBS 0.029836f
C118 VP.n62 VSUBS 0.038985f
C119 VP.n63 VSUBS 0.048131f
C120 VP.n64 VSUBS 0.055607f
C121 VP.n65 VSUBS 0.029836f
C122 VP.n66 VSUBS 0.029836f
C123 VP.n67 VSUBS 0.029836f
C124 VP.n68 VSUBS 0.055607f
C125 VP.n69 VSUBS 0.048131f
C126 VP.n70 VSUBS 0.038985f
C127 VP.n71 VSUBS 0.029836f
C128 VP.n72 VSUBS 0.029836f
C129 VP.n73 VSUBS 0.029836f
C130 VP.n74 VSUBS 0.034193f
C131 VP.n75 VSUBS 1.06899f
C132 VP.n76 VSUBS 0.049567f
C133 VP.n77 VSUBS 0.055607f
C134 VP.n78 VSUBS 0.029836f
C135 VP.n79 VSUBS 0.029836f
C136 VP.n80 VSUBS 0.029836f
C137 VP.n81 VSUBS 0.060106f
C138 VP.n82 VSUBS 0.040233f
C139 VP.n83 VSUBS 1.15727f
C140 VP.n84 VSUBS 0.045065f
C141 VTAIL.t12 VSUBS 0.356187f
C142 VTAIL.t15 VSUBS 0.356187f
C143 VTAIL.n0 VSUBS 2.74721f
C144 VTAIL.n1 VSUBS 0.970575f
C145 VTAIL.t3 VSUBS 3.59497f
C146 VTAIL.n2 VSUBS 1.13892f
C147 VTAIL.t0 VSUBS 0.356187f
C148 VTAIL.t8 VSUBS 0.356187f
C149 VTAIL.n3 VSUBS 2.74721f
C150 VTAIL.n4 VSUBS 1.07332f
C151 VTAIL.t6 VSUBS 0.356187f
C152 VTAIL.t7 VSUBS 0.356187f
C153 VTAIL.n5 VSUBS 2.74721f
C154 VTAIL.n6 VSUBS 2.89832f
C155 VTAIL.t10 VSUBS 0.356187f
C156 VTAIL.t11 VSUBS 0.356187f
C157 VTAIL.n7 VSUBS 2.74721f
C158 VTAIL.n8 VSUBS 2.89831f
C159 VTAIL.t18 VSUBS 0.356187f
C160 VTAIL.t14 VSUBS 0.356187f
C161 VTAIL.n9 VSUBS 2.74721f
C162 VTAIL.n10 VSUBS 1.07332f
C163 VTAIL.t17 VSUBS 3.59497f
C164 VTAIL.n11 VSUBS 1.13892f
C165 VTAIL.t1 VSUBS 0.356187f
C166 VTAIL.t5 VSUBS 0.356187f
C167 VTAIL.n12 VSUBS 2.74721f
C168 VTAIL.n13 VSUBS 1.01526f
C169 VTAIL.t2 VSUBS 0.356187f
C170 VTAIL.t4 VSUBS 0.356187f
C171 VTAIL.n14 VSUBS 2.74721f
C172 VTAIL.n15 VSUBS 1.07332f
C173 VTAIL.t9 VSUBS 3.59496f
C174 VTAIL.n16 VSUBS 2.8226f
C175 VTAIL.t16 VSUBS 3.59497f
C176 VTAIL.n17 VSUBS 2.8226f
C177 VTAIL.t13 VSUBS 0.356187f
C178 VTAIL.t19 VSUBS 0.356187f
C179 VTAIL.n18 VSUBS 2.74721f
C180 VTAIL.n19 VSUBS 0.918629f
C181 VDD2.t6 VSUBS 3.72751f
C182 VDD2.t5 VSUBS 0.347802f
C183 VDD2.t1 VSUBS 0.347802f
C184 VDD2.n0 VSUBS 2.85027f
C185 VDD2.n1 VSUBS 1.57152f
C186 VDD2.t7 VSUBS 0.347802f
C187 VDD2.t3 VSUBS 0.347802f
C188 VDD2.n2 VSUBS 2.87059f
C189 VDD2.n3 VSUBS 3.53538f
C190 VDD2.t9 VSUBS 3.70189f
C191 VDD2.n4 VSUBS 3.91542f
C192 VDD2.t0 VSUBS 0.347802f
C193 VDD2.t4 VSUBS 0.347802f
C194 VDD2.n5 VSUBS 2.85027f
C195 VDD2.n6 VSUBS 0.775846f
C196 VDD2.t2 VSUBS 0.347802f
C197 VDD2.t8 VSUBS 0.347802f
C198 VDD2.n7 VSUBS 2.87053f
C199 VN.n0 VSUBS 0.036886f
C200 VN.t3 VSUBS 2.87041f
C201 VN.n1 VSUBS 0.025327f
C202 VN.n2 VSUBS 0.027978f
C203 VN.t0 VSUBS 2.87041f
C204 VN.n3 VSUBS 0.052144f
C205 VN.n4 VSUBS 0.027978f
C206 VN.t6 VSUBS 2.87041f
C207 VN.n5 VSUBS 1.02881f
C208 VN.n6 VSUBS 0.027978f
C209 VN.n7 VSUBS 0.052144f
C210 VN.t7 VSUBS 3.04657f
C211 VN.n8 VSUBS 1.06837f
C212 VN.t4 VSUBS 2.87041f
C213 VN.n9 VSUBS 1.07011f
C214 VN.n10 VSUBS 0.032064f
C215 VN.n11 VSUBS 0.240125f
C216 VN.n12 VSUBS 0.027978f
C217 VN.n13 VSUBS 0.027978f
C218 VN.n14 VSUBS 0.036557f
C219 VN.n15 VSUBS 0.045133f
C220 VN.n16 VSUBS 0.052144f
C221 VN.n17 VSUBS 0.027978f
C222 VN.n18 VSUBS 0.027978f
C223 VN.n19 VSUBS 0.027978f
C224 VN.n20 VSUBS 0.052144f
C225 VN.n21 VSUBS 0.045133f
C226 VN.n22 VSUBS 0.036557f
C227 VN.n23 VSUBS 0.027978f
C228 VN.n24 VSUBS 0.027978f
C229 VN.n25 VSUBS 0.027978f
C230 VN.n26 VSUBS 0.032064f
C231 VN.n27 VSUBS 1.00241f
C232 VN.n28 VSUBS 0.04648f
C233 VN.n29 VSUBS 0.052144f
C234 VN.n30 VSUBS 0.027978f
C235 VN.n31 VSUBS 0.027978f
C236 VN.n32 VSUBS 0.027978f
C237 VN.n33 VSUBS 0.056363f
C238 VN.n34 VSUBS 0.037727f
C239 VN.n35 VSUBS 1.08519f
C240 VN.n36 VSUBS 0.042258f
C241 VN.n37 VSUBS 0.036886f
C242 VN.t9 VSUBS 2.87041f
C243 VN.n38 VSUBS 0.025327f
C244 VN.n39 VSUBS 0.027978f
C245 VN.t8 VSUBS 2.87041f
C246 VN.n40 VSUBS 0.052144f
C247 VN.n41 VSUBS 0.027978f
C248 VN.t1 VSUBS 2.87041f
C249 VN.n42 VSUBS 1.02881f
C250 VN.n43 VSUBS 0.027978f
C251 VN.n44 VSUBS 0.052144f
C252 VN.t2 VSUBS 3.04657f
C253 VN.n45 VSUBS 1.06837f
C254 VN.t5 VSUBS 2.87041f
C255 VN.n46 VSUBS 1.07011f
C256 VN.n47 VSUBS 0.032064f
C257 VN.n48 VSUBS 0.240125f
C258 VN.n49 VSUBS 0.027978f
C259 VN.n50 VSUBS 0.027978f
C260 VN.n51 VSUBS 0.036557f
C261 VN.n52 VSUBS 0.045133f
C262 VN.n53 VSUBS 0.052144f
C263 VN.n54 VSUBS 0.027978f
C264 VN.n55 VSUBS 0.027978f
C265 VN.n56 VSUBS 0.027978f
C266 VN.n57 VSUBS 0.052144f
C267 VN.n58 VSUBS 0.045133f
C268 VN.n59 VSUBS 0.036557f
C269 VN.n60 VSUBS 0.027978f
C270 VN.n61 VSUBS 0.027978f
C271 VN.n62 VSUBS 0.027978f
C272 VN.n63 VSUBS 0.032064f
C273 VN.n64 VSUBS 1.00241f
C274 VN.n65 VSUBS 0.04648f
C275 VN.n66 VSUBS 0.052144f
C276 VN.n67 VSUBS 0.027978f
C277 VN.n68 VSUBS 0.027978f
C278 VN.n69 VSUBS 0.027978f
C279 VN.n70 VSUBS 0.056363f
C280 VN.n71 VSUBS 0.037727f
C281 VN.n72 VSUBS 1.08519f
C282 VN.n73 VSUBS 1.78003f
C283 B.n0 VSUBS 0.005414f
C284 B.n1 VSUBS 0.005414f
C285 B.n2 VSUBS 0.008562f
C286 B.n3 VSUBS 0.008562f
C287 B.n4 VSUBS 0.008562f
C288 B.n5 VSUBS 0.008562f
C289 B.n6 VSUBS 0.008562f
C290 B.n7 VSUBS 0.008562f
C291 B.n8 VSUBS 0.008562f
C292 B.n9 VSUBS 0.008562f
C293 B.n10 VSUBS 0.008562f
C294 B.n11 VSUBS 0.008562f
C295 B.n12 VSUBS 0.008562f
C296 B.n13 VSUBS 0.008562f
C297 B.n14 VSUBS 0.008562f
C298 B.n15 VSUBS 0.008562f
C299 B.n16 VSUBS 0.008562f
C300 B.n17 VSUBS 0.008562f
C301 B.n18 VSUBS 0.008562f
C302 B.n19 VSUBS 0.008562f
C303 B.n20 VSUBS 0.008562f
C304 B.n21 VSUBS 0.008562f
C305 B.n22 VSUBS 0.008562f
C306 B.n23 VSUBS 0.008562f
C307 B.n24 VSUBS 0.008562f
C308 B.n25 VSUBS 0.008562f
C309 B.n26 VSUBS 0.008562f
C310 B.n27 VSUBS 0.008562f
C311 B.n28 VSUBS 0.008562f
C312 B.n29 VSUBS 0.020678f
C313 B.n30 VSUBS 0.008562f
C314 B.n31 VSUBS 0.008562f
C315 B.n32 VSUBS 0.008562f
C316 B.n33 VSUBS 0.008562f
C317 B.n34 VSUBS 0.008562f
C318 B.n35 VSUBS 0.008562f
C319 B.n36 VSUBS 0.008562f
C320 B.n37 VSUBS 0.008562f
C321 B.n38 VSUBS 0.008562f
C322 B.n39 VSUBS 0.008562f
C323 B.n40 VSUBS 0.008562f
C324 B.n41 VSUBS 0.008562f
C325 B.n42 VSUBS 0.008562f
C326 B.n43 VSUBS 0.008562f
C327 B.n44 VSUBS 0.008562f
C328 B.n45 VSUBS 0.008562f
C329 B.n46 VSUBS 0.008562f
C330 B.n47 VSUBS 0.008562f
C331 B.n48 VSUBS 0.008562f
C332 B.n49 VSUBS 0.008562f
C333 B.n50 VSUBS 0.008562f
C334 B.n51 VSUBS 0.008562f
C335 B.n52 VSUBS 0.008562f
C336 B.n53 VSUBS 0.008562f
C337 B.n54 VSUBS 0.008562f
C338 B.n55 VSUBS 0.008562f
C339 B.n56 VSUBS 0.005918f
C340 B.n57 VSUBS 0.008562f
C341 B.t11 VSUBS 0.672094f
C342 B.t10 VSUBS 0.69585f
C343 B.t9 VSUBS 2.02042f
C344 B.n58 VSUBS 0.358367f
C345 B.n59 VSUBS 0.086521f
C346 B.n60 VSUBS 0.019836f
C347 B.n61 VSUBS 0.008562f
C348 B.n62 VSUBS 0.008562f
C349 B.n63 VSUBS 0.008562f
C350 B.n64 VSUBS 0.008562f
C351 B.t8 VSUBS 0.672072f
C352 B.t7 VSUBS 0.695832f
C353 B.t6 VSUBS 2.02042f
C354 B.n65 VSUBS 0.358385f
C355 B.n66 VSUBS 0.086543f
C356 B.n67 VSUBS 0.008562f
C357 B.n68 VSUBS 0.008562f
C358 B.n69 VSUBS 0.008562f
C359 B.n70 VSUBS 0.008562f
C360 B.n71 VSUBS 0.008562f
C361 B.n72 VSUBS 0.008562f
C362 B.n73 VSUBS 0.008562f
C363 B.n74 VSUBS 0.008562f
C364 B.n75 VSUBS 0.008562f
C365 B.n76 VSUBS 0.008562f
C366 B.n77 VSUBS 0.008562f
C367 B.n78 VSUBS 0.008562f
C368 B.n79 VSUBS 0.008562f
C369 B.n80 VSUBS 0.008562f
C370 B.n81 VSUBS 0.008562f
C371 B.n82 VSUBS 0.008562f
C372 B.n83 VSUBS 0.008562f
C373 B.n84 VSUBS 0.008562f
C374 B.n85 VSUBS 0.008562f
C375 B.n86 VSUBS 0.008562f
C376 B.n87 VSUBS 0.008562f
C377 B.n88 VSUBS 0.008562f
C378 B.n89 VSUBS 0.008562f
C379 B.n90 VSUBS 0.008562f
C380 B.n91 VSUBS 0.008562f
C381 B.n92 VSUBS 0.008562f
C382 B.n93 VSUBS 0.019656f
C383 B.n94 VSUBS 0.008562f
C384 B.n95 VSUBS 0.008562f
C385 B.n96 VSUBS 0.008562f
C386 B.n97 VSUBS 0.008562f
C387 B.n98 VSUBS 0.008562f
C388 B.n99 VSUBS 0.008562f
C389 B.n100 VSUBS 0.008562f
C390 B.n101 VSUBS 0.008562f
C391 B.n102 VSUBS 0.008562f
C392 B.n103 VSUBS 0.008562f
C393 B.n104 VSUBS 0.008562f
C394 B.n105 VSUBS 0.008562f
C395 B.n106 VSUBS 0.008562f
C396 B.n107 VSUBS 0.008562f
C397 B.n108 VSUBS 0.008562f
C398 B.n109 VSUBS 0.008562f
C399 B.n110 VSUBS 0.008562f
C400 B.n111 VSUBS 0.008562f
C401 B.n112 VSUBS 0.008562f
C402 B.n113 VSUBS 0.008562f
C403 B.n114 VSUBS 0.008562f
C404 B.n115 VSUBS 0.008562f
C405 B.n116 VSUBS 0.008562f
C406 B.n117 VSUBS 0.008562f
C407 B.n118 VSUBS 0.008562f
C408 B.n119 VSUBS 0.008562f
C409 B.n120 VSUBS 0.008562f
C410 B.n121 VSUBS 0.008562f
C411 B.n122 VSUBS 0.008562f
C412 B.n123 VSUBS 0.008562f
C413 B.n124 VSUBS 0.008562f
C414 B.n125 VSUBS 0.008562f
C415 B.n126 VSUBS 0.008562f
C416 B.n127 VSUBS 0.008562f
C417 B.n128 VSUBS 0.008562f
C418 B.n129 VSUBS 0.008562f
C419 B.n130 VSUBS 0.008562f
C420 B.n131 VSUBS 0.008562f
C421 B.n132 VSUBS 0.008562f
C422 B.n133 VSUBS 0.008562f
C423 B.n134 VSUBS 0.008562f
C424 B.n135 VSUBS 0.008562f
C425 B.n136 VSUBS 0.008562f
C426 B.n137 VSUBS 0.008562f
C427 B.n138 VSUBS 0.008562f
C428 B.n139 VSUBS 0.008562f
C429 B.n140 VSUBS 0.008562f
C430 B.n141 VSUBS 0.008562f
C431 B.n142 VSUBS 0.008562f
C432 B.n143 VSUBS 0.008562f
C433 B.n144 VSUBS 0.008562f
C434 B.n145 VSUBS 0.008562f
C435 B.n146 VSUBS 0.008562f
C436 B.n147 VSUBS 0.008562f
C437 B.n148 VSUBS 0.020678f
C438 B.n149 VSUBS 0.008562f
C439 B.n150 VSUBS 0.008562f
C440 B.n151 VSUBS 0.008562f
C441 B.n152 VSUBS 0.008562f
C442 B.n153 VSUBS 0.008562f
C443 B.n154 VSUBS 0.008562f
C444 B.n155 VSUBS 0.008562f
C445 B.n156 VSUBS 0.008562f
C446 B.n157 VSUBS 0.008562f
C447 B.n158 VSUBS 0.008562f
C448 B.n159 VSUBS 0.008562f
C449 B.n160 VSUBS 0.008562f
C450 B.n161 VSUBS 0.008562f
C451 B.n162 VSUBS 0.008562f
C452 B.n163 VSUBS 0.008562f
C453 B.n164 VSUBS 0.008562f
C454 B.n165 VSUBS 0.008562f
C455 B.n166 VSUBS 0.008562f
C456 B.n167 VSUBS 0.008562f
C457 B.n168 VSUBS 0.008562f
C458 B.n169 VSUBS 0.008562f
C459 B.n170 VSUBS 0.008562f
C460 B.n171 VSUBS 0.008562f
C461 B.n172 VSUBS 0.008562f
C462 B.n173 VSUBS 0.008562f
C463 B.n174 VSUBS 0.008562f
C464 B.n175 VSUBS 0.005918f
C465 B.n176 VSUBS 0.008562f
C466 B.n177 VSUBS 0.008562f
C467 B.n178 VSUBS 0.008562f
C468 B.n179 VSUBS 0.008562f
C469 B.n180 VSUBS 0.008562f
C470 B.t4 VSUBS 0.672094f
C471 B.t5 VSUBS 0.69585f
C472 B.t3 VSUBS 2.02042f
C473 B.n181 VSUBS 0.358367f
C474 B.n182 VSUBS 0.086521f
C475 B.n183 VSUBS 0.008562f
C476 B.n184 VSUBS 0.008562f
C477 B.n185 VSUBS 0.008562f
C478 B.n186 VSUBS 0.008562f
C479 B.n187 VSUBS 0.008562f
C480 B.n188 VSUBS 0.008562f
C481 B.n189 VSUBS 0.008562f
C482 B.n190 VSUBS 0.008562f
C483 B.n191 VSUBS 0.008562f
C484 B.n192 VSUBS 0.008562f
C485 B.n193 VSUBS 0.008562f
C486 B.n194 VSUBS 0.008562f
C487 B.n195 VSUBS 0.008562f
C488 B.n196 VSUBS 0.008562f
C489 B.n197 VSUBS 0.008562f
C490 B.n198 VSUBS 0.008562f
C491 B.n199 VSUBS 0.008562f
C492 B.n200 VSUBS 0.008562f
C493 B.n201 VSUBS 0.008562f
C494 B.n202 VSUBS 0.008562f
C495 B.n203 VSUBS 0.008562f
C496 B.n204 VSUBS 0.008562f
C497 B.n205 VSUBS 0.008562f
C498 B.n206 VSUBS 0.008562f
C499 B.n207 VSUBS 0.008562f
C500 B.n208 VSUBS 0.008562f
C501 B.n209 VSUBS 0.020678f
C502 B.n210 VSUBS 0.008562f
C503 B.n211 VSUBS 0.008562f
C504 B.n212 VSUBS 0.008562f
C505 B.n213 VSUBS 0.008562f
C506 B.n214 VSUBS 0.008562f
C507 B.n215 VSUBS 0.008562f
C508 B.n216 VSUBS 0.008562f
C509 B.n217 VSUBS 0.008562f
C510 B.n218 VSUBS 0.008562f
C511 B.n219 VSUBS 0.008562f
C512 B.n220 VSUBS 0.008562f
C513 B.n221 VSUBS 0.008562f
C514 B.n222 VSUBS 0.008562f
C515 B.n223 VSUBS 0.008562f
C516 B.n224 VSUBS 0.008562f
C517 B.n225 VSUBS 0.008562f
C518 B.n226 VSUBS 0.008562f
C519 B.n227 VSUBS 0.008562f
C520 B.n228 VSUBS 0.008562f
C521 B.n229 VSUBS 0.008562f
C522 B.n230 VSUBS 0.008562f
C523 B.n231 VSUBS 0.008562f
C524 B.n232 VSUBS 0.008562f
C525 B.n233 VSUBS 0.008562f
C526 B.n234 VSUBS 0.008562f
C527 B.n235 VSUBS 0.008562f
C528 B.n236 VSUBS 0.008562f
C529 B.n237 VSUBS 0.008562f
C530 B.n238 VSUBS 0.008562f
C531 B.n239 VSUBS 0.008562f
C532 B.n240 VSUBS 0.008562f
C533 B.n241 VSUBS 0.008562f
C534 B.n242 VSUBS 0.008562f
C535 B.n243 VSUBS 0.008562f
C536 B.n244 VSUBS 0.008562f
C537 B.n245 VSUBS 0.008562f
C538 B.n246 VSUBS 0.008562f
C539 B.n247 VSUBS 0.008562f
C540 B.n248 VSUBS 0.008562f
C541 B.n249 VSUBS 0.008562f
C542 B.n250 VSUBS 0.008562f
C543 B.n251 VSUBS 0.008562f
C544 B.n252 VSUBS 0.008562f
C545 B.n253 VSUBS 0.008562f
C546 B.n254 VSUBS 0.008562f
C547 B.n255 VSUBS 0.008562f
C548 B.n256 VSUBS 0.008562f
C549 B.n257 VSUBS 0.008562f
C550 B.n258 VSUBS 0.008562f
C551 B.n259 VSUBS 0.008562f
C552 B.n260 VSUBS 0.008562f
C553 B.n261 VSUBS 0.008562f
C554 B.n262 VSUBS 0.008562f
C555 B.n263 VSUBS 0.008562f
C556 B.n264 VSUBS 0.008562f
C557 B.n265 VSUBS 0.008562f
C558 B.n266 VSUBS 0.008562f
C559 B.n267 VSUBS 0.008562f
C560 B.n268 VSUBS 0.008562f
C561 B.n269 VSUBS 0.008562f
C562 B.n270 VSUBS 0.008562f
C563 B.n271 VSUBS 0.008562f
C564 B.n272 VSUBS 0.008562f
C565 B.n273 VSUBS 0.008562f
C566 B.n274 VSUBS 0.008562f
C567 B.n275 VSUBS 0.008562f
C568 B.n276 VSUBS 0.008562f
C569 B.n277 VSUBS 0.008562f
C570 B.n278 VSUBS 0.008562f
C571 B.n279 VSUBS 0.008562f
C572 B.n280 VSUBS 0.008562f
C573 B.n281 VSUBS 0.008562f
C574 B.n282 VSUBS 0.008562f
C575 B.n283 VSUBS 0.008562f
C576 B.n284 VSUBS 0.008562f
C577 B.n285 VSUBS 0.008562f
C578 B.n286 VSUBS 0.008562f
C579 B.n287 VSUBS 0.008562f
C580 B.n288 VSUBS 0.008562f
C581 B.n289 VSUBS 0.008562f
C582 B.n290 VSUBS 0.008562f
C583 B.n291 VSUBS 0.008562f
C584 B.n292 VSUBS 0.008562f
C585 B.n293 VSUBS 0.008562f
C586 B.n294 VSUBS 0.008562f
C587 B.n295 VSUBS 0.008562f
C588 B.n296 VSUBS 0.008562f
C589 B.n297 VSUBS 0.008562f
C590 B.n298 VSUBS 0.008562f
C591 B.n299 VSUBS 0.008562f
C592 B.n300 VSUBS 0.008562f
C593 B.n301 VSUBS 0.008562f
C594 B.n302 VSUBS 0.008562f
C595 B.n303 VSUBS 0.008562f
C596 B.n304 VSUBS 0.008562f
C597 B.n305 VSUBS 0.008562f
C598 B.n306 VSUBS 0.008562f
C599 B.n307 VSUBS 0.008562f
C600 B.n308 VSUBS 0.008562f
C601 B.n309 VSUBS 0.008562f
C602 B.n310 VSUBS 0.008562f
C603 B.n311 VSUBS 0.008562f
C604 B.n312 VSUBS 0.008562f
C605 B.n313 VSUBS 0.008562f
C606 B.n314 VSUBS 0.019107f
C607 B.n315 VSUBS 0.019107f
C608 B.n316 VSUBS 0.020678f
C609 B.n317 VSUBS 0.008562f
C610 B.n318 VSUBS 0.008562f
C611 B.n319 VSUBS 0.008562f
C612 B.n320 VSUBS 0.008562f
C613 B.n321 VSUBS 0.008562f
C614 B.n322 VSUBS 0.008562f
C615 B.n323 VSUBS 0.008562f
C616 B.n324 VSUBS 0.008562f
C617 B.n325 VSUBS 0.008562f
C618 B.n326 VSUBS 0.008562f
C619 B.n327 VSUBS 0.008562f
C620 B.n328 VSUBS 0.008562f
C621 B.n329 VSUBS 0.008562f
C622 B.n330 VSUBS 0.008562f
C623 B.n331 VSUBS 0.008562f
C624 B.n332 VSUBS 0.008562f
C625 B.n333 VSUBS 0.008562f
C626 B.n334 VSUBS 0.008562f
C627 B.n335 VSUBS 0.008562f
C628 B.n336 VSUBS 0.008562f
C629 B.n337 VSUBS 0.008562f
C630 B.n338 VSUBS 0.008562f
C631 B.n339 VSUBS 0.008562f
C632 B.n340 VSUBS 0.008562f
C633 B.n341 VSUBS 0.008562f
C634 B.n342 VSUBS 0.008562f
C635 B.n343 VSUBS 0.008562f
C636 B.n344 VSUBS 0.008562f
C637 B.n345 VSUBS 0.008562f
C638 B.n346 VSUBS 0.008562f
C639 B.n347 VSUBS 0.008562f
C640 B.n348 VSUBS 0.008562f
C641 B.n349 VSUBS 0.008562f
C642 B.n350 VSUBS 0.008562f
C643 B.n351 VSUBS 0.008562f
C644 B.n352 VSUBS 0.008562f
C645 B.n353 VSUBS 0.008562f
C646 B.n354 VSUBS 0.008562f
C647 B.n355 VSUBS 0.008562f
C648 B.n356 VSUBS 0.008562f
C649 B.n357 VSUBS 0.008562f
C650 B.n358 VSUBS 0.008562f
C651 B.n359 VSUBS 0.008562f
C652 B.n360 VSUBS 0.008562f
C653 B.n361 VSUBS 0.008562f
C654 B.n362 VSUBS 0.008562f
C655 B.n363 VSUBS 0.008562f
C656 B.n364 VSUBS 0.008562f
C657 B.n365 VSUBS 0.008562f
C658 B.n366 VSUBS 0.008562f
C659 B.n367 VSUBS 0.008562f
C660 B.n368 VSUBS 0.008562f
C661 B.n369 VSUBS 0.008562f
C662 B.n370 VSUBS 0.008562f
C663 B.n371 VSUBS 0.008562f
C664 B.n372 VSUBS 0.008562f
C665 B.n373 VSUBS 0.008562f
C666 B.n374 VSUBS 0.008562f
C667 B.n375 VSUBS 0.008562f
C668 B.n376 VSUBS 0.008562f
C669 B.n377 VSUBS 0.008562f
C670 B.n378 VSUBS 0.008562f
C671 B.n379 VSUBS 0.008562f
C672 B.n380 VSUBS 0.008562f
C673 B.n381 VSUBS 0.008562f
C674 B.n382 VSUBS 0.008562f
C675 B.n383 VSUBS 0.008562f
C676 B.n384 VSUBS 0.008562f
C677 B.n385 VSUBS 0.008562f
C678 B.n386 VSUBS 0.008562f
C679 B.n387 VSUBS 0.008562f
C680 B.n388 VSUBS 0.008562f
C681 B.n389 VSUBS 0.008562f
C682 B.n390 VSUBS 0.008562f
C683 B.n391 VSUBS 0.008562f
C684 B.n392 VSUBS 0.008562f
C685 B.n393 VSUBS 0.008562f
C686 B.n394 VSUBS 0.008562f
C687 B.n395 VSUBS 0.008562f
C688 B.n396 VSUBS 0.008562f
C689 B.n397 VSUBS 0.005918f
C690 B.n398 VSUBS 0.019836f
C691 B.n399 VSUBS 0.006925f
C692 B.n400 VSUBS 0.008562f
C693 B.n401 VSUBS 0.008562f
C694 B.n402 VSUBS 0.008562f
C695 B.n403 VSUBS 0.008562f
C696 B.n404 VSUBS 0.008562f
C697 B.n405 VSUBS 0.008562f
C698 B.n406 VSUBS 0.008562f
C699 B.n407 VSUBS 0.008562f
C700 B.n408 VSUBS 0.008562f
C701 B.n409 VSUBS 0.008562f
C702 B.n410 VSUBS 0.008562f
C703 B.t1 VSUBS 0.672072f
C704 B.t2 VSUBS 0.695832f
C705 B.t0 VSUBS 2.02042f
C706 B.n411 VSUBS 0.358385f
C707 B.n412 VSUBS 0.086543f
C708 B.n413 VSUBS 0.019836f
C709 B.n414 VSUBS 0.006925f
C710 B.n415 VSUBS 0.008562f
C711 B.n416 VSUBS 0.008562f
C712 B.n417 VSUBS 0.008562f
C713 B.n418 VSUBS 0.008562f
C714 B.n419 VSUBS 0.008562f
C715 B.n420 VSUBS 0.008562f
C716 B.n421 VSUBS 0.008562f
C717 B.n422 VSUBS 0.008562f
C718 B.n423 VSUBS 0.008562f
C719 B.n424 VSUBS 0.008562f
C720 B.n425 VSUBS 0.008562f
C721 B.n426 VSUBS 0.008562f
C722 B.n427 VSUBS 0.008562f
C723 B.n428 VSUBS 0.008562f
C724 B.n429 VSUBS 0.008562f
C725 B.n430 VSUBS 0.008562f
C726 B.n431 VSUBS 0.008562f
C727 B.n432 VSUBS 0.008562f
C728 B.n433 VSUBS 0.008562f
C729 B.n434 VSUBS 0.008562f
C730 B.n435 VSUBS 0.008562f
C731 B.n436 VSUBS 0.008562f
C732 B.n437 VSUBS 0.008562f
C733 B.n438 VSUBS 0.008562f
C734 B.n439 VSUBS 0.008562f
C735 B.n440 VSUBS 0.008562f
C736 B.n441 VSUBS 0.008562f
C737 B.n442 VSUBS 0.008562f
C738 B.n443 VSUBS 0.008562f
C739 B.n444 VSUBS 0.008562f
C740 B.n445 VSUBS 0.008562f
C741 B.n446 VSUBS 0.008562f
C742 B.n447 VSUBS 0.008562f
C743 B.n448 VSUBS 0.008562f
C744 B.n449 VSUBS 0.008562f
C745 B.n450 VSUBS 0.008562f
C746 B.n451 VSUBS 0.008562f
C747 B.n452 VSUBS 0.008562f
C748 B.n453 VSUBS 0.008562f
C749 B.n454 VSUBS 0.008562f
C750 B.n455 VSUBS 0.008562f
C751 B.n456 VSUBS 0.008562f
C752 B.n457 VSUBS 0.008562f
C753 B.n458 VSUBS 0.008562f
C754 B.n459 VSUBS 0.008562f
C755 B.n460 VSUBS 0.008562f
C756 B.n461 VSUBS 0.008562f
C757 B.n462 VSUBS 0.008562f
C758 B.n463 VSUBS 0.008562f
C759 B.n464 VSUBS 0.008562f
C760 B.n465 VSUBS 0.008562f
C761 B.n466 VSUBS 0.008562f
C762 B.n467 VSUBS 0.008562f
C763 B.n468 VSUBS 0.008562f
C764 B.n469 VSUBS 0.008562f
C765 B.n470 VSUBS 0.008562f
C766 B.n471 VSUBS 0.008562f
C767 B.n472 VSUBS 0.008562f
C768 B.n473 VSUBS 0.008562f
C769 B.n474 VSUBS 0.008562f
C770 B.n475 VSUBS 0.008562f
C771 B.n476 VSUBS 0.008562f
C772 B.n477 VSUBS 0.008562f
C773 B.n478 VSUBS 0.008562f
C774 B.n479 VSUBS 0.008562f
C775 B.n480 VSUBS 0.008562f
C776 B.n481 VSUBS 0.008562f
C777 B.n482 VSUBS 0.008562f
C778 B.n483 VSUBS 0.008562f
C779 B.n484 VSUBS 0.008562f
C780 B.n485 VSUBS 0.008562f
C781 B.n486 VSUBS 0.008562f
C782 B.n487 VSUBS 0.008562f
C783 B.n488 VSUBS 0.008562f
C784 B.n489 VSUBS 0.008562f
C785 B.n490 VSUBS 0.008562f
C786 B.n491 VSUBS 0.008562f
C787 B.n492 VSUBS 0.008562f
C788 B.n493 VSUBS 0.008562f
C789 B.n494 VSUBS 0.008562f
C790 B.n495 VSUBS 0.008562f
C791 B.n496 VSUBS 0.008562f
C792 B.n497 VSUBS 0.020678f
C793 B.n498 VSUBS 0.019107f
C794 B.n499 VSUBS 0.019107f
C795 B.n500 VSUBS 0.008562f
C796 B.n501 VSUBS 0.008562f
C797 B.n502 VSUBS 0.008562f
C798 B.n503 VSUBS 0.008562f
C799 B.n504 VSUBS 0.008562f
C800 B.n505 VSUBS 0.008562f
C801 B.n506 VSUBS 0.008562f
C802 B.n507 VSUBS 0.008562f
C803 B.n508 VSUBS 0.008562f
C804 B.n509 VSUBS 0.008562f
C805 B.n510 VSUBS 0.008562f
C806 B.n511 VSUBS 0.008562f
C807 B.n512 VSUBS 0.008562f
C808 B.n513 VSUBS 0.008562f
C809 B.n514 VSUBS 0.008562f
C810 B.n515 VSUBS 0.008562f
C811 B.n516 VSUBS 0.008562f
C812 B.n517 VSUBS 0.008562f
C813 B.n518 VSUBS 0.008562f
C814 B.n519 VSUBS 0.008562f
C815 B.n520 VSUBS 0.008562f
C816 B.n521 VSUBS 0.008562f
C817 B.n522 VSUBS 0.008562f
C818 B.n523 VSUBS 0.008562f
C819 B.n524 VSUBS 0.008562f
C820 B.n525 VSUBS 0.008562f
C821 B.n526 VSUBS 0.008562f
C822 B.n527 VSUBS 0.008562f
C823 B.n528 VSUBS 0.008562f
C824 B.n529 VSUBS 0.008562f
C825 B.n530 VSUBS 0.008562f
C826 B.n531 VSUBS 0.008562f
C827 B.n532 VSUBS 0.008562f
C828 B.n533 VSUBS 0.008562f
C829 B.n534 VSUBS 0.008562f
C830 B.n535 VSUBS 0.008562f
C831 B.n536 VSUBS 0.008562f
C832 B.n537 VSUBS 0.008562f
C833 B.n538 VSUBS 0.008562f
C834 B.n539 VSUBS 0.008562f
C835 B.n540 VSUBS 0.008562f
C836 B.n541 VSUBS 0.008562f
C837 B.n542 VSUBS 0.008562f
C838 B.n543 VSUBS 0.008562f
C839 B.n544 VSUBS 0.008562f
C840 B.n545 VSUBS 0.008562f
C841 B.n546 VSUBS 0.008562f
C842 B.n547 VSUBS 0.008562f
C843 B.n548 VSUBS 0.008562f
C844 B.n549 VSUBS 0.008562f
C845 B.n550 VSUBS 0.008562f
C846 B.n551 VSUBS 0.008562f
C847 B.n552 VSUBS 0.008562f
C848 B.n553 VSUBS 0.008562f
C849 B.n554 VSUBS 0.008562f
C850 B.n555 VSUBS 0.008562f
C851 B.n556 VSUBS 0.008562f
C852 B.n557 VSUBS 0.008562f
C853 B.n558 VSUBS 0.008562f
C854 B.n559 VSUBS 0.008562f
C855 B.n560 VSUBS 0.008562f
C856 B.n561 VSUBS 0.008562f
C857 B.n562 VSUBS 0.008562f
C858 B.n563 VSUBS 0.008562f
C859 B.n564 VSUBS 0.008562f
C860 B.n565 VSUBS 0.008562f
C861 B.n566 VSUBS 0.008562f
C862 B.n567 VSUBS 0.008562f
C863 B.n568 VSUBS 0.008562f
C864 B.n569 VSUBS 0.008562f
C865 B.n570 VSUBS 0.008562f
C866 B.n571 VSUBS 0.008562f
C867 B.n572 VSUBS 0.008562f
C868 B.n573 VSUBS 0.008562f
C869 B.n574 VSUBS 0.008562f
C870 B.n575 VSUBS 0.008562f
C871 B.n576 VSUBS 0.008562f
C872 B.n577 VSUBS 0.008562f
C873 B.n578 VSUBS 0.008562f
C874 B.n579 VSUBS 0.008562f
C875 B.n580 VSUBS 0.008562f
C876 B.n581 VSUBS 0.008562f
C877 B.n582 VSUBS 0.008562f
C878 B.n583 VSUBS 0.008562f
C879 B.n584 VSUBS 0.008562f
C880 B.n585 VSUBS 0.008562f
C881 B.n586 VSUBS 0.008562f
C882 B.n587 VSUBS 0.008562f
C883 B.n588 VSUBS 0.008562f
C884 B.n589 VSUBS 0.008562f
C885 B.n590 VSUBS 0.008562f
C886 B.n591 VSUBS 0.008562f
C887 B.n592 VSUBS 0.008562f
C888 B.n593 VSUBS 0.008562f
C889 B.n594 VSUBS 0.008562f
C890 B.n595 VSUBS 0.008562f
C891 B.n596 VSUBS 0.008562f
C892 B.n597 VSUBS 0.008562f
C893 B.n598 VSUBS 0.008562f
C894 B.n599 VSUBS 0.008562f
C895 B.n600 VSUBS 0.008562f
C896 B.n601 VSUBS 0.008562f
C897 B.n602 VSUBS 0.008562f
C898 B.n603 VSUBS 0.008562f
C899 B.n604 VSUBS 0.008562f
C900 B.n605 VSUBS 0.008562f
C901 B.n606 VSUBS 0.008562f
C902 B.n607 VSUBS 0.008562f
C903 B.n608 VSUBS 0.008562f
C904 B.n609 VSUBS 0.008562f
C905 B.n610 VSUBS 0.008562f
C906 B.n611 VSUBS 0.008562f
C907 B.n612 VSUBS 0.008562f
C908 B.n613 VSUBS 0.008562f
C909 B.n614 VSUBS 0.008562f
C910 B.n615 VSUBS 0.008562f
C911 B.n616 VSUBS 0.008562f
C912 B.n617 VSUBS 0.008562f
C913 B.n618 VSUBS 0.008562f
C914 B.n619 VSUBS 0.008562f
C915 B.n620 VSUBS 0.008562f
C916 B.n621 VSUBS 0.008562f
C917 B.n622 VSUBS 0.008562f
C918 B.n623 VSUBS 0.008562f
C919 B.n624 VSUBS 0.008562f
C920 B.n625 VSUBS 0.008562f
C921 B.n626 VSUBS 0.008562f
C922 B.n627 VSUBS 0.008562f
C923 B.n628 VSUBS 0.008562f
C924 B.n629 VSUBS 0.008562f
C925 B.n630 VSUBS 0.008562f
C926 B.n631 VSUBS 0.008562f
C927 B.n632 VSUBS 0.008562f
C928 B.n633 VSUBS 0.008562f
C929 B.n634 VSUBS 0.008562f
C930 B.n635 VSUBS 0.008562f
C931 B.n636 VSUBS 0.008562f
C932 B.n637 VSUBS 0.008562f
C933 B.n638 VSUBS 0.008562f
C934 B.n639 VSUBS 0.008562f
C935 B.n640 VSUBS 0.008562f
C936 B.n641 VSUBS 0.008562f
C937 B.n642 VSUBS 0.008562f
C938 B.n643 VSUBS 0.008562f
C939 B.n644 VSUBS 0.008562f
C940 B.n645 VSUBS 0.008562f
C941 B.n646 VSUBS 0.008562f
C942 B.n647 VSUBS 0.008562f
C943 B.n648 VSUBS 0.008562f
C944 B.n649 VSUBS 0.008562f
C945 B.n650 VSUBS 0.008562f
C946 B.n651 VSUBS 0.008562f
C947 B.n652 VSUBS 0.008562f
C948 B.n653 VSUBS 0.008562f
C949 B.n654 VSUBS 0.008562f
C950 B.n655 VSUBS 0.008562f
C951 B.n656 VSUBS 0.008562f
C952 B.n657 VSUBS 0.008562f
C953 B.n658 VSUBS 0.008562f
C954 B.n659 VSUBS 0.008562f
C955 B.n660 VSUBS 0.02013f
C956 B.n661 VSUBS 0.019107f
C957 B.n662 VSUBS 0.020678f
C958 B.n663 VSUBS 0.008562f
C959 B.n664 VSUBS 0.008562f
C960 B.n665 VSUBS 0.008562f
C961 B.n666 VSUBS 0.008562f
C962 B.n667 VSUBS 0.008562f
C963 B.n668 VSUBS 0.008562f
C964 B.n669 VSUBS 0.008562f
C965 B.n670 VSUBS 0.008562f
C966 B.n671 VSUBS 0.008562f
C967 B.n672 VSUBS 0.008562f
C968 B.n673 VSUBS 0.008562f
C969 B.n674 VSUBS 0.008562f
C970 B.n675 VSUBS 0.008562f
C971 B.n676 VSUBS 0.008562f
C972 B.n677 VSUBS 0.008562f
C973 B.n678 VSUBS 0.008562f
C974 B.n679 VSUBS 0.008562f
C975 B.n680 VSUBS 0.008562f
C976 B.n681 VSUBS 0.008562f
C977 B.n682 VSUBS 0.008562f
C978 B.n683 VSUBS 0.008562f
C979 B.n684 VSUBS 0.008562f
C980 B.n685 VSUBS 0.008562f
C981 B.n686 VSUBS 0.008562f
C982 B.n687 VSUBS 0.008562f
C983 B.n688 VSUBS 0.008562f
C984 B.n689 VSUBS 0.008562f
C985 B.n690 VSUBS 0.008562f
C986 B.n691 VSUBS 0.008562f
C987 B.n692 VSUBS 0.008562f
C988 B.n693 VSUBS 0.008562f
C989 B.n694 VSUBS 0.008562f
C990 B.n695 VSUBS 0.008562f
C991 B.n696 VSUBS 0.008562f
C992 B.n697 VSUBS 0.008562f
C993 B.n698 VSUBS 0.008562f
C994 B.n699 VSUBS 0.008562f
C995 B.n700 VSUBS 0.008562f
C996 B.n701 VSUBS 0.008562f
C997 B.n702 VSUBS 0.008562f
C998 B.n703 VSUBS 0.008562f
C999 B.n704 VSUBS 0.008562f
C1000 B.n705 VSUBS 0.008562f
C1001 B.n706 VSUBS 0.008562f
C1002 B.n707 VSUBS 0.008562f
C1003 B.n708 VSUBS 0.008562f
C1004 B.n709 VSUBS 0.008562f
C1005 B.n710 VSUBS 0.008562f
C1006 B.n711 VSUBS 0.008562f
C1007 B.n712 VSUBS 0.008562f
C1008 B.n713 VSUBS 0.008562f
C1009 B.n714 VSUBS 0.008562f
C1010 B.n715 VSUBS 0.008562f
C1011 B.n716 VSUBS 0.008562f
C1012 B.n717 VSUBS 0.008562f
C1013 B.n718 VSUBS 0.008562f
C1014 B.n719 VSUBS 0.008562f
C1015 B.n720 VSUBS 0.008562f
C1016 B.n721 VSUBS 0.008562f
C1017 B.n722 VSUBS 0.008562f
C1018 B.n723 VSUBS 0.008562f
C1019 B.n724 VSUBS 0.008562f
C1020 B.n725 VSUBS 0.008562f
C1021 B.n726 VSUBS 0.008562f
C1022 B.n727 VSUBS 0.008562f
C1023 B.n728 VSUBS 0.008562f
C1024 B.n729 VSUBS 0.008562f
C1025 B.n730 VSUBS 0.008562f
C1026 B.n731 VSUBS 0.008562f
C1027 B.n732 VSUBS 0.008562f
C1028 B.n733 VSUBS 0.008562f
C1029 B.n734 VSUBS 0.008562f
C1030 B.n735 VSUBS 0.008562f
C1031 B.n736 VSUBS 0.008562f
C1032 B.n737 VSUBS 0.008562f
C1033 B.n738 VSUBS 0.008562f
C1034 B.n739 VSUBS 0.008562f
C1035 B.n740 VSUBS 0.008562f
C1036 B.n741 VSUBS 0.008562f
C1037 B.n742 VSUBS 0.008562f
C1038 B.n743 VSUBS 0.005918f
C1039 B.n744 VSUBS 0.019836f
C1040 B.n745 VSUBS 0.006925f
C1041 B.n746 VSUBS 0.008562f
C1042 B.n747 VSUBS 0.008562f
C1043 B.n748 VSUBS 0.008562f
C1044 B.n749 VSUBS 0.008562f
C1045 B.n750 VSUBS 0.008562f
C1046 B.n751 VSUBS 0.008562f
C1047 B.n752 VSUBS 0.008562f
C1048 B.n753 VSUBS 0.008562f
C1049 B.n754 VSUBS 0.008562f
C1050 B.n755 VSUBS 0.008562f
C1051 B.n756 VSUBS 0.008562f
C1052 B.n757 VSUBS 0.006925f
C1053 B.n758 VSUBS 0.008562f
C1054 B.n759 VSUBS 0.008562f
C1055 B.n760 VSUBS 0.008562f
C1056 B.n761 VSUBS 0.008562f
C1057 B.n762 VSUBS 0.008562f
C1058 B.n763 VSUBS 0.008562f
C1059 B.n764 VSUBS 0.008562f
C1060 B.n765 VSUBS 0.008562f
C1061 B.n766 VSUBS 0.008562f
C1062 B.n767 VSUBS 0.008562f
C1063 B.n768 VSUBS 0.008562f
C1064 B.n769 VSUBS 0.008562f
C1065 B.n770 VSUBS 0.008562f
C1066 B.n771 VSUBS 0.008562f
C1067 B.n772 VSUBS 0.008562f
C1068 B.n773 VSUBS 0.008562f
C1069 B.n774 VSUBS 0.008562f
C1070 B.n775 VSUBS 0.008562f
C1071 B.n776 VSUBS 0.008562f
C1072 B.n777 VSUBS 0.008562f
C1073 B.n778 VSUBS 0.008562f
C1074 B.n779 VSUBS 0.008562f
C1075 B.n780 VSUBS 0.008562f
C1076 B.n781 VSUBS 0.008562f
C1077 B.n782 VSUBS 0.008562f
C1078 B.n783 VSUBS 0.008562f
C1079 B.n784 VSUBS 0.008562f
C1080 B.n785 VSUBS 0.008562f
C1081 B.n786 VSUBS 0.008562f
C1082 B.n787 VSUBS 0.008562f
C1083 B.n788 VSUBS 0.008562f
C1084 B.n789 VSUBS 0.008562f
C1085 B.n790 VSUBS 0.008562f
C1086 B.n791 VSUBS 0.008562f
C1087 B.n792 VSUBS 0.008562f
C1088 B.n793 VSUBS 0.008562f
C1089 B.n794 VSUBS 0.008562f
C1090 B.n795 VSUBS 0.008562f
C1091 B.n796 VSUBS 0.008562f
C1092 B.n797 VSUBS 0.008562f
C1093 B.n798 VSUBS 0.008562f
C1094 B.n799 VSUBS 0.008562f
C1095 B.n800 VSUBS 0.008562f
C1096 B.n801 VSUBS 0.008562f
C1097 B.n802 VSUBS 0.008562f
C1098 B.n803 VSUBS 0.008562f
C1099 B.n804 VSUBS 0.008562f
C1100 B.n805 VSUBS 0.008562f
C1101 B.n806 VSUBS 0.008562f
C1102 B.n807 VSUBS 0.008562f
C1103 B.n808 VSUBS 0.008562f
C1104 B.n809 VSUBS 0.008562f
C1105 B.n810 VSUBS 0.008562f
C1106 B.n811 VSUBS 0.008562f
C1107 B.n812 VSUBS 0.008562f
C1108 B.n813 VSUBS 0.008562f
C1109 B.n814 VSUBS 0.008562f
C1110 B.n815 VSUBS 0.008562f
C1111 B.n816 VSUBS 0.008562f
C1112 B.n817 VSUBS 0.008562f
C1113 B.n818 VSUBS 0.008562f
C1114 B.n819 VSUBS 0.008562f
C1115 B.n820 VSUBS 0.008562f
C1116 B.n821 VSUBS 0.008562f
C1117 B.n822 VSUBS 0.008562f
C1118 B.n823 VSUBS 0.008562f
C1119 B.n824 VSUBS 0.008562f
C1120 B.n825 VSUBS 0.008562f
C1121 B.n826 VSUBS 0.008562f
C1122 B.n827 VSUBS 0.008562f
C1123 B.n828 VSUBS 0.008562f
C1124 B.n829 VSUBS 0.008562f
C1125 B.n830 VSUBS 0.008562f
C1126 B.n831 VSUBS 0.008562f
C1127 B.n832 VSUBS 0.008562f
C1128 B.n833 VSUBS 0.008562f
C1129 B.n834 VSUBS 0.008562f
C1130 B.n835 VSUBS 0.008562f
C1131 B.n836 VSUBS 0.008562f
C1132 B.n837 VSUBS 0.008562f
C1133 B.n838 VSUBS 0.008562f
C1134 B.n839 VSUBS 0.008562f
C1135 B.n840 VSUBS 0.020678f
C1136 B.n841 VSUBS 0.019107f
C1137 B.n842 VSUBS 0.019107f
C1138 B.n843 VSUBS 0.008562f
C1139 B.n844 VSUBS 0.008562f
C1140 B.n845 VSUBS 0.008562f
C1141 B.n846 VSUBS 0.008562f
C1142 B.n847 VSUBS 0.008562f
C1143 B.n848 VSUBS 0.008562f
C1144 B.n849 VSUBS 0.008562f
C1145 B.n850 VSUBS 0.008562f
C1146 B.n851 VSUBS 0.008562f
C1147 B.n852 VSUBS 0.008562f
C1148 B.n853 VSUBS 0.008562f
C1149 B.n854 VSUBS 0.008562f
C1150 B.n855 VSUBS 0.008562f
C1151 B.n856 VSUBS 0.008562f
C1152 B.n857 VSUBS 0.008562f
C1153 B.n858 VSUBS 0.008562f
C1154 B.n859 VSUBS 0.008562f
C1155 B.n860 VSUBS 0.008562f
C1156 B.n861 VSUBS 0.008562f
C1157 B.n862 VSUBS 0.008562f
C1158 B.n863 VSUBS 0.008562f
C1159 B.n864 VSUBS 0.008562f
C1160 B.n865 VSUBS 0.008562f
C1161 B.n866 VSUBS 0.008562f
C1162 B.n867 VSUBS 0.008562f
C1163 B.n868 VSUBS 0.008562f
C1164 B.n869 VSUBS 0.008562f
C1165 B.n870 VSUBS 0.008562f
C1166 B.n871 VSUBS 0.008562f
C1167 B.n872 VSUBS 0.008562f
C1168 B.n873 VSUBS 0.008562f
C1169 B.n874 VSUBS 0.008562f
C1170 B.n875 VSUBS 0.008562f
C1171 B.n876 VSUBS 0.008562f
C1172 B.n877 VSUBS 0.008562f
C1173 B.n878 VSUBS 0.008562f
C1174 B.n879 VSUBS 0.008562f
C1175 B.n880 VSUBS 0.008562f
C1176 B.n881 VSUBS 0.008562f
C1177 B.n882 VSUBS 0.008562f
C1178 B.n883 VSUBS 0.008562f
C1179 B.n884 VSUBS 0.008562f
C1180 B.n885 VSUBS 0.008562f
C1181 B.n886 VSUBS 0.008562f
C1182 B.n887 VSUBS 0.008562f
C1183 B.n888 VSUBS 0.008562f
C1184 B.n889 VSUBS 0.008562f
C1185 B.n890 VSUBS 0.008562f
C1186 B.n891 VSUBS 0.008562f
C1187 B.n892 VSUBS 0.008562f
C1188 B.n893 VSUBS 0.008562f
C1189 B.n894 VSUBS 0.008562f
C1190 B.n895 VSUBS 0.008562f
C1191 B.n896 VSUBS 0.008562f
C1192 B.n897 VSUBS 0.008562f
C1193 B.n898 VSUBS 0.008562f
C1194 B.n899 VSUBS 0.008562f
C1195 B.n900 VSUBS 0.008562f
C1196 B.n901 VSUBS 0.008562f
C1197 B.n902 VSUBS 0.008562f
C1198 B.n903 VSUBS 0.008562f
C1199 B.n904 VSUBS 0.008562f
C1200 B.n905 VSUBS 0.008562f
C1201 B.n906 VSUBS 0.008562f
C1202 B.n907 VSUBS 0.008562f
C1203 B.n908 VSUBS 0.008562f
C1204 B.n909 VSUBS 0.008562f
C1205 B.n910 VSUBS 0.008562f
C1206 B.n911 VSUBS 0.008562f
C1207 B.n912 VSUBS 0.008562f
C1208 B.n913 VSUBS 0.008562f
C1209 B.n914 VSUBS 0.008562f
C1210 B.n915 VSUBS 0.008562f
C1211 B.n916 VSUBS 0.008562f
C1212 B.n917 VSUBS 0.008562f
C1213 B.n918 VSUBS 0.008562f
C1214 B.n919 VSUBS 0.008562f
C1215 B.n920 VSUBS 0.008562f
C1216 B.n921 VSUBS 0.008562f
C1217 B.n922 VSUBS 0.008562f
C1218 B.n923 VSUBS 0.019386f
.ends

