* NGSPICE file created from diff_pair_sample_0771.ext - technology: sky130A

.subckt diff_pair_sample_0771 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=4.5747 pd=24.24 as=0 ps=0 w=11.73 l=2.95
X1 B.t8 B.t6 B.t7 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=4.5747 pd=24.24 as=0 ps=0 w=11.73 l=2.95
X2 VTAIL.t11 VN.t0 VDD2.t0 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=1.93545 pd=12.06 as=1.93545 ps=12.06 w=11.73 l=2.95
X3 VTAIL.t3 VP.t0 VDD1.t5 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=1.93545 pd=12.06 as=1.93545 ps=12.06 w=11.73 l=2.95
X4 B.t5 B.t3 B.t4 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=4.5747 pd=24.24 as=0 ps=0 w=11.73 l=2.95
X5 VDD2.t3 VN.t1 VTAIL.t10 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=1.93545 pd=12.06 as=4.5747 ps=24.24 w=11.73 l=2.95
X6 VTAIL.t9 VN.t2 VDD2.t5 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=1.93545 pd=12.06 as=1.93545 ps=12.06 w=11.73 l=2.95
X7 B.t2 B.t0 B.t1 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=4.5747 pd=24.24 as=0 ps=0 w=11.73 l=2.95
X8 VDD1.t4 VP.t1 VTAIL.t0 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=4.5747 pd=24.24 as=1.93545 ps=12.06 w=11.73 l=2.95
X9 VDD1.t3 VP.t2 VTAIL.t2 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=1.93545 pd=12.06 as=4.5747 ps=24.24 w=11.73 l=2.95
X10 VDD2.t2 VN.t3 VTAIL.t8 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=1.93545 pd=12.06 as=4.5747 ps=24.24 w=11.73 l=2.95
X11 VTAIL.t1 VP.t3 VDD1.t2 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=1.93545 pd=12.06 as=1.93545 ps=12.06 w=11.73 l=2.95
X12 VDD2.t1 VN.t4 VTAIL.t7 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=4.5747 pd=24.24 as=1.93545 ps=12.06 w=11.73 l=2.95
X13 VDD1.t1 VP.t4 VTAIL.t5 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=4.5747 pd=24.24 as=1.93545 ps=12.06 w=11.73 l=2.95
X14 VDD2.t4 VN.t5 VTAIL.t6 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=4.5747 pd=24.24 as=1.93545 ps=12.06 w=11.73 l=2.95
X15 VDD1.t0 VP.t5 VTAIL.t4 w_n3594_n3314# sky130_fd_pr__pfet_01v8 ad=1.93545 pd=12.06 as=4.5747 ps=24.24 w=11.73 l=2.95
R0 B.n399 B.n122 585
R1 B.n398 B.n397 585
R2 B.n396 B.n123 585
R3 B.n395 B.n394 585
R4 B.n393 B.n124 585
R5 B.n392 B.n391 585
R6 B.n390 B.n125 585
R7 B.n389 B.n388 585
R8 B.n387 B.n126 585
R9 B.n386 B.n385 585
R10 B.n384 B.n127 585
R11 B.n383 B.n382 585
R12 B.n381 B.n128 585
R13 B.n380 B.n379 585
R14 B.n378 B.n129 585
R15 B.n377 B.n376 585
R16 B.n375 B.n130 585
R17 B.n374 B.n373 585
R18 B.n372 B.n131 585
R19 B.n371 B.n370 585
R20 B.n369 B.n132 585
R21 B.n368 B.n367 585
R22 B.n366 B.n133 585
R23 B.n365 B.n364 585
R24 B.n363 B.n134 585
R25 B.n362 B.n361 585
R26 B.n360 B.n135 585
R27 B.n359 B.n358 585
R28 B.n357 B.n136 585
R29 B.n356 B.n355 585
R30 B.n354 B.n137 585
R31 B.n353 B.n352 585
R32 B.n351 B.n138 585
R33 B.n350 B.n349 585
R34 B.n348 B.n139 585
R35 B.n347 B.n346 585
R36 B.n345 B.n140 585
R37 B.n344 B.n343 585
R38 B.n342 B.n141 585
R39 B.n341 B.n340 585
R40 B.n339 B.n142 585
R41 B.n338 B.n337 585
R42 B.n333 B.n143 585
R43 B.n332 B.n331 585
R44 B.n330 B.n144 585
R45 B.n329 B.n328 585
R46 B.n327 B.n145 585
R47 B.n326 B.n325 585
R48 B.n324 B.n146 585
R49 B.n323 B.n322 585
R50 B.n320 B.n147 585
R51 B.n319 B.n318 585
R52 B.n317 B.n150 585
R53 B.n316 B.n315 585
R54 B.n314 B.n151 585
R55 B.n313 B.n312 585
R56 B.n311 B.n152 585
R57 B.n310 B.n309 585
R58 B.n308 B.n153 585
R59 B.n307 B.n306 585
R60 B.n305 B.n154 585
R61 B.n304 B.n303 585
R62 B.n302 B.n155 585
R63 B.n301 B.n300 585
R64 B.n299 B.n156 585
R65 B.n298 B.n297 585
R66 B.n296 B.n157 585
R67 B.n295 B.n294 585
R68 B.n293 B.n158 585
R69 B.n292 B.n291 585
R70 B.n290 B.n159 585
R71 B.n289 B.n288 585
R72 B.n287 B.n160 585
R73 B.n286 B.n285 585
R74 B.n284 B.n161 585
R75 B.n283 B.n282 585
R76 B.n281 B.n162 585
R77 B.n280 B.n279 585
R78 B.n278 B.n163 585
R79 B.n277 B.n276 585
R80 B.n275 B.n164 585
R81 B.n274 B.n273 585
R82 B.n272 B.n165 585
R83 B.n271 B.n270 585
R84 B.n269 B.n166 585
R85 B.n268 B.n267 585
R86 B.n266 B.n167 585
R87 B.n265 B.n264 585
R88 B.n263 B.n168 585
R89 B.n262 B.n261 585
R90 B.n260 B.n169 585
R91 B.n401 B.n400 585
R92 B.n402 B.n121 585
R93 B.n404 B.n403 585
R94 B.n405 B.n120 585
R95 B.n407 B.n406 585
R96 B.n408 B.n119 585
R97 B.n410 B.n409 585
R98 B.n411 B.n118 585
R99 B.n413 B.n412 585
R100 B.n414 B.n117 585
R101 B.n416 B.n415 585
R102 B.n417 B.n116 585
R103 B.n419 B.n418 585
R104 B.n420 B.n115 585
R105 B.n422 B.n421 585
R106 B.n423 B.n114 585
R107 B.n425 B.n424 585
R108 B.n426 B.n113 585
R109 B.n428 B.n427 585
R110 B.n429 B.n112 585
R111 B.n431 B.n430 585
R112 B.n432 B.n111 585
R113 B.n434 B.n433 585
R114 B.n435 B.n110 585
R115 B.n437 B.n436 585
R116 B.n438 B.n109 585
R117 B.n440 B.n439 585
R118 B.n441 B.n108 585
R119 B.n443 B.n442 585
R120 B.n444 B.n107 585
R121 B.n446 B.n445 585
R122 B.n447 B.n106 585
R123 B.n449 B.n448 585
R124 B.n450 B.n105 585
R125 B.n452 B.n451 585
R126 B.n453 B.n104 585
R127 B.n455 B.n454 585
R128 B.n456 B.n103 585
R129 B.n458 B.n457 585
R130 B.n459 B.n102 585
R131 B.n461 B.n460 585
R132 B.n462 B.n101 585
R133 B.n464 B.n463 585
R134 B.n465 B.n100 585
R135 B.n467 B.n466 585
R136 B.n468 B.n99 585
R137 B.n470 B.n469 585
R138 B.n471 B.n98 585
R139 B.n473 B.n472 585
R140 B.n474 B.n97 585
R141 B.n476 B.n475 585
R142 B.n477 B.n96 585
R143 B.n479 B.n478 585
R144 B.n480 B.n95 585
R145 B.n482 B.n481 585
R146 B.n483 B.n94 585
R147 B.n485 B.n484 585
R148 B.n486 B.n93 585
R149 B.n488 B.n487 585
R150 B.n489 B.n92 585
R151 B.n491 B.n490 585
R152 B.n492 B.n91 585
R153 B.n494 B.n493 585
R154 B.n495 B.n90 585
R155 B.n497 B.n496 585
R156 B.n498 B.n89 585
R157 B.n500 B.n499 585
R158 B.n501 B.n88 585
R159 B.n503 B.n502 585
R160 B.n504 B.n87 585
R161 B.n506 B.n505 585
R162 B.n507 B.n86 585
R163 B.n509 B.n508 585
R164 B.n510 B.n85 585
R165 B.n512 B.n511 585
R166 B.n513 B.n84 585
R167 B.n515 B.n514 585
R168 B.n516 B.n83 585
R169 B.n518 B.n517 585
R170 B.n519 B.n82 585
R171 B.n521 B.n520 585
R172 B.n522 B.n81 585
R173 B.n524 B.n523 585
R174 B.n525 B.n80 585
R175 B.n527 B.n526 585
R176 B.n528 B.n79 585
R177 B.n530 B.n529 585
R178 B.n531 B.n78 585
R179 B.n533 B.n532 585
R180 B.n534 B.n77 585
R181 B.n536 B.n535 585
R182 B.n537 B.n76 585
R183 B.n539 B.n538 585
R184 B.n540 B.n75 585
R185 B.n678 B.n25 585
R186 B.n677 B.n676 585
R187 B.n675 B.n26 585
R188 B.n674 B.n673 585
R189 B.n672 B.n27 585
R190 B.n671 B.n670 585
R191 B.n669 B.n28 585
R192 B.n668 B.n667 585
R193 B.n666 B.n29 585
R194 B.n665 B.n664 585
R195 B.n663 B.n30 585
R196 B.n662 B.n661 585
R197 B.n660 B.n31 585
R198 B.n659 B.n658 585
R199 B.n657 B.n32 585
R200 B.n656 B.n655 585
R201 B.n654 B.n33 585
R202 B.n653 B.n652 585
R203 B.n651 B.n34 585
R204 B.n650 B.n649 585
R205 B.n648 B.n35 585
R206 B.n647 B.n646 585
R207 B.n645 B.n36 585
R208 B.n644 B.n643 585
R209 B.n642 B.n37 585
R210 B.n641 B.n640 585
R211 B.n639 B.n38 585
R212 B.n638 B.n637 585
R213 B.n636 B.n39 585
R214 B.n635 B.n634 585
R215 B.n633 B.n40 585
R216 B.n632 B.n631 585
R217 B.n630 B.n41 585
R218 B.n629 B.n628 585
R219 B.n627 B.n42 585
R220 B.n626 B.n625 585
R221 B.n624 B.n43 585
R222 B.n623 B.n622 585
R223 B.n621 B.n44 585
R224 B.n620 B.n619 585
R225 B.n618 B.n45 585
R226 B.n616 B.n615 585
R227 B.n614 B.n48 585
R228 B.n613 B.n612 585
R229 B.n611 B.n49 585
R230 B.n610 B.n609 585
R231 B.n608 B.n50 585
R232 B.n607 B.n606 585
R233 B.n605 B.n51 585
R234 B.n604 B.n603 585
R235 B.n602 B.n601 585
R236 B.n600 B.n55 585
R237 B.n599 B.n598 585
R238 B.n597 B.n56 585
R239 B.n596 B.n595 585
R240 B.n594 B.n57 585
R241 B.n593 B.n592 585
R242 B.n591 B.n58 585
R243 B.n590 B.n589 585
R244 B.n588 B.n59 585
R245 B.n587 B.n586 585
R246 B.n585 B.n60 585
R247 B.n584 B.n583 585
R248 B.n582 B.n61 585
R249 B.n581 B.n580 585
R250 B.n579 B.n62 585
R251 B.n578 B.n577 585
R252 B.n576 B.n63 585
R253 B.n575 B.n574 585
R254 B.n573 B.n64 585
R255 B.n572 B.n571 585
R256 B.n570 B.n65 585
R257 B.n569 B.n568 585
R258 B.n567 B.n66 585
R259 B.n566 B.n565 585
R260 B.n564 B.n67 585
R261 B.n563 B.n562 585
R262 B.n561 B.n68 585
R263 B.n560 B.n559 585
R264 B.n558 B.n69 585
R265 B.n557 B.n556 585
R266 B.n555 B.n70 585
R267 B.n554 B.n553 585
R268 B.n552 B.n71 585
R269 B.n551 B.n550 585
R270 B.n549 B.n72 585
R271 B.n548 B.n547 585
R272 B.n546 B.n73 585
R273 B.n545 B.n544 585
R274 B.n543 B.n74 585
R275 B.n542 B.n541 585
R276 B.n680 B.n679 585
R277 B.n681 B.n24 585
R278 B.n683 B.n682 585
R279 B.n684 B.n23 585
R280 B.n686 B.n685 585
R281 B.n687 B.n22 585
R282 B.n689 B.n688 585
R283 B.n690 B.n21 585
R284 B.n692 B.n691 585
R285 B.n693 B.n20 585
R286 B.n695 B.n694 585
R287 B.n696 B.n19 585
R288 B.n698 B.n697 585
R289 B.n699 B.n18 585
R290 B.n701 B.n700 585
R291 B.n702 B.n17 585
R292 B.n704 B.n703 585
R293 B.n705 B.n16 585
R294 B.n707 B.n706 585
R295 B.n708 B.n15 585
R296 B.n710 B.n709 585
R297 B.n711 B.n14 585
R298 B.n713 B.n712 585
R299 B.n714 B.n13 585
R300 B.n716 B.n715 585
R301 B.n717 B.n12 585
R302 B.n719 B.n718 585
R303 B.n720 B.n11 585
R304 B.n722 B.n721 585
R305 B.n723 B.n10 585
R306 B.n725 B.n724 585
R307 B.n726 B.n9 585
R308 B.n728 B.n727 585
R309 B.n729 B.n8 585
R310 B.n731 B.n730 585
R311 B.n732 B.n7 585
R312 B.n734 B.n733 585
R313 B.n735 B.n6 585
R314 B.n737 B.n736 585
R315 B.n738 B.n5 585
R316 B.n740 B.n739 585
R317 B.n741 B.n4 585
R318 B.n743 B.n742 585
R319 B.n744 B.n3 585
R320 B.n746 B.n745 585
R321 B.n747 B.n0 585
R322 B.n2 B.n1 585
R323 B.n193 B.n192 585
R324 B.n194 B.n191 585
R325 B.n196 B.n195 585
R326 B.n197 B.n190 585
R327 B.n199 B.n198 585
R328 B.n200 B.n189 585
R329 B.n202 B.n201 585
R330 B.n203 B.n188 585
R331 B.n205 B.n204 585
R332 B.n206 B.n187 585
R333 B.n208 B.n207 585
R334 B.n209 B.n186 585
R335 B.n211 B.n210 585
R336 B.n212 B.n185 585
R337 B.n214 B.n213 585
R338 B.n215 B.n184 585
R339 B.n217 B.n216 585
R340 B.n218 B.n183 585
R341 B.n220 B.n219 585
R342 B.n221 B.n182 585
R343 B.n223 B.n222 585
R344 B.n224 B.n181 585
R345 B.n226 B.n225 585
R346 B.n227 B.n180 585
R347 B.n229 B.n228 585
R348 B.n230 B.n179 585
R349 B.n232 B.n231 585
R350 B.n233 B.n178 585
R351 B.n235 B.n234 585
R352 B.n236 B.n177 585
R353 B.n238 B.n237 585
R354 B.n239 B.n176 585
R355 B.n241 B.n240 585
R356 B.n242 B.n175 585
R357 B.n244 B.n243 585
R358 B.n245 B.n174 585
R359 B.n247 B.n246 585
R360 B.n248 B.n173 585
R361 B.n250 B.n249 585
R362 B.n251 B.n172 585
R363 B.n253 B.n252 585
R364 B.n254 B.n171 585
R365 B.n256 B.n255 585
R366 B.n257 B.n170 585
R367 B.n259 B.n258 585
R368 B.n258 B.n169 550.159
R369 B.n400 B.n399 550.159
R370 B.n542 B.n75 550.159
R371 B.n680 B.n25 550.159
R372 B.n148 B.t0 304.349
R373 B.n334 B.t3 304.349
R374 B.n52 B.t9 304.349
R375 B.n46 B.t6 304.349
R376 B.n749 B.n748 256.663
R377 B.n748 B.n747 235.042
R378 B.n748 B.n2 235.042
R379 B.n334 B.t4 174.077
R380 B.n52 B.t11 174.077
R381 B.n148 B.t1 174.064
R382 B.n46 B.t8 174.064
R383 B.n262 B.n169 163.367
R384 B.n263 B.n262 163.367
R385 B.n264 B.n263 163.367
R386 B.n264 B.n167 163.367
R387 B.n268 B.n167 163.367
R388 B.n269 B.n268 163.367
R389 B.n270 B.n269 163.367
R390 B.n270 B.n165 163.367
R391 B.n274 B.n165 163.367
R392 B.n275 B.n274 163.367
R393 B.n276 B.n275 163.367
R394 B.n276 B.n163 163.367
R395 B.n280 B.n163 163.367
R396 B.n281 B.n280 163.367
R397 B.n282 B.n281 163.367
R398 B.n282 B.n161 163.367
R399 B.n286 B.n161 163.367
R400 B.n287 B.n286 163.367
R401 B.n288 B.n287 163.367
R402 B.n288 B.n159 163.367
R403 B.n292 B.n159 163.367
R404 B.n293 B.n292 163.367
R405 B.n294 B.n293 163.367
R406 B.n294 B.n157 163.367
R407 B.n298 B.n157 163.367
R408 B.n299 B.n298 163.367
R409 B.n300 B.n299 163.367
R410 B.n300 B.n155 163.367
R411 B.n304 B.n155 163.367
R412 B.n305 B.n304 163.367
R413 B.n306 B.n305 163.367
R414 B.n306 B.n153 163.367
R415 B.n310 B.n153 163.367
R416 B.n311 B.n310 163.367
R417 B.n312 B.n311 163.367
R418 B.n312 B.n151 163.367
R419 B.n316 B.n151 163.367
R420 B.n317 B.n316 163.367
R421 B.n318 B.n317 163.367
R422 B.n318 B.n147 163.367
R423 B.n323 B.n147 163.367
R424 B.n324 B.n323 163.367
R425 B.n325 B.n324 163.367
R426 B.n325 B.n145 163.367
R427 B.n329 B.n145 163.367
R428 B.n330 B.n329 163.367
R429 B.n331 B.n330 163.367
R430 B.n331 B.n143 163.367
R431 B.n338 B.n143 163.367
R432 B.n339 B.n338 163.367
R433 B.n340 B.n339 163.367
R434 B.n340 B.n141 163.367
R435 B.n344 B.n141 163.367
R436 B.n345 B.n344 163.367
R437 B.n346 B.n345 163.367
R438 B.n346 B.n139 163.367
R439 B.n350 B.n139 163.367
R440 B.n351 B.n350 163.367
R441 B.n352 B.n351 163.367
R442 B.n352 B.n137 163.367
R443 B.n356 B.n137 163.367
R444 B.n357 B.n356 163.367
R445 B.n358 B.n357 163.367
R446 B.n358 B.n135 163.367
R447 B.n362 B.n135 163.367
R448 B.n363 B.n362 163.367
R449 B.n364 B.n363 163.367
R450 B.n364 B.n133 163.367
R451 B.n368 B.n133 163.367
R452 B.n369 B.n368 163.367
R453 B.n370 B.n369 163.367
R454 B.n370 B.n131 163.367
R455 B.n374 B.n131 163.367
R456 B.n375 B.n374 163.367
R457 B.n376 B.n375 163.367
R458 B.n376 B.n129 163.367
R459 B.n380 B.n129 163.367
R460 B.n381 B.n380 163.367
R461 B.n382 B.n381 163.367
R462 B.n382 B.n127 163.367
R463 B.n386 B.n127 163.367
R464 B.n387 B.n386 163.367
R465 B.n388 B.n387 163.367
R466 B.n388 B.n125 163.367
R467 B.n392 B.n125 163.367
R468 B.n393 B.n392 163.367
R469 B.n394 B.n393 163.367
R470 B.n394 B.n123 163.367
R471 B.n398 B.n123 163.367
R472 B.n399 B.n398 163.367
R473 B.n538 B.n75 163.367
R474 B.n538 B.n537 163.367
R475 B.n537 B.n536 163.367
R476 B.n536 B.n77 163.367
R477 B.n532 B.n77 163.367
R478 B.n532 B.n531 163.367
R479 B.n531 B.n530 163.367
R480 B.n530 B.n79 163.367
R481 B.n526 B.n79 163.367
R482 B.n526 B.n525 163.367
R483 B.n525 B.n524 163.367
R484 B.n524 B.n81 163.367
R485 B.n520 B.n81 163.367
R486 B.n520 B.n519 163.367
R487 B.n519 B.n518 163.367
R488 B.n518 B.n83 163.367
R489 B.n514 B.n83 163.367
R490 B.n514 B.n513 163.367
R491 B.n513 B.n512 163.367
R492 B.n512 B.n85 163.367
R493 B.n508 B.n85 163.367
R494 B.n508 B.n507 163.367
R495 B.n507 B.n506 163.367
R496 B.n506 B.n87 163.367
R497 B.n502 B.n87 163.367
R498 B.n502 B.n501 163.367
R499 B.n501 B.n500 163.367
R500 B.n500 B.n89 163.367
R501 B.n496 B.n89 163.367
R502 B.n496 B.n495 163.367
R503 B.n495 B.n494 163.367
R504 B.n494 B.n91 163.367
R505 B.n490 B.n91 163.367
R506 B.n490 B.n489 163.367
R507 B.n489 B.n488 163.367
R508 B.n488 B.n93 163.367
R509 B.n484 B.n93 163.367
R510 B.n484 B.n483 163.367
R511 B.n483 B.n482 163.367
R512 B.n482 B.n95 163.367
R513 B.n478 B.n95 163.367
R514 B.n478 B.n477 163.367
R515 B.n477 B.n476 163.367
R516 B.n476 B.n97 163.367
R517 B.n472 B.n97 163.367
R518 B.n472 B.n471 163.367
R519 B.n471 B.n470 163.367
R520 B.n470 B.n99 163.367
R521 B.n466 B.n99 163.367
R522 B.n466 B.n465 163.367
R523 B.n465 B.n464 163.367
R524 B.n464 B.n101 163.367
R525 B.n460 B.n101 163.367
R526 B.n460 B.n459 163.367
R527 B.n459 B.n458 163.367
R528 B.n458 B.n103 163.367
R529 B.n454 B.n103 163.367
R530 B.n454 B.n453 163.367
R531 B.n453 B.n452 163.367
R532 B.n452 B.n105 163.367
R533 B.n448 B.n105 163.367
R534 B.n448 B.n447 163.367
R535 B.n447 B.n446 163.367
R536 B.n446 B.n107 163.367
R537 B.n442 B.n107 163.367
R538 B.n442 B.n441 163.367
R539 B.n441 B.n440 163.367
R540 B.n440 B.n109 163.367
R541 B.n436 B.n109 163.367
R542 B.n436 B.n435 163.367
R543 B.n435 B.n434 163.367
R544 B.n434 B.n111 163.367
R545 B.n430 B.n111 163.367
R546 B.n430 B.n429 163.367
R547 B.n429 B.n428 163.367
R548 B.n428 B.n113 163.367
R549 B.n424 B.n113 163.367
R550 B.n424 B.n423 163.367
R551 B.n423 B.n422 163.367
R552 B.n422 B.n115 163.367
R553 B.n418 B.n115 163.367
R554 B.n418 B.n417 163.367
R555 B.n417 B.n416 163.367
R556 B.n416 B.n117 163.367
R557 B.n412 B.n117 163.367
R558 B.n412 B.n411 163.367
R559 B.n411 B.n410 163.367
R560 B.n410 B.n119 163.367
R561 B.n406 B.n119 163.367
R562 B.n406 B.n405 163.367
R563 B.n405 B.n404 163.367
R564 B.n404 B.n121 163.367
R565 B.n400 B.n121 163.367
R566 B.n676 B.n25 163.367
R567 B.n676 B.n675 163.367
R568 B.n675 B.n674 163.367
R569 B.n674 B.n27 163.367
R570 B.n670 B.n27 163.367
R571 B.n670 B.n669 163.367
R572 B.n669 B.n668 163.367
R573 B.n668 B.n29 163.367
R574 B.n664 B.n29 163.367
R575 B.n664 B.n663 163.367
R576 B.n663 B.n662 163.367
R577 B.n662 B.n31 163.367
R578 B.n658 B.n31 163.367
R579 B.n658 B.n657 163.367
R580 B.n657 B.n656 163.367
R581 B.n656 B.n33 163.367
R582 B.n652 B.n33 163.367
R583 B.n652 B.n651 163.367
R584 B.n651 B.n650 163.367
R585 B.n650 B.n35 163.367
R586 B.n646 B.n35 163.367
R587 B.n646 B.n645 163.367
R588 B.n645 B.n644 163.367
R589 B.n644 B.n37 163.367
R590 B.n640 B.n37 163.367
R591 B.n640 B.n639 163.367
R592 B.n639 B.n638 163.367
R593 B.n638 B.n39 163.367
R594 B.n634 B.n39 163.367
R595 B.n634 B.n633 163.367
R596 B.n633 B.n632 163.367
R597 B.n632 B.n41 163.367
R598 B.n628 B.n41 163.367
R599 B.n628 B.n627 163.367
R600 B.n627 B.n626 163.367
R601 B.n626 B.n43 163.367
R602 B.n622 B.n43 163.367
R603 B.n622 B.n621 163.367
R604 B.n621 B.n620 163.367
R605 B.n620 B.n45 163.367
R606 B.n615 B.n45 163.367
R607 B.n615 B.n614 163.367
R608 B.n614 B.n613 163.367
R609 B.n613 B.n49 163.367
R610 B.n609 B.n49 163.367
R611 B.n609 B.n608 163.367
R612 B.n608 B.n607 163.367
R613 B.n607 B.n51 163.367
R614 B.n603 B.n51 163.367
R615 B.n603 B.n602 163.367
R616 B.n602 B.n55 163.367
R617 B.n598 B.n55 163.367
R618 B.n598 B.n597 163.367
R619 B.n597 B.n596 163.367
R620 B.n596 B.n57 163.367
R621 B.n592 B.n57 163.367
R622 B.n592 B.n591 163.367
R623 B.n591 B.n590 163.367
R624 B.n590 B.n59 163.367
R625 B.n586 B.n59 163.367
R626 B.n586 B.n585 163.367
R627 B.n585 B.n584 163.367
R628 B.n584 B.n61 163.367
R629 B.n580 B.n61 163.367
R630 B.n580 B.n579 163.367
R631 B.n579 B.n578 163.367
R632 B.n578 B.n63 163.367
R633 B.n574 B.n63 163.367
R634 B.n574 B.n573 163.367
R635 B.n573 B.n572 163.367
R636 B.n572 B.n65 163.367
R637 B.n568 B.n65 163.367
R638 B.n568 B.n567 163.367
R639 B.n567 B.n566 163.367
R640 B.n566 B.n67 163.367
R641 B.n562 B.n67 163.367
R642 B.n562 B.n561 163.367
R643 B.n561 B.n560 163.367
R644 B.n560 B.n69 163.367
R645 B.n556 B.n69 163.367
R646 B.n556 B.n555 163.367
R647 B.n555 B.n554 163.367
R648 B.n554 B.n71 163.367
R649 B.n550 B.n71 163.367
R650 B.n550 B.n549 163.367
R651 B.n549 B.n548 163.367
R652 B.n548 B.n73 163.367
R653 B.n544 B.n73 163.367
R654 B.n544 B.n543 163.367
R655 B.n543 B.n542 163.367
R656 B.n681 B.n680 163.367
R657 B.n682 B.n681 163.367
R658 B.n682 B.n23 163.367
R659 B.n686 B.n23 163.367
R660 B.n687 B.n686 163.367
R661 B.n688 B.n687 163.367
R662 B.n688 B.n21 163.367
R663 B.n692 B.n21 163.367
R664 B.n693 B.n692 163.367
R665 B.n694 B.n693 163.367
R666 B.n694 B.n19 163.367
R667 B.n698 B.n19 163.367
R668 B.n699 B.n698 163.367
R669 B.n700 B.n699 163.367
R670 B.n700 B.n17 163.367
R671 B.n704 B.n17 163.367
R672 B.n705 B.n704 163.367
R673 B.n706 B.n705 163.367
R674 B.n706 B.n15 163.367
R675 B.n710 B.n15 163.367
R676 B.n711 B.n710 163.367
R677 B.n712 B.n711 163.367
R678 B.n712 B.n13 163.367
R679 B.n716 B.n13 163.367
R680 B.n717 B.n716 163.367
R681 B.n718 B.n717 163.367
R682 B.n718 B.n11 163.367
R683 B.n722 B.n11 163.367
R684 B.n723 B.n722 163.367
R685 B.n724 B.n723 163.367
R686 B.n724 B.n9 163.367
R687 B.n728 B.n9 163.367
R688 B.n729 B.n728 163.367
R689 B.n730 B.n729 163.367
R690 B.n730 B.n7 163.367
R691 B.n734 B.n7 163.367
R692 B.n735 B.n734 163.367
R693 B.n736 B.n735 163.367
R694 B.n736 B.n5 163.367
R695 B.n740 B.n5 163.367
R696 B.n741 B.n740 163.367
R697 B.n742 B.n741 163.367
R698 B.n742 B.n3 163.367
R699 B.n746 B.n3 163.367
R700 B.n747 B.n746 163.367
R701 B.n192 B.n2 163.367
R702 B.n192 B.n191 163.367
R703 B.n196 B.n191 163.367
R704 B.n197 B.n196 163.367
R705 B.n198 B.n197 163.367
R706 B.n198 B.n189 163.367
R707 B.n202 B.n189 163.367
R708 B.n203 B.n202 163.367
R709 B.n204 B.n203 163.367
R710 B.n204 B.n187 163.367
R711 B.n208 B.n187 163.367
R712 B.n209 B.n208 163.367
R713 B.n210 B.n209 163.367
R714 B.n210 B.n185 163.367
R715 B.n214 B.n185 163.367
R716 B.n215 B.n214 163.367
R717 B.n216 B.n215 163.367
R718 B.n216 B.n183 163.367
R719 B.n220 B.n183 163.367
R720 B.n221 B.n220 163.367
R721 B.n222 B.n221 163.367
R722 B.n222 B.n181 163.367
R723 B.n226 B.n181 163.367
R724 B.n227 B.n226 163.367
R725 B.n228 B.n227 163.367
R726 B.n228 B.n179 163.367
R727 B.n232 B.n179 163.367
R728 B.n233 B.n232 163.367
R729 B.n234 B.n233 163.367
R730 B.n234 B.n177 163.367
R731 B.n238 B.n177 163.367
R732 B.n239 B.n238 163.367
R733 B.n240 B.n239 163.367
R734 B.n240 B.n175 163.367
R735 B.n244 B.n175 163.367
R736 B.n245 B.n244 163.367
R737 B.n246 B.n245 163.367
R738 B.n246 B.n173 163.367
R739 B.n250 B.n173 163.367
R740 B.n251 B.n250 163.367
R741 B.n252 B.n251 163.367
R742 B.n252 B.n171 163.367
R743 B.n256 B.n171 163.367
R744 B.n257 B.n256 163.367
R745 B.n258 B.n257 163.367
R746 B.n335 B.t5 110.466
R747 B.n53 B.t10 110.466
R748 B.n149 B.t2 110.451
R749 B.n47 B.t7 110.451
R750 B.n149 B.n148 63.6126
R751 B.n335 B.n334 63.6126
R752 B.n53 B.n52 63.6126
R753 B.n47 B.n46 63.6126
R754 B.n321 B.n149 59.5399
R755 B.n336 B.n335 59.5399
R756 B.n54 B.n53 59.5399
R757 B.n617 B.n47 59.5399
R758 B.n401 B.n122 35.7468
R759 B.n679 B.n678 35.7468
R760 B.n541 B.n540 35.7468
R761 B.n260 B.n259 35.7468
R762 B B.n749 18.0485
R763 B.n679 B.n24 10.6151
R764 B.n683 B.n24 10.6151
R765 B.n684 B.n683 10.6151
R766 B.n685 B.n684 10.6151
R767 B.n685 B.n22 10.6151
R768 B.n689 B.n22 10.6151
R769 B.n690 B.n689 10.6151
R770 B.n691 B.n690 10.6151
R771 B.n691 B.n20 10.6151
R772 B.n695 B.n20 10.6151
R773 B.n696 B.n695 10.6151
R774 B.n697 B.n696 10.6151
R775 B.n697 B.n18 10.6151
R776 B.n701 B.n18 10.6151
R777 B.n702 B.n701 10.6151
R778 B.n703 B.n702 10.6151
R779 B.n703 B.n16 10.6151
R780 B.n707 B.n16 10.6151
R781 B.n708 B.n707 10.6151
R782 B.n709 B.n708 10.6151
R783 B.n709 B.n14 10.6151
R784 B.n713 B.n14 10.6151
R785 B.n714 B.n713 10.6151
R786 B.n715 B.n714 10.6151
R787 B.n715 B.n12 10.6151
R788 B.n719 B.n12 10.6151
R789 B.n720 B.n719 10.6151
R790 B.n721 B.n720 10.6151
R791 B.n721 B.n10 10.6151
R792 B.n725 B.n10 10.6151
R793 B.n726 B.n725 10.6151
R794 B.n727 B.n726 10.6151
R795 B.n727 B.n8 10.6151
R796 B.n731 B.n8 10.6151
R797 B.n732 B.n731 10.6151
R798 B.n733 B.n732 10.6151
R799 B.n733 B.n6 10.6151
R800 B.n737 B.n6 10.6151
R801 B.n738 B.n737 10.6151
R802 B.n739 B.n738 10.6151
R803 B.n739 B.n4 10.6151
R804 B.n743 B.n4 10.6151
R805 B.n744 B.n743 10.6151
R806 B.n745 B.n744 10.6151
R807 B.n745 B.n0 10.6151
R808 B.n678 B.n677 10.6151
R809 B.n677 B.n26 10.6151
R810 B.n673 B.n26 10.6151
R811 B.n673 B.n672 10.6151
R812 B.n672 B.n671 10.6151
R813 B.n671 B.n28 10.6151
R814 B.n667 B.n28 10.6151
R815 B.n667 B.n666 10.6151
R816 B.n666 B.n665 10.6151
R817 B.n665 B.n30 10.6151
R818 B.n661 B.n30 10.6151
R819 B.n661 B.n660 10.6151
R820 B.n660 B.n659 10.6151
R821 B.n659 B.n32 10.6151
R822 B.n655 B.n32 10.6151
R823 B.n655 B.n654 10.6151
R824 B.n654 B.n653 10.6151
R825 B.n653 B.n34 10.6151
R826 B.n649 B.n34 10.6151
R827 B.n649 B.n648 10.6151
R828 B.n648 B.n647 10.6151
R829 B.n647 B.n36 10.6151
R830 B.n643 B.n36 10.6151
R831 B.n643 B.n642 10.6151
R832 B.n642 B.n641 10.6151
R833 B.n641 B.n38 10.6151
R834 B.n637 B.n38 10.6151
R835 B.n637 B.n636 10.6151
R836 B.n636 B.n635 10.6151
R837 B.n635 B.n40 10.6151
R838 B.n631 B.n40 10.6151
R839 B.n631 B.n630 10.6151
R840 B.n630 B.n629 10.6151
R841 B.n629 B.n42 10.6151
R842 B.n625 B.n42 10.6151
R843 B.n625 B.n624 10.6151
R844 B.n624 B.n623 10.6151
R845 B.n623 B.n44 10.6151
R846 B.n619 B.n44 10.6151
R847 B.n619 B.n618 10.6151
R848 B.n616 B.n48 10.6151
R849 B.n612 B.n48 10.6151
R850 B.n612 B.n611 10.6151
R851 B.n611 B.n610 10.6151
R852 B.n610 B.n50 10.6151
R853 B.n606 B.n50 10.6151
R854 B.n606 B.n605 10.6151
R855 B.n605 B.n604 10.6151
R856 B.n601 B.n600 10.6151
R857 B.n600 B.n599 10.6151
R858 B.n599 B.n56 10.6151
R859 B.n595 B.n56 10.6151
R860 B.n595 B.n594 10.6151
R861 B.n594 B.n593 10.6151
R862 B.n593 B.n58 10.6151
R863 B.n589 B.n58 10.6151
R864 B.n589 B.n588 10.6151
R865 B.n588 B.n587 10.6151
R866 B.n587 B.n60 10.6151
R867 B.n583 B.n60 10.6151
R868 B.n583 B.n582 10.6151
R869 B.n582 B.n581 10.6151
R870 B.n581 B.n62 10.6151
R871 B.n577 B.n62 10.6151
R872 B.n577 B.n576 10.6151
R873 B.n576 B.n575 10.6151
R874 B.n575 B.n64 10.6151
R875 B.n571 B.n64 10.6151
R876 B.n571 B.n570 10.6151
R877 B.n570 B.n569 10.6151
R878 B.n569 B.n66 10.6151
R879 B.n565 B.n66 10.6151
R880 B.n565 B.n564 10.6151
R881 B.n564 B.n563 10.6151
R882 B.n563 B.n68 10.6151
R883 B.n559 B.n68 10.6151
R884 B.n559 B.n558 10.6151
R885 B.n558 B.n557 10.6151
R886 B.n557 B.n70 10.6151
R887 B.n553 B.n70 10.6151
R888 B.n553 B.n552 10.6151
R889 B.n552 B.n551 10.6151
R890 B.n551 B.n72 10.6151
R891 B.n547 B.n72 10.6151
R892 B.n547 B.n546 10.6151
R893 B.n546 B.n545 10.6151
R894 B.n545 B.n74 10.6151
R895 B.n541 B.n74 10.6151
R896 B.n540 B.n539 10.6151
R897 B.n539 B.n76 10.6151
R898 B.n535 B.n76 10.6151
R899 B.n535 B.n534 10.6151
R900 B.n534 B.n533 10.6151
R901 B.n533 B.n78 10.6151
R902 B.n529 B.n78 10.6151
R903 B.n529 B.n528 10.6151
R904 B.n528 B.n527 10.6151
R905 B.n527 B.n80 10.6151
R906 B.n523 B.n80 10.6151
R907 B.n523 B.n522 10.6151
R908 B.n522 B.n521 10.6151
R909 B.n521 B.n82 10.6151
R910 B.n517 B.n82 10.6151
R911 B.n517 B.n516 10.6151
R912 B.n516 B.n515 10.6151
R913 B.n515 B.n84 10.6151
R914 B.n511 B.n84 10.6151
R915 B.n511 B.n510 10.6151
R916 B.n510 B.n509 10.6151
R917 B.n509 B.n86 10.6151
R918 B.n505 B.n86 10.6151
R919 B.n505 B.n504 10.6151
R920 B.n504 B.n503 10.6151
R921 B.n503 B.n88 10.6151
R922 B.n499 B.n88 10.6151
R923 B.n499 B.n498 10.6151
R924 B.n498 B.n497 10.6151
R925 B.n497 B.n90 10.6151
R926 B.n493 B.n90 10.6151
R927 B.n493 B.n492 10.6151
R928 B.n492 B.n491 10.6151
R929 B.n491 B.n92 10.6151
R930 B.n487 B.n92 10.6151
R931 B.n487 B.n486 10.6151
R932 B.n486 B.n485 10.6151
R933 B.n485 B.n94 10.6151
R934 B.n481 B.n94 10.6151
R935 B.n481 B.n480 10.6151
R936 B.n480 B.n479 10.6151
R937 B.n479 B.n96 10.6151
R938 B.n475 B.n96 10.6151
R939 B.n475 B.n474 10.6151
R940 B.n474 B.n473 10.6151
R941 B.n473 B.n98 10.6151
R942 B.n469 B.n98 10.6151
R943 B.n469 B.n468 10.6151
R944 B.n468 B.n467 10.6151
R945 B.n467 B.n100 10.6151
R946 B.n463 B.n100 10.6151
R947 B.n463 B.n462 10.6151
R948 B.n462 B.n461 10.6151
R949 B.n461 B.n102 10.6151
R950 B.n457 B.n102 10.6151
R951 B.n457 B.n456 10.6151
R952 B.n456 B.n455 10.6151
R953 B.n455 B.n104 10.6151
R954 B.n451 B.n104 10.6151
R955 B.n451 B.n450 10.6151
R956 B.n450 B.n449 10.6151
R957 B.n449 B.n106 10.6151
R958 B.n445 B.n106 10.6151
R959 B.n445 B.n444 10.6151
R960 B.n444 B.n443 10.6151
R961 B.n443 B.n108 10.6151
R962 B.n439 B.n108 10.6151
R963 B.n439 B.n438 10.6151
R964 B.n438 B.n437 10.6151
R965 B.n437 B.n110 10.6151
R966 B.n433 B.n110 10.6151
R967 B.n433 B.n432 10.6151
R968 B.n432 B.n431 10.6151
R969 B.n431 B.n112 10.6151
R970 B.n427 B.n112 10.6151
R971 B.n427 B.n426 10.6151
R972 B.n426 B.n425 10.6151
R973 B.n425 B.n114 10.6151
R974 B.n421 B.n114 10.6151
R975 B.n421 B.n420 10.6151
R976 B.n420 B.n419 10.6151
R977 B.n419 B.n116 10.6151
R978 B.n415 B.n116 10.6151
R979 B.n415 B.n414 10.6151
R980 B.n414 B.n413 10.6151
R981 B.n413 B.n118 10.6151
R982 B.n409 B.n118 10.6151
R983 B.n409 B.n408 10.6151
R984 B.n408 B.n407 10.6151
R985 B.n407 B.n120 10.6151
R986 B.n403 B.n120 10.6151
R987 B.n403 B.n402 10.6151
R988 B.n402 B.n401 10.6151
R989 B.n193 B.n1 10.6151
R990 B.n194 B.n193 10.6151
R991 B.n195 B.n194 10.6151
R992 B.n195 B.n190 10.6151
R993 B.n199 B.n190 10.6151
R994 B.n200 B.n199 10.6151
R995 B.n201 B.n200 10.6151
R996 B.n201 B.n188 10.6151
R997 B.n205 B.n188 10.6151
R998 B.n206 B.n205 10.6151
R999 B.n207 B.n206 10.6151
R1000 B.n207 B.n186 10.6151
R1001 B.n211 B.n186 10.6151
R1002 B.n212 B.n211 10.6151
R1003 B.n213 B.n212 10.6151
R1004 B.n213 B.n184 10.6151
R1005 B.n217 B.n184 10.6151
R1006 B.n218 B.n217 10.6151
R1007 B.n219 B.n218 10.6151
R1008 B.n219 B.n182 10.6151
R1009 B.n223 B.n182 10.6151
R1010 B.n224 B.n223 10.6151
R1011 B.n225 B.n224 10.6151
R1012 B.n225 B.n180 10.6151
R1013 B.n229 B.n180 10.6151
R1014 B.n230 B.n229 10.6151
R1015 B.n231 B.n230 10.6151
R1016 B.n231 B.n178 10.6151
R1017 B.n235 B.n178 10.6151
R1018 B.n236 B.n235 10.6151
R1019 B.n237 B.n236 10.6151
R1020 B.n237 B.n176 10.6151
R1021 B.n241 B.n176 10.6151
R1022 B.n242 B.n241 10.6151
R1023 B.n243 B.n242 10.6151
R1024 B.n243 B.n174 10.6151
R1025 B.n247 B.n174 10.6151
R1026 B.n248 B.n247 10.6151
R1027 B.n249 B.n248 10.6151
R1028 B.n249 B.n172 10.6151
R1029 B.n253 B.n172 10.6151
R1030 B.n254 B.n253 10.6151
R1031 B.n255 B.n254 10.6151
R1032 B.n255 B.n170 10.6151
R1033 B.n259 B.n170 10.6151
R1034 B.n261 B.n260 10.6151
R1035 B.n261 B.n168 10.6151
R1036 B.n265 B.n168 10.6151
R1037 B.n266 B.n265 10.6151
R1038 B.n267 B.n266 10.6151
R1039 B.n267 B.n166 10.6151
R1040 B.n271 B.n166 10.6151
R1041 B.n272 B.n271 10.6151
R1042 B.n273 B.n272 10.6151
R1043 B.n273 B.n164 10.6151
R1044 B.n277 B.n164 10.6151
R1045 B.n278 B.n277 10.6151
R1046 B.n279 B.n278 10.6151
R1047 B.n279 B.n162 10.6151
R1048 B.n283 B.n162 10.6151
R1049 B.n284 B.n283 10.6151
R1050 B.n285 B.n284 10.6151
R1051 B.n285 B.n160 10.6151
R1052 B.n289 B.n160 10.6151
R1053 B.n290 B.n289 10.6151
R1054 B.n291 B.n290 10.6151
R1055 B.n291 B.n158 10.6151
R1056 B.n295 B.n158 10.6151
R1057 B.n296 B.n295 10.6151
R1058 B.n297 B.n296 10.6151
R1059 B.n297 B.n156 10.6151
R1060 B.n301 B.n156 10.6151
R1061 B.n302 B.n301 10.6151
R1062 B.n303 B.n302 10.6151
R1063 B.n303 B.n154 10.6151
R1064 B.n307 B.n154 10.6151
R1065 B.n308 B.n307 10.6151
R1066 B.n309 B.n308 10.6151
R1067 B.n309 B.n152 10.6151
R1068 B.n313 B.n152 10.6151
R1069 B.n314 B.n313 10.6151
R1070 B.n315 B.n314 10.6151
R1071 B.n315 B.n150 10.6151
R1072 B.n319 B.n150 10.6151
R1073 B.n320 B.n319 10.6151
R1074 B.n322 B.n146 10.6151
R1075 B.n326 B.n146 10.6151
R1076 B.n327 B.n326 10.6151
R1077 B.n328 B.n327 10.6151
R1078 B.n328 B.n144 10.6151
R1079 B.n332 B.n144 10.6151
R1080 B.n333 B.n332 10.6151
R1081 B.n337 B.n333 10.6151
R1082 B.n341 B.n142 10.6151
R1083 B.n342 B.n341 10.6151
R1084 B.n343 B.n342 10.6151
R1085 B.n343 B.n140 10.6151
R1086 B.n347 B.n140 10.6151
R1087 B.n348 B.n347 10.6151
R1088 B.n349 B.n348 10.6151
R1089 B.n349 B.n138 10.6151
R1090 B.n353 B.n138 10.6151
R1091 B.n354 B.n353 10.6151
R1092 B.n355 B.n354 10.6151
R1093 B.n355 B.n136 10.6151
R1094 B.n359 B.n136 10.6151
R1095 B.n360 B.n359 10.6151
R1096 B.n361 B.n360 10.6151
R1097 B.n361 B.n134 10.6151
R1098 B.n365 B.n134 10.6151
R1099 B.n366 B.n365 10.6151
R1100 B.n367 B.n366 10.6151
R1101 B.n367 B.n132 10.6151
R1102 B.n371 B.n132 10.6151
R1103 B.n372 B.n371 10.6151
R1104 B.n373 B.n372 10.6151
R1105 B.n373 B.n130 10.6151
R1106 B.n377 B.n130 10.6151
R1107 B.n378 B.n377 10.6151
R1108 B.n379 B.n378 10.6151
R1109 B.n379 B.n128 10.6151
R1110 B.n383 B.n128 10.6151
R1111 B.n384 B.n383 10.6151
R1112 B.n385 B.n384 10.6151
R1113 B.n385 B.n126 10.6151
R1114 B.n389 B.n126 10.6151
R1115 B.n390 B.n389 10.6151
R1116 B.n391 B.n390 10.6151
R1117 B.n391 B.n124 10.6151
R1118 B.n395 B.n124 10.6151
R1119 B.n396 B.n395 10.6151
R1120 B.n397 B.n396 10.6151
R1121 B.n397 B.n122 10.6151
R1122 B.n749 B.n0 8.11757
R1123 B.n749 B.n1 8.11757
R1124 B.n617 B.n616 6.5566
R1125 B.n604 B.n54 6.5566
R1126 B.n322 B.n321 6.5566
R1127 B.n337 B.n336 6.5566
R1128 B.n618 B.n617 4.05904
R1129 B.n601 B.n54 4.05904
R1130 B.n321 B.n320 4.05904
R1131 B.n336 B.n142 4.05904
R1132 VN.n33 VN.n18 161.3
R1133 VN.n32 VN.n31 161.3
R1134 VN.n30 VN.n19 161.3
R1135 VN.n29 VN.n28 161.3
R1136 VN.n27 VN.n20 161.3
R1137 VN.n26 VN.n25 161.3
R1138 VN.n24 VN.n21 161.3
R1139 VN.n15 VN.n0 161.3
R1140 VN.n14 VN.n13 161.3
R1141 VN.n12 VN.n1 161.3
R1142 VN.n11 VN.n10 161.3
R1143 VN.n9 VN.n2 161.3
R1144 VN.n8 VN.n7 161.3
R1145 VN.n6 VN.n3 161.3
R1146 VN.n5 VN.t5 128.292
R1147 VN.n23 VN.t1 128.292
R1148 VN.n17 VN.n16 109.288
R1149 VN.n35 VN.n34 109.288
R1150 VN.n4 VN.t0 95.8286
R1151 VN.n16 VN.t3 95.8286
R1152 VN.n22 VN.t2 95.8286
R1153 VN.n34 VN.t4 95.8286
R1154 VN.n5 VN.n4 61.6325
R1155 VN.n23 VN.n22 61.6325
R1156 VN.n10 VN.n9 51.1773
R1157 VN.n28 VN.n27 51.1773
R1158 VN VN.n35 50.0966
R1159 VN.n10 VN.n1 29.8095
R1160 VN.n28 VN.n19 29.8095
R1161 VN.n8 VN.n3 24.4675
R1162 VN.n9 VN.n8 24.4675
R1163 VN.n14 VN.n1 24.4675
R1164 VN.n15 VN.n14 24.4675
R1165 VN.n27 VN.n26 24.4675
R1166 VN.n26 VN.n21 24.4675
R1167 VN.n33 VN.n32 24.4675
R1168 VN.n32 VN.n19 24.4675
R1169 VN.n4 VN.n3 12.234
R1170 VN.n22 VN.n21 12.234
R1171 VN.n24 VN.n23 5.14959
R1172 VN.n6 VN.n5 5.14959
R1173 VN.n16 VN.n15 1.46852
R1174 VN.n34 VN.n33 1.46852
R1175 VN.n35 VN.n18 0.278367
R1176 VN.n17 VN.n0 0.278367
R1177 VN.n31 VN.n18 0.189894
R1178 VN.n31 VN.n30 0.189894
R1179 VN.n30 VN.n29 0.189894
R1180 VN.n29 VN.n20 0.189894
R1181 VN.n25 VN.n20 0.189894
R1182 VN.n25 VN.n24 0.189894
R1183 VN.n7 VN.n6 0.189894
R1184 VN.n7 VN.n2 0.189894
R1185 VN.n11 VN.n2 0.189894
R1186 VN.n12 VN.n11 0.189894
R1187 VN.n13 VN.n12 0.189894
R1188 VN.n13 VN.n0 0.189894
R1189 VN VN.n17 0.153454
R1190 VDD2.n1 VDD2.t4 78.5493
R1191 VDD2.n2 VDD2.t1 76.4842
R1192 VDD2.n1 VDD2.n0 74.3644
R1193 VDD2 VDD2.n3 74.3616
R1194 VDD2.n2 VDD2.n1 43.017
R1195 VDD2.n3 VDD2.t5 2.7716
R1196 VDD2.n3 VDD2.t3 2.7716
R1197 VDD2.n0 VDD2.t0 2.7716
R1198 VDD2.n0 VDD2.t2 2.7716
R1199 VDD2 VDD2.n2 2.17938
R1200 VTAIL.n7 VTAIL.t10 59.8054
R1201 VTAIL.n11 VTAIL.t8 59.8052
R1202 VTAIL.n2 VTAIL.t4 59.8052
R1203 VTAIL.n10 VTAIL.t2 59.8052
R1204 VTAIL.n9 VTAIL.n8 57.0343
R1205 VTAIL.n6 VTAIL.n5 57.0343
R1206 VTAIL.n1 VTAIL.n0 57.0341
R1207 VTAIL.n4 VTAIL.n3 57.0341
R1208 VTAIL.n6 VTAIL.n4 28.1341
R1209 VTAIL.n11 VTAIL.n10 25.3065
R1210 VTAIL.n7 VTAIL.n6 2.82809
R1211 VTAIL.n10 VTAIL.n9 2.82809
R1212 VTAIL.n4 VTAIL.n2 2.82809
R1213 VTAIL.n0 VTAIL.t6 2.7716
R1214 VTAIL.n0 VTAIL.t11 2.7716
R1215 VTAIL.n3 VTAIL.t0 2.7716
R1216 VTAIL.n3 VTAIL.t3 2.7716
R1217 VTAIL.n8 VTAIL.t5 2.7716
R1218 VTAIL.n8 VTAIL.t1 2.7716
R1219 VTAIL.n5 VTAIL.t7 2.7716
R1220 VTAIL.n5 VTAIL.t9 2.7716
R1221 VTAIL VTAIL.n11 2.063
R1222 VTAIL.n9 VTAIL.n7 1.88412
R1223 VTAIL.n2 VTAIL.n1 1.88412
R1224 VTAIL VTAIL.n1 0.765586
R1225 VP.n14 VP.n11 161.3
R1226 VP.n16 VP.n15 161.3
R1227 VP.n17 VP.n10 161.3
R1228 VP.n19 VP.n18 161.3
R1229 VP.n20 VP.n9 161.3
R1230 VP.n22 VP.n21 161.3
R1231 VP.n23 VP.n8 161.3
R1232 VP.n48 VP.n0 161.3
R1233 VP.n47 VP.n46 161.3
R1234 VP.n45 VP.n1 161.3
R1235 VP.n44 VP.n43 161.3
R1236 VP.n42 VP.n2 161.3
R1237 VP.n41 VP.n40 161.3
R1238 VP.n39 VP.n3 161.3
R1239 VP.n38 VP.n37 161.3
R1240 VP.n35 VP.n4 161.3
R1241 VP.n34 VP.n33 161.3
R1242 VP.n32 VP.n5 161.3
R1243 VP.n31 VP.n30 161.3
R1244 VP.n29 VP.n6 161.3
R1245 VP.n28 VP.n27 161.3
R1246 VP.n13 VP.t4 128.292
R1247 VP.n26 VP.n7 109.288
R1248 VP.n50 VP.n49 109.288
R1249 VP.n25 VP.n24 109.288
R1250 VP.n7 VP.t1 95.8286
R1251 VP.n36 VP.t0 95.8286
R1252 VP.n49 VP.t5 95.8286
R1253 VP.n24 VP.t2 95.8286
R1254 VP.n12 VP.t3 95.8286
R1255 VP.n13 VP.n12 61.6325
R1256 VP.n34 VP.n5 51.1773
R1257 VP.n43 VP.n42 51.1773
R1258 VP.n18 VP.n17 51.1773
R1259 VP.n26 VP.n25 49.8178
R1260 VP.n30 VP.n5 29.8095
R1261 VP.n43 VP.n1 29.8095
R1262 VP.n18 VP.n9 29.8095
R1263 VP.n29 VP.n28 24.4675
R1264 VP.n30 VP.n29 24.4675
R1265 VP.n35 VP.n34 24.4675
R1266 VP.n37 VP.n35 24.4675
R1267 VP.n41 VP.n3 24.4675
R1268 VP.n42 VP.n41 24.4675
R1269 VP.n47 VP.n1 24.4675
R1270 VP.n48 VP.n47 24.4675
R1271 VP.n22 VP.n9 24.4675
R1272 VP.n23 VP.n22 24.4675
R1273 VP.n16 VP.n11 24.4675
R1274 VP.n17 VP.n16 24.4675
R1275 VP.n37 VP.n36 12.234
R1276 VP.n36 VP.n3 12.234
R1277 VP.n12 VP.n11 12.234
R1278 VP.n14 VP.n13 5.14959
R1279 VP.n28 VP.n7 1.46852
R1280 VP.n49 VP.n48 1.46852
R1281 VP.n24 VP.n23 1.46852
R1282 VP.n25 VP.n8 0.278367
R1283 VP.n27 VP.n26 0.278367
R1284 VP.n50 VP.n0 0.278367
R1285 VP.n15 VP.n14 0.189894
R1286 VP.n15 VP.n10 0.189894
R1287 VP.n19 VP.n10 0.189894
R1288 VP.n20 VP.n19 0.189894
R1289 VP.n21 VP.n20 0.189894
R1290 VP.n21 VP.n8 0.189894
R1291 VP.n27 VP.n6 0.189894
R1292 VP.n31 VP.n6 0.189894
R1293 VP.n32 VP.n31 0.189894
R1294 VP.n33 VP.n32 0.189894
R1295 VP.n33 VP.n4 0.189894
R1296 VP.n38 VP.n4 0.189894
R1297 VP.n39 VP.n38 0.189894
R1298 VP.n40 VP.n39 0.189894
R1299 VP.n40 VP.n2 0.189894
R1300 VP.n44 VP.n2 0.189894
R1301 VP.n45 VP.n44 0.189894
R1302 VP.n46 VP.n45 0.189894
R1303 VP.n46 VP.n0 0.189894
R1304 VP VP.n50 0.153454
R1305 VDD1 VDD1.t1 78.6631
R1306 VDD1.n1 VDD1.t4 78.5493
R1307 VDD1.n1 VDD1.n0 74.3644
R1308 VDD1.n3 VDD1.n2 73.7129
R1309 VDD1.n3 VDD1.n1 45.0138
R1310 VDD1.n2 VDD1.t2 2.7716
R1311 VDD1.n2 VDD1.t3 2.7716
R1312 VDD1.n0 VDD1.t5 2.7716
R1313 VDD1.n0 VDD1.t0 2.7716
R1314 VDD1 VDD1.n3 0.649207
C0 VP VTAIL 7.00361f
C1 VP w_n3594_n3314# 7.3505f
C2 VDD1 VDD2 1.54329f
C3 VTAIL B 3.77068f
C4 w_n3594_n3314# B 10.084f
C5 VDD1 VN 0.151198f
C6 VP VDD2 0.487953f
C7 VDD2 B 2.24578f
C8 VTAIL w_n3594_n3314# 2.96553f
C9 VP VN 7.21583f
C10 VN B 1.2378f
C11 VTAIL VDD2 7.773049f
C12 VDD2 w_n3594_n3314# 2.45356f
C13 VTAIL VN 6.98935f
C14 VN w_n3594_n3314# 6.88487f
C15 VN VDD2 6.73234f
C16 VP VDD1 7.06602f
C17 VDD1 B 2.16329f
C18 VP B 2.01698f
C19 VTAIL VDD1 7.719471f
C20 VDD1 w_n3594_n3314# 2.35732f
C21 VDD2 VSUBS 2.002128f
C22 VDD1 VSUBS 2.51771f
C23 VTAIL VSUBS 1.255185f
C24 VN VSUBS 6.14347f
C25 VP VSUBS 3.1893f
C26 B VSUBS 4.962228f
C27 w_n3594_n3314# VSUBS 0.146678p
C28 VDD1.t1 VSUBS 2.69741f
C29 VDD1.t4 VSUBS 2.69596f
C30 VDD1.t5 VSUBS 0.263581f
C31 VDD1.t0 VSUBS 0.263581f
C32 VDD1.n0 VSUBS 2.0536f
C33 VDD1.n1 VSUBS 4.2187f
C34 VDD1.t2 VSUBS 0.263581f
C35 VDD1.t3 VSUBS 0.263581f
C36 VDD1.n2 VSUBS 2.04601f
C37 VDD1.n3 VSUBS 3.56201f
C38 VP.n0 VSUBS 0.041739f
C39 VP.t5 VSUBS 2.98289f
C40 VP.n1 VSUBS 0.063074f
C41 VP.n2 VSUBS 0.031659f
C42 VP.n3 VSUBS 0.044439f
C43 VP.n4 VSUBS 0.031659f
C44 VP.n5 VSUBS 0.030881f
C45 VP.n6 VSUBS 0.031659f
C46 VP.t1 VSUBS 2.98289f
C47 VP.n7 VSUBS 1.15854f
C48 VP.n8 VSUBS 0.041739f
C49 VP.t2 VSUBS 2.98289f
C50 VP.n9 VSUBS 0.063074f
C51 VP.n10 VSUBS 0.031659f
C52 VP.n11 VSUBS 0.044439f
C53 VP.t4 VSUBS 3.30422f
C54 VP.t3 VSUBS 2.98289f
C55 VP.n12 VSUBS 1.15228f
C56 VP.n13 VSUBS 1.11182f
C57 VP.n14 VSUBS 0.337611f
C58 VP.n15 VSUBS 0.031659f
C59 VP.n16 VSUBS 0.059004f
C60 VP.n17 VSUBS 0.057481f
C61 VP.n18 VSUBS 0.030881f
C62 VP.n19 VSUBS 0.031659f
C63 VP.n20 VSUBS 0.031659f
C64 VP.n21 VSUBS 0.031659f
C65 VP.n22 VSUBS 0.059004f
C66 VP.n23 VSUBS 0.031621f
C67 VP.n24 VSUBS 1.15854f
C68 VP.n25 VSUBS 1.76279f
C69 VP.n26 VSUBS 1.78564f
C70 VP.n27 VSUBS 0.041739f
C71 VP.n28 VSUBS 0.031621f
C72 VP.n29 VSUBS 0.059004f
C73 VP.n30 VSUBS 0.063074f
C74 VP.n31 VSUBS 0.031659f
C75 VP.n32 VSUBS 0.031659f
C76 VP.n33 VSUBS 0.031659f
C77 VP.n34 VSUBS 0.057481f
C78 VP.n35 VSUBS 0.059004f
C79 VP.t0 VSUBS 2.98289f
C80 VP.n36 VSUBS 1.05251f
C81 VP.n37 VSUBS 0.044439f
C82 VP.n38 VSUBS 0.031659f
C83 VP.n39 VSUBS 0.031659f
C84 VP.n40 VSUBS 0.031659f
C85 VP.n41 VSUBS 0.059004f
C86 VP.n42 VSUBS 0.057481f
C87 VP.n43 VSUBS 0.030881f
C88 VP.n44 VSUBS 0.031659f
C89 VP.n45 VSUBS 0.031659f
C90 VP.n46 VSUBS 0.031659f
C91 VP.n47 VSUBS 0.059004f
C92 VP.n48 VSUBS 0.031621f
C93 VP.n49 VSUBS 1.15854f
C94 VP.n50 VSUBS 0.061948f
C95 VTAIL.t6 VSUBS 0.274261f
C96 VTAIL.t11 VSUBS 0.274261f
C97 VTAIL.n0 VSUBS 1.96796f
C98 VTAIL.n1 VSUBS 0.929264f
C99 VTAIL.t4 VSUBS 2.60281f
C100 VTAIL.n2 VSUBS 1.23904f
C101 VTAIL.t0 VSUBS 0.274261f
C102 VTAIL.t3 VSUBS 0.274261f
C103 VTAIL.n3 VSUBS 1.96796f
C104 VTAIL.n4 VSUBS 2.85146f
C105 VTAIL.t7 VSUBS 0.274261f
C106 VTAIL.t9 VSUBS 0.274261f
C107 VTAIL.n5 VSUBS 1.96797f
C108 VTAIL.n6 VSUBS 2.85145f
C109 VTAIL.t10 VSUBS 2.60282f
C110 VTAIL.n7 VSUBS 1.23903f
C111 VTAIL.t5 VSUBS 0.274261f
C112 VTAIL.t1 VSUBS 0.274261f
C113 VTAIL.n8 VSUBS 1.96797f
C114 VTAIL.n9 VSUBS 1.12589f
C115 VTAIL.t2 VSUBS 2.60281f
C116 VTAIL.n10 VSUBS 2.69502f
C117 VTAIL.t8 VSUBS 2.60281f
C118 VTAIL.n11 VSUBS 2.62207f
C119 VDD2.t4 VSUBS 2.68269f
C120 VDD2.t0 VSUBS 0.262284f
C121 VDD2.t2 VSUBS 0.262284f
C122 VDD2.n0 VSUBS 2.04349f
C123 VDD2.n1 VSUBS 4.0473f
C124 VDD2.t1 VSUBS 2.66109f
C125 VDD2.n2 VSUBS 3.56248f
C126 VDD2.t5 VSUBS 0.262284f
C127 VDD2.t3 VSUBS 0.262284f
C128 VDD2.n3 VSUBS 2.04344f
C129 VN.n0 VSUBS 0.037742f
C130 VN.t3 VSUBS 2.69721f
C131 VN.n1 VSUBS 0.057034f
C132 VN.n2 VSUBS 0.028627f
C133 VN.n3 VSUBS 0.040183f
C134 VN.t5 VSUBS 2.98776f
C135 VN.t0 VSUBS 2.69721f
C136 VN.n4 VSUBS 1.04192f
C137 VN.n5 VSUBS 1.00534f
C138 VN.n6 VSUBS 0.305276f
C139 VN.n7 VSUBS 0.028627f
C140 VN.n8 VSUBS 0.053353f
C141 VN.n9 VSUBS 0.051976f
C142 VN.n10 VSUBS 0.027924f
C143 VN.n11 VSUBS 0.028627f
C144 VN.n12 VSUBS 0.028627f
C145 VN.n13 VSUBS 0.028627f
C146 VN.n14 VSUBS 0.053353f
C147 VN.n15 VSUBS 0.028593f
C148 VN.n16 VSUBS 1.04758f
C149 VN.n17 VSUBS 0.056015f
C150 VN.n18 VSUBS 0.037742f
C151 VN.t4 VSUBS 2.69721f
C152 VN.n19 VSUBS 0.057034f
C153 VN.n20 VSUBS 0.028627f
C154 VN.n21 VSUBS 0.040183f
C155 VN.t1 VSUBS 2.98776f
C156 VN.t2 VSUBS 2.69721f
C157 VN.n22 VSUBS 1.04192f
C158 VN.n23 VSUBS 1.00534f
C159 VN.n24 VSUBS 0.305276f
C160 VN.n25 VSUBS 0.028627f
C161 VN.n26 VSUBS 0.053353f
C162 VN.n27 VSUBS 0.051976f
C163 VN.n28 VSUBS 0.027924f
C164 VN.n29 VSUBS 0.028627f
C165 VN.n30 VSUBS 0.028627f
C166 VN.n31 VSUBS 0.028627f
C167 VN.n32 VSUBS 0.053353f
C168 VN.n33 VSUBS 0.028593f
C169 VN.n34 VSUBS 1.04758f
C170 VN.n35 VSUBS 1.60935f
C171 B.n0 VSUBS 0.007794f
C172 B.n1 VSUBS 0.007794f
C173 B.n2 VSUBS 0.011527f
C174 B.n3 VSUBS 0.008833f
C175 B.n4 VSUBS 0.008833f
C176 B.n5 VSUBS 0.008833f
C177 B.n6 VSUBS 0.008833f
C178 B.n7 VSUBS 0.008833f
C179 B.n8 VSUBS 0.008833f
C180 B.n9 VSUBS 0.008833f
C181 B.n10 VSUBS 0.008833f
C182 B.n11 VSUBS 0.008833f
C183 B.n12 VSUBS 0.008833f
C184 B.n13 VSUBS 0.008833f
C185 B.n14 VSUBS 0.008833f
C186 B.n15 VSUBS 0.008833f
C187 B.n16 VSUBS 0.008833f
C188 B.n17 VSUBS 0.008833f
C189 B.n18 VSUBS 0.008833f
C190 B.n19 VSUBS 0.008833f
C191 B.n20 VSUBS 0.008833f
C192 B.n21 VSUBS 0.008833f
C193 B.n22 VSUBS 0.008833f
C194 B.n23 VSUBS 0.008833f
C195 B.n24 VSUBS 0.008833f
C196 B.n25 VSUBS 0.022476f
C197 B.n26 VSUBS 0.008833f
C198 B.n27 VSUBS 0.008833f
C199 B.n28 VSUBS 0.008833f
C200 B.n29 VSUBS 0.008833f
C201 B.n30 VSUBS 0.008833f
C202 B.n31 VSUBS 0.008833f
C203 B.n32 VSUBS 0.008833f
C204 B.n33 VSUBS 0.008833f
C205 B.n34 VSUBS 0.008833f
C206 B.n35 VSUBS 0.008833f
C207 B.n36 VSUBS 0.008833f
C208 B.n37 VSUBS 0.008833f
C209 B.n38 VSUBS 0.008833f
C210 B.n39 VSUBS 0.008833f
C211 B.n40 VSUBS 0.008833f
C212 B.n41 VSUBS 0.008833f
C213 B.n42 VSUBS 0.008833f
C214 B.n43 VSUBS 0.008833f
C215 B.n44 VSUBS 0.008833f
C216 B.n45 VSUBS 0.008833f
C217 B.t7 VSUBS 0.481183f
C218 B.t8 VSUBS 0.510344f
C219 B.t6 VSUBS 2.00818f
C220 B.n46 VSUBS 0.276299f
C221 B.n47 VSUBS 0.092395f
C222 B.n48 VSUBS 0.008833f
C223 B.n49 VSUBS 0.008833f
C224 B.n50 VSUBS 0.008833f
C225 B.n51 VSUBS 0.008833f
C226 B.t10 VSUBS 0.481174f
C227 B.t11 VSUBS 0.510336f
C228 B.t9 VSUBS 2.00818f
C229 B.n52 VSUBS 0.276307f
C230 B.n53 VSUBS 0.092404f
C231 B.n54 VSUBS 0.020465f
C232 B.n55 VSUBS 0.008833f
C233 B.n56 VSUBS 0.008833f
C234 B.n57 VSUBS 0.008833f
C235 B.n58 VSUBS 0.008833f
C236 B.n59 VSUBS 0.008833f
C237 B.n60 VSUBS 0.008833f
C238 B.n61 VSUBS 0.008833f
C239 B.n62 VSUBS 0.008833f
C240 B.n63 VSUBS 0.008833f
C241 B.n64 VSUBS 0.008833f
C242 B.n65 VSUBS 0.008833f
C243 B.n66 VSUBS 0.008833f
C244 B.n67 VSUBS 0.008833f
C245 B.n68 VSUBS 0.008833f
C246 B.n69 VSUBS 0.008833f
C247 B.n70 VSUBS 0.008833f
C248 B.n71 VSUBS 0.008833f
C249 B.n72 VSUBS 0.008833f
C250 B.n73 VSUBS 0.008833f
C251 B.n74 VSUBS 0.008833f
C252 B.n75 VSUBS 0.021429f
C253 B.n76 VSUBS 0.008833f
C254 B.n77 VSUBS 0.008833f
C255 B.n78 VSUBS 0.008833f
C256 B.n79 VSUBS 0.008833f
C257 B.n80 VSUBS 0.008833f
C258 B.n81 VSUBS 0.008833f
C259 B.n82 VSUBS 0.008833f
C260 B.n83 VSUBS 0.008833f
C261 B.n84 VSUBS 0.008833f
C262 B.n85 VSUBS 0.008833f
C263 B.n86 VSUBS 0.008833f
C264 B.n87 VSUBS 0.008833f
C265 B.n88 VSUBS 0.008833f
C266 B.n89 VSUBS 0.008833f
C267 B.n90 VSUBS 0.008833f
C268 B.n91 VSUBS 0.008833f
C269 B.n92 VSUBS 0.008833f
C270 B.n93 VSUBS 0.008833f
C271 B.n94 VSUBS 0.008833f
C272 B.n95 VSUBS 0.008833f
C273 B.n96 VSUBS 0.008833f
C274 B.n97 VSUBS 0.008833f
C275 B.n98 VSUBS 0.008833f
C276 B.n99 VSUBS 0.008833f
C277 B.n100 VSUBS 0.008833f
C278 B.n101 VSUBS 0.008833f
C279 B.n102 VSUBS 0.008833f
C280 B.n103 VSUBS 0.008833f
C281 B.n104 VSUBS 0.008833f
C282 B.n105 VSUBS 0.008833f
C283 B.n106 VSUBS 0.008833f
C284 B.n107 VSUBS 0.008833f
C285 B.n108 VSUBS 0.008833f
C286 B.n109 VSUBS 0.008833f
C287 B.n110 VSUBS 0.008833f
C288 B.n111 VSUBS 0.008833f
C289 B.n112 VSUBS 0.008833f
C290 B.n113 VSUBS 0.008833f
C291 B.n114 VSUBS 0.008833f
C292 B.n115 VSUBS 0.008833f
C293 B.n116 VSUBS 0.008833f
C294 B.n117 VSUBS 0.008833f
C295 B.n118 VSUBS 0.008833f
C296 B.n119 VSUBS 0.008833f
C297 B.n120 VSUBS 0.008833f
C298 B.n121 VSUBS 0.008833f
C299 B.n122 VSUBS 0.021522f
C300 B.n123 VSUBS 0.008833f
C301 B.n124 VSUBS 0.008833f
C302 B.n125 VSUBS 0.008833f
C303 B.n126 VSUBS 0.008833f
C304 B.n127 VSUBS 0.008833f
C305 B.n128 VSUBS 0.008833f
C306 B.n129 VSUBS 0.008833f
C307 B.n130 VSUBS 0.008833f
C308 B.n131 VSUBS 0.008833f
C309 B.n132 VSUBS 0.008833f
C310 B.n133 VSUBS 0.008833f
C311 B.n134 VSUBS 0.008833f
C312 B.n135 VSUBS 0.008833f
C313 B.n136 VSUBS 0.008833f
C314 B.n137 VSUBS 0.008833f
C315 B.n138 VSUBS 0.008833f
C316 B.n139 VSUBS 0.008833f
C317 B.n140 VSUBS 0.008833f
C318 B.n141 VSUBS 0.008833f
C319 B.n142 VSUBS 0.006105f
C320 B.n143 VSUBS 0.008833f
C321 B.n144 VSUBS 0.008833f
C322 B.n145 VSUBS 0.008833f
C323 B.n146 VSUBS 0.008833f
C324 B.n147 VSUBS 0.008833f
C325 B.t2 VSUBS 0.481183f
C326 B.t1 VSUBS 0.510344f
C327 B.t0 VSUBS 2.00818f
C328 B.n148 VSUBS 0.276299f
C329 B.n149 VSUBS 0.092395f
C330 B.n150 VSUBS 0.008833f
C331 B.n151 VSUBS 0.008833f
C332 B.n152 VSUBS 0.008833f
C333 B.n153 VSUBS 0.008833f
C334 B.n154 VSUBS 0.008833f
C335 B.n155 VSUBS 0.008833f
C336 B.n156 VSUBS 0.008833f
C337 B.n157 VSUBS 0.008833f
C338 B.n158 VSUBS 0.008833f
C339 B.n159 VSUBS 0.008833f
C340 B.n160 VSUBS 0.008833f
C341 B.n161 VSUBS 0.008833f
C342 B.n162 VSUBS 0.008833f
C343 B.n163 VSUBS 0.008833f
C344 B.n164 VSUBS 0.008833f
C345 B.n165 VSUBS 0.008833f
C346 B.n166 VSUBS 0.008833f
C347 B.n167 VSUBS 0.008833f
C348 B.n168 VSUBS 0.008833f
C349 B.n169 VSUBS 0.022476f
C350 B.n170 VSUBS 0.008833f
C351 B.n171 VSUBS 0.008833f
C352 B.n172 VSUBS 0.008833f
C353 B.n173 VSUBS 0.008833f
C354 B.n174 VSUBS 0.008833f
C355 B.n175 VSUBS 0.008833f
C356 B.n176 VSUBS 0.008833f
C357 B.n177 VSUBS 0.008833f
C358 B.n178 VSUBS 0.008833f
C359 B.n179 VSUBS 0.008833f
C360 B.n180 VSUBS 0.008833f
C361 B.n181 VSUBS 0.008833f
C362 B.n182 VSUBS 0.008833f
C363 B.n183 VSUBS 0.008833f
C364 B.n184 VSUBS 0.008833f
C365 B.n185 VSUBS 0.008833f
C366 B.n186 VSUBS 0.008833f
C367 B.n187 VSUBS 0.008833f
C368 B.n188 VSUBS 0.008833f
C369 B.n189 VSUBS 0.008833f
C370 B.n190 VSUBS 0.008833f
C371 B.n191 VSUBS 0.008833f
C372 B.n192 VSUBS 0.008833f
C373 B.n193 VSUBS 0.008833f
C374 B.n194 VSUBS 0.008833f
C375 B.n195 VSUBS 0.008833f
C376 B.n196 VSUBS 0.008833f
C377 B.n197 VSUBS 0.008833f
C378 B.n198 VSUBS 0.008833f
C379 B.n199 VSUBS 0.008833f
C380 B.n200 VSUBS 0.008833f
C381 B.n201 VSUBS 0.008833f
C382 B.n202 VSUBS 0.008833f
C383 B.n203 VSUBS 0.008833f
C384 B.n204 VSUBS 0.008833f
C385 B.n205 VSUBS 0.008833f
C386 B.n206 VSUBS 0.008833f
C387 B.n207 VSUBS 0.008833f
C388 B.n208 VSUBS 0.008833f
C389 B.n209 VSUBS 0.008833f
C390 B.n210 VSUBS 0.008833f
C391 B.n211 VSUBS 0.008833f
C392 B.n212 VSUBS 0.008833f
C393 B.n213 VSUBS 0.008833f
C394 B.n214 VSUBS 0.008833f
C395 B.n215 VSUBS 0.008833f
C396 B.n216 VSUBS 0.008833f
C397 B.n217 VSUBS 0.008833f
C398 B.n218 VSUBS 0.008833f
C399 B.n219 VSUBS 0.008833f
C400 B.n220 VSUBS 0.008833f
C401 B.n221 VSUBS 0.008833f
C402 B.n222 VSUBS 0.008833f
C403 B.n223 VSUBS 0.008833f
C404 B.n224 VSUBS 0.008833f
C405 B.n225 VSUBS 0.008833f
C406 B.n226 VSUBS 0.008833f
C407 B.n227 VSUBS 0.008833f
C408 B.n228 VSUBS 0.008833f
C409 B.n229 VSUBS 0.008833f
C410 B.n230 VSUBS 0.008833f
C411 B.n231 VSUBS 0.008833f
C412 B.n232 VSUBS 0.008833f
C413 B.n233 VSUBS 0.008833f
C414 B.n234 VSUBS 0.008833f
C415 B.n235 VSUBS 0.008833f
C416 B.n236 VSUBS 0.008833f
C417 B.n237 VSUBS 0.008833f
C418 B.n238 VSUBS 0.008833f
C419 B.n239 VSUBS 0.008833f
C420 B.n240 VSUBS 0.008833f
C421 B.n241 VSUBS 0.008833f
C422 B.n242 VSUBS 0.008833f
C423 B.n243 VSUBS 0.008833f
C424 B.n244 VSUBS 0.008833f
C425 B.n245 VSUBS 0.008833f
C426 B.n246 VSUBS 0.008833f
C427 B.n247 VSUBS 0.008833f
C428 B.n248 VSUBS 0.008833f
C429 B.n249 VSUBS 0.008833f
C430 B.n250 VSUBS 0.008833f
C431 B.n251 VSUBS 0.008833f
C432 B.n252 VSUBS 0.008833f
C433 B.n253 VSUBS 0.008833f
C434 B.n254 VSUBS 0.008833f
C435 B.n255 VSUBS 0.008833f
C436 B.n256 VSUBS 0.008833f
C437 B.n257 VSUBS 0.008833f
C438 B.n258 VSUBS 0.021429f
C439 B.n259 VSUBS 0.021429f
C440 B.n260 VSUBS 0.022476f
C441 B.n261 VSUBS 0.008833f
C442 B.n262 VSUBS 0.008833f
C443 B.n263 VSUBS 0.008833f
C444 B.n264 VSUBS 0.008833f
C445 B.n265 VSUBS 0.008833f
C446 B.n266 VSUBS 0.008833f
C447 B.n267 VSUBS 0.008833f
C448 B.n268 VSUBS 0.008833f
C449 B.n269 VSUBS 0.008833f
C450 B.n270 VSUBS 0.008833f
C451 B.n271 VSUBS 0.008833f
C452 B.n272 VSUBS 0.008833f
C453 B.n273 VSUBS 0.008833f
C454 B.n274 VSUBS 0.008833f
C455 B.n275 VSUBS 0.008833f
C456 B.n276 VSUBS 0.008833f
C457 B.n277 VSUBS 0.008833f
C458 B.n278 VSUBS 0.008833f
C459 B.n279 VSUBS 0.008833f
C460 B.n280 VSUBS 0.008833f
C461 B.n281 VSUBS 0.008833f
C462 B.n282 VSUBS 0.008833f
C463 B.n283 VSUBS 0.008833f
C464 B.n284 VSUBS 0.008833f
C465 B.n285 VSUBS 0.008833f
C466 B.n286 VSUBS 0.008833f
C467 B.n287 VSUBS 0.008833f
C468 B.n288 VSUBS 0.008833f
C469 B.n289 VSUBS 0.008833f
C470 B.n290 VSUBS 0.008833f
C471 B.n291 VSUBS 0.008833f
C472 B.n292 VSUBS 0.008833f
C473 B.n293 VSUBS 0.008833f
C474 B.n294 VSUBS 0.008833f
C475 B.n295 VSUBS 0.008833f
C476 B.n296 VSUBS 0.008833f
C477 B.n297 VSUBS 0.008833f
C478 B.n298 VSUBS 0.008833f
C479 B.n299 VSUBS 0.008833f
C480 B.n300 VSUBS 0.008833f
C481 B.n301 VSUBS 0.008833f
C482 B.n302 VSUBS 0.008833f
C483 B.n303 VSUBS 0.008833f
C484 B.n304 VSUBS 0.008833f
C485 B.n305 VSUBS 0.008833f
C486 B.n306 VSUBS 0.008833f
C487 B.n307 VSUBS 0.008833f
C488 B.n308 VSUBS 0.008833f
C489 B.n309 VSUBS 0.008833f
C490 B.n310 VSUBS 0.008833f
C491 B.n311 VSUBS 0.008833f
C492 B.n312 VSUBS 0.008833f
C493 B.n313 VSUBS 0.008833f
C494 B.n314 VSUBS 0.008833f
C495 B.n315 VSUBS 0.008833f
C496 B.n316 VSUBS 0.008833f
C497 B.n317 VSUBS 0.008833f
C498 B.n318 VSUBS 0.008833f
C499 B.n319 VSUBS 0.008833f
C500 B.n320 VSUBS 0.006105f
C501 B.n321 VSUBS 0.020465f
C502 B.n322 VSUBS 0.007144f
C503 B.n323 VSUBS 0.008833f
C504 B.n324 VSUBS 0.008833f
C505 B.n325 VSUBS 0.008833f
C506 B.n326 VSUBS 0.008833f
C507 B.n327 VSUBS 0.008833f
C508 B.n328 VSUBS 0.008833f
C509 B.n329 VSUBS 0.008833f
C510 B.n330 VSUBS 0.008833f
C511 B.n331 VSUBS 0.008833f
C512 B.n332 VSUBS 0.008833f
C513 B.n333 VSUBS 0.008833f
C514 B.t5 VSUBS 0.481174f
C515 B.t4 VSUBS 0.510336f
C516 B.t3 VSUBS 2.00818f
C517 B.n334 VSUBS 0.276307f
C518 B.n335 VSUBS 0.092404f
C519 B.n336 VSUBS 0.020465f
C520 B.n337 VSUBS 0.007144f
C521 B.n338 VSUBS 0.008833f
C522 B.n339 VSUBS 0.008833f
C523 B.n340 VSUBS 0.008833f
C524 B.n341 VSUBS 0.008833f
C525 B.n342 VSUBS 0.008833f
C526 B.n343 VSUBS 0.008833f
C527 B.n344 VSUBS 0.008833f
C528 B.n345 VSUBS 0.008833f
C529 B.n346 VSUBS 0.008833f
C530 B.n347 VSUBS 0.008833f
C531 B.n348 VSUBS 0.008833f
C532 B.n349 VSUBS 0.008833f
C533 B.n350 VSUBS 0.008833f
C534 B.n351 VSUBS 0.008833f
C535 B.n352 VSUBS 0.008833f
C536 B.n353 VSUBS 0.008833f
C537 B.n354 VSUBS 0.008833f
C538 B.n355 VSUBS 0.008833f
C539 B.n356 VSUBS 0.008833f
C540 B.n357 VSUBS 0.008833f
C541 B.n358 VSUBS 0.008833f
C542 B.n359 VSUBS 0.008833f
C543 B.n360 VSUBS 0.008833f
C544 B.n361 VSUBS 0.008833f
C545 B.n362 VSUBS 0.008833f
C546 B.n363 VSUBS 0.008833f
C547 B.n364 VSUBS 0.008833f
C548 B.n365 VSUBS 0.008833f
C549 B.n366 VSUBS 0.008833f
C550 B.n367 VSUBS 0.008833f
C551 B.n368 VSUBS 0.008833f
C552 B.n369 VSUBS 0.008833f
C553 B.n370 VSUBS 0.008833f
C554 B.n371 VSUBS 0.008833f
C555 B.n372 VSUBS 0.008833f
C556 B.n373 VSUBS 0.008833f
C557 B.n374 VSUBS 0.008833f
C558 B.n375 VSUBS 0.008833f
C559 B.n376 VSUBS 0.008833f
C560 B.n377 VSUBS 0.008833f
C561 B.n378 VSUBS 0.008833f
C562 B.n379 VSUBS 0.008833f
C563 B.n380 VSUBS 0.008833f
C564 B.n381 VSUBS 0.008833f
C565 B.n382 VSUBS 0.008833f
C566 B.n383 VSUBS 0.008833f
C567 B.n384 VSUBS 0.008833f
C568 B.n385 VSUBS 0.008833f
C569 B.n386 VSUBS 0.008833f
C570 B.n387 VSUBS 0.008833f
C571 B.n388 VSUBS 0.008833f
C572 B.n389 VSUBS 0.008833f
C573 B.n390 VSUBS 0.008833f
C574 B.n391 VSUBS 0.008833f
C575 B.n392 VSUBS 0.008833f
C576 B.n393 VSUBS 0.008833f
C577 B.n394 VSUBS 0.008833f
C578 B.n395 VSUBS 0.008833f
C579 B.n396 VSUBS 0.008833f
C580 B.n397 VSUBS 0.008833f
C581 B.n398 VSUBS 0.008833f
C582 B.n399 VSUBS 0.022476f
C583 B.n400 VSUBS 0.021429f
C584 B.n401 VSUBS 0.022383f
C585 B.n402 VSUBS 0.008833f
C586 B.n403 VSUBS 0.008833f
C587 B.n404 VSUBS 0.008833f
C588 B.n405 VSUBS 0.008833f
C589 B.n406 VSUBS 0.008833f
C590 B.n407 VSUBS 0.008833f
C591 B.n408 VSUBS 0.008833f
C592 B.n409 VSUBS 0.008833f
C593 B.n410 VSUBS 0.008833f
C594 B.n411 VSUBS 0.008833f
C595 B.n412 VSUBS 0.008833f
C596 B.n413 VSUBS 0.008833f
C597 B.n414 VSUBS 0.008833f
C598 B.n415 VSUBS 0.008833f
C599 B.n416 VSUBS 0.008833f
C600 B.n417 VSUBS 0.008833f
C601 B.n418 VSUBS 0.008833f
C602 B.n419 VSUBS 0.008833f
C603 B.n420 VSUBS 0.008833f
C604 B.n421 VSUBS 0.008833f
C605 B.n422 VSUBS 0.008833f
C606 B.n423 VSUBS 0.008833f
C607 B.n424 VSUBS 0.008833f
C608 B.n425 VSUBS 0.008833f
C609 B.n426 VSUBS 0.008833f
C610 B.n427 VSUBS 0.008833f
C611 B.n428 VSUBS 0.008833f
C612 B.n429 VSUBS 0.008833f
C613 B.n430 VSUBS 0.008833f
C614 B.n431 VSUBS 0.008833f
C615 B.n432 VSUBS 0.008833f
C616 B.n433 VSUBS 0.008833f
C617 B.n434 VSUBS 0.008833f
C618 B.n435 VSUBS 0.008833f
C619 B.n436 VSUBS 0.008833f
C620 B.n437 VSUBS 0.008833f
C621 B.n438 VSUBS 0.008833f
C622 B.n439 VSUBS 0.008833f
C623 B.n440 VSUBS 0.008833f
C624 B.n441 VSUBS 0.008833f
C625 B.n442 VSUBS 0.008833f
C626 B.n443 VSUBS 0.008833f
C627 B.n444 VSUBS 0.008833f
C628 B.n445 VSUBS 0.008833f
C629 B.n446 VSUBS 0.008833f
C630 B.n447 VSUBS 0.008833f
C631 B.n448 VSUBS 0.008833f
C632 B.n449 VSUBS 0.008833f
C633 B.n450 VSUBS 0.008833f
C634 B.n451 VSUBS 0.008833f
C635 B.n452 VSUBS 0.008833f
C636 B.n453 VSUBS 0.008833f
C637 B.n454 VSUBS 0.008833f
C638 B.n455 VSUBS 0.008833f
C639 B.n456 VSUBS 0.008833f
C640 B.n457 VSUBS 0.008833f
C641 B.n458 VSUBS 0.008833f
C642 B.n459 VSUBS 0.008833f
C643 B.n460 VSUBS 0.008833f
C644 B.n461 VSUBS 0.008833f
C645 B.n462 VSUBS 0.008833f
C646 B.n463 VSUBS 0.008833f
C647 B.n464 VSUBS 0.008833f
C648 B.n465 VSUBS 0.008833f
C649 B.n466 VSUBS 0.008833f
C650 B.n467 VSUBS 0.008833f
C651 B.n468 VSUBS 0.008833f
C652 B.n469 VSUBS 0.008833f
C653 B.n470 VSUBS 0.008833f
C654 B.n471 VSUBS 0.008833f
C655 B.n472 VSUBS 0.008833f
C656 B.n473 VSUBS 0.008833f
C657 B.n474 VSUBS 0.008833f
C658 B.n475 VSUBS 0.008833f
C659 B.n476 VSUBS 0.008833f
C660 B.n477 VSUBS 0.008833f
C661 B.n478 VSUBS 0.008833f
C662 B.n479 VSUBS 0.008833f
C663 B.n480 VSUBS 0.008833f
C664 B.n481 VSUBS 0.008833f
C665 B.n482 VSUBS 0.008833f
C666 B.n483 VSUBS 0.008833f
C667 B.n484 VSUBS 0.008833f
C668 B.n485 VSUBS 0.008833f
C669 B.n486 VSUBS 0.008833f
C670 B.n487 VSUBS 0.008833f
C671 B.n488 VSUBS 0.008833f
C672 B.n489 VSUBS 0.008833f
C673 B.n490 VSUBS 0.008833f
C674 B.n491 VSUBS 0.008833f
C675 B.n492 VSUBS 0.008833f
C676 B.n493 VSUBS 0.008833f
C677 B.n494 VSUBS 0.008833f
C678 B.n495 VSUBS 0.008833f
C679 B.n496 VSUBS 0.008833f
C680 B.n497 VSUBS 0.008833f
C681 B.n498 VSUBS 0.008833f
C682 B.n499 VSUBS 0.008833f
C683 B.n500 VSUBS 0.008833f
C684 B.n501 VSUBS 0.008833f
C685 B.n502 VSUBS 0.008833f
C686 B.n503 VSUBS 0.008833f
C687 B.n504 VSUBS 0.008833f
C688 B.n505 VSUBS 0.008833f
C689 B.n506 VSUBS 0.008833f
C690 B.n507 VSUBS 0.008833f
C691 B.n508 VSUBS 0.008833f
C692 B.n509 VSUBS 0.008833f
C693 B.n510 VSUBS 0.008833f
C694 B.n511 VSUBS 0.008833f
C695 B.n512 VSUBS 0.008833f
C696 B.n513 VSUBS 0.008833f
C697 B.n514 VSUBS 0.008833f
C698 B.n515 VSUBS 0.008833f
C699 B.n516 VSUBS 0.008833f
C700 B.n517 VSUBS 0.008833f
C701 B.n518 VSUBS 0.008833f
C702 B.n519 VSUBS 0.008833f
C703 B.n520 VSUBS 0.008833f
C704 B.n521 VSUBS 0.008833f
C705 B.n522 VSUBS 0.008833f
C706 B.n523 VSUBS 0.008833f
C707 B.n524 VSUBS 0.008833f
C708 B.n525 VSUBS 0.008833f
C709 B.n526 VSUBS 0.008833f
C710 B.n527 VSUBS 0.008833f
C711 B.n528 VSUBS 0.008833f
C712 B.n529 VSUBS 0.008833f
C713 B.n530 VSUBS 0.008833f
C714 B.n531 VSUBS 0.008833f
C715 B.n532 VSUBS 0.008833f
C716 B.n533 VSUBS 0.008833f
C717 B.n534 VSUBS 0.008833f
C718 B.n535 VSUBS 0.008833f
C719 B.n536 VSUBS 0.008833f
C720 B.n537 VSUBS 0.008833f
C721 B.n538 VSUBS 0.008833f
C722 B.n539 VSUBS 0.008833f
C723 B.n540 VSUBS 0.021429f
C724 B.n541 VSUBS 0.022476f
C725 B.n542 VSUBS 0.022476f
C726 B.n543 VSUBS 0.008833f
C727 B.n544 VSUBS 0.008833f
C728 B.n545 VSUBS 0.008833f
C729 B.n546 VSUBS 0.008833f
C730 B.n547 VSUBS 0.008833f
C731 B.n548 VSUBS 0.008833f
C732 B.n549 VSUBS 0.008833f
C733 B.n550 VSUBS 0.008833f
C734 B.n551 VSUBS 0.008833f
C735 B.n552 VSUBS 0.008833f
C736 B.n553 VSUBS 0.008833f
C737 B.n554 VSUBS 0.008833f
C738 B.n555 VSUBS 0.008833f
C739 B.n556 VSUBS 0.008833f
C740 B.n557 VSUBS 0.008833f
C741 B.n558 VSUBS 0.008833f
C742 B.n559 VSUBS 0.008833f
C743 B.n560 VSUBS 0.008833f
C744 B.n561 VSUBS 0.008833f
C745 B.n562 VSUBS 0.008833f
C746 B.n563 VSUBS 0.008833f
C747 B.n564 VSUBS 0.008833f
C748 B.n565 VSUBS 0.008833f
C749 B.n566 VSUBS 0.008833f
C750 B.n567 VSUBS 0.008833f
C751 B.n568 VSUBS 0.008833f
C752 B.n569 VSUBS 0.008833f
C753 B.n570 VSUBS 0.008833f
C754 B.n571 VSUBS 0.008833f
C755 B.n572 VSUBS 0.008833f
C756 B.n573 VSUBS 0.008833f
C757 B.n574 VSUBS 0.008833f
C758 B.n575 VSUBS 0.008833f
C759 B.n576 VSUBS 0.008833f
C760 B.n577 VSUBS 0.008833f
C761 B.n578 VSUBS 0.008833f
C762 B.n579 VSUBS 0.008833f
C763 B.n580 VSUBS 0.008833f
C764 B.n581 VSUBS 0.008833f
C765 B.n582 VSUBS 0.008833f
C766 B.n583 VSUBS 0.008833f
C767 B.n584 VSUBS 0.008833f
C768 B.n585 VSUBS 0.008833f
C769 B.n586 VSUBS 0.008833f
C770 B.n587 VSUBS 0.008833f
C771 B.n588 VSUBS 0.008833f
C772 B.n589 VSUBS 0.008833f
C773 B.n590 VSUBS 0.008833f
C774 B.n591 VSUBS 0.008833f
C775 B.n592 VSUBS 0.008833f
C776 B.n593 VSUBS 0.008833f
C777 B.n594 VSUBS 0.008833f
C778 B.n595 VSUBS 0.008833f
C779 B.n596 VSUBS 0.008833f
C780 B.n597 VSUBS 0.008833f
C781 B.n598 VSUBS 0.008833f
C782 B.n599 VSUBS 0.008833f
C783 B.n600 VSUBS 0.008833f
C784 B.n601 VSUBS 0.006105f
C785 B.n602 VSUBS 0.008833f
C786 B.n603 VSUBS 0.008833f
C787 B.n604 VSUBS 0.007144f
C788 B.n605 VSUBS 0.008833f
C789 B.n606 VSUBS 0.008833f
C790 B.n607 VSUBS 0.008833f
C791 B.n608 VSUBS 0.008833f
C792 B.n609 VSUBS 0.008833f
C793 B.n610 VSUBS 0.008833f
C794 B.n611 VSUBS 0.008833f
C795 B.n612 VSUBS 0.008833f
C796 B.n613 VSUBS 0.008833f
C797 B.n614 VSUBS 0.008833f
C798 B.n615 VSUBS 0.008833f
C799 B.n616 VSUBS 0.007144f
C800 B.n617 VSUBS 0.020465f
C801 B.n618 VSUBS 0.006105f
C802 B.n619 VSUBS 0.008833f
C803 B.n620 VSUBS 0.008833f
C804 B.n621 VSUBS 0.008833f
C805 B.n622 VSUBS 0.008833f
C806 B.n623 VSUBS 0.008833f
C807 B.n624 VSUBS 0.008833f
C808 B.n625 VSUBS 0.008833f
C809 B.n626 VSUBS 0.008833f
C810 B.n627 VSUBS 0.008833f
C811 B.n628 VSUBS 0.008833f
C812 B.n629 VSUBS 0.008833f
C813 B.n630 VSUBS 0.008833f
C814 B.n631 VSUBS 0.008833f
C815 B.n632 VSUBS 0.008833f
C816 B.n633 VSUBS 0.008833f
C817 B.n634 VSUBS 0.008833f
C818 B.n635 VSUBS 0.008833f
C819 B.n636 VSUBS 0.008833f
C820 B.n637 VSUBS 0.008833f
C821 B.n638 VSUBS 0.008833f
C822 B.n639 VSUBS 0.008833f
C823 B.n640 VSUBS 0.008833f
C824 B.n641 VSUBS 0.008833f
C825 B.n642 VSUBS 0.008833f
C826 B.n643 VSUBS 0.008833f
C827 B.n644 VSUBS 0.008833f
C828 B.n645 VSUBS 0.008833f
C829 B.n646 VSUBS 0.008833f
C830 B.n647 VSUBS 0.008833f
C831 B.n648 VSUBS 0.008833f
C832 B.n649 VSUBS 0.008833f
C833 B.n650 VSUBS 0.008833f
C834 B.n651 VSUBS 0.008833f
C835 B.n652 VSUBS 0.008833f
C836 B.n653 VSUBS 0.008833f
C837 B.n654 VSUBS 0.008833f
C838 B.n655 VSUBS 0.008833f
C839 B.n656 VSUBS 0.008833f
C840 B.n657 VSUBS 0.008833f
C841 B.n658 VSUBS 0.008833f
C842 B.n659 VSUBS 0.008833f
C843 B.n660 VSUBS 0.008833f
C844 B.n661 VSUBS 0.008833f
C845 B.n662 VSUBS 0.008833f
C846 B.n663 VSUBS 0.008833f
C847 B.n664 VSUBS 0.008833f
C848 B.n665 VSUBS 0.008833f
C849 B.n666 VSUBS 0.008833f
C850 B.n667 VSUBS 0.008833f
C851 B.n668 VSUBS 0.008833f
C852 B.n669 VSUBS 0.008833f
C853 B.n670 VSUBS 0.008833f
C854 B.n671 VSUBS 0.008833f
C855 B.n672 VSUBS 0.008833f
C856 B.n673 VSUBS 0.008833f
C857 B.n674 VSUBS 0.008833f
C858 B.n675 VSUBS 0.008833f
C859 B.n676 VSUBS 0.008833f
C860 B.n677 VSUBS 0.008833f
C861 B.n678 VSUBS 0.022476f
C862 B.n679 VSUBS 0.021429f
C863 B.n680 VSUBS 0.021429f
C864 B.n681 VSUBS 0.008833f
C865 B.n682 VSUBS 0.008833f
C866 B.n683 VSUBS 0.008833f
C867 B.n684 VSUBS 0.008833f
C868 B.n685 VSUBS 0.008833f
C869 B.n686 VSUBS 0.008833f
C870 B.n687 VSUBS 0.008833f
C871 B.n688 VSUBS 0.008833f
C872 B.n689 VSUBS 0.008833f
C873 B.n690 VSUBS 0.008833f
C874 B.n691 VSUBS 0.008833f
C875 B.n692 VSUBS 0.008833f
C876 B.n693 VSUBS 0.008833f
C877 B.n694 VSUBS 0.008833f
C878 B.n695 VSUBS 0.008833f
C879 B.n696 VSUBS 0.008833f
C880 B.n697 VSUBS 0.008833f
C881 B.n698 VSUBS 0.008833f
C882 B.n699 VSUBS 0.008833f
C883 B.n700 VSUBS 0.008833f
C884 B.n701 VSUBS 0.008833f
C885 B.n702 VSUBS 0.008833f
C886 B.n703 VSUBS 0.008833f
C887 B.n704 VSUBS 0.008833f
C888 B.n705 VSUBS 0.008833f
C889 B.n706 VSUBS 0.008833f
C890 B.n707 VSUBS 0.008833f
C891 B.n708 VSUBS 0.008833f
C892 B.n709 VSUBS 0.008833f
C893 B.n710 VSUBS 0.008833f
C894 B.n711 VSUBS 0.008833f
C895 B.n712 VSUBS 0.008833f
C896 B.n713 VSUBS 0.008833f
C897 B.n714 VSUBS 0.008833f
C898 B.n715 VSUBS 0.008833f
C899 B.n716 VSUBS 0.008833f
C900 B.n717 VSUBS 0.008833f
C901 B.n718 VSUBS 0.008833f
C902 B.n719 VSUBS 0.008833f
C903 B.n720 VSUBS 0.008833f
C904 B.n721 VSUBS 0.008833f
C905 B.n722 VSUBS 0.008833f
C906 B.n723 VSUBS 0.008833f
C907 B.n724 VSUBS 0.008833f
C908 B.n725 VSUBS 0.008833f
C909 B.n726 VSUBS 0.008833f
C910 B.n727 VSUBS 0.008833f
C911 B.n728 VSUBS 0.008833f
C912 B.n729 VSUBS 0.008833f
C913 B.n730 VSUBS 0.008833f
C914 B.n731 VSUBS 0.008833f
C915 B.n732 VSUBS 0.008833f
C916 B.n733 VSUBS 0.008833f
C917 B.n734 VSUBS 0.008833f
C918 B.n735 VSUBS 0.008833f
C919 B.n736 VSUBS 0.008833f
C920 B.n737 VSUBS 0.008833f
C921 B.n738 VSUBS 0.008833f
C922 B.n739 VSUBS 0.008833f
C923 B.n740 VSUBS 0.008833f
C924 B.n741 VSUBS 0.008833f
C925 B.n742 VSUBS 0.008833f
C926 B.n743 VSUBS 0.008833f
C927 B.n744 VSUBS 0.008833f
C928 B.n745 VSUBS 0.008833f
C929 B.n746 VSUBS 0.008833f
C930 B.n747 VSUBS 0.011527f
C931 B.n748 VSUBS 0.012279f
C932 B.n749 VSUBS 0.024418f
.ends

