* NGSPICE file created from diff_pair_sample_1601.ext - technology: sky130A

.subckt diff_pair_sample_1601 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VP.t0 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4653 pd=3.15 as=0.4653 ps=3.15 w=2.82 l=3.65
X1 VDD2.t5 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4653 pd=3.15 as=1.0998 ps=6.42 w=2.82 l=3.65
X2 VDD1.t0 VP.t1 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0998 pd=6.42 as=0.4653 ps=3.15 w=2.82 l=3.65
X3 VDD1.t1 VP.t2 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4653 pd=3.15 as=1.0998 ps=6.42 w=2.82 l=3.65
X4 VDD1.t5 VP.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4653 pd=3.15 as=1.0998 ps=6.42 w=2.82 l=3.65
X5 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=1.0998 pd=6.42 as=0 ps=0 w=2.82 l=3.65
X6 VTAIL.t5 VP.t4 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=0.4653 pd=3.15 as=0.4653 ps=3.15 w=2.82 l=3.65
X7 VDD2.t4 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0998 pd=6.42 as=0.4653 ps=3.15 w=2.82 l=3.65
X8 VTAIL.t0 VN.t2 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4653 pd=3.15 as=0.4653 ps=3.15 w=2.82 l=3.65
X9 VDD1.t3 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0998 pd=6.42 as=0.4653 ps=3.15 w=2.82 l=3.65
X10 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4653 pd=3.15 as=1.0998 ps=6.42 w=2.82 l=3.65
X11 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=1.0998 pd=6.42 as=0 ps=0 w=2.82 l=3.65
X12 VTAIL.t11 VN.t4 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=0.4653 pd=3.15 as=0.4653 ps=3.15 w=2.82 l=3.65
X13 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0998 pd=6.42 as=0 ps=0 w=2.82 l=3.65
X14 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0998 pd=6.42 as=0 ps=0 w=2.82 l=3.65
X15 VDD2.t0 VN.t5 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.0998 pd=6.42 as=0.4653 ps=3.15 w=2.82 l=3.65
R0 VP.n16 VP.n13 161.3
R1 VP.n18 VP.n17 161.3
R2 VP.n19 VP.n12 161.3
R3 VP.n21 VP.n20 161.3
R4 VP.n22 VP.n11 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n10 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n55 VP.n54 161.3
R9 VP.n53 VP.n1 161.3
R10 VP.n52 VP.n51 161.3
R11 VP.n50 VP.n2 161.3
R12 VP.n49 VP.n48 161.3
R13 VP.n47 VP.n3 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n44 VP.n4 161.3
R16 VP.n43 VP.n42 161.3
R17 VP.n40 VP.n5 161.3
R18 VP.n39 VP.n38 161.3
R19 VP.n37 VP.n6 161.3
R20 VP.n36 VP.n35 161.3
R21 VP.n34 VP.n7 161.3
R22 VP.n33 VP.n32 161.3
R23 VP.n31 VP.n8 161.3
R24 VP.n30 VP.n29 78.9333
R25 VP.n56 VP.n0 78.9333
R26 VP.n28 VP.n9 78.9333
R27 VP.n15 VP.n14 62.5822
R28 VP.n48 VP.n2 56.5617
R29 VP.n35 VP.n6 56.5617
R30 VP.n20 VP.n11 56.5617
R31 VP.n15 VP.t5 52.2845
R32 VP.n30 VP.n28 45.9844
R33 VP.n33 VP.n8 24.5923
R34 VP.n34 VP.n33 24.5923
R35 VP.n35 VP.n34 24.5923
R36 VP.n39 VP.n6 24.5923
R37 VP.n40 VP.n39 24.5923
R38 VP.n42 VP.n40 24.5923
R39 VP.n46 VP.n4 24.5923
R40 VP.n47 VP.n46 24.5923
R41 VP.n48 VP.n47 24.5923
R42 VP.n52 VP.n2 24.5923
R43 VP.n53 VP.n52 24.5923
R44 VP.n54 VP.n53 24.5923
R45 VP.n24 VP.n11 24.5923
R46 VP.n25 VP.n24 24.5923
R47 VP.n26 VP.n25 24.5923
R48 VP.n18 VP.n13 24.5923
R49 VP.n19 VP.n18 24.5923
R50 VP.n20 VP.n19 24.5923
R51 VP.n29 VP.t1 18.6202
R52 VP.n41 VP.t0 18.6202
R53 VP.n0 VP.t3 18.6202
R54 VP.n9 VP.t2 18.6202
R55 VP.n14 VP.t4 18.6202
R56 VP.n42 VP.n41 12.2964
R57 VP.n41 VP.n4 12.2964
R58 VP.n14 VP.n13 12.2964
R59 VP.n29 VP.n8 11.3127
R60 VP.n54 VP.n0 11.3127
R61 VP.n26 VP.n9 11.3127
R62 VP.n16 VP.n15 3.10329
R63 VP.n28 VP.n27 0.354861
R64 VP.n31 VP.n30 0.354861
R65 VP.n56 VP.n55 0.354861
R66 VP VP.n56 0.267071
R67 VP.n17 VP.n16 0.189894
R68 VP.n17 VP.n12 0.189894
R69 VP.n21 VP.n12 0.189894
R70 VP.n22 VP.n21 0.189894
R71 VP.n23 VP.n22 0.189894
R72 VP.n23 VP.n10 0.189894
R73 VP.n27 VP.n10 0.189894
R74 VP.n32 VP.n31 0.189894
R75 VP.n32 VP.n7 0.189894
R76 VP.n36 VP.n7 0.189894
R77 VP.n37 VP.n36 0.189894
R78 VP.n38 VP.n37 0.189894
R79 VP.n38 VP.n5 0.189894
R80 VP.n43 VP.n5 0.189894
R81 VP.n44 VP.n43 0.189894
R82 VP.n45 VP.n44 0.189894
R83 VP.n45 VP.n3 0.189894
R84 VP.n49 VP.n3 0.189894
R85 VP.n50 VP.n49 0.189894
R86 VP.n51 VP.n50 0.189894
R87 VP.n51 VP.n1 0.189894
R88 VP.n55 VP.n1 0.189894
R89 VDD1 VDD1.t3 91.645
R90 VDD1.n1 VDD1.t0 91.5312
R91 VDD1.n1 VDD1.n0 82.7944
R92 VDD1.n3 VDD1.n2 81.9921
R93 VDD1.n3 VDD1.n1 39.5957
R94 VDD1.n2 VDD1.t4 7.02178
R95 VDD1.n2 VDD1.t1 7.02178
R96 VDD1.n0 VDD1.t2 7.02178
R97 VDD1.n0 VDD1.t5 7.02178
R98 VDD1 VDD1.n3 0.800069
R99 VTAIL.n7 VTAIL.t2 72.3347
R100 VTAIL.n11 VTAIL.t1 72.3345
R101 VTAIL.n2 VTAIL.t6 72.3345
R102 VTAIL.n10 VTAIL.t7 72.3345
R103 VTAIL.n9 VTAIL.n8 65.3134
R104 VTAIL.n6 VTAIL.n5 65.3134
R105 VTAIL.n1 VTAIL.n0 65.3132
R106 VTAIL.n4 VTAIL.n3 65.3132
R107 VTAIL.n6 VTAIL.n4 21.66
R108 VTAIL.n11 VTAIL.n10 18.2289
R109 VTAIL.n0 VTAIL.t10 7.02178
R110 VTAIL.n0 VTAIL.t11 7.02178
R111 VTAIL.n3 VTAIL.t8 7.02178
R112 VTAIL.n3 VTAIL.t9 7.02178
R113 VTAIL.n8 VTAIL.t4 7.02178
R114 VTAIL.n8 VTAIL.t5 7.02178
R115 VTAIL.n5 VTAIL.t3 7.02178
R116 VTAIL.n5 VTAIL.t0 7.02178
R117 VTAIL.n7 VTAIL.n6 3.43153
R118 VTAIL.n10 VTAIL.n9 3.43153
R119 VTAIL.n4 VTAIL.n2 3.43153
R120 VTAIL VTAIL.n11 2.51559
R121 VTAIL.n9 VTAIL.n7 2.18584
R122 VTAIL.n2 VTAIL.n1 2.18584
R123 VTAIL VTAIL.n1 0.916448
R124 B.n646 B.n645 585
R125 B.n647 B.n646 585
R126 B.n199 B.n121 585
R127 B.n198 B.n197 585
R128 B.n196 B.n195 585
R129 B.n194 B.n193 585
R130 B.n192 B.n191 585
R131 B.n190 B.n189 585
R132 B.n188 B.n187 585
R133 B.n186 B.n185 585
R134 B.n184 B.n183 585
R135 B.n182 B.n181 585
R136 B.n180 B.n179 585
R137 B.n178 B.n177 585
R138 B.n176 B.n175 585
R139 B.n174 B.n173 585
R140 B.n172 B.n171 585
R141 B.n170 B.n169 585
R142 B.n168 B.n167 585
R143 B.n166 B.n165 585
R144 B.n164 B.n163 585
R145 B.n162 B.n161 585
R146 B.n160 B.n159 585
R147 B.n158 B.n157 585
R148 B.n156 B.n155 585
R149 B.n153 B.n152 585
R150 B.n151 B.n150 585
R151 B.n149 B.n148 585
R152 B.n147 B.n146 585
R153 B.n145 B.n144 585
R154 B.n143 B.n142 585
R155 B.n141 B.n140 585
R156 B.n139 B.n138 585
R157 B.n137 B.n136 585
R158 B.n135 B.n134 585
R159 B.n133 B.n132 585
R160 B.n131 B.n130 585
R161 B.n129 B.n128 585
R162 B.n102 B.n101 585
R163 B.n650 B.n649 585
R164 B.n644 B.n122 585
R165 B.n122 B.n99 585
R166 B.n643 B.n98 585
R167 B.n654 B.n98 585
R168 B.n642 B.n97 585
R169 B.n655 B.n97 585
R170 B.n641 B.n96 585
R171 B.n656 B.n96 585
R172 B.n640 B.n639 585
R173 B.n639 B.n92 585
R174 B.n638 B.n91 585
R175 B.n662 B.n91 585
R176 B.n637 B.n90 585
R177 B.n663 B.n90 585
R178 B.n636 B.n89 585
R179 B.n664 B.n89 585
R180 B.n635 B.n634 585
R181 B.n634 B.n85 585
R182 B.n633 B.n84 585
R183 B.n670 B.n84 585
R184 B.n632 B.n83 585
R185 B.n671 B.n83 585
R186 B.n631 B.n82 585
R187 B.n672 B.n82 585
R188 B.n630 B.n629 585
R189 B.n629 B.n78 585
R190 B.n628 B.n77 585
R191 B.n678 B.n77 585
R192 B.n627 B.n76 585
R193 B.n679 B.n76 585
R194 B.n626 B.n75 585
R195 B.n680 B.n75 585
R196 B.n625 B.n624 585
R197 B.n624 B.n71 585
R198 B.n623 B.n70 585
R199 B.n686 B.n70 585
R200 B.n622 B.n69 585
R201 B.n687 B.n69 585
R202 B.n621 B.n68 585
R203 B.n688 B.n68 585
R204 B.n620 B.n619 585
R205 B.n619 B.n64 585
R206 B.n618 B.n63 585
R207 B.n694 B.n63 585
R208 B.n617 B.n62 585
R209 B.n695 B.n62 585
R210 B.n616 B.n61 585
R211 B.n696 B.n61 585
R212 B.n615 B.n614 585
R213 B.n614 B.n60 585
R214 B.n613 B.n56 585
R215 B.n702 B.n56 585
R216 B.n612 B.n55 585
R217 B.n703 B.n55 585
R218 B.n611 B.n54 585
R219 B.n704 B.n54 585
R220 B.n610 B.n609 585
R221 B.n609 B.n50 585
R222 B.n608 B.n49 585
R223 B.n710 B.n49 585
R224 B.n607 B.n48 585
R225 B.n711 B.n48 585
R226 B.n606 B.n47 585
R227 B.n712 B.n47 585
R228 B.n605 B.n604 585
R229 B.n604 B.n43 585
R230 B.n603 B.n42 585
R231 B.n718 B.n42 585
R232 B.n602 B.n41 585
R233 B.n719 B.n41 585
R234 B.n601 B.n40 585
R235 B.n720 B.n40 585
R236 B.n600 B.n599 585
R237 B.n599 B.n36 585
R238 B.n598 B.n35 585
R239 B.n726 B.n35 585
R240 B.n597 B.n34 585
R241 B.n727 B.n34 585
R242 B.n596 B.n33 585
R243 B.n728 B.n33 585
R244 B.n595 B.n594 585
R245 B.n594 B.n29 585
R246 B.n593 B.n28 585
R247 B.n734 B.n28 585
R248 B.n592 B.n27 585
R249 B.n735 B.n27 585
R250 B.n591 B.n26 585
R251 B.n736 B.n26 585
R252 B.n590 B.n589 585
R253 B.n589 B.n22 585
R254 B.n588 B.n21 585
R255 B.n742 B.n21 585
R256 B.n587 B.n20 585
R257 B.n743 B.n20 585
R258 B.n586 B.n19 585
R259 B.n744 B.n19 585
R260 B.n585 B.n584 585
R261 B.n584 B.n15 585
R262 B.n583 B.n14 585
R263 B.n750 B.n14 585
R264 B.n582 B.n13 585
R265 B.n751 B.n13 585
R266 B.n581 B.n12 585
R267 B.n752 B.n12 585
R268 B.n580 B.n579 585
R269 B.n579 B.n8 585
R270 B.n578 B.n7 585
R271 B.n758 B.n7 585
R272 B.n577 B.n6 585
R273 B.n759 B.n6 585
R274 B.n576 B.n5 585
R275 B.n760 B.n5 585
R276 B.n575 B.n574 585
R277 B.n574 B.n4 585
R278 B.n573 B.n200 585
R279 B.n573 B.n572 585
R280 B.n563 B.n201 585
R281 B.n202 B.n201 585
R282 B.n565 B.n564 585
R283 B.n566 B.n565 585
R284 B.n562 B.n207 585
R285 B.n207 B.n206 585
R286 B.n561 B.n560 585
R287 B.n560 B.n559 585
R288 B.n209 B.n208 585
R289 B.n210 B.n209 585
R290 B.n552 B.n551 585
R291 B.n553 B.n552 585
R292 B.n550 B.n215 585
R293 B.n215 B.n214 585
R294 B.n549 B.n548 585
R295 B.n548 B.n547 585
R296 B.n217 B.n216 585
R297 B.n218 B.n217 585
R298 B.n540 B.n539 585
R299 B.n541 B.n540 585
R300 B.n538 B.n223 585
R301 B.n223 B.n222 585
R302 B.n537 B.n536 585
R303 B.n536 B.n535 585
R304 B.n225 B.n224 585
R305 B.n226 B.n225 585
R306 B.n528 B.n527 585
R307 B.n529 B.n528 585
R308 B.n526 B.n231 585
R309 B.n231 B.n230 585
R310 B.n525 B.n524 585
R311 B.n524 B.n523 585
R312 B.n233 B.n232 585
R313 B.n234 B.n233 585
R314 B.n516 B.n515 585
R315 B.n517 B.n516 585
R316 B.n514 B.n239 585
R317 B.n239 B.n238 585
R318 B.n513 B.n512 585
R319 B.n512 B.n511 585
R320 B.n241 B.n240 585
R321 B.n242 B.n241 585
R322 B.n504 B.n503 585
R323 B.n505 B.n504 585
R324 B.n502 B.n247 585
R325 B.n247 B.n246 585
R326 B.n501 B.n500 585
R327 B.n500 B.n499 585
R328 B.n249 B.n248 585
R329 B.n250 B.n249 585
R330 B.n492 B.n491 585
R331 B.n493 B.n492 585
R332 B.n490 B.n255 585
R333 B.n255 B.n254 585
R334 B.n489 B.n488 585
R335 B.n488 B.n487 585
R336 B.n257 B.n256 585
R337 B.n480 B.n257 585
R338 B.n479 B.n478 585
R339 B.n481 B.n479 585
R340 B.n477 B.n262 585
R341 B.n262 B.n261 585
R342 B.n476 B.n475 585
R343 B.n475 B.n474 585
R344 B.n264 B.n263 585
R345 B.n265 B.n264 585
R346 B.n467 B.n466 585
R347 B.n468 B.n467 585
R348 B.n465 B.n270 585
R349 B.n270 B.n269 585
R350 B.n464 B.n463 585
R351 B.n463 B.n462 585
R352 B.n272 B.n271 585
R353 B.n273 B.n272 585
R354 B.n455 B.n454 585
R355 B.n456 B.n455 585
R356 B.n453 B.n278 585
R357 B.n278 B.n277 585
R358 B.n452 B.n451 585
R359 B.n451 B.n450 585
R360 B.n280 B.n279 585
R361 B.n281 B.n280 585
R362 B.n443 B.n442 585
R363 B.n444 B.n443 585
R364 B.n441 B.n286 585
R365 B.n286 B.n285 585
R366 B.n440 B.n439 585
R367 B.n439 B.n438 585
R368 B.n288 B.n287 585
R369 B.n289 B.n288 585
R370 B.n431 B.n430 585
R371 B.n432 B.n431 585
R372 B.n429 B.n294 585
R373 B.n294 B.n293 585
R374 B.n428 B.n427 585
R375 B.n427 B.n426 585
R376 B.n296 B.n295 585
R377 B.n297 B.n296 585
R378 B.n419 B.n418 585
R379 B.n420 B.n419 585
R380 B.n417 B.n302 585
R381 B.n302 B.n301 585
R382 B.n416 B.n415 585
R383 B.n415 B.n414 585
R384 B.n304 B.n303 585
R385 B.n305 B.n304 585
R386 B.n410 B.n409 585
R387 B.n308 B.n307 585
R388 B.n406 B.n405 585
R389 B.n407 B.n406 585
R390 B.n404 B.n327 585
R391 B.n403 B.n402 585
R392 B.n401 B.n400 585
R393 B.n399 B.n398 585
R394 B.n397 B.n396 585
R395 B.n395 B.n394 585
R396 B.n393 B.n392 585
R397 B.n391 B.n390 585
R398 B.n389 B.n388 585
R399 B.n387 B.n386 585
R400 B.n385 B.n384 585
R401 B.n383 B.n382 585
R402 B.n381 B.n380 585
R403 B.n379 B.n378 585
R404 B.n377 B.n376 585
R405 B.n375 B.n374 585
R406 B.n373 B.n372 585
R407 B.n371 B.n370 585
R408 B.n369 B.n368 585
R409 B.n367 B.n366 585
R410 B.n365 B.n364 585
R411 B.n362 B.n361 585
R412 B.n360 B.n359 585
R413 B.n358 B.n357 585
R414 B.n356 B.n355 585
R415 B.n354 B.n353 585
R416 B.n352 B.n351 585
R417 B.n350 B.n349 585
R418 B.n348 B.n347 585
R419 B.n346 B.n345 585
R420 B.n344 B.n343 585
R421 B.n342 B.n341 585
R422 B.n340 B.n339 585
R423 B.n338 B.n337 585
R424 B.n336 B.n335 585
R425 B.n334 B.n333 585
R426 B.n411 B.n306 585
R427 B.n306 B.n305 585
R428 B.n413 B.n412 585
R429 B.n414 B.n413 585
R430 B.n300 B.n299 585
R431 B.n301 B.n300 585
R432 B.n422 B.n421 585
R433 B.n421 B.n420 585
R434 B.n423 B.n298 585
R435 B.n298 B.n297 585
R436 B.n425 B.n424 585
R437 B.n426 B.n425 585
R438 B.n292 B.n291 585
R439 B.n293 B.n292 585
R440 B.n434 B.n433 585
R441 B.n433 B.n432 585
R442 B.n435 B.n290 585
R443 B.n290 B.n289 585
R444 B.n437 B.n436 585
R445 B.n438 B.n437 585
R446 B.n284 B.n283 585
R447 B.n285 B.n284 585
R448 B.n446 B.n445 585
R449 B.n445 B.n444 585
R450 B.n447 B.n282 585
R451 B.n282 B.n281 585
R452 B.n449 B.n448 585
R453 B.n450 B.n449 585
R454 B.n276 B.n275 585
R455 B.n277 B.n276 585
R456 B.n458 B.n457 585
R457 B.n457 B.n456 585
R458 B.n459 B.n274 585
R459 B.n274 B.n273 585
R460 B.n461 B.n460 585
R461 B.n462 B.n461 585
R462 B.n268 B.n267 585
R463 B.n269 B.n268 585
R464 B.n470 B.n469 585
R465 B.n469 B.n468 585
R466 B.n471 B.n266 585
R467 B.n266 B.n265 585
R468 B.n473 B.n472 585
R469 B.n474 B.n473 585
R470 B.n260 B.n259 585
R471 B.n261 B.n260 585
R472 B.n483 B.n482 585
R473 B.n482 B.n481 585
R474 B.n484 B.n258 585
R475 B.n480 B.n258 585
R476 B.n486 B.n485 585
R477 B.n487 B.n486 585
R478 B.n253 B.n252 585
R479 B.n254 B.n253 585
R480 B.n495 B.n494 585
R481 B.n494 B.n493 585
R482 B.n496 B.n251 585
R483 B.n251 B.n250 585
R484 B.n498 B.n497 585
R485 B.n499 B.n498 585
R486 B.n245 B.n244 585
R487 B.n246 B.n245 585
R488 B.n507 B.n506 585
R489 B.n506 B.n505 585
R490 B.n508 B.n243 585
R491 B.n243 B.n242 585
R492 B.n510 B.n509 585
R493 B.n511 B.n510 585
R494 B.n237 B.n236 585
R495 B.n238 B.n237 585
R496 B.n519 B.n518 585
R497 B.n518 B.n517 585
R498 B.n520 B.n235 585
R499 B.n235 B.n234 585
R500 B.n522 B.n521 585
R501 B.n523 B.n522 585
R502 B.n229 B.n228 585
R503 B.n230 B.n229 585
R504 B.n531 B.n530 585
R505 B.n530 B.n529 585
R506 B.n532 B.n227 585
R507 B.n227 B.n226 585
R508 B.n534 B.n533 585
R509 B.n535 B.n534 585
R510 B.n221 B.n220 585
R511 B.n222 B.n221 585
R512 B.n543 B.n542 585
R513 B.n542 B.n541 585
R514 B.n544 B.n219 585
R515 B.n219 B.n218 585
R516 B.n546 B.n545 585
R517 B.n547 B.n546 585
R518 B.n213 B.n212 585
R519 B.n214 B.n213 585
R520 B.n555 B.n554 585
R521 B.n554 B.n553 585
R522 B.n556 B.n211 585
R523 B.n211 B.n210 585
R524 B.n558 B.n557 585
R525 B.n559 B.n558 585
R526 B.n205 B.n204 585
R527 B.n206 B.n205 585
R528 B.n568 B.n567 585
R529 B.n567 B.n566 585
R530 B.n569 B.n203 585
R531 B.n203 B.n202 585
R532 B.n571 B.n570 585
R533 B.n572 B.n571 585
R534 B.n2 B.n0 585
R535 B.n4 B.n2 585
R536 B.n3 B.n1 585
R537 B.n759 B.n3 585
R538 B.n757 B.n756 585
R539 B.n758 B.n757 585
R540 B.n755 B.n9 585
R541 B.n9 B.n8 585
R542 B.n754 B.n753 585
R543 B.n753 B.n752 585
R544 B.n11 B.n10 585
R545 B.n751 B.n11 585
R546 B.n749 B.n748 585
R547 B.n750 B.n749 585
R548 B.n747 B.n16 585
R549 B.n16 B.n15 585
R550 B.n746 B.n745 585
R551 B.n745 B.n744 585
R552 B.n18 B.n17 585
R553 B.n743 B.n18 585
R554 B.n741 B.n740 585
R555 B.n742 B.n741 585
R556 B.n739 B.n23 585
R557 B.n23 B.n22 585
R558 B.n738 B.n737 585
R559 B.n737 B.n736 585
R560 B.n25 B.n24 585
R561 B.n735 B.n25 585
R562 B.n733 B.n732 585
R563 B.n734 B.n733 585
R564 B.n731 B.n30 585
R565 B.n30 B.n29 585
R566 B.n730 B.n729 585
R567 B.n729 B.n728 585
R568 B.n32 B.n31 585
R569 B.n727 B.n32 585
R570 B.n725 B.n724 585
R571 B.n726 B.n725 585
R572 B.n723 B.n37 585
R573 B.n37 B.n36 585
R574 B.n722 B.n721 585
R575 B.n721 B.n720 585
R576 B.n39 B.n38 585
R577 B.n719 B.n39 585
R578 B.n717 B.n716 585
R579 B.n718 B.n717 585
R580 B.n715 B.n44 585
R581 B.n44 B.n43 585
R582 B.n714 B.n713 585
R583 B.n713 B.n712 585
R584 B.n46 B.n45 585
R585 B.n711 B.n46 585
R586 B.n709 B.n708 585
R587 B.n710 B.n709 585
R588 B.n707 B.n51 585
R589 B.n51 B.n50 585
R590 B.n706 B.n705 585
R591 B.n705 B.n704 585
R592 B.n53 B.n52 585
R593 B.n703 B.n53 585
R594 B.n701 B.n700 585
R595 B.n702 B.n701 585
R596 B.n699 B.n57 585
R597 B.n60 B.n57 585
R598 B.n698 B.n697 585
R599 B.n697 B.n696 585
R600 B.n59 B.n58 585
R601 B.n695 B.n59 585
R602 B.n693 B.n692 585
R603 B.n694 B.n693 585
R604 B.n691 B.n65 585
R605 B.n65 B.n64 585
R606 B.n690 B.n689 585
R607 B.n689 B.n688 585
R608 B.n67 B.n66 585
R609 B.n687 B.n67 585
R610 B.n685 B.n684 585
R611 B.n686 B.n685 585
R612 B.n683 B.n72 585
R613 B.n72 B.n71 585
R614 B.n682 B.n681 585
R615 B.n681 B.n680 585
R616 B.n74 B.n73 585
R617 B.n679 B.n74 585
R618 B.n677 B.n676 585
R619 B.n678 B.n677 585
R620 B.n675 B.n79 585
R621 B.n79 B.n78 585
R622 B.n674 B.n673 585
R623 B.n673 B.n672 585
R624 B.n81 B.n80 585
R625 B.n671 B.n81 585
R626 B.n669 B.n668 585
R627 B.n670 B.n669 585
R628 B.n667 B.n86 585
R629 B.n86 B.n85 585
R630 B.n666 B.n665 585
R631 B.n665 B.n664 585
R632 B.n88 B.n87 585
R633 B.n663 B.n88 585
R634 B.n661 B.n660 585
R635 B.n662 B.n661 585
R636 B.n659 B.n93 585
R637 B.n93 B.n92 585
R638 B.n658 B.n657 585
R639 B.n657 B.n656 585
R640 B.n95 B.n94 585
R641 B.n655 B.n95 585
R642 B.n653 B.n652 585
R643 B.n654 B.n653 585
R644 B.n651 B.n100 585
R645 B.n100 B.n99 585
R646 B.n762 B.n761 585
R647 B.n761 B.n760 585
R648 B.n409 B.n306 473.281
R649 B.n649 B.n100 473.281
R650 B.n333 B.n304 473.281
R651 B.n646 B.n122 473.281
R652 B.n647 B.n120 256.663
R653 B.n647 B.n119 256.663
R654 B.n647 B.n118 256.663
R655 B.n647 B.n117 256.663
R656 B.n647 B.n116 256.663
R657 B.n647 B.n115 256.663
R658 B.n647 B.n114 256.663
R659 B.n647 B.n113 256.663
R660 B.n647 B.n112 256.663
R661 B.n647 B.n111 256.663
R662 B.n647 B.n110 256.663
R663 B.n647 B.n109 256.663
R664 B.n647 B.n108 256.663
R665 B.n647 B.n107 256.663
R666 B.n647 B.n106 256.663
R667 B.n647 B.n105 256.663
R668 B.n647 B.n104 256.663
R669 B.n647 B.n103 256.663
R670 B.n648 B.n647 256.663
R671 B.n408 B.n407 256.663
R672 B.n407 B.n309 256.663
R673 B.n407 B.n310 256.663
R674 B.n407 B.n311 256.663
R675 B.n407 B.n312 256.663
R676 B.n407 B.n313 256.663
R677 B.n407 B.n314 256.663
R678 B.n407 B.n315 256.663
R679 B.n407 B.n316 256.663
R680 B.n407 B.n317 256.663
R681 B.n407 B.n318 256.663
R682 B.n407 B.n319 256.663
R683 B.n407 B.n320 256.663
R684 B.n407 B.n321 256.663
R685 B.n407 B.n322 256.663
R686 B.n407 B.n323 256.663
R687 B.n407 B.n324 256.663
R688 B.n407 B.n325 256.663
R689 B.n407 B.n326 256.663
R690 B.n331 B.t10 227.844
R691 B.n328 B.t6 227.844
R692 B.n126 B.t17 227.844
R693 B.n123 B.t13 227.844
R694 B.n413 B.n306 163.367
R695 B.n413 B.n300 163.367
R696 B.n421 B.n300 163.367
R697 B.n421 B.n298 163.367
R698 B.n425 B.n298 163.367
R699 B.n425 B.n292 163.367
R700 B.n433 B.n292 163.367
R701 B.n433 B.n290 163.367
R702 B.n437 B.n290 163.367
R703 B.n437 B.n284 163.367
R704 B.n445 B.n284 163.367
R705 B.n445 B.n282 163.367
R706 B.n449 B.n282 163.367
R707 B.n449 B.n276 163.367
R708 B.n457 B.n276 163.367
R709 B.n457 B.n274 163.367
R710 B.n461 B.n274 163.367
R711 B.n461 B.n268 163.367
R712 B.n469 B.n268 163.367
R713 B.n469 B.n266 163.367
R714 B.n473 B.n266 163.367
R715 B.n473 B.n260 163.367
R716 B.n482 B.n260 163.367
R717 B.n482 B.n258 163.367
R718 B.n486 B.n258 163.367
R719 B.n486 B.n253 163.367
R720 B.n494 B.n253 163.367
R721 B.n494 B.n251 163.367
R722 B.n498 B.n251 163.367
R723 B.n498 B.n245 163.367
R724 B.n506 B.n245 163.367
R725 B.n506 B.n243 163.367
R726 B.n510 B.n243 163.367
R727 B.n510 B.n237 163.367
R728 B.n518 B.n237 163.367
R729 B.n518 B.n235 163.367
R730 B.n522 B.n235 163.367
R731 B.n522 B.n229 163.367
R732 B.n530 B.n229 163.367
R733 B.n530 B.n227 163.367
R734 B.n534 B.n227 163.367
R735 B.n534 B.n221 163.367
R736 B.n542 B.n221 163.367
R737 B.n542 B.n219 163.367
R738 B.n546 B.n219 163.367
R739 B.n546 B.n213 163.367
R740 B.n554 B.n213 163.367
R741 B.n554 B.n211 163.367
R742 B.n558 B.n211 163.367
R743 B.n558 B.n205 163.367
R744 B.n567 B.n205 163.367
R745 B.n567 B.n203 163.367
R746 B.n571 B.n203 163.367
R747 B.n571 B.n2 163.367
R748 B.n761 B.n2 163.367
R749 B.n761 B.n3 163.367
R750 B.n757 B.n3 163.367
R751 B.n757 B.n9 163.367
R752 B.n753 B.n9 163.367
R753 B.n753 B.n11 163.367
R754 B.n749 B.n11 163.367
R755 B.n749 B.n16 163.367
R756 B.n745 B.n16 163.367
R757 B.n745 B.n18 163.367
R758 B.n741 B.n18 163.367
R759 B.n741 B.n23 163.367
R760 B.n737 B.n23 163.367
R761 B.n737 B.n25 163.367
R762 B.n733 B.n25 163.367
R763 B.n733 B.n30 163.367
R764 B.n729 B.n30 163.367
R765 B.n729 B.n32 163.367
R766 B.n725 B.n32 163.367
R767 B.n725 B.n37 163.367
R768 B.n721 B.n37 163.367
R769 B.n721 B.n39 163.367
R770 B.n717 B.n39 163.367
R771 B.n717 B.n44 163.367
R772 B.n713 B.n44 163.367
R773 B.n713 B.n46 163.367
R774 B.n709 B.n46 163.367
R775 B.n709 B.n51 163.367
R776 B.n705 B.n51 163.367
R777 B.n705 B.n53 163.367
R778 B.n701 B.n53 163.367
R779 B.n701 B.n57 163.367
R780 B.n697 B.n57 163.367
R781 B.n697 B.n59 163.367
R782 B.n693 B.n59 163.367
R783 B.n693 B.n65 163.367
R784 B.n689 B.n65 163.367
R785 B.n689 B.n67 163.367
R786 B.n685 B.n67 163.367
R787 B.n685 B.n72 163.367
R788 B.n681 B.n72 163.367
R789 B.n681 B.n74 163.367
R790 B.n677 B.n74 163.367
R791 B.n677 B.n79 163.367
R792 B.n673 B.n79 163.367
R793 B.n673 B.n81 163.367
R794 B.n669 B.n81 163.367
R795 B.n669 B.n86 163.367
R796 B.n665 B.n86 163.367
R797 B.n665 B.n88 163.367
R798 B.n661 B.n88 163.367
R799 B.n661 B.n93 163.367
R800 B.n657 B.n93 163.367
R801 B.n657 B.n95 163.367
R802 B.n653 B.n95 163.367
R803 B.n653 B.n100 163.367
R804 B.n406 B.n308 163.367
R805 B.n406 B.n327 163.367
R806 B.n402 B.n401 163.367
R807 B.n398 B.n397 163.367
R808 B.n394 B.n393 163.367
R809 B.n390 B.n389 163.367
R810 B.n386 B.n385 163.367
R811 B.n382 B.n381 163.367
R812 B.n378 B.n377 163.367
R813 B.n374 B.n373 163.367
R814 B.n370 B.n369 163.367
R815 B.n366 B.n365 163.367
R816 B.n361 B.n360 163.367
R817 B.n357 B.n356 163.367
R818 B.n353 B.n352 163.367
R819 B.n349 B.n348 163.367
R820 B.n345 B.n344 163.367
R821 B.n341 B.n340 163.367
R822 B.n337 B.n336 163.367
R823 B.n415 B.n304 163.367
R824 B.n415 B.n302 163.367
R825 B.n419 B.n302 163.367
R826 B.n419 B.n296 163.367
R827 B.n427 B.n296 163.367
R828 B.n427 B.n294 163.367
R829 B.n431 B.n294 163.367
R830 B.n431 B.n288 163.367
R831 B.n439 B.n288 163.367
R832 B.n439 B.n286 163.367
R833 B.n443 B.n286 163.367
R834 B.n443 B.n280 163.367
R835 B.n451 B.n280 163.367
R836 B.n451 B.n278 163.367
R837 B.n455 B.n278 163.367
R838 B.n455 B.n272 163.367
R839 B.n463 B.n272 163.367
R840 B.n463 B.n270 163.367
R841 B.n467 B.n270 163.367
R842 B.n467 B.n264 163.367
R843 B.n475 B.n264 163.367
R844 B.n475 B.n262 163.367
R845 B.n479 B.n262 163.367
R846 B.n479 B.n257 163.367
R847 B.n488 B.n257 163.367
R848 B.n488 B.n255 163.367
R849 B.n492 B.n255 163.367
R850 B.n492 B.n249 163.367
R851 B.n500 B.n249 163.367
R852 B.n500 B.n247 163.367
R853 B.n504 B.n247 163.367
R854 B.n504 B.n241 163.367
R855 B.n512 B.n241 163.367
R856 B.n512 B.n239 163.367
R857 B.n516 B.n239 163.367
R858 B.n516 B.n233 163.367
R859 B.n524 B.n233 163.367
R860 B.n524 B.n231 163.367
R861 B.n528 B.n231 163.367
R862 B.n528 B.n225 163.367
R863 B.n536 B.n225 163.367
R864 B.n536 B.n223 163.367
R865 B.n540 B.n223 163.367
R866 B.n540 B.n217 163.367
R867 B.n548 B.n217 163.367
R868 B.n548 B.n215 163.367
R869 B.n552 B.n215 163.367
R870 B.n552 B.n209 163.367
R871 B.n560 B.n209 163.367
R872 B.n560 B.n207 163.367
R873 B.n565 B.n207 163.367
R874 B.n565 B.n201 163.367
R875 B.n573 B.n201 163.367
R876 B.n574 B.n573 163.367
R877 B.n574 B.n5 163.367
R878 B.n6 B.n5 163.367
R879 B.n7 B.n6 163.367
R880 B.n579 B.n7 163.367
R881 B.n579 B.n12 163.367
R882 B.n13 B.n12 163.367
R883 B.n14 B.n13 163.367
R884 B.n584 B.n14 163.367
R885 B.n584 B.n19 163.367
R886 B.n20 B.n19 163.367
R887 B.n21 B.n20 163.367
R888 B.n589 B.n21 163.367
R889 B.n589 B.n26 163.367
R890 B.n27 B.n26 163.367
R891 B.n28 B.n27 163.367
R892 B.n594 B.n28 163.367
R893 B.n594 B.n33 163.367
R894 B.n34 B.n33 163.367
R895 B.n35 B.n34 163.367
R896 B.n599 B.n35 163.367
R897 B.n599 B.n40 163.367
R898 B.n41 B.n40 163.367
R899 B.n42 B.n41 163.367
R900 B.n604 B.n42 163.367
R901 B.n604 B.n47 163.367
R902 B.n48 B.n47 163.367
R903 B.n49 B.n48 163.367
R904 B.n609 B.n49 163.367
R905 B.n609 B.n54 163.367
R906 B.n55 B.n54 163.367
R907 B.n56 B.n55 163.367
R908 B.n614 B.n56 163.367
R909 B.n614 B.n61 163.367
R910 B.n62 B.n61 163.367
R911 B.n63 B.n62 163.367
R912 B.n619 B.n63 163.367
R913 B.n619 B.n68 163.367
R914 B.n69 B.n68 163.367
R915 B.n70 B.n69 163.367
R916 B.n624 B.n70 163.367
R917 B.n624 B.n75 163.367
R918 B.n76 B.n75 163.367
R919 B.n77 B.n76 163.367
R920 B.n629 B.n77 163.367
R921 B.n629 B.n82 163.367
R922 B.n83 B.n82 163.367
R923 B.n84 B.n83 163.367
R924 B.n634 B.n84 163.367
R925 B.n634 B.n89 163.367
R926 B.n90 B.n89 163.367
R927 B.n91 B.n90 163.367
R928 B.n639 B.n91 163.367
R929 B.n639 B.n96 163.367
R930 B.n97 B.n96 163.367
R931 B.n98 B.n97 163.367
R932 B.n122 B.n98 163.367
R933 B.n128 B.n102 163.367
R934 B.n132 B.n131 163.367
R935 B.n136 B.n135 163.367
R936 B.n140 B.n139 163.367
R937 B.n144 B.n143 163.367
R938 B.n148 B.n147 163.367
R939 B.n152 B.n151 163.367
R940 B.n157 B.n156 163.367
R941 B.n161 B.n160 163.367
R942 B.n165 B.n164 163.367
R943 B.n169 B.n168 163.367
R944 B.n173 B.n172 163.367
R945 B.n177 B.n176 163.367
R946 B.n181 B.n180 163.367
R947 B.n185 B.n184 163.367
R948 B.n189 B.n188 163.367
R949 B.n193 B.n192 163.367
R950 B.n197 B.n196 163.367
R951 B.n646 B.n121 163.367
R952 B.n407 B.n305 161.706
R953 B.n647 B.n99 161.706
R954 B.n331 B.t12 154.733
R955 B.n123 B.t15 154.733
R956 B.n328 B.t9 154.732
R957 B.n126 B.t18 154.732
R958 B.n414 B.n305 92.4032
R959 B.n414 B.n301 92.4032
R960 B.n420 B.n301 92.4032
R961 B.n420 B.n297 92.4032
R962 B.n426 B.n297 92.4032
R963 B.n426 B.n293 92.4032
R964 B.n432 B.n293 92.4032
R965 B.n432 B.n289 92.4032
R966 B.n438 B.n289 92.4032
R967 B.n444 B.n285 92.4032
R968 B.n444 B.n281 92.4032
R969 B.n450 B.n281 92.4032
R970 B.n450 B.n277 92.4032
R971 B.n456 B.n277 92.4032
R972 B.n456 B.n273 92.4032
R973 B.n462 B.n273 92.4032
R974 B.n462 B.n269 92.4032
R975 B.n468 B.n269 92.4032
R976 B.n468 B.n265 92.4032
R977 B.n474 B.n265 92.4032
R978 B.n474 B.n261 92.4032
R979 B.n481 B.n261 92.4032
R980 B.n481 B.n480 92.4032
R981 B.n487 B.n254 92.4032
R982 B.n493 B.n254 92.4032
R983 B.n493 B.n250 92.4032
R984 B.n499 B.n250 92.4032
R985 B.n499 B.n246 92.4032
R986 B.n505 B.n246 92.4032
R987 B.n505 B.n242 92.4032
R988 B.n511 B.n242 92.4032
R989 B.n511 B.n238 92.4032
R990 B.n517 B.n238 92.4032
R991 B.n523 B.n234 92.4032
R992 B.n523 B.n230 92.4032
R993 B.n529 B.n230 92.4032
R994 B.n529 B.n226 92.4032
R995 B.n535 B.n226 92.4032
R996 B.n535 B.n222 92.4032
R997 B.n541 B.n222 92.4032
R998 B.n541 B.n218 92.4032
R999 B.n547 B.n218 92.4032
R1000 B.n547 B.n214 92.4032
R1001 B.n553 B.n214 92.4032
R1002 B.n559 B.n210 92.4032
R1003 B.n559 B.n206 92.4032
R1004 B.n566 B.n206 92.4032
R1005 B.n566 B.n202 92.4032
R1006 B.n572 B.n202 92.4032
R1007 B.n572 B.n4 92.4032
R1008 B.n760 B.n4 92.4032
R1009 B.n760 B.n759 92.4032
R1010 B.n759 B.n758 92.4032
R1011 B.n758 B.n8 92.4032
R1012 B.n752 B.n8 92.4032
R1013 B.n752 B.n751 92.4032
R1014 B.n751 B.n750 92.4032
R1015 B.n750 B.n15 92.4032
R1016 B.n744 B.n743 92.4032
R1017 B.n743 B.n742 92.4032
R1018 B.n742 B.n22 92.4032
R1019 B.n736 B.n22 92.4032
R1020 B.n736 B.n735 92.4032
R1021 B.n735 B.n734 92.4032
R1022 B.n734 B.n29 92.4032
R1023 B.n728 B.n29 92.4032
R1024 B.n728 B.n727 92.4032
R1025 B.n727 B.n726 92.4032
R1026 B.n726 B.n36 92.4032
R1027 B.n720 B.n719 92.4032
R1028 B.n719 B.n718 92.4032
R1029 B.n718 B.n43 92.4032
R1030 B.n712 B.n43 92.4032
R1031 B.n712 B.n711 92.4032
R1032 B.n711 B.n710 92.4032
R1033 B.n710 B.n50 92.4032
R1034 B.n704 B.n50 92.4032
R1035 B.n704 B.n703 92.4032
R1036 B.n703 B.n702 92.4032
R1037 B.n696 B.n60 92.4032
R1038 B.n696 B.n695 92.4032
R1039 B.n695 B.n694 92.4032
R1040 B.n694 B.n64 92.4032
R1041 B.n688 B.n64 92.4032
R1042 B.n688 B.n687 92.4032
R1043 B.n687 B.n686 92.4032
R1044 B.n686 B.n71 92.4032
R1045 B.n680 B.n71 92.4032
R1046 B.n680 B.n679 92.4032
R1047 B.n679 B.n678 92.4032
R1048 B.n678 B.n78 92.4032
R1049 B.n672 B.n78 92.4032
R1050 B.n672 B.n671 92.4032
R1051 B.n670 B.n85 92.4032
R1052 B.n664 B.n85 92.4032
R1053 B.n664 B.n663 92.4032
R1054 B.n663 B.n662 92.4032
R1055 B.n662 B.n92 92.4032
R1056 B.n656 B.n92 92.4032
R1057 B.n656 B.n655 92.4032
R1058 B.n655 B.n654 92.4032
R1059 B.n654 B.n99 92.4032
R1060 B.n487 B.t3 80.1734
R1061 B.n702 B.t1 80.1734
R1062 B.n332 B.t11 77.5452
R1063 B.n124 B.t16 77.5452
R1064 B.n329 B.t8 77.5434
R1065 B.n127 B.t19 77.5434
R1066 B.n517 B.t0 77.4557
R1067 B.n720 B.t5 77.4557
R1068 B.n332 B.n331 77.1884
R1069 B.n329 B.n328 77.1884
R1070 B.n127 B.n126 77.1884
R1071 B.n124 B.n123 77.1884
R1072 B.t7 B.n285 72.0203
R1073 B.n671 B.t14 72.0203
R1074 B.n409 B.n408 71.676
R1075 B.n327 B.n309 71.676
R1076 B.n401 B.n310 71.676
R1077 B.n397 B.n311 71.676
R1078 B.n393 B.n312 71.676
R1079 B.n389 B.n313 71.676
R1080 B.n385 B.n314 71.676
R1081 B.n381 B.n315 71.676
R1082 B.n377 B.n316 71.676
R1083 B.n373 B.n317 71.676
R1084 B.n369 B.n318 71.676
R1085 B.n365 B.n319 71.676
R1086 B.n360 B.n320 71.676
R1087 B.n356 B.n321 71.676
R1088 B.n352 B.n322 71.676
R1089 B.n348 B.n323 71.676
R1090 B.n344 B.n324 71.676
R1091 B.n340 B.n325 71.676
R1092 B.n336 B.n326 71.676
R1093 B.n649 B.n648 71.676
R1094 B.n128 B.n103 71.676
R1095 B.n132 B.n104 71.676
R1096 B.n136 B.n105 71.676
R1097 B.n140 B.n106 71.676
R1098 B.n144 B.n107 71.676
R1099 B.n148 B.n108 71.676
R1100 B.n152 B.n109 71.676
R1101 B.n157 B.n110 71.676
R1102 B.n161 B.n111 71.676
R1103 B.n165 B.n112 71.676
R1104 B.n169 B.n113 71.676
R1105 B.n173 B.n114 71.676
R1106 B.n177 B.n115 71.676
R1107 B.n181 B.n116 71.676
R1108 B.n185 B.n117 71.676
R1109 B.n189 B.n118 71.676
R1110 B.n193 B.n119 71.676
R1111 B.n197 B.n120 71.676
R1112 B.n121 B.n120 71.676
R1113 B.n196 B.n119 71.676
R1114 B.n192 B.n118 71.676
R1115 B.n188 B.n117 71.676
R1116 B.n184 B.n116 71.676
R1117 B.n180 B.n115 71.676
R1118 B.n176 B.n114 71.676
R1119 B.n172 B.n113 71.676
R1120 B.n168 B.n112 71.676
R1121 B.n164 B.n111 71.676
R1122 B.n160 B.n110 71.676
R1123 B.n156 B.n109 71.676
R1124 B.n151 B.n108 71.676
R1125 B.n147 B.n107 71.676
R1126 B.n143 B.n106 71.676
R1127 B.n139 B.n105 71.676
R1128 B.n135 B.n104 71.676
R1129 B.n131 B.n103 71.676
R1130 B.n648 B.n102 71.676
R1131 B.n408 B.n308 71.676
R1132 B.n402 B.n309 71.676
R1133 B.n398 B.n310 71.676
R1134 B.n394 B.n311 71.676
R1135 B.n390 B.n312 71.676
R1136 B.n386 B.n313 71.676
R1137 B.n382 B.n314 71.676
R1138 B.n378 B.n315 71.676
R1139 B.n374 B.n316 71.676
R1140 B.n370 B.n317 71.676
R1141 B.n366 B.n318 71.676
R1142 B.n361 B.n319 71.676
R1143 B.n357 B.n320 71.676
R1144 B.n353 B.n321 71.676
R1145 B.n349 B.n322 71.676
R1146 B.n345 B.n323 71.676
R1147 B.n341 B.n324 71.676
R1148 B.n337 B.n325 71.676
R1149 B.n333 B.n326 71.676
R1150 B.n363 B.n332 59.5399
R1151 B.n330 B.n329 59.5399
R1152 B.n154 B.n127 59.5399
R1153 B.n125 B.n124 59.5399
R1154 B.n553 B.t2 50.2785
R1155 B.n744 B.t4 50.2785
R1156 B.t2 B.n210 42.1253
R1157 B.t4 B.n15 42.1253
R1158 B.n651 B.n650 30.7517
R1159 B.n645 B.n644 30.7517
R1160 B.n334 B.n303 30.7517
R1161 B.n411 B.n410 30.7517
R1162 B.n438 B.t7 20.3835
R1163 B.t14 B.n670 20.3835
R1164 B B.n762 18.0485
R1165 B.t0 B.n234 14.948
R1166 B.t5 B.n36 14.948
R1167 B.n480 B.t3 12.2303
R1168 B.n60 B.t1 12.2303
R1169 B.n650 B.n101 10.6151
R1170 B.n129 B.n101 10.6151
R1171 B.n130 B.n129 10.6151
R1172 B.n133 B.n130 10.6151
R1173 B.n134 B.n133 10.6151
R1174 B.n137 B.n134 10.6151
R1175 B.n138 B.n137 10.6151
R1176 B.n141 B.n138 10.6151
R1177 B.n142 B.n141 10.6151
R1178 B.n145 B.n142 10.6151
R1179 B.n146 B.n145 10.6151
R1180 B.n149 B.n146 10.6151
R1181 B.n150 B.n149 10.6151
R1182 B.n153 B.n150 10.6151
R1183 B.n158 B.n155 10.6151
R1184 B.n159 B.n158 10.6151
R1185 B.n162 B.n159 10.6151
R1186 B.n163 B.n162 10.6151
R1187 B.n166 B.n163 10.6151
R1188 B.n167 B.n166 10.6151
R1189 B.n170 B.n167 10.6151
R1190 B.n171 B.n170 10.6151
R1191 B.n175 B.n174 10.6151
R1192 B.n178 B.n175 10.6151
R1193 B.n179 B.n178 10.6151
R1194 B.n182 B.n179 10.6151
R1195 B.n183 B.n182 10.6151
R1196 B.n186 B.n183 10.6151
R1197 B.n187 B.n186 10.6151
R1198 B.n190 B.n187 10.6151
R1199 B.n191 B.n190 10.6151
R1200 B.n194 B.n191 10.6151
R1201 B.n195 B.n194 10.6151
R1202 B.n198 B.n195 10.6151
R1203 B.n199 B.n198 10.6151
R1204 B.n645 B.n199 10.6151
R1205 B.n416 B.n303 10.6151
R1206 B.n417 B.n416 10.6151
R1207 B.n418 B.n417 10.6151
R1208 B.n418 B.n295 10.6151
R1209 B.n428 B.n295 10.6151
R1210 B.n429 B.n428 10.6151
R1211 B.n430 B.n429 10.6151
R1212 B.n430 B.n287 10.6151
R1213 B.n440 B.n287 10.6151
R1214 B.n441 B.n440 10.6151
R1215 B.n442 B.n441 10.6151
R1216 B.n442 B.n279 10.6151
R1217 B.n452 B.n279 10.6151
R1218 B.n453 B.n452 10.6151
R1219 B.n454 B.n453 10.6151
R1220 B.n454 B.n271 10.6151
R1221 B.n464 B.n271 10.6151
R1222 B.n465 B.n464 10.6151
R1223 B.n466 B.n465 10.6151
R1224 B.n466 B.n263 10.6151
R1225 B.n476 B.n263 10.6151
R1226 B.n477 B.n476 10.6151
R1227 B.n478 B.n477 10.6151
R1228 B.n478 B.n256 10.6151
R1229 B.n489 B.n256 10.6151
R1230 B.n490 B.n489 10.6151
R1231 B.n491 B.n490 10.6151
R1232 B.n491 B.n248 10.6151
R1233 B.n501 B.n248 10.6151
R1234 B.n502 B.n501 10.6151
R1235 B.n503 B.n502 10.6151
R1236 B.n503 B.n240 10.6151
R1237 B.n513 B.n240 10.6151
R1238 B.n514 B.n513 10.6151
R1239 B.n515 B.n514 10.6151
R1240 B.n515 B.n232 10.6151
R1241 B.n525 B.n232 10.6151
R1242 B.n526 B.n525 10.6151
R1243 B.n527 B.n526 10.6151
R1244 B.n527 B.n224 10.6151
R1245 B.n537 B.n224 10.6151
R1246 B.n538 B.n537 10.6151
R1247 B.n539 B.n538 10.6151
R1248 B.n539 B.n216 10.6151
R1249 B.n549 B.n216 10.6151
R1250 B.n550 B.n549 10.6151
R1251 B.n551 B.n550 10.6151
R1252 B.n551 B.n208 10.6151
R1253 B.n561 B.n208 10.6151
R1254 B.n562 B.n561 10.6151
R1255 B.n564 B.n562 10.6151
R1256 B.n564 B.n563 10.6151
R1257 B.n563 B.n200 10.6151
R1258 B.n575 B.n200 10.6151
R1259 B.n576 B.n575 10.6151
R1260 B.n577 B.n576 10.6151
R1261 B.n578 B.n577 10.6151
R1262 B.n580 B.n578 10.6151
R1263 B.n581 B.n580 10.6151
R1264 B.n582 B.n581 10.6151
R1265 B.n583 B.n582 10.6151
R1266 B.n585 B.n583 10.6151
R1267 B.n586 B.n585 10.6151
R1268 B.n587 B.n586 10.6151
R1269 B.n588 B.n587 10.6151
R1270 B.n590 B.n588 10.6151
R1271 B.n591 B.n590 10.6151
R1272 B.n592 B.n591 10.6151
R1273 B.n593 B.n592 10.6151
R1274 B.n595 B.n593 10.6151
R1275 B.n596 B.n595 10.6151
R1276 B.n597 B.n596 10.6151
R1277 B.n598 B.n597 10.6151
R1278 B.n600 B.n598 10.6151
R1279 B.n601 B.n600 10.6151
R1280 B.n602 B.n601 10.6151
R1281 B.n603 B.n602 10.6151
R1282 B.n605 B.n603 10.6151
R1283 B.n606 B.n605 10.6151
R1284 B.n607 B.n606 10.6151
R1285 B.n608 B.n607 10.6151
R1286 B.n610 B.n608 10.6151
R1287 B.n611 B.n610 10.6151
R1288 B.n612 B.n611 10.6151
R1289 B.n613 B.n612 10.6151
R1290 B.n615 B.n613 10.6151
R1291 B.n616 B.n615 10.6151
R1292 B.n617 B.n616 10.6151
R1293 B.n618 B.n617 10.6151
R1294 B.n620 B.n618 10.6151
R1295 B.n621 B.n620 10.6151
R1296 B.n622 B.n621 10.6151
R1297 B.n623 B.n622 10.6151
R1298 B.n625 B.n623 10.6151
R1299 B.n626 B.n625 10.6151
R1300 B.n627 B.n626 10.6151
R1301 B.n628 B.n627 10.6151
R1302 B.n630 B.n628 10.6151
R1303 B.n631 B.n630 10.6151
R1304 B.n632 B.n631 10.6151
R1305 B.n633 B.n632 10.6151
R1306 B.n635 B.n633 10.6151
R1307 B.n636 B.n635 10.6151
R1308 B.n637 B.n636 10.6151
R1309 B.n638 B.n637 10.6151
R1310 B.n640 B.n638 10.6151
R1311 B.n641 B.n640 10.6151
R1312 B.n642 B.n641 10.6151
R1313 B.n643 B.n642 10.6151
R1314 B.n644 B.n643 10.6151
R1315 B.n410 B.n307 10.6151
R1316 B.n405 B.n307 10.6151
R1317 B.n405 B.n404 10.6151
R1318 B.n404 B.n403 10.6151
R1319 B.n403 B.n400 10.6151
R1320 B.n400 B.n399 10.6151
R1321 B.n399 B.n396 10.6151
R1322 B.n396 B.n395 10.6151
R1323 B.n395 B.n392 10.6151
R1324 B.n392 B.n391 10.6151
R1325 B.n391 B.n388 10.6151
R1326 B.n388 B.n387 10.6151
R1327 B.n387 B.n384 10.6151
R1328 B.n384 B.n383 10.6151
R1329 B.n380 B.n379 10.6151
R1330 B.n379 B.n376 10.6151
R1331 B.n376 B.n375 10.6151
R1332 B.n375 B.n372 10.6151
R1333 B.n372 B.n371 10.6151
R1334 B.n371 B.n368 10.6151
R1335 B.n368 B.n367 10.6151
R1336 B.n367 B.n364 10.6151
R1337 B.n362 B.n359 10.6151
R1338 B.n359 B.n358 10.6151
R1339 B.n358 B.n355 10.6151
R1340 B.n355 B.n354 10.6151
R1341 B.n354 B.n351 10.6151
R1342 B.n351 B.n350 10.6151
R1343 B.n350 B.n347 10.6151
R1344 B.n347 B.n346 10.6151
R1345 B.n346 B.n343 10.6151
R1346 B.n343 B.n342 10.6151
R1347 B.n342 B.n339 10.6151
R1348 B.n339 B.n338 10.6151
R1349 B.n338 B.n335 10.6151
R1350 B.n335 B.n334 10.6151
R1351 B.n412 B.n411 10.6151
R1352 B.n412 B.n299 10.6151
R1353 B.n422 B.n299 10.6151
R1354 B.n423 B.n422 10.6151
R1355 B.n424 B.n423 10.6151
R1356 B.n424 B.n291 10.6151
R1357 B.n434 B.n291 10.6151
R1358 B.n435 B.n434 10.6151
R1359 B.n436 B.n435 10.6151
R1360 B.n436 B.n283 10.6151
R1361 B.n446 B.n283 10.6151
R1362 B.n447 B.n446 10.6151
R1363 B.n448 B.n447 10.6151
R1364 B.n448 B.n275 10.6151
R1365 B.n458 B.n275 10.6151
R1366 B.n459 B.n458 10.6151
R1367 B.n460 B.n459 10.6151
R1368 B.n460 B.n267 10.6151
R1369 B.n470 B.n267 10.6151
R1370 B.n471 B.n470 10.6151
R1371 B.n472 B.n471 10.6151
R1372 B.n472 B.n259 10.6151
R1373 B.n483 B.n259 10.6151
R1374 B.n484 B.n483 10.6151
R1375 B.n485 B.n484 10.6151
R1376 B.n485 B.n252 10.6151
R1377 B.n495 B.n252 10.6151
R1378 B.n496 B.n495 10.6151
R1379 B.n497 B.n496 10.6151
R1380 B.n497 B.n244 10.6151
R1381 B.n507 B.n244 10.6151
R1382 B.n508 B.n507 10.6151
R1383 B.n509 B.n508 10.6151
R1384 B.n509 B.n236 10.6151
R1385 B.n519 B.n236 10.6151
R1386 B.n520 B.n519 10.6151
R1387 B.n521 B.n520 10.6151
R1388 B.n521 B.n228 10.6151
R1389 B.n531 B.n228 10.6151
R1390 B.n532 B.n531 10.6151
R1391 B.n533 B.n532 10.6151
R1392 B.n533 B.n220 10.6151
R1393 B.n543 B.n220 10.6151
R1394 B.n544 B.n543 10.6151
R1395 B.n545 B.n544 10.6151
R1396 B.n545 B.n212 10.6151
R1397 B.n555 B.n212 10.6151
R1398 B.n556 B.n555 10.6151
R1399 B.n557 B.n556 10.6151
R1400 B.n557 B.n204 10.6151
R1401 B.n568 B.n204 10.6151
R1402 B.n569 B.n568 10.6151
R1403 B.n570 B.n569 10.6151
R1404 B.n570 B.n0 10.6151
R1405 B.n756 B.n1 10.6151
R1406 B.n756 B.n755 10.6151
R1407 B.n755 B.n754 10.6151
R1408 B.n754 B.n10 10.6151
R1409 B.n748 B.n10 10.6151
R1410 B.n748 B.n747 10.6151
R1411 B.n747 B.n746 10.6151
R1412 B.n746 B.n17 10.6151
R1413 B.n740 B.n17 10.6151
R1414 B.n740 B.n739 10.6151
R1415 B.n739 B.n738 10.6151
R1416 B.n738 B.n24 10.6151
R1417 B.n732 B.n24 10.6151
R1418 B.n732 B.n731 10.6151
R1419 B.n731 B.n730 10.6151
R1420 B.n730 B.n31 10.6151
R1421 B.n724 B.n31 10.6151
R1422 B.n724 B.n723 10.6151
R1423 B.n723 B.n722 10.6151
R1424 B.n722 B.n38 10.6151
R1425 B.n716 B.n38 10.6151
R1426 B.n716 B.n715 10.6151
R1427 B.n715 B.n714 10.6151
R1428 B.n714 B.n45 10.6151
R1429 B.n708 B.n45 10.6151
R1430 B.n708 B.n707 10.6151
R1431 B.n707 B.n706 10.6151
R1432 B.n706 B.n52 10.6151
R1433 B.n700 B.n52 10.6151
R1434 B.n700 B.n699 10.6151
R1435 B.n699 B.n698 10.6151
R1436 B.n698 B.n58 10.6151
R1437 B.n692 B.n58 10.6151
R1438 B.n692 B.n691 10.6151
R1439 B.n691 B.n690 10.6151
R1440 B.n690 B.n66 10.6151
R1441 B.n684 B.n66 10.6151
R1442 B.n684 B.n683 10.6151
R1443 B.n683 B.n682 10.6151
R1444 B.n682 B.n73 10.6151
R1445 B.n676 B.n73 10.6151
R1446 B.n676 B.n675 10.6151
R1447 B.n675 B.n674 10.6151
R1448 B.n674 B.n80 10.6151
R1449 B.n668 B.n80 10.6151
R1450 B.n668 B.n667 10.6151
R1451 B.n667 B.n666 10.6151
R1452 B.n666 B.n87 10.6151
R1453 B.n660 B.n87 10.6151
R1454 B.n660 B.n659 10.6151
R1455 B.n659 B.n658 10.6151
R1456 B.n658 B.n94 10.6151
R1457 B.n652 B.n94 10.6151
R1458 B.n652 B.n651 10.6151
R1459 B.n155 B.n154 6.5566
R1460 B.n171 B.n125 6.5566
R1461 B.n380 B.n330 6.5566
R1462 B.n364 B.n363 6.5566
R1463 B.n154 B.n153 4.05904
R1464 B.n174 B.n125 4.05904
R1465 B.n383 B.n330 4.05904
R1466 B.n363 B.n362 4.05904
R1467 B.n762 B.n0 2.81026
R1468 B.n762 B.n1 2.81026
R1469 VN.n38 VN.n37 161.3
R1470 VN.n36 VN.n21 161.3
R1471 VN.n35 VN.n34 161.3
R1472 VN.n33 VN.n22 161.3
R1473 VN.n32 VN.n31 161.3
R1474 VN.n30 VN.n23 161.3
R1475 VN.n29 VN.n28 161.3
R1476 VN.n27 VN.n24 161.3
R1477 VN.n18 VN.n17 161.3
R1478 VN.n16 VN.n1 161.3
R1479 VN.n15 VN.n14 161.3
R1480 VN.n13 VN.n2 161.3
R1481 VN.n12 VN.n11 161.3
R1482 VN.n10 VN.n3 161.3
R1483 VN.n9 VN.n8 161.3
R1484 VN.n7 VN.n4 161.3
R1485 VN.n19 VN.n0 78.9333
R1486 VN.n39 VN.n20 78.9333
R1487 VN.n6 VN.n5 62.5821
R1488 VN.n26 VN.n25 62.5821
R1489 VN.n11 VN.n2 56.5617
R1490 VN.n31 VN.n22 56.5617
R1491 VN.n26 VN.t3 52.2847
R1492 VN.n6 VN.t5 52.2847
R1493 VN VN.n39 46.1496
R1494 VN.n9 VN.n4 24.5923
R1495 VN.n10 VN.n9 24.5923
R1496 VN.n11 VN.n10 24.5923
R1497 VN.n15 VN.n2 24.5923
R1498 VN.n16 VN.n15 24.5923
R1499 VN.n17 VN.n16 24.5923
R1500 VN.n31 VN.n30 24.5923
R1501 VN.n30 VN.n29 24.5923
R1502 VN.n29 VN.n24 24.5923
R1503 VN.n37 VN.n36 24.5923
R1504 VN.n36 VN.n35 24.5923
R1505 VN.n35 VN.n22 24.5923
R1506 VN.n5 VN.t4 18.6202
R1507 VN.n0 VN.t0 18.6202
R1508 VN.n25 VN.t2 18.6202
R1509 VN.n20 VN.t1 18.6202
R1510 VN.n5 VN.n4 12.2964
R1511 VN.n25 VN.n24 12.2964
R1512 VN.n17 VN.n0 11.3127
R1513 VN.n37 VN.n20 11.3127
R1514 VN.n7 VN.n6 3.10331
R1515 VN.n27 VN.n26 3.1033
R1516 VN.n39 VN.n38 0.354861
R1517 VN.n19 VN.n18 0.354861
R1518 VN VN.n19 0.267071
R1519 VN.n38 VN.n21 0.189894
R1520 VN.n34 VN.n21 0.189894
R1521 VN.n34 VN.n33 0.189894
R1522 VN.n33 VN.n32 0.189894
R1523 VN.n32 VN.n23 0.189894
R1524 VN.n28 VN.n23 0.189894
R1525 VN.n28 VN.n27 0.189894
R1526 VN.n8 VN.n7 0.189894
R1527 VN.n8 VN.n3 0.189894
R1528 VN.n12 VN.n3 0.189894
R1529 VN.n13 VN.n12 0.189894
R1530 VN.n14 VN.n13 0.189894
R1531 VN.n14 VN.n1 0.189894
R1532 VN.n18 VN.n1 0.189894
R1533 VDD2.n1 VDD2.t0 91.5312
R1534 VDD2.n2 VDD2.t4 89.0135
R1535 VDD2.n1 VDD2.n0 82.7944
R1536 VDD2 VDD2.n3 82.7917
R1537 VDD2.n2 VDD2.n1 37.2972
R1538 VDD2.n3 VDD2.t3 7.02178
R1539 VDD2.n3 VDD2.t2 7.02178
R1540 VDD2.n0 VDD2.t1 7.02178
R1541 VDD2.n0 VDD2.t5 7.02178
R1542 VDD2 VDD2.n2 2.63197
C0 VP VDD2 0.553431f
C1 VDD1 VN 0.157943f
C2 VDD1 VTAIL 5.13082f
C3 VTAIL VN 3.10367f
C4 VDD1 VDD2 1.81662f
C5 VDD2 VN 1.97976f
C6 VTAIL VDD2 5.19106f
C7 VDD1 VP 2.37231f
C8 VP VN 6.24526f
C9 VP VTAIL 3.11785f
C10 VDD2 B 4.956527f
C11 VDD1 B 5.521129f
C12 VTAIL B 4.278261f
C13 VN B 15.00364f
C14 VP B 13.794811f
C15 VDD2.t0 B 0.347292f
C16 VDD2.t1 B 0.036348f
C17 VDD2.t5 B 0.036348f
C18 VDD2.n0 B 0.269641f
C19 VDD2.n1 B 1.79054f
C20 VDD2.t4 B 0.339421f
C21 VDD2.n2 B 1.51111f
C22 VDD2.t3 B 0.036348f
C23 VDD2.t2 B 0.036348f
C24 VDD2.n3 B 0.269623f
C25 VN.t0 B 0.547204f
C26 VN.n0 B 0.313922f
C27 VN.n1 B 0.021513f
C28 VN.n2 B 0.031868f
C29 VN.n3 B 0.021513f
C30 VN.n4 B 0.030046f
C31 VN.t4 B 0.547204f
C32 VN.n5 B 0.30127f
C33 VN.t5 B 0.799332f
C34 VN.n6 B 0.313094f
C35 VN.n7 B 0.268919f
C36 VN.n8 B 0.021513f
C37 VN.n9 B 0.039894f
C38 VN.n10 B 0.039894f
C39 VN.n11 B 0.030677f
C40 VN.n12 B 0.021513f
C41 VN.n13 B 0.021513f
C42 VN.n14 B 0.021513f
C43 VN.n15 B 0.039894f
C44 VN.n16 B 0.039894f
C45 VN.n17 B 0.029259f
C46 VN.n18 B 0.034716f
C47 VN.n19 B 0.058202f
C48 VN.t1 B 0.547204f
C49 VN.n20 B 0.313922f
C50 VN.n21 B 0.021513f
C51 VN.n22 B 0.031868f
C52 VN.n23 B 0.021513f
C53 VN.n24 B 0.030046f
C54 VN.t3 B 0.799332f
C55 VN.t2 B 0.547204f
C56 VN.n25 B 0.30127f
C57 VN.n26 B 0.313094f
C58 VN.n27 B 0.268919f
C59 VN.n28 B 0.021513f
C60 VN.n29 B 0.039894f
C61 VN.n30 B 0.039894f
C62 VN.n31 B 0.030677f
C63 VN.n32 B 0.021513f
C64 VN.n33 B 0.021513f
C65 VN.n34 B 0.021513f
C66 VN.n35 B 0.039894f
C67 VN.n36 B 0.039894f
C68 VN.n37 B 0.029259f
C69 VN.n38 B 0.034716f
C70 VN.n39 B 1.09934f
C71 VTAIL.t10 B 0.07506f
C72 VTAIL.t11 B 0.07506f
C73 VTAIL.n0 B 0.487565f
C74 VTAIL.n1 B 0.603162f
C75 VTAIL.t6 B 0.632363f
C76 VTAIL.n2 B 0.936044f
C77 VTAIL.t8 B 0.07506f
C78 VTAIL.t9 B 0.07506f
C79 VTAIL.n3 B 0.487565f
C80 VTAIL.n4 B 2.1051f
C81 VTAIL.t3 B 0.07506f
C82 VTAIL.t0 B 0.07506f
C83 VTAIL.n5 B 0.487567f
C84 VTAIL.n6 B 2.1051f
C85 VTAIL.t2 B 0.632365f
C86 VTAIL.n7 B 0.936041f
C87 VTAIL.t4 B 0.07506f
C88 VTAIL.t5 B 0.07506f
C89 VTAIL.n8 B 0.487567f
C90 VTAIL.n9 B 0.87613f
C91 VTAIL.t7 B 0.632363f
C92 VTAIL.n10 B 1.79263f
C93 VTAIL.t1 B 0.632363f
C94 VTAIL.n11 B 1.69322f
C95 VDD1.t3 B 0.495896f
C96 VDD1.t0 B 0.495165f
C97 VDD1.t2 B 0.051825f
C98 VDD1.t5 B 0.051825f
C99 VDD1.n0 B 0.384451f
C100 VDD1.n1 B 2.68413f
C101 VDD1.t4 B 0.051825f
C102 VDD1.t1 B 0.051825f
C103 VDD1.n2 B 0.379605f
C104 VDD1.n3 B 2.19204f
C105 VP.t3 B 0.690664f
C106 VP.n0 B 0.396222f
C107 VP.n1 B 0.027153f
C108 VP.n2 B 0.040222f
C109 VP.n3 B 0.027153f
C110 VP.n4 B 0.037924f
C111 VP.n5 B 0.027153f
C112 VP.n6 B 0.03872f
C113 VP.n7 B 0.027153f
C114 VP.n8 B 0.036929f
C115 VP.t2 B 0.690664f
C116 VP.n9 B 0.396222f
C117 VP.n10 B 0.027153f
C118 VP.n11 B 0.040222f
C119 VP.n12 B 0.027153f
C120 VP.n13 B 0.037924f
C121 VP.t5 B 1.00889f
C122 VP.t4 B 0.690664f
C123 VP.n14 B 0.380253f
C124 VP.n15 B 0.395178f
C125 VP.n16 B 0.339422f
C126 VP.n17 B 0.027153f
C127 VP.n18 B 0.050353f
C128 VP.n19 B 0.050353f
C129 VP.n20 B 0.03872f
C130 VP.n21 B 0.027153f
C131 VP.n22 B 0.027153f
C132 VP.n23 B 0.027153f
C133 VP.n24 B 0.050353f
C134 VP.n25 B 0.050353f
C135 VP.n26 B 0.036929f
C136 VP.n27 B 0.043817f
C137 VP.n28 B 1.37612f
C138 VP.t1 B 0.690664f
C139 VP.n29 B 0.396222f
C140 VP.n30 B 1.39741f
C141 VP.n31 B 0.043817f
C142 VP.n32 B 0.027153f
C143 VP.n33 B 0.050353f
C144 VP.n34 B 0.050353f
C145 VP.n35 B 0.040222f
C146 VP.n36 B 0.027153f
C147 VP.n37 B 0.027153f
C148 VP.n38 B 0.027153f
C149 VP.n39 B 0.050353f
C150 VP.n40 B 0.050353f
C151 VP.t0 B 0.690664f
C152 VP.n41 B 0.28594f
C153 VP.n42 B 0.037924f
C154 VP.n43 B 0.027153f
C155 VP.n44 B 0.027153f
C156 VP.n45 B 0.027153f
C157 VP.n46 B 0.050353f
C158 VP.n47 B 0.050353f
C159 VP.n48 B 0.03872f
C160 VP.n49 B 0.027153f
C161 VP.n50 B 0.027153f
C162 VP.n51 B 0.027153f
C163 VP.n52 B 0.050353f
C164 VP.n53 B 0.050353f
C165 VP.n54 B 0.036929f
C166 VP.n55 B 0.043817f
C167 VP.n56 B 0.073461f
.ends

