** sch_path: /home/lmadhu/openmpw/pdk_1/Project_gf180_tp/xschem/gmid_nfet.sch
**.subckt gmid_nfet
V1 vgs GND dc 3.3
.save i(v1)
V2 vgs vds dc 0
.save i(v2)
XM1 vds vgs GND GND nfet_03v3 L=0.28u W=1u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u'
+ pd='2*int((nf+1)/2) * (W/nf + 0.18u)' ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W'
+ sa=0 sb=0 sd=0 m=1
**** begin user architecture code
.lib /home/lmadhu/openmpw/pdk_1/gf180mcuA/libs.tech/ngspice/sm141064.ngspice typical

.include /home/lmadhu/openmpw/pdk_1/gf180mcuA/libs.tech/ngspice/design.ngspice
.param  sw_stat_mismatch = 0



*.dc v1 0 3.3 0.05
.save all
.control

run
*display
save @m.xm1.m0[gm]
save @m.xm1.m0[id]
save @m.xm1.m0[gds]
save @m.xm1.m0[vth]
save @m.xm1.m0[cgs]
save @m.xm1.m0[cgd]
save @m.xm1.m0[l]

let l_start = 0.5u
let l_stop  = 10u
let delta_l = 1u

let l_test = l_start
 while l_test le l_stop
  alter @m.xm1.m0[l] = l_test
  *op
  DC v1 0.01 3.3 0.01
  set filetype=binary
  write ./gmid/binary/data_L{$&l_test}.raw
   let l_test = l_test + delta_l
   let r = @m.xm1.m0[gm]/v2#branch
   let s = v2#branch/@m.xm1.m0[w]
   let gmd = @m.xm1.m0[gm]/1e-6
   let gain = abs(@m.xm1.m0[gm]/@m.xm1.m0[gds])
   let vov = vgs - @m.xm1.m0[vth]
   *plot r vs vov
   *plot gmd vs @m.xm1.m0[id]
 end
plot dc1.r dc2.r dc3.r dc4.r dc5.r dc6.r dc7.r
plot dc1.s vs dc1.r dc2.s vs dc2.r dc3.s vs dc3.r dc4.s vs dc4.r dc5.s vs dc5.r dc6.s vs dc6.r dc7.s
+ vs dc7.r retraceplot
plot dc1.gain vs dc1.r dc2.gain vs dc2.r dc3.gain vs dc3.r dc4.gain vs dc4.r dc5.gain vs dc5.r
+ dc6.gain vs dc6.r dc7.gain vs dc7.r
plot v2#branch
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
