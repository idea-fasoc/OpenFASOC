* NGSPICE file created from diff_pair_sample_1558.ext - technology: sky130A

.subckt diff_pair_sample_1558 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4164 pd=18.3 as=1.4454 ps=9.09 w=8.76 l=0.92
X1 VDD2.t5 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4164 pd=18.3 as=1.4454 ps=9.09 w=8.76 l=0.92
X2 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=3.4164 pd=18.3 as=0 ps=0 w=8.76 l=0.92
X3 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=3.4164 pd=18.3 as=0 ps=0 w=8.76 l=0.92
X4 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4164 pd=18.3 as=0 ps=0 w=8.76 l=0.92
X5 VTAIL.t7 VP.t1 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4454 pd=9.09 as=1.4454 ps=9.09 w=8.76 l=0.92
X6 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4164 pd=18.3 as=1.4454 ps=9.09 w=8.76 l=0.92
X7 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.4164 pd=18.3 as=0 ps=0 w=8.76 l=0.92
X8 VDD1.t3 VP.t2 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=3.4164 pd=18.3 as=1.4454 ps=9.09 w=8.76 l=0.92
X9 VTAIL.t6 VP.t3 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4454 pd=9.09 as=1.4454 ps=9.09 w=8.76 l=0.92
X10 VDD1.t1 VP.t4 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=1.4454 pd=9.09 as=3.4164 ps=18.3 w=8.76 l=0.92
X11 VDD2.t3 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4454 pd=9.09 as=3.4164 ps=18.3 w=8.76 l=0.92
X12 VTAIL.t3 VN.t3 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4454 pd=9.09 as=1.4454 ps=9.09 w=8.76 l=0.92
X13 VDD2.t1 VN.t4 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=1.4454 pd=9.09 as=3.4164 ps=18.3 w=8.76 l=0.92
X14 VTAIL.t4 VN.t5 VDD2.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4454 pd=9.09 as=1.4454 ps=9.09 w=8.76 l=0.92
X15 VDD1.t0 VP.t5 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4454 pd=9.09 as=3.4164 ps=18.3 w=8.76 l=0.92
R0 VP.n5 VP.t0 289.942
R1 VP.n12 VP.t2 272.173
R2 VP.n19 VP.t5 272.173
R3 VP.n9 VP.t4 272.173
R4 VP.n1 VP.t3 229.475
R5 VP.n4 VP.t1 229.475
R6 VP.n20 VP.n19 161.3
R7 VP.n7 VP.n6 161.3
R8 VP.n8 VP.n3 161.3
R9 VP.n10 VP.n9 161.3
R10 VP.n18 VP.n0 161.3
R11 VP.n17 VP.n16 161.3
R12 VP.n15 VP.n14 161.3
R13 VP.n13 VP.n2 161.3
R14 VP.n12 VP.n11 161.3
R15 VP.n14 VP.n13 52.6866
R16 VP.n18 VP.n17 52.6866
R17 VP.n8 VP.n7 52.6866
R18 VP.n6 VP.n5 43.4418
R19 VP.n5 VP.n4 42.5389
R20 VP.n11 VP.n10 39.6407
R21 VP.n14 VP.n1 12.2964
R22 VP.n17 VP.n1 12.2964
R23 VP.n7 VP.n4 12.2964
R24 VP.n13 VP.n12 5.84292
R25 VP.n19 VP.n18 5.84292
R26 VP.n9 VP.n8 5.84292
R27 VP.n6 VP.n3 0.189894
R28 VP.n10 VP.n3 0.189894
R29 VP.n11 VP.n2 0.189894
R30 VP.n15 VP.n2 0.189894
R31 VP.n16 VP.n15 0.189894
R32 VP.n16 VP.n0 0.189894
R33 VP.n20 VP.n0 0.189894
R34 VP VP.n20 0.0516364
R35 VTAIL.n194 VTAIL.n152 289.615
R36 VTAIL.n44 VTAIL.n2 289.615
R37 VTAIL.n146 VTAIL.n104 289.615
R38 VTAIL.n96 VTAIL.n54 289.615
R39 VTAIL.n169 VTAIL.n168 185
R40 VTAIL.n171 VTAIL.n170 185
R41 VTAIL.n164 VTAIL.n163 185
R42 VTAIL.n177 VTAIL.n176 185
R43 VTAIL.n179 VTAIL.n178 185
R44 VTAIL.n160 VTAIL.n159 185
R45 VTAIL.n185 VTAIL.n184 185
R46 VTAIL.n187 VTAIL.n186 185
R47 VTAIL.n156 VTAIL.n155 185
R48 VTAIL.n193 VTAIL.n192 185
R49 VTAIL.n195 VTAIL.n194 185
R50 VTAIL.n19 VTAIL.n18 185
R51 VTAIL.n21 VTAIL.n20 185
R52 VTAIL.n14 VTAIL.n13 185
R53 VTAIL.n27 VTAIL.n26 185
R54 VTAIL.n29 VTAIL.n28 185
R55 VTAIL.n10 VTAIL.n9 185
R56 VTAIL.n35 VTAIL.n34 185
R57 VTAIL.n37 VTAIL.n36 185
R58 VTAIL.n6 VTAIL.n5 185
R59 VTAIL.n43 VTAIL.n42 185
R60 VTAIL.n45 VTAIL.n44 185
R61 VTAIL.n147 VTAIL.n146 185
R62 VTAIL.n145 VTAIL.n144 185
R63 VTAIL.n108 VTAIL.n107 185
R64 VTAIL.n139 VTAIL.n138 185
R65 VTAIL.n137 VTAIL.n136 185
R66 VTAIL.n112 VTAIL.n111 185
R67 VTAIL.n131 VTAIL.n130 185
R68 VTAIL.n129 VTAIL.n128 185
R69 VTAIL.n116 VTAIL.n115 185
R70 VTAIL.n123 VTAIL.n122 185
R71 VTAIL.n121 VTAIL.n120 185
R72 VTAIL.n97 VTAIL.n96 185
R73 VTAIL.n95 VTAIL.n94 185
R74 VTAIL.n58 VTAIL.n57 185
R75 VTAIL.n89 VTAIL.n88 185
R76 VTAIL.n87 VTAIL.n86 185
R77 VTAIL.n62 VTAIL.n61 185
R78 VTAIL.n81 VTAIL.n80 185
R79 VTAIL.n79 VTAIL.n78 185
R80 VTAIL.n66 VTAIL.n65 185
R81 VTAIL.n73 VTAIL.n72 185
R82 VTAIL.n71 VTAIL.n70 185
R83 VTAIL.n69 VTAIL.t2 147.659
R84 VTAIL.n167 VTAIL.t11 147.659
R85 VTAIL.n17 VTAIL.t5 147.659
R86 VTAIL.n119 VTAIL.t10 147.659
R87 VTAIL.n170 VTAIL.n169 104.615
R88 VTAIL.n170 VTAIL.n163 104.615
R89 VTAIL.n177 VTAIL.n163 104.615
R90 VTAIL.n178 VTAIL.n177 104.615
R91 VTAIL.n178 VTAIL.n159 104.615
R92 VTAIL.n185 VTAIL.n159 104.615
R93 VTAIL.n186 VTAIL.n185 104.615
R94 VTAIL.n186 VTAIL.n155 104.615
R95 VTAIL.n193 VTAIL.n155 104.615
R96 VTAIL.n194 VTAIL.n193 104.615
R97 VTAIL.n20 VTAIL.n19 104.615
R98 VTAIL.n20 VTAIL.n13 104.615
R99 VTAIL.n27 VTAIL.n13 104.615
R100 VTAIL.n28 VTAIL.n27 104.615
R101 VTAIL.n28 VTAIL.n9 104.615
R102 VTAIL.n35 VTAIL.n9 104.615
R103 VTAIL.n36 VTAIL.n35 104.615
R104 VTAIL.n36 VTAIL.n5 104.615
R105 VTAIL.n43 VTAIL.n5 104.615
R106 VTAIL.n44 VTAIL.n43 104.615
R107 VTAIL.n146 VTAIL.n145 104.615
R108 VTAIL.n145 VTAIL.n107 104.615
R109 VTAIL.n138 VTAIL.n107 104.615
R110 VTAIL.n138 VTAIL.n137 104.615
R111 VTAIL.n137 VTAIL.n111 104.615
R112 VTAIL.n130 VTAIL.n111 104.615
R113 VTAIL.n130 VTAIL.n129 104.615
R114 VTAIL.n129 VTAIL.n115 104.615
R115 VTAIL.n122 VTAIL.n115 104.615
R116 VTAIL.n122 VTAIL.n121 104.615
R117 VTAIL.n96 VTAIL.n95 104.615
R118 VTAIL.n95 VTAIL.n57 104.615
R119 VTAIL.n88 VTAIL.n57 104.615
R120 VTAIL.n88 VTAIL.n87 104.615
R121 VTAIL.n87 VTAIL.n61 104.615
R122 VTAIL.n80 VTAIL.n61 104.615
R123 VTAIL.n80 VTAIL.n79 104.615
R124 VTAIL.n79 VTAIL.n65 104.615
R125 VTAIL.n72 VTAIL.n65 104.615
R126 VTAIL.n72 VTAIL.n71 104.615
R127 VTAIL.n169 VTAIL.t11 52.3082
R128 VTAIL.n19 VTAIL.t5 52.3082
R129 VTAIL.n121 VTAIL.t10 52.3082
R130 VTAIL.n71 VTAIL.t2 52.3082
R131 VTAIL.n103 VTAIL.n102 44.9321
R132 VTAIL.n53 VTAIL.n52 44.9321
R133 VTAIL.n1 VTAIL.n0 44.9319
R134 VTAIL.n51 VTAIL.n50 44.9319
R135 VTAIL.n199 VTAIL.n198 29.8581
R136 VTAIL.n49 VTAIL.n48 29.8581
R137 VTAIL.n151 VTAIL.n150 29.8581
R138 VTAIL.n101 VTAIL.n100 29.8581
R139 VTAIL.n53 VTAIL.n51 22.0738
R140 VTAIL.n199 VTAIL.n151 20.9962
R141 VTAIL.n168 VTAIL.n167 15.6677
R142 VTAIL.n18 VTAIL.n17 15.6677
R143 VTAIL.n120 VTAIL.n119 15.6677
R144 VTAIL.n70 VTAIL.n69 15.6677
R145 VTAIL.n171 VTAIL.n166 12.8005
R146 VTAIL.n21 VTAIL.n16 12.8005
R147 VTAIL.n123 VTAIL.n118 12.8005
R148 VTAIL.n73 VTAIL.n68 12.8005
R149 VTAIL.n172 VTAIL.n164 12.0247
R150 VTAIL.n22 VTAIL.n14 12.0247
R151 VTAIL.n124 VTAIL.n116 12.0247
R152 VTAIL.n74 VTAIL.n66 12.0247
R153 VTAIL.n176 VTAIL.n175 11.249
R154 VTAIL.n26 VTAIL.n25 11.249
R155 VTAIL.n128 VTAIL.n127 11.249
R156 VTAIL.n78 VTAIL.n77 11.249
R157 VTAIL.n179 VTAIL.n162 10.4732
R158 VTAIL.n29 VTAIL.n12 10.4732
R159 VTAIL.n131 VTAIL.n114 10.4732
R160 VTAIL.n81 VTAIL.n64 10.4732
R161 VTAIL.n180 VTAIL.n160 9.69747
R162 VTAIL.n30 VTAIL.n10 9.69747
R163 VTAIL.n132 VTAIL.n112 9.69747
R164 VTAIL.n82 VTAIL.n62 9.69747
R165 VTAIL.n198 VTAIL.n197 9.45567
R166 VTAIL.n48 VTAIL.n47 9.45567
R167 VTAIL.n150 VTAIL.n149 9.45567
R168 VTAIL.n100 VTAIL.n99 9.45567
R169 VTAIL.n191 VTAIL.n190 9.3005
R170 VTAIL.n154 VTAIL.n153 9.3005
R171 VTAIL.n197 VTAIL.n196 9.3005
R172 VTAIL.n158 VTAIL.n157 9.3005
R173 VTAIL.n183 VTAIL.n182 9.3005
R174 VTAIL.n181 VTAIL.n180 9.3005
R175 VTAIL.n162 VTAIL.n161 9.3005
R176 VTAIL.n175 VTAIL.n174 9.3005
R177 VTAIL.n173 VTAIL.n172 9.3005
R178 VTAIL.n166 VTAIL.n165 9.3005
R179 VTAIL.n189 VTAIL.n188 9.3005
R180 VTAIL.n41 VTAIL.n40 9.3005
R181 VTAIL.n4 VTAIL.n3 9.3005
R182 VTAIL.n47 VTAIL.n46 9.3005
R183 VTAIL.n8 VTAIL.n7 9.3005
R184 VTAIL.n33 VTAIL.n32 9.3005
R185 VTAIL.n31 VTAIL.n30 9.3005
R186 VTAIL.n12 VTAIL.n11 9.3005
R187 VTAIL.n25 VTAIL.n24 9.3005
R188 VTAIL.n23 VTAIL.n22 9.3005
R189 VTAIL.n16 VTAIL.n15 9.3005
R190 VTAIL.n39 VTAIL.n38 9.3005
R191 VTAIL.n106 VTAIL.n105 9.3005
R192 VTAIL.n143 VTAIL.n142 9.3005
R193 VTAIL.n141 VTAIL.n140 9.3005
R194 VTAIL.n110 VTAIL.n109 9.3005
R195 VTAIL.n135 VTAIL.n134 9.3005
R196 VTAIL.n133 VTAIL.n132 9.3005
R197 VTAIL.n114 VTAIL.n113 9.3005
R198 VTAIL.n127 VTAIL.n126 9.3005
R199 VTAIL.n125 VTAIL.n124 9.3005
R200 VTAIL.n118 VTAIL.n117 9.3005
R201 VTAIL.n149 VTAIL.n148 9.3005
R202 VTAIL.n56 VTAIL.n55 9.3005
R203 VTAIL.n99 VTAIL.n98 9.3005
R204 VTAIL.n93 VTAIL.n92 9.3005
R205 VTAIL.n91 VTAIL.n90 9.3005
R206 VTAIL.n60 VTAIL.n59 9.3005
R207 VTAIL.n85 VTAIL.n84 9.3005
R208 VTAIL.n83 VTAIL.n82 9.3005
R209 VTAIL.n64 VTAIL.n63 9.3005
R210 VTAIL.n77 VTAIL.n76 9.3005
R211 VTAIL.n75 VTAIL.n74 9.3005
R212 VTAIL.n68 VTAIL.n67 9.3005
R213 VTAIL.n184 VTAIL.n183 8.92171
R214 VTAIL.n198 VTAIL.n152 8.92171
R215 VTAIL.n34 VTAIL.n33 8.92171
R216 VTAIL.n48 VTAIL.n2 8.92171
R217 VTAIL.n150 VTAIL.n104 8.92171
R218 VTAIL.n136 VTAIL.n135 8.92171
R219 VTAIL.n100 VTAIL.n54 8.92171
R220 VTAIL.n86 VTAIL.n85 8.92171
R221 VTAIL.n187 VTAIL.n158 8.14595
R222 VTAIL.n196 VTAIL.n195 8.14595
R223 VTAIL.n37 VTAIL.n8 8.14595
R224 VTAIL.n46 VTAIL.n45 8.14595
R225 VTAIL.n148 VTAIL.n147 8.14595
R226 VTAIL.n139 VTAIL.n110 8.14595
R227 VTAIL.n98 VTAIL.n97 8.14595
R228 VTAIL.n89 VTAIL.n60 8.14595
R229 VTAIL.n188 VTAIL.n156 7.3702
R230 VTAIL.n192 VTAIL.n154 7.3702
R231 VTAIL.n38 VTAIL.n6 7.3702
R232 VTAIL.n42 VTAIL.n4 7.3702
R233 VTAIL.n144 VTAIL.n106 7.3702
R234 VTAIL.n140 VTAIL.n108 7.3702
R235 VTAIL.n94 VTAIL.n56 7.3702
R236 VTAIL.n90 VTAIL.n58 7.3702
R237 VTAIL.n191 VTAIL.n156 6.59444
R238 VTAIL.n192 VTAIL.n191 6.59444
R239 VTAIL.n41 VTAIL.n6 6.59444
R240 VTAIL.n42 VTAIL.n41 6.59444
R241 VTAIL.n144 VTAIL.n143 6.59444
R242 VTAIL.n143 VTAIL.n108 6.59444
R243 VTAIL.n94 VTAIL.n93 6.59444
R244 VTAIL.n93 VTAIL.n58 6.59444
R245 VTAIL.n188 VTAIL.n187 5.81868
R246 VTAIL.n195 VTAIL.n154 5.81868
R247 VTAIL.n38 VTAIL.n37 5.81868
R248 VTAIL.n45 VTAIL.n4 5.81868
R249 VTAIL.n147 VTAIL.n106 5.81868
R250 VTAIL.n140 VTAIL.n139 5.81868
R251 VTAIL.n97 VTAIL.n56 5.81868
R252 VTAIL.n90 VTAIL.n89 5.81868
R253 VTAIL.n184 VTAIL.n158 5.04292
R254 VTAIL.n196 VTAIL.n152 5.04292
R255 VTAIL.n34 VTAIL.n8 5.04292
R256 VTAIL.n46 VTAIL.n2 5.04292
R257 VTAIL.n148 VTAIL.n104 5.04292
R258 VTAIL.n136 VTAIL.n110 5.04292
R259 VTAIL.n98 VTAIL.n54 5.04292
R260 VTAIL.n86 VTAIL.n60 5.04292
R261 VTAIL.n167 VTAIL.n165 4.38563
R262 VTAIL.n17 VTAIL.n15 4.38563
R263 VTAIL.n119 VTAIL.n117 4.38563
R264 VTAIL.n69 VTAIL.n67 4.38563
R265 VTAIL.n183 VTAIL.n160 4.26717
R266 VTAIL.n33 VTAIL.n10 4.26717
R267 VTAIL.n135 VTAIL.n112 4.26717
R268 VTAIL.n85 VTAIL.n62 4.26717
R269 VTAIL.n180 VTAIL.n179 3.49141
R270 VTAIL.n30 VTAIL.n29 3.49141
R271 VTAIL.n132 VTAIL.n131 3.49141
R272 VTAIL.n82 VTAIL.n81 3.49141
R273 VTAIL.n176 VTAIL.n162 2.71565
R274 VTAIL.n26 VTAIL.n12 2.71565
R275 VTAIL.n128 VTAIL.n114 2.71565
R276 VTAIL.n78 VTAIL.n64 2.71565
R277 VTAIL.n0 VTAIL.t0 2.26077
R278 VTAIL.n0 VTAIL.t4 2.26077
R279 VTAIL.n50 VTAIL.t9 2.26077
R280 VTAIL.n50 VTAIL.t6 2.26077
R281 VTAIL.n102 VTAIL.t8 2.26077
R282 VTAIL.n102 VTAIL.t7 2.26077
R283 VTAIL.n52 VTAIL.t1 2.26077
R284 VTAIL.n52 VTAIL.t3 2.26077
R285 VTAIL.n175 VTAIL.n164 1.93989
R286 VTAIL.n25 VTAIL.n14 1.93989
R287 VTAIL.n127 VTAIL.n116 1.93989
R288 VTAIL.n77 VTAIL.n66 1.93989
R289 VTAIL.n172 VTAIL.n171 1.16414
R290 VTAIL.n22 VTAIL.n21 1.16414
R291 VTAIL.n124 VTAIL.n123 1.16414
R292 VTAIL.n74 VTAIL.n73 1.16414
R293 VTAIL.n101 VTAIL.n53 1.07809
R294 VTAIL.n151 VTAIL.n103 1.07809
R295 VTAIL.n51 VTAIL.n49 1.07809
R296 VTAIL.n103 VTAIL.n101 1.00912
R297 VTAIL.n49 VTAIL.n1 1.00912
R298 VTAIL VTAIL.n199 0.7505
R299 VTAIL.n168 VTAIL.n166 0.388379
R300 VTAIL.n18 VTAIL.n16 0.388379
R301 VTAIL.n120 VTAIL.n118 0.388379
R302 VTAIL.n70 VTAIL.n68 0.388379
R303 VTAIL VTAIL.n1 0.328086
R304 VTAIL.n173 VTAIL.n165 0.155672
R305 VTAIL.n174 VTAIL.n173 0.155672
R306 VTAIL.n174 VTAIL.n161 0.155672
R307 VTAIL.n181 VTAIL.n161 0.155672
R308 VTAIL.n182 VTAIL.n181 0.155672
R309 VTAIL.n182 VTAIL.n157 0.155672
R310 VTAIL.n189 VTAIL.n157 0.155672
R311 VTAIL.n190 VTAIL.n189 0.155672
R312 VTAIL.n190 VTAIL.n153 0.155672
R313 VTAIL.n197 VTAIL.n153 0.155672
R314 VTAIL.n23 VTAIL.n15 0.155672
R315 VTAIL.n24 VTAIL.n23 0.155672
R316 VTAIL.n24 VTAIL.n11 0.155672
R317 VTAIL.n31 VTAIL.n11 0.155672
R318 VTAIL.n32 VTAIL.n31 0.155672
R319 VTAIL.n32 VTAIL.n7 0.155672
R320 VTAIL.n39 VTAIL.n7 0.155672
R321 VTAIL.n40 VTAIL.n39 0.155672
R322 VTAIL.n40 VTAIL.n3 0.155672
R323 VTAIL.n47 VTAIL.n3 0.155672
R324 VTAIL.n149 VTAIL.n105 0.155672
R325 VTAIL.n142 VTAIL.n105 0.155672
R326 VTAIL.n142 VTAIL.n141 0.155672
R327 VTAIL.n141 VTAIL.n109 0.155672
R328 VTAIL.n134 VTAIL.n109 0.155672
R329 VTAIL.n134 VTAIL.n133 0.155672
R330 VTAIL.n133 VTAIL.n113 0.155672
R331 VTAIL.n126 VTAIL.n113 0.155672
R332 VTAIL.n126 VTAIL.n125 0.155672
R333 VTAIL.n125 VTAIL.n117 0.155672
R334 VTAIL.n99 VTAIL.n55 0.155672
R335 VTAIL.n92 VTAIL.n55 0.155672
R336 VTAIL.n92 VTAIL.n91 0.155672
R337 VTAIL.n91 VTAIL.n59 0.155672
R338 VTAIL.n84 VTAIL.n59 0.155672
R339 VTAIL.n84 VTAIL.n83 0.155672
R340 VTAIL.n83 VTAIL.n63 0.155672
R341 VTAIL.n76 VTAIL.n63 0.155672
R342 VTAIL.n76 VTAIL.n75 0.155672
R343 VTAIL.n75 VTAIL.n67 0.155672
R344 VDD1.n42 VDD1.n0 289.615
R345 VDD1.n89 VDD1.n47 289.615
R346 VDD1.n43 VDD1.n42 185
R347 VDD1.n41 VDD1.n40 185
R348 VDD1.n4 VDD1.n3 185
R349 VDD1.n35 VDD1.n34 185
R350 VDD1.n33 VDD1.n32 185
R351 VDD1.n8 VDD1.n7 185
R352 VDD1.n27 VDD1.n26 185
R353 VDD1.n25 VDD1.n24 185
R354 VDD1.n12 VDD1.n11 185
R355 VDD1.n19 VDD1.n18 185
R356 VDD1.n17 VDD1.n16 185
R357 VDD1.n64 VDD1.n63 185
R358 VDD1.n66 VDD1.n65 185
R359 VDD1.n59 VDD1.n58 185
R360 VDD1.n72 VDD1.n71 185
R361 VDD1.n74 VDD1.n73 185
R362 VDD1.n55 VDD1.n54 185
R363 VDD1.n80 VDD1.n79 185
R364 VDD1.n82 VDD1.n81 185
R365 VDD1.n51 VDD1.n50 185
R366 VDD1.n88 VDD1.n87 185
R367 VDD1.n90 VDD1.n89 185
R368 VDD1.n15 VDD1.t5 147.659
R369 VDD1.n62 VDD1.t3 147.659
R370 VDD1.n42 VDD1.n41 104.615
R371 VDD1.n41 VDD1.n3 104.615
R372 VDD1.n34 VDD1.n3 104.615
R373 VDD1.n34 VDD1.n33 104.615
R374 VDD1.n33 VDD1.n7 104.615
R375 VDD1.n26 VDD1.n7 104.615
R376 VDD1.n26 VDD1.n25 104.615
R377 VDD1.n25 VDD1.n11 104.615
R378 VDD1.n18 VDD1.n11 104.615
R379 VDD1.n18 VDD1.n17 104.615
R380 VDD1.n65 VDD1.n64 104.615
R381 VDD1.n65 VDD1.n58 104.615
R382 VDD1.n72 VDD1.n58 104.615
R383 VDD1.n73 VDD1.n72 104.615
R384 VDD1.n73 VDD1.n54 104.615
R385 VDD1.n80 VDD1.n54 104.615
R386 VDD1.n81 VDD1.n80 104.615
R387 VDD1.n81 VDD1.n50 104.615
R388 VDD1.n88 VDD1.n50 104.615
R389 VDD1.n89 VDD1.n88 104.615
R390 VDD1.n95 VDD1.n94 61.8248
R391 VDD1.n97 VDD1.n96 61.6109
R392 VDD1.n17 VDD1.t5 52.3082
R393 VDD1.n64 VDD1.t3 52.3082
R394 VDD1 VDD1.n46 47.4032
R395 VDD1.n95 VDD1.n93 47.2897
R396 VDD1.n97 VDD1.n95 35.891
R397 VDD1.n16 VDD1.n15 15.6677
R398 VDD1.n63 VDD1.n62 15.6677
R399 VDD1.n19 VDD1.n14 12.8005
R400 VDD1.n66 VDD1.n61 12.8005
R401 VDD1.n20 VDD1.n12 12.0247
R402 VDD1.n67 VDD1.n59 12.0247
R403 VDD1.n24 VDD1.n23 11.249
R404 VDD1.n71 VDD1.n70 11.249
R405 VDD1.n27 VDD1.n10 10.4732
R406 VDD1.n74 VDD1.n57 10.4732
R407 VDD1.n28 VDD1.n8 9.69747
R408 VDD1.n75 VDD1.n55 9.69747
R409 VDD1.n46 VDD1.n45 9.45567
R410 VDD1.n93 VDD1.n92 9.45567
R411 VDD1.n2 VDD1.n1 9.3005
R412 VDD1.n45 VDD1.n44 9.3005
R413 VDD1.n39 VDD1.n38 9.3005
R414 VDD1.n37 VDD1.n36 9.3005
R415 VDD1.n6 VDD1.n5 9.3005
R416 VDD1.n31 VDD1.n30 9.3005
R417 VDD1.n29 VDD1.n28 9.3005
R418 VDD1.n10 VDD1.n9 9.3005
R419 VDD1.n23 VDD1.n22 9.3005
R420 VDD1.n21 VDD1.n20 9.3005
R421 VDD1.n14 VDD1.n13 9.3005
R422 VDD1.n86 VDD1.n85 9.3005
R423 VDD1.n49 VDD1.n48 9.3005
R424 VDD1.n92 VDD1.n91 9.3005
R425 VDD1.n53 VDD1.n52 9.3005
R426 VDD1.n78 VDD1.n77 9.3005
R427 VDD1.n76 VDD1.n75 9.3005
R428 VDD1.n57 VDD1.n56 9.3005
R429 VDD1.n70 VDD1.n69 9.3005
R430 VDD1.n68 VDD1.n67 9.3005
R431 VDD1.n61 VDD1.n60 9.3005
R432 VDD1.n84 VDD1.n83 9.3005
R433 VDD1.n46 VDD1.n0 8.92171
R434 VDD1.n32 VDD1.n31 8.92171
R435 VDD1.n79 VDD1.n78 8.92171
R436 VDD1.n93 VDD1.n47 8.92171
R437 VDD1.n44 VDD1.n43 8.14595
R438 VDD1.n35 VDD1.n6 8.14595
R439 VDD1.n82 VDD1.n53 8.14595
R440 VDD1.n91 VDD1.n90 8.14595
R441 VDD1.n40 VDD1.n2 7.3702
R442 VDD1.n36 VDD1.n4 7.3702
R443 VDD1.n83 VDD1.n51 7.3702
R444 VDD1.n87 VDD1.n49 7.3702
R445 VDD1.n40 VDD1.n39 6.59444
R446 VDD1.n39 VDD1.n4 6.59444
R447 VDD1.n86 VDD1.n51 6.59444
R448 VDD1.n87 VDD1.n86 6.59444
R449 VDD1.n43 VDD1.n2 5.81868
R450 VDD1.n36 VDD1.n35 5.81868
R451 VDD1.n83 VDD1.n82 5.81868
R452 VDD1.n90 VDD1.n49 5.81868
R453 VDD1.n44 VDD1.n0 5.04292
R454 VDD1.n32 VDD1.n6 5.04292
R455 VDD1.n79 VDD1.n53 5.04292
R456 VDD1.n91 VDD1.n47 5.04292
R457 VDD1.n15 VDD1.n13 4.38563
R458 VDD1.n62 VDD1.n60 4.38563
R459 VDD1.n31 VDD1.n8 4.26717
R460 VDD1.n78 VDD1.n55 4.26717
R461 VDD1.n28 VDD1.n27 3.49141
R462 VDD1.n75 VDD1.n74 3.49141
R463 VDD1.n24 VDD1.n10 2.71565
R464 VDD1.n71 VDD1.n57 2.71565
R465 VDD1.n96 VDD1.t4 2.26077
R466 VDD1.n96 VDD1.t1 2.26077
R467 VDD1.n94 VDD1.t2 2.26077
R468 VDD1.n94 VDD1.t0 2.26077
R469 VDD1.n23 VDD1.n12 1.93989
R470 VDD1.n70 VDD1.n59 1.93989
R471 VDD1.n20 VDD1.n19 1.16414
R472 VDD1.n67 VDD1.n66 1.16414
R473 VDD1.n16 VDD1.n14 0.388379
R474 VDD1.n63 VDD1.n61 0.388379
R475 VDD1 VDD1.n97 0.211707
R476 VDD1.n45 VDD1.n1 0.155672
R477 VDD1.n38 VDD1.n1 0.155672
R478 VDD1.n38 VDD1.n37 0.155672
R479 VDD1.n37 VDD1.n5 0.155672
R480 VDD1.n30 VDD1.n5 0.155672
R481 VDD1.n30 VDD1.n29 0.155672
R482 VDD1.n29 VDD1.n9 0.155672
R483 VDD1.n22 VDD1.n9 0.155672
R484 VDD1.n22 VDD1.n21 0.155672
R485 VDD1.n21 VDD1.n13 0.155672
R486 VDD1.n68 VDD1.n60 0.155672
R487 VDD1.n69 VDD1.n68 0.155672
R488 VDD1.n69 VDD1.n56 0.155672
R489 VDD1.n76 VDD1.n56 0.155672
R490 VDD1.n77 VDD1.n76 0.155672
R491 VDD1.n77 VDD1.n52 0.155672
R492 VDD1.n84 VDD1.n52 0.155672
R493 VDD1.n85 VDD1.n84 0.155672
R494 VDD1.n85 VDD1.n48 0.155672
R495 VDD1.n92 VDD1.n48 0.155672
R496 B.n564 B.n563 585
R497 B.n230 B.n82 585
R498 B.n229 B.n228 585
R499 B.n227 B.n226 585
R500 B.n225 B.n224 585
R501 B.n223 B.n222 585
R502 B.n221 B.n220 585
R503 B.n219 B.n218 585
R504 B.n217 B.n216 585
R505 B.n215 B.n214 585
R506 B.n213 B.n212 585
R507 B.n211 B.n210 585
R508 B.n209 B.n208 585
R509 B.n207 B.n206 585
R510 B.n205 B.n204 585
R511 B.n203 B.n202 585
R512 B.n201 B.n200 585
R513 B.n199 B.n198 585
R514 B.n197 B.n196 585
R515 B.n195 B.n194 585
R516 B.n193 B.n192 585
R517 B.n191 B.n190 585
R518 B.n189 B.n188 585
R519 B.n187 B.n186 585
R520 B.n185 B.n184 585
R521 B.n183 B.n182 585
R522 B.n181 B.n180 585
R523 B.n179 B.n178 585
R524 B.n177 B.n176 585
R525 B.n175 B.n174 585
R526 B.n173 B.n172 585
R527 B.n171 B.n170 585
R528 B.n169 B.n168 585
R529 B.n167 B.n166 585
R530 B.n165 B.n164 585
R531 B.n163 B.n162 585
R532 B.n161 B.n160 585
R533 B.n159 B.n158 585
R534 B.n157 B.n156 585
R535 B.n155 B.n154 585
R536 B.n153 B.n152 585
R537 B.n151 B.n150 585
R538 B.n149 B.n148 585
R539 B.n147 B.n146 585
R540 B.n145 B.n144 585
R541 B.n143 B.n142 585
R542 B.n141 B.n140 585
R543 B.n139 B.n138 585
R544 B.n137 B.n136 585
R545 B.n135 B.n134 585
R546 B.n133 B.n132 585
R547 B.n131 B.n130 585
R548 B.n129 B.n128 585
R549 B.n127 B.n126 585
R550 B.n125 B.n124 585
R551 B.n123 B.n122 585
R552 B.n121 B.n120 585
R553 B.n119 B.n118 585
R554 B.n117 B.n116 585
R555 B.n115 B.n114 585
R556 B.n113 B.n112 585
R557 B.n111 B.n110 585
R558 B.n109 B.n108 585
R559 B.n107 B.n106 585
R560 B.n105 B.n104 585
R561 B.n103 B.n102 585
R562 B.n101 B.n100 585
R563 B.n99 B.n98 585
R564 B.n97 B.n96 585
R565 B.n95 B.n94 585
R566 B.n93 B.n92 585
R567 B.n91 B.n90 585
R568 B.n46 B.n45 585
R569 B.n569 B.n568 585
R570 B.n562 B.n83 585
R571 B.n83 B.n43 585
R572 B.n561 B.n42 585
R573 B.n573 B.n42 585
R574 B.n560 B.n41 585
R575 B.n574 B.n41 585
R576 B.n559 B.n40 585
R577 B.n575 B.n40 585
R578 B.n558 B.n557 585
R579 B.n557 B.n36 585
R580 B.n556 B.n35 585
R581 B.n581 B.n35 585
R582 B.n555 B.n34 585
R583 B.n582 B.n34 585
R584 B.n554 B.n33 585
R585 B.n583 B.n33 585
R586 B.n553 B.n552 585
R587 B.n552 B.n29 585
R588 B.n551 B.n28 585
R589 B.n589 B.n28 585
R590 B.n550 B.n27 585
R591 B.n590 B.n27 585
R592 B.n549 B.n26 585
R593 B.n591 B.n26 585
R594 B.n548 B.n547 585
R595 B.n547 B.n25 585
R596 B.n546 B.n21 585
R597 B.n597 B.n21 585
R598 B.n545 B.n20 585
R599 B.n598 B.n20 585
R600 B.n544 B.n19 585
R601 B.n599 B.n19 585
R602 B.n543 B.n542 585
R603 B.n542 B.n15 585
R604 B.n541 B.n14 585
R605 B.n605 B.n14 585
R606 B.n540 B.n13 585
R607 B.n606 B.n13 585
R608 B.n539 B.n12 585
R609 B.n607 B.n12 585
R610 B.n538 B.n537 585
R611 B.n537 B.n8 585
R612 B.n536 B.n7 585
R613 B.n613 B.n7 585
R614 B.n535 B.n6 585
R615 B.n614 B.n6 585
R616 B.n534 B.n5 585
R617 B.n615 B.n5 585
R618 B.n533 B.n532 585
R619 B.n532 B.n4 585
R620 B.n531 B.n231 585
R621 B.n531 B.n530 585
R622 B.n521 B.n232 585
R623 B.n233 B.n232 585
R624 B.n523 B.n522 585
R625 B.n524 B.n523 585
R626 B.n520 B.n238 585
R627 B.n238 B.n237 585
R628 B.n519 B.n518 585
R629 B.n518 B.n517 585
R630 B.n240 B.n239 585
R631 B.n241 B.n240 585
R632 B.n510 B.n509 585
R633 B.n511 B.n510 585
R634 B.n508 B.n246 585
R635 B.n246 B.n245 585
R636 B.n507 B.n506 585
R637 B.n506 B.n505 585
R638 B.n248 B.n247 585
R639 B.n498 B.n248 585
R640 B.n497 B.n496 585
R641 B.n499 B.n497 585
R642 B.n495 B.n253 585
R643 B.n253 B.n252 585
R644 B.n494 B.n493 585
R645 B.n493 B.n492 585
R646 B.n255 B.n254 585
R647 B.n256 B.n255 585
R648 B.n485 B.n484 585
R649 B.n486 B.n485 585
R650 B.n483 B.n261 585
R651 B.n261 B.n260 585
R652 B.n482 B.n481 585
R653 B.n481 B.n480 585
R654 B.n263 B.n262 585
R655 B.n264 B.n263 585
R656 B.n473 B.n472 585
R657 B.n474 B.n473 585
R658 B.n471 B.n269 585
R659 B.n269 B.n268 585
R660 B.n470 B.n469 585
R661 B.n469 B.n468 585
R662 B.n271 B.n270 585
R663 B.n272 B.n271 585
R664 B.n464 B.n463 585
R665 B.n275 B.n274 585
R666 B.n460 B.n459 585
R667 B.n461 B.n460 585
R668 B.n458 B.n312 585
R669 B.n457 B.n456 585
R670 B.n455 B.n454 585
R671 B.n453 B.n452 585
R672 B.n451 B.n450 585
R673 B.n449 B.n448 585
R674 B.n447 B.n446 585
R675 B.n445 B.n444 585
R676 B.n443 B.n442 585
R677 B.n441 B.n440 585
R678 B.n439 B.n438 585
R679 B.n437 B.n436 585
R680 B.n435 B.n434 585
R681 B.n433 B.n432 585
R682 B.n431 B.n430 585
R683 B.n429 B.n428 585
R684 B.n427 B.n426 585
R685 B.n425 B.n424 585
R686 B.n423 B.n422 585
R687 B.n421 B.n420 585
R688 B.n419 B.n418 585
R689 B.n417 B.n416 585
R690 B.n415 B.n414 585
R691 B.n413 B.n412 585
R692 B.n411 B.n410 585
R693 B.n409 B.n408 585
R694 B.n407 B.n406 585
R695 B.n405 B.n404 585
R696 B.n403 B.n402 585
R697 B.n400 B.n399 585
R698 B.n398 B.n397 585
R699 B.n396 B.n395 585
R700 B.n394 B.n393 585
R701 B.n392 B.n391 585
R702 B.n390 B.n389 585
R703 B.n388 B.n387 585
R704 B.n386 B.n385 585
R705 B.n384 B.n383 585
R706 B.n382 B.n381 585
R707 B.n379 B.n378 585
R708 B.n377 B.n376 585
R709 B.n375 B.n374 585
R710 B.n373 B.n372 585
R711 B.n371 B.n370 585
R712 B.n369 B.n368 585
R713 B.n367 B.n366 585
R714 B.n365 B.n364 585
R715 B.n363 B.n362 585
R716 B.n361 B.n360 585
R717 B.n359 B.n358 585
R718 B.n357 B.n356 585
R719 B.n355 B.n354 585
R720 B.n353 B.n352 585
R721 B.n351 B.n350 585
R722 B.n349 B.n348 585
R723 B.n347 B.n346 585
R724 B.n345 B.n344 585
R725 B.n343 B.n342 585
R726 B.n341 B.n340 585
R727 B.n339 B.n338 585
R728 B.n337 B.n336 585
R729 B.n335 B.n334 585
R730 B.n333 B.n332 585
R731 B.n331 B.n330 585
R732 B.n329 B.n328 585
R733 B.n327 B.n326 585
R734 B.n325 B.n324 585
R735 B.n323 B.n322 585
R736 B.n321 B.n320 585
R737 B.n319 B.n318 585
R738 B.n317 B.n311 585
R739 B.n461 B.n311 585
R740 B.n465 B.n273 585
R741 B.n273 B.n272 585
R742 B.n467 B.n466 585
R743 B.n468 B.n467 585
R744 B.n267 B.n266 585
R745 B.n268 B.n267 585
R746 B.n476 B.n475 585
R747 B.n475 B.n474 585
R748 B.n477 B.n265 585
R749 B.n265 B.n264 585
R750 B.n479 B.n478 585
R751 B.n480 B.n479 585
R752 B.n259 B.n258 585
R753 B.n260 B.n259 585
R754 B.n488 B.n487 585
R755 B.n487 B.n486 585
R756 B.n489 B.n257 585
R757 B.n257 B.n256 585
R758 B.n491 B.n490 585
R759 B.n492 B.n491 585
R760 B.n251 B.n250 585
R761 B.n252 B.n251 585
R762 B.n501 B.n500 585
R763 B.n500 B.n499 585
R764 B.n502 B.n249 585
R765 B.n498 B.n249 585
R766 B.n504 B.n503 585
R767 B.n505 B.n504 585
R768 B.n244 B.n243 585
R769 B.n245 B.n244 585
R770 B.n513 B.n512 585
R771 B.n512 B.n511 585
R772 B.n514 B.n242 585
R773 B.n242 B.n241 585
R774 B.n516 B.n515 585
R775 B.n517 B.n516 585
R776 B.n236 B.n235 585
R777 B.n237 B.n236 585
R778 B.n526 B.n525 585
R779 B.n525 B.n524 585
R780 B.n527 B.n234 585
R781 B.n234 B.n233 585
R782 B.n529 B.n528 585
R783 B.n530 B.n529 585
R784 B.n2 B.n0 585
R785 B.n4 B.n2 585
R786 B.n3 B.n1 585
R787 B.n614 B.n3 585
R788 B.n612 B.n611 585
R789 B.n613 B.n612 585
R790 B.n610 B.n9 585
R791 B.n9 B.n8 585
R792 B.n609 B.n608 585
R793 B.n608 B.n607 585
R794 B.n11 B.n10 585
R795 B.n606 B.n11 585
R796 B.n604 B.n603 585
R797 B.n605 B.n604 585
R798 B.n602 B.n16 585
R799 B.n16 B.n15 585
R800 B.n601 B.n600 585
R801 B.n600 B.n599 585
R802 B.n18 B.n17 585
R803 B.n598 B.n18 585
R804 B.n596 B.n595 585
R805 B.n597 B.n596 585
R806 B.n594 B.n22 585
R807 B.n25 B.n22 585
R808 B.n593 B.n592 585
R809 B.n592 B.n591 585
R810 B.n24 B.n23 585
R811 B.n590 B.n24 585
R812 B.n588 B.n587 585
R813 B.n589 B.n588 585
R814 B.n586 B.n30 585
R815 B.n30 B.n29 585
R816 B.n585 B.n584 585
R817 B.n584 B.n583 585
R818 B.n32 B.n31 585
R819 B.n582 B.n32 585
R820 B.n580 B.n579 585
R821 B.n581 B.n580 585
R822 B.n578 B.n37 585
R823 B.n37 B.n36 585
R824 B.n577 B.n576 585
R825 B.n576 B.n575 585
R826 B.n39 B.n38 585
R827 B.n574 B.n39 585
R828 B.n572 B.n571 585
R829 B.n573 B.n572 585
R830 B.n570 B.n44 585
R831 B.n44 B.n43 585
R832 B.n617 B.n616 585
R833 B.n616 B.n615 585
R834 B.n463 B.n273 449.257
R835 B.n568 B.n44 449.257
R836 B.n311 B.n271 449.257
R837 B.n564 B.n83 449.257
R838 B.n315 B.t13 431.825
R839 B.n313 B.t17 431.825
R840 B.n87 B.t10 431.825
R841 B.n84 B.t6 431.825
R842 B.n566 B.n565 256.663
R843 B.n566 B.n81 256.663
R844 B.n566 B.n80 256.663
R845 B.n566 B.n79 256.663
R846 B.n566 B.n78 256.663
R847 B.n566 B.n77 256.663
R848 B.n566 B.n76 256.663
R849 B.n566 B.n75 256.663
R850 B.n566 B.n74 256.663
R851 B.n566 B.n73 256.663
R852 B.n566 B.n72 256.663
R853 B.n566 B.n71 256.663
R854 B.n566 B.n70 256.663
R855 B.n566 B.n69 256.663
R856 B.n566 B.n68 256.663
R857 B.n566 B.n67 256.663
R858 B.n566 B.n66 256.663
R859 B.n566 B.n65 256.663
R860 B.n566 B.n64 256.663
R861 B.n566 B.n63 256.663
R862 B.n566 B.n62 256.663
R863 B.n566 B.n61 256.663
R864 B.n566 B.n60 256.663
R865 B.n566 B.n59 256.663
R866 B.n566 B.n58 256.663
R867 B.n566 B.n57 256.663
R868 B.n566 B.n56 256.663
R869 B.n566 B.n55 256.663
R870 B.n566 B.n54 256.663
R871 B.n566 B.n53 256.663
R872 B.n566 B.n52 256.663
R873 B.n566 B.n51 256.663
R874 B.n566 B.n50 256.663
R875 B.n566 B.n49 256.663
R876 B.n566 B.n48 256.663
R877 B.n566 B.n47 256.663
R878 B.n567 B.n566 256.663
R879 B.n462 B.n461 256.663
R880 B.n461 B.n276 256.663
R881 B.n461 B.n277 256.663
R882 B.n461 B.n278 256.663
R883 B.n461 B.n279 256.663
R884 B.n461 B.n280 256.663
R885 B.n461 B.n281 256.663
R886 B.n461 B.n282 256.663
R887 B.n461 B.n283 256.663
R888 B.n461 B.n284 256.663
R889 B.n461 B.n285 256.663
R890 B.n461 B.n286 256.663
R891 B.n461 B.n287 256.663
R892 B.n461 B.n288 256.663
R893 B.n461 B.n289 256.663
R894 B.n461 B.n290 256.663
R895 B.n461 B.n291 256.663
R896 B.n461 B.n292 256.663
R897 B.n461 B.n293 256.663
R898 B.n461 B.n294 256.663
R899 B.n461 B.n295 256.663
R900 B.n461 B.n296 256.663
R901 B.n461 B.n297 256.663
R902 B.n461 B.n298 256.663
R903 B.n461 B.n299 256.663
R904 B.n461 B.n300 256.663
R905 B.n461 B.n301 256.663
R906 B.n461 B.n302 256.663
R907 B.n461 B.n303 256.663
R908 B.n461 B.n304 256.663
R909 B.n461 B.n305 256.663
R910 B.n461 B.n306 256.663
R911 B.n461 B.n307 256.663
R912 B.n461 B.n308 256.663
R913 B.n461 B.n309 256.663
R914 B.n461 B.n310 256.663
R915 B.n315 B.t16 250.794
R916 B.n84 B.t8 250.794
R917 B.n313 B.t19 250.794
R918 B.n87 B.t11 250.794
R919 B.n316 B.t15 226.552
R920 B.n85 B.t9 226.552
R921 B.n314 B.t18 226.552
R922 B.n88 B.t12 226.552
R923 B.n467 B.n273 163.367
R924 B.n467 B.n267 163.367
R925 B.n475 B.n267 163.367
R926 B.n475 B.n265 163.367
R927 B.n479 B.n265 163.367
R928 B.n479 B.n259 163.367
R929 B.n487 B.n259 163.367
R930 B.n487 B.n257 163.367
R931 B.n491 B.n257 163.367
R932 B.n491 B.n251 163.367
R933 B.n500 B.n251 163.367
R934 B.n500 B.n249 163.367
R935 B.n504 B.n249 163.367
R936 B.n504 B.n244 163.367
R937 B.n512 B.n244 163.367
R938 B.n512 B.n242 163.367
R939 B.n516 B.n242 163.367
R940 B.n516 B.n236 163.367
R941 B.n525 B.n236 163.367
R942 B.n525 B.n234 163.367
R943 B.n529 B.n234 163.367
R944 B.n529 B.n2 163.367
R945 B.n616 B.n2 163.367
R946 B.n616 B.n3 163.367
R947 B.n612 B.n3 163.367
R948 B.n612 B.n9 163.367
R949 B.n608 B.n9 163.367
R950 B.n608 B.n11 163.367
R951 B.n604 B.n11 163.367
R952 B.n604 B.n16 163.367
R953 B.n600 B.n16 163.367
R954 B.n600 B.n18 163.367
R955 B.n596 B.n18 163.367
R956 B.n596 B.n22 163.367
R957 B.n592 B.n22 163.367
R958 B.n592 B.n24 163.367
R959 B.n588 B.n24 163.367
R960 B.n588 B.n30 163.367
R961 B.n584 B.n30 163.367
R962 B.n584 B.n32 163.367
R963 B.n580 B.n32 163.367
R964 B.n580 B.n37 163.367
R965 B.n576 B.n37 163.367
R966 B.n576 B.n39 163.367
R967 B.n572 B.n39 163.367
R968 B.n572 B.n44 163.367
R969 B.n460 B.n275 163.367
R970 B.n460 B.n312 163.367
R971 B.n456 B.n455 163.367
R972 B.n452 B.n451 163.367
R973 B.n448 B.n447 163.367
R974 B.n444 B.n443 163.367
R975 B.n440 B.n439 163.367
R976 B.n436 B.n435 163.367
R977 B.n432 B.n431 163.367
R978 B.n428 B.n427 163.367
R979 B.n424 B.n423 163.367
R980 B.n420 B.n419 163.367
R981 B.n416 B.n415 163.367
R982 B.n412 B.n411 163.367
R983 B.n408 B.n407 163.367
R984 B.n404 B.n403 163.367
R985 B.n399 B.n398 163.367
R986 B.n395 B.n394 163.367
R987 B.n391 B.n390 163.367
R988 B.n387 B.n386 163.367
R989 B.n383 B.n382 163.367
R990 B.n378 B.n377 163.367
R991 B.n374 B.n373 163.367
R992 B.n370 B.n369 163.367
R993 B.n366 B.n365 163.367
R994 B.n362 B.n361 163.367
R995 B.n358 B.n357 163.367
R996 B.n354 B.n353 163.367
R997 B.n350 B.n349 163.367
R998 B.n346 B.n345 163.367
R999 B.n342 B.n341 163.367
R1000 B.n338 B.n337 163.367
R1001 B.n334 B.n333 163.367
R1002 B.n330 B.n329 163.367
R1003 B.n326 B.n325 163.367
R1004 B.n322 B.n321 163.367
R1005 B.n318 B.n311 163.367
R1006 B.n469 B.n271 163.367
R1007 B.n469 B.n269 163.367
R1008 B.n473 B.n269 163.367
R1009 B.n473 B.n263 163.367
R1010 B.n481 B.n263 163.367
R1011 B.n481 B.n261 163.367
R1012 B.n485 B.n261 163.367
R1013 B.n485 B.n255 163.367
R1014 B.n493 B.n255 163.367
R1015 B.n493 B.n253 163.367
R1016 B.n497 B.n253 163.367
R1017 B.n497 B.n248 163.367
R1018 B.n506 B.n248 163.367
R1019 B.n506 B.n246 163.367
R1020 B.n510 B.n246 163.367
R1021 B.n510 B.n240 163.367
R1022 B.n518 B.n240 163.367
R1023 B.n518 B.n238 163.367
R1024 B.n523 B.n238 163.367
R1025 B.n523 B.n232 163.367
R1026 B.n531 B.n232 163.367
R1027 B.n532 B.n531 163.367
R1028 B.n532 B.n5 163.367
R1029 B.n6 B.n5 163.367
R1030 B.n7 B.n6 163.367
R1031 B.n537 B.n7 163.367
R1032 B.n537 B.n12 163.367
R1033 B.n13 B.n12 163.367
R1034 B.n14 B.n13 163.367
R1035 B.n542 B.n14 163.367
R1036 B.n542 B.n19 163.367
R1037 B.n20 B.n19 163.367
R1038 B.n21 B.n20 163.367
R1039 B.n547 B.n21 163.367
R1040 B.n547 B.n26 163.367
R1041 B.n27 B.n26 163.367
R1042 B.n28 B.n27 163.367
R1043 B.n552 B.n28 163.367
R1044 B.n552 B.n33 163.367
R1045 B.n34 B.n33 163.367
R1046 B.n35 B.n34 163.367
R1047 B.n557 B.n35 163.367
R1048 B.n557 B.n40 163.367
R1049 B.n41 B.n40 163.367
R1050 B.n42 B.n41 163.367
R1051 B.n83 B.n42 163.367
R1052 B.n90 B.n46 163.367
R1053 B.n94 B.n93 163.367
R1054 B.n98 B.n97 163.367
R1055 B.n102 B.n101 163.367
R1056 B.n106 B.n105 163.367
R1057 B.n110 B.n109 163.367
R1058 B.n114 B.n113 163.367
R1059 B.n118 B.n117 163.367
R1060 B.n122 B.n121 163.367
R1061 B.n126 B.n125 163.367
R1062 B.n130 B.n129 163.367
R1063 B.n134 B.n133 163.367
R1064 B.n138 B.n137 163.367
R1065 B.n142 B.n141 163.367
R1066 B.n146 B.n145 163.367
R1067 B.n150 B.n149 163.367
R1068 B.n154 B.n153 163.367
R1069 B.n158 B.n157 163.367
R1070 B.n162 B.n161 163.367
R1071 B.n166 B.n165 163.367
R1072 B.n170 B.n169 163.367
R1073 B.n174 B.n173 163.367
R1074 B.n178 B.n177 163.367
R1075 B.n182 B.n181 163.367
R1076 B.n186 B.n185 163.367
R1077 B.n190 B.n189 163.367
R1078 B.n194 B.n193 163.367
R1079 B.n198 B.n197 163.367
R1080 B.n202 B.n201 163.367
R1081 B.n206 B.n205 163.367
R1082 B.n210 B.n209 163.367
R1083 B.n214 B.n213 163.367
R1084 B.n218 B.n217 163.367
R1085 B.n222 B.n221 163.367
R1086 B.n226 B.n225 163.367
R1087 B.n228 B.n82 163.367
R1088 B.n461 B.n272 86.9973
R1089 B.n566 B.n43 86.9973
R1090 B.n463 B.n462 71.676
R1091 B.n312 B.n276 71.676
R1092 B.n455 B.n277 71.676
R1093 B.n451 B.n278 71.676
R1094 B.n447 B.n279 71.676
R1095 B.n443 B.n280 71.676
R1096 B.n439 B.n281 71.676
R1097 B.n435 B.n282 71.676
R1098 B.n431 B.n283 71.676
R1099 B.n427 B.n284 71.676
R1100 B.n423 B.n285 71.676
R1101 B.n419 B.n286 71.676
R1102 B.n415 B.n287 71.676
R1103 B.n411 B.n288 71.676
R1104 B.n407 B.n289 71.676
R1105 B.n403 B.n290 71.676
R1106 B.n398 B.n291 71.676
R1107 B.n394 B.n292 71.676
R1108 B.n390 B.n293 71.676
R1109 B.n386 B.n294 71.676
R1110 B.n382 B.n295 71.676
R1111 B.n377 B.n296 71.676
R1112 B.n373 B.n297 71.676
R1113 B.n369 B.n298 71.676
R1114 B.n365 B.n299 71.676
R1115 B.n361 B.n300 71.676
R1116 B.n357 B.n301 71.676
R1117 B.n353 B.n302 71.676
R1118 B.n349 B.n303 71.676
R1119 B.n345 B.n304 71.676
R1120 B.n341 B.n305 71.676
R1121 B.n337 B.n306 71.676
R1122 B.n333 B.n307 71.676
R1123 B.n329 B.n308 71.676
R1124 B.n325 B.n309 71.676
R1125 B.n321 B.n310 71.676
R1126 B.n568 B.n567 71.676
R1127 B.n90 B.n47 71.676
R1128 B.n94 B.n48 71.676
R1129 B.n98 B.n49 71.676
R1130 B.n102 B.n50 71.676
R1131 B.n106 B.n51 71.676
R1132 B.n110 B.n52 71.676
R1133 B.n114 B.n53 71.676
R1134 B.n118 B.n54 71.676
R1135 B.n122 B.n55 71.676
R1136 B.n126 B.n56 71.676
R1137 B.n130 B.n57 71.676
R1138 B.n134 B.n58 71.676
R1139 B.n138 B.n59 71.676
R1140 B.n142 B.n60 71.676
R1141 B.n146 B.n61 71.676
R1142 B.n150 B.n62 71.676
R1143 B.n154 B.n63 71.676
R1144 B.n158 B.n64 71.676
R1145 B.n162 B.n65 71.676
R1146 B.n166 B.n66 71.676
R1147 B.n170 B.n67 71.676
R1148 B.n174 B.n68 71.676
R1149 B.n178 B.n69 71.676
R1150 B.n182 B.n70 71.676
R1151 B.n186 B.n71 71.676
R1152 B.n190 B.n72 71.676
R1153 B.n194 B.n73 71.676
R1154 B.n198 B.n74 71.676
R1155 B.n202 B.n75 71.676
R1156 B.n206 B.n76 71.676
R1157 B.n210 B.n77 71.676
R1158 B.n214 B.n78 71.676
R1159 B.n218 B.n79 71.676
R1160 B.n222 B.n80 71.676
R1161 B.n226 B.n81 71.676
R1162 B.n565 B.n82 71.676
R1163 B.n565 B.n564 71.676
R1164 B.n228 B.n81 71.676
R1165 B.n225 B.n80 71.676
R1166 B.n221 B.n79 71.676
R1167 B.n217 B.n78 71.676
R1168 B.n213 B.n77 71.676
R1169 B.n209 B.n76 71.676
R1170 B.n205 B.n75 71.676
R1171 B.n201 B.n74 71.676
R1172 B.n197 B.n73 71.676
R1173 B.n193 B.n72 71.676
R1174 B.n189 B.n71 71.676
R1175 B.n185 B.n70 71.676
R1176 B.n181 B.n69 71.676
R1177 B.n177 B.n68 71.676
R1178 B.n173 B.n67 71.676
R1179 B.n169 B.n66 71.676
R1180 B.n165 B.n65 71.676
R1181 B.n161 B.n64 71.676
R1182 B.n157 B.n63 71.676
R1183 B.n153 B.n62 71.676
R1184 B.n149 B.n61 71.676
R1185 B.n145 B.n60 71.676
R1186 B.n141 B.n59 71.676
R1187 B.n137 B.n58 71.676
R1188 B.n133 B.n57 71.676
R1189 B.n129 B.n56 71.676
R1190 B.n125 B.n55 71.676
R1191 B.n121 B.n54 71.676
R1192 B.n117 B.n53 71.676
R1193 B.n113 B.n52 71.676
R1194 B.n109 B.n51 71.676
R1195 B.n105 B.n50 71.676
R1196 B.n101 B.n49 71.676
R1197 B.n97 B.n48 71.676
R1198 B.n93 B.n47 71.676
R1199 B.n567 B.n46 71.676
R1200 B.n462 B.n275 71.676
R1201 B.n456 B.n276 71.676
R1202 B.n452 B.n277 71.676
R1203 B.n448 B.n278 71.676
R1204 B.n444 B.n279 71.676
R1205 B.n440 B.n280 71.676
R1206 B.n436 B.n281 71.676
R1207 B.n432 B.n282 71.676
R1208 B.n428 B.n283 71.676
R1209 B.n424 B.n284 71.676
R1210 B.n420 B.n285 71.676
R1211 B.n416 B.n286 71.676
R1212 B.n412 B.n287 71.676
R1213 B.n408 B.n288 71.676
R1214 B.n404 B.n289 71.676
R1215 B.n399 B.n290 71.676
R1216 B.n395 B.n291 71.676
R1217 B.n391 B.n292 71.676
R1218 B.n387 B.n293 71.676
R1219 B.n383 B.n294 71.676
R1220 B.n378 B.n295 71.676
R1221 B.n374 B.n296 71.676
R1222 B.n370 B.n297 71.676
R1223 B.n366 B.n298 71.676
R1224 B.n362 B.n299 71.676
R1225 B.n358 B.n300 71.676
R1226 B.n354 B.n301 71.676
R1227 B.n350 B.n302 71.676
R1228 B.n346 B.n303 71.676
R1229 B.n342 B.n304 71.676
R1230 B.n338 B.n305 71.676
R1231 B.n334 B.n306 71.676
R1232 B.n330 B.n307 71.676
R1233 B.n326 B.n308 71.676
R1234 B.n322 B.n309 71.676
R1235 B.n318 B.n310 71.676
R1236 B.n380 B.n316 59.5399
R1237 B.n401 B.n314 59.5399
R1238 B.n89 B.n88 59.5399
R1239 B.n86 B.n85 59.5399
R1240 B.n468 B.n272 53.2958
R1241 B.n468 B.n268 53.2958
R1242 B.n474 B.n268 53.2958
R1243 B.n474 B.n264 53.2958
R1244 B.n480 B.n264 53.2958
R1245 B.n486 B.n260 53.2958
R1246 B.n486 B.n256 53.2958
R1247 B.n492 B.n256 53.2958
R1248 B.n492 B.n252 53.2958
R1249 B.n499 B.n252 53.2958
R1250 B.n499 B.n498 53.2958
R1251 B.n505 B.n245 53.2958
R1252 B.n511 B.n245 53.2958
R1253 B.n517 B.n241 53.2958
R1254 B.n517 B.n237 53.2958
R1255 B.n524 B.n237 53.2958
R1256 B.n530 B.n233 53.2958
R1257 B.n530 B.n4 53.2958
R1258 B.n615 B.n4 53.2958
R1259 B.n615 B.n614 53.2958
R1260 B.n614 B.n613 53.2958
R1261 B.n613 B.n8 53.2958
R1262 B.n607 B.n606 53.2958
R1263 B.n606 B.n605 53.2958
R1264 B.n605 B.n15 53.2958
R1265 B.n599 B.n598 53.2958
R1266 B.n598 B.n597 53.2958
R1267 B.n591 B.n25 53.2958
R1268 B.n591 B.n590 53.2958
R1269 B.n590 B.n589 53.2958
R1270 B.n589 B.n29 53.2958
R1271 B.n583 B.n29 53.2958
R1272 B.n583 B.n582 53.2958
R1273 B.n581 B.n36 53.2958
R1274 B.n575 B.n36 53.2958
R1275 B.n575 B.n574 53.2958
R1276 B.n574 B.n573 53.2958
R1277 B.n573 B.n43 53.2958
R1278 B.n511 B.t3 47.0258
R1279 B.n599 B.t4 47.0258
R1280 B.n505 B.t1 42.3233
R1281 B.n597 B.t5 42.3233
R1282 B.t14 B.n260 36.0532
R1283 B.n582 B.t7 36.0532
R1284 B.n524 B.t2 29.7832
R1285 B.n607 B.t0 29.7832
R1286 B.n570 B.n569 29.1907
R1287 B.n317 B.n270 29.1907
R1288 B.n465 B.n464 29.1907
R1289 B.n563 B.n562 29.1907
R1290 B.n316 B.n315 24.2429
R1291 B.n314 B.n313 24.2429
R1292 B.n88 B.n87 24.2429
R1293 B.n85 B.n84 24.2429
R1294 B.t2 B.n233 23.5131
R1295 B.t0 B.n8 23.5131
R1296 B B.n617 18.0485
R1297 B.n480 B.t14 17.2431
R1298 B.t7 B.n581 17.2431
R1299 B.n498 B.t1 10.9731
R1300 B.n25 B.t5 10.9731
R1301 B.n569 B.n45 10.6151
R1302 B.n91 B.n45 10.6151
R1303 B.n92 B.n91 10.6151
R1304 B.n95 B.n92 10.6151
R1305 B.n96 B.n95 10.6151
R1306 B.n99 B.n96 10.6151
R1307 B.n100 B.n99 10.6151
R1308 B.n103 B.n100 10.6151
R1309 B.n104 B.n103 10.6151
R1310 B.n107 B.n104 10.6151
R1311 B.n108 B.n107 10.6151
R1312 B.n111 B.n108 10.6151
R1313 B.n112 B.n111 10.6151
R1314 B.n115 B.n112 10.6151
R1315 B.n116 B.n115 10.6151
R1316 B.n119 B.n116 10.6151
R1317 B.n120 B.n119 10.6151
R1318 B.n123 B.n120 10.6151
R1319 B.n124 B.n123 10.6151
R1320 B.n127 B.n124 10.6151
R1321 B.n128 B.n127 10.6151
R1322 B.n131 B.n128 10.6151
R1323 B.n132 B.n131 10.6151
R1324 B.n135 B.n132 10.6151
R1325 B.n136 B.n135 10.6151
R1326 B.n139 B.n136 10.6151
R1327 B.n140 B.n139 10.6151
R1328 B.n143 B.n140 10.6151
R1329 B.n144 B.n143 10.6151
R1330 B.n147 B.n144 10.6151
R1331 B.n148 B.n147 10.6151
R1332 B.n152 B.n151 10.6151
R1333 B.n155 B.n152 10.6151
R1334 B.n156 B.n155 10.6151
R1335 B.n159 B.n156 10.6151
R1336 B.n160 B.n159 10.6151
R1337 B.n163 B.n160 10.6151
R1338 B.n164 B.n163 10.6151
R1339 B.n167 B.n164 10.6151
R1340 B.n168 B.n167 10.6151
R1341 B.n172 B.n171 10.6151
R1342 B.n175 B.n172 10.6151
R1343 B.n176 B.n175 10.6151
R1344 B.n179 B.n176 10.6151
R1345 B.n180 B.n179 10.6151
R1346 B.n183 B.n180 10.6151
R1347 B.n184 B.n183 10.6151
R1348 B.n187 B.n184 10.6151
R1349 B.n188 B.n187 10.6151
R1350 B.n191 B.n188 10.6151
R1351 B.n192 B.n191 10.6151
R1352 B.n195 B.n192 10.6151
R1353 B.n196 B.n195 10.6151
R1354 B.n199 B.n196 10.6151
R1355 B.n200 B.n199 10.6151
R1356 B.n203 B.n200 10.6151
R1357 B.n204 B.n203 10.6151
R1358 B.n207 B.n204 10.6151
R1359 B.n208 B.n207 10.6151
R1360 B.n211 B.n208 10.6151
R1361 B.n212 B.n211 10.6151
R1362 B.n215 B.n212 10.6151
R1363 B.n216 B.n215 10.6151
R1364 B.n219 B.n216 10.6151
R1365 B.n220 B.n219 10.6151
R1366 B.n223 B.n220 10.6151
R1367 B.n224 B.n223 10.6151
R1368 B.n227 B.n224 10.6151
R1369 B.n229 B.n227 10.6151
R1370 B.n230 B.n229 10.6151
R1371 B.n563 B.n230 10.6151
R1372 B.n470 B.n270 10.6151
R1373 B.n471 B.n470 10.6151
R1374 B.n472 B.n471 10.6151
R1375 B.n472 B.n262 10.6151
R1376 B.n482 B.n262 10.6151
R1377 B.n483 B.n482 10.6151
R1378 B.n484 B.n483 10.6151
R1379 B.n484 B.n254 10.6151
R1380 B.n494 B.n254 10.6151
R1381 B.n495 B.n494 10.6151
R1382 B.n496 B.n495 10.6151
R1383 B.n496 B.n247 10.6151
R1384 B.n507 B.n247 10.6151
R1385 B.n508 B.n507 10.6151
R1386 B.n509 B.n508 10.6151
R1387 B.n509 B.n239 10.6151
R1388 B.n519 B.n239 10.6151
R1389 B.n520 B.n519 10.6151
R1390 B.n522 B.n520 10.6151
R1391 B.n522 B.n521 10.6151
R1392 B.n521 B.n231 10.6151
R1393 B.n533 B.n231 10.6151
R1394 B.n534 B.n533 10.6151
R1395 B.n535 B.n534 10.6151
R1396 B.n536 B.n535 10.6151
R1397 B.n538 B.n536 10.6151
R1398 B.n539 B.n538 10.6151
R1399 B.n540 B.n539 10.6151
R1400 B.n541 B.n540 10.6151
R1401 B.n543 B.n541 10.6151
R1402 B.n544 B.n543 10.6151
R1403 B.n545 B.n544 10.6151
R1404 B.n546 B.n545 10.6151
R1405 B.n548 B.n546 10.6151
R1406 B.n549 B.n548 10.6151
R1407 B.n550 B.n549 10.6151
R1408 B.n551 B.n550 10.6151
R1409 B.n553 B.n551 10.6151
R1410 B.n554 B.n553 10.6151
R1411 B.n555 B.n554 10.6151
R1412 B.n556 B.n555 10.6151
R1413 B.n558 B.n556 10.6151
R1414 B.n559 B.n558 10.6151
R1415 B.n560 B.n559 10.6151
R1416 B.n561 B.n560 10.6151
R1417 B.n562 B.n561 10.6151
R1418 B.n464 B.n274 10.6151
R1419 B.n459 B.n274 10.6151
R1420 B.n459 B.n458 10.6151
R1421 B.n458 B.n457 10.6151
R1422 B.n457 B.n454 10.6151
R1423 B.n454 B.n453 10.6151
R1424 B.n453 B.n450 10.6151
R1425 B.n450 B.n449 10.6151
R1426 B.n449 B.n446 10.6151
R1427 B.n446 B.n445 10.6151
R1428 B.n445 B.n442 10.6151
R1429 B.n442 B.n441 10.6151
R1430 B.n441 B.n438 10.6151
R1431 B.n438 B.n437 10.6151
R1432 B.n437 B.n434 10.6151
R1433 B.n434 B.n433 10.6151
R1434 B.n433 B.n430 10.6151
R1435 B.n430 B.n429 10.6151
R1436 B.n429 B.n426 10.6151
R1437 B.n426 B.n425 10.6151
R1438 B.n425 B.n422 10.6151
R1439 B.n422 B.n421 10.6151
R1440 B.n421 B.n418 10.6151
R1441 B.n418 B.n417 10.6151
R1442 B.n417 B.n414 10.6151
R1443 B.n414 B.n413 10.6151
R1444 B.n413 B.n410 10.6151
R1445 B.n410 B.n409 10.6151
R1446 B.n409 B.n406 10.6151
R1447 B.n406 B.n405 10.6151
R1448 B.n405 B.n402 10.6151
R1449 B.n400 B.n397 10.6151
R1450 B.n397 B.n396 10.6151
R1451 B.n396 B.n393 10.6151
R1452 B.n393 B.n392 10.6151
R1453 B.n392 B.n389 10.6151
R1454 B.n389 B.n388 10.6151
R1455 B.n388 B.n385 10.6151
R1456 B.n385 B.n384 10.6151
R1457 B.n384 B.n381 10.6151
R1458 B.n379 B.n376 10.6151
R1459 B.n376 B.n375 10.6151
R1460 B.n375 B.n372 10.6151
R1461 B.n372 B.n371 10.6151
R1462 B.n371 B.n368 10.6151
R1463 B.n368 B.n367 10.6151
R1464 B.n367 B.n364 10.6151
R1465 B.n364 B.n363 10.6151
R1466 B.n363 B.n360 10.6151
R1467 B.n360 B.n359 10.6151
R1468 B.n359 B.n356 10.6151
R1469 B.n356 B.n355 10.6151
R1470 B.n355 B.n352 10.6151
R1471 B.n352 B.n351 10.6151
R1472 B.n351 B.n348 10.6151
R1473 B.n348 B.n347 10.6151
R1474 B.n347 B.n344 10.6151
R1475 B.n344 B.n343 10.6151
R1476 B.n343 B.n340 10.6151
R1477 B.n340 B.n339 10.6151
R1478 B.n339 B.n336 10.6151
R1479 B.n336 B.n335 10.6151
R1480 B.n335 B.n332 10.6151
R1481 B.n332 B.n331 10.6151
R1482 B.n331 B.n328 10.6151
R1483 B.n328 B.n327 10.6151
R1484 B.n327 B.n324 10.6151
R1485 B.n324 B.n323 10.6151
R1486 B.n323 B.n320 10.6151
R1487 B.n320 B.n319 10.6151
R1488 B.n319 B.n317 10.6151
R1489 B.n466 B.n465 10.6151
R1490 B.n466 B.n266 10.6151
R1491 B.n476 B.n266 10.6151
R1492 B.n477 B.n476 10.6151
R1493 B.n478 B.n477 10.6151
R1494 B.n478 B.n258 10.6151
R1495 B.n488 B.n258 10.6151
R1496 B.n489 B.n488 10.6151
R1497 B.n490 B.n489 10.6151
R1498 B.n490 B.n250 10.6151
R1499 B.n501 B.n250 10.6151
R1500 B.n502 B.n501 10.6151
R1501 B.n503 B.n502 10.6151
R1502 B.n503 B.n243 10.6151
R1503 B.n513 B.n243 10.6151
R1504 B.n514 B.n513 10.6151
R1505 B.n515 B.n514 10.6151
R1506 B.n515 B.n235 10.6151
R1507 B.n526 B.n235 10.6151
R1508 B.n527 B.n526 10.6151
R1509 B.n528 B.n527 10.6151
R1510 B.n528 B.n0 10.6151
R1511 B.n611 B.n1 10.6151
R1512 B.n611 B.n610 10.6151
R1513 B.n610 B.n609 10.6151
R1514 B.n609 B.n10 10.6151
R1515 B.n603 B.n10 10.6151
R1516 B.n603 B.n602 10.6151
R1517 B.n602 B.n601 10.6151
R1518 B.n601 B.n17 10.6151
R1519 B.n595 B.n17 10.6151
R1520 B.n595 B.n594 10.6151
R1521 B.n594 B.n593 10.6151
R1522 B.n593 B.n23 10.6151
R1523 B.n587 B.n23 10.6151
R1524 B.n587 B.n586 10.6151
R1525 B.n586 B.n585 10.6151
R1526 B.n585 B.n31 10.6151
R1527 B.n579 B.n31 10.6151
R1528 B.n579 B.n578 10.6151
R1529 B.n578 B.n577 10.6151
R1530 B.n577 B.n38 10.6151
R1531 B.n571 B.n38 10.6151
R1532 B.n571 B.n570 10.6151
R1533 B.n148 B.n89 9.36635
R1534 B.n171 B.n86 9.36635
R1535 B.n402 B.n401 9.36635
R1536 B.n380 B.n379 9.36635
R1537 B.t3 B.n241 6.27054
R1538 B.t4 B.n15 6.27054
R1539 B.n617 B.n0 2.81026
R1540 B.n617 B.n1 2.81026
R1541 B.n151 B.n89 1.24928
R1542 B.n168 B.n86 1.24928
R1543 B.n401 B.n400 1.24928
R1544 B.n381 B.n380 1.24928
R1545 VN.n2 VN.t1 289.942
R1546 VN.n10 VN.t2 289.942
R1547 VN.n6 VN.t4 272.173
R1548 VN.n14 VN.t0 272.173
R1549 VN.n1 VN.t5 229.475
R1550 VN.n9 VN.t3 229.475
R1551 VN.n7 VN.n6 161.3
R1552 VN.n15 VN.n14 161.3
R1553 VN.n13 VN.n8 161.3
R1554 VN.n12 VN.n11 161.3
R1555 VN.n5 VN.n0 161.3
R1556 VN.n4 VN.n3 161.3
R1557 VN.n5 VN.n4 52.6866
R1558 VN.n13 VN.n12 52.6866
R1559 VN.n11 VN.n10 43.4418
R1560 VN.n3 VN.n2 43.4418
R1561 VN.n2 VN.n1 42.5389
R1562 VN.n10 VN.n9 42.5389
R1563 VN VN.n15 40.0213
R1564 VN.n4 VN.n1 12.2964
R1565 VN.n12 VN.n9 12.2964
R1566 VN.n6 VN.n5 5.84292
R1567 VN.n14 VN.n13 5.84292
R1568 VN.n15 VN.n8 0.189894
R1569 VN.n11 VN.n8 0.189894
R1570 VN.n3 VN.n0 0.189894
R1571 VN.n7 VN.n0 0.189894
R1572 VN VN.n7 0.0516364
R1573 VDD2.n91 VDD2.n49 289.615
R1574 VDD2.n42 VDD2.n0 289.615
R1575 VDD2.n92 VDD2.n91 185
R1576 VDD2.n90 VDD2.n89 185
R1577 VDD2.n53 VDD2.n52 185
R1578 VDD2.n84 VDD2.n83 185
R1579 VDD2.n82 VDD2.n81 185
R1580 VDD2.n57 VDD2.n56 185
R1581 VDD2.n76 VDD2.n75 185
R1582 VDD2.n74 VDD2.n73 185
R1583 VDD2.n61 VDD2.n60 185
R1584 VDD2.n68 VDD2.n67 185
R1585 VDD2.n66 VDD2.n65 185
R1586 VDD2.n17 VDD2.n16 185
R1587 VDD2.n19 VDD2.n18 185
R1588 VDD2.n12 VDD2.n11 185
R1589 VDD2.n25 VDD2.n24 185
R1590 VDD2.n27 VDD2.n26 185
R1591 VDD2.n8 VDD2.n7 185
R1592 VDD2.n33 VDD2.n32 185
R1593 VDD2.n35 VDD2.n34 185
R1594 VDD2.n4 VDD2.n3 185
R1595 VDD2.n41 VDD2.n40 185
R1596 VDD2.n43 VDD2.n42 185
R1597 VDD2.n64 VDD2.t5 147.659
R1598 VDD2.n15 VDD2.t4 147.659
R1599 VDD2.n91 VDD2.n90 104.615
R1600 VDD2.n90 VDD2.n52 104.615
R1601 VDD2.n83 VDD2.n52 104.615
R1602 VDD2.n83 VDD2.n82 104.615
R1603 VDD2.n82 VDD2.n56 104.615
R1604 VDD2.n75 VDD2.n56 104.615
R1605 VDD2.n75 VDD2.n74 104.615
R1606 VDD2.n74 VDD2.n60 104.615
R1607 VDD2.n67 VDD2.n60 104.615
R1608 VDD2.n67 VDD2.n66 104.615
R1609 VDD2.n18 VDD2.n17 104.615
R1610 VDD2.n18 VDD2.n11 104.615
R1611 VDD2.n25 VDD2.n11 104.615
R1612 VDD2.n26 VDD2.n25 104.615
R1613 VDD2.n26 VDD2.n7 104.615
R1614 VDD2.n33 VDD2.n7 104.615
R1615 VDD2.n34 VDD2.n33 104.615
R1616 VDD2.n34 VDD2.n3 104.615
R1617 VDD2.n41 VDD2.n3 104.615
R1618 VDD2.n42 VDD2.n41 104.615
R1619 VDD2.n48 VDD2.n47 61.8248
R1620 VDD2 VDD2.n97 61.8221
R1621 VDD2.n66 VDD2.t5 52.3082
R1622 VDD2.n17 VDD2.t4 52.3082
R1623 VDD2.n48 VDD2.n46 47.2897
R1624 VDD2.n96 VDD2.n95 46.5369
R1625 VDD2.n96 VDD2.n48 34.7692
R1626 VDD2.n65 VDD2.n64 15.6677
R1627 VDD2.n16 VDD2.n15 15.6677
R1628 VDD2.n68 VDD2.n63 12.8005
R1629 VDD2.n19 VDD2.n14 12.8005
R1630 VDD2.n69 VDD2.n61 12.0247
R1631 VDD2.n20 VDD2.n12 12.0247
R1632 VDD2.n73 VDD2.n72 11.249
R1633 VDD2.n24 VDD2.n23 11.249
R1634 VDD2.n76 VDD2.n59 10.4732
R1635 VDD2.n27 VDD2.n10 10.4732
R1636 VDD2.n77 VDD2.n57 9.69747
R1637 VDD2.n28 VDD2.n8 9.69747
R1638 VDD2.n95 VDD2.n94 9.45567
R1639 VDD2.n46 VDD2.n45 9.45567
R1640 VDD2.n51 VDD2.n50 9.3005
R1641 VDD2.n94 VDD2.n93 9.3005
R1642 VDD2.n88 VDD2.n87 9.3005
R1643 VDD2.n86 VDD2.n85 9.3005
R1644 VDD2.n55 VDD2.n54 9.3005
R1645 VDD2.n80 VDD2.n79 9.3005
R1646 VDD2.n78 VDD2.n77 9.3005
R1647 VDD2.n59 VDD2.n58 9.3005
R1648 VDD2.n72 VDD2.n71 9.3005
R1649 VDD2.n70 VDD2.n69 9.3005
R1650 VDD2.n63 VDD2.n62 9.3005
R1651 VDD2.n39 VDD2.n38 9.3005
R1652 VDD2.n2 VDD2.n1 9.3005
R1653 VDD2.n45 VDD2.n44 9.3005
R1654 VDD2.n6 VDD2.n5 9.3005
R1655 VDD2.n31 VDD2.n30 9.3005
R1656 VDD2.n29 VDD2.n28 9.3005
R1657 VDD2.n10 VDD2.n9 9.3005
R1658 VDD2.n23 VDD2.n22 9.3005
R1659 VDD2.n21 VDD2.n20 9.3005
R1660 VDD2.n14 VDD2.n13 9.3005
R1661 VDD2.n37 VDD2.n36 9.3005
R1662 VDD2.n95 VDD2.n49 8.92171
R1663 VDD2.n81 VDD2.n80 8.92171
R1664 VDD2.n32 VDD2.n31 8.92171
R1665 VDD2.n46 VDD2.n0 8.92171
R1666 VDD2.n93 VDD2.n92 8.14595
R1667 VDD2.n84 VDD2.n55 8.14595
R1668 VDD2.n35 VDD2.n6 8.14595
R1669 VDD2.n44 VDD2.n43 8.14595
R1670 VDD2.n89 VDD2.n51 7.3702
R1671 VDD2.n85 VDD2.n53 7.3702
R1672 VDD2.n36 VDD2.n4 7.3702
R1673 VDD2.n40 VDD2.n2 7.3702
R1674 VDD2.n89 VDD2.n88 6.59444
R1675 VDD2.n88 VDD2.n53 6.59444
R1676 VDD2.n39 VDD2.n4 6.59444
R1677 VDD2.n40 VDD2.n39 6.59444
R1678 VDD2.n92 VDD2.n51 5.81868
R1679 VDD2.n85 VDD2.n84 5.81868
R1680 VDD2.n36 VDD2.n35 5.81868
R1681 VDD2.n43 VDD2.n2 5.81868
R1682 VDD2.n93 VDD2.n49 5.04292
R1683 VDD2.n81 VDD2.n55 5.04292
R1684 VDD2.n32 VDD2.n6 5.04292
R1685 VDD2.n44 VDD2.n0 5.04292
R1686 VDD2.n64 VDD2.n62 4.38563
R1687 VDD2.n15 VDD2.n13 4.38563
R1688 VDD2.n80 VDD2.n57 4.26717
R1689 VDD2.n31 VDD2.n8 4.26717
R1690 VDD2.n77 VDD2.n76 3.49141
R1691 VDD2.n28 VDD2.n27 3.49141
R1692 VDD2.n73 VDD2.n59 2.71565
R1693 VDD2.n24 VDD2.n10 2.71565
R1694 VDD2.n97 VDD2.t2 2.26077
R1695 VDD2.n97 VDD2.t3 2.26077
R1696 VDD2.n47 VDD2.t0 2.26077
R1697 VDD2.n47 VDD2.t1 2.26077
R1698 VDD2.n72 VDD2.n61 1.93989
R1699 VDD2.n23 VDD2.n12 1.93989
R1700 VDD2.n69 VDD2.n68 1.16414
R1701 VDD2.n20 VDD2.n19 1.16414
R1702 VDD2 VDD2.n96 0.866879
R1703 VDD2.n65 VDD2.n63 0.388379
R1704 VDD2.n16 VDD2.n14 0.388379
R1705 VDD2.n94 VDD2.n50 0.155672
R1706 VDD2.n87 VDD2.n50 0.155672
R1707 VDD2.n87 VDD2.n86 0.155672
R1708 VDD2.n86 VDD2.n54 0.155672
R1709 VDD2.n79 VDD2.n54 0.155672
R1710 VDD2.n79 VDD2.n78 0.155672
R1711 VDD2.n78 VDD2.n58 0.155672
R1712 VDD2.n71 VDD2.n58 0.155672
R1713 VDD2.n71 VDD2.n70 0.155672
R1714 VDD2.n70 VDD2.n62 0.155672
R1715 VDD2.n21 VDD2.n13 0.155672
R1716 VDD2.n22 VDD2.n21 0.155672
R1717 VDD2.n22 VDD2.n9 0.155672
R1718 VDD2.n29 VDD2.n9 0.155672
R1719 VDD2.n30 VDD2.n29 0.155672
R1720 VDD2.n30 VDD2.n5 0.155672
R1721 VDD2.n37 VDD2.n5 0.155672
R1722 VDD2.n38 VDD2.n37 0.155672
R1723 VDD2.n38 VDD2.n1 0.155672
R1724 VDD2.n45 VDD2.n1 0.155672
C0 VN VTAIL 3.55537f
C1 VTAIL VDD1 7.14815f
C2 VN VDD1 0.148755f
C3 VTAIL VP 3.56979f
C4 VN VP 4.69028f
C5 VTAIL VDD2 7.18609f
C6 VP VDD1 3.84423f
C7 VN VDD2 3.68016f
C8 VDD2 VDD1 0.790006f
C9 VP VDD2 0.316044f
C10 VDD2 B 4.090711f
C11 VDD1 B 4.114464f
C12 VTAIL B 5.376605f
C13 VN B 7.909971f
C14 VP B 6.204378f
C15 VDD2.n0 B 0.032528f
C16 VDD2.n1 B 0.022706f
C17 VDD2.n2 B 0.012201f
C18 VDD2.n3 B 0.028839f
C19 VDD2.n4 B 0.012919f
C20 VDD2.n5 B 0.022706f
C21 VDD2.n6 B 0.012201f
C22 VDD2.n7 B 0.028839f
C23 VDD2.n8 B 0.012919f
C24 VDD2.n9 B 0.022706f
C25 VDD2.n10 B 0.012201f
C26 VDD2.n11 B 0.028839f
C27 VDD2.n12 B 0.012919f
C28 VDD2.n13 B 0.827913f
C29 VDD2.n14 B 0.012201f
C30 VDD2.t4 B 0.047076f
C31 VDD2.n15 B 0.112591f
C32 VDD2.n16 B 0.017036f
C33 VDD2.n17 B 0.02163f
C34 VDD2.n18 B 0.028839f
C35 VDD2.n19 B 0.012919f
C36 VDD2.n20 B 0.012201f
C37 VDD2.n21 B 0.022706f
C38 VDD2.n22 B 0.022706f
C39 VDD2.n23 B 0.012201f
C40 VDD2.n24 B 0.012919f
C41 VDD2.n25 B 0.028839f
C42 VDD2.n26 B 0.028839f
C43 VDD2.n27 B 0.012919f
C44 VDD2.n28 B 0.012201f
C45 VDD2.n29 B 0.022706f
C46 VDD2.n30 B 0.022706f
C47 VDD2.n31 B 0.012201f
C48 VDD2.n32 B 0.012919f
C49 VDD2.n33 B 0.028839f
C50 VDD2.n34 B 0.028839f
C51 VDD2.n35 B 0.012919f
C52 VDD2.n36 B 0.012201f
C53 VDD2.n37 B 0.022706f
C54 VDD2.n38 B 0.022706f
C55 VDD2.n39 B 0.012201f
C56 VDD2.n40 B 0.012919f
C57 VDD2.n41 B 0.028839f
C58 VDD2.n42 B 0.063516f
C59 VDD2.n43 B 0.012919f
C60 VDD2.n44 B 0.012201f
C61 VDD2.n45 B 0.048762f
C62 VDD2.n46 B 0.052793f
C63 VDD2.t0 B 0.157181f
C64 VDD2.t1 B 0.157181f
C65 VDD2.n47 B 1.36222f
C66 VDD2.n48 B 1.59561f
C67 VDD2.n49 B 0.032528f
C68 VDD2.n50 B 0.022706f
C69 VDD2.n51 B 0.012201f
C70 VDD2.n52 B 0.028839f
C71 VDD2.n53 B 0.012919f
C72 VDD2.n54 B 0.022706f
C73 VDD2.n55 B 0.012201f
C74 VDD2.n56 B 0.028839f
C75 VDD2.n57 B 0.012919f
C76 VDD2.n58 B 0.022706f
C77 VDD2.n59 B 0.012201f
C78 VDD2.n60 B 0.028839f
C79 VDD2.n61 B 0.012919f
C80 VDD2.n62 B 0.827913f
C81 VDD2.n63 B 0.012201f
C82 VDD2.t5 B 0.047076f
C83 VDD2.n64 B 0.112591f
C84 VDD2.n65 B 0.017036f
C85 VDD2.n66 B 0.02163f
C86 VDD2.n67 B 0.028839f
C87 VDD2.n68 B 0.012919f
C88 VDD2.n69 B 0.012201f
C89 VDD2.n70 B 0.022706f
C90 VDD2.n71 B 0.022706f
C91 VDD2.n72 B 0.012201f
C92 VDD2.n73 B 0.012919f
C93 VDD2.n74 B 0.028839f
C94 VDD2.n75 B 0.028839f
C95 VDD2.n76 B 0.012919f
C96 VDD2.n77 B 0.012201f
C97 VDD2.n78 B 0.022706f
C98 VDD2.n79 B 0.022706f
C99 VDD2.n80 B 0.012201f
C100 VDD2.n81 B 0.012919f
C101 VDD2.n82 B 0.028839f
C102 VDD2.n83 B 0.028839f
C103 VDD2.n84 B 0.012919f
C104 VDD2.n85 B 0.012201f
C105 VDD2.n86 B 0.022706f
C106 VDD2.n87 B 0.022706f
C107 VDD2.n88 B 0.012201f
C108 VDD2.n89 B 0.012919f
C109 VDD2.n90 B 0.028839f
C110 VDD2.n91 B 0.063516f
C111 VDD2.n92 B 0.012919f
C112 VDD2.n93 B 0.012201f
C113 VDD2.n94 B 0.048762f
C114 VDD2.n95 B 0.051243f
C115 VDD2.n96 B 1.67702f
C116 VDD2.t2 B 0.157181f
C117 VDD2.t3 B 0.157181f
C118 VDD2.n97 B 1.3622f
C119 VN.n0 B 0.04206f
C120 VN.t5 B 0.913813f
C121 VN.n1 B 0.395108f
C122 VN.t1 B 0.998043f
C123 VN.n2 B 0.40673f
C124 VN.n3 B 0.178248f
C125 VN.n4 B 0.055459f
C126 VN.n5 B 0.014189f
C127 VN.t4 B 0.972733f
C128 VN.n6 B 0.401456f
C129 VN.n7 B 0.032595f
C130 VN.n8 B 0.04206f
C131 VN.t3 B 0.913813f
C132 VN.n9 B 0.395108f
C133 VN.t2 B 0.998043f
C134 VN.n10 B 0.40673f
C135 VN.n11 B 0.178248f
C136 VN.n12 B 0.055459f
C137 VN.n13 B 0.014189f
C138 VN.t0 B 0.972733f
C139 VN.n14 B 0.401456f
C140 VN.n15 B 1.60119f
C141 VDD1.n0 B 0.03228f
C142 VDD1.n1 B 0.022533f
C143 VDD1.n2 B 0.012108f
C144 VDD1.n3 B 0.028619f
C145 VDD1.n4 B 0.01282f
C146 VDD1.n5 B 0.022533f
C147 VDD1.n6 B 0.012108f
C148 VDD1.n7 B 0.028619f
C149 VDD1.n8 B 0.01282f
C150 VDD1.n9 B 0.022533f
C151 VDD1.n10 B 0.012108f
C152 VDD1.n11 B 0.028619f
C153 VDD1.n12 B 0.01282f
C154 VDD1.n13 B 0.821591f
C155 VDD1.n14 B 0.012108f
C156 VDD1.t5 B 0.046717f
C157 VDD1.n15 B 0.111731f
C158 VDD1.n16 B 0.016906f
C159 VDD1.n17 B 0.021464f
C160 VDD1.n18 B 0.028619f
C161 VDD1.n19 B 0.01282f
C162 VDD1.n20 B 0.012108f
C163 VDD1.n21 B 0.022533f
C164 VDD1.n22 B 0.022533f
C165 VDD1.n23 B 0.012108f
C166 VDD1.n24 B 0.01282f
C167 VDD1.n25 B 0.028619f
C168 VDD1.n26 B 0.028619f
C169 VDD1.n27 B 0.01282f
C170 VDD1.n28 B 0.012108f
C171 VDD1.n29 B 0.022533f
C172 VDD1.n30 B 0.022533f
C173 VDD1.n31 B 0.012108f
C174 VDD1.n32 B 0.01282f
C175 VDD1.n33 B 0.028619f
C176 VDD1.n34 B 0.028619f
C177 VDD1.n35 B 0.01282f
C178 VDD1.n36 B 0.012108f
C179 VDD1.n37 B 0.022533f
C180 VDD1.n38 B 0.022533f
C181 VDD1.n39 B 0.012108f
C182 VDD1.n40 B 0.01282f
C183 VDD1.n41 B 0.028619f
C184 VDD1.n42 B 0.063031f
C185 VDD1.n43 B 0.01282f
C186 VDD1.n44 B 0.012108f
C187 VDD1.n45 B 0.04839f
C188 VDD1.n46 B 0.052756f
C189 VDD1.n47 B 0.03228f
C190 VDD1.n48 B 0.022533f
C191 VDD1.n49 B 0.012108f
C192 VDD1.n50 B 0.028619f
C193 VDD1.n51 B 0.01282f
C194 VDD1.n52 B 0.022533f
C195 VDD1.n53 B 0.012108f
C196 VDD1.n54 B 0.028619f
C197 VDD1.n55 B 0.01282f
C198 VDD1.n56 B 0.022533f
C199 VDD1.n57 B 0.012108f
C200 VDD1.n58 B 0.028619f
C201 VDD1.n59 B 0.01282f
C202 VDD1.n60 B 0.821591f
C203 VDD1.n61 B 0.012108f
C204 VDD1.t3 B 0.046717f
C205 VDD1.n62 B 0.111731f
C206 VDD1.n63 B 0.016906f
C207 VDD1.n64 B 0.021464f
C208 VDD1.n65 B 0.028619f
C209 VDD1.n66 B 0.01282f
C210 VDD1.n67 B 0.012108f
C211 VDD1.n68 B 0.022533f
C212 VDD1.n69 B 0.022533f
C213 VDD1.n70 B 0.012108f
C214 VDD1.n71 B 0.01282f
C215 VDD1.n72 B 0.028619f
C216 VDD1.n73 B 0.028619f
C217 VDD1.n74 B 0.01282f
C218 VDD1.n75 B 0.012108f
C219 VDD1.n76 B 0.022533f
C220 VDD1.n77 B 0.022533f
C221 VDD1.n78 B 0.012108f
C222 VDD1.n79 B 0.01282f
C223 VDD1.n80 B 0.028619f
C224 VDD1.n81 B 0.028619f
C225 VDD1.n82 B 0.01282f
C226 VDD1.n83 B 0.012108f
C227 VDD1.n84 B 0.022533f
C228 VDD1.n85 B 0.022533f
C229 VDD1.n86 B 0.012108f
C230 VDD1.n87 B 0.01282f
C231 VDD1.n88 B 0.028619f
C232 VDD1.n89 B 0.063031f
C233 VDD1.n90 B 0.01282f
C234 VDD1.n91 B 0.012108f
C235 VDD1.n92 B 0.04839f
C236 VDD1.n93 B 0.05239f
C237 VDD1.t2 B 0.155981f
C238 VDD1.t0 B 0.155981f
C239 VDD1.n94 B 1.35181f
C240 VDD1.n95 B 1.65628f
C241 VDD1.t4 B 0.155981f
C242 VDD1.t1 B 0.155981f
C243 VDD1.n96 B 1.3508f
C244 VDD1.n97 B 1.86379f
C245 VTAIL.t0 B 0.169012f
C246 VTAIL.t4 B 0.169012f
C247 VTAIL.n0 B 1.38864f
C248 VTAIL.n1 B 0.353588f
C249 VTAIL.n2 B 0.034977f
C250 VTAIL.n3 B 0.024415f
C251 VTAIL.n4 B 0.01312f
C252 VTAIL.n5 B 0.03101f
C253 VTAIL.n6 B 0.013891f
C254 VTAIL.n7 B 0.024415f
C255 VTAIL.n8 B 0.01312f
C256 VTAIL.n9 B 0.03101f
C257 VTAIL.n10 B 0.013891f
C258 VTAIL.n11 B 0.024415f
C259 VTAIL.n12 B 0.01312f
C260 VTAIL.n13 B 0.03101f
C261 VTAIL.n14 B 0.013891f
C262 VTAIL.n15 B 0.890226f
C263 VTAIL.n16 B 0.01312f
C264 VTAIL.t5 B 0.05062f
C265 VTAIL.n17 B 0.121065f
C266 VTAIL.n18 B 0.018319f
C267 VTAIL.n19 B 0.023257f
C268 VTAIL.n20 B 0.03101f
C269 VTAIL.n21 B 0.013891f
C270 VTAIL.n22 B 0.01312f
C271 VTAIL.n23 B 0.024415f
C272 VTAIL.n24 B 0.024415f
C273 VTAIL.n25 B 0.01312f
C274 VTAIL.n26 B 0.013891f
C275 VTAIL.n27 B 0.03101f
C276 VTAIL.n28 B 0.03101f
C277 VTAIL.n29 B 0.013891f
C278 VTAIL.n30 B 0.01312f
C279 VTAIL.n31 B 0.024415f
C280 VTAIL.n32 B 0.024415f
C281 VTAIL.n33 B 0.01312f
C282 VTAIL.n34 B 0.013891f
C283 VTAIL.n35 B 0.03101f
C284 VTAIL.n36 B 0.03101f
C285 VTAIL.n37 B 0.013891f
C286 VTAIL.n38 B 0.01312f
C287 VTAIL.n39 B 0.024415f
C288 VTAIL.n40 B 0.024415f
C289 VTAIL.n41 B 0.01312f
C290 VTAIL.n42 B 0.013891f
C291 VTAIL.n43 B 0.03101f
C292 VTAIL.n44 B 0.068297f
C293 VTAIL.n45 B 0.013891f
C294 VTAIL.n46 B 0.01312f
C295 VTAIL.n47 B 0.052432f
C296 VTAIL.n48 B 0.038207f
C297 VTAIL.n49 B 0.182722f
C298 VTAIL.t9 B 0.169012f
C299 VTAIL.t6 B 0.169012f
C300 VTAIL.n50 B 1.38864f
C301 VTAIL.n51 B 1.42854f
C302 VTAIL.t1 B 0.169012f
C303 VTAIL.t3 B 0.169012f
C304 VTAIL.n52 B 1.38865f
C305 VTAIL.n53 B 1.42853f
C306 VTAIL.n54 B 0.034977f
C307 VTAIL.n55 B 0.024415f
C308 VTAIL.n56 B 0.01312f
C309 VTAIL.n57 B 0.03101f
C310 VTAIL.n58 B 0.013891f
C311 VTAIL.n59 B 0.024415f
C312 VTAIL.n60 B 0.01312f
C313 VTAIL.n61 B 0.03101f
C314 VTAIL.n62 B 0.013891f
C315 VTAIL.n63 B 0.024415f
C316 VTAIL.n64 B 0.01312f
C317 VTAIL.n65 B 0.03101f
C318 VTAIL.n66 B 0.013891f
C319 VTAIL.n67 B 0.890226f
C320 VTAIL.n68 B 0.01312f
C321 VTAIL.t2 B 0.05062f
C322 VTAIL.n69 B 0.121065f
C323 VTAIL.n70 B 0.018319f
C324 VTAIL.n71 B 0.023257f
C325 VTAIL.n72 B 0.03101f
C326 VTAIL.n73 B 0.013891f
C327 VTAIL.n74 B 0.01312f
C328 VTAIL.n75 B 0.024415f
C329 VTAIL.n76 B 0.024415f
C330 VTAIL.n77 B 0.01312f
C331 VTAIL.n78 B 0.013891f
C332 VTAIL.n79 B 0.03101f
C333 VTAIL.n80 B 0.03101f
C334 VTAIL.n81 B 0.013891f
C335 VTAIL.n82 B 0.01312f
C336 VTAIL.n83 B 0.024415f
C337 VTAIL.n84 B 0.024415f
C338 VTAIL.n85 B 0.01312f
C339 VTAIL.n86 B 0.013891f
C340 VTAIL.n87 B 0.03101f
C341 VTAIL.n88 B 0.03101f
C342 VTAIL.n89 B 0.013891f
C343 VTAIL.n90 B 0.01312f
C344 VTAIL.n91 B 0.024415f
C345 VTAIL.n92 B 0.024415f
C346 VTAIL.n93 B 0.01312f
C347 VTAIL.n94 B 0.013891f
C348 VTAIL.n95 B 0.03101f
C349 VTAIL.n96 B 0.068297f
C350 VTAIL.n97 B 0.013891f
C351 VTAIL.n98 B 0.01312f
C352 VTAIL.n99 B 0.052432f
C353 VTAIL.n100 B 0.038207f
C354 VTAIL.n101 B 0.182722f
C355 VTAIL.t8 B 0.169012f
C356 VTAIL.t7 B 0.169012f
C357 VTAIL.n102 B 1.38865f
C358 VTAIL.n103 B 0.412582f
C359 VTAIL.n104 B 0.034977f
C360 VTAIL.n105 B 0.024415f
C361 VTAIL.n106 B 0.01312f
C362 VTAIL.n107 B 0.03101f
C363 VTAIL.n108 B 0.013891f
C364 VTAIL.n109 B 0.024415f
C365 VTAIL.n110 B 0.01312f
C366 VTAIL.n111 B 0.03101f
C367 VTAIL.n112 B 0.013891f
C368 VTAIL.n113 B 0.024415f
C369 VTAIL.n114 B 0.01312f
C370 VTAIL.n115 B 0.03101f
C371 VTAIL.n116 B 0.013891f
C372 VTAIL.n117 B 0.890226f
C373 VTAIL.n118 B 0.01312f
C374 VTAIL.t10 B 0.05062f
C375 VTAIL.n119 B 0.121065f
C376 VTAIL.n120 B 0.018319f
C377 VTAIL.n121 B 0.023257f
C378 VTAIL.n122 B 0.03101f
C379 VTAIL.n123 B 0.013891f
C380 VTAIL.n124 B 0.01312f
C381 VTAIL.n125 B 0.024415f
C382 VTAIL.n126 B 0.024415f
C383 VTAIL.n127 B 0.01312f
C384 VTAIL.n128 B 0.013891f
C385 VTAIL.n129 B 0.03101f
C386 VTAIL.n130 B 0.03101f
C387 VTAIL.n131 B 0.013891f
C388 VTAIL.n132 B 0.01312f
C389 VTAIL.n133 B 0.024415f
C390 VTAIL.n134 B 0.024415f
C391 VTAIL.n135 B 0.01312f
C392 VTAIL.n136 B 0.013891f
C393 VTAIL.n137 B 0.03101f
C394 VTAIL.n138 B 0.03101f
C395 VTAIL.n139 B 0.013891f
C396 VTAIL.n140 B 0.01312f
C397 VTAIL.n141 B 0.024415f
C398 VTAIL.n142 B 0.024415f
C399 VTAIL.n143 B 0.01312f
C400 VTAIL.n144 B 0.013891f
C401 VTAIL.n145 B 0.03101f
C402 VTAIL.n146 B 0.068297f
C403 VTAIL.n147 B 0.013891f
C404 VTAIL.n148 B 0.01312f
C405 VTAIL.n149 B 0.052432f
C406 VTAIL.n150 B 0.038207f
C407 VTAIL.n151 B 1.1139f
C408 VTAIL.n152 B 0.034977f
C409 VTAIL.n153 B 0.024415f
C410 VTAIL.n154 B 0.01312f
C411 VTAIL.n155 B 0.03101f
C412 VTAIL.n156 B 0.013891f
C413 VTAIL.n157 B 0.024415f
C414 VTAIL.n158 B 0.01312f
C415 VTAIL.n159 B 0.03101f
C416 VTAIL.n160 B 0.013891f
C417 VTAIL.n161 B 0.024415f
C418 VTAIL.n162 B 0.01312f
C419 VTAIL.n163 B 0.03101f
C420 VTAIL.n164 B 0.013891f
C421 VTAIL.n165 B 0.890226f
C422 VTAIL.n166 B 0.01312f
C423 VTAIL.t11 B 0.05062f
C424 VTAIL.n167 B 0.121065f
C425 VTAIL.n168 B 0.018319f
C426 VTAIL.n169 B 0.023257f
C427 VTAIL.n170 B 0.03101f
C428 VTAIL.n171 B 0.013891f
C429 VTAIL.n172 B 0.01312f
C430 VTAIL.n173 B 0.024415f
C431 VTAIL.n174 B 0.024415f
C432 VTAIL.n175 B 0.01312f
C433 VTAIL.n176 B 0.013891f
C434 VTAIL.n177 B 0.03101f
C435 VTAIL.n178 B 0.03101f
C436 VTAIL.n179 B 0.013891f
C437 VTAIL.n180 B 0.01312f
C438 VTAIL.n181 B 0.024415f
C439 VTAIL.n182 B 0.024415f
C440 VTAIL.n183 B 0.01312f
C441 VTAIL.n184 B 0.013891f
C442 VTAIL.n185 B 0.03101f
C443 VTAIL.n186 B 0.03101f
C444 VTAIL.n187 B 0.013891f
C445 VTAIL.n188 B 0.01312f
C446 VTAIL.n189 B 0.024415f
C447 VTAIL.n190 B 0.024415f
C448 VTAIL.n191 B 0.01312f
C449 VTAIL.n192 B 0.013891f
C450 VTAIL.n193 B 0.03101f
C451 VTAIL.n194 B 0.068297f
C452 VTAIL.n195 B 0.013891f
C453 VTAIL.n196 B 0.01312f
C454 VTAIL.n197 B 0.052432f
C455 VTAIL.n198 B 0.038207f
C456 VTAIL.n199 B 1.08813f
C457 VP.n0 B 0.042621f
C458 VP.t3 B 0.92599f
C459 VP.n1 B 0.359891f
C460 VP.n2 B 0.042621f
C461 VP.n3 B 0.042621f
C462 VP.t4 B 0.985696f
C463 VP.t1 B 0.92599f
C464 VP.n4 B 0.400373f
C465 VP.t0 B 1.01134f
C466 VP.n5 B 0.41215f
C467 VP.n6 B 0.180623f
C468 VP.n7 B 0.056198f
C469 VP.n8 B 0.014378f
C470 VP.n9 B 0.406805f
C471 VP.n10 B 1.59444f
C472 VP.n11 B 1.6332f
C473 VP.t2 B 0.985696f
C474 VP.n12 B 0.406805f
C475 VP.n13 B 0.014378f
C476 VP.n14 B 0.056198f
C477 VP.n15 B 0.042621f
C478 VP.n16 B 0.042621f
C479 VP.n17 B 0.056198f
C480 VP.n18 B 0.014378f
C481 VP.t5 B 0.985696f
C482 VP.n19 B 0.406805f
C483 VP.n20 B 0.03303f
.ends

