* NGSPICE file created from diff_pair_sample_0463.ext - technology: sky130A

.subckt diff_pair_sample_0463 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t14 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=7.2774 pd=38.1 as=3.0789 ps=18.99 w=18.66 l=3.25
X1 B.t11 B.t9 B.t10 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=7.2774 pd=38.1 as=0 ps=0 w=18.66 l=3.25
X2 VDD2.t9 VN.t0 VTAIL.t7 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=7.2774 pd=38.1 as=3.0789 ps=18.99 w=18.66 l=3.25
X3 VTAIL.t19 VP.t1 VDD1.t8 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
X4 VTAIL.t9 VN.t1 VDD2.t8 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
X5 VDD1.t7 VP.t2 VTAIL.t13 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=7.2774 pd=38.1 as=3.0789 ps=18.99 w=18.66 l=3.25
X6 VDD1.t6 VP.t3 VTAIL.t10 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=7.2774 ps=38.1 w=18.66 l=3.25
X7 VTAIL.t18 VP.t4 VDD1.t5 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
X8 B.t8 B.t6 B.t7 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=7.2774 pd=38.1 as=0 ps=0 w=18.66 l=3.25
X9 VTAIL.t6 VN.t2 VDD2.t7 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
X10 VDD2.t6 VN.t3 VTAIL.t8 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=7.2774 ps=38.1 w=18.66 l=3.25
X11 VDD2.t5 VN.t4 VTAIL.t5 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
X12 VTAIL.t4 VN.t5 VDD2.t4 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
X13 VTAIL.t16 VP.t5 VDD1.t4 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
X14 VDD1.t3 VP.t6 VTAIL.t17 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
X15 VDD1.t2 VP.t7 VTAIL.t11 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
X16 VTAIL.t15 VP.t8 VDD1.t1 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
X17 VDD2.t3 VN.t6 VTAIL.t3 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=7.2774 ps=38.1 w=18.66 l=3.25
X18 B.t5 B.t3 B.t4 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=7.2774 pd=38.1 as=0 ps=0 w=18.66 l=3.25
X19 VDD1.t0 VP.t9 VTAIL.t12 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=7.2774 ps=38.1 w=18.66 l=3.25
X20 VTAIL.t2 VN.t7 VDD2.t2 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
X21 VDD2.t1 VN.t8 VTAIL.t1 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=7.2774 pd=38.1 as=3.0789 ps=18.99 w=18.66 l=3.25
X22 B.t2 B.t0 B.t1 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=7.2774 pd=38.1 as=0 ps=0 w=18.66 l=3.25
X23 VDD2.t0 VN.t9 VTAIL.t0 w_n5266_n4700# sky130_fd_pr__pfet_01v8 ad=3.0789 pd=18.99 as=3.0789 ps=18.99 w=18.66 l=3.25
R0 VP.n30 VP.t2 171.821
R1 VP.n32 VP.n31 161.3
R2 VP.n33 VP.n28 161.3
R3 VP.n35 VP.n34 161.3
R4 VP.n36 VP.n27 161.3
R5 VP.n38 VP.n37 161.3
R6 VP.n39 VP.n26 161.3
R7 VP.n41 VP.n40 161.3
R8 VP.n43 VP.n42 161.3
R9 VP.n44 VP.n24 161.3
R10 VP.n46 VP.n45 161.3
R11 VP.n47 VP.n23 161.3
R12 VP.n49 VP.n48 161.3
R13 VP.n50 VP.n22 161.3
R14 VP.n52 VP.n51 161.3
R15 VP.n54 VP.n53 161.3
R16 VP.n55 VP.n20 161.3
R17 VP.n57 VP.n56 161.3
R18 VP.n58 VP.n19 161.3
R19 VP.n60 VP.n59 161.3
R20 VP.n61 VP.n18 161.3
R21 VP.n63 VP.n62 161.3
R22 VP.n109 VP.n108 161.3
R23 VP.n107 VP.n1 161.3
R24 VP.n106 VP.n105 161.3
R25 VP.n104 VP.n2 161.3
R26 VP.n103 VP.n102 161.3
R27 VP.n101 VP.n3 161.3
R28 VP.n100 VP.n99 161.3
R29 VP.n98 VP.n97 161.3
R30 VP.n96 VP.n5 161.3
R31 VP.n95 VP.n94 161.3
R32 VP.n93 VP.n6 161.3
R33 VP.n92 VP.n91 161.3
R34 VP.n90 VP.n7 161.3
R35 VP.n89 VP.n88 161.3
R36 VP.n87 VP.n86 161.3
R37 VP.n85 VP.n9 161.3
R38 VP.n84 VP.n83 161.3
R39 VP.n82 VP.n10 161.3
R40 VP.n81 VP.n80 161.3
R41 VP.n79 VP.n11 161.3
R42 VP.n78 VP.n77 161.3
R43 VP.n76 VP.n75 161.3
R44 VP.n74 VP.n13 161.3
R45 VP.n73 VP.n72 161.3
R46 VP.n71 VP.n14 161.3
R47 VP.n70 VP.n69 161.3
R48 VP.n68 VP.n15 161.3
R49 VP.n67 VP.n66 161.3
R50 VP.n16 VP.t0 138.371
R51 VP.n12 VP.t5 138.371
R52 VP.n8 VP.t6 138.371
R53 VP.n4 VP.t8 138.371
R54 VP.n0 VP.t3 138.371
R55 VP.n17 VP.t9 138.371
R56 VP.n21 VP.t4 138.371
R57 VP.n25 VP.t7 138.371
R58 VP.n29 VP.t1 138.371
R59 VP.n65 VP.n16 70.0803
R60 VP.n110 VP.n0 70.0803
R61 VP.n64 VP.n17 70.0803
R62 VP.n65 VP.n64 61.8783
R63 VP.n30 VP.n29 58.1016
R64 VP.n69 VP.n14 52.2023
R65 VP.n106 VP.n2 52.2023
R66 VP.n60 VP.n19 52.2023
R67 VP.n80 VP.n10 44.4521
R68 VP.n95 VP.n6 44.4521
R69 VP.n49 VP.n23 44.4521
R70 VP.n34 VP.n27 44.4521
R71 VP.n84 VP.n10 36.702
R72 VP.n91 VP.n6 36.702
R73 VP.n45 VP.n23 36.702
R74 VP.n38 VP.n27 36.702
R75 VP.n73 VP.n14 28.9518
R76 VP.n102 VP.n2 28.9518
R77 VP.n56 VP.n19 28.9518
R78 VP.n68 VP.n67 24.5923
R79 VP.n69 VP.n68 24.5923
R80 VP.n74 VP.n73 24.5923
R81 VP.n75 VP.n74 24.5923
R82 VP.n79 VP.n78 24.5923
R83 VP.n80 VP.n79 24.5923
R84 VP.n85 VP.n84 24.5923
R85 VP.n86 VP.n85 24.5923
R86 VP.n90 VP.n89 24.5923
R87 VP.n91 VP.n90 24.5923
R88 VP.n96 VP.n95 24.5923
R89 VP.n97 VP.n96 24.5923
R90 VP.n101 VP.n100 24.5923
R91 VP.n102 VP.n101 24.5923
R92 VP.n107 VP.n106 24.5923
R93 VP.n108 VP.n107 24.5923
R94 VP.n61 VP.n60 24.5923
R95 VP.n62 VP.n61 24.5923
R96 VP.n50 VP.n49 24.5923
R97 VP.n51 VP.n50 24.5923
R98 VP.n55 VP.n54 24.5923
R99 VP.n56 VP.n55 24.5923
R100 VP.n39 VP.n38 24.5923
R101 VP.n40 VP.n39 24.5923
R102 VP.n44 VP.n43 24.5923
R103 VP.n45 VP.n44 24.5923
R104 VP.n33 VP.n32 24.5923
R105 VP.n34 VP.n33 24.5923
R106 VP.n67 VP.n16 20.1658
R107 VP.n108 VP.n0 20.1658
R108 VP.n62 VP.n17 20.1658
R109 VP.n78 VP.n12 16.2311
R110 VP.n97 VP.n4 16.2311
R111 VP.n51 VP.n21 16.2311
R112 VP.n32 VP.n29 16.2311
R113 VP.n86 VP.n8 12.2964
R114 VP.n89 VP.n8 12.2964
R115 VP.n40 VP.n25 12.2964
R116 VP.n43 VP.n25 12.2964
R117 VP.n75 VP.n12 8.36172
R118 VP.n100 VP.n4 8.36172
R119 VP.n54 VP.n21 8.36172
R120 VP.n31 VP.n30 3.88974
R121 VP.n64 VP.n63 0.354861
R122 VP.n66 VP.n65 0.354861
R123 VP.n110 VP.n109 0.354861
R124 VP VP.n110 0.267071
R125 VP.n31 VP.n28 0.189894
R126 VP.n35 VP.n28 0.189894
R127 VP.n36 VP.n35 0.189894
R128 VP.n37 VP.n36 0.189894
R129 VP.n37 VP.n26 0.189894
R130 VP.n41 VP.n26 0.189894
R131 VP.n42 VP.n41 0.189894
R132 VP.n42 VP.n24 0.189894
R133 VP.n46 VP.n24 0.189894
R134 VP.n47 VP.n46 0.189894
R135 VP.n48 VP.n47 0.189894
R136 VP.n48 VP.n22 0.189894
R137 VP.n52 VP.n22 0.189894
R138 VP.n53 VP.n52 0.189894
R139 VP.n53 VP.n20 0.189894
R140 VP.n57 VP.n20 0.189894
R141 VP.n58 VP.n57 0.189894
R142 VP.n59 VP.n58 0.189894
R143 VP.n59 VP.n18 0.189894
R144 VP.n63 VP.n18 0.189894
R145 VP.n66 VP.n15 0.189894
R146 VP.n70 VP.n15 0.189894
R147 VP.n71 VP.n70 0.189894
R148 VP.n72 VP.n71 0.189894
R149 VP.n72 VP.n13 0.189894
R150 VP.n76 VP.n13 0.189894
R151 VP.n77 VP.n76 0.189894
R152 VP.n77 VP.n11 0.189894
R153 VP.n81 VP.n11 0.189894
R154 VP.n82 VP.n81 0.189894
R155 VP.n83 VP.n82 0.189894
R156 VP.n83 VP.n9 0.189894
R157 VP.n87 VP.n9 0.189894
R158 VP.n88 VP.n87 0.189894
R159 VP.n88 VP.n7 0.189894
R160 VP.n92 VP.n7 0.189894
R161 VP.n93 VP.n92 0.189894
R162 VP.n94 VP.n93 0.189894
R163 VP.n94 VP.n5 0.189894
R164 VP.n98 VP.n5 0.189894
R165 VP.n99 VP.n98 0.189894
R166 VP.n99 VP.n3 0.189894
R167 VP.n103 VP.n3 0.189894
R168 VP.n104 VP.n103 0.189894
R169 VP.n105 VP.n104 0.189894
R170 VP.n105 VP.n1 0.189894
R171 VP.n109 VP.n1 0.189894
R172 VTAIL.n11 VTAIL.t8 54.7593
R173 VTAIL.n17 VTAIL.t3 54.7591
R174 VTAIL.n2 VTAIL.t10 54.7591
R175 VTAIL.n16 VTAIL.t12 54.7591
R176 VTAIL.n15 VTAIL.n14 53.0174
R177 VTAIL.n13 VTAIL.n12 53.0174
R178 VTAIL.n10 VTAIL.n9 53.0174
R179 VTAIL.n8 VTAIL.n7 53.0174
R180 VTAIL.n19 VTAIL.n18 53.0171
R181 VTAIL.n1 VTAIL.n0 53.0171
R182 VTAIL.n4 VTAIL.n3 53.0171
R183 VTAIL.n6 VTAIL.n5 53.0171
R184 VTAIL.n8 VTAIL.n6 34.6255
R185 VTAIL.n17 VTAIL.n16 31.5393
R186 VTAIL.n10 VTAIL.n8 3.08671
R187 VTAIL.n11 VTAIL.n10 3.08671
R188 VTAIL.n15 VTAIL.n13 3.08671
R189 VTAIL.n16 VTAIL.n15 3.08671
R190 VTAIL.n6 VTAIL.n4 3.08671
R191 VTAIL.n4 VTAIL.n2 3.08671
R192 VTAIL.n19 VTAIL.n17 3.08671
R193 VTAIL VTAIL.n1 2.37334
R194 VTAIL.n13 VTAIL.n11 2.01343
R195 VTAIL.n2 VTAIL.n1 2.01343
R196 VTAIL.n18 VTAIL.t5 1.74246
R197 VTAIL.n18 VTAIL.t2 1.74246
R198 VTAIL.n0 VTAIL.t1 1.74246
R199 VTAIL.n0 VTAIL.t4 1.74246
R200 VTAIL.n3 VTAIL.t17 1.74246
R201 VTAIL.n3 VTAIL.t15 1.74246
R202 VTAIL.n5 VTAIL.t14 1.74246
R203 VTAIL.n5 VTAIL.t16 1.74246
R204 VTAIL.n14 VTAIL.t11 1.74246
R205 VTAIL.n14 VTAIL.t18 1.74246
R206 VTAIL.n12 VTAIL.t13 1.74246
R207 VTAIL.n12 VTAIL.t19 1.74246
R208 VTAIL.n9 VTAIL.t0 1.74246
R209 VTAIL.n9 VTAIL.t9 1.74246
R210 VTAIL.n7 VTAIL.t7 1.74246
R211 VTAIL.n7 VTAIL.t6 1.74246
R212 VTAIL VTAIL.n19 0.713862
R213 VDD1.n1 VDD1.t7 74.5243
R214 VDD1.n3 VDD1.t9 74.5241
R215 VDD1.n5 VDD1.n4 71.9552
R216 VDD1.n1 VDD1.n0 69.6962
R217 VDD1.n7 VDD1.n6 69.696
R218 VDD1.n3 VDD1.n2 69.6959
R219 VDD1.n7 VDD1.n5 56.5871
R220 VDD1 VDD1.n7 2.25697
R221 VDD1.n6 VDD1.t5 1.74246
R222 VDD1.n6 VDD1.t0 1.74246
R223 VDD1.n0 VDD1.t8 1.74246
R224 VDD1.n0 VDD1.t2 1.74246
R225 VDD1.n4 VDD1.t1 1.74246
R226 VDD1.n4 VDD1.t6 1.74246
R227 VDD1.n2 VDD1.t4 1.74246
R228 VDD1.n2 VDD1.t3 1.74246
R229 VDD1 VDD1.n1 0.830241
R230 VDD1.n5 VDD1.n3 0.716706
R231 B.n805 B.n804 585
R232 B.n806 B.n107 585
R233 B.n808 B.n807 585
R234 B.n809 B.n106 585
R235 B.n811 B.n810 585
R236 B.n812 B.n105 585
R237 B.n814 B.n813 585
R238 B.n815 B.n104 585
R239 B.n817 B.n816 585
R240 B.n818 B.n103 585
R241 B.n820 B.n819 585
R242 B.n821 B.n102 585
R243 B.n823 B.n822 585
R244 B.n824 B.n101 585
R245 B.n826 B.n825 585
R246 B.n827 B.n100 585
R247 B.n829 B.n828 585
R248 B.n830 B.n99 585
R249 B.n832 B.n831 585
R250 B.n833 B.n98 585
R251 B.n835 B.n834 585
R252 B.n836 B.n97 585
R253 B.n838 B.n837 585
R254 B.n839 B.n96 585
R255 B.n841 B.n840 585
R256 B.n842 B.n95 585
R257 B.n844 B.n843 585
R258 B.n845 B.n94 585
R259 B.n847 B.n846 585
R260 B.n848 B.n93 585
R261 B.n850 B.n849 585
R262 B.n851 B.n92 585
R263 B.n853 B.n852 585
R264 B.n854 B.n91 585
R265 B.n856 B.n855 585
R266 B.n857 B.n90 585
R267 B.n859 B.n858 585
R268 B.n860 B.n89 585
R269 B.n862 B.n861 585
R270 B.n863 B.n88 585
R271 B.n865 B.n864 585
R272 B.n866 B.n87 585
R273 B.n868 B.n867 585
R274 B.n869 B.n86 585
R275 B.n871 B.n870 585
R276 B.n872 B.n85 585
R277 B.n874 B.n873 585
R278 B.n875 B.n84 585
R279 B.n877 B.n876 585
R280 B.n878 B.n83 585
R281 B.n880 B.n879 585
R282 B.n881 B.n82 585
R283 B.n883 B.n882 585
R284 B.n884 B.n81 585
R285 B.n886 B.n885 585
R286 B.n887 B.n80 585
R287 B.n889 B.n888 585
R288 B.n890 B.n79 585
R289 B.n892 B.n891 585
R290 B.n893 B.n78 585
R291 B.n895 B.n894 585
R292 B.n897 B.n75 585
R293 B.n899 B.n898 585
R294 B.n900 B.n74 585
R295 B.n902 B.n901 585
R296 B.n903 B.n73 585
R297 B.n905 B.n904 585
R298 B.n906 B.n72 585
R299 B.n908 B.n907 585
R300 B.n909 B.n71 585
R301 B.n911 B.n910 585
R302 B.n913 B.n912 585
R303 B.n914 B.n67 585
R304 B.n916 B.n915 585
R305 B.n917 B.n66 585
R306 B.n919 B.n918 585
R307 B.n920 B.n65 585
R308 B.n922 B.n921 585
R309 B.n923 B.n64 585
R310 B.n925 B.n924 585
R311 B.n926 B.n63 585
R312 B.n928 B.n927 585
R313 B.n929 B.n62 585
R314 B.n931 B.n930 585
R315 B.n932 B.n61 585
R316 B.n934 B.n933 585
R317 B.n935 B.n60 585
R318 B.n937 B.n936 585
R319 B.n938 B.n59 585
R320 B.n940 B.n939 585
R321 B.n941 B.n58 585
R322 B.n943 B.n942 585
R323 B.n944 B.n57 585
R324 B.n946 B.n945 585
R325 B.n947 B.n56 585
R326 B.n949 B.n948 585
R327 B.n950 B.n55 585
R328 B.n952 B.n951 585
R329 B.n953 B.n54 585
R330 B.n955 B.n954 585
R331 B.n956 B.n53 585
R332 B.n958 B.n957 585
R333 B.n959 B.n52 585
R334 B.n961 B.n960 585
R335 B.n962 B.n51 585
R336 B.n964 B.n963 585
R337 B.n965 B.n50 585
R338 B.n967 B.n966 585
R339 B.n968 B.n49 585
R340 B.n970 B.n969 585
R341 B.n971 B.n48 585
R342 B.n973 B.n972 585
R343 B.n974 B.n47 585
R344 B.n976 B.n975 585
R345 B.n977 B.n46 585
R346 B.n979 B.n978 585
R347 B.n980 B.n45 585
R348 B.n982 B.n981 585
R349 B.n983 B.n44 585
R350 B.n985 B.n984 585
R351 B.n986 B.n43 585
R352 B.n988 B.n987 585
R353 B.n989 B.n42 585
R354 B.n991 B.n990 585
R355 B.n992 B.n41 585
R356 B.n994 B.n993 585
R357 B.n995 B.n40 585
R358 B.n997 B.n996 585
R359 B.n998 B.n39 585
R360 B.n1000 B.n999 585
R361 B.n1001 B.n38 585
R362 B.n1003 B.n1002 585
R363 B.n803 B.n108 585
R364 B.n802 B.n801 585
R365 B.n800 B.n109 585
R366 B.n799 B.n798 585
R367 B.n797 B.n110 585
R368 B.n796 B.n795 585
R369 B.n794 B.n111 585
R370 B.n793 B.n792 585
R371 B.n791 B.n112 585
R372 B.n790 B.n789 585
R373 B.n788 B.n113 585
R374 B.n787 B.n786 585
R375 B.n785 B.n114 585
R376 B.n784 B.n783 585
R377 B.n782 B.n115 585
R378 B.n781 B.n780 585
R379 B.n779 B.n116 585
R380 B.n778 B.n777 585
R381 B.n776 B.n117 585
R382 B.n775 B.n774 585
R383 B.n773 B.n118 585
R384 B.n772 B.n771 585
R385 B.n770 B.n119 585
R386 B.n769 B.n768 585
R387 B.n767 B.n120 585
R388 B.n766 B.n765 585
R389 B.n764 B.n121 585
R390 B.n763 B.n762 585
R391 B.n761 B.n122 585
R392 B.n760 B.n759 585
R393 B.n758 B.n123 585
R394 B.n757 B.n756 585
R395 B.n755 B.n124 585
R396 B.n754 B.n753 585
R397 B.n752 B.n125 585
R398 B.n751 B.n750 585
R399 B.n749 B.n126 585
R400 B.n748 B.n747 585
R401 B.n746 B.n127 585
R402 B.n745 B.n744 585
R403 B.n743 B.n128 585
R404 B.n742 B.n741 585
R405 B.n740 B.n129 585
R406 B.n739 B.n738 585
R407 B.n737 B.n130 585
R408 B.n736 B.n735 585
R409 B.n734 B.n131 585
R410 B.n733 B.n732 585
R411 B.n731 B.n132 585
R412 B.n730 B.n729 585
R413 B.n728 B.n133 585
R414 B.n727 B.n726 585
R415 B.n725 B.n134 585
R416 B.n724 B.n723 585
R417 B.n722 B.n135 585
R418 B.n721 B.n720 585
R419 B.n719 B.n136 585
R420 B.n718 B.n717 585
R421 B.n716 B.n137 585
R422 B.n715 B.n714 585
R423 B.n713 B.n138 585
R424 B.n712 B.n711 585
R425 B.n710 B.n139 585
R426 B.n709 B.n708 585
R427 B.n707 B.n140 585
R428 B.n706 B.n705 585
R429 B.n704 B.n141 585
R430 B.n703 B.n702 585
R431 B.n701 B.n142 585
R432 B.n700 B.n699 585
R433 B.n698 B.n143 585
R434 B.n697 B.n696 585
R435 B.n695 B.n144 585
R436 B.n694 B.n693 585
R437 B.n692 B.n145 585
R438 B.n691 B.n690 585
R439 B.n689 B.n146 585
R440 B.n688 B.n687 585
R441 B.n686 B.n147 585
R442 B.n685 B.n684 585
R443 B.n683 B.n148 585
R444 B.n682 B.n681 585
R445 B.n680 B.n149 585
R446 B.n679 B.n678 585
R447 B.n677 B.n150 585
R448 B.n676 B.n675 585
R449 B.n674 B.n151 585
R450 B.n673 B.n672 585
R451 B.n671 B.n152 585
R452 B.n670 B.n669 585
R453 B.n668 B.n153 585
R454 B.n667 B.n666 585
R455 B.n665 B.n154 585
R456 B.n664 B.n663 585
R457 B.n662 B.n155 585
R458 B.n661 B.n660 585
R459 B.n659 B.n156 585
R460 B.n658 B.n657 585
R461 B.n656 B.n157 585
R462 B.n655 B.n654 585
R463 B.n653 B.n158 585
R464 B.n652 B.n651 585
R465 B.n650 B.n159 585
R466 B.n649 B.n648 585
R467 B.n647 B.n160 585
R468 B.n646 B.n645 585
R469 B.n644 B.n161 585
R470 B.n643 B.n642 585
R471 B.n641 B.n162 585
R472 B.n640 B.n639 585
R473 B.n638 B.n163 585
R474 B.n637 B.n636 585
R475 B.n635 B.n164 585
R476 B.n634 B.n633 585
R477 B.n632 B.n165 585
R478 B.n631 B.n630 585
R479 B.n629 B.n166 585
R480 B.n628 B.n627 585
R481 B.n626 B.n167 585
R482 B.n625 B.n624 585
R483 B.n623 B.n168 585
R484 B.n622 B.n621 585
R485 B.n620 B.n169 585
R486 B.n619 B.n618 585
R487 B.n617 B.n170 585
R488 B.n616 B.n615 585
R489 B.n614 B.n171 585
R490 B.n613 B.n612 585
R491 B.n611 B.n172 585
R492 B.n610 B.n609 585
R493 B.n608 B.n173 585
R494 B.n607 B.n606 585
R495 B.n605 B.n174 585
R496 B.n604 B.n603 585
R497 B.n602 B.n175 585
R498 B.n601 B.n600 585
R499 B.n599 B.n176 585
R500 B.n598 B.n597 585
R501 B.n596 B.n177 585
R502 B.n595 B.n594 585
R503 B.n593 B.n178 585
R504 B.n592 B.n591 585
R505 B.n590 B.n179 585
R506 B.n391 B.n390 585
R507 B.n392 B.n249 585
R508 B.n394 B.n393 585
R509 B.n395 B.n248 585
R510 B.n397 B.n396 585
R511 B.n398 B.n247 585
R512 B.n400 B.n399 585
R513 B.n401 B.n246 585
R514 B.n403 B.n402 585
R515 B.n404 B.n245 585
R516 B.n406 B.n405 585
R517 B.n407 B.n244 585
R518 B.n409 B.n408 585
R519 B.n410 B.n243 585
R520 B.n412 B.n411 585
R521 B.n413 B.n242 585
R522 B.n415 B.n414 585
R523 B.n416 B.n241 585
R524 B.n418 B.n417 585
R525 B.n419 B.n240 585
R526 B.n421 B.n420 585
R527 B.n422 B.n239 585
R528 B.n424 B.n423 585
R529 B.n425 B.n238 585
R530 B.n427 B.n426 585
R531 B.n428 B.n237 585
R532 B.n430 B.n429 585
R533 B.n431 B.n236 585
R534 B.n433 B.n432 585
R535 B.n434 B.n235 585
R536 B.n436 B.n435 585
R537 B.n437 B.n234 585
R538 B.n439 B.n438 585
R539 B.n440 B.n233 585
R540 B.n442 B.n441 585
R541 B.n443 B.n232 585
R542 B.n445 B.n444 585
R543 B.n446 B.n231 585
R544 B.n448 B.n447 585
R545 B.n449 B.n230 585
R546 B.n451 B.n450 585
R547 B.n452 B.n229 585
R548 B.n454 B.n453 585
R549 B.n455 B.n228 585
R550 B.n457 B.n456 585
R551 B.n458 B.n227 585
R552 B.n460 B.n459 585
R553 B.n461 B.n226 585
R554 B.n463 B.n462 585
R555 B.n464 B.n225 585
R556 B.n466 B.n465 585
R557 B.n467 B.n224 585
R558 B.n469 B.n468 585
R559 B.n470 B.n223 585
R560 B.n472 B.n471 585
R561 B.n473 B.n222 585
R562 B.n475 B.n474 585
R563 B.n476 B.n221 585
R564 B.n478 B.n477 585
R565 B.n479 B.n220 585
R566 B.n481 B.n480 585
R567 B.n483 B.n217 585
R568 B.n485 B.n484 585
R569 B.n486 B.n216 585
R570 B.n488 B.n487 585
R571 B.n489 B.n215 585
R572 B.n491 B.n490 585
R573 B.n492 B.n214 585
R574 B.n494 B.n493 585
R575 B.n495 B.n213 585
R576 B.n497 B.n496 585
R577 B.n499 B.n498 585
R578 B.n500 B.n209 585
R579 B.n502 B.n501 585
R580 B.n503 B.n208 585
R581 B.n505 B.n504 585
R582 B.n506 B.n207 585
R583 B.n508 B.n507 585
R584 B.n509 B.n206 585
R585 B.n511 B.n510 585
R586 B.n512 B.n205 585
R587 B.n514 B.n513 585
R588 B.n515 B.n204 585
R589 B.n517 B.n516 585
R590 B.n518 B.n203 585
R591 B.n520 B.n519 585
R592 B.n521 B.n202 585
R593 B.n523 B.n522 585
R594 B.n524 B.n201 585
R595 B.n526 B.n525 585
R596 B.n527 B.n200 585
R597 B.n529 B.n528 585
R598 B.n530 B.n199 585
R599 B.n532 B.n531 585
R600 B.n533 B.n198 585
R601 B.n535 B.n534 585
R602 B.n536 B.n197 585
R603 B.n538 B.n537 585
R604 B.n539 B.n196 585
R605 B.n541 B.n540 585
R606 B.n542 B.n195 585
R607 B.n544 B.n543 585
R608 B.n545 B.n194 585
R609 B.n547 B.n546 585
R610 B.n548 B.n193 585
R611 B.n550 B.n549 585
R612 B.n551 B.n192 585
R613 B.n553 B.n552 585
R614 B.n554 B.n191 585
R615 B.n556 B.n555 585
R616 B.n557 B.n190 585
R617 B.n559 B.n558 585
R618 B.n560 B.n189 585
R619 B.n562 B.n561 585
R620 B.n563 B.n188 585
R621 B.n565 B.n564 585
R622 B.n566 B.n187 585
R623 B.n568 B.n567 585
R624 B.n569 B.n186 585
R625 B.n571 B.n570 585
R626 B.n572 B.n185 585
R627 B.n574 B.n573 585
R628 B.n575 B.n184 585
R629 B.n577 B.n576 585
R630 B.n578 B.n183 585
R631 B.n580 B.n579 585
R632 B.n581 B.n182 585
R633 B.n583 B.n582 585
R634 B.n584 B.n181 585
R635 B.n586 B.n585 585
R636 B.n587 B.n180 585
R637 B.n589 B.n588 585
R638 B.n389 B.n250 585
R639 B.n388 B.n387 585
R640 B.n386 B.n251 585
R641 B.n385 B.n384 585
R642 B.n383 B.n252 585
R643 B.n382 B.n381 585
R644 B.n380 B.n253 585
R645 B.n379 B.n378 585
R646 B.n377 B.n254 585
R647 B.n376 B.n375 585
R648 B.n374 B.n255 585
R649 B.n373 B.n372 585
R650 B.n371 B.n256 585
R651 B.n370 B.n369 585
R652 B.n368 B.n257 585
R653 B.n367 B.n366 585
R654 B.n365 B.n258 585
R655 B.n364 B.n363 585
R656 B.n362 B.n259 585
R657 B.n361 B.n360 585
R658 B.n359 B.n260 585
R659 B.n358 B.n357 585
R660 B.n356 B.n261 585
R661 B.n355 B.n354 585
R662 B.n353 B.n262 585
R663 B.n352 B.n351 585
R664 B.n350 B.n263 585
R665 B.n349 B.n348 585
R666 B.n347 B.n264 585
R667 B.n346 B.n345 585
R668 B.n344 B.n265 585
R669 B.n343 B.n342 585
R670 B.n341 B.n266 585
R671 B.n340 B.n339 585
R672 B.n338 B.n267 585
R673 B.n337 B.n336 585
R674 B.n335 B.n268 585
R675 B.n334 B.n333 585
R676 B.n332 B.n269 585
R677 B.n331 B.n330 585
R678 B.n329 B.n270 585
R679 B.n328 B.n327 585
R680 B.n326 B.n271 585
R681 B.n325 B.n324 585
R682 B.n323 B.n272 585
R683 B.n322 B.n321 585
R684 B.n320 B.n273 585
R685 B.n319 B.n318 585
R686 B.n317 B.n274 585
R687 B.n316 B.n315 585
R688 B.n314 B.n275 585
R689 B.n313 B.n312 585
R690 B.n311 B.n276 585
R691 B.n310 B.n309 585
R692 B.n308 B.n277 585
R693 B.n307 B.n306 585
R694 B.n305 B.n278 585
R695 B.n304 B.n303 585
R696 B.n302 B.n279 585
R697 B.n301 B.n300 585
R698 B.n299 B.n280 585
R699 B.n298 B.n297 585
R700 B.n296 B.n281 585
R701 B.n295 B.n294 585
R702 B.n293 B.n282 585
R703 B.n292 B.n291 585
R704 B.n290 B.n283 585
R705 B.n289 B.n288 585
R706 B.n287 B.n284 585
R707 B.n286 B.n285 585
R708 B.n2 B.n0 585
R709 B.n1109 B.n1 585
R710 B.n1108 B.n1107 585
R711 B.n1106 B.n3 585
R712 B.n1105 B.n1104 585
R713 B.n1103 B.n4 585
R714 B.n1102 B.n1101 585
R715 B.n1100 B.n5 585
R716 B.n1099 B.n1098 585
R717 B.n1097 B.n6 585
R718 B.n1096 B.n1095 585
R719 B.n1094 B.n7 585
R720 B.n1093 B.n1092 585
R721 B.n1091 B.n8 585
R722 B.n1090 B.n1089 585
R723 B.n1088 B.n9 585
R724 B.n1087 B.n1086 585
R725 B.n1085 B.n10 585
R726 B.n1084 B.n1083 585
R727 B.n1082 B.n11 585
R728 B.n1081 B.n1080 585
R729 B.n1079 B.n12 585
R730 B.n1078 B.n1077 585
R731 B.n1076 B.n13 585
R732 B.n1075 B.n1074 585
R733 B.n1073 B.n14 585
R734 B.n1072 B.n1071 585
R735 B.n1070 B.n15 585
R736 B.n1069 B.n1068 585
R737 B.n1067 B.n16 585
R738 B.n1066 B.n1065 585
R739 B.n1064 B.n17 585
R740 B.n1063 B.n1062 585
R741 B.n1061 B.n18 585
R742 B.n1060 B.n1059 585
R743 B.n1058 B.n19 585
R744 B.n1057 B.n1056 585
R745 B.n1055 B.n20 585
R746 B.n1054 B.n1053 585
R747 B.n1052 B.n21 585
R748 B.n1051 B.n1050 585
R749 B.n1049 B.n22 585
R750 B.n1048 B.n1047 585
R751 B.n1046 B.n23 585
R752 B.n1045 B.n1044 585
R753 B.n1043 B.n24 585
R754 B.n1042 B.n1041 585
R755 B.n1040 B.n25 585
R756 B.n1039 B.n1038 585
R757 B.n1037 B.n26 585
R758 B.n1036 B.n1035 585
R759 B.n1034 B.n27 585
R760 B.n1033 B.n1032 585
R761 B.n1031 B.n28 585
R762 B.n1030 B.n1029 585
R763 B.n1028 B.n29 585
R764 B.n1027 B.n1026 585
R765 B.n1025 B.n30 585
R766 B.n1024 B.n1023 585
R767 B.n1022 B.n31 585
R768 B.n1021 B.n1020 585
R769 B.n1019 B.n32 585
R770 B.n1018 B.n1017 585
R771 B.n1016 B.n33 585
R772 B.n1015 B.n1014 585
R773 B.n1013 B.n34 585
R774 B.n1012 B.n1011 585
R775 B.n1010 B.n35 585
R776 B.n1009 B.n1008 585
R777 B.n1007 B.n36 585
R778 B.n1006 B.n1005 585
R779 B.n1004 B.n37 585
R780 B.n1111 B.n1110 585
R781 B.n390 B.n389 545.355
R782 B.n1002 B.n37 545.355
R783 B.n588 B.n179 545.355
R784 B.n804 B.n803 545.355
R785 B.n210 B.t9 347.226
R786 B.n218 B.t6 347.226
R787 B.n68 B.t3 347.226
R788 B.n76 B.t0 347.226
R789 B.n210 B.t11 181.389
R790 B.n76 B.t1 181.389
R791 B.n218 B.t8 181.365
R792 B.n68 B.t4 181.365
R793 B.n389 B.n388 163.367
R794 B.n388 B.n251 163.367
R795 B.n384 B.n251 163.367
R796 B.n384 B.n383 163.367
R797 B.n383 B.n382 163.367
R798 B.n382 B.n253 163.367
R799 B.n378 B.n253 163.367
R800 B.n378 B.n377 163.367
R801 B.n377 B.n376 163.367
R802 B.n376 B.n255 163.367
R803 B.n372 B.n255 163.367
R804 B.n372 B.n371 163.367
R805 B.n371 B.n370 163.367
R806 B.n370 B.n257 163.367
R807 B.n366 B.n257 163.367
R808 B.n366 B.n365 163.367
R809 B.n365 B.n364 163.367
R810 B.n364 B.n259 163.367
R811 B.n360 B.n259 163.367
R812 B.n360 B.n359 163.367
R813 B.n359 B.n358 163.367
R814 B.n358 B.n261 163.367
R815 B.n354 B.n261 163.367
R816 B.n354 B.n353 163.367
R817 B.n353 B.n352 163.367
R818 B.n352 B.n263 163.367
R819 B.n348 B.n263 163.367
R820 B.n348 B.n347 163.367
R821 B.n347 B.n346 163.367
R822 B.n346 B.n265 163.367
R823 B.n342 B.n265 163.367
R824 B.n342 B.n341 163.367
R825 B.n341 B.n340 163.367
R826 B.n340 B.n267 163.367
R827 B.n336 B.n267 163.367
R828 B.n336 B.n335 163.367
R829 B.n335 B.n334 163.367
R830 B.n334 B.n269 163.367
R831 B.n330 B.n269 163.367
R832 B.n330 B.n329 163.367
R833 B.n329 B.n328 163.367
R834 B.n328 B.n271 163.367
R835 B.n324 B.n271 163.367
R836 B.n324 B.n323 163.367
R837 B.n323 B.n322 163.367
R838 B.n322 B.n273 163.367
R839 B.n318 B.n273 163.367
R840 B.n318 B.n317 163.367
R841 B.n317 B.n316 163.367
R842 B.n316 B.n275 163.367
R843 B.n312 B.n275 163.367
R844 B.n312 B.n311 163.367
R845 B.n311 B.n310 163.367
R846 B.n310 B.n277 163.367
R847 B.n306 B.n277 163.367
R848 B.n306 B.n305 163.367
R849 B.n305 B.n304 163.367
R850 B.n304 B.n279 163.367
R851 B.n300 B.n279 163.367
R852 B.n300 B.n299 163.367
R853 B.n299 B.n298 163.367
R854 B.n298 B.n281 163.367
R855 B.n294 B.n281 163.367
R856 B.n294 B.n293 163.367
R857 B.n293 B.n292 163.367
R858 B.n292 B.n283 163.367
R859 B.n288 B.n283 163.367
R860 B.n288 B.n287 163.367
R861 B.n287 B.n286 163.367
R862 B.n286 B.n2 163.367
R863 B.n1110 B.n2 163.367
R864 B.n1110 B.n1109 163.367
R865 B.n1109 B.n1108 163.367
R866 B.n1108 B.n3 163.367
R867 B.n1104 B.n3 163.367
R868 B.n1104 B.n1103 163.367
R869 B.n1103 B.n1102 163.367
R870 B.n1102 B.n5 163.367
R871 B.n1098 B.n5 163.367
R872 B.n1098 B.n1097 163.367
R873 B.n1097 B.n1096 163.367
R874 B.n1096 B.n7 163.367
R875 B.n1092 B.n7 163.367
R876 B.n1092 B.n1091 163.367
R877 B.n1091 B.n1090 163.367
R878 B.n1090 B.n9 163.367
R879 B.n1086 B.n9 163.367
R880 B.n1086 B.n1085 163.367
R881 B.n1085 B.n1084 163.367
R882 B.n1084 B.n11 163.367
R883 B.n1080 B.n11 163.367
R884 B.n1080 B.n1079 163.367
R885 B.n1079 B.n1078 163.367
R886 B.n1078 B.n13 163.367
R887 B.n1074 B.n13 163.367
R888 B.n1074 B.n1073 163.367
R889 B.n1073 B.n1072 163.367
R890 B.n1072 B.n15 163.367
R891 B.n1068 B.n15 163.367
R892 B.n1068 B.n1067 163.367
R893 B.n1067 B.n1066 163.367
R894 B.n1066 B.n17 163.367
R895 B.n1062 B.n17 163.367
R896 B.n1062 B.n1061 163.367
R897 B.n1061 B.n1060 163.367
R898 B.n1060 B.n19 163.367
R899 B.n1056 B.n19 163.367
R900 B.n1056 B.n1055 163.367
R901 B.n1055 B.n1054 163.367
R902 B.n1054 B.n21 163.367
R903 B.n1050 B.n21 163.367
R904 B.n1050 B.n1049 163.367
R905 B.n1049 B.n1048 163.367
R906 B.n1048 B.n23 163.367
R907 B.n1044 B.n23 163.367
R908 B.n1044 B.n1043 163.367
R909 B.n1043 B.n1042 163.367
R910 B.n1042 B.n25 163.367
R911 B.n1038 B.n25 163.367
R912 B.n1038 B.n1037 163.367
R913 B.n1037 B.n1036 163.367
R914 B.n1036 B.n27 163.367
R915 B.n1032 B.n27 163.367
R916 B.n1032 B.n1031 163.367
R917 B.n1031 B.n1030 163.367
R918 B.n1030 B.n29 163.367
R919 B.n1026 B.n29 163.367
R920 B.n1026 B.n1025 163.367
R921 B.n1025 B.n1024 163.367
R922 B.n1024 B.n31 163.367
R923 B.n1020 B.n31 163.367
R924 B.n1020 B.n1019 163.367
R925 B.n1019 B.n1018 163.367
R926 B.n1018 B.n33 163.367
R927 B.n1014 B.n33 163.367
R928 B.n1014 B.n1013 163.367
R929 B.n1013 B.n1012 163.367
R930 B.n1012 B.n35 163.367
R931 B.n1008 B.n35 163.367
R932 B.n1008 B.n1007 163.367
R933 B.n1007 B.n1006 163.367
R934 B.n1006 B.n37 163.367
R935 B.n390 B.n249 163.367
R936 B.n394 B.n249 163.367
R937 B.n395 B.n394 163.367
R938 B.n396 B.n395 163.367
R939 B.n396 B.n247 163.367
R940 B.n400 B.n247 163.367
R941 B.n401 B.n400 163.367
R942 B.n402 B.n401 163.367
R943 B.n402 B.n245 163.367
R944 B.n406 B.n245 163.367
R945 B.n407 B.n406 163.367
R946 B.n408 B.n407 163.367
R947 B.n408 B.n243 163.367
R948 B.n412 B.n243 163.367
R949 B.n413 B.n412 163.367
R950 B.n414 B.n413 163.367
R951 B.n414 B.n241 163.367
R952 B.n418 B.n241 163.367
R953 B.n419 B.n418 163.367
R954 B.n420 B.n419 163.367
R955 B.n420 B.n239 163.367
R956 B.n424 B.n239 163.367
R957 B.n425 B.n424 163.367
R958 B.n426 B.n425 163.367
R959 B.n426 B.n237 163.367
R960 B.n430 B.n237 163.367
R961 B.n431 B.n430 163.367
R962 B.n432 B.n431 163.367
R963 B.n432 B.n235 163.367
R964 B.n436 B.n235 163.367
R965 B.n437 B.n436 163.367
R966 B.n438 B.n437 163.367
R967 B.n438 B.n233 163.367
R968 B.n442 B.n233 163.367
R969 B.n443 B.n442 163.367
R970 B.n444 B.n443 163.367
R971 B.n444 B.n231 163.367
R972 B.n448 B.n231 163.367
R973 B.n449 B.n448 163.367
R974 B.n450 B.n449 163.367
R975 B.n450 B.n229 163.367
R976 B.n454 B.n229 163.367
R977 B.n455 B.n454 163.367
R978 B.n456 B.n455 163.367
R979 B.n456 B.n227 163.367
R980 B.n460 B.n227 163.367
R981 B.n461 B.n460 163.367
R982 B.n462 B.n461 163.367
R983 B.n462 B.n225 163.367
R984 B.n466 B.n225 163.367
R985 B.n467 B.n466 163.367
R986 B.n468 B.n467 163.367
R987 B.n468 B.n223 163.367
R988 B.n472 B.n223 163.367
R989 B.n473 B.n472 163.367
R990 B.n474 B.n473 163.367
R991 B.n474 B.n221 163.367
R992 B.n478 B.n221 163.367
R993 B.n479 B.n478 163.367
R994 B.n480 B.n479 163.367
R995 B.n480 B.n217 163.367
R996 B.n485 B.n217 163.367
R997 B.n486 B.n485 163.367
R998 B.n487 B.n486 163.367
R999 B.n487 B.n215 163.367
R1000 B.n491 B.n215 163.367
R1001 B.n492 B.n491 163.367
R1002 B.n493 B.n492 163.367
R1003 B.n493 B.n213 163.367
R1004 B.n497 B.n213 163.367
R1005 B.n498 B.n497 163.367
R1006 B.n498 B.n209 163.367
R1007 B.n502 B.n209 163.367
R1008 B.n503 B.n502 163.367
R1009 B.n504 B.n503 163.367
R1010 B.n504 B.n207 163.367
R1011 B.n508 B.n207 163.367
R1012 B.n509 B.n508 163.367
R1013 B.n510 B.n509 163.367
R1014 B.n510 B.n205 163.367
R1015 B.n514 B.n205 163.367
R1016 B.n515 B.n514 163.367
R1017 B.n516 B.n515 163.367
R1018 B.n516 B.n203 163.367
R1019 B.n520 B.n203 163.367
R1020 B.n521 B.n520 163.367
R1021 B.n522 B.n521 163.367
R1022 B.n522 B.n201 163.367
R1023 B.n526 B.n201 163.367
R1024 B.n527 B.n526 163.367
R1025 B.n528 B.n527 163.367
R1026 B.n528 B.n199 163.367
R1027 B.n532 B.n199 163.367
R1028 B.n533 B.n532 163.367
R1029 B.n534 B.n533 163.367
R1030 B.n534 B.n197 163.367
R1031 B.n538 B.n197 163.367
R1032 B.n539 B.n538 163.367
R1033 B.n540 B.n539 163.367
R1034 B.n540 B.n195 163.367
R1035 B.n544 B.n195 163.367
R1036 B.n545 B.n544 163.367
R1037 B.n546 B.n545 163.367
R1038 B.n546 B.n193 163.367
R1039 B.n550 B.n193 163.367
R1040 B.n551 B.n550 163.367
R1041 B.n552 B.n551 163.367
R1042 B.n552 B.n191 163.367
R1043 B.n556 B.n191 163.367
R1044 B.n557 B.n556 163.367
R1045 B.n558 B.n557 163.367
R1046 B.n558 B.n189 163.367
R1047 B.n562 B.n189 163.367
R1048 B.n563 B.n562 163.367
R1049 B.n564 B.n563 163.367
R1050 B.n564 B.n187 163.367
R1051 B.n568 B.n187 163.367
R1052 B.n569 B.n568 163.367
R1053 B.n570 B.n569 163.367
R1054 B.n570 B.n185 163.367
R1055 B.n574 B.n185 163.367
R1056 B.n575 B.n574 163.367
R1057 B.n576 B.n575 163.367
R1058 B.n576 B.n183 163.367
R1059 B.n580 B.n183 163.367
R1060 B.n581 B.n580 163.367
R1061 B.n582 B.n581 163.367
R1062 B.n582 B.n181 163.367
R1063 B.n586 B.n181 163.367
R1064 B.n587 B.n586 163.367
R1065 B.n588 B.n587 163.367
R1066 B.n592 B.n179 163.367
R1067 B.n593 B.n592 163.367
R1068 B.n594 B.n593 163.367
R1069 B.n594 B.n177 163.367
R1070 B.n598 B.n177 163.367
R1071 B.n599 B.n598 163.367
R1072 B.n600 B.n599 163.367
R1073 B.n600 B.n175 163.367
R1074 B.n604 B.n175 163.367
R1075 B.n605 B.n604 163.367
R1076 B.n606 B.n605 163.367
R1077 B.n606 B.n173 163.367
R1078 B.n610 B.n173 163.367
R1079 B.n611 B.n610 163.367
R1080 B.n612 B.n611 163.367
R1081 B.n612 B.n171 163.367
R1082 B.n616 B.n171 163.367
R1083 B.n617 B.n616 163.367
R1084 B.n618 B.n617 163.367
R1085 B.n618 B.n169 163.367
R1086 B.n622 B.n169 163.367
R1087 B.n623 B.n622 163.367
R1088 B.n624 B.n623 163.367
R1089 B.n624 B.n167 163.367
R1090 B.n628 B.n167 163.367
R1091 B.n629 B.n628 163.367
R1092 B.n630 B.n629 163.367
R1093 B.n630 B.n165 163.367
R1094 B.n634 B.n165 163.367
R1095 B.n635 B.n634 163.367
R1096 B.n636 B.n635 163.367
R1097 B.n636 B.n163 163.367
R1098 B.n640 B.n163 163.367
R1099 B.n641 B.n640 163.367
R1100 B.n642 B.n641 163.367
R1101 B.n642 B.n161 163.367
R1102 B.n646 B.n161 163.367
R1103 B.n647 B.n646 163.367
R1104 B.n648 B.n647 163.367
R1105 B.n648 B.n159 163.367
R1106 B.n652 B.n159 163.367
R1107 B.n653 B.n652 163.367
R1108 B.n654 B.n653 163.367
R1109 B.n654 B.n157 163.367
R1110 B.n658 B.n157 163.367
R1111 B.n659 B.n658 163.367
R1112 B.n660 B.n659 163.367
R1113 B.n660 B.n155 163.367
R1114 B.n664 B.n155 163.367
R1115 B.n665 B.n664 163.367
R1116 B.n666 B.n665 163.367
R1117 B.n666 B.n153 163.367
R1118 B.n670 B.n153 163.367
R1119 B.n671 B.n670 163.367
R1120 B.n672 B.n671 163.367
R1121 B.n672 B.n151 163.367
R1122 B.n676 B.n151 163.367
R1123 B.n677 B.n676 163.367
R1124 B.n678 B.n677 163.367
R1125 B.n678 B.n149 163.367
R1126 B.n682 B.n149 163.367
R1127 B.n683 B.n682 163.367
R1128 B.n684 B.n683 163.367
R1129 B.n684 B.n147 163.367
R1130 B.n688 B.n147 163.367
R1131 B.n689 B.n688 163.367
R1132 B.n690 B.n689 163.367
R1133 B.n690 B.n145 163.367
R1134 B.n694 B.n145 163.367
R1135 B.n695 B.n694 163.367
R1136 B.n696 B.n695 163.367
R1137 B.n696 B.n143 163.367
R1138 B.n700 B.n143 163.367
R1139 B.n701 B.n700 163.367
R1140 B.n702 B.n701 163.367
R1141 B.n702 B.n141 163.367
R1142 B.n706 B.n141 163.367
R1143 B.n707 B.n706 163.367
R1144 B.n708 B.n707 163.367
R1145 B.n708 B.n139 163.367
R1146 B.n712 B.n139 163.367
R1147 B.n713 B.n712 163.367
R1148 B.n714 B.n713 163.367
R1149 B.n714 B.n137 163.367
R1150 B.n718 B.n137 163.367
R1151 B.n719 B.n718 163.367
R1152 B.n720 B.n719 163.367
R1153 B.n720 B.n135 163.367
R1154 B.n724 B.n135 163.367
R1155 B.n725 B.n724 163.367
R1156 B.n726 B.n725 163.367
R1157 B.n726 B.n133 163.367
R1158 B.n730 B.n133 163.367
R1159 B.n731 B.n730 163.367
R1160 B.n732 B.n731 163.367
R1161 B.n732 B.n131 163.367
R1162 B.n736 B.n131 163.367
R1163 B.n737 B.n736 163.367
R1164 B.n738 B.n737 163.367
R1165 B.n738 B.n129 163.367
R1166 B.n742 B.n129 163.367
R1167 B.n743 B.n742 163.367
R1168 B.n744 B.n743 163.367
R1169 B.n744 B.n127 163.367
R1170 B.n748 B.n127 163.367
R1171 B.n749 B.n748 163.367
R1172 B.n750 B.n749 163.367
R1173 B.n750 B.n125 163.367
R1174 B.n754 B.n125 163.367
R1175 B.n755 B.n754 163.367
R1176 B.n756 B.n755 163.367
R1177 B.n756 B.n123 163.367
R1178 B.n760 B.n123 163.367
R1179 B.n761 B.n760 163.367
R1180 B.n762 B.n761 163.367
R1181 B.n762 B.n121 163.367
R1182 B.n766 B.n121 163.367
R1183 B.n767 B.n766 163.367
R1184 B.n768 B.n767 163.367
R1185 B.n768 B.n119 163.367
R1186 B.n772 B.n119 163.367
R1187 B.n773 B.n772 163.367
R1188 B.n774 B.n773 163.367
R1189 B.n774 B.n117 163.367
R1190 B.n778 B.n117 163.367
R1191 B.n779 B.n778 163.367
R1192 B.n780 B.n779 163.367
R1193 B.n780 B.n115 163.367
R1194 B.n784 B.n115 163.367
R1195 B.n785 B.n784 163.367
R1196 B.n786 B.n785 163.367
R1197 B.n786 B.n113 163.367
R1198 B.n790 B.n113 163.367
R1199 B.n791 B.n790 163.367
R1200 B.n792 B.n791 163.367
R1201 B.n792 B.n111 163.367
R1202 B.n796 B.n111 163.367
R1203 B.n797 B.n796 163.367
R1204 B.n798 B.n797 163.367
R1205 B.n798 B.n109 163.367
R1206 B.n802 B.n109 163.367
R1207 B.n803 B.n802 163.367
R1208 B.n1002 B.n1001 163.367
R1209 B.n1001 B.n1000 163.367
R1210 B.n1000 B.n39 163.367
R1211 B.n996 B.n39 163.367
R1212 B.n996 B.n995 163.367
R1213 B.n995 B.n994 163.367
R1214 B.n994 B.n41 163.367
R1215 B.n990 B.n41 163.367
R1216 B.n990 B.n989 163.367
R1217 B.n989 B.n988 163.367
R1218 B.n988 B.n43 163.367
R1219 B.n984 B.n43 163.367
R1220 B.n984 B.n983 163.367
R1221 B.n983 B.n982 163.367
R1222 B.n982 B.n45 163.367
R1223 B.n978 B.n45 163.367
R1224 B.n978 B.n977 163.367
R1225 B.n977 B.n976 163.367
R1226 B.n976 B.n47 163.367
R1227 B.n972 B.n47 163.367
R1228 B.n972 B.n971 163.367
R1229 B.n971 B.n970 163.367
R1230 B.n970 B.n49 163.367
R1231 B.n966 B.n49 163.367
R1232 B.n966 B.n965 163.367
R1233 B.n965 B.n964 163.367
R1234 B.n964 B.n51 163.367
R1235 B.n960 B.n51 163.367
R1236 B.n960 B.n959 163.367
R1237 B.n959 B.n958 163.367
R1238 B.n958 B.n53 163.367
R1239 B.n954 B.n53 163.367
R1240 B.n954 B.n953 163.367
R1241 B.n953 B.n952 163.367
R1242 B.n952 B.n55 163.367
R1243 B.n948 B.n55 163.367
R1244 B.n948 B.n947 163.367
R1245 B.n947 B.n946 163.367
R1246 B.n946 B.n57 163.367
R1247 B.n942 B.n57 163.367
R1248 B.n942 B.n941 163.367
R1249 B.n941 B.n940 163.367
R1250 B.n940 B.n59 163.367
R1251 B.n936 B.n59 163.367
R1252 B.n936 B.n935 163.367
R1253 B.n935 B.n934 163.367
R1254 B.n934 B.n61 163.367
R1255 B.n930 B.n61 163.367
R1256 B.n930 B.n929 163.367
R1257 B.n929 B.n928 163.367
R1258 B.n928 B.n63 163.367
R1259 B.n924 B.n63 163.367
R1260 B.n924 B.n923 163.367
R1261 B.n923 B.n922 163.367
R1262 B.n922 B.n65 163.367
R1263 B.n918 B.n65 163.367
R1264 B.n918 B.n917 163.367
R1265 B.n917 B.n916 163.367
R1266 B.n916 B.n67 163.367
R1267 B.n912 B.n67 163.367
R1268 B.n912 B.n911 163.367
R1269 B.n911 B.n71 163.367
R1270 B.n907 B.n71 163.367
R1271 B.n907 B.n906 163.367
R1272 B.n906 B.n905 163.367
R1273 B.n905 B.n73 163.367
R1274 B.n901 B.n73 163.367
R1275 B.n901 B.n900 163.367
R1276 B.n900 B.n899 163.367
R1277 B.n899 B.n75 163.367
R1278 B.n894 B.n75 163.367
R1279 B.n894 B.n893 163.367
R1280 B.n893 B.n892 163.367
R1281 B.n892 B.n79 163.367
R1282 B.n888 B.n79 163.367
R1283 B.n888 B.n887 163.367
R1284 B.n887 B.n886 163.367
R1285 B.n886 B.n81 163.367
R1286 B.n882 B.n81 163.367
R1287 B.n882 B.n881 163.367
R1288 B.n881 B.n880 163.367
R1289 B.n880 B.n83 163.367
R1290 B.n876 B.n83 163.367
R1291 B.n876 B.n875 163.367
R1292 B.n875 B.n874 163.367
R1293 B.n874 B.n85 163.367
R1294 B.n870 B.n85 163.367
R1295 B.n870 B.n869 163.367
R1296 B.n869 B.n868 163.367
R1297 B.n868 B.n87 163.367
R1298 B.n864 B.n87 163.367
R1299 B.n864 B.n863 163.367
R1300 B.n863 B.n862 163.367
R1301 B.n862 B.n89 163.367
R1302 B.n858 B.n89 163.367
R1303 B.n858 B.n857 163.367
R1304 B.n857 B.n856 163.367
R1305 B.n856 B.n91 163.367
R1306 B.n852 B.n91 163.367
R1307 B.n852 B.n851 163.367
R1308 B.n851 B.n850 163.367
R1309 B.n850 B.n93 163.367
R1310 B.n846 B.n93 163.367
R1311 B.n846 B.n845 163.367
R1312 B.n845 B.n844 163.367
R1313 B.n844 B.n95 163.367
R1314 B.n840 B.n95 163.367
R1315 B.n840 B.n839 163.367
R1316 B.n839 B.n838 163.367
R1317 B.n838 B.n97 163.367
R1318 B.n834 B.n97 163.367
R1319 B.n834 B.n833 163.367
R1320 B.n833 B.n832 163.367
R1321 B.n832 B.n99 163.367
R1322 B.n828 B.n99 163.367
R1323 B.n828 B.n827 163.367
R1324 B.n827 B.n826 163.367
R1325 B.n826 B.n101 163.367
R1326 B.n822 B.n101 163.367
R1327 B.n822 B.n821 163.367
R1328 B.n821 B.n820 163.367
R1329 B.n820 B.n103 163.367
R1330 B.n816 B.n103 163.367
R1331 B.n816 B.n815 163.367
R1332 B.n815 B.n814 163.367
R1333 B.n814 B.n105 163.367
R1334 B.n810 B.n105 163.367
R1335 B.n810 B.n809 163.367
R1336 B.n809 B.n808 163.367
R1337 B.n808 B.n107 163.367
R1338 B.n804 B.n107 163.367
R1339 B.n211 B.t10 111.96
R1340 B.n77 B.t2 111.96
R1341 B.n219 B.t7 111.936
R1342 B.n69 B.t5 111.936
R1343 B.n211 B.n210 69.4308
R1344 B.n219 B.n218 69.4308
R1345 B.n69 B.n68 69.4308
R1346 B.n77 B.n76 69.4308
R1347 B.n212 B.n211 59.5399
R1348 B.n482 B.n219 59.5399
R1349 B.n70 B.n69 59.5399
R1350 B.n896 B.n77 59.5399
R1351 B.n1004 B.n1003 35.4346
R1352 B.n805 B.n108 35.4346
R1353 B.n590 B.n589 35.4346
R1354 B.n391 B.n250 35.4346
R1355 B B.n1111 18.0485
R1356 B.n1003 B.n38 10.6151
R1357 B.n999 B.n38 10.6151
R1358 B.n999 B.n998 10.6151
R1359 B.n998 B.n997 10.6151
R1360 B.n997 B.n40 10.6151
R1361 B.n993 B.n40 10.6151
R1362 B.n993 B.n992 10.6151
R1363 B.n992 B.n991 10.6151
R1364 B.n991 B.n42 10.6151
R1365 B.n987 B.n42 10.6151
R1366 B.n987 B.n986 10.6151
R1367 B.n986 B.n985 10.6151
R1368 B.n985 B.n44 10.6151
R1369 B.n981 B.n44 10.6151
R1370 B.n981 B.n980 10.6151
R1371 B.n980 B.n979 10.6151
R1372 B.n979 B.n46 10.6151
R1373 B.n975 B.n46 10.6151
R1374 B.n975 B.n974 10.6151
R1375 B.n974 B.n973 10.6151
R1376 B.n973 B.n48 10.6151
R1377 B.n969 B.n48 10.6151
R1378 B.n969 B.n968 10.6151
R1379 B.n968 B.n967 10.6151
R1380 B.n967 B.n50 10.6151
R1381 B.n963 B.n50 10.6151
R1382 B.n963 B.n962 10.6151
R1383 B.n962 B.n961 10.6151
R1384 B.n961 B.n52 10.6151
R1385 B.n957 B.n52 10.6151
R1386 B.n957 B.n956 10.6151
R1387 B.n956 B.n955 10.6151
R1388 B.n955 B.n54 10.6151
R1389 B.n951 B.n54 10.6151
R1390 B.n951 B.n950 10.6151
R1391 B.n950 B.n949 10.6151
R1392 B.n949 B.n56 10.6151
R1393 B.n945 B.n56 10.6151
R1394 B.n945 B.n944 10.6151
R1395 B.n944 B.n943 10.6151
R1396 B.n943 B.n58 10.6151
R1397 B.n939 B.n58 10.6151
R1398 B.n939 B.n938 10.6151
R1399 B.n938 B.n937 10.6151
R1400 B.n937 B.n60 10.6151
R1401 B.n933 B.n60 10.6151
R1402 B.n933 B.n932 10.6151
R1403 B.n932 B.n931 10.6151
R1404 B.n931 B.n62 10.6151
R1405 B.n927 B.n62 10.6151
R1406 B.n927 B.n926 10.6151
R1407 B.n926 B.n925 10.6151
R1408 B.n925 B.n64 10.6151
R1409 B.n921 B.n64 10.6151
R1410 B.n921 B.n920 10.6151
R1411 B.n920 B.n919 10.6151
R1412 B.n919 B.n66 10.6151
R1413 B.n915 B.n66 10.6151
R1414 B.n915 B.n914 10.6151
R1415 B.n914 B.n913 10.6151
R1416 B.n910 B.n909 10.6151
R1417 B.n909 B.n908 10.6151
R1418 B.n908 B.n72 10.6151
R1419 B.n904 B.n72 10.6151
R1420 B.n904 B.n903 10.6151
R1421 B.n903 B.n902 10.6151
R1422 B.n902 B.n74 10.6151
R1423 B.n898 B.n74 10.6151
R1424 B.n898 B.n897 10.6151
R1425 B.n895 B.n78 10.6151
R1426 B.n891 B.n78 10.6151
R1427 B.n891 B.n890 10.6151
R1428 B.n890 B.n889 10.6151
R1429 B.n889 B.n80 10.6151
R1430 B.n885 B.n80 10.6151
R1431 B.n885 B.n884 10.6151
R1432 B.n884 B.n883 10.6151
R1433 B.n883 B.n82 10.6151
R1434 B.n879 B.n82 10.6151
R1435 B.n879 B.n878 10.6151
R1436 B.n878 B.n877 10.6151
R1437 B.n877 B.n84 10.6151
R1438 B.n873 B.n84 10.6151
R1439 B.n873 B.n872 10.6151
R1440 B.n872 B.n871 10.6151
R1441 B.n871 B.n86 10.6151
R1442 B.n867 B.n86 10.6151
R1443 B.n867 B.n866 10.6151
R1444 B.n866 B.n865 10.6151
R1445 B.n865 B.n88 10.6151
R1446 B.n861 B.n88 10.6151
R1447 B.n861 B.n860 10.6151
R1448 B.n860 B.n859 10.6151
R1449 B.n859 B.n90 10.6151
R1450 B.n855 B.n90 10.6151
R1451 B.n855 B.n854 10.6151
R1452 B.n854 B.n853 10.6151
R1453 B.n853 B.n92 10.6151
R1454 B.n849 B.n92 10.6151
R1455 B.n849 B.n848 10.6151
R1456 B.n848 B.n847 10.6151
R1457 B.n847 B.n94 10.6151
R1458 B.n843 B.n94 10.6151
R1459 B.n843 B.n842 10.6151
R1460 B.n842 B.n841 10.6151
R1461 B.n841 B.n96 10.6151
R1462 B.n837 B.n96 10.6151
R1463 B.n837 B.n836 10.6151
R1464 B.n836 B.n835 10.6151
R1465 B.n835 B.n98 10.6151
R1466 B.n831 B.n98 10.6151
R1467 B.n831 B.n830 10.6151
R1468 B.n830 B.n829 10.6151
R1469 B.n829 B.n100 10.6151
R1470 B.n825 B.n100 10.6151
R1471 B.n825 B.n824 10.6151
R1472 B.n824 B.n823 10.6151
R1473 B.n823 B.n102 10.6151
R1474 B.n819 B.n102 10.6151
R1475 B.n819 B.n818 10.6151
R1476 B.n818 B.n817 10.6151
R1477 B.n817 B.n104 10.6151
R1478 B.n813 B.n104 10.6151
R1479 B.n813 B.n812 10.6151
R1480 B.n812 B.n811 10.6151
R1481 B.n811 B.n106 10.6151
R1482 B.n807 B.n106 10.6151
R1483 B.n807 B.n806 10.6151
R1484 B.n806 B.n805 10.6151
R1485 B.n591 B.n590 10.6151
R1486 B.n591 B.n178 10.6151
R1487 B.n595 B.n178 10.6151
R1488 B.n596 B.n595 10.6151
R1489 B.n597 B.n596 10.6151
R1490 B.n597 B.n176 10.6151
R1491 B.n601 B.n176 10.6151
R1492 B.n602 B.n601 10.6151
R1493 B.n603 B.n602 10.6151
R1494 B.n603 B.n174 10.6151
R1495 B.n607 B.n174 10.6151
R1496 B.n608 B.n607 10.6151
R1497 B.n609 B.n608 10.6151
R1498 B.n609 B.n172 10.6151
R1499 B.n613 B.n172 10.6151
R1500 B.n614 B.n613 10.6151
R1501 B.n615 B.n614 10.6151
R1502 B.n615 B.n170 10.6151
R1503 B.n619 B.n170 10.6151
R1504 B.n620 B.n619 10.6151
R1505 B.n621 B.n620 10.6151
R1506 B.n621 B.n168 10.6151
R1507 B.n625 B.n168 10.6151
R1508 B.n626 B.n625 10.6151
R1509 B.n627 B.n626 10.6151
R1510 B.n627 B.n166 10.6151
R1511 B.n631 B.n166 10.6151
R1512 B.n632 B.n631 10.6151
R1513 B.n633 B.n632 10.6151
R1514 B.n633 B.n164 10.6151
R1515 B.n637 B.n164 10.6151
R1516 B.n638 B.n637 10.6151
R1517 B.n639 B.n638 10.6151
R1518 B.n639 B.n162 10.6151
R1519 B.n643 B.n162 10.6151
R1520 B.n644 B.n643 10.6151
R1521 B.n645 B.n644 10.6151
R1522 B.n645 B.n160 10.6151
R1523 B.n649 B.n160 10.6151
R1524 B.n650 B.n649 10.6151
R1525 B.n651 B.n650 10.6151
R1526 B.n651 B.n158 10.6151
R1527 B.n655 B.n158 10.6151
R1528 B.n656 B.n655 10.6151
R1529 B.n657 B.n656 10.6151
R1530 B.n657 B.n156 10.6151
R1531 B.n661 B.n156 10.6151
R1532 B.n662 B.n661 10.6151
R1533 B.n663 B.n662 10.6151
R1534 B.n663 B.n154 10.6151
R1535 B.n667 B.n154 10.6151
R1536 B.n668 B.n667 10.6151
R1537 B.n669 B.n668 10.6151
R1538 B.n669 B.n152 10.6151
R1539 B.n673 B.n152 10.6151
R1540 B.n674 B.n673 10.6151
R1541 B.n675 B.n674 10.6151
R1542 B.n675 B.n150 10.6151
R1543 B.n679 B.n150 10.6151
R1544 B.n680 B.n679 10.6151
R1545 B.n681 B.n680 10.6151
R1546 B.n681 B.n148 10.6151
R1547 B.n685 B.n148 10.6151
R1548 B.n686 B.n685 10.6151
R1549 B.n687 B.n686 10.6151
R1550 B.n687 B.n146 10.6151
R1551 B.n691 B.n146 10.6151
R1552 B.n692 B.n691 10.6151
R1553 B.n693 B.n692 10.6151
R1554 B.n693 B.n144 10.6151
R1555 B.n697 B.n144 10.6151
R1556 B.n698 B.n697 10.6151
R1557 B.n699 B.n698 10.6151
R1558 B.n699 B.n142 10.6151
R1559 B.n703 B.n142 10.6151
R1560 B.n704 B.n703 10.6151
R1561 B.n705 B.n704 10.6151
R1562 B.n705 B.n140 10.6151
R1563 B.n709 B.n140 10.6151
R1564 B.n710 B.n709 10.6151
R1565 B.n711 B.n710 10.6151
R1566 B.n711 B.n138 10.6151
R1567 B.n715 B.n138 10.6151
R1568 B.n716 B.n715 10.6151
R1569 B.n717 B.n716 10.6151
R1570 B.n717 B.n136 10.6151
R1571 B.n721 B.n136 10.6151
R1572 B.n722 B.n721 10.6151
R1573 B.n723 B.n722 10.6151
R1574 B.n723 B.n134 10.6151
R1575 B.n727 B.n134 10.6151
R1576 B.n728 B.n727 10.6151
R1577 B.n729 B.n728 10.6151
R1578 B.n729 B.n132 10.6151
R1579 B.n733 B.n132 10.6151
R1580 B.n734 B.n733 10.6151
R1581 B.n735 B.n734 10.6151
R1582 B.n735 B.n130 10.6151
R1583 B.n739 B.n130 10.6151
R1584 B.n740 B.n739 10.6151
R1585 B.n741 B.n740 10.6151
R1586 B.n741 B.n128 10.6151
R1587 B.n745 B.n128 10.6151
R1588 B.n746 B.n745 10.6151
R1589 B.n747 B.n746 10.6151
R1590 B.n747 B.n126 10.6151
R1591 B.n751 B.n126 10.6151
R1592 B.n752 B.n751 10.6151
R1593 B.n753 B.n752 10.6151
R1594 B.n753 B.n124 10.6151
R1595 B.n757 B.n124 10.6151
R1596 B.n758 B.n757 10.6151
R1597 B.n759 B.n758 10.6151
R1598 B.n759 B.n122 10.6151
R1599 B.n763 B.n122 10.6151
R1600 B.n764 B.n763 10.6151
R1601 B.n765 B.n764 10.6151
R1602 B.n765 B.n120 10.6151
R1603 B.n769 B.n120 10.6151
R1604 B.n770 B.n769 10.6151
R1605 B.n771 B.n770 10.6151
R1606 B.n771 B.n118 10.6151
R1607 B.n775 B.n118 10.6151
R1608 B.n776 B.n775 10.6151
R1609 B.n777 B.n776 10.6151
R1610 B.n777 B.n116 10.6151
R1611 B.n781 B.n116 10.6151
R1612 B.n782 B.n781 10.6151
R1613 B.n783 B.n782 10.6151
R1614 B.n783 B.n114 10.6151
R1615 B.n787 B.n114 10.6151
R1616 B.n788 B.n787 10.6151
R1617 B.n789 B.n788 10.6151
R1618 B.n789 B.n112 10.6151
R1619 B.n793 B.n112 10.6151
R1620 B.n794 B.n793 10.6151
R1621 B.n795 B.n794 10.6151
R1622 B.n795 B.n110 10.6151
R1623 B.n799 B.n110 10.6151
R1624 B.n800 B.n799 10.6151
R1625 B.n801 B.n800 10.6151
R1626 B.n801 B.n108 10.6151
R1627 B.n392 B.n391 10.6151
R1628 B.n393 B.n392 10.6151
R1629 B.n393 B.n248 10.6151
R1630 B.n397 B.n248 10.6151
R1631 B.n398 B.n397 10.6151
R1632 B.n399 B.n398 10.6151
R1633 B.n399 B.n246 10.6151
R1634 B.n403 B.n246 10.6151
R1635 B.n404 B.n403 10.6151
R1636 B.n405 B.n404 10.6151
R1637 B.n405 B.n244 10.6151
R1638 B.n409 B.n244 10.6151
R1639 B.n410 B.n409 10.6151
R1640 B.n411 B.n410 10.6151
R1641 B.n411 B.n242 10.6151
R1642 B.n415 B.n242 10.6151
R1643 B.n416 B.n415 10.6151
R1644 B.n417 B.n416 10.6151
R1645 B.n417 B.n240 10.6151
R1646 B.n421 B.n240 10.6151
R1647 B.n422 B.n421 10.6151
R1648 B.n423 B.n422 10.6151
R1649 B.n423 B.n238 10.6151
R1650 B.n427 B.n238 10.6151
R1651 B.n428 B.n427 10.6151
R1652 B.n429 B.n428 10.6151
R1653 B.n429 B.n236 10.6151
R1654 B.n433 B.n236 10.6151
R1655 B.n434 B.n433 10.6151
R1656 B.n435 B.n434 10.6151
R1657 B.n435 B.n234 10.6151
R1658 B.n439 B.n234 10.6151
R1659 B.n440 B.n439 10.6151
R1660 B.n441 B.n440 10.6151
R1661 B.n441 B.n232 10.6151
R1662 B.n445 B.n232 10.6151
R1663 B.n446 B.n445 10.6151
R1664 B.n447 B.n446 10.6151
R1665 B.n447 B.n230 10.6151
R1666 B.n451 B.n230 10.6151
R1667 B.n452 B.n451 10.6151
R1668 B.n453 B.n452 10.6151
R1669 B.n453 B.n228 10.6151
R1670 B.n457 B.n228 10.6151
R1671 B.n458 B.n457 10.6151
R1672 B.n459 B.n458 10.6151
R1673 B.n459 B.n226 10.6151
R1674 B.n463 B.n226 10.6151
R1675 B.n464 B.n463 10.6151
R1676 B.n465 B.n464 10.6151
R1677 B.n465 B.n224 10.6151
R1678 B.n469 B.n224 10.6151
R1679 B.n470 B.n469 10.6151
R1680 B.n471 B.n470 10.6151
R1681 B.n471 B.n222 10.6151
R1682 B.n475 B.n222 10.6151
R1683 B.n476 B.n475 10.6151
R1684 B.n477 B.n476 10.6151
R1685 B.n477 B.n220 10.6151
R1686 B.n481 B.n220 10.6151
R1687 B.n484 B.n483 10.6151
R1688 B.n484 B.n216 10.6151
R1689 B.n488 B.n216 10.6151
R1690 B.n489 B.n488 10.6151
R1691 B.n490 B.n489 10.6151
R1692 B.n490 B.n214 10.6151
R1693 B.n494 B.n214 10.6151
R1694 B.n495 B.n494 10.6151
R1695 B.n496 B.n495 10.6151
R1696 B.n500 B.n499 10.6151
R1697 B.n501 B.n500 10.6151
R1698 B.n501 B.n208 10.6151
R1699 B.n505 B.n208 10.6151
R1700 B.n506 B.n505 10.6151
R1701 B.n507 B.n506 10.6151
R1702 B.n507 B.n206 10.6151
R1703 B.n511 B.n206 10.6151
R1704 B.n512 B.n511 10.6151
R1705 B.n513 B.n512 10.6151
R1706 B.n513 B.n204 10.6151
R1707 B.n517 B.n204 10.6151
R1708 B.n518 B.n517 10.6151
R1709 B.n519 B.n518 10.6151
R1710 B.n519 B.n202 10.6151
R1711 B.n523 B.n202 10.6151
R1712 B.n524 B.n523 10.6151
R1713 B.n525 B.n524 10.6151
R1714 B.n525 B.n200 10.6151
R1715 B.n529 B.n200 10.6151
R1716 B.n530 B.n529 10.6151
R1717 B.n531 B.n530 10.6151
R1718 B.n531 B.n198 10.6151
R1719 B.n535 B.n198 10.6151
R1720 B.n536 B.n535 10.6151
R1721 B.n537 B.n536 10.6151
R1722 B.n537 B.n196 10.6151
R1723 B.n541 B.n196 10.6151
R1724 B.n542 B.n541 10.6151
R1725 B.n543 B.n542 10.6151
R1726 B.n543 B.n194 10.6151
R1727 B.n547 B.n194 10.6151
R1728 B.n548 B.n547 10.6151
R1729 B.n549 B.n548 10.6151
R1730 B.n549 B.n192 10.6151
R1731 B.n553 B.n192 10.6151
R1732 B.n554 B.n553 10.6151
R1733 B.n555 B.n554 10.6151
R1734 B.n555 B.n190 10.6151
R1735 B.n559 B.n190 10.6151
R1736 B.n560 B.n559 10.6151
R1737 B.n561 B.n560 10.6151
R1738 B.n561 B.n188 10.6151
R1739 B.n565 B.n188 10.6151
R1740 B.n566 B.n565 10.6151
R1741 B.n567 B.n566 10.6151
R1742 B.n567 B.n186 10.6151
R1743 B.n571 B.n186 10.6151
R1744 B.n572 B.n571 10.6151
R1745 B.n573 B.n572 10.6151
R1746 B.n573 B.n184 10.6151
R1747 B.n577 B.n184 10.6151
R1748 B.n578 B.n577 10.6151
R1749 B.n579 B.n578 10.6151
R1750 B.n579 B.n182 10.6151
R1751 B.n583 B.n182 10.6151
R1752 B.n584 B.n583 10.6151
R1753 B.n585 B.n584 10.6151
R1754 B.n585 B.n180 10.6151
R1755 B.n589 B.n180 10.6151
R1756 B.n387 B.n250 10.6151
R1757 B.n387 B.n386 10.6151
R1758 B.n386 B.n385 10.6151
R1759 B.n385 B.n252 10.6151
R1760 B.n381 B.n252 10.6151
R1761 B.n381 B.n380 10.6151
R1762 B.n380 B.n379 10.6151
R1763 B.n379 B.n254 10.6151
R1764 B.n375 B.n254 10.6151
R1765 B.n375 B.n374 10.6151
R1766 B.n374 B.n373 10.6151
R1767 B.n373 B.n256 10.6151
R1768 B.n369 B.n256 10.6151
R1769 B.n369 B.n368 10.6151
R1770 B.n368 B.n367 10.6151
R1771 B.n367 B.n258 10.6151
R1772 B.n363 B.n258 10.6151
R1773 B.n363 B.n362 10.6151
R1774 B.n362 B.n361 10.6151
R1775 B.n361 B.n260 10.6151
R1776 B.n357 B.n260 10.6151
R1777 B.n357 B.n356 10.6151
R1778 B.n356 B.n355 10.6151
R1779 B.n355 B.n262 10.6151
R1780 B.n351 B.n262 10.6151
R1781 B.n351 B.n350 10.6151
R1782 B.n350 B.n349 10.6151
R1783 B.n349 B.n264 10.6151
R1784 B.n345 B.n264 10.6151
R1785 B.n345 B.n344 10.6151
R1786 B.n344 B.n343 10.6151
R1787 B.n343 B.n266 10.6151
R1788 B.n339 B.n266 10.6151
R1789 B.n339 B.n338 10.6151
R1790 B.n338 B.n337 10.6151
R1791 B.n337 B.n268 10.6151
R1792 B.n333 B.n268 10.6151
R1793 B.n333 B.n332 10.6151
R1794 B.n332 B.n331 10.6151
R1795 B.n331 B.n270 10.6151
R1796 B.n327 B.n270 10.6151
R1797 B.n327 B.n326 10.6151
R1798 B.n326 B.n325 10.6151
R1799 B.n325 B.n272 10.6151
R1800 B.n321 B.n272 10.6151
R1801 B.n321 B.n320 10.6151
R1802 B.n320 B.n319 10.6151
R1803 B.n319 B.n274 10.6151
R1804 B.n315 B.n274 10.6151
R1805 B.n315 B.n314 10.6151
R1806 B.n314 B.n313 10.6151
R1807 B.n313 B.n276 10.6151
R1808 B.n309 B.n276 10.6151
R1809 B.n309 B.n308 10.6151
R1810 B.n308 B.n307 10.6151
R1811 B.n307 B.n278 10.6151
R1812 B.n303 B.n278 10.6151
R1813 B.n303 B.n302 10.6151
R1814 B.n302 B.n301 10.6151
R1815 B.n301 B.n280 10.6151
R1816 B.n297 B.n280 10.6151
R1817 B.n297 B.n296 10.6151
R1818 B.n296 B.n295 10.6151
R1819 B.n295 B.n282 10.6151
R1820 B.n291 B.n282 10.6151
R1821 B.n291 B.n290 10.6151
R1822 B.n290 B.n289 10.6151
R1823 B.n289 B.n284 10.6151
R1824 B.n285 B.n284 10.6151
R1825 B.n285 B.n0 10.6151
R1826 B.n1107 B.n1 10.6151
R1827 B.n1107 B.n1106 10.6151
R1828 B.n1106 B.n1105 10.6151
R1829 B.n1105 B.n4 10.6151
R1830 B.n1101 B.n4 10.6151
R1831 B.n1101 B.n1100 10.6151
R1832 B.n1100 B.n1099 10.6151
R1833 B.n1099 B.n6 10.6151
R1834 B.n1095 B.n6 10.6151
R1835 B.n1095 B.n1094 10.6151
R1836 B.n1094 B.n1093 10.6151
R1837 B.n1093 B.n8 10.6151
R1838 B.n1089 B.n8 10.6151
R1839 B.n1089 B.n1088 10.6151
R1840 B.n1088 B.n1087 10.6151
R1841 B.n1087 B.n10 10.6151
R1842 B.n1083 B.n10 10.6151
R1843 B.n1083 B.n1082 10.6151
R1844 B.n1082 B.n1081 10.6151
R1845 B.n1081 B.n12 10.6151
R1846 B.n1077 B.n12 10.6151
R1847 B.n1077 B.n1076 10.6151
R1848 B.n1076 B.n1075 10.6151
R1849 B.n1075 B.n14 10.6151
R1850 B.n1071 B.n14 10.6151
R1851 B.n1071 B.n1070 10.6151
R1852 B.n1070 B.n1069 10.6151
R1853 B.n1069 B.n16 10.6151
R1854 B.n1065 B.n16 10.6151
R1855 B.n1065 B.n1064 10.6151
R1856 B.n1064 B.n1063 10.6151
R1857 B.n1063 B.n18 10.6151
R1858 B.n1059 B.n18 10.6151
R1859 B.n1059 B.n1058 10.6151
R1860 B.n1058 B.n1057 10.6151
R1861 B.n1057 B.n20 10.6151
R1862 B.n1053 B.n20 10.6151
R1863 B.n1053 B.n1052 10.6151
R1864 B.n1052 B.n1051 10.6151
R1865 B.n1051 B.n22 10.6151
R1866 B.n1047 B.n22 10.6151
R1867 B.n1047 B.n1046 10.6151
R1868 B.n1046 B.n1045 10.6151
R1869 B.n1045 B.n24 10.6151
R1870 B.n1041 B.n24 10.6151
R1871 B.n1041 B.n1040 10.6151
R1872 B.n1040 B.n1039 10.6151
R1873 B.n1039 B.n26 10.6151
R1874 B.n1035 B.n26 10.6151
R1875 B.n1035 B.n1034 10.6151
R1876 B.n1034 B.n1033 10.6151
R1877 B.n1033 B.n28 10.6151
R1878 B.n1029 B.n28 10.6151
R1879 B.n1029 B.n1028 10.6151
R1880 B.n1028 B.n1027 10.6151
R1881 B.n1027 B.n30 10.6151
R1882 B.n1023 B.n30 10.6151
R1883 B.n1023 B.n1022 10.6151
R1884 B.n1022 B.n1021 10.6151
R1885 B.n1021 B.n32 10.6151
R1886 B.n1017 B.n32 10.6151
R1887 B.n1017 B.n1016 10.6151
R1888 B.n1016 B.n1015 10.6151
R1889 B.n1015 B.n34 10.6151
R1890 B.n1011 B.n34 10.6151
R1891 B.n1011 B.n1010 10.6151
R1892 B.n1010 B.n1009 10.6151
R1893 B.n1009 B.n36 10.6151
R1894 B.n1005 B.n36 10.6151
R1895 B.n1005 B.n1004 10.6151
R1896 B.n913 B.n70 9.36635
R1897 B.n896 B.n895 9.36635
R1898 B.n482 B.n481 9.36635
R1899 B.n499 B.n212 9.36635
R1900 B.n1111 B.n0 2.81026
R1901 B.n1111 B.n1 2.81026
R1902 B.n910 B.n70 1.24928
R1903 B.n897 B.n896 1.24928
R1904 B.n483 B.n482 1.24928
R1905 B.n496 B.n212 1.24928
R1906 VN.n61 VN.t3 171.821
R1907 VN.n13 VN.t8 171.821
R1908 VN.n94 VN.n93 161.3
R1909 VN.n92 VN.n49 161.3
R1910 VN.n91 VN.n90 161.3
R1911 VN.n89 VN.n50 161.3
R1912 VN.n88 VN.n87 161.3
R1913 VN.n86 VN.n51 161.3
R1914 VN.n85 VN.n84 161.3
R1915 VN.n83 VN.n82 161.3
R1916 VN.n81 VN.n53 161.3
R1917 VN.n80 VN.n79 161.3
R1918 VN.n78 VN.n54 161.3
R1919 VN.n77 VN.n76 161.3
R1920 VN.n75 VN.n55 161.3
R1921 VN.n74 VN.n73 161.3
R1922 VN.n72 VN.n71 161.3
R1923 VN.n70 VN.n57 161.3
R1924 VN.n69 VN.n68 161.3
R1925 VN.n67 VN.n58 161.3
R1926 VN.n66 VN.n65 161.3
R1927 VN.n64 VN.n59 161.3
R1928 VN.n63 VN.n62 161.3
R1929 VN.n46 VN.n45 161.3
R1930 VN.n44 VN.n1 161.3
R1931 VN.n43 VN.n42 161.3
R1932 VN.n41 VN.n2 161.3
R1933 VN.n40 VN.n39 161.3
R1934 VN.n38 VN.n3 161.3
R1935 VN.n37 VN.n36 161.3
R1936 VN.n35 VN.n34 161.3
R1937 VN.n33 VN.n5 161.3
R1938 VN.n32 VN.n31 161.3
R1939 VN.n30 VN.n6 161.3
R1940 VN.n29 VN.n28 161.3
R1941 VN.n27 VN.n7 161.3
R1942 VN.n26 VN.n25 161.3
R1943 VN.n24 VN.n23 161.3
R1944 VN.n22 VN.n9 161.3
R1945 VN.n21 VN.n20 161.3
R1946 VN.n19 VN.n10 161.3
R1947 VN.n18 VN.n17 161.3
R1948 VN.n16 VN.n11 161.3
R1949 VN.n15 VN.n14 161.3
R1950 VN.n12 VN.t5 138.371
R1951 VN.n8 VN.t4 138.371
R1952 VN.n4 VN.t7 138.371
R1953 VN.n0 VN.t6 138.371
R1954 VN.n60 VN.t1 138.371
R1955 VN.n56 VN.t9 138.371
R1956 VN.n52 VN.t2 138.371
R1957 VN.n48 VN.t0 138.371
R1958 VN.n47 VN.n0 70.0803
R1959 VN.n95 VN.n48 70.0803
R1960 VN VN.n95 62.0436
R1961 VN.n13 VN.n12 58.1015
R1962 VN.n61 VN.n60 58.1015
R1963 VN.n43 VN.n2 52.2023
R1964 VN.n91 VN.n50 52.2023
R1965 VN.n17 VN.n10 44.4521
R1966 VN.n32 VN.n6 44.4521
R1967 VN.n65 VN.n58 44.4521
R1968 VN.n80 VN.n54 44.4521
R1969 VN.n21 VN.n10 36.702
R1970 VN.n28 VN.n6 36.702
R1971 VN.n69 VN.n58 36.702
R1972 VN.n76 VN.n54 36.702
R1973 VN.n39 VN.n2 28.9518
R1974 VN.n87 VN.n50 28.9518
R1975 VN.n16 VN.n15 24.5923
R1976 VN.n17 VN.n16 24.5923
R1977 VN.n22 VN.n21 24.5923
R1978 VN.n23 VN.n22 24.5923
R1979 VN.n27 VN.n26 24.5923
R1980 VN.n28 VN.n27 24.5923
R1981 VN.n33 VN.n32 24.5923
R1982 VN.n34 VN.n33 24.5923
R1983 VN.n38 VN.n37 24.5923
R1984 VN.n39 VN.n38 24.5923
R1985 VN.n44 VN.n43 24.5923
R1986 VN.n45 VN.n44 24.5923
R1987 VN.n65 VN.n64 24.5923
R1988 VN.n64 VN.n63 24.5923
R1989 VN.n76 VN.n75 24.5923
R1990 VN.n75 VN.n74 24.5923
R1991 VN.n71 VN.n70 24.5923
R1992 VN.n70 VN.n69 24.5923
R1993 VN.n87 VN.n86 24.5923
R1994 VN.n86 VN.n85 24.5923
R1995 VN.n82 VN.n81 24.5923
R1996 VN.n81 VN.n80 24.5923
R1997 VN.n93 VN.n92 24.5923
R1998 VN.n92 VN.n91 24.5923
R1999 VN.n45 VN.n0 20.1658
R2000 VN.n93 VN.n48 20.1658
R2001 VN.n15 VN.n12 16.2311
R2002 VN.n34 VN.n4 16.2311
R2003 VN.n63 VN.n60 16.2311
R2004 VN.n82 VN.n52 16.2311
R2005 VN.n23 VN.n8 12.2964
R2006 VN.n26 VN.n8 12.2964
R2007 VN.n74 VN.n56 12.2964
R2008 VN.n71 VN.n56 12.2964
R2009 VN.n37 VN.n4 8.36172
R2010 VN.n85 VN.n52 8.36172
R2011 VN.n14 VN.n13 3.88977
R2012 VN.n62 VN.n61 3.88977
R2013 VN.n95 VN.n94 0.354861
R2014 VN.n47 VN.n46 0.354861
R2015 VN VN.n47 0.267071
R2016 VN.n94 VN.n49 0.189894
R2017 VN.n90 VN.n49 0.189894
R2018 VN.n90 VN.n89 0.189894
R2019 VN.n89 VN.n88 0.189894
R2020 VN.n88 VN.n51 0.189894
R2021 VN.n84 VN.n51 0.189894
R2022 VN.n84 VN.n83 0.189894
R2023 VN.n83 VN.n53 0.189894
R2024 VN.n79 VN.n53 0.189894
R2025 VN.n79 VN.n78 0.189894
R2026 VN.n78 VN.n77 0.189894
R2027 VN.n77 VN.n55 0.189894
R2028 VN.n73 VN.n55 0.189894
R2029 VN.n73 VN.n72 0.189894
R2030 VN.n72 VN.n57 0.189894
R2031 VN.n68 VN.n57 0.189894
R2032 VN.n68 VN.n67 0.189894
R2033 VN.n67 VN.n66 0.189894
R2034 VN.n66 VN.n59 0.189894
R2035 VN.n62 VN.n59 0.189894
R2036 VN.n14 VN.n11 0.189894
R2037 VN.n18 VN.n11 0.189894
R2038 VN.n19 VN.n18 0.189894
R2039 VN.n20 VN.n19 0.189894
R2040 VN.n20 VN.n9 0.189894
R2041 VN.n24 VN.n9 0.189894
R2042 VN.n25 VN.n24 0.189894
R2043 VN.n25 VN.n7 0.189894
R2044 VN.n29 VN.n7 0.189894
R2045 VN.n30 VN.n29 0.189894
R2046 VN.n31 VN.n30 0.189894
R2047 VN.n31 VN.n5 0.189894
R2048 VN.n35 VN.n5 0.189894
R2049 VN.n36 VN.n35 0.189894
R2050 VN.n36 VN.n3 0.189894
R2051 VN.n40 VN.n3 0.189894
R2052 VN.n41 VN.n40 0.189894
R2053 VN.n42 VN.n41 0.189894
R2054 VN.n42 VN.n1 0.189894
R2055 VN.n46 VN.n1 0.189894
R2056 VDD2.n1 VDD2.t1 74.5241
R2057 VDD2.n3 VDD2.n2 71.9552
R2058 VDD2 VDD2.n7 71.9524
R2059 VDD2.n4 VDD2.t9 71.4381
R2060 VDD2.n6 VDD2.n5 69.6962
R2061 VDD2.n1 VDD2.n0 69.6959
R2062 VDD2.n4 VDD2.n3 54.461
R2063 VDD2.n6 VDD2.n4 3.08671
R2064 VDD2.n7 VDD2.t8 1.74246
R2065 VDD2.n7 VDD2.t6 1.74246
R2066 VDD2.n5 VDD2.t7 1.74246
R2067 VDD2.n5 VDD2.t0 1.74246
R2068 VDD2.n2 VDD2.t2 1.74246
R2069 VDD2.n2 VDD2.t3 1.74246
R2070 VDD2.n0 VDD2.t4 1.74246
R2071 VDD2.n0 VDD2.t5 1.74246
R2072 VDD2 VDD2.n6 0.830241
R2073 VDD2.n3 VDD2.n1 0.716706
C0 VDD1 B 3.26721f
C1 VN B 1.53126f
C2 VTAIL VP 17.606302f
C3 w_n5266_n4700# VP 12.2553f
C4 w_n5266_n4700# VTAIL 4.20802f
C5 VDD2 VDD1 2.59735f
C6 VDD2 VN 16.979301f
C7 VP B 2.6911f
C8 VTAIL B 5.537f
C9 w_n5266_n4700# B 13.5069f
C10 VN VDD1 0.155031f
C11 VDD2 VP 0.667138f
C12 VDD2 VTAIL 13.467501f
C13 w_n5266_n4700# VDD2 3.66803f
C14 VP VDD1 17.486599f
C15 VTAIL VDD1 13.4128f
C16 VDD2 B 3.41044f
C17 VN VP 10.580299f
C18 VTAIL VN 17.592001f
C19 w_n5266_n4700# VDD1 3.4907f
C20 w_n5266_n4700# VN 11.5677f
C21 VDD2 VSUBS 2.53586f
C22 VDD1 VSUBS 2.397904f
C23 VTAIL VSUBS 1.686384f
C24 VN VSUBS 8.99858f
C25 VP VSUBS 5.316225f
C26 B VSUBS 6.734859f
C27 w_n5266_n4700# VSUBS 0.3025p
C28 VDD2.t1 VSUBS 4.62185f
C29 VDD2.t4 VSUBS 0.422817f
C30 VDD2.t5 VSUBS 0.422817f
C31 VDD2.n0 VSUBS 3.53275f
C32 VDD2.n1 VSUBS 1.83973f
C33 VDD2.t2 VSUBS 0.422817f
C34 VDD2.t3 VSUBS 0.422817f
C35 VDD2.n2 VSUBS 3.56632f
C36 VDD2.n3 VSUBS 4.52111f
C37 VDD2.t9 VSUBS 4.58195f
C38 VDD2.n4 VSUBS 4.80937f
C39 VDD2.t7 VSUBS 0.422817f
C40 VDD2.t0 VSUBS 0.422817f
C41 VDD2.n5 VSUBS 3.53276f
C42 VDD2.n6 VSUBS 0.925177f
C43 VDD2.t8 VSUBS 0.422817f
C44 VDD2.t6 VSUBS 0.422817f
C45 VDD2.n7 VSUBS 3.56625f
C46 VN.t6 VSUBS 3.68281f
C47 VN.n0 VSUBS 1.36323f
C48 VN.n1 VSUBS 0.022063f
C49 VN.n2 VSUBS 0.022232f
C50 VN.n3 VSUBS 0.022063f
C51 VN.t7 VSUBS 3.68281f
C52 VN.n4 VSUBS 1.27013f
C53 VN.n5 VSUBS 0.022063f
C54 VN.n6 VSUBS 0.018274f
C55 VN.n7 VSUBS 0.022063f
C56 VN.t4 VSUBS 3.68281f
C57 VN.n8 VSUBS 1.27013f
C58 VN.n9 VSUBS 0.022063f
C59 VN.n10 VSUBS 0.018274f
C60 VN.n11 VSUBS 0.022063f
C61 VN.t5 VSUBS 3.68281f
C62 VN.n12 VSUBS 1.34586f
C63 VN.t8 VSUBS 3.96136f
C64 VN.n13 VSUBS 1.29209f
C65 VN.n14 VSUBS 0.255165f
C66 VN.n15 VSUBS 0.034047f
C67 VN.n16 VSUBS 0.040915f
C68 VN.n17 VSUBS 0.042539f
C69 VN.n18 VSUBS 0.022063f
C70 VN.n19 VSUBS 0.022063f
C71 VN.n20 VSUBS 0.022063f
C72 VN.n21 VSUBS 0.044247f
C73 VN.n22 VSUBS 0.040915f
C74 VN.n23 VSUBS 0.030815f
C75 VN.n24 VSUBS 0.022063f
C76 VN.n25 VSUBS 0.022063f
C77 VN.n26 VSUBS 0.030815f
C78 VN.n27 VSUBS 0.040915f
C79 VN.n28 VSUBS 0.044247f
C80 VN.n29 VSUBS 0.022063f
C81 VN.n30 VSUBS 0.022063f
C82 VN.n31 VSUBS 0.022063f
C83 VN.n32 VSUBS 0.042539f
C84 VN.n33 VSUBS 0.040915f
C85 VN.n34 VSUBS 0.034047f
C86 VN.n35 VSUBS 0.022063f
C87 VN.n36 VSUBS 0.022063f
C88 VN.n37 VSUBS 0.027584f
C89 VN.n38 VSUBS 0.040915f
C90 VN.n39 VSUBS 0.043408f
C91 VN.n40 VSUBS 0.022063f
C92 VN.n41 VSUBS 0.022063f
C93 VN.n42 VSUBS 0.022063f
C94 VN.n43 VSUBS 0.039419f
C95 VN.n44 VSUBS 0.040915f
C96 VN.n45 VSUBS 0.037279f
C97 VN.n46 VSUBS 0.035604f
C98 VN.n47 VSUBS 0.047624f
C99 VN.t0 VSUBS 3.68281f
C100 VN.n48 VSUBS 1.36323f
C101 VN.n49 VSUBS 0.022063f
C102 VN.n50 VSUBS 0.022232f
C103 VN.n51 VSUBS 0.022063f
C104 VN.t2 VSUBS 3.68281f
C105 VN.n52 VSUBS 1.27013f
C106 VN.n53 VSUBS 0.022063f
C107 VN.n54 VSUBS 0.018274f
C108 VN.n55 VSUBS 0.022063f
C109 VN.t9 VSUBS 3.68281f
C110 VN.n56 VSUBS 1.27013f
C111 VN.n57 VSUBS 0.022063f
C112 VN.n58 VSUBS 0.018274f
C113 VN.n59 VSUBS 0.022063f
C114 VN.t1 VSUBS 3.68281f
C115 VN.n60 VSUBS 1.34586f
C116 VN.t3 VSUBS 3.96136f
C117 VN.n61 VSUBS 1.29209f
C118 VN.n62 VSUBS 0.255165f
C119 VN.n63 VSUBS 0.034047f
C120 VN.n64 VSUBS 0.040915f
C121 VN.n65 VSUBS 0.042539f
C122 VN.n66 VSUBS 0.022063f
C123 VN.n67 VSUBS 0.022063f
C124 VN.n68 VSUBS 0.022063f
C125 VN.n69 VSUBS 0.044247f
C126 VN.n70 VSUBS 0.040915f
C127 VN.n71 VSUBS 0.030815f
C128 VN.n72 VSUBS 0.022063f
C129 VN.n73 VSUBS 0.022063f
C130 VN.n74 VSUBS 0.030815f
C131 VN.n75 VSUBS 0.040915f
C132 VN.n76 VSUBS 0.044247f
C133 VN.n77 VSUBS 0.022063f
C134 VN.n78 VSUBS 0.022063f
C135 VN.n79 VSUBS 0.022063f
C136 VN.n80 VSUBS 0.042539f
C137 VN.n81 VSUBS 0.040915f
C138 VN.n82 VSUBS 0.034047f
C139 VN.n83 VSUBS 0.022063f
C140 VN.n84 VSUBS 0.022063f
C141 VN.n85 VSUBS 0.027584f
C142 VN.n86 VSUBS 0.040915f
C143 VN.n87 VSUBS 0.043408f
C144 VN.n88 VSUBS 0.022063f
C145 VN.n89 VSUBS 0.022063f
C146 VN.n90 VSUBS 0.022063f
C147 VN.n91 VSUBS 0.039419f
C148 VN.n92 VSUBS 0.040915f
C149 VN.n93 VSUBS 0.037279f
C150 VN.n94 VSUBS 0.035604f
C151 VN.n95 VSUBS 1.68724f
C152 B.n0 VSUBS 0.004861f
C153 B.n1 VSUBS 0.004861f
C154 B.n2 VSUBS 0.007687f
C155 B.n3 VSUBS 0.007687f
C156 B.n4 VSUBS 0.007687f
C157 B.n5 VSUBS 0.007687f
C158 B.n6 VSUBS 0.007687f
C159 B.n7 VSUBS 0.007687f
C160 B.n8 VSUBS 0.007687f
C161 B.n9 VSUBS 0.007687f
C162 B.n10 VSUBS 0.007687f
C163 B.n11 VSUBS 0.007687f
C164 B.n12 VSUBS 0.007687f
C165 B.n13 VSUBS 0.007687f
C166 B.n14 VSUBS 0.007687f
C167 B.n15 VSUBS 0.007687f
C168 B.n16 VSUBS 0.007687f
C169 B.n17 VSUBS 0.007687f
C170 B.n18 VSUBS 0.007687f
C171 B.n19 VSUBS 0.007687f
C172 B.n20 VSUBS 0.007687f
C173 B.n21 VSUBS 0.007687f
C174 B.n22 VSUBS 0.007687f
C175 B.n23 VSUBS 0.007687f
C176 B.n24 VSUBS 0.007687f
C177 B.n25 VSUBS 0.007687f
C178 B.n26 VSUBS 0.007687f
C179 B.n27 VSUBS 0.007687f
C180 B.n28 VSUBS 0.007687f
C181 B.n29 VSUBS 0.007687f
C182 B.n30 VSUBS 0.007687f
C183 B.n31 VSUBS 0.007687f
C184 B.n32 VSUBS 0.007687f
C185 B.n33 VSUBS 0.007687f
C186 B.n34 VSUBS 0.007687f
C187 B.n35 VSUBS 0.007687f
C188 B.n36 VSUBS 0.007687f
C189 B.n37 VSUBS 0.01839f
C190 B.n38 VSUBS 0.007687f
C191 B.n39 VSUBS 0.007687f
C192 B.n40 VSUBS 0.007687f
C193 B.n41 VSUBS 0.007687f
C194 B.n42 VSUBS 0.007687f
C195 B.n43 VSUBS 0.007687f
C196 B.n44 VSUBS 0.007687f
C197 B.n45 VSUBS 0.007687f
C198 B.n46 VSUBS 0.007687f
C199 B.n47 VSUBS 0.007687f
C200 B.n48 VSUBS 0.007687f
C201 B.n49 VSUBS 0.007687f
C202 B.n50 VSUBS 0.007687f
C203 B.n51 VSUBS 0.007687f
C204 B.n52 VSUBS 0.007687f
C205 B.n53 VSUBS 0.007687f
C206 B.n54 VSUBS 0.007687f
C207 B.n55 VSUBS 0.007687f
C208 B.n56 VSUBS 0.007687f
C209 B.n57 VSUBS 0.007687f
C210 B.n58 VSUBS 0.007687f
C211 B.n59 VSUBS 0.007687f
C212 B.n60 VSUBS 0.007687f
C213 B.n61 VSUBS 0.007687f
C214 B.n62 VSUBS 0.007687f
C215 B.n63 VSUBS 0.007687f
C216 B.n64 VSUBS 0.007687f
C217 B.n65 VSUBS 0.007687f
C218 B.n66 VSUBS 0.007687f
C219 B.n67 VSUBS 0.007687f
C220 B.t5 VSUBS 0.693549f
C221 B.t4 VSUBS 0.720801f
C222 B.t3 VSUBS 2.9954f
C223 B.n68 VSUBS 0.431444f
C224 B.n69 VSUBS 0.082153f
C225 B.n70 VSUBS 0.017811f
C226 B.n71 VSUBS 0.007687f
C227 B.n72 VSUBS 0.007687f
C228 B.n73 VSUBS 0.007687f
C229 B.n74 VSUBS 0.007687f
C230 B.n75 VSUBS 0.007687f
C231 B.t2 VSUBS 0.693522f
C232 B.t1 VSUBS 0.720781f
C233 B.t0 VSUBS 2.9954f
C234 B.n76 VSUBS 0.431464f
C235 B.n77 VSUBS 0.082179f
C236 B.n78 VSUBS 0.007687f
C237 B.n79 VSUBS 0.007687f
C238 B.n80 VSUBS 0.007687f
C239 B.n81 VSUBS 0.007687f
C240 B.n82 VSUBS 0.007687f
C241 B.n83 VSUBS 0.007687f
C242 B.n84 VSUBS 0.007687f
C243 B.n85 VSUBS 0.007687f
C244 B.n86 VSUBS 0.007687f
C245 B.n87 VSUBS 0.007687f
C246 B.n88 VSUBS 0.007687f
C247 B.n89 VSUBS 0.007687f
C248 B.n90 VSUBS 0.007687f
C249 B.n91 VSUBS 0.007687f
C250 B.n92 VSUBS 0.007687f
C251 B.n93 VSUBS 0.007687f
C252 B.n94 VSUBS 0.007687f
C253 B.n95 VSUBS 0.007687f
C254 B.n96 VSUBS 0.007687f
C255 B.n97 VSUBS 0.007687f
C256 B.n98 VSUBS 0.007687f
C257 B.n99 VSUBS 0.007687f
C258 B.n100 VSUBS 0.007687f
C259 B.n101 VSUBS 0.007687f
C260 B.n102 VSUBS 0.007687f
C261 B.n103 VSUBS 0.007687f
C262 B.n104 VSUBS 0.007687f
C263 B.n105 VSUBS 0.007687f
C264 B.n106 VSUBS 0.007687f
C265 B.n107 VSUBS 0.007687f
C266 B.n108 VSUBS 0.019227f
C267 B.n109 VSUBS 0.007687f
C268 B.n110 VSUBS 0.007687f
C269 B.n111 VSUBS 0.007687f
C270 B.n112 VSUBS 0.007687f
C271 B.n113 VSUBS 0.007687f
C272 B.n114 VSUBS 0.007687f
C273 B.n115 VSUBS 0.007687f
C274 B.n116 VSUBS 0.007687f
C275 B.n117 VSUBS 0.007687f
C276 B.n118 VSUBS 0.007687f
C277 B.n119 VSUBS 0.007687f
C278 B.n120 VSUBS 0.007687f
C279 B.n121 VSUBS 0.007687f
C280 B.n122 VSUBS 0.007687f
C281 B.n123 VSUBS 0.007687f
C282 B.n124 VSUBS 0.007687f
C283 B.n125 VSUBS 0.007687f
C284 B.n126 VSUBS 0.007687f
C285 B.n127 VSUBS 0.007687f
C286 B.n128 VSUBS 0.007687f
C287 B.n129 VSUBS 0.007687f
C288 B.n130 VSUBS 0.007687f
C289 B.n131 VSUBS 0.007687f
C290 B.n132 VSUBS 0.007687f
C291 B.n133 VSUBS 0.007687f
C292 B.n134 VSUBS 0.007687f
C293 B.n135 VSUBS 0.007687f
C294 B.n136 VSUBS 0.007687f
C295 B.n137 VSUBS 0.007687f
C296 B.n138 VSUBS 0.007687f
C297 B.n139 VSUBS 0.007687f
C298 B.n140 VSUBS 0.007687f
C299 B.n141 VSUBS 0.007687f
C300 B.n142 VSUBS 0.007687f
C301 B.n143 VSUBS 0.007687f
C302 B.n144 VSUBS 0.007687f
C303 B.n145 VSUBS 0.007687f
C304 B.n146 VSUBS 0.007687f
C305 B.n147 VSUBS 0.007687f
C306 B.n148 VSUBS 0.007687f
C307 B.n149 VSUBS 0.007687f
C308 B.n150 VSUBS 0.007687f
C309 B.n151 VSUBS 0.007687f
C310 B.n152 VSUBS 0.007687f
C311 B.n153 VSUBS 0.007687f
C312 B.n154 VSUBS 0.007687f
C313 B.n155 VSUBS 0.007687f
C314 B.n156 VSUBS 0.007687f
C315 B.n157 VSUBS 0.007687f
C316 B.n158 VSUBS 0.007687f
C317 B.n159 VSUBS 0.007687f
C318 B.n160 VSUBS 0.007687f
C319 B.n161 VSUBS 0.007687f
C320 B.n162 VSUBS 0.007687f
C321 B.n163 VSUBS 0.007687f
C322 B.n164 VSUBS 0.007687f
C323 B.n165 VSUBS 0.007687f
C324 B.n166 VSUBS 0.007687f
C325 B.n167 VSUBS 0.007687f
C326 B.n168 VSUBS 0.007687f
C327 B.n169 VSUBS 0.007687f
C328 B.n170 VSUBS 0.007687f
C329 B.n171 VSUBS 0.007687f
C330 B.n172 VSUBS 0.007687f
C331 B.n173 VSUBS 0.007687f
C332 B.n174 VSUBS 0.007687f
C333 B.n175 VSUBS 0.007687f
C334 B.n176 VSUBS 0.007687f
C335 B.n177 VSUBS 0.007687f
C336 B.n178 VSUBS 0.007687f
C337 B.n179 VSUBS 0.01839f
C338 B.n180 VSUBS 0.007687f
C339 B.n181 VSUBS 0.007687f
C340 B.n182 VSUBS 0.007687f
C341 B.n183 VSUBS 0.007687f
C342 B.n184 VSUBS 0.007687f
C343 B.n185 VSUBS 0.007687f
C344 B.n186 VSUBS 0.007687f
C345 B.n187 VSUBS 0.007687f
C346 B.n188 VSUBS 0.007687f
C347 B.n189 VSUBS 0.007687f
C348 B.n190 VSUBS 0.007687f
C349 B.n191 VSUBS 0.007687f
C350 B.n192 VSUBS 0.007687f
C351 B.n193 VSUBS 0.007687f
C352 B.n194 VSUBS 0.007687f
C353 B.n195 VSUBS 0.007687f
C354 B.n196 VSUBS 0.007687f
C355 B.n197 VSUBS 0.007687f
C356 B.n198 VSUBS 0.007687f
C357 B.n199 VSUBS 0.007687f
C358 B.n200 VSUBS 0.007687f
C359 B.n201 VSUBS 0.007687f
C360 B.n202 VSUBS 0.007687f
C361 B.n203 VSUBS 0.007687f
C362 B.n204 VSUBS 0.007687f
C363 B.n205 VSUBS 0.007687f
C364 B.n206 VSUBS 0.007687f
C365 B.n207 VSUBS 0.007687f
C366 B.n208 VSUBS 0.007687f
C367 B.n209 VSUBS 0.007687f
C368 B.t10 VSUBS 0.693522f
C369 B.t11 VSUBS 0.720781f
C370 B.t9 VSUBS 2.9954f
C371 B.n210 VSUBS 0.431464f
C372 B.n211 VSUBS 0.082179f
C373 B.n212 VSUBS 0.017811f
C374 B.n213 VSUBS 0.007687f
C375 B.n214 VSUBS 0.007687f
C376 B.n215 VSUBS 0.007687f
C377 B.n216 VSUBS 0.007687f
C378 B.n217 VSUBS 0.007687f
C379 B.t7 VSUBS 0.693549f
C380 B.t8 VSUBS 0.720801f
C381 B.t6 VSUBS 2.9954f
C382 B.n218 VSUBS 0.431444f
C383 B.n219 VSUBS 0.082153f
C384 B.n220 VSUBS 0.007687f
C385 B.n221 VSUBS 0.007687f
C386 B.n222 VSUBS 0.007687f
C387 B.n223 VSUBS 0.007687f
C388 B.n224 VSUBS 0.007687f
C389 B.n225 VSUBS 0.007687f
C390 B.n226 VSUBS 0.007687f
C391 B.n227 VSUBS 0.007687f
C392 B.n228 VSUBS 0.007687f
C393 B.n229 VSUBS 0.007687f
C394 B.n230 VSUBS 0.007687f
C395 B.n231 VSUBS 0.007687f
C396 B.n232 VSUBS 0.007687f
C397 B.n233 VSUBS 0.007687f
C398 B.n234 VSUBS 0.007687f
C399 B.n235 VSUBS 0.007687f
C400 B.n236 VSUBS 0.007687f
C401 B.n237 VSUBS 0.007687f
C402 B.n238 VSUBS 0.007687f
C403 B.n239 VSUBS 0.007687f
C404 B.n240 VSUBS 0.007687f
C405 B.n241 VSUBS 0.007687f
C406 B.n242 VSUBS 0.007687f
C407 B.n243 VSUBS 0.007687f
C408 B.n244 VSUBS 0.007687f
C409 B.n245 VSUBS 0.007687f
C410 B.n246 VSUBS 0.007687f
C411 B.n247 VSUBS 0.007687f
C412 B.n248 VSUBS 0.007687f
C413 B.n249 VSUBS 0.007687f
C414 B.n250 VSUBS 0.01839f
C415 B.n251 VSUBS 0.007687f
C416 B.n252 VSUBS 0.007687f
C417 B.n253 VSUBS 0.007687f
C418 B.n254 VSUBS 0.007687f
C419 B.n255 VSUBS 0.007687f
C420 B.n256 VSUBS 0.007687f
C421 B.n257 VSUBS 0.007687f
C422 B.n258 VSUBS 0.007687f
C423 B.n259 VSUBS 0.007687f
C424 B.n260 VSUBS 0.007687f
C425 B.n261 VSUBS 0.007687f
C426 B.n262 VSUBS 0.007687f
C427 B.n263 VSUBS 0.007687f
C428 B.n264 VSUBS 0.007687f
C429 B.n265 VSUBS 0.007687f
C430 B.n266 VSUBS 0.007687f
C431 B.n267 VSUBS 0.007687f
C432 B.n268 VSUBS 0.007687f
C433 B.n269 VSUBS 0.007687f
C434 B.n270 VSUBS 0.007687f
C435 B.n271 VSUBS 0.007687f
C436 B.n272 VSUBS 0.007687f
C437 B.n273 VSUBS 0.007687f
C438 B.n274 VSUBS 0.007687f
C439 B.n275 VSUBS 0.007687f
C440 B.n276 VSUBS 0.007687f
C441 B.n277 VSUBS 0.007687f
C442 B.n278 VSUBS 0.007687f
C443 B.n279 VSUBS 0.007687f
C444 B.n280 VSUBS 0.007687f
C445 B.n281 VSUBS 0.007687f
C446 B.n282 VSUBS 0.007687f
C447 B.n283 VSUBS 0.007687f
C448 B.n284 VSUBS 0.007687f
C449 B.n285 VSUBS 0.007687f
C450 B.n286 VSUBS 0.007687f
C451 B.n287 VSUBS 0.007687f
C452 B.n288 VSUBS 0.007687f
C453 B.n289 VSUBS 0.007687f
C454 B.n290 VSUBS 0.007687f
C455 B.n291 VSUBS 0.007687f
C456 B.n292 VSUBS 0.007687f
C457 B.n293 VSUBS 0.007687f
C458 B.n294 VSUBS 0.007687f
C459 B.n295 VSUBS 0.007687f
C460 B.n296 VSUBS 0.007687f
C461 B.n297 VSUBS 0.007687f
C462 B.n298 VSUBS 0.007687f
C463 B.n299 VSUBS 0.007687f
C464 B.n300 VSUBS 0.007687f
C465 B.n301 VSUBS 0.007687f
C466 B.n302 VSUBS 0.007687f
C467 B.n303 VSUBS 0.007687f
C468 B.n304 VSUBS 0.007687f
C469 B.n305 VSUBS 0.007687f
C470 B.n306 VSUBS 0.007687f
C471 B.n307 VSUBS 0.007687f
C472 B.n308 VSUBS 0.007687f
C473 B.n309 VSUBS 0.007687f
C474 B.n310 VSUBS 0.007687f
C475 B.n311 VSUBS 0.007687f
C476 B.n312 VSUBS 0.007687f
C477 B.n313 VSUBS 0.007687f
C478 B.n314 VSUBS 0.007687f
C479 B.n315 VSUBS 0.007687f
C480 B.n316 VSUBS 0.007687f
C481 B.n317 VSUBS 0.007687f
C482 B.n318 VSUBS 0.007687f
C483 B.n319 VSUBS 0.007687f
C484 B.n320 VSUBS 0.007687f
C485 B.n321 VSUBS 0.007687f
C486 B.n322 VSUBS 0.007687f
C487 B.n323 VSUBS 0.007687f
C488 B.n324 VSUBS 0.007687f
C489 B.n325 VSUBS 0.007687f
C490 B.n326 VSUBS 0.007687f
C491 B.n327 VSUBS 0.007687f
C492 B.n328 VSUBS 0.007687f
C493 B.n329 VSUBS 0.007687f
C494 B.n330 VSUBS 0.007687f
C495 B.n331 VSUBS 0.007687f
C496 B.n332 VSUBS 0.007687f
C497 B.n333 VSUBS 0.007687f
C498 B.n334 VSUBS 0.007687f
C499 B.n335 VSUBS 0.007687f
C500 B.n336 VSUBS 0.007687f
C501 B.n337 VSUBS 0.007687f
C502 B.n338 VSUBS 0.007687f
C503 B.n339 VSUBS 0.007687f
C504 B.n340 VSUBS 0.007687f
C505 B.n341 VSUBS 0.007687f
C506 B.n342 VSUBS 0.007687f
C507 B.n343 VSUBS 0.007687f
C508 B.n344 VSUBS 0.007687f
C509 B.n345 VSUBS 0.007687f
C510 B.n346 VSUBS 0.007687f
C511 B.n347 VSUBS 0.007687f
C512 B.n348 VSUBS 0.007687f
C513 B.n349 VSUBS 0.007687f
C514 B.n350 VSUBS 0.007687f
C515 B.n351 VSUBS 0.007687f
C516 B.n352 VSUBS 0.007687f
C517 B.n353 VSUBS 0.007687f
C518 B.n354 VSUBS 0.007687f
C519 B.n355 VSUBS 0.007687f
C520 B.n356 VSUBS 0.007687f
C521 B.n357 VSUBS 0.007687f
C522 B.n358 VSUBS 0.007687f
C523 B.n359 VSUBS 0.007687f
C524 B.n360 VSUBS 0.007687f
C525 B.n361 VSUBS 0.007687f
C526 B.n362 VSUBS 0.007687f
C527 B.n363 VSUBS 0.007687f
C528 B.n364 VSUBS 0.007687f
C529 B.n365 VSUBS 0.007687f
C530 B.n366 VSUBS 0.007687f
C531 B.n367 VSUBS 0.007687f
C532 B.n368 VSUBS 0.007687f
C533 B.n369 VSUBS 0.007687f
C534 B.n370 VSUBS 0.007687f
C535 B.n371 VSUBS 0.007687f
C536 B.n372 VSUBS 0.007687f
C537 B.n373 VSUBS 0.007687f
C538 B.n374 VSUBS 0.007687f
C539 B.n375 VSUBS 0.007687f
C540 B.n376 VSUBS 0.007687f
C541 B.n377 VSUBS 0.007687f
C542 B.n378 VSUBS 0.007687f
C543 B.n379 VSUBS 0.007687f
C544 B.n380 VSUBS 0.007687f
C545 B.n381 VSUBS 0.007687f
C546 B.n382 VSUBS 0.007687f
C547 B.n383 VSUBS 0.007687f
C548 B.n384 VSUBS 0.007687f
C549 B.n385 VSUBS 0.007687f
C550 B.n386 VSUBS 0.007687f
C551 B.n387 VSUBS 0.007687f
C552 B.n388 VSUBS 0.007687f
C553 B.n389 VSUBS 0.01839f
C554 B.n390 VSUBS 0.019595f
C555 B.n391 VSUBS 0.019595f
C556 B.n392 VSUBS 0.007687f
C557 B.n393 VSUBS 0.007687f
C558 B.n394 VSUBS 0.007687f
C559 B.n395 VSUBS 0.007687f
C560 B.n396 VSUBS 0.007687f
C561 B.n397 VSUBS 0.007687f
C562 B.n398 VSUBS 0.007687f
C563 B.n399 VSUBS 0.007687f
C564 B.n400 VSUBS 0.007687f
C565 B.n401 VSUBS 0.007687f
C566 B.n402 VSUBS 0.007687f
C567 B.n403 VSUBS 0.007687f
C568 B.n404 VSUBS 0.007687f
C569 B.n405 VSUBS 0.007687f
C570 B.n406 VSUBS 0.007687f
C571 B.n407 VSUBS 0.007687f
C572 B.n408 VSUBS 0.007687f
C573 B.n409 VSUBS 0.007687f
C574 B.n410 VSUBS 0.007687f
C575 B.n411 VSUBS 0.007687f
C576 B.n412 VSUBS 0.007687f
C577 B.n413 VSUBS 0.007687f
C578 B.n414 VSUBS 0.007687f
C579 B.n415 VSUBS 0.007687f
C580 B.n416 VSUBS 0.007687f
C581 B.n417 VSUBS 0.007687f
C582 B.n418 VSUBS 0.007687f
C583 B.n419 VSUBS 0.007687f
C584 B.n420 VSUBS 0.007687f
C585 B.n421 VSUBS 0.007687f
C586 B.n422 VSUBS 0.007687f
C587 B.n423 VSUBS 0.007687f
C588 B.n424 VSUBS 0.007687f
C589 B.n425 VSUBS 0.007687f
C590 B.n426 VSUBS 0.007687f
C591 B.n427 VSUBS 0.007687f
C592 B.n428 VSUBS 0.007687f
C593 B.n429 VSUBS 0.007687f
C594 B.n430 VSUBS 0.007687f
C595 B.n431 VSUBS 0.007687f
C596 B.n432 VSUBS 0.007687f
C597 B.n433 VSUBS 0.007687f
C598 B.n434 VSUBS 0.007687f
C599 B.n435 VSUBS 0.007687f
C600 B.n436 VSUBS 0.007687f
C601 B.n437 VSUBS 0.007687f
C602 B.n438 VSUBS 0.007687f
C603 B.n439 VSUBS 0.007687f
C604 B.n440 VSUBS 0.007687f
C605 B.n441 VSUBS 0.007687f
C606 B.n442 VSUBS 0.007687f
C607 B.n443 VSUBS 0.007687f
C608 B.n444 VSUBS 0.007687f
C609 B.n445 VSUBS 0.007687f
C610 B.n446 VSUBS 0.007687f
C611 B.n447 VSUBS 0.007687f
C612 B.n448 VSUBS 0.007687f
C613 B.n449 VSUBS 0.007687f
C614 B.n450 VSUBS 0.007687f
C615 B.n451 VSUBS 0.007687f
C616 B.n452 VSUBS 0.007687f
C617 B.n453 VSUBS 0.007687f
C618 B.n454 VSUBS 0.007687f
C619 B.n455 VSUBS 0.007687f
C620 B.n456 VSUBS 0.007687f
C621 B.n457 VSUBS 0.007687f
C622 B.n458 VSUBS 0.007687f
C623 B.n459 VSUBS 0.007687f
C624 B.n460 VSUBS 0.007687f
C625 B.n461 VSUBS 0.007687f
C626 B.n462 VSUBS 0.007687f
C627 B.n463 VSUBS 0.007687f
C628 B.n464 VSUBS 0.007687f
C629 B.n465 VSUBS 0.007687f
C630 B.n466 VSUBS 0.007687f
C631 B.n467 VSUBS 0.007687f
C632 B.n468 VSUBS 0.007687f
C633 B.n469 VSUBS 0.007687f
C634 B.n470 VSUBS 0.007687f
C635 B.n471 VSUBS 0.007687f
C636 B.n472 VSUBS 0.007687f
C637 B.n473 VSUBS 0.007687f
C638 B.n474 VSUBS 0.007687f
C639 B.n475 VSUBS 0.007687f
C640 B.n476 VSUBS 0.007687f
C641 B.n477 VSUBS 0.007687f
C642 B.n478 VSUBS 0.007687f
C643 B.n479 VSUBS 0.007687f
C644 B.n480 VSUBS 0.007687f
C645 B.n481 VSUBS 0.007235f
C646 B.n482 VSUBS 0.017811f
C647 B.n483 VSUBS 0.004296f
C648 B.n484 VSUBS 0.007687f
C649 B.n485 VSUBS 0.007687f
C650 B.n486 VSUBS 0.007687f
C651 B.n487 VSUBS 0.007687f
C652 B.n488 VSUBS 0.007687f
C653 B.n489 VSUBS 0.007687f
C654 B.n490 VSUBS 0.007687f
C655 B.n491 VSUBS 0.007687f
C656 B.n492 VSUBS 0.007687f
C657 B.n493 VSUBS 0.007687f
C658 B.n494 VSUBS 0.007687f
C659 B.n495 VSUBS 0.007687f
C660 B.n496 VSUBS 0.004296f
C661 B.n497 VSUBS 0.007687f
C662 B.n498 VSUBS 0.007687f
C663 B.n499 VSUBS 0.007235f
C664 B.n500 VSUBS 0.007687f
C665 B.n501 VSUBS 0.007687f
C666 B.n502 VSUBS 0.007687f
C667 B.n503 VSUBS 0.007687f
C668 B.n504 VSUBS 0.007687f
C669 B.n505 VSUBS 0.007687f
C670 B.n506 VSUBS 0.007687f
C671 B.n507 VSUBS 0.007687f
C672 B.n508 VSUBS 0.007687f
C673 B.n509 VSUBS 0.007687f
C674 B.n510 VSUBS 0.007687f
C675 B.n511 VSUBS 0.007687f
C676 B.n512 VSUBS 0.007687f
C677 B.n513 VSUBS 0.007687f
C678 B.n514 VSUBS 0.007687f
C679 B.n515 VSUBS 0.007687f
C680 B.n516 VSUBS 0.007687f
C681 B.n517 VSUBS 0.007687f
C682 B.n518 VSUBS 0.007687f
C683 B.n519 VSUBS 0.007687f
C684 B.n520 VSUBS 0.007687f
C685 B.n521 VSUBS 0.007687f
C686 B.n522 VSUBS 0.007687f
C687 B.n523 VSUBS 0.007687f
C688 B.n524 VSUBS 0.007687f
C689 B.n525 VSUBS 0.007687f
C690 B.n526 VSUBS 0.007687f
C691 B.n527 VSUBS 0.007687f
C692 B.n528 VSUBS 0.007687f
C693 B.n529 VSUBS 0.007687f
C694 B.n530 VSUBS 0.007687f
C695 B.n531 VSUBS 0.007687f
C696 B.n532 VSUBS 0.007687f
C697 B.n533 VSUBS 0.007687f
C698 B.n534 VSUBS 0.007687f
C699 B.n535 VSUBS 0.007687f
C700 B.n536 VSUBS 0.007687f
C701 B.n537 VSUBS 0.007687f
C702 B.n538 VSUBS 0.007687f
C703 B.n539 VSUBS 0.007687f
C704 B.n540 VSUBS 0.007687f
C705 B.n541 VSUBS 0.007687f
C706 B.n542 VSUBS 0.007687f
C707 B.n543 VSUBS 0.007687f
C708 B.n544 VSUBS 0.007687f
C709 B.n545 VSUBS 0.007687f
C710 B.n546 VSUBS 0.007687f
C711 B.n547 VSUBS 0.007687f
C712 B.n548 VSUBS 0.007687f
C713 B.n549 VSUBS 0.007687f
C714 B.n550 VSUBS 0.007687f
C715 B.n551 VSUBS 0.007687f
C716 B.n552 VSUBS 0.007687f
C717 B.n553 VSUBS 0.007687f
C718 B.n554 VSUBS 0.007687f
C719 B.n555 VSUBS 0.007687f
C720 B.n556 VSUBS 0.007687f
C721 B.n557 VSUBS 0.007687f
C722 B.n558 VSUBS 0.007687f
C723 B.n559 VSUBS 0.007687f
C724 B.n560 VSUBS 0.007687f
C725 B.n561 VSUBS 0.007687f
C726 B.n562 VSUBS 0.007687f
C727 B.n563 VSUBS 0.007687f
C728 B.n564 VSUBS 0.007687f
C729 B.n565 VSUBS 0.007687f
C730 B.n566 VSUBS 0.007687f
C731 B.n567 VSUBS 0.007687f
C732 B.n568 VSUBS 0.007687f
C733 B.n569 VSUBS 0.007687f
C734 B.n570 VSUBS 0.007687f
C735 B.n571 VSUBS 0.007687f
C736 B.n572 VSUBS 0.007687f
C737 B.n573 VSUBS 0.007687f
C738 B.n574 VSUBS 0.007687f
C739 B.n575 VSUBS 0.007687f
C740 B.n576 VSUBS 0.007687f
C741 B.n577 VSUBS 0.007687f
C742 B.n578 VSUBS 0.007687f
C743 B.n579 VSUBS 0.007687f
C744 B.n580 VSUBS 0.007687f
C745 B.n581 VSUBS 0.007687f
C746 B.n582 VSUBS 0.007687f
C747 B.n583 VSUBS 0.007687f
C748 B.n584 VSUBS 0.007687f
C749 B.n585 VSUBS 0.007687f
C750 B.n586 VSUBS 0.007687f
C751 B.n587 VSUBS 0.007687f
C752 B.n588 VSUBS 0.019595f
C753 B.n589 VSUBS 0.019595f
C754 B.n590 VSUBS 0.01839f
C755 B.n591 VSUBS 0.007687f
C756 B.n592 VSUBS 0.007687f
C757 B.n593 VSUBS 0.007687f
C758 B.n594 VSUBS 0.007687f
C759 B.n595 VSUBS 0.007687f
C760 B.n596 VSUBS 0.007687f
C761 B.n597 VSUBS 0.007687f
C762 B.n598 VSUBS 0.007687f
C763 B.n599 VSUBS 0.007687f
C764 B.n600 VSUBS 0.007687f
C765 B.n601 VSUBS 0.007687f
C766 B.n602 VSUBS 0.007687f
C767 B.n603 VSUBS 0.007687f
C768 B.n604 VSUBS 0.007687f
C769 B.n605 VSUBS 0.007687f
C770 B.n606 VSUBS 0.007687f
C771 B.n607 VSUBS 0.007687f
C772 B.n608 VSUBS 0.007687f
C773 B.n609 VSUBS 0.007687f
C774 B.n610 VSUBS 0.007687f
C775 B.n611 VSUBS 0.007687f
C776 B.n612 VSUBS 0.007687f
C777 B.n613 VSUBS 0.007687f
C778 B.n614 VSUBS 0.007687f
C779 B.n615 VSUBS 0.007687f
C780 B.n616 VSUBS 0.007687f
C781 B.n617 VSUBS 0.007687f
C782 B.n618 VSUBS 0.007687f
C783 B.n619 VSUBS 0.007687f
C784 B.n620 VSUBS 0.007687f
C785 B.n621 VSUBS 0.007687f
C786 B.n622 VSUBS 0.007687f
C787 B.n623 VSUBS 0.007687f
C788 B.n624 VSUBS 0.007687f
C789 B.n625 VSUBS 0.007687f
C790 B.n626 VSUBS 0.007687f
C791 B.n627 VSUBS 0.007687f
C792 B.n628 VSUBS 0.007687f
C793 B.n629 VSUBS 0.007687f
C794 B.n630 VSUBS 0.007687f
C795 B.n631 VSUBS 0.007687f
C796 B.n632 VSUBS 0.007687f
C797 B.n633 VSUBS 0.007687f
C798 B.n634 VSUBS 0.007687f
C799 B.n635 VSUBS 0.007687f
C800 B.n636 VSUBS 0.007687f
C801 B.n637 VSUBS 0.007687f
C802 B.n638 VSUBS 0.007687f
C803 B.n639 VSUBS 0.007687f
C804 B.n640 VSUBS 0.007687f
C805 B.n641 VSUBS 0.007687f
C806 B.n642 VSUBS 0.007687f
C807 B.n643 VSUBS 0.007687f
C808 B.n644 VSUBS 0.007687f
C809 B.n645 VSUBS 0.007687f
C810 B.n646 VSUBS 0.007687f
C811 B.n647 VSUBS 0.007687f
C812 B.n648 VSUBS 0.007687f
C813 B.n649 VSUBS 0.007687f
C814 B.n650 VSUBS 0.007687f
C815 B.n651 VSUBS 0.007687f
C816 B.n652 VSUBS 0.007687f
C817 B.n653 VSUBS 0.007687f
C818 B.n654 VSUBS 0.007687f
C819 B.n655 VSUBS 0.007687f
C820 B.n656 VSUBS 0.007687f
C821 B.n657 VSUBS 0.007687f
C822 B.n658 VSUBS 0.007687f
C823 B.n659 VSUBS 0.007687f
C824 B.n660 VSUBS 0.007687f
C825 B.n661 VSUBS 0.007687f
C826 B.n662 VSUBS 0.007687f
C827 B.n663 VSUBS 0.007687f
C828 B.n664 VSUBS 0.007687f
C829 B.n665 VSUBS 0.007687f
C830 B.n666 VSUBS 0.007687f
C831 B.n667 VSUBS 0.007687f
C832 B.n668 VSUBS 0.007687f
C833 B.n669 VSUBS 0.007687f
C834 B.n670 VSUBS 0.007687f
C835 B.n671 VSUBS 0.007687f
C836 B.n672 VSUBS 0.007687f
C837 B.n673 VSUBS 0.007687f
C838 B.n674 VSUBS 0.007687f
C839 B.n675 VSUBS 0.007687f
C840 B.n676 VSUBS 0.007687f
C841 B.n677 VSUBS 0.007687f
C842 B.n678 VSUBS 0.007687f
C843 B.n679 VSUBS 0.007687f
C844 B.n680 VSUBS 0.007687f
C845 B.n681 VSUBS 0.007687f
C846 B.n682 VSUBS 0.007687f
C847 B.n683 VSUBS 0.007687f
C848 B.n684 VSUBS 0.007687f
C849 B.n685 VSUBS 0.007687f
C850 B.n686 VSUBS 0.007687f
C851 B.n687 VSUBS 0.007687f
C852 B.n688 VSUBS 0.007687f
C853 B.n689 VSUBS 0.007687f
C854 B.n690 VSUBS 0.007687f
C855 B.n691 VSUBS 0.007687f
C856 B.n692 VSUBS 0.007687f
C857 B.n693 VSUBS 0.007687f
C858 B.n694 VSUBS 0.007687f
C859 B.n695 VSUBS 0.007687f
C860 B.n696 VSUBS 0.007687f
C861 B.n697 VSUBS 0.007687f
C862 B.n698 VSUBS 0.007687f
C863 B.n699 VSUBS 0.007687f
C864 B.n700 VSUBS 0.007687f
C865 B.n701 VSUBS 0.007687f
C866 B.n702 VSUBS 0.007687f
C867 B.n703 VSUBS 0.007687f
C868 B.n704 VSUBS 0.007687f
C869 B.n705 VSUBS 0.007687f
C870 B.n706 VSUBS 0.007687f
C871 B.n707 VSUBS 0.007687f
C872 B.n708 VSUBS 0.007687f
C873 B.n709 VSUBS 0.007687f
C874 B.n710 VSUBS 0.007687f
C875 B.n711 VSUBS 0.007687f
C876 B.n712 VSUBS 0.007687f
C877 B.n713 VSUBS 0.007687f
C878 B.n714 VSUBS 0.007687f
C879 B.n715 VSUBS 0.007687f
C880 B.n716 VSUBS 0.007687f
C881 B.n717 VSUBS 0.007687f
C882 B.n718 VSUBS 0.007687f
C883 B.n719 VSUBS 0.007687f
C884 B.n720 VSUBS 0.007687f
C885 B.n721 VSUBS 0.007687f
C886 B.n722 VSUBS 0.007687f
C887 B.n723 VSUBS 0.007687f
C888 B.n724 VSUBS 0.007687f
C889 B.n725 VSUBS 0.007687f
C890 B.n726 VSUBS 0.007687f
C891 B.n727 VSUBS 0.007687f
C892 B.n728 VSUBS 0.007687f
C893 B.n729 VSUBS 0.007687f
C894 B.n730 VSUBS 0.007687f
C895 B.n731 VSUBS 0.007687f
C896 B.n732 VSUBS 0.007687f
C897 B.n733 VSUBS 0.007687f
C898 B.n734 VSUBS 0.007687f
C899 B.n735 VSUBS 0.007687f
C900 B.n736 VSUBS 0.007687f
C901 B.n737 VSUBS 0.007687f
C902 B.n738 VSUBS 0.007687f
C903 B.n739 VSUBS 0.007687f
C904 B.n740 VSUBS 0.007687f
C905 B.n741 VSUBS 0.007687f
C906 B.n742 VSUBS 0.007687f
C907 B.n743 VSUBS 0.007687f
C908 B.n744 VSUBS 0.007687f
C909 B.n745 VSUBS 0.007687f
C910 B.n746 VSUBS 0.007687f
C911 B.n747 VSUBS 0.007687f
C912 B.n748 VSUBS 0.007687f
C913 B.n749 VSUBS 0.007687f
C914 B.n750 VSUBS 0.007687f
C915 B.n751 VSUBS 0.007687f
C916 B.n752 VSUBS 0.007687f
C917 B.n753 VSUBS 0.007687f
C918 B.n754 VSUBS 0.007687f
C919 B.n755 VSUBS 0.007687f
C920 B.n756 VSUBS 0.007687f
C921 B.n757 VSUBS 0.007687f
C922 B.n758 VSUBS 0.007687f
C923 B.n759 VSUBS 0.007687f
C924 B.n760 VSUBS 0.007687f
C925 B.n761 VSUBS 0.007687f
C926 B.n762 VSUBS 0.007687f
C927 B.n763 VSUBS 0.007687f
C928 B.n764 VSUBS 0.007687f
C929 B.n765 VSUBS 0.007687f
C930 B.n766 VSUBS 0.007687f
C931 B.n767 VSUBS 0.007687f
C932 B.n768 VSUBS 0.007687f
C933 B.n769 VSUBS 0.007687f
C934 B.n770 VSUBS 0.007687f
C935 B.n771 VSUBS 0.007687f
C936 B.n772 VSUBS 0.007687f
C937 B.n773 VSUBS 0.007687f
C938 B.n774 VSUBS 0.007687f
C939 B.n775 VSUBS 0.007687f
C940 B.n776 VSUBS 0.007687f
C941 B.n777 VSUBS 0.007687f
C942 B.n778 VSUBS 0.007687f
C943 B.n779 VSUBS 0.007687f
C944 B.n780 VSUBS 0.007687f
C945 B.n781 VSUBS 0.007687f
C946 B.n782 VSUBS 0.007687f
C947 B.n783 VSUBS 0.007687f
C948 B.n784 VSUBS 0.007687f
C949 B.n785 VSUBS 0.007687f
C950 B.n786 VSUBS 0.007687f
C951 B.n787 VSUBS 0.007687f
C952 B.n788 VSUBS 0.007687f
C953 B.n789 VSUBS 0.007687f
C954 B.n790 VSUBS 0.007687f
C955 B.n791 VSUBS 0.007687f
C956 B.n792 VSUBS 0.007687f
C957 B.n793 VSUBS 0.007687f
C958 B.n794 VSUBS 0.007687f
C959 B.n795 VSUBS 0.007687f
C960 B.n796 VSUBS 0.007687f
C961 B.n797 VSUBS 0.007687f
C962 B.n798 VSUBS 0.007687f
C963 B.n799 VSUBS 0.007687f
C964 B.n800 VSUBS 0.007687f
C965 B.n801 VSUBS 0.007687f
C966 B.n802 VSUBS 0.007687f
C967 B.n803 VSUBS 0.01839f
C968 B.n804 VSUBS 0.019595f
C969 B.n805 VSUBS 0.018757f
C970 B.n806 VSUBS 0.007687f
C971 B.n807 VSUBS 0.007687f
C972 B.n808 VSUBS 0.007687f
C973 B.n809 VSUBS 0.007687f
C974 B.n810 VSUBS 0.007687f
C975 B.n811 VSUBS 0.007687f
C976 B.n812 VSUBS 0.007687f
C977 B.n813 VSUBS 0.007687f
C978 B.n814 VSUBS 0.007687f
C979 B.n815 VSUBS 0.007687f
C980 B.n816 VSUBS 0.007687f
C981 B.n817 VSUBS 0.007687f
C982 B.n818 VSUBS 0.007687f
C983 B.n819 VSUBS 0.007687f
C984 B.n820 VSUBS 0.007687f
C985 B.n821 VSUBS 0.007687f
C986 B.n822 VSUBS 0.007687f
C987 B.n823 VSUBS 0.007687f
C988 B.n824 VSUBS 0.007687f
C989 B.n825 VSUBS 0.007687f
C990 B.n826 VSUBS 0.007687f
C991 B.n827 VSUBS 0.007687f
C992 B.n828 VSUBS 0.007687f
C993 B.n829 VSUBS 0.007687f
C994 B.n830 VSUBS 0.007687f
C995 B.n831 VSUBS 0.007687f
C996 B.n832 VSUBS 0.007687f
C997 B.n833 VSUBS 0.007687f
C998 B.n834 VSUBS 0.007687f
C999 B.n835 VSUBS 0.007687f
C1000 B.n836 VSUBS 0.007687f
C1001 B.n837 VSUBS 0.007687f
C1002 B.n838 VSUBS 0.007687f
C1003 B.n839 VSUBS 0.007687f
C1004 B.n840 VSUBS 0.007687f
C1005 B.n841 VSUBS 0.007687f
C1006 B.n842 VSUBS 0.007687f
C1007 B.n843 VSUBS 0.007687f
C1008 B.n844 VSUBS 0.007687f
C1009 B.n845 VSUBS 0.007687f
C1010 B.n846 VSUBS 0.007687f
C1011 B.n847 VSUBS 0.007687f
C1012 B.n848 VSUBS 0.007687f
C1013 B.n849 VSUBS 0.007687f
C1014 B.n850 VSUBS 0.007687f
C1015 B.n851 VSUBS 0.007687f
C1016 B.n852 VSUBS 0.007687f
C1017 B.n853 VSUBS 0.007687f
C1018 B.n854 VSUBS 0.007687f
C1019 B.n855 VSUBS 0.007687f
C1020 B.n856 VSUBS 0.007687f
C1021 B.n857 VSUBS 0.007687f
C1022 B.n858 VSUBS 0.007687f
C1023 B.n859 VSUBS 0.007687f
C1024 B.n860 VSUBS 0.007687f
C1025 B.n861 VSUBS 0.007687f
C1026 B.n862 VSUBS 0.007687f
C1027 B.n863 VSUBS 0.007687f
C1028 B.n864 VSUBS 0.007687f
C1029 B.n865 VSUBS 0.007687f
C1030 B.n866 VSUBS 0.007687f
C1031 B.n867 VSUBS 0.007687f
C1032 B.n868 VSUBS 0.007687f
C1033 B.n869 VSUBS 0.007687f
C1034 B.n870 VSUBS 0.007687f
C1035 B.n871 VSUBS 0.007687f
C1036 B.n872 VSUBS 0.007687f
C1037 B.n873 VSUBS 0.007687f
C1038 B.n874 VSUBS 0.007687f
C1039 B.n875 VSUBS 0.007687f
C1040 B.n876 VSUBS 0.007687f
C1041 B.n877 VSUBS 0.007687f
C1042 B.n878 VSUBS 0.007687f
C1043 B.n879 VSUBS 0.007687f
C1044 B.n880 VSUBS 0.007687f
C1045 B.n881 VSUBS 0.007687f
C1046 B.n882 VSUBS 0.007687f
C1047 B.n883 VSUBS 0.007687f
C1048 B.n884 VSUBS 0.007687f
C1049 B.n885 VSUBS 0.007687f
C1050 B.n886 VSUBS 0.007687f
C1051 B.n887 VSUBS 0.007687f
C1052 B.n888 VSUBS 0.007687f
C1053 B.n889 VSUBS 0.007687f
C1054 B.n890 VSUBS 0.007687f
C1055 B.n891 VSUBS 0.007687f
C1056 B.n892 VSUBS 0.007687f
C1057 B.n893 VSUBS 0.007687f
C1058 B.n894 VSUBS 0.007687f
C1059 B.n895 VSUBS 0.007235f
C1060 B.n896 VSUBS 0.017811f
C1061 B.n897 VSUBS 0.004296f
C1062 B.n898 VSUBS 0.007687f
C1063 B.n899 VSUBS 0.007687f
C1064 B.n900 VSUBS 0.007687f
C1065 B.n901 VSUBS 0.007687f
C1066 B.n902 VSUBS 0.007687f
C1067 B.n903 VSUBS 0.007687f
C1068 B.n904 VSUBS 0.007687f
C1069 B.n905 VSUBS 0.007687f
C1070 B.n906 VSUBS 0.007687f
C1071 B.n907 VSUBS 0.007687f
C1072 B.n908 VSUBS 0.007687f
C1073 B.n909 VSUBS 0.007687f
C1074 B.n910 VSUBS 0.004296f
C1075 B.n911 VSUBS 0.007687f
C1076 B.n912 VSUBS 0.007687f
C1077 B.n913 VSUBS 0.007235f
C1078 B.n914 VSUBS 0.007687f
C1079 B.n915 VSUBS 0.007687f
C1080 B.n916 VSUBS 0.007687f
C1081 B.n917 VSUBS 0.007687f
C1082 B.n918 VSUBS 0.007687f
C1083 B.n919 VSUBS 0.007687f
C1084 B.n920 VSUBS 0.007687f
C1085 B.n921 VSUBS 0.007687f
C1086 B.n922 VSUBS 0.007687f
C1087 B.n923 VSUBS 0.007687f
C1088 B.n924 VSUBS 0.007687f
C1089 B.n925 VSUBS 0.007687f
C1090 B.n926 VSUBS 0.007687f
C1091 B.n927 VSUBS 0.007687f
C1092 B.n928 VSUBS 0.007687f
C1093 B.n929 VSUBS 0.007687f
C1094 B.n930 VSUBS 0.007687f
C1095 B.n931 VSUBS 0.007687f
C1096 B.n932 VSUBS 0.007687f
C1097 B.n933 VSUBS 0.007687f
C1098 B.n934 VSUBS 0.007687f
C1099 B.n935 VSUBS 0.007687f
C1100 B.n936 VSUBS 0.007687f
C1101 B.n937 VSUBS 0.007687f
C1102 B.n938 VSUBS 0.007687f
C1103 B.n939 VSUBS 0.007687f
C1104 B.n940 VSUBS 0.007687f
C1105 B.n941 VSUBS 0.007687f
C1106 B.n942 VSUBS 0.007687f
C1107 B.n943 VSUBS 0.007687f
C1108 B.n944 VSUBS 0.007687f
C1109 B.n945 VSUBS 0.007687f
C1110 B.n946 VSUBS 0.007687f
C1111 B.n947 VSUBS 0.007687f
C1112 B.n948 VSUBS 0.007687f
C1113 B.n949 VSUBS 0.007687f
C1114 B.n950 VSUBS 0.007687f
C1115 B.n951 VSUBS 0.007687f
C1116 B.n952 VSUBS 0.007687f
C1117 B.n953 VSUBS 0.007687f
C1118 B.n954 VSUBS 0.007687f
C1119 B.n955 VSUBS 0.007687f
C1120 B.n956 VSUBS 0.007687f
C1121 B.n957 VSUBS 0.007687f
C1122 B.n958 VSUBS 0.007687f
C1123 B.n959 VSUBS 0.007687f
C1124 B.n960 VSUBS 0.007687f
C1125 B.n961 VSUBS 0.007687f
C1126 B.n962 VSUBS 0.007687f
C1127 B.n963 VSUBS 0.007687f
C1128 B.n964 VSUBS 0.007687f
C1129 B.n965 VSUBS 0.007687f
C1130 B.n966 VSUBS 0.007687f
C1131 B.n967 VSUBS 0.007687f
C1132 B.n968 VSUBS 0.007687f
C1133 B.n969 VSUBS 0.007687f
C1134 B.n970 VSUBS 0.007687f
C1135 B.n971 VSUBS 0.007687f
C1136 B.n972 VSUBS 0.007687f
C1137 B.n973 VSUBS 0.007687f
C1138 B.n974 VSUBS 0.007687f
C1139 B.n975 VSUBS 0.007687f
C1140 B.n976 VSUBS 0.007687f
C1141 B.n977 VSUBS 0.007687f
C1142 B.n978 VSUBS 0.007687f
C1143 B.n979 VSUBS 0.007687f
C1144 B.n980 VSUBS 0.007687f
C1145 B.n981 VSUBS 0.007687f
C1146 B.n982 VSUBS 0.007687f
C1147 B.n983 VSUBS 0.007687f
C1148 B.n984 VSUBS 0.007687f
C1149 B.n985 VSUBS 0.007687f
C1150 B.n986 VSUBS 0.007687f
C1151 B.n987 VSUBS 0.007687f
C1152 B.n988 VSUBS 0.007687f
C1153 B.n989 VSUBS 0.007687f
C1154 B.n990 VSUBS 0.007687f
C1155 B.n991 VSUBS 0.007687f
C1156 B.n992 VSUBS 0.007687f
C1157 B.n993 VSUBS 0.007687f
C1158 B.n994 VSUBS 0.007687f
C1159 B.n995 VSUBS 0.007687f
C1160 B.n996 VSUBS 0.007687f
C1161 B.n997 VSUBS 0.007687f
C1162 B.n998 VSUBS 0.007687f
C1163 B.n999 VSUBS 0.007687f
C1164 B.n1000 VSUBS 0.007687f
C1165 B.n1001 VSUBS 0.007687f
C1166 B.n1002 VSUBS 0.019595f
C1167 B.n1003 VSUBS 0.019595f
C1168 B.n1004 VSUBS 0.01839f
C1169 B.n1005 VSUBS 0.007687f
C1170 B.n1006 VSUBS 0.007687f
C1171 B.n1007 VSUBS 0.007687f
C1172 B.n1008 VSUBS 0.007687f
C1173 B.n1009 VSUBS 0.007687f
C1174 B.n1010 VSUBS 0.007687f
C1175 B.n1011 VSUBS 0.007687f
C1176 B.n1012 VSUBS 0.007687f
C1177 B.n1013 VSUBS 0.007687f
C1178 B.n1014 VSUBS 0.007687f
C1179 B.n1015 VSUBS 0.007687f
C1180 B.n1016 VSUBS 0.007687f
C1181 B.n1017 VSUBS 0.007687f
C1182 B.n1018 VSUBS 0.007687f
C1183 B.n1019 VSUBS 0.007687f
C1184 B.n1020 VSUBS 0.007687f
C1185 B.n1021 VSUBS 0.007687f
C1186 B.n1022 VSUBS 0.007687f
C1187 B.n1023 VSUBS 0.007687f
C1188 B.n1024 VSUBS 0.007687f
C1189 B.n1025 VSUBS 0.007687f
C1190 B.n1026 VSUBS 0.007687f
C1191 B.n1027 VSUBS 0.007687f
C1192 B.n1028 VSUBS 0.007687f
C1193 B.n1029 VSUBS 0.007687f
C1194 B.n1030 VSUBS 0.007687f
C1195 B.n1031 VSUBS 0.007687f
C1196 B.n1032 VSUBS 0.007687f
C1197 B.n1033 VSUBS 0.007687f
C1198 B.n1034 VSUBS 0.007687f
C1199 B.n1035 VSUBS 0.007687f
C1200 B.n1036 VSUBS 0.007687f
C1201 B.n1037 VSUBS 0.007687f
C1202 B.n1038 VSUBS 0.007687f
C1203 B.n1039 VSUBS 0.007687f
C1204 B.n1040 VSUBS 0.007687f
C1205 B.n1041 VSUBS 0.007687f
C1206 B.n1042 VSUBS 0.007687f
C1207 B.n1043 VSUBS 0.007687f
C1208 B.n1044 VSUBS 0.007687f
C1209 B.n1045 VSUBS 0.007687f
C1210 B.n1046 VSUBS 0.007687f
C1211 B.n1047 VSUBS 0.007687f
C1212 B.n1048 VSUBS 0.007687f
C1213 B.n1049 VSUBS 0.007687f
C1214 B.n1050 VSUBS 0.007687f
C1215 B.n1051 VSUBS 0.007687f
C1216 B.n1052 VSUBS 0.007687f
C1217 B.n1053 VSUBS 0.007687f
C1218 B.n1054 VSUBS 0.007687f
C1219 B.n1055 VSUBS 0.007687f
C1220 B.n1056 VSUBS 0.007687f
C1221 B.n1057 VSUBS 0.007687f
C1222 B.n1058 VSUBS 0.007687f
C1223 B.n1059 VSUBS 0.007687f
C1224 B.n1060 VSUBS 0.007687f
C1225 B.n1061 VSUBS 0.007687f
C1226 B.n1062 VSUBS 0.007687f
C1227 B.n1063 VSUBS 0.007687f
C1228 B.n1064 VSUBS 0.007687f
C1229 B.n1065 VSUBS 0.007687f
C1230 B.n1066 VSUBS 0.007687f
C1231 B.n1067 VSUBS 0.007687f
C1232 B.n1068 VSUBS 0.007687f
C1233 B.n1069 VSUBS 0.007687f
C1234 B.n1070 VSUBS 0.007687f
C1235 B.n1071 VSUBS 0.007687f
C1236 B.n1072 VSUBS 0.007687f
C1237 B.n1073 VSUBS 0.007687f
C1238 B.n1074 VSUBS 0.007687f
C1239 B.n1075 VSUBS 0.007687f
C1240 B.n1076 VSUBS 0.007687f
C1241 B.n1077 VSUBS 0.007687f
C1242 B.n1078 VSUBS 0.007687f
C1243 B.n1079 VSUBS 0.007687f
C1244 B.n1080 VSUBS 0.007687f
C1245 B.n1081 VSUBS 0.007687f
C1246 B.n1082 VSUBS 0.007687f
C1247 B.n1083 VSUBS 0.007687f
C1248 B.n1084 VSUBS 0.007687f
C1249 B.n1085 VSUBS 0.007687f
C1250 B.n1086 VSUBS 0.007687f
C1251 B.n1087 VSUBS 0.007687f
C1252 B.n1088 VSUBS 0.007687f
C1253 B.n1089 VSUBS 0.007687f
C1254 B.n1090 VSUBS 0.007687f
C1255 B.n1091 VSUBS 0.007687f
C1256 B.n1092 VSUBS 0.007687f
C1257 B.n1093 VSUBS 0.007687f
C1258 B.n1094 VSUBS 0.007687f
C1259 B.n1095 VSUBS 0.007687f
C1260 B.n1096 VSUBS 0.007687f
C1261 B.n1097 VSUBS 0.007687f
C1262 B.n1098 VSUBS 0.007687f
C1263 B.n1099 VSUBS 0.007687f
C1264 B.n1100 VSUBS 0.007687f
C1265 B.n1101 VSUBS 0.007687f
C1266 B.n1102 VSUBS 0.007687f
C1267 B.n1103 VSUBS 0.007687f
C1268 B.n1104 VSUBS 0.007687f
C1269 B.n1105 VSUBS 0.007687f
C1270 B.n1106 VSUBS 0.007687f
C1271 B.n1107 VSUBS 0.007687f
C1272 B.n1108 VSUBS 0.007687f
C1273 B.n1109 VSUBS 0.007687f
C1274 B.n1110 VSUBS 0.007687f
C1275 B.n1111 VSUBS 0.017407f
C1276 VDD1.t7 VSUBS 4.6212f
C1277 VDD1.t8 VSUBS 0.422755f
C1278 VDD1.t2 VSUBS 0.422755f
C1279 VDD1.n0 VSUBS 3.53224f
C1280 VDD1.n1 VSUBS 1.84899f
C1281 VDD1.t9 VSUBS 4.62117f
C1282 VDD1.t4 VSUBS 0.422755f
C1283 VDD1.t3 VSUBS 0.422755f
C1284 VDD1.n2 VSUBS 3.53224f
C1285 VDD1.n3 VSUBS 1.83946f
C1286 VDD1.t1 VSUBS 0.422755f
C1287 VDD1.t6 VSUBS 0.422755f
C1288 VDD1.n4 VSUBS 3.5658f
C1289 VDD1.n5 VSUBS 4.68921f
C1290 VDD1.t5 VSUBS 0.422755f
C1291 VDD1.t0 VSUBS 0.422755f
C1292 VDD1.n6 VSUBS 3.53223f
C1293 VDD1.n7 VSUBS 4.85033f
C1294 VTAIL.t1 VSUBS 0.407036f
C1295 VTAIL.t4 VSUBS 0.407036f
C1296 VTAIL.n0 VSUBS 3.23194f
C1297 VTAIL.n1 VSUBS 1.06389f
C1298 VTAIL.t10 VSUBS 4.21684f
C1299 VTAIL.n2 VSUBS 1.25253f
C1300 VTAIL.t17 VSUBS 0.407036f
C1301 VTAIL.t15 VSUBS 0.407036f
C1302 VTAIL.n3 VSUBS 3.23194f
C1303 VTAIL.n4 VSUBS 1.2228f
C1304 VTAIL.t14 VSUBS 0.407036f
C1305 VTAIL.t16 VSUBS 0.407036f
C1306 VTAIL.n5 VSUBS 3.23194f
C1307 VTAIL.n6 VSUBS 3.30306f
C1308 VTAIL.t7 VSUBS 0.407036f
C1309 VTAIL.t6 VSUBS 0.407036f
C1310 VTAIL.n7 VSUBS 3.23194f
C1311 VTAIL.n8 VSUBS 3.30306f
C1312 VTAIL.t0 VSUBS 0.407036f
C1313 VTAIL.t9 VSUBS 0.407036f
C1314 VTAIL.n9 VSUBS 3.23194f
C1315 VTAIL.n10 VSUBS 1.22279f
C1316 VTAIL.t8 VSUBS 4.21687f
C1317 VTAIL.n11 VSUBS 1.2525f
C1318 VTAIL.t13 VSUBS 0.407036f
C1319 VTAIL.t19 VSUBS 0.407036f
C1320 VTAIL.n12 VSUBS 3.23194f
C1321 VTAIL.n13 VSUBS 1.12733f
C1322 VTAIL.t11 VSUBS 0.407036f
C1323 VTAIL.t18 VSUBS 0.407036f
C1324 VTAIL.n14 VSUBS 3.23194f
C1325 VTAIL.n15 VSUBS 1.22279f
C1326 VTAIL.t12 VSUBS 4.21684f
C1327 VTAIL.n16 VSUBS 3.15375f
C1328 VTAIL.t3 VSUBS 4.21684f
C1329 VTAIL.n17 VSUBS 3.15375f
C1330 VTAIL.t5 VSUBS 0.407036f
C1331 VTAIL.t2 VSUBS 0.407036f
C1332 VTAIL.n18 VSUBS 3.23194f
C1333 VTAIL.n19 VSUBS 1.01175f
C1334 VP.t3 VSUBS 3.93783f
C1335 VP.n0 VSUBS 1.45762f
C1336 VP.n1 VSUBS 0.023591f
C1337 VP.n2 VSUBS 0.023772f
C1338 VP.n3 VSUBS 0.023591f
C1339 VP.t8 VSUBS 3.93783f
C1340 VP.n4 VSUBS 1.35808f
C1341 VP.n5 VSUBS 0.023591f
C1342 VP.n6 VSUBS 0.019539f
C1343 VP.n7 VSUBS 0.023591f
C1344 VP.t6 VSUBS 3.93783f
C1345 VP.n8 VSUBS 1.35808f
C1346 VP.n9 VSUBS 0.023591f
C1347 VP.n10 VSUBS 0.019539f
C1348 VP.n11 VSUBS 0.023591f
C1349 VP.t5 VSUBS 3.93783f
C1350 VP.n12 VSUBS 1.35808f
C1351 VP.n13 VSUBS 0.023591f
C1352 VP.n14 VSUBS 0.023772f
C1353 VP.n15 VSUBS 0.023591f
C1354 VP.t0 VSUBS 3.93783f
C1355 VP.n16 VSUBS 1.45762f
C1356 VP.t9 VSUBS 3.93783f
C1357 VP.n17 VSUBS 1.45762f
C1358 VP.n18 VSUBS 0.023591f
C1359 VP.n19 VSUBS 0.023772f
C1360 VP.n20 VSUBS 0.023591f
C1361 VP.t4 VSUBS 3.93783f
C1362 VP.n21 VSUBS 1.35808f
C1363 VP.n22 VSUBS 0.023591f
C1364 VP.n23 VSUBS 0.019539f
C1365 VP.n24 VSUBS 0.023591f
C1366 VP.t7 VSUBS 3.93783f
C1367 VP.n25 VSUBS 1.35808f
C1368 VP.n26 VSUBS 0.023591f
C1369 VP.n27 VSUBS 0.019539f
C1370 VP.n28 VSUBS 0.023591f
C1371 VP.t1 VSUBS 3.93783f
C1372 VP.n29 VSUBS 1.43906f
C1373 VP.t2 VSUBS 4.23567f
C1374 VP.n30 VSUBS 1.38156f
C1375 VP.n31 VSUBS 0.272834f
C1376 VP.n32 VSUBS 0.036405f
C1377 VP.n33 VSUBS 0.043748f
C1378 VP.n34 VSUBS 0.045484f
C1379 VP.n35 VSUBS 0.023591f
C1380 VP.n36 VSUBS 0.023591f
C1381 VP.n37 VSUBS 0.023591f
C1382 VP.n38 VSUBS 0.047311f
C1383 VP.n39 VSUBS 0.043748f
C1384 VP.n40 VSUBS 0.032949f
C1385 VP.n41 VSUBS 0.023591f
C1386 VP.n42 VSUBS 0.023591f
C1387 VP.n43 VSUBS 0.032949f
C1388 VP.n44 VSUBS 0.043748f
C1389 VP.n45 VSUBS 0.047311f
C1390 VP.n46 VSUBS 0.023591f
C1391 VP.n47 VSUBS 0.023591f
C1392 VP.n48 VSUBS 0.023591f
C1393 VP.n49 VSUBS 0.045484f
C1394 VP.n50 VSUBS 0.043748f
C1395 VP.n51 VSUBS 0.036405f
C1396 VP.n52 VSUBS 0.023591f
C1397 VP.n53 VSUBS 0.023591f
C1398 VP.n54 VSUBS 0.029493f
C1399 VP.n55 VSUBS 0.043748f
C1400 VP.n56 VSUBS 0.046414f
C1401 VP.n57 VSUBS 0.023591f
C1402 VP.n58 VSUBS 0.023591f
C1403 VP.n59 VSUBS 0.023591f
C1404 VP.n60 VSUBS 0.042148f
C1405 VP.n61 VSUBS 0.043748f
C1406 VP.n62 VSUBS 0.03986f
C1407 VP.n63 VSUBS 0.03807f
C1408 VP.n64 VSUBS 1.79507f
C1409 VP.n65 VSUBS 1.80881f
C1410 VP.n66 VSUBS 0.03807f
C1411 VP.n67 VSUBS 0.03986f
C1412 VP.n68 VSUBS 0.043748f
C1413 VP.n69 VSUBS 0.042148f
C1414 VP.n70 VSUBS 0.023591f
C1415 VP.n71 VSUBS 0.023591f
C1416 VP.n72 VSUBS 0.023591f
C1417 VP.n73 VSUBS 0.046414f
C1418 VP.n74 VSUBS 0.043748f
C1419 VP.n75 VSUBS 0.029493f
C1420 VP.n76 VSUBS 0.023591f
C1421 VP.n77 VSUBS 0.023591f
C1422 VP.n78 VSUBS 0.036405f
C1423 VP.n79 VSUBS 0.043748f
C1424 VP.n80 VSUBS 0.045484f
C1425 VP.n81 VSUBS 0.023591f
C1426 VP.n82 VSUBS 0.023591f
C1427 VP.n83 VSUBS 0.023591f
C1428 VP.n84 VSUBS 0.047311f
C1429 VP.n85 VSUBS 0.043748f
C1430 VP.n86 VSUBS 0.032949f
C1431 VP.n87 VSUBS 0.023591f
C1432 VP.n88 VSUBS 0.023591f
C1433 VP.n89 VSUBS 0.032949f
C1434 VP.n90 VSUBS 0.043748f
C1435 VP.n91 VSUBS 0.047311f
C1436 VP.n92 VSUBS 0.023591f
C1437 VP.n93 VSUBS 0.023591f
C1438 VP.n94 VSUBS 0.023591f
C1439 VP.n95 VSUBS 0.045484f
C1440 VP.n96 VSUBS 0.043748f
C1441 VP.n97 VSUBS 0.036405f
C1442 VP.n98 VSUBS 0.023591f
C1443 VP.n99 VSUBS 0.023591f
C1444 VP.n100 VSUBS 0.029493f
C1445 VP.n101 VSUBS 0.043748f
C1446 VP.n102 VSUBS 0.046414f
C1447 VP.n103 VSUBS 0.023591f
C1448 VP.n104 VSUBS 0.023591f
C1449 VP.n105 VSUBS 0.023591f
C1450 VP.n106 VSUBS 0.042148f
C1451 VP.n107 VSUBS 0.043748f
C1452 VP.n108 VSUBS 0.03986f
C1453 VP.n109 VSUBS 0.03807f
C1454 VP.n110 VSUBS 0.050921f
.ends

