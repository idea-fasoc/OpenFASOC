* NGSPICE file created from diff_pair_sample_1155.ext - technology: sky130A

.subckt diff_pair_sample_1155 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=4.914 pd=25.98 as=2.079 ps=12.93 w=12.6 l=0.41
X1 VDD1.t5 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=4.914 pd=25.98 as=2.079 ps=12.93 w=12.6 l=0.41
X2 VTAIL.t10 VN.t1 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.079 pd=12.93 as=2.079 ps=12.93 w=12.6 l=0.41
X3 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.914 pd=25.98 as=0 ps=0 w=12.6 l=0.41
X4 VTAIL.t1 VP.t1 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.079 pd=12.93 as=2.079 ps=12.93 w=12.6 l=0.41
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.914 pd=25.98 as=0 ps=0 w=12.6 l=0.41
X6 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.914 pd=25.98 as=0 ps=0 w=12.6 l=0.41
X7 VDD1.t3 VP.t2 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.079 pd=12.93 as=4.914 ps=25.98 w=12.6 l=0.41
X8 VDD2.t3 VN.t2 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=2.079 pd=12.93 as=4.914 ps=25.98 w=12.6 l=0.41
X9 VTAIL.t8 VN.t3 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.079 pd=12.93 as=2.079 ps=12.93 w=12.6 l=0.41
X10 VDD1.t2 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.079 pd=12.93 as=4.914 ps=25.98 w=12.6 l=0.41
X11 VDD2.t1 VN.t4 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=4.914 pd=25.98 as=2.079 ps=12.93 w=12.6 l=0.41
X12 VDD1.t1 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=4.914 pd=25.98 as=2.079 ps=12.93 w=12.6 l=0.41
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.914 pd=25.98 as=0 ps=0 w=12.6 l=0.41
X14 VDD2.t0 VN.t5 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.079 pd=12.93 as=4.914 ps=25.98 w=12.6 l=0.41
X15 VTAIL.t0 VP.t5 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.079 pd=12.93 as=2.079 ps=12.93 w=12.6 l=0.41
R0 VN.n0 VN.t4 860.577
R1 VN.n4 VN.t2 860.577
R2 VN.n2 VN.t5 841.558
R3 VN.n6 VN.t0 841.558
R4 VN.n1 VN.t1 836.447
R5 VN.n5 VN.t3 836.447
R6 VN.n3 VN.n2 161.3
R7 VN.n7 VN.n6 161.3
R8 VN.n7 VN.n4 71.3843
R9 VN.n3 VN.n0 71.3843
R10 VN.n2 VN.n1 43.0884
R11 VN.n6 VN.n5 43.0884
R12 VN VN.n7 40.9872
R13 VN.n5 VN.n4 18.9966
R14 VN.n1 VN.n0 18.9966
R15 VN VN.n3 0.0516364
R16 VTAIL.n286 VTAIL.n285 289.615
R17 VTAIL.n70 VTAIL.n69 289.615
R18 VTAIL.n216 VTAIL.n215 289.615
R19 VTAIL.n144 VTAIL.n143 289.615
R20 VTAIL.n240 VTAIL.n239 185
R21 VTAIL.n245 VTAIL.n244 185
R22 VTAIL.n247 VTAIL.n246 185
R23 VTAIL.n236 VTAIL.n235 185
R24 VTAIL.n253 VTAIL.n252 185
R25 VTAIL.n255 VTAIL.n254 185
R26 VTAIL.n232 VTAIL.n231 185
R27 VTAIL.n261 VTAIL.n260 185
R28 VTAIL.n263 VTAIL.n262 185
R29 VTAIL.n228 VTAIL.n227 185
R30 VTAIL.n269 VTAIL.n268 185
R31 VTAIL.n271 VTAIL.n270 185
R32 VTAIL.n224 VTAIL.n223 185
R33 VTAIL.n277 VTAIL.n276 185
R34 VTAIL.n279 VTAIL.n278 185
R35 VTAIL.n220 VTAIL.n219 185
R36 VTAIL.n285 VTAIL.n284 185
R37 VTAIL.n24 VTAIL.n23 185
R38 VTAIL.n29 VTAIL.n28 185
R39 VTAIL.n31 VTAIL.n30 185
R40 VTAIL.n20 VTAIL.n19 185
R41 VTAIL.n37 VTAIL.n36 185
R42 VTAIL.n39 VTAIL.n38 185
R43 VTAIL.n16 VTAIL.n15 185
R44 VTAIL.n45 VTAIL.n44 185
R45 VTAIL.n47 VTAIL.n46 185
R46 VTAIL.n12 VTAIL.n11 185
R47 VTAIL.n53 VTAIL.n52 185
R48 VTAIL.n55 VTAIL.n54 185
R49 VTAIL.n8 VTAIL.n7 185
R50 VTAIL.n61 VTAIL.n60 185
R51 VTAIL.n63 VTAIL.n62 185
R52 VTAIL.n4 VTAIL.n3 185
R53 VTAIL.n69 VTAIL.n68 185
R54 VTAIL.n215 VTAIL.n214 185
R55 VTAIL.n150 VTAIL.n149 185
R56 VTAIL.n209 VTAIL.n208 185
R57 VTAIL.n207 VTAIL.n206 185
R58 VTAIL.n154 VTAIL.n153 185
R59 VTAIL.n201 VTAIL.n200 185
R60 VTAIL.n199 VTAIL.n198 185
R61 VTAIL.n158 VTAIL.n157 185
R62 VTAIL.n193 VTAIL.n192 185
R63 VTAIL.n191 VTAIL.n190 185
R64 VTAIL.n162 VTAIL.n161 185
R65 VTAIL.n185 VTAIL.n184 185
R66 VTAIL.n183 VTAIL.n182 185
R67 VTAIL.n166 VTAIL.n165 185
R68 VTAIL.n177 VTAIL.n176 185
R69 VTAIL.n175 VTAIL.n174 185
R70 VTAIL.n170 VTAIL.n169 185
R71 VTAIL.n143 VTAIL.n142 185
R72 VTAIL.n78 VTAIL.n77 185
R73 VTAIL.n137 VTAIL.n136 185
R74 VTAIL.n135 VTAIL.n134 185
R75 VTAIL.n82 VTAIL.n81 185
R76 VTAIL.n129 VTAIL.n128 185
R77 VTAIL.n127 VTAIL.n126 185
R78 VTAIL.n86 VTAIL.n85 185
R79 VTAIL.n121 VTAIL.n120 185
R80 VTAIL.n119 VTAIL.n118 185
R81 VTAIL.n90 VTAIL.n89 185
R82 VTAIL.n113 VTAIL.n112 185
R83 VTAIL.n111 VTAIL.n110 185
R84 VTAIL.n94 VTAIL.n93 185
R85 VTAIL.n105 VTAIL.n104 185
R86 VTAIL.n103 VTAIL.n102 185
R87 VTAIL.n98 VTAIL.n97 185
R88 VTAIL.n241 VTAIL.t6 147.659
R89 VTAIL.n25 VTAIL.t2 147.659
R90 VTAIL.n171 VTAIL.t4 147.659
R91 VTAIL.n99 VTAIL.t7 147.659
R92 VTAIL.n245 VTAIL.n239 104.615
R93 VTAIL.n246 VTAIL.n245 104.615
R94 VTAIL.n246 VTAIL.n235 104.615
R95 VTAIL.n253 VTAIL.n235 104.615
R96 VTAIL.n254 VTAIL.n253 104.615
R97 VTAIL.n254 VTAIL.n231 104.615
R98 VTAIL.n261 VTAIL.n231 104.615
R99 VTAIL.n262 VTAIL.n261 104.615
R100 VTAIL.n262 VTAIL.n227 104.615
R101 VTAIL.n269 VTAIL.n227 104.615
R102 VTAIL.n270 VTAIL.n269 104.615
R103 VTAIL.n270 VTAIL.n223 104.615
R104 VTAIL.n277 VTAIL.n223 104.615
R105 VTAIL.n278 VTAIL.n277 104.615
R106 VTAIL.n278 VTAIL.n219 104.615
R107 VTAIL.n285 VTAIL.n219 104.615
R108 VTAIL.n29 VTAIL.n23 104.615
R109 VTAIL.n30 VTAIL.n29 104.615
R110 VTAIL.n30 VTAIL.n19 104.615
R111 VTAIL.n37 VTAIL.n19 104.615
R112 VTAIL.n38 VTAIL.n37 104.615
R113 VTAIL.n38 VTAIL.n15 104.615
R114 VTAIL.n45 VTAIL.n15 104.615
R115 VTAIL.n46 VTAIL.n45 104.615
R116 VTAIL.n46 VTAIL.n11 104.615
R117 VTAIL.n53 VTAIL.n11 104.615
R118 VTAIL.n54 VTAIL.n53 104.615
R119 VTAIL.n54 VTAIL.n7 104.615
R120 VTAIL.n61 VTAIL.n7 104.615
R121 VTAIL.n62 VTAIL.n61 104.615
R122 VTAIL.n62 VTAIL.n3 104.615
R123 VTAIL.n69 VTAIL.n3 104.615
R124 VTAIL.n215 VTAIL.n149 104.615
R125 VTAIL.n208 VTAIL.n149 104.615
R126 VTAIL.n208 VTAIL.n207 104.615
R127 VTAIL.n207 VTAIL.n153 104.615
R128 VTAIL.n200 VTAIL.n153 104.615
R129 VTAIL.n200 VTAIL.n199 104.615
R130 VTAIL.n199 VTAIL.n157 104.615
R131 VTAIL.n192 VTAIL.n157 104.615
R132 VTAIL.n192 VTAIL.n191 104.615
R133 VTAIL.n191 VTAIL.n161 104.615
R134 VTAIL.n184 VTAIL.n161 104.615
R135 VTAIL.n184 VTAIL.n183 104.615
R136 VTAIL.n183 VTAIL.n165 104.615
R137 VTAIL.n176 VTAIL.n165 104.615
R138 VTAIL.n176 VTAIL.n175 104.615
R139 VTAIL.n175 VTAIL.n169 104.615
R140 VTAIL.n143 VTAIL.n77 104.615
R141 VTAIL.n136 VTAIL.n77 104.615
R142 VTAIL.n136 VTAIL.n135 104.615
R143 VTAIL.n135 VTAIL.n81 104.615
R144 VTAIL.n128 VTAIL.n81 104.615
R145 VTAIL.n128 VTAIL.n127 104.615
R146 VTAIL.n127 VTAIL.n85 104.615
R147 VTAIL.n120 VTAIL.n85 104.615
R148 VTAIL.n120 VTAIL.n119 104.615
R149 VTAIL.n119 VTAIL.n89 104.615
R150 VTAIL.n112 VTAIL.n89 104.615
R151 VTAIL.n112 VTAIL.n111 104.615
R152 VTAIL.n111 VTAIL.n93 104.615
R153 VTAIL.n104 VTAIL.n93 104.615
R154 VTAIL.n104 VTAIL.n103 104.615
R155 VTAIL.n103 VTAIL.n97 104.615
R156 VTAIL.t6 VTAIL.n239 52.3082
R157 VTAIL.t2 VTAIL.n23 52.3082
R158 VTAIL.t4 VTAIL.n169 52.3082
R159 VTAIL.t7 VTAIL.n97 52.3082
R160 VTAIL.n147 VTAIL.n146 46.8569
R161 VTAIL.n75 VTAIL.n74 46.8569
R162 VTAIL.n1 VTAIL.n0 46.8559
R163 VTAIL.n73 VTAIL.n72 46.8559
R164 VTAIL.n287 VTAIL.n286 34.1247
R165 VTAIL.n71 VTAIL.n70 34.1247
R166 VTAIL.n217 VTAIL.n216 34.1247
R167 VTAIL.n145 VTAIL.n144 34.1247
R168 VTAIL.n75 VTAIL.n73 24.5048
R169 VTAIL.n287 VTAIL.n217 23.8669
R170 VTAIL.n241 VTAIL.n240 15.6677
R171 VTAIL.n25 VTAIL.n24 15.6677
R172 VTAIL.n171 VTAIL.n170 15.6677
R173 VTAIL.n99 VTAIL.n98 15.6677
R174 VTAIL.n244 VTAIL.n243 12.8005
R175 VTAIL.n284 VTAIL.n218 12.8005
R176 VTAIL.n28 VTAIL.n27 12.8005
R177 VTAIL.n68 VTAIL.n2 12.8005
R178 VTAIL.n214 VTAIL.n148 12.8005
R179 VTAIL.n174 VTAIL.n173 12.8005
R180 VTAIL.n142 VTAIL.n76 12.8005
R181 VTAIL.n102 VTAIL.n101 12.8005
R182 VTAIL.n247 VTAIL.n238 12.0247
R183 VTAIL.n283 VTAIL.n220 12.0247
R184 VTAIL.n31 VTAIL.n22 12.0247
R185 VTAIL.n67 VTAIL.n4 12.0247
R186 VTAIL.n213 VTAIL.n150 12.0247
R187 VTAIL.n177 VTAIL.n168 12.0247
R188 VTAIL.n141 VTAIL.n78 12.0247
R189 VTAIL.n105 VTAIL.n96 12.0247
R190 VTAIL.n248 VTAIL.n236 11.249
R191 VTAIL.n280 VTAIL.n279 11.249
R192 VTAIL.n32 VTAIL.n20 11.249
R193 VTAIL.n64 VTAIL.n63 11.249
R194 VTAIL.n210 VTAIL.n209 11.249
R195 VTAIL.n178 VTAIL.n166 11.249
R196 VTAIL.n138 VTAIL.n137 11.249
R197 VTAIL.n106 VTAIL.n94 11.249
R198 VTAIL.n252 VTAIL.n251 10.4732
R199 VTAIL.n276 VTAIL.n222 10.4732
R200 VTAIL.n36 VTAIL.n35 10.4732
R201 VTAIL.n60 VTAIL.n6 10.4732
R202 VTAIL.n206 VTAIL.n152 10.4732
R203 VTAIL.n182 VTAIL.n181 10.4732
R204 VTAIL.n134 VTAIL.n80 10.4732
R205 VTAIL.n110 VTAIL.n109 10.4732
R206 VTAIL.n255 VTAIL.n234 9.69747
R207 VTAIL.n275 VTAIL.n224 9.69747
R208 VTAIL.n39 VTAIL.n18 9.69747
R209 VTAIL.n59 VTAIL.n8 9.69747
R210 VTAIL.n205 VTAIL.n154 9.69747
R211 VTAIL.n185 VTAIL.n164 9.69747
R212 VTAIL.n133 VTAIL.n82 9.69747
R213 VTAIL.n113 VTAIL.n92 9.69747
R214 VTAIL.n282 VTAIL.n218 9.45567
R215 VTAIL.n66 VTAIL.n2 9.45567
R216 VTAIL.n212 VTAIL.n148 9.45567
R217 VTAIL.n140 VTAIL.n76 9.45567
R218 VTAIL.n265 VTAIL.n264 9.3005
R219 VTAIL.n267 VTAIL.n266 9.3005
R220 VTAIL.n226 VTAIL.n225 9.3005
R221 VTAIL.n273 VTAIL.n272 9.3005
R222 VTAIL.n275 VTAIL.n274 9.3005
R223 VTAIL.n222 VTAIL.n221 9.3005
R224 VTAIL.n281 VTAIL.n280 9.3005
R225 VTAIL.n283 VTAIL.n282 9.3005
R226 VTAIL.n259 VTAIL.n258 9.3005
R227 VTAIL.n257 VTAIL.n256 9.3005
R228 VTAIL.n234 VTAIL.n233 9.3005
R229 VTAIL.n251 VTAIL.n250 9.3005
R230 VTAIL.n249 VTAIL.n248 9.3005
R231 VTAIL.n238 VTAIL.n237 9.3005
R232 VTAIL.n243 VTAIL.n242 9.3005
R233 VTAIL.n230 VTAIL.n229 9.3005
R234 VTAIL.n49 VTAIL.n48 9.3005
R235 VTAIL.n51 VTAIL.n50 9.3005
R236 VTAIL.n10 VTAIL.n9 9.3005
R237 VTAIL.n57 VTAIL.n56 9.3005
R238 VTAIL.n59 VTAIL.n58 9.3005
R239 VTAIL.n6 VTAIL.n5 9.3005
R240 VTAIL.n65 VTAIL.n64 9.3005
R241 VTAIL.n67 VTAIL.n66 9.3005
R242 VTAIL.n43 VTAIL.n42 9.3005
R243 VTAIL.n41 VTAIL.n40 9.3005
R244 VTAIL.n18 VTAIL.n17 9.3005
R245 VTAIL.n35 VTAIL.n34 9.3005
R246 VTAIL.n33 VTAIL.n32 9.3005
R247 VTAIL.n22 VTAIL.n21 9.3005
R248 VTAIL.n27 VTAIL.n26 9.3005
R249 VTAIL.n14 VTAIL.n13 9.3005
R250 VTAIL.n213 VTAIL.n212 9.3005
R251 VTAIL.n211 VTAIL.n210 9.3005
R252 VTAIL.n152 VTAIL.n151 9.3005
R253 VTAIL.n205 VTAIL.n204 9.3005
R254 VTAIL.n203 VTAIL.n202 9.3005
R255 VTAIL.n156 VTAIL.n155 9.3005
R256 VTAIL.n197 VTAIL.n196 9.3005
R257 VTAIL.n195 VTAIL.n194 9.3005
R258 VTAIL.n160 VTAIL.n159 9.3005
R259 VTAIL.n189 VTAIL.n188 9.3005
R260 VTAIL.n187 VTAIL.n186 9.3005
R261 VTAIL.n164 VTAIL.n163 9.3005
R262 VTAIL.n181 VTAIL.n180 9.3005
R263 VTAIL.n179 VTAIL.n178 9.3005
R264 VTAIL.n168 VTAIL.n167 9.3005
R265 VTAIL.n173 VTAIL.n172 9.3005
R266 VTAIL.n125 VTAIL.n124 9.3005
R267 VTAIL.n84 VTAIL.n83 9.3005
R268 VTAIL.n131 VTAIL.n130 9.3005
R269 VTAIL.n133 VTAIL.n132 9.3005
R270 VTAIL.n80 VTAIL.n79 9.3005
R271 VTAIL.n139 VTAIL.n138 9.3005
R272 VTAIL.n141 VTAIL.n140 9.3005
R273 VTAIL.n123 VTAIL.n122 9.3005
R274 VTAIL.n88 VTAIL.n87 9.3005
R275 VTAIL.n117 VTAIL.n116 9.3005
R276 VTAIL.n115 VTAIL.n114 9.3005
R277 VTAIL.n92 VTAIL.n91 9.3005
R278 VTAIL.n109 VTAIL.n108 9.3005
R279 VTAIL.n107 VTAIL.n106 9.3005
R280 VTAIL.n96 VTAIL.n95 9.3005
R281 VTAIL.n101 VTAIL.n100 9.3005
R282 VTAIL.n256 VTAIL.n232 8.92171
R283 VTAIL.n272 VTAIL.n271 8.92171
R284 VTAIL.n40 VTAIL.n16 8.92171
R285 VTAIL.n56 VTAIL.n55 8.92171
R286 VTAIL.n202 VTAIL.n201 8.92171
R287 VTAIL.n186 VTAIL.n162 8.92171
R288 VTAIL.n130 VTAIL.n129 8.92171
R289 VTAIL.n114 VTAIL.n90 8.92171
R290 VTAIL.n260 VTAIL.n259 8.14595
R291 VTAIL.n268 VTAIL.n226 8.14595
R292 VTAIL.n44 VTAIL.n43 8.14595
R293 VTAIL.n52 VTAIL.n10 8.14595
R294 VTAIL.n198 VTAIL.n156 8.14595
R295 VTAIL.n190 VTAIL.n189 8.14595
R296 VTAIL.n126 VTAIL.n84 8.14595
R297 VTAIL.n118 VTAIL.n117 8.14595
R298 VTAIL.n263 VTAIL.n230 7.3702
R299 VTAIL.n267 VTAIL.n228 7.3702
R300 VTAIL.n47 VTAIL.n14 7.3702
R301 VTAIL.n51 VTAIL.n12 7.3702
R302 VTAIL.n197 VTAIL.n158 7.3702
R303 VTAIL.n193 VTAIL.n160 7.3702
R304 VTAIL.n125 VTAIL.n86 7.3702
R305 VTAIL.n121 VTAIL.n88 7.3702
R306 VTAIL.n264 VTAIL.n263 6.59444
R307 VTAIL.n264 VTAIL.n228 6.59444
R308 VTAIL.n48 VTAIL.n47 6.59444
R309 VTAIL.n48 VTAIL.n12 6.59444
R310 VTAIL.n194 VTAIL.n158 6.59444
R311 VTAIL.n194 VTAIL.n193 6.59444
R312 VTAIL.n122 VTAIL.n86 6.59444
R313 VTAIL.n122 VTAIL.n121 6.59444
R314 VTAIL.n260 VTAIL.n230 5.81868
R315 VTAIL.n268 VTAIL.n267 5.81868
R316 VTAIL.n44 VTAIL.n14 5.81868
R317 VTAIL.n52 VTAIL.n51 5.81868
R318 VTAIL.n198 VTAIL.n197 5.81868
R319 VTAIL.n190 VTAIL.n160 5.81868
R320 VTAIL.n126 VTAIL.n125 5.81868
R321 VTAIL.n118 VTAIL.n88 5.81868
R322 VTAIL.n259 VTAIL.n232 5.04292
R323 VTAIL.n271 VTAIL.n226 5.04292
R324 VTAIL.n43 VTAIL.n16 5.04292
R325 VTAIL.n55 VTAIL.n10 5.04292
R326 VTAIL.n201 VTAIL.n156 5.04292
R327 VTAIL.n189 VTAIL.n162 5.04292
R328 VTAIL.n129 VTAIL.n84 5.04292
R329 VTAIL.n117 VTAIL.n90 5.04292
R330 VTAIL.n242 VTAIL.n241 4.38563
R331 VTAIL.n26 VTAIL.n25 4.38563
R332 VTAIL.n172 VTAIL.n171 4.38563
R333 VTAIL.n100 VTAIL.n99 4.38563
R334 VTAIL.n256 VTAIL.n255 4.26717
R335 VTAIL.n272 VTAIL.n224 4.26717
R336 VTAIL.n40 VTAIL.n39 4.26717
R337 VTAIL.n56 VTAIL.n8 4.26717
R338 VTAIL.n202 VTAIL.n154 4.26717
R339 VTAIL.n186 VTAIL.n185 4.26717
R340 VTAIL.n130 VTAIL.n82 4.26717
R341 VTAIL.n114 VTAIL.n113 4.26717
R342 VTAIL.n252 VTAIL.n234 3.49141
R343 VTAIL.n276 VTAIL.n275 3.49141
R344 VTAIL.n36 VTAIL.n18 3.49141
R345 VTAIL.n60 VTAIL.n59 3.49141
R346 VTAIL.n206 VTAIL.n205 3.49141
R347 VTAIL.n182 VTAIL.n164 3.49141
R348 VTAIL.n134 VTAIL.n133 3.49141
R349 VTAIL.n110 VTAIL.n92 3.49141
R350 VTAIL.n251 VTAIL.n236 2.71565
R351 VTAIL.n279 VTAIL.n222 2.71565
R352 VTAIL.n35 VTAIL.n20 2.71565
R353 VTAIL.n63 VTAIL.n6 2.71565
R354 VTAIL.n209 VTAIL.n152 2.71565
R355 VTAIL.n181 VTAIL.n166 2.71565
R356 VTAIL.n137 VTAIL.n80 2.71565
R357 VTAIL.n109 VTAIL.n94 2.71565
R358 VTAIL.n248 VTAIL.n247 1.93989
R359 VTAIL.n280 VTAIL.n220 1.93989
R360 VTAIL.n32 VTAIL.n31 1.93989
R361 VTAIL.n64 VTAIL.n4 1.93989
R362 VTAIL.n210 VTAIL.n150 1.93989
R363 VTAIL.n178 VTAIL.n177 1.93989
R364 VTAIL.n138 VTAIL.n78 1.93989
R365 VTAIL.n106 VTAIL.n105 1.93989
R366 VTAIL.n0 VTAIL.t11 1.57193
R367 VTAIL.n0 VTAIL.t10 1.57193
R368 VTAIL.n72 VTAIL.t3 1.57193
R369 VTAIL.n72 VTAIL.t0 1.57193
R370 VTAIL.n146 VTAIL.t5 1.57193
R371 VTAIL.n146 VTAIL.t1 1.57193
R372 VTAIL.n74 VTAIL.t9 1.57193
R373 VTAIL.n74 VTAIL.t8 1.57193
R374 VTAIL.n244 VTAIL.n238 1.16414
R375 VTAIL.n284 VTAIL.n283 1.16414
R376 VTAIL.n28 VTAIL.n22 1.16414
R377 VTAIL.n68 VTAIL.n67 1.16414
R378 VTAIL.n214 VTAIL.n213 1.16414
R379 VTAIL.n174 VTAIL.n168 1.16414
R380 VTAIL.n142 VTAIL.n141 1.16414
R381 VTAIL.n102 VTAIL.n96 1.16414
R382 VTAIL.n147 VTAIL.n145 0.789293
R383 VTAIL.n71 VTAIL.n1 0.789293
R384 VTAIL.n145 VTAIL.n75 0.638431
R385 VTAIL.n217 VTAIL.n147 0.638431
R386 VTAIL.n73 VTAIL.n71 0.638431
R387 VTAIL VTAIL.n287 0.420759
R388 VTAIL.n243 VTAIL.n240 0.388379
R389 VTAIL.n286 VTAIL.n218 0.388379
R390 VTAIL.n27 VTAIL.n24 0.388379
R391 VTAIL.n70 VTAIL.n2 0.388379
R392 VTAIL.n216 VTAIL.n148 0.388379
R393 VTAIL.n173 VTAIL.n170 0.388379
R394 VTAIL.n144 VTAIL.n76 0.388379
R395 VTAIL.n101 VTAIL.n98 0.388379
R396 VTAIL VTAIL.n1 0.218172
R397 VTAIL.n242 VTAIL.n237 0.155672
R398 VTAIL.n249 VTAIL.n237 0.155672
R399 VTAIL.n250 VTAIL.n249 0.155672
R400 VTAIL.n250 VTAIL.n233 0.155672
R401 VTAIL.n257 VTAIL.n233 0.155672
R402 VTAIL.n258 VTAIL.n257 0.155672
R403 VTAIL.n258 VTAIL.n229 0.155672
R404 VTAIL.n265 VTAIL.n229 0.155672
R405 VTAIL.n266 VTAIL.n265 0.155672
R406 VTAIL.n266 VTAIL.n225 0.155672
R407 VTAIL.n273 VTAIL.n225 0.155672
R408 VTAIL.n274 VTAIL.n273 0.155672
R409 VTAIL.n274 VTAIL.n221 0.155672
R410 VTAIL.n281 VTAIL.n221 0.155672
R411 VTAIL.n282 VTAIL.n281 0.155672
R412 VTAIL.n26 VTAIL.n21 0.155672
R413 VTAIL.n33 VTAIL.n21 0.155672
R414 VTAIL.n34 VTAIL.n33 0.155672
R415 VTAIL.n34 VTAIL.n17 0.155672
R416 VTAIL.n41 VTAIL.n17 0.155672
R417 VTAIL.n42 VTAIL.n41 0.155672
R418 VTAIL.n42 VTAIL.n13 0.155672
R419 VTAIL.n49 VTAIL.n13 0.155672
R420 VTAIL.n50 VTAIL.n49 0.155672
R421 VTAIL.n50 VTAIL.n9 0.155672
R422 VTAIL.n57 VTAIL.n9 0.155672
R423 VTAIL.n58 VTAIL.n57 0.155672
R424 VTAIL.n58 VTAIL.n5 0.155672
R425 VTAIL.n65 VTAIL.n5 0.155672
R426 VTAIL.n66 VTAIL.n65 0.155672
R427 VTAIL.n212 VTAIL.n211 0.155672
R428 VTAIL.n211 VTAIL.n151 0.155672
R429 VTAIL.n204 VTAIL.n151 0.155672
R430 VTAIL.n204 VTAIL.n203 0.155672
R431 VTAIL.n203 VTAIL.n155 0.155672
R432 VTAIL.n196 VTAIL.n155 0.155672
R433 VTAIL.n196 VTAIL.n195 0.155672
R434 VTAIL.n195 VTAIL.n159 0.155672
R435 VTAIL.n188 VTAIL.n159 0.155672
R436 VTAIL.n188 VTAIL.n187 0.155672
R437 VTAIL.n187 VTAIL.n163 0.155672
R438 VTAIL.n180 VTAIL.n163 0.155672
R439 VTAIL.n180 VTAIL.n179 0.155672
R440 VTAIL.n179 VTAIL.n167 0.155672
R441 VTAIL.n172 VTAIL.n167 0.155672
R442 VTAIL.n140 VTAIL.n139 0.155672
R443 VTAIL.n139 VTAIL.n79 0.155672
R444 VTAIL.n132 VTAIL.n79 0.155672
R445 VTAIL.n132 VTAIL.n131 0.155672
R446 VTAIL.n131 VTAIL.n83 0.155672
R447 VTAIL.n124 VTAIL.n83 0.155672
R448 VTAIL.n124 VTAIL.n123 0.155672
R449 VTAIL.n123 VTAIL.n87 0.155672
R450 VTAIL.n116 VTAIL.n87 0.155672
R451 VTAIL.n116 VTAIL.n115 0.155672
R452 VTAIL.n115 VTAIL.n91 0.155672
R453 VTAIL.n108 VTAIL.n91 0.155672
R454 VTAIL.n108 VTAIL.n107 0.155672
R455 VTAIL.n107 VTAIL.n95 0.155672
R456 VTAIL.n100 VTAIL.n95 0.155672
R457 VDD2.n139 VDD2.n138 289.615
R458 VDD2.n68 VDD2.n67 289.615
R459 VDD2.n138 VDD2.n137 185
R460 VDD2.n73 VDD2.n72 185
R461 VDD2.n132 VDD2.n131 185
R462 VDD2.n130 VDD2.n129 185
R463 VDD2.n77 VDD2.n76 185
R464 VDD2.n124 VDD2.n123 185
R465 VDD2.n122 VDD2.n121 185
R466 VDD2.n81 VDD2.n80 185
R467 VDD2.n116 VDD2.n115 185
R468 VDD2.n114 VDD2.n113 185
R469 VDD2.n85 VDD2.n84 185
R470 VDD2.n108 VDD2.n107 185
R471 VDD2.n106 VDD2.n105 185
R472 VDD2.n89 VDD2.n88 185
R473 VDD2.n100 VDD2.n99 185
R474 VDD2.n98 VDD2.n97 185
R475 VDD2.n93 VDD2.n92 185
R476 VDD2.n22 VDD2.n21 185
R477 VDD2.n27 VDD2.n26 185
R478 VDD2.n29 VDD2.n28 185
R479 VDD2.n18 VDD2.n17 185
R480 VDD2.n35 VDD2.n34 185
R481 VDD2.n37 VDD2.n36 185
R482 VDD2.n14 VDD2.n13 185
R483 VDD2.n43 VDD2.n42 185
R484 VDD2.n45 VDD2.n44 185
R485 VDD2.n10 VDD2.n9 185
R486 VDD2.n51 VDD2.n50 185
R487 VDD2.n53 VDD2.n52 185
R488 VDD2.n6 VDD2.n5 185
R489 VDD2.n59 VDD2.n58 185
R490 VDD2.n61 VDD2.n60 185
R491 VDD2.n2 VDD2.n1 185
R492 VDD2.n67 VDD2.n66 185
R493 VDD2.n23 VDD2.t1 147.659
R494 VDD2.n94 VDD2.t5 147.659
R495 VDD2.n138 VDD2.n72 104.615
R496 VDD2.n131 VDD2.n72 104.615
R497 VDD2.n131 VDD2.n130 104.615
R498 VDD2.n130 VDD2.n76 104.615
R499 VDD2.n123 VDD2.n76 104.615
R500 VDD2.n123 VDD2.n122 104.615
R501 VDD2.n122 VDD2.n80 104.615
R502 VDD2.n115 VDD2.n80 104.615
R503 VDD2.n115 VDD2.n114 104.615
R504 VDD2.n114 VDD2.n84 104.615
R505 VDD2.n107 VDD2.n84 104.615
R506 VDD2.n107 VDD2.n106 104.615
R507 VDD2.n106 VDD2.n88 104.615
R508 VDD2.n99 VDD2.n88 104.615
R509 VDD2.n99 VDD2.n98 104.615
R510 VDD2.n98 VDD2.n92 104.615
R511 VDD2.n27 VDD2.n21 104.615
R512 VDD2.n28 VDD2.n27 104.615
R513 VDD2.n28 VDD2.n17 104.615
R514 VDD2.n35 VDD2.n17 104.615
R515 VDD2.n36 VDD2.n35 104.615
R516 VDD2.n36 VDD2.n13 104.615
R517 VDD2.n43 VDD2.n13 104.615
R518 VDD2.n44 VDD2.n43 104.615
R519 VDD2.n44 VDD2.n9 104.615
R520 VDD2.n51 VDD2.n9 104.615
R521 VDD2.n52 VDD2.n51 104.615
R522 VDD2.n52 VDD2.n5 104.615
R523 VDD2.n59 VDD2.n5 104.615
R524 VDD2.n60 VDD2.n59 104.615
R525 VDD2.n60 VDD2.n1 104.615
R526 VDD2.n67 VDD2.n1 104.615
R527 VDD2.n70 VDD2.n69 63.6388
R528 VDD2 VDD2.n141 63.636
R529 VDD2.t5 VDD2.n92 52.3082
R530 VDD2.t1 VDD2.n21 52.3082
R531 VDD2.n70 VDD2.n68 51.2266
R532 VDD2.n140 VDD2.n139 50.8035
R533 VDD2.n140 VDD2.n70 36.6506
R534 VDD2.n94 VDD2.n93 15.6677
R535 VDD2.n23 VDD2.n22 15.6677
R536 VDD2.n137 VDD2.n71 12.8005
R537 VDD2.n97 VDD2.n96 12.8005
R538 VDD2.n26 VDD2.n25 12.8005
R539 VDD2.n66 VDD2.n0 12.8005
R540 VDD2.n136 VDD2.n73 12.0247
R541 VDD2.n100 VDD2.n91 12.0247
R542 VDD2.n29 VDD2.n20 12.0247
R543 VDD2.n65 VDD2.n2 12.0247
R544 VDD2.n133 VDD2.n132 11.249
R545 VDD2.n101 VDD2.n89 11.249
R546 VDD2.n30 VDD2.n18 11.249
R547 VDD2.n62 VDD2.n61 11.249
R548 VDD2.n129 VDD2.n75 10.4732
R549 VDD2.n105 VDD2.n104 10.4732
R550 VDD2.n34 VDD2.n33 10.4732
R551 VDD2.n58 VDD2.n4 10.4732
R552 VDD2.n128 VDD2.n77 9.69747
R553 VDD2.n108 VDD2.n87 9.69747
R554 VDD2.n37 VDD2.n16 9.69747
R555 VDD2.n57 VDD2.n6 9.69747
R556 VDD2.n135 VDD2.n71 9.45567
R557 VDD2.n64 VDD2.n0 9.45567
R558 VDD2.n120 VDD2.n119 9.3005
R559 VDD2.n79 VDD2.n78 9.3005
R560 VDD2.n126 VDD2.n125 9.3005
R561 VDD2.n128 VDD2.n127 9.3005
R562 VDD2.n75 VDD2.n74 9.3005
R563 VDD2.n134 VDD2.n133 9.3005
R564 VDD2.n136 VDD2.n135 9.3005
R565 VDD2.n118 VDD2.n117 9.3005
R566 VDD2.n83 VDD2.n82 9.3005
R567 VDD2.n112 VDD2.n111 9.3005
R568 VDD2.n110 VDD2.n109 9.3005
R569 VDD2.n87 VDD2.n86 9.3005
R570 VDD2.n104 VDD2.n103 9.3005
R571 VDD2.n102 VDD2.n101 9.3005
R572 VDD2.n91 VDD2.n90 9.3005
R573 VDD2.n96 VDD2.n95 9.3005
R574 VDD2.n47 VDD2.n46 9.3005
R575 VDD2.n49 VDD2.n48 9.3005
R576 VDD2.n8 VDD2.n7 9.3005
R577 VDD2.n55 VDD2.n54 9.3005
R578 VDD2.n57 VDD2.n56 9.3005
R579 VDD2.n4 VDD2.n3 9.3005
R580 VDD2.n63 VDD2.n62 9.3005
R581 VDD2.n65 VDD2.n64 9.3005
R582 VDD2.n41 VDD2.n40 9.3005
R583 VDD2.n39 VDD2.n38 9.3005
R584 VDD2.n16 VDD2.n15 9.3005
R585 VDD2.n33 VDD2.n32 9.3005
R586 VDD2.n31 VDD2.n30 9.3005
R587 VDD2.n20 VDD2.n19 9.3005
R588 VDD2.n25 VDD2.n24 9.3005
R589 VDD2.n12 VDD2.n11 9.3005
R590 VDD2.n125 VDD2.n124 8.92171
R591 VDD2.n109 VDD2.n85 8.92171
R592 VDD2.n38 VDD2.n14 8.92171
R593 VDD2.n54 VDD2.n53 8.92171
R594 VDD2.n121 VDD2.n79 8.14595
R595 VDD2.n113 VDD2.n112 8.14595
R596 VDD2.n42 VDD2.n41 8.14595
R597 VDD2.n50 VDD2.n8 8.14595
R598 VDD2.n120 VDD2.n81 7.3702
R599 VDD2.n116 VDD2.n83 7.3702
R600 VDD2.n45 VDD2.n12 7.3702
R601 VDD2.n49 VDD2.n10 7.3702
R602 VDD2.n117 VDD2.n81 6.59444
R603 VDD2.n117 VDD2.n116 6.59444
R604 VDD2.n46 VDD2.n45 6.59444
R605 VDD2.n46 VDD2.n10 6.59444
R606 VDD2.n121 VDD2.n120 5.81868
R607 VDD2.n113 VDD2.n83 5.81868
R608 VDD2.n42 VDD2.n12 5.81868
R609 VDD2.n50 VDD2.n49 5.81868
R610 VDD2.n124 VDD2.n79 5.04292
R611 VDD2.n112 VDD2.n85 5.04292
R612 VDD2.n41 VDD2.n14 5.04292
R613 VDD2.n53 VDD2.n8 5.04292
R614 VDD2.n24 VDD2.n23 4.38563
R615 VDD2.n95 VDD2.n94 4.38563
R616 VDD2.n125 VDD2.n77 4.26717
R617 VDD2.n109 VDD2.n108 4.26717
R618 VDD2.n38 VDD2.n37 4.26717
R619 VDD2.n54 VDD2.n6 4.26717
R620 VDD2.n129 VDD2.n128 3.49141
R621 VDD2.n105 VDD2.n87 3.49141
R622 VDD2.n34 VDD2.n16 3.49141
R623 VDD2.n58 VDD2.n57 3.49141
R624 VDD2.n132 VDD2.n75 2.71565
R625 VDD2.n104 VDD2.n89 2.71565
R626 VDD2.n33 VDD2.n18 2.71565
R627 VDD2.n61 VDD2.n4 2.71565
R628 VDD2.n133 VDD2.n73 1.93989
R629 VDD2.n101 VDD2.n100 1.93989
R630 VDD2.n30 VDD2.n29 1.93989
R631 VDD2.n62 VDD2.n2 1.93989
R632 VDD2.n141 VDD2.t2 1.57193
R633 VDD2.n141 VDD2.t3 1.57193
R634 VDD2.n69 VDD2.t4 1.57193
R635 VDD2.n69 VDD2.t0 1.57193
R636 VDD2.n137 VDD2.n136 1.16414
R637 VDD2.n97 VDD2.n91 1.16414
R638 VDD2.n26 VDD2.n20 1.16414
R639 VDD2.n66 VDD2.n65 1.16414
R640 VDD2 VDD2.n140 0.537138
R641 VDD2.n139 VDD2.n71 0.388379
R642 VDD2.n96 VDD2.n93 0.388379
R643 VDD2.n25 VDD2.n22 0.388379
R644 VDD2.n68 VDD2.n0 0.388379
R645 VDD2.n135 VDD2.n134 0.155672
R646 VDD2.n134 VDD2.n74 0.155672
R647 VDD2.n127 VDD2.n74 0.155672
R648 VDD2.n127 VDD2.n126 0.155672
R649 VDD2.n126 VDD2.n78 0.155672
R650 VDD2.n119 VDD2.n78 0.155672
R651 VDD2.n119 VDD2.n118 0.155672
R652 VDD2.n118 VDD2.n82 0.155672
R653 VDD2.n111 VDD2.n82 0.155672
R654 VDD2.n111 VDD2.n110 0.155672
R655 VDD2.n110 VDD2.n86 0.155672
R656 VDD2.n103 VDD2.n86 0.155672
R657 VDD2.n103 VDD2.n102 0.155672
R658 VDD2.n102 VDD2.n90 0.155672
R659 VDD2.n95 VDD2.n90 0.155672
R660 VDD2.n24 VDD2.n19 0.155672
R661 VDD2.n31 VDD2.n19 0.155672
R662 VDD2.n32 VDD2.n31 0.155672
R663 VDD2.n32 VDD2.n15 0.155672
R664 VDD2.n39 VDD2.n15 0.155672
R665 VDD2.n40 VDD2.n39 0.155672
R666 VDD2.n40 VDD2.n11 0.155672
R667 VDD2.n47 VDD2.n11 0.155672
R668 VDD2.n48 VDD2.n47 0.155672
R669 VDD2.n48 VDD2.n7 0.155672
R670 VDD2.n55 VDD2.n7 0.155672
R671 VDD2.n56 VDD2.n55 0.155672
R672 VDD2.n56 VDD2.n3 0.155672
R673 VDD2.n63 VDD2.n3 0.155672
R674 VDD2.n64 VDD2.n63 0.155672
R675 B.n362 B.t10 949.688
R676 B.n359 B.t6 949.688
R677 B.n85 B.t17 949.688
R678 B.n83 B.t13 949.688
R679 B.n629 B.n628 585
R680 B.n277 B.n82 585
R681 B.n276 B.n275 585
R682 B.n274 B.n273 585
R683 B.n272 B.n271 585
R684 B.n270 B.n269 585
R685 B.n268 B.n267 585
R686 B.n266 B.n265 585
R687 B.n264 B.n263 585
R688 B.n262 B.n261 585
R689 B.n260 B.n259 585
R690 B.n258 B.n257 585
R691 B.n256 B.n255 585
R692 B.n254 B.n253 585
R693 B.n252 B.n251 585
R694 B.n250 B.n249 585
R695 B.n248 B.n247 585
R696 B.n246 B.n245 585
R697 B.n244 B.n243 585
R698 B.n242 B.n241 585
R699 B.n240 B.n239 585
R700 B.n238 B.n237 585
R701 B.n236 B.n235 585
R702 B.n234 B.n233 585
R703 B.n232 B.n231 585
R704 B.n230 B.n229 585
R705 B.n228 B.n227 585
R706 B.n226 B.n225 585
R707 B.n224 B.n223 585
R708 B.n222 B.n221 585
R709 B.n220 B.n219 585
R710 B.n218 B.n217 585
R711 B.n216 B.n215 585
R712 B.n214 B.n213 585
R713 B.n212 B.n211 585
R714 B.n210 B.n209 585
R715 B.n208 B.n207 585
R716 B.n206 B.n205 585
R717 B.n204 B.n203 585
R718 B.n202 B.n201 585
R719 B.n200 B.n199 585
R720 B.n198 B.n197 585
R721 B.n196 B.n195 585
R722 B.n193 B.n192 585
R723 B.n191 B.n190 585
R724 B.n189 B.n188 585
R725 B.n187 B.n186 585
R726 B.n185 B.n184 585
R727 B.n183 B.n182 585
R728 B.n181 B.n180 585
R729 B.n179 B.n178 585
R730 B.n177 B.n176 585
R731 B.n175 B.n174 585
R732 B.n172 B.n171 585
R733 B.n170 B.n169 585
R734 B.n168 B.n167 585
R735 B.n166 B.n165 585
R736 B.n164 B.n163 585
R737 B.n162 B.n161 585
R738 B.n160 B.n159 585
R739 B.n158 B.n157 585
R740 B.n156 B.n155 585
R741 B.n154 B.n153 585
R742 B.n152 B.n151 585
R743 B.n150 B.n149 585
R744 B.n148 B.n147 585
R745 B.n146 B.n145 585
R746 B.n144 B.n143 585
R747 B.n142 B.n141 585
R748 B.n140 B.n139 585
R749 B.n138 B.n137 585
R750 B.n136 B.n135 585
R751 B.n134 B.n133 585
R752 B.n132 B.n131 585
R753 B.n130 B.n129 585
R754 B.n128 B.n127 585
R755 B.n126 B.n125 585
R756 B.n124 B.n123 585
R757 B.n122 B.n121 585
R758 B.n120 B.n119 585
R759 B.n118 B.n117 585
R760 B.n116 B.n115 585
R761 B.n114 B.n113 585
R762 B.n112 B.n111 585
R763 B.n110 B.n109 585
R764 B.n108 B.n107 585
R765 B.n106 B.n105 585
R766 B.n104 B.n103 585
R767 B.n102 B.n101 585
R768 B.n100 B.n99 585
R769 B.n98 B.n97 585
R770 B.n96 B.n95 585
R771 B.n94 B.n93 585
R772 B.n92 B.n91 585
R773 B.n90 B.n89 585
R774 B.n88 B.n87 585
R775 B.n627 B.n34 585
R776 B.n632 B.n34 585
R777 B.n626 B.n33 585
R778 B.n633 B.n33 585
R779 B.n625 B.n624 585
R780 B.n624 B.n29 585
R781 B.n623 B.n28 585
R782 B.n639 B.n28 585
R783 B.n622 B.n27 585
R784 B.n640 B.n27 585
R785 B.n621 B.n26 585
R786 B.n641 B.n26 585
R787 B.n620 B.n619 585
R788 B.n619 B.n22 585
R789 B.n618 B.n21 585
R790 B.n647 B.n21 585
R791 B.n617 B.n20 585
R792 B.n648 B.n20 585
R793 B.n616 B.n19 585
R794 B.n649 B.n19 585
R795 B.n615 B.n614 585
R796 B.n614 B.n15 585
R797 B.n613 B.n14 585
R798 B.n655 B.n14 585
R799 B.n612 B.n13 585
R800 B.n656 B.n13 585
R801 B.n611 B.n12 585
R802 B.n657 B.n12 585
R803 B.n610 B.n609 585
R804 B.n609 B.n11 585
R805 B.n608 B.n7 585
R806 B.n663 B.n7 585
R807 B.n607 B.n6 585
R808 B.n664 B.n6 585
R809 B.n606 B.n5 585
R810 B.n665 B.n5 585
R811 B.n605 B.n604 585
R812 B.n604 B.n4 585
R813 B.n603 B.n278 585
R814 B.n603 B.n602 585
R815 B.n592 B.n279 585
R816 B.n595 B.n279 585
R817 B.n594 B.n593 585
R818 B.n596 B.n594 585
R819 B.n591 B.n283 585
R820 B.n287 B.n283 585
R821 B.n590 B.n589 585
R822 B.n589 B.n588 585
R823 B.n285 B.n284 585
R824 B.n286 B.n285 585
R825 B.n581 B.n580 585
R826 B.n582 B.n581 585
R827 B.n579 B.n292 585
R828 B.n292 B.n291 585
R829 B.n578 B.n577 585
R830 B.n577 B.n576 585
R831 B.n294 B.n293 585
R832 B.n295 B.n294 585
R833 B.n569 B.n568 585
R834 B.n570 B.n569 585
R835 B.n567 B.n299 585
R836 B.n303 B.n299 585
R837 B.n566 B.n565 585
R838 B.n565 B.n564 585
R839 B.n301 B.n300 585
R840 B.n302 B.n301 585
R841 B.n557 B.n556 585
R842 B.n558 B.n557 585
R843 B.n555 B.n308 585
R844 B.n308 B.n307 585
R845 B.n550 B.n549 585
R846 B.n548 B.n358 585
R847 B.n547 B.n357 585
R848 B.n552 B.n357 585
R849 B.n546 B.n545 585
R850 B.n544 B.n543 585
R851 B.n542 B.n541 585
R852 B.n540 B.n539 585
R853 B.n538 B.n537 585
R854 B.n536 B.n535 585
R855 B.n534 B.n533 585
R856 B.n532 B.n531 585
R857 B.n530 B.n529 585
R858 B.n528 B.n527 585
R859 B.n526 B.n525 585
R860 B.n524 B.n523 585
R861 B.n522 B.n521 585
R862 B.n520 B.n519 585
R863 B.n518 B.n517 585
R864 B.n516 B.n515 585
R865 B.n514 B.n513 585
R866 B.n512 B.n511 585
R867 B.n510 B.n509 585
R868 B.n508 B.n507 585
R869 B.n506 B.n505 585
R870 B.n504 B.n503 585
R871 B.n502 B.n501 585
R872 B.n500 B.n499 585
R873 B.n498 B.n497 585
R874 B.n496 B.n495 585
R875 B.n494 B.n493 585
R876 B.n492 B.n491 585
R877 B.n490 B.n489 585
R878 B.n488 B.n487 585
R879 B.n486 B.n485 585
R880 B.n484 B.n483 585
R881 B.n482 B.n481 585
R882 B.n480 B.n479 585
R883 B.n478 B.n477 585
R884 B.n476 B.n475 585
R885 B.n474 B.n473 585
R886 B.n472 B.n471 585
R887 B.n470 B.n469 585
R888 B.n468 B.n467 585
R889 B.n466 B.n465 585
R890 B.n464 B.n463 585
R891 B.n462 B.n461 585
R892 B.n460 B.n459 585
R893 B.n458 B.n457 585
R894 B.n456 B.n455 585
R895 B.n454 B.n453 585
R896 B.n452 B.n451 585
R897 B.n450 B.n449 585
R898 B.n448 B.n447 585
R899 B.n446 B.n445 585
R900 B.n444 B.n443 585
R901 B.n442 B.n441 585
R902 B.n440 B.n439 585
R903 B.n438 B.n437 585
R904 B.n436 B.n435 585
R905 B.n434 B.n433 585
R906 B.n432 B.n431 585
R907 B.n430 B.n429 585
R908 B.n428 B.n427 585
R909 B.n426 B.n425 585
R910 B.n424 B.n423 585
R911 B.n422 B.n421 585
R912 B.n420 B.n419 585
R913 B.n418 B.n417 585
R914 B.n416 B.n415 585
R915 B.n414 B.n413 585
R916 B.n412 B.n411 585
R917 B.n410 B.n409 585
R918 B.n408 B.n407 585
R919 B.n406 B.n405 585
R920 B.n404 B.n403 585
R921 B.n402 B.n401 585
R922 B.n400 B.n399 585
R923 B.n398 B.n397 585
R924 B.n396 B.n395 585
R925 B.n394 B.n393 585
R926 B.n392 B.n391 585
R927 B.n390 B.n389 585
R928 B.n388 B.n387 585
R929 B.n386 B.n385 585
R930 B.n384 B.n383 585
R931 B.n382 B.n381 585
R932 B.n380 B.n379 585
R933 B.n378 B.n377 585
R934 B.n376 B.n375 585
R935 B.n374 B.n373 585
R936 B.n372 B.n371 585
R937 B.n370 B.n369 585
R938 B.n368 B.n367 585
R939 B.n366 B.n365 585
R940 B.n310 B.n309 585
R941 B.n554 B.n553 585
R942 B.n553 B.n552 585
R943 B.n306 B.n305 585
R944 B.n307 B.n306 585
R945 B.n560 B.n559 585
R946 B.n559 B.n558 585
R947 B.n561 B.n304 585
R948 B.n304 B.n302 585
R949 B.n563 B.n562 585
R950 B.n564 B.n563 585
R951 B.n298 B.n297 585
R952 B.n303 B.n298 585
R953 B.n572 B.n571 585
R954 B.n571 B.n570 585
R955 B.n573 B.n296 585
R956 B.n296 B.n295 585
R957 B.n575 B.n574 585
R958 B.n576 B.n575 585
R959 B.n290 B.n289 585
R960 B.n291 B.n290 585
R961 B.n584 B.n583 585
R962 B.n583 B.n582 585
R963 B.n585 B.n288 585
R964 B.n288 B.n286 585
R965 B.n587 B.n586 585
R966 B.n588 B.n587 585
R967 B.n282 B.n281 585
R968 B.n287 B.n282 585
R969 B.n598 B.n597 585
R970 B.n597 B.n596 585
R971 B.n599 B.n280 585
R972 B.n595 B.n280 585
R973 B.n601 B.n600 585
R974 B.n602 B.n601 585
R975 B.n2 B.n0 585
R976 B.n4 B.n2 585
R977 B.n3 B.n1 585
R978 B.n664 B.n3 585
R979 B.n662 B.n661 585
R980 B.n663 B.n662 585
R981 B.n660 B.n8 585
R982 B.n11 B.n8 585
R983 B.n659 B.n658 585
R984 B.n658 B.n657 585
R985 B.n10 B.n9 585
R986 B.n656 B.n10 585
R987 B.n654 B.n653 585
R988 B.n655 B.n654 585
R989 B.n652 B.n16 585
R990 B.n16 B.n15 585
R991 B.n651 B.n650 585
R992 B.n650 B.n649 585
R993 B.n18 B.n17 585
R994 B.n648 B.n18 585
R995 B.n646 B.n645 585
R996 B.n647 B.n646 585
R997 B.n644 B.n23 585
R998 B.n23 B.n22 585
R999 B.n643 B.n642 585
R1000 B.n642 B.n641 585
R1001 B.n25 B.n24 585
R1002 B.n640 B.n25 585
R1003 B.n638 B.n637 585
R1004 B.n639 B.n638 585
R1005 B.n636 B.n30 585
R1006 B.n30 B.n29 585
R1007 B.n635 B.n634 585
R1008 B.n634 B.n633 585
R1009 B.n32 B.n31 585
R1010 B.n632 B.n32 585
R1011 B.n667 B.n666 585
R1012 B.n666 B.n665 585
R1013 B.n550 B.n306 497.305
R1014 B.n87 B.n32 497.305
R1015 B.n553 B.n308 497.305
R1016 B.n629 B.n34 497.305
R1017 B.n362 B.t12 306.521
R1018 B.n83 B.t15 306.521
R1019 B.n359 B.t9 306.521
R1020 B.n85 B.t18 306.521
R1021 B.n363 B.t11 292.17
R1022 B.n84 B.t16 292.17
R1023 B.n360 B.t8 292.168
R1024 B.n86 B.t19 292.168
R1025 B.n631 B.n630 256.663
R1026 B.n631 B.n81 256.663
R1027 B.n631 B.n80 256.663
R1028 B.n631 B.n79 256.663
R1029 B.n631 B.n78 256.663
R1030 B.n631 B.n77 256.663
R1031 B.n631 B.n76 256.663
R1032 B.n631 B.n75 256.663
R1033 B.n631 B.n74 256.663
R1034 B.n631 B.n73 256.663
R1035 B.n631 B.n72 256.663
R1036 B.n631 B.n71 256.663
R1037 B.n631 B.n70 256.663
R1038 B.n631 B.n69 256.663
R1039 B.n631 B.n68 256.663
R1040 B.n631 B.n67 256.663
R1041 B.n631 B.n66 256.663
R1042 B.n631 B.n65 256.663
R1043 B.n631 B.n64 256.663
R1044 B.n631 B.n63 256.663
R1045 B.n631 B.n62 256.663
R1046 B.n631 B.n61 256.663
R1047 B.n631 B.n60 256.663
R1048 B.n631 B.n59 256.663
R1049 B.n631 B.n58 256.663
R1050 B.n631 B.n57 256.663
R1051 B.n631 B.n56 256.663
R1052 B.n631 B.n55 256.663
R1053 B.n631 B.n54 256.663
R1054 B.n631 B.n53 256.663
R1055 B.n631 B.n52 256.663
R1056 B.n631 B.n51 256.663
R1057 B.n631 B.n50 256.663
R1058 B.n631 B.n49 256.663
R1059 B.n631 B.n48 256.663
R1060 B.n631 B.n47 256.663
R1061 B.n631 B.n46 256.663
R1062 B.n631 B.n45 256.663
R1063 B.n631 B.n44 256.663
R1064 B.n631 B.n43 256.663
R1065 B.n631 B.n42 256.663
R1066 B.n631 B.n41 256.663
R1067 B.n631 B.n40 256.663
R1068 B.n631 B.n39 256.663
R1069 B.n631 B.n38 256.663
R1070 B.n631 B.n37 256.663
R1071 B.n631 B.n36 256.663
R1072 B.n631 B.n35 256.663
R1073 B.n552 B.n551 256.663
R1074 B.n552 B.n311 256.663
R1075 B.n552 B.n312 256.663
R1076 B.n552 B.n313 256.663
R1077 B.n552 B.n314 256.663
R1078 B.n552 B.n315 256.663
R1079 B.n552 B.n316 256.663
R1080 B.n552 B.n317 256.663
R1081 B.n552 B.n318 256.663
R1082 B.n552 B.n319 256.663
R1083 B.n552 B.n320 256.663
R1084 B.n552 B.n321 256.663
R1085 B.n552 B.n322 256.663
R1086 B.n552 B.n323 256.663
R1087 B.n552 B.n324 256.663
R1088 B.n552 B.n325 256.663
R1089 B.n552 B.n326 256.663
R1090 B.n552 B.n327 256.663
R1091 B.n552 B.n328 256.663
R1092 B.n552 B.n329 256.663
R1093 B.n552 B.n330 256.663
R1094 B.n552 B.n331 256.663
R1095 B.n552 B.n332 256.663
R1096 B.n552 B.n333 256.663
R1097 B.n552 B.n334 256.663
R1098 B.n552 B.n335 256.663
R1099 B.n552 B.n336 256.663
R1100 B.n552 B.n337 256.663
R1101 B.n552 B.n338 256.663
R1102 B.n552 B.n339 256.663
R1103 B.n552 B.n340 256.663
R1104 B.n552 B.n341 256.663
R1105 B.n552 B.n342 256.663
R1106 B.n552 B.n343 256.663
R1107 B.n552 B.n344 256.663
R1108 B.n552 B.n345 256.663
R1109 B.n552 B.n346 256.663
R1110 B.n552 B.n347 256.663
R1111 B.n552 B.n348 256.663
R1112 B.n552 B.n349 256.663
R1113 B.n552 B.n350 256.663
R1114 B.n552 B.n351 256.663
R1115 B.n552 B.n352 256.663
R1116 B.n552 B.n353 256.663
R1117 B.n552 B.n354 256.663
R1118 B.n552 B.n355 256.663
R1119 B.n552 B.n356 256.663
R1120 B.n559 B.n306 163.367
R1121 B.n559 B.n304 163.367
R1122 B.n563 B.n304 163.367
R1123 B.n563 B.n298 163.367
R1124 B.n571 B.n298 163.367
R1125 B.n571 B.n296 163.367
R1126 B.n575 B.n296 163.367
R1127 B.n575 B.n290 163.367
R1128 B.n583 B.n290 163.367
R1129 B.n583 B.n288 163.367
R1130 B.n587 B.n288 163.367
R1131 B.n587 B.n282 163.367
R1132 B.n597 B.n282 163.367
R1133 B.n597 B.n280 163.367
R1134 B.n601 B.n280 163.367
R1135 B.n601 B.n2 163.367
R1136 B.n666 B.n2 163.367
R1137 B.n666 B.n3 163.367
R1138 B.n662 B.n3 163.367
R1139 B.n662 B.n8 163.367
R1140 B.n658 B.n8 163.367
R1141 B.n658 B.n10 163.367
R1142 B.n654 B.n10 163.367
R1143 B.n654 B.n16 163.367
R1144 B.n650 B.n16 163.367
R1145 B.n650 B.n18 163.367
R1146 B.n646 B.n18 163.367
R1147 B.n646 B.n23 163.367
R1148 B.n642 B.n23 163.367
R1149 B.n642 B.n25 163.367
R1150 B.n638 B.n25 163.367
R1151 B.n638 B.n30 163.367
R1152 B.n634 B.n30 163.367
R1153 B.n634 B.n32 163.367
R1154 B.n358 B.n357 163.367
R1155 B.n545 B.n357 163.367
R1156 B.n543 B.n542 163.367
R1157 B.n539 B.n538 163.367
R1158 B.n535 B.n534 163.367
R1159 B.n531 B.n530 163.367
R1160 B.n527 B.n526 163.367
R1161 B.n523 B.n522 163.367
R1162 B.n519 B.n518 163.367
R1163 B.n515 B.n514 163.367
R1164 B.n511 B.n510 163.367
R1165 B.n507 B.n506 163.367
R1166 B.n503 B.n502 163.367
R1167 B.n499 B.n498 163.367
R1168 B.n495 B.n494 163.367
R1169 B.n491 B.n490 163.367
R1170 B.n487 B.n486 163.367
R1171 B.n483 B.n482 163.367
R1172 B.n479 B.n478 163.367
R1173 B.n475 B.n474 163.367
R1174 B.n471 B.n470 163.367
R1175 B.n467 B.n466 163.367
R1176 B.n463 B.n462 163.367
R1177 B.n459 B.n458 163.367
R1178 B.n455 B.n454 163.367
R1179 B.n451 B.n450 163.367
R1180 B.n447 B.n446 163.367
R1181 B.n443 B.n442 163.367
R1182 B.n439 B.n438 163.367
R1183 B.n435 B.n434 163.367
R1184 B.n431 B.n430 163.367
R1185 B.n427 B.n426 163.367
R1186 B.n423 B.n422 163.367
R1187 B.n419 B.n418 163.367
R1188 B.n415 B.n414 163.367
R1189 B.n411 B.n410 163.367
R1190 B.n407 B.n406 163.367
R1191 B.n403 B.n402 163.367
R1192 B.n399 B.n398 163.367
R1193 B.n395 B.n394 163.367
R1194 B.n391 B.n390 163.367
R1195 B.n387 B.n386 163.367
R1196 B.n383 B.n382 163.367
R1197 B.n379 B.n378 163.367
R1198 B.n375 B.n374 163.367
R1199 B.n371 B.n370 163.367
R1200 B.n367 B.n366 163.367
R1201 B.n553 B.n310 163.367
R1202 B.n557 B.n308 163.367
R1203 B.n557 B.n301 163.367
R1204 B.n565 B.n301 163.367
R1205 B.n565 B.n299 163.367
R1206 B.n569 B.n299 163.367
R1207 B.n569 B.n294 163.367
R1208 B.n577 B.n294 163.367
R1209 B.n577 B.n292 163.367
R1210 B.n581 B.n292 163.367
R1211 B.n581 B.n285 163.367
R1212 B.n589 B.n285 163.367
R1213 B.n589 B.n283 163.367
R1214 B.n594 B.n283 163.367
R1215 B.n594 B.n279 163.367
R1216 B.n603 B.n279 163.367
R1217 B.n604 B.n603 163.367
R1218 B.n604 B.n5 163.367
R1219 B.n6 B.n5 163.367
R1220 B.n7 B.n6 163.367
R1221 B.n609 B.n7 163.367
R1222 B.n609 B.n12 163.367
R1223 B.n13 B.n12 163.367
R1224 B.n14 B.n13 163.367
R1225 B.n614 B.n14 163.367
R1226 B.n614 B.n19 163.367
R1227 B.n20 B.n19 163.367
R1228 B.n21 B.n20 163.367
R1229 B.n619 B.n21 163.367
R1230 B.n619 B.n26 163.367
R1231 B.n27 B.n26 163.367
R1232 B.n28 B.n27 163.367
R1233 B.n624 B.n28 163.367
R1234 B.n624 B.n33 163.367
R1235 B.n34 B.n33 163.367
R1236 B.n91 B.n90 163.367
R1237 B.n95 B.n94 163.367
R1238 B.n99 B.n98 163.367
R1239 B.n103 B.n102 163.367
R1240 B.n107 B.n106 163.367
R1241 B.n111 B.n110 163.367
R1242 B.n115 B.n114 163.367
R1243 B.n119 B.n118 163.367
R1244 B.n123 B.n122 163.367
R1245 B.n127 B.n126 163.367
R1246 B.n131 B.n130 163.367
R1247 B.n135 B.n134 163.367
R1248 B.n139 B.n138 163.367
R1249 B.n143 B.n142 163.367
R1250 B.n147 B.n146 163.367
R1251 B.n151 B.n150 163.367
R1252 B.n155 B.n154 163.367
R1253 B.n159 B.n158 163.367
R1254 B.n163 B.n162 163.367
R1255 B.n167 B.n166 163.367
R1256 B.n171 B.n170 163.367
R1257 B.n176 B.n175 163.367
R1258 B.n180 B.n179 163.367
R1259 B.n184 B.n183 163.367
R1260 B.n188 B.n187 163.367
R1261 B.n192 B.n191 163.367
R1262 B.n197 B.n196 163.367
R1263 B.n201 B.n200 163.367
R1264 B.n205 B.n204 163.367
R1265 B.n209 B.n208 163.367
R1266 B.n213 B.n212 163.367
R1267 B.n217 B.n216 163.367
R1268 B.n221 B.n220 163.367
R1269 B.n225 B.n224 163.367
R1270 B.n229 B.n228 163.367
R1271 B.n233 B.n232 163.367
R1272 B.n237 B.n236 163.367
R1273 B.n241 B.n240 163.367
R1274 B.n245 B.n244 163.367
R1275 B.n249 B.n248 163.367
R1276 B.n253 B.n252 163.367
R1277 B.n257 B.n256 163.367
R1278 B.n261 B.n260 163.367
R1279 B.n265 B.n264 163.367
R1280 B.n269 B.n268 163.367
R1281 B.n273 B.n272 163.367
R1282 B.n275 B.n82 163.367
R1283 B.n551 B.n550 71.676
R1284 B.n545 B.n311 71.676
R1285 B.n542 B.n312 71.676
R1286 B.n538 B.n313 71.676
R1287 B.n534 B.n314 71.676
R1288 B.n530 B.n315 71.676
R1289 B.n526 B.n316 71.676
R1290 B.n522 B.n317 71.676
R1291 B.n518 B.n318 71.676
R1292 B.n514 B.n319 71.676
R1293 B.n510 B.n320 71.676
R1294 B.n506 B.n321 71.676
R1295 B.n502 B.n322 71.676
R1296 B.n498 B.n323 71.676
R1297 B.n494 B.n324 71.676
R1298 B.n490 B.n325 71.676
R1299 B.n486 B.n326 71.676
R1300 B.n482 B.n327 71.676
R1301 B.n478 B.n328 71.676
R1302 B.n474 B.n329 71.676
R1303 B.n470 B.n330 71.676
R1304 B.n466 B.n331 71.676
R1305 B.n462 B.n332 71.676
R1306 B.n458 B.n333 71.676
R1307 B.n454 B.n334 71.676
R1308 B.n450 B.n335 71.676
R1309 B.n446 B.n336 71.676
R1310 B.n442 B.n337 71.676
R1311 B.n438 B.n338 71.676
R1312 B.n434 B.n339 71.676
R1313 B.n430 B.n340 71.676
R1314 B.n426 B.n341 71.676
R1315 B.n422 B.n342 71.676
R1316 B.n418 B.n343 71.676
R1317 B.n414 B.n344 71.676
R1318 B.n410 B.n345 71.676
R1319 B.n406 B.n346 71.676
R1320 B.n402 B.n347 71.676
R1321 B.n398 B.n348 71.676
R1322 B.n394 B.n349 71.676
R1323 B.n390 B.n350 71.676
R1324 B.n386 B.n351 71.676
R1325 B.n382 B.n352 71.676
R1326 B.n378 B.n353 71.676
R1327 B.n374 B.n354 71.676
R1328 B.n370 B.n355 71.676
R1329 B.n366 B.n356 71.676
R1330 B.n87 B.n35 71.676
R1331 B.n91 B.n36 71.676
R1332 B.n95 B.n37 71.676
R1333 B.n99 B.n38 71.676
R1334 B.n103 B.n39 71.676
R1335 B.n107 B.n40 71.676
R1336 B.n111 B.n41 71.676
R1337 B.n115 B.n42 71.676
R1338 B.n119 B.n43 71.676
R1339 B.n123 B.n44 71.676
R1340 B.n127 B.n45 71.676
R1341 B.n131 B.n46 71.676
R1342 B.n135 B.n47 71.676
R1343 B.n139 B.n48 71.676
R1344 B.n143 B.n49 71.676
R1345 B.n147 B.n50 71.676
R1346 B.n151 B.n51 71.676
R1347 B.n155 B.n52 71.676
R1348 B.n159 B.n53 71.676
R1349 B.n163 B.n54 71.676
R1350 B.n167 B.n55 71.676
R1351 B.n171 B.n56 71.676
R1352 B.n176 B.n57 71.676
R1353 B.n180 B.n58 71.676
R1354 B.n184 B.n59 71.676
R1355 B.n188 B.n60 71.676
R1356 B.n192 B.n61 71.676
R1357 B.n197 B.n62 71.676
R1358 B.n201 B.n63 71.676
R1359 B.n205 B.n64 71.676
R1360 B.n209 B.n65 71.676
R1361 B.n213 B.n66 71.676
R1362 B.n217 B.n67 71.676
R1363 B.n221 B.n68 71.676
R1364 B.n225 B.n69 71.676
R1365 B.n229 B.n70 71.676
R1366 B.n233 B.n71 71.676
R1367 B.n237 B.n72 71.676
R1368 B.n241 B.n73 71.676
R1369 B.n245 B.n74 71.676
R1370 B.n249 B.n75 71.676
R1371 B.n253 B.n76 71.676
R1372 B.n257 B.n77 71.676
R1373 B.n261 B.n78 71.676
R1374 B.n265 B.n79 71.676
R1375 B.n269 B.n80 71.676
R1376 B.n273 B.n81 71.676
R1377 B.n630 B.n82 71.676
R1378 B.n630 B.n629 71.676
R1379 B.n275 B.n81 71.676
R1380 B.n272 B.n80 71.676
R1381 B.n268 B.n79 71.676
R1382 B.n264 B.n78 71.676
R1383 B.n260 B.n77 71.676
R1384 B.n256 B.n76 71.676
R1385 B.n252 B.n75 71.676
R1386 B.n248 B.n74 71.676
R1387 B.n244 B.n73 71.676
R1388 B.n240 B.n72 71.676
R1389 B.n236 B.n71 71.676
R1390 B.n232 B.n70 71.676
R1391 B.n228 B.n69 71.676
R1392 B.n224 B.n68 71.676
R1393 B.n220 B.n67 71.676
R1394 B.n216 B.n66 71.676
R1395 B.n212 B.n65 71.676
R1396 B.n208 B.n64 71.676
R1397 B.n204 B.n63 71.676
R1398 B.n200 B.n62 71.676
R1399 B.n196 B.n61 71.676
R1400 B.n191 B.n60 71.676
R1401 B.n187 B.n59 71.676
R1402 B.n183 B.n58 71.676
R1403 B.n179 B.n57 71.676
R1404 B.n175 B.n56 71.676
R1405 B.n170 B.n55 71.676
R1406 B.n166 B.n54 71.676
R1407 B.n162 B.n53 71.676
R1408 B.n158 B.n52 71.676
R1409 B.n154 B.n51 71.676
R1410 B.n150 B.n50 71.676
R1411 B.n146 B.n49 71.676
R1412 B.n142 B.n48 71.676
R1413 B.n138 B.n47 71.676
R1414 B.n134 B.n46 71.676
R1415 B.n130 B.n45 71.676
R1416 B.n126 B.n44 71.676
R1417 B.n122 B.n43 71.676
R1418 B.n118 B.n42 71.676
R1419 B.n114 B.n41 71.676
R1420 B.n110 B.n40 71.676
R1421 B.n106 B.n39 71.676
R1422 B.n102 B.n38 71.676
R1423 B.n98 B.n37 71.676
R1424 B.n94 B.n36 71.676
R1425 B.n90 B.n35 71.676
R1426 B.n551 B.n358 71.676
R1427 B.n543 B.n311 71.676
R1428 B.n539 B.n312 71.676
R1429 B.n535 B.n313 71.676
R1430 B.n531 B.n314 71.676
R1431 B.n527 B.n315 71.676
R1432 B.n523 B.n316 71.676
R1433 B.n519 B.n317 71.676
R1434 B.n515 B.n318 71.676
R1435 B.n511 B.n319 71.676
R1436 B.n507 B.n320 71.676
R1437 B.n503 B.n321 71.676
R1438 B.n499 B.n322 71.676
R1439 B.n495 B.n323 71.676
R1440 B.n491 B.n324 71.676
R1441 B.n487 B.n325 71.676
R1442 B.n483 B.n326 71.676
R1443 B.n479 B.n327 71.676
R1444 B.n475 B.n328 71.676
R1445 B.n471 B.n329 71.676
R1446 B.n467 B.n330 71.676
R1447 B.n463 B.n331 71.676
R1448 B.n459 B.n332 71.676
R1449 B.n455 B.n333 71.676
R1450 B.n451 B.n334 71.676
R1451 B.n447 B.n335 71.676
R1452 B.n443 B.n336 71.676
R1453 B.n439 B.n337 71.676
R1454 B.n435 B.n338 71.676
R1455 B.n431 B.n339 71.676
R1456 B.n427 B.n340 71.676
R1457 B.n423 B.n341 71.676
R1458 B.n419 B.n342 71.676
R1459 B.n415 B.n343 71.676
R1460 B.n411 B.n344 71.676
R1461 B.n407 B.n345 71.676
R1462 B.n403 B.n346 71.676
R1463 B.n399 B.n347 71.676
R1464 B.n395 B.n348 71.676
R1465 B.n391 B.n349 71.676
R1466 B.n387 B.n350 71.676
R1467 B.n383 B.n351 71.676
R1468 B.n379 B.n352 71.676
R1469 B.n375 B.n353 71.676
R1470 B.n371 B.n354 71.676
R1471 B.n367 B.n355 71.676
R1472 B.n356 B.n310 71.676
R1473 B.n552 B.n307 68.3082
R1474 B.n632 B.n631 68.3082
R1475 B.n364 B.n363 59.5399
R1476 B.n361 B.n360 59.5399
R1477 B.n173 B.n86 59.5399
R1478 B.n194 B.n84 59.5399
R1479 B.n558 B.n307 41.8467
R1480 B.n558 B.n302 41.8467
R1481 B.n564 B.n302 41.8467
R1482 B.n564 B.n303 41.8467
R1483 B.n570 B.n295 41.8467
R1484 B.n576 B.n295 41.8467
R1485 B.n576 B.n291 41.8467
R1486 B.n582 B.n291 41.8467
R1487 B.n588 B.n286 41.8467
R1488 B.n588 B.n287 41.8467
R1489 B.n596 B.n595 41.8467
R1490 B.n602 B.n4 41.8467
R1491 B.n665 B.n4 41.8467
R1492 B.n665 B.n664 41.8467
R1493 B.n664 B.n663 41.8467
R1494 B.n657 B.n11 41.8467
R1495 B.n656 B.n655 41.8467
R1496 B.n655 B.n15 41.8467
R1497 B.n649 B.n648 41.8467
R1498 B.n648 B.n647 41.8467
R1499 B.n647 B.n22 41.8467
R1500 B.n641 B.n22 41.8467
R1501 B.n640 B.n639 41.8467
R1502 B.n639 B.n29 41.8467
R1503 B.n633 B.n29 41.8467
R1504 B.n633 B.n632 41.8467
R1505 B.n582 B.t3 40.0005
R1506 B.n649 B.t4 40.0005
R1507 B.n596 B.t0 36.3082
R1508 B.n657 B.t1 36.3082
R1509 B.n88 B.n31 32.3127
R1510 B.n628 B.n627 32.3127
R1511 B.n555 B.n554 32.3127
R1512 B.n549 B.n305 32.3127
R1513 B.n602 B.t2 28.9236
R1514 B.n663 B.t5 28.9236
R1515 B.n303 B.t7 24.0005
R1516 B.t14 B.n640 24.0005
R1517 B B.n667 18.0485
R1518 B.n570 B.t7 17.8467
R1519 B.n641 B.t14 17.8467
R1520 B.n363 B.n362 14.352
R1521 B.n360 B.n359 14.352
R1522 B.n86 B.n85 14.352
R1523 B.n84 B.n83 14.352
R1524 B.n595 B.t2 12.9236
R1525 B.n11 B.t5 12.9236
R1526 B.n89 B.n88 10.6151
R1527 B.n92 B.n89 10.6151
R1528 B.n93 B.n92 10.6151
R1529 B.n96 B.n93 10.6151
R1530 B.n97 B.n96 10.6151
R1531 B.n100 B.n97 10.6151
R1532 B.n101 B.n100 10.6151
R1533 B.n104 B.n101 10.6151
R1534 B.n105 B.n104 10.6151
R1535 B.n108 B.n105 10.6151
R1536 B.n109 B.n108 10.6151
R1537 B.n112 B.n109 10.6151
R1538 B.n113 B.n112 10.6151
R1539 B.n116 B.n113 10.6151
R1540 B.n117 B.n116 10.6151
R1541 B.n120 B.n117 10.6151
R1542 B.n121 B.n120 10.6151
R1543 B.n124 B.n121 10.6151
R1544 B.n125 B.n124 10.6151
R1545 B.n128 B.n125 10.6151
R1546 B.n129 B.n128 10.6151
R1547 B.n132 B.n129 10.6151
R1548 B.n133 B.n132 10.6151
R1549 B.n136 B.n133 10.6151
R1550 B.n137 B.n136 10.6151
R1551 B.n140 B.n137 10.6151
R1552 B.n141 B.n140 10.6151
R1553 B.n144 B.n141 10.6151
R1554 B.n145 B.n144 10.6151
R1555 B.n148 B.n145 10.6151
R1556 B.n149 B.n148 10.6151
R1557 B.n152 B.n149 10.6151
R1558 B.n153 B.n152 10.6151
R1559 B.n156 B.n153 10.6151
R1560 B.n157 B.n156 10.6151
R1561 B.n160 B.n157 10.6151
R1562 B.n161 B.n160 10.6151
R1563 B.n164 B.n161 10.6151
R1564 B.n165 B.n164 10.6151
R1565 B.n168 B.n165 10.6151
R1566 B.n169 B.n168 10.6151
R1567 B.n172 B.n169 10.6151
R1568 B.n177 B.n174 10.6151
R1569 B.n178 B.n177 10.6151
R1570 B.n181 B.n178 10.6151
R1571 B.n182 B.n181 10.6151
R1572 B.n185 B.n182 10.6151
R1573 B.n186 B.n185 10.6151
R1574 B.n189 B.n186 10.6151
R1575 B.n190 B.n189 10.6151
R1576 B.n193 B.n190 10.6151
R1577 B.n198 B.n195 10.6151
R1578 B.n199 B.n198 10.6151
R1579 B.n202 B.n199 10.6151
R1580 B.n203 B.n202 10.6151
R1581 B.n206 B.n203 10.6151
R1582 B.n207 B.n206 10.6151
R1583 B.n210 B.n207 10.6151
R1584 B.n211 B.n210 10.6151
R1585 B.n214 B.n211 10.6151
R1586 B.n215 B.n214 10.6151
R1587 B.n218 B.n215 10.6151
R1588 B.n219 B.n218 10.6151
R1589 B.n222 B.n219 10.6151
R1590 B.n223 B.n222 10.6151
R1591 B.n226 B.n223 10.6151
R1592 B.n227 B.n226 10.6151
R1593 B.n230 B.n227 10.6151
R1594 B.n231 B.n230 10.6151
R1595 B.n234 B.n231 10.6151
R1596 B.n235 B.n234 10.6151
R1597 B.n238 B.n235 10.6151
R1598 B.n239 B.n238 10.6151
R1599 B.n242 B.n239 10.6151
R1600 B.n243 B.n242 10.6151
R1601 B.n246 B.n243 10.6151
R1602 B.n247 B.n246 10.6151
R1603 B.n250 B.n247 10.6151
R1604 B.n251 B.n250 10.6151
R1605 B.n254 B.n251 10.6151
R1606 B.n255 B.n254 10.6151
R1607 B.n258 B.n255 10.6151
R1608 B.n259 B.n258 10.6151
R1609 B.n262 B.n259 10.6151
R1610 B.n263 B.n262 10.6151
R1611 B.n266 B.n263 10.6151
R1612 B.n267 B.n266 10.6151
R1613 B.n270 B.n267 10.6151
R1614 B.n271 B.n270 10.6151
R1615 B.n274 B.n271 10.6151
R1616 B.n276 B.n274 10.6151
R1617 B.n277 B.n276 10.6151
R1618 B.n628 B.n277 10.6151
R1619 B.n556 B.n555 10.6151
R1620 B.n556 B.n300 10.6151
R1621 B.n566 B.n300 10.6151
R1622 B.n567 B.n566 10.6151
R1623 B.n568 B.n567 10.6151
R1624 B.n568 B.n293 10.6151
R1625 B.n578 B.n293 10.6151
R1626 B.n579 B.n578 10.6151
R1627 B.n580 B.n579 10.6151
R1628 B.n580 B.n284 10.6151
R1629 B.n590 B.n284 10.6151
R1630 B.n591 B.n590 10.6151
R1631 B.n593 B.n591 10.6151
R1632 B.n593 B.n592 10.6151
R1633 B.n592 B.n278 10.6151
R1634 B.n605 B.n278 10.6151
R1635 B.n606 B.n605 10.6151
R1636 B.n607 B.n606 10.6151
R1637 B.n608 B.n607 10.6151
R1638 B.n610 B.n608 10.6151
R1639 B.n611 B.n610 10.6151
R1640 B.n612 B.n611 10.6151
R1641 B.n613 B.n612 10.6151
R1642 B.n615 B.n613 10.6151
R1643 B.n616 B.n615 10.6151
R1644 B.n617 B.n616 10.6151
R1645 B.n618 B.n617 10.6151
R1646 B.n620 B.n618 10.6151
R1647 B.n621 B.n620 10.6151
R1648 B.n622 B.n621 10.6151
R1649 B.n623 B.n622 10.6151
R1650 B.n625 B.n623 10.6151
R1651 B.n626 B.n625 10.6151
R1652 B.n627 B.n626 10.6151
R1653 B.n549 B.n548 10.6151
R1654 B.n548 B.n547 10.6151
R1655 B.n547 B.n546 10.6151
R1656 B.n546 B.n544 10.6151
R1657 B.n544 B.n541 10.6151
R1658 B.n541 B.n540 10.6151
R1659 B.n540 B.n537 10.6151
R1660 B.n537 B.n536 10.6151
R1661 B.n536 B.n533 10.6151
R1662 B.n533 B.n532 10.6151
R1663 B.n532 B.n529 10.6151
R1664 B.n529 B.n528 10.6151
R1665 B.n528 B.n525 10.6151
R1666 B.n525 B.n524 10.6151
R1667 B.n524 B.n521 10.6151
R1668 B.n521 B.n520 10.6151
R1669 B.n520 B.n517 10.6151
R1670 B.n517 B.n516 10.6151
R1671 B.n516 B.n513 10.6151
R1672 B.n513 B.n512 10.6151
R1673 B.n512 B.n509 10.6151
R1674 B.n509 B.n508 10.6151
R1675 B.n508 B.n505 10.6151
R1676 B.n505 B.n504 10.6151
R1677 B.n504 B.n501 10.6151
R1678 B.n501 B.n500 10.6151
R1679 B.n500 B.n497 10.6151
R1680 B.n497 B.n496 10.6151
R1681 B.n496 B.n493 10.6151
R1682 B.n493 B.n492 10.6151
R1683 B.n492 B.n489 10.6151
R1684 B.n489 B.n488 10.6151
R1685 B.n488 B.n485 10.6151
R1686 B.n485 B.n484 10.6151
R1687 B.n484 B.n481 10.6151
R1688 B.n481 B.n480 10.6151
R1689 B.n480 B.n477 10.6151
R1690 B.n477 B.n476 10.6151
R1691 B.n476 B.n473 10.6151
R1692 B.n473 B.n472 10.6151
R1693 B.n472 B.n469 10.6151
R1694 B.n469 B.n468 10.6151
R1695 B.n465 B.n464 10.6151
R1696 B.n464 B.n461 10.6151
R1697 B.n461 B.n460 10.6151
R1698 B.n460 B.n457 10.6151
R1699 B.n457 B.n456 10.6151
R1700 B.n456 B.n453 10.6151
R1701 B.n453 B.n452 10.6151
R1702 B.n452 B.n449 10.6151
R1703 B.n449 B.n448 10.6151
R1704 B.n445 B.n444 10.6151
R1705 B.n444 B.n441 10.6151
R1706 B.n441 B.n440 10.6151
R1707 B.n440 B.n437 10.6151
R1708 B.n437 B.n436 10.6151
R1709 B.n436 B.n433 10.6151
R1710 B.n433 B.n432 10.6151
R1711 B.n432 B.n429 10.6151
R1712 B.n429 B.n428 10.6151
R1713 B.n428 B.n425 10.6151
R1714 B.n425 B.n424 10.6151
R1715 B.n424 B.n421 10.6151
R1716 B.n421 B.n420 10.6151
R1717 B.n420 B.n417 10.6151
R1718 B.n417 B.n416 10.6151
R1719 B.n416 B.n413 10.6151
R1720 B.n413 B.n412 10.6151
R1721 B.n412 B.n409 10.6151
R1722 B.n409 B.n408 10.6151
R1723 B.n408 B.n405 10.6151
R1724 B.n405 B.n404 10.6151
R1725 B.n404 B.n401 10.6151
R1726 B.n401 B.n400 10.6151
R1727 B.n400 B.n397 10.6151
R1728 B.n397 B.n396 10.6151
R1729 B.n396 B.n393 10.6151
R1730 B.n393 B.n392 10.6151
R1731 B.n392 B.n389 10.6151
R1732 B.n389 B.n388 10.6151
R1733 B.n388 B.n385 10.6151
R1734 B.n385 B.n384 10.6151
R1735 B.n384 B.n381 10.6151
R1736 B.n381 B.n380 10.6151
R1737 B.n380 B.n377 10.6151
R1738 B.n377 B.n376 10.6151
R1739 B.n376 B.n373 10.6151
R1740 B.n373 B.n372 10.6151
R1741 B.n372 B.n369 10.6151
R1742 B.n369 B.n368 10.6151
R1743 B.n368 B.n365 10.6151
R1744 B.n365 B.n309 10.6151
R1745 B.n554 B.n309 10.6151
R1746 B.n560 B.n305 10.6151
R1747 B.n561 B.n560 10.6151
R1748 B.n562 B.n561 10.6151
R1749 B.n562 B.n297 10.6151
R1750 B.n572 B.n297 10.6151
R1751 B.n573 B.n572 10.6151
R1752 B.n574 B.n573 10.6151
R1753 B.n574 B.n289 10.6151
R1754 B.n584 B.n289 10.6151
R1755 B.n585 B.n584 10.6151
R1756 B.n586 B.n585 10.6151
R1757 B.n586 B.n281 10.6151
R1758 B.n598 B.n281 10.6151
R1759 B.n599 B.n598 10.6151
R1760 B.n600 B.n599 10.6151
R1761 B.n600 B.n0 10.6151
R1762 B.n661 B.n1 10.6151
R1763 B.n661 B.n660 10.6151
R1764 B.n660 B.n659 10.6151
R1765 B.n659 B.n9 10.6151
R1766 B.n653 B.n9 10.6151
R1767 B.n653 B.n652 10.6151
R1768 B.n652 B.n651 10.6151
R1769 B.n651 B.n17 10.6151
R1770 B.n645 B.n17 10.6151
R1771 B.n645 B.n644 10.6151
R1772 B.n644 B.n643 10.6151
R1773 B.n643 B.n24 10.6151
R1774 B.n637 B.n24 10.6151
R1775 B.n637 B.n636 10.6151
R1776 B.n636 B.n635 10.6151
R1777 B.n635 B.n31 10.6151
R1778 B.n173 B.n172 9.36635
R1779 B.n195 B.n194 9.36635
R1780 B.n468 B.n361 9.36635
R1781 B.n445 B.n364 9.36635
R1782 B.n287 B.t0 5.53896
R1783 B.t1 B.n656 5.53896
R1784 B.n667 B.n0 2.81026
R1785 B.n667 B.n1 2.81026
R1786 B.t3 B.n286 1.84665
R1787 B.t4 B.n15 1.84665
R1788 B.n174 B.n173 1.24928
R1789 B.n194 B.n193 1.24928
R1790 B.n465 B.n361 1.24928
R1791 B.n448 B.n364 1.24928
R1792 VP.n1 VP.t0 860.577
R1793 VP.n8 VP.t3 841.558
R1794 VP.n6 VP.t4 841.558
R1795 VP.n3 VP.t2 841.558
R1796 VP.n7 VP.t5 836.447
R1797 VP.n2 VP.t1 836.447
R1798 VP.n9 VP.n8 161.3
R1799 VP.n4 VP.n3 161.3
R1800 VP.n7 VP.n0 161.3
R1801 VP.n6 VP.n5 161.3
R1802 VP.n4 VP.n1 71.3843
R1803 VP.n7 VP.n6 43.0884
R1804 VP.n8 VP.n7 43.0884
R1805 VP.n3 VP.n2 43.0884
R1806 VP.n5 VP.n4 40.6066
R1807 VP.n2 VP.n1 18.9966
R1808 VP.n5 VP.n0 0.189894
R1809 VP.n9 VP.n0 0.189894
R1810 VP VP.n9 0.0516364
R1811 VDD1.n68 VDD1.n67 289.615
R1812 VDD1.n137 VDD1.n136 289.615
R1813 VDD1.n67 VDD1.n66 185
R1814 VDD1.n2 VDD1.n1 185
R1815 VDD1.n61 VDD1.n60 185
R1816 VDD1.n59 VDD1.n58 185
R1817 VDD1.n6 VDD1.n5 185
R1818 VDD1.n53 VDD1.n52 185
R1819 VDD1.n51 VDD1.n50 185
R1820 VDD1.n10 VDD1.n9 185
R1821 VDD1.n45 VDD1.n44 185
R1822 VDD1.n43 VDD1.n42 185
R1823 VDD1.n14 VDD1.n13 185
R1824 VDD1.n37 VDD1.n36 185
R1825 VDD1.n35 VDD1.n34 185
R1826 VDD1.n18 VDD1.n17 185
R1827 VDD1.n29 VDD1.n28 185
R1828 VDD1.n27 VDD1.n26 185
R1829 VDD1.n22 VDD1.n21 185
R1830 VDD1.n91 VDD1.n90 185
R1831 VDD1.n96 VDD1.n95 185
R1832 VDD1.n98 VDD1.n97 185
R1833 VDD1.n87 VDD1.n86 185
R1834 VDD1.n104 VDD1.n103 185
R1835 VDD1.n106 VDD1.n105 185
R1836 VDD1.n83 VDD1.n82 185
R1837 VDD1.n112 VDD1.n111 185
R1838 VDD1.n114 VDD1.n113 185
R1839 VDD1.n79 VDD1.n78 185
R1840 VDD1.n120 VDD1.n119 185
R1841 VDD1.n122 VDD1.n121 185
R1842 VDD1.n75 VDD1.n74 185
R1843 VDD1.n128 VDD1.n127 185
R1844 VDD1.n130 VDD1.n129 185
R1845 VDD1.n71 VDD1.n70 185
R1846 VDD1.n136 VDD1.n135 185
R1847 VDD1.n92 VDD1.t1 147.659
R1848 VDD1.n23 VDD1.t5 147.659
R1849 VDD1.n67 VDD1.n1 104.615
R1850 VDD1.n60 VDD1.n1 104.615
R1851 VDD1.n60 VDD1.n59 104.615
R1852 VDD1.n59 VDD1.n5 104.615
R1853 VDD1.n52 VDD1.n5 104.615
R1854 VDD1.n52 VDD1.n51 104.615
R1855 VDD1.n51 VDD1.n9 104.615
R1856 VDD1.n44 VDD1.n9 104.615
R1857 VDD1.n44 VDD1.n43 104.615
R1858 VDD1.n43 VDD1.n13 104.615
R1859 VDD1.n36 VDD1.n13 104.615
R1860 VDD1.n36 VDD1.n35 104.615
R1861 VDD1.n35 VDD1.n17 104.615
R1862 VDD1.n28 VDD1.n17 104.615
R1863 VDD1.n28 VDD1.n27 104.615
R1864 VDD1.n27 VDD1.n21 104.615
R1865 VDD1.n96 VDD1.n90 104.615
R1866 VDD1.n97 VDD1.n96 104.615
R1867 VDD1.n97 VDD1.n86 104.615
R1868 VDD1.n104 VDD1.n86 104.615
R1869 VDD1.n105 VDD1.n104 104.615
R1870 VDD1.n105 VDD1.n82 104.615
R1871 VDD1.n112 VDD1.n82 104.615
R1872 VDD1.n113 VDD1.n112 104.615
R1873 VDD1.n113 VDD1.n78 104.615
R1874 VDD1.n120 VDD1.n78 104.615
R1875 VDD1.n121 VDD1.n120 104.615
R1876 VDD1.n121 VDD1.n74 104.615
R1877 VDD1.n128 VDD1.n74 104.615
R1878 VDD1.n129 VDD1.n128 104.615
R1879 VDD1.n129 VDD1.n70 104.615
R1880 VDD1.n136 VDD1.n70 104.615
R1881 VDD1.n139 VDD1.n138 63.6388
R1882 VDD1.n141 VDD1.n140 63.5347
R1883 VDD1.t5 VDD1.n21 52.3082
R1884 VDD1.t1 VDD1.n90 52.3082
R1885 VDD1 VDD1.n68 51.3402
R1886 VDD1.n139 VDD1.n137 51.2266
R1887 VDD1.n141 VDD1.n139 37.5526
R1888 VDD1.n23 VDD1.n22 15.6677
R1889 VDD1.n92 VDD1.n91 15.6677
R1890 VDD1.n66 VDD1.n0 12.8005
R1891 VDD1.n26 VDD1.n25 12.8005
R1892 VDD1.n95 VDD1.n94 12.8005
R1893 VDD1.n135 VDD1.n69 12.8005
R1894 VDD1.n65 VDD1.n2 12.0247
R1895 VDD1.n29 VDD1.n20 12.0247
R1896 VDD1.n98 VDD1.n89 12.0247
R1897 VDD1.n134 VDD1.n71 12.0247
R1898 VDD1.n62 VDD1.n61 11.249
R1899 VDD1.n30 VDD1.n18 11.249
R1900 VDD1.n99 VDD1.n87 11.249
R1901 VDD1.n131 VDD1.n130 11.249
R1902 VDD1.n58 VDD1.n4 10.4732
R1903 VDD1.n34 VDD1.n33 10.4732
R1904 VDD1.n103 VDD1.n102 10.4732
R1905 VDD1.n127 VDD1.n73 10.4732
R1906 VDD1.n57 VDD1.n6 9.69747
R1907 VDD1.n37 VDD1.n16 9.69747
R1908 VDD1.n106 VDD1.n85 9.69747
R1909 VDD1.n126 VDD1.n75 9.69747
R1910 VDD1.n64 VDD1.n0 9.45567
R1911 VDD1.n133 VDD1.n69 9.45567
R1912 VDD1.n49 VDD1.n48 9.3005
R1913 VDD1.n8 VDD1.n7 9.3005
R1914 VDD1.n55 VDD1.n54 9.3005
R1915 VDD1.n57 VDD1.n56 9.3005
R1916 VDD1.n4 VDD1.n3 9.3005
R1917 VDD1.n63 VDD1.n62 9.3005
R1918 VDD1.n65 VDD1.n64 9.3005
R1919 VDD1.n47 VDD1.n46 9.3005
R1920 VDD1.n12 VDD1.n11 9.3005
R1921 VDD1.n41 VDD1.n40 9.3005
R1922 VDD1.n39 VDD1.n38 9.3005
R1923 VDD1.n16 VDD1.n15 9.3005
R1924 VDD1.n33 VDD1.n32 9.3005
R1925 VDD1.n31 VDD1.n30 9.3005
R1926 VDD1.n20 VDD1.n19 9.3005
R1927 VDD1.n25 VDD1.n24 9.3005
R1928 VDD1.n116 VDD1.n115 9.3005
R1929 VDD1.n118 VDD1.n117 9.3005
R1930 VDD1.n77 VDD1.n76 9.3005
R1931 VDD1.n124 VDD1.n123 9.3005
R1932 VDD1.n126 VDD1.n125 9.3005
R1933 VDD1.n73 VDD1.n72 9.3005
R1934 VDD1.n132 VDD1.n131 9.3005
R1935 VDD1.n134 VDD1.n133 9.3005
R1936 VDD1.n110 VDD1.n109 9.3005
R1937 VDD1.n108 VDD1.n107 9.3005
R1938 VDD1.n85 VDD1.n84 9.3005
R1939 VDD1.n102 VDD1.n101 9.3005
R1940 VDD1.n100 VDD1.n99 9.3005
R1941 VDD1.n89 VDD1.n88 9.3005
R1942 VDD1.n94 VDD1.n93 9.3005
R1943 VDD1.n81 VDD1.n80 9.3005
R1944 VDD1.n54 VDD1.n53 8.92171
R1945 VDD1.n38 VDD1.n14 8.92171
R1946 VDD1.n107 VDD1.n83 8.92171
R1947 VDD1.n123 VDD1.n122 8.92171
R1948 VDD1.n50 VDD1.n8 8.14595
R1949 VDD1.n42 VDD1.n41 8.14595
R1950 VDD1.n111 VDD1.n110 8.14595
R1951 VDD1.n119 VDD1.n77 8.14595
R1952 VDD1.n49 VDD1.n10 7.3702
R1953 VDD1.n45 VDD1.n12 7.3702
R1954 VDD1.n114 VDD1.n81 7.3702
R1955 VDD1.n118 VDD1.n79 7.3702
R1956 VDD1.n46 VDD1.n10 6.59444
R1957 VDD1.n46 VDD1.n45 6.59444
R1958 VDD1.n115 VDD1.n114 6.59444
R1959 VDD1.n115 VDD1.n79 6.59444
R1960 VDD1.n50 VDD1.n49 5.81868
R1961 VDD1.n42 VDD1.n12 5.81868
R1962 VDD1.n111 VDD1.n81 5.81868
R1963 VDD1.n119 VDD1.n118 5.81868
R1964 VDD1.n53 VDD1.n8 5.04292
R1965 VDD1.n41 VDD1.n14 5.04292
R1966 VDD1.n110 VDD1.n83 5.04292
R1967 VDD1.n122 VDD1.n77 5.04292
R1968 VDD1.n93 VDD1.n92 4.38563
R1969 VDD1.n24 VDD1.n23 4.38563
R1970 VDD1.n54 VDD1.n6 4.26717
R1971 VDD1.n38 VDD1.n37 4.26717
R1972 VDD1.n107 VDD1.n106 4.26717
R1973 VDD1.n123 VDD1.n75 4.26717
R1974 VDD1.n58 VDD1.n57 3.49141
R1975 VDD1.n34 VDD1.n16 3.49141
R1976 VDD1.n103 VDD1.n85 3.49141
R1977 VDD1.n127 VDD1.n126 3.49141
R1978 VDD1.n61 VDD1.n4 2.71565
R1979 VDD1.n33 VDD1.n18 2.71565
R1980 VDD1.n102 VDD1.n87 2.71565
R1981 VDD1.n130 VDD1.n73 2.71565
R1982 VDD1.n62 VDD1.n2 1.93989
R1983 VDD1.n30 VDD1.n29 1.93989
R1984 VDD1.n99 VDD1.n98 1.93989
R1985 VDD1.n131 VDD1.n71 1.93989
R1986 VDD1.n140 VDD1.t4 1.57193
R1987 VDD1.n140 VDD1.t3 1.57193
R1988 VDD1.n138 VDD1.t0 1.57193
R1989 VDD1.n138 VDD1.t2 1.57193
R1990 VDD1.n66 VDD1.n65 1.16414
R1991 VDD1.n26 VDD1.n20 1.16414
R1992 VDD1.n95 VDD1.n89 1.16414
R1993 VDD1.n135 VDD1.n134 1.16414
R1994 VDD1.n68 VDD1.n0 0.388379
R1995 VDD1.n25 VDD1.n22 0.388379
R1996 VDD1.n94 VDD1.n91 0.388379
R1997 VDD1.n137 VDD1.n69 0.388379
R1998 VDD1.n64 VDD1.n63 0.155672
R1999 VDD1.n63 VDD1.n3 0.155672
R2000 VDD1.n56 VDD1.n3 0.155672
R2001 VDD1.n56 VDD1.n55 0.155672
R2002 VDD1.n55 VDD1.n7 0.155672
R2003 VDD1.n48 VDD1.n7 0.155672
R2004 VDD1.n48 VDD1.n47 0.155672
R2005 VDD1.n47 VDD1.n11 0.155672
R2006 VDD1.n40 VDD1.n11 0.155672
R2007 VDD1.n40 VDD1.n39 0.155672
R2008 VDD1.n39 VDD1.n15 0.155672
R2009 VDD1.n32 VDD1.n15 0.155672
R2010 VDD1.n32 VDD1.n31 0.155672
R2011 VDD1.n31 VDD1.n19 0.155672
R2012 VDD1.n24 VDD1.n19 0.155672
R2013 VDD1.n93 VDD1.n88 0.155672
R2014 VDD1.n100 VDD1.n88 0.155672
R2015 VDD1.n101 VDD1.n100 0.155672
R2016 VDD1.n101 VDD1.n84 0.155672
R2017 VDD1.n108 VDD1.n84 0.155672
R2018 VDD1.n109 VDD1.n108 0.155672
R2019 VDD1.n109 VDD1.n80 0.155672
R2020 VDD1.n116 VDD1.n80 0.155672
R2021 VDD1.n117 VDD1.n116 0.155672
R2022 VDD1.n117 VDD1.n76 0.155672
R2023 VDD1.n124 VDD1.n76 0.155672
R2024 VDD1.n125 VDD1.n124 0.155672
R2025 VDD1.n125 VDD1.n72 0.155672
R2026 VDD1.n132 VDD1.n72 0.155672
R2027 VDD1.n133 VDD1.n132 0.155672
R2028 VDD1 VDD1.n141 0.101793
C0 VP VTAIL 2.9762f
C1 VTAIL VDD2 12.838201f
C2 VP VDD1 3.51872f
C3 VDD1 VDD2 0.608284f
C4 VTAIL VN 2.96146f
C5 VDD1 VN 0.148061f
C6 VP VDD2 0.273618f
C7 VTAIL VDD1 12.807799f
C8 VP VN 4.90654f
C9 VDD2 VN 3.39836f
C10 VDD2 B 4.378258f
C11 VDD1 B 4.357642f
C12 VTAIL B 6.310402f
C13 VN B 7.15885f
C14 VP B 4.927495f
C15 VDD1.n0 B 0.014504f
C16 VDD1.n1 B 0.032781f
C17 VDD1.n2 B 0.014685f
C18 VDD1.n3 B 0.02581f
C19 VDD1.n4 B 0.013869f
C20 VDD1.n5 B 0.032781f
C21 VDD1.n6 B 0.014685f
C22 VDD1.n7 B 0.02581f
C23 VDD1.n8 B 0.013869f
C24 VDD1.n9 B 0.032781f
C25 VDD1.n10 B 0.014685f
C26 VDD1.n11 B 0.02581f
C27 VDD1.n12 B 0.013869f
C28 VDD1.n13 B 0.032781f
C29 VDD1.n14 B 0.014685f
C30 VDD1.n15 B 0.02581f
C31 VDD1.n16 B 0.013869f
C32 VDD1.n17 B 0.032781f
C33 VDD1.n18 B 0.014685f
C34 VDD1.n19 B 0.02581f
C35 VDD1.n20 B 0.013869f
C36 VDD1.n21 B 0.024586f
C37 VDD1.n22 B 0.019365f
C38 VDD1.t5 B 0.05384f
C39 VDD1.n23 B 0.152805f
C40 VDD1.n24 B 1.39532f
C41 VDD1.n25 B 0.013869f
C42 VDD1.n26 B 0.014685f
C43 VDD1.n27 B 0.032781f
C44 VDD1.n28 B 0.032781f
C45 VDD1.n29 B 0.014685f
C46 VDD1.n30 B 0.013869f
C47 VDD1.n31 B 0.02581f
C48 VDD1.n32 B 0.02581f
C49 VDD1.n33 B 0.013869f
C50 VDD1.n34 B 0.014685f
C51 VDD1.n35 B 0.032781f
C52 VDD1.n36 B 0.032781f
C53 VDD1.n37 B 0.014685f
C54 VDD1.n38 B 0.013869f
C55 VDD1.n39 B 0.02581f
C56 VDD1.n40 B 0.02581f
C57 VDD1.n41 B 0.013869f
C58 VDD1.n42 B 0.014685f
C59 VDD1.n43 B 0.032781f
C60 VDD1.n44 B 0.032781f
C61 VDD1.n45 B 0.014685f
C62 VDD1.n46 B 0.013869f
C63 VDD1.n47 B 0.02581f
C64 VDD1.n48 B 0.02581f
C65 VDD1.n49 B 0.013869f
C66 VDD1.n50 B 0.014685f
C67 VDD1.n51 B 0.032781f
C68 VDD1.n52 B 0.032781f
C69 VDD1.n53 B 0.014685f
C70 VDD1.n54 B 0.013869f
C71 VDD1.n55 B 0.02581f
C72 VDD1.n56 B 0.02581f
C73 VDD1.n57 B 0.013869f
C74 VDD1.n58 B 0.014685f
C75 VDD1.n59 B 0.032781f
C76 VDD1.n60 B 0.032781f
C77 VDD1.n61 B 0.014685f
C78 VDD1.n62 B 0.013869f
C79 VDD1.n63 B 0.02581f
C80 VDD1.n64 B 0.063888f
C81 VDD1.n65 B 0.013869f
C82 VDD1.n66 B 0.014685f
C83 VDD1.n67 B 0.064807f
C84 VDD1.n68 B 0.072431f
C85 VDD1.n69 B 0.014504f
C86 VDD1.n70 B 0.032781f
C87 VDD1.n71 B 0.014685f
C88 VDD1.n72 B 0.02581f
C89 VDD1.n73 B 0.013869f
C90 VDD1.n74 B 0.032781f
C91 VDD1.n75 B 0.014685f
C92 VDD1.n76 B 0.02581f
C93 VDD1.n77 B 0.013869f
C94 VDD1.n78 B 0.032781f
C95 VDD1.n79 B 0.014685f
C96 VDD1.n80 B 0.02581f
C97 VDD1.n81 B 0.013869f
C98 VDD1.n82 B 0.032781f
C99 VDD1.n83 B 0.014685f
C100 VDD1.n84 B 0.02581f
C101 VDD1.n85 B 0.013869f
C102 VDD1.n86 B 0.032781f
C103 VDD1.n87 B 0.014685f
C104 VDD1.n88 B 0.02581f
C105 VDD1.n89 B 0.013869f
C106 VDD1.n90 B 0.024586f
C107 VDD1.n91 B 0.019365f
C108 VDD1.t1 B 0.05384f
C109 VDD1.n92 B 0.152805f
C110 VDD1.n93 B 1.39532f
C111 VDD1.n94 B 0.013869f
C112 VDD1.n95 B 0.014685f
C113 VDD1.n96 B 0.032781f
C114 VDD1.n97 B 0.032781f
C115 VDD1.n98 B 0.014685f
C116 VDD1.n99 B 0.013869f
C117 VDD1.n100 B 0.02581f
C118 VDD1.n101 B 0.02581f
C119 VDD1.n102 B 0.013869f
C120 VDD1.n103 B 0.014685f
C121 VDD1.n104 B 0.032781f
C122 VDD1.n105 B 0.032781f
C123 VDD1.n106 B 0.014685f
C124 VDD1.n107 B 0.013869f
C125 VDD1.n108 B 0.02581f
C126 VDD1.n109 B 0.02581f
C127 VDD1.n110 B 0.013869f
C128 VDD1.n111 B 0.014685f
C129 VDD1.n112 B 0.032781f
C130 VDD1.n113 B 0.032781f
C131 VDD1.n114 B 0.014685f
C132 VDD1.n115 B 0.013869f
C133 VDD1.n116 B 0.02581f
C134 VDD1.n117 B 0.02581f
C135 VDD1.n118 B 0.013869f
C136 VDD1.n119 B 0.014685f
C137 VDD1.n120 B 0.032781f
C138 VDD1.n121 B 0.032781f
C139 VDD1.n122 B 0.014685f
C140 VDD1.n123 B 0.013869f
C141 VDD1.n124 B 0.02581f
C142 VDD1.n125 B 0.02581f
C143 VDD1.n126 B 0.013869f
C144 VDD1.n127 B 0.014685f
C145 VDD1.n128 B 0.032781f
C146 VDD1.n129 B 0.032781f
C147 VDD1.n130 B 0.014685f
C148 VDD1.n131 B 0.013869f
C149 VDD1.n132 B 0.02581f
C150 VDD1.n133 B 0.063888f
C151 VDD1.n134 B 0.013869f
C152 VDD1.n135 B 0.014685f
C153 VDD1.n136 B 0.064807f
C154 VDD1.n137 B 0.072153f
C155 VDD1.t0 B 0.256983f
C156 VDD1.t2 B 0.256983f
C157 VDD1.n138 B 2.30588f
C158 VDD1.n139 B 1.88689f
C159 VDD1.t4 B 0.256983f
C160 VDD1.t3 B 0.256983f
C161 VDD1.n140 B 2.30541f
C162 VDD1.n141 B 2.28286f
C163 VP.n0 B 0.054899f
C164 VP.t4 B 0.809961f
C165 VP.t0 B 0.817141f
C166 VP.n1 B 0.318045f
C167 VP.t1 B 0.808052f
C168 VP.n2 B 0.334344f
C169 VP.t2 B 0.809961f
C170 VP.n3 B 0.324819f
C171 VP.n4 B 2.26327f
C172 VP.n5 B 2.18942f
C173 VP.n6 B 0.324819f
C174 VP.t5 B 0.808052f
C175 VP.n7 B 0.334344f
C176 VP.t3 B 0.809961f
C177 VP.n8 B 0.324819f
C178 VP.n9 B 0.042545f
C179 VDD2.n0 B 0.0145f
C180 VDD2.n1 B 0.032772f
C181 VDD2.n2 B 0.014681f
C182 VDD2.n3 B 0.025802f
C183 VDD2.n4 B 0.013865f
C184 VDD2.n5 B 0.032772f
C185 VDD2.n6 B 0.014681f
C186 VDD2.n7 B 0.025802f
C187 VDD2.n8 B 0.013865f
C188 VDD2.n9 B 0.032772f
C189 VDD2.n10 B 0.014681f
C190 VDD2.n11 B 0.025802f
C191 VDD2.n12 B 0.013865f
C192 VDD2.n13 B 0.032772f
C193 VDD2.n14 B 0.014681f
C194 VDD2.n15 B 0.025802f
C195 VDD2.n16 B 0.013865f
C196 VDD2.n17 B 0.032772f
C197 VDD2.n18 B 0.014681f
C198 VDD2.n19 B 0.025802f
C199 VDD2.n20 B 0.013865f
C200 VDD2.n21 B 0.024579f
C201 VDD2.n22 B 0.019359f
C202 VDD2.t1 B 0.053824f
C203 VDD2.n23 B 0.152761f
C204 VDD2.n24 B 1.39492f
C205 VDD2.n25 B 0.013865f
C206 VDD2.n26 B 0.014681f
C207 VDD2.n27 B 0.032772f
C208 VDD2.n28 B 0.032772f
C209 VDD2.n29 B 0.014681f
C210 VDD2.n30 B 0.013865f
C211 VDD2.n31 B 0.025802f
C212 VDD2.n32 B 0.025802f
C213 VDD2.n33 B 0.013865f
C214 VDD2.n34 B 0.014681f
C215 VDD2.n35 B 0.032772f
C216 VDD2.n36 B 0.032772f
C217 VDD2.n37 B 0.014681f
C218 VDD2.n38 B 0.013865f
C219 VDD2.n39 B 0.025802f
C220 VDD2.n40 B 0.025802f
C221 VDD2.n41 B 0.013865f
C222 VDD2.n42 B 0.014681f
C223 VDD2.n43 B 0.032772f
C224 VDD2.n44 B 0.032772f
C225 VDD2.n45 B 0.014681f
C226 VDD2.n46 B 0.013865f
C227 VDD2.n47 B 0.025802f
C228 VDD2.n48 B 0.025802f
C229 VDD2.n49 B 0.013865f
C230 VDD2.n50 B 0.014681f
C231 VDD2.n51 B 0.032772f
C232 VDD2.n52 B 0.032772f
C233 VDD2.n53 B 0.014681f
C234 VDD2.n54 B 0.013865f
C235 VDD2.n55 B 0.025802f
C236 VDD2.n56 B 0.025802f
C237 VDD2.n57 B 0.013865f
C238 VDD2.n58 B 0.014681f
C239 VDD2.n59 B 0.032772f
C240 VDD2.n60 B 0.032772f
C241 VDD2.n61 B 0.014681f
C242 VDD2.n62 B 0.013865f
C243 VDD2.n63 B 0.025802f
C244 VDD2.n64 B 0.06387f
C245 VDD2.n65 B 0.013865f
C246 VDD2.n66 B 0.014681f
C247 VDD2.n67 B 0.064788f
C248 VDD2.n68 B 0.072132f
C249 VDD2.t4 B 0.256909f
C250 VDD2.t0 B 0.256909f
C251 VDD2.n69 B 2.30522f
C252 VDD2.n70 B 1.81348f
C253 VDD2.n71 B 0.0145f
C254 VDD2.n72 B 0.032772f
C255 VDD2.n73 B 0.014681f
C256 VDD2.n74 B 0.025802f
C257 VDD2.n75 B 0.013865f
C258 VDD2.n76 B 0.032772f
C259 VDD2.n77 B 0.014681f
C260 VDD2.n78 B 0.025802f
C261 VDD2.n79 B 0.013865f
C262 VDD2.n80 B 0.032772f
C263 VDD2.n81 B 0.014681f
C264 VDD2.n82 B 0.025802f
C265 VDD2.n83 B 0.013865f
C266 VDD2.n84 B 0.032772f
C267 VDD2.n85 B 0.014681f
C268 VDD2.n86 B 0.025802f
C269 VDD2.n87 B 0.013865f
C270 VDD2.n88 B 0.032772f
C271 VDD2.n89 B 0.014681f
C272 VDD2.n90 B 0.025802f
C273 VDD2.n91 B 0.013865f
C274 VDD2.n92 B 0.024579f
C275 VDD2.n93 B 0.019359f
C276 VDD2.t5 B 0.053824f
C277 VDD2.n94 B 0.152761f
C278 VDD2.n95 B 1.39492f
C279 VDD2.n96 B 0.013865f
C280 VDD2.n97 B 0.014681f
C281 VDD2.n98 B 0.032772f
C282 VDD2.n99 B 0.032772f
C283 VDD2.n100 B 0.014681f
C284 VDD2.n101 B 0.013865f
C285 VDD2.n102 B 0.025802f
C286 VDD2.n103 B 0.025802f
C287 VDD2.n104 B 0.013865f
C288 VDD2.n105 B 0.014681f
C289 VDD2.n106 B 0.032772f
C290 VDD2.n107 B 0.032772f
C291 VDD2.n108 B 0.014681f
C292 VDD2.n109 B 0.013865f
C293 VDD2.n110 B 0.025802f
C294 VDD2.n111 B 0.025802f
C295 VDD2.n112 B 0.013865f
C296 VDD2.n113 B 0.014681f
C297 VDD2.n114 B 0.032772f
C298 VDD2.n115 B 0.032772f
C299 VDD2.n116 B 0.014681f
C300 VDD2.n117 B 0.013865f
C301 VDD2.n118 B 0.025802f
C302 VDD2.n119 B 0.025802f
C303 VDD2.n120 B 0.013865f
C304 VDD2.n121 B 0.014681f
C305 VDD2.n122 B 0.032772f
C306 VDD2.n123 B 0.032772f
C307 VDD2.n124 B 0.014681f
C308 VDD2.n125 B 0.013865f
C309 VDD2.n126 B 0.025802f
C310 VDD2.n127 B 0.025802f
C311 VDD2.n128 B 0.013865f
C312 VDD2.n129 B 0.014681f
C313 VDD2.n130 B 0.032772f
C314 VDD2.n131 B 0.032772f
C315 VDD2.n132 B 0.014681f
C316 VDD2.n133 B 0.013865f
C317 VDD2.n134 B 0.025802f
C318 VDD2.n135 B 0.06387f
C319 VDD2.n136 B 0.013865f
C320 VDD2.n137 B 0.014681f
C321 VDD2.n138 B 0.064788f
C322 VDD2.n139 B 0.071403f
C323 VDD2.n140 B 2.07879f
C324 VDD2.t2 B 0.256909f
C325 VDD2.t3 B 0.256909f
C326 VDD2.n141 B 2.30519f
C327 VTAIL.t11 B 0.264631f
C328 VTAIL.t10 B 0.264631f
C329 VTAIL.n0 B 2.3005f
C330 VTAIL.n1 B 0.335197f
C331 VTAIL.n2 B 0.014936f
C332 VTAIL.n3 B 0.033757f
C333 VTAIL.n4 B 0.015122f
C334 VTAIL.n5 B 0.026578f
C335 VTAIL.n6 B 0.014282f
C336 VTAIL.n7 B 0.033757f
C337 VTAIL.n8 B 0.015122f
C338 VTAIL.n9 B 0.026578f
C339 VTAIL.n10 B 0.014282f
C340 VTAIL.n11 B 0.033757f
C341 VTAIL.n12 B 0.015122f
C342 VTAIL.n13 B 0.026578f
C343 VTAIL.n14 B 0.014282f
C344 VTAIL.n15 B 0.033757f
C345 VTAIL.n16 B 0.015122f
C346 VTAIL.n17 B 0.026578f
C347 VTAIL.n18 B 0.014282f
C348 VTAIL.n19 B 0.033757f
C349 VTAIL.n20 B 0.015122f
C350 VTAIL.n21 B 0.026578f
C351 VTAIL.n22 B 0.014282f
C352 VTAIL.n23 B 0.025317f
C353 VTAIL.n24 B 0.019941f
C354 VTAIL.t2 B 0.055442f
C355 VTAIL.n25 B 0.157352f
C356 VTAIL.n26 B 1.43684f
C357 VTAIL.n27 B 0.014282f
C358 VTAIL.n28 B 0.015122f
C359 VTAIL.n29 B 0.033757f
C360 VTAIL.n30 B 0.033757f
C361 VTAIL.n31 B 0.015122f
C362 VTAIL.n32 B 0.014282f
C363 VTAIL.n33 B 0.026578f
C364 VTAIL.n34 B 0.026578f
C365 VTAIL.n35 B 0.014282f
C366 VTAIL.n36 B 0.015122f
C367 VTAIL.n37 B 0.033757f
C368 VTAIL.n38 B 0.033757f
C369 VTAIL.n39 B 0.015122f
C370 VTAIL.n40 B 0.014282f
C371 VTAIL.n41 B 0.026578f
C372 VTAIL.n42 B 0.026578f
C373 VTAIL.n43 B 0.014282f
C374 VTAIL.n44 B 0.015122f
C375 VTAIL.n45 B 0.033757f
C376 VTAIL.n46 B 0.033757f
C377 VTAIL.n47 B 0.015122f
C378 VTAIL.n48 B 0.014282f
C379 VTAIL.n49 B 0.026578f
C380 VTAIL.n50 B 0.026578f
C381 VTAIL.n51 B 0.014282f
C382 VTAIL.n52 B 0.015122f
C383 VTAIL.n53 B 0.033757f
C384 VTAIL.n54 B 0.033757f
C385 VTAIL.n55 B 0.015122f
C386 VTAIL.n56 B 0.014282f
C387 VTAIL.n57 B 0.026578f
C388 VTAIL.n58 B 0.026578f
C389 VTAIL.n59 B 0.014282f
C390 VTAIL.n60 B 0.015122f
C391 VTAIL.n61 B 0.033757f
C392 VTAIL.n62 B 0.033757f
C393 VTAIL.n63 B 0.015122f
C394 VTAIL.n64 B 0.014282f
C395 VTAIL.n65 B 0.026578f
C396 VTAIL.n66 B 0.06579f
C397 VTAIL.n67 B 0.014282f
C398 VTAIL.n68 B 0.015122f
C399 VTAIL.n69 B 0.066735f
C400 VTAIL.n70 B 0.055225f
C401 VTAIL.n71 B 0.146935f
C402 VTAIL.t3 B 0.264631f
C403 VTAIL.t0 B 0.264631f
C404 VTAIL.n72 B 2.3005f
C405 VTAIL.n73 B 1.70414f
C406 VTAIL.t9 B 0.264631f
C407 VTAIL.t8 B 0.264631f
C408 VTAIL.n74 B 2.3005f
C409 VTAIL.n75 B 1.70415f
C410 VTAIL.n76 B 0.014936f
C411 VTAIL.n77 B 0.033757f
C412 VTAIL.n78 B 0.015122f
C413 VTAIL.n79 B 0.026578f
C414 VTAIL.n80 B 0.014282f
C415 VTAIL.n81 B 0.033757f
C416 VTAIL.n82 B 0.015122f
C417 VTAIL.n83 B 0.026578f
C418 VTAIL.n84 B 0.014282f
C419 VTAIL.n85 B 0.033757f
C420 VTAIL.n86 B 0.015122f
C421 VTAIL.n87 B 0.026578f
C422 VTAIL.n88 B 0.014282f
C423 VTAIL.n89 B 0.033757f
C424 VTAIL.n90 B 0.015122f
C425 VTAIL.n91 B 0.026578f
C426 VTAIL.n92 B 0.014282f
C427 VTAIL.n93 B 0.033757f
C428 VTAIL.n94 B 0.015122f
C429 VTAIL.n95 B 0.026578f
C430 VTAIL.n96 B 0.014282f
C431 VTAIL.n97 B 0.025317f
C432 VTAIL.n98 B 0.019941f
C433 VTAIL.t7 B 0.055442f
C434 VTAIL.n99 B 0.157352f
C435 VTAIL.n100 B 1.43684f
C436 VTAIL.n101 B 0.014282f
C437 VTAIL.n102 B 0.015122f
C438 VTAIL.n103 B 0.033757f
C439 VTAIL.n104 B 0.033757f
C440 VTAIL.n105 B 0.015122f
C441 VTAIL.n106 B 0.014282f
C442 VTAIL.n107 B 0.026578f
C443 VTAIL.n108 B 0.026578f
C444 VTAIL.n109 B 0.014282f
C445 VTAIL.n110 B 0.015122f
C446 VTAIL.n111 B 0.033757f
C447 VTAIL.n112 B 0.033757f
C448 VTAIL.n113 B 0.015122f
C449 VTAIL.n114 B 0.014282f
C450 VTAIL.n115 B 0.026578f
C451 VTAIL.n116 B 0.026578f
C452 VTAIL.n117 B 0.014282f
C453 VTAIL.n118 B 0.015122f
C454 VTAIL.n119 B 0.033757f
C455 VTAIL.n120 B 0.033757f
C456 VTAIL.n121 B 0.015122f
C457 VTAIL.n122 B 0.014282f
C458 VTAIL.n123 B 0.026578f
C459 VTAIL.n124 B 0.026578f
C460 VTAIL.n125 B 0.014282f
C461 VTAIL.n126 B 0.015122f
C462 VTAIL.n127 B 0.033757f
C463 VTAIL.n128 B 0.033757f
C464 VTAIL.n129 B 0.015122f
C465 VTAIL.n130 B 0.014282f
C466 VTAIL.n131 B 0.026578f
C467 VTAIL.n132 B 0.026578f
C468 VTAIL.n133 B 0.014282f
C469 VTAIL.n134 B 0.015122f
C470 VTAIL.n135 B 0.033757f
C471 VTAIL.n136 B 0.033757f
C472 VTAIL.n137 B 0.015122f
C473 VTAIL.n138 B 0.014282f
C474 VTAIL.n139 B 0.026578f
C475 VTAIL.n140 B 0.06579f
C476 VTAIL.n141 B 0.014282f
C477 VTAIL.n142 B 0.015122f
C478 VTAIL.n143 B 0.066735f
C479 VTAIL.n144 B 0.055225f
C480 VTAIL.n145 B 0.146935f
C481 VTAIL.t5 B 0.264631f
C482 VTAIL.t1 B 0.264631f
C483 VTAIL.n146 B 2.3005f
C484 VTAIL.n147 B 0.371193f
C485 VTAIL.n148 B 0.014936f
C486 VTAIL.n149 B 0.033757f
C487 VTAIL.n150 B 0.015122f
C488 VTAIL.n151 B 0.026578f
C489 VTAIL.n152 B 0.014282f
C490 VTAIL.n153 B 0.033757f
C491 VTAIL.n154 B 0.015122f
C492 VTAIL.n155 B 0.026578f
C493 VTAIL.n156 B 0.014282f
C494 VTAIL.n157 B 0.033757f
C495 VTAIL.n158 B 0.015122f
C496 VTAIL.n159 B 0.026578f
C497 VTAIL.n160 B 0.014282f
C498 VTAIL.n161 B 0.033757f
C499 VTAIL.n162 B 0.015122f
C500 VTAIL.n163 B 0.026578f
C501 VTAIL.n164 B 0.014282f
C502 VTAIL.n165 B 0.033757f
C503 VTAIL.n166 B 0.015122f
C504 VTAIL.n167 B 0.026578f
C505 VTAIL.n168 B 0.014282f
C506 VTAIL.n169 B 0.025317f
C507 VTAIL.n170 B 0.019941f
C508 VTAIL.t4 B 0.055442f
C509 VTAIL.n171 B 0.157352f
C510 VTAIL.n172 B 1.43684f
C511 VTAIL.n173 B 0.014282f
C512 VTAIL.n174 B 0.015122f
C513 VTAIL.n175 B 0.033757f
C514 VTAIL.n176 B 0.033757f
C515 VTAIL.n177 B 0.015122f
C516 VTAIL.n178 B 0.014282f
C517 VTAIL.n179 B 0.026578f
C518 VTAIL.n180 B 0.026578f
C519 VTAIL.n181 B 0.014282f
C520 VTAIL.n182 B 0.015122f
C521 VTAIL.n183 B 0.033757f
C522 VTAIL.n184 B 0.033757f
C523 VTAIL.n185 B 0.015122f
C524 VTAIL.n186 B 0.014282f
C525 VTAIL.n187 B 0.026578f
C526 VTAIL.n188 B 0.026578f
C527 VTAIL.n189 B 0.014282f
C528 VTAIL.n190 B 0.015122f
C529 VTAIL.n191 B 0.033757f
C530 VTAIL.n192 B 0.033757f
C531 VTAIL.n193 B 0.015122f
C532 VTAIL.n194 B 0.014282f
C533 VTAIL.n195 B 0.026578f
C534 VTAIL.n196 B 0.026578f
C535 VTAIL.n197 B 0.014282f
C536 VTAIL.n198 B 0.015122f
C537 VTAIL.n199 B 0.033757f
C538 VTAIL.n200 B 0.033757f
C539 VTAIL.n201 B 0.015122f
C540 VTAIL.n202 B 0.014282f
C541 VTAIL.n203 B 0.026578f
C542 VTAIL.n204 B 0.026578f
C543 VTAIL.n205 B 0.014282f
C544 VTAIL.n206 B 0.015122f
C545 VTAIL.n207 B 0.033757f
C546 VTAIL.n208 B 0.033757f
C547 VTAIL.n209 B 0.015122f
C548 VTAIL.n210 B 0.014282f
C549 VTAIL.n211 B 0.026578f
C550 VTAIL.n212 B 0.06579f
C551 VTAIL.n213 B 0.014282f
C552 VTAIL.n214 B 0.015122f
C553 VTAIL.n215 B 0.066735f
C554 VTAIL.n216 B 0.055225f
C555 VTAIL.n217 B 1.42526f
C556 VTAIL.n218 B 0.014936f
C557 VTAIL.n219 B 0.033757f
C558 VTAIL.n220 B 0.015122f
C559 VTAIL.n221 B 0.026578f
C560 VTAIL.n222 B 0.014282f
C561 VTAIL.n223 B 0.033757f
C562 VTAIL.n224 B 0.015122f
C563 VTAIL.n225 B 0.026578f
C564 VTAIL.n226 B 0.014282f
C565 VTAIL.n227 B 0.033757f
C566 VTAIL.n228 B 0.015122f
C567 VTAIL.n229 B 0.026578f
C568 VTAIL.n230 B 0.014282f
C569 VTAIL.n231 B 0.033757f
C570 VTAIL.n232 B 0.015122f
C571 VTAIL.n233 B 0.026578f
C572 VTAIL.n234 B 0.014282f
C573 VTAIL.n235 B 0.033757f
C574 VTAIL.n236 B 0.015122f
C575 VTAIL.n237 B 0.026578f
C576 VTAIL.n238 B 0.014282f
C577 VTAIL.n239 B 0.025317f
C578 VTAIL.n240 B 0.019941f
C579 VTAIL.t6 B 0.055442f
C580 VTAIL.n241 B 0.157352f
C581 VTAIL.n242 B 1.43684f
C582 VTAIL.n243 B 0.014282f
C583 VTAIL.n244 B 0.015122f
C584 VTAIL.n245 B 0.033757f
C585 VTAIL.n246 B 0.033757f
C586 VTAIL.n247 B 0.015122f
C587 VTAIL.n248 B 0.014282f
C588 VTAIL.n249 B 0.026578f
C589 VTAIL.n250 B 0.026578f
C590 VTAIL.n251 B 0.014282f
C591 VTAIL.n252 B 0.015122f
C592 VTAIL.n253 B 0.033757f
C593 VTAIL.n254 B 0.033757f
C594 VTAIL.n255 B 0.015122f
C595 VTAIL.n256 B 0.014282f
C596 VTAIL.n257 B 0.026578f
C597 VTAIL.n258 B 0.026578f
C598 VTAIL.n259 B 0.014282f
C599 VTAIL.n260 B 0.015122f
C600 VTAIL.n261 B 0.033757f
C601 VTAIL.n262 B 0.033757f
C602 VTAIL.n263 B 0.015122f
C603 VTAIL.n264 B 0.014282f
C604 VTAIL.n265 B 0.026578f
C605 VTAIL.n266 B 0.026578f
C606 VTAIL.n267 B 0.014282f
C607 VTAIL.n268 B 0.015122f
C608 VTAIL.n269 B 0.033757f
C609 VTAIL.n270 B 0.033757f
C610 VTAIL.n271 B 0.015122f
C611 VTAIL.n272 B 0.014282f
C612 VTAIL.n273 B 0.026578f
C613 VTAIL.n274 B 0.026578f
C614 VTAIL.n275 B 0.014282f
C615 VTAIL.n276 B 0.015122f
C616 VTAIL.n277 B 0.033757f
C617 VTAIL.n278 B 0.033757f
C618 VTAIL.n279 B 0.015122f
C619 VTAIL.n280 B 0.014282f
C620 VTAIL.n281 B 0.026578f
C621 VTAIL.n282 B 0.06579f
C622 VTAIL.n283 B 0.014282f
C623 VTAIL.n284 B 0.015122f
C624 VTAIL.n285 B 0.066735f
C625 VTAIL.n286 B 0.055225f
C626 VTAIL.n287 B 1.40662f
C627 VN.t4 B 0.804527f
C628 VN.n0 B 0.313135f
C629 VN.t1 B 0.795578f
C630 VN.n1 B 0.329183f
C631 VN.t5 B 0.797457f
C632 VN.n2 B 0.319805f
C633 VN.n3 B 0.162588f
C634 VN.t2 B 0.804527f
C635 VN.n4 B 0.313135f
C636 VN.t0 B 0.797457f
C637 VN.t3 B 0.795578f
C638 VN.n5 B 0.329183f
C639 VN.n6 B 0.319805f
C640 VN.n7 B 2.26389f
.ends

