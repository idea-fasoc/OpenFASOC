* NGSPICE file created from diff_pair_sample_0800.ext - technology: sky130A

.subckt diff_pair_sample_0800 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t0 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=4.9647 pd=26.24 as=2.10045 ps=13.06 w=12.73 l=3.61
X1 B.t11 B.t9 B.t10 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=4.9647 pd=26.24 as=0 ps=0 w=12.73 l=3.61
X2 B.t8 B.t6 B.t7 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=4.9647 pd=26.24 as=0 ps=0 w=12.73 l=3.61
X3 VDD1.t1 VP.t1 VTAIL.t6 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=2.10045 pd=13.06 as=4.9647 ps=26.24 w=12.73 l=3.61
X4 B.t5 B.t3 B.t4 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=4.9647 pd=26.24 as=0 ps=0 w=12.73 l=3.61
X5 VTAIL.t5 VP.t2 VDD1.t2 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=4.9647 pd=26.24 as=2.10045 ps=13.06 w=12.73 l=3.61
X6 VDD2.t3 VN.t0 VTAIL.t2 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=2.10045 pd=13.06 as=4.9647 ps=26.24 w=12.73 l=3.61
X7 B.t2 B.t0 B.t1 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=4.9647 pd=26.24 as=0 ps=0 w=12.73 l=3.61
X8 VDD1.t3 VP.t3 VTAIL.t4 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=2.10045 pd=13.06 as=4.9647 ps=26.24 w=12.73 l=3.61
X9 VTAIL.t3 VN.t1 VDD2.t2 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=4.9647 pd=26.24 as=2.10045 ps=13.06 w=12.73 l=3.61
X10 VDD2.t1 VN.t2 VTAIL.t0 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=2.10045 pd=13.06 as=4.9647 ps=26.24 w=12.73 l=3.61
X11 VTAIL.t1 VN.t3 VDD2.t0 w_n3334_n3514# sky130_fd_pr__pfet_01v8 ad=4.9647 pd=26.24 as=2.10045 ps=13.06 w=12.73 l=3.61
R0 VP.n19 VP.n18 161.3
R1 VP.n17 VP.n1 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n14 VP.n2 161.3
R4 VP.n13 VP.n12 161.3
R5 VP.n11 VP.n3 161.3
R6 VP.n10 VP.n9 161.3
R7 VP.n8 VP.n4 161.3
R8 VP.n5 VP.t0 119.895
R9 VP.n5 VP.t3 118.65
R10 VP.n6 VP.t2 84.9847
R11 VP.n0 VP.t1 84.9847
R12 VP.n7 VP.n6 79.3019
R13 VP.n20 VP.n0 79.3019
R14 VP.n12 VP.n2 56.5193
R15 VP.n7 VP.n5 52.1546
R16 VP.n10 VP.n4 24.4675
R17 VP.n11 VP.n10 24.4675
R18 VP.n12 VP.n11 24.4675
R19 VP.n16 VP.n2 24.4675
R20 VP.n17 VP.n16 24.4675
R21 VP.n18 VP.n17 24.4675
R22 VP.n6 VP.n4 10.766
R23 VP.n18 VP.n0 10.766
R24 VP.n8 VP.n7 0.354971
R25 VP.n20 VP.n19 0.354971
R26 VP VP.n20 0.26696
R27 VP.n9 VP.n8 0.189894
R28 VP.n9 VP.n3 0.189894
R29 VP.n13 VP.n3 0.189894
R30 VP.n14 VP.n13 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n15 VP.n1 0.189894
R33 VP.n19 VP.n1 0.189894
R34 VDD1 VDD1.n1 116.281
R35 VDD1 VDD1.n0 70.936
R36 VDD1.n0 VDD1.t0 2.55392
R37 VDD1.n0 VDD1.t3 2.55392
R38 VDD1.n1 VDD1.t2 2.55392
R39 VDD1.n1 VDD1.t1 2.55392
R40 VTAIL.n554 VTAIL.n490 756.745
R41 VTAIL.n64 VTAIL.n0 756.745
R42 VTAIL.n134 VTAIL.n70 756.745
R43 VTAIL.n204 VTAIL.n140 756.745
R44 VTAIL.n484 VTAIL.n420 756.745
R45 VTAIL.n414 VTAIL.n350 756.745
R46 VTAIL.n344 VTAIL.n280 756.745
R47 VTAIL.n274 VTAIL.n210 756.745
R48 VTAIL.n513 VTAIL.n512 585
R49 VTAIL.n510 VTAIL.n509 585
R50 VTAIL.n519 VTAIL.n518 585
R51 VTAIL.n521 VTAIL.n520 585
R52 VTAIL.n506 VTAIL.n505 585
R53 VTAIL.n527 VTAIL.n526 585
R54 VTAIL.n530 VTAIL.n529 585
R55 VTAIL.n528 VTAIL.n502 585
R56 VTAIL.n535 VTAIL.n501 585
R57 VTAIL.n537 VTAIL.n536 585
R58 VTAIL.n539 VTAIL.n538 585
R59 VTAIL.n498 VTAIL.n497 585
R60 VTAIL.n545 VTAIL.n544 585
R61 VTAIL.n547 VTAIL.n546 585
R62 VTAIL.n494 VTAIL.n493 585
R63 VTAIL.n553 VTAIL.n552 585
R64 VTAIL.n555 VTAIL.n554 585
R65 VTAIL.n23 VTAIL.n22 585
R66 VTAIL.n20 VTAIL.n19 585
R67 VTAIL.n29 VTAIL.n28 585
R68 VTAIL.n31 VTAIL.n30 585
R69 VTAIL.n16 VTAIL.n15 585
R70 VTAIL.n37 VTAIL.n36 585
R71 VTAIL.n40 VTAIL.n39 585
R72 VTAIL.n38 VTAIL.n12 585
R73 VTAIL.n45 VTAIL.n11 585
R74 VTAIL.n47 VTAIL.n46 585
R75 VTAIL.n49 VTAIL.n48 585
R76 VTAIL.n8 VTAIL.n7 585
R77 VTAIL.n55 VTAIL.n54 585
R78 VTAIL.n57 VTAIL.n56 585
R79 VTAIL.n4 VTAIL.n3 585
R80 VTAIL.n63 VTAIL.n62 585
R81 VTAIL.n65 VTAIL.n64 585
R82 VTAIL.n93 VTAIL.n92 585
R83 VTAIL.n90 VTAIL.n89 585
R84 VTAIL.n99 VTAIL.n98 585
R85 VTAIL.n101 VTAIL.n100 585
R86 VTAIL.n86 VTAIL.n85 585
R87 VTAIL.n107 VTAIL.n106 585
R88 VTAIL.n110 VTAIL.n109 585
R89 VTAIL.n108 VTAIL.n82 585
R90 VTAIL.n115 VTAIL.n81 585
R91 VTAIL.n117 VTAIL.n116 585
R92 VTAIL.n119 VTAIL.n118 585
R93 VTAIL.n78 VTAIL.n77 585
R94 VTAIL.n125 VTAIL.n124 585
R95 VTAIL.n127 VTAIL.n126 585
R96 VTAIL.n74 VTAIL.n73 585
R97 VTAIL.n133 VTAIL.n132 585
R98 VTAIL.n135 VTAIL.n134 585
R99 VTAIL.n163 VTAIL.n162 585
R100 VTAIL.n160 VTAIL.n159 585
R101 VTAIL.n169 VTAIL.n168 585
R102 VTAIL.n171 VTAIL.n170 585
R103 VTAIL.n156 VTAIL.n155 585
R104 VTAIL.n177 VTAIL.n176 585
R105 VTAIL.n180 VTAIL.n179 585
R106 VTAIL.n178 VTAIL.n152 585
R107 VTAIL.n185 VTAIL.n151 585
R108 VTAIL.n187 VTAIL.n186 585
R109 VTAIL.n189 VTAIL.n188 585
R110 VTAIL.n148 VTAIL.n147 585
R111 VTAIL.n195 VTAIL.n194 585
R112 VTAIL.n197 VTAIL.n196 585
R113 VTAIL.n144 VTAIL.n143 585
R114 VTAIL.n203 VTAIL.n202 585
R115 VTAIL.n205 VTAIL.n204 585
R116 VTAIL.n485 VTAIL.n484 585
R117 VTAIL.n483 VTAIL.n482 585
R118 VTAIL.n424 VTAIL.n423 585
R119 VTAIL.n477 VTAIL.n476 585
R120 VTAIL.n475 VTAIL.n474 585
R121 VTAIL.n428 VTAIL.n427 585
R122 VTAIL.n469 VTAIL.n468 585
R123 VTAIL.n467 VTAIL.n466 585
R124 VTAIL.n465 VTAIL.n431 585
R125 VTAIL.n435 VTAIL.n432 585
R126 VTAIL.n460 VTAIL.n459 585
R127 VTAIL.n458 VTAIL.n457 585
R128 VTAIL.n437 VTAIL.n436 585
R129 VTAIL.n452 VTAIL.n451 585
R130 VTAIL.n450 VTAIL.n449 585
R131 VTAIL.n441 VTAIL.n440 585
R132 VTAIL.n444 VTAIL.n443 585
R133 VTAIL.n415 VTAIL.n414 585
R134 VTAIL.n413 VTAIL.n412 585
R135 VTAIL.n354 VTAIL.n353 585
R136 VTAIL.n407 VTAIL.n406 585
R137 VTAIL.n405 VTAIL.n404 585
R138 VTAIL.n358 VTAIL.n357 585
R139 VTAIL.n399 VTAIL.n398 585
R140 VTAIL.n397 VTAIL.n396 585
R141 VTAIL.n395 VTAIL.n361 585
R142 VTAIL.n365 VTAIL.n362 585
R143 VTAIL.n390 VTAIL.n389 585
R144 VTAIL.n388 VTAIL.n387 585
R145 VTAIL.n367 VTAIL.n366 585
R146 VTAIL.n382 VTAIL.n381 585
R147 VTAIL.n380 VTAIL.n379 585
R148 VTAIL.n371 VTAIL.n370 585
R149 VTAIL.n374 VTAIL.n373 585
R150 VTAIL.n345 VTAIL.n344 585
R151 VTAIL.n343 VTAIL.n342 585
R152 VTAIL.n284 VTAIL.n283 585
R153 VTAIL.n337 VTAIL.n336 585
R154 VTAIL.n335 VTAIL.n334 585
R155 VTAIL.n288 VTAIL.n287 585
R156 VTAIL.n329 VTAIL.n328 585
R157 VTAIL.n327 VTAIL.n326 585
R158 VTAIL.n325 VTAIL.n291 585
R159 VTAIL.n295 VTAIL.n292 585
R160 VTAIL.n320 VTAIL.n319 585
R161 VTAIL.n318 VTAIL.n317 585
R162 VTAIL.n297 VTAIL.n296 585
R163 VTAIL.n312 VTAIL.n311 585
R164 VTAIL.n310 VTAIL.n309 585
R165 VTAIL.n301 VTAIL.n300 585
R166 VTAIL.n304 VTAIL.n303 585
R167 VTAIL.n275 VTAIL.n274 585
R168 VTAIL.n273 VTAIL.n272 585
R169 VTAIL.n214 VTAIL.n213 585
R170 VTAIL.n267 VTAIL.n266 585
R171 VTAIL.n265 VTAIL.n264 585
R172 VTAIL.n218 VTAIL.n217 585
R173 VTAIL.n259 VTAIL.n258 585
R174 VTAIL.n257 VTAIL.n256 585
R175 VTAIL.n255 VTAIL.n221 585
R176 VTAIL.n225 VTAIL.n222 585
R177 VTAIL.n250 VTAIL.n249 585
R178 VTAIL.n248 VTAIL.n247 585
R179 VTAIL.n227 VTAIL.n226 585
R180 VTAIL.n242 VTAIL.n241 585
R181 VTAIL.n240 VTAIL.n239 585
R182 VTAIL.n231 VTAIL.n230 585
R183 VTAIL.n234 VTAIL.n233 585
R184 VTAIL.t0 VTAIL.n511 329.036
R185 VTAIL.t3 VTAIL.n21 329.036
R186 VTAIL.t6 VTAIL.n91 329.036
R187 VTAIL.t5 VTAIL.n161 329.036
R188 VTAIL.t4 VTAIL.n442 329.036
R189 VTAIL.t7 VTAIL.n372 329.036
R190 VTAIL.t2 VTAIL.n302 329.036
R191 VTAIL.t1 VTAIL.n232 329.036
R192 VTAIL.n512 VTAIL.n509 171.744
R193 VTAIL.n519 VTAIL.n509 171.744
R194 VTAIL.n520 VTAIL.n519 171.744
R195 VTAIL.n520 VTAIL.n505 171.744
R196 VTAIL.n527 VTAIL.n505 171.744
R197 VTAIL.n529 VTAIL.n527 171.744
R198 VTAIL.n529 VTAIL.n528 171.744
R199 VTAIL.n528 VTAIL.n501 171.744
R200 VTAIL.n537 VTAIL.n501 171.744
R201 VTAIL.n538 VTAIL.n537 171.744
R202 VTAIL.n538 VTAIL.n497 171.744
R203 VTAIL.n545 VTAIL.n497 171.744
R204 VTAIL.n546 VTAIL.n545 171.744
R205 VTAIL.n546 VTAIL.n493 171.744
R206 VTAIL.n553 VTAIL.n493 171.744
R207 VTAIL.n554 VTAIL.n553 171.744
R208 VTAIL.n22 VTAIL.n19 171.744
R209 VTAIL.n29 VTAIL.n19 171.744
R210 VTAIL.n30 VTAIL.n29 171.744
R211 VTAIL.n30 VTAIL.n15 171.744
R212 VTAIL.n37 VTAIL.n15 171.744
R213 VTAIL.n39 VTAIL.n37 171.744
R214 VTAIL.n39 VTAIL.n38 171.744
R215 VTAIL.n38 VTAIL.n11 171.744
R216 VTAIL.n47 VTAIL.n11 171.744
R217 VTAIL.n48 VTAIL.n47 171.744
R218 VTAIL.n48 VTAIL.n7 171.744
R219 VTAIL.n55 VTAIL.n7 171.744
R220 VTAIL.n56 VTAIL.n55 171.744
R221 VTAIL.n56 VTAIL.n3 171.744
R222 VTAIL.n63 VTAIL.n3 171.744
R223 VTAIL.n64 VTAIL.n63 171.744
R224 VTAIL.n92 VTAIL.n89 171.744
R225 VTAIL.n99 VTAIL.n89 171.744
R226 VTAIL.n100 VTAIL.n99 171.744
R227 VTAIL.n100 VTAIL.n85 171.744
R228 VTAIL.n107 VTAIL.n85 171.744
R229 VTAIL.n109 VTAIL.n107 171.744
R230 VTAIL.n109 VTAIL.n108 171.744
R231 VTAIL.n108 VTAIL.n81 171.744
R232 VTAIL.n117 VTAIL.n81 171.744
R233 VTAIL.n118 VTAIL.n117 171.744
R234 VTAIL.n118 VTAIL.n77 171.744
R235 VTAIL.n125 VTAIL.n77 171.744
R236 VTAIL.n126 VTAIL.n125 171.744
R237 VTAIL.n126 VTAIL.n73 171.744
R238 VTAIL.n133 VTAIL.n73 171.744
R239 VTAIL.n134 VTAIL.n133 171.744
R240 VTAIL.n162 VTAIL.n159 171.744
R241 VTAIL.n169 VTAIL.n159 171.744
R242 VTAIL.n170 VTAIL.n169 171.744
R243 VTAIL.n170 VTAIL.n155 171.744
R244 VTAIL.n177 VTAIL.n155 171.744
R245 VTAIL.n179 VTAIL.n177 171.744
R246 VTAIL.n179 VTAIL.n178 171.744
R247 VTAIL.n178 VTAIL.n151 171.744
R248 VTAIL.n187 VTAIL.n151 171.744
R249 VTAIL.n188 VTAIL.n187 171.744
R250 VTAIL.n188 VTAIL.n147 171.744
R251 VTAIL.n195 VTAIL.n147 171.744
R252 VTAIL.n196 VTAIL.n195 171.744
R253 VTAIL.n196 VTAIL.n143 171.744
R254 VTAIL.n203 VTAIL.n143 171.744
R255 VTAIL.n204 VTAIL.n203 171.744
R256 VTAIL.n484 VTAIL.n483 171.744
R257 VTAIL.n483 VTAIL.n423 171.744
R258 VTAIL.n476 VTAIL.n423 171.744
R259 VTAIL.n476 VTAIL.n475 171.744
R260 VTAIL.n475 VTAIL.n427 171.744
R261 VTAIL.n468 VTAIL.n427 171.744
R262 VTAIL.n468 VTAIL.n467 171.744
R263 VTAIL.n467 VTAIL.n431 171.744
R264 VTAIL.n435 VTAIL.n431 171.744
R265 VTAIL.n459 VTAIL.n435 171.744
R266 VTAIL.n459 VTAIL.n458 171.744
R267 VTAIL.n458 VTAIL.n436 171.744
R268 VTAIL.n451 VTAIL.n436 171.744
R269 VTAIL.n451 VTAIL.n450 171.744
R270 VTAIL.n450 VTAIL.n440 171.744
R271 VTAIL.n443 VTAIL.n440 171.744
R272 VTAIL.n414 VTAIL.n413 171.744
R273 VTAIL.n413 VTAIL.n353 171.744
R274 VTAIL.n406 VTAIL.n353 171.744
R275 VTAIL.n406 VTAIL.n405 171.744
R276 VTAIL.n405 VTAIL.n357 171.744
R277 VTAIL.n398 VTAIL.n357 171.744
R278 VTAIL.n398 VTAIL.n397 171.744
R279 VTAIL.n397 VTAIL.n361 171.744
R280 VTAIL.n365 VTAIL.n361 171.744
R281 VTAIL.n389 VTAIL.n365 171.744
R282 VTAIL.n389 VTAIL.n388 171.744
R283 VTAIL.n388 VTAIL.n366 171.744
R284 VTAIL.n381 VTAIL.n366 171.744
R285 VTAIL.n381 VTAIL.n380 171.744
R286 VTAIL.n380 VTAIL.n370 171.744
R287 VTAIL.n373 VTAIL.n370 171.744
R288 VTAIL.n344 VTAIL.n343 171.744
R289 VTAIL.n343 VTAIL.n283 171.744
R290 VTAIL.n336 VTAIL.n283 171.744
R291 VTAIL.n336 VTAIL.n335 171.744
R292 VTAIL.n335 VTAIL.n287 171.744
R293 VTAIL.n328 VTAIL.n287 171.744
R294 VTAIL.n328 VTAIL.n327 171.744
R295 VTAIL.n327 VTAIL.n291 171.744
R296 VTAIL.n295 VTAIL.n291 171.744
R297 VTAIL.n319 VTAIL.n295 171.744
R298 VTAIL.n319 VTAIL.n318 171.744
R299 VTAIL.n318 VTAIL.n296 171.744
R300 VTAIL.n311 VTAIL.n296 171.744
R301 VTAIL.n311 VTAIL.n310 171.744
R302 VTAIL.n310 VTAIL.n300 171.744
R303 VTAIL.n303 VTAIL.n300 171.744
R304 VTAIL.n274 VTAIL.n273 171.744
R305 VTAIL.n273 VTAIL.n213 171.744
R306 VTAIL.n266 VTAIL.n213 171.744
R307 VTAIL.n266 VTAIL.n265 171.744
R308 VTAIL.n265 VTAIL.n217 171.744
R309 VTAIL.n258 VTAIL.n217 171.744
R310 VTAIL.n258 VTAIL.n257 171.744
R311 VTAIL.n257 VTAIL.n221 171.744
R312 VTAIL.n225 VTAIL.n221 171.744
R313 VTAIL.n249 VTAIL.n225 171.744
R314 VTAIL.n249 VTAIL.n248 171.744
R315 VTAIL.n248 VTAIL.n226 171.744
R316 VTAIL.n241 VTAIL.n226 171.744
R317 VTAIL.n241 VTAIL.n240 171.744
R318 VTAIL.n240 VTAIL.n230 171.744
R319 VTAIL.n233 VTAIL.n230 171.744
R320 VTAIL.n512 VTAIL.t0 85.8723
R321 VTAIL.n22 VTAIL.t3 85.8723
R322 VTAIL.n92 VTAIL.t6 85.8723
R323 VTAIL.n162 VTAIL.t5 85.8723
R324 VTAIL.n443 VTAIL.t4 85.8723
R325 VTAIL.n373 VTAIL.t7 85.8723
R326 VTAIL.n303 VTAIL.t2 85.8723
R327 VTAIL.n233 VTAIL.t1 85.8723
R328 VTAIL.n559 VTAIL.n558 30.052
R329 VTAIL.n69 VTAIL.n68 30.052
R330 VTAIL.n139 VTAIL.n138 30.052
R331 VTAIL.n209 VTAIL.n208 30.052
R332 VTAIL.n489 VTAIL.n488 30.052
R333 VTAIL.n419 VTAIL.n418 30.052
R334 VTAIL.n349 VTAIL.n348 30.052
R335 VTAIL.n279 VTAIL.n278 30.052
R336 VTAIL.n559 VTAIL.n489 26.7376
R337 VTAIL.n279 VTAIL.n209 26.7376
R338 VTAIL.n536 VTAIL.n535 13.1884
R339 VTAIL.n46 VTAIL.n45 13.1884
R340 VTAIL.n116 VTAIL.n115 13.1884
R341 VTAIL.n186 VTAIL.n185 13.1884
R342 VTAIL.n466 VTAIL.n465 13.1884
R343 VTAIL.n396 VTAIL.n395 13.1884
R344 VTAIL.n326 VTAIL.n325 13.1884
R345 VTAIL.n256 VTAIL.n255 13.1884
R346 VTAIL.n534 VTAIL.n502 12.8005
R347 VTAIL.n539 VTAIL.n500 12.8005
R348 VTAIL.n44 VTAIL.n12 12.8005
R349 VTAIL.n49 VTAIL.n10 12.8005
R350 VTAIL.n114 VTAIL.n82 12.8005
R351 VTAIL.n119 VTAIL.n80 12.8005
R352 VTAIL.n184 VTAIL.n152 12.8005
R353 VTAIL.n189 VTAIL.n150 12.8005
R354 VTAIL.n469 VTAIL.n430 12.8005
R355 VTAIL.n464 VTAIL.n432 12.8005
R356 VTAIL.n399 VTAIL.n360 12.8005
R357 VTAIL.n394 VTAIL.n362 12.8005
R358 VTAIL.n329 VTAIL.n290 12.8005
R359 VTAIL.n324 VTAIL.n292 12.8005
R360 VTAIL.n259 VTAIL.n220 12.8005
R361 VTAIL.n254 VTAIL.n222 12.8005
R362 VTAIL.n531 VTAIL.n530 12.0247
R363 VTAIL.n540 VTAIL.n498 12.0247
R364 VTAIL.n41 VTAIL.n40 12.0247
R365 VTAIL.n50 VTAIL.n8 12.0247
R366 VTAIL.n111 VTAIL.n110 12.0247
R367 VTAIL.n120 VTAIL.n78 12.0247
R368 VTAIL.n181 VTAIL.n180 12.0247
R369 VTAIL.n190 VTAIL.n148 12.0247
R370 VTAIL.n470 VTAIL.n428 12.0247
R371 VTAIL.n461 VTAIL.n460 12.0247
R372 VTAIL.n400 VTAIL.n358 12.0247
R373 VTAIL.n391 VTAIL.n390 12.0247
R374 VTAIL.n330 VTAIL.n288 12.0247
R375 VTAIL.n321 VTAIL.n320 12.0247
R376 VTAIL.n260 VTAIL.n218 12.0247
R377 VTAIL.n251 VTAIL.n250 12.0247
R378 VTAIL.n526 VTAIL.n504 11.249
R379 VTAIL.n544 VTAIL.n543 11.249
R380 VTAIL.n36 VTAIL.n14 11.249
R381 VTAIL.n54 VTAIL.n53 11.249
R382 VTAIL.n106 VTAIL.n84 11.249
R383 VTAIL.n124 VTAIL.n123 11.249
R384 VTAIL.n176 VTAIL.n154 11.249
R385 VTAIL.n194 VTAIL.n193 11.249
R386 VTAIL.n474 VTAIL.n473 11.249
R387 VTAIL.n457 VTAIL.n434 11.249
R388 VTAIL.n404 VTAIL.n403 11.249
R389 VTAIL.n387 VTAIL.n364 11.249
R390 VTAIL.n334 VTAIL.n333 11.249
R391 VTAIL.n317 VTAIL.n294 11.249
R392 VTAIL.n264 VTAIL.n263 11.249
R393 VTAIL.n247 VTAIL.n224 11.249
R394 VTAIL.n513 VTAIL.n511 10.7239
R395 VTAIL.n23 VTAIL.n21 10.7239
R396 VTAIL.n93 VTAIL.n91 10.7239
R397 VTAIL.n163 VTAIL.n161 10.7239
R398 VTAIL.n444 VTAIL.n442 10.7239
R399 VTAIL.n374 VTAIL.n372 10.7239
R400 VTAIL.n304 VTAIL.n302 10.7239
R401 VTAIL.n234 VTAIL.n232 10.7239
R402 VTAIL.n525 VTAIL.n506 10.4732
R403 VTAIL.n547 VTAIL.n496 10.4732
R404 VTAIL.n35 VTAIL.n16 10.4732
R405 VTAIL.n57 VTAIL.n6 10.4732
R406 VTAIL.n105 VTAIL.n86 10.4732
R407 VTAIL.n127 VTAIL.n76 10.4732
R408 VTAIL.n175 VTAIL.n156 10.4732
R409 VTAIL.n197 VTAIL.n146 10.4732
R410 VTAIL.n477 VTAIL.n426 10.4732
R411 VTAIL.n456 VTAIL.n437 10.4732
R412 VTAIL.n407 VTAIL.n356 10.4732
R413 VTAIL.n386 VTAIL.n367 10.4732
R414 VTAIL.n337 VTAIL.n286 10.4732
R415 VTAIL.n316 VTAIL.n297 10.4732
R416 VTAIL.n267 VTAIL.n216 10.4732
R417 VTAIL.n246 VTAIL.n227 10.4732
R418 VTAIL.n522 VTAIL.n521 9.69747
R419 VTAIL.n548 VTAIL.n494 9.69747
R420 VTAIL.n32 VTAIL.n31 9.69747
R421 VTAIL.n58 VTAIL.n4 9.69747
R422 VTAIL.n102 VTAIL.n101 9.69747
R423 VTAIL.n128 VTAIL.n74 9.69747
R424 VTAIL.n172 VTAIL.n171 9.69747
R425 VTAIL.n198 VTAIL.n144 9.69747
R426 VTAIL.n478 VTAIL.n424 9.69747
R427 VTAIL.n453 VTAIL.n452 9.69747
R428 VTAIL.n408 VTAIL.n354 9.69747
R429 VTAIL.n383 VTAIL.n382 9.69747
R430 VTAIL.n338 VTAIL.n284 9.69747
R431 VTAIL.n313 VTAIL.n312 9.69747
R432 VTAIL.n268 VTAIL.n214 9.69747
R433 VTAIL.n243 VTAIL.n242 9.69747
R434 VTAIL.n558 VTAIL.n557 9.45567
R435 VTAIL.n68 VTAIL.n67 9.45567
R436 VTAIL.n138 VTAIL.n137 9.45567
R437 VTAIL.n208 VTAIL.n207 9.45567
R438 VTAIL.n488 VTAIL.n487 9.45567
R439 VTAIL.n418 VTAIL.n417 9.45567
R440 VTAIL.n348 VTAIL.n347 9.45567
R441 VTAIL.n278 VTAIL.n277 9.45567
R442 VTAIL.n492 VTAIL.n491 9.3005
R443 VTAIL.n551 VTAIL.n550 9.3005
R444 VTAIL.n549 VTAIL.n548 9.3005
R445 VTAIL.n496 VTAIL.n495 9.3005
R446 VTAIL.n543 VTAIL.n542 9.3005
R447 VTAIL.n541 VTAIL.n540 9.3005
R448 VTAIL.n500 VTAIL.n499 9.3005
R449 VTAIL.n515 VTAIL.n514 9.3005
R450 VTAIL.n517 VTAIL.n516 9.3005
R451 VTAIL.n508 VTAIL.n507 9.3005
R452 VTAIL.n523 VTAIL.n522 9.3005
R453 VTAIL.n525 VTAIL.n524 9.3005
R454 VTAIL.n504 VTAIL.n503 9.3005
R455 VTAIL.n532 VTAIL.n531 9.3005
R456 VTAIL.n534 VTAIL.n533 9.3005
R457 VTAIL.n557 VTAIL.n556 9.3005
R458 VTAIL.n2 VTAIL.n1 9.3005
R459 VTAIL.n61 VTAIL.n60 9.3005
R460 VTAIL.n59 VTAIL.n58 9.3005
R461 VTAIL.n6 VTAIL.n5 9.3005
R462 VTAIL.n53 VTAIL.n52 9.3005
R463 VTAIL.n51 VTAIL.n50 9.3005
R464 VTAIL.n10 VTAIL.n9 9.3005
R465 VTAIL.n25 VTAIL.n24 9.3005
R466 VTAIL.n27 VTAIL.n26 9.3005
R467 VTAIL.n18 VTAIL.n17 9.3005
R468 VTAIL.n33 VTAIL.n32 9.3005
R469 VTAIL.n35 VTAIL.n34 9.3005
R470 VTAIL.n14 VTAIL.n13 9.3005
R471 VTAIL.n42 VTAIL.n41 9.3005
R472 VTAIL.n44 VTAIL.n43 9.3005
R473 VTAIL.n67 VTAIL.n66 9.3005
R474 VTAIL.n72 VTAIL.n71 9.3005
R475 VTAIL.n131 VTAIL.n130 9.3005
R476 VTAIL.n129 VTAIL.n128 9.3005
R477 VTAIL.n76 VTAIL.n75 9.3005
R478 VTAIL.n123 VTAIL.n122 9.3005
R479 VTAIL.n121 VTAIL.n120 9.3005
R480 VTAIL.n80 VTAIL.n79 9.3005
R481 VTAIL.n95 VTAIL.n94 9.3005
R482 VTAIL.n97 VTAIL.n96 9.3005
R483 VTAIL.n88 VTAIL.n87 9.3005
R484 VTAIL.n103 VTAIL.n102 9.3005
R485 VTAIL.n105 VTAIL.n104 9.3005
R486 VTAIL.n84 VTAIL.n83 9.3005
R487 VTAIL.n112 VTAIL.n111 9.3005
R488 VTAIL.n114 VTAIL.n113 9.3005
R489 VTAIL.n137 VTAIL.n136 9.3005
R490 VTAIL.n142 VTAIL.n141 9.3005
R491 VTAIL.n201 VTAIL.n200 9.3005
R492 VTAIL.n199 VTAIL.n198 9.3005
R493 VTAIL.n146 VTAIL.n145 9.3005
R494 VTAIL.n193 VTAIL.n192 9.3005
R495 VTAIL.n191 VTAIL.n190 9.3005
R496 VTAIL.n150 VTAIL.n149 9.3005
R497 VTAIL.n165 VTAIL.n164 9.3005
R498 VTAIL.n167 VTAIL.n166 9.3005
R499 VTAIL.n158 VTAIL.n157 9.3005
R500 VTAIL.n173 VTAIL.n172 9.3005
R501 VTAIL.n175 VTAIL.n174 9.3005
R502 VTAIL.n154 VTAIL.n153 9.3005
R503 VTAIL.n182 VTAIL.n181 9.3005
R504 VTAIL.n184 VTAIL.n183 9.3005
R505 VTAIL.n207 VTAIL.n206 9.3005
R506 VTAIL.n446 VTAIL.n445 9.3005
R507 VTAIL.n448 VTAIL.n447 9.3005
R508 VTAIL.n439 VTAIL.n438 9.3005
R509 VTAIL.n454 VTAIL.n453 9.3005
R510 VTAIL.n456 VTAIL.n455 9.3005
R511 VTAIL.n434 VTAIL.n433 9.3005
R512 VTAIL.n462 VTAIL.n461 9.3005
R513 VTAIL.n464 VTAIL.n463 9.3005
R514 VTAIL.n487 VTAIL.n486 9.3005
R515 VTAIL.n422 VTAIL.n421 9.3005
R516 VTAIL.n481 VTAIL.n480 9.3005
R517 VTAIL.n479 VTAIL.n478 9.3005
R518 VTAIL.n426 VTAIL.n425 9.3005
R519 VTAIL.n473 VTAIL.n472 9.3005
R520 VTAIL.n471 VTAIL.n470 9.3005
R521 VTAIL.n430 VTAIL.n429 9.3005
R522 VTAIL.n376 VTAIL.n375 9.3005
R523 VTAIL.n378 VTAIL.n377 9.3005
R524 VTAIL.n369 VTAIL.n368 9.3005
R525 VTAIL.n384 VTAIL.n383 9.3005
R526 VTAIL.n386 VTAIL.n385 9.3005
R527 VTAIL.n364 VTAIL.n363 9.3005
R528 VTAIL.n392 VTAIL.n391 9.3005
R529 VTAIL.n394 VTAIL.n393 9.3005
R530 VTAIL.n417 VTAIL.n416 9.3005
R531 VTAIL.n352 VTAIL.n351 9.3005
R532 VTAIL.n411 VTAIL.n410 9.3005
R533 VTAIL.n409 VTAIL.n408 9.3005
R534 VTAIL.n356 VTAIL.n355 9.3005
R535 VTAIL.n403 VTAIL.n402 9.3005
R536 VTAIL.n401 VTAIL.n400 9.3005
R537 VTAIL.n360 VTAIL.n359 9.3005
R538 VTAIL.n306 VTAIL.n305 9.3005
R539 VTAIL.n308 VTAIL.n307 9.3005
R540 VTAIL.n299 VTAIL.n298 9.3005
R541 VTAIL.n314 VTAIL.n313 9.3005
R542 VTAIL.n316 VTAIL.n315 9.3005
R543 VTAIL.n294 VTAIL.n293 9.3005
R544 VTAIL.n322 VTAIL.n321 9.3005
R545 VTAIL.n324 VTAIL.n323 9.3005
R546 VTAIL.n347 VTAIL.n346 9.3005
R547 VTAIL.n282 VTAIL.n281 9.3005
R548 VTAIL.n341 VTAIL.n340 9.3005
R549 VTAIL.n339 VTAIL.n338 9.3005
R550 VTAIL.n286 VTAIL.n285 9.3005
R551 VTAIL.n333 VTAIL.n332 9.3005
R552 VTAIL.n331 VTAIL.n330 9.3005
R553 VTAIL.n290 VTAIL.n289 9.3005
R554 VTAIL.n236 VTAIL.n235 9.3005
R555 VTAIL.n238 VTAIL.n237 9.3005
R556 VTAIL.n229 VTAIL.n228 9.3005
R557 VTAIL.n244 VTAIL.n243 9.3005
R558 VTAIL.n246 VTAIL.n245 9.3005
R559 VTAIL.n224 VTAIL.n223 9.3005
R560 VTAIL.n252 VTAIL.n251 9.3005
R561 VTAIL.n254 VTAIL.n253 9.3005
R562 VTAIL.n277 VTAIL.n276 9.3005
R563 VTAIL.n212 VTAIL.n211 9.3005
R564 VTAIL.n271 VTAIL.n270 9.3005
R565 VTAIL.n269 VTAIL.n268 9.3005
R566 VTAIL.n216 VTAIL.n215 9.3005
R567 VTAIL.n263 VTAIL.n262 9.3005
R568 VTAIL.n261 VTAIL.n260 9.3005
R569 VTAIL.n220 VTAIL.n219 9.3005
R570 VTAIL.n518 VTAIL.n508 8.92171
R571 VTAIL.n552 VTAIL.n551 8.92171
R572 VTAIL.n28 VTAIL.n18 8.92171
R573 VTAIL.n62 VTAIL.n61 8.92171
R574 VTAIL.n98 VTAIL.n88 8.92171
R575 VTAIL.n132 VTAIL.n131 8.92171
R576 VTAIL.n168 VTAIL.n158 8.92171
R577 VTAIL.n202 VTAIL.n201 8.92171
R578 VTAIL.n482 VTAIL.n481 8.92171
R579 VTAIL.n449 VTAIL.n439 8.92171
R580 VTAIL.n412 VTAIL.n411 8.92171
R581 VTAIL.n379 VTAIL.n369 8.92171
R582 VTAIL.n342 VTAIL.n341 8.92171
R583 VTAIL.n309 VTAIL.n299 8.92171
R584 VTAIL.n272 VTAIL.n271 8.92171
R585 VTAIL.n239 VTAIL.n229 8.92171
R586 VTAIL.n517 VTAIL.n510 8.14595
R587 VTAIL.n555 VTAIL.n492 8.14595
R588 VTAIL.n27 VTAIL.n20 8.14595
R589 VTAIL.n65 VTAIL.n2 8.14595
R590 VTAIL.n97 VTAIL.n90 8.14595
R591 VTAIL.n135 VTAIL.n72 8.14595
R592 VTAIL.n167 VTAIL.n160 8.14595
R593 VTAIL.n205 VTAIL.n142 8.14595
R594 VTAIL.n485 VTAIL.n422 8.14595
R595 VTAIL.n448 VTAIL.n441 8.14595
R596 VTAIL.n415 VTAIL.n352 8.14595
R597 VTAIL.n378 VTAIL.n371 8.14595
R598 VTAIL.n345 VTAIL.n282 8.14595
R599 VTAIL.n308 VTAIL.n301 8.14595
R600 VTAIL.n275 VTAIL.n212 8.14595
R601 VTAIL.n238 VTAIL.n231 8.14595
R602 VTAIL.n514 VTAIL.n513 7.3702
R603 VTAIL.n556 VTAIL.n490 7.3702
R604 VTAIL.n24 VTAIL.n23 7.3702
R605 VTAIL.n66 VTAIL.n0 7.3702
R606 VTAIL.n94 VTAIL.n93 7.3702
R607 VTAIL.n136 VTAIL.n70 7.3702
R608 VTAIL.n164 VTAIL.n163 7.3702
R609 VTAIL.n206 VTAIL.n140 7.3702
R610 VTAIL.n486 VTAIL.n420 7.3702
R611 VTAIL.n445 VTAIL.n444 7.3702
R612 VTAIL.n416 VTAIL.n350 7.3702
R613 VTAIL.n375 VTAIL.n374 7.3702
R614 VTAIL.n346 VTAIL.n280 7.3702
R615 VTAIL.n305 VTAIL.n304 7.3702
R616 VTAIL.n276 VTAIL.n210 7.3702
R617 VTAIL.n235 VTAIL.n234 7.3702
R618 VTAIL.n558 VTAIL.n490 6.59444
R619 VTAIL.n68 VTAIL.n0 6.59444
R620 VTAIL.n138 VTAIL.n70 6.59444
R621 VTAIL.n208 VTAIL.n140 6.59444
R622 VTAIL.n488 VTAIL.n420 6.59444
R623 VTAIL.n418 VTAIL.n350 6.59444
R624 VTAIL.n348 VTAIL.n280 6.59444
R625 VTAIL.n278 VTAIL.n210 6.59444
R626 VTAIL.n514 VTAIL.n510 5.81868
R627 VTAIL.n556 VTAIL.n555 5.81868
R628 VTAIL.n24 VTAIL.n20 5.81868
R629 VTAIL.n66 VTAIL.n65 5.81868
R630 VTAIL.n94 VTAIL.n90 5.81868
R631 VTAIL.n136 VTAIL.n135 5.81868
R632 VTAIL.n164 VTAIL.n160 5.81868
R633 VTAIL.n206 VTAIL.n205 5.81868
R634 VTAIL.n486 VTAIL.n485 5.81868
R635 VTAIL.n445 VTAIL.n441 5.81868
R636 VTAIL.n416 VTAIL.n415 5.81868
R637 VTAIL.n375 VTAIL.n371 5.81868
R638 VTAIL.n346 VTAIL.n345 5.81868
R639 VTAIL.n305 VTAIL.n301 5.81868
R640 VTAIL.n276 VTAIL.n275 5.81868
R641 VTAIL.n235 VTAIL.n231 5.81868
R642 VTAIL.n518 VTAIL.n517 5.04292
R643 VTAIL.n552 VTAIL.n492 5.04292
R644 VTAIL.n28 VTAIL.n27 5.04292
R645 VTAIL.n62 VTAIL.n2 5.04292
R646 VTAIL.n98 VTAIL.n97 5.04292
R647 VTAIL.n132 VTAIL.n72 5.04292
R648 VTAIL.n168 VTAIL.n167 5.04292
R649 VTAIL.n202 VTAIL.n142 5.04292
R650 VTAIL.n482 VTAIL.n422 5.04292
R651 VTAIL.n449 VTAIL.n448 5.04292
R652 VTAIL.n412 VTAIL.n352 5.04292
R653 VTAIL.n379 VTAIL.n378 5.04292
R654 VTAIL.n342 VTAIL.n282 5.04292
R655 VTAIL.n309 VTAIL.n308 5.04292
R656 VTAIL.n272 VTAIL.n212 5.04292
R657 VTAIL.n239 VTAIL.n238 5.04292
R658 VTAIL.n521 VTAIL.n508 4.26717
R659 VTAIL.n551 VTAIL.n494 4.26717
R660 VTAIL.n31 VTAIL.n18 4.26717
R661 VTAIL.n61 VTAIL.n4 4.26717
R662 VTAIL.n101 VTAIL.n88 4.26717
R663 VTAIL.n131 VTAIL.n74 4.26717
R664 VTAIL.n171 VTAIL.n158 4.26717
R665 VTAIL.n201 VTAIL.n144 4.26717
R666 VTAIL.n481 VTAIL.n424 4.26717
R667 VTAIL.n452 VTAIL.n439 4.26717
R668 VTAIL.n411 VTAIL.n354 4.26717
R669 VTAIL.n382 VTAIL.n369 4.26717
R670 VTAIL.n341 VTAIL.n284 4.26717
R671 VTAIL.n312 VTAIL.n299 4.26717
R672 VTAIL.n271 VTAIL.n214 4.26717
R673 VTAIL.n242 VTAIL.n229 4.26717
R674 VTAIL.n522 VTAIL.n506 3.49141
R675 VTAIL.n548 VTAIL.n547 3.49141
R676 VTAIL.n32 VTAIL.n16 3.49141
R677 VTAIL.n58 VTAIL.n57 3.49141
R678 VTAIL.n102 VTAIL.n86 3.49141
R679 VTAIL.n128 VTAIL.n127 3.49141
R680 VTAIL.n172 VTAIL.n156 3.49141
R681 VTAIL.n198 VTAIL.n197 3.49141
R682 VTAIL.n478 VTAIL.n477 3.49141
R683 VTAIL.n453 VTAIL.n437 3.49141
R684 VTAIL.n408 VTAIL.n407 3.49141
R685 VTAIL.n383 VTAIL.n367 3.49141
R686 VTAIL.n338 VTAIL.n337 3.49141
R687 VTAIL.n313 VTAIL.n297 3.49141
R688 VTAIL.n268 VTAIL.n267 3.49141
R689 VTAIL.n243 VTAIL.n227 3.49141
R690 VTAIL.n349 VTAIL.n279 3.39705
R691 VTAIL.n489 VTAIL.n419 3.39705
R692 VTAIL.n209 VTAIL.n139 3.39705
R693 VTAIL.n526 VTAIL.n525 2.71565
R694 VTAIL.n544 VTAIL.n496 2.71565
R695 VTAIL.n36 VTAIL.n35 2.71565
R696 VTAIL.n54 VTAIL.n6 2.71565
R697 VTAIL.n106 VTAIL.n105 2.71565
R698 VTAIL.n124 VTAIL.n76 2.71565
R699 VTAIL.n176 VTAIL.n175 2.71565
R700 VTAIL.n194 VTAIL.n146 2.71565
R701 VTAIL.n474 VTAIL.n426 2.71565
R702 VTAIL.n457 VTAIL.n456 2.71565
R703 VTAIL.n404 VTAIL.n356 2.71565
R704 VTAIL.n387 VTAIL.n386 2.71565
R705 VTAIL.n334 VTAIL.n286 2.71565
R706 VTAIL.n317 VTAIL.n316 2.71565
R707 VTAIL.n264 VTAIL.n216 2.71565
R708 VTAIL.n247 VTAIL.n246 2.71565
R709 VTAIL.n515 VTAIL.n511 2.41282
R710 VTAIL.n25 VTAIL.n21 2.41282
R711 VTAIL.n95 VTAIL.n91 2.41282
R712 VTAIL.n165 VTAIL.n161 2.41282
R713 VTAIL.n446 VTAIL.n442 2.41282
R714 VTAIL.n376 VTAIL.n372 2.41282
R715 VTAIL.n306 VTAIL.n302 2.41282
R716 VTAIL.n236 VTAIL.n232 2.41282
R717 VTAIL.n530 VTAIL.n504 1.93989
R718 VTAIL.n543 VTAIL.n498 1.93989
R719 VTAIL.n40 VTAIL.n14 1.93989
R720 VTAIL.n53 VTAIL.n8 1.93989
R721 VTAIL.n110 VTAIL.n84 1.93989
R722 VTAIL.n123 VTAIL.n78 1.93989
R723 VTAIL.n180 VTAIL.n154 1.93989
R724 VTAIL.n193 VTAIL.n148 1.93989
R725 VTAIL.n473 VTAIL.n428 1.93989
R726 VTAIL.n460 VTAIL.n434 1.93989
R727 VTAIL.n403 VTAIL.n358 1.93989
R728 VTAIL.n390 VTAIL.n364 1.93989
R729 VTAIL.n333 VTAIL.n288 1.93989
R730 VTAIL.n320 VTAIL.n294 1.93989
R731 VTAIL.n263 VTAIL.n218 1.93989
R732 VTAIL.n250 VTAIL.n224 1.93989
R733 VTAIL VTAIL.n69 1.75697
R734 VTAIL VTAIL.n559 1.64059
R735 VTAIL.n531 VTAIL.n502 1.16414
R736 VTAIL.n540 VTAIL.n539 1.16414
R737 VTAIL.n41 VTAIL.n12 1.16414
R738 VTAIL.n50 VTAIL.n49 1.16414
R739 VTAIL.n111 VTAIL.n82 1.16414
R740 VTAIL.n120 VTAIL.n119 1.16414
R741 VTAIL.n181 VTAIL.n152 1.16414
R742 VTAIL.n190 VTAIL.n189 1.16414
R743 VTAIL.n470 VTAIL.n469 1.16414
R744 VTAIL.n461 VTAIL.n432 1.16414
R745 VTAIL.n400 VTAIL.n399 1.16414
R746 VTAIL.n391 VTAIL.n362 1.16414
R747 VTAIL.n330 VTAIL.n329 1.16414
R748 VTAIL.n321 VTAIL.n292 1.16414
R749 VTAIL.n260 VTAIL.n259 1.16414
R750 VTAIL.n251 VTAIL.n222 1.16414
R751 VTAIL.n419 VTAIL.n349 0.470328
R752 VTAIL.n139 VTAIL.n69 0.470328
R753 VTAIL.n535 VTAIL.n534 0.388379
R754 VTAIL.n536 VTAIL.n500 0.388379
R755 VTAIL.n45 VTAIL.n44 0.388379
R756 VTAIL.n46 VTAIL.n10 0.388379
R757 VTAIL.n115 VTAIL.n114 0.388379
R758 VTAIL.n116 VTAIL.n80 0.388379
R759 VTAIL.n185 VTAIL.n184 0.388379
R760 VTAIL.n186 VTAIL.n150 0.388379
R761 VTAIL.n466 VTAIL.n430 0.388379
R762 VTAIL.n465 VTAIL.n464 0.388379
R763 VTAIL.n396 VTAIL.n360 0.388379
R764 VTAIL.n395 VTAIL.n394 0.388379
R765 VTAIL.n326 VTAIL.n290 0.388379
R766 VTAIL.n325 VTAIL.n324 0.388379
R767 VTAIL.n256 VTAIL.n220 0.388379
R768 VTAIL.n255 VTAIL.n254 0.388379
R769 VTAIL.n516 VTAIL.n515 0.155672
R770 VTAIL.n516 VTAIL.n507 0.155672
R771 VTAIL.n523 VTAIL.n507 0.155672
R772 VTAIL.n524 VTAIL.n523 0.155672
R773 VTAIL.n524 VTAIL.n503 0.155672
R774 VTAIL.n532 VTAIL.n503 0.155672
R775 VTAIL.n533 VTAIL.n532 0.155672
R776 VTAIL.n533 VTAIL.n499 0.155672
R777 VTAIL.n541 VTAIL.n499 0.155672
R778 VTAIL.n542 VTAIL.n541 0.155672
R779 VTAIL.n542 VTAIL.n495 0.155672
R780 VTAIL.n549 VTAIL.n495 0.155672
R781 VTAIL.n550 VTAIL.n549 0.155672
R782 VTAIL.n550 VTAIL.n491 0.155672
R783 VTAIL.n557 VTAIL.n491 0.155672
R784 VTAIL.n26 VTAIL.n25 0.155672
R785 VTAIL.n26 VTAIL.n17 0.155672
R786 VTAIL.n33 VTAIL.n17 0.155672
R787 VTAIL.n34 VTAIL.n33 0.155672
R788 VTAIL.n34 VTAIL.n13 0.155672
R789 VTAIL.n42 VTAIL.n13 0.155672
R790 VTAIL.n43 VTAIL.n42 0.155672
R791 VTAIL.n43 VTAIL.n9 0.155672
R792 VTAIL.n51 VTAIL.n9 0.155672
R793 VTAIL.n52 VTAIL.n51 0.155672
R794 VTAIL.n52 VTAIL.n5 0.155672
R795 VTAIL.n59 VTAIL.n5 0.155672
R796 VTAIL.n60 VTAIL.n59 0.155672
R797 VTAIL.n60 VTAIL.n1 0.155672
R798 VTAIL.n67 VTAIL.n1 0.155672
R799 VTAIL.n96 VTAIL.n95 0.155672
R800 VTAIL.n96 VTAIL.n87 0.155672
R801 VTAIL.n103 VTAIL.n87 0.155672
R802 VTAIL.n104 VTAIL.n103 0.155672
R803 VTAIL.n104 VTAIL.n83 0.155672
R804 VTAIL.n112 VTAIL.n83 0.155672
R805 VTAIL.n113 VTAIL.n112 0.155672
R806 VTAIL.n113 VTAIL.n79 0.155672
R807 VTAIL.n121 VTAIL.n79 0.155672
R808 VTAIL.n122 VTAIL.n121 0.155672
R809 VTAIL.n122 VTAIL.n75 0.155672
R810 VTAIL.n129 VTAIL.n75 0.155672
R811 VTAIL.n130 VTAIL.n129 0.155672
R812 VTAIL.n130 VTAIL.n71 0.155672
R813 VTAIL.n137 VTAIL.n71 0.155672
R814 VTAIL.n166 VTAIL.n165 0.155672
R815 VTAIL.n166 VTAIL.n157 0.155672
R816 VTAIL.n173 VTAIL.n157 0.155672
R817 VTAIL.n174 VTAIL.n173 0.155672
R818 VTAIL.n174 VTAIL.n153 0.155672
R819 VTAIL.n182 VTAIL.n153 0.155672
R820 VTAIL.n183 VTAIL.n182 0.155672
R821 VTAIL.n183 VTAIL.n149 0.155672
R822 VTAIL.n191 VTAIL.n149 0.155672
R823 VTAIL.n192 VTAIL.n191 0.155672
R824 VTAIL.n192 VTAIL.n145 0.155672
R825 VTAIL.n199 VTAIL.n145 0.155672
R826 VTAIL.n200 VTAIL.n199 0.155672
R827 VTAIL.n200 VTAIL.n141 0.155672
R828 VTAIL.n207 VTAIL.n141 0.155672
R829 VTAIL.n487 VTAIL.n421 0.155672
R830 VTAIL.n480 VTAIL.n421 0.155672
R831 VTAIL.n480 VTAIL.n479 0.155672
R832 VTAIL.n479 VTAIL.n425 0.155672
R833 VTAIL.n472 VTAIL.n425 0.155672
R834 VTAIL.n472 VTAIL.n471 0.155672
R835 VTAIL.n471 VTAIL.n429 0.155672
R836 VTAIL.n463 VTAIL.n429 0.155672
R837 VTAIL.n463 VTAIL.n462 0.155672
R838 VTAIL.n462 VTAIL.n433 0.155672
R839 VTAIL.n455 VTAIL.n433 0.155672
R840 VTAIL.n455 VTAIL.n454 0.155672
R841 VTAIL.n454 VTAIL.n438 0.155672
R842 VTAIL.n447 VTAIL.n438 0.155672
R843 VTAIL.n447 VTAIL.n446 0.155672
R844 VTAIL.n417 VTAIL.n351 0.155672
R845 VTAIL.n410 VTAIL.n351 0.155672
R846 VTAIL.n410 VTAIL.n409 0.155672
R847 VTAIL.n409 VTAIL.n355 0.155672
R848 VTAIL.n402 VTAIL.n355 0.155672
R849 VTAIL.n402 VTAIL.n401 0.155672
R850 VTAIL.n401 VTAIL.n359 0.155672
R851 VTAIL.n393 VTAIL.n359 0.155672
R852 VTAIL.n393 VTAIL.n392 0.155672
R853 VTAIL.n392 VTAIL.n363 0.155672
R854 VTAIL.n385 VTAIL.n363 0.155672
R855 VTAIL.n385 VTAIL.n384 0.155672
R856 VTAIL.n384 VTAIL.n368 0.155672
R857 VTAIL.n377 VTAIL.n368 0.155672
R858 VTAIL.n377 VTAIL.n376 0.155672
R859 VTAIL.n347 VTAIL.n281 0.155672
R860 VTAIL.n340 VTAIL.n281 0.155672
R861 VTAIL.n340 VTAIL.n339 0.155672
R862 VTAIL.n339 VTAIL.n285 0.155672
R863 VTAIL.n332 VTAIL.n285 0.155672
R864 VTAIL.n332 VTAIL.n331 0.155672
R865 VTAIL.n331 VTAIL.n289 0.155672
R866 VTAIL.n323 VTAIL.n289 0.155672
R867 VTAIL.n323 VTAIL.n322 0.155672
R868 VTAIL.n322 VTAIL.n293 0.155672
R869 VTAIL.n315 VTAIL.n293 0.155672
R870 VTAIL.n315 VTAIL.n314 0.155672
R871 VTAIL.n314 VTAIL.n298 0.155672
R872 VTAIL.n307 VTAIL.n298 0.155672
R873 VTAIL.n307 VTAIL.n306 0.155672
R874 VTAIL.n277 VTAIL.n211 0.155672
R875 VTAIL.n270 VTAIL.n211 0.155672
R876 VTAIL.n270 VTAIL.n269 0.155672
R877 VTAIL.n269 VTAIL.n215 0.155672
R878 VTAIL.n262 VTAIL.n215 0.155672
R879 VTAIL.n262 VTAIL.n261 0.155672
R880 VTAIL.n261 VTAIL.n219 0.155672
R881 VTAIL.n253 VTAIL.n219 0.155672
R882 VTAIL.n253 VTAIL.n252 0.155672
R883 VTAIL.n252 VTAIL.n223 0.155672
R884 VTAIL.n245 VTAIL.n223 0.155672
R885 VTAIL.n245 VTAIL.n244 0.155672
R886 VTAIL.n244 VTAIL.n228 0.155672
R887 VTAIL.n237 VTAIL.n228 0.155672
R888 VTAIL.n237 VTAIL.n236 0.155672
R889 B.n535 B.n76 585
R890 B.n537 B.n536 585
R891 B.n538 B.n75 585
R892 B.n540 B.n539 585
R893 B.n541 B.n74 585
R894 B.n543 B.n542 585
R895 B.n544 B.n73 585
R896 B.n546 B.n545 585
R897 B.n547 B.n72 585
R898 B.n549 B.n548 585
R899 B.n550 B.n71 585
R900 B.n552 B.n551 585
R901 B.n553 B.n70 585
R902 B.n555 B.n554 585
R903 B.n556 B.n69 585
R904 B.n558 B.n557 585
R905 B.n559 B.n68 585
R906 B.n561 B.n560 585
R907 B.n562 B.n67 585
R908 B.n564 B.n563 585
R909 B.n565 B.n66 585
R910 B.n567 B.n566 585
R911 B.n568 B.n65 585
R912 B.n570 B.n569 585
R913 B.n571 B.n64 585
R914 B.n573 B.n572 585
R915 B.n574 B.n63 585
R916 B.n576 B.n575 585
R917 B.n577 B.n62 585
R918 B.n579 B.n578 585
R919 B.n580 B.n61 585
R920 B.n582 B.n581 585
R921 B.n583 B.n60 585
R922 B.n585 B.n584 585
R923 B.n586 B.n59 585
R924 B.n588 B.n587 585
R925 B.n589 B.n58 585
R926 B.n591 B.n590 585
R927 B.n592 B.n57 585
R928 B.n594 B.n593 585
R929 B.n595 B.n56 585
R930 B.n597 B.n596 585
R931 B.n598 B.n55 585
R932 B.n600 B.n599 585
R933 B.n602 B.n601 585
R934 B.n603 B.n51 585
R935 B.n605 B.n604 585
R936 B.n606 B.n50 585
R937 B.n608 B.n607 585
R938 B.n609 B.n49 585
R939 B.n611 B.n610 585
R940 B.n612 B.n48 585
R941 B.n614 B.n613 585
R942 B.n616 B.n45 585
R943 B.n618 B.n617 585
R944 B.n619 B.n44 585
R945 B.n621 B.n620 585
R946 B.n622 B.n43 585
R947 B.n624 B.n623 585
R948 B.n625 B.n42 585
R949 B.n627 B.n626 585
R950 B.n628 B.n41 585
R951 B.n630 B.n629 585
R952 B.n631 B.n40 585
R953 B.n633 B.n632 585
R954 B.n634 B.n39 585
R955 B.n636 B.n635 585
R956 B.n637 B.n38 585
R957 B.n639 B.n638 585
R958 B.n640 B.n37 585
R959 B.n642 B.n641 585
R960 B.n643 B.n36 585
R961 B.n645 B.n644 585
R962 B.n646 B.n35 585
R963 B.n648 B.n647 585
R964 B.n649 B.n34 585
R965 B.n651 B.n650 585
R966 B.n652 B.n33 585
R967 B.n654 B.n653 585
R968 B.n655 B.n32 585
R969 B.n657 B.n656 585
R970 B.n658 B.n31 585
R971 B.n660 B.n659 585
R972 B.n661 B.n30 585
R973 B.n663 B.n662 585
R974 B.n664 B.n29 585
R975 B.n666 B.n665 585
R976 B.n667 B.n28 585
R977 B.n669 B.n668 585
R978 B.n670 B.n27 585
R979 B.n672 B.n671 585
R980 B.n673 B.n26 585
R981 B.n675 B.n674 585
R982 B.n676 B.n25 585
R983 B.n678 B.n677 585
R984 B.n679 B.n24 585
R985 B.n681 B.n680 585
R986 B.n534 B.n533 585
R987 B.n532 B.n77 585
R988 B.n531 B.n530 585
R989 B.n529 B.n78 585
R990 B.n528 B.n527 585
R991 B.n526 B.n79 585
R992 B.n525 B.n524 585
R993 B.n523 B.n80 585
R994 B.n522 B.n521 585
R995 B.n520 B.n81 585
R996 B.n519 B.n518 585
R997 B.n517 B.n82 585
R998 B.n516 B.n515 585
R999 B.n514 B.n83 585
R1000 B.n513 B.n512 585
R1001 B.n511 B.n84 585
R1002 B.n510 B.n509 585
R1003 B.n508 B.n85 585
R1004 B.n507 B.n506 585
R1005 B.n505 B.n86 585
R1006 B.n504 B.n503 585
R1007 B.n502 B.n87 585
R1008 B.n501 B.n500 585
R1009 B.n499 B.n88 585
R1010 B.n498 B.n497 585
R1011 B.n496 B.n89 585
R1012 B.n495 B.n494 585
R1013 B.n493 B.n90 585
R1014 B.n492 B.n491 585
R1015 B.n490 B.n91 585
R1016 B.n489 B.n488 585
R1017 B.n487 B.n92 585
R1018 B.n486 B.n485 585
R1019 B.n484 B.n93 585
R1020 B.n483 B.n482 585
R1021 B.n481 B.n94 585
R1022 B.n480 B.n479 585
R1023 B.n478 B.n95 585
R1024 B.n477 B.n476 585
R1025 B.n475 B.n96 585
R1026 B.n474 B.n473 585
R1027 B.n472 B.n97 585
R1028 B.n471 B.n470 585
R1029 B.n469 B.n98 585
R1030 B.n468 B.n467 585
R1031 B.n466 B.n99 585
R1032 B.n465 B.n464 585
R1033 B.n463 B.n100 585
R1034 B.n462 B.n461 585
R1035 B.n460 B.n101 585
R1036 B.n459 B.n458 585
R1037 B.n457 B.n102 585
R1038 B.n456 B.n455 585
R1039 B.n454 B.n103 585
R1040 B.n453 B.n452 585
R1041 B.n451 B.n104 585
R1042 B.n450 B.n449 585
R1043 B.n448 B.n105 585
R1044 B.n447 B.n446 585
R1045 B.n445 B.n106 585
R1046 B.n444 B.n443 585
R1047 B.n442 B.n107 585
R1048 B.n441 B.n440 585
R1049 B.n439 B.n108 585
R1050 B.n438 B.n437 585
R1051 B.n436 B.n109 585
R1052 B.n435 B.n434 585
R1053 B.n433 B.n110 585
R1054 B.n432 B.n431 585
R1055 B.n430 B.n111 585
R1056 B.n429 B.n428 585
R1057 B.n427 B.n112 585
R1058 B.n426 B.n425 585
R1059 B.n424 B.n113 585
R1060 B.n423 B.n422 585
R1061 B.n421 B.n114 585
R1062 B.n420 B.n419 585
R1063 B.n418 B.n115 585
R1064 B.n417 B.n416 585
R1065 B.n415 B.n116 585
R1066 B.n414 B.n413 585
R1067 B.n412 B.n117 585
R1068 B.n411 B.n410 585
R1069 B.n409 B.n118 585
R1070 B.n408 B.n407 585
R1071 B.n406 B.n119 585
R1072 B.n405 B.n404 585
R1073 B.n258 B.n257 585
R1074 B.n259 B.n172 585
R1075 B.n261 B.n260 585
R1076 B.n262 B.n171 585
R1077 B.n264 B.n263 585
R1078 B.n265 B.n170 585
R1079 B.n267 B.n266 585
R1080 B.n268 B.n169 585
R1081 B.n270 B.n269 585
R1082 B.n271 B.n168 585
R1083 B.n273 B.n272 585
R1084 B.n274 B.n167 585
R1085 B.n276 B.n275 585
R1086 B.n277 B.n166 585
R1087 B.n279 B.n278 585
R1088 B.n280 B.n165 585
R1089 B.n282 B.n281 585
R1090 B.n283 B.n164 585
R1091 B.n285 B.n284 585
R1092 B.n286 B.n163 585
R1093 B.n288 B.n287 585
R1094 B.n289 B.n162 585
R1095 B.n291 B.n290 585
R1096 B.n292 B.n161 585
R1097 B.n294 B.n293 585
R1098 B.n295 B.n160 585
R1099 B.n297 B.n296 585
R1100 B.n298 B.n159 585
R1101 B.n300 B.n299 585
R1102 B.n301 B.n158 585
R1103 B.n303 B.n302 585
R1104 B.n304 B.n157 585
R1105 B.n306 B.n305 585
R1106 B.n307 B.n156 585
R1107 B.n309 B.n308 585
R1108 B.n310 B.n155 585
R1109 B.n312 B.n311 585
R1110 B.n313 B.n154 585
R1111 B.n315 B.n314 585
R1112 B.n316 B.n153 585
R1113 B.n318 B.n317 585
R1114 B.n319 B.n152 585
R1115 B.n321 B.n320 585
R1116 B.n322 B.n149 585
R1117 B.n325 B.n324 585
R1118 B.n326 B.n148 585
R1119 B.n328 B.n327 585
R1120 B.n329 B.n147 585
R1121 B.n331 B.n330 585
R1122 B.n332 B.n146 585
R1123 B.n334 B.n333 585
R1124 B.n335 B.n145 585
R1125 B.n337 B.n336 585
R1126 B.n339 B.n338 585
R1127 B.n340 B.n141 585
R1128 B.n342 B.n341 585
R1129 B.n343 B.n140 585
R1130 B.n345 B.n344 585
R1131 B.n346 B.n139 585
R1132 B.n348 B.n347 585
R1133 B.n349 B.n138 585
R1134 B.n351 B.n350 585
R1135 B.n352 B.n137 585
R1136 B.n354 B.n353 585
R1137 B.n355 B.n136 585
R1138 B.n357 B.n356 585
R1139 B.n358 B.n135 585
R1140 B.n360 B.n359 585
R1141 B.n361 B.n134 585
R1142 B.n363 B.n362 585
R1143 B.n364 B.n133 585
R1144 B.n366 B.n365 585
R1145 B.n367 B.n132 585
R1146 B.n369 B.n368 585
R1147 B.n370 B.n131 585
R1148 B.n372 B.n371 585
R1149 B.n373 B.n130 585
R1150 B.n375 B.n374 585
R1151 B.n376 B.n129 585
R1152 B.n378 B.n377 585
R1153 B.n379 B.n128 585
R1154 B.n381 B.n380 585
R1155 B.n382 B.n127 585
R1156 B.n384 B.n383 585
R1157 B.n385 B.n126 585
R1158 B.n387 B.n386 585
R1159 B.n388 B.n125 585
R1160 B.n390 B.n389 585
R1161 B.n391 B.n124 585
R1162 B.n393 B.n392 585
R1163 B.n394 B.n123 585
R1164 B.n396 B.n395 585
R1165 B.n397 B.n122 585
R1166 B.n399 B.n398 585
R1167 B.n400 B.n121 585
R1168 B.n402 B.n401 585
R1169 B.n403 B.n120 585
R1170 B.n256 B.n173 585
R1171 B.n255 B.n254 585
R1172 B.n253 B.n174 585
R1173 B.n252 B.n251 585
R1174 B.n250 B.n175 585
R1175 B.n249 B.n248 585
R1176 B.n247 B.n176 585
R1177 B.n246 B.n245 585
R1178 B.n244 B.n177 585
R1179 B.n243 B.n242 585
R1180 B.n241 B.n178 585
R1181 B.n240 B.n239 585
R1182 B.n238 B.n179 585
R1183 B.n237 B.n236 585
R1184 B.n235 B.n180 585
R1185 B.n234 B.n233 585
R1186 B.n232 B.n181 585
R1187 B.n231 B.n230 585
R1188 B.n229 B.n182 585
R1189 B.n228 B.n227 585
R1190 B.n226 B.n183 585
R1191 B.n225 B.n224 585
R1192 B.n223 B.n184 585
R1193 B.n222 B.n221 585
R1194 B.n220 B.n185 585
R1195 B.n219 B.n218 585
R1196 B.n217 B.n186 585
R1197 B.n216 B.n215 585
R1198 B.n214 B.n187 585
R1199 B.n213 B.n212 585
R1200 B.n211 B.n188 585
R1201 B.n210 B.n209 585
R1202 B.n208 B.n189 585
R1203 B.n207 B.n206 585
R1204 B.n205 B.n190 585
R1205 B.n204 B.n203 585
R1206 B.n202 B.n191 585
R1207 B.n201 B.n200 585
R1208 B.n199 B.n192 585
R1209 B.n198 B.n197 585
R1210 B.n196 B.n193 585
R1211 B.n195 B.n194 585
R1212 B.n2 B.n0 585
R1213 B.n745 B.n1 585
R1214 B.n744 B.n743 585
R1215 B.n742 B.n3 585
R1216 B.n741 B.n740 585
R1217 B.n739 B.n4 585
R1218 B.n738 B.n737 585
R1219 B.n736 B.n5 585
R1220 B.n735 B.n734 585
R1221 B.n733 B.n6 585
R1222 B.n732 B.n731 585
R1223 B.n730 B.n7 585
R1224 B.n729 B.n728 585
R1225 B.n727 B.n8 585
R1226 B.n726 B.n725 585
R1227 B.n724 B.n9 585
R1228 B.n723 B.n722 585
R1229 B.n721 B.n10 585
R1230 B.n720 B.n719 585
R1231 B.n718 B.n11 585
R1232 B.n717 B.n716 585
R1233 B.n715 B.n12 585
R1234 B.n714 B.n713 585
R1235 B.n712 B.n13 585
R1236 B.n711 B.n710 585
R1237 B.n709 B.n14 585
R1238 B.n708 B.n707 585
R1239 B.n706 B.n15 585
R1240 B.n705 B.n704 585
R1241 B.n703 B.n16 585
R1242 B.n702 B.n701 585
R1243 B.n700 B.n17 585
R1244 B.n699 B.n698 585
R1245 B.n697 B.n18 585
R1246 B.n696 B.n695 585
R1247 B.n694 B.n19 585
R1248 B.n693 B.n692 585
R1249 B.n691 B.n20 585
R1250 B.n690 B.n689 585
R1251 B.n688 B.n21 585
R1252 B.n687 B.n686 585
R1253 B.n685 B.n22 585
R1254 B.n684 B.n683 585
R1255 B.n682 B.n23 585
R1256 B.n747 B.n746 585
R1257 B.n258 B.n173 487.695
R1258 B.n680 B.n23 487.695
R1259 B.n404 B.n403 487.695
R1260 B.n535 B.n534 487.695
R1261 B.n142 B.t2 465.159
R1262 B.n52 B.t10 465.159
R1263 B.n150 B.t8 465.159
R1264 B.n46 B.t4 465.159
R1265 B.n143 B.t1 388.747
R1266 B.n53 B.t11 388.747
R1267 B.n151 B.t7 388.747
R1268 B.n47 B.t5 388.747
R1269 B.n142 B.t0 294.175
R1270 B.n150 B.t6 294.175
R1271 B.n46 B.t3 294.175
R1272 B.n52 B.t9 294.175
R1273 B.n254 B.n173 163.367
R1274 B.n254 B.n253 163.367
R1275 B.n253 B.n252 163.367
R1276 B.n252 B.n175 163.367
R1277 B.n248 B.n175 163.367
R1278 B.n248 B.n247 163.367
R1279 B.n247 B.n246 163.367
R1280 B.n246 B.n177 163.367
R1281 B.n242 B.n177 163.367
R1282 B.n242 B.n241 163.367
R1283 B.n241 B.n240 163.367
R1284 B.n240 B.n179 163.367
R1285 B.n236 B.n179 163.367
R1286 B.n236 B.n235 163.367
R1287 B.n235 B.n234 163.367
R1288 B.n234 B.n181 163.367
R1289 B.n230 B.n181 163.367
R1290 B.n230 B.n229 163.367
R1291 B.n229 B.n228 163.367
R1292 B.n228 B.n183 163.367
R1293 B.n224 B.n183 163.367
R1294 B.n224 B.n223 163.367
R1295 B.n223 B.n222 163.367
R1296 B.n222 B.n185 163.367
R1297 B.n218 B.n185 163.367
R1298 B.n218 B.n217 163.367
R1299 B.n217 B.n216 163.367
R1300 B.n216 B.n187 163.367
R1301 B.n212 B.n187 163.367
R1302 B.n212 B.n211 163.367
R1303 B.n211 B.n210 163.367
R1304 B.n210 B.n189 163.367
R1305 B.n206 B.n189 163.367
R1306 B.n206 B.n205 163.367
R1307 B.n205 B.n204 163.367
R1308 B.n204 B.n191 163.367
R1309 B.n200 B.n191 163.367
R1310 B.n200 B.n199 163.367
R1311 B.n199 B.n198 163.367
R1312 B.n198 B.n193 163.367
R1313 B.n194 B.n193 163.367
R1314 B.n194 B.n2 163.367
R1315 B.n746 B.n2 163.367
R1316 B.n746 B.n745 163.367
R1317 B.n745 B.n744 163.367
R1318 B.n744 B.n3 163.367
R1319 B.n740 B.n3 163.367
R1320 B.n740 B.n739 163.367
R1321 B.n739 B.n738 163.367
R1322 B.n738 B.n5 163.367
R1323 B.n734 B.n5 163.367
R1324 B.n734 B.n733 163.367
R1325 B.n733 B.n732 163.367
R1326 B.n732 B.n7 163.367
R1327 B.n728 B.n7 163.367
R1328 B.n728 B.n727 163.367
R1329 B.n727 B.n726 163.367
R1330 B.n726 B.n9 163.367
R1331 B.n722 B.n9 163.367
R1332 B.n722 B.n721 163.367
R1333 B.n721 B.n720 163.367
R1334 B.n720 B.n11 163.367
R1335 B.n716 B.n11 163.367
R1336 B.n716 B.n715 163.367
R1337 B.n715 B.n714 163.367
R1338 B.n714 B.n13 163.367
R1339 B.n710 B.n13 163.367
R1340 B.n710 B.n709 163.367
R1341 B.n709 B.n708 163.367
R1342 B.n708 B.n15 163.367
R1343 B.n704 B.n15 163.367
R1344 B.n704 B.n703 163.367
R1345 B.n703 B.n702 163.367
R1346 B.n702 B.n17 163.367
R1347 B.n698 B.n17 163.367
R1348 B.n698 B.n697 163.367
R1349 B.n697 B.n696 163.367
R1350 B.n696 B.n19 163.367
R1351 B.n692 B.n19 163.367
R1352 B.n692 B.n691 163.367
R1353 B.n691 B.n690 163.367
R1354 B.n690 B.n21 163.367
R1355 B.n686 B.n21 163.367
R1356 B.n686 B.n685 163.367
R1357 B.n685 B.n684 163.367
R1358 B.n684 B.n23 163.367
R1359 B.n259 B.n258 163.367
R1360 B.n260 B.n259 163.367
R1361 B.n260 B.n171 163.367
R1362 B.n264 B.n171 163.367
R1363 B.n265 B.n264 163.367
R1364 B.n266 B.n265 163.367
R1365 B.n266 B.n169 163.367
R1366 B.n270 B.n169 163.367
R1367 B.n271 B.n270 163.367
R1368 B.n272 B.n271 163.367
R1369 B.n272 B.n167 163.367
R1370 B.n276 B.n167 163.367
R1371 B.n277 B.n276 163.367
R1372 B.n278 B.n277 163.367
R1373 B.n278 B.n165 163.367
R1374 B.n282 B.n165 163.367
R1375 B.n283 B.n282 163.367
R1376 B.n284 B.n283 163.367
R1377 B.n284 B.n163 163.367
R1378 B.n288 B.n163 163.367
R1379 B.n289 B.n288 163.367
R1380 B.n290 B.n289 163.367
R1381 B.n290 B.n161 163.367
R1382 B.n294 B.n161 163.367
R1383 B.n295 B.n294 163.367
R1384 B.n296 B.n295 163.367
R1385 B.n296 B.n159 163.367
R1386 B.n300 B.n159 163.367
R1387 B.n301 B.n300 163.367
R1388 B.n302 B.n301 163.367
R1389 B.n302 B.n157 163.367
R1390 B.n306 B.n157 163.367
R1391 B.n307 B.n306 163.367
R1392 B.n308 B.n307 163.367
R1393 B.n308 B.n155 163.367
R1394 B.n312 B.n155 163.367
R1395 B.n313 B.n312 163.367
R1396 B.n314 B.n313 163.367
R1397 B.n314 B.n153 163.367
R1398 B.n318 B.n153 163.367
R1399 B.n319 B.n318 163.367
R1400 B.n320 B.n319 163.367
R1401 B.n320 B.n149 163.367
R1402 B.n325 B.n149 163.367
R1403 B.n326 B.n325 163.367
R1404 B.n327 B.n326 163.367
R1405 B.n327 B.n147 163.367
R1406 B.n331 B.n147 163.367
R1407 B.n332 B.n331 163.367
R1408 B.n333 B.n332 163.367
R1409 B.n333 B.n145 163.367
R1410 B.n337 B.n145 163.367
R1411 B.n338 B.n337 163.367
R1412 B.n338 B.n141 163.367
R1413 B.n342 B.n141 163.367
R1414 B.n343 B.n342 163.367
R1415 B.n344 B.n343 163.367
R1416 B.n344 B.n139 163.367
R1417 B.n348 B.n139 163.367
R1418 B.n349 B.n348 163.367
R1419 B.n350 B.n349 163.367
R1420 B.n350 B.n137 163.367
R1421 B.n354 B.n137 163.367
R1422 B.n355 B.n354 163.367
R1423 B.n356 B.n355 163.367
R1424 B.n356 B.n135 163.367
R1425 B.n360 B.n135 163.367
R1426 B.n361 B.n360 163.367
R1427 B.n362 B.n361 163.367
R1428 B.n362 B.n133 163.367
R1429 B.n366 B.n133 163.367
R1430 B.n367 B.n366 163.367
R1431 B.n368 B.n367 163.367
R1432 B.n368 B.n131 163.367
R1433 B.n372 B.n131 163.367
R1434 B.n373 B.n372 163.367
R1435 B.n374 B.n373 163.367
R1436 B.n374 B.n129 163.367
R1437 B.n378 B.n129 163.367
R1438 B.n379 B.n378 163.367
R1439 B.n380 B.n379 163.367
R1440 B.n380 B.n127 163.367
R1441 B.n384 B.n127 163.367
R1442 B.n385 B.n384 163.367
R1443 B.n386 B.n385 163.367
R1444 B.n386 B.n125 163.367
R1445 B.n390 B.n125 163.367
R1446 B.n391 B.n390 163.367
R1447 B.n392 B.n391 163.367
R1448 B.n392 B.n123 163.367
R1449 B.n396 B.n123 163.367
R1450 B.n397 B.n396 163.367
R1451 B.n398 B.n397 163.367
R1452 B.n398 B.n121 163.367
R1453 B.n402 B.n121 163.367
R1454 B.n403 B.n402 163.367
R1455 B.n404 B.n119 163.367
R1456 B.n408 B.n119 163.367
R1457 B.n409 B.n408 163.367
R1458 B.n410 B.n409 163.367
R1459 B.n410 B.n117 163.367
R1460 B.n414 B.n117 163.367
R1461 B.n415 B.n414 163.367
R1462 B.n416 B.n415 163.367
R1463 B.n416 B.n115 163.367
R1464 B.n420 B.n115 163.367
R1465 B.n421 B.n420 163.367
R1466 B.n422 B.n421 163.367
R1467 B.n422 B.n113 163.367
R1468 B.n426 B.n113 163.367
R1469 B.n427 B.n426 163.367
R1470 B.n428 B.n427 163.367
R1471 B.n428 B.n111 163.367
R1472 B.n432 B.n111 163.367
R1473 B.n433 B.n432 163.367
R1474 B.n434 B.n433 163.367
R1475 B.n434 B.n109 163.367
R1476 B.n438 B.n109 163.367
R1477 B.n439 B.n438 163.367
R1478 B.n440 B.n439 163.367
R1479 B.n440 B.n107 163.367
R1480 B.n444 B.n107 163.367
R1481 B.n445 B.n444 163.367
R1482 B.n446 B.n445 163.367
R1483 B.n446 B.n105 163.367
R1484 B.n450 B.n105 163.367
R1485 B.n451 B.n450 163.367
R1486 B.n452 B.n451 163.367
R1487 B.n452 B.n103 163.367
R1488 B.n456 B.n103 163.367
R1489 B.n457 B.n456 163.367
R1490 B.n458 B.n457 163.367
R1491 B.n458 B.n101 163.367
R1492 B.n462 B.n101 163.367
R1493 B.n463 B.n462 163.367
R1494 B.n464 B.n463 163.367
R1495 B.n464 B.n99 163.367
R1496 B.n468 B.n99 163.367
R1497 B.n469 B.n468 163.367
R1498 B.n470 B.n469 163.367
R1499 B.n470 B.n97 163.367
R1500 B.n474 B.n97 163.367
R1501 B.n475 B.n474 163.367
R1502 B.n476 B.n475 163.367
R1503 B.n476 B.n95 163.367
R1504 B.n480 B.n95 163.367
R1505 B.n481 B.n480 163.367
R1506 B.n482 B.n481 163.367
R1507 B.n482 B.n93 163.367
R1508 B.n486 B.n93 163.367
R1509 B.n487 B.n486 163.367
R1510 B.n488 B.n487 163.367
R1511 B.n488 B.n91 163.367
R1512 B.n492 B.n91 163.367
R1513 B.n493 B.n492 163.367
R1514 B.n494 B.n493 163.367
R1515 B.n494 B.n89 163.367
R1516 B.n498 B.n89 163.367
R1517 B.n499 B.n498 163.367
R1518 B.n500 B.n499 163.367
R1519 B.n500 B.n87 163.367
R1520 B.n504 B.n87 163.367
R1521 B.n505 B.n504 163.367
R1522 B.n506 B.n505 163.367
R1523 B.n506 B.n85 163.367
R1524 B.n510 B.n85 163.367
R1525 B.n511 B.n510 163.367
R1526 B.n512 B.n511 163.367
R1527 B.n512 B.n83 163.367
R1528 B.n516 B.n83 163.367
R1529 B.n517 B.n516 163.367
R1530 B.n518 B.n517 163.367
R1531 B.n518 B.n81 163.367
R1532 B.n522 B.n81 163.367
R1533 B.n523 B.n522 163.367
R1534 B.n524 B.n523 163.367
R1535 B.n524 B.n79 163.367
R1536 B.n528 B.n79 163.367
R1537 B.n529 B.n528 163.367
R1538 B.n530 B.n529 163.367
R1539 B.n530 B.n77 163.367
R1540 B.n534 B.n77 163.367
R1541 B.n680 B.n679 163.367
R1542 B.n679 B.n678 163.367
R1543 B.n678 B.n25 163.367
R1544 B.n674 B.n25 163.367
R1545 B.n674 B.n673 163.367
R1546 B.n673 B.n672 163.367
R1547 B.n672 B.n27 163.367
R1548 B.n668 B.n27 163.367
R1549 B.n668 B.n667 163.367
R1550 B.n667 B.n666 163.367
R1551 B.n666 B.n29 163.367
R1552 B.n662 B.n29 163.367
R1553 B.n662 B.n661 163.367
R1554 B.n661 B.n660 163.367
R1555 B.n660 B.n31 163.367
R1556 B.n656 B.n31 163.367
R1557 B.n656 B.n655 163.367
R1558 B.n655 B.n654 163.367
R1559 B.n654 B.n33 163.367
R1560 B.n650 B.n33 163.367
R1561 B.n650 B.n649 163.367
R1562 B.n649 B.n648 163.367
R1563 B.n648 B.n35 163.367
R1564 B.n644 B.n35 163.367
R1565 B.n644 B.n643 163.367
R1566 B.n643 B.n642 163.367
R1567 B.n642 B.n37 163.367
R1568 B.n638 B.n37 163.367
R1569 B.n638 B.n637 163.367
R1570 B.n637 B.n636 163.367
R1571 B.n636 B.n39 163.367
R1572 B.n632 B.n39 163.367
R1573 B.n632 B.n631 163.367
R1574 B.n631 B.n630 163.367
R1575 B.n630 B.n41 163.367
R1576 B.n626 B.n41 163.367
R1577 B.n626 B.n625 163.367
R1578 B.n625 B.n624 163.367
R1579 B.n624 B.n43 163.367
R1580 B.n620 B.n43 163.367
R1581 B.n620 B.n619 163.367
R1582 B.n619 B.n618 163.367
R1583 B.n618 B.n45 163.367
R1584 B.n613 B.n45 163.367
R1585 B.n613 B.n612 163.367
R1586 B.n612 B.n611 163.367
R1587 B.n611 B.n49 163.367
R1588 B.n607 B.n49 163.367
R1589 B.n607 B.n606 163.367
R1590 B.n606 B.n605 163.367
R1591 B.n605 B.n51 163.367
R1592 B.n601 B.n51 163.367
R1593 B.n601 B.n600 163.367
R1594 B.n600 B.n55 163.367
R1595 B.n596 B.n55 163.367
R1596 B.n596 B.n595 163.367
R1597 B.n595 B.n594 163.367
R1598 B.n594 B.n57 163.367
R1599 B.n590 B.n57 163.367
R1600 B.n590 B.n589 163.367
R1601 B.n589 B.n588 163.367
R1602 B.n588 B.n59 163.367
R1603 B.n584 B.n59 163.367
R1604 B.n584 B.n583 163.367
R1605 B.n583 B.n582 163.367
R1606 B.n582 B.n61 163.367
R1607 B.n578 B.n61 163.367
R1608 B.n578 B.n577 163.367
R1609 B.n577 B.n576 163.367
R1610 B.n576 B.n63 163.367
R1611 B.n572 B.n63 163.367
R1612 B.n572 B.n571 163.367
R1613 B.n571 B.n570 163.367
R1614 B.n570 B.n65 163.367
R1615 B.n566 B.n65 163.367
R1616 B.n566 B.n565 163.367
R1617 B.n565 B.n564 163.367
R1618 B.n564 B.n67 163.367
R1619 B.n560 B.n67 163.367
R1620 B.n560 B.n559 163.367
R1621 B.n559 B.n558 163.367
R1622 B.n558 B.n69 163.367
R1623 B.n554 B.n69 163.367
R1624 B.n554 B.n553 163.367
R1625 B.n553 B.n552 163.367
R1626 B.n552 B.n71 163.367
R1627 B.n548 B.n71 163.367
R1628 B.n548 B.n547 163.367
R1629 B.n547 B.n546 163.367
R1630 B.n546 B.n73 163.367
R1631 B.n542 B.n73 163.367
R1632 B.n542 B.n541 163.367
R1633 B.n541 B.n540 163.367
R1634 B.n540 B.n75 163.367
R1635 B.n536 B.n75 163.367
R1636 B.n536 B.n535 163.367
R1637 B.n143 B.n142 76.4126
R1638 B.n151 B.n150 76.4126
R1639 B.n47 B.n46 76.4126
R1640 B.n53 B.n52 76.4126
R1641 B.n144 B.n143 59.5399
R1642 B.n323 B.n151 59.5399
R1643 B.n615 B.n47 59.5399
R1644 B.n54 B.n53 59.5399
R1645 B.n682 B.n681 31.6883
R1646 B.n533 B.n76 31.6883
R1647 B.n405 B.n120 31.6883
R1648 B.n257 B.n256 31.6883
R1649 B B.n747 18.0485
R1650 B.n681 B.n24 10.6151
R1651 B.n677 B.n24 10.6151
R1652 B.n677 B.n676 10.6151
R1653 B.n676 B.n675 10.6151
R1654 B.n675 B.n26 10.6151
R1655 B.n671 B.n26 10.6151
R1656 B.n671 B.n670 10.6151
R1657 B.n670 B.n669 10.6151
R1658 B.n669 B.n28 10.6151
R1659 B.n665 B.n28 10.6151
R1660 B.n665 B.n664 10.6151
R1661 B.n664 B.n663 10.6151
R1662 B.n663 B.n30 10.6151
R1663 B.n659 B.n30 10.6151
R1664 B.n659 B.n658 10.6151
R1665 B.n658 B.n657 10.6151
R1666 B.n657 B.n32 10.6151
R1667 B.n653 B.n32 10.6151
R1668 B.n653 B.n652 10.6151
R1669 B.n652 B.n651 10.6151
R1670 B.n651 B.n34 10.6151
R1671 B.n647 B.n34 10.6151
R1672 B.n647 B.n646 10.6151
R1673 B.n646 B.n645 10.6151
R1674 B.n645 B.n36 10.6151
R1675 B.n641 B.n36 10.6151
R1676 B.n641 B.n640 10.6151
R1677 B.n640 B.n639 10.6151
R1678 B.n639 B.n38 10.6151
R1679 B.n635 B.n38 10.6151
R1680 B.n635 B.n634 10.6151
R1681 B.n634 B.n633 10.6151
R1682 B.n633 B.n40 10.6151
R1683 B.n629 B.n40 10.6151
R1684 B.n629 B.n628 10.6151
R1685 B.n628 B.n627 10.6151
R1686 B.n627 B.n42 10.6151
R1687 B.n623 B.n42 10.6151
R1688 B.n623 B.n622 10.6151
R1689 B.n622 B.n621 10.6151
R1690 B.n621 B.n44 10.6151
R1691 B.n617 B.n44 10.6151
R1692 B.n617 B.n616 10.6151
R1693 B.n614 B.n48 10.6151
R1694 B.n610 B.n48 10.6151
R1695 B.n610 B.n609 10.6151
R1696 B.n609 B.n608 10.6151
R1697 B.n608 B.n50 10.6151
R1698 B.n604 B.n50 10.6151
R1699 B.n604 B.n603 10.6151
R1700 B.n603 B.n602 10.6151
R1701 B.n599 B.n598 10.6151
R1702 B.n598 B.n597 10.6151
R1703 B.n597 B.n56 10.6151
R1704 B.n593 B.n56 10.6151
R1705 B.n593 B.n592 10.6151
R1706 B.n592 B.n591 10.6151
R1707 B.n591 B.n58 10.6151
R1708 B.n587 B.n58 10.6151
R1709 B.n587 B.n586 10.6151
R1710 B.n586 B.n585 10.6151
R1711 B.n585 B.n60 10.6151
R1712 B.n581 B.n60 10.6151
R1713 B.n581 B.n580 10.6151
R1714 B.n580 B.n579 10.6151
R1715 B.n579 B.n62 10.6151
R1716 B.n575 B.n62 10.6151
R1717 B.n575 B.n574 10.6151
R1718 B.n574 B.n573 10.6151
R1719 B.n573 B.n64 10.6151
R1720 B.n569 B.n64 10.6151
R1721 B.n569 B.n568 10.6151
R1722 B.n568 B.n567 10.6151
R1723 B.n567 B.n66 10.6151
R1724 B.n563 B.n66 10.6151
R1725 B.n563 B.n562 10.6151
R1726 B.n562 B.n561 10.6151
R1727 B.n561 B.n68 10.6151
R1728 B.n557 B.n68 10.6151
R1729 B.n557 B.n556 10.6151
R1730 B.n556 B.n555 10.6151
R1731 B.n555 B.n70 10.6151
R1732 B.n551 B.n70 10.6151
R1733 B.n551 B.n550 10.6151
R1734 B.n550 B.n549 10.6151
R1735 B.n549 B.n72 10.6151
R1736 B.n545 B.n72 10.6151
R1737 B.n545 B.n544 10.6151
R1738 B.n544 B.n543 10.6151
R1739 B.n543 B.n74 10.6151
R1740 B.n539 B.n74 10.6151
R1741 B.n539 B.n538 10.6151
R1742 B.n538 B.n537 10.6151
R1743 B.n537 B.n76 10.6151
R1744 B.n406 B.n405 10.6151
R1745 B.n407 B.n406 10.6151
R1746 B.n407 B.n118 10.6151
R1747 B.n411 B.n118 10.6151
R1748 B.n412 B.n411 10.6151
R1749 B.n413 B.n412 10.6151
R1750 B.n413 B.n116 10.6151
R1751 B.n417 B.n116 10.6151
R1752 B.n418 B.n417 10.6151
R1753 B.n419 B.n418 10.6151
R1754 B.n419 B.n114 10.6151
R1755 B.n423 B.n114 10.6151
R1756 B.n424 B.n423 10.6151
R1757 B.n425 B.n424 10.6151
R1758 B.n425 B.n112 10.6151
R1759 B.n429 B.n112 10.6151
R1760 B.n430 B.n429 10.6151
R1761 B.n431 B.n430 10.6151
R1762 B.n431 B.n110 10.6151
R1763 B.n435 B.n110 10.6151
R1764 B.n436 B.n435 10.6151
R1765 B.n437 B.n436 10.6151
R1766 B.n437 B.n108 10.6151
R1767 B.n441 B.n108 10.6151
R1768 B.n442 B.n441 10.6151
R1769 B.n443 B.n442 10.6151
R1770 B.n443 B.n106 10.6151
R1771 B.n447 B.n106 10.6151
R1772 B.n448 B.n447 10.6151
R1773 B.n449 B.n448 10.6151
R1774 B.n449 B.n104 10.6151
R1775 B.n453 B.n104 10.6151
R1776 B.n454 B.n453 10.6151
R1777 B.n455 B.n454 10.6151
R1778 B.n455 B.n102 10.6151
R1779 B.n459 B.n102 10.6151
R1780 B.n460 B.n459 10.6151
R1781 B.n461 B.n460 10.6151
R1782 B.n461 B.n100 10.6151
R1783 B.n465 B.n100 10.6151
R1784 B.n466 B.n465 10.6151
R1785 B.n467 B.n466 10.6151
R1786 B.n467 B.n98 10.6151
R1787 B.n471 B.n98 10.6151
R1788 B.n472 B.n471 10.6151
R1789 B.n473 B.n472 10.6151
R1790 B.n473 B.n96 10.6151
R1791 B.n477 B.n96 10.6151
R1792 B.n478 B.n477 10.6151
R1793 B.n479 B.n478 10.6151
R1794 B.n479 B.n94 10.6151
R1795 B.n483 B.n94 10.6151
R1796 B.n484 B.n483 10.6151
R1797 B.n485 B.n484 10.6151
R1798 B.n485 B.n92 10.6151
R1799 B.n489 B.n92 10.6151
R1800 B.n490 B.n489 10.6151
R1801 B.n491 B.n490 10.6151
R1802 B.n491 B.n90 10.6151
R1803 B.n495 B.n90 10.6151
R1804 B.n496 B.n495 10.6151
R1805 B.n497 B.n496 10.6151
R1806 B.n497 B.n88 10.6151
R1807 B.n501 B.n88 10.6151
R1808 B.n502 B.n501 10.6151
R1809 B.n503 B.n502 10.6151
R1810 B.n503 B.n86 10.6151
R1811 B.n507 B.n86 10.6151
R1812 B.n508 B.n507 10.6151
R1813 B.n509 B.n508 10.6151
R1814 B.n509 B.n84 10.6151
R1815 B.n513 B.n84 10.6151
R1816 B.n514 B.n513 10.6151
R1817 B.n515 B.n514 10.6151
R1818 B.n515 B.n82 10.6151
R1819 B.n519 B.n82 10.6151
R1820 B.n520 B.n519 10.6151
R1821 B.n521 B.n520 10.6151
R1822 B.n521 B.n80 10.6151
R1823 B.n525 B.n80 10.6151
R1824 B.n526 B.n525 10.6151
R1825 B.n527 B.n526 10.6151
R1826 B.n527 B.n78 10.6151
R1827 B.n531 B.n78 10.6151
R1828 B.n532 B.n531 10.6151
R1829 B.n533 B.n532 10.6151
R1830 B.n257 B.n172 10.6151
R1831 B.n261 B.n172 10.6151
R1832 B.n262 B.n261 10.6151
R1833 B.n263 B.n262 10.6151
R1834 B.n263 B.n170 10.6151
R1835 B.n267 B.n170 10.6151
R1836 B.n268 B.n267 10.6151
R1837 B.n269 B.n268 10.6151
R1838 B.n269 B.n168 10.6151
R1839 B.n273 B.n168 10.6151
R1840 B.n274 B.n273 10.6151
R1841 B.n275 B.n274 10.6151
R1842 B.n275 B.n166 10.6151
R1843 B.n279 B.n166 10.6151
R1844 B.n280 B.n279 10.6151
R1845 B.n281 B.n280 10.6151
R1846 B.n281 B.n164 10.6151
R1847 B.n285 B.n164 10.6151
R1848 B.n286 B.n285 10.6151
R1849 B.n287 B.n286 10.6151
R1850 B.n287 B.n162 10.6151
R1851 B.n291 B.n162 10.6151
R1852 B.n292 B.n291 10.6151
R1853 B.n293 B.n292 10.6151
R1854 B.n293 B.n160 10.6151
R1855 B.n297 B.n160 10.6151
R1856 B.n298 B.n297 10.6151
R1857 B.n299 B.n298 10.6151
R1858 B.n299 B.n158 10.6151
R1859 B.n303 B.n158 10.6151
R1860 B.n304 B.n303 10.6151
R1861 B.n305 B.n304 10.6151
R1862 B.n305 B.n156 10.6151
R1863 B.n309 B.n156 10.6151
R1864 B.n310 B.n309 10.6151
R1865 B.n311 B.n310 10.6151
R1866 B.n311 B.n154 10.6151
R1867 B.n315 B.n154 10.6151
R1868 B.n316 B.n315 10.6151
R1869 B.n317 B.n316 10.6151
R1870 B.n317 B.n152 10.6151
R1871 B.n321 B.n152 10.6151
R1872 B.n322 B.n321 10.6151
R1873 B.n324 B.n148 10.6151
R1874 B.n328 B.n148 10.6151
R1875 B.n329 B.n328 10.6151
R1876 B.n330 B.n329 10.6151
R1877 B.n330 B.n146 10.6151
R1878 B.n334 B.n146 10.6151
R1879 B.n335 B.n334 10.6151
R1880 B.n336 B.n335 10.6151
R1881 B.n340 B.n339 10.6151
R1882 B.n341 B.n340 10.6151
R1883 B.n341 B.n140 10.6151
R1884 B.n345 B.n140 10.6151
R1885 B.n346 B.n345 10.6151
R1886 B.n347 B.n346 10.6151
R1887 B.n347 B.n138 10.6151
R1888 B.n351 B.n138 10.6151
R1889 B.n352 B.n351 10.6151
R1890 B.n353 B.n352 10.6151
R1891 B.n353 B.n136 10.6151
R1892 B.n357 B.n136 10.6151
R1893 B.n358 B.n357 10.6151
R1894 B.n359 B.n358 10.6151
R1895 B.n359 B.n134 10.6151
R1896 B.n363 B.n134 10.6151
R1897 B.n364 B.n363 10.6151
R1898 B.n365 B.n364 10.6151
R1899 B.n365 B.n132 10.6151
R1900 B.n369 B.n132 10.6151
R1901 B.n370 B.n369 10.6151
R1902 B.n371 B.n370 10.6151
R1903 B.n371 B.n130 10.6151
R1904 B.n375 B.n130 10.6151
R1905 B.n376 B.n375 10.6151
R1906 B.n377 B.n376 10.6151
R1907 B.n377 B.n128 10.6151
R1908 B.n381 B.n128 10.6151
R1909 B.n382 B.n381 10.6151
R1910 B.n383 B.n382 10.6151
R1911 B.n383 B.n126 10.6151
R1912 B.n387 B.n126 10.6151
R1913 B.n388 B.n387 10.6151
R1914 B.n389 B.n388 10.6151
R1915 B.n389 B.n124 10.6151
R1916 B.n393 B.n124 10.6151
R1917 B.n394 B.n393 10.6151
R1918 B.n395 B.n394 10.6151
R1919 B.n395 B.n122 10.6151
R1920 B.n399 B.n122 10.6151
R1921 B.n400 B.n399 10.6151
R1922 B.n401 B.n400 10.6151
R1923 B.n401 B.n120 10.6151
R1924 B.n256 B.n255 10.6151
R1925 B.n255 B.n174 10.6151
R1926 B.n251 B.n174 10.6151
R1927 B.n251 B.n250 10.6151
R1928 B.n250 B.n249 10.6151
R1929 B.n249 B.n176 10.6151
R1930 B.n245 B.n176 10.6151
R1931 B.n245 B.n244 10.6151
R1932 B.n244 B.n243 10.6151
R1933 B.n243 B.n178 10.6151
R1934 B.n239 B.n178 10.6151
R1935 B.n239 B.n238 10.6151
R1936 B.n238 B.n237 10.6151
R1937 B.n237 B.n180 10.6151
R1938 B.n233 B.n180 10.6151
R1939 B.n233 B.n232 10.6151
R1940 B.n232 B.n231 10.6151
R1941 B.n231 B.n182 10.6151
R1942 B.n227 B.n182 10.6151
R1943 B.n227 B.n226 10.6151
R1944 B.n226 B.n225 10.6151
R1945 B.n225 B.n184 10.6151
R1946 B.n221 B.n184 10.6151
R1947 B.n221 B.n220 10.6151
R1948 B.n220 B.n219 10.6151
R1949 B.n219 B.n186 10.6151
R1950 B.n215 B.n186 10.6151
R1951 B.n215 B.n214 10.6151
R1952 B.n214 B.n213 10.6151
R1953 B.n213 B.n188 10.6151
R1954 B.n209 B.n188 10.6151
R1955 B.n209 B.n208 10.6151
R1956 B.n208 B.n207 10.6151
R1957 B.n207 B.n190 10.6151
R1958 B.n203 B.n190 10.6151
R1959 B.n203 B.n202 10.6151
R1960 B.n202 B.n201 10.6151
R1961 B.n201 B.n192 10.6151
R1962 B.n197 B.n192 10.6151
R1963 B.n197 B.n196 10.6151
R1964 B.n196 B.n195 10.6151
R1965 B.n195 B.n0 10.6151
R1966 B.n743 B.n1 10.6151
R1967 B.n743 B.n742 10.6151
R1968 B.n742 B.n741 10.6151
R1969 B.n741 B.n4 10.6151
R1970 B.n737 B.n4 10.6151
R1971 B.n737 B.n736 10.6151
R1972 B.n736 B.n735 10.6151
R1973 B.n735 B.n6 10.6151
R1974 B.n731 B.n6 10.6151
R1975 B.n731 B.n730 10.6151
R1976 B.n730 B.n729 10.6151
R1977 B.n729 B.n8 10.6151
R1978 B.n725 B.n8 10.6151
R1979 B.n725 B.n724 10.6151
R1980 B.n724 B.n723 10.6151
R1981 B.n723 B.n10 10.6151
R1982 B.n719 B.n10 10.6151
R1983 B.n719 B.n718 10.6151
R1984 B.n718 B.n717 10.6151
R1985 B.n717 B.n12 10.6151
R1986 B.n713 B.n12 10.6151
R1987 B.n713 B.n712 10.6151
R1988 B.n712 B.n711 10.6151
R1989 B.n711 B.n14 10.6151
R1990 B.n707 B.n14 10.6151
R1991 B.n707 B.n706 10.6151
R1992 B.n706 B.n705 10.6151
R1993 B.n705 B.n16 10.6151
R1994 B.n701 B.n16 10.6151
R1995 B.n701 B.n700 10.6151
R1996 B.n700 B.n699 10.6151
R1997 B.n699 B.n18 10.6151
R1998 B.n695 B.n18 10.6151
R1999 B.n695 B.n694 10.6151
R2000 B.n694 B.n693 10.6151
R2001 B.n693 B.n20 10.6151
R2002 B.n689 B.n20 10.6151
R2003 B.n689 B.n688 10.6151
R2004 B.n688 B.n687 10.6151
R2005 B.n687 B.n22 10.6151
R2006 B.n683 B.n22 10.6151
R2007 B.n683 B.n682 10.6151
R2008 B.n615 B.n614 6.5566
R2009 B.n602 B.n54 6.5566
R2010 B.n324 B.n323 6.5566
R2011 B.n336 B.n144 6.5566
R2012 B.n616 B.n615 4.05904
R2013 B.n599 B.n54 4.05904
R2014 B.n323 B.n322 4.05904
R2015 B.n339 B.n144 4.05904
R2016 B.n747 B.n0 2.81026
R2017 B.n747 B.n1 2.81026
R2018 VN.n1 VN.t0 119.895
R2019 VN.n0 VN.t1 119.895
R2020 VN.n0 VN.t2 118.65
R2021 VN.n1 VN.t3 118.65
R2022 VN VN.n1 52.32
R2023 VN VN.n0 2.08893
R2024 VDD2.n2 VDD2.n0 115.757
R2025 VDD2.n2 VDD2.n1 70.8778
R2026 VDD2.n1 VDD2.t0 2.55392
R2027 VDD2.n1 VDD2.t3 2.55392
R2028 VDD2.n0 VDD2.t2 2.55392
R2029 VDD2.n0 VDD2.t1 2.55392
R2030 VDD2 VDD2.n2 0.0586897
C0 VN VP 7.05245f
C1 B VN 1.30891f
C2 VDD1 VP 5.58754f
C3 B VDD1 1.46029f
C4 VDD2 VTAIL 5.89436f
C5 VTAIL w_n3334_n3514# 4.16762f
C6 VN VDD1 0.150065f
C7 VDD2 w_n3334_n3514# 1.7427f
C8 VTAIL VP 5.32286f
C9 B VTAIL 5.60919f
C10 VDD2 VP 0.458725f
C11 VP w_n3334_n3514# 6.27094f
C12 B VDD2 1.52916f
C13 B w_n3334_n3514# 10.6923f
C14 VTAIL VN 5.30876f
C15 VTAIL VDD1 5.83338f
C16 B VP 2.02909f
C17 VDD2 VN 5.27987f
C18 VN w_n3334_n3514# 5.83978f
C19 VDD2 VDD1 1.27025f
C20 VDD1 w_n3334_n3514# 1.66431f
C21 VDD2 VSUBS 1.130199f
C22 VDD1 VSUBS 6.41322f
C23 VTAIL VSUBS 1.376579f
C24 VN VSUBS 6.03758f
C25 VP VSUBS 2.851126f
C26 B VSUBS 5.207374f
C27 w_n3334_n3514# VSUBS 0.144069p
C28 VDD2.t2 VSUBS 0.273554f
C29 VDD2.t1 VSUBS 0.273554f
C30 VDD2.n0 VSUBS 2.96651f
C31 VDD2.t0 VSUBS 0.273554f
C32 VDD2.t3 VSUBS 0.273554f
C33 VDD2.n1 VSUBS 2.14608f
C34 VDD2.n2 VSUBS 4.68973f
C35 VN.t2 VSUBS 3.80254f
C36 VN.t1 VSUBS 3.81646f
C37 VN.n0 VSUBS 2.2711f
C38 VN.t0 VSUBS 3.81646f
C39 VN.t3 VSUBS 3.80254f
C40 VN.n1 VSUBS 4.04743f
C41 B.n0 VSUBS 0.004343f
C42 B.n1 VSUBS 0.004343f
C43 B.n2 VSUBS 0.006868f
C44 B.n3 VSUBS 0.006868f
C45 B.n4 VSUBS 0.006868f
C46 B.n5 VSUBS 0.006868f
C47 B.n6 VSUBS 0.006868f
C48 B.n7 VSUBS 0.006868f
C49 B.n8 VSUBS 0.006868f
C50 B.n9 VSUBS 0.006868f
C51 B.n10 VSUBS 0.006868f
C52 B.n11 VSUBS 0.006868f
C53 B.n12 VSUBS 0.006868f
C54 B.n13 VSUBS 0.006868f
C55 B.n14 VSUBS 0.006868f
C56 B.n15 VSUBS 0.006868f
C57 B.n16 VSUBS 0.006868f
C58 B.n17 VSUBS 0.006868f
C59 B.n18 VSUBS 0.006868f
C60 B.n19 VSUBS 0.006868f
C61 B.n20 VSUBS 0.006868f
C62 B.n21 VSUBS 0.006868f
C63 B.n22 VSUBS 0.006868f
C64 B.n23 VSUBS 0.015481f
C65 B.n24 VSUBS 0.006868f
C66 B.n25 VSUBS 0.006868f
C67 B.n26 VSUBS 0.006868f
C68 B.n27 VSUBS 0.006868f
C69 B.n28 VSUBS 0.006868f
C70 B.n29 VSUBS 0.006868f
C71 B.n30 VSUBS 0.006868f
C72 B.n31 VSUBS 0.006868f
C73 B.n32 VSUBS 0.006868f
C74 B.n33 VSUBS 0.006868f
C75 B.n34 VSUBS 0.006868f
C76 B.n35 VSUBS 0.006868f
C77 B.n36 VSUBS 0.006868f
C78 B.n37 VSUBS 0.006868f
C79 B.n38 VSUBS 0.006868f
C80 B.n39 VSUBS 0.006868f
C81 B.n40 VSUBS 0.006868f
C82 B.n41 VSUBS 0.006868f
C83 B.n42 VSUBS 0.006868f
C84 B.n43 VSUBS 0.006868f
C85 B.n44 VSUBS 0.006868f
C86 B.n45 VSUBS 0.006868f
C87 B.t5 VSUBS 0.223073f
C88 B.t4 VSUBS 0.264351f
C89 B.t3 VSUBS 2.09001f
C90 B.n46 VSUBS 0.421618f
C91 B.n47 VSUBS 0.261077f
C92 B.n48 VSUBS 0.006868f
C93 B.n49 VSUBS 0.006868f
C94 B.n50 VSUBS 0.006868f
C95 B.n51 VSUBS 0.006868f
C96 B.t11 VSUBS 0.223076f
C97 B.t10 VSUBS 0.264353f
C98 B.t9 VSUBS 2.09001f
C99 B.n52 VSUBS 0.421615f
C100 B.n53 VSUBS 0.261074f
C101 B.n54 VSUBS 0.015913f
C102 B.n55 VSUBS 0.006868f
C103 B.n56 VSUBS 0.006868f
C104 B.n57 VSUBS 0.006868f
C105 B.n58 VSUBS 0.006868f
C106 B.n59 VSUBS 0.006868f
C107 B.n60 VSUBS 0.006868f
C108 B.n61 VSUBS 0.006868f
C109 B.n62 VSUBS 0.006868f
C110 B.n63 VSUBS 0.006868f
C111 B.n64 VSUBS 0.006868f
C112 B.n65 VSUBS 0.006868f
C113 B.n66 VSUBS 0.006868f
C114 B.n67 VSUBS 0.006868f
C115 B.n68 VSUBS 0.006868f
C116 B.n69 VSUBS 0.006868f
C117 B.n70 VSUBS 0.006868f
C118 B.n71 VSUBS 0.006868f
C119 B.n72 VSUBS 0.006868f
C120 B.n73 VSUBS 0.006868f
C121 B.n74 VSUBS 0.006868f
C122 B.n75 VSUBS 0.006868f
C123 B.n76 VSUBS 0.015196f
C124 B.n77 VSUBS 0.006868f
C125 B.n78 VSUBS 0.006868f
C126 B.n79 VSUBS 0.006868f
C127 B.n80 VSUBS 0.006868f
C128 B.n81 VSUBS 0.006868f
C129 B.n82 VSUBS 0.006868f
C130 B.n83 VSUBS 0.006868f
C131 B.n84 VSUBS 0.006868f
C132 B.n85 VSUBS 0.006868f
C133 B.n86 VSUBS 0.006868f
C134 B.n87 VSUBS 0.006868f
C135 B.n88 VSUBS 0.006868f
C136 B.n89 VSUBS 0.006868f
C137 B.n90 VSUBS 0.006868f
C138 B.n91 VSUBS 0.006868f
C139 B.n92 VSUBS 0.006868f
C140 B.n93 VSUBS 0.006868f
C141 B.n94 VSUBS 0.006868f
C142 B.n95 VSUBS 0.006868f
C143 B.n96 VSUBS 0.006868f
C144 B.n97 VSUBS 0.006868f
C145 B.n98 VSUBS 0.006868f
C146 B.n99 VSUBS 0.006868f
C147 B.n100 VSUBS 0.006868f
C148 B.n101 VSUBS 0.006868f
C149 B.n102 VSUBS 0.006868f
C150 B.n103 VSUBS 0.006868f
C151 B.n104 VSUBS 0.006868f
C152 B.n105 VSUBS 0.006868f
C153 B.n106 VSUBS 0.006868f
C154 B.n107 VSUBS 0.006868f
C155 B.n108 VSUBS 0.006868f
C156 B.n109 VSUBS 0.006868f
C157 B.n110 VSUBS 0.006868f
C158 B.n111 VSUBS 0.006868f
C159 B.n112 VSUBS 0.006868f
C160 B.n113 VSUBS 0.006868f
C161 B.n114 VSUBS 0.006868f
C162 B.n115 VSUBS 0.006868f
C163 B.n116 VSUBS 0.006868f
C164 B.n117 VSUBS 0.006868f
C165 B.n118 VSUBS 0.006868f
C166 B.n119 VSUBS 0.006868f
C167 B.n120 VSUBS 0.016032f
C168 B.n121 VSUBS 0.006868f
C169 B.n122 VSUBS 0.006868f
C170 B.n123 VSUBS 0.006868f
C171 B.n124 VSUBS 0.006868f
C172 B.n125 VSUBS 0.006868f
C173 B.n126 VSUBS 0.006868f
C174 B.n127 VSUBS 0.006868f
C175 B.n128 VSUBS 0.006868f
C176 B.n129 VSUBS 0.006868f
C177 B.n130 VSUBS 0.006868f
C178 B.n131 VSUBS 0.006868f
C179 B.n132 VSUBS 0.006868f
C180 B.n133 VSUBS 0.006868f
C181 B.n134 VSUBS 0.006868f
C182 B.n135 VSUBS 0.006868f
C183 B.n136 VSUBS 0.006868f
C184 B.n137 VSUBS 0.006868f
C185 B.n138 VSUBS 0.006868f
C186 B.n139 VSUBS 0.006868f
C187 B.n140 VSUBS 0.006868f
C188 B.n141 VSUBS 0.006868f
C189 B.t1 VSUBS 0.223076f
C190 B.t2 VSUBS 0.264353f
C191 B.t0 VSUBS 2.09001f
C192 B.n142 VSUBS 0.421615f
C193 B.n143 VSUBS 0.261074f
C194 B.n144 VSUBS 0.015913f
C195 B.n145 VSUBS 0.006868f
C196 B.n146 VSUBS 0.006868f
C197 B.n147 VSUBS 0.006868f
C198 B.n148 VSUBS 0.006868f
C199 B.n149 VSUBS 0.006868f
C200 B.t7 VSUBS 0.223073f
C201 B.t8 VSUBS 0.264351f
C202 B.t6 VSUBS 2.09001f
C203 B.n150 VSUBS 0.421618f
C204 B.n151 VSUBS 0.261077f
C205 B.n152 VSUBS 0.006868f
C206 B.n153 VSUBS 0.006868f
C207 B.n154 VSUBS 0.006868f
C208 B.n155 VSUBS 0.006868f
C209 B.n156 VSUBS 0.006868f
C210 B.n157 VSUBS 0.006868f
C211 B.n158 VSUBS 0.006868f
C212 B.n159 VSUBS 0.006868f
C213 B.n160 VSUBS 0.006868f
C214 B.n161 VSUBS 0.006868f
C215 B.n162 VSUBS 0.006868f
C216 B.n163 VSUBS 0.006868f
C217 B.n164 VSUBS 0.006868f
C218 B.n165 VSUBS 0.006868f
C219 B.n166 VSUBS 0.006868f
C220 B.n167 VSUBS 0.006868f
C221 B.n168 VSUBS 0.006868f
C222 B.n169 VSUBS 0.006868f
C223 B.n170 VSUBS 0.006868f
C224 B.n171 VSUBS 0.006868f
C225 B.n172 VSUBS 0.006868f
C226 B.n173 VSUBS 0.015481f
C227 B.n174 VSUBS 0.006868f
C228 B.n175 VSUBS 0.006868f
C229 B.n176 VSUBS 0.006868f
C230 B.n177 VSUBS 0.006868f
C231 B.n178 VSUBS 0.006868f
C232 B.n179 VSUBS 0.006868f
C233 B.n180 VSUBS 0.006868f
C234 B.n181 VSUBS 0.006868f
C235 B.n182 VSUBS 0.006868f
C236 B.n183 VSUBS 0.006868f
C237 B.n184 VSUBS 0.006868f
C238 B.n185 VSUBS 0.006868f
C239 B.n186 VSUBS 0.006868f
C240 B.n187 VSUBS 0.006868f
C241 B.n188 VSUBS 0.006868f
C242 B.n189 VSUBS 0.006868f
C243 B.n190 VSUBS 0.006868f
C244 B.n191 VSUBS 0.006868f
C245 B.n192 VSUBS 0.006868f
C246 B.n193 VSUBS 0.006868f
C247 B.n194 VSUBS 0.006868f
C248 B.n195 VSUBS 0.006868f
C249 B.n196 VSUBS 0.006868f
C250 B.n197 VSUBS 0.006868f
C251 B.n198 VSUBS 0.006868f
C252 B.n199 VSUBS 0.006868f
C253 B.n200 VSUBS 0.006868f
C254 B.n201 VSUBS 0.006868f
C255 B.n202 VSUBS 0.006868f
C256 B.n203 VSUBS 0.006868f
C257 B.n204 VSUBS 0.006868f
C258 B.n205 VSUBS 0.006868f
C259 B.n206 VSUBS 0.006868f
C260 B.n207 VSUBS 0.006868f
C261 B.n208 VSUBS 0.006868f
C262 B.n209 VSUBS 0.006868f
C263 B.n210 VSUBS 0.006868f
C264 B.n211 VSUBS 0.006868f
C265 B.n212 VSUBS 0.006868f
C266 B.n213 VSUBS 0.006868f
C267 B.n214 VSUBS 0.006868f
C268 B.n215 VSUBS 0.006868f
C269 B.n216 VSUBS 0.006868f
C270 B.n217 VSUBS 0.006868f
C271 B.n218 VSUBS 0.006868f
C272 B.n219 VSUBS 0.006868f
C273 B.n220 VSUBS 0.006868f
C274 B.n221 VSUBS 0.006868f
C275 B.n222 VSUBS 0.006868f
C276 B.n223 VSUBS 0.006868f
C277 B.n224 VSUBS 0.006868f
C278 B.n225 VSUBS 0.006868f
C279 B.n226 VSUBS 0.006868f
C280 B.n227 VSUBS 0.006868f
C281 B.n228 VSUBS 0.006868f
C282 B.n229 VSUBS 0.006868f
C283 B.n230 VSUBS 0.006868f
C284 B.n231 VSUBS 0.006868f
C285 B.n232 VSUBS 0.006868f
C286 B.n233 VSUBS 0.006868f
C287 B.n234 VSUBS 0.006868f
C288 B.n235 VSUBS 0.006868f
C289 B.n236 VSUBS 0.006868f
C290 B.n237 VSUBS 0.006868f
C291 B.n238 VSUBS 0.006868f
C292 B.n239 VSUBS 0.006868f
C293 B.n240 VSUBS 0.006868f
C294 B.n241 VSUBS 0.006868f
C295 B.n242 VSUBS 0.006868f
C296 B.n243 VSUBS 0.006868f
C297 B.n244 VSUBS 0.006868f
C298 B.n245 VSUBS 0.006868f
C299 B.n246 VSUBS 0.006868f
C300 B.n247 VSUBS 0.006868f
C301 B.n248 VSUBS 0.006868f
C302 B.n249 VSUBS 0.006868f
C303 B.n250 VSUBS 0.006868f
C304 B.n251 VSUBS 0.006868f
C305 B.n252 VSUBS 0.006868f
C306 B.n253 VSUBS 0.006868f
C307 B.n254 VSUBS 0.006868f
C308 B.n255 VSUBS 0.006868f
C309 B.n256 VSUBS 0.015481f
C310 B.n257 VSUBS 0.016032f
C311 B.n258 VSUBS 0.016032f
C312 B.n259 VSUBS 0.006868f
C313 B.n260 VSUBS 0.006868f
C314 B.n261 VSUBS 0.006868f
C315 B.n262 VSUBS 0.006868f
C316 B.n263 VSUBS 0.006868f
C317 B.n264 VSUBS 0.006868f
C318 B.n265 VSUBS 0.006868f
C319 B.n266 VSUBS 0.006868f
C320 B.n267 VSUBS 0.006868f
C321 B.n268 VSUBS 0.006868f
C322 B.n269 VSUBS 0.006868f
C323 B.n270 VSUBS 0.006868f
C324 B.n271 VSUBS 0.006868f
C325 B.n272 VSUBS 0.006868f
C326 B.n273 VSUBS 0.006868f
C327 B.n274 VSUBS 0.006868f
C328 B.n275 VSUBS 0.006868f
C329 B.n276 VSUBS 0.006868f
C330 B.n277 VSUBS 0.006868f
C331 B.n278 VSUBS 0.006868f
C332 B.n279 VSUBS 0.006868f
C333 B.n280 VSUBS 0.006868f
C334 B.n281 VSUBS 0.006868f
C335 B.n282 VSUBS 0.006868f
C336 B.n283 VSUBS 0.006868f
C337 B.n284 VSUBS 0.006868f
C338 B.n285 VSUBS 0.006868f
C339 B.n286 VSUBS 0.006868f
C340 B.n287 VSUBS 0.006868f
C341 B.n288 VSUBS 0.006868f
C342 B.n289 VSUBS 0.006868f
C343 B.n290 VSUBS 0.006868f
C344 B.n291 VSUBS 0.006868f
C345 B.n292 VSUBS 0.006868f
C346 B.n293 VSUBS 0.006868f
C347 B.n294 VSUBS 0.006868f
C348 B.n295 VSUBS 0.006868f
C349 B.n296 VSUBS 0.006868f
C350 B.n297 VSUBS 0.006868f
C351 B.n298 VSUBS 0.006868f
C352 B.n299 VSUBS 0.006868f
C353 B.n300 VSUBS 0.006868f
C354 B.n301 VSUBS 0.006868f
C355 B.n302 VSUBS 0.006868f
C356 B.n303 VSUBS 0.006868f
C357 B.n304 VSUBS 0.006868f
C358 B.n305 VSUBS 0.006868f
C359 B.n306 VSUBS 0.006868f
C360 B.n307 VSUBS 0.006868f
C361 B.n308 VSUBS 0.006868f
C362 B.n309 VSUBS 0.006868f
C363 B.n310 VSUBS 0.006868f
C364 B.n311 VSUBS 0.006868f
C365 B.n312 VSUBS 0.006868f
C366 B.n313 VSUBS 0.006868f
C367 B.n314 VSUBS 0.006868f
C368 B.n315 VSUBS 0.006868f
C369 B.n316 VSUBS 0.006868f
C370 B.n317 VSUBS 0.006868f
C371 B.n318 VSUBS 0.006868f
C372 B.n319 VSUBS 0.006868f
C373 B.n320 VSUBS 0.006868f
C374 B.n321 VSUBS 0.006868f
C375 B.n322 VSUBS 0.004747f
C376 B.n323 VSUBS 0.015913f
C377 B.n324 VSUBS 0.005555f
C378 B.n325 VSUBS 0.006868f
C379 B.n326 VSUBS 0.006868f
C380 B.n327 VSUBS 0.006868f
C381 B.n328 VSUBS 0.006868f
C382 B.n329 VSUBS 0.006868f
C383 B.n330 VSUBS 0.006868f
C384 B.n331 VSUBS 0.006868f
C385 B.n332 VSUBS 0.006868f
C386 B.n333 VSUBS 0.006868f
C387 B.n334 VSUBS 0.006868f
C388 B.n335 VSUBS 0.006868f
C389 B.n336 VSUBS 0.005555f
C390 B.n337 VSUBS 0.006868f
C391 B.n338 VSUBS 0.006868f
C392 B.n339 VSUBS 0.004747f
C393 B.n340 VSUBS 0.006868f
C394 B.n341 VSUBS 0.006868f
C395 B.n342 VSUBS 0.006868f
C396 B.n343 VSUBS 0.006868f
C397 B.n344 VSUBS 0.006868f
C398 B.n345 VSUBS 0.006868f
C399 B.n346 VSUBS 0.006868f
C400 B.n347 VSUBS 0.006868f
C401 B.n348 VSUBS 0.006868f
C402 B.n349 VSUBS 0.006868f
C403 B.n350 VSUBS 0.006868f
C404 B.n351 VSUBS 0.006868f
C405 B.n352 VSUBS 0.006868f
C406 B.n353 VSUBS 0.006868f
C407 B.n354 VSUBS 0.006868f
C408 B.n355 VSUBS 0.006868f
C409 B.n356 VSUBS 0.006868f
C410 B.n357 VSUBS 0.006868f
C411 B.n358 VSUBS 0.006868f
C412 B.n359 VSUBS 0.006868f
C413 B.n360 VSUBS 0.006868f
C414 B.n361 VSUBS 0.006868f
C415 B.n362 VSUBS 0.006868f
C416 B.n363 VSUBS 0.006868f
C417 B.n364 VSUBS 0.006868f
C418 B.n365 VSUBS 0.006868f
C419 B.n366 VSUBS 0.006868f
C420 B.n367 VSUBS 0.006868f
C421 B.n368 VSUBS 0.006868f
C422 B.n369 VSUBS 0.006868f
C423 B.n370 VSUBS 0.006868f
C424 B.n371 VSUBS 0.006868f
C425 B.n372 VSUBS 0.006868f
C426 B.n373 VSUBS 0.006868f
C427 B.n374 VSUBS 0.006868f
C428 B.n375 VSUBS 0.006868f
C429 B.n376 VSUBS 0.006868f
C430 B.n377 VSUBS 0.006868f
C431 B.n378 VSUBS 0.006868f
C432 B.n379 VSUBS 0.006868f
C433 B.n380 VSUBS 0.006868f
C434 B.n381 VSUBS 0.006868f
C435 B.n382 VSUBS 0.006868f
C436 B.n383 VSUBS 0.006868f
C437 B.n384 VSUBS 0.006868f
C438 B.n385 VSUBS 0.006868f
C439 B.n386 VSUBS 0.006868f
C440 B.n387 VSUBS 0.006868f
C441 B.n388 VSUBS 0.006868f
C442 B.n389 VSUBS 0.006868f
C443 B.n390 VSUBS 0.006868f
C444 B.n391 VSUBS 0.006868f
C445 B.n392 VSUBS 0.006868f
C446 B.n393 VSUBS 0.006868f
C447 B.n394 VSUBS 0.006868f
C448 B.n395 VSUBS 0.006868f
C449 B.n396 VSUBS 0.006868f
C450 B.n397 VSUBS 0.006868f
C451 B.n398 VSUBS 0.006868f
C452 B.n399 VSUBS 0.006868f
C453 B.n400 VSUBS 0.006868f
C454 B.n401 VSUBS 0.006868f
C455 B.n402 VSUBS 0.006868f
C456 B.n403 VSUBS 0.016032f
C457 B.n404 VSUBS 0.015481f
C458 B.n405 VSUBS 0.015481f
C459 B.n406 VSUBS 0.006868f
C460 B.n407 VSUBS 0.006868f
C461 B.n408 VSUBS 0.006868f
C462 B.n409 VSUBS 0.006868f
C463 B.n410 VSUBS 0.006868f
C464 B.n411 VSUBS 0.006868f
C465 B.n412 VSUBS 0.006868f
C466 B.n413 VSUBS 0.006868f
C467 B.n414 VSUBS 0.006868f
C468 B.n415 VSUBS 0.006868f
C469 B.n416 VSUBS 0.006868f
C470 B.n417 VSUBS 0.006868f
C471 B.n418 VSUBS 0.006868f
C472 B.n419 VSUBS 0.006868f
C473 B.n420 VSUBS 0.006868f
C474 B.n421 VSUBS 0.006868f
C475 B.n422 VSUBS 0.006868f
C476 B.n423 VSUBS 0.006868f
C477 B.n424 VSUBS 0.006868f
C478 B.n425 VSUBS 0.006868f
C479 B.n426 VSUBS 0.006868f
C480 B.n427 VSUBS 0.006868f
C481 B.n428 VSUBS 0.006868f
C482 B.n429 VSUBS 0.006868f
C483 B.n430 VSUBS 0.006868f
C484 B.n431 VSUBS 0.006868f
C485 B.n432 VSUBS 0.006868f
C486 B.n433 VSUBS 0.006868f
C487 B.n434 VSUBS 0.006868f
C488 B.n435 VSUBS 0.006868f
C489 B.n436 VSUBS 0.006868f
C490 B.n437 VSUBS 0.006868f
C491 B.n438 VSUBS 0.006868f
C492 B.n439 VSUBS 0.006868f
C493 B.n440 VSUBS 0.006868f
C494 B.n441 VSUBS 0.006868f
C495 B.n442 VSUBS 0.006868f
C496 B.n443 VSUBS 0.006868f
C497 B.n444 VSUBS 0.006868f
C498 B.n445 VSUBS 0.006868f
C499 B.n446 VSUBS 0.006868f
C500 B.n447 VSUBS 0.006868f
C501 B.n448 VSUBS 0.006868f
C502 B.n449 VSUBS 0.006868f
C503 B.n450 VSUBS 0.006868f
C504 B.n451 VSUBS 0.006868f
C505 B.n452 VSUBS 0.006868f
C506 B.n453 VSUBS 0.006868f
C507 B.n454 VSUBS 0.006868f
C508 B.n455 VSUBS 0.006868f
C509 B.n456 VSUBS 0.006868f
C510 B.n457 VSUBS 0.006868f
C511 B.n458 VSUBS 0.006868f
C512 B.n459 VSUBS 0.006868f
C513 B.n460 VSUBS 0.006868f
C514 B.n461 VSUBS 0.006868f
C515 B.n462 VSUBS 0.006868f
C516 B.n463 VSUBS 0.006868f
C517 B.n464 VSUBS 0.006868f
C518 B.n465 VSUBS 0.006868f
C519 B.n466 VSUBS 0.006868f
C520 B.n467 VSUBS 0.006868f
C521 B.n468 VSUBS 0.006868f
C522 B.n469 VSUBS 0.006868f
C523 B.n470 VSUBS 0.006868f
C524 B.n471 VSUBS 0.006868f
C525 B.n472 VSUBS 0.006868f
C526 B.n473 VSUBS 0.006868f
C527 B.n474 VSUBS 0.006868f
C528 B.n475 VSUBS 0.006868f
C529 B.n476 VSUBS 0.006868f
C530 B.n477 VSUBS 0.006868f
C531 B.n478 VSUBS 0.006868f
C532 B.n479 VSUBS 0.006868f
C533 B.n480 VSUBS 0.006868f
C534 B.n481 VSUBS 0.006868f
C535 B.n482 VSUBS 0.006868f
C536 B.n483 VSUBS 0.006868f
C537 B.n484 VSUBS 0.006868f
C538 B.n485 VSUBS 0.006868f
C539 B.n486 VSUBS 0.006868f
C540 B.n487 VSUBS 0.006868f
C541 B.n488 VSUBS 0.006868f
C542 B.n489 VSUBS 0.006868f
C543 B.n490 VSUBS 0.006868f
C544 B.n491 VSUBS 0.006868f
C545 B.n492 VSUBS 0.006868f
C546 B.n493 VSUBS 0.006868f
C547 B.n494 VSUBS 0.006868f
C548 B.n495 VSUBS 0.006868f
C549 B.n496 VSUBS 0.006868f
C550 B.n497 VSUBS 0.006868f
C551 B.n498 VSUBS 0.006868f
C552 B.n499 VSUBS 0.006868f
C553 B.n500 VSUBS 0.006868f
C554 B.n501 VSUBS 0.006868f
C555 B.n502 VSUBS 0.006868f
C556 B.n503 VSUBS 0.006868f
C557 B.n504 VSUBS 0.006868f
C558 B.n505 VSUBS 0.006868f
C559 B.n506 VSUBS 0.006868f
C560 B.n507 VSUBS 0.006868f
C561 B.n508 VSUBS 0.006868f
C562 B.n509 VSUBS 0.006868f
C563 B.n510 VSUBS 0.006868f
C564 B.n511 VSUBS 0.006868f
C565 B.n512 VSUBS 0.006868f
C566 B.n513 VSUBS 0.006868f
C567 B.n514 VSUBS 0.006868f
C568 B.n515 VSUBS 0.006868f
C569 B.n516 VSUBS 0.006868f
C570 B.n517 VSUBS 0.006868f
C571 B.n518 VSUBS 0.006868f
C572 B.n519 VSUBS 0.006868f
C573 B.n520 VSUBS 0.006868f
C574 B.n521 VSUBS 0.006868f
C575 B.n522 VSUBS 0.006868f
C576 B.n523 VSUBS 0.006868f
C577 B.n524 VSUBS 0.006868f
C578 B.n525 VSUBS 0.006868f
C579 B.n526 VSUBS 0.006868f
C580 B.n527 VSUBS 0.006868f
C581 B.n528 VSUBS 0.006868f
C582 B.n529 VSUBS 0.006868f
C583 B.n530 VSUBS 0.006868f
C584 B.n531 VSUBS 0.006868f
C585 B.n532 VSUBS 0.006868f
C586 B.n533 VSUBS 0.016318f
C587 B.n534 VSUBS 0.015481f
C588 B.n535 VSUBS 0.016032f
C589 B.n536 VSUBS 0.006868f
C590 B.n537 VSUBS 0.006868f
C591 B.n538 VSUBS 0.006868f
C592 B.n539 VSUBS 0.006868f
C593 B.n540 VSUBS 0.006868f
C594 B.n541 VSUBS 0.006868f
C595 B.n542 VSUBS 0.006868f
C596 B.n543 VSUBS 0.006868f
C597 B.n544 VSUBS 0.006868f
C598 B.n545 VSUBS 0.006868f
C599 B.n546 VSUBS 0.006868f
C600 B.n547 VSUBS 0.006868f
C601 B.n548 VSUBS 0.006868f
C602 B.n549 VSUBS 0.006868f
C603 B.n550 VSUBS 0.006868f
C604 B.n551 VSUBS 0.006868f
C605 B.n552 VSUBS 0.006868f
C606 B.n553 VSUBS 0.006868f
C607 B.n554 VSUBS 0.006868f
C608 B.n555 VSUBS 0.006868f
C609 B.n556 VSUBS 0.006868f
C610 B.n557 VSUBS 0.006868f
C611 B.n558 VSUBS 0.006868f
C612 B.n559 VSUBS 0.006868f
C613 B.n560 VSUBS 0.006868f
C614 B.n561 VSUBS 0.006868f
C615 B.n562 VSUBS 0.006868f
C616 B.n563 VSUBS 0.006868f
C617 B.n564 VSUBS 0.006868f
C618 B.n565 VSUBS 0.006868f
C619 B.n566 VSUBS 0.006868f
C620 B.n567 VSUBS 0.006868f
C621 B.n568 VSUBS 0.006868f
C622 B.n569 VSUBS 0.006868f
C623 B.n570 VSUBS 0.006868f
C624 B.n571 VSUBS 0.006868f
C625 B.n572 VSUBS 0.006868f
C626 B.n573 VSUBS 0.006868f
C627 B.n574 VSUBS 0.006868f
C628 B.n575 VSUBS 0.006868f
C629 B.n576 VSUBS 0.006868f
C630 B.n577 VSUBS 0.006868f
C631 B.n578 VSUBS 0.006868f
C632 B.n579 VSUBS 0.006868f
C633 B.n580 VSUBS 0.006868f
C634 B.n581 VSUBS 0.006868f
C635 B.n582 VSUBS 0.006868f
C636 B.n583 VSUBS 0.006868f
C637 B.n584 VSUBS 0.006868f
C638 B.n585 VSUBS 0.006868f
C639 B.n586 VSUBS 0.006868f
C640 B.n587 VSUBS 0.006868f
C641 B.n588 VSUBS 0.006868f
C642 B.n589 VSUBS 0.006868f
C643 B.n590 VSUBS 0.006868f
C644 B.n591 VSUBS 0.006868f
C645 B.n592 VSUBS 0.006868f
C646 B.n593 VSUBS 0.006868f
C647 B.n594 VSUBS 0.006868f
C648 B.n595 VSUBS 0.006868f
C649 B.n596 VSUBS 0.006868f
C650 B.n597 VSUBS 0.006868f
C651 B.n598 VSUBS 0.006868f
C652 B.n599 VSUBS 0.004747f
C653 B.n600 VSUBS 0.006868f
C654 B.n601 VSUBS 0.006868f
C655 B.n602 VSUBS 0.005555f
C656 B.n603 VSUBS 0.006868f
C657 B.n604 VSUBS 0.006868f
C658 B.n605 VSUBS 0.006868f
C659 B.n606 VSUBS 0.006868f
C660 B.n607 VSUBS 0.006868f
C661 B.n608 VSUBS 0.006868f
C662 B.n609 VSUBS 0.006868f
C663 B.n610 VSUBS 0.006868f
C664 B.n611 VSUBS 0.006868f
C665 B.n612 VSUBS 0.006868f
C666 B.n613 VSUBS 0.006868f
C667 B.n614 VSUBS 0.005555f
C668 B.n615 VSUBS 0.015913f
C669 B.n616 VSUBS 0.004747f
C670 B.n617 VSUBS 0.006868f
C671 B.n618 VSUBS 0.006868f
C672 B.n619 VSUBS 0.006868f
C673 B.n620 VSUBS 0.006868f
C674 B.n621 VSUBS 0.006868f
C675 B.n622 VSUBS 0.006868f
C676 B.n623 VSUBS 0.006868f
C677 B.n624 VSUBS 0.006868f
C678 B.n625 VSUBS 0.006868f
C679 B.n626 VSUBS 0.006868f
C680 B.n627 VSUBS 0.006868f
C681 B.n628 VSUBS 0.006868f
C682 B.n629 VSUBS 0.006868f
C683 B.n630 VSUBS 0.006868f
C684 B.n631 VSUBS 0.006868f
C685 B.n632 VSUBS 0.006868f
C686 B.n633 VSUBS 0.006868f
C687 B.n634 VSUBS 0.006868f
C688 B.n635 VSUBS 0.006868f
C689 B.n636 VSUBS 0.006868f
C690 B.n637 VSUBS 0.006868f
C691 B.n638 VSUBS 0.006868f
C692 B.n639 VSUBS 0.006868f
C693 B.n640 VSUBS 0.006868f
C694 B.n641 VSUBS 0.006868f
C695 B.n642 VSUBS 0.006868f
C696 B.n643 VSUBS 0.006868f
C697 B.n644 VSUBS 0.006868f
C698 B.n645 VSUBS 0.006868f
C699 B.n646 VSUBS 0.006868f
C700 B.n647 VSUBS 0.006868f
C701 B.n648 VSUBS 0.006868f
C702 B.n649 VSUBS 0.006868f
C703 B.n650 VSUBS 0.006868f
C704 B.n651 VSUBS 0.006868f
C705 B.n652 VSUBS 0.006868f
C706 B.n653 VSUBS 0.006868f
C707 B.n654 VSUBS 0.006868f
C708 B.n655 VSUBS 0.006868f
C709 B.n656 VSUBS 0.006868f
C710 B.n657 VSUBS 0.006868f
C711 B.n658 VSUBS 0.006868f
C712 B.n659 VSUBS 0.006868f
C713 B.n660 VSUBS 0.006868f
C714 B.n661 VSUBS 0.006868f
C715 B.n662 VSUBS 0.006868f
C716 B.n663 VSUBS 0.006868f
C717 B.n664 VSUBS 0.006868f
C718 B.n665 VSUBS 0.006868f
C719 B.n666 VSUBS 0.006868f
C720 B.n667 VSUBS 0.006868f
C721 B.n668 VSUBS 0.006868f
C722 B.n669 VSUBS 0.006868f
C723 B.n670 VSUBS 0.006868f
C724 B.n671 VSUBS 0.006868f
C725 B.n672 VSUBS 0.006868f
C726 B.n673 VSUBS 0.006868f
C727 B.n674 VSUBS 0.006868f
C728 B.n675 VSUBS 0.006868f
C729 B.n676 VSUBS 0.006868f
C730 B.n677 VSUBS 0.006868f
C731 B.n678 VSUBS 0.006868f
C732 B.n679 VSUBS 0.006868f
C733 B.n680 VSUBS 0.016032f
C734 B.n681 VSUBS 0.016032f
C735 B.n682 VSUBS 0.015481f
C736 B.n683 VSUBS 0.006868f
C737 B.n684 VSUBS 0.006868f
C738 B.n685 VSUBS 0.006868f
C739 B.n686 VSUBS 0.006868f
C740 B.n687 VSUBS 0.006868f
C741 B.n688 VSUBS 0.006868f
C742 B.n689 VSUBS 0.006868f
C743 B.n690 VSUBS 0.006868f
C744 B.n691 VSUBS 0.006868f
C745 B.n692 VSUBS 0.006868f
C746 B.n693 VSUBS 0.006868f
C747 B.n694 VSUBS 0.006868f
C748 B.n695 VSUBS 0.006868f
C749 B.n696 VSUBS 0.006868f
C750 B.n697 VSUBS 0.006868f
C751 B.n698 VSUBS 0.006868f
C752 B.n699 VSUBS 0.006868f
C753 B.n700 VSUBS 0.006868f
C754 B.n701 VSUBS 0.006868f
C755 B.n702 VSUBS 0.006868f
C756 B.n703 VSUBS 0.006868f
C757 B.n704 VSUBS 0.006868f
C758 B.n705 VSUBS 0.006868f
C759 B.n706 VSUBS 0.006868f
C760 B.n707 VSUBS 0.006868f
C761 B.n708 VSUBS 0.006868f
C762 B.n709 VSUBS 0.006868f
C763 B.n710 VSUBS 0.006868f
C764 B.n711 VSUBS 0.006868f
C765 B.n712 VSUBS 0.006868f
C766 B.n713 VSUBS 0.006868f
C767 B.n714 VSUBS 0.006868f
C768 B.n715 VSUBS 0.006868f
C769 B.n716 VSUBS 0.006868f
C770 B.n717 VSUBS 0.006868f
C771 B.n718 VSUBS 0.006868f
C772 B.n719 VSUBS 0.006868f
C773 B.n720 VSUBS 0.006868f
C774 B.n721 VSUBS 0.006868f
C775 B.n722 VSUBS 0.006868f
C776 B.n723 VSUBS 0.006868f
C777 B.n724 VSUBS 0.006868f
C778 B.n725 VSUBS 0.006868f
C779 B.n726 VSUBS 0.006868f
C780 B.n727 VSUBS 0.006868f
C781 B.n728 VSUBS 0.006868f
C782 B.n729 VSUBS 0.006868f
C783 B.n730 VSUBS 0.006868f
C784 B.n731 VSUBS 0.006868f
C785 B.n732 VSUBS 0.006868f
C786 B.n733 VSUBS 0.006868f
C787 B.n734 VSUBS 0.006868f
C788 B.n735 VSUBS 0.006868f
C789 B.n736 VSUBS 0.006868f
C790 B.n737 VSUBS 0.006868f
C791 B.n738 VSUBS 0.006868f
C792 B.n739 VSUBS 0.006868f
C793 B.n740 VSUBS 0.006868f
C794 B.n741 VSUBS 0.006868f
C795 B.n742 VSUBS 0.006868f
C796 B.n743 VSUBS 0.006868f
C797 B.n744 VSUBS 0.006868f
C798 B.n745 VSUBS 0.006868f
C799 B.n746 VSUBS 0.006868f
C800 B.n747 VSUBS 0.015552f
C801 VTAIL.n0 VSUBS 0.025743f
C802 VTAIL.n1 VSUBS 0.024174f
C803 VTAIL.n2 VSUBS 0.01299f
C804 VTAIL.n3 VSUBS 0.030704f
C805 VTAIL.n4 VSUBS 0.013754f
C806 VTAIL.n5 VSUBS 0.024174f
C807 VTAIL.n6 VSUBS 0.01299f
C808 VTAIL.n7 VSUBS 0.030704f
C809 VTAIL.n8 VSUBS 0.013754f
C810 VTAIL.n9 VSUBS 0.024174f
C811 VTAIL.n10 VSUBS 0.01299f
C812 VTAIL.n11 VSUBS 0.030704f
C813 VTAIL.n12 VSUBS 0.013754f
C814 VTAIL.n13 VSUBS 0.024174f
C815 VTAIL.n14 VSUBS 0.01299f
C816 VTAIL.n15 VSUBS 0.030704f
C817 VTAIL.n16 VSUBS 0.013754f
C818 VTAIL.n17 VSUBS 0.024174f
C819 VTAIL.n18 VSUBS 0.01299f
C820 VTAIL.n19 VSUBS 0.030704f
C821 VTAIL.n20 VSUBS 0.013754f
C822 VTAIL.n21 VSUBS 0.19836f
C823 VTAIL.t3 VSUBS 0.06622f
C824 VTAIL.n22 VSUBS 0.023028f
C825 VTAIL.n23 VSUBS 0.023097f
C826 VTAIL.n24 VSUBS 0.01299f
C827 VTAIL.n25 VSUBS 1.26506f
C828 VTAIL.n26 VSUBS 0.024174f
C829 VTAIL.n27 VSUBS 0.01299f
C830 VTAIL.n28 VSUBS 0.013754f
C831 VTAIL.n29 VSUBS 0.030704f
C832 VTAIL.n30 VSUBS 0.030704f
C833 VTAIL.n31 VSUBS 0.013754f
C834 VTAIL.n32 VSUBS 0.01299f
C835 VTAIL.n33 VSUBS 0.024174f
C836 VTAIL.n34 VSUBS 0.024174f
C837 VTAIL.n35 VSUBS 0.01299f
C838 VTAIL.n36 VSUBS 0.013754f
C839 VTAIL.n37 VSUBS 0.030704f
C840 VTAIL.n38 VSUBS 0.030704f
C841 VTAIL.n39 VSUBS 0.030704f
C842 VTAIL.n40 VSUBS 0.013754f
C843 VTAIL.n41 VSUBS 0.01299f
C844 VTAIL.n42 VSUBS 0.024174f
C845 VTAIL.n43 VSUBS 0.024174f
C846 VTAIL.n44 VSUBS 0.01299f
C847 VTAIL.n45 VSUBS 0.013372f
C848 VTAIL.n46 VSUBS 0.013372f
C849 VTAIL.n47 VSUBS 0.030704f
C850 VTAIL.n48 VSUBS 0.030704f
C851 VTAIL.n49 VSUBS 0.013754f
C852 VTAIL.n50 VSUBS 0.01299f
C853 VTAIL.n51 VSUBS 0.024174f
C854 VTAIL.n52 VSUBS 0.024174f
C855 VTAIL.n53 VSUBS 0.01299f
C856 VTAIL.n54 VSUBS 0.013754f
C857 VTAIL.n55 VSUBS 0.030704f
C858 VTAIL.n56 VSUBS 0.030704f
C859 VTAIL.n57 VSUBS 0.013754f
C860 VTAIL.n58 VSUBS 0.01299f
C861 VTAIL.n59 VSUBS 0.024174f
C862 VTAIL.n60 VSUBS 0.024174f
C863 VTAIL.n61 VSUBS 0.01299f
C864 VTAIL.n62 VSUBS 0.013754f
C865 VTAIL.n63 VSUBS 0.030704f
C866 VTAIL.n64 VSUBS 0.071542f
C867 VTAIL.n65 VSUBS 0.013754f
C868 VTAIL.n66 VSUBS 0.01299f
C869 VTAIL.n67 VSUBS 0.052244f
C870 VTAIL.n68 VSUBS 0.035739f
C871 VTAIL.n69 VSUBS 0.192013f
C872 VTAIL.n70 VSUBS 0.025743f
C873 VTAIL.n71 VSUBS 0.024174f
C874 VTAIL.n72 VSUBS 0.01299f
C875 VTAIL.n73 VSUBS 0.030704f
C876 VTAIL.n74 VSUBS 0.013754f
C877 VTAIL.n75 VSUBS 0.024174f
C878 VTAIL.n76 VSUBS 0.01299f
C879 VTAIL.n77 VSUBS 0.030704f
C880 VTAIL.n78 VSUBS 0.013754f
C881 VTAIL.n79 VSUBS 0.024174f
C882 VTAIL.n80 VSUBS 0.01299f
C883 VTAIL.n81 VSUBS 0.030704f
C884 VTAIL.n82 VSUBS 0.013754f
C885 VTAIL.n83 VSUBS 0.024174f
C886 VTAIL.n84 VSUBS 0.01299f
C887 VTAIL.n85 VSUBS 0.030704f
C888 VTAIL.n86 VSUBS 0.013754f
C889 VTAIL.n87 VSUBS 0.024174f
C890 VTAIL.n88 VSUBS 0.01299f
C891 VTAIL.n89 VSUBS 0.030704f
C892 VTAIL.n90 VSUBS 0.013754f
C893 VTAIL.n91 VSUBS 0.19836f
C894 VTAIL.t6 VSUBS 0.06622f
C895 VTAIL.n92 VSUBS 0.023028f
C896 VTAIL.n93 VSUBS 0.023097f
C897 VTAIL.n94 VSUBS 0.01299f
C898 VTAIL.n95 VSUBS 1.26506f
C899 VTAIL.n96 VSUBS 0.024174f
C900 VTAIL.n97 VSUBS 0.01299f
C901 VTAIL.n98 VSUBS 0.013754f
C902 VTAIL.n99 VSUBS 0.030704f
C903 VTAIL.n100 VSUBS 0.030704f
C904 VTAIL.n101 VSUBS 0.013754f
C905 VTAIL.n102 VSUBS 0.01299f
C906 VTAIL.n103 VSUBS 0.024174f
C907 VTAIL.n104 VSUBS 0.024174f
C908 VTAIL.n105 VSUBS 0.01299f
C909 VTAIL.n106 VSUBS 0.013754f
C910 VTAIL.n107 VSUBS 0.030704f
C911 VTAIL.n108 VSUBS 0.030704f
C912 VTAIL.n109 VSUBS 0.030704f
C913 VTAIL.n110 VSUBS 0.013754f
C914 VTAIL.n111 VSUBS 0.01299f
C915 VTAIL.n112 VSUBS 0.024174f
C916 VTAIL.n113 VSUBS 0.024174f
C917 VTAIL.n114 VSUBS 0.01299f
C918 VTAIL.n115 VSUBS 0.013372f
C919 VTAIL.n116 VSUBS 0.013372f
C920 VTAIL.n117 VSUBS 0.030704f
C921 VTAIL.n118 VSUBS 0.030704f
C922 VTAIL.n119 VSUBS 0.013754f
C923 VTAIL.n120 VSUBS 0.01299f
C924 VTAIL.n121 VSUBS 0.024174f
C925 VTAIL.n122 VSUBS 0.024174f
C926 VTAIL.n123 VSUBS 0.01299f
C927 VTAIL.n124 VSUBS 0.013754f
C928 VTAIL.n125 VSUBS 0.030704f
C929 VTAIL.n126 VSUBS 0.030704f
C930 VTAIL.n127 VSUBS 0.013754f
C931 VTAIL.n128 VSUBS 0.01299f
C932 VTAIL.n129 VSUBS 0.024174f
C933 VTAIL.n130 VSUBS 0.024174f
C934 VTAIL.n131 VSUBS 0.01299f
C935 VTAIL.n132 VSUBS 0.013754f
C936 VTAIL.n133 VSUBS 0.030704f
C937 VTAIL.n134 VSUBS 0.071542f
C938 VTAIL.n135 VSUBS 0.013754f
C939 VTAIL.n136 VSUBS 0.01299f
C940 VTAIL.n137 VSUBS 0.052244f
C941 VTAIL.n138 VSUBS 0.035739f
C942 VTAIL.n139 VSUBS 0.319764f
C943 VTAIL.n140 VSUBS 0.025743f
C944 VTAIL.n141 VSUBS 0.024174f
C945 VTAIL.n142 VSUBS 0.01299f
C946 VTAIL.n143 VSUBS 0.030704f
C947 VTAIL.n144 VSUBS 0.013754f
C948 VTAIL.n145 VSUBS 0.024174f
C949 VTAIL.n146 VSUBS 0.01299f
C950 VTAIL.n147 VSUBS 0.030704f
C951 VTAIL.n148 VSUBS 0.013754f
C952 VTAIL.n149 VSUBS 0.024174f
C953 VTAIL.n150 VSUBS 0.01299f
C954 VTAIL.n151 VSUBS 0.030704f
C955 VTAIL.n152 VSUBS 0.013754f
C956 VTAIL.n153 VSUBS 0.024174f
C957 VTAIL.n154 VSUBS 0.01299f
C958 VTAIL.n155 VSUBS 0.030704f
C959 VTAIL.n156 VSUBS 0.013754f
C960 VTAIL.n157 VSUBS 0.024174f
C961 VTAIL.n158 VSUBS 0.01299f
C962 VTAIL.n159 VSUBS 0.030704f
C963 VTAIL.n160 VSUBS 0.013754f
C964 VTAIL.n161 VSUBS 0.19836f
C965 VTAIL.t5 VSUBS 0.06622f
C966 VTAIL.n162 VSUBS 0.023028f
C967 VTAIL.n163 VSUBS 0.023097f
C968 VTAIL.n164 VSUBS 0.01299f
C969 VTAIL.n165 VSUBS 1.26506f
C970 VTAIL.n166 VSUBS 0.024174f
C971 VTAIL.n167 VSUBS 0.01299f
C972 VTAIL.n168 VSUBS 0.013754f
C973 VTAIL.n169 VSUBS 0.030704f
C974 VTAIL.n170 VSUBS 0.030704f
C975 VTAIL.n171 VSUBS 0.013754f
C976 VTAIL.n172 VSUBS 0.01299f
C977 VTAIL.n173 VSUBS 0.024174f
C978 VTAIL.n174 VSUBS 0.024174f
C979 VTAIL.n175 VSUBS 0.01299f
C980 VTAIL.n176 VSUBS 0.013754f
C981 VTAIL.n177 VSUBS 0.030704f
C982 VTAIL.n178 VSUBS 0.030704f
C983 VTAIL.n179 VSUBS 0.030704f
C984 VTAIL.n180 VSUBS 0.013754f
C985 VTAIL.n181 VSUBS 0.01299f
C986 VTAIL.n182 VSUBS 0.024174f
C987 VTAIL.n183 VSUBS 0.024174f
C988 VTAIL.n184 VSUBS 0.01299f
C989 VTAIL.n185 VSUBS 0.013372f
C990 VTAIL.n186 VSUBS 0.013372f
C991 VTAIL.n187 VSUBS 0.030704f
C992 VTAIL.n188 VSUBS 0.030704f
C993 VTAIL.n189 VSUBS 0.013754f
C994 VTAIL.n190 VSUBS 0.01299f
C995 VTAIL.n191 VSUBS 0.024174f
C996 VTAIL.n192 VSUBS 0.024174f
C997 VTAIL.n193 VSUBS 0.01299f
C998 VTAIL.n194 VSUBS 0.013754f
C999 VTAIL.n195 VSUBS 0.030704f
C1000 VTAIL.n196 VSUBS 0.030704f
C1001 VTAIL.n197 VSUBS 0.013754f
C1002 VTAIL.n198 VSUBS 0.01299f
C1003 VTAIL.n199 VSUBS 0.024174f
C1004 VTAIL.n200 VSUBS 0.024174f
C1005 VTAIL.n201 VSUBS 0.01299f
C1006 VTAIL.n202 VSUBS 0.013754f
C1007 VTAIL.n203 VSUBS 0.030704f
C1008 VTAIL.n204 VSUBS 0.071542f
C1009 VTAIL.n205 VSUBS 0.013754f
C1010 VTAIL.n206 VSUBS 0.01299f
C1011 VTAIL.n207 VSUBS 0.052244f
C1012 VTAIL.n208 VSUBS 0.035739f
C1013 VTAIL.n209 VSUBS 1.73092f
C1014 VTAIL.n210 VSUBS 0.025743f
C1015 VTAIL.n211 VSUBS 0.024174f
C1016 VTAIL.n212 VSUBS 0.01299f
C1017 VTAIL.n213 VSUBS 0.030704f
C1018 VTAIL.n214 VSUBS 0.013754f
C1019 VTAIL.n215 VSUBS 0.024174f
C1020 VTAIL.n216 VSUBS 0.01299f
C1021 VTAIL.n217 VSUBS 0.030704f
C1022 VTAIL.n218 VSUBS 0.013754f
C1023 VTAIL.n219 VSUBS 0.024174f
C1024 VTAIL.n220 VSUBS 0.01299f
C1025 VTAIL.n221 VSUBS 0.030704f
C1026 VTAIL.n222 VSUBS 0.013754f
C1027 VTAIL.n223 VSUBS 0.024174f
C1028 VTAIL.n224 VSUBS 0.01299f
C1029 VTAIL.n225 VSUBS 0.030704f
C1030 VTAIL.n226 VSUBS 0.030704f
C1031 VTAIL.n227 VSUBS 0.013754f
C1032 VTAIL.n228 VSUBS 0.024174f
C1033 VTAIL.n229 VSUBS 0.01299f
C1034 VTAIL.n230 VSUBS 0.030704f
C1035 VTAIL.n231 VSUBS 0.013754f
C1036 VTAIL.n232 VSUBS 0.19836f
C1037 VTAIL.t1 VSUBS 0.06622f
C1038 VTAIL.n233 VSUBS 0.023028f
C1039 VTAIL.n234 VSUBS 0.023097f
C1040 VTAIL.n235 VSUBS 0.01299f
C1041 VTAIL.n236 VSUBS 1.26506f
C1042 VTAIL.n237 VSUBS 0.024174f
C1043 VTAIL.n238 VSUBS 0.01299f
C1044 VTAIL.n239 VSUBS 0.013754f
C1045 VTAIL.n240 VSUBS 0.030704f
C1046 VTAIL.n241 VSUBS 0.030704f
C1047 VTAIL.n242 VSUBS 0.013754f
C1048 VTAIL.n243 VSUBS 0.01299f
C1049 VTAIL.n244 VSUBS 0.024174f
C1050 VTAIL.n245 VSUBS 0.024174f
C1051 VTAIL.n246 VSUBS 0.01299f
C1052 VTAIL.n247 VSUBS 0.013754f
C1053 VTAIL.n248 VSUBS 0.030704f
C1054 VTAIL.n249 VSUBS 0.030704f
C1055 VTAIL.n250 VSUBS 0.013754f
C1056 VTAIL.n251 VSUBS 0.01299f
C1057 VTAIL.n252 VSUBS 0.024174f
C1058 VTAIL.n253 VSUBS 0.024174f
C1059 VTAIL.n254 VSUBS 0.01299f
C1060 VTAIL.n255 VSUBS 0.013372f
C1061 VTAIL.n256 VSUBS 0.013372f
C1062 VTAIL.n257 VSUBS 0.030704f
C1063 VTAIL.n258 VSUBS 0.030704f
C1064 VTAIL.n259 VSUBS 0.013754f
C1065 VTAIL.n260 VSUBS 0.01299f
C1066 VTAIL.n261 VSUBS 0.024174f
C1067 VTAIL.n262 VSUBS 0.024174f
C1068 VTAIL.n263 VSUBS 0.01299f
C1069 VTAIL.n264 VSUBS 0.013754f
C1070 VTAIL.n265 VSUBS 0.030704f
C1071 VTAIL.n266 VSUBS 0.030704f
C1072 VTAIL.n267 VSUBS 0.013754f
C1073 VTAIL.n268 VSUBS 0.01299f
C1074 VTAIL.n269 VSUBS 0.024174f
C1075 VTAIL.n270 VSUBS 0.024174f
C1076 VTAIL.n271 VSUBS 0.01299f
C1077 VTAIL.n272 VSUBS 0.013754f
C1078 VTAIL.n273 VSUBS 0.030704f
C1079 VTAIL.n274 VSUBS 0.071542f
C1080 VTAIL.n275 VSUBS 0.013754f
C1081 VTAIL.n276 VSUBS 0.01299f
C1082 VTAIL.n277 VSUBS 0.052244f
C1083 VTAIL.n278 VSUBS 0.035739f
C1084 VTAIL.n279 VSUBS 1.73092f
C1085 VTAIL.n280 VSUBS 0.025743f
C1086 VTAIL.n281 VSUBS 0.024174f
C1087 VTAIL.n282 VSUBS 0.01299f
C1088 VTAIL.n283 VSUBS 0.030704f
C1089 VTAIL.n284 VSUBS 0.013754f
C1090 VTAIL.n285 VSUBS 0.024174f
C1091 VTAIL.n286 VSUBS 0.01299f
C1092 VTAIL.n287 VSUBS 0.030704f
C1093 VTAIL.n288 VSUBS 0.013754f
C1094 VTAIL.n289 VSUBS 0.024174f
C1095 VTAIL.n290 VSUBS 0.01299f
C1096 VTAIL.n291 VSUBS 0.030704f
C1097 VTAIL.n292 VSUBS 0.013754f
C1098 VTAIL.n293 VSUBS 0.024174f
C1099 VTAIL.n294 VSUBS 0.01299f
C1100 VTAIL.n295 VSUBS 0.030704f
C1101 VTAIL.n296 VSUBS 0.030704f
C1102 VTAIL.n297 VSUBS 0.013754f
C1103 VTAIL.n298 VSUBS 0.024174f
C1104 VTAIL.n299 VSUBS 0.01299f
C1105 VTAIL.n300 VSUBS 0.030704f
C1106 VTAIL.n301 VSUBS 0.013754f
C1107 VTAIL.n302 VSUBS 0.19836f
C1108 VTAIL.t2 VSUBS 0.06622f
C1109 VTAIL.n303 VSUBS 0.023028f
C1110 VTAIL.n304 VSUBS 0.023097f
C1111 VTAIL.n305 VSUBS 0.01299f
C1112 VTAIL.n306 VSUBS 1.26506f
C1113 VTAIL.n307 VSUBS 0.024174f
C1114 VTAIL.n308 VSUBS 0.01299f
C1115 VTAIL.n309 VSUBS 0.013754f
C1116 VTAIL.n310 VSUBS 0.030704f
C1117 VTAIL.n311 VSUBS 0.030704f
C1118 VTAIL.n312 VSUBS 0.013754f
C1119 VTAIL.n313 VSUBS 0.01299f
C1120 VTAIL.n314 VSUBS 0.024174f
C1121 VTAIL.n315 VSUBS 0.024174f
C1122 VTAIL.n316 VSUBS 0.01299f
C1123 VTAIL.n317 VSUBS 0.013754f
C1124 VTAIL.n318 VSUBS 0.030704f
C1125 VTAIL.n319 VSUBS 0.030704f
C1126 VTAIL.n320 VSUBS 0.013754f
C1127 VTAIL.n321 VSUBS 0.01299f
C1128 VTAIL.n322 VSUBS 0.024174f
C1129 VTAIL.n323 VSUBS 0.024174f
C1130 VTAIL.n324 VSUBS 0.01299f
C1131 VTAIL.n325 VSUBS 0.013372f
C1132 VTAIL.n326 VSUBS 0.013372f
C1133 VTAIL.n327 VSUBS 0.030704f
C1134 VTAIL.n328 VSUBS 0.030704f
C1135 VTAIL.n329 VSUBS 0.013754f
C1136 VTAIL.n330 VSUBS 0.01299f
C1137 VTAIL.n331 VSUBS 0.024174f
C1138 VTAIL.n332 VSUBS 0.024174f
C1139 VTAIL.n333 VSUBS 0.01299f
C1140 VTAIL.n334 VSUBS 0.013754f
C1141 VTAIL.n335 VSUBS 0.030704f
C1142 VTAIL.n336 VSUBS 0.030704f
C1143 VTAIL.n337 VSUBS 0.013754f
C1144 VTAIL.n338 VSUBS 0.01299f
C1145 VTAIL.n339 VSUBS 0.024174f
C1146 VTAIL.n340 VSUBS 0.024174f
C1147 VTAIL.n341 VSUBS 0.01299f
C1148 VTAIL.n342 VSUBS 0.013754f
C1149 VTAIL.n343 VSUBS 0.030704f
C1150 VTAIL.n344 VSUBS 0.071542f
C1151 VTAIL.n345 VSUBS 0.013754f
C1152 VTAIL.n346 VSUBS 0.01299f
C1153 VTAIL.n347 VSUBS 0.052244f
C1154 VTAIL.n348 VSUBS 0.035739f
C1155 VTAIL.n349 VSUBS 0.319764f
C1156 VTAIL.n350 VSUBS 0.025743f
C1157 VTAIL.n351 VSUBS 0.024174f
C1158 VTAIL.n352 VSUBS 0.01299f
C1159 VTAIL.n353 VSUBS 0.030704f
C1160 VTAIL.n354 VSUBS 0.013754f
C1161 VTAIL.n355 VSUBS 0.024174f
C1162 VTAIL.n356 VSUBS 0.01299f
C1163 VTAIL.n357 VSUBS 0.030704f
C1164 VTAIL.n358 VSUBS 0.013754f
C1165 VTAIL.n359 VSUBS 0.024174f
C1166 VTAIL.n360 VSUBS 0.01299f
C1167 VTAIL.n361 VSUBS 0.030704f
C1168 VTAIL.n362 VSUBS 0.013754f
C1169 VTAIL.n363 VSUBS 0.024174f
C1170 VTAIL.n364 VSUBS 0.01299f
C1171 VTAIL.n365 VSUBS 0.030704f
C1172 VTAIL.n366 VSUBS 0.030704f
C1173 VTAIL.n367 VSUBS 0.013754f
C1174 VTAIL.n368 VSUBS 0.024174f
C1175 VTAIL.n369 VSUBS 0.01299f
C1176 VTAIL.n370 VSUBS 0.030704f
C1177 VTAIL.n371 VSUBS 0.013754f
C1178 VTAIL.n372 VSUBS 0.19836f
C1179 VTAIL.t7 VSUBS 0.06622f
C1180 VTAIL.n373 VSUBS 0.023028f
C1181 VTAIL.n374 VSUBS 0.023097f
C1182 VTAIL.n375 VSUBS 0.01299f
C1183 VTAIL.n376 VSUBS 1.26506f
C1184 VTAIL.n377 VSUBS 0.024174f
C1185 VTAIL.n378 VSUBS 0.01299f
C1186 VTAIL.n379 VSUBS 0.013754f
C1187 VTAIL.n380 VSUBS 0.030704f
C1188 VTAIL.n381 VSUBS 0.030704f
C1189 VTAIL.n382 VSUBS 0.013754f
C1190 VTAIL.n383 VSUBS 0.01299f
C1191 VTAIL.n384 VSUBS 0.024174f
C1192 VTAIL.n385 VSUBS 0.024174f
C1193 VTAIL.n386 VSUBS 0.01299f
C1194 VTAIL.n387 VSUBS 0.013754f
C1195 VTAIL.n388 VSUBS 0.030704f
C1196 VTAIL.n389 VSUBS 0.030704f
C1197 VTAIL.n390 VSUBS 0.013754f
C1198 VTAIL.n391 VSUBS 0.01299f
C1199 VTAIL.n392 VSUBS 0.024174f
C1200 VTAIL.n393 VSUBS 0.024174f
C1201 VTAIL.n394 VSUBS 0.01299f
C1202 VTAIL.n395 VSUBS 0.013372f
C1203 VTAIL.n396 VSUBS 0.013372f
C1204 VTAIL.n397 VSUBS 0.030704f
C1205 VTAIL.n398 VSUBS 0.030704f
C1206 VTAIL.n399 VSUBS 0.013754f
C1207 VTAIL.n400 VSUBS 0.01299f
C1208 VTAIL.n401 VSUBS 0.024174f
C1209 VTAIL.n402 VSUBS 0.024174f
C1210 VTAIL.n403 VSUBS 0.01299f
C1211 VTAIL.n404 VSUBS 0.013754f
C1212 VTAIL.n405 VSUBS 0.030704f
C1213 VTAIL.n406 VSUBS 0.030704f
C1214 VTAIL.n407 VSUBS 0.013754f
C1215 VTAIL.n408 VSUBS 0.01299f
C1216 VTAIL.n409 VSUBS 0.024174f
C1217 VTAIL.n410 VSUBS 0.024174f
C1218 VTAIL.n411 VSUBS 0.01299f
C1219 VTAIL.n412 VSUBS 0.013754f
C1220 VTAIL.n413 VSUBS 0.030704f
C1221 VTAIL.n414 VSUBS 0.071542f
C1222 VTAIL.n415 VSUBS 0.013754f
C1223 VTAIL.n416 VSUBS 0.01299f
C1224 VTAIL.n417 VSUBS 0.052244f
C1225 VTAIL.n418 VSUBS 0.035739f
C1226 VTAIL.n419 VSUBS 0.319764f
C1227 VTAIL.n420 VSUBS 0.025743f
C1228 VTAIL.n421 VSUBS 0.024174f
C1229 VTAIL.n422 VSUBS 0.01299f
C1230 VTAIL.n423 VSUBS 0.030704f
C1231 VTAIL.n424 VSUBS 0.013754f
C1232 VTAIL.n425 VSUBS 0.024174f
C1233 VTAIL.n426 VSUBS 0.01299f
C1234 VTAIL.n427 VSUBS 0.030704f
C1235 VTAIL.n428 VSUBS 0.013754f
C1236 VTAIL.n429 VSUBS 0.024174f
C1237 VTAIL.n430 VSUBS 0.01299f
C1238 VTAIL.n431 VSUBS 0.030704f
C1239 VTAIL.n432 VSUBS 0.013754f
C1240 VTAIL.n433 VSUBS 0.024174f
C1241 VTAIL.n434 VSUBS 0.01299f
C1242 VTAIL.n435 VSUBS 0.030704f
C1243 VTAIL.n436 VSUBS 0.030704f
C1244 VTAIL.n437 VSUBS 0.013754f
C1245 VTAIL.n438 VSUBS 0.024174f
C1246 VTAIL.n439 VSUBS 0.01299f
C1247 VTAIL.n440 VSUBS 0.030704f
C1248 VTAIL.n441 VSUBS 0.013754f
C1249 VTAIL.n442 VSUBS 0.19836f
C1250 VTAIL.t4 VSUBS 0.06622f
C1251 VTAIL.n443 VSUBS 0.023028f
C1252 VTAIL.n444 VSUBS 0.023097f
C1253 VTAIL.n445 VSUBS 0.01299f
C1254 VTAIL.n446 VSUBS 1.26506f
C1255 VTAIL.n447 VSUBS 0.024174f
C1256 VTAIL.n448 VSUBS 0.01299f
C1257 VTAIL.n449 VSUBS 0.013754f
C1258 VTAIL.n450 VSUBS 0.030704f
C1259 VTAIL.n451 VSUBS 0.030704f
C1260 VTAIL.n452 VSUBS 0.013754f
C1261 VTAIL.n453 VSUBS 0.01299f
C1262 VTAIL.n454 VSUBS 0.024174f
C1263 VTAIL.n455 VSUBS 0.024174f
C1264 VTAIL.n456 VSUBS 0.01299f
C1265 VTAIL.n457 VSUBS 0.013754f
C1266 VTAIL.n458 VSUBS 0.030704f
C1267 VTAIL.n459 VSUBS 0.030704f
C1268 VTAIL.n460 VSUBS 0.013754f
C1269 VTAIL.n461 VSUBS 0.01299f
C1270 VTAIL.n462 VSUBS 0.024174f
C1271 VTAIL.n463 VSUBS 0.024174f
C1272 VTAIL.n464 VSUBS 0.01299f
C1273 VTAIL.n465 VSUBS 0.013372f
C1274 VTAIL.n466 VSUBS 0.013372f
C1275 VTAIL.n467 VSUBS 0.030704f
C1276 VTAIL.n468 VSUBS 0.030704f
C1277 VTAIL.n469 VSUBS 0.013754f
C1278 VTAIL.n470 VSUBS 0.01299f
C1279 VTAIL.n471 VSUBS 0.024174f
C1280 VTAIL.n472 VSUBS 0.024174f
C1281 VTAIL.n473 VSUBS 0.01299f
C1282 VTAIL.n474 VSUBS 0.013754f
C1283 VTAIL.n475 VSUBS 0.030704f
C1284 VTAIL.n476 VSUBS 0.030704f
C1285 VTAIL.n477 VSUBS 0.013754f
C1286 VTAIL.n478 VSUBS 0.01299f
C1287 VTAIL.n479 VSUBS 0.024174f
C1288 VTAIL.n480 VSUBS 0.024174f
C1289 VTAIL.n481 VSUBS 0.01299f
C1290 VTAIL.n482 VSUBS 0.013754f
C1291 VTAIL.n483 VSUBS 0.030704f
C1292 VTAIL.n484 VSUBS 0.071542f
C1293 VTAIL.n485 VSUBS 0.013754f
C1294 VTAIL.n486 VSUBS 0.01299f
C1295 VTAIL.n487 VSUBS 0.052244f
C1296 VTAIL.n488 VSUBS 0.035739f
C1297 VTAIL.n489 VSUBS 1.73092f
C1298 VTAIL.n490 VSUBS 0.025743f
C1299 VTAIL.n491 VSUBS 0.024174f
C1300 VTAIL.n492 VSUBS 0.01299f
C1301 VTAIL.n493 VSUBS 0.030704f
C1302 VTAIL.n494 VSUBS 0.013754f
C1303 VTAIL.n495 VSUBS 0.024174f
C1304 VTAIL.n496 VSUBS 0.01299f
C1305 VTAIL.n497 VSUBS 0.030704f
C1306 VTAIL.n498 VSUBS 0.013754f
C1307 VTAIL.n499 VSUBS 0.024174f
C1308 VTAIL.n500 VSUBS 0.01299f
C1309 VTAIL.n501 VSUBS 0.030704f
C1310 VTAIL.n502 VSUBS 0.013754f
C1311 VTAIL.n503 VSUBS 0.024174f
C1312 VTAIL.n504 VSUBS 0.01299f
C1313 VTAIL.n505 VSUBS 0.030704f
C1314 VTAIL.n506 VSUBS 0.013754f
C1315 VTAIL.n507 VSUBS 0.024174f
C1316 VTAIL.n508 VSUBS 0.01299f
C1317 VTAIL.n509 VSUBS 0.030704f
C1318 VTAIL.n510 VSUBS 0.013754f
C1319 VTAIL.n511 VSUBS 0.19836f
C1320 VTAIL.t0 VSUBS 0.06622f
C1321 VTAIL.n512 VSUBS 0.023028f
C1322 VTAIL.n513 VSUBS 0.023097f
C1323 VTAIL.n514 VSUBS 0.01299f
C1324 VTAIL.n515 VSUBS 1.26506f
C1325 VTAIL.n516 VSUBS 0.024174f
C1326 VTAIL.n517 VSUBS 0.01299f
C1327 VTAIL.n518 VSUBS 0.013754f
C1328 VTAIL.n519 VSUBS 0.030704f
C1329 VTAIL.n520 VSUBS 0.030704f
C1330 VTAIL.n521 VSUBS 0.013754f
C1331 VTAIL.n522 VSUBS 0.01299f
C1332 VTAIL.n523 VSUBS 0.024174f
C1333 VTAIL.n524 VSUBS 0.024174f
C1334 VTAIL.n525 VSUBS 0.01299f
C1335 VTAIL.n526 VSUBS 0.013754f
C1336 VTAIL.n527 VSUBS 0.030704f
C1337 VTAIL.n528 VSUBS 0.030704f
C1338 VTAIL.n529 VSUBS 0.030704f
C1339 VTAIL.n530 VSUBS 0.013754f
C1340 VTAIL.n531 VSUBS 0.01299f
C1341 VTAIL.n532 VSUBS 0.024174f
C1342 VTAIL.n533 VSUBS 0.024174f
C1343 VTAIL.n534 VSUBS 0.01299f
C1344 VTAIL.n535 VSUBS 0.013372f
C1345 VTAIL.n536 VSUBS 0.013372f
C1346 VTAIL.n537 VSUBS 0.030704f
C1347 VTAIL.n538 VSUBS 0.030704f
C1348 VTAIL.n539 VSUBS 0.013754f
C1349 VTAIL.n540 VSUBS 0.01299f
C1350 VTAIL.n541 VSUBS 0.024174f
C1351 VTAIL.n542 VSUBS 0.024174f
C1352 VTAIL.n543 VSUBS 0.01299f
C1353 VTAIL.n544 VSUBS 0.013754f
C1354 VTAIL.n545 VSUBS 0.030704f
C1355 VTAIL.n546 VSUBS 0.030704f
C1356 VTAIL.n547 VSUBS 0.013754f
C1357 VTAIL.n548 VSUBS 0.01299f
C1358 VTAIL.n549 VSUBS 0.024174f
C1359 VTAIL.n550 VSUBS 0.024174f
C1360 VTAIL.n551 VSUBS 0.01299f
C1361 VTAIL.n552 VSUBS 0.013754f
C1362 VTAIL.n553 VSUBS 0.030704f
C1363 VTAIL.n554 VSUBS 0.071542f
C1364 VTAIL.n555 VSUBS 0.013754f
C1365 VTAIL.n556 VSUBS 0.01299f
C1366 VTAIL.n557 VSUBS 0.052244f
C1367 VTAIL.n558 VSUBS 0.035739f
C1368 VTAIL.n559 VSUBS 1.5941f
C1369 VDD1.t0 VSUBS 0.275964f
C1370 VDD1.t3 VSUBS 0.275964f
C1371 VDD1.n0 VSUBS 2.16568f
C1372 VDD1.t2 VSUBS 0.275964f
C1373 VDD1.t1 VSUBS 0.275964f
C1374 VDD1.n1 VSUBS 3.01964f
C1375 VP.t1 VSUBS 3.81847f
C1376 VP.n0 VSUBS 1.45738f
C1377 VP.n1 VSUBS 0.030446f
C1378 VP.n2 VSUBS 0.044446f
C1379 VP.n3 VSUBS 0.030446f
C1380 VP.n4 VSUBS 0.041056f
C1381 VP.t0 VSUBS 4.27813f
C1382 VP.t3 VSUBS 4.26254f
C1383 VP.n5 VSUBS 4.52483f
C1384 VP.t2 VSUBS 3.81847f
C1385 VP.n6 VSUBS 1.45738f
C1386 VP.n7 VSUBS 1.85447f
C1387 VP.n8 VSUBS 0.04914f
C1388 VP.n9 VSUBS 0.030446f
C1389 VP.n10 VSUBS 0.056745f
C1390 VP.n11 VSUBS 0.056745f
C1391 VP.n12 VSUBS 0.044446f
C1392 VP.n13 VSUBS 0.030446f
C1393 VP.n14 VSUBS 0.030446f
C1394 VP.n15 VSUBS 0.030446f
C1395 VP.n16 VSUBS 0.056745f
C1396 VP.n17 VSUBS 0.056745f
C1397 VP.n18 VSUBS 0.041056f
C1398 VP.n19 VSUBS 0.04914f
C1399 VP.n20 VSUBS 0.082484f
.ends

