* NGSPICE file created from diff_pair_sample_0912.ext - technology: sky130A

.subckt diff_pair_sample_0912 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t11 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.3315 ps=2.48 w=0.85 l=1.79
X1 VDD2.t4 VN.t1 VTAIL.t8 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0.14025 ps=1.18 w=0.85 l=1.79
X2 B.t11 B.t9 B.t10 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0 ps=0 w=0.85 l=1.79
X3 VDD1.t5 VP.t0 VTAIL.t4 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.3315 ps=2.48 w=0.85 l=1.79
X4 B.t8 B.t6 B.t7 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0 ps=0 w=0.85 l=1.79
X5 VDD1.t4 VP.t1 VTAIL.t5 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0.14025 ps=1.18 w=0.85 l=1.79
X6 VDD2.t3 VN.t2 VTAIL.t9 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.3315 ps=2.48 w=0.85 l=1.79
X7 VDD2.t2 VN.t3 VTAIL.t10 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0.14025 ps=1.18 w=0.85 l=1.79
X8 VTAIL.t7 VN.t4 VDD2.t1 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.14025 ps=1.18 w=0.85 l=1.79
X9 VDD1.t3 VP.t2 VTAIL.t1 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0.14025 ps=1.18 w=0.85 l=1.79
X10 VTAIL.t6 VN.t5 VDD2.t0 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.14025 ps=1.18 w=0.85 l=1.79
X11 VTAIL.t2 VP.t3 VDD1.t2 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.14025 ps=1.18 w=0.85 l=1.79
X12 VDD1.t1 VP.t4 VTAIL.t3 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.3315 ps=2.48 w=0.85 l=1.79
X13 VTAIL.t0 VP.t5 VDD1.t0 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.14025 pd=1.18 as=0.14025 ps=1.18 w=0.85 l=1.79
X14 B.t5 B.t3 B.t4 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0 ps=0 w=0.85 l=1.79
X15 B.t2 B.t0 B.t1 w_n2666_n1138# sky130_fd_pr__pfet_01v8 ad=0.3315 pd=2.48 as=0 ps=0 w=0.85 l=1.79
R0 VN.n11 VN.n10 179.895
R1 VN.n23 VN.n22 179.895
R2 VN.n21 VN.n12 161.3
R3 VN.n20 VN.n19 161.3
R4 VN.n18 VN.n13 161.3
R5 VN.n17 VN.n16 161.3
R6 VN.n9 VN.n0 161.3
R7 VN.n8 VN.n7 161.3
R8 VN.n6 VN.n1 161.3
R9 VN.n5 VN.n4 161.3
R10 VN.n2 VN.t1 47.3648
R11 VN.n14 VN.t2 47.3648
R12 VN.n8 VN.n1 46.321
R13 VN.n20 VN.n13 46.321
R14 VN.n15 VN.n14 44.4801
R15 VN.n3 VN.n2 44.4801
R16 VN VN.n23 37.366
R17 VN.n4 VN.n1 34.6658
R18 VN.n16 VN.n13 34.6658
R19 VN.n4 VN.n3 24.4675
R20 VN.n9 VN.n8 24.4675
R21 VN.n16 VN.n15 24.4675
R22 VN.n21 VN.n20 24.4675
R23 VN.n17 VN.n14 12.138
R24 VN.n5 VN.n2 12.138
R25 VN.n3 VN.t5 11.4446
R26 VN.n10 VN.t0 11.4446
R27 VN.n15 VN.t4 11.4446
R28 VN.n22 VN.t3 11.4446
R29 VN.n10 VN.n9 5.87258
R30 VN.n22 VN.n21 5.87258
R31 VN.n23 VN.n12 0.189894
R32 VN.n19 VN.n12 0.189894
R33 VN.n19 VN.n18 0.189894
R34 VN.n18 VN.n17 0.189894
R35 VN.n6 VN.n5 0.189894
R36 VN.n7 VN.n6 0.189894
R37 VN.n7 VN.n0 0.189894
R38 VN.n11 VN.n0 0.189894
R39 VN VN.n11 0.0516364
R40 VTAIL.n10 VTAIL.t3 658.787
R41 VTAIL.n7 VTAIL.t9 658.787
R42 VTAIL.n11 VTAIL.t11 658.785
R43 VTAIL.n2 VTAIL.t4 658.785
R44 VTAIL.n9 VTAIL.n8 620.544
R45 VTAIL.n6 VTAIL.n5 620.544
R46 VTAIL.n1 VTAIL.n0 620.544
R47 VTAIL.n4 VTAIL.n3 620.544
R48 VTAIL.n0 VTAIL.t8 38.2417
R49 VTAIL.n0 VTAIL.t6 38.2417
R50 VTAIL.n3 VTAIL.t5 38.2417
R51 VTAIL.n3 VTAIL.t2 38.2417
R52 VTAIL.n8 VTAIL.t1 38.2417
R53 VTAIL.n8 VTAIL.t0 38.2417
R54 VTAIL.n5 VTAIL.t10 38.2417
R55 VTAIL.n5 VTAIL.t7 38.2417
R56 VTAIL.n6 VTAIL.n4 16.7548
R57 VTAIL.n11 VTAIL.n10 14.9272
R58 VTAIL.n7 VTAIL.n6 1.82809
R59 VTAIL.n10 VTAIL.n9 1.82809
R60 VTAIL.n4 VTAIL.n2 1.82809
R61 VTAIL.n9 VTAIL.n7 1.38412
R62 VTAIL.n2 VTAIL.n1 1.38412
R63 VTAIL VTAIL.n11 1.313
R64 VTAIL VTAIL.n1 0.515586
R65 VDD2.n1 VDD2.t4 676.779
R66 VDD2.n2 VDD2.t2 675.465
R67 VDD2.n1 VDD2.n0 637.625
R68 VDD2 VDD2.n3 637.622
R69 VDD2.n3 VDD2.t1 38.2417
R70 VDD2.n3 VDD2.t3 38.2417
R71 VDD2.n0 VDD2.t0 38.2417
R72 VDD2.n0 VDD2.t5 38.2417
R73 VDD2.n2 VDD2.n1 30.3877
R74 VDD2 VDD2.n2 1.42938
R75 B.n74 B.t2 690.538
R76 B.n82 B.t8 690.538
R77 B.n24 B.t10 690.538
R78 B.n30 B.t4 690.538
R79 B.n75 B.t1 649.423
R80 B.n83 B.t7 649.423
R81 B.n25 B.t11 649.423
R82 B.n31 B.t5 649.423
R83 B.n295 B.n294 585
R84 B.n296 B.n35 585
R85 B.n298 B.n297 585
R86 B.n299 B.n34 585
R87 B.n301 B.n300 585
R88 B.n302 B.n33 585
R89 B.n304 B.n303 585
R90 B.n305 B.n32 585
R91 B.n307 B.n306 585
R92 B.n309 B.n29 585
R93 B.n311 B.n310 585
R94 B.n312 B.n28 585
R95 B.n314 B.n313 585
R96 B.n315 B.n27 585
R97 B.n317 B.n316 585
R98 B.n318 B.n26 585
R99 B.n320 B.n319 585
R100 B.n321 B.n23 585
R101 B.n324 B.n323 585
R102 B.n325 B.n22 585
R103 B.n327 B.n326 585
R104 B.n328 B.n21 585
R105 B.n330 B.n329 585
R106 B.n331 B.n20 585
R107 B.n333 B.n332 585
R108 B.n334 B.n19 585
R109 B.n336 B.n335 585
R110 B.n293 B.n36 585
R111 B.n292 B.n291 585
R112 B.n290 B.n37 585
R113 B.n289 B.n288 585
R114 B.n287 B.n38 585
R115 B.n286 B.n285 585
R116 B.n284 B.n39 585
R117 B.n283 B.n282 585
R118 B.n281 B.n40 585
R119 B.n280 B.n279 585
R120 B.n278 B.n41 585
R121 B.n277 B.n276 585
R122 B.n275 B.n42 585
R123 B.n274 B.n273 585
R124 B.n272 B.n43 585
R125 B.n271 B.n270 585
R126 B.n269 B.n44 585
R127 B.n268 B.n267 585
R128 B.n266 B.n45 585
R129 B.n265 B.n264 585
R130 B.n263 B.n46 585
R131 B.n262 B.n261 585
R132 B.n260 B.n47 585
R133 B.n259 B.n258 585
R134 B.n257 B.n48 585
R135 B.n256 B.n255 585
R136 B.n254 B.n49 585
R137 B.n253 B.n252 585
R138 B.n251 B.n50 585
R139 B.n250 B.n249 585
R140 B.n248 B.n51 585
R141 B.n247 B.n246 585
R142 B.n245 B.n52 585
R143 B.n244 B.n243 585
R144 B.n242 B.n53 585
R145 B.n241 B.n240 585
R146 B.n239 B.n54 585
R147 B.n238 B.n237 585
R148 B.n236 B.n55 585
R149 B.n235 B.n234 585
R150 B.n233 B.n56 585
R151 B.n232 B.n231 585
R152 B.n230 B.n57 585
R153 B.n229 B.n228 585
R154 B.n227 B.n58 585
R155 B.n226 B.n225 585
R156 B.n224 B.n59 585
R157 B.n223 B.n222 585
R158 B.n221 B.n60 585
R159 B.n220 B.n219 585
R160 B.n218 B.n61 585
R161 B.n217 B.n216 585
R162 B.n215 B.n62 585
R163 B.n214 B.n213 585
R164 B.n212 B.n63 585
R165 B.n211 B.n210 585
R166 B.n209 B.n64 585
R167 B.n208 B.n207 585
R168 B.n206 B.n65 585
R169 B.n205 B.n204 585
R170 B.n203 B.n66 585
R171 B.n202 B.n201 585
R172 B.n200 B.n67 585
R173 B.n199 B.n198 585
R174 B.n197 B.n68 585
R175 B.n196 B.n195 585
R176 B.n194 B.n69 585
R177 B.n152 B.n87 585
R178 B.n154 B.n153 585
R179 B.n155 B.n86 585
R180 B.n157 B.n156 585
R181 B.n158 B.n85 585
R182 B.n160 B.n159 585
R183 B.n161 B.n84 585
R184 B.n163 B.n162 585
R185 B.n164 B.n81 585
R186 B.n167 B.n166 585
R187 B.n168 B.n80 585
R188 B.n170 B.n169 585
R189 B.n171 B.n79 585
R190 B.n173 B.n172 585
R191 B.n174 B.n78 585
R192 B.n176 B.n175 585
R193 B.n177 B.n77 585
R194 B.n179 B.n178 585
R195 B.n181 B.n180 585
R196 B.n182 B.n73 585
R197 B.n184 B.n183 585
R198 B.n185 B.n72 585
R199 B.n187 B.n186 585
R200 B.n188 B.n71 585
R201 B.n190 B.n189 585
R202 B.n191 B.n70 585
R203 B.n193 B.n192 585
R204 B.n151 B.n150 585
R205 B.n149 B.n88 585
R206 B.n148 B.n147 585
R207 B.n146 B.n89 585
R208 B.n145 B.n144 585
R209 B.n143 B.n90 585
R210 B.n142 B.n141 585
R211 B.n140 B.n91 585
R212 B.n139 B.n138 585
R213 B.n137 B.n92 585
R214 B.n136 B.n135 585
R215 B.n134 B.n93 585
R216 B.n133 B.n132 585
R217 B.n131 B.n94 585
R218 B.n130 B.n129 585
R219 B.n128 B.n95 585
R220 B.n127 B.n126 585
R221 B.n125 B.n96 585
R222 B.n124 B.n123 585
R223 B.n122 B.n97 585
R224 B.n121 B.n120 585
R225 B.n119 B.n98 585
R226 B.n118 B.n117 585
R227 B.n116 B.n99 585
R228 B.n115 B.n114 585
R229 B.n113 B.n100 585
R230 B.n112 B.n111 585
R231 B.n110 B.n101 585
R232 B.n109 B.n108 585
R233 B.n107 B.n102 585
R234 B.n106 B.n105 585
R235 B.n104 B.n103 585
R236 B.n2 B.n0 585
R237 B.n385 B.n1 585
R238 B.n384 B.n383 585
R239 B.n382 B.n3 585
R240 B.n381 B.n380 585
R241 B.n379 B.n4 585
R242 B.n378 B.n377 585
R243 B.n376 B.n5 585
R244 B.n375 B.n374 585
R245 B.n373 B.n6 585
R246 B.n372 B.n371 585
R247 B.n370 B.n7 585
R248 B.n369 B.n368 585
R249 B.n367 B.n8 585
R250 B.n366 B.n365 585
R251 B.n364 B.n9 585
R252 B.n363 B.n362 585
R253 B.n361 B.n10 585
R254 B.n360 B.n359 585
R255 B.n358 B.n11 585
R256 B.n357 B.n356 585
R257 B.n355 B.n12 585
R258 B.n354 B.n353 585
R259 B.n352 B.n13 585
R260 B.n351 B.n350 585
R261 B.n349 B.n14 585
R262 B.n348 B.n347 585
R263 B.n346 B.n15 585
R264 B.n345 B.n344 585
R265 B.n343 B.n16 585
R266 B.n342 B.n341 585
R267 B.n340 B.n17 585
R268 B.n339 B.n338 585
R269 B.n337 B.n18 585
R270 B.n387 B.n386 585
R271 B.n150 B.n87 526.135
R272 B.n337 B.n336 526.135
R273 B.n192 B.n69 526.135
R274 B.n294 B.n293 526.135
R275 B.n74 B.t0 207.748
R276 B.n82 B.t6 207.748
R277 B.n24 B.t9 207.748
R278 B.n30 B.t3 207.748
R279 B.n150 B.n149 163.367
R280 B.n149 B.n148 163.367
R281 B.n148 B.n89 163.367
R282 B.n144 B.n89 163.367
R283 B.n144 B.n143 163.367
R284 B.n143 B.n142 163.367
R285 B.n142 B.n91 163.367
R286 B.n138 B.n91 163.367
R287 B.n138 B.n137 163.367
R288 B.n137 B.n136 163.367
R289 B.n136 B.n93 163.367
R290 B.n132 B.n93 163.367
R291 B.n132 B.n131 163.367
R292 B.n131 B.n130 163.367
R293 B.n130 B.n95 163.367
R294 B.n126 B.n95 163.367
R295 B.n126 B.n125 163.367
R296 B.n125 B.n124 163.367
R297 B.n124 B.n97 163.367
R298 B.n120 B.n97 163.367
R299 B.n120 B.n119 163.367
R300 B.n119 B.n118 163.367
R301 B.n118 B.n99 163.367
R302 B.n114 B.n99 163.367
R303 B.n114 B.n113 163.367
R304 B.n113 B.n112 163.367
R305 B.n112 B.n101 163.367
R306 B.n108 B.n101 163.367
R307 B.n108 B.n107 163.367
R308 B.n107 B.n106 163.367
R309 B.n106 B.n103 163.367
R310 B.n103 B.n2 163.367
R311 B.n386 B.n2 163.367
R312 B.n386 B.n385 163.367
R313 B.n385 B.n384 163.367
R314 B.n384 B.n3 163.367
R315 B.n380 B.n3 163.367
R316 B.n380 B.n379 163.367
R317 B.n379 B.n378 163.367
R318 B.n378 B.n5 163.367
R319 B.n374 B.n5 163.367
R320 B.n374 B.n373 163.367
R321 B.n373 B.n372 163.367
R322 B.n372 B.n7 163.367
R323 B.n368 B.n7 163.367
R324 B.n368 B.n367 163.367
R325 B.n367 B.n366 163.367
R326 B.n366 B.n9 163.367
R327 B.n362 B.n9 163.367
R328 B.n362 B.n361 163.367
R329 B.n361 B.n360 163.367
R330 B.n360 B.n11 163.367
R331 B.n356 B.n11 163.367
R332 B.n356 B.n355 163.367
R333 B.n355 B.n354 163.367
R334 B.n354 B.n13 163.367
R335 B.n350 B.n13 163.367
R336 B.n350 B.n349 163.367
R337 B.n349 B.n348 163.367
R338 B.n348 B.n15 163.367
R339 B.n344 B.n15 163.367
R340 B.n344 B.n343 163.367
R341 B.n343 B.n342 163.367
R342 B.n342 B.n17 163.367
R343 B.n338 B.n17 163.367
R344 B.n338 B.n337 163.367
R345 B.n154 B.n87 163.367
R346 B.n155 B.n154 163.367
R347 B.n156 B.n155 163.367
R348 B.n156 B.n85 163.367
R349 B.n160 B.n85 163.367
R350 B.n161 B.n160 163.367
R351 B.n162 B.n161 163.367
R352 B.n162 B.n81 163.367
R353 B.n167 B.n81 163.367
R354 B.n168 B.n167 163.367
R355 B.n169 B.n168 163.367
R356 B.n169 B.n79 163.367
R357 B.n173 B.n79 163.367
R358 B.n174 B.n173 163.367
R359 B.n175 B.n174 163.367
R360 B.n175 B.n77 163.367
R361 B.n179 B.n77 163.367
R362 B.n180 B.n179 163.367
R363 B.n180 B.n73 163.367
R364 B.n184 B.n73 163.367
R365 B.n185 B.n184 163.367
R366 B.n186 B.n185 163.367
R367 B.n186 B.n71 163.367
R368 B.n190 B.n71 163.367
R369 B.n191 B.n190 163.367
R370 B.n192 B.n191 163.367
R371 B.n196 B.n69 163.367
R372 B.n197 B.n196 163.367
R373 B.n198 B.n197 163.367
R374 B.n198 B.n67 163.367
R375 B.n202 B.n67 163.367
R376 B.n203 B.n202 163.367
R377 B.n204 B.n203 163.367
R378 B.n204 B.n65 163.367
R379 B.n208 B.n65 163.367
R380 B.n209 B.n208 163.367
R381 B.n210 B.n209 163.367
R382 B.n210 B.n63 163.367
R383 B.n214 B.n63 163.367
R384 B.n215 B.n214 163.367
R385 B.n216 B.n215 163.367
R386 B.n216 B.n61 163.367
R387 B.n220 B.n61 163.367
R388 B.n221 B.n220 163.367
R389 B.n222 B.n221 163.367
R390 B.n222 B.n59 163.367
R391 B.n226 B.n59 163.367
R392 B.n227 B.n226 163.367
R393 B.n228 B.n227 163.367
R394 B.n228 B.n57 163.367
R395 B.n232 B.n57 163.367
R396 B.n233 B.n232 163.367
R397 B.n234 B.n233 163.367
R398 B.n234 B.n55 163.367
R399 B.n238 B.n55 163.367
R400 B.n239 B.n238 163.367
R401 B.n240 B.n239 163.367
R402 B.n240 B.n53 163.367
R403 B.n244 B.n53 163.367
R404 B.n245 B.n244 163.367
R405 B.n246 B.n245 163.367
R406 B.n246 B.n51 163.367
R407 B.n250 B.n51 163.367
R408 B.n251 B.n250 163.367
R409 B.n252 B.n251 163.367
R410 B.n252 B.n49 163.367
R411 B.n256 B.n49 163.367
R412 B.n257 B.n256 163.367
R413 B.n258 B.n257 163.367
R414 B.n258 B.n47 163.367
R415 B.n262 B.n47 163.367
R416 B.n263 B.n262 163.367
R417 B.n264 B.n263 163.367
R418 B.n264 B.n45 163.367
R419 B.n268 B.n45 163.367
R420 B.n269 B.n268 163.367
R421 B.n270 B.n269 163.367
R422 B.n270 B.n43 163.367
R423 B.n274 B.n43 163.367
R424 B.n275 B.n274 163.367
R425 B.n276 B.n275 163.367
R426 B.n276 B.n41 163.367
R427 B.n280 B.n41 163.367
R428 B.n281 B.n280 163.367
R429 B.n282 B.n281 163.367
R430 B.n282 B.n39 163.367
R431 B.n286 B.n39 163.367
R432 B.n287 B.n286 163.367
R433 B.n288 B.n287 163.367
R434 B.n288 B.n37 163.367
R435 B.n292 B.n37 163.367
R436 B.n293 B.n292 163.367
R437 B.n336 B.n19 163.367
R438 B.n332 B.n19 163.367
R439 B.n332 B.n331 163.367
R440 B.n331 B.n330 163.367
R441 B.n330 B.n21 163.367
R442 B.n326 B.n21 163.367
R443 B.n326 B.n325 163.367
R444 B.n325 B.n324 163.367
R445 B.n324 B.n23 163.367
R446 B.n319 B.n23 163.367
R447 B.n319 B.n318 163.367
R448 B.n318 B.n317 163.367
R449 B.n317 B.n27 163.367
R450 B.n313 B.n27 163.367
R451 B.n313 B.n312 163.367
R452 B.n312 B.n311 163.367
R453 B.n311 B.n29 163.367
R454 B.n306 B.n29 163.367
R455 B.n306 B.n305 163.367
R456 B.n305 B.n304 163.367
R457 B.n304 B.n33 163.367
R458 B.n300 B.n33 163.367
R459 B.n300 B.n299 163.367
R460 B.n299 B.n298 163.367
R461 B.n298 B.n35 163.367
R462 B.n294 B.n35 163.367
R463 B.n76 B.n75 59.5399
R464 B.n165 B.n83 59.5399
R465 B.n322 B.n25 59.5399
R466 B.n308 B.n31 59.5399
R467 B.n75 B.n74 41.1157
R468 B.n83 B.n82 41.1157
R469 B.n25 B.n24 41.1157
R470 B.n31 B.n30 41.1157
R471 B.n335 B.n18 34.1859
R472 B.n295 B.n36 34.1859
R473 B.n194 B.n193 34.1859
R474 B.n152 B.n151 34.1859
R475 B B.n387 18.0485
R476 B.n335 B.n334 10.6151
R477 B.n334 B.n333 10.6151
R478 B.n333 B.n20 10.6151
R479 B.n329 B.n20 10.6151
R480 B.n329 B.n328 10.6151
R481 B.n328 B.n327 10.6151
R482 B.n327 B.n22 10.6151
R483 B.n323 B.n22 10.6151
R484 B.n321 B.n320 10.6151
R485 B.n320 B.n26 10.6151
R486 B.n316 B.n26 10.6151
R487 B.n316 B.n315 10.6151
R488 B.n315 B.n314 10.6151
R489 B.n314 B.n28 10.6151
R490 B.n310 B.n28 10.6151
R491 B.n310 B.n309 10.6151
R492 B.n307 B.n32 10.6151
R493 B.n303 B.n32 10.6151
R494 B.n303 B.n302 10.6151
R495 B.n302 B.n301 10.6151
R496 B.n301 B.n34 10.6151
R497 B.n297 B.n34 10.6151
R498 B.n297 B.n296 10.6151
R499 B.n296 B.n295 10.6151
R500 B.n195 B.n194 10.6151
R501 B.n195 B.n68 10.6151
R502 B.n199 B.n68 10.6151
R503 B.n200 B.n199 10.6151
R504 B.n201 B.n200 10.6151
R505 B.n201 B.n66 10.6151
R506 B.n205 B.n66 10.6151
R507 B.n206 B.n205 10.6151
R508 B.n207 B.n206 10.6151
R509 B.n207 B.n64 10.6151
R510 B.n211 B.n64 10.6151
R511 B.n212 B.n211 10.6151
R512 B.n213 B.n212 10.6151
R513 B.n213 B.n62 10.6151
R514 B.n217 B.n62 10.6151
R515 B.n218 B.n217 10.6151
R516 B.n219 B.n218 10.6151
R517 B.n219 B.n60 10.6151
R518 B.n223 B.n60 10.6151
R519 B.n224 B.n223 10.6151
R520 B.n225 B.n224 10.6151
R521 B.n225 B.n58 10.6151
R522 B.n229 B.n58 10.6151
R523 B.n230 B.n229 10.6151
R524 B.n231 B.n230 10.6151
R525 B.n231 B.n56 10.6151
R526 B.n235 B.n56 10.6151
R527 B.n236 B.n235 10.6151
R528 B.n237 B.n236 10.6151
R529 B.n237 B.n54 10.6151
R530 B.n241 B.n54 10.6151
R531 B.n242 B.n241 10.6151
R532 B.n243 B.n242 10.6151
R533 B.n243 B.n52 10.6151
R534 B.n247 B.n52 10.6151
R535 B.n248 B.n247 10.6151
R536 B.n249 B.n248 10.6151
R537 B.n249 B.n50 10.6151
R538 B.n253 B.n50 10.6151
R539 B.n254 B.n253 10.6151
R540 B.n255 B.n254 10.6151
R541 B.n255 B.n48 10.6151
R542 B.n259 B.n48 10.6151
R543 B.n260 B.n259 10.6151
R544 B.n261 B.n260 10.6151
R545 B.n261 B.n46 10.6151
R546 B.n265 B.n46 10.6151
R547 B.n266 B.n265 10.6151
R548 B.n267 B.n266 10.6151
R549 B.n267 B.n44 10.6151
R550 B.n271 B.n44 10.6151
R551 B.n272 B.n271 10.6151
R552 B.n273 B.n272 10.6151
R553 B.n273 B.n42 10.6151
R554 B.n277 B.n42 10.6151
R555 B.n278 B.n277 10.6151
R556 B.n279 B.n278 10.6151
R557 B.n279 B.n40 10.6151
R558 B.n283 B.n40 10.6151
R559 B.n284 B.n283 10.6151
R560 B.n285 B.n284 10.6151
R561 B.n285 B.n38 10.6151
R562 B.n289 B.n38 10.6151
R563 B.n290 B.n289 10.6151
R564 B.n291 B.n290 10.6151
R565 B.n291 B.n36 10.6151
R566 B.n153 B.n152 10.6151
R567 B.n153 B.n86 10.6151
R568 B.n157 B.n86 10.6151
R569 B.n158 B.n157 10.6151
R570 B.n159 B.n158 10.6151
R571 B.n159 B.n84 10.6151
R572 B.n163 B.n84 10.6151
R573 B.n164 B.n163 10.6151
R574 B.n166 B.n80 10.6151
R575 B.n170 B.n80 10.6151
R576 B.n171 B.n170 10.6151
R577 B.n172 B.n171 10.6151
R578 B.n172 B.n78 10.6151
R579 B.n176 B.n78 10.6151
R580 B.n177 B.n176 10.6151
R581 B.n178 B.n177 10.6151
R582 B.n182 B.n181 10.6151
R583 B.n183 B.n182 10.6151
R584 B.n183 B.n72 10.6151
R585 B.n187 B.n72 10.6151
R586 B.n188 B.n187 10.6151
R587 B.n189 B.n188 10.6151
R588 B.n189 B.n70 10.6151
R589 B.n193 B.n70 10.6151
R590 B.n151 B.n88 10.6151
R591 B.n147 B.n88 10.6151
R592 B.n147 B.n146 10.6151
R593 B.n146 B.n145 10.6151
R594 B.n145 B.n90 10.6151
R595 B.n141 B.n90 10.6151
R596 B.n141 B.n140 10.6151
R597 B.n140 B.n139 10.6151
R598 B.n139 B.n92 10.6151
R599 B.n135 B.n92 10.6151
R600 B.n135 B.n134 10.6151
R601 B.n134 B.n133 10.6151
R602 B.n133 B.n94 10.6151
R603 B.n129 B.n94 10.6151
R604 B.n129 B.n128 10.6151
R605 B.n128 B.n127 10.6151
R606 B.n127 B.n96 10.6151
R607 B.n123 B.n96 10.6151
R608 B.n123 B.n122 10.6151
R609 B.n122 B.n121 10.6151
R610 B.n121 B.n98 10.6151
R611 B.n117 B.n98 10.6151
R612 B.n117 B.n116 10.6151
R613 B.n116 B.n115 10.6151
R614 B.n115 B.n100 10.6151
R615 B.n111 B.n100 10.6151
R616 B.n111 B.n110 10.6151
R617 B.n110 B.n109 10.6151
R618 B.n109 B.n102 10.6151
R619 B.n105 B.n102 10.6151
R620 B.n105 B.n104 10.6151
R621 B.n104 B.n0 10.6151
R622 B.n383 B.n1 10.6151
R623 B.n383 B.n382 10.6151
R624 B.n382 B.n381 10.6151
R625 B.n381 B.n4 10.6151
R626 B.n377 B.n4 10.6151
R627 B.n377 B.n376 10.6151
R628 B.n376 B.n375 10.6151
R629 B.n375 B.n6 10.6151
R630 B.n371 B.n6 10.6151
R631 B.n371 B.n370 10.6151
R632 B.n370 B.n369 10.6151
R633 B.n369 B.n8 10.6151
R634 B.n365 B.n8 10.6151
R635 B.n365 B.n364 10.6151
R636 B.n364 B.n363 10.6151
R637 B.n363 B.n10 10.6151
R638 B.n359 B.n10 10.6151
R639 B.n359 B.n358 10.6151
R640 B.n358 B.n357 10.6151
R641 B.n357 B.n12 10.6151
R642 B.n353 B.n12 10.6151
R643 B.n353 B.n352 10.6151
R644 B.n352 B.n351 10.6151
R645 B.n351 B.n14 10.6151
R646 B.n347 B.n14 10.6151
R647 B.n347 B.n346 10.6151
R648 B.n346 B.n345 10.6151
R649 B.n345 B.n16 10.6151
R650 B.n341 B.n16 10.6151
R651 B.n341 B.n340 10.6151
R652 B.n340 B.n339 10.6151
R653 B.n339 B.n18 10.6151
R654 B.n322 B.n321 6.5566
R655 B.n309 B.n308 6.5566
R656 B.n166 B.n165 6.5566
R657 B.n178 B.n76 6.5566
R658 B.n323 B.n322 4.05904
R659 B.n308 B.n307 4.05904
R660 B.n165 B.n164 4.05904
R661 B.n181 B.n76 4.05904
R662 B.n387 B.n0 2.81026
R663 B.n387 B.n1 2.81026
R664 VP.n18 VP.n17 179.895
R665 VP.n33 VP.n32 179.895
R666 VP.n16 VP.n15 179.895
R667 VP.n10 VP.n9 161.3
R668 VP.n11 VP.n6 161.3
R669 VP.n13 VP.n12 161.3
R670 VP.n14 VP.n5 161.3
R671 VP.n31 VP.n0 161.3
R672 VP.n30 VP.n29 161.3
R673 VP.n28 VP.n1 161.3
R674 VP.n27 VP.n26 161.3
R675 VP.n25 VP.n2 161.3
R676 VP.n24 VP.n23 161.3
R677 VP.n22 VP.n3 161.3
R678 VP.n21 VP.n20 161.3
R679 VP.n19 VP.n4 161.3
R680 VP.n7 VP.t2 47.3648
R681 VP.n20 VP.n3 46.321
R682 VP.n30 VP.n1 46.321
R683 VP.n13 VP.n6 46.321
R684 VP.n8 VP.n7 44.4801
R685 VP.n17 VP.n16 36.9854
R686 VP.n24 VP.n3 34.6658
R687 VP.n26 VP.n1 34.6658
R688 VP.n9 VP.n6 34.6658
R689 VP.n20 VP.n19 24.4675
R690 VP.n25 VP.n24 24.4675
R691 VP.n26 VP.n25 24.4675
R692 VP.n31 VP.n30 24.4675
R693 VP.n14 VP.n13 24.4675
R694 VP.n9 VP.n8 24.4675
R695 VP.n10 VP.n7 12.138
R696 VP.n25 VP.t3 11.4446
R697 VP.n18 VP.t1 11.4446
R698 VP.n32 VP.t0 11.4446
R699 VP.n8 VP.t5 11.4446
R700 VP.n15 VP.t4 11.4446
R701 VP.n19 VP.n18 5.87258
R702 VP.n32 VP.n31 5.87258
R703 VP.n15 VP.n14 5.87258
R704 VP.n11 VP.n10 0.189894
R705 VP.n12 VP.n11 0.189894
R706 VP.n12 VP.n5 0.189894
R707 VP.n16 VP.n5 0.189894
R708 VP.n17 VP.n4 0.189894
R709 VP.n21 VP.n4 0.189894
R710 VP.n22 VP.n21 0.189894
R711 VP.n23 VP.n22 0.189894
R712 VP.n23 VP.n2 0.189894
R713 VP.n27 VP.n2 0.189894
R714 VP.n28 VP.n27 0.189894
R715 VP.n29 VP.n28 0.189894
R716 VP.n29 VP.n0 0.189894
R717 VP.n33 VP.n0 0.189894
R718 VP VP.n33 0.0516364
R719 VDD1 VDD1.t3 676.894
R720 VDD1.n1 VDD1.t4 676.779
R721 VDD1.n1 VDD1.n0 637.625
R722 VDD1.n3 VDD1.n2 637.223
R723 VDD1.n2 VDD1.t0 38.2417
R724 VDD1.n2 VDD1.t1 38.2417
R725 VDD1.n0 VDD1.t2 38.2417
R726 VDD1.n0 VDD1.t5 38.2417
R727 VDD1.n3 VDD1.n1 31.8845
R728 VDD1 VDD1.n3 0.399207
C0 VN VDD2 0.788052f
C1 VDD1 VN 0.157575f
C2 VP VN 4.08202f
C3 VDD1 VDD2 1.11428f
C4 VTAIL VN 1.50575f
C5 VP VDD2 0.398039f
C6 B VN 0.820338f
C7 VN w_n2666_n1138# 4.6189f
C8 VTAIL VDD2 3.13118f
C9 VDD1 VP 1.02581f
C10 VDD1 VTAIL 3.0833f
C11 B VDD2 1.06931f
C12 w_n2666_n1138# VDD2 1.34952f
C13 VTAIL VP 1.51988f
C14 VDD1 B 1.01407f
C15 VDD1 w_n2666_n1138# 1.29153f
C16 VP B 1.38662f
C17 VP w_n2666_n1138# 4.95305f
C18 VTAIL B 0.872287f
C19 VTAIL w_n2666_n1138# 1.21966f
C20 B w_n2666_n1138# 5.47081f
C21 VDD2 VSUBS 0.811623f
C22 VDD1 VSUBS 1.15859f
C23 VTAIL VSUBS 0.35475f
C24 VN VSUBS 4.65758f
C25 VP VSUBS 1.721095f
C26 B VSUBS 2.733161f
C27 w_n2666_n1138# VSUBS 39.190197f
C28 VDD1.t3 VSUBS 0.062775f
C29 VDD1.t4 VSUBS 0.062726f
C30 VDD1.t2 VSUBS 0.012036f
C31 VDD1.t5 VSUBS 0.012036f
C32 VDD1.n0 VSUBS 0.032668f
C33 VDD1.n1 VSUBS 1.35314f
C34 VDD1.t0 VSUBS 0.012036f
C35 VDD1.t1 VSUBS 0.012036f
C36 VDD1.n2 VSUBS 0.032501f
C37 VDD1.n3 VSUBS 1.18263f
C38 VP.n0 VSUBS 0.059287f
C39 VP.t0 VSUBS 0.153662f
C40 VP.n1 VSUBS 0.050727f
C41 VP.n2 VSUBS 0.059287f
C42 VP.t3 VSUBS 0.153662f
C43 VP.n3 VSUBS 0.050727f
C44 VP.n4 VSUBS 0.059287f
C45 VP.t1 VSUBS 0.153662f
C46 VP.n5 VSUBS 0.059287f
C47 VP.t4 VSUBS 0.153662f
C48 VP.n6 VSUBS 0.050727f
C49 VP.t2 VSUBS 0.472413f
C50 VP.n7 VSUBS 0.220291f
C51 VP.t5 VSUBS 0.153662f
C52 VP.n8 VSUBS 0.29874f
C53 VP.n9 VSUBS 0.119801f
C54 VP.n10 VSUBS 0.438043f
C55 VP.n11 VSUBS 0.059287f
C56 VP.n12 VSUBS 0.059287f
C57 VP.n13 VSUBS 0.113066f
C58 VP.n14 VSUBS 0.069036f
C59 VP.n15 VSUBS 0.278003f
C60 VP.n16 VSUBS 1.97588f
C61 VP.n17 VSUBS 2.03351f
C62 VP.n18 VSUBS 0.278003f
C63 VP.n19 VSUBS 0.069036f
C64 VP.n20 VSUBS 0.113066f
C65 VP.n21 VSUBS 0.059287f
C66 VP.n22 VSUBS 0.059287f
C67 VP.n23 VSUBS 0.059287f
C68 VP.n24 VSUBS 0.119801f
C69 VP.n25 VSUBS 0.194763f
C70 VP.n26 VSUBS 0.119801f
C71 VP.n27 VSUBS 0.059287f
C72 VP.n28 VSUBS 0.059287f
C73 VP.n29 VSUBS 0.059287f
C74 VP.n30 VSUBS 0.113066f
C75 VP.n31 VSUBS 0.069036f
C76 VP.n32 VSUBS 0.278003f
C77 VP.n33 VSUBS 0.061991f
C78 B.n0 VSUBS 0.006648f
C79 B.n1 VSUBS 0.006648f
C80 B.n2 VSUBS 0.010512f
C81 B.n3 VSUBS 0.010512f
C82 B.n4 VSUBS 0.010512f
C83 B.n5 VSUBS 0.010512f
C84 B.n6 VSUBS 0.010512f
C85 B.n7 VSUBS 0.010512f
C86 B.n8 VSUBS 0.010512f
C87 B.n9 VSUBS 0.010512f
C88 B.n10 VSUBS 0.010512f
C89 B.n11 VSUBS 0.010512f
C90 B.n12 VSUBS 0.010512f
C91 B.n13 VSUBS 0.010512f
C92 B.n14 VSUBS 0.010512f
C93 B.n15 VSUBS 0.010512f
C94 B.n16 VSUBS 0.010512f
C95 B.n17 VSUBS 0.010512f
C96 B.n18 VSUBS 0.024847f
C97 B.n19 VSUBS 0.010512f
C98 B.n20 VSUBS 0.010512f
C99 B.n21 VSUBS 0.010512f
C100 B.n22 VSUBS 0.010512f
C101 B.n23 VSUBS 0.010512f
C102 B.t11 VSUBS 0.024603f
C103 B.t10 VSUBS 0.027287f
C104 B.t9 VSUBS 0.118148f
C105 B.n24 VSUBS 0.073564f
C106 B.n25 VSUBS 0.060059f
C107 B.n26 VSUBS 0.010512f
C108 B.n27 VSUBS 0.010512f
C109 B.n28 VSUBS 0.010512f
C110 B.n29 VSUBS 0.010512f
C111 B.t5 VSUBS 0.024603f
C112 B.t4 VSUBS 0.027287f
C113 B.t3 VSUBS 0.118148f
C114 B.n30 VSUBS 0.073564f
C115 B.n31 VSUBS 0.060059f
C116 B.n32 VSUBS 0.010512f
C117 B.n33 VSUBS 0.010512f
C118 B.n34 VSUBS 0.010512f
C119 B.n35 VSUBS 0.010512f
C120 B.n36 VSUBS 0.026034f
C121 B.n37 VSUBS 0.010512f
C122 B.n38 VSUBS 0.010512f
C123 B.n39 VSUBS 0.010512f
C124 B.n40 VSUBS 0.010512f
C125 B.n41 VSUBS 0.010512f
C126 B.n42 VSUBS 0.010512f
C127 B.n43 VSUBS 0.010512f
C128 B.n44 VSUBS 0.010512f
C129 B.n45 VSUBS 0.010512f
C130 B.n46 VSUBS 0.010512f
C131 B.n47 VSUBS 0.010512f
C132 B.n48 VSUBS 0.010512f
C133 B.n49 VSUBS 0.010512f
C134 B.n50 VSUBS 0.010512f
C135 B.n51 VSUBS 0.010512f
C136 B.n52 VSUBS 0.010512f
C137 B.n53 VSUBS 0.010512f
C138 B.n54 VSUBS 0.010512f
C139 B.n55 VSUBS 0.010512f
C140 B.n56 VSUBS 0.010512f
C141 B.n57 VSUBS 0.010512f
C142 B.n58 VSUBS 0.010512f
C143 B.n59 VSUBS 0.010512f
C144 B.n60 VSUBS 0.010512f
C145 B.n61 VSUBS 0.010512f
C146 B.n62 VSUBS 0.010512f
C147 B.n63 VSUBS 0.010512f
C148 B.n64 VSUBS 0.010512f
C149 B.n65 VSUBS 0.010512f
C150 B.n66 VSUBS 0.010512f
C151 B.n67 VSUBS 0.010512f
C152 B.n68 VSUBS 0.010512f
C153 B.n69 VSUBS 0.024847f
C154 B.n70 VSUBS 0.010512f
C155 B.n71 VSUBS 0.010512f
C156 B.n72 VSUBS 0.010512f
C157 B.n73 VSUBS 0.010512f
C158 B.t1 VSUBS 0.024603f
C159 B.t2 VSUBS 0.027287f
C160 B.t0 VSUBS 0.118148f
C161 B.n74 VSUBS 0.073564f
C162 B.n75 VSUBS 0.060059f
C163 B.n76 VSUBS 0.024356f
C164 B.n77 VSUBS 0.010512f
C165 B.n78 VSUBS 0.010512f
C166 B.n79 VSUBS 0.010512f
C167 B.n80 VSUBS 0.010512f
C168 B.n81 VSUBS 0.010512f
C169 B.t7 VSUBS 0.024603f
C170 B.t8 VSUBS 0.027287f
C171 B.t6 VSUBS 0.118148f
C172 B.n82 VSUBS 0.073564f
C173 B.n83 VSUBS 0.060059f
C174 B.n84 VSUBS 0.010512f
C175 B.n85 VSUBS 0.010512f
C176 B.n86 VSUBS 0.010512f
C177 B.n87 VSUBS 0.02586f
C178 B.n88 VSUBS 0.010512f
C179 B.n89 VSUBS 0.010512f
C180 B.n90 VSUBS 0.010512f
C181 B.n91 VSUBS 0.010512f
C182 B.n92 VSUBS 0.010512f
C183 B.n93 VSUBS 0.010512f
C184 B.n94 VSUBS 0.010512f
C185 B.n95 VSUBS 0.010512f
C186 B.n96 VSUBS 0.010512f
C187 B.n97 VSUBS 0.010512f
C188 B.n98 VSUBS 0.010512f
C189 B.n99 VSUBS 0.010512f
C190 B.n100 VSUBS 0.010512f
C191 B.n101 VSUBS 0.010512f
C192 B.n102 VSUBS 0.010512f
C193 B.n103 VSUBS 0.010512f
C194 B.n104 VSUBS 0.010512f
C195 B.n105 VSUBS 0.010512f
C196 B.n106 VSUBS 0.010512f
C197 B.n107 VSUBS 0.010512f
C198 B.n108 VSUBS 0.010512f
C199 B.n109 VSUBS 0.010512f
C200 B.n110 VSUBS 0.010512f
C201 B.n111 VSUBS 0.010512f
C202 B.n112 VSUBS 0.010512f
C203 B.n113 VSUBS 0.010512f
C204 B.n114 VSUBS 0.010512f
C205 B.n115 VSUBS 0.010512f
C206 B.n116 VSUBS 0.010512f
C207 B.n117 VSUBS 0.010512f
C208 B.n118 VSUBS 0.010512f
C209 B.n119 VSUBS 0.010512f
C210 B.n120 VSUBS 0.010512f
C211 B.n121 VSUBS 0.010512f
C212 B.n122 VSUBS 0.010512f
C213 B.n123 VSUBS 0.010512f
C214 B.n124 VSUBS 0.010512f
C215 B.n125 VSUBS 0.010512f
C216 B.n126 VSUBS 0.010512f
C217 B.n127 VSUBS 0.010512f
C218 B.n128 VSUBS 0.010512f
C219 B.n129 VSUBS 0.010512f
C220 B.n130 VSUBS 0.010512f
C221 B.n131 VSUBS 0.010512f
C222 B.n132 VSUBS 0.010512f
C223 B.n133 VSUBS 0.010512f
C224 B.n134 VSUBS 0.010512f
C225 B.n135 VSUBS 0.010512f
C226 B.n136 VSUBS 0.010512f
C227 B.n137 VSUBS 0.010512f
C228 B.n138 VSUBS 0.010512f
C229 B.n139 VSUBS 0.010512f
C230 B.n140 VSUBS 0.010512f
C231 B.n141 VSUBS 0.010512f
C232 B.n142 VSUBS 0.010512f
C233 B.n143 VSUBS 0.010512f
C234 B.n144 VSUBS 0.010512f
C235 B.n145 VSUBS 0.010512f
C236 B.n146 VSUBS 0.010512f
C237 B.n147 VSUBS 0.010512f
C238 B.n148 VSUBS 0.010512f
C239 B.n149 VSUBS 0.010512f
C240 B.n150 VSUBS 0.024847f
C241 B.n151 VSUBS 0.024847f
C242 B.n152 VSUBS 0.02586f
C243 B.n153 VSUBS 0.010512f
C244 B.n154 VSUBS 0.010512f
C245 B.n155 VSUBS 0.010512f
C246 B.n156 VSUBS 0.010512f
C247 B.n157 VSUBS 0.010512f
C248 B.n158 VSUBS 0.010512f
C249 B.n159 VSUBS 0.010512f
C250 B.n160 VSUBS 0.010512f
C251 B.n161 VSUBS 0.010512f
C252 B.n162 VSUBS 0.010512f
C253 B.n163 VSUBS 0.010512f
C254 B.n164 VSUBS 0.007266f
C255 B.n165 VSUBS 0.024356f
C256 B.n166 VSUBS 0.008503f
C257 B.n167 VSUBS 0.010512f
C258 B.n168 VSUBS 0.010512f
C259 B.n169 VSUBS 0.010512f
C260 B.n170 VSUBS 0.010512f
C261 B.n171 VSUBS 0.010512f
C262 B.n172 VSUBS 0.010512f
C263 B.n173 VSUBS 0.010512f
C264 B.n174 VSUBS 0.010512f
C265 B.n175 VSUBS 0.010512f
C266 B.n176 VSUBS 0.010512f
C267 B.n177 VSUBS 0.010512f
C268 B.n178 VSUBS 0.008503f
C269 B.n179 VSUBS 0.010512f
C270 B.n180 VSUBS 0.010512f
C271 B.n181 VSUBS 0.007266f
C272 B.n182 VSUBS 0.010512f
C273 B.n183 VSUBS 0.010512f
C274 B.n184 VSUBS 0.010512f
C275 B.n185 VSUBS 0.010512f
C276 B.n186 VSUBS 0.010512f
C277 B.n187 VSUBS 0.010512f
C278 B.n188 VSUBS 0.010512f
C279 B.n189 VSUBS 0.010512f
C280 B.n190 VSUBS 0.010512f
C281 B.n191 VSUBS 0.010512f
C282 B.n192 VSUBS 0.02586f
C283 B.n193 VSUBS 0.02586f
C284 B.n194 VSUBS 0.024847f
C285 B.n195 VSUBS 0.010512f
C286 B.n196 VSUBS 0.010512f
C287 B.n197 VSUBS 0.010512f
C288 B.n198 VSUBS 0.010512f
C289 B.n199 VSUBS 0.010512f
C290 B.n200 VSUBS 0.010512f
C291 B.n201 VSUBS 0.010512f
C292 B.n202 VSUBS 0.010512f
C293 B.n203 VSUBS 0.010512f
C294 B.n204 VSUBS 0.010512f
C295 B.n205 VSUBS 0.010512f
C296 B.n206 VSUBS 0.010512f
C297 B.n207 VSUBS 0.010512f
C298 B.n208 VSUBS 0.010512f
C299 B.n209 VSUBS 0.010512f
C300 B.n210 VSUBS 0.010512f
C301 B.n211 VSUBS 0.010512f
C302 B.n212 VSUBS 0.010512f
C303 B.n213 VSUBS 0.010512f
C304 B.n214 VSUBS 0.010512f
C305 B.n215 VSUBS 0.010512f
C306 B.n216 VSUBS 0.010512f
C307 B.n217 VSUBS 0.010512f
C308 B.n218 VSUBS 0.010512f
C309 B.n219 VSUBS 0.010512f
C310 B.n220 VSUBS 0.010512f
C311 B.n221 VSUBS 0.010512f
C312 B.n222 VSUBS 0.010512f
C313 B.n223 VSUBS 0.010512f
C314 B.n224 VSUBS 0.010512f
C315 B.n225 VSUBS 0.010512f
C316 B.n226 VSUBS 0.010512f
C317 B.n227 VSUBS 0.010512f
C318 B.n228 VSUBS 0.010512f
C319 B.n229 VSUBS 0.010512f
C320 B.n230 VSUBS 0.010512f
C321 B.n231 VSUBS 0.010512f
C322 B.n232 VSUBS 0.010512f
C323 B.n233 VSUBS 0.010512f
C324 B.n234 VSUBS 0.010512f
C325 B.n235 VSUBS 0.010512f
C326 B.n236 VSUBS 0.010512f
C327 B.n237 VSUBS 0.010512f
C328 B.n238 VSUBS 0.010512f
C329 B.n239 VSUBS 0.010512f
C330 B.n240 VSUBS 0.010512f
C331 B.n241 VSUBS 0.010512f
C332 B.n242 VSUBS 0.010512f
C333 B.n243 VSUBS 0.010512f
C334 B.n244 VSUBS 0.010512f
C335 B.n245 VSUBS 0.010512f
C336 B.n246 VSUBS 0.010512f
C337 B.n247 VSUBS 0.010512f
C338 B.n248 VSUBS 0.010512f
C339 B.n249 VSUBS 0.010512f
C340 B.n250 VSUBS 0.010512f
C341 B.n251 VSUBS 0.010512f
C342 B.n252 VSUBS 0.010512f
C343 B.n253 VSUBS 0.010512f
C344 B.n254 VSUBS 0.010512f
C345 B.n255 VSUBS 0.010512f
C346 B.n256 VSUBS 0.010512f
C347 B.n257 VSUBS 0.010512f
C348 B.n258 VSUBS 0.010512f
C349 B.n259 VSUBS 0.010512f
C350 B.n260 VSUBS 0.010512f
C351 B.n261 VSUBS 0.010512f
C352 B.n262 VSUBS 0.010512f
C353 B.n263 VSUBS 0.010512f
C354 B.n264 VSUBS 0.010512f
C355 B.n265 VSUBS 0.010512f
C356 B.n266 VSUBS 0.010512f
C357 B.n267 VSUBS 0.010512f
C358 B.n268 VSUBS 0.010512f
C359 B.n269 VSUBS 0.010512f
C360 B.n270 VSUBS 0.010512f
C361 B.n271 VSUBS 0.010512f
C362 B.n272 VSUBS 0.010512f
C363 B.n273 VSUBS 0.010512f
C364 B.n274 VSUBS 0.010512f
C365 B.n275 VSUBS 0.010512f
C366 B.n276 VSUBS 0.010512f
C367 B.n277 VSUBS 0.010512f
C368 B.n278 VSUBS 0.010512f
C369 B.n279 VSUBS 0.010512f
C370 B.n280 VSUBS 0.010512f
C371 B.n281 VSUBS 0.010512f
C372 B.n282 VSUBS 0.010512f
C373 B.n283 VSUBS 0.010512f
C374 B.n284 VSUBS 0.010512f
C375 B.n285 VSUBS 0.010512f
C376 B.n286 VSUBS 0.010512f
C377 B.n287 VSUBS 0.010512f
C378 B.n288 VSUBS 0.010512f
C379 B.n289 VSUBS 0.010512f
C380 B.n290 VSUBS 0.010512f
C381 B.n291 VSUBS 0.010512f
C382 B.n292 VSUBS 0.010512f
C383 B.n293 VSUBS 0.024847f
C384 B.n294 VSUBS 0.02586f
C385 B.n295 VSUBS 0.024673f
C386 B.n296 VSUBS 0.010512f
C387 B.n297 VSUBS 0.010512f
C388 B.n298 VSUBS 0.010512f
C389 B.n299 VSUBS 0.010512f
C390 B.n300 VSUBS 0.010512f
C391 B.n301 VSUBS 0.010512f
C392 B.n302 VSUBS 0.010512f
C393 B.n303 VSUBS 0.010512f
C394 B.n304 VSUBS 0.010512f
C395 B.n305 VSUBS 0.010512f
C396 B.n306 VSUBS 0.010512f
C397 B.n307 VSUBS 0.007266f
C398 B.n308 VSUBS 0.024356f
C399 B.n309 VSUBS 0.008503f
C400 B.n310 VSUBS 0.010512f
C401 B.n311 VSUBS 0.010512f
C402 B.n312 VSUBS 0.010512f
C403 B.n313 VSUBS 0.010512f
C404 B.n314 VSUBS 0.010512f
C405 B.n315 VSUBS 0.010512f
C406 B.n316 VSUBS 0.010512f
C407 B.n317 VSUBS 0.010512f
C408 B.n318 VSUBS 0.010512f
C409 B.n319 VSUBS 0.010512f
C410 B.n320 VSUBS 0.010512f
C411 B.n321 VSUBS 0.008503f
C412 B.n322 VSUBS 0.024356f
C413 B.n323 VSUBS 0.007266f
C414 B.n324 VSUBS 0.010512f
C415 B.n325 VSUBS 0.010512f
C416 B.n326 VSUBS 0.010512f
C417 B.n327 VSUBS 0.010512f
C418 B.n328 VSUBS 0.010512f
C419 B.n329 VSUBS 0.010512f
C420 B.n330 VSUBS 0.010512f
C421 B.n331 VSUBS 0.010512f
C422 B.n332 VSUBS 0.010512f
C423 B.n333 VSUBS 0.010512f
C424 B.n334 VSUBS 0.010512f
C425 B.n335 VSUBS 0.02586f
C426 B.n336 VSUBS 0.02586f
C427 B.n337 VSUBS 0.024847f
C428 B.n338 VSUBS 0.010512f
C429 B.n339 VSUBS 0.010512f
C430 B.n340 VSUBS 0.010512f
C431 B.n341 VSUBS 0.010512f
C432 B.n342 VSUBS 0.010512f
C433 B.n343 VSUBS 0.010512f
C434 B.n344 VSUBS 0.010512f
C435 B.n345 VSUBS 0.010512f
C436 B.n346 VSUBS 0.010512f
C437 B.n347 VSUBS 0.010512f
C438 B.n348 VSUBS 0.010512f
C439 B.n349 VSUBS 0.010512f
C440 B.n350 VSUBS 0.010512f
C441 B.n351 VSUBS 0.010512f
C442 B.n352 VSUBS 0.010512f
C443 B.n353 VSUBS 0.010512f
C444 B.n354 VSUBS 0.010512f
C445 B.n355 VSUBS 0.010512f
C446 B.n356 VSUBS 0.010512f
C447 B.n357 VSUBS 0.010512f
C448 B.n358 VSUBS 0.010512f
C449 B.n359 VSUBS 0.010512f
C450 B.n360 VSUBS 0.010512f
C451 B.n361 VSUBS 0.010512f
C452 B.n362 VSUBS 0.010512f
C453 B.n363 VSUBS 0.010512f
C454 B.n364 VSUBS 0.010512f
C455 B.n365 VSUBS 0.010512f
C456 B.n366 VSUBS 0.010512f
C457 B.n367 VSUBS 0.010512f
C458 B.n368 VSUBS 0.010512f
C459 B.n369 VSUBS 0.010512f
C460 B.n370 VSUBS 0.010512f
C461 B.n371 VSUBS 0.010512f
C462 B.n372 VSUBS 0.010512f
C463 B.n373 VSUBS 0.010512f
C464 B.n374 VSUBS 0.010512f
C465 B.n375 VSUBS 0.010512f
C466 B.n376 VSUBS 0.010512f
C467 B.n377 VSUBS 0.010512f
C468 B.n378 VSUBS 0.010512f
C469 B.n379 VSUBS 0.010512f
C470 B.n380 VSUBS 0.010512f
C471 B.n381 VSUBS 0.010512f
C472 B.n382 VSUBS 0.010512f
C473 B.n383 VSUBS 0.010512f
C474 B.n384 VSUBS 0.010512f
C475 B.n385 VSUBS 0.010512f
C476 B.n386 VSUBS 0.010512f
C477 B.n387 VSUBS 0.023804f
C478 VDD2.t4 VSUBS 0.064095f
C479 VDD2.t0 VSUBS 0.012299f
C480 VDD2.t5 VSUBS 0.012299f
C481 VDD2.n0 VSUBS 0.033381f
C482 VDD2.n1 VSUBS 1.31445f
C483 VDD2.t2 VSUBS 0.063669f
C484 VDD2.n2 VSUBS 1.16505f
C485 VDD2.t1 VSUBS 0.012299f
C486 VDD2.t3 VSUBS 0.012299f
C487 VDD2.n3 VSUBS 0.033379f
C488 VTAIL.t8 VSUBS 0.017544f
C489 VTAIL.t6 VSUBS 0.017544f
C490 VTAIL.n0 VSUBS 0.042509f
C491 VTAIL.n1 VSUBS 0.315188f
C492 VTAIL.t4 VSUBS 0.08613f
C493 VTAIL.n2 VSUBS 0.429878f
C494 VTAIL.t5 VSUBS 0.017544f
C495 VTAIL.t2 VSUBS 0.017544f
C496 VTAIL.n3 VSUBS 0.042509f
C497 VTAIL.n4 VSUBS 1.0333f
C498 VTAIL.t10 VSUBS 0.017544f
C499 VTAIL.t7 VSUBS 0.017544f
C500 VTAIL.n5 VSUBS 0.042509f
C501 VTAIL.n6 VSUBS 1.0333f
C502 VTAIL.t9 VSUBS 0.08613f
C503 VTAIL.n7 VSUBS 0.429878f
C504 VTAIL.t1 VSUBS 0.017544f
C505 VTAIL.t0 VSUBS 0.017544f
C506 VTAIL.n8 VSUBS 0.042509f
C507 VTAIL.n9 VSUBS 0.425651f
C508 VTAIL.t3 VSUBS 0.08613f
C509 VTAIL.n10 VSUBS 0.883715f
C510 VTAIL.t11 VSUBS 0.08613f
C511 VTAIL.n11 VSUBS 0.840364f
C512 VN.n0 VSUBS 0.056167f
C513 VN.t0 VSUBS 0.145574f
C514 VN.n1 VSUBS 0.048058f
C515 VN.t1 VSUBS 0.447549f
C516 VN.n2 VSUBS 0.208696f
C517 VN.t5 VSUBS 0.145574f
C518 VN.n3 VSUBS 0.283016f
C519 VN.n4 VSUBS 0.113496f
C520 VN.n5 VSUBS 0.414987f
C521 VN.n6 VSUBS 0.056167f
C522 VN.n7 VSUBS 0.056167f
C523 VN.n8 VSUBS 0.107115f
C524 VN.n9 VSUBS 0.065403f
C525 VN.n10 VSUBS 0.263371f
C526 VN.n11 VSUBS 0.058728f
C527 VN.n12 VSUBS 0.056167f
C528 VN.t3 VSUBS 0.145574f
C529 VN.n13 VSUBS 0.048058f
C530 VN.t2 VSUBS 0.447549f
C531 VN.n14 VSUBS 0.208696f
C532 VN.t4 VSUBS 0.145574f
C533 VN.n15 VSUBS 0.283016f
C534 VN.n16 VSUBS 0.113496f
C535 VN.n17 VSUBS 0.414987f
C536 VN.n18 VSUBS 0.056167f
C537 VN.n19 VSUBS 0.056167f
C538 VN.n20 VSUBS 0.107115f
C539 VN.n21 VSUBS 0.065403f
C540 VN.n22 VSUBS 0.263371f
C541 VN.n23 VSUBS 1.90907f
.ends

