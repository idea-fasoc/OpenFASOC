* NGSPICE file created from diff_pair_sample_0689.ext - technology: sky130A

.subckt diff_pair_sample_0689 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=4.7541 pd=25.16 as=0 ps=0 w=12.19 l=1.75
X1 VTAIL.t19 VP.t0 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X2 VTAIL.t9 VN.t0 VDD2.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X3 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7541 pd=25.16 as=0 ps=0 w=12.19 l=1.75
X4 VTAIL.t18 VP.t1 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X5 VDD1.t7 VP.t2 VTAIL.t17 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7541 pd=25.16 as=2.01135 ps=12.52 w=12.19 l=1.75
X6 VTAIL.t16 VP.t3 VDD1.t0 B.t9 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X7 VDD2.t8 VN.t1 VTAIL.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=4.7541 pd=25.16 as=2.01135 ps=12.52 w=12.19 l=1.75
X8 VTAIL.t2 VN.t2 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X9 VTAIL.t0 VN.t3 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X10 VTAIL.t4 VN.t4 VDD2.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X11 VDD2.t4 VN.t5 VTAIL.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7541 pd=25.16 as=2.01135 ps=12.52 w=12.19 l=1.75
X12 VDD2.t3 VN.t6 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=4.7541 ps=25.16 w=12.19 l=1.75
X13 VDD2.t2 VN.t7 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=4.7541 ps=25.16 w=12.19 l=1.75
X14 VDD1.t1 VP.t4 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=4.7541 ps=25.16 w=12.19 l=1.75
X15 VDD1.t8 VP.t5 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X16 VDD1.t5 VP.t6 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X17 VDD1.t6 VP.t7 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=4.7541 ps=25.16 w=12.19 l=1.75
X18 VDD1.t9 VP.t8 VTAIL.t11 B.t8 sky130_fd_pr__nfet_01v8 ad=4.7541 pd=25.16 as=2.01135 ps=12.52 w=12.19 l=1.75
X19 VDD2.t1 VN.t8 VTAIL.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X20 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.7541 pd=25.16 as=0 ps=0 w=12.19 l=1.75
X21 VDD2.t0 VN.t9 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X22 VTAIL.t10 VP.t9 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=2.01135 pd=12.52 as=2.01135 ps=12.52 w=12.19 l=1.75
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7541 pd=25.16 as=0 ps=0 w=12.19 l=1.75
R0 B.n843 B.n842 585
R1 B.n321 B.n130 585
R2 B.n320 B.n319 585
R3 B.n318 B.n317 585
R4 B.n316 B.n315 585
R5 B.n314 B.n313 585
R6 B.n312 B.n311 585
R7 B.n310 B.n309 585
R8 B.n308 B.n307 585
R9 B.n306 B.n305 585
R10 B.n304 B.n303 585
R11 B.n302 B.n301 585
R12 B.n300 B.n299 585
R13 B.n298 B.n297 585
R14 B.n296 B.n295 585
R15 B.n294 B.n293 585
R16 B.n292 B.n291 585
R17 B.n290 B.n289 585
R18 B.n288 B.n287 585
R19 B.n286 B.n285 585
R20 B.n284 B.n283 585
R21 B.n282 B.n281 585
R22 B.n280 B.n279 585
R23 B.n278 B.n277 585
R24 B.n276 B.n275 585
R25 B.n274 B.n273 585
R26 B.n272 B.n271 585
R27 B.n270 B.n269 585
R28 B.n268 B.n267 585
R29 B.n266 B.n265 585
R30 B.n264 B.n263 585
R31 B.n262 B.n261 585
R32 B.n260 B.n259 585
R33 B.n258 B.n257 585
R34 B.n256 B.n255 585
R35 B.n254 B.n253 585
R36 B.n252 B.n251 585
R37 B.n250 B.n249 585
R38 B.n248 B.n247 585
R39 B.n246 B.n245 585
R40 B.n244 B.n243 585
R41 B.n242 B.n241 585
R42 B.n240 B.n239 585
R43 B.n238 B.n237 585
R44 B.n236 B.n235 585
R45 B.n234 B.n233 585
R46 B.n232 B.n231 585
R47 B.n230 B.n229 585
R48 B.n228 B.n227 585
R49 B.n226 B.n225 585
R50 B.n224 B.n223 585
R51 B.n222 B.n221 585
R52 B.n220 B.n219 585
R53 B.n218 B.n217 585
R54 B.n216 B.n215 585
R55 B.n214 B.n213 585
R56 B.n212 B.n211 585
R57 B.n210 B.n209 585
R58 B.n208 B.n207 585
R59 B.n206 B.n205 585
R60 B.n204 B.n203 585
R61 B.n202 B.n201 585
R62 B.n200 B.n199 585
R63 B.n198 B.n197 585
R64 B.n196 B.n195 585
R65 B.n194 B.n193 585
R66 B.n192 B.n191 585
R67 B.n190 B.n189 585
R68 B.n188 B.n187 585
R69 B.n186 B.n185 585
R70 B.n184 B.n183 585
R71 B.n182 B.n181 585
R72 B.n180 B.n179 585
R73 B.n178 B.n177 585
R74 B.n176 B.n175 585
R75 B.n174 B.n173 585
R76 B.n172 B.n171 585
R77 B.n170 B.n169 585
R78 B.n168 B.n167 585
R79 B.n166 B.n165 585
R80 B.n164 B.n163 585
R81 B.n162 B.n161 585
R82 B.n160 B.n159 585
R83 B.n158 B.n157 585
R84 B.n156 B.n155 585
R85 B.n154 B.n153 585
R86 B.n152 B.n151 585
R87 B.n150 B.n149 585
R88 B.n148 B.n147 585
R89 B.n146 B.n145 585
R90 B.n144 B.n143 585
R91 B.n142 B.n141 585
R92 B.n140 B.n139 585
R93 B.n138 B.n137 585
R94 B.n841 B.n83 585
R95 B.n846 B.n83 585
R96 B.n840 B.n82 585
R97 B.n847 B.n82 585
R98 B.n839 B.n838 585
R99 B.n838 B.n78 585
R100 B.n837 B.n77 585
R101 B.n853 B.n77 585
R102 B.n836 B.n76 585
R103 B.n854 B.n76 585
R104 B.n835 B.n75 585
R105 B.n855 B.n75 585
R106 B.n834 B.n833 585
R107 B.n833 B.n74 585
R108 B.n832 B.n70 585
R109 B.n861 B.n70 585
R110 B.n831 B.n69 585
R111 B.n862 B.n69 585
R112 B.n830 B.n68 585
R113 B.n863 B.n68 585
R114 B.n829 B.n828 585
R115 B.n828 B.n64 585
R116 B.n827 B.n63 585
R117 B.n869 B.n63 585
R118 B.n826 B.n62 585
R119 B.n870 B.n62 585
R120 B.n825 B.n61 585
R121 B.n871 B.n61 585
R122 B.n824 B.n823 585
R123 B.n823 B.n57 585
R124 B.n822 B.n56 585
R125 B.n877 B.n56 585
R126 B.n821 B.n55 585
R127 B.n878 B.n55 585
R128 B.n820 B.n54 585
R129 B.n879 B.n54 585
R130 B.n819 B.n818 585
R131 B.n818 B.n50 585
R132 B.n817 B.n49 585
R133 B.n885 B.n49 585
R134 B.n816 B.n48 585
R135 B.n886 B.n48 585
R136 B.n815 B.n47 585
R137 B.n887 B.n47 585
R138 B.n814 B.n813 585
R139 B.n813 B.n43 585
R140 B.n812 B.n42 585
R141 B.n893 B.n42 585
R142 B.n811 B.n41 585
R143 B.n894 B.n41 585
R144 B.n810 B.n40 585
R145 B.n895 B.n40 585
R146 B.n809 B.n808 585
R147 B.n808 B.n36 585
R148 B.n807 B.n35 585
R149 B.n901 B.n35 585
R150 B.n806 B.n34 585
R151 B.n902 B.n34 585
R152 B.n805 B.n33 585
R153 B.n903 B.n33 585
R154 B.n804 B.n803 585
R155 B.n803 B.n29 585
R156 B.n802 B.n28 585
R157 B.n909 B.n28 585
R158 B.n801 B.n27 585
R159 B.n910 B.n27 585
R160 B.n800 B.n26 585
R161 B.n911 B.n26 585
R162 B.n799 B.n798 585
R163 B.n798 B.n25 585
R164 B.n797 B.n21 585
R165 B.n917 B.n21 585
R166 B.n796 B.n20 585
R167 B.n918 B.n20 585
R168 B.n795 B.n19 585
R169 B.n919 B.n19 585
R170 B.n794 B.n793 585
R171 B.n793 B.n15 585
R172 B.n792 B.n14 585
R173 B.n925 B.n14 585
R174 B.n791 B.n13 585
R175 B.n926 B.n13 585
R176 B.n790 B.n12 585
R177 B.n927 B.n12 585
R178 B.n789 B.n788 585
R179 B.n788 B.n8 585
R180 B.n787 B.n7 585
R181 B.n933 B.n7 585
R182 B.n786 B.n6 585
R183 B.n934 B.n6 585
R184 B.n785 B.n5 585
R185 B.n935 B.n5 585
R186 B.n784 B.n783 585
R187 B.n783 B.n4 585
R188 B.n782 B.n322 585
R189 B.n782 B.n781 585
R190 B.n772 B.n323 585
R191 B.n324 B.n323 585
R192 B.n774 B.n773 585
R193 B.n775 B.n774 585
R194 B.n771 B.n328 585
R195 B.n332 B.n328 585
R196 B.n770 B.n769 585
R197 B.n769 B.n768 585
R198 B.n330 B.n329 585
R199 B.n331 B.n330 585
R200 B.n761 B.n760 585
R201 B.n762 B.n761 585
R202 B.n759 B.n337 585
R203 B.n337 B.n336 585
R204 B.n758 B.n757 585
R205 B.n757 B.n756 585
R206 B.n339 B.n338 585
R207 B.n749 B.n339 585
R208 B.n748 B.n747 585
R209 B.n750 B.n748 585
R210 B.n746 B.n344 585
R211 B.n344 B.n343 585
R212 B.n745 B.n744 585
R213 B.n744 B.n743 585
R214 B.n346 B.n345 585
R215 B.n347 B.n346 585
R216 B.n736 B.n735 585
R217 B.n737 B.n736 585
R218 B.n734 B.n351 585
R219 B.n355 B.n351 585
R220 B.n733 B.n732 585
R221 B.n732 B.n731 585
R222 B.n353 B.n352 585
R223 B.n354 B.n353 585
R224 B.n724 B.n723 585
R225 B.n725 B.n724 585
R226 B.n722 B.n360 585
R227 B.n360 B.n359 585
R228 B.n721 B.n720 585
R229 B.n720 B.n719 585
R230 B.n362 B.n361 585
R231 B.n363 B.n362 585
R232 B.n712 B.n711 585
R233 B.n713 B.n712 585
R234 B.n710 B.n368 585
R235 B.n368 B.n367 585
R236 B.n709 B.n708 585
R237 B.n708 B.n707 585
R238 B.n370 B.n369 585
R239 B.n371 B.n370 585
R240 B.n700 B.n699 585
R241 B.n701 B.n700 585
R242 B.n698 B.n376 585
R243 B.n376 B.n375 585
R244 B.n697 B.n696 585
R245 B.n696 B.n695 585
R246 B.n378 B.n377 585
R247 B.n379 B.n378 585
R248 B.n688 B.n687 585
R249 B.n689 B.n688 585
R250 B.n686 B.n384 585
R251 B.n384 B.n383 585
R252 B.n685 B.n684 585
R253 B.n684 B.n683 585
R254 B.n386 B.n385 585
R255 B.n387 B.n386 585
R256 B.n676 B.n675 585
R257 B.n677 B.n676 585
R258 B.n674 B.n392 585
R259 B.n392 B.n391 585
R260 B.n673 B.n672 585
R261 B.n672 B.n671 585
R262 B.n394 B.n393 585
R263 B.n664 B.n394 585
R264 B.n663 B.n662 585
R265 B.n665 B.n663 585
R266 B.n661 B.n399 585
R267 B.n399 B.n398 585
R268 B.n660 B.n659 585
R269 B.n659 B.n658 585
R270 B.n401 B.n400 585
R271 B.n402 B.n401 585
R272 B.n651 B.n650 585
R273 B.n652 B.n651 585
R274 B.n649 B.n407 585
R275 B.n407 B.n406 585
R276 B.n644 B.n643 585
R277 B.n642 B.n456 585
R278 B.n641 B.n455 585
R279 B.n646 B.n455 585
R280 B.n640 B.n639 585
R281 B.n638 B.n637 585
R282 B.n636 B.n635 585
R283 B.n634 B.n633 585
R284 B.n632 B.n631 585
R285 B.n630 B.n629 585
R286 B.n628 B.n627 585
R287 B.n626 B.n625 585
R288 B.n624 B.n623 585
R289 B.n622 B.n621 585
R290 B.n620 B.n619 585
R291 B.n618 B.n617 585
R292 B.n616 B.n615 585
R293 B.n614 B.n613 585
R294 B.n612 B.n611 585
R295 B.n610 B.n609 585
R296 B.n608 B.n607 585
R297 B.n606 B.n605 585
R298 B.n604 B.n603 585
R299 B.n602 B.n601 585
R300 B.n600 B.n599 585
R301 B.n598 B.n597 585
R302 B.n596 B.n595 585
R303 B.n594 B.n593 585
R304 B.n592 B.n591 585
R305 B.n590 B.n589 585
R306 B.n588 B.n587 585
R307 B.n586 B.n585 585
R308 B.n584 B.n583 585
R309 B.n582 B.n581 585
R310 B.n580 B.n579 585
R311 B.n578 B.n577 585
R312 B.n576 B.n575 585
R313 B.n574 B.n573 585
R314 B.n572 B.n571 585
R315 B.n570 B.n569 585
R316 B.n568 B.n567 585
R317 B.n566 B.n565 585
R318 B.n564 B.n563 585
R319 B.n561 B.n560 585
R320 B.n559 B.n558 585
R321 B.n557 B.n556 585
R322 B.n555 B.n554 585
R323 B.n553 B.n552 585
R324 B.n551 B.n550 585
R325 B.n549 B.n548 585
R326 B.n547 B.n546 585
R327 B.n545 B.n544 585
R328 B.n543 B.n542 585
R329 B.n540 B.n539 585
R330 B.n538 B.n537 585
R331 B.n536 B.n535 585
R332 B.n534 B.n533 585
R333 B.n532 B.n531 585
R334 B.n530 B.n529 585
R335 B.n528 B.n527 585
R336 B.n526 B.n525 585
R337 B.n524 B.n523 585
R338 B.n522 B.n521 585
R339 B.n520 B.n519 585
R340 B.n518 B.n517 585
R341 B.n516 B.n515 585
R342 B.n514 B.n513 585
R343 B.n512 B.n511 585
R344 B.n510 B.n509 585
R345 B.n508 B.n507 585
R346 B.n506 B.n505 585
R347 B.n504 B.n503 585
R348 B.n502 B.n501 585
R349 B.n500 B.n499 585
R350 B.n498 B.n497 585
R351 B.n496 B.n495 585
R352 B.n494 B.n493 585
R353 B.n492 B.n491 585
R354 B.n490 B.n489 585
R355 B.n488 B.n487 585
R356 B.n486 B.n485 585
R357 B.n484 B.n483 585
R358 B.n482 B.n481 585
R359 B.n480 B.n479 585
R360 B.n478 B.n477 585
R361 B.n476 B.n475 585
R362 B.n474 B.n473 585
R363 B.n472 B.n471 585
R364 B.n470 B.n469 585
R365 B.n468 B.n467 585
R366 B.n466 B.n465 585
R367 B.n464 B.n463 585
R368 B.n462 B.n461 585
R369 B.n409 B.n408 585
R370 B.n648 B.n647 585
R371 B.n647 B.n646 585
R372 B.n405 B.n404 585
R373 B.n406 B.n405 585
R374 B.n654 B.n653 585
R375 B.n653 B.n652 585
R376 B.n655 B.n403 585
R377 B.n403 B.n402 585
R378 B.n657 B.n656 585
R379 B.n658 B.n657 585
R380 B.n397 B.n396 585
R381 B.n398 B.n397 585
R382 B.n667 B.n666 585
R383 B.n666 B.n665 585
R384 B.n668 B.n395 585
R385 B.n664 B.n395 585
R386 B.n670 B.n669 585
R387 B.n671 B.n670 585
R388 B.n390 B.n389 585
R389 B.n391 B.n390 585
R390 B.n679 B.n678 585
R391 B.n678 B.n677 585
R392 B.n680 B.n388 585
R393 B.n388 B.n387 585
R394 B.n682 B.n681 585
R395 B.n683 B.n682 585
R396 B.n382 B.n381 585
R397 B.n383 B.n382 585
R398 B.n691 B.n690 585
R399 B.n690 B.n689 585
R400 B.n692 B.n380 585
R401 B.n380 B.n379 585
R402 B.n694 B.n693 585
R403 B.n695 B.n694 585
R404 B.n374 B.n373 585
R405 B.n375 B.n374 585
R406 B.n703 B.n702 585
R407 B.n702 B.n701 585
R408 B.n704 B.n372 585
R409 B.n372 B.n371 585
R410 B.n706 B.n705 585
R411 B.n707 B.n706 585
R412 B.n366 B.n365 585
R413 B.n367 B.n366 585
R414 B.n715 B.n714 585
R415 B.n714 B.n713 585
R416 B.n716 B.n364 585
R417 B.n364 B.n363 585
R418 B.n718 B.n717 585
R419 B.n719 B.n718 585
R420 B.n358 B.n357 585
R421 B.n359 B.n358 585
R422 B.n727 B.n726 585
R423 B.n726 B.n725 585
R424 B.n728 B.n356 585
R425 B.n356 B.n354 585
R426 B.n730 B.n729 585
R427 B.n731 B.n730 585
R428 B.n350 B.n349 585
R429 B.n355 B.n350 585
R430 B.n739 B.n738 585
R431 B.n738 B.n737 585
R432 B.n740 B.n348 585
R433 B.n348 B.n347 585
R434 B.n742 B.n741 585
R435 B.n743 B.n742 585
R436 B.n342 B.n341 585
R437 B.n343 B.n342 585
R438 B.n752 B.n751 585
R439 B.n751 B.n750 585
R440 B.n753 B.n340 585
R441 B.n749 B.n340 585
R442 B.n755 B.n754 585
R443 B.n756 B.n755 585
R444 B.n335 B.n334 585
R445 B.n336 B.n335 585
R446 B.n764 B.n763 585
R447 B.n763 B.n762 585
R448 B.n765 B.n333 585
R449 B.n333 B.n331 585
R450 B.n767 B.n766 585
R451 B.n768 B.n767 585
R452 B.n327 B.n326 585
R453 B.n332 B.n327 585
R454 B.n777 B.n776 585
R455 B.n776 B.n775 585
R456 B.n778 B.n325 585
R457 B.n325 B.n324 585
R458 B.n780 B.n779 585
R459 B.n781 B.n780 585
R460 B.n2 B.n0 585
R461 B.n4 B.n2 585
R462 B.n3 B.n1 585
R463 B.n934 B.n3 585
R464 B.n932 B.n931 585
R465 B.n933 B.n932 585
R466 B.n930 B.n9 585
R467 B.n9 B.n8 585
R468 B.n929 B.n928 585
R469 B.n928 B.n927 585
R470 B.n11 B.n10 585
R471 B.n926 B.n11 585
R472 B.n924 B.n923 585
R473 B.n925 B.n924 585
R474 B.n922 B.n16 585
R475 B.n16 B.n15 585
R476 B.n921 B.n920 585
R477 B.n920 B.n919 585
R478 B.n18 B.n17 585
R479 B.n918 B.n18 585
R480 B.n916 B.n915 585
R481 B.n917 B.n916 585
R482 B.n914 B.n22 585
R483 B.n25 B.n22 585
R484 B.n913 B.n912 585
R485 B.n912 B.n911 585
R486 B.n24 B.n23 585
R487 B.n910 B.n24 585
R488 B.n908 B.n907 585
R489 B.n909 B.n908 585
R490 B.n906 B.n30 585
R491 B.n30 B.n29 585
R492 B.n905 B.n904 585
R493 B.n904 B.n903 585
R494 B.n32 B.n31 585
R495 B.n902 B.n32 585
R496 B.n900 B.n899 585
R497 B.n901 B.n900 585
R498 B.n898 B.n37 585
R499 B.n37 B.n36 585
R500 B.n897 B.n896 585
R501 B.n896 B.n895 585
R502 B.n39 B.n38 585
R503 B.n894 B.n39 585
R504 B.n892 B.n891 585
R505 B.n893 B.n892 585
R506 B.n890 B.n44 585
R507 B.n44 B.n43 585
R508 B.n889 B.n888 585
R509 B.n888 B.n887 585
R510 B.n46 B.n45 585
R511 B.n886 B.n46 585
R512 B.n884 B.n883 585
R513 B.n885 B.n884 585
R514 B.n882 B.n51 585
R515 B.n51 B.n50 585
R516 B.n881 B.n880 585
R517 B.n880 B.n879 585
R518 B.n53 B.n52 585
R519 B.n878 B.n53 585
R520 B.n876 B.n875 585
R521 B.n877 B.n876 585
R522 B.n874 B.n58 585
R523 B.n58 B.n57 585
R524 B.n873 B.n872 585
R525 B.n872 B.n871 585
R526 B.n60 B.n59 585
R527 B.n870 B.n60 585
R528 B.n868 B.n867 585
R529 B.n869 B.n868 585
R530 B.n866 B.n65 585
R531 B.n65 B.n64 585
R532 B.n865 B.n864 585
R533 B.n864 B.n863 585
R534 B.n67 B.n66 585
R535 B.n862 B.n67 585
R536 B.n860 B.n859 585
R537 B.n861 B.n860 585
R538 B.n858 B.n71 585
R539 B.n74 B.n71 585
R540 B.n857 B.n856 585
R541 B.n856 B.n855 585
R542 B.n73 B.n72 585
R543 B.n854 B.n73 585
R544 B.n852 B.n851 585
R545 B.n853 B.n852 585
R546 B.n850 B.n79 585
R547 B.n79 B.n78 585
R548 B.n849 B.n848 585
R549 B.n848 B.n847 585
R550 B.n81 B.n80 585
R551 B.n846 B.n81 585
R552 B.n937 B.n936 585
R553 B.n936 B.n935 585
R554 B.n644 B.n405 463.671
R555 B.n137 B.n81 463.671
R556 B.n647 B.n407 463.671
R557 B.n843 B.n83 463.671
R558 B.n459 B.t10 374.137
R559 B.n457 B.t18 374.137
R560 B.n134 B.t14 374.137
R561 B.n131 B.t21 374.137
R562 B.n459 B.t13 326.033
R563 B.n131 B.t22 326.033
R564 B.n457 B.t20 326.033
R565 B.n134 B.t16 326.033
R566 B.n460 B.t12 285.693
R567 B.n132 B.t23 285.693
R568 B.n458 B.t19 285.692
R569 B.n135 B.t17 285.692
R570 B.n845 B.n844 256.663
R571 B.n845 B.n129 256.663
R572 B.n845 B.n128 256.663
R573 B.n845 B.n127 256.663
R574 B.n845 B.n126 256.663
R575 B.n845 B.n125 256.663
R576 B.n845 B.n124 256.663
R577 B.n845 B.n123 256.663
R578 B.n845 B.n122 256.663
R579 B.n845 B.n121 256.663
R580 B.n845 B.n120 256.663
R581 B.n845 B.n119 256.663
R582 B.n845 B.n118 256.663
R583 B.n845 B.n117 256.663
R584 B.n845 B.n116 256.663
R585 B.n845 B.n115 256.663
R586 B.n845 B.n114 256.663
R587 B.n845 B.n113 256.663
R588 B.n845 B.n112 256.663
R589 B.n845 B.n111 256.663
R590 B.n845 B.n110 256.663
R591 B.n845 B.n109 256.663
R592 B.n845 B.n108 256.663
R593 B.n845 B.n107 256.663
R594 B.n845 B.n106 256.663
R595 B.n845 B.n105 256.663
R596 B.n845 B.n104 256.663
R597 B.n845 B.n103 256.663
R598 B.n845 B.n102 256.663
R599 B.n845 B.n101 256.663
R600 B.n845 B.n100 256.663
R601 B.n845 B.n99 256.663
R602 B.n845 B.n98 256.663
R603 B.n845 B.n97 256.663
R604 B.n845 B.n96 256.663
R605 B.n845 B.n95 256.663
R606 B.n845 B.n94 256.663
R607 B.n845 B.n93 256.663
R608 B.n845 B.n92 256.663
R609 B.n845 B.n91 256.663
R610 B.n845 B.n90 256.663
R611 B.n845 B.n89 256.663
R612 B.n845 B.n88 256.663
R613 B.n845 B.n87 256.663
R614 B.n845 B.n86 256.663
R615 B.n845 B.n85 256.663
R616 B.n845 B.n84 256.663
R617 B.n646 B.n645 256.663
R618 B.n646 B.n410 256.663
R619 B.n646 B.n411 256.663
R620 B.n646 B.n412 256.663
R621 B.n646 B.n413 256.663
R622 B.n646 B.n414 256.663
R623 B.n646 B.n415 256.663
R624 B.n646 B.n416 256.663
R625 B.n646 B.n417 256.663
R626 B.n646 B.n418 256.663
R627 B.n646 B.n419 256.663
R628 B.n646 B.n420 256.663
R629 B.n646 B.n421 256.663
R630 B.n646 B.n422 256.663
R631 B.n646 B.n423 256.663
R632 B.n646 B.n424 256.663
R633 B.n646 B.n425 256.663
R634 B.n646 B.n426 256.663
R635 B.n646 B.n427 256.663
R636 B.n646 B.n428 256.663
R637 B.n646 B.n429 256.663
R638 B.n646 B.n430 256.663
R639 B.n646 B.n431 256.663
R640 B.n646 B.n432 256.663
R641 B.n646 B.n433 256.663
R642 B.n646 B.n434 256.663
R643 B.n646 B.n435 256.663
R644 B.n646 B.n436 256.663
R645 B.n646 B.n437 256.663
R646 B.n646 B.n438 256.663
R647 B.n646 B.n439 256.663
R648 B.n646 B.n440 256.663
R649 B.n646 B.n441 256.663
R650 B.n646 B.n442 256.663
R651 B.n646 B.n443 256.663
R652 B.n646 B.n444 256.663
R653 B.n646 B.n445 256.663
R654 B.n646 B.n446 256.663
R655 B.n646 B.n447 256.663
R656 B.n646 B.n448 256.663
R657 B.n646 B.n449 256.663
R658 B.n646 B.n450 256.663
R659 B.n646 B.n451 256.663
R660 B.n646 B.n452 256.663
R661 B.n646 B.n453 256.663
R662 B.n646 B.n454 256.663
R663 B.n653 B.n405 163.367
R664 B.n653 B.n403 163.367
R665 B.n657 B.n403 163.367
R666 B.n657 B.n397 163.367
R667 B.n666 B.n397 163.367
R668 B.n666 B.n395 163.367
R669 B.n670 B.n395 163.367
R670 B.n670 B.n390 163.367
R671 B.n678 B.n390 163.367
R672 B.n678 B.n388 163.367
R673 B.n682 B.n388 163.367
R674 B.n682 B.n382 163.367
R675 B.n690 B.n382 163.367
R676 B.n690 B.n380 163.367
R677 B.n694 B.n380 163.367
R678 B.n694 B.n374 163.367
R679 B.n702 B.n374 163.367
R680 B.n702 B.n372 163.367
R681 B.n706 B.n372 163.367
R682 B.n706 B.n366 163.367
R683 B.n714 B.n366 163.367
R684 B.n714 B.n364 163.367
R685 B.n718 B.n364 163.367
R686 B.n718 B.n358 163.367
R687 B.n726 B.n358 163.367
R688 B.n726 B.n356 163.367
R689 B.n730 B.n356 163.367
R690 B.n730 B.n350 163.367
R691 B.n738 B.n350 163.367
R692 B.n738 B.n348 163.367
R693 B.n742 B.n348 163.367
R694 B.n742 B.n342 163.367
R695 B.n751 B.n342 163.367
R696 B.n751 B.n340 163.367
R697 B.n755 B.n340 163.367
R698 B.n755 B.n335 163.367
R699 B.n763 B.n335 163.367
R700 B.n763 B.n333 163.367
R701 B.n767 B.n333 163.367
R702 B.n767 B.n327 163.367
R703 B.n776 B.n327 163.367
R704 B.n776 B.n325 163.367
R705 B.n780 B.n325 163.367
R706 B.n780 B.n2 163.367
R707 B.n936 B.n2 163.367
R708 B.n936 B.n3 163.367
R709 B.n932 B.n3 163.367
R710 B.n932 B.n9 163.367
R711 B.n928 B.n9 163.367
R712 B.n928 B.n11 163.367
R713 B.n924 B.n11 163.367
R714 B.n924 B.n16 163.367
R715 B.n920 B.n16 163.367
R716 B.n920 B.n18 163.367
R717 B.n916 B.n18 163.367
R718 B.n916 B.n22 163.367
R719 B.n912 B.n22 163.367
R720 B.n912 B.n24 163.367
R721 B.n908 B.n24 163.367
R722 B.n908 B.n30 163.367
R723 B.n904 B.n30 163.367
R724 B.n904 B.n32 163.367
R725 B.n900 B.n32 163.367
R726 B.n900 B.n37 163.367
R727 B.n896 B.n37 163.367
R728 B.n896 B.n39 163.367
R729 B.n892 B.n39 163.367
R730 B.n892 B.n44 163.367
R731 B.n888 B.n44 163.367
R732 B.n888 B.n46 163.367
R733 B.n884 B.n46 163.367
R734 B.n884 B.n51 163.367
R735 B.n880 B.n51 163.367
R736 B.n880 B.n53 163.367
R737 B.n876 B.n53 163.367
R738 B.n876 B.n58 163.367
R739 B.n872 B.n58 163.367
R740 B.n872 B.n60 163.367
R741 B.n868 B.n60 163.367
R742 B.n868 B.n65 163.367
R743 B.n864 B.n65 163.367
R744 B.n864 B.n67 163.367
R745 B.n860 B.n67 163.367
R746 B.n860 B.n71 163.367
R747 B.n856 B.n71 163.367
R748 B.n856 B.n73 163.367
R749 B.n852 B.n73 163.367
R750 B.n852 B.n79 163.367
R751 B.n848 B.n79 163.367
R752 B.n848 B.n81 163.367
R753 B.n456 B.n455 163.367
R754 B.n639 B.n455 163.367
R755 B.n637 B.n636 163.367
R756 B.n633 B.n632 163.367
R757 B.n629 B.n628 163.367
R758 B.n625 B.n624 163.367
R759 B.n621 B.n620 163.367
R760 B.n617 B.n616 163.367
R761 B.n613 B.n612 163.367
R762 B.n609 B.n608 163.367
R763 B.n605 B.n604 163.367
R764 B.n601 B.n600 163.367
R765 B.n597 B.n596 163.367
R766 B.n593 B.n592 163.367
R767 B.n589 B.n588 163.367
R768 B.n585 B.n584 163.367
R769 B.n581 B.n580 163.367
R770 B.n577 B.n576 163.367
R771 B.n573 B.n572 163.367
R772 B.n569 B.n568 163.367
R773 B.n565 B.n564 163.367
R774 B.n560 B.n559 163.367
R775 B.n556 B.n555 163.367
R776 B.n552 B.n551 163.367
R777 B.n548 B.n547 163.367
R778 B.n544 B.n543 163.367
R779 B.n539 B.n538 163.367
R780 B.n535 B.n534 163.367
R781 B.n531 B.n530 163.367
R782 B.n527 B.n526 163.367
R783 B.n523 B.n522 163.367
R784 B.n519 B.n518 163.367
R785 B.n515 B.n514 163.367
R786 B.n511 B.n510 163.367
R787 B.n507 B.n506 163.367
R788 B.n503 B.n502 163.367
R789 B.n499 B.n498 163.367
R790 B.n495 B.n494 163.367
R791 B.n491 B.n490 163.367
R792 B.n487 B.n486 163.367
R793 B.n483 B.n482 163.367
R794 B.n479 B.n478 163.367
R795 B.n475 B.n474 163.367
R796 B.n471 B.n470 163.367
R797 B.n467 B.n466 163.367
R798 B.n463 B.n462 163.367
R799 B.n647 B.n409 163.367
R800 B.n651 B.n407 163.367
R801 B.n651 B.n401 163.367
R802 B.n659 B.n401 163.367
R803 B.n659 B.n399 163.367
R804 B.n663 B.n399 163.367
R805 B.n663 B.n394 163.367
R806 B.n672 B.n394 163.367
R807 B.n672 B.n392 163.367
R808 B.n676 B.n392 163.367
R809 B.n676 B.n386 163.367
R810 B.n684 B.n386 163.367
R811 B.n684 B.n384 163.367
R812 B.n688 B.n384 163.367
R813 B.n688 B.n378 163.367
R814 B.n696 B.n378 163.367
R815 B.n696 B.n376 163.367
R816 B.n700 B.n376 163.367
R817 B.n700 B.n370 163.367
R818 B.n708 B.n370 163.367
R819 B.n708 B.n368 163.367
R820 B.n712 B.n368 163.367
R821 B.n712 B.n362 163.367
R822 B.n720 B.n362 163.367
R823 B.n720 B.n360 163.367
R824 B.n724 B.n360 163.367
R825 B.n724 B.n353 163.367
R826 B.n732 B.n353 163.367
R827 B.n732 B.n351 163.367
R828 B.n736 B.n351 163.367
R829 B.n736 B.n346 163.367
R830 B.n744 B.n346 163.367
R831 B.n744 B.n344 163.367
R832 B.n748 B.n344 163.367
R833 B.n748 B.n339 163.367
R834 B.n757 B.n339 163.367
R835 B.n757 B.n337 163.367
R836 B.n761 B.n337 163.367
R837 B.n761 B.n330 163.367
R838 B.n769 B.n330 163.367
R839 B.n769 B.n328 163.367
R840 B.n774 B.n328 163.367
R841 B.n774 B.n323 163.367
R842 B.n782 B.n323 163.367
R843 B.n783 B.n782 163.367
R844 B.n783 B.n5 163.367
R845 B.n6 B.n5 163.367
R846 B.n7 B.n6 163.367
R847 B.n788 B.n7 163.367
R848 B.n788 B.n12 163.367
R849 B.n13 B.n12 163.367
R850 B.n14 B.n13 163.367
R851 B.n793 B.n14 163.367
R852 B.n793 B.n19 163.367
R853 B.n20 B.n19 163.367
R854 B.n21 B.n20 163.367
R855 B.n798 B.n21 163.367
R856 B.n798 B.n26 163.367
R857 B.n27 B.n26 163.367
R858 B.n28 B.n27 163.367
R859 B.n803 B.n28 163.367
R860 B.n803 B.n33 163.367
R861 B.n34 B.n33 163.367
R862 B.n35 B.n34 163.367
R863 B.n808 B.n35 163.367
R864 B.n808 B.n40 163.367
R865 B.n41 B.n40 163.367
R866 B.n42 B.n41 163.367
R867 B.n813 B.n42 163.367
R868 B.n813 B.n47 163.367
R869 B.n48 B.n47 163.367
R870 B.n49 B.n48 163.367
R871 B.n818 B.n49 163.367
R872 B.n818 B.n54 163.367
R873 B.n55 B.n54 163.367
R874 B.n56 B.n55 163.367
R875 B.n823 B.n56 163.367
R876 B.n823 B.n61 163.367
R877 B.n62 B.n61 163.367
R878 B.n63 B.n62 163.367
R879 B.n828 B.n63 163.367
R880 B.n828 B.n68 163.367
R881 B.n69 B.n68 163.367
R882 B.n70 B.n69 163.367
R883 B.n833 B.n70 163.367
R884 B.n833 B.n75 163.367
R885 B.n76 B.n75 163.367
R886 B.n77 B.n76 163.367
R887 B.n838 B.n77 163.367
R888 B.n838 B.n82 163.367
R889 B.n83 B.n82 163.367
R890 B.n141 B.n140 163.367
R891 B.n145 B.n144 163.367
R892 B.n149 B.n148 163.367
R893 B.n153 B.n152 163.367
R894 B.n157 B.n156 163.367
R895 B.n161 B.n160 163.367
R896 B.n165 B.n164 163.367
R897 B.n169 B.n168 163.367
R898 B.n173 B.n172 163.367
R899 B.n177 B.n176 163.367
R900 B.n181 B.n180 163.367
R901 B.n185 B.n184 163.367
R902 B.n189 B.n188 163.367
R903 B.n193 B.n192 163.367
R904 B.n197 B.n196 163.367
R905 B.n201 B.n200 163.367
R906 B.n205 B.n204 163.367
R907 B.n209 B.n208 163.367
R908 B.n213 B.n212 163.367
R909 B.n217 B.n216 163.367
R910 B.n221 B.n220 163.367
R911 B.n225 B.n224 163.367
R912 B.n229 B.n228 163.367
R913 B.n233 B.n232 163.367
R914 B.n237 B.n236 163.367
R915 B.n241 B.n240 163.367
R916 B.n245 B.n244 163.367
R917 B.n249 B.n248 163.367
R918 B.n253 B.n252 163.367
R919 B.n257 B.n256 163.367
R920 B.n261 B.n260 163.367
R921 B.n265 B.n264 163.367
R922 B.n269 B.n268 163.367
R923 B.n273 B.n272 163.367
R924 B.n277 B.n276 163.367
R925 B.n281 B.n280 163.367
R926 B.n285 B.n284 163.367
R927 B.n289 B.n288 163.367
R928 B.n293 B.n292 163.367
R929 B.n297 B.n296 163.367
R930 B.n301 B.n300 163.367
R931 B.n305 B.n304 163.367
R932 B.n309 B.n308 163.367
R933 B.n313 B.n312 163.367
R934 B.n317 B.n316 163.367
R935 B.n319 B.n130 163.367
R936 B.n645 B.n644 71.676
R937 B.n639 B.n410 71.676
R938 B.n636 B.n411 71.676
R939 B.n632 B.n412 71.676
R940 B.n628 B.n413 71.676
R941 B.n624 B.n414 71.676
R942 B.n620 B.n415 71.676
R943 B.n616 B.n416 71.676
R944 B.n612 B.n417 71.676
R945 B.n608 B.n418 71.676
R946 B.n604 B.n419 71.676
R947 B.n600 B.n420 71.676
R948 B.n596 B.n421 71.676
R949 B.n592 B.n422 71.676
R950 B.n588 B.n423 71.676
R951 B.n584 B.n424 71.676
R952 B.n580 B.n425 71.676
R953 B.n576 B.n426 71.676
R954 B.n572 B.n427 71.676
R955 B.n568 B.n428 71.676
R956 B.n564 B.n429 71.676
R957 B.n559 B.n430 71.676
R958 B.n555 B.n431 71.676
R959 B.n551 B.n432 71.676
R960 B.n547 B.n433 71.676
R961 B.n543 B.n434 71.676
R962 B.n538 B.n435 71.676
R963 B.n534 B.n436 71.676
R964 B.n530 B.n437 71.676
R965 B.n526 B.n438 71.676
R966 B.n522 B.n439 71.676
R967 B.n518 B.n440 71.676
R968 B.n514 B.n441 71.676
R969 B.n510 B.n442 71.676
R970 B.n506 B.n443 71.676
R971 B.n502 B.n444 71.676
R972 B.n498 B.n445 71.676
R973 B.n494 B.n446 71.676
R974 B.n490 B.n447 71.676
R975 B.n486 B.n448 71.676
R976 B.n482 B.n449 71.676
R977 B.n478 B.n450 71.676
R978 B.n474 B.n451 71.676
R979 B.n470 B.n452 71.676
R980 B.n466 B.n453 71.676
R981 B.n462 B.n454 71.676
R982 B.n137 B.n84 71.676
R983 B.n141 B.n85 71.676
R984 B.n145 B.n86 71.676
R985 B.n149 B.n87 71.676
R986 B.n153 B.n88 71.676
R987 B.n157 B.n89 71.676
R988 B.n161 B.n90 71.676
R989 B.n165 B.n91 71.676
R990 B.n169 B.n92 71.676
R991 B.n173 B.n93 71.676
R992 B.n177 B.n94 71.676
R993 B.n181 B.n95 71.676
R994 B.n185 B.n96 71.676
R995 B.n189 B.n97 71.676
R996 B.n193 B.n98 71.676
R997 B.n197 B.n99 71.676
R998 B.n201 B.n100 71.676
R999 B.n205 B.n101 71.676
R1000 B.n209 B.n102 71.676
R1001 B.n213 B.n103 71.676
R1002 B.n217 B.n104 71.676
R1003 B.n221 B.n105 71.676
R1004 B.n225 B.n106 71.676
R1005 B.n229 B.n107 71.676
R1006 B.n233 B.n108 71.676
R1007 B.n237 B.n109 71.676
R1008 B.n241 B.n110 71.676
R1009 B.n245 B.n111 71.676
R1010 B.n249 B.n112 71.676
R1011 B.n253 B.n113 71.676
R1012 B.n257 B.n114 71.676
R1013 B.n261 B.n115 71.676
R1014 B.n265 B.n116 71.676
R1015 B.n269 B.n117 71.676
R1016 B.n273 B.n118 71.676
R1017 B.n277 B.n119 71.676
R1018 B.n281 B.n120 71.676
R1019 B.n285 B.n121 71.676
R1020 B.n289 B.n122 71.676
R1021 B.n293 B.n123 71.676
R1022 B.n297 B.n124 71.676
R1023 B.n301 B.n125 71.676
R1024 B.n305 B.n126 71.676
R1025 B.n309 B.n127 71.676
R1026 B.n313 B.n128 71.676
R1027 B.n317 B.n129 71.676
R1028 B.n844 B.n130 71.676
R1029 B.n844 B.n843 71.676
R1030 B.n319 B.n129 71.676
R1031 B.n316 B.n128 71.676
R1032 B.n312 B.n127 71.676
R1033 B.n308 B.n126 71.676
R1034 B.n304 B.n125 71.676
R1035 B.n300 B.n124 71.676
R1036 B.n296 B.n123 71.676
R1037 B.n292 B.n122 71.676
R1038 B.n288 B.n121 71.676
R1039 B.n284 B.n120 71.676
R1040 B.n280 B.n119 71.676
R1041 B.n276 B.n118 71.676
R1042 B.n272 B.n117 71.676
R1043 B.n268 B.n116 71.676
R1044 B.n264 B.n115 71.676
R1045 B.n260 B.n114 71.676
R1046 B.n256 B.n113 71.676
R1047 B.n252 B.n112 71.676
R1048 B.n248 B.n111 71.676
R1049 B.n244 B.n110 71.676
R1050 B.n240 B.n109 71.676
R1051 B.n236 B.n108 71.676
R1052 B.n232 B.n107 71.676
R1053 B.n228 B.n106 71.676
R1054 B.n224 B.n105 71.676
R1055 B.n220 B.n104 71.676
R1056 B.n216 B.n103 71.676
R1057 B.n212 B.n102 71.676
R1058 B.n208 B.n101 71.676
R1059 B.n204 B.n100 71.676
R1060 B.n200 B.n99 71.676
R1061 B.n196 B.n98 71.676
R1062 B.n192 B.n97 71.676
R1063 B.n188 B.n96 71.676
R1064 B.n184 B.n95 71.676
R1065 B.n180 B.n94 71.676
R1066 B.n176 B.n93 71.676
R1067 B.n172 B.n92 71.676
R1068 B.n168 B.n91 71.676
R1069 B.n164 B.n90 71.676
R1070 B.n160 B.n89 71.676
R1071 B.n156 B.n88 71.676
R1072 B.n152 B.n87 71.676
R1073 B.n148 B.n86 71.676
R1074 B.n144 B.n85 71.676
R1075 B.n140 B.n84 71.676
R1076 B.n645 B.n456 71.676
R1077 B.n637 B.n410 71.676
R1078 B.n633 B.n411 71.676
R1079 B.n629 B.n412 71.676
R1080 B.n625 B.n413 71.676
R1081 B.n621 B.n414 71.676
R1082 B.n617 B.n415 71.676
R1083 B.n613 B.n416 71.676
R1084 B.n609 B.n417 71.676
R1085 B.n605 B.n418 71.676
R1086 B.n601 B.n419 71.676
R1087 B.n597 B.n420 71.676
R1088 B.n593 B.n421 71.676
R1089 B.n589 B.n422 71.676
R1090 B.n585 B.n423 71.676
R1091 B.n581 B.n424 71.676
R1092 B.n577 B.n425 71.676
R1093 B.n573 B.n426 71.676
R1094 B.n569 B.n427 71.676
R1095 B.n565 B.n428 71.676
R1096 B.n560 B.n429 71.676
R1097 B.n556 B.n430 71.676
R1098 B.n552 B.n431 71.676
R1099 B.n548 B.n432 71.676
R1100 B.n544 B.n433 71.676
R1101 B.n539 B.n434 71.676
R1102 B.n535 B.n435 71.676
R1103 B.n531 B.n436 71.676
R1104 B.n527 B.n437 71.676
R1105 B.n523 B.n438 71.676
R1106 B.n519 B.n439 71.676
R1107 B.n515 B.n440 71.676
R1108 B.n511 B.n441 71.676
R1109 B.n507 B.n442 71.676
R1110 B.n503 B.n443 71.676
R1111 B.n499 B.n444 71.676
R1112 B.n495 B.n445 71.676
R1113 B.n491 B.n446 71.676
R1114 B.n487 B.n447 71.676
R1115 B.n483 B.n448 71.676
R1116 B.n479 B.n449 71.676
R1117 B.n475 B.n450 71.676
R1118 B.n471 B.n451 71.676
R1119 B.n467 B.n452 71.676
R1120 B.n463 B.n453 71.676
R1121 B.n454 B.n409 71.676
R1122 B.n646 B.n406 69.9117
R1123 B.n846 B.n845 69.9117
R1124 B.n541 B.n460 59.5399
R1125 B.n562 B.n458 59.5399
R1126 B.n136 B.n135 59.5399
R1127 B.n133 B.n132 59.5399
R1128 B.n652 B.n406 42.829
R1129 B.n652 B.n402 42.829
R1130 B.n658 B.n402 42.829
R1131 B.n658 B.n398 42.829
R1132 B.n665 B.n398 42.829
R1133 B.n665 B.n664 42.829
R1134 B.n671 B.n391 42.829
R1135 B.n677 B.n391 42.829
R1136 B.n677 B.n387 42.829
R1137 B.n683 B.n387 42.829
R1138 B.n683 B.n383 42.829
R1139 B.n689 B.n383 42.829
R1140 B.n689 B.n379 42.829
R1141 B.n695 B.n379 42.829
R1142 B.n701 B.n375 42.829
R1143 B.n701 B.n371 42.829
R1144 B.n707 B.n371 42.829
R1145 B.n707 B.n367 42.829
R1146 B.n713 B.n367 42.829
R1147 B.n719 B.n363 42.829
R1148 B.n719 B.n359 42.829
R1149 B.n725 B.n359 42.829
R1150 B.n725 B.n354 42.829
R1151 B.n731 B.n354 42.829
R1152 B.n731 B.n355 42.829
R1153 B.n737 B.n347 42.829
R1154 B.n743 B.n347 42.829
R1155 B.n743 B.n343 42.829
R1156 B.n750 B.n343 42.829
R1157 B.n750 B.n749 42.829
R1158 B.n756 B.n336 42.829
R1159 B.n762 B.n336 42.829
R1160 B.n762 B.n331 42.829
R1161 B.n768 B.n331 42.829
R1162 B.n768 B.n332 42.829
R1163 B.n775 B.n324 42.829
R1164 B.n781 B.n324 42.829
R1165 B.n781 B.n4 42.829
R1166 B.n935 B.n4 42.829
R1167 B.n935 B.n934 42.829
R1168 B.n934 B.n933 42.829
R1169 B.n933 B.n8 42.829
R1170 B.n927 B.n8 42.829
R1171 B.n926 B.n925 42.829
R1172 B.n925 B.n15 42.829
R1173 B.n919 B.n15 42.829
R1174 B.n919 B.n918 42.829
R1175 B.n918 B.n917 42.829
R1176 B.n911 B.n25 42.829
R1177 B.n911 B.n910 42.829
R1178 B.n910 B.n909 42.829
R1179 B.n909 B.n29 42.829
R1180 B.n903 B.n29 42.829
R1181 B.n902 B.n901 42.829
R1182 B.n901 B.n36 42.829
R1183 B.n895 B.n36 42.829
R1184 B.n895 B.n894 42.829
R1185 B.n894 B.n893 42.829
R1186 B.n893 B.n43 42.829
R1187 B.n887 B.n886 42.829
R1188 B.n886 B.n885 42.829
R1189 B.n885 B.n50 42.829
R1190 B.n879 B.n50 42.829
R1191 B.n879 B.n878 42.829
R1192 B.n877 B.n57 42.829
R1193 B.n871 B.n57 42.829
R1194 B.n871 B.n870 42.829
R1195 B.n870 B.n869 42.829
R1196 B.n869 B.n64 42.829
R1197 B.n863 B.n64 42.829
R1198 B.n863 B.n862 42.829
R1199 B.n862 B.n861 42.829
R1200 B.n855 B.n74 42.829
R1201 B.n855 B.n854 42.829
R1202 B.n854 B.n853 42.829
R1203 B.n853 B.n78 42.829
R1204 B.n847 B.n78 42.829
R1205 B.n847 B.n846 42.829
R1206 B.n713 B.t6 42.1992
R1207 B.n887 B.t3 42.1992
R1208 B.n460 B.n459 40.3399
R1209 B.n458 B.n457 40.3399
R1210 B.n135 B.n134 40.3399
R1211 B.n132 B.n131 40.3399
R1212 B.n737 B.t1 38.4202
R1213 B.n903 B.t2 38.4202
R1214 B.n695 B.t8 37.1605
R1215 B.t5 B.n877 37.1605
R1216 B.n756 B.t9 33.3815
R1217 B.n917 B.t0 33.3815
R1218 B.n138 B.n80 30.1273
R1219 B.n649 B.n648 30.1273
R1220 B.n643 B.n404 30.1273
R1221 B.n842 B.n841 30.1273
R1222 B.n775 B.t4 28.3429
R1223 B.n927 B.t7 28.3429
R1224 B.n664 B.t11 23.3042
R1225 B.n74 B.t15 23.3042
R1226 B.n671 B.t11 19.5253
R1227 B.n861 B.t15 19.5253
R1228 B B.n937 18.0485
R1229 B.n332 B.t4 14.4866
R1230 B.t7 B.n926 14.4866
R1231 B.n139 B.n138 10.6151
R1232 B.n142 B.n139 10.6151
R1233 B.n143 B.n142 10.6151
R1234 B.n146 B.n143 10.6151
R1235 B.n147 B.n146 10.6151
R1236 B.n150 B.n147 10.6151
R1237 B.n151 B.n150 10.6151
R1238 B.n154 B.n151 10.6151
R1239 B.n155 B.n154 10.6151
R1240 B.n158 B.n155 10.6151
R1241 B.n159 B.n158 10.6151
R1242 B.n162 B.n159 10.6151
R1243 B.n163 B.n162 10.6151
R1244 B.n166 B.n163 10.6151
R1245 B.n167 B.n166 10.6151
R1246 B.n170 B.n167 10.6151
R1247 B.n171 B.n170 10.6151
R1248 B.n174 B.n171 10.6151
R1249 B.n175 B.n174 10.6151
R1250 B.n178 B.n175 10.6151
R1251 B.n179 B.n178 10.6151
R1252 B.n182 B.n179 10.6151
R1253 B.n183 B.n182 10.6151
R1254 B.n186 B.n183 10.6151
R1255 B.n187 B.n186 10.6151
R1256 B.n190 B.n187 10.6151
R1257 B.n191 B.n190 10.6151
R1258 B.n194 B.n191 10.6151
R1259 B.n195 B.n194 10.6151
R1260 B.n198 B.n195 10.6151
R1261 B.n199 B.n198 10.6151
R1262 B.n202 B.n199 10.6151
R1263 B.n203 B.n202 10.6151
R1264 B.n206 B.n203 10.6151
R1265 B.n207 B.n206 10.6151
R1266 B.n210 B.n207 10.6151
R1267 B.n211 B.n210 10.6151
R1268 B.n214 B.n211 10.6151
R1269 B.n215 B.n214 10.6151
R1270 B.n218 B.n215 10.6151
R1271 B.n219 B.n218 10.6151
R1272 B.n223 B.n222 10.6151
R1273 B.n226 B.n223 10.6151
R1274 B.n227 B.n226 10.6151
R1275 B.n230 B.n227 10.6151
R1276 B.n231 B.n230 10.6151
R1277 B.n234 B.n231 10.6151
R1278 B.n235 B.n234 10.6151
R1279 B.n238 B.n235 10.6151
R1280 B.n239 B.n238 10.6151
R1281 B.n243 B.n242 10.6151
R1282 B.n246 B.n243 10.6151
R1283 B.n247 B.n246 10.6151
R1284 B.n250 B.n247 10.6151
R1285 B.n251 B.n250 10.6151
R1286 B.n254 B.n251 10.6151
R1287 B.n255 B.n254 10.6151
R1288 B.n258 B.n255 10.6151
R1289 B.n259 B.n258 10.6151
R1290 B.n262 B.n259 10.6151
R1291 B.n263 B.n262 10.6151
R1292 B.n266 B.n263 10.6151
R1293 B.n267 B.n266 10.6151
R1294 B.n270 B.n267 10.6151
R1295 B.n271 B.n270 10.6151
R1296 B.n274 B.n271 10.6151
R1297 B.n275 B.n274 10.6151
R1298 B.n278 B.n275 10.6151
R1299 B.n279 B.n278 10.6151
R1300 B.n282 B.n279 10.6151
R1301 B.n283 B.n282 10.6151
R1302 B.n286 B.n283 10.6151
R1303 B.n287 B.n286 10.6151
R1304 B.n290 B.n287 10.6151
R1305 B.n291 B.n290 10.6151
R1306 B.n294 B.n291 10.6151
R1307 B.n295 B.n294 10.6151
R1308 B.n298 B.n295 10.6151
R1309 B.n299 B.n298 10.6151
R1310 B.n302 B.n299 10.6151
R1311 B.n303 B.n302 10.6151
R1312 B.n306 B.n303 10.6151
R1313 B.n307 B.n306 10.6151
R1314 B.n310 B.n307 10.6151
R1315 B.n311 B.n310 10.6151
R1316 B.n314 B.n311 10.6151
R1317 B.n315 B.n314 10.6151
R1318 B.n318 B.n315 10.6151
R1319 B.n320 B.n318 10.6151
R1320 B.n321 B.n320 10.6151
R1321 B.n842 B.n321 10.6151
R1322 B.n650 B.n649 10.6151
R1323 B.n650 B.n400 10.6151
R1324 B.n660 B.n400 10.6151
R1325 B.n661 B.n660 10.6151
R1326 B.n662 B.n661 10.6151
R1327 B.n662 B.n393 10.6151
R1328 B.n673 B.n393 10.6151
R1329 B.n674 B.n673 10.6151
R1330 B.n675 B.n674 10.6151
R1331 B.n675 B.n385 10.6151
R1332 B.n685 B.n385 10.6151
R1333 B.n686 B.n685 10.6151
R1334 B.n687 B.n686 10.6151
R1335 B.n687 B.n377 10.6151
R1336 B.n697 B.n377 10.6151
R1337 B.n698 B.n697 10.6151
R1338 B.n699 B.n698 10.6151
R1339 B.n699 B.n369 10.6151
R1340 B.n709 B.n369 10.6151
R1341 B.n710 B.n709 10.6151
R1342 B.n711 B.n710 10.6151
R1343 B.n711 B.n361 10.6151
R1344 B.n721 B.n361 10.6151
R1345 B.n722 B.n721 10.6151
R1346 B.n723 B.n722 10.6151
R1347 B.n723 B.n352 10.6151
R1348 B.n733 B.n352 10.6151
R1349 B.n734 B.n733 10.6151
R1350 B.n735 B.n734 10.6151
R1351 B.n735 B.n345 10.6151
R1352 B.n745 B.n345 10.6151
R1353 B.n746 B.n745 10.6151
R1354 B.n747 B.n746 10.6151
R1355 B.n747 B.n338 10.6151
R1356 B.n758 B.n338 10.6151
R1357 B.n759 B.n758 10.6151
R1358 B.n760 B.n759 10.6151
R1359 B.n760 B.n329 10.6151
R1360 B.n770 B.n329 10.6151
R1361 B.n771 B.n770 10.6151
R1362 B.n773 B.n771 10.6151
R1363 B.n773 B.n772 10.6151
R1364 B.n772 B.n322 10.6151
R1365 B.n784 B.n322 10.6151
R1366 B.n785 B.n784 10.6151
R1367 B.n786 B.n785 10.6151
R1368 B.n787 B.n786 10.6151
R1369 B.n789 B.n787 10.6151
R1370 B.n790 B.n789 10.6151
R1371 B.n791 B.n790 10.6151
R1372 B.n792 B.n791 10.6151
R1373 B.n794 B.n792 10.6151
R1374 B.n795 B.n794 10.6151
R1375 B.n796 B.n795 10.6151
R1376 B.n797 B.n796 10.6151
R1377 B.n799 B.n797 10.6151
R1378 B.n800 B.n799 10.6151
R1379 B.n801 B.n800 10.6151
R1380 B.n802 B.n801 10.6151
R1381 B.n804 B.n802 10.6151
R1382 B.n805 B.n804 10.6151
R1383 B.n806 B.n805 10.6151
R1384 B.n807 B.n806 10.6151
R1385 B.n809 B.n807 10.6151
R1386 B.n810 B.n809 10.6151
R1387 B.n811 B.n810 10.6151
R1388 B.n812 B.n811 10.6151
R1389 B.n814 B.n812 10.6151
R1390 B.n815 B.n814 10.6151
R1391 B.n816 B.n815 10.6151
R1392 B.n817 B.n816 10.6151
R1393 B.n819 B.n817 10.6151
R1394 B.n820 B.n819 10.6151
R1395 B.n821 B.n820 10.6151
R1396 B.n822 B.n821 10.6151
R1397 B.n824 B.n822 10.6151
R1398 B.n825 B.n824 10.6151
R1399 B.n826 B.n825 10.6151
R1400 B.n827 B.n826 10.6151
R1401 B.n829 B.n827 10.6151
R1402 B.n830 B.n829 10.6151
R1403 B.n831 B.n830 10.6151
R1404 B.n832 B.n831 10.6151
R1405 B.n834 B.n832 10.6151
R1406 B.n835 B.n834 10.6151
R1407 B.n836 B.n835 10.6151
R1408 B.n837 B.n836 10.6151
R1409 B.n839 B.n837 10.6151
R1410 B.n840 B.n839 10.6151
R1411 B.n841 B.n840 10.6151
R1412 B.n643 B.n642 10.6151
R1413 B.n642 B.n641 10.6151
R1414 B.n641 B.n640 10.6151
R1415 B.n640 B.n638 10.6151
R1416 B.n638 B.n635 10.6151
R1417 B.n635 B.n634 10.6151
R1418 B.n634 B.n631 10.6151
R1419 B.n631 B.n630 10.6151
R1420 B.n630 B.n627 10.6151
R1421 B.n627 B.n626 10.6151
R1422 B.n626 B.n623 10.6151
R1423 B.n623 B.n622 10.6151
R1424 B.n622 B.n619 10.6151
R1425 B.n619 B.n618 10.6151
R1426 B.n618 B.n615 10.6151
R1427 B.n615 B.n614 10.6151
R1428 B.n614 B.n611 10.6151
R1429 B.n611 B.n610 10.6151
R1430 B.n610 B.n607 10.6151
R1431 B.n607 B.n606 10.6151
R1432 B.n606 B.n603 10.6151
R1433 B.n603 B.n602 10.6151
R1434 B.n602 B.n599 10.6151
R1435 B.n599 B.n598 10.6151
R1436 B.n598 B.n595 10.6151
R1437 B.n595 B.n594 10.6151
R1438 B.n594 B.n591 10.6151
R1439 B.n591 B.n590 10.6151
R1440 B.n590 B.n587 10.6151
R1441 B.n587 B.n586 10.6151
R1442 B.n586 B.n583 10.6151
R1443 B.n583 B.n582 10.6151
R1444 B.n582 B.n579 10.6151
R1445 B.n579 B.n578 10.6151
R1446 B.n578 B.n575 10.6151
R1447 B.n575 B.n574 10.6151
R1448 B.n574 B.n571 10.6151
R1449 B.n571 B.n570 10.6151
R1450 B.n570 B.n567 10.6151
R1451 B.n567 B.n566 10.6151
R1452 B.n566 B.n563 10.6151
R1453 B.n561 B.n558 10.6151
R1454 B.n558 B.n557 10.6151
R1455 B.n557 B.n554 10.6151
R1456 B.n554 B.n553 10.6151
R1457 B.n553 B.n550 10.6151
R1458 B.n550 B.n549 10.6151
R1459 B.n549 B.n546 10.6151
R1460 B.n546 B.n545 10.6151
R1461 B.n545 B.n542 10.6151
R1462 B.n540 B.n537 10.6151
R1463 B.n537 B.n536 10.6151
R1464 B.n536 B.n533 10.6151
R1465 B.n533 B.n532 10.6151
R1466 B.n532 B.n529 10.6151
R1467 B.n529 B.n528 10.6151
R1468 B.n528 B.n525 10.6151
R1469 B.n525 B.n524 10.6151
R1470 B.n524 B.n521 10.6151
R1471 B.n521 B.n520 10.6151
R1472 B.n520 B.n517 10.6151
R1473 B.n517 B.n516 10.6151
R1474 B.n516 B.n513 10.6151
R1475 B.n513 B.n512 10.6151
R1476 B.n512 B.n509 10.6151
R1477 B.n509 B.n508 10.6151
R1478 B.n508 B.n505 10.6151
R1479 B.n505 B.n504 10.6151
R1480 B.n504 B.n501 10.6151
R1481 B.n501 B.n500 10.6151
R1482 B.n500 B.n497 10.6151
R1483 B.n497 B.n496 10.6151
R1484 B.n496 B.n493 10.6151
R1485 B.n493 B.n492 10.6151
R1486 B.n492 B.n489 10.6151
R1487 B.n489 B.n488 10.6151
R1488 B.n488 B.n485 10.6151
R1489 B.n485 B.n484 10.6151
R1490 B.n484 B.n481 10.6151
R1491 B.n481 B.n480 10.6151
R1492 B.n480 B.n477 10.6151
R1493 B.n477 B.n476 10.6151
R1494 B.n476 B.n473 10.6151
R1495 B.n473 B.n472 10.6151
R1496 B.n472 B.n469 10.6151
R1497 B.n469 B.n468 10.6151
R1498 B.n468 B.n465 10.6151
R1499 B.n465 B.n464 10.6151
R1500 B.n464 B.n461 10.6151
R1501 B.n461 B.n408 10.6151
R1502 B.n648 B.n408 10.6151
R1503 B.n654 B.n404 10.6151
R1504 B.n655 B.n654 10.6151
R1505 B.n656 B.n655 10.6151
R1506 B.n656 B.n396 10.6151
R1507 B.n667 B.n396 10.6151
R1508 B.n668 B.n667 10.6151
R1509 B.n669 B.n668 10.6151
R1510 B.n669 B.n389 10.6151
R1511 B.n679 B.n389 10.6151
R1512 B.n680 B.n679 10.6151
R1513 B.n681 B.n680 10.6151
R1514 B.n681 B.n381 10.6151
R1515 B.n691 B.n381 10.6151
R1516 B.n692 B.n691 10.6151
R1517 B.n693 B.n692 10.6151
R1518 B.n693 B.n373 10.6151
R1519 B.n703 B.n373 10.6151
R1520 B.n704 B.n703 10.6151
R1521 B.n705 B.n704 10.6151
R1522 B.n705 B.n365 10.6151
R1523 B.n715 B.n365 10.6151
R1524 B.n716 B.n715 10.6151
R1525 B.n717 B.n716 10.6151
R1526 B.n717 B.n357 10.6151
R1527 B.n727 B.n357 10.6151
R1528 B.n728 B.n727 10.6151
R1529 B.n729 B.n728 10.6151
R1530 B.n729 B.n349 10.6151
R1531 B.n739 B.n349 10.6151
R1532 B.n740 B.n739 10.6151
R1533 B.n741 B.n740 10.6151
R1534 B.n741 B.n341 10.6151
R1535 B.n752 B.n341 10.6151
R1536 B.n753 B.n752 10.6151
R1537 B.n754 B.n753 10.6151
R1538 B.n754 B.n334 10.6151
R1539 B.n764 B.n334 10.6151
R1540 B.n765 B.n764 10.6151
R1541 B.n766 B.n765 10.6151
R1542 B.n766 B.n326 10.6151
R1543 B.n777 B.n326 10.6151
R1544 B.n778 B.n777 10.6151
R1545 B.n779 B.n778 10.6151
R1546 B.n779 B.n0 10.6151
R1547 B.n931 B.n1 10.6151
R1548 B.n931 B.n930 10.6151
R1549 B.n930 B.n929 10.6151
R1550 B.n929 B.n10 10.6151
R1551 B.n923 B.n10 10.6151
R1552 B.n923 B.n922 10.6151
R1553 B.n922 B.n921 10.6151
R1554 B.n921 B.n17 10.6151
R1555 B.n915 B.n17 10.6151
R1556 B.n915 B.n914 10.6151
R1557 B.n914 B.n913 10.6151
R1558 B.n913 B.n23 10.6151
R1559 B.n907 B.n23 10.6151
R1560 B.n907 B.n906 10.6151
R1561 B.n906 B.n905 10.6151
R1562 B.n905 B.n31 10.6151
R1563 B.n899 B.n31 10.6151
R1564 B.n899 B.n898 10.6151
R1565 B.n898 B.n897 10.6151
R1566 B.n897 B.n38 10.6151
R1567 B.n891 B.n38 10.6151
R1568 B.n891 B.n890 10.6151
R1569 B.n890 B.n889 10.6151
R1570 B.n889 B.n45 10.6151
R1571 B.n883 B.n45 10.6151
R1572 B.n883 B.n882 10.6151
R1573 B.n882 B.n881 10.6151
R1574 B.n881 B.n52 10.6151
R1575 B.n875 B.n52 10.6151
R1576 B.n875 B.n874 10.6151
R1577 B.n874 B.n873 10.6151
R1578 B.n873 B.n59 10.6151
R1579 B.n867 B.n59 10.6151
R1580 B.n867 B.n866 10.6151
R1581 B.n866 B.n865 10.6151
R1582 B.n865 B.n66 10.6151
R1583 B.n859 B.n66 10.6151
R1584 B.n859 B.n858 10.6151
R1585 B.n858 B.n857 10.6151
R1586 B.n857 B.n72 10.6151
R1587 B.n851 B.n72 10.6151
R1588 B.n851 B.n850 10.6151
R1589 B.n850 B.n849 10.6151
R1590 B.n849 B.n80 10.6151
R1591 B.n749 B.t9 9.44797
R1592 B.n25 B.t0 9.44797
R1593 B.n219 B.n136 9.36635
R1594 B.n242 B.n133 9.36635
R1595 B.n563 B.n562 9.36635
R1596 B.n541 B.n540 9.36635
R1597 B.t8 B.n375 5.66898
R1598 B.n878 B.t5 5.66898
R1599 B.n355 B.t1 4.40932
R1600 B.t2 B.n902 4.40932
R1601 B.n937 B.n0 2.81026
R1602 B.n937 B.n1 2.81026
R1603 B.n222 B.n136 1.24928
R1604 B.n239 B.n133 1.24928
R1605 B.n562 B.n561 1.24928
R1606 B.n542 B.n541 1.24928
R1607 B.t6 B.n363 0.630331
R1608 B.t3 B.n43 0.630331
R1609 VP.n16 VP.t2 200.19
R1610 VP.n41 VP.n40 177.939
R1611 VP.n70 VP.n69 177.939
R1612 VP.n39 VP.n38 177.939
R1613 VP.n55 VP.t5 167.875
R1614 VP.n41 VP.t8 167.875
R1615 VP.n48 VP.t9 167.875
R1616 VP.n62 VP.t3 167.875
R1617 VP.n69 VP.t7 167.875
R1618 VP.n24 VP.t6 167.875
R1619 VP.n38 VP.t4 167.875
R1620 VP.n31 VP.t1 167.875
R1621 VP.n17 VP.t0 167.875
R1622 VP.n18 VP.n15 161.3
R1623 VP.n20 VP.n19 161.3
R1624 VP.n21 VP.n14 161.3
R1625 VP.n23 VP.n22 161.3
R1626 VP.n24 VP.n13 161.3
R1627 VP.n26 VP.n25 161.3
R1628 VP.n27 VP.n12 161.3
R1629 VP.n29 VP.n28 161.3
R1630 VP.n30 VP.n11 161.3
R1631 VP.n33 VP.n32 161.3
R1632 VP.n34 VP.n10 161.3
R1633 VP.n36 VP.n35 161.3
R1634 VP.n37 VP.n9 161.3
R1635 VP.n68 VP.n0 161.3
R1636 VP.n67 VP.n66 161.3
R1637 VP.n65 VP.n1 161.3
R1638 VP.n64 VP.n63 161.3
R1639 VP.n61 VP.n2 161.3
R1640 VP.n60 VP.n59 161.3
R1641 VP.n58 VP.n3 161.3
R1642 VP.n57 VP.n56 161.3
R1643 VP.n55 VP.n4 161.3
R1644 VP.n54 VP.n53 161.3
R1645 VP.n52 VP.n5 161.3
R1646 VP.n51 VP.n50 161.3
R1647 VP.n49 VP.n6 161.3
R1648 VP.n47 VP.n46 161.3
R1649 VP.n45 VP.n7 161.3
R1650 VP.n44 VP.n43 161.3
R1651 VP.n42 VP.n8 161.3
R1652 VP.n17 VP.n16 63.3281
R1653 VP.n43 VP.n7 52.1486
R1654 VP.n67 VP.n1 52.1486
R1655 VP.n36 VP.n10 52.1486
R1656 VP.n40 VP.n39 48.5914
R1657 VP.n50 VP.n5 44.3785
R1658 VP.n60 VP.n3 44.3785
R1659 VP.n29 VP.n12 44.3785
R1660 VP.n19 VP.n14 44.3785
R1661 VP.n54 VP.n5 36.6083
R1662 VP.n56 VP.n3 36.6083
R1663 VP.n25 VP.n12 36.6083
R1664 VP.n23 VP.n14 36.6083
R1665 VP.n47 VP.n7 28.8382
R1666 VP.n63 VP.n1 28.8382
R1667 VP.n32 VP.n10 28.8382
R1668 VP.n43 VP.n42 24.4675
R1669 VP.n50 VP.n49 24.4675
R1670 VP.n55 VP.n54 24.4675
R1671 VP.n56 VP.n55 24.4675
R1672 VP.n61 VP.n60 24.4675
R1673 VP.n68 VP.n67 24.4675
R1674 VP.n37 VP.n36 24.4675
R1675 VP.n30 VP.n29 24.4675
R1676 VP.n24 VP.n23 24.4675
R1677 VP.n25 VP.n24 24.4675
R1678 VP.n19 VP.n18 24.4675
R1679 VP.n48 VP.n47 20.5528
R1680 VP.n63 VP.n62 20.5528
R1681 VP.n32 VP.n31 20.5528
R1682 VP.n16 VP.n15 18.0704
R1683 VP.n42 VP.n41 7.82994
R1684 VP.n69 VP.n68 7.82994
R1685 VP.n38 VP.n37 7.82994
R1686 VP.n49 VP.n48 3.91522
R1687 VP.n62 VP.n61 3.91522
R1688 VP.n31 VP.n30 3.91522
R1689 VP.n18 VP.n17 3.91522
R1690 VP.n20 VP.n15 0.189894
R1691 VP.n21 VP.n20 0.189894
R1692 VP.n22 VP.n21 0.189894
R1693 VP.n22 VP.n13 0.189894
R1694 VP.n26 VP.n13 0.189894
R1695 VP.n27 VP.n26 0.189894
R1696 VP.n28 VP.n27 0.189894
R1697 VP.n28 VP.n11 0.189894
R1698 VP.n33 VP.n11 0.189894
R1699 VP.n34 VP.n33 0.189894
R1700 VP.n35 VP.n34 0.189894
R1701 VP.n35 VP.n9 0.189894
R1702 VP.n39 VP.n9 0.189894
R1703 VP.n40 VP.n8 0.189894
R1704 VP.n44 VP.n8 0.189894
R1705 VP.n45 VP.n44 0.189894
R1706 VP.n46 VP.n45 0.189894
R1707 VP.n46 VP.n6 0.189894
R1708 VP.n51 VP.n6 0.189894
R1709 VP.n52 VP.n51 0.189894
R1710 VP.n53 VP.n52 0.189894
R1711 VP.n53 VP.n4 0.189894
R1712 VP.n57 VP.n4 0.189894
R1713 VP.n58 VP.n57 0.189894
R1714 VP.n59 VP.n58 0.189894
R1715 VP.n59 VP.n2 0.189894
R1716 VP.n64 VP.n2 0.189894
R1717 VP.n65 VP.n64 0.189894
R1718 VP.n66 VP.n65 0.189894
R1719 VP.n66 VP.n0 0.189894
R1720 VP.n70 VP.n0 0.189894
R1721 VP VP.n70 0.0516364
R1722 VDD1.n60 VDD1.n0 289.615
R1723 VDD1.n127 VDD1.n67 289.615
R1724 VDD1.n61 VDD1.n60 185
R1725 VDD1.n59 VDD1.n58 185
R1726 VDD1.n4 VDD1.n3 185
R1727 VDD1.n53 VDD1.n52 185
R1728 VDD1.n51 VDD1.n50 185
R1729 VDD1.n8 VDD1.n7 185
R1730 VDD1.n45 VDD1.n44 185
R1731 VDD1.n43 VDD1.n10 185
R1732 VDD1.n42 VDD1.n41 185
R1733 VDD1.n13 VDD1.n11 185
R1734 VDD1.n36 VDD1.n35 185
R1735 VDD1.n34 VDD1.n33 185
R1736 VDD1.n17 VDD1.n16 185
R1737 VDD1.n28 VDD1.n27 185
R1738 VDD1.n26 VDD1.n25 185
R1739 VDD1.n21 VDD1.n20 185
R1740 VDD1.n87 VDD1.n86 185
R1741 VDD1.n92 VDD1.n91 185
R1742 VDD1.n94 VDD1.n93 185
R1743 VDD1.n83 VDD1.n82 185
R1744 VDD1.n100 VDD1.n99 185
R1745 VDD1.n102 VDD1.n101 185
R1746 VDD1.n79 VDD1.n78 185
R1747 VDD1.n109 VDD1.n108 185
R1748 VDD1.n110 VDD1.n77 185
R1749 VDD1.n112 VDD1.n111 185
R1750 VDD1.n75 VDD1.n74 185
R1751 VDD1.n118 VDD1.n117 185
R1752 VDD1.n120 VDD1.n119 185
R1753 VDD1.n71 VDD1.n70 185
R1754 VDD1.n126 VDD1.n125 185
R1755 VDD1.n128 VDD1.n127 185
R1756 VDD1.n22 VDD1.t7 149.524
R1757 VDD1.n88 VDD1.t9 149.524
R1758 VDD1.n60 VDD1.n59 104.615
R1759 VDD1.n59 VDD1.n3 104.615
R1760 VDD1.n52 VDD1.n3 104.615
R1761 VDD1.n52 VDD1.n51 104.615
R1762 VDD1.n51 VDD1.n7 104.615
R1763 VDD1.n44 VDD1.n7 104.615
R1764 VDD1.n44 VDD1.n43 104.615
R1765 VDD1.n43 VDD1.n42 104.615
R1766 VDD1.n42 VDD1.n11 104.615
R1767 VDD1.n35 VDD1.n11 104.615
R1768 VDD1.n35 VDD1.n34 104.615
R1769 VDD1.n34 VDD1.n16 104.615
R1770 VDD1.n27 VDD1.n16 104.615
R1771 VDD1.n27 VDD1.n26 104.615
R1772 VDD1.n26 VDD1.n20 104.615
R1773 VDD1.n92 VDD1.n86 104.615
R1774 VDD1.n93 VDD1.n92 104.615
R1775 VDD1.n93 VDD1.n82 104.615
R1776 VDD1.n100 VDD1.n82 104.615
R1777 VDD1.n101 VDD1.n100 104.615
R1778 VDD1.n101 VDD1.n78 104.615
R1779 VDD1.n109 VDD1.n78 104.615
R1780 VDD1.n110 VDD1.n109 104.615
R1781 VDD1.n111 VDD1.n110 104.615
R1782 VDD1.n111 VDD1.n74 104.615
R1783 VDD1.n118 VDD1.n74 104.615
R1784 VDD1.n119 VDD1.n118 104.615
R1785 VDD1.n119 VDD1.n70 104.615
R1786 VDD1.n126 VDD1.n70 104.615
R1787 VDD1.n127 VDD1.n126 104.615
R1788 VDD1.n135 VDD1.n134 64.5268
R1789 VDD1.n66 VDD1.n65 63.2375
R1790 VDD1.n137 VDD1.n136 63.2374
R1791 VDD1.n133 VDD1.n132 63.2374
R1792 VDD1.t7 VDD1.n20 52.3082
R1793 VDD1.t9 VDD1.n86 52.3082
R1794 VDD1.n66 VDD1.n64 52.0148
R1795 VDD1.n133 VDD1.n131 52.0148
R1796 VDD1.n137 VDD1.n135 44.2207
R1797 VDD1.n45 VDD1.n10 13.1884
R1798 VDD1.n112 VDD1.n77 13.1884
R1799 VDD1.n46 VDD1.n8 12.8005
R1800 VDD1.n41 VDD1.n12 12.8005
R1801 VDD1.n108 VDD1.n107 12.8005
R1802 VDD1.n113 VDD1.n75 12.8005
R1803 VDD1.n50 VDD1.n49 12.0247
R1804 VDD1.n40 VDD1.n13 12.0247
R1805 VDD1.n106 VDD1.n79 12.0247
R1806 VDD1.n117 VDD1.n116 12.0247
R1807 VDD1.n53 VDD1.n6 11.249
R1808 VDD1.n37 VDD1.n36 11.249
R1809 VDD1.n103 VDD1.n102 11.249
R1810 VDD1.n120 VDD1.n73 11.249
R1811 VDD1.n54 VDD1.n4 10.4732
R1812 VDD1.n33 VDD1.n15 10.4732
R1813 VDD1.n99 VDD1.n81 10.4732
R1814 VDD1.n121 VDD1.n71 10.4732
R1815 VDD1.n22 VDD1.n21 10.2747
R1816 VDD1.n88 VDD1.n87 10.2747
R1817 VDD1.n58 VDD1.n57 9.69747
R1818 VDD1.n32 VDD1.n17 9.69747
R1819 VDD1.n98 VDD1.n83 9.69747
R1820 VDD1.n125 VDD1.n124 9.69747
R1821 VDD1.n64 VDD1.n63 9.45567
R1822 VDD1.n131 VDD1.n130 9.45567
R1823 VDD1.n24 VDD1.n23 9.3005
R1824 VDD1.n19 VDD1.n18 9.3005
R1825 VDD1.n30 VDD1.n29 9.3005
R1826 VDD1.n32 VDD1.n31 9.3005
R1827 VDD1.n15 VDD1.n14 9.3005
R1828 VDD1.n38 VDD1.n37 9.3005
R1829 VDD1.n40 VDD1.n39 9.3005
R1830 VDD1.n12 VDD1.n9 9.3005
R1831 VDD1.n63 VDD1.n62 9.3005
R1832 VDD1.n2 VDD1.n1 9.3005
R1833 VDD1.n57 VDD1.n56 9.3005
R1834 VDD1.n55 VDD1.n54 9.3005
R1835 VDD1.n6 VDD1.n5 9.3005
R1836 VDD1.n49 VDD1.n48 9.3005
R1837 VDD1.n47 VDD1.n46 9.3005
R1838 VDD1.n130 VDD1.n129 9.3005
R1839 VDD1.n69 VDD1.n68 9.3005
R1840 VDD1.n124 VDD1.n123 9.3005
R1841 VDD1.n122 VDD1.n121 9.3005
R1842 VDD1.n73 VDD1.n72 9.3005
R1843 VDD1.n116 VDD1.n115 9.3005
R1844 VDD1.n114 VDD1.n113 9.3005
R1845 VDD1.n90 VDD1.n89 9.3005
R1846 VDD1.n85 VDD1.n84 9.3005
R1847 VDD1.n96 VDD1.n95 9.3005
R1848 VDD1.n98 VDD1.n97 9.3005
R1849 VDD1.n81 VDD1.n80 9.3005
R1850 VDD1.n104 VDD1.n103 9.3005
R1851 VDD1.n106 VDD1.n105 9.3005
R1852 VDD1.n107 VDD1.n76 9.3005
R1853 VDD1.n61 VDD1.n2 8.92171
R1854 VDD1.n29 VDD1.n28 8.92171
R1855 VDD1.n95 VDD1.n94 8.92171
R1856 VDD1.n128 VDD1.n69 8.92171
R1857 VDD1.n62 VDD1.n0 8.14595
R1858 VDD1.n25 VDD1.n19 8.14595
R1859 VDD1.n91 VDD1.n85 8.14595
R1860 VDD1.n129 VDD1.n67 8.14595
R1861 VDD1.n24 VDD1.n21 7.3702
R1862 VDD1.n90 VDD1.n87 7.3702
R1863 VDD1.n64 VDD1.n0 5.81868
R1864 VDD1.n25 VDD1.n24 5.81868
R1865 VDD1.n91 VDD1.n90 5.81868
R1866 VDD1.n131 VDD1.n67 5.81868
R1867 VDD1.n62 VDD1.n61 5.04292
R1868 VDD1.n28 VDD1.n19 5.04292
R1869 VDD1.n94 VDD1.n85 5.04292
R1870 VDD1.n129 VDD1.n128 5.04292
R1871 VDD1.n58 VDD1.n2 4.26717
R1872 VDD1.n29 VDD1.n17 4.26717
R1873 VDD1.n95 VDD1.n83 4.26717
R1874 VDD1.n125 VDD1.n69 4.26717
R1875 VDD1.n57 VDD1.n4 3.49141
R1876 VDD1.n33 VDD1.n32 3.49141
R1877 VDD1.n99 VDD1.n98 3.49141
R1878 VDD1.n124 VDD1.n71 3.49141
R1879 VDD1.n23 VDD1.n22 2.84303
R1880 VDD1.n89 VDD1.n88 2.84303
R1881 VDD1.n54 VDD1.n53 2.71565
R1882 VDD1.n36 VDD1.n15 2.71565
R1883 VDD1.n102 VDD1.n81 2.71565
R1884 VDD1.n121 VDD1.n120 2.71565
R1885 VDD1.n50 VDD1.n6 1.93989
R1886 VDD1.n37 VDD1.n13 1.93989
R1887 VDD1.n103 VDD1.n79 1.93989
R1888 VDD1.n117 VDD1.n73 1.93989
R1889 VDD1.n136 VDD1.t3 1.62478
R1890 VDD1.n136 VDD1.t1 1.62478
R1891 VDD1.n65 VDD1.t2 1.62478
R1892 VDD1.n65 VDD1.t5 1.62478
R1893 VDD1.n134 VDD1.t0 1.62478
R1894 VDD1.n134 VDD1.t6 1.62478
R1895 VDD1.n132 VDD1.t4 1.62478
R1896 VDD1.n132 VDD1.t8 1.62478
R1897 VDD1 VDD1.n137 1.28714
R1898 VDD1.n49 VDD1.n8 1.16414
R1899 VDD1.n41 VDD1.n40 1.16414
R1900 VDD1.n108 VDD1.n106 1.16414
R1901 VDD1.n116 VDD1.n75 1.16414
R1902 VDD1 VDD1.n66 0.506965
R1903 VDD1.n135 VDD1.n133 0.39343
R1904 VDD1.n46 VDD1.n45 0.388379
R1905 VDD1.n12 VDD1.n10 0.388379
R1906 VDD1.n107 VDD1.n77 0.388379
R1907 VDD1.n113 VDD1.n112 0.388379
R1908 VDD1.n63 VDD1.n1 0.155672
R1909 VDD1.n56 VDD1.n1 0.155672
R1910 VDD1.n56 VDD1.n55 0.155672
R1911 VDD1.n55 VDD1.n5 0.155672
R1912 VDD1.n48 VDD1.n5 0.155672
R1913 VDD1.n48 VDD1.n47 0.155672
R1914 VDD1.n47 VDD1.n9 0.155672
R1915 VDD1.n39 VDD1.n9 0.155672
R1916 VDD1.n39 VDD1.n38 0.155672
R1917 VDD1.n38 VDD1.n14 0.155672
R1918 VDD1.n31 VDD1.n14 0.155672
R1919 VDD1.n31 VDD1.n30 0.155672
R1920 VDD1.n30 VDD1.n18 0.155672
R1921 VDD1.n23 VDD1.n18 0.155672
R1922 VDD1.n89 VDD1.n84 0.155672
R1923 VDD1.n96 VDD1.n84 0.155672
R1924 VDD1.n97 VDD1.n96 0.155672
R1925 VDD1.n97 VDD1.n80 0.155672
R1926 VDD1.n104 VDD1.n80 0.155672
R1927 VDD1.n105 VDD1.n104 0.155672
R1928 VDD1.n105 VDD1.n76 0.155672
R1929 VDD1.n114 VDD1.n76 0.155672
R1930 VDD1.n115 VDD1.n114 0.155672
R1931 VDD1.n115 VDD1.n72 0.155672
R1932 VDD1.n122 VDD1.n72 0.155672
R1933 VDD1.n123 VDD1.n122 0.155672
R1934 VDD1.n123 VDD1.n68 0.155672
R1935 VDD1.n130 VDD1.n68 0.155672
R1936 VTAIL.n272 VTAIL.n212 289.615
R1937 VTAIL.n62 VTAIL.n2 289.615
R1938 VTAIL.n206 VTAIL.n146 289.615
R1939 VTAIL.n136 VTAIL.n76 289.615
R1940 VTAIL.n232 VTAIL.n231 185
R1941 VTAIL.n237 VTAIL.n236 185
R1942 VTAIL.n239 VTAIL.n238 185
R1943 VTAIL.n228 VTAIL.n227 185
R1944 VTAIL.n245 VTAIL.n244 185
R1945 VTAIL.n247 VTAIL.n246 185
R1946 VTAIL.n224 VTAIL.n223 185
R1947 VTAIL.n254 VTAIL.n253 185
R1948 VTAIL.n255 VTAIL.n222 185
R1949 VTAIL.n257 VTAIL.n256 185
R1950 VTAIL.n220 VTAIL.n219 185
R1951 VTAIL.n263 VTAIL.n262 185
R1952 VTAIL.n265 VTAIL.n264 185
R1953 VTAIL.n216 VTAIL.n215 185
R1954 VTAIL.n271 VTAIL.n270 185
R1955 VTAIL.n273 VTAIL.n272 185
R1956 VTAIL.n22 VTAIL.n21 185
R1957 VTAIL.n27 VTAIL.n26 185
R1958 VTAIL.n29 VTAIL.n28 185
R1959 VTAIL.n18 VTAIL.n17 185
R1960 VTAIL.n35 VTAIL.n34 185
R1961 VTAIL.n37 VTAIL.n36 185
R1962 VTAIL.n14 VTAIL.n13 185
R1963 VTAIL.n44 VTAIL.n43 185
R1964 VTAIL.n45 VTAIL.n12 185
R1965 VTAIL.n47 VTAIL.n46 185
R1966 VTAIL.n10 VTAIL.n9 185
R1967 VTAIL.n53 VTAIL.n52 185
R1968 VTAIL.n55 VTAIL.n54 185
R1969 VTAIL.n6 VTAIL.n5 185
R1970 VTAIL.n61 VTAIL.n60 185
R1971 VTAIL.n63 VTAIL.n62 185
R1972 VTAIL.n207 VTAIL.n206 185
R1973 VTAIL.n205 VTAIL.n204 185
R1974 VTAIL.n150 VTAIL.n149 185
R1975 VTAIL.n199 VTAIL.n198 185
R1976 VTAIL.n197 VTAIL.n196 185
R1977 VTAIL.n154 VTAIL.n153 185
R1978 VTAIL.n191 VTAIL.n190 185
R1979 VTAIL.n189 VTAIL.n156 185
R1980 VTAIL.n188 VTAIL.n187 185
R1981 VTAIL.n159 VTAIL.n157 185
R1982 VTAIL.n182 VTAIL.n181 185
R1983 VTAIL.n180 VTAIL.n179 185
R1984 VTAIL.n163 VTAIL.n162 185
R1985 VTAIL.n174 VTAIL.n173 185
R1986 VTAIL.n172 VTAIL.n171 185
R1987 VTAIL.n167 VTAIL.n166 185
R1988 VTAIL.n137 VTAIL.n136 185
R1989 VTAIL.n135 VTAIL.n134 185
R1990 VTAIL.n80 VTAIL.n79 185
R1991 VTAIL.n129 VTAIL.n128 185
R1992 VTAIL.n127 VTAIL.n126 185
R1993 VTAIL.n84 VTAIL.n83 185
R1994 VTAIL.n121 VTAIL.n120 185
R1995 VTAIL.n119 VTAIL.n86 185
R1996 VTAIL.n118 VTAIL.n117 185
R1997 VTAIL.n89 VTAIL.n87 185
R1998 VTAIL.n112 VTAIL.n111 185
R1999 VTAIL.n110 VTAIL.n109 185
R2000 VTAIL.n93 VTAIL.n92 185
R2001 VTAIL.n104 VTAIL.n103 185
R2002 VTAIL.n102 VTAIL.n101 185
R2003 VTAIL.n97 VTAIL.n96 185
R2004 VTAIL.n233 VTAIL.t8 149.524
R2005 VTAIL.n23 VTAIL.t12 149.524
R2006 VTAIL.n168 VTAIL.t15 149.524
R2007 VTAIL.n98 VTAIL.t3 149.524
R2008 VTAIL.n237 VTAIL.n231 104.615
R2009 VTAIL.n238 VTAIL.n237 104.615
R2010 VTAIL.n238 VTAIL.n227 104.615
R2011 VTAIL.n245 VTAIL.n227 104.615
R2012 VTAIL.n246 VTAIL.n245 104.615
R2013 VTAIL.n246 VTAIL.n223 104.615
R2014 VTAIL.n254 VTAIL.n223 104.615
R2015 VTAIL.n255 VTAIL.n254 104.615
R2016 VTAIL.n256 VTAIL.n255 104.615
R2017 VTAIL.n256 VTAIL.n219 104.615
R2018 VTAIL.n263 VTAIL.n219 104.615
R2019 VTAIL.n264 VTAIL.n263 104.615
R2020 VTAIL.n264 VTAIL.n215 104.615
R2021 VTAIL.n271 VTAIL.n215 104.615
R2022 VTAIL.n272 VTAIL.n271 104.615
R2023 VTAIL.n27 VTAIL.n21 104.615
R2024 VTAIL.n28 VTAIL.n27 104.615
R2025 VTAIL.n28 VTAIL.n17 104.615
R2026 VTAIL.n35 VTAIL.n17 104.615
R2027 VTAIL.n36 VTAIL.n35 104.615
R2028 VTAIL.n36 VTAIL.n13 104.615
R2029 VTAIL.n44 VTAIL.n13 104.615
R2030 VTAIL.n45 VTAIL.n44 104.615
R2031 VTAIL.n46 VTAIL.n45 104.615
R2032 VTAIL.n46 VTAIL.n9 104.615
R2033 VTAIL.n53 VTAIL.n9 104.615
R2034 VTAIL.n54 VTAIL.n53 104.615
R2035 VTAIL.n54 VTAIL.n5 104.615
R2036 VTAIL.n61 VTAIL.n5 104.615
R2037 VTAIL.n62 VTAIL.n61 104.615
R2038 VTAIL.n206 VTAIL.n205 104.615
R2039 VTAIL.n205 VTAIL.n149 104.615
R2040 VTAIL.n198 VTAIL.n149 104.615
R2041 VTAIL.n198 VTAIL.n197 104.615
R2042 VTAIL.n197 VTAIL.n153 104.615
R2043 VTAIL.n190 VTAIL.n153 104.615
R2044 VTAIL.n190 VTAIL.n189 104.615
R2045 VTAIL.n189 VTAIL.n188 104.615
R2046 VTAIL.n188 VTAIL.n157 104.615
R2047 VTAIL.n181 VTAIL.n157 104.615
R2048 VTAIL.n181 VTAIL.n180 104.615
R2049 VTAIL.n180 VTAIL.n162 104.615
R2050 VTAIL.n173 VTAIL.n162 104.615
R2051 VTAIL.n173 VTAIL.n172 104.615
R2052 VTAIL.n172 VTAIL.n166 104.615
R2053 VTAIL.n136 VTAIL.n135 104.615
R2054 VTAIL.n135 VTAIL.n79 104.615
R2055 VTAIL.n128 VTAIL.n79 104.615
R2056 VTAIL.n128 VTAIL.n127 104.615
R2057 VTAIL.n127 VTAIL.n83 104.615
R2058 VTAIL.n120 VTAIL.n83 104.615
R2059 VTAIL.n120 VTAIL.n119 104.615
R2060 VTAIL.n119 VTAIL.n118 104.615
R2061 VTAIL.n118 VTAIL.n87 104.615
R2062 VTAIL.n111 VTAIL.n87 104.615
R2063 VTAIL.n111 VTAIL.n110 104.615
R2064 VTAIL.n110 VTAIL.n92 104.615
R2065 VTAIL.n103 VTAIL.n92 104.615
R2066 VTAIL.n103 VTAIL.n102 104.615
R2067 VTAIL.n102 VTAIL.n96 104.615
R2068 VTAIL.t8 VTAIL.n231 52.3082
R2069 VTAIL.t12 VTAIL.n21 52.3082
R2070 VTAIL.t15 VTAIL.n166 52.3082
R2071 VTAIL.t3 VTAIL.n96 52.3082
R2072 VTAIL.n145 VTAIL.n144 46.5587
R2073 VTAIL.n143 VTAIL.n142 46.5587
R2074 VTAIL.n75 VTAIL.n74 46.5587
R2075 VTAIL.n73 VTAIL.n72 46.5587
R2076 VTAIL.n279 VTAIL.n278 46.5586
R2077 VTAIL.n1 VTAIL.n0 46.5586
R2078 VTAIL.n69 VTAIL.n68 46.5586
R2079 VTAIL.n71 VTAIL.n70 46.5586
R2080 VTAIL.n277 VTAIL.n276 33.5429
R2081 VTAIL.n67 VTAIL.n66 33.5429
R2082 VTAIL.n211 VTAIL.n210 33.5429
R2083 VTAIL.n141 VTAIL.n140 33.5429
R2084 VTAIL.n73 VTAIL.n71 26.4617
R2085 VTAIL.n277 VTAIL.n211 24.6686
R2086 VTAIL.n257 VTAIL.n222 13.1884
R2087 VTAIL.n47 VTAIL.n12 13.1884
R2088 VTAIL.n191 VTAIL.n156 13.1884
R2089 VTAIL.n121 VTAIL.n86 13.1884
R2090 VTAIL.n253 VTAIL.n252 12.8005
R2091 VTAIL.n258 VTAIL.n220 12.8005
R2092 VTAIL.n43 VTAIL.n42 12.8005
R2093 VTAIL.n48 VTAIL.n10 12.8005
R2094 VTAIL.n192 VTAIL.n154 12.8005
R2095 VTAIL.n187 VTAIL.n158 12.8005
R2096 VTAIL.n122 VTAIL.n84 12.8005
R2097 VTAIL.n117 VTAIL.n88 12.8005
R2098 VTAIL.n251 VTAIL.n224 12.0247
R2099 VTAIL.n262 VTAIL.n261 12.0247
R2100 VTAIL.n41 VTAIL.n14 12.0247
R2101 VTAIL.n52 VTAIL.n51 12.0247
R2102 VTAIL.n196 VTAIL.n195 12.0247
R2103 VTAIL.n186 VTAIL.n159 12.0247
R2104 VTAIL.n126 VTAIL.n125 12.0247
R2105 VTAIL.n116 VTAIL.n89 12.0247
R2106 VTAIL.n248 VTAIL.n247 11.249
R2107 VTAIL.n265 VTAIL.n218 11.249
R2108 VTAIL.n38 VTAIL.n37 11.249
R2109 VTAIL.n55 VTAIL.n8 11.249
R2110 VTAIL.n199 VTAIL.n152 11.249
R2111 VTAIL.n183 VTAIL.n182 11.249
R2112 VTAIL.n129 VTAIL.n82 11.249
R2113 VTAIL.n113 VTAIL.n112 11.249
R2114 VTAIL.n244 VTAIL.n226 10.4732
R2115 VTAIL.n266 VTAIL.n216 10.4732
R2116 VTAIL.n34 VTAIL.n16 10.4732
R2117 VTAIL.n56 VTAIL.n6 10.4732
R2118 VTAIL.n200 VTAIL.n150 10.4732
R2119 VTAIL.n179 VTAIL.n161 10.4732
R2120 VTAIL.n130 VTAIL.n80 10.4732
R2121 VTAIL.n109 VTAIL.n91 10.4732
R2122 VTAIL.n233 VTAIL.n232 10.2747
R2123 VTAIL.n23 VTAIL.n22 10.2747
R2124 VTAIL.n168 VTAIL.n167 10.2747
R2125 VTAIL.n98 VTAIL.n97 10.2747
R2126 VTAIL.n243 VTAIL.n228 9.69747
R2127 VTAIL.n270 VTAIL.n269 9.69747
R2128 VTAIL.n33 VTAIL.n18 9.69747
R2129 VTAIL.n60 VTAIL.n59 9.69747
R2130 VTAIL.n204 VTAIL.n203 9.69747
R2131 VTAIL.n178 VTAIL.n163 9.69747
R2132 VTAIL.n134 VTAIL.n133 9.69747
R2133 VTAIL.n108 VTAIL.n93 9.69747
R2134 VTAIL.n276 VTAIL.n275 9.45567
R2135 VTAIL.n66 VTAIL.n65 9.45567
R2136 VTAIL.n210 VTAIL.n209 9.45567
R2137 VTAIL.n140 VTAIL.n139 9.45567
R2138 VTAIL.n275 VTAIL.n274 9.3005
R2139 VTAIL.n214 VTAIL.n213 9.3005
R2140 VTAIL.n269 VTAIL.n268 9.3005
R2141 VTAIL.n267 VTAIL.n266 9.3005
R2142 VTAIL.n218 VTAIL.n217 9.3005
R2143 VTAIL.n261 VTAIL.n260 9.3005
R2144 VTAIL.n259 VTAIL.n258 9.3005
R2145 VTAIL.n235 VTAIL.n234 9.3005
R2146 VTAIL.n230 VTAIL.n229 9.3005
R2147 VTAIL.n241 VTAIL.n240 9.3005
R2148 VTAIL.n243 VTAIL.n242 9.3005
R2149 VTAIL.n226 VTAIL.n225 9.3005
R2150 VTAIL.n249 VTAIL.n248 9.3005
R2151 VTAIL.n251 VTAIL.n250 9.3005
R2152 VTAIL.n252 VTAIL.n221 9.3005
R2153 VTAIL.n65 VTAIL.n64 9.3005
R2154 VTAIL.n4 VTAIL.n3 9.3005
R2155 VTAIL.n59 VTAIL.n58 9.3005
R2156 VTAIL.n57 VTAIL.n56 9.3005
R2157 VTAIL.n8 VTAIL.n7 9.3005
R2158 VTAIL.n51 VTAIL.n50 9.3005
R2159 VTAIL.n49 VTAIL.n48 9.3005
R2160 VTAIL.n25 VTAIL.n24 9.3005
R2161 VTAIL.n20 VTAIL.n19 9.3005
R2162 VTAIL.n31 VTAIL.n30 9.3005
R2163 VTAIL.n33 VTAIL.n32 9.3005
R2164 VTAIL.n16 VTAIL.n15 9.3005
R2165 VTAIL.n39 VTAIL.n38 9.3005
R2166 VTAIL.n41 VTAIL.n40 9.3005
R2167 VTAIL.n42 VTAIL.n11 9.3005
R2168 VTAIL.n170 VTAIL.n169 9.3005
R2169 VTAIL.n165 VTAIL.n164 9.3005
R2170 VTAIL.n176 VTAIL.n175 9.3005
R2171 VTAIL.n178 VTAIL.n177 9.3005
R2172 VTAIL.n161 VTAIL.n160 9.3005
R2173 VTAIL.n184 VTAIL.n183 9.3005
R2174 VTAIL.n186 VTAIL.n185 9.3005
R2175 VTAIL.n158 VTAIL.n155 9.3005
R2176 VTAIL.n209 VTAIL.n208 9.3005
R2177 VTAIL.n148 VTAIL.n147 9.3005
R2178 VTAIL.n203 VTAIL.n202 9.3005
R2179 VTAIL.n201 VTAIL.n200 9.3005
R2180 VTAIL.n152 VTAIL.n151 9.3005
R2181 VTAIL.n195 VTAIL.n194 9.3005
R2182 VTAIL.n193 VTAIL.n192 9.3005
R2183 VTAIL.n100 VTAIL.n99 9.3005
R2184 VTAIL.n95 VTAIL.n94 9.3005
R2185 VTAIL.n106 VTAIL.n105 9.3005
R2186 VTAIL.n108 VTAIL.n107 9.3005
R2187 VTAIL.n91 VTAIL.n90 9.3005
R2188 VTAIL.n114 VTAIL.n113 9.3005
R2189 VTAIL.n116 VTAIL.n115 9.3005
R2190 VTAIL.n88 VTAIL.n85 9.3005
R2191 VTAIL.n139 VTAIL.n138 9.3005
R2192 VTAIL.n78 VTAIL.n77 9.3005
R2193 VTAIL.n133 VTAIL.n132 9.3005
R2194 VTAIL.n131 VTAIL.n130 9.3005
R2195 VTAIL.n82 VTAIL.n81 9.3005
R2196 VTAIL.n125 VTAIL.n124 9.3005
R2197 VTAIL.n123 VTAIL.n122 9.3005
R2198 VTAIL.n240 VTAIL.n239 8.92171
R2199 VTAIL.n273 VTAIL.n214 8.92171
R2200 VTAIL.n30 VTAIL.n29 8.92171
R2201 VTAIL.n63 VTAIL.n4 8.92171
R2202 VTAIL.n207 VTAIL.n148 8.92171
R2203 VTAIL.n175 VTAIL.n174 8.92171
R2204 VTAIL.n137 VTAIL.n78 8.92171
R2205 VTAIL.n105 VTAIL.n104 8.92171
R2206 VTAIL.n236 VTAIL.n230 8.14595
R2207 VTAIL.n274 VTAIL.n212 8.14595
R2208 VTAIL.n26 VTAIL.n20 8.14595
R2209 VTAIL.n64 VTAIL.n2 8.14595
R2210 VTAIL.n208 VTAIL.n146 8.14595
R2211 VTAIL.n171 VTAIL.n165 8.14595
R2212 VTAIL.n138 VTAIL.n76 8.14595
R2213 VTAIL.n101 VTAIL.n95 8.14595
R2214 VTAIL.n235 VTAIL.n232 7.3702
R2215 VTAIL.n25 VTAIL.n22 7.3702
R2216 VTAIL.n170 VTAIL.n167 7.3702
R2217 VTAIL.n100 VTAIL.n97 7.3702
R2218 VTAIL.n236 VTAIL.n235 5.81868
R2219 VTAIL.n276 VTAIL.n212 5.81868
R2220 VTAIL.n26 VTAIL.n25 5.81868
R2221 VTAIL.n66 VTAIL.n2 5.81868
R2222 VTAIL.n210 VTAIL.n146 5.81868
R2223 VTAIL.n171 VTAIL.n170 5.81868
R2224 VTAIL.n140 VTAIL.n76 5.81868
R2225 VTAIL.n101 VTAIL.n100 5.81868
R2226 VTAIL.n239 VTAIL.n230 5.04292
R2227 VTAIL.n274 VTAIL.n273 5.04292
R2228 VTAIL.n29 VTAIL.n20 5.04292
R2229 VTAIL.n64 VTAIL.n63 5.04292
R2230 VTAIL.n208 VTAIL.n207 5.04292
R2231 VTAIL.n174 VTAIL.n165 5.04292
R2232 VTAIL.n138 VTAIL.n137 5.04292
R2233 VTAIL.n104 VTAIL.n95 5.04292
R2234 VTAIL.n240 VTAIL.n228 4.26717
R2235 VTAIL.n270 VTAIL.n214 4.26717
R2236 VTAIL.n30 VTAIL.n18 4.26717
R2237 VTAIL.n60 VTAIL.n4 4.26717
R2238 VTAIL.n204 VTAIL.n148 4.26717
R2239 VTAIL.n175 VTAIL.n163 4.26717
R2240 VTAIL.n134 VTAIL.n78 4.26717
R2241 VTAIL.n105 VTAIL.n93 4.26717
R2242 VTAIL.n244 VTAIL.n243 3.49141
R2243 VTAIL.n269 VTAIL.n216 3.49141
R2244 VTAIL.n34 VTAIL.n33 3.49141
R2245 VTAIL.n59 VTAIL.n6 3.49141
R2246 VTAIL.n203 VTAIL.n150 3.49141
R2247 VTAIL.n179 VTAIL.n178 3.49141
R2248 VTAIL.n133 VTAIL.n80 3.49141
R2249 VTAIL.n109 VTAIL.n108 3.49141
R2250 VTAIL.n234 VTAIL.n233 2.84303
R2251 VTAIL.n24 VTAIL.n23 2.84303
R2252 VTAIL.n169 VTAIL.n168 2.84303
R2253 VTAIL.n99 VTAIL.n98 2.84303
R2254 VTAIL.n247 VTAIL.n226 2.71565
R2255 VTAIL.n266 VTAIL.n265 2.71565
R2256 VTAIL.n37 VTAIL.n16 2.71565
R2257 VTAIL.n56 VTAIL.n55 2.71565
R2258 VTAIL.n200 VTAIL.n199 2.71565
R2259 VTAIL.n182 VTAIL.n161 2.71565
R2260 VTAIL.n130 VTAIL.n129 2.71565
R2261 VTAIL.n112 VTAIL.n91 2.71565
R2262 VTAIL.n248 VTAIL.n224 1.93989
R2263 VTAIL.n262 VTAIL.n218 1.93989
R2264 VTAIL.n38 VTAIL.n14 1.93989
R2265 VTAIL.n52 VTAIL.n8 1.93989
R2266 VTAIL.n196 VTAIL.n152 1.93989
R2267 VTAIL.n183 VTAIL.n159 1.93989
R2268 VTAIL.n126 VTAIL.n82 1.93989
R2269 VTAIL.n113 VTAIL.n89 1.93989
R2270 VTAIL.n75 VTAIL.n73 1.7936
R2271 VTAIL.n141 VTAIL.n75 1.7936
R2272 VTAIL.n145 VTAIL.n143 1.7936
R2273 VTAIL.n211 VTAIL.n145 1.7936
R2274 VTAIL.n71 VTAIL.n69 1.7936
R2275 VTAIL.n69 VTAIL.n67 1.7936
R2276 VTAIL.n279 VTAIL.n277 1.7936
R2277 VTAIL.n278 VTAIL.t1 1.62478
R2278 VTAIL.n278 VTAIL.t2 1.62478
R2279 VTAIL.n0 VTAIL.t6 1.62478
R2280 VTAIL.n0 VTAIL.t0 1.62478
R2281 VTAIL.n68 VTAIL.t14 1.62478
R2282 VTAIL.n68 VTAIL.t16 1.62478
R2283 VTAIL.n70 VTAIL.t11 1.62478
R2284 VTAIL.n70 VTAIL.t10 1.62478
R2285 VTAIL.n144 VTAIL.t13 1.62478
R2286 VTAIL.n144 VTAIL.t18 1.62478
R2287 VTAIL.n142 VTAIL.t17 1.62478
R2288 VTAIL.n142 VTAIL.t19 1.62478
R2289 VTAIL.n74 VTAIL.t5 1.62478
R2290 VTAIL.n74 VTAIL.t9 1.62478
R2291 VTAIL.n72 VTAIL.t7 1.62478
R2292 VTAIL.n72 VTAIL.t4 1.62478
R2293 VTAIL VTAIL.n1 1.40352
R2294 VTAIL.n143 VTAIL.n141 1.36688
R2295 VTAIL.n67 VTAIL.n1 1.36688
R2296 VTAIL.n253 VTAIL.n251 1.16414
R2297 VTAIL.n261 VTAIL.n220 1.16414
R2298 VTAIL.n43 VTAIL.n41 1.16414
R2299 VTAIL.n51 VTAIL.n10 1.16414
R2300 VTAIL.n195 VTAIL.n154 1.16414
R2301 VTAIL.n187 VTAIL.n186 1.16414
R2302 VTAIL.n125 VTAIL.n84 1.16414
R2303 VTAIL.n117 VTAIL.n116 1.16414
R2304 VTAIL VTAIL.n279 0.390586
R2305 VTAIL.n252 VTAIL.n222 0.388379
R2306 VTAIL.n258 VTAIL.n257 0.388379
R2307 VTAIL.n42 VTAIL.n12 0.388379
R2308 VTAIL.n48 VTAIL.n47 0.388379
R2309 VTAIL.n192 VTAIL.n191 0.388379
R2310 VTAIL.n158 VTAIL.n156 0.388379
R2311 VTAIL.n122 VTAIL.n121 0.388379
R2312 VTAIL.n88 VTAIL.n86 0.388379
R2313 VTAIL.n234 VTAIL.n229 0.155672
R2314 VTAIL.n241 VTAIL.n229 0.155672
R2315 VTAIL.n242 VTAIL.n241 0.155672
R2316 VTAIL.n242 VTAIL.n225 0.155672
R2317 VTAIL.n249 VTAIL.n225 0.155672
R2318 VTAIL.n250 VTAIL.n249 0.155672
R2319 VTAIL.n250 VTAIL.n221 0.155672
R2320 VTAIL.n259 VTAIL.n221 0.155672
R2321 VTAIL.n260 VTAIL.n259 0.155672
R2322 VTAIL.n260 VTAIL.n217 0.155672
R2323 VTAIL.n267 VTAIL.n217 0.155672
R2324 VTAIL.n268 VTAIL.n267 0.155672
R2325 VTAIL.n268 VTAIL.n213 0.155672
R2326 VTAIL.n275 VTAIL.n213 0.155672
R2327 VTAIL.n24 VTAIL.n19 0.155672
R2328 VTAIL.n31 VTAIL.n19 0.155672
R2329 VTAIL.n32 VTAIL.n31 0.155672
R2330 VTAIL.n32 VTAIL.n15 0.155672
R2331 VTAIL.n39 VTAIL.n15 0.155672
R2332 VTAIL.n40 VTAIL.n39 0.155672
R2333 VTAIL.n40 VTAIL.n11 0.155672
R2334 VTAIL.n49 VTAIL.n11 0.155672
R2335 VTAIL.n50 VTAIL.n49 0.155672
R2336 VTAIL.n50 VTAIL.n7 0.155672
R2337 VTAIL.n57 VTAIL.n7 0.155672
R2338 VTAIL.n58 VTAIL.n57 0.155672
R2339 VTAIL.n58 VTAIL.n3 0.155672
R2340 VTAIL.n65 VTAIL.n3 0.155672
R2341 VTAIL.n209 VTAIL.n147 0.155672
R2342 VTAIL.n202 VTAIL.n147 0.155672
R2343 VTAIL.n202 VTAIL.n201 0.155672
R2344 VTAIL.n201 VTAIL.n151 0.155672
R2345 VTAIL.n194 VTAIL.n151 0.155672
R2346 VTAIL.n194 VTAIL.n193 0.155672
R2347 VTAIL.n193 VTAIL.n155 0.155672
R2348 VTAIL.n185 VTAIL.n155 0.155672
R2349 VTAIL.n185 VTAIL.n184 0.155672
R2350 VTAIL.n184 VTAIL.n160 0.155672
R2351 VTAIL.n177 VTAIL.n160 0.155672
R2352 VTAIL.n177 VTAIL.n176 0.155672
R2353 VTAIL.n176 VTAIL.n164 0.155672
R2354 VTAIL.n169 VTAIL.n164 0.155672
R2355 VTAIL.n139 VTAIL.n77 0.155672
R2356 VTAIL.n132 VTAIL.n77 0.155672
R2357 VTAIL.n132 VTAIL.n131 0.155672
R2358 VTAIL.n131 VTAIL.n81 0.155672
R2359 VTAIL.n124 VTAIL.n81 0.155672
R2360 VTAIL.n124 VTAIL.n123 0.155672
R2361 VTAIL.n123 VTAIL.n85 0.155672
R2362 VTAIL.n115 VTAIL.n85 0.155672
R2363 VTAIL.n115 VTAIL.n114 0.155672
R2364 VTAIL.n114 VTAIL.n90 0.155672
R2365 VTAIL.n107 VTAIL.n90 0.155672
R2366 VTAIL.n107 VTAIL.n106 0.155672
R2367 VTAIL.n106 VTAIL.n94 0.155672
R2368 VTAIL.n99 VTAIL.n94 0.155672
R2369 VN.n7 VN.t5 200.19
R2370 VN.n38 VN.t7 200.19
R2371 VN.n30 VN.n29 177.939
R2372 VN.n61 VN.n60 177.939
R2373 VN.n15 VN.t8 167.875
R2374 VN.n8 VN.t3 167.875
R2375 VN.n22 VN.t2 167.875
R2376 VN.n29 VN.t6 167.875
R2377 VN.n46 VN.t9 167.875
R2378 VN.n39 VN.t0 167.875
R2379 VN.n53 VN.t4 167.875
R2380 VN.n60 VN.t1 167.875
R2381 VN.n59 VN.n31 161.3
R2382 VN.n58 VN.n57 161.3
R2383 VN.n56 VN.n32 161.3
R2384 VN.n55 VN.n54 161.3
R2385 VN.n52 VN.n33 161.3
R2386 VN.n51 VN.n50 161.3
R2387 VN.n49 VN.n34 161.3
R2388 VN.n48 VN.n47 161.3
R2389 VN.n46 VN.n35 161.3
R2390 VN.n45 VN.n44 161.3
R2391 VN.n43 VN.n36 161.3
R2392 VN.n42 VN.n41 161.3
R2393 VN.n40 VN.n37 161.3
R2394 VN.n28 VN.n0 161.3
R2395 VN.n27 VN.n26 161.3
R2396 VN.n25 VN.n1 161.3
R2397 VN.n24 VN.n23 161.3
R2398 VN.n21 VN.n2 161.3
R2399 VN.n20 VN.n19 161.3
R2400 VN.n18 VN.n3 161.3
R2401 VN.n17 VN.n16 161.3
R2402 VN.n15 VN.n4 161.3
R2403 VN.n14 VN.n13 161.3
R2404 VN.n12 VN.n5 161.3
R2405 VN.n11 VN.n10 161.3
R2406 VN.n9 VN.n6 161.3
R2407 VN.n8 VN.n7 63.3281
R2408 VN.n39 VN.n38 63.3281
R2409 VN.n27 VN.n1 52.1486
R2410 VN.n58 VN.n32 52.1486
R2411 VN VN.n61 48.9721
R2412 VN.n10 VN.n5 44.3785
R2413 VN.n20 VN.n3 44.3785
R2414 VN.n41 VN.n36 44.3785
R2415 VN.n51 VN.n34 44.3785
R2416 VN.n14 VN.n5 36.6083
R2417 VN.n16 VN.n3 36.6083
R2418 VN.n45 VN.n36 36.6083
R2419 VN.n47 VN.n34 36.6083
R2420 VN.n23 VN.n1 28.8382
R2421 VN.n54 VN.n32 28.8382
R2422 VN.n10 VN.n9 24.4675
R2423 VN.n15 VN.n14 24.4675
R2424 VN.n16 VN.n15 24.4675
R2425 VN.n21 VN.n20 24.4675
R2426 VN.n28 VN.n27 24.4675
R2427 VN.n41 VN.n40 24.4675
R2428 VN.n47 VN.n46 24.4675
R2429 VN.n46 VN.n45 24.4675
R2430 VN.n52 VN.n51 24.4675
R2431 VN.n59 VN.n58 24.4675
R2432 VN.n23 VN.n22 20.5528
R2433 VN.n54 VN.n53 20.5528
R2434 VN.n38 VN.n37 18.0704
R2435 VN.n7 VN.n6 18.0704
R2436 VN.n29 VN.n28 7.82994
R2437 VN.n60 VN.n59 7.82994
R2438 VN.n9 VN.n8 3.91522
R2439 VN.n22 VN.n21 3.91522
R2440 VN.n40 VN.n39 3.91522
R2441 VN.n53 VN.n52 3.91522
R2442 VN.n61 VN.n31 0.189894
R2443 VN.n57 VN.n31 0.189894
R2444 VN.n57 VN.n56 0.189894
R2445 VN.n56 VN.n55 0.189894
R2446 VN.n55 VN.n33 0.189894
R2447 VN.n50 VN.n33 0.189894
R2448 VN.n50 VN.n49 0.189894
R2449 VN.n49 VN.n48 0.189894
R2450 VN.n48 VN.n35 0.189894
R2451 VN.n44 VN.n35 0.189894
R2452 VN.n44 VN.n43 0.189894
R2453 VN.n43 VN.n42 0.189894
R2454 VN.n42 VN.n37 0.189894
R2455 VN.n11 VN.n6 0.189894
R2456 VN.n12 VN.n11 0.189894
R2457 VN.n13 VN.n12 0.189894
R2458 VN.n13 VN.n4 0.189894
R2459 VN.n17 VN.n4 0.189894
R2460 VN.n18 VN.n17 0.189894
R2461 VN.n19 VN.n18 0.189894
R2462 VN.n19 VN.n2 0.189894
R2463 VN.n24 VN.n2 0.189894
R2464 VN.n25 VN.n24 0.189894
R2465 VN.n26 VN.n25 0.189894
R2466 VN.n26 VN.n0 0.189894
R2467 VN.n30 VN.n0 0.189894
R2468 VN VN.n30 0.0516364
R2469 VDD2.n129 VDD2.n69 289.615
R2470 VDD2.n60 VDD2.n0 289.615
R2471 VDD2.n130 VDD2.n129 185
R2472 VDD2.n128 VDD2.n127 185
R2473 VDD2.n73 VDD2.n72 185
R2474 VDD2.n122 VDD2.n121 185
R2475 VDD2.n120 VDD2.n119 185
R2476 VDD2.n77 VDD2.n76 185
R2477 VDD2.n114 VDD2.n113 185
R2478 VDD2.n112 VDD2.n79 185
R2479 VDD2.n111 VDD2.n110 185
R2480 VDD2.n82 VDD2.n80 185
R2481 VDD2.n105 VDD2.n104 185
R2482 VDD2.n103 VDD2.n102 185
R2483 VDD2.n86 VDD2.n85 185
R2484 VDD2.n97 VDD2.n96 185
R2485 VDD2.n95 VDD2.n94 185
R2486 VDD2.n90 VDD2.n89 185
R2487 VDD2.n20 VDD2.n19 185
R2488 VDD2.n25 VDD2.n24 185
R2489 VDD2.n27 VDD2.n26 185
R2490 VDD2.n16 VDD2.n15 185
R2491 VDD2.n33 VDD2.n32 185
R2492 VDD2.n35 VDD2.n34 185
R2493 VDD2.n12 VDD2.n11 185
R2494 VDD2.n42 VDD2.n41 185
R2495 VDD2.n43 VDD2.n10 185
R2496 VDD2.n45 VDD2.n44 185
R2497 VDD2.n8 VDD2.n7 185
R2498 VDD2.n51 VDD2.n50 185
R2499 VDD2.n53 VDD2.n52 185
R2500 VDD2.n4 VDD2.n3 185
R2501 VDD2.n59 VDD2.n58 185
R2502 VDD2.n61 VDD2.n60 185
R2503 VDD2.n91 VDD2.t8 149.524
R2504 VDD2.n21 VDD2.t4 149.524
R2505 VDD2.n129 VDD2.n128 104.615
R2506 VDD2.n128 VDD2.n72 104.615
R2507 VDD2.n121 VDD2.n72 104.615
R2508 VDD2.n121 VDD2.n120 104.615
R2509 VDD2.n120 VDD2.n76 104.615
R2510 VDD2.n113 VDD2.n76 104.615
R2511 VDD2.n113 VDD2.n112 104.615
R2512 VDD2.n112 VDD2.n111 104.615
R2513 VDD2.n111 VDD2.n80 104.615
R2514 VDD2.n104 VDD2.n80 104.615
R2515 VDD2.n104 VDD2.n103 104.615
R2516 VDD2.n103 VDD2.n85 104.615
R2517 VDD2.n96 VDD2.n85 104.615
R2518 VDD2.n96 VDD2.n95 104.615
R2519 VDD2.n95 VDD2.n89 104.615
R2520 VDD2.n25 VDD2.n19 104.615
R2521 VDD2.n26 VDD2.n25 104.615
R2522 VDD2.n26 VDD2.n15 104.615
R2523 VDD2.n33 VDD2.n15 104.615
R2524 VDD2.n34 VDD2.n33 104.615
R2525 VDD2.n34 VDD2.n11 104.615
R2526 VDD2.n42 VDD2.n11 104.615
R2527 VDD2.n43 VDD2.n42 104.615
R2528 VDD2.n44 VDD2.n43 104.615
R2529 VDD2.n44 VDD2.n7 104.615
R2530 VDD2.n51 VDD2.n7 104.615
R2531 VDD2.n52 VDD2.n51 104.615
R2532 VDD2.n52 VDD2.n3 104.615
R2533 VDD2.n59 VDD2.n3 104.615
R2534 VDD2.n60 VDD2.n59 104.615
R2535 VDD2.n68 VDD2.n67 64.5268
R2536 VDD2 VDD2.n137 64.524
R2537 VDD2.n136 VDD2.n135 63.2375
R2538 VDD2.n66 VDD2.n65 63.2374
R2539 VDD2.t8 VDD2.n89 52.3082
R2540 VDD2.t4 VDD2.n19 52.3082
R2541 VDD2.n66 VDD2.n64 52.0148
R2542 VDD2.n134 VDD2.n133 50.2217
R2543 VDD2.n134 VDD2.n68 42.7412
R2544 VDD2.n114 VDD2.n79 13.1884
R2545 VDD2.n45 VDD2.n10 13.1884
R2546 VDD2.n115 VDD2.n77 12.8005
R2547 VDD2.n110 VDD2.n81 12.8005
R2548 VDD2.n41 VDD2.n40 12.8005
R2549 VDD2.n46 VDD2.n8 12.8005
R2550 VDD2.n119 VDD2.n118 12.0247
R2551 VDD2.n109 VDD2.n82 12.0247
R2552 VDD2.n39 VDD2.n12 12.0247
R2553 VDD2.n50 VDD2.n49 12.0247
R2554 VDD2.n122 VDD2.n75 11.249
R2555 VDD2.n106 VDD2.n105 11.249
R2556 VDD2.n36 VDD2.n35 11.249
R2557 VDD2.n53 VDD2.n6 11.249
R2558 VDD2.n123 VDD2.n73 10.4732
R2559 VDD2.n102 VDD2.n84 10.4732
R2560 VDD2.n32 VDD2.n14 10.4732
R2561 VDD2.n54 VDD2.n4 10.4732
R2562 VDD2.n91 VDD2.n90 10.2747
R2563 VDD2.n21 VDD2.n20 10.2747
R2564 VDD2.n127 VDD2.n126 9.69747
R2565 VDD2.n101 VDD2.n86 9.69747
R2566 VDD2.n31 VDD2.n16 9.69747
R2567 VDD2.n58 VDD2.n57 9.69747
R2568 VDD2.n133 VDD2.n132 9.45567
R2569 VDD2.n64 VDD2.n63 9.45567
R2570 VDD2.n93 VDD2.n92 9.3005
R2571 VDD2.n88 VDD2.n87 9.3005
R2572 VDD2.n99 VDD2.n98 9.3005
R2573 VDD2.n101 VDD2.n100 9.3005
R2574 VDD2.n84 VDD2.n83 9.3005
R2575 VDD2.n107 VDD2.n106 9.3005
R2576 VDD2.n109 VDD2.n108 9.3005
R2577 VDD2.n81 VDD2.n78 9.3005
R2578 VDD2.n132 VDD2.n131 9.3005
R2579 VDD2.n71 VDD2.n70 9.3005
R2580 VDD2.n126 VDD2.n125 9.3005
R2581 VDD2.n124 VDD2.n123 9.3005
R2582 VDD2.n75 VDD2.n74 9.3005
R2583 VDD2.n118 VDD2.n117 9.3005
R2584 VDD2.n116 VDD2.n115 9.3005
R2585 VDD2.n63 VDD2.n62 9.3005
R2586 VDD2.n2 VDD2.n1 9.3005
R2587 VDD2.n57 VDD2.n56 9.3005
R2588 VDD2.n55 VDD2.n54 9.3005
R2589 VDD2.n6 VDD2.n5 9.3005
R2590 VDD2.n49 VDD2.n48 9.3005
R2591 VDD2.n47 VDD2.n46 9.3005
R2592 VDD2.n23 VDD2.n22 9.3005
R2593 VDD2.n18 VDD2.n17 9.3005
R2594 VDD2.n29 VDD2.n28 9.3005
R2595 VDD2.n31 VDD2.n30 9.3005
R2596 VDD2.n14 VDD2.n13 9.3005
R2597 VDD2.n37 VDD2.n36 9.3005
R2598 VDD2.n39 VDD2.n38 9.3005
R2599 VDD2.n40 VDD2.n9 9.3005
R2600 VDD2.n130 VDD2.n71 8.92171
R2601 VDD2.n98 VDD2.n97 8.92171
R2602 VDD2.n28 VDD2.n27 8.92171
R2603 VDD2.n61 VDD2.n2 8.92171
R2604 VDD2.n131 VDD2.n69 8.14595
R2605 VDD2.n94 VDD2.n88 8.14595
R2606 VDD2.n24 VDD2.n18 8.14595
R2607 VDD2.n62 VDD2.n0 8.14595
R2608 VDD2.n93 VDD2.n90 7.3702
R2609 VDD2.n23 VDD2.n20 7.3702
R2610 VDD2.n133 VDD2.n69 5.81868
R2611 VDD2.n94 VDD2.n93 5.81868
R2612 VDD2.n24 VDD2.n23 5.81868
R2613 VDD2.n64 VDD2.n0 5.81868
R2614 VDD2.n131 VDD2.n130 5.04292
R2615 VDD2.n97 VDD2.n88 5.04292
R2616 VDD2.n27 VDD2.n18 5.04292
R2617 VDD2.n62 VDD2.n61 5.04292
R2618 VDD2.n127 VDD2.n71 4.26717
R2619 VDD2.n98 VDD2.n86 4.26717
R2620 VDD2.n28 VDD2.n16 4.26717
R2621 VDD2.n58 VDD2.n2 4.26717
R2622 VDD2.n126 VDD2.n73 3.49141
R2623 VDD2.n102 VDD2.n101 3.49141
R2624 VDD2.n32 VDD2.n31 3.49141
R2625 VDD2.n57 VDD2.n4 3.49141
R2626 VDD2.n92 VDD2.n91 2.84303
R2627 VDD2.n22 VDD2.n21 2.84303
R2628 VDD2.n123 VDD2.n122 2.71565
R2629 VDD2.n105 VDD2.n84 2.71565
R2630 VDD2.n35 VDD2.n14 2.71565
R2631 VDD2.n54 VDD2.n53 2.71565
R2632 VDD2.n119 VDD2.n75 1.93989
R2633 VDD2.n106 VDD2.n82 1.93989
R2634 VDD2.n36 VDD2.n12 1.93989
R2635 VDD2.n50 VDD2.n6 1.93989
R2636 VDD2.n136 VDD2.n134 1.7936
R2637 VDD2.n137 VDD2.t9 1.62478
R2638 VDD2.n137 VDD2.t2 1.62478
R2639 VDD2.n135 VDD2.t5 1.62478
R2640 VDD2.n135 VDD2.t0 1.62478
R2641 VDD2.n67 VDD2.t7 1.62478
R2642 VDD2.n67 VDD2.t3 1.62478
R2643 VDD2.n65 VDD2.t6 1.62478
R2644 VDD2.n65 VDD2.t1 1.62478
R2645 VDD2.n118 VDD2.n77 1.16414
R2646 VDD2.n110 VDD2.n109 1.16414
R2647 VDD2.n41 VDD2.n39 1.16414
R2648 VDD2.n49 VDD2.n8 1.16414
R2649 VDD2 VDD2.n136 0.506965
R2650 VDD2.n68 VDD2.n66 0.39343
R2651 VDD2.n115 VDD2.n114 0.388379
R2652 VDD2.n81 VDD2.n79 0.388379
R2653 VDD2.n40 VDD2.n10 0.388379
R2654 VDD2.n46 VDD2.n45 0.388379
R2655 VDD2.n132 VDD2.n70 0.155672
R2656 VDD2.n125 VDD2.n70 0.155672
R2657 VDD2.n125 VDD2.n124 0.155672
R2658 VDD2.n124 VDD2.n74 0.155672
R2659 VDD2.n117 VDD2.n74 0.155672
R2660 VDD2.n117 VDD2.n116 0.155672
R2661 VDD2.n116 VDD2.n78 0.155672
R2662 VDD2.n108 VDD2.n78 0.155672
R2663 VDD2.n108 VDD2.n107 0.155672
R2664 VDD2.n107 VDD2.n83 0.155672
R2665 VDD2.n100 VDD2.n83 0.155672
R2666 VDD2.n100 VDD2.n99 0.155672
R2667 VDD2.n99 VDD2.n87 0.155672
R2668 VDD2.n92 VDD2.n87 0.155672
R2669 VDD2.n22 VDD2.n17 0.155672
R2670 VDD2.n29 VDD2.n17 0.155672
R2671 VDD2.n30 VDD2.n29 0.155672
R2672 VDD2.n30 VDD2.n13 0.155672
R2673 VDD2.n37 VDD2.n13 0.155672
R2674 VDD2.n38 VDD2.n37 0.155672
R2675 VDD2.n38 VDD2.n9 0.155672
R2676 VDD2.n47 VDD2.n9 0.155672
R2677 VDD2.n48 VDD2.n47 0.155672
R2678 VDD2.n48 VDD2.n5 0.155672
R2679 VDD2.n55 VDD2.n5 0.155672
R2680 VDD2.n56 VDD2.n55 0.155672
R2681 VDD2.n56 VDD2.n1 0.155672
R2682 VDD2.n63 VDD2.n1 0.155672
C0 VN VDD2 9.84891f
C1 VTAIL VDD2 10.7667f
C2 VN VDD1 0.151243f
C3 VTAIL VDD1 10.7227f
C4 VDD1 VDD2 1.62039f
C5 VP VN 7.177751f
C6 VP VTAIL 10.141901f
C7 VP VDD2 0.475062f
C8 VN VTAIL 10.127501f
C9 VP VDD1 10.1687f
C10 VDD2 B 6.233392f
C11 VDD1 B 6.213834f
C12 VTAIL B 7.586165f
C13 VN B 14.15492f
C14 VP B 12.566099f
C15 VDD2.n0 B 0.032386f
C16 VDD2.n1 B 0.022292f
C17 VDD2.n2 B 0.011979f
C18 VDD2.n3 B 0.028314f
C19 VDD2.n4 B 0.012684f
C20 VDD2.n5 B 0.022292f
C21 VDD2.n6 B 0.011979f
C22 VDD2.n7 B 0.028314f
C23 VDD2.n8 B 0.012684f
C24 VDD2.n9 B 0.022292f
C25 VDD2.n10 B 0.012331f
C26 VDD2.n11 B 0.028314f
C27 VDD2.n12 B 0.012684f
C28 VDD2.n13 B 0.022292f
C29 VDD2.n14 B 0.011979f
C30 VDD2.n15 B 0.028314f
C31 VDD2.n16 B 0.012684f
C32 VDD2.n17 B 0.022292f
C33 VDD2.n18 B 0.011979f
C34 VDD2.n19 B 0.021235f
C35 VDD2.n20 B 0.020015f
C36 VDD2.t4 B 0.047843f
C37 VDD2.n21 B 0.16235f
C38 VDD2.n22 B 1.14344f
C39 VDD2.n23 B 0.011979f
C40 VDD2.n24 B 0.012684f
C41 VDD2.n25 B 0.028314f
C42 VDD2.n26 B 0.028314f
C43 VDD2.n27 B 0.012684f
C44 VDD2.n28 B 0.011979f
C45 VDD2.n29 B 0.022292f
C46 VDD2.n30 B 0.022292f
C47 VDD2.n31 B 0.011979f
C48 VDD2.n32 B 0.012684f
C49 VDD2.n33 B 0.028314f
C50 VDD2.n34 B 0.028314f
C51 VDD2.n35 B 0.012684f
C52 VDD2.n36 B 0.011979f
C53 VDD2.n37 B 0.022292f
C54 VDD2.n38 B 0.022292f
C55 VDD2.n39 B 0.011979f
C56 VDD2.n40 B 0.011979f
C57 VDD2.n41 B 0.012684f
C58 VDD2.n42 B 0.028314f
C59 VDD2.n43 B 0.028314f
C60 VDD2.n44 B 0.028314f
C61 VDD2.n45 B 0.012331f
C62 VDD2.n46 B 0.011979f
C63 VDD2.n47 B 0.022292f
C64 VDD2.n48 B 0.022292f
C65 VDD2.n49 B 0.011979f
C66 VDD2.n50 B 0.012684f
C67 VDD2.n51 B 0.028314f
C68 VDD2.n52 B 0.028314f
C69 VDD2.n53 B 0.012684f
C70 VDD2.n54 B 0.011979f
C71 VDD2.n55 B 0.022292f
C72 VDD2.n56 B 0.022292f
C73 VDD2.n57 B 0.011979f
C74 VDD2.n58 B 0.012684f
C75 VDD2.n59 B 0.028314f
C76 VDD2.n60 B 0.063156f
C77 VDD2.n61 B 0.012684f
C78 VDD2.n62 B 0.011979f
C79 VDD2.n63 B 0.053659f
C80 VDD2.n64 B 0.056932f
C81 VDD2.t6 B 0.214738f
C82 VDD2.t1 B 0.214738f
C83 VDD2.n65 B 1.91633f
C84 VDD2.n66 B 0.508979f
C85 VDD2.t7 B 0.214738f
C86 VDD2.t3 B 0.214738f
C87 VDD2.n67 B 1.92461f
C88 VDD2.n68 B 2.204f
C89 VDD2.n69 B 0.032386f
C90 VDD2.n70 B 0.022292f
C91 VDD2.n71 B 0.011979f
C92 VDD2.n72 B 0.028314f
C93 VDD2.n73 B 0.012684f
C94 VDD2.n74 B 0.022292f
C95 VDD2.n75 B 0.011979f
C96 VDD2.n76 B 0.028314f
C97 VDD2.n77 B 0.012684f
C98 VDD2.n78 B 0.022292f
C99 VDD2.n79 B 0.012331f
C100 VDD2.n80 B 0.028314f
C101 VDD2.n81 B 0.011979f
C102 VDD2.n82 B 0.012684f
C103 VDD2.n83 B 0.022292f
C104 VDD2.n84 B 0.011979f
C105 VDD2.n85 B 0.028314f
C106 VDD2.n86 B 0.012684f
C107 VDD2.n87 B 0.022292f
C108 VDD2.n88 B 0.011979f
C109 VDD2.n89 B 0.021235f
C110 VDD2.n90 B 0.020015f
C111 VDD2.t8 B 0.047843f
C112 VDD2.n91 B 0.16235f
C113 VDD2.n92 B 1.14344f
C114 VDD2.n93 B 0.011979f
C115 VDD2.n94 B 0.012684f
C116 VDD2.n95 B 0.028314f
C117 VDD2.n96 B 0.028314f
C118 VDD2.n97 B 0.012684f
C119 VDD2.n98 B 0.011979f
C120 VDD2.n99 B 0.022292f
C121 VDD2.n100 B 0.022292f
C122 VDD2.n101 B 0.011979f
C123 VDD2.n102 B 0.012684f
C124 VDD2.n103 B 0.028314f
C125 VDD2.n104 B 0.028314f
C126 VDD2.n105 B 0.012684f
C127 VDD2.n106 B 0.011979f
C128 VDD2.n107 B 0.022292f
C129 VDD2.n108 B 0.022292f
C130 VDD2.n109 B 0.011979f
C131 VDD2.n110 B 0.012684f
C132 VDD2.n111 B 0.028314f
C133 VDD2.n112 B 0.028314f
C134 VDD2.n113 B 0.028314f
C135 VDD2.n114 B 0.012331f
C136 VDD2.n115 B 0.011979f
C137 VDD2.n116 B 0.022292f
C138 VDD2.n117 B 0.022292f
C139 VDD2.n118 B 0.011979f
C140 VDD2.n119 B 0.012684f
C141 VDD2.n120 B 0.028314f
C142 VDD2.n121 B 0.028314f
C143 VDD2.n122 B 0.012684f
C144 VDD2.n123 B 0.011979f
C145 VDD2.n124 B 0.022292f
C146 VDD2.n125 B 0.022292f
C147 VDD2.n126 B 0.011979f
C148 VDD2.n127 B 0.012684f
C149 VDD2.n128 B 0.028314f
C150 VDD2.n129 B 0.063156f
C151 VDD2.n130 B 0.012684f
C152 VDD2.n131 B 0.011979f
C153 VDD2.n132 B 0.053659f
C154 VDD2.n133 B 0.05097f
C155 VDD2.n134 B 2.29713f
C156 VDD2.t5 B 0.214738f
C157 VDD2.t0 B 0.214738f
C158 VDD2.n135 B 1.91634f
C159 VDD2.n136 B 0.348829f
C160 VDD2.t9 B 0.214738f
C161 VDD2.t2 B 0.214738f
C162 VDD2.n137 B 1.92458f
C163 VN.n0 B 0.02731f
C164 VN.t6 B 1.58806f
C165 VN.n1 B 0.027585f
C166 VN.n2 B 0.02731f
C167 VN.t2 B 1.58806f
C168 VN.n3 B 0.022644f
C169 VN.n4 B 0.02731f
C170 VN.t8 B 1.58806f
C171 VN.n5 B 0.022644f
C172 VN.n6 B 0.177148f
C173 VN.t3 B 1.58806f
C174 VN.t5 B 1.69934f
C175 VN.n7 B 0.636712f
C176 VN.n8 B 0.618991f
C177 VN.n9 B 0.029791f
C178 VN.n10 B 0.052927f
C179 VN.n11 B 0.02731f
C180 VN.n12 B 0.02731f
C181 VN.n13 B 0.02731f
C182 VN.n14 B 0.055065f
C183 VN.n15 B 0.595136f
C184 VN.n16 B 0.055065f
C185 VN.n17 B 0.02731f
C186 VN.n18 B 0.02731f
C187 VN.n19 B 0.02731f
C188 VN.n20 B 0.052927f
C189 VN.n21 B 0.029791f
C190 VN.n22 B 0.569366f
C191 VN.n23 B 0.05f
C192 VN.n24 B 0.02731f
C193 VN.n25 B 0.02731f
C194 VN.n26 B 0.02731f
C195 VN.n27 B 0.04903f
C196 VN.n28 B 0.033812f
C197 VN.n29 B 0.634186f
C198 VN.n30 B 0.02785f
C199 VN.n31 B 0.02731f
C200 VN.t1 B 1.58806f
C201 VN.n32 B 0.027585f
C202 VN.n33 B 0.02731f
C203 VN.t4 B 1.58806f
C204 VN.n34 B 0.022644f
C205 VN.n35 B 0.02731f
C206 VN.t9 B 1.58806f
C207 VN.n36 B 0.022644f
C208 VN.n37 B 0.177148f
C209 VN.t0 B 1.58806f
C210 VN.t7 B 1.69934f
C211 VN.n38 B 0.636712f
C212 VN.n39 B 0.618991f
C213 VN.n40 B 0.029791f
C214 VN.n41 B 0.052927f
C215 VN.n42 B 0.02731f
C216 VN.n43 B 0.02731f
C217 VN.n44 B 0.02731f
C218 VN.n45 B 0.055065f
C219 VN.n46 B 0.595136f
C220 VN.n47 B 0.055065f
C221 VN.n48 B 0.02731f
C222 VN.n49 B 0.02731f
C223 VN.n50 B 0.02731f
C224 VN.n51 B 0.052927f
C225 VN.n52 B 0.029791f
C226 VN.n53 B 0.569366f
C227 VN.n54 B 0.05f
C228 VN.n55 B 0.02731f
C229 VN.n56 B 0.02731f
C230 VN.n57 B 0.02731f
C231 VN.n58 B 0.04903f
C232 VN.n59 B 0.033812f
C233 VN.n60 B 0.634186f
C234 VN.n61 B 1.44634f
C235 VTAIL.t6 B 0.235205f
C236 VTAIL.t0 B 0.235205f
C237 VTAIL.n0 B 2.02858f
C238 VTAIL.n1 B 0.45626f
C239 VTAIL.n2 B 0.035473f
C240 VTAIL.n3 B 0.024417f
C241 VTAIL.n4 B 0.01312f
C242 VTAIL.n5 B 0.031012f
C243 VTAIL.n6 B 0.013892f
C244 VTAIL.n7 B 0.024417f
C245 VTAIL.n8 B 0.01312f
C246 VTAIL.n9 B 0.031012f
C247 VTAIL.n10 B 0.013892f
C248 VTAIL.n11 B 0.024417f
C249 VTAIL.n12 B 0.013506f
C250 VTAIL.n13 B 0.031012f
C251 VTAIL.n14 B 0.013892f
C252 VTAIL.n15 B 0.024417f
C253 VTAIL.n16 B 0.01312f
C254 VTAIL.n17 B 0.031012f
C255 VTAIL.n18 B 0.013892f
C256 VTAIL.n19 B 0.024417f
C257 VTAIL.n20 B 0.01312f
C258 VTAIL.n21 B 0.023259f
C259 VTAIL.n22 B 0.021923f
C260 VTAIL.t12 B 0.052403f
C261 VTAIL.n23 B 0.177823f
C262 VTAIL.n24 B 1.25242f
C263 VTAIL.n25 B 0.01312f
C264 VTAIL.n26 B 0.013892f
C265 VTAIL.n27 B 0.031012f
C266 VTAIL.n28 B 0.031012f
C267 VTAIL.n29 B 0.013892f
C268 VTAIL.n30 B 0.01312f
C269 VTAIL.n31 B 0.024417f
C270 VTAIL.n32 B 0.024417f
C271 VTAIL.n33 B 0.01312f
C272 VTAIL.n34 B 0.013892f
C273 VTAIL.n35 B 0.031012f
C274 VTAIL.n36 B 0.031012f
C275 VTAIL.n37 B 0.013892f
C276 VTAIL.n38 B 0.01312f
C277 VTAIL.n39 B 0.024417f
C278 VTAIL.n40 B 0.024417f
C279 VTAIL.n41 B 0.01312f
C280 VTAIL.n42 B 0.01312f
C281 VTAIL.n43 B 0.013892f
C282 VTAIL.n44 B 0.031012f
C283 VTAIL.n45 B 0.031012f
C284 VTAIL.n46 B 0.031012f
C285 VTAIL.n47 B 0.013506f
C286 VTAIL.n48 B 0.01312f
C287 VTAIL.n49 B 0.024417f
C288 VTAIL.n50 B 0.024417f
C289 VTAIL.n51 B 0.01312f
C290 VTAIL.n52 B 0.013892f
C291 VTAIL.n53 B 0.031012f
C292 VTAIL.n54 B 0.031012f
C293 VTAIL.n55 B 0.013892f
C294 VTAIL.n56 B 0.01312f
C295 VTAIL.n57 B 0.024417f
C296 VTAIL.n58 B 0.024417f
C297 VTAIL.n59 B 0.01312f
C298 VTAIL.n60 B 0.013892f
C299 VTAIL.n61 B 0.031012f
C300 VTAIL.n62 B 0.069175f
C301 VTAIL.n63 B 0.013892f
C302 VTAIL.n64 B 0.01312f
C303 VTAIL.n65 B 0.058773f
C304 VTAIL.n66 B 0.038986f
C305 VTAIL.n67 B 0.270749f
C306 VTAIL.t14 B 0.235205f
C307 VTAIL.t16 B 0.235205f
C308 VTAIL.n68 B 2.02858f
C309 VTAIL.n69 B 0.520523f
C310 VTAIL.t11 B 0.235205f
C311 VTAIL.t10 B 0.235205f
C312 VTAIL.n70 B 2.02858f
C313 VTAIL.n71 B 1.82005f
C314 VTAIL.t7 B 0.235205f
C315 VTAIL.t4 B 0.235205f
C316 VTAIL.n72 B 2.02859f
C317 VTAIL.n73 B 1.82004f
C318 VTAIL.t5 B 0.235205f
C319 VTAIL.t9 B 0.235205f
C320 VTAIL.n74 B 2.02859f
C321 VTAIL.n75 B 0.520512f
C322 VTAIL.n76 B 0.035473f
C323 VTAIL.n77 B 0.024417f
C324 VTAIL.n78 B 0.01312f
C325 VTAIL.n79 B 0.031012f
C326 VTAIL.n80 B 0.013892f
C327 VTAIL.n81 B 0.024417f
C328 VTAIL.n82 B 0.01312f
C329 VTAIL.n83 B 0.031012f
C330 VTAIL.n84 B 0.013892f
C331 VTAIL.n85 B 0.024417f
C332 VTAIL.n86 B 0.013506f
C333 VTAIL.n87 B 0.031012f
C334 VTAIL.n88 B 0.01312f
C335 VTAIL.n89 B 0.013892f
C336 VTAIL.n90 B 0.024417f
C337 VTAIL.n91 B 0.01312f
C338 VTAIL.n92 B 0.031012f
C339 VTAIL.n93 B 0.013892f
C340 VTAIL.n94 B 0.024417f
C341 VTAIL.n95 B 0.01312f
C342 VTAIL.n96 B 0.023259f
C343 VTAIL.n97 B 0.021923f
C344 VTAIL.t3 B 0.052403f
C345 VTAIL.n98 B 0.177823f
C346 VTAIL.n99 B 1.25242f
C347 VTAIL.n100 B 0.01312f
C348 VTAIL.n101 B 0.013892f
C349 VTAIL.n102 B 0.031012f
C350 VTAIL.n103 B 0.031012f
C351 VTAIL.n104 B 0.013892f
C352 VTAIL.n105 B 0.01312f
C353 VTAIL.n106 B 0.024417f
C354 VTAIL.n107 B 0.024417f
C355 VTAIL.n108 B 0.01312f
C356 VTAIL.n109 B 0.013892f
C357 VTAIL.n110 B 0.031012f
C358 VTAIL.n111 B 0.031012f
C359 VTAIL.n112 B 0.013892f
C360 VTAIL.n113 B 0.01312f
C361 VTAIL.n114 B 0.024417f
C362 VTAIL.n115 B 0.024417f
C363 VTAIL.n116 B 0.01312f
C364 VTAIL.n117 B 0.013892f
C365 VTAIL.n118 B 0.031012f
C366 VTAIL.n119 B 0.031012f
C367 VTAIL.n120 B 0.031012f
C368 VTAIL.n121 B 0.013506f
C369 VTAIL.n122 B 0.01312f
C370 VTAIL.n123 B 0.024417f
C371 VTAIL.n124 B 0.024417f
C372 VTAIL.n125 B 0.01312f
C373 VTAIL.n126 B 0.013892f
C374 VTAIL.n127 B 0.031012f
C375 VTAIL.n128 B 0.031012f
C376 VTAIL.n129 B 0.013892f
C377 VTAIL.n130 B 0.01312f
C378 VTAIL.n131 B 0.024417f
C379 VTAIL.n132 B 0.024417f
C380 VTAIL.n133 B 0.01312f
C381 VTAIL.n134 B 0.013892f
C382 VTAIL.n135 B 0.031012f
C383 VTAIL.n136 B 0.069175f
C384 VTAIL.n137 B 0.013892f
C385 VTAIL.n138 B 0.01312f
C386 VTAIL.n139 B 0.058773f
C387 VTAIL.n140 B 0.038986f
C388 VTAIL.n141 B 0.270749f
C389 VTAIL.t17 B 0.235205f
C390 VTAIL.t19 B 0.235205f
C391 VTAIL.n142 B 2.02859f
C392 VTAIL.n143 B 0.486939f
C393 VTAIL.t13 B 0.235205f
C394 VTAIL.t18 B 0.235205f
C395 VTAIL.n144 B 2.02859f
C396 VTAIL.n145 B 0.520512f
C397 VTAIL.n146 B 0.035473f
C398 VTAIL.n147 B 0.024417f
C399 VTAIL.n148 B 0.01312f
C400 VTAIL.n149 B 0.031012f
C401 VTAIL.n150 B 0.013892f
C402 VTAIL.n151 B 0.024417f
C403 VTAIL.n152 B 0.01312f
C404 VTAIL.n153 B 0.031012f
C405 VTAIL.n154 B 0.013892f
C406 VTAIL.n155 B 0.024417f
C407 VTAIL.n156 B 0.013506f
C408 VTAIL.n157 B 0.031012f
C409 VTAIL.n158 B 0.01312f
C410 VTAIL.n159 B 0.013892f
C411 VTAIL.n160 B 0.024417f
C412 VTAIL.n161 B 0.01312f
C413 VTAIL.n162 B 0.031012f
C414 VTAIL.n163 B 0.013892f
C415 VTAIL.n164 B 0.024417f
C416 VTAIL.n165 B 0.01312f
C417 VTAIL.n166 B 0.023259f
C418 VTAIL.n167 B 0.021923f
C419 VTAIL.t15 B 0.052403f
C420 VTAIL.n168 B 0.177823f
C421 VTAIL.n169 B 1.25242f
C422 VTAIL.n170 B 0.01312f
C423 VTAIL.n171 B 0.013892f
C424 VTAIL.n172 B 0.031012f
C425 VTAIL.n173 B 0.031012f
C426 VTAIL.n174 B 0.013892f
C427 VTAIL.n175 B 0.01312f
C428 VTAIL.n176 B 0.024417f
C429 VTAIL.n177 B 0.024417f
C430 VTAIL.n178 B 0.01312f
C431 VTAIL.n179 B 0.013892f
C432 VTAIL.n180 B 0.031012f
C433 VTAIL.n181 B 0.031012f
C434 VTAIL.n182 B 0.013892f
C435 VTAIL.n183 B 0.01312f
C436 VTAIL.n184 B 0.024417f
C437 VTAIL.n185 B 0.024417f
C438 VTAIL.n186 B 0.01312f
C439 VTAIL.n187 B 0.013892f
C440 VTAIL.n188 B 0.031012f
C441 VTAIL.n189 B 0.031012f
C442 VTAIL.n190 B 0.031012f
C443 VTAIL.n191 B 0.013506f
C444 VTAIL.n192 B 0.01312f
C445 VTAIL.n193 B 0.024417f
C446 VTAIL.n194 B 0.024417f
C447 VTAIL.n195 B 0.01312f
C448 VTAIL.n196 B 0.013892f
C449 VTAIL.n197 B 0.031012f
C450 VTAIL.n198 B 0.031012f
C451 VTAIL.n199 B 0.013892f
C452 VTAIL.n200 B 0.01312f
C453 VTAIL.n201 B 0.024417f
C454 VTAIL.n202 B 0.024417f
C455 VTAIL.n203 B 0.01312f
C456 VTAIL.n204 B 0.013892f
C457 VTAIL.n205 B 0.031012f
C458 VTAIL.n206 B 0.069175f
C459 VTAIL.n207 B 0.013892f
C460 VTAIL.n208 B 0.01312f
C461 VTAIL.n209 B 0.058773f
C462 VTAIL.n210 B 0.038986f
C463 VTAIL.n211 B 1.46278f
C464 VTAIL.n212 B 0.035473f
C465 VTAIL.n213 B 0.024417f
C466 VTAIL.n214 B 0.01312f
C467 VTAIL.n215 B 0.031012f
C468 VTAIL.n216 B 0.013892f
C469 VTAIL.n217 B 0.024417f
C470 VTAIL.n218 B 0.01312f
C471 VTAIL.n219 B 0.031012f
C472 VTAIL.n220 B 0.013892f
C473 VTAIL.n221 B 0.024417f
C474 VTAIL.n222 B 0.013506f
C475 VTAIL.n223 B 0.031012f
C476 VTAIL.n224 B 0.013892f
C477 VTAIL.n225 B 0.024417f
C478 VTAIL.n226 B 0.01312f
C479 VTAIL.n227 B 0.031012f
C480 VTAIL.n228 B 0.013892f
C481 VTAIL.n229 B 0.024417f
C482 VTAIL.n230 B 0.01312f
C483 VTAIL.n231 B 0.023259f
C484 VTAIL.n232 B 0.021923f
C485 VTAIL.t8 B 0.052403f
C486 VTAIL.n233 B 0.177823f
C487 VTAIL.n234 B 1.25242f
C488 VTAIL.n235 B 0.01312f
C489 VTAIL.n236 B 0.013892f
C490 VTAIL.n237 B 0.031012f
C491 VTAIL.n238 B 0.031012f
C492 VTAIL.n239 B 0.013892f
C493 VTAIL.n240 B 0.01312f
C494 VTAIL.n241 B 0.024417f
C495 VTAIL.n242 B 0.024417f
C496 VTAIL.n243 B 0.01312f
C497 VTAIL.n244 B 0.013892f
C498 VTAIL.n245 B 0.031012f
C499 VTAIL.n246 B 0.031012f
C500 VTAIL.n247 B 0.013892f
C501 VTAIL.n248 B 0.01312f
C502 VTAIL.n249 B 0.024417f
C503 VTAIL.n250 B 0.024417f
C504 VTAIL.n251 B 0.01312f
C505 VTAIL.n252 B 0.01312f
C506 VTAIL.n253 B 0.013892f
C507 VTAIL.n254 B 0.031012f
C508 VTAIL.n255 B 0.031012f
C509 VTAIL.n256 B 0.031012f
C510 VTAIL.n257 B 0.013506f
C511 VTAIL.n258 B 0.01312f
C512 VTAIL.n259 B 0.024417f
C513 VTAIL.n260 B 0.024417f
C514 VTAIL.n261 B 0.01312f
C515 VTAIL.n262 B 0.013892f
C516 VTAIL.n263 B 0.031012f
C517 VTAIL.n264 B 0.031012f
C518 VTAIL.n265 B 0.013892f
C519 VTAIL.n266 B 0.01312f
C520 VTAIL.n267 B 0.024417f
C521 VTAIL.n268 B 0.024417f
C522 VTAIL.n269 B 0.01312f
C523 VTAIL.n270 B 0.013892f
C524 VTAIL.n271 B 0.031012f
C525 VTAIL.n272 B 0.069175f
C526 VTAIL.n273 B 0.013892f
C527 VTAIL.n274 B 0.01312f
C528 VTAIL.n275 B 0.058773f
C529 VTAIL.n276 B 0.038986f
C530 VTAIL.n277 B 1.46278f
C531 VTAIL.t1 B 0.235205f
C532 VTAIL.t2 B 0.235205f
C533 VTAIL.n278 B 2.02858f
C534 VTAIL.n279 B 0.410139f
C535 VDD1.n0 B 0.032727f
C536 VDD1.n1 B 0.022527f
C537 VDD1.n2 B 0.012105f
C538 VDD1.n3 B 0.028611f
C539 VDD1.n4 B 0.012817f
C540 VDD1.n5 B 0.022527f
C541 VDD1.n6 B 0.012105f
C542 VDD1.n7 B 0.028611f
C543 VDD1.n8 B 0.012817f
C544 VDD1.n9 B 0.022527f
C545 VDD1.n10 B 0.012461f
C546 VDD1.n11 B 0.028611f
C547 VDD1.n12 B 0.012105f
C548 VDD1.n13 B 0.012817f
C549 VDD1.n14 B 0.022527f
C550 VDD1.n15 B 0.012105f
C551 VDD1.n16 B 0.028611f
C552 VDD1.n17 B 0.012817f
C553 VDD1.n18 B 0.022527f
C554 VDD1.n19 B 0.012105f
C555 VDD1.n20 B 0.021459f
C556 VDD1.n21 B 0.020226f
C557 VDD1.t7 B 0.048346f
C558 VDD1.n22 B 0.164058f
C559 VDD1.n23 B 1.15547f
C560 VDD1.n24 B 0.012105f
C561 VDD1.n25 B 0.012817f
C562 VDD1.n26 B 0.028611f
C563 VDD1.n27 B 0.028611f
C564 VDD1.n28 B 0.012817f
C565 VDD1.n29 B 0.012105f
C566 VDD1.n30 B 0.022527f
C567 VDD1.n31 B 0.022527f
C568 VDD1.n32 B 0.012105f
C569 VDD1.n33 B 0.012817f
C570 VDD1.n34 B 0.028611f
C571 VDD1.n35 B 0.028611f
C572 VDD1.n36 B 0.012817f
C573 VDD1.n37 B 0.012105f
C574 VDD1.n38 B 0.022527f
C575 VDD1.n39 B 0.022527f
C576 VDD1.n40 B 0.012105f
C577 VDD1.n41 B 0.012817f
C578 VDD1.n42 B 0.028611f
C579 VDD1.n43 B 0.028611f
C580 VDD1.n44 B 0.028611f
C581 VDD1.n45 B 0.012461f
C582 VDD1.n46 B 0.012105f
C583 VDD1.n47 B 0.022527f
C584 VDD1.n48 B 0.022527f
C585 VDD1.n49 B 0.012105f
C586 VDD1.n50 B 0.012817f
C587 VDD1.n51 B 0.028611f
C588 VDD1.n52 B 0.028611f
C589 VDD1.n53 B 0.012817f
C590 VDD1.n54 B 0.012105f
C591 VDD1.n55 B 0.022527f
C592 VDD1.n56 B 0.022527f
C593 VDD1.n57 B 0.012105f
C594 VDD1.n58 B 0.012817f
C595 VDD1.n59 B 0.028611f
C596 VDD1.n60 B 0.06382f
C597 VDD1.n61 B 0.012817f
C598 VDD1.n62 B 0.012105f
C599 VDD1.n63 B 0.054224f
C600 VDD1.n64 B 0.057531f
C601 VDD1.t2 B 0.216998f
C602 VDD1.t5 B 0.216998f
C603 VDD1.n65 B 1.9365f
C604 VDD1.n66 B 0.52124f
C605 VDD1.n67 B 0.032727f
C606 VDD1.n68 B 0.022527f
C607 VDD1.n69 B 0.012105f
C608 VDD1.n70 B 0.028611f
C609 VDD1.n71 B 0.012817f
C610 VDD1.n72 B 0.022527f
C611 VDD1.n73 B 0.012105f
C612 VDD1.n74 B 0.028611f
C613 VDD1.n75 B 0.012817f
C614 VDD1.n76 B 0.022527f
C615 VDD1.n77 B 0.012461f
C616 VDD1.n78 B 0.028611f
C617 VDD1.n79 B 0.012817f
C618 VDD1.n80 B 0.022527f
C619 VDD1.n81 B 0.012105f
C620 VDD1.n82 B 0.028611f
C621 VDD1.n83 B 0.012817f
C622 VDD1.n84 B 0.022527f
C623 VDD1.n85 B 0.012105f
C624 VDD1.n86 B 0.021459f
C625 VDD1.n87 B 0.020226f
C626 VDD1.t9 B 0.048346f
C627 VDD1.n88 B 0.164058f
C628 VDD1.n89 B 1.15547f
C629 VDD1.n90 B 0.012105f
C630 VDD1.n91 B 0.012817f
C631 VDD1.n92 B 0.028611f
C632 VDD1.n93 B 0.028611f
C633 VDD1.n94 B 0.012817f
C634 VDD1.n95 B 0.012105f
C635 VDD1.n96 B 0.022527f
C636 VDD1.n97 B 0.022527f
C637 VDD1.n98 B 0.012105f
C638 VDD1.n99 B 0.012817f
C639 VDD1.n100 B 0.028611f
C640 VDD1.n101 B 0.028611f
C641 VDD1.n102 B 0.012817f
C642 VDD1.n103 B 0.012105f
C643 VDD1.n104 B 0.022527f
C644 VDD1.n105 B 0.022527f
C645 VDD1.n106 B 0.012105f
C646 VDD1.n107 B 0.012105f
C647 VDD1.n108 B 0.012817f
C648 VDD1.n109 B 0.028611f
C649 VDD1.n110 B 0.028611f
C650 VDD1.n111 B 0.028611f
C651 VDD1.n112 B 0.012461f
C652 VDD1.n113 B 0.012105f
C653 VDD1.n114 B 0.022527f
C654 VDD1.n115 B 0.022527f
C655 VDD1.n116 B 0.012105f
C656 VDD1.n117 B 0.012817f
C657 VDD1.n118 B 0.028611f
C658 VDD1.n119 B 0.028611f
C659 VDD1.n120 B 0.012817f
C660 VDD1.n121 B 0.012105f
C661 VDD1.n122 B 0.022527f
C662 VDD1.n123 B 0.022527f
C663 VDD1.n124 B 0.012105f
C664 VDD1.n125 B 0.012817f
C665 VDD1.n126 B 0.028611f
C666 VDD1.n127 B 0.06382f
C667 VDD1.n128 B 0.012817f
C668 VDD1.n129 B 0.012105f
C669 VDD1.n130 B 0.054224f
C670 VDD1.n131 B 0.057531f
C671 VDD1.t4 B 0.216998f
C672 VDD1.t8 B 0.216998f
C673 VDD1.n132 B 1.9365f
C674 VDD1.n133 B 0.514336f
C675 VDD1.t0 B 0.216998f
C676 VDD1.t6 B 0.216998f
C677 VDD1.n134 B 1.94487f
C678 VDD1.n135 B 2.31989f
C679 VDD1.t3 B 0.216998f
C680 VDD1.t1 B 0.216998f
C681 VDD1.n136 B 1.9365f
C682 VDD1.n137 B 2.55526f
C683 VP.n0 B 0.027753f
C684 VP.t7 B 1.61379f
C685 VP.n1 B 0.028032f
C686 VP.n2 B 0.027753f
C687 VP.t3 B 1.61379f
C688 VP.n3 B 0.023011f
C689 VP.n4 B 0.027753f
C690 VP.t5 B 1.61379f
C691 VP.n5 B 0.023011f
C692 VP.n6 B 0.027753f
C693 VP.t9 B 1.61379f
C694 VP.n7 B 0.028032f
C695 VP.n8 B 0.027753f
C696 VP.t8 B 1.61379f
C697 VP.n9 B 0.027753f
C698 VP.t4 B 1.61379f
C699 VP.n10 B 0.028032f
C700 VP.n11 B 0.027753f
C701 VP.t1 B 1.61379f
C702 VP.n12 B 0.023011f
C703 VP.n13 B 0.027753f
C704 VP.t6 B 1.61379f
C705 VP.n14 B 0.023011f
C706 VP.n15 B 0.180018f
C707 VP.t0 B 1.61379f
C708 VP.t2 B 1.72687f
C709 VP.n16 B 0.647026f
C710 VP.n17 B 0.629019f
C711 VP.n18 B 0.030274f
C712 VP.n19 B 0.053784f
C713 VP.n20 B 0.027753f
C714 VP.n21 B 0.027753f
C715 VP.n22 B 0.027753f
C716 VP.n23 B 0.055957f
C717 VP.n24 B 0.604777f
C718 VP.n25 B 0.055957f
C719 VP.n26 B 0.027753f
C720 VP.n27 B 0.027753f
C721 VP.n28 B 0.027753f
C722 VP.n29 B 0.053784f
C723 VP.n30 B 0.030274f
C724 VP.n31 B 0.57859f
C725 VP.n32 B 0.05081f
C726 VP.n33 B 0.027753f
C727 VP.n34 B 0.027753f
C728 VP.n35 B 0.027753f
C729 VP.n36 B 0.049824f
C730 VP.n37 B 0.034359f
C731 VP.n38 B 0.64446f
C732 VP.n39 B 1.4517f
C733 VP.n40 B 1.47223f
C734 VP.n41 B 0.64446f
C735 VP.n42 B 0.034359f
C736 VP.n43 B 0.049824f
C737 VP.n44 B 0.027753f
C738 VP.n45 B 0.027753f
C739 VP.n46 B 0.027753f
C740 VP.n47 B 0.05081f
C741 VP.n48 B 0.57859f
C742 VP.n49 B 0.030274f
C743 VP.n50 B 0.053784f
C744 VP.n51 B 0.027753f
C745 VP.n52 B 0.027753f
C746 VP.n53 B 0.027753f
C747 VP.n54 B 0.055957f
C748 VP.n55 B 0.604777f
C749 VP.n56 B 0.055957f
C750 VP.n57 B 0.027753f
C751 VP.n58 B 0.027753f
C752 VP.n59 B 0.027753f
C753 VP.n60 B 0.053784f
C754 VP.n61 B 0.030274f
C755 VP.n62 B 0.57859f
C756 VP.n63 B 0.05081f
C757 VP.n64 B 0.027753f
C758 VP.n65 B 0.027753f
C759 VP.n66 B 0.027753f
C760 VP.n67 B 0.049824f
C761 VP.n68 B 0.034359f
C762 VP.n69 B 0.64446f
C763 VP.n70 B 0.028302f
.ends

