* NGSPICE file created from diff_pair_sample_1437.ext - technology: sky130A

.subckt diff_pair_sample_1437 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=0 ps=0 w=3.18 l=2.72
X1 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=1.2402 ps=7.14 w=3.18 l=2.72
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=0 ps=0 w=3.18 l=2.72
X3 VDD1.t1 VP.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=1.2402 ps=7.14 w=3.18 l=2.72
X4 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=1.2402 ps=7.14 w=3.18 l=2.72
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=0 ps=0 w=3.18 l=2.72
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=0 ps=0 w=3.18 l=2.72
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2402 pd=7.14 as=1.2402 ps=7.14 w=3.18 l=2.72
R0 B.n345 B.n75 585
R1 B.n75 B.n50 585
R2 B.n347 B.n346 585
R3 B.n349 B.n74 585
R4 B.n352 B.n351 585
R5 B.n353 B.n73 585
R6 B.n355 B.n354 585
R7 B.n357 B.n72 585
R8 B.n360 B.n359 585
R9 B.n361 B.n71 585
R10 B.n363 B.n362 585
R11 B.n365 B.n70 585
R12 B.n368 B.n367 585
R13 B.n369 B.n69 585
R14 B.n371 B.n370 585
R15 B.n373 B.n68 585
R16 B.n376 B.n375 585
R17 B.n378 B.n65 585
R18 B.n380 B.n379 585
R19 B.n382 B.n64 585
R20 B.n385 B.n384 585
R21 B.n386 B.n63 585
R22 B.n388 B.n387 585
R23 B.n390 B.n62 585
R24 B.n393 B.n392 585
R25 B.n394 B.n59 585
R26 B.n397 B.n396 585
R27 B.n399 B.n58 585
R28 B.n402 B.n401 585
R29 B.n403 B.n57 585
R30 B.n405 B.n404 585
R31 B.n407 B.n56 585
R32 B.n410 B.n409 585
R33 B.n411 B.n55 585
R34 B.n413 B.n412 585
R35 B.n415 B.n54 585
R36 B.n418 B.n417 585
R37 B.n419 B.n53 585
R38 B.n421 B.n420 585
R39 B.n423 B.n52 585
R40 B.n426 B.n425 585
R41 B.n427 B.n51 585
R42 B.n344 B.n49 585
R43 B.n430 B.n49 585
R44 B.n343 B.n48 585
R45 B.n431 B.n48 585
R46 B.n342 B.n47 585
R47 B.n432 B.n47 585
R48 B.n341 B.n340 585
R49 B.n340 B.n43 585
R50 B.n339 B.n42 585
R51 B.n438 B.n42 585
R52 B.n338 B.n41 585
R53 B.n439 B.n41 585
R54 B.n337 B.n40 585
R55 B.n440 B.n40 585
R56 B.n336 B.n335 585
R57 B.n335 B.n39 585
R58 B.n334 B.n35 585
R59 B.n446 B.n35 585
R60 B.n333 B.n34 585
R61 B.n447 B.n34 585
R62 B.n332 B.n33 585
R63 B.n448 B.n33 585
R64 B.n331 B.n330 585
R65 B.n330 B.n29 585
R66 B.n329 B.n28 585
R67 B.n454 B.n28 585
R68 B.n328 B.n27 585
R69 B.n455 B.n27 585
R70 B.n327 B.n26 585
R71 B.n456 B.n26 585
R72 B.n326 B.n325 585
R73 B.n325 B.n22 585
R74 B.n324 B.n21 585
R75 B.n462 B.n21 585
R76 B.n323 B.n20 585
R77 B.n463 B.n20 585
R78 B.n322 B.n19 585
R79 B.n464 B.n19 585
R80 B.n321 B.n320 585
R81 B.n320 B.n18 585
R82 B.n319 B.n14 585
R83 B.n470 B.n14 585
R84 B.n318 B.n13 585
R85 B.n471 B.n13 585
R86 B.n317 B.n12 585
R87 B.n472 B.n12 585
R88 B.n316 B.n315 585
R89 B.n315 B.n8 585
R90 B.n314 B.n7 585
R91 B.n478 B.n7 585
R92 B.n313 B.n6 585
R93 B.n479 B.n6 585
R94 B.n312 B.n5 585
R95 B.n480 B.n5 585
R96 B.n311 B.n310 585
R97 B.n310 B.n4 585
R98 B.n309 B.n76 585
R99 B.n309 B.n308 585
R100 B.n299 B.n77 585
R101 B.n78 B.n77 585
R102 B.n301 B.n300 585
R103 B.n302 B.n301 585
R104 B.n298 B.n83 585
R105 B.n83 B.n82 585
R106 B.n297 B.n296 585
R107 B.n296 B.n295 585
R108 B.n85 B.n84 585
R109 B.n288 B.n85 585
R110 B.n287 B.n286 585
R111 B.n289 B.n287 585
R112 B.n285 B.n90 585
R113 B.n90 B.n89 585
R114 B.n284 B.n283 585
R115 B.n283 B.n282 585
R116 B.n92 B.n91 585
R117 B.n93 B.n92 585
R118 B.n275 B.n274 585
R119 B.n276 B.n275 585
R120 B.n273 B.n98 585
R121 B.n98 B.n97 585
R122 B.n272 B.n271 585
R123 B.n271 B.n270 585
R124 B.n100 B.n99 585
R125 B.n101 B.n100 585
R126 B.n263 B.n262 585
R127 B.n264 B.n263 585
R128 B.n261 B.n106 585
R129 B.n106 B.n105 585
R130 B.n260 B.n259 585
R131 B.n259 B.n258 585
R132 B.n108 B.n107 585
R133 B.n251 B.n108 585
R134 B.n250 B.n249 585
R135 B.n252 B.n250 585
R136 B.n248 B.n113 585
R137 B.n113 B.n112 585
R138 B.n247 B.n246 585
R139 B.n246 B.n245 585
R140 B.n115 B.n114 585
R141 B.n116 B.n115 585
R142 B.n238 B.n237 585
R143 B.n239 B.n238 585
R144 B.n236 B.n121 585
R145 B.n121 B.n120 585
R146 B.n235 B.n234 585
R147 B.n234 B.n233 585
R148 B.n230 B.n125 585
R149 B.n229 B.n228 585
R150 B.n226 B.n126 585
R151 B.n226 B.n124 585
R152 B.n225 B.n224 585
R153 B.n223 B.n222 585
R154 B.n221 B.n128 585
R155 B.n219 B.n218 585
R156 B.n217 B.n129 585
R157 B.n216 B.n215 585
R158 B.n213 B.n130 585
R159 B.n211 B.n210 585
R160 B.n209 B.n131 585
R161 B.n208 B.n207 585
R162 B.n205 B.n132 585
R163 B.n203 B.n202 585
R164 B.n201 B.n133 585
R165 B.n199 B.n198 585
R166 B.n196 B.n136 585
R167 B.n194 B.n193 585
R168 B.n192 B.n137 585
R169 B.n191 B.n190 585
R170 B.n188 B.n138 585
R171 B.n186 B.n185 585
R172 B.n184 B.n139 585
R173 B.n183 B.n182 585
R174 B.n180 B.n179 585
R175 B.n178 B.n177 585
R176 B.n176 B.n144 585
R177 B.n174 B.n173 585
R178 B.n172 B.n145 585
R179 B.n171 B.n170 585
R180 B.n168 B.n146 585
R181 B.n166 B.n165 585
R182 B.n164 B.n147 585
R183 B.n163 B.n162 585
R184 B.n160 B.n148 585
R185 B.n158 B.n157 585
R186 B.n156 B.n149 585
R187 B.n155 B.n154 585
R188 B.n152 B.n150 585
R189 B.n123 B.n122 585
R190 B.n232 B.n231 585
R191 B.n233 B.n232 585
R192 B.n119 B.n118 585
R193 B.n120 B.n119 585
R194 B.n241 B.n240 585
R195 B.n240 B.n239 585
R196 B.n242 B.n117 585
R197 B.n117 B.n116 585
R198 B.n244 B.n243 585
R199 B.n245 B.n244 585
R200 B.n111 B.n110 585
R201 B.n112 B.n111 585
R202 B.n254 B.n253 585
R203 B.n253 B.n252 585
R204 B.n255 B.n109 585
R205 B.n251 B.n109 585
R206 B.n257 B.n256 585
R207 B.n258 B.n257 585
R208 B.n104 B.n103 585
R209 B.n105 B.n104 585
R210 B.n266 B.n265 585
R211 B.n265 B.n264 585
R212 B.n267 B.n102 585
R213 B.n102 B.n101 585
R214 B.n269 B.n268 585
R215 B.n270 B.n269 585
R216 B.n96 B.n95 585
R217 B.n97 B.n96 585
R218 B.n278 B.n277 585
R219 B.n277 B.n276 585
R220 B.n279 B.n94 585
R221 B.n94 B.n93 585
R222 B.n281 B.n280 585
R223 B.n282 B.n281 585
R224 B.n88 B.n87 585
R225 B.n89 B.n88 585
R226 B.n291 B.n290 585
R227 B.n290 B.n289 585
R228 B.n292 B.n86 585
R229 B.n288 B.n86 585
R230 B.n294 B.n293 585
R231 B.n295 B.n294 585
R232 B.n81 B.n80 585
R233 B.n82 B.n81 585
R234 B.n304 B.n303 585
R235 B.n303 B.n302 585
R236 B.n305 B.n79 585
R237 B.n79 B.n78 585
R238 B.n307 B.n306 585
R239 B.n308 B.n307 585
R240 B.n2 B.n0 585
R241 B.n4 B.n2 585
R242 B.n3 B.n1 585
R243 B.n479 B.n3 585
R244 B.n477 B.n476 585
R245 B.n478 B.n477 585
R246 B.n475 B.n9 585
R247 B.n9 B.n8 585
R248 B.n474 B.n473 585
R249 B.n473 B.n472 585
R250 B.n11 B.n10 585
R251 B.n471 B.n11 585
R252 B.n469 B.n468 585
R253 B.n470 B.n469 585
R254 B.n467 B.n15 585
R255 B.n18 B.n15 585
R256 B.n466 B.n465 585
R257 B.n465 B.n464 585
R258 B.n17 B.n16 585
R259 B.n463 B.n17 585
R260 B.n461 B.n460 585
R261 B.n462 B.n461 585
R262 B.n459 B.n23 585
R263 B.n23 B.n22 585
R264 B.n458 B.n457 585
R265 B.n457 B.n456 585
R266 B.n25 B.n24 585
R267 B.n455 B.n25 585
R268 B.n453 B.n452 585
R269 B.n454 B.n453 585
R270 B.n451 B.n30 585
R271 B.n30 B.n29 585
R272 B.n450 B.n449 585
R273 B.n449 B.n448 585
R274 B.n32 B.n31 585
R275 B.n447 B.n32 585
R276 B.n445 B.n444 585
R277 B.n446 B.n445 585
R278 B.n443 B.n36 585
R279 B.n39 B.n36 585
R280 B.n442 B.n441 585
R281 B.n441 B.n440 585
R282 B.n38 B.n37 585
R283 B.n439 B.n38 585
R284 B.n437 B.n436 585
R285 B.n438 B.n437 585
R286 B.n435 B.n44 585
R287 B.n44 B.n43 585
R288 B.n434 B.n433 585
R289 B.n433 B.n432 585
R290 B.n46 B.n45 585
R291 B.n431 B.n46 585
R292 B.n429 B.n428 585
R293 B.n430 B.n429 585
R294 B.n482 B.n481 585
R295 B.n481 B.n480 585
R296 B.n232 B.n125 502.111
R297 B.n429 B.n51 502.111
R298 B.n234 B.n123 502.111
R299 B.n75 B.n49 502.111
R300 B.n348 B.n50 256.663
R301 B.n350 B.n50 256.663
R302 B.n356 B.n50 256.663
R303 B.n358 B.n50 256.663
R304 B.n364 B.n50 256.663
R305 B.n366 B.n50 256.663
R306 B.n372 B.n50 256.663
R307 B.n374 B.n50 256.663
R308 B.n381 B.n50 256.663
R309 B.n383 B.n50 256.663
R310 B.n389 B.n50 256.663
R311 B.n391 B.n50 256.663
R312 B.n398 B.n50 256.663
R313 B.n400 B.n50 256.663
R314 B.n406 B.n50 256.663
R315 B.n408 B.n50 256.663
R316 B.n414 B.n50 256.663
R317 B.n416 B.n50 256.663
R318 B.n422 B.n50 256.663
R319 B.n424 B.n50 256.663
R320 B.n227 B.n124 256.663
R321 B.n127 B.n124 256.663
R322 B.n220 B.n124 256.663
R323 B.n214 B.n124 256.663
R324 B.n212 B.n124 256.663
R325 B.n206 B.n124 256.663
R326 B.n204 B.n124 256.663
R327 B.n197 B.n124 256.663
R328 B.n195 B.n124 256.663
R329 B.n189 B.n124 256.663
R330 B.n187 B.n124 256.663
R331 B.n181 B.n124 256.663
R332 B.n143 B.n124 256.663
R333 B.n175 B.n124 256.663
R334 B.n169 B.n124 256.663
R335 B.n167 B.n124 256.663
R336 B.n161 B.n124 256.663
R337 B.n159 B.n124 256.663
R338 B.n153 B.n124 256.663
R339 B.n151 B.n124 256.663
R340 B.n140 B.t2 236.397
R341 B.n134 B.t13 236.397
R342 B.n60 B.t10 236.397
R343 B.n66 B.t6 236.397
R344 B.n140 B.t5 190.942
R345 B.n66 B.t8 190.942
R346 B.n134 B.t15 190.942
R347 B.n60 B.t11 190.942
R348 B.n233 B.n124 165.228
R349 B.n430 B.n50 165.228
R350 B.n232 B.n119 163.367
R351 B.n240 B.n119 163.367
R352 B.n240 B.n117 163.367
R353 B.n244 B.n117 163.367
R354 B.n244 B.n111 163.367
R355 B.n253 B.n111 163.367
R356 B.n253 B.n109 163.367
R357 B.n257 B.n109 163.367
R358 B.n257 B.n104 163.367
R359 B.n265 B.n104 163.367
R360 B.n265 B.n102 163.367
R361 B.n269 B.n102 163.367
R362 B.n269 B.n96 163.367
R363 B.n277 B.n96 163.367
R364 B.n277 B.n94 163.367
R365 B.n281 B.n94 163.367
R366 B.n281 B.n88 163.367
R367 B.n290 B.n88 163.367
R368 B.n290 B.n86 163.367
R369 B.n294 B.n86 163.367
R370 B.n294 B.n81 163.367
R371 B.n303 B.n81 163.367
R372 B.n303 B.n79 163.367
R373 B.n307 B.n79 163.367
R374 B.n307 B.n2 163.367
R375 B.n481 B.n2 163.367
R376 B.n481 B.n3 163.367
R377 B.n477 B.n3 163.367
R378 B.n477 B.n9 163.367
R379 B.n473 B.n9 163.367
R380 B.n473 B.n11 163.367
R381 B.n469 B.n11 163.367
R382 B.n469 B.n15 163.367
R383 B.n465 B.n15 163.367
R384 B.n465 B.n17 163.367
R385 B.n461 B.n17 163.367
R386 B.n461 B.n23 163.367
R387 B.n457 B.n23 163.367
R388 B.n457 B.n25 163.367
R389 B.n453 B.n25 163.367
R390 B.n453 B.n30 163.367
R391 B.n449 B.n30 163.367
R392 B.n449 B.n32 163.367
R393 B.n445 B.n32 163.367
R394 B.n445 B.n36 163.367
R395 B.n441 B.n36 163.367
R396 B.n441 B.n38 163.367
R397 B.n437 B.n38 163.367
R398 B.n437 B.n44 163.367
R399 B.n433 B.n44 163.367
R400 B.n433 B.n46 163.367
R401 B.n429 B.n46 163.367
R402 B.n228 B.n226 163.367
R403 B.n226 B.n225 163.367
R404 B.n222 B.n221 163.367
R405 B.n219 B.n129 163.367
R406 B.n215 B.n213 163.367
R407 B.n211 B.n131 163.367
R408 B.n207 B.n205 163.367
R409 B.n203 B.n133 163.367
R410 B.n198 B.n196 163.367
R411 B.n194 B.n137 163.367
R412 B.n190 B.n188 163.367
R413 B.n186 B.n139 163.367
R414 B.n182 B.n180 163.367
R415 B.n177 B.n176 163.367
R416 B.n174 B.n145 163.367
R417 B.n170 B.n168 163.367
R418 B.n166 B.n147 163.367
R419 B.n162 B.n160 163.367
R420 B.n158 B.n149 163.367
R421 B.n154 B.n152 163.367
R422 B.n234 B.n121 163.367
R423 B.n238 B.n121 163.367
R424 B.n238 B.n115 163.367
R425 B.n246 B.n115 163.367
R426 B.n246 B.n113 163.367
R427 B.n250 B.n113 163.367
R428 B.n250 B.n108 163.367
R429 B.n259 B.n108 163.367
R430 B.n259 B.n106 163.367
R431 B.n263 B.n106 163.367
R432 B.n263 B.n100 163.367
R433 B.n271 B.n100 163.367
R434 B.n271 B.n98 163.367
R435 B.n275 B.n98 163.367
R436 B.n275 B.n92 163.367
R437 B.n283 B.n92 163.367
R438 B.n283 B.n90 163.367
R439 B.n287 B.n90 163.367
R440 B.n287 B.n85 163.367
R441 B.n296 B.n85 163.367
R442 B.n296 B.n83 163.367
R443 B.n301 B.n83 163.367
R444 B.n301 B.n77 163.367
R445 B.n309 B.n77 163.367
R446 B.n310 B.n309 163.367
R447 B.n310 B.n5 163.367
R448 B.n6 B.n5 163.367
R449 B.n7 B.n6 163.367
R450 B.n315 B.n7 163.367
R451 B.n315 B.n12 163.367
R452 B.n13 B.n12 163.367
R453 B.n14 B.n13 163.367
R454 B.n320 B.n14 163.367
R455 B.n320 B.n19 163.367
R456 B.n20 B.n19 163.367
R457 B.n21 B.n20 163.367
R458 B.n325 B.n21 163.367
R459 B.n325 B.n26 163.367
R460 B.n27 B.n26 163.367
R461 B.n28 B.n27 163.367
R462 B.n330 B.n28 163.367
R463 B.n330 B.n33 163.367
R464 B.n34 B.n33 163.367
R465 B.n35 B.n34 163.367
R466 B.n335 B.n35 163.367
R467 B.n335 B.n40 163.367
R468 B.n41 B.n40 163.367
R469 B.n42 B.n41 163.367
R470 B.n340 B.n42 163.367
R471 B.n340 B.n47 163.367
R472 B.n48 B.n47 163.367
R473 B.n49 B.n48 163.367
R474 B.n425 B.n423 163.367
R475 B.n421 B.n53 163.367
R476 B.n417 B.n415 163.367
R477 B.n413 B.n55 163.367
R478 B.n409 B.n407 163.367
R479 B.n405 B.n57 163.367
R480 B.n401 B.n399 163.367
R481 B.n397 B.n59 163.367
R482 B.n392 B.n390 163.367
R483 B.n388 B.n63 163.367
R484 B.n384 B.n382 163.367
R485 B.n380 B.n65 163.367
R486 B.n375 B.n373 163.367
R487 B.n371 B.n69 163.367
R488 B.n367 B.n365 163.367
R489 B.n363 B.n71 163.367
R490 B.n359 B.n357 163.367
R491 B.n355 B.n73 163.367
R492 B.n351 B.n349 163.367
R493 B.n347 B.n75 163.367
R494 B.n141 B.t4 131.792
R495 B.n67 B.t9 131.792
R496 B.n135 B.t14 131.792
R497 B.n61 B.t12 131.792
R498 B.n233 B.n120 88.4689
R499 B.n239 B.n120 88.4689
R500 B.n239 B.n116 88.4689
R501 B.n245 B.n116 88.4689
R502 B.n245 B.n112 88.4689
R503 B.n252 B.n112 88.4689
R504 B.n252 B.n251 88.4689
R505 B.n258 B.n105 88.4689
R506 B.n264 B.n105 88.4689
R507 B.n264 B.n101 88.4689
R508 B.n270 B.n101 88.4689
R509 B.n270 B.n97 88.4689
R510 B.n276 B.n97 88.4689
R511 B.n276 B.n93 88.4689
R512 B.n282 B.n93 88.4689
R513 B.n282 B.n89 88.4689
R514 B.n289 B.n89 88.4689
R515 B.n289 B.n288 88.4689
R516 B.n295 B.n82 88.4689
R517 B.n302 B.n82 88.4689
R518 B.n302 B.n78 88.4689
R519 B.n308 B.n78 88.4689
R520 B.n308 B.n4 88.4689
R521 B.n480 B.n4 88.4689
R522 B.n480 B.n479 88.4689
R523 B.n479 B.n478 88.4689
R524 B.n478 B.n8 88.4689
R525 B.n472 B.n8 88.4689
R526 B.n472 B.n471 88.4689
R527 B.n471 B.n470 88.4689
R528 B.n464 B.n18 88.4689
R529 B.n464 B.n463 88.4689
R530 B.n463 B.n462 88.4689
R531 B.n462 B.n22 88.4689
R532 B.n456 B.n22 88.4689
R533 B.n456 B.n455 88.4689
R534 B.n455 B.n454 88.4689
R535 B.n454 B.n29 88.4689
R536 B.n448 B.n29 88.4689
R537 B.n448 B.n447 88.4689
R538 B.n447 B.n446 88.4689
R539 B.n440 B.n39 88.4689
R540 B.n440 B.n439 88.4689
R541 B.n439 B.n438 88.4689
R542 B.n438 B.n43 88.4689
R543 B.n432 B.n43 88.4689
R544 B.n432 B.n431 88.4689
R545 B.n431 B.n430 88.4689
R546 B.n288 B.t1 80.6628
R547 B.n18 B.t0 80.6628
R548 B.n227 B.n125 71.676
R549 B.n225 B.n127 71.676
R550 B.n221 B.n220 71.676
R551 B.n214 B.n129 71.676
R552 B.n213 B.n212 71.676
R553 B.n206 B.n131 71.676
R554 B.n205 B.n204 71.676
R555 B.n197 B.n133 71.676
R556 B.n196 B.n195 71.676
R557 B.n189 B.n137 71.676
R558 B.n188 B.n187 71.676
R559 B.n181 B.n139 71.676
R560 B.n180 B.n143 71.676
R561 B.n176 B.n175 71.676
R562 B.n169 B.n145 71.676
R563 B.n168 B.n167 71.676
R564 B.n161 B.n147 71.676
R565 B.n160 B.n159 71.676
R566 B.n153 B.n149 71.676
R567 B.n152 B.n151 71.676
R568 B.n424 B.n51 71.676
R569 B.n423 B.n422 71.676
R570 B.n416 B.n53 71.676
R571 B.n415 B.n414 71.676
R572 B.n408 B.n55 71.676
R573 B.n407 B.n406 71.676
R574 B.n400 B.n57 71.676
R575 B.n399 B.n398 71.676
R576 B.n391 B.n59 71.676
R577 B.n390 B.n389 71.676
R578 B.n383 B.n63 71.676
R579 B.n382 B.n381 71.676
R580 B.n374 B.n65 71.676
R581 B.n373 B.n372 71.676
R582 B.n366 B.n69 71.676
R583 B.n365 B.n364 71.676
R584 B.n358 B.n71 71.676
R585 B.n357 B.n356 71.676
R586 B.n350 B.n73 71.676
R587 B.n349 B.n348 71.676
R588 B.n348 B.n347 71.676
R589 B.n351 B.n350 71.676
R590 B.n356 B.n355 71.676
R591 B.n359 B.n358 71.676
R592 B.n364 B.n363 71.676
R593 B.n367 B.n366 71.676
R594 B.n372 B.n371 71.676
R595 B.n375 B.n374 71.676
R596 B.n381 B.n380 71.676
R597 B.n384 B.n383 71.676
R598 B.n389 B.n388 71.676
R599 B.n392 B.n391 71.676
R600 B.n398 B.n397 71.676
R601 B.n401 B.n400 71.676
R602 B.n406 B.n405 71.676
R603 B.n409 B.n408 71.676
R604 B.n414 B.n413 71.676
R605 B.n417 B.n416 71.676
R606 B.n422 B.n421 71.676
R607 B.n425 B.n424 71.676
R608 B.n228 B.n227 71.676
R609 B.n222 B.n127 71.676
R610 B.n220 B.n219 71.676
R611 B.n215 B.n214 71.676
R612 B.n212 B.n211 71.676
R613 B.n207 B.n206 71.676
R614 B.n204 B.n203 71.676
R615 B.n198 B.n197 71.676
R616 B.n195 B.n194 71.676
R617 B.n190 B.n189 71.676
R618 B.n187 B.n186 71.676
R619 B.n182 B.n181 71.676
R620 B.n177 B.n143 71.676
R621 B.n175 B.n174 71.676
R622 B.n170 B.n169 71.676
R623 B.n167 B.n166 71.676
R624 B.n162 B.n161 71.676
R625 B.n159 B.n158 71.676
R626 B.n154 B.n153 71.676
R627 B.n151 B.n123 71.676
R628 B.n251 B.t3 65.0508
R629 B.n39 B.t7 65.0508
R630 B.n142 B.n141 59.5399
R631 B.n200 B.n135 59.5399
R632 B.n395 B.n61 59.5399
R633 B.n377 B.n67 59.5399
R634 B.n141 B.n140 59.152
R635 B.n135 B.n134 59.152
R636 B.n61 B.n60 59.152
R637 B.n67 B.n66 59.152
R638 B.n428 B.n427 32.6249
R639 B.n345 B.n344 32.6249
R640 B.n235 B.n122 32.6249
R641 B.n231 B.n230 32.6249
R642 B.n258 B.t3 23.4186
R643 B.n446 B.t7 23.4186
R644 B B.n482 18.0485
R645 B.n427 B.n426 10.6151
R646 B.n426 B.n52 10.6151
R647 B.n420 B.n52 10.6151
R648 B.n420 B.n419 10.6151
R649 B.n419 B.n418 10.6151
R650 B.n418 B.n54 10.6151
R651 B.n412 B.n54 10.6151
R652 B.n412 B.n411 10.6151
R653 B.n411 B.n410 10.6151
R654 B.n410 B.n56 10.6151
R655 B.n404 B.n56 10.6151
R656 B.n404 B.n403 10.6151
R657 B.n403 B.n402 10.6151
R658 B.n402 B.n58 10.6151
R659 B.n396 B.n58 10.6151
R660 B.n394 B.n393 10.6151
R661 B.n393 B.n62 10.6151
R662 B.n387 B.n62 10.6151
R663 B.n387 B.n386 10.6151
R664 B.n386 B.n385 10.6151
R665 B.n385 B.n64 10.6151
R666 B.n379 B.n64 10.6151
R667 B.n379 B.n378 10.6151
R668 B.n376 B.n68 10.6151
R669 B.n370 B.n68 10.6151
R670 B.n370 B.n369 10.6151
R671 B.n369 B.n368 10.6151
R672 B.n368 B.n70 10.6151
R673 B.n362 B.n70 10.6151
R674 B.n362 B.n361 10.6151
R675 B.n361 B.n360 10.6151
R676 B.n360 B.n72 10.6151
R677 B.n354 B.n72 10.6151
R678 B.n354 B.n353 10.6151
R679 B.n353 B.n352 10.6151
R680 B.n352 B.n74 10.6151
R681 B.n346 B.n74 10.6151
R682 B.n346 B.n345 10.6151
R683 B.n236 B.n235 10.6151
R684 B.n237 B.n236 10.6151
R685 B.n237 B.n114 10.6151
R686 B.n247 B.n114 10.6151
R687 B.n248 B.n247 10.6151
R688 B.n249 B.n248 10.6151
R689 B.n249 B.n107 10.6151
R690 B.n260 B.n107 10.6151
R691 B.n261 B.n260 10.6151
R692 B.n262 B.n261 10.6151
R693 B.n262 B.n99 10.6151
R694 B.n272 B.n99 10.6151
R695 B.n273 B.n272 10.6151
R696 B.n274 B.n273 10.6151
R697 B.n274 B.n91 10.6151
R698 B.n284 B.n91 10.6151
R699 B.n285 B.n284 10.6151
R700 B.n286 B.n285 10.6151
R701 B.n286 B.n84 10.6151
R702 B.n297 B.n84 10.6151
R703 B.n298 B.n297 10.6151
R704 B.n300 B.n298 10.6151
R705 B.n300 B.n299 10.6151
R706 B.n299 B.n76 10.6151
R707 B.n311 B.n76 10.6151
R708 B.n312 B.n311 10.6151
R709 B.n313 B.n312 10.6151
R710 B.n314 B.n313 10.6151
R711 B.n316 B.n314 10.6151
R712 B.n317 B.n316 10.6151
R713 B.n318 B.n317 10.6151
R714 B.n319 B.n318 10.6151
R715 B.n321 B.n319 10.6151
R716 B.n322 B.n321 10.6151
R717 B.n323 B.n322 10.6151
R718 B.n324 B.n323 10.6151
R719 B.n326 B.n324 10.6151
R720 B.n327 B.n326 10.6151
R721 B.n328 B.n327 10.6151
R722 B.n329 B.n328 10.6151
R723 B.n331 B.n329 10.6151
R724 B.n332 B.n331 10.6151
R725 B.n333 B.n332 10.6151
R726 B.n334 B.n333 10.6151
R727 B.n336 B.n334 10.6151
R728 B.n337 B.n336 10.6151
R729 B.n338 B.n337 10.6151
R730 B.n339 B.n338 10.6151
R731 B.n341 B.n339 10.6151
R732 B.n342 B.n341 10.6151
R733 B.n343 B.n342 10.6151
R734 B.n344 B.n343 10.6151
R735 B.n230 B.n229 10.6151
R736 B.n229 B.n126 10.6151
R737 B.n224 B.n126 10.6151
R738 B.n224 B.n223 10.6151
R739 B.n223 B.n128 10.6151
R740 B.n218 B.n128 10.6151
R741 B.n218 B.n217 10.6151
R742 B.n217 B.n216 10.6151
R743 B.n216 B.n130 10.6151
R744 B.n210 B.n130 10.6151
R745 B.n210 B.n209 10.6151
R746 B.n209 B.n208 10.6151
R747 B.n208 B.n132 10.6151
R748 B.n202 B.n132 10.6151
R749 B.n202 B.n201 10.6151
R750 B.n199 B.n136 10.6151
R751 B.n193 B.n136 10.6151
R752 B.n193 B.n192 10.6151
R753 B.n192 B.n191 10.6151
R754 B.n191 B.n138 10.6151
R755 B.n185 B.n138 10.6151
R756 B.n185 B.n184 10.6151
R757 B.n184 B.n183 10.6151
R758 B.n179 B.n178 10.6151
R759 B.n178 B.n144 10.6151
R760 B.n173 B.n144 10.6151
R761 B.n173 B.n172 10.6151
R762 B.n172 B.n171 10.6151
R763 B.n171 B.n146 10.6151
R764 B.n165 B.n146 10.6151
R765 B.n165 B.n164 10.6151
R766 B.n164 B.n163 10.6151
R767 B.n163 B.n148 10.6151
R768 B.n157 B.n148 10.6151
R769 B.n157 B.n156 10.6151
R770 B.n156 B.n155 10.6151
R771 B.n155 B.n150 10.6151
R772 B.n150 B.n122 10.6151
R773 B.n231 B.n118 10.6151
R774 B.n241 B.n118 10.6151
R775 B.n242 B.n241 10.6151
R776 B.n243 B.n242 10.6151
R777 B.n243 B.n110 10.6151
R778 B.n254 B.n110 10.6151
R779 B.n255 B.n254 10.6151
R780 B.n256 B.n255 10.6151
R781 B.n256 B.n103 10.6151
R782 B.n266 B.n103 10.6151
R783 B.n267 B.n266 10.6151
R784 B.n268 B.n267 10.6151
R785 B.n268 B.n95 10.6151
R786 B.n278 B.n95 10.6151
R787 B.n279 B.n278 10.6151
R788 B.n280 B.n279 10.6151
R789 B.n280 B.n87 10.6151
R790 B.n291 B.n87 10.6151
R791 B.n292 B.n291 10.6151
R792 B.n293 B.n292 10.6151
R793 B.n293 B.n80 10.6151
R794 B.n304 B.n80 10.6151
R795 B.n305 B.n304 10.6151
R796 B.n306 B.n305 10.6151
R797 B.n306 B.n0 10.6151
R798 B.n476 B.n1 10.6151
R799 B.n476 B.n475 10.6151
R800 B.n475 B.n474 10.6151
R801 B.n474 B.n10 10.6151
R802 B.n468 B.n10 10.6151
R803 B.n468 B.n467 10.6151
R804 B.n467 B.n466 10.6151
R805 B.n466 B.n16 10.6151
R806 B.n460 B.n16 10.6151
R807 B.n460 B.n459 10.6151
R808 B.n459 B.n458 10.6151
R809 B.n458 B.n24 10.6151
R810 B.n452 B.n24 10.6151
R811 B.n452 B.n451 10.6151
R812 B.n451 B.n450 10.6151
R813 B.n450 B.n31 10.6151
R814 B.n444 B.n31 10.6151
R815 B.n444 B.n443 10.6151
R816 B.n443 B.n442 10.6151
R817 B.n442 B.n37 10.6151
R818 B.n436 B.n37 10.6151
R819 B.n436 B.n435 10.6151
R820 B.n435 B.n434 10.6151
R821 B.n434 B.n45 10.6151
R822 B.n428 B.n45 10.6151
R823 B.n295 B.t1 7.80653
R824 B.n470 B.t0 7.80653
R825 B.n395 B.n394 6.5566
R826 B.n378 B.n377 6.5566
R827 B.n200 B.n199 6.5566
R828 B.n183 B.n142 6.5566
R829 B.n396 B.n395 4.05904
R830 B.n377 B.n376 4.05904
R831 B.n201 B.n200 4.05904
R832 B.n179 B.n142 4.05904
R833 B.n482 B.n0 2.81026
R834 B.n482 B.n1 2.81026
R835 VN VN.t1 107.609
R836 VN VN.t0 69.7453
R837 VTAIL.n58 VTAIL.n48 289.615
R838 VTAIL.n10 VTAIL.n0 289.615
R839 VTAIL.n42 VTAIL.n32 289.615
R840 VTAIL.n26 VTAIL.n16 289.615
R841 VTAIL.n52 VTAIL.n51 185
R842 VTAIL.n57 VTAIL.n56 185
R843 VTAIL.n59 VTAIL.n58 185
R844 VTAIL.n4 VTAIL.n3 185
R845 VTAIL.n9 VTAIL.n8 185
R846 VTAIL.n11 VTAIL.n10 185
R847 VTAIL.n43 VTAIL.n42 185
R848 VTAIL.n41 VTAIL.n40 185
R849 VTAIL.n36 VTAIL.n35 185
R850 VTAIL.n27 VTAIL.n26 185
R851 VTAIL.n25 VTAIL.n24 185
R852 VTAIL.n20 VTAIL.n19 185
R853 VTAIL.n53 VTAIL.t2 148.606
R854 VTAIL.n5 VTAIL.t0 148.606
R855 VTAIL.n37 VTAIL.t1 148.606
R856 VTAIL.n21 VTAIL.t3 148.606
R857 VTAIL.n57 VTAIL.n51 104.615
R858 VTAIL.n58 VTAIL.n57 104.615
R859 VTAIL.n9 VTAIL.n3 104.615
R860 VTAIL.n10 VTAIL.n9 104.615
R861 VTAIL.n42 VTAIL.n41 104.615
R862 VTAIL.n41 VTAIL.n35 104.615
R863 VTAIL.n26 VTAIL.n25 104.615
R864 VTAIL.n25 VTAIL.n19 104.615
R865 VTAIL.t2 VTAIL.n51 52.3082
R866 VTAIL.t0 VTAIL.n3 52.3082
R867 VTAIL.t1 VTAIL.n35 52.3082
R868 VTAIL.t3 VTAIL.n19 52.3082
R869 VTAIL.n63 VTAIL.n62 33.349
R870 VTAIL.n15 VTAIL.n14 33.349
R871 VTAIL.n47 VTAIL.n46 33.349
R872 VTAIL.n31 VTAIL.n30 33.349
R873 VTAIL.n31 VTAIL.n15 20.3669
R874 VTAIL.n63 VTAIL.n47 17.7376
R875 VTAIL.n53 VTAIL.n52 15.5966
R876 VTAIL.n5 VTAIL.n4 15.5966
R877 VTAIL.n37 VTAIL.n36 15.5966
R878 VTAIL.n21 VTAIL.n20 15.5966
R879 VTAIL.n56 VTAIL.n55 12.8005
R880 VTAIL.n8 VTAIL.n7 12.8005
R881 VTAIL.n40 VTAIL.n39 12.8005
R882 VTAIL.n24 VTAIL.n23 12.8005
R883 VTAIL.n59 VTAIL.n50 12.0247
R884 VTAIL.n11 VTAIL.n2 12.0247
R885 VTAIL.n43 VTAIL.n34 12.0247
R886 VTAIL.n27 VTAIL.n18 12.0247
R887 VTAIL.n60 VTAIL.n48 11.249
R888 VTAIL.n12 VTAIL.n0 11.249
R889 VTAIL.n44 VTAIL.n32 11.249
R890 VTAIL.n28 VTAIL.n16 11.249
R891 VTAIL.n62 VTAIL.n61 9.45567
R892 VTAIL.n14 VTAIL.n13 9.45567
R893 VTAIL.n46 VTAIL.n45 9.45567
R894 VTAIL.n30 VTAIL.n29 9.45567
R895 VTAIL.n61 VTAIL.n60 9.3005
R896 VTAIL.n50 VTAIL.n49 9.3005
R897 VTAIL.n55 VTAIL.n54 9.3005
R898 VTAIL.n13 VTAIL.n12 9.3005
R899 VTAIL.n2 VTAIL.n1 9.3005
R900 VTAIL.n7 VTAIL.n6 9.3005
R901 VTAIL.n45 VTAIL.n44 9.3005
R902 VTAIL.n34 VTAIL.n33 9.3005
R903 VTAIL.n39 VTAIL.n38 9.3005
R904 VTAIL.n29 VTAIL.n28 9.3005
R905 VTAIL.n18 VTAIL.n17 9.3005
R906 VTAIL.n23 VTAIL.n22 9.3005
R907 VTAIL.n54 VTAIL.n53 4.46457
R908 VTAIL.n6 VTAIL.n5 4.46457
R909 VTAIL.n38 VTAIL.n37 4.46457
R910 VTAIL.n22 VTAIL.n21 4.46457
R911 VTAIL.n62 VTAIL.n48 2.71565
R912 VTAIL.n14 VTAIL.n0 2.71565
R913 VTAIL.n46 VTAIL.n32 2.71565
R914 VTAIL.n30 VTAIL.n16 2.71565
R915 VTAIL.n60 VTAIL.n59 1.93989
R916 VTAIL.n12 VTAIL.n11 1.93989
R917 VTAIL.n44 VTAIL.n43 1.93989
R918 VTAIL.n28 VTAIL.n27 1.93989
R919 VTAIL.n47 VTAIL.n31 1.78498
R920 VTAIL VTAIL.n15 1.18584
R921 VTAIL.n56 VTAIL.n50 1.16414
R922 VTAIL.n8 VTAIL.n2 1.16414
R923 VTAIL.n40 VTAIL.n34 1.16414
R924 VTAIL.n24 VTAIL.n18 1.16414
R925 VTAIL VTAIL.n63 0.599638
R926 VTAIL.n55 VTAIL.n52 0.388379
R927 VTAIL.n7 VTAIL.n4 0.388379
R928 VTAIL.n39 VTAIL.n36 0.388379
R929 VTAIL.n23 VTAIL.n20 0.388379
R930 VTAIL.n54 VTAIL.n49 0.155672
R931 VTAIL.n61 VTAIL.n49 0.155672
R932 VTAIL.n6 VTAIL.n1 0.155672
R933 VTAIL.n13 VTAIL.n1 0.155672
R934 VTAIL.n45 VTAIL.n33 0.155672
R935 VTAIL.n38 VTAIL.n33 0.155672
R936 VTAIL.n29 VTAIL.n17 0.155672
R937 VTAIL.n22 VTAIL.n17 0.155672
R938 VDD2.n25 VDD2.n15 289.615
R939 VDD2.n10 VDD2.n0 289.615
R940 VDD2.n26 VDD2.n25 185
R941 VDD2.n24 VDD2.n23 185
R942 VDD2.n19 VDD2.n18 185
R943 VDD2.n4 VDD2.n3 185
R944 VDD2.n9 VDD2.n8 185
R945 VDD2.n11 VDD2.n10 185
R946 VDD2.n20 VDD2.t0 148.606
R947 VDD2.n5 VDD2.t1 148.606
R948 VDD2.n25 VDD2.n24 104.615
R949 VDD2.n24 VDD2.n18 104.615
R950 VDD2.n9 VDD2.n3 104.615
R951 VDD2.n10 VDD2.n9 104.615
R952 VDD2.n30 VDD2.n14 81.6872
R953 VDD2.t0 VDD2.n18 52.3082
R954 VDD2.t1 VDD2.n3 52.3082
R955 VDD2.n30 VDD2.n29 50.0278
R956 VDD2.n20 VDD2.n19 15.5966
R957 VDD2.n5 VDD2.n4 15.5966
R958 VDD2.n23 VDD2.n22 12.8005
R959 VDD2.n8 VDD2.n7 12.8005
R960 VDD2.n26 VDD2.n17 12.0247
R961 VDD2.n11 VDD2.n2 12.0247
R962 VDD2.n27 VDD2.n15 11.249
R963 VDD2.n12 VDD2.n0 11.249
R964 VDD2.n29 VDD2.n28 9.45567
R965 VDD2.n14 VDD2.n13 9.45567
R966 VDD2.n28 VDD2.n27 9.3005
R967 VDD2.n17 VDD2.n16 9.3005
R968 VDD2.n22 VDD2.n21 9.3005
R969 VDD2.n13 VDD2.n12 9.3005
R970 VDD2.n2 VDD2.n1 9.3005
R971 VDD2.n7 VDD2.n6 9.3005
R972 VDD2.n21 VDD2.n20 4.46457
R973 VDD2.n6 VDD2.n5 4.46457
R974 VDD2.n29 VDD2.n15 2.71565
R975 VDD2.n14 VDD2.n0 2.71565
R976 VDD2.n27 VDD2.n26 1.93989
R977 VDD2.n12 VDD2.n11 1.93989
R978 VDD2.n23 VDD2.n17 1.16414
R979 VDD2.n8 VDD2.n2 1.16414
R980 VDD2 VDD2.n30 0.716017
R981 VDD2.n22 VDD2.n19 0.388379
R982 VDD2.n7 VDD2.n4 0.388379
R983 VDD2.n28 VDD2.n16 0.155672
R984 VDD2.n21 VDD2.n16 0.155672
R985 VDD2.n6 VDD2.n1 0.155672
R986 VDD2.n13 VDD2.n1 0.155672
R987 VP.n0 VP.t1 107.608
R988 VP.n0 VP.t0 69.314
R989 VP VP.n0 0.431812
R990 VDD1.n10 VDD1.n0 289.615
R991 VDD1.n25 VDD1.n15 289.615
R992 VDD1.n11 VDD1.n10 185
R993 VDD1.n9 VDD1.n8 185
R994 VDD1.n4 VDD1.n3 185
R995 VDD1.n19 VDD1.n18 185
R996 VDD1.n24 VDD1.n23 185
R997 VDD1.n26 VDD1.n25 185
R998 VDD1.n5 VDD1.t0 148.606
R999 VDD1.n20 VDD1.t1 148.606
R1000 VDD1.n10 VDD1.n9 104.615
R1001 VDD1.n9 VDD1.n3 104.615
R1002 VDD1.n24 VDD1.n18 104.615
R1003 VDD1.n25 VDD1.n24 104.615
R1004 VDD1 VDD1.n29 82.8694
R1005 VDD1.t0 VDD1.n3 52.3082
R1006 VDD1.t1 VDD1.n18 52.3082
R1007 VDD1 VDD1.n14 50.7433
R1008 VDD1.n5 VDD1.n4 15.5966
R1009 VDD1.n20 VDD1.n19 15.5966
R1010 VDD1.n8 VDD1.n7 12.8005
R1011 VDD1.n23 VDD1.n22 12.8005
R1012 VDD1.n11 VDD1.n2 12.0247
R1013 VDD1.n26 VDD1.n17 12.0247
R1014 VDD1.n12 VDD1.n0 11.249
R1015 VDD1.n27 VDD1.n15 11.249
R1016 VDD1.n14 VDD1.n13 9.45567
R1017 VDD1.n29 VDD1.n28 9.45567
R1018 VDD1.n13 VDD1.n12 9.3005
R1019 VDD1.n2 VDD1.n1 9.3005
R1020 VDD1.n7 VDD1.n6 9.3005
R1021 VDD1.n28 VDD1.n27 9.3005
R1022 VDD1.n17 VDD1.n16 9.3005
R1023 VDD1.n22 VDD1.n21 9.3005
R1024 VDD1.n6 VDD1.n5 4.46457
R1025 VDD1.n21 VDD1.n20 4.46457
R1026 VDD1.n14 VDD1.n0 2.71565
R1027 VDD1.n29 VDD1.n15 2.71565
R1028 VDD1.n12 VDD1.n11 1.93989
R1029 VDD1.n27 VDD1.n26 1.93989
R1030 VDD1.n8 VDD1.n2 1.16414
R1031 VDD1.n23 VDD1.n17 1.16414
R1032 VDD1.n7 VDD1.n4 0.388379
R1033 VDD1.n22 VDD1.n19 0.388379
R1034 VDD1.n13 VDD1.n1 0.155672
R1035 VDD1.n6 VDD1.n1 0.155672
R1036 VDD1.n21 VDD1.n16 0.155672
R1037 VDD1.n28 VDD1.n16 0.155672
C0 VN VP 3.8846f
C1 VN VTAIL 1.13738f
C2 VN VDD1 0.153427f
C3 VP VDD2 0.343176f
C4 VDD2 VTAIL 2.82544f
C5 VDD1 VDD2 0.688113f
C6 VN VDD2 0.929697f
C7 VP VTAIL 1.15153f
C8 VP VDD1 1.11792f
C9 VDD1 VTAIL 2.77193f
C10 VDD2 B 2.848755f
C11 VDD1 B 4.45471f
C12 VTAIL B 3.553789f
C13 VN B 7.80048f
C14 VP B 5.779329f
C15 VDD1.n0 B 0.021365f
C16 VDD1.n1 B 0.015966f
C17 VDD1.n2 B 0.00858f
C18 VDD1.n3 B 0.015209f
C19 VDD1.n4 B 0.011825f
C20 VDD1.t0 B 0.034104f
C21 VDD1.n5 B 0.058789f
C22 VDD1.n6 B 0.170744f
C23 VDD1.n7 B 0.00858f
C24 VDD1.n8 B 0.009084f
C25 VDD1.n9 B 0.020279f
C26 VDD1.n10 B 0.041995f
C27 VDD1.n11 B 0.009084f
C28 VDD1.n12 B 0.00858f
C29 VDD1.n13 B 0.038214f
C30 VDD1.n14 B 0.035319f
C31 VDD1.n15 B 0.021365f
C32 VDD1.n16 B 0.015966f
C33 VDD1.n17 B 0.00858f
C34 VDD1.n18 B 0.015209f
C35 VDD1.n19 B 0.011825f
C36 VDD1.t1 B 0.034104f
C37 VDD1.n20 B 0.058789f
C38 VDD1.n21 B 0.170744f
C39 VDD1.n22 B 0.00858f
C40 VDD1.n23 B 0.009084f
C41 VDD1.n24 B 0.020279f
C42 VDD1.n25 B 0.041995f
C43 VDD1.n26 B 0.009084f
C44 VDD1.n27 B 0.00858f
C45 VDD1.n28 B 0.038214f
C46 VDD1.n29 B 0.313565f
C47 VP.t0 B 0.773691f
C48 VP.t1 B 1.18813f
C49 VP.n0 B 1.87143f
C50 VDD2.n0 B 0.021824f
C51 VDD2.n1 B 0.01631f
C52 VDD2.n2 B 0.008764f
C53 VDD2.n3 B 0.015536f
C54 VDD2.n4 B 0.012079f
C55 VDD2.t1 B 0.034838f
C56 VDD2.n5 B 0.060054f
C57 VDD2.n6 B 0.174417f
C58 VDD2.n7 B 0.008764f
C59 VDD2.n8 B 0.00928f
C60 VDD2.n9 B 0.020715f
C61 VDD2.n10 B 0.042899f
C62 VDD2.n11 B 0.00928f
C63 VDD2.n12 B 0.008764f
C64 VDD2.n13 B 0.039036f
C65 VDD2.n14 B 0.293659f
C66 VDD2.n15 B 0.021824f
C67 VDD2.n16 B 0.01631f
C68 VDD2.n17 B 0.008764f
C69 VDD2.n18 B 0.015536f
C70 VDD2.n19 B 0.012079f
C71 VDD2.t0 B 0.034838f
C72 VDD2.n20 B 0.060054f
C73 VDD2.n21 B 0.174417f
C74 VDD2.n22 B 0.008764f
C75 VDD2.n23 B 0.00928f
C76 VDD2.n24 B 0.020715f
C77 VDD2.n25 B 0.042899f
C78 VDD2.n26 B 0.00928f
C79 VDD2.n27 B 0.008764f
C80 VDD2.n28 B 0.039036f
C81 VDD2.n29 B 0.035095f
C82 VDD2.n30 B 1.39898f
C83 VTAIL.n0 B 0.025724f
C84 VTAIL.n1 B 0.019224f
C85 VTAIL.n2 B 0.01033f
C86 VTAIL.n3 B 0.018313f
C87 VTAIL.n4 B 0.014238f
C88 VTAIL.t0 B 0.041063f
C89 VTAIL.n5 B 0.070785f
C90 VTAIL.n6 B 0.205585f
C91 VTAIL.n7 B 0.01033f
C92 VTAIL.n8 B 0.010938f
C93 VTAIL.n9 B 0.024417f
C94 VTAIL.n10 B 0.050565f
C95 VTAIL.n11 B 0.010938f
C96 VTAIL.n12 B 0.01033f
C97 VTAIL.n13 B 0.046011f
C98 VTAIL.n14 B 0.028105f
C99 VTAIL.n15 B 0.847426f
C100 VTAIL.n16 B 0.025724f
C101 VTAIL.n17 B 0.019224f
C102 VTAIL.n18 B 0.01033f
C103 VTAIL.n19 B 0.018313f
C104 VTAIL.n20 B 0.014238f
C105 VTAIL.t3 B 0.041063f
C106 VTAIL.n21 B 0.070785f
C107 VTAIL.n22 B 0.205585f
C108 VTAIL.n23 B 0.01033f
C109 VTAIL.n24 B 0.010938f
C110 VTAIL.n25 B 0.024417f
C111 VTAIL.n26 B 0.050565f
C112 VTAIL.n27 B 0.010938f
C113 VTAIL.n28 B 0.01033f
C114 VTAIL.n29 B 0.046011f
C115 VTAIL.n30 B 0.028105f
C116 VTAIL.n31 B 0.884539f
C117 VTAIL.n32 B 0.025724f
C118 VTAIL.n33 B 0.019224f
C119 VTAIL.n34 B 0.01033f
C120 VTAIL.n35 B 0.018313f
C121 VTAIL.n36 B 0.014238f
C122 VTAIL.t1 B 0.041063f
C123 VTAIL.n37 B 0.070785f
C124 VTAIL.n38 B 0.205585f
C125 VTAIL.n39 B 0.01033f
C126 VTAIL.n40 B 0.010938f
C127 VTAIL.n41 B 0.024417f
C128 VTAIL.n42 B 0.050565f
C129 VTAIL.n43 B 0.010938f
C130 VTAIL.n44 B 0.01033f
C131 VTAIL.n45 B 0.046011f
C132 VTAIL.n46 B 0.028105f
C133 VTAIL.n47 B 0.721668f
C134 VTAIL.n48 B 0.025724f
C135 VTAIL.n49 B 0.019224f
C136 VTAIL.n50 B 0.01033f
C137 VTAIL.n51 B 0.018313f
C138 VTAIL.n52 B 0.014238f
C139 VTAIL.t2 B 0.041063f
C140 VTAIL.n53 B 0.070785f
C141 VTAIL.n54 B 0.205585f
C142 VTAIL.n55 B 0.01033f
C143 VTAIL.n56 B 0.010938f
C144 VTAIL.n57 B 0.024417f
C145 VTAIL.n58 B 0.050565f
C146 VTAIL.n59 B 0.010938f
C147 VTAIL.n60 B 0.01033f
C148 VTAIL.n61 B 0.046011f
C149 VTAIL.n62 B 0.028105f
C150 VTAIL.n63 B 0.648243f
C151 VN.t0 B 0.768545f
C152 VN.t1 B 1.18013f
.ends

