* NGSPICE file created from diff_pair_sample_0495.ext - technology: sky130A

.subckt diff_pair_sample_0495 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t1 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
X1 VTAIL.t9 VP.t0 VDD1.t9 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
X2 VTAIL.t6 VP.t1 VDD1.t8 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
X3 VDD1.t7 VP.t2 VTAIL.t8 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=5.655 ps=29.78 w=14.5 l=1.81
X4 VDD1.t6 VP.t3 VTAIL.t3 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=5.655 ps=29.78 w=14.5 l=1.81
X5 VTAIL.t18 VN.t1 VDD2.t9 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
X6 B.t11 B.t9 B.t10 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=5.655 pd=29.78 as=0 ps=0 w=14.5 l=1.81
X7 B.t8 B.t6 B.t7 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=5.655 pd=29.78 as=0 ps=0 w=14.5 l=1.81
X8 B.t5 B.t3 B.t4 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=5.655 pd=29.78 as=0 ps=0 w=14.5 l=1.81
X9 VDD2.t3 VN.t2 VTAIL.t17 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=5.655 ps=29.78 w=14.5 l=1.81
X10 VDD1.t5 VP.t4 VTAIL.t7 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
X11 VDD2.t4 VN.t3 VTAIL.t16 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=5.655 pd=29.78 as=2.3925 ps=14.83 w=14.5 l=1.81
X12 VTAIL.t2 VP.t5 VDD1.t4 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
X13 VDD1.t3 VP.t6 VTAIL.t5 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=5.655 pd=29.78 as=2.3925 ps=14.83 w=14.5 l=1.81
X14 VDD2.t8 VN.t4 VTAIL.t15 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=5.655 pd=29.78 as=2.3925 ps=14.83 w=14.5 l=1.81
X15 VDD1.t2 VP.t7 VTAIL.t0 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=5.655 pd=29.78 as=2.3925 ps=14.83 w=14.5 l=1.81
X16 VTAIL.t4 VP.t8 VDD1.t1 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
X17 VDD2.t5 VN.t5 VTAIL.t14 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
X18 B.t2 B.t0 B.t1 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=5.655 pd=29.78 as=0 ps=0 w=14.5 l=1.81
X19 VDD1.t0 VP.t9 VTAIL.t1 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
X20 VDD2.t0 VN.t6 VTAIL.t13 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
X21 VTAIL.t12 VN.t7 VDD2.t6 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
X22 VDD2.t2 VN.t8 VTAIL.t11 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=5.655 ps=29.78 w=14.5 l=1.81
X23 VTAIL.t10 VN.t9 VDD2.t7 w_n3538_n3868# sky130_fd_pr__pfet_01v8 ad=2.3925 pd=14.83 as=2.3925 ps=14.83 w=14.5 l=1.81
R0 VN.n7 VN.t3 226.022
R1 VN.n39 VN.t2 226.022
R2 VN.n8 VN.t9 193.066
R3 VN.n15 VN.t5 193.066
R4 VN.n22 VN.t1 193.066
R5 VN.n30 VN.t8 193.066
R6 VN.n40 VN.t0 193.066
R7 VN.n47 VN.t6 193.066
R8 VN.n54 VN.t7 193.066
R9 VN.n62 VN.t4 193.066
R10 VN.n31 VN.n30 184.417
R11 VN.n63 VN.n62 184.417
R12 VN.n61 VN.n32 161.3
R13 VN.n60 VN.n59 161.3
R14 VN.n58 VN.n33 161.3
R15 VN.n57 VN.n56 161.3
R16 VN.n55 VN.n34 161.3
R17 VN.n53 VN.n52 161.3
R18 VN.n51 VN.n35 161.3
R19 VN.n50 VN.n49 161.3
R20 VN.n48 VN.n36 161.3
R21 VN.n46 VN.n45 161.3
R22 VN.n44 VN.n37 161.3
R23 VN.n43 VN.n42 161.3
R24 VN.n41 VN.n38 161.3
R25 VN.n29 VN.n0 161.3
R26 VN.n28 VN.n27 161.3
R27 VN.n26 VN.n1 161.3
R28 VN.n25 VN.n24 161.3
R29 VN.n23 VN.n2 161.3
R30 VN.n21 VN.n20 161.3
R31 VN.n19 VN.n3 161.3
R32 VN.n18 VN.n17 161.3
R33 VN.n16 VN.n4 161.3
R34 VN.n14 VN.n13 161.3
R35 VN.n12 VN.n5 161.3
R36 VN.n11 VN.n10 161.3
R37 VN.n9 VN.n6 161.3
R38 VN.n10 VN.n5 56.5617
R39 VN.n17 VN.n3 56.5617
R40 VN.n42 VN.n37 56.5617
R41 VN.n49 VN.n35 56.5617
R42 VN VN.n63 50.9645
R43 VN.n8 VN.n7 50.6216
R44 VN.n40 VN.n39 50.6216
R45 VN.n24 VN.n1 44.4521
R46 VN.n56 VN.n33 44.4521
R47 VN.n28 VN.n1 36.702
R48 VN.n60 VN.n33 36.702
R49 VN.n10 VN.n9 24.5923
R50 VN.n14 VN.n5 24.5923
R51 VN.n17 VN.n16 24.5923
R52 VN.n21 VN.n3 24.5923
R53 VN.n24 VN.n23 24.5923
R54 VN.n29 VN.n28 24.5923
R55 VN.n42 VN.n41 24.5923
R56 VN.n49 VN.n48 24.5923
R57 VN.n46 VN.n37 24.5923
R58 VN.n56 VN.n55 24.5923
R59 VN.n53 VN.n35 24.5923
R60 VN.n61 VN.n60 24.5923
R61 VN.n9 VN.n8 19.1821
R62 VN.n22 VN.n21 19.1821
R63 VN.n41 VN.n40 19.1821
R64 VN.n54 VN.n53 19.1821
R65 VN.n39 VN.n38 12.4384
R66 VN.n7 VN.n6 12.4384
R67 VN.n15 VN.n14 12.2964
R68 VN.n16 VN.n15 12.2964
R69 VN.n48 VN.n47 12.2964
R70 VN.n47 VN.n46 12.2964
R71 VN.n23 VN.n22 5.4107
R72 VN.n55 VN.n54 5.4107
R73 VN.n30 VN.n29 1.47601
R74 VN.n62 VN.n61 1.47601
R75 VN.n63 VN.n32 0.189894
R76 VN.n59 VN.n32 0.189894
R77 VN.n59 VN.n58 0.189894
R78 VN.n58 VN.n57 0.189894
R79 VN.n57 VN.n34 0.189894
R80 VN.n52 VN.n34 0.189894
R81 VN.n52 VN.n51 0.189894
R82 VN.n51 VN.n50 0.189894
R83 VN.n50 VN.n36 0.189894
R84 VN.n45 VN.n36 0.189894
R85 VN.n45 VN.n44 0.189894
R86 VN.n44 VN.n43 0.189894
R87 VN.n43 VN.n38 0.189894
R88 VN.n11 VN.n6 0.189894
R89 VN.n12 VN.n11 0.189894
R90 VN.n13 VN.n12 0.189894
R91 VN.n13 VN.n4 0.189894
R92 VN.n18 VN.n4 0.189894
R93 VN.n19 VN.n18 0.189894
R94 VN.n20 VN.n19 0.189894
R95 VN.n20 VN.n2 0.189894
R96 VN.n25 VN.n2 0.189894
R97 VN.n26 VN.n25 0.189894
R98 VN.n27 VN.n26 0.189894
R99 VN.n27 VN.n0 0.189894
R100 VN.n31 VN.n0 0.189894
R101 VN VN.n31 0.0516364
R102 VDD2.n1 VDD2.t4 79.3956
R103 VDD2.n4 VDD2.t8 77.5509
R104 VDD2.n3 VDD2.n2 76.6373
R105 VDD2 VDD2.n7 76.6345
R106 VDD2.n6 VDD2.n5 75.3093
R107 VDD2.n1 VDD2.n0 75.309
R108 VDD2.n4 VDD2.n3 44.9782
R109 VDD2.n7 VDD2.t1 2.24222
R110 VDD2.n7 VDD2.t3 2.24222
R111 VDD2.n5 VDD2.t6 2.24222
R112 VDD2.n5 VDD2.t0 2.24222
R113 VDD2.n2 VDD2.t9 2.24222
R114 VDD2.n2 VDD2.t2 2.24222
R115 VDD2.n0 VDD2.t7 2.24222
R116 VDD2.n0 VDD2.t5 2.24222
R117 VDD2.n6 VDD2.n4 1.84533
R118 VDD2 VDD2.n6 0.519897
R119 VDD2.n3 VDD2.n1 0.406361
R120 VTAIL.n11 VTAIL.t17 60.8721
R121 VTAIL.n17 VTAIL.t11 60.872
R122 VTAIL.n2 VTAIL.t8 60.872
R123 VTAIL.n16 VTAIL.t3 60.872
R124 VTAIL.n15 VTAIL.n14 58.6305
R125 VTAIL.n13 VTAIL.n12 58.6305
R126 VTAIL.n10 VTAIL.n9 58.6305
R127 VTAIL.n8 VTAIL.n7 58.6305
R128 VTAIL.n19 VTAIL.n18 58.6302
R129 VTAIL.n1 VTAIL.n0 58.6302
R130 VTAIL.n4 VTAIL.n3 58.6302
R131 VTAIL.n6 VTAIL.n5 58.6302
R132 VTAIL.n8 VTAIL.n6 28.5565
R133 VTAIL.n17 VTAIL.n16 26.7117
R134 VTAIL.n18 VTAIL.t14 2.24222
R135 VTAIL.n18 VTAIL.t18 2.24222
R136 VTAIL.n0 VTAIL.t16 2.24222
R137 VTAIL.n0 VTAIL.t10 2.24222
R138 VTAIL.n3 VTAIL.t7 2.24222
R139 VTAIL.n3 VTAIL.t4 2.24222
R140 VTAIL.n5 VTAIL.t0 2.24222
R141 VTAIL.n5 VTAIL.t9 2.24222
R142 VTAIL.n14 VTAIL.t1 2.24222
R143 VTAIL.n14 VTAIL.t2 2.24222
R144 VTAIL.n12 VTAIL.t5 2.24222
R145 VTAIL.n12 VTAIL.t6 2.24222
R146 VTAIL.n9 VTAIL.t13 2.24222
R147 VTAIL.n9 VTAIL.t19 2.24222
R148 VTAIL.n7 VTAIL.t15 2.24222
R149 VTAIL.n7 VTAIL.t12 2.24222
R150 VTAIL.n10 VTAIL.n8 1.84533
R151 VTAIL.n11 VTAIL.n10 1.84533
R152 VTAIL.n15 VTAIL.n13 1.84533
R153 VTAIL.n16 VTAIL.n15 1.84533
R154 VTAIL.n6 VTAIL.n4 1.84533
R155 VTAIL.n4 VTAIL.n2 1.84533
R156 VTAIL.n19 VTAIL.n17 1.84533
R157 VTAIL VTAIL.n1 1.44231
R158 VTAIL.n13 VTAIL.n11 1.39274
R159 VTAIL.n2 VTAIL.n1 1.39274
R160 VTAIL VTAIL.n19 0.403517
R161 VP.n17 VP.t6 226.022
R162 VP.n9 VP.t7 193.066
R163 VP.n51 VP.t0 193.066
R164 VP.n58 VP.t4 193.066
R165 VP.n65 VP.t8 193.066
R166 VP.n73 VP.t2 193.066
R167 VP.n40 VP.t3 193.066
R168 VP.n32 VP.t5 193.066
R169 VP.n25 VP.t9 193.066
R170 VP.n18 VP.t1 193.066
R171 VP.n42 VP.n9 184.417
R172 VP.n74 VP.n73 184.417
R173 VP.n41 VP.n40 184.417
R174 VP.n19 VP.n16 161.3
R175 VP.n21 VP.n20 161.3
R176 VP.n22 VP.n15 161.3
R177 VP.n24 VP.n23 161.3
R178 VP.n26 VP.n14 161.3
R179 VP.n28 VP.n27 161.3
R180 VP.n29 VP.n13 161.3
R181 VP.n31 VP.n30 161.3
R182 VP.n33 VP.n12 161.3
R183 VP.n35 VP.n34 161.3
R184 VP.n36 VP.n11 161.3
R185 VP.n38 VP.n37 161.3
R186 VP.n39 VP.n10 161.3
R187 VP.n72 VP.n0 161.3
R188 VP.n71 VP.n70 161.3
R189 VP.n69 VP.n1 161.3
R190 VP.n68 VP.n67 161.3
R191 VP.n66 VP.n2 161.3
R192 VP.n64 VP.n63 161.3
R193 VP.n62 VP.n3 161.3
R194 VP.n61 VP.n60 161.3
R195 VP.n59 VP.n4 161.3
R196 VP.n57 VP.n56 161.3
R197 VP.n55 VP.n5 161.3
R198 VP.n54 VP.n53 161.3
R199 VP.n52 VP.n6 161.3
R200 VP.n50 VP.n49 161.3
R201 VP.n48 VP.n7 161.3
R202 VP.n47 VP.n46 161.3
R203 VP.n45 VP.n8 161.3
R204 VP.n44 VP.n43 161.3
R205 VP.n53 VP.n5 56.5617
R206 VP.n60 VP.n3 56.5617
R207 VP.n27 VP.n13 56.5617
R208 VP.n20 VP.n15 56.5617
R209 VP.n18 VP.n17 50.6216
R210 VP.n42 VP.n41 50.5838
R211 VP.n46 VP.n7 44.4521
R212 VP.n67 VP.n1 44.4521
R213 VP.n34 VP.n11 44.4521
R214 VP.n46 VP.n45 36.702
R215 VP.n71 VP.n1 36.702
R216 VP.n38 VP.n11 36.702
R217 VP.n45 VP.n44 24.5923
R218 VP.n50 VP.n7 24.5923
R219 VP.n53 VP.n52 24.5923
R220 VP.n57 VP.n5 24.5923
R221 VP.n60 VP.n59 24.5923
R222 VP.n64 VP.n3 24.5923
R223 VP.n67 VP.n66 24.5923
R224 VP.n72 VP.n71 24.5923
R225 VP.n39 VP.n38 24.5923
R226 VP.n31 VP.n13 24.5923
R227 VP.n34 VP.n33 24.5923
R228 VP.n24 VP.n15 24.5923
R229 VP.n27 VP.n26 24.5923
R230 VP.n20 VP.n19 24.5923
R231 VP.n52 VP.n51 19.1821
R232 VP.n65 VP.n64 19.1821
R233 VP.n32 VP.n31 19.1821
R234 VP.n19 VP.n18 19.1821
R235 VP.n17 VP.n16 12.4384
R236 VP.n58 VP.n57 12.2964
R237 VP.n59 VP.n58 12.2964
R238 VP.n25 VP.n24 12.2964
R239 VP.n26 VP.n25 12.2964
R240 VP.n51 VP.n50 5.4107
R241 VP.n66 VP.n65 5.4107
R242 VP.n33 VP.n32 5.4107
R243 VP.n44 VP.n9 1.47601
R244 VP.n73 VP.n72 1.47601
R245 VP.n40 VP.n39 1.47601
R246 VP.n21 VP.n16 0.189894
R247 VP.n22 VP.n21 0.189894
R248 VP.n23 VP.n22 0.189894
R249 VP.n23 VP.n14 0.189894
R250 VP.n28 VP.n14 0.189894
R251 VP.n29 VP.n28 0.189894
R252 VP.n30 VP.n29 0.189894
R253 VP.n30 VP.n12 0.189894
R254 VP.n35 VP.n12 0.189894
R255 VP.n36 VP.n35 0.189894
R256 VP.n37 VP.n36 0.189894
R257 VP.n37 VP.n10 0.189894
R258 VP.n41 VP.n10 0.189894
R259 VP.n43 VP.n42 0.189894
R260 VP.n43 VP.n8 0.189894
R261 VP.n47 VP.n8 0.189894
R262 VP.n48 VP.n47 0.189894
R263 VP.n49 VP.n48 0.189894
R264 VP.n49 VP.n6 0.189894
R265 VP.n54 VP.n6 0.189894
R266 VP.n55 VP.n54 0.189894
R267 VP.n56 VP.n55 0.189894
R268 VP.n56 VP.n4 0.189894
R269 VP.n61 VP.n4 0.189894
R270 VP.n62 VP.n61 0.189894
R271 VP.n63 VP.n62 0.189894
R272 VP.n63 VP.n2 0.189894
R273 VP.n68 VP.n2 0.189894
R274 VP.n69 VP.n68 0.189894
R275 VP.n70 VP.n69 0.189894
R276 VP.n70 VP.n0 0.189894
R277 VP.n74 VP.n0 0.189894
R278 VP VP.n74 0.0516364
R279 VDD1.n1 VDD1.t3 79.3957
R280 VDD1.n3 VDD1.t2 79.3956
R281 VDD1.n5 VDD1.n4 76.6373
R282 VDD1.n1 VDD1.n0 75.3093
R283 VDD1.n7 VDD1.n6 75.3091
R284 VDD1.n3 VDD1.n2 75.309
R285 VDD1.n7 VDD1.n5 46.4837
R286 VDD1.n6 VDD1.t4 2.24222
R287 VDD1.n6 VDD1.t6 2.24222
R288 VDD1.n0 VDD1.t8 2.24222
R289 VDD1.n0 VDD1.t0 2.24222
R290 VDD1.n4 VDD1.t1 2.24222
R291 VDD1.n4 VDD1.t7 2.24222
R292 VDD1.n2 VDD1.t9 2.24222
R293 VDD1.n2 VDD1.t5 2.24222
R294 VDD1 VDD1.n7 1.32593
R295 VDD1 VDD1.n1 0.519897
R296 VDD1.n5 VDD1.n3 0.406361
R297 B.n583 B.n582 585
R298 B.n584 B.n83 585
R299 B.n586 B.n585 585
R300 B.n587 B.n82 585
R301 B.n589 B.n588 585
R302 B.n590 B.n81 585
R303 B.n592 B.n591 585
R304 B.n593 B.n80 585
R305 B.n595 B.n594 585
R306 B.n596 B.n79 585
R307 B.n598 B.n597 585
R308 B.n599 B.n78 585
R309 B.n601 B.n600 585
R310 B.n602 B.n77 585
R311 B.n604 B.n603 585
R312 B.n605 B.n76 585
R313 B.n607 B.n606 585
R314 B.n608 B.n75 585
R315 B.n610 B.n609 585
R316 B.n611 B.n74 585
R317 B.n613 B.n612 585
R318 B.n614 B.n73 585
R319 B.n616 B.n615 585
R320 B.n617 B.n72 585
R321 B.n619 B.n618 585
R322 B.n620 B.n71 585
R323 B.n622 B.n621 585
R324 B.n623 B.n70 585
R325 B.n625 B.n624 585
R326 B.n626 B.n69 585
R327 B.n628 B.n627 585
R328 B.n629 B.n68 585
R329 B.n631 B.n630 585
R330 B.n632 B.n67 585
R331 B.n634 B.n633 585
R332 B.n635 B.n66 585
R333 B.n637 B.n636 585
R334 B.n638 B.n65 585
R335 B.n640 B.n639 585
R336 B.n641 B.n64 585
R337 B.n643 B.n642 585
R338 B.n644 B.n63 585
R339 B.n646 B.n645 585
R340 B.n647 B.n62 585
R341 B.n649 B.n648 585
R342 B.n650 B.n61 585
R343 B.n652 B.n651 585
R344 B.n653 B.n57 585
R345 B.n655 B.n654 585
R346 B.n656 B.n56 585
R347 B.n658 B.n657 585
R348 B.n659 B.n55 585
R349 B.n661 B.n660 585
R350 B.n662 B.n54 585
R351 B.n664 B.n663 585
R352 B.n665 B.n53 585
R353 B.n667 B.n666 585
R354 B.n668 B.n52 585
R355 B.n670 B.n669 585
R356 B.n672 B.n49 585
R357 B.n674 B.n673 585
R358 B.n675 B.n48 585
R359 B.n677 B.n676 585
R360 B.n678 B.n47 585
R361 B.n680 B.n679 585
R362 B.n681 B.n46 585
R363 B.n683 B.n682 585
R364 B.n684 B.n45 585
R365 B.n686 B.n685 585
R366 B.n687 B.n44 585
R367 B.n689 B.n688 585
R368 B.n690 B.n43 585
R369 B.n692 B.n691 585
R370 B.n693 B.n42 585
R371 B.n695 B.n694 585
R372 B.n696 B.n41 585
R373 B.n698 B.n697 585
R374 B.n699 B.n40 585
R375 B.n701 B.n700 585
R376 B.n702 B.n39 585
R377 B.n704 B.n703 585
R378 B.n705 B.n38 585
R379 B.n707 B.n706 585
R380 B.n708 B.n37 585
R381 B.n710 B.n709 585
R382 B.n711 B.n36 585
R383 B.n713 B.n712 585
R384 B.n714 B.n35 585
R385 B.n716 B.n715 585
R386 B.n717 B.n34 585
R387 B.n719 B.n718 585
R388 B.n720 B.n33 585
R389 B.n722 B.n721 585
R390 B.n723 B.n32 585
R391 B.n725 B.n724 585
R392 B.n726 B.n31 585
R393 B.n728 B.n727 585
R394 B.n729 B.n30 585
R395 B.n731 B.n730 585
R396 B.n732 B.n29 585
R397 B.n734 B.n733 585
R398 B.n735 B.n28 585
R399 B.n737 B.n736 585
R400 B.n738 B.n27 585
R401 B.n740 B.n739 585
R402 B.n741 B.n26 585
R403 B.n743 B.n742 585
R404 B.n744 B.n25 585
R405 B.n581 B.n84 585
R406 B.n580 B.n579 585
R407 B.n578 B.n85 585
R408 B.n577 B.n576 585
R409 B.n575 B.n86 585
R410 B.n574 B.n573 585
R411 B.n572 B.n87 585
R412 B.n571 B.n570 585
R413 B.n569 B.n88 585
R414 B.n568 B.n567 585
R415 B.n566 B.n89 585
R416 B.n565 B.n564 585
R417 B.n563 B.n90 585
R418 B.n562 B.n561 585
R419 B.n560 B.n91 585
R420 B.n559 B.n558 585
R421 B.n557 B.n92 585
R422 B.n556 B.n555 585
R423 B.n554 B.n93 585
R424 B.n553 B.n552 585
R425 B.n551 B.n94 585
R426 B.n550 B.n549 585
R427 B.n548 B.n95 585
R428 B.n547 B.n546 585
R429 B.n545 B.n96 585
R430 B.n544 B.n543 585
R431 B.n542 B.n97 585
R432 B.n541 B.n540 585
R433 B.n539 B.n98 585
R434 B.n538 B.n537 585
R435 B.n536 B.n99 585
R436 B.n535 B.n534 585
R437 B.n533 B.n100 585
R438 B.n532 B.n531 585
R439 B.n530 B.n101 585
R440 B.n529 B.n528 585
R441 B.n527 B.n102 585
R442 B.n526 B.n525 585
R443 B.n524 B.n103 585
R444 B.n523 B.n522 585
R445 B.n521 B.n104 585
R446 B.n520 B.n519 585
R447 B.n518 B.n105 585
R448 B.n517 B.n516 585
R449 B.n515 B.n106 585
R450 B.n514 B.n513 585
R451 B.n512 B.n107 585
R452 B.n511 B.n510 585
R453 B.n509 B.n108 585
R454 B.n508 B.n507 585
R455 B.n506 B.n109 585
R456 B.n505 B.n504 585
R457 B.n503 B.n110 585
R458 B.n502 B.n501 585
R459 B.n500 B.n111 585
R460 B.n499 B.n498 585
R461 B.n497 B.n112 585
R462 B.n496 B.n495 585
R463 B.n494 B.n113 585
R464 B.n493 B.n492 585
R465 B.n491 B.n114 585
R466 B.n490 B.n489 585
R467 B.n488 B.n115 585
R468 B.n487 B.n486 585
R469 B.n485 B.n116 585
R470 B.n484 B.n483 585
R471 B.n482 B.n117 585
R472 B.n481 B.n480 585
R473 B.n479 B.n118 585
R474 B.n478 B.n477 585
R475 B.n476 B.n119 585
R476 B.n475 B.n474 585
R477 B.n473 B.n120 585
R478 B.n472 B.n471 585
R479 B.n470 B.n121 585
R480 B.n469 B.n468 585
R481 B.n467 B.n122 585
R482 B.n466 B.n465 585
R483 B.n464 B.n123 585
R484 B.n463 B.n462 585
R485 B.n461 B.n124 585
R486 B.n460 B.n459 585
R487 B.n458 B.n125 585
R488 B.n457 B.n456 585
R489 B.n455 B.n126 585
R490 B.n454 B.n453 585
R491 B.n452 B.n127 585
R492 B.n451 B.n450 585
R493 B.n449 B.n128 585
R494 B.n448 B.n447 585
R495 B.n446 B.n129 585
R496 B.n445 B.n444 585
R497 B.n443 B.n130 585
R498 B.n280 B.n279 585
R499 B.n281 B.n188 585
R500 B.n283 B.n282 585
R501 B.n284 B.n187 585
R502 B.n286 B.n285 585
R503 B.n287 B.n186 585
R504 B.n289 B.n288 585
R505 B.n290 B.n185 585
R506 B.n292 B.n291 585
R507 B.n293 B.n184 585
R508 B.n295 B.n294 585
R509 B.n296 B.n183 585
R510 B.n298 B.n297 585
R511 B.n299 B.n182 585
R512 B.n301 B.n300 585
R513 B.n302 B.n181 585
R514 B.n304 B.n303 585
R515 B.n305 B.n180 585
R516 B.n307 B.n306 585
R517 B.n308 B.n179 585
R518 B.n310 B.n309 585
R519 B.n311 B.n178 585
R520 B.n313 B.n312 585
R521 B.n314 B.n177 585
R522 B.n316 B.n315 585
R523 B.n317 B.n176 585
R524 B.n319 B.n318 585
R525 B.n320 B.n175 585
R526 B.n322 B.n321 585
R527 B.n323 B.n174 585
R528 B.n325 B.n324 585
R529 B.n326 B.n173 585
R530 B.n328 B.n327 585
R531 B.n329 B.n172 585
R532 B.n331 B.n330 585
R533 B.n332 B.n171 585
R534 B.n334 B.n333 585
R535 B.n335 B.n170 585
R536 B.n337 B.n336 585
R537 B.n338 B.n169 585
R538 B.n340 B.n339 585
R539 B.n341 B.n168 585
R540 B.n343 B.n342 585
R541 B.n344 B.n167 585
R542 B.n346 B.n345 585
R543 B.n347 B.n166 585
R544 B.n349 B.n348 585
R545 B.n350 B.n165 585
R546 B.n352 B.n351 585
R547 B.n354 B.n162 585
R548 B.n356 B.n355 585
R549 B.n357 B.n161 585
R550 B.n359 B.n358 585
R551 B.n360 B.n160 585
R552 B.n362 B.n361 585
R553 B.n363 B.n159 585
R554 B.n365 B.n364 585
R555 B.n366 B.n158 585
R556 B.n368 B.n367 585
R557 B.n370 B.n369 585
R558 B.n371 B.n154 585
R559 B.n373 B.n372 585
R560 B.n374 B.n153 585
R561 B.n376 B.n375 585
R562 B.n377 B.n152 585
R563 B.n379 B.n378 585
R564 B.n380 B.n151 585
R565 B.n382 B.n381 585
R566 B.n383 B.n150 585
R567 B.n385 B.n384 585
R568 B.n386 B.n149 585
R569 B.n388 B.n387 585
R570 B.n389 B.n148 585
R571 B.n391 B.n390 585
R572 B.n392 B.n147 585
R573 B.n394 B.n393 585
R574 B.n395 B.n146 585
R575 B.n397 B.n396 585
R576 B.n398 B.n145 585
R577 B.n400 B.n399 585
R578 B.n401 B.n144 585
R579 B.n403 B.n402 585
R580 B.n404 B.n143 585
R581 B.n406 B.n405 585
R582 B.n407 B.n142 585
R583 B.n409 B.n408 585
R584 B.n410 B.n141 585
R585 B.n412 B.n411 585
R586 B.n413 B.n140 585
R587 B.n415 B.n414 585
R588 B.n416 B.n139 585
R589 B.n418 B.n417 585
R590 B.n419 B.n138 585
R591 B.n421 B.n420 585
R592 B.n422 B.n137 585
R593 B.n424 B.n423 585
R594 B.n425 B.n136 585
R595 B.n427 B.n426 585
R596 B.n428 B.n135 585
R597 B.n430 B.n429 585
R598 B.n431 B.n134 585
R599 B.n433 B.n432 585
R600 B.n434 B.n133 585
R601 B.n436 B.n435 585
R602 B.n437 B.n132 585
R603 B.n439 B.n438 585
R604 B.n440 B.n131 585
R605 B.n442 B.n441 585
R606 B.n278 B.n189 585
R607 B.n277 B.n276 585
R608 B.n275 B.n190 585
R609 B.n274 B.n273 585
R610 B.n272 B.n191 585
R611 B.n271 B.n270 585
R612 B.n269 B.n192 585
R613 B.n268 B.n267 585
R614 B.n266 B.n193 585
R615 B.n265 B.n264 585
R616 B.n263 B.n194 585
R617 B.n262 B.n261 585
R618 B.n260 B.n195 585
R619 B.n259 B.n258 585
R620 B.n257 B.n196 585
R621 B.n256 B.n255 585
R622 B.n254 B.n197 585
R623 B.n253 B.n252 585
R624 B.n251 B.n198 585
R625 B.n250 B.n249 585
R626 B.n248 B.n199 585
R627 B.n247 B.n246 585
R628 B.n245 B.n200 585
R629 B.n244 B.n243 585
R630 B.n242 B.n201 585
R631 B.n241 B.n240 585
R632 B.n239 B.n202 585
R633 B.n238 B.n237 585
R634 B.n236 B.n203 585
R635 B.n235 B.n234 585
R636 B.n233 B.n204 585
R637 B.n232 B.n231 585
R638 B.n230 B.n205 585
R639 B.n229 B.n228 585
R640 B.n227 B.n206 585
R641 B.n226 B.n225 585
R642 B.n224 B.n207 585
R643 B.n223 B.n222 585
R644 B.n221 B.n208 585
R645 B.n220 B.n219 585
R646 B.n218 B.n209 585
R647 B.n217 B.n216 585
R648 B.n215 B.n210 585
R649 B.n214 B.n213 585
R650 B.n212 B.n211 585
R651 B.n2 B.n0 585
R652 B.n813 B.n1 585
R653 B.n812 B.n811 585
R654 B.n810 B.n3 585
R655 B.n809 B.n808 585
R656 B.n807 B.n4 585
R657 B.n806 B.n805 585
R658 B.n804 B.n5 585
R659 B.n803 B.n802 585
R660 B.n801 B.n6 585
R661 B.n800 B.n799 585
R662 B.n798 B.n7 585
R663 B.n797 B.n796 585
R664 B.n795 B.n8 585
R665 B.n794 B.n793 585
R666 B.n792 B.n9 585
R667 B.n791 B.n790 585
R668 B.n789 B.n10 585
R669 B.n788 B.n787 585
R670 B.n786 B.n11 585
R671 B.n785 B.n784 585
R672 B.n783 B.n12 585
R673 B.n782 B.n781 585
R674 B.n780 B.n13 585
R675 B.n779 B.n778 585
R676 B.n777 B.n14 585
R677 B.n776 B.n775 585
R678 B.n774 B.n15 585
R679 B.n773 B.n772 585
R680 B.n771 B.n16 585
R681 B.n770 B.n769 585
R682 B.n768 B.n17 585
R683 B.n767 B.n766 585
R684 B.n765 B.n18 585
R685 B.n764 B.n763 585
R686 B.n762 B.n19 585
R687 B.n761 B.n760 585
R688 B.n759 B.n20 585
R689 B.n758 B.n757 585
R690 B.n756 B.n21 585
R691 B.n755 B.n754 585
R692 B.n753 B.n22 585
R693 B.n752 B.n751 585
R694 B.n750 B.n23 585
R695 B.n749 B.n748 585
R696 B.n747 B.n24 585
R697 B.n746 B.n745 585
R698 B.n815 B.n814 585
R699 B.n279 B.n278 439.647
R700 B.n746 B.n25 439.647
R701 B.n441 B.n130 439.647
R702 B.n583 B.n84 439.647
R703 B.n155 B.t9 399.5
R704 B.n163 B.t0 399.5
R705 B.n50 B.t3 399.5
R706 B.n58 B.t6 399.5
R707 B.n278 B.n277 163.367
R708 B.n277 B.n190 163.367
R709 B.n273 B.n190 163.367
R710 B.n273 B.n272 163.367
R711 B.n272 B.n271 163.367
R712 B.n271 B.n192 163.367
R713 B.n267 B.n192 163.367
R714 B.n267 B.n266 163.367
R715 B.n266 B.n265 163.367
R716 B.n265 B.n194 163.367
R717 B.n261 B.n194 163.367
R718 B.n261 B.n260 163.367
R719 B.n260 B.n259 163.367
R720 B.n259 B.n196 163.367
R721 B.n255 B.n196 163.367
R722 B.n255 B.n254 163.367
R723 B.n254 B.n253 163.367
R724 B.n253 B.n198 163.367
R725 B.n249 B.n198 163.367
R726 B.n249 B.n248 163.367
R727 B.n248 B.n247 163.367
R728 B.n247 B.n200 163.367
R729 B.n243 B.n200 163.367
R730 B.n243 B.n242 163.367
R731 B.n242 B.n241 163.367
R732 B.n241 B.n202 163.367
R733 B.n237 B.n202 163.367
R734 B.n237 B.n236 163.367
R735 B.n236 B.n235 163.367
R736 B.n235 B.n204 163.367
R737 B.n231 B.n204 163.367
R738 B.n231 B.n230 163.367
R739 B.n230 B.n229 163.367
R740 B.n229 B.n206 163.367
R741 B.n225 B.n206 163.367
R742 B.n225 B.n224 163.367
R743 B.n224 B.n223 163.367
R744 B.n223 B.n208 163.367
R745 B.n219 B.n208 163.367
R746 B.n219 B.n218 163.367
R747 B.n218 B.n217 163.367
R748 B.n217 B.n210 163.367
R749 B.n213 B.n210 163.367
R750 B.n213 B.n212 163.367
R751 B.n212 B.n2 163.367
R752 B.n814 B.n2 163.367
R753 B.n814 B.n813 163.367
R754 B.n813 B.n812 163.367
R755 B.n812 B.n3 163.367
R756 B.n808 B.n3 163.367
R757 B.n808 B.n807 163.367
R758 B.n807 B.n806 163.367
R759 B.n806 B.n5 163.367
R760 B.n802 B.n5 163.367
R761 B.n802 B.n801 163.367
R762 B.n801 B.n800 163.367
R763 B.n800 B.n7 163.367
R764 B.n796 B.n7 163.367
R765 B.n796 B.n795 163.367
R766 B.n795 B.n794 163.367
R767 B.n794 B.n9 163.367
R768 B.n790 B.n9 163.367
R769 B.n790 B.n789 163.367
R770 B.n789 B.n788 163.367
R771 B.n788 B.n11 163.367
R772 B.n784 B.n11 163.367
R773 B.n784 B.n783 163.367
R774 B.n783 B.n782 163.367
R775 B.n782 B.n13 163.367
R776 B.n778 B.n13 163.367
R777 B.n778 B.n777 163.367
R778 B.n777 B.n776 163.367
R779 B.n776 B.n15 163.367
R780 B.n772 B.n15 163.367
R781 B.n772 B.n771 163.367
R782 B.n771 B.n770 163.367
R783 B.n770 B.n17 163.367
R784 B.n766 B.n17 163.367
R785 B.n766 B.n765 163.367
R786 B.n765 B.n764 163.367
R787 B.n764 B.n19 163.367
R788 B.n760 B.n19 163.367
R789 B.n760 B.n759 163.367
R790 B.n759 B.n758 163.367
R791 B.n758 B.n21 163.367
R792 B.n754 B.n21 163.367
R793 B.n754 B.n753 163.367
R794 B.n753 B.n752 163.367
R795 B.n752 B.n23 163.367
R796 B.n748 B.n23 163.367
R797 B.n748 B.n747 163.367
R798 B.n747 B.n746 163.367
R799 B.n279 B.n188 163.367
R800 B.n283 B.n188 163.367
R801 B.n284 B.n283 163.367
R802 B.n285 B.n284 163.367
R803 B.n285 B.n186 163.367
R804 B.n289 B.n186 163.367
R805 B.n290 B.n289 163.367
R806 B.n291 B.n290 163.367
R807 B.n291 B.n184 163.367
R808 B.n295 B.n184 163.367
R809 B.n296 B.n295 163.367
R810 B.n297 B.n296 163.367
R811 B.n297 B.n182 163.367
R812 B.n301 B.n182 163.367
R813 B.n302 B.n301 163.367
R814 B.n303 B.n302 163.367
R815 B.n303 B.n180 163.367
R816 B.n307 B.n180 163.367
R817 B.n308 B.n307 163.367
R818 B.n309 B.n308 163.367
R819 B.n309 B.n178 163.367
R820 B.n313 B.n178 163.367
R821 B.n314 B.n313 163.367
R822 B.n315 B.n314 163.367
R823 B.n315 B.n176 163.367
R824 B.n319 B.n176 163.367
R825 B.n320 B.n319 163.367
R826 B.n321 B.n320 163.367
R827 B.n321 B.n174 163.367
R828 B.n325 B.n174 163.367
R829 B.n326 B.n325 163.367
R830 B.n327 B.n326 163.367
R831 B.n327 B.n172 163.367
R832 B.n331 B.n172 163.367
R833 B.n332 B.n331 163.367
R834 B.n333 B.n332 163.367
R835 B.n333 B.n170 163.367
R836 B.n337 B.n170 163.367
R837 B.n338 B.n337 163.367
R838 B.n339 B.n338 163.367
R839 B.n339 B.n168 163.367
R840 B.n343 B.n168 163.367
R841 B.n344 B.n343 163.367
R842 B.n345 B.n344 163.367
R843 B.n345 B.n166 163.367
R844 B.n349 B.n166 163.367
R845 B.n350 B.n349 163.367
R846 B.n351 B.n350 163.367
R847 B.n351 B.n162 163.367
R848 B.n356 B.n162 163.367
R849 B.n357 B.n356 163.367
R850 B.n358 B.n357 163.367
R851 B.n358 B.n160 163.367
R852 B.n362 B.n160 163.367
R853 B.n363 B.n362 163.367
R854 B.n364 B.n363 163.367
R855 B.n364 B.n158 163.367
R856 B.n368 B.n158 163.367
R857 B.n369 B.n368 163.367
R858 B.n369 B.n154 163.367
R859 B.n373 B.n154 163.367
R860 B.n374 B.n373 163.367
R861 B.n375 B.n374 163.367
R862 B.n375 B.n152 163.367
R863 B.n379 B.n152 163.367
R864 B.n380 B.n379 163.367
R865 B.n381 B.n380 163.367
R866 B.n381 B.n150 163.367
R867 B.n385 B.n150 163.367
R868 B.n386 B.n385 163.367
R869 B.n387 B.n386 163.367
R870 B.n387 B.n148 163.367
R871 B.n391 B.n148 163.367
R872 B.n392 B.n391 163.367
R873 B.n393 B.n392 163.367
R874 B.n393 B.n146 163.367
R875 B.n397 B.n146 163.367
R876 B.n398 B.n397 163.367
R877 B.n399 B.n398 163.367
R878 B.n399 B.n144 163.367
R879 B.n403 B.n144 163.367
R880 B.n404 B.n403 163.367
R881 B.n405 B.n404 163.367
R882 B.n405 B.n142 163.367
R883 B.n409 B.n142 163.367
R884 B.n410 B.n409 163.367
R885 B.n411 B.n410 163.367
R886 B.n411 B.n140 163.367
R887 B.n415 B.n140 163.367
R888 B.n416 B.n415 163.367
R889 B.n417 B.n416 163.367
R890 B.n417 B.n138 163.367
R891 B.n421 B.n138 163.367
R892 B.n422 B.n421 163.367
R893 B.n423 B.n422 163.367
R894 B.n423 B.n136 163.367
R895 B.n427 B.n136 163.367
R896 B.n428 B.n427 163.367
R897 B.n429 B.n428 163.367
R898 B.n429 B.n134 163.367
R899 B.n433 B.n134 163.367
R900 B.n434 B.n433 163.367
R901 B.n435 B.n434 163.367
R902 B.n435 B.n132 163.367
R903 B.n439 B.n132 163.367
R904 B.n440 B.n439 163.367
R905 B.n441 B.n440 163.367
R906 B.n445 B.n130 163.367
R907 B.n446 B.n445 163.367
R908 B.n447 B.n446 163.367
R909 B.n447 B.n128 163.367
R910 B.n451 B.n128 163.367
R911 B.n452 B.n451 163.367
R912 B.n453 B.n452 163.367
R913 B.n453 B.n126 163.367
R914 B.n457 B.n126 163.367
R915 B.n458 B.n457 163.367
R916 B.n459 B.n458 163.367
R917 B.n459 B.n124 163.367
R918 B.n463 B.n124 163.367
R919 B.n464 B.n463 163.367
R920 B.n465 B.n464 163.367
R921 B.n465 B.n122 163.367
R922 B.n469 B.n122 163.367
R923 B.n470 B.n469 163.367
R924 B.n471 B.n470 163.367
R925 B.n471 B.n120 163.367
R926 B.n475 B.n120 163.367
R927 B.n476 B.n475 163.367
R928 B.n477 B.n476 163.367
R929 B.n477 B.n118 163.367
R930 B.n481 B.n118 163.367
R931 B.n482 B.n481 163.367
R932 B.n483 B.n482 163.367
R933 B.n483 B.n116 163.367
R934 B.n487 B.n116 163.367
R935 B.n488 B.n487 163.367
R936 B.n489 B.n488 163.367
R937 B.n489 B.n114 163.367
R938 B.n493 B.n114 163.367
R939 B.n494 B.n493 163.367
R940 B.n495 B.n494 163.367
R941 B.n495 B.n112 163.367
R942 B.n499 B.n112 163.367
R943 B.n500 B.n499 163.367
R944 B.n501 B.n500 163.367
R945 B.n501 B.n110 163.367
R946 B.n505 B.n110 163.367
R947 B.n506 B.n505 163.367
R948 B.n507 B.n506 163.367
R949 B.n507 B.n108 163.367
R950 B.n511 B.n108 163.367
R951 B.n512 B.n511 163.367
R952 B.n513 B.n512 163.367
R953 B.n513 B.n106 163.367
R954 B.n517 B.n106 163.367
R955 B.n518 B.n517 163.367
R956 B.n519 B.n518 163.367
R957 B.n519 B.n104 163.367
R958 B.n523 B.n104 163.367
R959 B.n524 B.n523 163.367
R960 B.n525 B.n524 163.367
R961 B.n525 B.n102 163.367
R962 B.n529 B.n102 163.367
R963 B.n530 B.n529 163.367
R964 B.n531 B.n530 163.367
R965 B.n531 B.n100 163.367
R966 B.n535 B.n100 163.367
R967 B.n536 B.n535 163.367
R968 B.n537 B.n536 163.367
R969 B.n537 B.n98 163.367
R970 B.n541 B.n98 163.367
R971 B.n542 B.n541 163.367
R972 B.n543 B.n542 163.367
R973 B.n543 B.n96 163.367
R974 B.n547 B.n96 163.367
R975 B.n548 B.n547 163.367
R976 B.n549 B.n548 163.367
R977 B.n549 B.n94 163.367
R978 B.n553 B.n94 163.367
R979 B.n554 B.n553 163.367
R980 B.n555 B.n554 163.367
R981 B.n555 B.n92 163.367
R982 B.n559 B.n92 163.367
R983 B.n560 B.n559 163.367
R984 B.n561 B.n560 163.367
R985 B.n561 B.n90 163.367
R986 B.n565 B.n90 163.367
R987 B.n566 B.n565 163.367
R988 B.n567 B.n566 163.367
R989 B.n567 B.n88 163.367
R990 B.n571 B.n88 163.367
R991 B.n572 B.n571 163.367
R992 B.n573 B.n572 163.367
R993 B.n573 B.n86 163.367
R994 B.n577 B.n86 163.367
R995 B.n578 B.n577 163.367
R996 B.n579 B.n578 163.367
R997 B.n579 B.n84 163.367
R998 B.n742 B.n25 163.367
R999 B.n742 B.n741 163.367
R1000 B.n741 B.n740 163.367
R1001 B.n740 B.n27 163.367
R1002 B.n736 B.n27 163.367
R1003 B.n736 B.n735 163.367
R1004 B.n735 B.n734 163.367
R1005 B.n734 B.n29 163.367
R1006 B.n730 B.n29 163.367
R1007 B.n730 B.n729 163.367
R1008 B.n729 B.n728 163.367
R1009 B.n728 B.n31 163.367
R1010 B.n724 B.n31 163.367
R1011 B.n724 B.n723 163.367
R1012 B.n723 B.n722 163.367
R1013 B.n722 B.n33 163.367
R1014 B.n718 B.n33 163.367
R1015 B.n718 B.n717 163.367
R1016 B.n717 B.n716 163.367
R1017 B.n716 B.n35 163.367
R1018 B.n712 B.n35 163.367
R1019 B.n712 B.n711 163.367
R1020 B.n711 B.n710 163.367
R1021 B.n710 B.n37 163.367
R1022 B.n706 B.n37 163.367
R1023 B.n706 B.n705 163.367
R1024 B.n705 B.n704 163.367
R1025 B.n704 B.n39 163.367
R1026 B.n700 B.n39 163.367
R1027 B.n700 B.n699 163.367
R1028 B.n699 B.n698 163.367
R1029 B.n698 B.n41 163.367
R1030 B.n694 B.n41 163.367
R1031 B.n694 B.n693 163.367
R1032 B.n693 B.n692 163.367
R1033 B.n692 B.n43 163.367
R1034 B.n688 B.n43 163.367
R1035 B.n688 B.n687 163.367
R1036 B.n687 B.n686 163.367
R1037 B.n686 B.n45 163.367
R1038 B.n682 B.n45 163.367
R1039 B.n682 B.n681 163.367
R1040 B.n681 B.n680 163.367
R1041 B.n680 B.n47 163.367
R1042 B.n676 B.n47 163.367
R1043 B.n676 B.n675 163.367
R1044 B.n675 B.n674 163.367
R1045 B.n674 B.n49 163.367
R1046 B.n669 B.n49 163.367
R1047 B.n669 B.n668 163.367
R1048 B.n668 B.n667 163.367
R1049 B.n667 B.n53 163.367
R1050 B.n663 B.n53 163.367
R1051 B.n663 B.n662 163.367
R1052 B.n662 B.n661 163.367
R1053 B.n661 B.n55 163.367
R1054 B.n657 B.n55 163.367
R1055 B.n657 B.n656 163.367
R1056 B.n656 B.n655 163.367
R1057 B.n655 B.n57 163.367
R1058 B.n651 B.n57 163.367
R1059 B.n651 B.n650 163.367
R1060 B.n650 B.n649 163.367
R1061 B.n649 B.n62 163.367
R1062 B.n645 B.n62 163.367
R1063 B.n645 B.n644 163.367
R1064 B.n644 B.n643 163.367
R1065 B.n643 B.n64 163.367
R1066 B.n639 B.n64 163.367
R1067 B.n639 B.n638 163.367
R1068 B.n638 B.n637 163.367
R1069 B.n637 B.n66 163.367
R1070 B.n633 B.n66 163.367
R1071 B.n633 B.n632 163.367
R1072 B.n632 B.n631 163.367
R1073 B.n631 B.n68 163.367
R1074 B.n627 B.n68 163.367
R1075 B.n627 B.n626 163.367
R1076 B.n626 B.n625 163.367
R1077 B.n625 B.n70 163.367
R1078 B.n621 B.n70 163.367
R1079 B.n621 B.n620 163.367
R1080 B.n620 B.n619 163.367
R1081 B.n619 B.n72 163.367
R1082 B.n615 B.n72 163.367
R1083 B.n615 B.n614 163.367
R1084 B.n614 B.n613 163.367
R1085 B.n613 B.n74 163.367
R1086 B.n609 B.n74 163.367
R1087 B.n609 B.n608 163.367
R1088 B.n608 B.n607 163.367
R1089 B.n607 B.n76 163.367
R1090 B.n603 B.n76 163.367
R1091 B.n603 B.n602 163.367
R1092 B.n602 B.n601 163.367
R1093 B.n601 B.n78 163.367
R1094 B.n597 B.n78 163.367
R1095 B.n597 B.n596 163.367
R1096 B.n596 B.n595 163.367
R1097 B.n595 B.n80 163.367
R1098 B.n591 B.n80 163.367
R1099 B.n591 B.n590 163.367
R1100 B.n590 B.n589 163.367
R1101 B.n589 B.n82 163.367
R1102 B.n585 B.n82 163.367
R1103 B.n585 B.n584 163.367
R1104 B.n584 B.n583 163.367
R1105 B.n155 B.t11 152.405
R1106 B.n58 B.t7 152.405
R1107 B.n163 B.t2 152.387
R1108 B.n50 B.t4 152.387
R1109 B.n156 B.t10 110.903
R1110 B.n59 B.t8 110.903
R1111 B.n164 B.t1 110.885
R1112 B.n51 B.t5 110.885
R1113 B.n157 B.n156 59.5399
R1114 B.n353 B.n164 59.5399
R1115 B.n671 B.n51 59.5399
R1116 B.n60 B.n59 59.5399
R1117 B.n156 B.n155 41.5035
R1118 B.n164 B.n163 41.5035
R1119 B.n51 B.n50 41.5035
R1120 B.n59 B.n58 41.5035
R1121 B.n582 B.n581 28.5664
R1122 B.n745 B.n744 28.5664
R1123 B.n443 B.n442 28.5664
R1124 B.n280 B.n189 28.5664
R1125 B B.n815 18.0485
R1126 B.n744 B.n743 10.6151
R1127 B.n743 B.n26 10.6151
R1128 B.n739 B.n26 10.6151
R1129 B.n739 B.n738 10.6151
R1130 B.n738 B.n737 10.6151
R1131 B.n737 B.n28 10.6151
R1132 B.n733 B.n28 10.6151
R1133 B.n733 B.n732 10.6151
R1134 B.n732 B.n731 10.6151
R1135 B.n731 B.n30 10.6151
R1136 B.n727 B.n30 10.6151
R1137 B.n727 B.n726 10.6151
R1138 B.n726 B.n725 10.6151
R1139 B.n725 B.n32 10.6151
R1140 B.n721 B.n32 10.6151
R1141 B.n721 B.n720 10.6151
R1142 B.n720 B.n719 10.6151
R1143 B.n719 B.n34 10.6151
R1144 B.n715 B.n34 10.6151
R1145 B.n715 B.n714 10.6151
R1146 B.n714 B.n713 10.6151
R1147 B.n713 B.n36 10.6151
R1148 B.n709 B.n36 10.6151
R1149 B.n709 B.n708 10.6151
R1150 B.n708 B.n707 10.6151
R1151 B.n707 B.n38 10.6151
R1152 B.n703 B.n38 10.6151
R1153 B.n703 B.n702 10.6151
R1154 B.n702 B.n701 10.6151
R1155 B.n701 B.n40 10.6151
R1156 B.n697 B.n40 10.6151
R1157 B.n697 B.n696 10.6151
R1158 B.n696 B.n695 10.6151
R1159 B.n695 B.n42 10.6151
R1160 B.n691 B.n42 10.6151
R1161 B.n691 B.n690 10.6151
R1162 B.n690 B.n689 10.6151
R1163 B.n689 B.n44 10.6151
R1164 B.n685 B.n44 10.6151
R1165 B.n685 B.n684 10.6151
R1166 B.n684 B.n683 10.6151
R1167 B.n683 B.n46 10.6151
R1168 B.n679 B.n46 10.6151
R1169 B.n679 B.n678 10.6151
R1170 B.n678 B.n677 10.6151
R1171 B.n677 B.n48 10.6151
R1172 B.n673 B.n48 10.6151
R1173 B.n673 B.n672 10.6151
R1174 B.n670 B.n52 10.6151
R1175 B.n666 B.n52 10.6151
R1176 B.n666 B.n665 10.6151
R1177 B.n665 B.n664 10.6151
R1178 B.n664 B.n54 10.6151
R1179 B.n660 B.n54 10.6151
R1180 B.n660 B.n659 10.6151
R1181 B.n659 B.n658 10.6151
R1182 B.n658 B.n56 10.6151
R1183 B.n654 B.n653 10.6151
R1184 B.n653 B.n652 10.6151
R1185 B.n652 B.n61 10.6151
R1186 B.n648 B.n61 10.6151
R1187 B.n648 B.n647 10.6151
R1188 B.n647 B.n646 10.6151
R1189 B.n646 B.n63 10.6151
R1190 B.n642 B.n63 10.6151
R1191 B.n642 B.n641 10.6151
R1192 B.n641 B.n640 10.6151
R1193 B.n640 B.n65 10.6151
R1194 B.n636 B.n65 10.6151
R1195 B.n636 B.n635 10.6151
R1196 B.n635 B.n634 10.6151
R1197 B.n634 B.n67 10.6151
R1198 B.n630 B.n67 10.6151
R1199 B.n630 B.n629 10.6151
R1200 B.n629 B.n628 10.6151
R1201 B.n628 B.n69 10.6151
R1202 B.n624 B.n69 10.6151
R1203 B.n624 B.n623 10.6151
R1204 B.n623 B.n622 10.6151
R1205 B.n622 B.n71 10.6151
R1206 B.n618 B.n71 10.6151
R1207 B.n618 B.n617 10.6151
R1208 B.n617 B.n616 10.6151
R1209 B.n616 B.n73 10.6151
R1210 B.n612 B.n73 10.6151
R1211 B.n612 B.n611 10.6151
R1212 B.n611 B.n610 10.6151
R1213 B.n610 B.n75 10.6151
R1214 B.n606 B.n75 10.6151
R1215 B.n606 B.n605 10.6151
R1216 B.n605 B.n604 10.6151
R1217 B.n604 B.n77 10.6151
R1218 B.n600 B.n77 10.6151
R1219 B.n600 B.n599 10.6151
R1220 B.n599 B.n598 10.6151
R1221 B.n598 B.n79 10.6151
R1222 B.n594 B.n79 10.6151
R1223 B.n594 B.n593 10.6151
R1224 B.n593 B.n592 10.6151
R1225 B.n592 B.n81 10.6151
R1226 B.n588 B.n81 10.6151
R1227 B.n588 B.n587 10.6151
R1228 B.n587 B.n586 10.6151
R1229 B.n586 B.n83 10.6151
R1230 B.n582 B.n83 10.6151
R1231 B.n444 B.n443 10.6151
R1232 B.n444 B.n129 10.6151
R1233 B.n448 B.n129 10.6151
R1234 B.n449 B.n448 10.6151
R1235 B.n450 B.n449 10.6151
R1236 B.n450 B.n127 10.6151
R1237 B.n454 B.n127 10.6151
R1238 B.n455 B.n454 10.6151
R1239 B.n456 B.n455 10.6151
R1240 B.n456 B.n125 10.6151
R1241 B.n460 B.n125 10.6151
R1242 B.n461 B.n460 10.6151
R1243 B.n462 B.n461 10.6151
R1244 B.n462 B.n123 10.6151
R1245 B.n466 B.n123 10.6151
R1246 B.n467 B.n466 10.6151
R1247 B.n468 B.n467 10.6151
R1248 B.n468 B.n121 10.6151
R1249 B.n472 B.n121 10.6151
R1250 B.n473 B.n472 10.6151
R1251 B.n474 B.n473 10.6151
R1252 B.n474 B.n119 10.6151
R1253 B.n478 B.n119 10.6151
R1254 B.n479 B.n478 10.6151
R1255 B.n480 B.n479 10.6151
R1256 B.n480 B.n117 10.6151
R1257 B.n484 B.n117 10.6151
R1258 B.n485 B.n484 10.6151
R1259 B.n486 B.n485 10.6151
R1260 B.n486 B.n115 10.6151
R1261 B.n490 B.n115 10.6151
R1262 B.n491 B.n490 10.6151
R1263 B.n492 B.n491 10.6151
R1264 B.n492 B.n113 10.6151
R1265 B.n496 B.n113 10.6151
R1266 B.n497 B.n496 10.6151
R1267 B.n498 B.n497 10.6151
R1268 B.n498 B.n111 10.6151
R1269 B.n502 B.n111 10.6151
R1270 B.n503 B.n502 10.6151
R1271 B.n504 B.n503 10.6151
R1272 B.n504 B.n109 10.6151
R1273 B.n508 B.n109 10.6151
R1274 B.n509 B.n508 10.6151
R1275 B.n510 B.n509 10.6151
R1276 B.n510 B.n107 10.6151
R1277 B.n514 B.n107 10.6151
R1278 B.n515 B.n514 10.6151
R1279 B.n516 B.n515 10.6151
R1280 B.n516 B.n105 10.6151
R1281 B.n520 B.n105 10.6151
R1282 B.n521 B.n520 10.6151
R1283 B.n522 B.n521 10.6151
R1284 B.n522 B.n103 10.6151
R1285 B.n526 B.n103 10.6151
R1286 B.n527 B.n526 10.6151
R1287 B.n528 B.n527 10.6151
R1288 B.n528 B.n101 10.6151
R1289 B.n532 B.n101 10.6151
R1290 B.n533 B.n532 10.6151
R1291 B.n534 B.n533 10.6151
R1292 B.n534 B.n99 10.6151
R1293 B.n538 B.n99 10.6151
R1294 B.n539 B.n538 10.6151
R1295 B.n540 B.n539 10.6151
R1296 B.n540 B.n97 10.6151
R1297 B.n544 B.n97 10.6151
R1298 B.n545 B.n544 10.6151
R1299 B.n546 B.n545 10.6151
R1300 B.n546 B.n95 10.6151
R1301 B.n550 B.n95 10.6151
R1302 B.n551 B.n550 10.6151
R1303 B.n552 B.n551 10.6151
R1304 B.n552 B.n93 10.6151
R1305 B.n556 B.n93 10.6151
R1306 B.n557 B.n556 10.6151
R1307 B.n558 B.n557 10.6151
R1308 B.n558 B.n91 10.6151
R1309 B.n562 B.n91 10.6151
R1310 B.n563 B.n562 10.6151
R1311 B.n564 B.n563 10.6151
R1312 B.n564 B.n89 10.6151
R1313 B.n568 B.n89 10.6151
R1314 B.n569 B.n568 10.6151
R1315 B.n570 B.n569 10.6151
R1316 B.n570 B.n87 10.6151
R1317 B.n574 B.n87 10.6151
R1318 B.n575 B.n574 10.6151
R1319 B.n576 B.n575 10.6151
R1320 B.n576 B.n85 10.6151
R1321 B.n580 B.n85 10.6151
R1322 B.n581 B.n580 10.6151
R1323 B.n281 B.n280 10.6151
R1324 B.n282 B.n281 10.6151
R1325 B.n282 B.n187 10.6151
R1326 B.n286 B.n187 10.6151
R1327 B.n287 B.n286 10.6151
R1328 B.n288 B.n287 10.6151
R1329 B.n288 B.n185 10.6151
R1330 B.n292 B.n185 10.6151
R1331 B.n293 B.n292 10.6151
R1332 B.n294 B.n293 10.6151
R1333 B.n294 B.n183 10.6151
R1334 B.n298 B.n183 10.6151
R1335 B.n299 B.n298 10.6151
R1336 B.n300 B.n299 10.6151
R1337 B.n300 B.n181 10.6151
R1338 B.n304 B.n181 10.6151
R1339 B.n305 B.n304 10.6151
R1340 B.n306 B.n305 10.6151
R1341 B.n306 B.n179 10.6151
R1342 B.n310 B.n179 10.6151
R1343 B.n311 B.n310 10.6151
R1344 B.n312 B.n311 10.6151
R1345 B.n312 B.n177 10.6151
R1346 B.n316 B.n177 10.6151
R1347 B.n317 B.n316 10.6151
R1348 B.n318 B.n317 10.6151
R1349 B.n318 B.n175 10.6151
R1350 B.n322 B.n175 10.6151
R1351 B.n323 B.n322 10.6151
R1352 B.n324 B.n323 10.6151
R1353 B.n324 B.n173 10.6151
R1354 B.n328 B.n173 10.6151
R1355 B.n329 B.n328 10.6151
R1356 B.n330 B.n329 10.6151
R1357 B.n330 B.n171 10.6151
R1358 B.n334 B.n171 10.6151
R1359 B.n335 B.n334 10.6151
R1360 B.n336 B.n335 10.6151
R1361 B.n336 B.n169 10.6151
R1362 B.n340 B.n169 10.6151
R1363 B.n341 B.n340 10.6151
R1364 B.n342 B.n341 10.6151
R1365 B.n342 B.n167 10.6151
R1366 B.n346 B.n167 10.6151
R1367 B.n347 B.n346 10.6151
R1368 B.n348 B.n347 10.6151
R1369 B.n348 B.n165 10.6151
R1370 B.n352 B.n165 10.6151
R1371 B.n355 B.n354 10.6151
R1372 B.n355 B.n161 10.6151
R1373 B.n359 B.n161 10.6151
R1374 B.n360 B.n359 10.6151
R1375 B.n361 B.n360 10.6151
R1376 B.n361 B.n159 10.6151
R1377 B.n365 B.n159 10.6151
R1378 B.n366 B.n365 10.6151
R1379 B.n367 B.n366 10.6151
R1380 B.n371 B.n370 10.6151
R1381 B.n372 B.n371 10.6151
R1382 B.n372 B.n153 10.6151
R1383 B.n376 B.n153 10.6151
R1384 B.n377 B.n376 10.6151
R1385 B.n378 B.n377 10.6151
R1386 B.n378 B.n151 10.6151
R1387 B.n382 B.n151 10.6151
R1388 B.n383 B.n382 10.6151
R1389 B.n384 B.n383 10.6151
R1390 B.n384 B.n149 10.6151
R1391 B.n388 B.n149 10.6151
R1392 B.n389 B.n388 10.6151
R1393 B.n390 B.n389 10.6151
R1394 B.n390 B.n147 10.6151
R1395 B.n394 B.n147 10.6151
R1396 B.n395 B.n394 10.6151
R1397 B.n396 B.n395 10.6151
R1398 B.n396 B.n145 10.6151
R1399 B.n400 B.n145 10.6151
R1400 B.n401 B.n400 10.6151
R1401 B.n402 B.n401 10.6151
R1402 B.n402 B.n143 10.6151
R1403 B.n406 B.n143 10.6151
R1404 B.n407 B.n406 10.6151
R1405 B.n408 B.n407 10.6151
R1406 B.n408 B.n141 10.6151
R1407 B.n412 B.n141 10.6151
R1408 B.n413 B.n412 10.6151
R1409 B.n414 B.n413 10.6151
R1410 B.n414 B.n139 10.6151
R1411 B.n418 B.n139 10.6151
R1412 B.n419 B.n418 10.6151
R1413 B.n420 B.n419 10.6151
R1414 B.n420 B.n137 10.6151
R1415 B.n424 B.n137 10.6151
R1416 B.n425 B.n424 10.6151
R1417 B.n426 B.n425 10.6151
R1418 B.n426 B.n135 10.6151
R1419 B.n430 B.n135 10.6151
R1420 B.n431 B.n430 10.6151
R1421 B.n432 B.n431 10.6151
R1422 B.n432 B.n133 10.6151
R1423 B.n436 B.n133 10.6151
R1424 B.n437 B.n436 10.6151
R1425 B.n438 B.n437 10.6151
R1426 B.n438 B.n131 10.6151
R1427 B.n442 B.n131 10.6151
R1428 B.n276 B.n189 10.6151
R1429 B.n276 B.n275 10.6151
R1430 B.n275 B.n274 10.6151
R1431 B.n274 B.n191 10.6151
R1432 B.n270 B.n191 10.6151
R1433 B.n270 B.n269 10.6151
R1434 B.n269 B.n268 10.6151
R1435 B.n268 B.n193 10.6151
R1436 B.n264 B.n193 10.6151
R1437 B.n264 B.n263 10.6151
R1438 B.n263 B.n262 10.6151
R1439 B.n262 B.n195 10.6151
R1440 B.n258 B.n195 10.6151
R1441 B.n258 B.n257 10.6151
R1442 B.n257 B.n256 10.6151
R1443 B.n256 B.n197 10.6151
R1444 B.n252 B.n197 10.6151
R1445 B.n252 B.n251 10.6151
R1446 B.n251 B.n250 10.6151
R1447 B.n250 B.n199 10.6151
R1448 B.n246 B.n199 10.6151
R1449 B.n246 B.n245 10.6151
R1450 B.n245 B.n244 10.6151
R1451 B.n244 B.n201 10.6151
R1452 B.n240 B.n201 10.6151
R1453 B.n240 B.n239 10.6151
R1454 B.n239 B.n238 10.6151
R1455 B.n238 B.n203 10.6151
R1456 B.n234 B.n203 10.6151
R1457 B.n234 B.n233 10.6151
R1458 B.n233 B.n232 10.6151
R1459 B.n232 B.n205 10.6151
R1460 B.n228 B.n205 10.6151
R1461 B.n228 B.n227 10.6151
R1462 B.n227 B.n226 10.6151
R1463 B.n226 B.n207 10.6151
R1464 B.n222 B.n207 10.6151
R1465 B.n222 B.n221 10.6151
R1466 B.n221 B.n220 10.6151
R1467 B.n220 B.n209 10.6151
R1468 B.n216 B.n209 10.6151
R1469 B.n216 B.n215 10.6151
R1470 B.n215 B.n214 10.6151
R1471 B.n214 B.n211 10.6151
R1472 B.n211 B.n0 10.6151
R1473 B.n811 B.n1 10.6151
R1474 B.n811 B.n810 10.6151
R1475 B.n810 B.n809 10.6151
R1476 B.n809 B.n4 10.6151
R1477 B.n805 B.n4 10.6151
R1478 B.n805 B.n804 10.6151
R1479 B.n804 B.n803 10.6151
R1480 B.n803 B.n6 10.6151
R1481 B.n799 B.n6 10.6151
R1482 B.n799 B.n798 10.6151
R1483 B.n798 B.n797 10.6151
R1484 B.n797 B.n8 10.6151
R1485 B.n793 B.n8 10.6151
R1486 B.n793 B.n792 10.6151
R1487 B.n792 B.n791 10.6151
R1488 B.n791 B.n10 10.6151
R1489 B.n787 B.n10 10.6151
R1490 B.n787 B.n786 10.6151
R1491 B.n786 B.n785 10.6151
R1492 B.n785 B.n12 10.6151
R1493 B.n781 B.n12 10.6151
R1494 B.n781 B.n780 10.6151
R1495 B.n780 B.n779 10.6151
R1496 B.n779 B.n14 10.6151
R1497 B.n775 B.n14 10.6151
R1498 B.n775 B.n774 10.6151
R1499 B.n774 B.n773 10.6151
R1500 B.n773 B.n16 10.6151
R1501 B.n769 B.n16 10.6151
R1502 B.n769 B.n768 10.6151
R1503 B.n768 B.n767 10.6151
R1504 B.n767 B.n18 10.6151
R1505 B.n763 B.n18 10.6151
R1506 B.n763 B.n762 10.6151
R1507 B.n762 B.n761 10.6151
R1508 B.n761 B.n20 10.6151
R1509 B.n757 B.n20 10.6151
R1510 B.n757 B.n756 10.6151
R1511 B.n756 B.n755 10.6151
R1512 B.n755 B.n22 10.6151
R1513 B.n751 B.n22 10.6151
R1514 B.n751 B.n750 10.6151
R1515 B.n750 B.n749 10.6151
R1516 B.n749 B.n24 10.6151
R1517 B.n745 B.n24 10.6151
R1518 B.n672 B.n671 9.36635
R1519 B.n654 B.n60 9.36635
R1520 B.n353 B.n352 9.36635
R1521 B.n370 B.n157 9.36635
R1522 B.n815 B.n0 2.81026
R1523 B.n815 B.n1 2.81026
R1524 B.n671 B.n670 1.24928
R1525 B.n60 B.n56 1.24928
R1526 B.n354 B.n353 1.24928
R1527 B.n367 B.n157 1.24928
C0 VDD2 VP 0.483364f
C1 w_n3538_n3868# VDD1 2.66317f
C2 VDD2 VTAIL 12.000401f
C3 VDD1 VN 0.151803f
C4 B VDD2 2.44744f
C5 w_n3538_n3868# VP 7.82482f
C6 VP VN 7.69191f
C7 w_n3538_n3868# VTAIL 3.46958f
C8 VTAIL VN 11.9433f
C9 B w_n3538_n3868# 9.91927f
C10 B VN 1.1148f
C11 VDD1 VP 12.059099f
C12 VDD1 VTAIL 11.956599f
C13 w_n3538_n3868# VDD2 2.76576f
C14 B VDD1 2.36029f
C15 VDD2 VN 11.7321f
C16 VP VTAIL 11.957701f
C17 B VP 1.88091f
C18 B VTAIL 3.89768f
C19 w_n3538_n3868# VN 7.36662f
C20 VDD2 VDD1 1.66038f
C21 VDD2 VSUBS 1.888763f
C22 VDD1 VSUBS 1.700292f
C23 VTAIL VSUBS 1.199991f
C24 VN VSUBS 6.51086f
C25 VP VSUBS 3.307476f
C26 B VSUBS 4.5972f
C27 w_n3538_n3868# VSUBS 0.167913p
C28 B.n0 VSUBS 0.005297f
C29 B.n1 VSUBS 0.005297f
C30 B.n2 VSUBS 0.008376f
C31 B.n3 VSUBS 0.008376f
C32 B.n4 VSUBS 0.008376f
C33 B.n5 VSUBS 0.008376f
C34 B.n6 VSUBS 0.008376f
C35 B.n7 VSUBS 0.008376f
C36 B.n8 VSUBS 0.008376f
C37 B.n9 VSUBS 0.008376f
C38 B.n10 VSUBS 0.008376f
C39 B.n11 VSUBS 0.008376f
C40 B.n12 VSUBS 0.008376f
C41 B.n13 VSUBS 0.008376f
C42 B.n14 VSUBS 0.008376f
C43 B.n15 VSUBS 0.008376f
C44 B.n16 VSUBS 0.008376f
C45 B.n17 VSUBS 0.008376f
C46 B.n18 VSUBS 0.008376f
C47 B.n19 VSUBS 0.008376f
C48 B.n20 VSUBS 0.008376f
C49 B.n21 VSUBS 0.008376f
C50 B.n22 VSUBS 0.008376f
C51 B.n23 VSUBS 0.008376f
C52 B.n24 VSUBS 0.008376f
C53 B.n25 VSUBS 0.018633f
C54 B.n26 VSUBS 0.008376f
C55 B.n27 VSUBS 0.008376f
C56 B.n28 VSUBS 0.008376f
C57 B.n29 VSUBS 0.008376f
C58 B.n30 VSUBS 0.008376f
C59 B.n31 VSUBS 0.008376f
C60 B.n32 VSUBS 0.008376f
C61 B.n33 VSUBS 0.008376f
C62 B.n34 VSUBS 0.008376f
C63 B.n35 VSUBS 0.008376f
C64 B.n36 VSUBS 0.008376f
C65 B.n37 VSUBS 0.008376f
C66 B.n38 VSUBS 0.008376f
C67 B.n39 VSUBS 0.008376f
C68 B.n40 VSUBS 0.008376f
C69 B.n41 VSUBS 0.008376f
C70 B.n42 VSUBS 0.008376f
C71 B.n43 VSUBS 0.008376f
C72 B.n44 VSUBS 0.008376f
C73 B.n45 VSUBS 0.008376f
C74 B.n46 VSUBS 0.008376f
C75 B.n47 VSUBS 0.008376f
C76 B.n48 VSUBS 0.008376f
C77 B.n49 VSUBS 0.008376f
C78 B.t5 VSUBS 0.575928f
C79 B.t4 VSUBS 0.595052f
C80 B.t3 VSUBS 1.37557f
C81 B.n50 VSUBS 0.280271f
C82 B.n51 VSUBS 0.082166f
C83 B.n52 VSUBS 0.008376f
C84 B.n53 VSUBS 0.008376f
C85 B.n54 VSUBS 0.008376f
C86 B.n55 VSUBS 0.008376f
C87 B.n56 VSUBS 0.004681f
C88 B.n57 VSUBS 0.008376f
C89 B.t8 VSUBS 0.575913f
C90 B.t7 VSUBS 0.595039f
C91 B.t6 VSUBS 1.37557f
C92 B.n58 VSUBS 0.280285f
C93 B.n59 VSUBS 0.082181f
C94 B.n60 VSUBS 0.019407f
C95 B.n61 VSUBS 0.008376f
C96 B.n62 VSUBS 0.008376f
C97 B.n63 VSUBS 0.008376f
C98 B.n64 VSUBS 0.008376f
C99 B.n65 VSUBS 0.008376f
C100 B.n66 VSUBS 0.008376f
C101 B.n67 VSUBS 0.008376f
C102 B.n68 VSUBS 0.008376f
C103 B.n69 VSUBS 0.008376f
C104 B.n70 VSUBS 0.008376f
C105 B.n71 VSUBS 0.008376f
C106 B.n72 VSUBS 0.008376f
C107 B.n73 VSUBS 0.008376f
C108 B.n74 VSUBS 0.008376f
C109 B.n75 VSUBS 0.008376f
C110 B.n76 VSUBS 0.008376f
C111 B.n77 VSUBS 0.008376f
C112 B.n78 VSUBS 0.008376f
C113 B.n79 VSUBS 0.008376f
C114 B.n80 VSUBS 0.008376f
C115 B.n81 VSUBS 0.008376f
C116 B.n82 VSUBS 0.008376f
C117 B.n83 VSUBS 0.008376f
C118 B.n84 VSUBS 0.017336f
C119 B.n85 VSUBS 0.008376f
C120 B.n86 VSUBS 0.008376f
C121 B.n87 VSUBS 0.008376f
C122 B.n88 VSUBS 0.008376f
C123 B.n89 VSUBS 0.008376f
C124 B.n90 VSUBS 0.008376f
C125 B.n91 VSUBS 0.008376f
C126 B.n92 VSUBS 0.008376f
C127 B.n93 VSUBS 0.008376f
C128 B.n94 VSUBS 0.008376f
C129 B.n95 VSUBS 0.008376f
C130 B.n96 VSUBS 0.008376f
C131 B.n97 VSUBS 0.008376f
C132 B.n98 VSUBS 0.008376f
C133 B.n99 VSUBS 0.008376f
C134 B.n100 VSUBS 0.008376f
C135 B.n101 VSUBS 0.008376f
C136 B.n102 VSUBS 0.008376f
C137 B.n103 VSUBS 0.008376f
C138 B.n104 VSUBS 0.008376f
C139 B.n105 VSUBS 0.008376f
C140 B.n106 VSUBS 0.008376f
C141 B.n107 VSUBS 0.008376f
C142 B.n108 VSUBS 0.008376f
C143 B.n109 VSUBS 0.008376f
C144 B.n110 VSUBS 0.008376f
C145 B.n111 VSUBS 0.008376f
C146 B.n112 VSUBS 0.008376f
C147 B.n113 VSUBS 0.008376f
C148 B.n114 VSUBS 0.008376f
C149 B.n115 VSUBS 0.008376f
C150 B.n116 VSUBS 0.008376f
C151 B.n117 VSUBS 0.008376f
C152 B.n118 VSUBS 0.008376f
C153 B.n119 VSUBS 0.008376f
C154 B.n120 VSUBS 0.008376f
C155 B.n121 VSUBS 0.008376f
C156 B.n122 VSUBS 0.008376f
C157 B.n123 VSUBS 0.008376f
C158 B.n124 VSUBS 0.008376f
C159 B.n125 VSUBS 0.008376f
C160 B.n126 VSUBS 0.008376f
C161 B.n127 VSUBS 0.008376f
C162 B.n128 VSUBS 0.008376f
C163 B.n129 VSUBS 0.008376f
C164 B.n130 VSUBS 0.017336f
C165 B.n131 VSUBS 0.008376f
C166 B.n132 VSUBS 0.008376f
C167 B.n133 VSUBS 0.008376f
C168 B.n134 VSUBS 0.008376f
C169 B.n135 VSUBS 0.008376f
C170 B.n136 VSUBS 0.008376f
C171 B.n137 VSUBS 0.008376f
C172 B.n138 VSUBS 0.008376f
C173 B.n139 VSUBS 0.008376f
C174 B.n140 VSUBS 0.008376f
C175 B.n141 VSUBS 0.008376f
C176 B.n142 VSUBS 0.008376f
C177 B.n143 VSUBS 0.008376f
C178 B.n144 VSUBS 0.008376f
C179 B.n145 VSUBS 0.008376f
C180 B.n146 VSUBS 0.008376f
C181 B.n147 VSUBS 0.008376f
C182 B.n148 VSUBS 0.008376f
C183 B.n149 VSUBS 0.008376f
C184 B.n150 VSUBS 0.008376f
C185 B.n151 VSUBS 0.008376f
C186 B.n152 VSUBS 0.008376f
C187 B.n153 VSUBS 0.008376f
C188 B.n154 VSUBS 0.008376f
C189 B.t10 VSUBS 0.575913f
C190 B.t11 VSUBS 0.595039f
C191 B.t9 VSUBS 1.37557f
C192 B.n155 VSUBS 0.280285f
C193 B.n156 VSUBS 0.082181f
C194 B.n157 VSUBS 0.019407f
C195 B.n158 VSUBS 0.008376f
C196 B.n159 VSUBS 0.008376f
C197 B.n160 VSUBS 0.008376f
C198 B.n161 VSUBS 0.008376f
C199 B.n162 VSUBS 0.008376f
C200 B.t1 VSUBS 0.575928f
C201 B.t2 VSUBS 0.595052f
C202 B.t0 VSUBS 1.37557f
C203 B.n163 VSUBS 0.280271f
C204 B.n164 VSUBS 0.082166f
C205 B.n165 VSUBS 0.008376f
C206 B.n166 VSUBS 0.008376f
C207 B.n167 VSUBS 0.008376f
C208 B.n168 VSUBS 0.008376f
C209 B.n169 VSUBS 0.008376f
C210 B.n170 VSUBS 0.008376f
C211 B.n171 VSUBS 0.008376f
C212 B.n172 VSUBS 0.008376f
C213 B.n173 VSUBS 0.008376f
C214 B.n174 VSUBS 0.008376f
C215 B.n175 VSUBS 0.008376f
C216 B.n176 VSUBS 0.008376f
C217 B.n177 VSUBS 0.008376f
C218 B.n178 VSUBS 0.008376f
C219 B.n179 VSUBS 0.008376f
C220 B.n180 VSUBS 0.008376f
C221 B.n181 VSUBS 0.008376f
C222 B.n182 VSUBS 0.008376f
C223 B.n183 VSUBS 0.008376f
C224 B.n184 VSUBS 0.008376f
C225 B.n185 VSUBS 0.008376f
C226 B.n186 VSUBS 0.008376f
C227 B.n187 VSUBS 0.008376f
C228 B.n188 VSUBS 0.008376f
C229 B.n189 VSUBS 0.017336f
C230 B.n190 VSUBS 0.008376f
C231 B.n191 VSUBS 0.008376f
C232 B.n192 VSUBS 0.008376f
C233 B.n193 VSUBS 0.008376f
C234 B.n194 VSUBS 0.008376f
C235 B.n195 VSUBS 0.008376f
C236 B.n196 VSUBS 0.008376f
C237 B.n197 VSUBS 0.008376f
C238 B.n198 VSUBS 0.008376f
C239 B.n199 VSUBS 0.008376f
C240 B.n200 VSUBS 0.008376f
C241 B.n201 VSUBS 0.008376f
C242 B.n202 VSUBS 0.008376f
C243 B.n203 VSUBS 0.008376f
C244 B.n204 VSUBS 0.008376f
C245 B.n205 VSUBS 0.008376f
C246 B.n206 VSUBS 0.008376f
C247 B.n207 VSUBS 0.008376f
C248 B.n208 VSUBS 0.008376f
C249 B.n209 VSUBS 0.008376f
C250 B.n210 VSUBS 0.008376f
C251 B.n211 VSUBS 0.008376f
C252 B.n212 VSUBS 0.008376f
C253 B.n213 VSUBS 0.008376f
C254 B.n214 VSUBS 0.008376f
C255 B.n215 VSUBS 0.008376f
C256 B.n216 VSUBS 0.008376f
C257 B.n217 VSUBS 0.008376f
C258 B.n218 VSUBS 0.008376f
C259 B.n219 VSUBS 0.008376f
C260 B.n220 VSUBS 0.008376f
C261 B.n221 VSUBS 0.008376f
C262 B.n222 VSUBS 0.008376f
C263 B.n223 VSUBS 0.008376f
C264 B.n224 VSUBS 0.008376f
C265 B.n225 VSUBS 0.008376f
C266 B.n226 VSUBS 0.008376f
C267 B.n227 VSUBS 0.008376f
C268 B.n228 VSUBS 0.008376f
C269 B.n229 VSUBS 0.008376f
C270 B.n230 VSUBS 0.008376f
C271 B.n231 VSUBS 0.008376f
C272 B.n232 VSUBS 0.008376f
C273 B.n233 VSUBS 0.008376f
C274 B.n234 VSUBS 0.008376f
C275 B.n235 VSUBS 0.008376f
C276 B.n236 VSUBS 0.008376f
C277 B.n237 VSUBS 0.008376f
C278 B.n238 VSUBS 0.008376f
C279 B.n239 VSUBS 0.008376f
C280 B.n240 VSUBS 0.008376f
C281 B.n241 VSUBS 0.008376f
C282 B.n242 VSUBS 0.008376f
C283 B.n243 VSUBS 0.008376f
C284 B.n244 VSUBS 0.008376f
C285 B.n245 VSUBS 0.008376f
C286 B.n246 VSUBS 0.008376f
C287 B.n247 VSUBS 0.008376f
C288 B.n248 VSUBS 0.008376f
C289 B.n249 VSUBS 0.008376f
C290 B.n250 VSUBS 0.008376f
C291 B.n251 VSUBS 0.008376f
C292 B.n252 VSUBS 0.008376f
C293 B.n253 VSUBS 0.008376f
C294 B.n254 VSUBS 0.008376f
C295 B.n255 VSUBS 0.008376f
C296 B.n256 VSUBS 0.008376f
C297 B.n257 VSUBS 0.008376f
C298 B.n258 VSUBS 0.008376f
C299 B.n259 VSUBS 0.008376f
C300 B.n260 VSUBS 0.008376f
C301 B.n261 VSUBS 0.008376f
C302 B.n262 VSUBS 0.008376f
C303 B.n263 VSUBS 0.008376f
C304 B.n264 VSUBS 0.008376f
C305 B.n265 VSUBS 0.008376f
C306 B.n266 VSUBS 0.008376f
C307 B.n267 VSUBS 0.008376f
C308 B.n268 VSUBS 0.008376f
C309 B.n269 VSUBS 0.008376f
C310 B.n270 VSUBS 0.008376f
C311 B.n271 VSUBS 0.008376f
C312 B.n272 VSUBS 0.008376f
C313 B.n273 VSUBS 0.008376f
C314 B.n274 VSUBS 0.008376f
C315 B.n275 VSUBS 0.008376f
C316 B.n276 VSUBS 0.008376f
C317 B.n277 VSUBS 0.008376f
C318 B.n278 VSUBS 0.017336f
C319 B.n279 VSUBS 0.018633f
C320 B.n280 VSUBS 0.018633f
C321 B.n281 VSUBS 0.008376f
C322 B.n282 VSUBS 0.008376f
C323 B.n283 VSUBS 0.008376f
C324 B.n284 VSUBS 0.008376f
C325 B.n285 VSUBS 0.008376f
C326 B.n286 VSUBS 0.008376f
C327 B.n287 VSUBS 0.008376f
C328 B.n288 VSUBS 0.008376f
C329 B.n289 VSUBS 0.008376f
C330 B.n290 VSUBS 0.008376f
C331 B.n291 VSUBS 0.008376f
C332 B.n292 VSUBS 0.008376f
C333 B.n293 VSUBS 0.008376f
C334 B.n294 VSUBS 0.008376f
C335 B.n295 VSUBS 0.008376f
C336 B.n296 VSUBS 0.008376f
C337 B.n297 VSUBS 0.008376f
C338 B.n298 VSUBS 0.008376f
C339 B.n299 VSUBS 0.008376f
C340 B.n300 VSUBS 0.008376f
C341 B.n301 VSUBS 0.008376f
C342 B.n302 VSUBS 0.008376f
C343 B.n303 VSUBS 0.008376f
C344 B.n304 VSUBS 0.008376f
C345 B.n305 VSUBS 0.008376f
C346 B.n306 VSUBS 0.008376f
C347 B.n307 VSUBS 0.008376f
C348 B.n308 VSUBS 0.008376f
C349 B.n309 VSUBS 0.008376f
C350 B.n310 VSUBS 0.008376f
C351 B.n311 VSUBS 0.008376f
C352 B.n312 VSUBS 0.008376f
C353 B.n313 VSUBS 0.008376f
C354 B.n314 VSUBS 0.008376f
C355 B.n315 VSUBS 0.008376f
C356 B.n316 VSUBS 0.008376f
C357 B.n317 VSUBS 0.008376f
C358 B.n318 VSUBS 0.008376f
C359 B.n319 VSUBS 0.008376f
C360 B.n320 VSUBS 0.008376f
C361 B.n321 VSUBS 0.008376f
C362 B.n322 VSUBS 0.008376f
C363 B.n323 VSUBS 0.008376f
C364 B.n324 VSUBS 0.008376f
C365 B.n325 VSUBS 0.008376f
C366 B.n326 VSUBS 0.008376f
C367 B.n327 VSUBS 0.008376f
C368 B.n328 VSUBS 0.008376f
C369 B.n329 VSUBS 0.008376f
C370 B.n330 VSUBS 0.008376f
C371 B.n331 VSUBS 0.008376f
C372 B.n332 VSUBS 0.008376f
C373 B.n333 VSUBS 0.008376f
C374 B.n334 VSUBS 0.008376f
C375 B.n335 VSUBS 0.008376f
C376 B.n336 VSUBS 0.008376f
C377 B.n337 VSUBS 0.008376f
C378 B.n338 VSUBS 0.008376f
C379 B.n339 VSUBS 0.008376f
C380 B.n340 VSUBS 0.008376f
C381 B.n341 VSUBS 0.008376f
C382 B.n342 VSUBS 0.008376f
C383 B.n343 VSUBS 0.008376f
C384 B.n344 VSUBS 0.008376f
C385 B.n345 VSUBS 0.008376f
C386 B.n346 VSUBS 0.008376f
C387 B.n347 VSUBS 0.008376f
C388 B.n348 VSUBS 0.008376f
C389 B.n349 VSUBS 0.008376f
C390 B.n350 VSUBS 0.008376f
C391 B.n351 VSUBS 0.008376f
C392 B.n352 VSUBS 0.007883f
C393 B.n353 VSUBS 0.019407f
C394 B.n354 VSUBS 0.004681f
C395 B.n355 VSUBS 0.008376f
C396 B.n356 VSUBS 0.008376f
C397 B.n357 VSUBS 0.008376f
C398 B.n358 VSUBS 0.008376f
C399 B.n359 VSUBS 0.008376f
C400 B.n360 VSUBS 0.008376f
C401 B.n361 VSUBS 0.008376f
C402 B.n362 VSUBS 0.008376f
C403 B.n363 VSUBS 0.008376f
C404 B.n364 VSUBS 0.008376f
C405 B.n365 VSUBS 0.008376f
C406 B.n366 VSUBS 0.008376f
C407 B.n367 VSUBS 0.004681f
C408 B.n368 VSUBS 0.008376f
C409 B.n369 VSUBS 0.008376f
C410 B.n370 VSUBS 0.007883f
C411 B.n371 VSUBS 0.008376f
C412 B.n372 VSUBS 0.008376f
C413 B.n373 VSUBS 0.008376f
C414 B.n374 VSUBS 0.008376f
C415 B.n375 VSUBS 0.008376f
C416 B.n376 VSUBS 0.008376f
C417 B.n377 VSUBS 0.008376f
C418 B.n378 VSUBS 0.008376f
C419 B.n379 VSUBS 0.008376f
C420 B.n380 VSUBS 0.008376f
C421 B.n381 VSUBS 0.008376f
C422 B.n382 VSUBS 0.008376f
C423 B.n383 VSUBS 0.008376f
C424 B.n384 VSUBS 0.008376f
C425 B.n385 VSUBS 0.008376f
C426 B.n386 VSUBS 0.008376f
C427 B.n387 VSUBS 0.008376f
C428 B.n388 VSUBS 0.008376f
C429 B.n389 VSUBS 0.008376f
C430 B.n390 VSUBS 0.008376f
C431 B.n391 VSUBS 0.008376f
C432 B.n392 VSUBS 0.008376f
C433 B.n393 VSUBS 0.008376f
C434 B.n394 VSUBS 0.008376f
C435 B.n395 VSUBS 0.008376f
C436 B.n396 VSUBS 0.008376f
C437 B.n397 VSUBS 0.008376f
C438 B.n398 VSUBS 0.008376f
C439 B.n399 VSUBS 0.008376f
C440 B.n400 VSUBS 0.008376f
C441 B.n401 VSUBS 0.008376f
C442 B.n402 VSUBS 0.008376f
C443 B.n403 VSUBS 0.008376f
C444 B.n404 VSUBS 0.008376f
C445 B.n405 VSUBS 0.008376f
C446 B.n406 VSUBS 0.008376f
C447 B.n407 VSUBS 0.008376f
C448 B.n408 VSUBS 0.008376f
C449 B.n409 VSUBS 0.008376f
C450 B.n410 VSUBS 0.008376f
C451 B.n411 VSUBS 0.008376f
C452 B.n412 VSUBS 0.008376f
C453 B.n413 VSUBS 0.008376f
C454 B.n414 VSUBS 0.008376f
C455 B.n415 VSUBS 0.008376f
C456 B.n416 VSUBS 0.008376f
C457 B.n417 VSUBS 0.008376f
C458 B.n418 VSUBS 0.008376f
C459 B.n419 VSUBS 0.008376f
C460 B.n420 VSUBS 0.008376f
C461 B.n421 VSUBS 0.008376f
C462 B.n422 VSUBS 0.008376f
C463 B.n423 VSUBS 0.008376f
C464 B.n424 VSUBS 0.008376f
C465 B.n425 VSUBS 0.008376f
C466 B.n426 VSUBS 0.008376f
C467 B.n427 VSUBS 0.008376f
C468 B.n428 VSUBS 0.008376f
C469 B.n429 VSUBS 0.008376f
C470 B.n430 VSUBS 0.008376f
C471 B.n431 VSUBS 0.008376f
C472 B.n432 VSUBS 0.008376f
C473 B.n433 VSUBS 0.008376f
C474 B.n434 VSUBS 0.008376f
C475 B.n435 VSUBS 0.008376f
C476 B.n436 VSUBS 0.008376f
C477 B.n437 VSUBS 0.008376f
C478 B.n438 VSUBS 0.008376f
C479 B.n439 VSUBS 0.008376f
C480 B.n440 VSUBS 0.008376f
C481 B.n441 VSUBS 0.018633f
C482 B.n442 VSUBS 0.018633f
C483 B.n443 VSUBS 0.017336f
C484 B.n444 VSUBS 0.008376f
C485 B.n445 VSUBS 0.008376f
C486 B.n446 VSUBS 0.008376f
C487 B.n447 VSUBS 0.008376f
C488 B.n448 VSUBS 0.008376f
C489 B.n449 VSUBS 0.008376f
C490 B.n450 VSUBS 0.008376f
C491 B.n451 VSUBS 0.008376f
C492 B.n452 VSUBS 0.008376f
C493 B.n453 VSUBS 0.008376f
C494 B.n454 VSUBS 0.008376f
C495 B.n455 VSUBS 0.008376f
C496 B.n456 VSUBS 0.008376f
C497 B.n457 VSUBS 0.008376f
C498 B.n458 VSUBS 0.008376f
C499 B.n459 VSUBS 0.008376f
C500 B.n460 VSUBS 0.008376f
C501 B.n461 VSUBS 0.008376f
C502 B.n462 VSUBS 0.008376f
C503 B.n463 VSUBS 0.008376f
C504 B.n464 VSUBS 0.008376f
C505 B.n465 VSUBS 0.008376f
C506 B.n466 VSUBS 0.008376f
C507 B.n467 VSUBS 0.008376f
C508 B.n468 VSUBS 0.008376f
C509 B.n469 VSUBS 0.008376f
C510 B.n470 VSUBS 0.008376f
C511 B.n471 VSUBS 0.008376f
C512 B.n472 VSUBS 0.008376f
C513 B.n473 VSUBS 0.008376f
C514 B.n474 VSUBS 0.008376f
C515 B.n475 VSUBS 0.008376f
C516 B.n476 VSUBS 0.008376f
C517 B.n477 VSUBS 0.008376f
C518 B.n478 VSUBS 0.008376f
C519 B.n479 VSUBS 0.008376f
C520 B.n480 VSUBS 0.008376f
C521 B.n481 VSUBS 0.008376f
C522 B.n482 VSUBS 0.008376f
C523 B.n483 VSUBS 0.008376f
C524 B.n484 VSUBS 0.008376f
C525 B.n485 VSUBS 0.008376f
C526 B.n486 VSUBS 0.008376f
C527 B.n487 VSUBS 0.008376f
C528 B.n488 VSUBS 0.008376f
C529 B.n489 VSUBS 0.008376f
C530 B.n490 VSUBS 0.008376f
C531 B.n491 VSUBS 0.008376f
C532 B.n492 VSUBS 0.008376f
C533 B.n493 VSUBS 0.008376f
C534 B.n494 VSUBS 0.008376f
C535 B.n495 VSUBS 0.008376f
C536 B.n496 VSUBS 0.008376f
C537 B.n497 VSUBS 0.008376f
C538 B.n498 VSUBS 0.008376f
C539 B.n499 VSUBS 0.008376f
C540 B.n500 VSUBS 0.008376f
C541 B.n501 VSUBS 0.008376f
C542 B.n502 VSUBS 0.008376f
C543 B.n503 VSUBS 0.008376f
C544 B.n504 VSUBS 0.008376f
C545 B.n505 VSUBS 0.008376f
C546 B.n506 VSUBS 0.008376f
C547 B.n507 VSUBS 0.008376f
C548 B.n508 VSUBS 0.008376f
C549 B.n509 VSUBS 0.008376f
C550 B.n510 VSUBS 0.008376f
C551 B.n511 VSUBS 0.008376f
C552 B.n512 VSUBS 0.008376f
C553 B.n513 VSUBS 0.008376f
C554 B.n514 VSUBS 0.008376f
C555 B.n515 VSUBS 0.008376f
C556 B.n516 VSUBS 0.008376f
C557 B.n517 VSUBS 0.008376f
C558 B.n518 VSUBS 0.008376f
C559 B.n519 VSUBS 0.008376f
C560 B.n520 VSUBS 0.008376f
C561 B.n521 VSUBS 0.008376f
C562 B.n522 VSUBS 0.008376f
C563 B.n523 VSUBS 0.008376f
C564 B.n524 VSUBS 0.008376f
C565 B.n525 VSUBS 0.008376f
C566 B.n526 VSUBS 0.008376f
C567 B.n527 VSUBS 0.008376f
C568 B.n528 VSUBS 0.008376f
C569 B.n529 VSUBS 0.008376f
C570 B.n530 VSUBS 0.008376f
C571 B.n531 VSUBS 0.008376f
C572 B.n532 VSUBS 0.008376f
C573 B.n533 VSUBS 0.008376f
C574 B.n534 VSUBS 0.008376f
C575 B.n535 VSUBS 0.008376f
C576 B.n536 VSUBS 0.008376f
C577 B.n537 VSUBS 0.008376f
C578 B.n538 VSUBS 0.008376f
C579 B.n539 VSUBS 0.008376f
C580 B.n540 VSUBS 0.008376f
C581 B.n541 VSUBS 0.008376f
C582 B.n542 VSUBS 0.008376f
C583 B.n543 VSUBS 0.008376f
C584 B.n544 VSUBS 0.008376f
C585 B.n545 VSUBS 0.008376f
C586 B.n546 VSUBS 0.008376f
C587 B.n547 VSUBS 0.008376f
C588 B.n548 VSUBS 0.008376f
C589 B.n549 VSUBS 0.008376f
C590 B.n550 VSUBS 0.008376f
C591 B.n551 VSUBS 0.008376f
C592 B.n552 VSUBS 0.008376f
C593 B.n553 VSUBS 0.008376f
C594 B.n554 VSUBS 0.008376f
C595 B.n555 VSUBS 0.008376f
C596 B.n556 VSUBS 0.008376f
C597 B.n557 VSUBS 0.008376f
C598 B.n558 VSUBS 0.008376f
C599 B.n559 VSUBS 0.008376f
C600 B.n560 VSUBS 0.008376f
C601 B.n561 VSUBS 0.008376f
C602 B.n562 VSUBS 0.008376f
C603 B.n563 VSUBS 0.008376f
C604 B.n564 VSUBS 0.008376f
C605 B.n565 VSUBS 0.008376f
C606 B.n566 VSUBS 0.008376f
C607 B.n567 VSUBS 0.008376f
C608 B.n568 VSUBS 0.008376f
C609 B.n569 VSUBS 0.008376f
C610 B.n570 VSUBS 0.008376f
C611 B.n571 VSUBS 0.008376f
C612 B.n572 VSUBS 0.008376f
C613 B.n573 VSUBS 0.008376f
C614 B.n574 VSUBS 0.008376f
C615 B.n575 VSUBS 0.008376f
C616 B.n576 VSUBS 0.008376f
C617 B.n577 VSUBS 0.008376f
C618 B.n578 VSUBS 0.008376f
C619 B.n579 VSUBS 0.008376f
C620 B.n580 VSUBS 0.008376f
C621 B.n581 VSUBS 0.018467f
C622 B.n582 VSUBS 0.017501f
C623 B.n583 VSUBS 0.018633f
C624 B.n584 VSUBS 0.008376f
C625 B.n585 VSUBS 0.008376f
C626 B.n586 VSUBS 0.008376f
C627 B.n587 VSUBS 0.008376f
C628 B.n588 VSUBS 0.008376f
C629 B.n589 VSUBS 0.008376f
C630 B.n590 VSUBS 0.008376f
C631 B.n591 VSUBS 0.008376f
C632 B.n592 VSUBS 0.008376f
C633 B.n593 VSUBS 0.008376f
C634 B.n594 VSUBS 0.008376f
C635 B.n595 VSUBS 0.008376f
C636 B.n596 VSUBS 0.008376f
C637 B.n597 VSUBS 0.008376f
C638 B.n598 VSUBS 0.008376f
C639 B.n599 VSUBS 0.008376f
C640 B.n600 VSUBS 0.008376f
C641 B.n601 VSUBS 0.008376f
C642 B.n602 VSUBS 0.008376f
C643 B.n603 VSUBS 0.008376f
C644 B.n604 VSUBS 0.008376f
C645 B.n605 VSUBS 0.008376f
C646 B.n606 VSUBS 0.008376f
C647 B.n607 VSUBS 0.008376f
C648 B.n608 VSUBS 0.008376f
C649 B.n609 VSUBS 0.008376f
C650 B.n610 VSUBS 0.008376f
C651 B.n611 VSUBS 0.008376f
C652 B.n612 VSUBS 0.008376f
C653 B.n613 VSUBS 0.008376f
C654 B.n614 VSUBS 0.008376f
C655 B.n615 VSUBS 0.008376f
C656 B.n616 VSUBS 0.008376f
C657 B.n617 VSUBS 0.008376f
C658 B.n618 VSUBS 0.008376f
C659 B.n619 VSUBS 0.008376f
C660 B.n620 VSUBS 0.008376f
C661 B.n621 VSUBS 0.008376f
C662 B.n622 VSUBS 0.008376f
C663 B.n623 VSUBS 0.008376f
C664 B.n624 VSUBS 0.008376f
C665 B.n625 VSUBS 0.008376f
C666 B.n626 VSUBS 0.008376f
C667 B.n627 VSUBS 0.008376f
C668 B.n628 VSUBS 0.008376f
C669 B.n629 VSUBS 0.008376f
C670 B.n630 VSUBS 0.008376f
C671 B.n631 VSUBS 0.008376f
C672 B.n632 VSUBS 0.008376f
C673 B.n633 VSUBS 0.008376f
C674 B.n634 VSUBS 0.008376f
C675 B.n635 VSUBS 0.008376f
C676 B.n636 VSUBS 0.008376f
C677 B.n637 VSUBS 0.008376f
C678 B.n638 VSUBS 0.008376f
C679 B.n639 VSUBS 0.008376f
C680 B.n640 VSUBS 0.008376f
C681 B.n641 VSUBS 0.008376f
C682 B.n642 VSUBS 0.008376f
C683 B.n643 VSUBS 0.008376f
C684 B.n644 VSUBS 0.008376f
C685 B.n645 VSUBS 0.008376f
C686 B.n646 VSUBS 0.008376f
C687 B.n647 VSUBS 0.008376f
C688 B.n648 VSUBS 0.008376f
C689 B.n649 VSUBS 0.008376f
C690 B.n650 VSUBS 0.008376f
C691 B.n651 VSUBS 0.008376f
C692 B.n652 VSUBS 0.008376f
C693 B.n653 VSUBS 0.008376f
C694 B.n654 VSUBS 0.007883f
C695 B.n655 VSUBS 0.008376f
C696 B.n656 VSUBS 0.008376f
C697 B.n657 VSUBS 0.008376f
C698 B.n658 VSUBS 0.008376f
C699 B.n659 VSUBS 0.008376f
C700 B.n660 VSUBS 0.008376f
C701 B.n661 VSUBS 0.008376f
C702 B.n662 VSUBS 0.008376f
C703 B.n663 VSUBS 0.008376f
C704 B.n664 VSUBS 0.008376f
C705 B.n665 VSUBS 0.008376f
C706 B.n666 VSUBS 0.008376f
C707 B.n667 VSUBS 0.008376f
C708 B.n668 VSUBS 0.008376f
C709 B.n669 VSUBS 0.008376f
C710 B.n670 VSUBS 0.004681f
C711 B.n671 VSUBS 0.019407f
C712 B.n672 VSUBS 0.007883f
C713 B.n673 VSUBS 0.008376f
C714 B.n674 VSUBS 0.008376f
C715 B.n675 VSUBS 0.008376f
C716 B.n676 VSUBS 0.008376f
C717 B.n677 VSUBS 0.008376f
C718 B.n678 VSUBS 0.008376f
C719 B.n679 VSUBS 0.008376f
C720 B.n680 VSUBS 0.008376f
C721 B.n681 VSUBS 0.008376f
C722 B.n682 VSUBS 0.008376f
C723 B.n683 VSUBS 0.008376f
C724 B.n684 VSUBS 0.008376f
C725 B.n685 VSUBS 0.008376f
C726 B.n686 VSUBS 0.008376f
C727 B.n687 VSUBS 0.008376f
C728 B.n688 VSUBS 0.008376f
C729 B.n689 VSUBS 0.008376f
C730 B.n690 VSUBS 0.008376f
C731 B.n691 VSUBS 0.008376f
C732 B.n692 VSUBS 0.008376f
C733 B.n693 VSUBS 0.008376f
C734 B.n694 VSUBS 0.008376f
C735 B.n695 VSUBS 0.008376f
C736 B.n696 VSUBS 0.008376f
C737 B.n697 VSUBS 0.008376f
C738 B.n698 VSUBS 0.008376f
C739 B.n699 VSUBS 0.008376f
C740 B.n700 VSUBS 0.008376f
C741 B.n701 VSUBS 0.008376f
C742 B.n702 VSUBS 0.008376f
C743 B.n703 VSUBS 0.008376f
C744 B.n704 VSUBS 0.008376f
C745 B.n705 VSUBS 0.008376f
C746 B.n706 VSUBS 0.008376f
C747 B.n707 VSUBS 0.008376f
C748 B.n708 VSUBS 0.008376f
C749 B.n709 VSUBS 0.008376f
C750 B.n710 VSUBS 0.008376f
C751 B.n711 VSUBS 0.008376f
C752 B.n712 VSUBS 0.008376f
C753 B.n713 VSUBS 0.008376f
C754 B.n714 VSUBS 0.008376f
C755 B.n715 VSUBS 0.008376f
C756 B.n716 VSUBS 0.008376f
C757 B.n717 VSUBS 0.008376f
C758 B.n718 VSUBS 0.008376f
C759 B.n719 VSUBS 0.008376f
C760 B.n720 VSUBS 0.008376f
C761 B.n721 VSUBS 0.008376f
C762 B.n722 VSUBS 0.008376f
C763 B.n723 VSUBS 0.008376f
C764 B.n724 VSUBS 0.008376f
C765 B.n725 VSUBS 0.008376f
C766 B.n726 VSUBS 0.008376f
C767 B.n727 VSUBS 0.008376f
C768 B.n728 VSUBS 0.008376f
C769 B.n729 VSUBS 0.008376f
C770 B.n730 VSUBS 0.008376f
C771 B.n731 VSUBS 0.008376f
C772 B.n732 VSUBS 0.008376f
C773 B.n733 VSUBS 0.008376f
C774 B.n734 VSUBS 0.008376f
C775 B.n735 VSUBS 0.008376f
C776 B.n736 VSUBS 0.008376f
C777 B.n737 VSUBS 0.008376f
C778 B.n738 VSUBS 0.008376f
C779 B.n739 VSUBS 0.008376f
C780 B.n740 VSUBS 0.008376f
C781 B.n741 VSUBS 0.008376f
C782 B.n742 VSUBS 0.008376f
C783 B.n743 VSUBS 0.008376f
C784 B.n744 VSUBS 0.018633f
C785 B.n745 VSUBS 0.017336f
C786 B.n746 VSUBS 0.017336f
C787 B.n747 VSUBS 0.008376f
C788 B.n748 VSUBS 0.008376f
C789 B.n749 VSUBS 0.008376f
C790 B.n750 VSUBS 0.008376f
C791 B.n751 VSUBS 0.008376f
C792 B.n752 VSUBS 0.008376f
C793 B.n753 VSUBS 0.008376f
C794 B.n754 VSUBS 0.008376f
C795 B.n755 VSUBS 0.008376f
C796 B.n756 VSUBS 0.008376f
C797 B.n757 VSUBS 0.008376f
C798 B.n758 VSUBS 0.008376f
C799 B.n759 VSUBS 0.008376f
C800 B.n760 VSUBS 0.008376f
C801 B.n761 VSUBS 0.008376f
C802 B.n762 VSUBS 0.008376f
C803 B.n763 VSUBS 0.008376f
C804 B.n764 VSUBS 0.008376f
C805 B.n765 VSUBS 0.008376f
C806 B.n766 VSUBS 0.008376f
C807 B.n767 VSUBS 0.008376f
C808 B.n768 VSUBS 0.008376f
C809 B.n769 VSUBS 0.008376f
C810 B.n770 VSUBS 0.008376f
C811 B.n771 VSUBS 0.008376f
C812 B.n772 VSUBS 0.008376f
C813 B.n773 VSUBS 0.008376f
C814 B.n774 VSUBS 0.008376f
C815 B.n775 VSUBS 0.008376f
C816 B.n776 VSUBS 0.008376f
C817 B.n777 VSUBS 0.008376f
C818 B.n778 VSUBS 0.008376f
C819 B.n779 VSUBS 0.008376f
C820 B.n780 VSUBS 0.008376f
C821 B.n781 VSUBS 0.008376f
C822 B.n782 VSUBS 0.008376f
C823 B.n783 VSUBS 0.008376f
C824 B.n784 VSUBS 0.008376f
C825 B.n785 VSUBS 0.008376f
C826 B.n786 VSUBS 0.008376f
C827 B.n787 VSUBS 0.008376f
C828 B.n788 VSUBS 0.008376f
C829 B.n789 VSUBS 0.008376f
C830 B.n790 VSUBS 0.008376f
C831 B.n791 VSUBS 0.008376f
C832 B.n792 VSUBS 0.008376f
C833 B.n793 VSUBS 0.008376f
C834 B.n794 VSUBS 0.008376f
C835 B.n795 VSUBS 0.008376f
C836 B.n796 VSUBS 0.008376f
C837 B.n797 VSUBS 0.008376f
C838 B.n798 VSUBS 0.008376f
C839 B.n799 VSUBS 0.008376f
C840 B.n800 VSUBS 0.008376f
C841 B.n801 VSUBS 0.008376f
C842 B.n802 VSUBS 0.008376f
C843 B.n803 VSUBS 0.008376f
C844 B.n804 VSUBS 0.008376f
C845 B.n805 VSUBS 0.008376f
C846 B.n806 VSUBS 0.008376f
C847 B.n807 VSUBS 0.008376f
C848 B.n808 VSUBS 0.008376f
C849 B.n809 VSUBS 0.008376f
C850 B.n810 VSUBS 0.008376f
C851 B.n811 VSUBS 0.008376f
C852 B.n812 VSUBS 0.008376f
C853 B.n813 VSUBS 0.008376f
C854 B.n814 VSUBS 0.008376f
C855 B.n815 VSUBS 0.018966f
C856 VDD1.t3 VSUBS 3.31521f
C857 VDD1.t8 VSUBS 0.311923f
C858 VDD1.t0 VSUBS 0.311923f
C859 VDD1.n0 VSUBS 2.53564f
C860 VDD1.n1 VSUBS 1.45455f
C861 VDD1.t2 VSUBS 3.3152f
C862 VDD1.t9 VSUBS 0.311923f
C863 VDD1.t5 VSUBS 0.311923f
C864 VDD1.n2 VSUBS 2.53564f
C865 VDD1.n3 VSUBS 1.44616f
C866 VDD1.t1 VSUBS 0.311923f
C867 VDD1.t7 VSUBS 0.311923f
C868 VDD1.n4 VSUBS 2.54936f
C869 VDD1.n5 VSUBS 3.27071f
C870 VDD1.t4 VSUBS 0.311923f
C871 VDD1.t6 VSUBS 0.311923f
C872 VDD1.n6 VSUBS 2.53563f
C873 VDD1.n7 VSUBS 3.58468f
C874 VP.n0 VSUBS 0.033445f
C875 VP.t2 VSUBS 2.40332f
C876 VP.n1 VSUBS 0.0277f
C877 VP.n2 VSUBS 0.033445f
C878 VP.t8 VSUBS 2.40332f
C879 VP.n3 VSUBS 0.04214f
C880 VP.n4 VSUBS 0.033445f
C881 VP.t4 VSUBS 2.40332f
C882 VP.n5 VSUBS 0.055094f
C883 VP.n6 VSUBS 0.033445f
C884 VP.t0 VSUBS 2.40332f
C885 VP.n7 VSUBS 0.064482f
C886 VP.n8 VSUBS 0.033445f
C887 VP.t7 VSUBS 2.40332f
C888 VP.n9 VSUBS 0.923029f
C889 VP.n10 VSUBS 0.033445f
C890 VP.t3 VSUBS 2.40332f
C891 VP.n11 VSUBS 0.0277f
C892 VP.n12 VSUBS 0.033445f
C893 VP.t5 VSUBS 2.40332f
C894 VP.n13 VSUBS 0.04214f
C895 VP.n14 VSUBS 0.033445f
C896 VP.t9 VSUBS 2.40332f
C897 VP.n15 VSUBS 0.055094f
C898 VP.n16 VSUBS 0.245428f
C899 VP.t1 VSUBS 2.40332f
C900 VP.t6 VSUBS 2.55029f
C901 VP.n17 VSUBS 0.930478f
C902 VP.n18 VSUBS 0.933479f
C903 VP.n19 VSUBS 0.055284f
C904 VP.n20 VSUBS 0.04214f
C905 VP.n21 VSUBS 0.033445f
C906 VP.n22 VSUBS 0.033445f
C907 VP.n23 VSUBS 0.033445f
C908 VP.n24 VSUBS 0.046711f
C909 VP.n25 VSUBS 0.850573f
C910 VP.n26 VSUBS 0.046711f
C911 VP.n27 VSUBS 0.055094f
C912 VP.n28 VSUBS 0.033445f
C913 VP.n29 VSUBS 0.033445f
C914 VP.n30 VSUBS 0.033445f
C915 VP.n31 VSUBS 0.055284f
C916 VP.n32 VSUBS 0.850573f
C917 VP.n33 VSUBS 0.038138f
C918 VP.n34 VSUBS 0.064482f
C919 VP.n35 VSUBS 0.033445f
C920 VP.n36 VSUBS 0.033445f
C921 VP.n37 VSUBS 0.033445f
C922 VP.n38 VSUBS 0.067071f
C923 VP.n39 VSUBS 0.033239f
C924 VP.n40 VSUBS 0.923029f
C925 VP.n41 VSUBS 1.86054f
C926 VP.n42 VSUBS 1.88437f
C927 VP.n43 VSUBS 0.033445f
C928 VP.n44 VSUBS 0.033239f
C929 VP.n45 VSUBS 0.067071f
C930 VP.n46 VSUBS 0.0277f
C931 VP.n47 VSUBS 0.033445f
C932 VP.n48 VSUBS 0.033445f
C933 VP.n49 VSUBS 0.033445f
C934 VP.n50 VSUBS 0.038138f
C935 VP.n51 VSUBS 0.850573f
C936 VP.n52 VSUBS 0.055284f
C937 VP.n53 VSUBS 0.04214f
C938 VP.n54 VSUBS 0.033445f
C939 VP.n55 VSUBS 0.033445f
C940 VP.n56 VSUBS 0.033445f
C941 VP.n57 VSUBS 0.046711f
C942 VP.n58 VSUBS 0.850573f
C943 VP.n59 VSUBS 0.046711f
C944 VP.n60 VSUBS 0.055094f
C945 VP.n61 VSUBS 0.033445f
C946 VP.n62 VSUBS 0.033445f
C947 VP.n63 VSUBS 0.033445f
C948 VP.n64 VSUBS 0.055284f
C949 VP.n65 VSUBS 0.850573f
C950 VP.n66 VSUBS 0.038138f
C951 VP.n67 VSUBS 0.064482f
C952 VP.n68 VSUBS 0.033445f
C953 VP.n69 VSUBS 0.033445f
C954 VP.n70 VSUBS 0.033445f
C955 VP.n71 VSUBS 0.067071f
C956 VP.n72 VSUBS 0.033239f
C957 VP.n73 VSUBS 0.923029f
C958 VP.n74 VSUBS 0.036302f
C959 VTAIL.t16 VSUBS 0.317608f
C960 VTAIL.t10 VSUBS 0.317608f
C961 VTAIL.n0 VSUBS 2.43805f
C962 VTAIL.n1 VSUBS 0.870018f
C963 VTAIL.t8 VSUBS 3.19425f
C964 VTAIL.n2 VSUBS 1.01601f
C965 VTAIL.t7 VSUBS 0.317608f
C966 VTAIL.t4 VSUBS 0.317608f
C967 VTAIL.n3 VSUBS 2.43805f
C968 VTAIL.n4 VSUBS 0.946436f
C969 VTAIL.t0 VSUBS 0.317608f
C970 VTAIL.t9 VSUBS 0.317608f
C971 VTAIL.n5 VSUBS 2.43805f
C972 VTAIL.n6 VSUBS 2.60417f
C973 VTAIL.t15 VSUBS 0.317608f
C974 VTAIL.t12 VSUBS 0.317608f
C975 VTAIL.n7 VSUBS 2.43805f
C976 VTAIL.n8 VSUBS 2.60416f
C977 VTAIL.t13 VSUBS 0.317608f
C978 VTAIL.t19 VSUBS 0.317608f
C979 VTAIL.n9 VSUBS 2.43805f
C980 VTAIL.n10 VSUBS 0.946431f
C981 VTAIL.t17 VSUBS 3.19427f
C982 VTAIL.n11 VSUBS 1.01599f
C983 VTAIL.t5 VSUBS 0.317608f
C984 VTAIL.t6 VSUBS 0.317608f
C985 VTAIL.n12 VSUBS 2.43805f
C986 VTAIL.n13 VSUBS 0.906009f
C987 VTAIL.t1 VSUBS 0.317608f
C988 VTAIL.t2 VSUBS 0.317608f
C989 VTAIL.n14 VSUBS 2.43805f
C990 VTAIL.n15 VSUBS 0.946431f
C991 VTAIL.t3 VSUBS 3.19425f
C992 VTAIL.n16 VSUBS 2.5494f
C993 VTAIL.t11 VSUBS 3.19425f
C994 VTAIL.n17 VSUBS 2.5494f
C995 VTAIL.t14 VSUBS 0.317608f
C996 VTAIL.t18 VSUBS 0.317608f
C997 VTAIL.n18 VSUBS 2.43805f
C998 VTAIL.n19 VSUBS 0.81766f
C999 VDD2.t4 VSUBS 3.29247f
C1000 VDD2.t7 VSUBS 0.309785f
C1001 VDD2.t5 VSUBS 0.309785f
C1002 VDD2.n0 VSUBS 2.51826f
C1003 VDD2.n1 VSUBS 1.43625f
C1004 VDD2.t9 VSUBS 0.309785f
C1005 VDD2.t2 VSUBS 0.309785f
C1006 VDD2.n2 VSUBS 2.53188f
C1007 VDD2.n3 VSUBS 3.13406f
C1008 VDD2.t8 VSUBS 3.27488f
C1009 VDD2.n4 VSUBS 3.54727f
C1010 VDD2.t6 VSUBS 0.309785f
C1011 VDD2.t0 VSUBS 0.309785f
C1012 VDD2.n5 VSUBS 2.51826f
C1013 VDD2.n6 VSUBS 0.704147f
C1014 VDD2.t1 VSUBS 0.309785f
C1015 VDD2.t3 VSUBS 0.309785f
C1016 VDD2.n7 VSUBS 2.53183f
C1017 VN.n0 VSUBS 0.032646f
C1018 VN.t8 VSUBS 2.34591f
C1019 VN.n1 VSUBS 0.027039f
C1020 VN.n2 VSUBS 0.032646f
C1021 VN.t1 VSUBS 2.34591f
C1022 VN.n3 VSUBS 0.041133f
C1023 VN.n4 VSUBS 0.032646f
C1024 VN.t5 VSUBS 2.34591f
C1025 VN.n5 VSUBS 0.053778f
C1026 VN.n6 VSUBS 0.239566f
C1027 VN.t9 VSUBS 2.34591f
C1028 VN.t3 VSUBS 2.48937f
C1029 VN.n7 VSUBS 0.908253f
C1030 VN.n8 VSUBS 0.911181f
C1031 VN.n9 VSUBS 0.053963f
C1032 VN.n10 VSUBS 0.041133f
C1033 VN.n11 VSUBS 0.032646f
C1034 VN.n12 VSUBS 0.032646f
C1035 VN.n13 VSUBS 0.032646f
C1036 VN.n14 VSUBS 0.045595f
C1037 VN.n15 VSUBS 0.830256f
C1038 VN.n16 VSUBS 0.045595f
C1039 VN.n17 VSUBS 0.053778f
C1040 VN.n18 VSUBS 0.032646f
C1041 VN.n19 VSUBS 0.032646f
C1042 VN.n20 VSUBS 0.032646f
C1043 VN.n21 VSUBS 0.053963f
C1044 VN.n22 VSUBS 0.830256f
C1045 VN.n23 VSUBS 0.037227f
C1046 VN.n24 VSUBS 0.062942f
C1047 VN.n25 VSUBS 0.032646f
C1048 VN.n26 VSUBS 0.032646f
C1049 VN.n27 VSUBS 0.032646f
C1050 VN.n28 VSUBS 0.065469f
C1051 VN.n29 VSUBS 0.032445f
C1052 VN.n30 VSUBS 0.900981f
C1053 VN.n31 VSUBS 0.035435f
C1054 VN.n32 VSUBS 0.032646f
C1055 VN.t4 VSUBS 2.34591f
C1056 VN.n33 VSUBS 0.027039f
C1057 VN.n34 VSUBS 0.032646f
C1058 VN.t7 VSUBS 2.34591f
C1059 VN.n35 VSUBS 0.041133f
C1060 VN.n36 VSUBS 0.032646f
C1061 VN.t6 VSUBS 2.34591f
C1062 VN.n37 VSUBS 0.053778f
C1063 VN.n38 VSUBS 0.239566f
C1064 VN.t0 VSUBS 2.34591f
C1065 VN.t2 VSUBS 2.48937f
C1066 VN.n39 VSUBS 0.908253f
C1067 VN.n40 VSUBS 0.911181f
C1068 VN.n41 VSUBS 0.053963f
C1069 VN.n42 VSUBS 0.041133f
C1070 VN.n43 VSUBS 0.032646f
C1071 VN.n44 VSUBS 0.032646f
C1072 VN.n45 VSUBS 0.032646f
C1073 VN.n46 VSUBS 0.045595f
C1074 VN.n47 VSUBS 0.830256f
C1075 VN.n48 VSUBS 0.045595f
C1076 VN.n49 VSUBS 0.053778f
C1077 VN.n50 VSUBS 0.032646f
C1078 VN.n51 VSUBS 0.032646f
C1079 VN.n52 VSUBS 0.032646f
C1080 VN.n53 VSUBS 0.053963f
C1081 VN.n54 VSUBS 0.830256f
C1082 VN.n55 VSUBS 0.037227f
C1083 VN.n56 VSUBS 0.062942f
C1084 VN.n57 VSUBS 0.032646f
C1085 VN.n58 VSUBS 0.032646f
C1086 VN.n59 VSUBS 0.032646f
C1087 VN.n60 VSUBS 0.065469f
C1088 VN.n61 VSUBS 0.032445f
C1089 VN.n62 VSUBS 0.900981f
C1090 VN.n63 VSUBS 1.83731f
.ends

