* NGSPICE file created from diff_pair_sample_0715.ext - technology: sky130A

.subckt diff_pair_sample_0715 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=1.14
X1 VTAIL.t7 VN.t0 VDD2.t2 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=1.14
X2 B.t8 B.t6 B.t7 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=1.14
X3 B.t5 B.t3 B.t4 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=1.14
X4 B.t2 B.t0 B.t1 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0 ps=0 w=3.95 l=1.14
X5 VDD2.t1 VN.t1 VTAIL.t6 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=1.14
X6 VTAIL.t5 VN.t2 VDD2.t3 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=1.14
X7 VDD2.t0 VN.t3 VTAIL.t4 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=1.14
X8 VTAIL.t3 VP.t0 VDD1.t3 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=1.14
X9 VTAIL.t2 VP.t1 VDD1.t2 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=1.5405 pd=8.68 as=0.65175 ps=4.28 w=3.95 l=1.14
X10 VDD1.t1 VP.t2 VTAIL.t0 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=1.14
X11 VDD1.t0 VP.t3 VTAIL.t1 w_n1852_n1758# sky130_fd_pr__pfet_01v8 ad=0.65175 pd=4.28 as=1.5405 ps=8.68 w=3.95 l=1.14
R0 B.n262 B.n39 585
R1 B.n264 B.n263 585
R2 B.n265 B.n38 585
R3 B.n267 B.n266 585
R4 B.n268 B.n37 585
R5 B.n270 B.n269 585
R6 B.n271 B.n36 585
R7 B.n273 B.n272 585
R8 B.n274 B.n35 585
R9 B.n276 B.n275 585
R10 B.n277 B.n34 585
R11 B.n279 B.n278 585
R12 B.n280 B.n33 585
R13 B.n282 B.n281 585
R14 B.n283 B.n32 585
R15 B.n285 B.n284 585
R16 B.n286 B.n31 585
R17 B.n288 B.n287 585
R18 B.n290 B.n289 585
R19 B.n291 B.n27 585
R20 B.n293 B.n292 585
R21 B.n294 B.n26 585
R22 B.n296 B.n295 585
R23 B.n297 B.n25 585
R24 B.n299 B.n298 585
R25 B.n300 B.n24 585
R26 B.n302 B.n301 585
R27 B.n304 B.n21 585
R28 B.n306 B.n305 585
R29 B.n307 B.n20 585
R30 B.n309 B.n308 585
R31 B.n310 B.n19 585
R32 B.n312 B.n311 585
R33 B.n313 B.n18 585
R34 B.n315 B.n314 585
R35 B.n316 B.n17 585
R36 B.n318 B.n317 585
R37 B.n319 B.n16 585
R38 B.n321 B.n320 585
R39 B.n322 B.n15 585
R40 B.n324 B.n323 585
R41 B.n325 B.n14 585
R42 B.n327 B.n326 585
R43 B.n328 B.n13 585
R44 B.n330 B.n329 585
R45 B.n261 B.n260 585
R46 B.n259 B.n40 585
R47 B.n258 B.n257 585
R48 B.n256 B.n41 585
R49 B.n255 B.n254 585
R50 B.n253 B.n42 585
R51 B.n252 B.n251 585
R52 B.n250 B.n43 585
R53 B.n249 B.n248 585
R54 B.n247 B.n44 585
R55 B.n246 B.n245 585
R56 B.n244 B.n45 585
R57 B.n243 B.n242 585
R58 B.n241 B.n46 585
R59 B.n240 B.n239 585
R60 B.n238 B.n47 585
R61 B.n237 B.n236 585
R62 B.n235 B.n48 585
R63 B.n234 B.n233 585
R64 B.n232 B.n49 585
R65 B.n231 B.n230 585
R66 B.n229 B.n50 585
R67 B.n228 B.n227 585
R68 B.n226 B.n51 585
R69 B.n225 B.n224 585
R70 B.n223 B.n52 585
R71 B.n222 B.n221 585
R72 B.n220 B.n53 585
R73 B.n219 B.n218 585
R74 B.n217 B.n54 585
R75 B.n216 B.n215 585
R76 B.n214 B.n55 585
R77 B.n213 B.n212 585
R78 B.n211 B.n56 585
R79 B.n210 B.n209 585
R80 B.n208 B.n57 585
R81 B.n207 B.n206 585
R82 B.n205 B.n58 585
R83 B.n204 B.n203 585
R84 B.n202 B.n59 585
R85 B.n201 B.n200 585
R86 B.n199 B.n60 585
R87 B.n198 B.n197 585
R88 B.n129 B.n128 585
R89 B.n130 B.n87 585
R90 B.n132 B.n131 585
R91 B.n133 B.n86 585
R92 B.n135 B.n134 585
R93 B.n136 B.n85 585
R94 B.n138 B.n137 585
R95 B.n139 B.n84 585
R96 B.n141 B.n140 585
R97 B.n142 B.n83 585
R98 B.n144 B.n143 585
R99 B.n145 B.n82 585
R100 B.n147 B.n146 585
R101 B.n148 B.n81 585
R102 B.n150 B.n149 585
R103 B.n151 B.n80 585
R104 B.n153 B.n152 585
R105 B.n154 B.n77 585
R106 B.n157 B.n156 585
R107 B.n158 B.n76 585
R108 B.n160 B.n159 585
R109 B.n161 B.n75 585
R110 B.n163 B.n162 585
R111 B.n164 B.n74 585
R112 B.n166 B.n165 585
R113 B.n167 B.n73 585
R114 B.n169 B.n168 585
R115 B.n171 B.n170 585
R116 B.n172 B.n69 585
R117 B.n174 B.n173 585
R118 B.n175 B.n68 585
R119 B.n177 B.n176 585
R120 B.n178 B.n67 585
R121 B.n180 B.n179 585
R122 B.n181 B.n66 585
R123 B.n183 B.n182 585
R124 B.n184 B.n65 585
R125 B.n186 B.n185 585
R126 B.n187 B.n64 585
R127 B.n189 B.n188 585
R128 B.n190 B.n63 585
R129 B.n192 B.n191 585
R130 B.n193 B.n62 585
R131 B.n195 B.n194 585
R132 B.n196 B.n61 585
R133 B.n127 B.n88 585
R134 B.n126 B.n125 585
R135 B.n124 B.n89 585
R136 B.n123 B.n122 585
R137 B.n121 B.n90 585
R138 B.n120 B.n119 585
R139 B.n118 B.n91 585
R140 B.n117 B.n116 585
R141 B.n115 B.n92 585
R142 B.n114 B.n113 585
R143 B.n112 B.n93 585
R144 B.n111 B.n110 585
R145 B.n109 B.n94 585
R146 B.n108 B.n107 585
R147 B.n106 B.n95 585
R148 B.n105 B.n104 585
R149 B.n103 B.n96 585
R150 B.n102 B.n101 585
R151 B.n100 B.n97 585
R152 B.n99 B.n98 585
R153 B.n2 B.n0 585
R154 B.n361 B.n1 585
R155 B.n360 B.n359 585
R156 B.n358 B.n3 585
R157 B.n357 B.n356 585
R158 B.n355 B.n4 585
R159 B.n354 B.n353 585
R160 B.n352 B.n5 585
R161 B.n351 B.n350 585
R162 B.n349 B.n6 585
R163 B.n348 B.n347 585
R164 B.n346 B.n7 585
R165 B.n345 B.n344 585
R166 B.n343 B.n8 585
R167 B.n342 B.n341 585
R168 B.n340 B.n9 585
R169 B.n339 B.n338 585
R170 B.n337 B.n10 585
R171 B.n336 B.n335 585
R172 B.n334 B.n11 585
R173 B.n333 B.n332 585
R174 B.n331 B.n12 585
R175 B.n363 B.n362 585
R176 B.n128 B.n127 550.159
R177 B.n331 B.n330 550.159
R178 B.n198 B.n61 550.159
R179 B.n260 B.n39 550.159
R180 B.n70 B.t0 287.296
R181 B.n78 B.t9 287.296
R182 B.n22 B.t6 287.296
R183 B.n28 B.t3 287.296
R184 B.n70 B.t2 263.168
R185 B.n28 B.t4 263.168
R186 B.n78 B.t11 263.168
R187 B.n22 B.t7 263.168
R188 B.n71 B.t1 234.66
R189 B.n29 B.t5 234.66
R190 B.n79 B.t10 234.66
R191 B.n23 B.t8 234.66
R192 B.n127 B.n126 163.367
R193 B.n126 B.n89 163.367
R194 B.n122 B.n89 163.367
R195 B.n122 B.n121 163.367
R196 B.n121 B.n120 163.367
R197 B.n120 B.n91 163.367
R198 B.n116 B.n91 163.367
R199 B.n116 B.n115 163.367
R200 B.n115 B.n114 163.367
R201 B.n114 B.n93 163.367
R202 B.n110 B.n93 163.367
R203 B.n110 B.n109 163.367
R204 B.n109 B.n108 163.367
R205 B.n108 B.n95 163.367
R206 B.n104 B.n95 163.367
R207 B.n104 B.n103 163.367
R208 B.n103 B.n102 163.367
R209 B.n102 B.n97 163.367
R210 B.n98 B.n97 163.367
R211 B.n98 B.n2 163.367
R212 B.n362 B.n2 163.367
R213 B.n362 B.n361 163.367
R214 B.n361 B.n360 163.367
R215 B.n360 B.n3 163.367
R216 B.n356 B.n3 163.367
R217 B.n356 B.n355 163.367
R218 B.n355 B.n354 163.367
R219 B.n354 B.n5 163.367
R220 B.n350 B.n5 163.367
R221 B.n350 B.n349 163.367
R222 B.n349 B.n348 163.367
R223 B.n348 B.n7 163.367
R224 B.n344 B.n7 163.367
R225 B.n344 B.n343 163.367
R226 B.n343 B.n342 163.367
R227 B.n342 B.n9 163.367
R228 B.n338 B.n9 163.367
R229 B.n338 B.n337 163.367
R230 B.n337 B.n336 163.367
R231 B.n336 B.n11 163.367
R232 B.n332 B.n11 163.367
R233 B.n332 B.n331 163.367
R234 B.n128 B.n87 163.367
R235 B.n132 B.n87 163.367
R236 B.n133 B.n132 163.367
R237 B.n134 B.n133 163.367
R238 B.n134 B.n85 163.367
R239 B.n138 B.n85 163.367
R240 B.n139 B.n138 163.367
R241 B.n140 B.n139 163.367
R242 B.n140 B.n83 163.367
R243 B.n144 B.n83 163.367
R244 B.n145 B.n144 163.367
R245 B.n146 B.n145 163.367
R246 B.n146 B.n81 163.367
R247 B.n150 B.n81 163.367
R248 B.n151 B.n150 163.367
R249 B.n152 B.n151 163.367
R250 B.n152 B.n77 163.367
R251 B.n157 B.n77 163.367
R252 B.n158 B.n157 163.367
R253 B.n159 B.n158 163.367
R254 B.n159 B.n75 163.367
R255 B.n163 B.n75 163.367
R256 B.n164 B.n163 163.367
R257 B.n165 B.n164 163.367
R258 B.n165 B.n73 163.367
R259 B.n169 B.n73 163.367
R260 B.n170 B.n169 163.367
R261 B.n170 B.n69 163.367
R262 B.n174 B.n69 163.367
R263 B.n175 B.n174 163.367
R264 B.n176 B.n175 163.367
R265 B.n176 B.n67 163.367
R266 B.n180 B.n67 163.367
R267 B.n181 B.n180 163.367
R268 B.n182 B.n181 163.367
R269 B.n182 B.n65 163.367
R270 B.n186 B.n65 163.367
R271 B.n187 B.n186 163.367
R272 B.n188 B.n187 163.367
R273 B.n188 B.n63 163.367
R274 B.n192 B.n63 163.367
R275 B.n193 B.n192 163.367
R276 B.n194 B.n193 163.367
R277 B.n194 B.n61 163.367
R278 B.n199 B.n198 163.367
R279 B.n200 B.n199 163.367
R280 B.n200 B.n59 163.367
R281 B.n204 B.n59 163.367
R282 B.n205 B.n204 163.367
R283 B.n206 B.n205 163.367
R284 B.n206 B.n57 163.367
R285 B.n210 B.n57 163.367
R286 B.n211 B.n210 163.367
R287 B.n212 B.n211 163.367
R288 B.n212 B.n55 163.367
R289 B.n216 B.n55 163.367
R290 B.n217 B.n216 163.367
R291 B.n218 B.n217 163.367
R292 B.n218 B.n53 163.367
R293 B.n222 B.n53 163.367
R294 B.n223 B.n222 163.367
R295 B.n224 B.n223 163.367
R296 B.n224 B.n51 163.367
R297 B.n228 B.n51 163.367
R298 B.n229 B.n228 163.367
R299 B.n230 B.n229 163.367
R300 B.n230 B.n49 163.367
R301 B.n234 B.n49 163.367
R302 B.n235 B.n234 163.367
R303 B.n236 B.n235 163.367
R304 B.n236 B.n47 163.367
R305 B.n240 B.n47 163.367
R306 B.n241 B.n240 163.367
R307 B.n242 B.n241 163.367
R308 B.n242 B.n45 163.367
R309 B.n246 B.n45 163.367
R310 B.n247 B.n246 163.367
R311 B.n248 B.n247 163.367
R312 B.n248 B.n43 163.367
R313 B.n252 B.n43 163.367
R314 B.n253 B.n252 163.367
R315 B.n254 B.n253 163.367
R316 B.n254 B.n41 163.367
R317 B.n258 B.n41 163.367
R318 B.n259 B.n258 163.367
R319 B.n260 B.n259 163.367
R320 B.n330 B.n13 163.367
R321 B.n326 B.n13 163.367
R322 B.n326 B.n325 163.367
R323 B.n325 B.n324 163.367
R324 B.n324 B.n15 163.367
R325 B.n320 B.n15 163.367
R326 B.n320 B.n319 163.367
R327 B.n319 B.n318 163.367
R328 B.n318 B.n17 163.367
R329 B.n314 B.n17 163.367
R330 B.n314 B.n313 163.367
R331 B.n313 B.n312 163.367
R332 B.n312 B.n19 163.367
R333 B.n308 B.n19 163.367
R334 B.n308 B.n307 163.367
R335 B.n307 B.n306 163.367
R336 B.n306 B.n21 163.367
R337 B.n301 B.n21 163.367
R338 B.n301 B.n300 163.367
R339 B.n300 B.n299 163.367
R340 B.n299 B.n25 163.367
R341 B.n295 B.n25 163.367
R342 B.n295 B.n294 163.367
R343 B.n294 B.n293 163.367
R344 B.n293 B.n27 163.367
R345 B.n289 B.n27 163.367
R346 B.n289 B.n288 163.367
R347 B.n288 B.n31 163.367
R348 B.n284 B.n31 163.367
R349 B.n284 B.n283 163.367
R350 B.n283 B.n282 163.367
R351 B.n282 B.n33 163.367
R352 B.n278 B.n33 163.367
R353 B.n278 B.n277 163.367
R354 B.n277 B.n276 163.367
R355 B.n276 B.n35 163.367
R356 B.n272 B.n35 163.367
R357 B.n272 B.n271 163.367
R358 B.n271 B.n270 163.367
R359 B.n270 B.n37 163.367
R360 B.n266 B.n37 163.367
R361 B.n266 B.n265 163.367
R362 B.n265 B.n264 163.367
R363 B.n264 B.n39 163.367
R364 B.n72 B.n71 59.5399
R365 B.n155 B.n79 59.5399
R366 B.n303 B.n23 59.5399
R367 B.n30 B.n29 59.5399
R368 B.n329 B.n12 35.7468
R369 B.n197 B.n196 35.7468
R370 B.n129 B.n88 35.7468
R371 B.n262 B.n261 35.7468
R372 B.n71 B.n70 28.5096
R373 B.n79 B.n78 28.5096
R374 B.n23 B.n22 28.5096
R375 B.n29 B.n28 28.5096
R376 B B.n363 18.0485
R377 B.n329 B.n328 10.6151
R378 B.n328 B.n327 10.6151
R379 B.n327 B.n14 10.6151
R380 B.n323 B.n14 10.6151
R381 B.n323 B.n322 10.6151
R382 B.n322 B.n321 10.6151
R383 B.n321 B.n16 10.6151
R384 B.n317 B.n16 10.6151
R385 B.n317 B.n316 10.6151
R386 B.n316 B.n315 10.6151
R387 B.n315 B.n18 10.6151
R388 B.n311 B.n18 10.6151
R389 B.n311 B.n310 10.6151
R390 B.n310 B.n309 10.6151
R391 B.n309 B.n20 10.6151
R392 B.n305 B.n20 10.6151
R393 B.n305 B.n304 10.6151
R394 B.n302 B.n24 10.6151
R395 B.n298 B.n24 10.6151
R396 B.n298 B.n297 10.6151
R397 B.n297 B.n296 10.6151
R398 B.n296 B.n26 10.6151
R399 B.n292 B.n26 10.6151
R400 B.n292 B.n291 10.6151
R401 B.n291 B.n290 10.6151
R402 B.n287 B.n286 10.6151
R403 B.n286 B.n285 10.6151
R404 B.n285 B.n32 10.6151
R405 B.n281 B.n32 10.6151
R406 B.n281 B.n280 10.6151
R407 B.n280 B.n279 10.6151
R408 B.n279 B.n34 10.6151
R409 B.n275 B.n34 10.6151
R410 B.n275 B.n274 10.6151
R411 B.n274 B.n273 10.6151
R412 B.n273 B.n36 10.6151
R413 B.n269 B.n36 10.6151
R414 B.n269 B.n268 10.6151
R415 B.n268 B.n267 10.6151
R416 B.n267 B.n38 10.6151
R417 B.n263 B.n38 10.6151
R418 B.n263 B.n262 10.6151
R419 B.n197 B.n60 10.6151
R420 B.n201 B.n60 10.6151
R421 B.n202 B.n201 10.6151
R422 B.n203 B.n202 10.6151
R423 B.n203 B.n58 10.6151
R424 B.n207 B.n58 10.6151
R425 B.n208 B.n207 10.6151
R426 B.n209 B.n208 10.6151
R427 B.n209 B.n56 10.6151
R428 B.n213 B.n56 10.6151
R429 B.n214 B.n213 10.6151
R430 B.n215 B.n214 10.6151
R431 B.n215 B.n54 10.6151
R432 B.n219 B.n54 10.6151
R433 B.n220 B.n219 10.6151
R434 B.n221 B.n220 10.6151
R435 B.n221 B.n52 10.6151
R436 B.n225 B.n52 10.6151
R437 B.n226 B.n225 10.6151
R438 B.n227 B.n226 10.6151
R439 B.n227 B.n50 10.6151
R440 B.n231 B.n50 10.6151
R441 B.n232 B.n231 10.6151
R442 B.n233 B.n232 10.6151
R443 B.n233 B.n48 10.6151
R444 B.n237 B.n48 10.6151
R445 B.n238 B.n237 10.6151
R446 B.n239 B.n238 10.6151
R447 B.n239 B.n46 10.6151
R448 B.n243 B.n46 10.6151
R449 B.n244 B.n243 10.6151
R450 B.n245 B.n244 10.6151
R451 B.n245 B.n44 10.6151
R452 B.n249 B.n44 10.6151
R453 B.n250 B.n249 10.6151
R454 B.n251 B.n250 10.6151
R455 B.n251 B.n42 10.6151
R456 B.n255 B.n42 10.6151
R457 B.n256 B.n255 10.6151
R458 B.n257 B.n256 10.6151
R459 B.n257 B.n40 10.6151
R460 B.n261 B.n40 10.6151
R461 B.n130 B.n129 10.6151
R462 B.n131 B.n130 10.6151
R463 B.n131 B.n86 10.6151
R464 B.n135 B.n86 10.6151
R465 B.n136 B.n135 10.6151
R466 B.n137 B.n136 10.6151
R467 B.n137 B.n84 10.6151
R468 B.n141 B.n84 10.6151
R469 B.n142 B.n141 10.6151
R470 B.n143 B.n142 10.6151
R471 B.n143 B.n82 10.6151
R472 B.n147 B.n82 10.6151
R473 B.n148 B.n147 10.6151
R474 B.n149 B.n148 10.6151
R475 B.n149 B.n80 10.6151
R476 B.n153 B.n80 10.6151
R477 B.n154 B.n153 10.6151
R478 B.n156 B.n76 10.6151
R479 B.n160 B.n76 10.6151
R480 B.n161 B.n160 10.6151
R481 B.n162 B.n161 10.6151
R482 B.n162 B.n74 10.6151
R483 B.n166 B.n74 10.6151
R484 B.n167 B.n166 10.6151
R485 B.n168 B.n167 10.6151
R486 B.n172 B.n171 10.6151
R487 B.n173 B.n172 10.6151
R488 B.n173 B.n68 10.6151
R489 B.n177 B.n68 10.6151
R490 B.n178 B.n177 10.6151
R491 B.n179 B.n178 10.6151
R492 B.n179 B.n66 10.6151
R493 B.n183 B.n66 10.6151
R494 B.n184 B.n183 10.6151
R495 B.n185 B.n184 10.6151
R496 B.n185 B.n64 10.6151
R497 B.n189 B.n64 10.6151
R498 B.n190 B.n189 10.6151
R499 B.n191 B.n190 10.6151
R500 B.n191 B.n62 10.6151
R501 B.n195 B.n62 10.6151
R502 B.n196 B.n195 10.6151
R503 B.n125 B.n88 10.6151
R504 B.n125 B.n124 10.6151
R505 B.n124 B.n123 10.6151
R506 B.n123 B.n90 10.6151
R507 B.n119 B.n90 10.6151
R508 B.n119 B.n118 10.6151
R509 B.n118 B.n117 10.6151
R510 B.n117 B.n92 10.6151
R511 B.n113 B.n92 10.6151
R512 B.n113 B.n112 10.6151
R513 B.n112 B.n111 10.6151
R514 B.n111 B.n94 10.6151
R515 B.n107 B.n94 10.6151
R516 B.n107 B.n106 10.6151
R517 B.n106 B.n105 10.6151
R518 B.n105 B.n96 10.6151
R519 B.n101 B.n96 10.6151
R520 B.n101 B.n100 10.6151
R521 B.n100 B.n99 10.6151
R522 B.n99 B.n0 10.6151
R523 B.n359 B.n1 10.6151
R524 B.n359 B.n358 10.6151
R525 B.n358 B.n357 10.6151
R526 B.n357 B.n4 10.6151
R527 B.n353 B.n4 10.6151
R528 B.n353 B.n352 10.6151
R529 B.n352 B.n351 10.6151
R530 B.n351 B.n6 10.6151
R531 B.n347 B.n6 10.6151
R532 B.n347 B.n346 10.6151
R533 B.n346 B.n345 10.6151
R534 B.n345 B.n8 10.6151
R535 B.n341 B.n8 10.6151
R536 B.n341 B.n340 10.6151
R537 B.n340 B.n339 10.6151
R538 B.n339 B.n10 10.6151
R539 B.n335 B.n10 10.6151
R540 B.n335 B.n334 10.6151
R541 B.n334 B.n333 10.6151
R542 B.n333 B.n12 10.6151
R543 B.n303 B.n302 6.5566
R544 B.n290 B.n30 6.5566
R545 B.n156 B.n155 6.5566
R546 B.n168 B.n72 6.5566
R547 B.n304 B.n303 4.05904
R548 B.n287 B.n30 4.05904
R549 B.n155 B.n154 4.05904
R550 B.n171 B.n72 4.05904
R551 B.n363 B.n0 2.81026
R552 B.n363 B.n1 2.81026
R553 VN.n0 VN.t0 136.782
R554 VN.n1 VN.t1 136.782
R555 VN.n1 VN.t2 136.695
R556 VN.n0 VN.t3 136.695
R557 VN VN.n1 67.3796
R558 VN VN.n0 31.2622
R559 VDD2.n2 VDD2.n0 146.624
R560 VDD2.n2 VDD2.n1 115.701
R561 VDD2.n1 VDD2.t3 8.22961
R562 VDD2.n1 VDD2.t1 8.22961
R563 VDD2.n0 VDD2.t2 8.22961
R564 VDD2.n0 VDD2.t0 8.22961
R565 VDD2 VDD2.n2 0.0586897
R566 VTAIL.n154 VTAIL.n140 756.745
R567 VTAIL.n14 VTAIL.n0 756.745
R568 VTAIL.n34 VTAIL.n20 756.745
R569 VTAIL.n54 VTAIL.n40 756.745
R570 VTAIL.n134 VTAIL.n120 756.745
R571 VTAIL.n114 VTAIL.n100 756.745
R572 VTAIL.n94 VTAIL.n80 756.745
R573 VTAIL.n74 VTAIL.n60 756.745
R574 VTAIL.n147 VTAIL.n146 585
R575 VTAIL.n144 VTAIL.n143 585
R576 VTAIL.n153 VTAIL.n152 585
R577 VTAIL.n155 VTAIL.n154 585
R578 VTAIL.n7 VTAIL.n6 585
R579 VTAIL.n4 VTAIL.n3 585
R580 VTAIL.n13 VTAIL.n12 585
R581 VTAIL.n15 VTAIL.n14 585
R582 VTAIL.n27 VTAIL.n26 585
R583 VTAIL.n24 VTAIL.n23 585
R584 VTAIL.n33 VTAIL.n32 585
R585 VTAIL.n35 VTAIL.n34 585
R586 VTAIL.n47 VTAIL.n46 585
R587 VTAIL.n44 VTAIL.n43 585
R588 VTAIL.n53 VTAIL.n52 585
R589 VTAIL.n55 VTAIL.n54 585
R590 VTAIL.n135 VTAIL.n134 585
R591 VTAIL.n133 VTAIL.n132 585
R592 VTAIL.n124 VTAIL.n123 585
R593 VTAIL.n127 VTAIL.n126 585
R594 VTAIL.n115 VTAIL.n114 585
R595 VTAIL.n113 VTAIL.n112 585
R596 VTAIL.n104 VTAIL.n103 585
R597 VTAIL.n107 VTAIL.n106 585
R598 VTAIL.n95 VTAIL.n94 585
R599 VTAIL.n93 VTAIL.n92 585
R600 VTAIL.n84 VTAIL.n83 585
R601 VTAIL.n87 VTAIL.n86 585
R602 VTAIL.n75 VTAIL.n74 585
R603 VTAIL.n73 VTAIL.n72 585
R604 VTAIL.n64 VTAIL.n63 585
R605 VTAIL.n67 VTAIL.n66 585
R606 VTAIL.t4 VTAIL.n145 330.707
R607 VTAIL.t7 VTAIL.n5 330.707
R608 VTAIL.t1 VTAIL.n25 330.707
R609 VTAIL.t2 VTAIL.n45 330.707
R610 VTAIL.t0 VTAIL.n125 330.707
R611 VTAIL.t3 VTAIL.n105 330.707
R612 VTAIL.t6 VTAIL.n85 330.707
R613 VTAIL.t5 VTAIL.n65 330.707
R614 VTAIL.n146 VTAIL.n143 171.744
R615 VTAIL.n153 VTAIL.n143 171.744
R616 VTAIL.n154 VTAIL.n153 171.744
R617 VTAIL.n6 VTAIL.n3 171.744
R618 VTAIL.n13 VTAIL.n3 171.744
R619 VTAIL.n14 VTAIL.n13 171.744
R620 VTAIL.n26 VTAIL.n23 171.744
R621 VTAIL.n33 VTAIL.n23 171.744
R622 VTAIL.n34 VTAIL.n33 171.744
R623 VTAIL.n46 VTAIL.n43 171.744
R624 VTAIL.n53 VTAIL.n43 171.744
R625 VTAIL.n54 VTAIL.n53 171.744
R626 VTAIL.n134 VTAIL.n133 171.744
R627 VTAIL.n133 VTAIL.n123 171.744
R628 VTAIL.n126 VTAIL.n123 171.744
R629 VTAIL.n114 VTAIL.n113 171.744
R630 VTAIL.n113 VTAIL.n103 171.744
R631 VTAIL.n106 VTAIL.n103 171.744
R632 VTAIL.n94 VTAIL.n93 171.744
R633 VTAIL.n93 VTAIL.n83 171.744
R634 VTAIL.n86 VTAIL.n83 171.744
R635 VTAIL.n74 VTAIL.n73 171.744
R636 VTAIL.n73 VTAIL.n63 171.744
R637 VTAIL.n66 VTAIL.n63 171.744
R638 VTAIL.n146 VTAIL.t4 85.8723
R639 VTAIL.n6 VTAIL.t7 85.8723
R640 VTAIL.n26 VTAIL.t1 85.8723
R641 VTAIL.n46 VTAIL.t2 85.8723
R642 VTAIL.n126 VTAIL.t0 85.8723
R643 VTAIL.n106 VTAIL.t3 85.8723
R644 VTAIL.n86 VTAIL.t6 85.8723
R645 VTAIL.n66 VTAIL.t5 85.8723
R646 VTAIL.n159 VTAIL.n158 34.3187
R647 VTAIL.n19 VTAIL.n18 34.3187
R648 VTAIL.n39 VTAIL.n38 34.3187
R649 VTAIL.n59 VTAIL.n58 34.3187
R650 VTAIL.n139 VTAIL.n138 34.3187
R651 VTAIL.n119 VTAIL.n118 34.3187
R652 VTAIL.n99 VTAIL.n98 34.3187
R653 VTAIL.n79 VTAIL.n78 34.3187
R654 VTAIL.n159 VTAIL.n139 17.0393
R655 VTAIL.n79 VTAIL.n59 17.0393
R656 VTAIL.n147 VTAIL.n145 16.3201
R657 VTAIL.n7 VTAIL.n5 16.3201
R658 VTAIL.n27 VTAIL.n25 16.3201
R659 VTAIL.n47 VTAIL.n45 16.3201
R660 VTAIL.n127 VTAIL.n125 16.3201
R661 VTAIL.n107 VTAIL.n105 16.3201
R662 VTAIL.n87 VTAIL.n85 16.3201
R663 VTAIL.n67 VTAIL.n65 16.3201
R664 VTAIL.n148 VTAIL.n144 12.8005
R665 VTAIL.n8 VTAIL.n4 12.8005
R666 VTAIL.n28 VTAIL.n24 12.8005
R667 VTAIL.n48 VTAIL.n44 12.8005
R668 VTAIL.n128 VTAIL.n124 12.8005
R669 VTAIL.n108 VTAIL.n104 12.8005
R670 VTAIL.n88 VTAIL.n84 12.8005
R671 VTAIL.n68 VTAIL.n64 12.8005
R672 VTAIL.n152 VTAIL.n151 12.0247
R673 VTAIL.n12 VTAIL.n11 12.0247
R674 VTAIL.n32 VTAIL.n31 12.0247
R675 VTAIL.n52 VTAIL.n51 12.0247
R676 VTAIL.n132 VTAIL.n131 12.0247
R677 VTAIL.n112 VTAIL.n111 12.0247
R678 VTAIL.n92 VTAIL.n91 12.0247
R679 VTAIL.n72 VTAIL.n71 12.0247
R680 VTAIL.n155 VTAIL.n142 11.249
R681 VTAIL.n15 VTAIL.n2 11.249
R682 VTAIL.n35 VTAIL.n22 11.249
R683 VTAIL.n55 VTAIL.n42 11.249
R684 VTAIL.n135 VTAIL.n122 11.249
R685 VTAIL.n115 VTAIL.n102 11.249
R686 VTAIL.n95 VTAIL.n82 11.249
R687 VTAIL.n75 VTAIL.n62 11.249
R688 VTAIL.n156 VTAIL.n140 10.4732
R689 VTAIL.n16 VTAIL.n0 10.4732
R690 VTAIL.n36 VTAIL.n20 10.4732
R691 VTAIL.n56 VTAIL.n40 10.4732
R692 VTAIL.n136 VTAIL.n120 10.4732
R693 VTAIL.n116 VTAIL.n100 10.4732
R694 VTAIL.n96 VTAIL.n80 10.4732
R695 VTAIL.n76 VTAIL.n60 10.4732
R696 VTAIL.n158 VTAIL.n157 9.45567
R697 VTAIL.n18 VTAIL.n17 9.45567
R698 VTAIL.n38 VTAIL.n37 9.45567
R699 VTAIL.n58 VTAIL.n57 9.45567
R700 VTAIL.n138 VTAIL.n137 9.45567
R701 VTAIL.n118 VTAIL.n117 9.45567
R702 VTAIL.n98 VTAIL.n97 9.45567
R703 VTAIL.n78 VTAIL.n77 9.45567
R704 VTAIL.n157 VTAIL.n156 9.3005
R705 VTAIL.n142 VTAIL.n141 9.3005
R706 VTAIL.n151 VTAIL.n150 9.3005
R707 VTAIL.n149 VTAIL.n148 9.3005
R708 VTAIL.n17 VTAIL.n16 9.3005
R709 VTAIL.n2 VTAIL.n1 9.3005
R710 VTAIL.n11 VTAIL.n10 9.3005
R711 VTAIL.n9 VTAIL.n8 9.3005
R712 VTAIL.n37 VTAIL.n36 9.3005
R713 VTAIL.n22 VTAIL.n21 9.3005
R714 VTAIL.n31 VTAIL.n30 9.3005
R715 VTAIL.n29 VTAIL.n28 9.3005
R716 VTAIL.n57 VTAIL.n56 9.3005
R717 VTAIL.n42 VTAIL.n41 9.3005
R718 VTAIL.n51 VTAIL.n50 9.3005
R719 VTAIL.n49 VTAIL.n48 9.3005
R720 VTAIL.n137 VTAIL.n136 9.3005
R721 VTAIL.n122 VTAIL.n121 9.3005
R722 VTAIL.n131 VTAIL.n130 9.3005
R723 VTAIL.n129 VTAIL.n128 9.3005
R724 VTAIL.n117 VTAIL.n116 9.3005
R725 VTAIL.n102 VTAIL.n101 9.3005
R726 VTAIL.n111 VTAIL.n110 9.3005
R727 VTAIL.n109 VTAIL.n108 9.3005
R728 VTAIL.n97 VTAIL.n96 9.3005
R729 VTAIL.n82 VTAIL.n81 9.3005
R730 VTAIL.n91 VTAIL.n90 9.3005
R731 VTAIL.n89 VTAIL.n88 9.3005
R732 VTAIL.n77 VTAIL.n76 9.3005
R733 VTAIL.n62 VTAIL.n61 9.3005
R734 VTAIL.n71 VTAIL.n70 9.3005
R735 VTAIL.n69 VTAIL.n68 9.3005
R736 VTAIL.n149 VTAIL.n145 3.78097
R737 VTAIL.n9 VTAIL.n5 3.78097
R738 VTAIL.n29 VTAIL.n25 3.78097
R739 VTAIL.n49 VTAIL.n45 3.78097
R740 VTAIL.n129 VTAIL.n125 3.78097
R741 VTAIL.n109 VTAIL.n105 3.78097
R742 VTAIL.n89 VTAIL.n85 3.78097
R743 VTAIL.n69 VTAIL.n65 3.78097
R744 VTAIL.n158 VTAIL.n140 3.49141
R745 VTAIL.n18 VTAIL.n0 3.49141
R746 VTAIL.n38 VTAIL.n20 3.49141
R747 VTAIL.n58 VTAIL.n40 3.49141
R748 VTAIL.n138 VTAIL.n120 3.49141
R749 VTAIL.n118 VTAIL.n100 3.49141
R750 VTAIL.n98 VTAIL.n80 3.49141
R751 VTAIL.n78 VTAIL.n60 3.49141
R752 VTAIL.n156 VTAIL.n155 2.71565
R753 VTAIL.n16 VTAIL.n15 2.71565
R754 VTAIL.n36 VTAIL.n35 2.71565
R755 VTAIL.n56 VTAIL.n55 2.71565
R756 VTAIL.n136 VTAIL.n135 2.71565
R757 VTAIL.n116 VTAIL.n115 2.71565
R758 VTAIL.n96 VTAIL.n95 2.71565
R759 VTAIL.n76 VTAIL.n75 2.71565
R760 VTAIL.n152 VTAIL.n142 1.93989
R761 VTAIL.n12 VTAIL.n2 1.93989
R762 VTAIL.n32 VTAIL.n22 1.93989
R763 VTAIL.n52 VTAIL.n42 1.93989
R764 VTAIL.n132 VTAIL.n122 1.93989
R765 VTAIL.n112 VTAIL.n102 1.93989
R766 VTAIL.n92 VTAIL.n82 1.93989
R767 VTAIL.n72 VTAIL.n62 1.93989
R768 VTAIL.n99 VTAIL.n79 1.26774
R769 VTAIL.n139 VTAIL.n119 1.26774
R770 VTAIL.n59 VTAIL.n39 1.26774
R771 VTAIL.n151 VTAIL.n144 1.16414
R772 VTAIL.n11 VTAIL.n4 1.16414
R773 VTAIL.n31 VTAIL.n24 1.16414
R774 VTAIL.n51 VTAIL.n44 1.16414
R775 VTAIL.n131 VTAIL.n124 1.16414
R776 VTAIL.n111 VTAIL.n104 1.16414
R777 VTAIL.n91 VTAIL.n84 1.16414
R778 VTAIL.n71 VTAIL.n64 1.16414
R779 VTAIL VTAIL.n19 0.69231
R780 VTAIL VTAIL.n159 0.575931
R781 VTAIL.n119 VTAIL.n99 0.470328
R782 VTAIL.n39 VTAIL.n19 0.470328
R783 VTAIL.n148 VTAIL.n147 0.388379
R784 VTAIL.n8 VTAIL.n7 0.388379
R785 VTAIL.n28 VTAIL.n27 0.388379
R786 VTAIL.n48 VTAIL.n47 0.388379
R787 VTAIL.n128 VTAIL.n127 0.388379
R788 VTAIL.n108 VTAIL.n107 0.388379
R789 VTAIL.n88 VTAIL.n87 0.388379
R790 VTAIL.n68 VTAIL.n67 0.388379
R791 VTAIL.n150 VTAIL.n149 0.155672
R792 VTAIL.n150 VTAIL.n141 0.155672
R793 VTAIL.n157 VTAIL.n141 0.155672
R794 VTAIL.n10 VTAIL.n9 0.155672
R795 VTAIL.n10 VTAIL.n1 0.155672
R796 VTAIL.n17 VTAIL.n1 0.155672
R797 VTAIL.n30 VTAIL.n29 0.155672
R798 VTAIL.n30 VTAIL.n21 0.155672
R799 VTAIL.n37 VTAIL.n21 0.155672
R800 VTAIL.n50 VTAIL.n49 0.155672
R801 VTAIL.n50 VTAIL.n41 0.155672
R802 VTAIL.n57 VTAIL.n41 0.155672
R803 VTAIL.n137 VTAIL.n121 0.155672
R804 VTAIL.n130 VTAIL.n121 0.155672
R805 VTAIL.n130 VTAIL.n129 0.155672
R806 VTAIL.n117 VTAIL.n101 0.155672
R807 VTAIL.n110 VTAIL.n101 0.155672
R808 VTAIL.n110 VTAIL.n109 0.155672
R809 VTAIL.n97 VTAIL.n81 0.155672
R810 VTAIL.n90 VTAIL.n81 0.155672
R811 VTAIL.n90 VTAIL.n89 0.155672
R812 VTAIL.n77 VTAIL.n61 0.155672
R813 VTAIL.n70 VTAIL.n61 0.155672
R814 VTAIL.n70 VTAIL.n69 0.155672
R815 VP.n0 VP.t0 136.782
R816 VP.n0 VP.t2 136.695
R817 VP.n2 VP.t1 118.175
R818 VP.n3 VP.t3 118.175
R819 VP.n4 VP.n3 80.6037
R820 VP.n2 VP.n1 80.6037
R821 VP.n1 VP.n0 67.0941
R822 VP.n3 VP.n2 48.2005
R823 VP.n4 VP.n1 0.380177
R824 VP VP.n4 0.146778
R825 VDD1 VDD1.n1 147.149
R826 VDD1 VDD1.n0 115.76
R827 VDD1.n0 VDD1.t3 8.22961
R828 VDD1.n0 VDD1.t1 8.22961
R829 VDD1.n1 VDD1.t2 8.22961
R830 VDD1.n1 VDD1.t0 8.22961
C0 w_n1852_n1758# VDD1 0.945071f
C1 VN VP 3.64988f
C2 VP VDD2 0.306181f
C3 VTAIL w_n1852_n1758# 2.06964f
C4 VN B 0.734598f
C5 B VDD2 0.815316f
C6 VN VDD1 0.152086f
C7 VDD2 VDD1 0.672052f
C8 VN VTAIL 1.55937f
C9 VTAIL VDD2 3.11737f
C10 VN w_n1852_n1758# 2.69526f
C11 B VP 1.11655f
C12 w_n1852_n1758# VDD2 0.968471f
C13 VP VDD1 1.61432f
C14 VTAIL VP 1.57348f
C15 B VDD1 0.786858f
C16 VN VDD2 1.46099f
C17 VTAIL B 1.79953f
C18 w_n1852_n1758# VP 2.9287f
C19 VTAIL VDD1 3.07295f
C20 w_n1852_n1758# B 5.1935f
C21 VDD2 VSUBS 0.492952f
C22 VDD1 VSUBS 2.704642f
C23 VTAIL VSUBS 0.431516f
C24 VN VSUBS 3.99471f
C25 VP VSUBS 1.130676f
C26 B VSUBS 2.218568f
C27 w_n1852_n1758# VSUBS 41.0033f
C28 VDD1.t3 VSUBS 0.056034f
C29 VDD1.t1 VSUBS 0.056034f
C30 VDD1.n0 VSUBS 0.326375f
C31 VDD1.t2 VSUBS 0.056034f
C32 VDD1.t0 VSUBS 0.056034f
C33 VDD1.n1 VSUBS 0.508207f
C34 VP.t2 VSUBS 0.613775f
C35 VP.t0 VSUBS 0.614004f
C36 VP.n0 VSUBS 1.31171f
C37 VP.n1 VSUBS 2.11572f
C38 VP.t1 VSUBS 0.573436f
C39 VP.n2 VSUBS 0.297742f
C40 VP.t3 VSUBS 0.573436f
C41 VP.n3 VSUBS 0.297742f
C42 VP.n4 VSUBS 0.054792f
C43 VTAIL.n0 VSUBS 0.019318f
C44 VTAIL.n1 VSUBS 0.017717f
C45 VTAIL.n2 VSUBS 0.00952f
C46 VTAIL.n3 VSUBS 0.022503f
C47 VTAIL.n4 VSUBS 0.01008f
C48 VTAIL.n5 VSUBS 0.068715f
C49 VTAIL.t7 VSUBS 0.049791f
C50 VTAIL.n6 VSUBS 0.016877f
C51 VTAIL.n7 VSUBS 0.014154f
C52 VTAIL.n8 VSUBS 0.00952f
C53 VTAIL.n9 VSUBS 0.239002f
C54 VTAIL.n10 VSUBS 0.017717f
C55 VTAIL.n11 VSUBS 0.00952f
C56 VTAIL.n12 VSUBS 0.01008f
C57 VTAIL.n13 VSUBS 0.022503f
C58 VTAIL.n14 VSUBS 0.053969f
C59 VTAIL.n15 VSUBS 0.01008f
C60 VTAIL.n16 VSUBS 0.00952f
C61 VTAIL.n17 VSUBS 0.043615f
C62 VTAIL.n18 VSUBS 0.027197f
C63 VTAIL.n19 VSUBS 0.082953f
C64 VTAIL.n20 VSUBS 0.019318f
C65 VTAIL.n21 VSUBS 0.017717f
C66 VTAIL.n22 VSUBS 0.00952f
C67 VTAIL.n23 VSUBS 0.022503f
C68 VTAIL.n24 VSUBS 0.01008f
C69 VTAIL.n25 VSUBS 0.068715f
C70 VTAIL.t1 VSUBS 0.049791f
C71 VTAIL.n26 VSUBS 0.016877f
C72 VTAIL.n27 VSUBS 0.014154f
C73 VTAIL.n28 VSUBS 0.00952f
C74 VTAIL.n29 VSUBS 0.239002f
C75 VTAIL.n30 VSUBS 0.017717f
C76 VTAIL.n31 VSUBS 0.00952f
C77 VTAIL.n32 VSUBS 0.01008f
C78 VTAIL.n33 VSUBS 0.022503f
C79 VTAIL.n34 VSUBS 0.053969f
C80 VTAIL.n35 VSUBS 0.01008f
C81 VTAIL.n36 VSUBS 0.00952f
C82 VTAIL.n37 VSUBS 0.043615f
C83 VTAIL.n38 VSUBS 0.027197f
C84 VTAIL.n39 VSUBS 0.115804f
C85 VTAIL.n40 VSUBS 0.019318f
C86 VTAIL.n41 VSUBS 0.017717f
C87 VTAIL.n42 VSUBS 0.00952f
C88 VTAIL.n43 VSUBS 0.022503f
C89 VTAIL.n44 VSUBS 0.01008f
C90 VTAIL.n45 VSUBS 0.068715f
C91 VTAIL.t2 VSUBS 0.049791f
C92 VTAIL.n46 VSUBS 0.016877f
C93 VTAIL.n47 VSUBS 0.014154f
C94 VTAIL.n48 VSUBS 0.00952f
C95 VTAIL.n49 VSUBS 0.239002f
C96 VTAIL.n50 VSUBS 0.017717f
C97 VTAIL.n51 VSUBS 0.00952f
C98 VTAIL.n52 VSUBS 0.01008f
C99 VTAIL.n53 VSUBS 0.022503f
C100 VTAIL.n54 VSUBS 0.053969f
C101 VTAIL.n55 VSUBS 0.01008f
C102 VTAIL.n56 VSUBS 0.00952f
C103 VTAIL.n57 VSUBS 0.043615f
C104 VTAIL.n58 VSUBS 0.027197f
C105 VTAIL.n59 VSUBS 0.596391f
C106 VTAIL.n60 VSUBS 0.019318f
C107 VTAIL.n61 VSUBS 0.017717f
C108 VTAIL.n62 VSUBS 0.00952f
C109 VTAIL.n63 VSUBS 0.022503f
C110 VTAIL.n64 VSUBS 0.01008f
C111 VTAIL.n65 VSUBS 0.068715f
C112 VTAIL.t5 VSUBS 0.049791f
C113 VTAIL.n66 VSUBS 0.016877f
C114 VTAIL.n67 VSUBS 0.014154f
C115 VTAIL.n68 VSUBS 0.00952f
C116 VTAIL.n69 VSUBS 0.239002f
C117 VTAIL.n70 VSUBS 0.017717f
C118 VTAIL.n71 VSUBS 0.00952f
C119 VTAIL.n72 VSUBS 0.01008f
C120 VTAIL.n73 VSUBS 0.022503f
C121 VTAIL.n74 VSUBS 0.053969f
C122 VTAIL.n75 VSUBS 0.01008f
C123 VTAIL.n76 VSUBS 0.00952f
C124 VTAIL.n77 VSUBS 0.043615f
C125 VTAIL.n78 VSUBS 0.027197f
C126 VTAIL.n79 VSUBS 0.596391f
C127 VTAIL.n80 VSUBS 0.019318f
C128 VTAIL.n81 VSUBS 0.017717f
C129 VTAIL.n82 VSUBS 0.00952f
C130 VTAIL.n83 VSUBS 0.022503f
C131 VTAIL.n84 VSUBS 0.01008f
C132 VTAIL.n85 VSUBS 0.068715f
C133 VTAIL.t6 VSUBS 0.049791f
C134 VTAIL.n86 VSUBS 0.016877f
C135 VTAIL.n87 VSUBS 0.014154f
C136 VTAIL.n88 VSUBS 0.00952f
C137 VTAIL.n89 VSUBS 0.239002f
C138 VTAIL.n90 VSUBS 0.017717f
C139 VTAIL.n91 VSUBS 0.00952f
C140 VTAIL.n92 VSUBS 0.01008f
C141 VTAIL.n93 VSUBS 0.022503f
C142 VTAIL.n94 VSUBS 0.053969f
C143 VTAIL.n95 VSUBS 0.01008f
C144 VTAIL.n96 VSUBS 0.00952f
C145 VTAIL.n97 VSUBS 0.043615f
C146 VTAIL.n98 VSUBS 0.027197f
C147 VTAIL.n99 VSUBS 0.115804f
C148 VTAIL.n100 VSUBS 0.019318f
C149 VTAIL.n101 VSUBS 0.017717f
C150 VTAIL.n102 VSUBS 0.00952f
C151 VTAIL.n103 VSUBS 0.022503f
C152 VTAIL.n104 VSUBS 0.01008f
C153 VTAIL.n105 VSUBS 0.068715f
C154 VTAIL.t3 VSUBS 0.049791f
C155 VTAIL.n106 VSUBS 0.016877f
C156 VTAIL.n107 VSUBS 0.014154f
C157 VTAIL.n108 VSUBS 0.00952f
C158 VTAIL.n109 VSUBS 0.239002f
C159 VTAIL.n110 VSUBS 0.017717f
C160 VTAIL.n111 VSUBS 0.00952f
C161 VTAIL.n112 VSUBS 0.01008f
C162 VTAIL.n113 VSUBS 0.022503f
C163 VTAIL.n114 VSUBS 0.053969f
C164 VTAIL.n115 VSUBS 0.01008f
C165 VTAIL.n116 VSUBS 0.00952f
C166 VTAIL.n117 VSUBS 0.043615f
C167 VTAIL.n118 VSUBS 0.027197f
C168 VTAIL.n119 VSUBS 0.115804f
C169 VTAIL.n120 VSUBS 0.019318f
C170 VTAIL.n121 VSUBS 0.017717f
C171 VTAIL.n122 VSUBS 0.00952f
C172 VTAIL.n123 VSUBS 0.022503f
C173 VTAIL.n124 VSUBS 0.01008f
C174 VTAIL.n125 VSUBS 0.068715f
C175 VTAIL.t0 VSUBS 0.049791f
C176 VTAIL.n126 VSUBS 0.016877f
C177 VTAIL.n127 VSUBS 0.014154f
C178 VTAIL.n128 VSUBS 0.00952f
C179 VTAIL.n129 VSUBS 0.239002f
C180 VTAIL.n130 VSUBS 0.017717f
C181 VTAIL.n131 VSUBS 0.00952f
C182 VTAIL.n132 VSUBS 0.01008f
C183 VTAIL.n133 VSUBS 0.022503f
C184 VTAIL.n134 VSUBS 0.053969f
C185 VTAIL.n135 VSUBS 0.01008f
C186 VTAIL.n136 VSUBS 0.00952f
C187 VTAIL.n137 VSUBS 0.043615f
C188 VTAIL.n138 VSUBS 0.027197f
C189 VTAIL.n139 VSUBS 0.596391f
C190 VTAIL.n140 VSUBS 0.019318f
C191 VTAIL.n141 VSUBS 0.017717f
C192 VTAIL.n142 VSUBS 0.00952f
C193 VTAIL.n143 VSUBS 0.022503f
C194 VTAIL.n144 VSUBS 0.01008f
C195 VTAIL.n145 VSUBS 0.068715f
C196 VTAIL.t4 VSUBS 0.049791f
C197 VTAIL.n146 VSUBS 0.016877f
C198 VTAIL.n147 VSUBS 0.014154f
C199 VTAIL.n148 VSUBS 0.00952f
C200 VTAIL.n149 VSUBS 0.239002f
C201 VTAIL.n150 VSUBS 0.017717f
C202 VTAIL.n151 VSUBS 0.00952f
C203 VTAIL.n152 VSUBS 0.01008f
C204 VTAIL.n153 VSUBS 0.022503f
C205 VTAIL.n154 VSUBS 0.053969f
C206 VTAIL.n155 VSUBS 0.01008f
C207 VTAIL.n156 VSUBS 0.00952f
C208 VTAIL.n157 VSUBS 0.043615f
C209 VTAIL.n158 VSUBS 0.027197f
C210 VTAIL.n159 VSUBS 0.556897f
C211 VDD2.t2 VSUBS 0.057259f
C212 VDD2.t0 VSUBS 0.057259f
C213 VDD2.n0 VSUBS 0.508925f
C214 VDD2.t3 VSUBS 0.057259f
C215 VDD2.t1 VSUBS 0.057259f
C216 VDD2.n1 VSUBS 0.333336f
C217 VDD2.n2 VSUBS 1.94985f
C218 VN.t0 VSUBS 0.589614f
C219 VN.t3 VSUBS 0.589394f
C220 VN.n0 VSUBS 0.495302f
C221 VN.t1 VSUBS 0.589614f
C222 VN.t2 VSUBS 0.589394f
C223 VN.n1 VSUBS 1.27528f
C224 B.n0 VSUBS 0.004645f
C225 B.n1 VSUBS 0.004645f
C226 B.n2 VSUBS 0.007346f
C227 B.n3 VSUBS 0.007346f
C228 B.n4 VSUBS 0.007346f
C229 B.n5 VSUBS 0.007346f
C230 B.n6 VSUBS 0.007346f
C231 B.n7 VSUBS 0.007346f
C232 B.n8 VSUBS 0.007346f
C233 B.n9 VSUBS 0.007346f
C234 B.n10 VSUBS 0.007346f
C235 B.n11 VSUBS 0.007346f
C236 B.n12 VSUBS 0.017977f
C237 B.n13 VSUBS 0.007346f
C238 B.n14 VSUBS 0.007346f
C239 B.n15 VSUBS 0.007346f
C240 B.n16 VSUBS 0.007346f
C241 B.n17 VSUBS 0.007346f
C242 B.n18 VSUBS 0.007346f
C243 B.n19 VSUBS 0.007346f
C244 B.n20 VSUBS 0.007346f
C245 B.n21 VSUBS 0.007346f
C246 B.t8 VSUBS 0.060042f
C247 B.t7 VSUBS 0.071248f
C248 B.t6 VSUBS 0.218583f
C249 B.n22 VSUBS 0.129469f
C250 B.n23 VSUBS 0.113916f
C251 B.n24 VSUBS 0.007346f
C252 B.n25 VSUBS 0.007346f
C253 B.n26 VSUBS 0.007346f
C254 B.n27 VSUBS 0.007346f
C255 B.t5 VSUBS 0.060043f
C256 B.t4 VSUBS 0.071249f
C257 B.t3 VSUBS 0.218583f
C258 B.n28 VSUBS 0.129468f
C259 B.n29 VSUBS 0.113915f
C260 B.n30 VSUBS 0.01702f
C261 B.n31 VSUBS 0.007346f
C262 B.n32 VSUBS 0.007346f
C263 B.n33 VSUBS 0.007346f
C264 B.n34 VSUBS 0.007346f
C265 B.n35 VSUBS 0.007346f
C266 B.n36 VSUBS 0.007346f
C267 B.n37 VSUBS 0.007346f
C268 B.n38 VSUBS 0.007346f
C269 B.n39 VSUBS 0.018538f
C270 B.n40 VSUBS 0.007346f
C271 B.n41 VSUBS 0.007346f
C272 B.n42 VSUBS 0.007346f
C273 B.n43 VSUBS 0.007346f
C274 B.n44 VSUBS 0.007346f
C275 B.n45 VSUBS 0.007346f
C276 B.n46 VSUBS 0.007346f
C277 B.n47 VSUBS 0.007346f
C278 B.n48 VSUBS 0.007346f
C279 B.n49 VSUBS 0.007346f
C280 B.n50 VSUBS 0.007346f
C281 B.n51 VSUBS 0.007346f
C282 B.n52 VSUBS 0.007346f
C283 B.n53 VSUBS 0.007346f
C284 B.n54 VSUBS 0.007346f
C285 B.n55 VSUBS 0.007346f
C286 B.n56 VSUBS 0.007346f
C287 B.n57 VSUBS 0.007346f
C288 B.n58 VSUBS 0.007346f
C289 B.n59 VSUBS 0.007346f
C290 B.n60 VSUBS 0.007346f
C291 B.n61 VSUBS 0.018538f
C292 B.n62 VSUBS 0.007346f
C293 B.n63 VSUBS 0.007346f
C294 B.n64 VSUBS 0.007346f
C295 B.n65 VSUBS 0.007346f
C296 B.n66 VSUBS 0.007346f
C297 B.n67 VSUBS 0.007346f
C298 B.n68 VSUBS 0.007346f
C299 B.n69 VSUBS 0.007346f
C300 B.t1 VSUBS 0.060043f
C301 B.t2 VSUBS 0.071249f
C302 B.t0 VSUBS 0.218583f
C303 B.n70 VSUBS 0.129468f
C304 B.n71 VSUBS 0.113915f
C305 B.n72 VSUBS 0.01702f
C306 B.n73 VSUBS 0.007346f
C307 B.n74 VSUBS 0.007346f
C308 B.n75 VSUBS 0.007346f
C309 B.n76 VSUBS 0.007346f
C310 B.n77 VSUBS 0.007346f
C311 B.t10 VSUBS 0.060042f
C312 B.t11 VSUBS 0.071248f
C313 B.t9 VSUBS 0.218583f
C314 B.n78 VSUBS 0.129469f
C315 B.n79 VSUBS 0.113916f
C316 B.n80 VSUBS 0.007346f
C317 B.n81 VSUBS 0.007346f
C318 B.n82 VSUBS 0.007346f
C319 B.n83 VSUBS 0.007346f
C320 B.n84 VSUBS 0.007346f
C321 B.n85 VSUBS 0.007346f
C322 B.n86 VSUBS 0.007346f
C323 B.n87 VSUBS 0.007346f
C324 B.n88 VSUBS 0.017977f
C325 B.n89 VSUBS 0.007346f
C326 B.n90 VSUBS 0.007346f
C327 B.n91 VSUBS 0.007346f
C328 B.n92 VSUBS 0.007346f
C329 B.n93 VSUBS 0.007346f
C330 B.n94 VSUBS 0.007346f
C331 B.n95 VSUBS 0.007346f
C332 B.n96 VSUBS 0.007346f
C333 B.n97 VSUBS 0.007346f
C334 B.n98 VSUBS 0.007346f
C335 B.n99 VSUBS 0.007346f
C336 B.n100 VSUBS 0.007346f
C337 B.n101 VSUBS 0.007346f
C338 B.n102 VSUBS 0.007346f
C339 B.n103 VSUBS 0.007346f
C340 B.n104 VSUBS 0.007346f
C341 B.n105 VSUBS 0.007346f
C342 B.n106 VSUBS 0.007346f
C343 B.n107 VSUBS 0.007346f
C344 B.n108 VSUBS 0.007346f
C345 B.n109 VSUBS 0.007346f
C346 B.n110 VSUBS 0.007346f
C347 B.n111 VSUBS 0.007346f
C348 B.n112 VSUBS 0.007346f
C349 B.n113 VSUBS 0.007346f
C350 B.n114 VSUBS 0.007346f
C351 B.n115 VSUBS 0.007346f
C352 B.n116 VSUBS 0.007346f
C353 B.n117 VSUBS 0.007346f
C354 B.n118 VSUBS 0.007346f
C355 B.n119 VSUBS 0.007346f
C356 B.n120 VSUBS 0.007346f
C357 B.n121 VSUBS 0.007346f
C358 B.n122 VSUBS 0.007346f
C359 B.n123 VSUBS 0.007346f
C360 B.n124 VSUBS 0.007346f
C361 B.n125 VSUBS 0.007346f
C362 B.n126 VSUBS 0.007346f
C363 B.n127 VSUBS 0.017977f
C364 B.n128 VSUBS 0.018538f
C365 B.n129 VSUBS 0.018538f
C366 B.n130 VSUBS 0.007346f
C367 B.n131 VSUBS 0.007346f
C368 B.n132 VSUBS 0.007346f
C369 B.n133 VSUBS 0.007346f
C370 B.n134 VSUBS 0.007346f
C371 B.n135 VSUBS 0.007346f
C372 B.n136 VSUBS 0.007346f
C373 B.n137 VSUBS 0.007346f
C374 B.n138 VSUBS 0.007346f
C375 B.n139 VSUBS 0.007346f
C376 B.n140 VSUBS 0.007346f
C377 B.n141 VSUBS 0.007346f
C378 B.n142 VSUBS 0.007346f
C379 B.n143 VSUBS 0.007346f
C380 B.n144 VSUBS 0.007346f
C381 B.n145 VSUBS 0.007346f
C382 B.n146 VSUBS 0.007346f
C383 B.n147 VSUBS 0.007346f
C384 B.n148 VSUBS 0.007346f
C385 B.n149 VSUBS 0.007346f
C386 B.n150 VSUBS 0.007346f
C387 B.n151 VSUBS 0.007346f
C388 B.n152 VSUBS 0.007346f
C389 B.n153 VSUBS 0.007346f
C390 B.n154 VSUBS 0.005077f
C391 B.n155 VSUBS 0.01702f
C392 B.n156 VSUBS 0.005942f
C393 B.n157 VSUBS 0.007346f
C394 B.n158 VSUBS 0.007346f
C395 B.n159 VSUBS 0.007346f
C396 B.n160 VSUBS 0.007346f
C397 B.n161 VSUBS 0.007346f
C398 B.n162 VSUBS 0.007346f
C399 B.n163 VSUBS 0.007346f
C400 B.n164 VSUBS 0.007346f
C401 B.n165 VSUBS 0.007346f
C402 B.n166 VSUBS 0.007346f
C403 B.n167 VSUBS 0.007346f
C404 B.n168 VSUBS 0.005942f
C405 B.n169 VSUBS 0.007346f
C406 B.n170 VSUBS 0.007346f
C407 B.n171 VSUBS 0.005077f
C408 B.n172 VSUBS 0.007346f
C409 B.n173 VSUBS 0.007346f
C410 B.n174 VSUBS 0.007346f
C411 B.n175 VSUBS 0.007346f
C412 B.n176 VSUBS 0.007346f
C413 B.n177 VSUBS 0.007346f
C414 B.n178 VSUBS 0.007346f
C415 B.n179 VSUBS 0.007346f
C416 B.n180 VSUBS 0.007346f
C417 B.n181 VSUBS 0.007346f
C418 B.n182 VSUBS 0.007346f
C419 B.n183 VSUBS 0.007346f
C420 B.n184 VSUBS 0.007346f
C421 B.n185 VSUBS 0.007346f
C422 B.n186 VSUBS 0.007346f
C423 B.n187 VSUBS 0.007346f
C424 B.n188 VSUBS 0.007346f
C425 B.n189 VSUBS 0.007346f
C426 B.n190 VSUBS 0.007346f
C427 B.n191 VSUBS 0.007346f
C428 B.n192 VSUBS 0.007346f
C429 B.n193 VSUBS 0.007346f
C430 B.n194 VSUBS 0.007346f
C431 B.n195 VSUBS 0.007346f
C432 B.n196 VSUBS 0.018538f
C433 B.n197 VSUBS 0.017977f
C434 B.n198 VSUBS 0.017977f
C435 B.n199 VSUBS 0.007346f
C436 B.n200 VSUBS 0.007346f
C437 B.n201 VSUBS 0.007346f
C438 B.n202 VSUBS 0.007346f
C439 B.n203 VSUBS 0.007346f
C440 B.n204 VSUBS 0.007346f
C441 B.n205 VSUBS 0.007346f
C442 B.n206 VSUBS 0.007346f
C443 B.n207 VSUBS 0.007346f
C444 B.n208 VSUBS 0.007346f
C445 B.n209 VSUBS 0.007346f
C446 B.n210 VSUBS 0.007346f
C447 B.n211 VSUBS 0.007346f
C448 B.n212 VSUBS 0.007346f
C449 B.n213 VSUBS 0.007346f
C450 B.n214 VSUBS 0.007346f
C451 B.n215 VSUBS 0.007346f
C452 B.n216 VSUBS 0.007346f
C453 B.n217 VSUBS 0.007346f
C454 B.n218 VSUBS 0.007346f
C455 B.n219 VSUBS 0.007346f
C456 B.n220 VSUBS 0.007346f
C457 B.n221 VSUBS 0.007346f
C458 B.n222 VSUBS 0.007346f
C459 B.n223 VSUBS 0.007346f
C460 B.n224 VSUBS 0.007346f
C461 B.n225 VSUBS 0.007346f
C462 B.n226 VSUBS 0.007346f
C463 B.n227 VSUBS 0.007346f
C464 B.n228 VSUBS 0.007346f
C465 B.n229 VSUBS 0.007346f
C466 B.n230 VSUBS 0.007346f
C467 B.n231 VSUBS 0.007346f
C468 B.n232 VSUBS 0.007346f
C469 B.n233 VSUBS 0.007346f
C470 B.n234 VSUBS 0.007346f
C471 B.n235 VSUBS 0.007346f
C472 B.n236 VSUBS 0.007346f
C473 B.n237 VSUBS 0.007346f
C474 B.n238 VSUBS 0.007346f
C475 B.n239 VSUBS 0.007346f
C476 B.n240 VSUBS 0.007346f
C477 B.n241 VSUBS 0.007346f
C478 B.n242 VSUBS 0.007346f
C479 B.n243 VSUBS 0.007346f
C480 B.n244 VSUBS 0.007346f
C481 B.n245 VSUBS 0.007346f
C482 B.n246 VSUBS 0.007346f
C483 B.n247 VSUBS 0.007346f
C484 B.n248 VSUBS 0.007346f
C485 B.n249 VSUBS 0.007346f
C486 B.n250 VSUBS 0.007346f
C487 B.n251 VSUBS 0.007346f
C488 B.n252 VSUBS 0.007346f
C489 B.n253 VSUBS 0.007346f
C490 B.n254 VSUBS 0.007346f
C491 B.n255 VSUBS 0.007346f
C492 B.n256 VSUBS 0.007346f
C493 B.n257 VSUBS 0.007346f
C494 B.n258 VSUBS 0.007346f
C495 B.n259 VSUBS 0.007346f
C496 B.n260 VSUBS 0.017977f
C497 B.n261 VSUBS 0.01877f
C498 B.n262 VSUBS 0.017745f
C499 B.n263 VSUBS 0.007346f
C500 B.n264 VSUBS 0.007346f
C501 B.n265 VSUBS 0.007346f
C502 B.n266 VSUBS 0.007346f
C503 B.n267 VSUBS 0.007346f
C504 B.n268 VSUBS 0.007346f
C505 B.n269 VSUBS 0.007346f
C506 B.n270 VSUBS 0.007346f
C507 B.n271 VSUBS 0.007346f
C508 B.n272 VSUBS 0.007346f
C509 B.n273 VSUBS 0.007346f
C510 B.n274 VSUBS 0.007346f
C511 B.n275 VSUBS 0.007346f
C512 B.n276 VSUBS 0.007346f
C513 B.n277 VSUBS 0.007346f
C514 B.n278 VSUBS 0.007346f
C515 B.n279 VSUBS 0.007346f
C516 B.n280 VSUBS 0.007346f
C517 B.n281 VSUBS 0.007346f
C518 B.n282 VSUBS 0.007346f
C519 B.n283 VSUBS 0.007346f
C520 B.n284 VSUBS 0.007346f
C521 B.n285 VSUBS 0.007346f
C522 B.n286 VSUBS 0.007346f
C523 B.n287 VSUBS 0.005077f
C524 B.n288 VSUBS 0.007346f
C525 B.n289 VSUBS 0.007346f
C526 B.n290 VSUBS 0.005942f
C527 B.n291 VSUBS 0.007346f
C528 B.n292 VSUBS 0.007346f
C529 B.n293 VSUBS 0.007346f
C530 B.n294 VSUBS 0.007346f
C531 B.n295 VSUBS 0.007346f
C532 B.n296 VSUBS 0.007346f
C533 B.n297 VSUBS 0.007346f
C534 B.n298 VSUBS 0.007346f
C535 B.n299 VSUBS 0.007346f
C536 B.n300 VSUBS 0.007346f
C537 B.n301 VSUBS 0.007346f
C538 B.n302 VSUBS 0.005942f
C539 B.n303 VSUBS 0.01702f
C540 B.n304 VSUBS 0.005077f
C541 B.n305 VSUBS 0.007346f
C542 B.n306 VSUBS 0.007346f
C543 B.n307 VSUBS 0.007346f
C544 B.n308 VSUBS 0.007346f
C545 B.n309 VSUBS 0.007346f
C546 B.n310 VSUBS 0.007346f
C547 B.n311 VSUBS 0.007346f
C548 B.n312 VSUBS 0.007346f
C549 B.n313 VSUBS 0.007346f
C550 B.n314 VSUBS 0.007346f
C551 B.n315 VSUBS 0.007346f
C552 B.n316 VSUBS 0.007346f
C553 B.n317 VSUBS 0.007346f
C554 B.n318 VSUBS 0.007346f
C555 B.n319 VSUBS 0.007346f
C556 B.n320 VSUBS 0.007346f
C557 B.n321 VSUBS 0.007346f
C558 B.n322 VSUBS 0.007346f
C559 B.n323 VSUBS 0.007346f
C560 B.n324 VSUBS 0.007346f
C561 B.n325 VSUBS 0.007346f
C562 B.n326 VSUBS 0.007346f
C563 B.n327 VSUBS 0.007346f
C564 B.n328 VSUBS 0.007346f
C565 B.n329 VSUBS 0.018538f
C566 B.n330 VSUBS 0.018538f
C567 B.n331 VSUBS 0.017977f
C568 B.n332 VSUBS 0.007346f
C569 B.n333 VSUBS 0.007346f
C570 B.n334 VSUBS 0.007346f
C571 B.n335 VSUBS 0.007346f
C572 B.n336 VSUBS 0.007346f
C573 B.n337 VSUBS 0.007346f
C574 B.n338 VSUBS 0.007346f
C575 B.n339 VSUBS 0.007346f
C576 B.n340 VSUBS 0.007346f
C577 B.n341 VSUBS 0.007346f
C578 B.n342 VSUBS 0.007346f
C579 B.n343 VSUBS 0.007346f
C580 B.n344 VSUBS 0.007346f
C581 B.n345 VSUBS 0.007346f
C582 B.n346 VSUBS 0.007346f
C583 B.n347 VSUBS 0.007346f
C584 B.n348 VSUBS 0.007346f
C585 B.n349 VSUBS 0.007346f
C586 B.n350 VSUBS 0.007346f
C587 B.n351 VSUBS 0.007346f
C588 B.n352 VSUBS 0.007346f
C589 B.n353 VSUBS 0.007346f
C590 B.n354 VSUBS 0.007346f
C591 B.n355 VSUBS 0.007346f
C592 B.n356 VSUBS 0.007346f
C593 B.n357 VSUBS 0.007346f
C594 B.n358 VSUBS 0.007346f
C595 B.n359 VSUBS 0.007346f
C596 B.n360 VSUBS 0.007346f
C597 B.n361 VSUBS 0.007346f
C598 B.n362 VSUBS 0.007346f
C599 B.n363 VSUBS 0.016634f
.ends

