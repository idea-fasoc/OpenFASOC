* NGSPICE file created from diff_pair_sample_1783.ext - technology: sky130A

.subckt diff_pair_sample_1783 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=3.15645 pd=19.46 as=7.4607 ps=39.04 w=19.13 l=0.68
X1 VTAIL.t7 VP.t1 VDD1.t2 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=7.4607 pd=39.04 as=3.15645 ps=19.46 w=19.13 l=0.68
X2 VTAIL.t2 VN.t0 VDD2.t3 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=7.4607 pd=39.04 as=3.15645 ps=19.46 w=19.13 l=0.68
X3 B.t11 B.t9 B.t10 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=7.4607 pd=39.04 as=0 ps=0 w=19.13 l=0.68
X4 VTAIL.t4 VP.t2 VDD1.t1 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=7.4607 pd=39.04 as=3.15645 ps=19.46 w=19.13 l=0.68
X5 B.t8 B.t6 B.t7 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=7.4607 pd=39.04 as=0 ps=0 w=19.13 l=0.68
X6 VDD2.t2 VN.t1 VTAIL.t1 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=3.15645 pd=19.46 as=7.4607 ps=39.04 w=19.13 l=0.68
X7 B.t5 B.t3 B.t4 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=7.4607 pd=39.04 as=0 ps=0 w=19.13 l=0.68
X8 VTAIL.t0 VN.t2 VDD2.t1 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=7.4607 pd=39.04 as=3.15645 ps=19.46 w=19.13 l=0.68
X9 VDD2.t0 VN.t3 VTAIL.t3 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=3.15645 pd=19.46 as=7.4607 ps=39.04 w=19.13 l=0.68
X10 VDD1.t0 VP.t3 VTAIL.t6 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=3.15645 pd=19.46 as=7.4607 ps=39.04 w=19.13 l=0.68
X11 B.t2 B.t0 B.t1 w_n1576_n4794# sky130_fd_pr__pfet_01v8 ad=7.4607 pd=39.04 as=0 ps=0 w=19.13 l=0.68
R0 VP.n1 VP.t2 757.11
R1 VP.n1 VP.t0 757.061
R2 VP.n3 VP.t1 736.114
R3 VP.n5 VP.t3 736.114
R4 VP.n6 VP.n5 161.3
R5 VP.n4 VP.n0 161.3
R6 VP.n3 VP.n2 161.3
R7 VP.n2 VP.n1 90.3969
R8 VP.n4 VP.n3 24.1005
R9 VP.n5 VP.n4 24.1005
R10 VP.n2 VP.n0 0.189894
R11 VP.n6 VP.n0 0.189894
R12 VP VP.n6 0.0516364
R13 VTAIL.n5 VTAIL.t4 56.2873
R14 VTAIL.n4 VTAIL.t1 56.2873
R15 VTAIL.n3 VTAIL.t2 56.2873
R16 VTAIL.n7 VTAIL.t3 56.2871
R17 VTAIL.n0 VTAIL.t0 56.2871
R18 VTAIL.n1 VTAIL.t6 56.2871
R19 VTAIL.n2 VTAIL.t7 56.2871
R20 VTAIL.n6 VTAIL.t5 56.2871
R21 VTAIL.n7 VTAIL.n6 29.7289
R22 VTAIL.n3 VTAIL.n2 29.7289
R23 VTAIL.n4 VTAIL.n3 0.87119
R24 VTAIL.n6 VTAIL.n5 0.87119
R25 VTAIL.n2 VTAIL.n1 0.87119
R26 VTAIL VTAIL.n0 0.494034
R27 VTAIL.n5 VTAIL.n4 0.470328
R28 VTAIL.n1 VTAIL.n0 0.470328
R29 VTAIL VTAIL.n7 0.377655
R30 VDD1 VDD1.n1 114.609
R31 VDD1 VDD1.n0 71.325
R32 VDD1.n0 VDD1.t1 1.69966
R33 VDD1.n0 VDD1.t3 1.69966
R34 VDD1.n1 VDD1.t2 1.69966
R35 VDD1.n1 VDD1.t0 1.69966
R36 VN.n0 VN.t2 757.11
R37 VN.n1 VN.t1 757.11
R38 VN.n0 VN.t3 757.061
R39 VN.n1 VN.t0 757.061
R40 VN VN.n1 90.7776
R41 VN VN.n0 44.7132
R42 VDD2.n2 VDD2.n0 114.084
R43 VDD2.n2 VDD2.n1 71.2668
R44 VDD2.n1 VDD2.t3 1.69966
R45 VDD2.n1 VDD2.t2 1.69966
R46 VDD2.n0 VDD2.t1 1.69966
R47 VDD2.n0 VDD2.t0 1.69966
R48 VDD2 VDD2.n2 0.0586897
R49 B.n132 B.t9 881.208
R50 B.n138 B.t3 881.208
R51 B.n42 B.t6 881.208
R52 B.n50 B.t0 881.208
R53 B.n461 B.n82 585
R54 B.n463 B.n462 585
R55 B.n464 B.n81 585
R56 B.n466 B.n465 585
R57 B.n467 B.n80 585
R58 B.n469 B.n468 585
R59 B.n470 B.n79 585
R60 B.n472 B.n471 585
R61 B.n473 B.n78 585
R62 B.n475 B.n474 585
R63 B.n476 B.n77 585
R64 B.n478 B.n477 585
R65 B.n479 B.n76 585
R66 B.n481 B.n480 585
R67 B.n482 B.n75 585
R68 B.n484 B.n483 585
R69 B.n485 B.n74 585
R70 B.n487 B.n486 585
R71 B.n488 B.n73 585
R72 B.n490 B.n489 585
R73 B.n491 B.n72 585
R74 B.n493 B.n492 585
R75 B.n494 B.n71 585
R76 B.n496 B.n495 585
R77 B.n497 B.n70 585
R78 B.n499 B.n498 585
R79 B.n500 B.n69 585
R80 B.n502 B.n501 585
R81 B.n503 B.n68 585
R82 B.n505 B.n504 585
R83 B.n506 B.n67 585
R84 B.n508 B.n507 585
R85 B.n509 B.n66 585
R86 B.n511 B.n510 585
R87 B.n512 B.n65 585
R88 B.n514 B.n513 585
R89 B.n515 B.n64 585
R90 B.n517 B.n516 585
R91 B.n518 B.n63 585
R92 B.n520 B.n519 585
R93 B.n521 B.n62 585
R94 B.n523 B.n522 585
R95 B.n524 B.n61 585
R96 B.n526 B.n525 585
R97 B.n527 B.n60 585
R98 B.n529 B.n528 585
R99 B.n530 B.n59 585
R100 B.n532 B.n531 585
R101 B.n533 B.n58 585
R102 B.n535 B.n534 585
R103 B.n536 B.n57 585
R104 B.n538 B.n537 585
R105 B.n539 B.n56 585
R106 B.n541 B.n540 585
R107 B.n542 B.n55 585
R108 B.n544 B.n543 585
R109 B.n545 B.n54 585
R110 B.n547 B.n546 585
R111 B.n548 B.n53 585
R112 B.n550 B.n549 585
R113 B.n551 B.n52 585
R114 B.n553 B.n552 585
R115 B.n554 B.n49 585
R116 B.n557 B.n556 585
R117 B.n558 B.n48 585
R118 B.n560 B.n559 585
R119 B.n561 B.n47 585
R120 B.n563 B.n562 585
R121 B.n564 B.n46 585
R122 B.n566 B.n565 585
R123 B.n567 B.n45 585
R124 B.n569 B.n568 585
R125 B.n571 B.n570 585
R126 B.n572 B.n41 585
R127 B.n574 B.n573 585
R128 B.n575 B.n40 585
R129 B.n577 B.n576 585
R130 B.n578 B.n39 585
R131 B.n580 B.n579 585
R132 B.n581 B.n38 585
R133 B.n583 B.n582 585
R134 B.n584 B.n37 585
R135 B.n586 B.n585 585
R136 B.n587 B.n36 585
R137 B.n589 B.n588 585
R138 B.n590 B.n35 585
R139 B.n592 B.n591 585
R140 B.n593 B.n34 585
R141 B.n595 B.n594 585
R142 B.n596 B.n33 585
R143 B.n598 B.n597 585
R144 B.n599 B.n32 585
R145 B.n601 B.n600 585
R146 B.n602 B.n31 585
R147 B.n604 B.n603 585
R148 B.n605 B.n30 585
R149 B.n607 B.n606 585
R150 B.n608 B.n29 585
R151 B.n610 B.n609 585
R152 B.n611 B.n28 585
R153 B.n613 B.n612 585
R154 B.n614 B.n27 585
R155 B.n616 B.n615 585
R156 B.n617 B.n26 585
R157 B.n619 B.n618 585
R158 B.n620 B.n25 585
R159 B.n622 B.n621 585
R160 B.n623 B.n24 585
R161 B.n625 B.n624 585
R162 B.n626 B.n23 585
R163 B.n628 B.n627 585
R164 B.n629 B.n22 585
R165 B.n631 B.n630 585
R166 B.n632 B.n21 585
R167 B.n634 B.n633 585
R168 B.n635 B.n20 585
R169 B.n637 B.n636 585
R170 B.n638 B.n19 585
R171 B.n640 B.n639 585
R172 B.n641 B.n18 585
R173 B.n643 B.n642 585
R174 B.n644 B.n17 585
R175 B.n646 B.n645 585
R176 B.n647 B.n16 585
R177 B.n649 B.n648 585
R178 B.n650 B.n15 585
R179 B.n652 B.n651 585
R180 B.n653 B.n14 585
R181 B.n655 B.n654 585
R182 B.n656 B.n13 585
R183 B.n658 B.n657 585
R184 B.n659 B.n12 585
R185 B.n661 B.n660 585
R186 B.n662 B.n11 585
R187 B.n664 B.n663 585
R188 B.n460 B.n459 585
R189 B.n458 B.n83 585
R190 B.n457 B.n456 585
R191 B.n455 B.n84 585
R192 B.n454 B.n453 585
R193 B.n452 B.n85 585
R194 B.n451 B.n450 585
R195 B.n449 B.n86 585
R196 B.n448 B.n447 585
R197 B.n446 B.n87 585
R198 B.n445 B.n444 585
R199 B.n443 B.n88 585
R200 B.n442 B.n441 585
R201 B.n440 B.n89 585
R202 B.n439 B.n438 585
R203 B.n437 B.n90 585
R204 B.n436 B.n435 585
R205 B.n434 B.n91 585
R206 B.n433 B.n432 585
R207 B.n431 B.n92 585
R208 B.n430 B.n429 585
R209 B.n428 B.n93 585
R210 B.n427 B.n426 585
R211 B.n425 B.n94 585
R212 B.n424 B.n423 585
R213 B.n422 B.n95 585
R214 B.n421 B.n420 585
R215 B.n419 B.n96 585
R216 B.n418 B.n417 585
R217 B.n416 B.n97 585
R218 B.n415 B.n414 585
R219 B.n413 B.n98 585
R220 B.n412 B.n411 585
R221 B.n410 B.n99 585
R222 B.n409 B.n408 585
R223 B.n205 B.n204 585
R224 B.n206 B.n171 585
R225 B.n208 B.n207 585
R226 B.n209 B.n170 585
R227 B.n211 B.n210 585
R228 B.n212 B.n169 585
R229 B.n214 B.n213 585
R230 B.n215 B.n168 585
R231 B.n217 B.n216 585
R232 B.n218 B.n167 585
R233 B.n220 B.n219 585
R234 B.n221 B.n166 585
R235 B.n223 B.n222 585
R236 B.n224 B.n165 585
R237 B.n226 B.n225 585
R238 B.n227 B.n164 585
R239 B.n229 B.n228 585
R240 B.n230 B.n163 585
R241 B.n232 B.n231 585
R242 B.n233 B.n162 585
R243 B.n235 B.n234 585
R244 B.n236 B.n161 585
R245 B.n238 B.n237 585
R246 B.n239 B.n160 585
R247 B.n241 B.n240 585
R248 B.n242 B.n159 585
R249 B.n244 B.n243 585
R250 B.n245 B.n158 585
R251 B.n247 B.n246 585
R252 B.n248 B.n157 585
R253 B.n250 B.n249 585
R254 B.n251 B.n156 585
R255 B.n253 B.n252 585
R256 B.n254 B.n155 585
R257 B.n256 B.n255 585
R258 B.n257 B.n154 585
R259 B.n259 B.n258 585
R260 B.n260 B.n153 585
R261 B.n262 B.n261 585
R262 B.n263 B.n152 585
R263 B.n265 B.n264 585
R264 B.n266 B.n151 585
R265 B.n268 B.n267 585
R266 B.n269 B.n150 585
R267 B.n271 B.n270 585
R268 B.n272 B.n149 585
R269 B.n274 B.n273 585
R270 B.n275 B.n148 585
R271 B.n277 B.n276 585
R272 B.n278 B.n147 585
R273 B.n280 B.n279 585
R274 B.n281 B.n146 585
R275 B.n283 B.n282 585
R276 B.n284 B.n145 585
R277 B.n286 B.n285 585
R278 B.n287 B.n144 585
R279 B.n289 B.n288 585
R280 B.n290 B.n143 585
R281 B.n292 B.n291 585
R282 B.n293 B.n142 585
R283 B.n295 B.n294 585
R284 B.n296 B.n141 585
R285 B.n298 B.n297 585
R286 B.n300 B.n299 585
R287 B.n301 B.n137 585
R288 B.n303 B.n302 585
R289 B.n304 B.n136 585
R290 B.n306 B.n305 585
R291 B.n307 B.n135 585
R292 B.n309 B.n308 585
R293 B.n310 B.n134 585
R294 B.n312 B.n311 585
R295 B.n314 B.n131 585
R296 B.n316 B.n315 585
R297 B.n317 B.n130 585
R298 B.n319 B.n318 585
R299 B.n320 B.n129 585
R300 B.n322 B.n321 585
R301 B.n323 B.n128 585
R302 B.n325 B.n324 585
R303 B.n326 B.n127 585
R304 B.n328 B.n327 585
R305 B.n329 B.n126 585
R306 B.n331 B.n330 585
R307 B.n332 B.n125 585
R308 B.n334 B.n333 585
R309 B.n335 B.n124 585
R310 B.n337 B.n336 585
R311 B.n338 B.n123 585
R312 B.n340 B.n339 585
R313 B.n341 B.n122 585
R314 B.n343 B.n342 585
R315 B.n344 B.n121 585
R316 B.n346 B.n345 585
R317 B.n347 B.n120 585
R318 B.n349 B.n348 585
R319 B.n350 B.n119 585
R320 B.n352 B.n351 585
R321 B.n353 B.n118 585
R322 B.n355 B.n354 585
R323 B.n356 B.n117 585
R324 B.n358 B.n357 585
R325 B.n359 B.n116 585
R326 B.n361 B.n360 585
R327 B.n362 B.n115 585
R328 B.n364 B.n363 585
R329 B.n365 B.n114 585
R330 B.n367 B.n366 585
R331 B.n368 B.n113 585
R332 B.n370 B.n369 585
R333 B.n371 B.n112 585
R334 B.n373 B.n372 585
R335 B.n374 B.n111 585
R336 B.n376 B.n375 585
R337 B.n377 B.n110 585
R338 B.n379 B.n378 585
R339 B.n380 B.n109 585
R340 B.n382 B.n381 585
R341 B.n383 B.n108 585
R342 B.n385 B.n384 585
R343 B.n386 B.n107 585
R344 B.n388 B.n387 585
R345 B.n389 B.n106 585
R346 B.n391 B.n390 585
R347 B.n392 B.n105 585
R348 B.n394 B.n393 585
R349 B.n395 B.n104 585
R350 B.n397 B.n396 585
R351 B.n398 B.n103 585
R352 B.n400 B.n399 585
R353 B.n401 B.n102 585
R354 B.n403 B.n402 585
R355 B.n404 B.n101 585
R356 B.n406 B.n405 585
R357 B.n407 B.n100 585
R358 B.n203 B.n172 585
R359 B.n202 B.n201 585
R360 B.n200 B.n173 585
R361 B.n199 B.n198 585
R362 B.n197 B.n174 585
R363 B.n196 B.n195 585
R364 B.n194 B.n175 585
R365 B.n193 B.n192 585
R366 B.n191 B.n176 585
R367 B.n190 B.n189 585
R368 B.n188 B.n177 585
R369 B.n187 B.n186 585
R370 B.n185 B.n178 585
R371 B.n184 B.n183 585
R372 B.n182 B.n179 585
R373 B.n181 B.n180 585
R374 B.n2 B.n0 585
R375 B.n689 B.n1 585
R376 B.n688 B.n687 585
R377 B.n686 B.n3 585
R378 B.n685 B.n684 585
R379 B.n683 B.n4 585
R380 B.n682 B.n681 585
R381 B.n680 B.n5 585
R382 B.n679 B.n678 585
R383 B.n677 B.n6 585
R384 B.n676 B.n675 585
R385 B.n674 B.n7 585
R386 B.n673 B.n672 585
R387 B.n671 B.n8 585
R388 B.n670 B.n669 585
R389 B.n668 B.n9 585
R390 B.n667 B.n666 585
R391 B.n665 B.n10 585
R392 B.n691 B.n690 585
R393 B.n204 B.n203 482.89
R394 B.n665 B.n664 482.89
R395 B.n408 B.n407 482.89
R396 B.n461 B.n460 482.89
R397 B.n203 B.n202 163.367
R398 B.n202 B.n173 163.367
R399 B.n198 B.n173 163.367
R400 B.n198 B.n197 163.367
R401 B.n197 B.n196 163.367
R402 B.n196 B.n175 163.367
R403 B.n192 B.n175 163.367
R404 B.n192 B.n191 163.367
R405 B.n191 B.n190 163.367
R406 B.n190 B.n177 163.367
R407 B.n186 B.n177 163.367
R408 B.n186 B.n185 163.367
R409 B.n185 B.n184 163.367
R410 B.n184 B.n179 163.367
R411 B.n180 B.n179 163.367
R412 B.n180 B.n2 163.367
R413 B.n690 B.n2 163.367
R414 B.n690 B.n689 163.367
R415 B.n689 B.n688 163.367
R416 B.n688 B.n3 163.367
R417 B.n684 B.n3 163.367
R418 B.n684 B.n683 163.367
R419 B.n683 B.n682 163.367
R420 B.n682 B.n5 163.367
R421 B.n678 B.n5 163.367
R422 B.n678 B.n677 163.367
R423 B.n677 B.n676 163.367
R424 B.n676 B.n7 163.367
R425 B.n672 B.n7 163.367
R426 B.n672 B.n671 163.367
R427 B.n671 B.n670 163.367
R428 B.n670 B.n9 163.367
R429 B.n666 B.n9 163.367
R430 B.n666 B.n665 163.367
R431 B.n204 B.n171 163.367
R432 B.n208 B.n171 163.367
R433 B.n209 B.n208 163.367
R434 B.n210 B.n209 163.367
R435 B.n210 B.n169 163.367
R436 B.n214 B.n169 163.367
R437 B.n215 B.n214 163.367
R438 B.n216 B.n215 163.367
R439 B.n216 B.n167 163.367
R440 B.n220 B.n167 163.367
R441 B.n221 B.n220 163.367
R442 B.n222 B.n221 163.367
R443 B.n222 B.n165 163.367
R444 B.n226 B.n165 163.367
R445 B.n227 B.n226 163.367
R446 B.n228 B.n227 163.367
R447 B.n228 B.n163 163.367
R448 B.n232 B.n163 163.367
R449 B.n233 B.n232 163.367
R450 B.n234 B.n233 163.367
R451 B.n234 B.n161 163.367
R452 B.n238 B.n161 163.367
R453 B.n239 B.n238 163.367
R454 B.n240 B.n239 163.367
R455 B.n240 B.n159 163.367
R456 B.n244 B.n159 163.367
R457 B.n245 B.n244 163.367
R458 B.n246 B.n245 163.367
R459 B.n246 B.n157 163.367
R460 B.n250 B.n157 163.367
R461 B.n251 B.n250 163.367
R462 B.n252 B.n251 163.367
R463 B.n252 B.n155 163.367
R464 B.n256 B.n155 163.367
R465 B.n257 B.n256 163.367
R466 B.n258 B.n257 163.367
R467 B.n258 B.n153 163.367
R468 B.n262 B.n153 163.367
R469 B.n263 B.n262 163.367
R470 B.n264 B.n263 163.367
R471 B.n264 B.n151 163.367
R472 B.n268 B.n151 163.367
R473 B.n269 B.n268 163.367
R474 B.n270 B.n269 163.367
R475 B.n270 B.n149 163.367
R476 B.n274 B.n149 163.367
R477 B.n275 B.n274 163.367
R478 B.n276 B.n275 163.367
R479 B.n276 B.n147 163.367
R480 B.n280 B.n147 163.367
R481 B.n281 B.n280 163.367
R482 B.n282 B.n281 163.367
R483 B.n282 B.n145 163.367
R484 B.n286 B.n145 163.367
R485 B.n287 B.n286 163.367
R486 B.n288 B.n287 163.367
R487 B.n288 B.n143 163.367
R488 B.n292 B.n143 163.367
R489 B.n293 B.n292 163.367
R490 B.n294 B.n293 163.367
R491 B.n294 B.n141 163.367
R492 B.n298 B.n141 163.367
R493 B.n299 B.n298 163.367
R494 B.n299 B.n137 163.367
R495 B.n303 B.n137 163.367
R496 B.n304 B.n303 163.367
R497 B.n305 B.n304 163.367
R498 B.n305 B.n135 163.367
R499 B.n309 B.n135 163.367
R500 B.n310 B.n309 163.367
R501 B.n311 B.n310 163.367
R502 B.n311 B.n131 163.367
R503 B.n316 B.n131 163.367
R504 B.n317 B.n316 163.367
R505 B.n318 B.n317 163.367
R506 B.n318 B.n129 163.367
R507 B.n322 B.n129 163.367
R508 B.n323 B.n322 163.367
R509 B.n324 B.n323 163.367
R510 B.n324 B.n127 163.367
R511 B.n328 B.n127 163.367
R512 B.n329 B.n328 163.367
R513 B.n330 B.n329 163.367
R514 B.n330 B.n125 163.367
R515 B.n334 B.n125 163.367
R516 B.n335 B.n334 163.367
R517 B.n336 B.n335 163.367
R518 B.n336 B.n123 163.367
R519 B.n340 B.n123 163.367
R520 B.n341 B.n340 163.367
R521 B.n342 B.n341 163.367
R522 B.n342 B.n121 163.367
R523 B.n346 B.n121 163.367
R524 B.n347 B.n346 163.367
R525 B.n348 B.n347 163.367
R526 B.n348 B.n119 163.367
R527 B.n352 B.n119 163.367
R528 B.n353 B.n352 163.367
R529 B.n354 B.n353 163.367
R530 B.n354 B.n117 163.367
R531 B.n358 B.n117 163.367
R532 B.n359 B.n358 163.367
R533 B.n360 B.n359 163.367
R534 B.n360 B.n115 163.367
R535 B.n364 B.n115 163.367
R536 B.n365 B.n364 163.367
R537 B.n366 B.n365 163.367
R538 B.n366 B.n113 163.367
R539 B.n370 B.n113 163.367
R540 B.n371 B.n370 163.367
R541 B.n372 B.n371 163.367
R542 B.n372 B.n111 163.367
R543 B.n376 B.n111 163.367
R544 B.n377 B.n376 163.367
R545 B.n378 B.n377 163.367
R546 B.n378 B.n109 163.367
R547 B.n382 B.n109 163.367
R548 B.n383 B.n382 163.367
R549 B.n384 B.n383 163.367
R550 B.n384 B.n107 163.367
R551 B.n388 B.n107 163.367
R552 B.n389 B.n388 163.367
R553 B.n390 B.n389 163.367
R554 B.n390 B.n105 163.367
R555 B.n394 B.n105 163.367
R556 B.n395 B.n394 163.367
R557 B.n396 B.n395 163.367
R558 B.n396 B.n103 163.367
R559 B.n400 B.n103 163.367
R560 B.n401 B.n400 163.367
R561 B.n402 B.n401 163.367
R562 B.n402 B.n101 163.367
R563 B.n406 B.n101 163.367
R564 B.n407 B.n406 163.367
R565 B.n408 B.n99 163.367
R566 B.n412 B.n99 163.367
R567 B.n413 B.n412 163.367
R568 B.n414 B.n413 163.367
R569 B.n414 B.n97 163.367
R570 B.n418 B.n97 163.367
R571 B.n419 B.n418 163.367
R572 B.n420 B.n419 163.367
R573 B.n420 B.n95 163.367
R574 B.n424 B.n95 163.367
R575 B.n425 B.n424 163.367
R576 B.n426 B.n425 163.367
R577 B.n426 B.n93 163.367
R578 B.n430 B.n93 163.367
R579 B.n431 B.n430 163.367
R580 B.n432 B.n431 163.367
R581 B.n432 B.n91 163.367
R582 B.n436 B.n91 163.367
R583 B.n437 B.n436 163.367
R584 B.n438 B.n437 163.367
R585 B.n438 B.n89 163.367
R586 B.n442 B.n89 163.367
R587 B.n443 B.n442 163.367
R588 B.n444 B.n443 163.367
R589 B.n444 B.n87 163.367
R590 B.n448 B.n87 163.367
R591 B.n449 B.n448 163.367
R592 B.n450 B.n449 163.367
R593 B.n450 B.n85 163.367
R594 B.n454 B.n85 163.367
R595 B.n455 B.n454 163.367
R596 B.n456 B.n455 163.367
R597 B.n456 B.n83 163.367
R598 B.n460 B.n83 163.367
R599 B.n664 B.n11 163.367
R600 B.n660 B.n11 163.367
R601 B.n660 B.n659 163.367
R602 B.n659 B.n658 163.367
R603 B.n658 B.n13 163.367
R604 B.n654 B.n13 163.367
R605 B.n654 B.n653 163.367
R606 B.n653 B.n652 163.367
R607 B.n652 B.n15 163.367
R608 B.n648 B.n15 163.367
R609 B.n648 B.n647 163.367
R610 B.n647 B.n646 163.367
R611 B.n646 B.n17 163.367
R612 B.n642 B.n17 163.367
R613 B.n642 B.n641 163.367
R614 B.n641 B.n640 163.367
R615 B.n640 B.n19 163.367
R616 B.n636 B.n19 163.367
R617 B.n636 B.n635 163.367
R618 B.n635 B.n634 163.367
R619 B.n634 B.n21 163.367
R620 B.n630 B.n21 163.367
R621 B.n630 B.n629 163.367
R622 B.n629 B.n628 163.367
R623 B.n628 B.n23 163.367
R624 B.n624 B.n23 163.367
R625 B.n624 B.n623 163.367
R626 B.n623 B.n622 163.367
R627 B.n622 B.n25 163.367
R628 B.n618 B.n25 163.367
R629 B.n618 B.n617 163.367
R630 B.n617 B.n616 163.367
R631 B.n616 B.n27 163.367
R632 B.n612 B.n27 163.367
R633 B.n612 B.n611 163.367
R634 B.n611 B.n610 163.367
R635 B.n610 B.n29 163.367
R636 B.n606 B.n29 163.367
R637 B.n606 B.n605 163.367
R638 B.n605 B.n604 163.367
R639 B.n604 B.n31 163.367
R640 B.n600 B.n31 163.367
R641 B.n600 B.n599 163.367
R642 B.n599 B.n598 163.367
R643 B.n598 B.n33 163.367
R644 B.n594 B.n33 163.367
R645 B.n594 B.n593 163.367
R646 B.n593 B.n592 163.367
R647 B.n592 B.n35 163.367
R648 B.n588 B.n35 163.367
R649 B.n588 B.n587 163.367
R650 B.n587 B.n586 163.367
R651 B.n586 B.n37 163.367
R652 B.n582 B.n37 163.367
R653 B.n582 B.n581 163.367
R654 B.n581 B.n580 163.367
R655 B.n580 B.n39 163.367
R656 B.n576 B.n39 163.367
R657 B.n576 B.n575 163.367
R658 B.n575 B.n574 163.367
R659 B.n574 B.n41 163.367
R660 B.n570 B.n41 163.367
R661 B.n570 B.n569 163.367
R662 B.n569 B.n45 163.367
R663 B.n565 B.n45 163.367
R664 B.n565 B.n564 163.367
R665 B.n564 B.n563 163.367
R666 B.n563 B.n47 163.367
R667 B.n559 B.n47 163.367
R668 B.n559 B.n558 163.367
R669 B.n558 B.n557 163.367
R670 B.n557 B.n49 163.367
R671 B.n552 B.n49 163.367
R672 B.n552 B.n551 163.367
R673 B.n551 B.n550 163.367
R674 B.n550 B.n53 163.367
R675 B.n546 B.n53 163.367
R676 B.n546 B.n545 163.367
R677 B.n545 B.n544 163.367
R678 B.n544 B.n55 163.367
R679 B.n540 B.n55 163.367
R680 B.n540 B.n539 163.367
R681 B.n539 B.n538 163.367
R682 B.n538 B.n57 163.367
R683 B.n534 B.n57 163.367
R684 B.n534 B.n533 163.367
R685 B.n533 B.n532 163.367
R686 B.n532 B.n59 163.367
R687 B.n528 B.n59 163.367
R688 B.n528 B.n527 163.367
R689 B.n527 B.n526 163.367
R690 B.n526 B.n61 163.367
R691 B.n522 B.n61 163.367
R692 B.n522 B.n521 163.367
R693 B.n521 B.n520 163.367
R694 B.n520 B.n63 163.367
R695 B.n516 B.n63 163.367
R696 B.n516 B.n515 163.367
R697 B.n515 B.n514 163.367
R698 B.n514 B.n65 163.367
R699 B.n510 B.n65 163.367
R700 B.n510 B.n509 163.367
R701 B.n509 B.n508 163.367
R702 B.n508 B.n67 163.367
R703 B.n504 B.n67 163.367
R704 B.n504 B.n503 163.367
R705 B.n503 B.n502 163.367
R706 B.n502 B.n69 163.367
R707 B.n498 B.n69 163.367
R708 B.n498 B.n497 163.367
R709 B.n497 B.n496 163.367
R710 B.n496 B.n71 163.367
R711 B.n492 B.n71 163.367
R712 B.n492 B.n491 163.367
R713 B.n491 B.n490 163.367
R714 B.n490 B.n73 163.367
R715 B.n486 B.n73 163.367
R716 B.n486 B.n485 163.367
R717 B.n485 B.n484 163.367
R718 B.n484 B.n75 163.367
R719 B.n480 B.n75 163.367
R720 B.n480 B.n479 163.367
R721 B.n479 B.n478 163.367
R722 B.n478 B.n77 163.367
R723 B.n474 B.n77 163.367
R724 B.n474 B.n473 163.367
R725 B.n473 B.n472 163.367
R726 B.n472 B.n79 163.367
R727 B.n468 B.n79 163.367
R728 B.n468 B.n467 163.367
R729 B.n467 B.n466 163.367
R730 B.n466 B.n81 163.367
R731 B.n462 B.n81 163.367
R732 B.n462 B.n461 163.367
R733 B.n132 B.t11 127.433
R734 B.n50 B.t1 127.433
R735 B.n138 B.t5 127.407
R736 B.n42 B.t7 127.407
R737 B.n133 B.t10 107.844
R738 B.n51 B.t2 107.844
R739 B.n139 B.t4 107.82
R740 B.n43 B.t8 107.82
R741 B.n313 B.n133 59.5399
R742 B.n140 B.n139 59.5399
R743 B.n44 B.n43 59.5399
R744 B.n555 B.n51 59.5399
R745 B.n663 B.n10 31.3761
R746 B.n459 B.n82 31.3761
R747 B.n409 B.n100 31.3761
R748 B.n205 B.n172 31.3761
R749 B.n133 B.n132 19.5884
R750 B.n139 B.n138 19.5884
R751 B.n43 B.n42 19.5884
R752 B.n51 B.n50 19.5884
R753 B B.n691 18.0485
R754 B.n663 B.n662 10.6151
R755 B.n662 B.n661 10.6151
R756 B.n661 B.n12 10.6151
R757 B.n657 B.n12 10.6151
R758 B.n657 B.n656 10.6151
R759 B.n656 B.n655 10.6151
R760 B.n655 B.n14 10.6151
R761 B.n651 B.n14 10.6151
R762 B.n651 B.n650 10.6151
R763 B.n650 B.n649 10.6151
R764 B.n649 B.n16 10.6151
R765 B.n645 B.n16 10.6151
R766 B.n645 B.n644 10.6151
R767 B.n644 B.n643 10.6151
R768 B.n643 B.n18 10.6151
R769 B.n639 B.n18 10.6151
R770 B.n639 B.n638 10.6151
R771 B.n638 B.n637 10.6151
R772 B.n637 B.n20 10.6151
R773 B.n633 B.n20 10.6151
R774 B.n633 B.n632 10.6151
R775 B.n632 B.n631 10.6151
R776 B.n631 B.n22 10.6151
R777 B.n627 B.n22 10.6151
R778 B.n627 B.n626 10.6151
R779 B.n626 B.n625 10.6151
R780 B.n625 B.n24 10.6151
R781 B.n621 B.n24 10.6151
R782 B.n621 B.n620 10.6151
R783 B.n620 B.n619 10.6151
R784 B.n619 B.n26 10.6151
R785 B.n615 B.n26 10.6151
R786 B.n615 B.n614 10.6151
R787 B.n614 B.n613 10.6151
R788 B.n613 B.n28 10.6151
R789 B.n609 B.n28 10.6151
R790 B.n609 B.n608 10.6151
R791 B.n608 B.n607 10.6151
R792 B.n607 B.n30 10.6151
R793 B.n603 B.n30 10.6151
R794 B.n603 B.n602 10.6151
R795 B.n602 B.n601 10.6151
R796 B.n601 B.n32 10.6151
R797 B.n597 B.n32 10.6151
R798 B.n597 B.n596 10.6151
R799 B.n596 B.n595 10.6151
R800 B.n595 B.n34 10.6151
R801 B.n591 B.n34 10.6151
R802 B.n591 B.n590 10.6151
R803 B.n590 B.n589 10.6151
R804 B.n589 B.n36 10.6151
R805 B.n585 B.n36 10.6151
R806 B.n585 B.n584 10.6151
R807 B.n584 B.n583 10.6151
R808 B.n583 B.n38 10.6151
R809 B.n579 B.n38 10.6151
R810 B.n579 B.n578 10.6151
R811 B.n578 B.n577 10.6151
R812 B.n577 B.n40 10.6151
R813 B.n573 B.n40 10.6151
R814 B.n573 B.n572 10.6151
R815 B.n572 B.n571 10.6151
R816 B.n568 B.n567 10.6151
R817 B.n567 B.n566 10.6151
R818 B.n566 B.n46 10.6151
R819 B.n562 B.n46 10.6151
R820 B.n562 B.n561 10.6151
R821 B.n561 B.n560 10.6151
R822 B.n560 B.n48 10.6151
R823 B.n556 B.n48 10.6151
R824 B.n554 B.n553 10.6151
R825 B.n553 B.n52 10.6151
R826 B.n549 B.n52 10.6151
R827 B.n549 B.n548 10.6151
R828 B.n548 B.n547 10.6151
R829 B.n547 B.n54 10.6151
R830 B.n543 B.n54 10.6151
R831 B.n543 B.n542 10.6151
R832 B.n542 B.n541 10.6151
R833 B.n541 B.n56 10.6151
R834 B.n537 B.n56 10.6151
R835 B.n537 B.n536 10.6151
R836 B.n536 B.n535 10.6151
R837 B.n535 B.n58 10.6151
R838 B.n531 B.n58 10.6151
R839 B.n531 B.n530 10.6151
R840 B.n530 B.n529 10.6151
R841 B.n529 B.n60 10.6151
R842 B.n525 B.n60 10.6151
R843 B.n525 B.n524 10.6151
R844 B.n524 B.n523 10.6151
R845 B.n523 B.n62 10.6151
R846 B.n519 B.n62 10.6151
R847 B.n519 B.n518 10.6151
R848 B.n518 B.n517 10.6151
R849 B.n517 B.n64 10.6151
R850 B.n513 B.n64 10.6151
R851 B.n513 B.n512 10.6151
R852 B.n512 B.n511 10.6151
R853 B.n511 B.n66 10.6151
R854 B.n507 B.n66 10.6151
R855 B.n507 B.n506 10.6151
R856 B.n506 B.n505 10.6151
R857 B.n505 B.n68 10.6151
R858 B.n501 B.n68 10.6151
R859 B.n501 B.n500 10.6151
R860 B.n500 B.n499 10.6151
R861 B.n499 B.n70 10.6151
R862 B.n495 B.n70 10.6151
R863 B.n495 B.n494 10.6151
R864 B.n494 B.n493 10.6151
R865 B.n493 B.n72 10.6151
R866 B.n489 B.n72 10.6151
R867 B.n489 B.n488 10.6151
R868 B.n488 B.n487 10.6151
R869 B.n487 B.n74 10.6151
R870 B.n483 B.n74 10.6151
R871 B.n483 B.n482 10.6151
R872 B.n482 B.n481 10.6151
R873 B.n481 B.n76 10.6151
R874 B.n477 B.n76 10.6151
R875 B.n477 B.n476 10.6151
R876 B.n476 B.n475 10.6151
R877 B.n475 B.n78 10.6151
R878 B.n471 B.n78 10.6151
R879 B.n471 B.n470 10.6151
R880 B.n470 B.n469 10.6151
R881 B.n469 B.n80 10.6151
R882 B.n465 B.n80 10.6151
R883 B.n465 B.n464 10.6151
R884 B.n464 B.n463 10.6151
R885 B.n463 B.n82 10.6151
R886 B.n410 B.n409 10.6151
R887 B.n411 B.n410 10.6151
R888 B.n411 B.n98 10.6151
R889 B.n415 B.n98 10.6151
R890 B.n416 B.n415 10.6151
R891 B.n417 B.n416 10.6151
R892 B.n417 B.n96 10.6151
R893 B.n421 B.n96 10.6151
R894 B.n422 B.n421 10.6151
R895 B.n423 B.n422 10.6151
R896 B.n423 B.n94 10.6151
R897 B.n427 B.n94 10.6151
R898 B.n428 B.n427 10.6151
R899 B.n429 B.n428 10.6151
R900 B.n429 B.n92 10.6151
R901 B.n433 B.n92 10.6151
R902 B.n434 B.n433 10.6151
R903 B.n435 B.n434 10.6151
R904 B.n435 B.n90 10.6151
R905 B.n439 B.n90 10.6151
R906 B.n440 B.n439 10.6151
R907 B.n441 B.n440 10.6151
R908 B.n441 B.n88 10.6151
R909 B.n445 B.n88 10.6151
R910 B.n446 B.n445 10.6151
R911 B.n447 B.n446 10.6151
R912 B.n447 B.n86 10.6151
R913 B.n451 B.n86 10.6151
R914 B.n452 B.n451 10.6151
R915 B.n453 B.n452 10.6151
R916 B.n453 B.n84 10.6151
R917 B.n457 B.n84 10.6151
R918 B.n458 B.n457 10.6151
R919 B.n459 B.n458 10.6151
R920 B.n206 B.n205 10.6151
R921 B.n207 B.n206 10.6151
R922 B.n207 B.n170 10.6151
R923 B.n211 B.n170 10.6151
R924 B.n212 B.n211 10.6151
R925 B.n213 B.n212 10.6151
R926 B.n213 B.n168 10.6151
R927 B.n217 B.n168 10.6151
R928 B.n218 B.n217 10.6151
R929 B.n219 B.n218 10.6151
R930 B.n219 B.n166 10.6151
R931 B.n223 B.n166 10.6151
R932 B.n224 B.n223 10.6151
R933 B.n225 B.n224 10.6151
R934 B.n225 B.n164 10.6151
R935 B.n229 B.n164 10.6151
R936 B.n230 B.n229 10.6151
R937 B.n231 B.n230 10.6151
R938 B.n231 B.n162 10.6151
R939 B.n235 B.n162 10.6151
R940 B.n236 B.n235 10.6151
R941 B.n237 B.n236 10.6151
R942 B.n237 B.n160 10.6151
R943 B.n241 B.n160 10.6151
R944 B.n242 B.n241 10.6151
R945 B.n243 B.n242 10.6151
R946 B.n243 B.n158 10.6151
R947 B.n247 B.n158 10.6151
R948 B.n248 B.n247 10.6151
R949 B.n249 B.n248 10.6151
R950 B.n249 B.n156 10.6151
R951 B.n253 B.n156 10.6151
R952 B.n254 B.n253 10.6151
R953 B.n255 B.n254 10.6151
R954 B.n255 B.n154 10.6151
R955 B.n259 B.n154 10.6151
R956 B.n260 B.n259 10.6151
R957 B.n261 B.n260 10.6151
R958 B.n261 B.n152 10.6151
R959 B.n265 B.n152 10.6151
R960 B.n266 B.n265 10.6151
R961 B.n267 B.n266 10.6151
R962 B.n267 B.n150 10.6151
R963 B.n271 B.n150 10.6151
R964 B.n272 B.n271 10.6151
R965 B.n273 B.n272 10.6151
R966 B.n273 B.n148 10.6151
R967 B.n277 B.n148 10.6151
R968 B.n278 B.n277 10.6151
R969 B.n279 B.n278 10.6151
R970 B.n279 B.n146 10.6151
R971 B.n283 B.n146 10.6151
R972 B.n284 B.n283 10.6151
R973 B.n285 B.n284 10.6151
R974 B.n285 B.n144 10.6151
R975 B.n289 B.n144 10.6151
R976 B.n290 B.n289 10.6151
R977 B.n291 B.n290 10.6151
R978 B.n291 B.n142 10.6151
R979 B.n295 B.n142 10.6151
R980 B.n296 B.n295 10.6151
R981 B.n297 B.n296 10.6151
R982 B.n301 B.n300 10.6151
R983 B.n302 B.n301 10.6151
R984 B.n302 B.n136 10.6151
R985 B.n306 B.n136 10.6151
R986 B.n307 B.n306 10.6151
R987 B.n308 B.n307 10.6151
R988 B.n308 B.n134 10.6151
R989 B.n312 B.n134 10.6151
R990 B.n315 B.n314 10.6151
R991 B.n315 B.n130 10.6151
R992 B.n319 B.n130 10.6151
R993 B.n320 B.n319 10.6151
R994 B.n321 B.n320 10.6151
R995 B.n321 B.n128 10.6151
R996 B.n325 B.n128 10.6151
R997 B.n326 B.n325 10.6151
R998 B.n327 B.n326 10.6151
R999 B.n327 B.n126 10.6151
R1000 B.n331 B.n126 10.6151
R1001 B.n332 B.n331 10.6151
R1002 B.n333 B.n332 10.6151
R1003 B.n333 B.n124 10.6151
R1004 B.n337 B.n124 10.6151
R1005 B.n338 B.n337 10.6151
R1006 B.n339 B.n338 10.6151
R1007 B.n339 B.n122 10.6151
R1008 B.n343 B.n122 10.6151
R1009 B.n344 B.n343 10.6151
R1010 B.n345 B.n344 10.6151
R1011 B.n345 B.n120 10.6151
R1012 B.n349 B.n120 10.6151
R1013 B.n350 B.n349 10.6151
R1014 B.n351 B.n350 10.6151
R1015 B.n351 B.n118 10.6151
R1016 B.n355 B.n118 10.6151
R1017 B.n356 B.n355 10.6151
R1018 B.n357 B.n356 10.6151
R1019 B.n357 B.n116 10.6151
R1020 B.n361 B.n116 10.6151
R1021 B.n362 B.n361 10.6151
R1022 B.n363 B.n362 10.6151
R1023 B.n363 B.n114 10.6151
R1024 B.n367 B.n114 10.6151
R1025 B.n368 B.n367 10.6151
R1026 B.n369 B.n368 10.6151
R1027 B.n369 B.n112 10.6151
R1028 B.n373 B.n112 10.6151
R1029 B.n374 B.n373 10.6151
R1030 B.n375 B.n374 10.6151
R1031 B.n375 B.n110 10.6151
R1032 B.n379 B.n110 10.6151
R1033 B.n380 B.n379 10.6151
R1034 B.n381 B.n380 10.6151
R1035 B.n381 B.n108 10.6151
R1036 B.n385 B.n108 10.6151
R1037 B.n386 B.n385 10.6151
R1038 B.n387 B.n386 10.6151
R1039 B.n387 B.n106 10.6151
R1040 B.n391 B.n106 10.6151
R1041 B.n392 B.n391 10.6151
R1042 B.n393 B.n392 10.6151
R1043 B.n393 B.n104 10.6151
R1044 B.n397 B.n104 10.6151
R1045 B.n398 B.n397 10.6151
R1046 B.n399 B.n398 10.6151
R1047 B.n399 B.n102 10.6151
R1048 B.n403 B.n102 10.6151
R1049 B.n404 B.n403 10.6151
R1050 B.n405 B.n404 10.6151
R1051 B.n405 B.n100 10.6151
R1052 B.n201 B.n172 10.6151
R1053 B.n201 B.n200 10.6151
R1054 B.n200 B.n199 10.6151
R1055 B.n199 B.n174 10.6151
R1056 B.n195 B.n174 10.6151
R1057 B.n195 B.n194 10.6151
R1058 B.n194 B.n193 10.6151
R1059 B.n193 B.n176 10.6151
R1060 B.n189 B.n176 10.6151
R1061 B.n189 B.n188 10.6151
R1062 B.n188 B.n187 10.6151
R1063 B.n187 B.n178 10.6151
R1064 B.n183 B.n178 10.6151
R1065 B.n183 B.n182 10.6151
R1066 B.n182 B.n181 10.6151
R1067 B.n181 B.n0 10.6151
R1068 B.n687 B.n1 10.6151
R1069 B.n687 B.n686 10.6151
R1070 B.n686 B.n685 10.6151
R1071 B.n685 B.n4 10.6151
R1072 B.n681 B.n4 10.6151
R1073 B.n681 B.n680 10.6151
R1074 B.n680 B.n679 10.6151
R1075 B.n679 B.n6 10.6151
R1076 B.n675 B.n6 10.6151
R1077 B.n675 B.n674 10.6151
R1078 B.n674 B.n673 10.6151
R1079 B.n673 B.n8 10.6151
R1080 B.n669 B.n8 10.6151
R1081 B.n669 B.n668 10.6151
R1082 B.n668 B.n667 10.6151
R1083 B.n667 B.n10 10.6151
R1084 B.n568 B.n44 6.5566
R1085 B.n556 B.n555 6.5566
R1086 B.n300 B.n140 6.5566
R1087 B.n313 B.n312 6.5566
R1088 B.n571 B.n44 4.05904
R1089 B.n555 B.n554 4.05904
R1090 B.n297 B.n140 4.05904
R1091 B.n314 B.n313 4.05904
R1092 B.n691 B.n0 2.81026
R1093 B.n691 B.n1 2.81026
C0 VTAIL B 5.71759f
C1 w_n1576_n4794# VDD2 1.26174f
C2 w_n1576_n4794# VP 2.65455f
C3 VN VDD2 4.8071f
C4 VDD1 w_n1576_n4794# 1.24762f
C5 VN VP 6.13059f
C6 VDD1 VN 0.147071f
C7 VTAIL VDD2 10.1113f
C8 B VDD2 1.13586f
C9 VTAIL VP 4.13114f
C10 VDD1 VTAIL 10.070001f
C11 B VP 1.14539f
C12 VDD1 B 1.11461f
C13 w_n1576_n4794# VN 2.4568f
C14 VP VDD2 0.271938f
C15 VDD1 VDD2 0.561847f
C16 VTAIL w_n1576_n4794# 5.93415f
C17 VDD1 VP 4.93172f
C18 B w_n1576_n4794# 8.88196f
C19 VTAIL VN 4.11703f
C20 B VN 0.826178f
C21 VDD2 VSUBS 0.847906f
C22 VDD1 VSUBS 6.029587f
C23 VTAIL VSUBS 1.142922f
C24 VN VSUBS 6.500411f
C25 VP VSUBS 1.542894f
C26 B VSUBS 3.205618f
C27 w_n1576_n4794# VSUBS 92.3095f
C28 B.n0 VSUBS 0.00486f
C29 B.n1 VSUBS 0.00486f
C30 B.n2 VSUBS 0.007686f
C31 B.n3 VSUBS 0.007686f
C32 B.n4 VSUBS 0.007686f
C33 B.n5 VSUBS 0.007686f
C34 B.n6 VSUBS 0.007686f
C35 B.n7 VSUBS 0.007686f
C36 B.n8 VSUBS 0.007686f
C37 B.n9 VSUBS 0.007686f
C38 B.n10 VSUBS 0.016955f
C39 B.n11 VSUBS 0.007686f
C40 B.n12 VSUBS 0.007686f
C41 B.n13 VSUBS 0.007686f
C42 B.n14 VSUBS 0.007686f
C43 B.n15 VSUBS 0.007686f
C44 B.n16 VSUBS 0.007686f
C45 B.n17 VSUBS 0.007686f
C46 B.n18 VSUBS 0.007686f
C47 B.n19 VSUBS 0.007686f
C48 B.n20 VSUBS 0.007686f
C49 B.n21 VSUBS 0.007686f
C50 B.n22 VSUBS 0.007686f
C51 B.n23 VSUBS 0.007686f
C52 B.n24 VSUBS 0.007686f
C53 B.n25 VSUBS 0.007686f
C54 B.n26 VSUBS 0.007686f
C55 B.n27 VSUBS 0.007686f
C56 B.n28 VSUBS 0.007686f
C57 B.n29 VSUBS 0.007686f
C58 B.n30 VSUBS 0.007686f
C59 B.n31 VSUBS 0.007686f
C60 B.n32 VSUBS 0.007686f
C61 B.n33 VSUBS 0.007686f
C62 B.n34 VSUBS 0.007686f
C63 B.n35 VSUBS 0.007686f
C64 B.n36 VSUBS 0.007686f
C65 B.n37 VSUBS 0.007686f
C66 B.n38 VSUBS 0.007686f
C67 B.n39 VSUBS 0.007686f
C68 B.n40 VSUBS 0.007686f
C69 B.n41 VSUBS 0.007686f
C70 B.t8 VSUBS 0.712045f
C71 B.t7 VSUBS 0.7212f
C72 B.t6 VSUBS 0.573064f
C73 B.n42 VSUBS 0.209775f
C74 B.n43 VSUBS 0.070511f
C75 B.n44 VSUBS 0.017808f
C76 B.n45 VSUBS 0.007686f
C77 B.n46 VSUBS 0.007686f
C78 B.n47 VSUBS 0.007686f
C79 B.n48 VSUBS 0.007686f
C80 B.n49 VSUBS 0.007686f
C81 B.t2 VSUBS 0.712016f
C82 B.t1 VSUBS 0.721174f
C83 B.t0 VSUBS 0.573064f
C84 B.n50 VSUBS 0.209802f
C85 B.n51 VSUBS 0.07054f
C86 B.n52 VSUBS 0.007686f
C87 B.n53 VSUBS 0.007686f
C88 B.n54 VSUBS 0.007686f
C89 B.n55 VSUBS 0.007686f
C90 B.n56 VSUBS 0.007686f
C91 B.n57 VSUBS 0.007686f
C92 B.n58 VSUBS 0.007686f
C93 B.n59 VSUBS 0.007686f
C94 B.n60 VSUBS 0.007686f
C95 B.n61 VSUBS 0.007686f
C96 B.n62 VSUBS 0.007686f
C97 B.n63 VSUBS 0.007686f
C98 B.n64 VSUBS 0.007686f
C99 B.n65 VSUBS 0.007686f
C100 B.n66 VSUBS 0.007686f
C101 B.n67 VSUBS 0.007686f
C102 B.n68 VSUBS 0.007686f
C103 B.n69 VSUBS 0.007686f
C104 B.n70 VSUBS 0.007686f
C105 B.n71 VSUBS 0.007686f
C106 B.n72 VSUBS 0.007686f
C107 B.n73 VSUBS 0.007686f
C108 B.n74 VSUBS 0.007686f
C109 B.n75 VSUBS 0.007686f
C110 B.n76 VSUBS 0.007686f
C111 B.n77 VSUBS 0.007686f
C112 B.n78 VSUBS 0.007686f
C113 B.n79 VSUBS 0.007686f
C114 B.n80 VSUBS 0.007686f
C115 B.n81 VSUBS 0.007686f
C116 B.n82 VSUBS 0.01714f
C117 B.n83 VSUBS 0.007686f
C118 B.n84 VSUBS 0.007686f
C119 B.n85 VSUBS 0.007686f
C120 B.n86 VSUBS 0.007686f
C121 B.n87 VSUBS 0.007686f
C122 B.n88 VSUBS 0.007686f
C123 B.n89 VSUBS 0.007686f
C124 B.n90 VSUBS 0.007686f
C125 B.n91 VSUBS 0.007686f
C126 B.n92 VSUBS 0.007686f
C127 B.n93 VSUBS 0.007686f
C128 B.n94 VSUBS 0.007686f
C129 B.n95 VSUBS 0.007686f
C130 B.n96 VSUBS 0.007686f
C131 B.n97 VSUBS 0.007686f
C132 B.n98 VSUBS 0.007686f
C133 B.n99 VSUBS 0.007686f
C134 B.n100 VSUBS 0.018085f
C135 B.n101 VSUBS 0.007686f
C136 B.n102 VSUBS 0.007686f
C137 B.n103 VSUBS 0.007686f
C138 B.n104 VSUBS 0.007686f
C139 B.n105 VSUBS 0.007686f
C140 B.n106 VSUBS 0.007686f
C141 B.n107 VSUBS 0.007686f
C142 B.n108 VSUBS 0.007686f
C143 B.n109 VSUBS 0.007686f
C144 B.n110 VSUBS 0.007686f
C145 B.n111 VSUBS 0.007686f
C146 B.n112 VSUBS 0.007686f
C147 B.n113 VSUBS 0.007686f
C148 B.n114 VSUBS 0.007686f
C149 B.n115 VSUBS 0.007686f
C150 B.n116 VSUBS 0.007686f
C151 B.n117 VSUBS 0.007686f
C152 B.n118 VSUBS 0.007686f
C153 B.n119 VSUBS 0.007686f
C154 B.n120 VSUBS 0.007686f
C155 B.n121 VSUBS 0.007686f
C156 B.n122 VSUBS 0.007686f
C157 B.n123 VSUBS 0.007686f
C158 B.n124 VSUBS 0.007686f
C159 B.n125 VSUBS 0.007686f
C160 B.n126 VSUBS 0.007686f
C161 B.n127 VSUBS 0.007686f
C162 B.n128 VSUBS 0.007686f
C163 B.n129 VSUBS 0.007686f
C164 B.n130 VSUBS 0.007686f
C165 B.n131 VSUBS 0.007686f
C166 B.t10 VSUBS 0.712016f
C167 B.t11 VSUBS 0.721174f
C168 B.t9 VSUBS 0.573064f
C169 B.n132 VSUBS 0.209802f
C170 B.n133 VSUBS 0.07054f
C171 B.n134 VSUBS 0.007686f
C172 B.n135 VSUBS 0.007686f
C173 B.n136 VSUBS 0.007686f
C174 B.n137 VSUBS 0.007686f
C175 B.t4 VSUBS 0.712045f
C176 B.t5 VSUBS 0.7212f
C177 B.t3 VSUBS 0.573064f
C178 B.n138 VSUBS 0.209775f
C179 B.n139 VSUBS 0.070511f
C180 B.n140 VSUBS 0.017808f
C181 B.n141 VSUBS 0.007686f
C182 B.n142 VSUBS 0.007686f
C183 B.n143 VSUBS 0.007686f
C184 B.n144 VSUBS 0.007686f
C185 B.n145 VSUBS 0.007686f
C186 B.n146 VSUBS 0.007686f
C187 B.n147 VSUBS 0.007686f
C188 B.n148 VSUBS 0.007686f
C189 B.n149 VSUBS 0.007686f
C190 B.n150 VSUBS 0.007686f
C191 B.n151 VSUBS 0.007686f
C192 B.n152 VSUBS 0.007686f
C193 B.n153 VSUBS 0.007686f
C194 B.n154 VSUBS 0.007686f
C195 B.n155 VSUBS 0.007686f
C196 B.n156 VSUBS 0.007686f
C197 B.n157 VSUBS 0.007686f
C198 B.n158 VSUBS 0.007686f
C199 B.n159 VSUBS 0.007686f
C200 B.n160 VSUBS 0.007686f
C201 B.n161 VSUBS 0.007686f
C202 B.n162 VSUBS 0.007686f
C203 B.n163 VSUBS 0.007686f
C204 B.n164 VSUBS 0.007686f
C205 B.n165 VSUBS 0.007686f
C206 B.n166 VSUBS 0.007686f
C207 B.n167 VSUBS 0.007686f
C208 B.n168 VSUBS 0.007686f
C209 B.n169 VSUBS 0.007686f
C210 B.n170 VSUBS 0.007686f
C211 B.n171 VSUBS 0.007686f
C212 B.n172 VSUBS 0.016955f
C213 B.n173 VSUBS 0.007686f
C214 B.n174 VSUBS 0.007686f
C215 B.n175 VSUBS 0.007686f
C216 B.n176 VSUBS 0.007686f
C217 B.n177 VSUBS 0.007686f
C218 B.n178 VSUBS 0.007686f
C219 B.n179 VSUBS 0.007686f
C220 B.n180 VSUBS 0.007686f
C221 B.n181 VSUBS 0.007686f
C222 B.n182 VSUBS 0.007686f
C223 B.n183 VSUBS 0.007686f
C224 B.n184 VSUBS 0.007686f
C225 B.n185 VSUBS 0.007686f
C226 B.n186 VSUBS 0.007686f
C227 B.n187 VSUBS 0.007686f
C228 B.n188 VSUBS 0.007686f
C229 B.n189 VSUBS 0.007686f
C230 B.n190 VSUBS 0.007686f
C231 B.n191 VSUBS 0.007686f
C232 B.n192 VSUBS 0.007686f
C233 B.n193 VSUBS 0.007686f
C234 B.n194 VSUBS 0.007686f
C235 B.n195 VSUBS 0.007686f
C236 B.n196 VSUBS 0.007686f
C237 B.n197 VSUBS 0.007686f
C238 B.n198 VSUBS 0.007686f
C239 B.n199 VSUBS 0.007686f
C240 B.n200 VSUBS 0.007686f
C241 B.n201 VSUBS 0.007686f
C242 B.n202 VSUBS 0.007686f
C243 B.n203 VSUBS 0.016955f
C244 B.n204 VSUBS 0.018085f
C245 B.n205 VSUBS 0.018085f
C246 B.n206 VSUBS 0.007686f
C247 B.n207 VSUBS 0.007686f
C248 B.n208 VSUBS 0.007686f
C249 B.n209 VSUBS 0.007686f
C250 B.n210 VSUBS 0.007686f
C251 B.n211 VSUBS 0.007686f
C252 B.n212 VSUBS 0.007686f
C253 B.n213 VSUBS 0.007686f
C254 B.n214 VSUBS 0.007686f
C255 B.n215 VSUBS 0.007686f
C256 B.n216 VSUBS 0.007686f
C257 B.n217 VSUBS 0.007686f
C258 B.n218 VSUBS 0.007686f
C259 B.n219 VSUBS 0.007686f
C260 B.n220 VSUBS 0.007686f
C261 B.n221 VSUBS 0.007686f
C262 B.n222 VSUBS 0.007686f
C263 B.n223 VSUBS 0.007686f
C264 B.n224 VSUBS 0.007686f
C265 B.n225 VSUBS 0.007686f
C266 B.n226 VSUBS 0.007686f
C267 B.n227 VSUBS 0.007686f
C268 B.n228 VSUBS 0.007686f
C269 B.n229 VSUBS 0.007686f
C270 B.n230 VSUBS 0.007686f
C271 B.n231 VSUBS 0.007686f
C272 B.n232 VSUBS 0.007686f
C273 B.n233 VSUBS 0.007686f
C274 B.n234 VSUBS 0.007686f
C275 B.n235 VSUBS 0.007686f
C276 B.n236 VSUBS 0.007686f
C277 B.n237 VSUBS 0.007686f
C278 B.n238 VSUBS 0.007686f
C279 B.n239 VSUBS 0.007686f
C280 B.n240 VSUBS 0.007686f
C281 B.n241 VSUBS 0.007686f
C282 B.n242 VSUBS 0.007686f
C283 B.n243 VSUBS 0.007686f
C284 B.n244 VSUBS 0.007686f
C285 B.n245 VSUBS 0.007686f
C286 B.n246 VSUBS 0.007686f
C287 B.n247 VSUBS 0.007686f
C288 B.n248 VSUBS 0.007686f
C289 B.n249 VSUBS 0.007686f
C290 B.n250 VSUBS 0.007686f
C291 B.n251 VSUBS 0.007686f
C292 B.n252 VSUBS 0.007686f
C293 B.n253 VSUBS 0.007686f
C294 B.n254 VSUBS 0.007686f
C295 B.n255 VSUBS 0.007686f
C296 B.n256 VSUBS 0.007686f
C297 B.n257 VSUBS 0.007686f
C298 B.n258 VSUBS 0.007686f
C299 B.n259 VSUBS 0.007686f
C300 B.n260 VSUBS 0.007686f
C301 B.n261 VSUBS 0.007686f
C302 B.n262 VSUBS 0.007686f
C303 B.n263 VSUBS 0.007686f
C304 B.n264 VSUBS 0.007686f
C305 B.n265 VSUBS 0.007686f
C306 B.n266 VSUBS 0.007686f
C307 B.n267 VSUBS 0.007686f
C308 B.n268 VSUBS 0.007686f
C309 B.n269 VSUBS 0.007686f
C310 B.n270 VSUBS 0.007686f
C311 B.n271 VSUBS 0.007686f
C312 B.n272 VSUBS 0.007686f
C313 B.n273 VSUBS 0.007686f
C314 B.n274 VSUBS 0.007686f
C315 B.n275 VSUBS 0.007686f
C316 B.n276 VSUBS 0.007686f
C317 B.n277 VSUBS 0.007686f
C318 B.n278 VSUBS 0.007686f
C319 B.n279 VSUBS 0.007686f
C320 B.n280 VSUBS 0.007686f
C321 B.n281 VSUBS 0.007686f
C322 B.n282 VSUBS 0.007686f
C323 B.n283 VSUBS 0.007686f
C324 B.n284 VSUBS 0.007686f
C325 B.n285 VSUBS 0.007686f
C326 B.n286 VSUBS 0.007686f
C327 B.n287 VSUBS 0.007686f
C328 B.n288 VSUBS 0.007686f
C329 B.n289 VSUBS 0.007686f
C330 B.n290 VSUBS 0.007686f
C331 B.n291 VSUBS 0.007686f
C332 B.n292 VSUBS 0.007686f
C333 B.n293 VSUBS 0.007686f
C334 B.n294 VSUBS 0.007686f
C335 B.n295 VSUBS 0.007686f
C336 B.n296 VSUBS 0.007686f
C337 B.n297 VSUBS 0.005313f
C338 B.n298 VSUBS 0.007686f
C339 B.n299 VSUBS 0.007686f
C340 B.n300 VSUBS 0.006217f
C341 B.n301 VSUBS 0.007686f
C342 B.n302 VSUBS 0.007686f
C343 B.n303 VSUBS 0.007686f
C344 B.n304 VSUBS 0.007686f
C345 B.n305 VSUBS 0.007686f
C346 B.n306 VSUBS 0.007686f
C347 B.n307 VSUBS 0.007686f
C348 B.n308 VSUBS 0.007686f
C349 B.n309 VSUBS 0.007686f
C350 B.n310 VSUBS 0.007686f
C351 B.n311 VSUBS 0.007686f
C352 B.n312 VSUBS 0.006217f
C353 B.n313 VSUBS 0.017808f
C354 B.n314 VSUBS 0.005313f
C355 B.n315 VSUBS 0.007686f
C356 B.n316 VSUBS 0.007686f
C357 B.n317 VSUBS 0.007686f
C358 B.n318 VSUBS 0.007686f
C359 B.n319 VSUBS 0.007686f
C360 B.n320 VSUBS 0.007686f
C361 B.n321 VSUBS 0.007686f
C362 B.n322 VSUBS 0.007686f
C363 B.n323 VSUBS 0.007686f
C364 B.n324 VSUBS 0.007686f
C365 B.n325 VSUBS 0.007686f
C366 B.n326 VSUBS 0.007686f
C367 B.n327 VSUBS 0.007686f
C368 B.n328 VSUBS 0.007686f
C369 B.n329 VSUBS 0.007686f
C370 B.n330 VSUBS 0.007686f
C371 B.n331 VSUBS 0.007686f
C372 B.n332 VSUBS 0.007686f
C373 B.n333 VSUBS 0.007686f
C374 B.n334 VSUBS 0.007686f
C375 B.n335 VSUBS 0.007686f
C376 B.n336 VSUBS 0.007686f
C377 B.n337 VSUBS 0.007686f
C378 B.n338 VSUBS 0.007686f
C379 B.n339 VSUBS 0.007686f
C380 B.n340 VSUBS 0.007686f
C381 B.n341 VSUBS 0.007686f
C382 B.n342 VSUBS 0.007686f
C383 B.n343 VSUBS 0.007686f
C384 B.n344 VSUBS 0.007686f
C385 B.n345 VSUBS 0.007686f
C386 B.n346 VSUBS 0.007686f
C387 B.n347 VSUBS 0.007686f
C388 B.n348 VSUBS 0.007686f
C389 B.n349 VSUBS 0.007686f
C390 B.n350 VSUBS 0.007686f
C391 B.n351 VSUBS 0.007686f
C392 B.n352 VSUBS 0.007686f
C393 B.n353 VSUBS 0.007686f
C394 B.n354 VSUBS 0.007686f
C395 B.n355 VSUBS 0.007686f
C396 B.n356 VSUBS 0.007686f
C397 B.n357 VSUBS 0.007686f
C398 B.n358 VSUBS 0.007686f
C399 B.n359 VSUBS 0.007686f
C400 B.n360 VSUBS 0.007686f
C401 B.n361 VSUBS 0.007686f
C402 B.n362 VSUBS 0.007686f
C403 B.n363 VSUBS 0.007686f
C404 B.n364 VSUBS 0.007686f
C405 B.n365 VSUBS 0.007686f
C406 B.n366 VSUBS 0.007686f
C407 B.n367 VSUBS 0.007686f
C408 B.n368 VSUBS 0.007686f
C409 B.n369 VSUBS 0.007686f
C410 B.n370 VSUBS 0.007686f
C411 B.n371 VSUBS 0.007686f
C412 B.n372 VSUBS 0.007686f
C413 B.n373 VSUBS 0.007686f
C414 B.n374 VSUBS 0.007686f
C415 B.n375 VSUBS 0.007686f
C416 B.n376 VSUBS 0.007686f
C417 B.n377 VSUBS 0.007686f
C418 B.n378 VSUBS 0.007686f
C419 B.n379 VSUBS 0.007686f
C420 B.n380 VSUBS 0.007686f
C421 B.n381 VSUBS 0.007686f
C422 B.n382 VSUBS 0.007686f
C423 B.n383 VSUBS 0.007686f
C424 B.n384 VSUBS 0.007686f
C425 B.n385 VSUBS 0.007686f
C426 B.n386 VSUBS 0.007686f
C427 B.n387 VSUBS 0.007686f
C428 B.n388 VSUBS 0.007686f
C429 B.n389 VSUBS 0.007686f
C430 B.n390 VSUBS 0.007686f
C431 B.n391 VSUBS 0.007686f
C432 B.n392 VSUBS 0.007686f
C433 B.n393 VSUBS 0.007686f
C434 B.n394 VSUBS 0.007686f
C435 B.n395 VSUBS 0.007686f
C436 B.n396 VSUBS 0.007686f
C437 B.n397 VSUBS 0.007686f
C438 B.n398 VSUBS 0.007686f
C439 B.n399 VSUBS 0.007686f
C440 B.n400 VSUBS 0.007686f
C441 B.n401 VSUBS 0.007686f
C442 B.n402 VSUBS 0.007686f
C443 B.n403 VSUBS 0.007686f
C444 B.n404 VSUBS 0.007686f
C445 B.n405 VSUBS 0.007686f
C446 B.n406 VSUBS 0.007686f
C447 B.n407 VSUBS 0.018085f
C448 B.n408 VSUBS 0.016955f
C449 B.n409 VSUBS 0.016955f
C450 B.n410 VSUBS 0.007686f
C451 B.n411 VSUBS 0.007686f
C452 B.n412 VSUBS 0.007686f
C453 B.n413 VSUBS 0.007686f
C454 B.n414 VSUBS 0.007686f
C455 B.n415 VSUBS 0.007686f
C456 B.n416 VSUBS 0.007686f
C457 B.n417 VSUBS 0.007686f
C458 B.n418 VSUBS 0.007686f
C459 B.n419 VSUBS 0.007686f
C460 B.n420 VSUBS 0.007686f
C461 B.n421 VSUBS 0.007686f
C462 B.n422 VSUBS 0.007686f
C463 B.n423 VSUBS 0.007686f
C464 B.n424 VSUBS 0.007686f
C465 B.n425 VSUBS 0.007686f
C466 B.n426 VSUBS 0.007686f
C467 B.n427 VSUBS 0.007686f
C468 B.n428 VSUBS 0.007686f
C469 B.n429 VSUBS 0.007686f
C470 B.n430 VSUBS 0.007686f
C471 B.n431 VSUBS 0.007686f
C472 B.n432 VSUBS 0.007686f
C473 B.n433 VSUBS 0.007686f
C474 B.n434 VSUBS 0.007686f
C475 B.n435 VSUBS 0.007686f
C476 B.n436 VSUBS 0.007686f
C477 B.n437 VSUBS 0.007686f
C478 B.n438 VSUBS 0.007686f
C479 B.n439 VSUBS 0.007686f
C480 B.n440 VSUBS 0.007686f
C481 B.n441 VSUBS 0.007686f
C482 B.n442 VSUBS 0.007686f
C483 B.n443 VSUBS 0.007686f
C484 B.n444 VSUBS 0.007686f
C485 B.n445 VSUBS 0.007686f
C486 B.n446 VSUBS 0.007686f
C487 B.n447 VSUBS 0.007686f
C488 B.n448 VSUBS 0.007686f
C489 B.n449 VSUBS 0.007686f
C490 B.n450 VSUBS 0.007686f
C491 B.n451 VSUBS 0.007686f
C492 B.n452 VSUBS 0.007686f
C493 B.n453 VSUBS 0.007686f
C494 B.n454 VSUBS 0.007686f
C495 B.n455 VSUBS 0.007686f
C496 B.n456 VSUBS 0.007686f
C497 B.n457 VSUBS 0.007686f
C498 B.n458 VSUBS 0.007686f
C499 B.n459 VSUBS 0.0179f
C500 B.n460 VSUBS 0.016955f
C501 B.n461 VSUBS 0.018085f
C502 B.n462 VSUBS 0.007686f
C503 B.n463 VSUBS 0.007686f
C504 B.n464 VSUBS 0.007686f
C505 B.n465 VSUBS 0.007686f
C506 B.n466 VSUBS 0.007686f
C507 B.n467 VSUBS 0.007686f
C508 B.n468 VSUBS 0.007686f
C509 B.n469 VSUBS 0.007686f
C510 B.n470 VSUBS 0.007686f
C511 B.n471 VSUBS 0.007686f
C512 B.n472 VSUBS 0.007686f
C513 B.n473 VSUBS 0.007686f
C514 B.n474 VSUBS 0.007686f
C515 B.n475 VSUBS 0.007686f
C516 B.n476 VSUBS 0.007686f
C517 B.n477 VSUBS 0.007686f
C518 B.n478 VSUBS 0.007686f
C519 B.n479 VSUBS 0.007686f
C520 B.n480 VSUBS 0.007686f
C521 B.n481 VSUBS 0.007686f
C522 B.n482 VSUBS 0.007686f
C523 B.n483 VSUBS 0.007686f
C524 B.n484 VSUBS 0.007686f
C525 B.n485 VSUBS 0.007686f
C526 B.n486 VSUBS 0.007686f
C527 B.n487 VSUBS 0.007686f
C528 B.n488 VSUBS 0.007686f
C529 B.n489 VSUBS 0.007686f
C530 B.n490 VSUBS 0.007686f
C531 B.n491 VSUBS 0.007686f
C532 B.n492 VSUBS 0.007686f
C533 B.n493 VSUBS 0.007686f
C534 B.n494 VSUBS 0.007686f
C535 B.n495 VSUBS 0.007686f
C536 B.n496 VSUBS 0.007686f
C537 B.n497 VSUBS 0.007686f
C538 B.n498 VSUBS 0.007686f
C539 B.n499 VSUBS 0.007686f
C540 B.n500 VSUBS 0.007686f
C541 B.n501 VSUBS 0.007686f
C542 B.n502 VSUBS 0.007686f
C543 B.n503 VSUBS 0.007686f
C544 B.n504 VSUBS 0.007686f
C545 B.n505 VSUBS 0.007686f
C546 B.n506 VSUBS 0.007686f
C547 B.n507 VSUBS 0.007686f
C548 B.n508 VSUBS 0.007686f
C549 B.n509 VSUBS 0.007686f
C550 B.n510 VSUBS 0.007686f
C551 B.n511 VSUBS 0.007686f
C552 B.n512 VSUBS 0.007686f
C553 B.n513 VSUBS 0.007686f
C554 B.n514 VSUBS 0.007686f
C555 B.n515 VSUBS 0.007686f
C556 B.n516 VSUBS 0.007686f
C557 B.n517 VSUBS 0.007686f
C558 B.n518 VSUBS 0.007686f
C559 B.n519 VSUBS 0.007686f
C560 B.n520 VSUBS 0.007686f
C561 B.n521 VSUBS 0.007686f
C562 B.n522 VSUBS 0.007686f
C563 B.n523 VSUBS 0.007686f
C564 B.n524 VSUBS 0.007686f
C565 B.n525 VSUBS 0.007686f
C566 B.n526 VSUBS 0.007686f
C567 B.n527 VSUBS 0.007686f
C568 B.n528 VSUBS 0.007686f
C569 B.n529 VSUBS 0.007686f
C570 B.n530 VSUBS 0.007686f
C571 B.n531 VSUBS 0.007686f
C572 B.n532 VSUBS 0.007686f
C573 B.n533 VSUBS 0.007686f
C574 B.n534 VSUBS 0.007686f
C575 B.n535 VSUBS 0.007686f
C576 B.n536 VSUBS 0.007686f
C577 B.n537 VSUBS 0.007686f
C578 B.n538 VSUBS 0.007686f
C579 B.n539 VSUBS 0.007686f
C580 B.n540 VSUBS 0.007686f
C581 B.n541 VSUBS 0.007686f
C582 B.n542 VSUBS 0.007686f
C583 B.n543 VSUBS 0.007686f
C584 B.n544 VSUBS 0.007686f
C585 B.n545 VSUBS 0.007686f
C586 B.n546 VSUBS 0.007686f
C587 B.n547 VSUBS 0.007686f
C588 B.n548 VSUBS 0.007686f
C589 B.n549 VSUBS 0.007686f
C590 B.n550 VSUBS 0.007686f
C591 B.n551 VSUBS 0.007686f
C592 B.n552 VSUBS 0.007686f
C593 B.n553 VSUBS 0.007686f
C594 B.n554 VSUBS 0.005313f
C595 B.n555 VSUBS 0.017808f
C596 B.n556 VSUBS 0.006217f
C597 B.n557 VSUBS 0.007686f
C598 B.n558 VSUBS 0.007686f
C599 B.n559 VSUBS 0.007686f
C600 B.n560 VSUBS 0.007686f
C601 B.n561 VSUBS 0.007686f
C602 B.n562 VSUBS 0.007686f
C603 B.n563 VSUBS 0.007686f
C604 B.n564 VSUBS 0.007686f
C605 B.n565 VSUBS 0.007686f
C606 B.n566 VSUBS 0.007686f
C607 B.n567 VSUBS 0.007686f
C608 B.n568 VSUBS 0.006217f
C609 B.n569 VSUBS 0.007686f
C610 B.n570 VSUBS 0.007686f
C611 B.n571 VSUBS 0.005313f
C612 B.n572 VSUBS 0.007686f
C613 B.n573 VSUBS 0.007686f
C614 B.n574 VSUBS 0.007686f
C615 B.n575 VSUBS 0.007686f
C616 B.n576 VSUBS 0.007686f
C617 B.n577 VSUBS 0.007686f
C618 B.n578 VSUBS 0.007686f
C619 B.n579 VSUBS 0.007686f
C620 B.n580 VSUBS 0.007686f
C621 B.n581 VSUBS 0.007686f
C622 B.n582 VSUBS 0.007686f
C623 B.n583 VSUBS 0.007686f
C624 B.n584 VSUBS 0.007686f
C625 B.n585 VSUBS 0.007686f
C626 B.n586 VSUBS 0.007686f
C627 B.n587 VSUBS 0.007686f
C628 B.n588 VSUBS 0.007686f
C629 B.n589 VSUBS 0.007686f
C630 B.n590 VSUBS 0.007686f
C631 B.n591 VSUBS 0.007686f
C632 B.n592 VSUBS 0.007686f
C633 B.n593 VSUBS 0.007686f
C634 B.n594 VSUBS 0.007686f
C635 B.n595 VSUBS 0.007686f
C636 B.n596 VSUBS 0.007686f
C637 B.n597 VSUBS 0.007686f
C638 B.n598 VSUBS 0.007686f
C639 B.n599 VSUBS 0.007686f
C640 B.n600 VSUBS 0.007686f
C641 B.n601 VSUBS 0.007686f
C642 B.n602 VSUBS 0.007686f
C643 B.n603 VSUBS 0.007686f
C644 B.n604 VSUBS 0.007686f
C645 B.n605 VSUBS 0.007686f
C646 B.n606 VSUBS 0.007686f
C647 B.n607 VSUBS 0.007686f
C648 B.n608 VSUBS 0.007686f
C649 B.n609 VSUBS 0.007686f
C650 B.n610 VSUBS 0.007686f
C651 B.n611 VSUBS 0.007686f
C652 B.n612 VSUBS 0.007686f
C653 B.n613 VSUBS 0.007686f
C654 B.n614 VSUBS 0.007686f
C655 B.n615 VSUBS 0.007686f
C656 B.n616 VSUBS 0.007686f
C657 B.n617 VSUBS 0.007686f
C658 B.n618 VSUBS 0.007686f
C659 B.n619 VSUBS 0.007686f
C660 B.n620 VSUBS 0.007686f
C661 B.n621 VSUBS 0.007686f
C662 B.n622 VSUBS 0.007686f
C663 B.n623 VSUBS 0.007686f
C664 B.n624 VSUBS 0.007686f
C665 B.n625 VSUBS 0.007686f
C666 B.n626 VSUBS 0.007686f
C667 B.n627 VSUBS 0.007686f
C668 B.n628 VSUBS 0.007686f
C669 B.n629 VSUBS 0.007686f
C670 B.n630 VSUBS 0.007686f
C671 B.n631 VSUBS 0.007686f
C672 B.n632 VSUBS 0.007686f
C673 B.n633 VSUBS 0.007686f
C674 B.n634 VSUBS 0.007686f
C675 B.n635 VSUBS 0.007686f
C676 B.n636 VSUBS 0.007686f
C677 B.n637 VSUBS 0.007686f
C678 B.n638 VSUBS 0.007686f
C679 B.n639 VSUBS 0.007686f
C680 B.n640 VSUBS 0.007686f
C681 B.n641 VSUBS 0.007686f
C682 B.n642 VSUBS 0.007686f
C683 B.n643 VSUBS 0.007686f
C684 B.n644 VSUBS 0.007686f
C685 B.n645 VSUBS 0.007686f
C686 B.n646 VSUBS 0.007686f
C687 B.n647 VSUBS 0.007686f
C688 B.n648 VSUBS 0.007686f
C689 B.n649 VSUBS 0.007686f
C690 B.n650 VSUBS 0.007686f
C691 B.n651 VSUBS 0.007686f
C692 B.n652 VSUBS 0.007686f
C693 B.n653 VSUBS 0.007686f
C694 B.n654 VSUBS 0.007686f
C695 B.n655 VSUBS 0.007686f
C696 B.n656 VSUBS 0.007686f
C697 B.n657 VSUBS 0.007686f
C698 B.n658 VSUBS 0.007686f
C699 B.n659 VSUBS 0.007686f
C700 B.n660 VSUBS 0.007686f
C701 B.n661 VSUBS 0.007686f
C702 B.n662 VSUBS 0.007686f
C703 B.n663 VSUBS 0.018085f
C704 B.n664 VSUBS 0.018085f
C705 B.n665 VSUBS 0.016955f
C706 B.n666 VSUBS 0.007686f
C707 B.n667 VSUBS 0.007686f
C708 B.n668 VSUBS 0.007686f
C709 B.n669 VSUBS 0.007686f
C710 B.n670 VSUBS 0.007686f
C711 B.n671 VSUBS 0.007686f
C712 B.n672 VSUBS 0.007686f
C713 B.n673 VSUBS 0.007686f
C714 B.n674 VSUBS 0.007686f
C715 B.n675 VSUBS 0.007686f
C716 B.n676 VSUBS 0.007686f
C717 B.n677 VSUBS 0.007686f
C718 B.n678 VSUBS 0.007686f
C719 B.n679 VSUBS 0.007686f
C720 B.n680 VSUBS 0.007686f
C721 B.n681 VSUBS 0.007686f
C722 B.n682 VSUBS 0.007686f
C723 B.n683 VSUBS 0.007686f
C724 B.n684 VSUBS 0.007686f
C725 B.n685 VSUBS 0.007686f
C726 B.n686 VSUBS 0.007686f
C727 B.n687 VSUBS 0.007686f
C728 B.n688 VSUBS 0.007686f
C729 B.n689 VSUBS 0.007686f
C730 B.n690 VSUBS 0.007686f
C731 B.n691 VSUBS 0.017404f
C732 VDD2.t1 VSUBS 0.430511f
C733 VDD2.t0 VSUBS 0.430511f
C734 VDD2.n0 VSUBS 4.54891f
C735 VDD2.t3 VSUBS 0.430511f
C736 VDD2.t2 VSUBS 0.430511f
C737 VDD2.n1 VSUBS 3.62751f
C738 VDD2.n2 VSUBS 4.91552f
C739 VN.t2 VSUBS 2.1436f
C740 VN.t3 VSUBS 2.14354f
C741 VN.n0 VSUBS 1.55094f
C742 VN.t1 VSUBS 2.1436f
C743 VN.t0 VSUBS 2.14354f
C744 VN.n1 VSUBS 3.01719f
C745 VDD1.t1 VSUBS 0.430362f
C746 VDD1.t3 VSUBS 0.430362f
C747 VDD1.n0 VSUBS 3.62677f
C748 VDD1.t2 VSUBS 0.430362f
C749 VDD1.t0 VSUBS 0.430362f
C750 VDD1.n1 VSUBS 4.57585f
C751 VTAIL.t0 VSUBS 3.52647f
C752 VTAIL.n0 VSUBS 0.689353f
C753 VTAIL.t6 VSUBS 3.52647f
C754 VTAIL.n1 VSUBS 0.71641f
C755 VTAIL.t7 VSUBS 3.52647f
C756 VTAIL.n2 VSUBS 2.23065f
C757 VTAIL.t2 VSUBS 3.5265f
C758 VTAIL.n3 VSUBS 2.23062f
C759 VTAIL.t1 VSUBS 3.5265f
C760 VTAIL.n4 VSUBS 0.716378f
C761 VTAIL.t4 VSUBS 3.5265f
C762 VTAIL.n5 VSUBS 0.716378f
C763 VTAIL.t5 VSUBS 3.52647f
C764 VTAIL.n6 VSUBS 2.23065f
C765 VTAIL.t3 VSUBS 3.52647f
C766 VTAIL.n7 VSUBS 2.19525f
C767 VP.n0 VSUBS 0.058812f
C768 VP.t0 VSUBS 2.19041f
C769 VP.t2 VSUBS 2.19047f
C770 VP.n1 VSUBS 3.05762f
C771 VP.n2 VSUBS 4.27182f
C772 VP.t1 VSUBS 2.16794f
C773 VP.n3 VSUBS 0.807966f
C774 VP.n4 VSUBS 0.013346f
C775 VP.t3 VSUBS 2.16794f
C776 VP.n5 VSUBS 0.807966f
C777 VP.n6 VSUBS 0.045577f
.ends

