* NGSPICE file created from diff_pair_sample_0146.ext - technology: sky130A

.subckt diff_pair_sample_0146 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6596 pd=40.06 as=0 ps=0 w=19.64 l=1.36
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=7.6596 pd=40.06 as=0 ps=0 w=19.64 l=1.36
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6596 pd=40.06 as=0 ps=0 w=19.64 l=1.36
X3 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=7.6596 pd=40.06 as=7.6596 ps=40.06 w=19.64 l=1.36
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.6596 pd=40.06 as=7.6596 ps=40.06 w=19.64 l=1.36
X5 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.6596 pd=40.06 as=7.6596 ps=40.06 w=19.64 l=1.36
X6 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.6596 pd=40.06 as=7.6596 ps=40.06 w=19.64 l=1.36
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.6596 pd=40.06 as=0 ps=0 w=19.64 l=1.36
R0 B.n573 B.n572 585
R1 B.n575 B.n110 585
R2 B.n578 B.n577 585
R3 B.n579 B.n109 585
R4 B.n581 B.n580 585
R5 B.n583 B.n108 585
R6 B.n586 B.n585 585
R7 B.n587 B.n107 585
R8 B.n589 B.n588 585
R9 B.n591 B.n106 585
R10 B.n594 B.n593 585
R11 B.n595 B.n105 585
R12 B.n597 B.n596 585
R13 B.n599 B.n104 585
R14 B.n602 B.n601 585
R15 B.n603 B.n103 585
R16 B.n605 B.n604 585
R17 B.n607 B.n102 585
R18 B.n610 B.n609 585
R19 B.n611 B.n101 585
R20 B.n613 B.n612 585
R21 B.n615 B.n100 585
R22 B.n618 B.n617 585
R23 B.n619 B.n99 585
R24 B.n621 B.n620 585
R25 B.n623 B.n98 585
R26 B.n626 B.n625 585
R27 B.n627 B.n97 585
R28 B.n629 B.n628 585
R29 B.n631 B.n96 585
R30 B.n634 B.n633 585
R31 B.n635 B.n95 585
R32 B.n637 B.n636 585
R33 B.n639 B.n94 585
R34 B.n642 B.n641 585
R35 B.n643 B.n93 585
R36 B.n645 B.n644 585
R37 B.n647 B.n92 585
R38 B.n650 B.n649 585
R39 B.n651 B.n91 585
R40 B.n653 B.n652 585
R41 B.n655 B.n90 585
R42 B.n658 B.n657 585
R43 B.n659 B.n89 585
R44 B.n661 B.n660 585
R45 B.n663 B.n88 585
R46 B.n666 B.n665 585
R47 B.n667 B.n87 585
R48 B.n669 B.n668 585
R49 B.n671 B.n86 585
R50 B.n674 B.n673 585
R51 B.n675 B.n85 585
R52 B.n677 B.n676 585
R53 B.n679 B.n84 585
R54 B.n682 B.n681 585
R55 B.n683 B.n83 585
R56 B.n685 B.n684 585
R57 B.n687 B.n82 585
R58 B.n690 B.n689 585
R59 B.n691 B.n81 585
R60 B.n693 B.n692 585
R61 B.n695 B.n80 585
R62 B.n697 B.n696 585
R63 B.n699 B.n698 585
R64 B.n702 B.n701 585
R65 B.n703 B.n75 585
R66 B.n705 B.n704 585
R67 B.n707 B.n74 585
R68 B.n710 B.n709 585
R69 B.n711 B.n73 585
R70 B.n713 B.n712 585
R71 B.n715 B.n72 585
R72 B.n718 B.n717 585
R73 B.n719 B.n69 585
R74 B.n722 B.n721 585
R75 B.n724 B.n68 585
R76 B.n727 B.n726 585
R77 B.n728 B.n67 585
R78 B.n730 B.n729 585
R79 B.n732 B.n66 585
R80 B.n735 B.n734 585
R81 B.n736 B.n65 585
R82 B.n738 B.n737 585
R83 B.n740 B.n64 585
R84 B.n743 B.n742 585
R85 B.n744 B.n63 585
R86 B.n746 B.n745 585
R87 B.n748 B.n62 585
R88 B.n751 B.n750 585
R89 B.n752 B.n61 585
R90 B.n754 B.n753 585
R91 B.n756 B.n60 585
R92 B.n759 B.n758 585
R93 B.n760 B.n59 585
R94 B.n762 B.n761 585
R95 B.n764 B.n58 585
R96 B.n767 B.n766 585
R97 B.n768 B.n57 585
R98 B.n770 B.n769 585
R99 B.n772 B.n56 585
R100 B.n775 B.n774 585
R101 B.n776 B.n55 585
R102 B.n778 B.n777 585
R103 B.n780 B.n54 585
R104 B.n783 B.n782 585
R105 B.n784 B.n53 585
R106 B.n786 B.n785 585
R107 B.n788 B.n52 585
R108 B.n791 B.n790 585
R109 B.n792 B.n51 585
R110 B.n794 B.n793 585
R111 B.n796 B.n50 585
R112 B.n799 B.n798 585
R113 B.n800 B.n49 585
R114 B.n802 B.n801 585
R115 B.n804 B.n48 585
R116 B.n807 B.n806 585
R117 B.n808 B.n47 585
R118 B.n810 B.n809 585
R119 B.n812 B.n46 585
R120 B.n815 B.n814 585
R121 B.n816 B.n45 585
R122 B.n818 B.n817 585
R123 B.n820 B.n44 585
R124 B.n823 B.n822 585
R125 B.n824 B.n43 585
R126 B.n826 B.n825 585
R127 B.n828 B.n42 585
R128 B.n831 B.n830 585
R129 B.n832 B.n41 585
R130 B.n834 B.n833 585
R131 B.n836 B.n40 585
R132 B.n839 B.n838 585
R133 B.n840 B.n39 585
R134 B.n842 B.n841 585
R135 B.n844 B.n38 585
R136 B.n847 B.n846 585
R137 B.n848 B.n37 585
R138 B.n571 B.n35 585
R139 B.n851 B.n35 585
R140 B.n570 B.n34 585
R141 B.n852 B.n34 585
R142 B.n569 B.n33 585
R143 B.n853 B.n33 585
R144 B.n568 B.n567 585
R145 B.n567 B.n29 585
R146 B.n566 B.n28 585
R147 B.n859 B.n28 585
R148 B.n565 B.n27 585
R149 B.n860 B.n27 585
R150 B.n564 B.n26 585
R151 B.n861 B.n26 585
R152 B.n563 B.n562 585
R153 B.n562 B.n22 585
R154 B.n561 B.n21 585
R155 B.n867 B.n21 585
R156 B.n560 B.n20 585
R157 B.n868 B.n20 585
R158 B.n559 B.n19 585
R159 B.n869 B.n19 585
R160 B.n558 B.n557 585
R161 B.n557 B.n15 585
R162 B.n556 B.n14 585
R163 B.n875 B.n14 585
R164 B.n555 B.n13 585
R165 B.n876 B.n13 585
R166 B.n554 B.n12 585
R167 B.n877 B.n12 585
R168 B.n553 B.n552 585
R169 B.n552 B.n8 585
R170 B.n551 B.n7 585
R171 B.n883 B.n7 585
R172 B.n550 B.n6 585
R173 B.n884 B.n6 585
R174 B.n549 B.n5 585
R175 B.n885 B.n5 585
R176 B.n548 B.n547 585
R177 B.n547 B.n4 585
R178 B.n546 B.n111 585
R179 B.n546 B.n545 585
R180 B.n536 B.n112 585
R181 B.n113 B.n112 585
R182 B.n538 B.n537 585
R183 B.n539 B.n538 585
R184 B.n535 B.n117 585
R185 B.n121 B.n117 585
R186 B.n534 B.n533 585
R187 B.n533 B.n532 585
R188 B.n119 B.n118 585
R189 B.n120 B.n119 585
R190 B.n525 B.n524 585
R191 B.n526 B.n525 585
R192 B.n523 B.n126 585
R193 B.n126 B.n125 585
R194 B.n522 B.n521 585
R195 B.n521 B.n520 585
R196 B.n128 B.n127 585
R197 B.n129 B.n128 585
R198 B.n513 B.n512 585
R199 B.n514 B.n513 585
R200 B.n511 B.n133 585
R201 B.n137 B.n133 585
R202 B.n510 B.n509 585
R203 B.n509 B.n508 585
R204 B.n135 B.n134 585
R205 B.n136 B.n135 585
R206 B.n501 B.n500 585
R207 B.n502 B.n501 585
R208 B.n499 B.n142 585
R209 B.n142 B.n141 585
R210 B.n498 B.n497 585
R211 B.n497 B.n496 585
R212 B.n493 B.n146 585
R213 B.n492 B.n491 585
R214 B.n489 B.n147 585
R215 B.n489 B.n145 585
R216 B.n488 B.n487 585
R217 B.n486 B.n485 585
R218 B.n484 B.n149 585
R219 B.n482 B.n481 585
R220 B.n480 B.n150 585
R221 B.n479 B.n478 585
R222 B.n476 B.n151 585
R223 B.n474 B.n473 585
R224 B.n472 B.n152 585
R225 B.n471 B.n470 585
R226 B.n468 B.n153 585
R227 B.n466 B.n465 585
R228 B.n464 B.n154 585
R229 B.n463 B.n462 585
R230 B.n460 B.n155 585
R231 B.n458 B.n457 585
R232 B.n456 B.n156 585
R233 B.n455 B.n454 585
R234 B.n452 B.n157 585
R235 B.n450 B.n449 585
R236 B.n448 B.n158 585
R237 B.n447 B.n446 585
R238 B.n444 B.n159 585
R239 B.n442 B.n441 585
R240 B.n440 B.n160 585
R241 B.n439 B.n438 585
R242 B.n436 B.n161 585
R243 B.n434 B.n433 585
R244 B.n432 B.n162 585
R245 B.n431 B.n430 585
R246 B.n428 B.n163 585
R247 B.n426 B.n425 585
R248 B.n424 B.n164 585
R249 B.n423 B.n422 585
R250 B.n420 B.n165 585
R251 B.n418 B.n417 585
R252 B.n416 B.n166 585
R253 B.n415 B.n414 585
R254 B.n412 B.n167 585
R255 B.n410 B.n409 585
R256 B.n408 B.n168 585
R257 B.n407 B.n406 585
R258 B.n404 B.n169 585
R259 B.n402 B.n401 585
R260 B.n400 B.n170 585
R261 B.n399 B.n398 585
R262 B.n396 B.n171 585
R263 B.n394 B.n393 585
R264 B.n392 B.n172 585
R265 B.n391 B.n390 585
R266 B.n388 B.n173 585
R267 B.n386 B.n385 585
R268 B.n384 B.n174 585
R269 B.n383 B.n382 585
R270 B.n380 B.n175 585
R271 B.n378 B.n377 585
R272 B.n376 B.n176 585
R273 B.n375 B.n374 585
R274 B.n372 B.n177 585
R275 B.n370 B.n369 585
R276 B.n368 B.n178 585
R277 B.n366 B.n365 585
R278 B.n363 B.n181 585
R279 B.n361 B.n360 585
R280 B.n359 B.n182 585
R281 B.n358 B.n357 585
R282 B.n355 B.n183 585
R283 B.n353 B.n352 585
R284 B.n351 B.n184 585
R285 B.n350 B.n349 585
R286 B.n347 B.n185 585
R287 B.n345 B.n344 585
R288 B.n343 B.n186 585
R289 B.n342 B.n341 585
R290 B.n339 B.n190 585
R291 B.n337 B.n336 585
R292 B.n335 B.n191 585
R293 B.n334 B.n333 585
R294 B.n331 B.n192 585
R295 B.n329 B.n328 585
R296 B.n327 B.n193 585
R297 B.n326 B.n325 585
R298 B.n323 B.n194 585
R299 B.n321 B.n320 585
R300 B.n319 B.n195 585
R301 B.n318 B.n317 585
R302 B.n315 B.n196 585
R303 B.n313 B.n312 585
R304 B.n311 B.n197 585
R305 B.n310 B.n309 585
R306 B.n307 B.n198 585
R307 B.n305 B.n304 585
R308 B.n303 B.n199 585
R309 B.n302 B.n301 585
R310 B.n299 B.n200 585
R311 B.n297 B.n296 585
R312 B.n295 B.n201 585
R313 B.n294 B.n293 585
R314 B.n291 B.n202 585
R315 B.n289 B.n288 585
R316 B.n287 B.n203 585
R317 B.n286 B.n285 585
R318 B.n283 B.n204 585
R319 B.n281 B.n280 585
R320 B.n279 B.n205 585
R321 B.n278 B.n277 585
R322 B.n275 B.n206 585
R323 B.n273 B.n272 585
R324 B.n271 B.n207 585
R325 B.n270 B.n269 585
R326 B.n267 B.n208 585
R327 B.n265 B.n264 585
R328 B.n263 B.n209 585
R329 B.n262 B.n261 585
R330 B.n259 B.n210 585
R331 B.n257 B.n256 585
R332 B.n255 B.n211 585
R333 B.n254 B.n253 585
R334 B.n251 B.n212 585
R335 B.n249 B.n248 585
R336 B.n247 B.n213 585
R337 B.n246 B.n245 585
R338 B.n243 B.n214 585
R339 B.n241 B.n240 585
R340 B.n239 B.n215 585
R341 B.n238 B.n237 585
R342 B.n235 B.n216 585
R343 B.n233 B.n232 585
R344 B.n231 B.n217 585
R345 B.n230 B.n229 585
R346 B.n227 B.n218 585
R347 B.n225 B.n224 585
R348 B.n223 B.n219 585
R349 B.n222 B.n221 585
R350 B.n144 B.n143 585
R351 B.n145 B.n144 585
R352 B.n495 B.n494 585
R353 B.n496 B.n495 585
R354 B.n140 B.n139 585
R355 B.n141 B.n140 585
R356 B.n504 B.n503 585
R357 B.n503 B.n502 585
R358 B.n505 B.n138 585
R359 B.n138 B.n136 585
R360 B.n507 B.n506 585
R361 B.n508 B.n507 585
R362 B.n132 B.n131 585
R363 B.n137 B.n132 585
R364 B.n516 B.n515 585
R365 B.n515 B.n514 585
R366 B.n517 B.n130 585
R367 B.n130 B.n129 585
R368 B.n519 B.n518 585
R369 B.n520 B.n519 585
R370 B.n124 B.n123 585
R371 B.n125 B.n124 585
R372 B.n528 B.n527 585
R373 B.n527 B.n526 585
R374 B.n529 B.n122 585
R375 B.n122 B.n120 585
R376 B.n531 B.n530 585
R377 B.n532 B.n531 585
R378 B.n116 B.n115 585
R379 B.n121 B.n116 585
R380 B.n541 B.n540 585
R381 B.n540 B.n539 585
R382 B.n542 B.n114 585
R383 B.n114 B.n113 585
R384 B.n544 B.n543 585
R385 B.n545 B.n544 585
R386 B.n2 B.n0 585
R387 B.n4 B.n2 585
R388 B.n3 B.n1 585
R389 B.n884 B.n3 585
R390 B.n882 B.n881 585
R391 B.n883 B.n882 585
R392 B.n880 B.n9 585
R393 B.n9 B.n8 585
R394 B.n879 B.n878 585
R395 B.n878 B.n877 585
R396 B.n11 B.n10 585
R397 B.n876 B.n11 585
R398 B.n874 B.n873 585
R399 B.n875 B.n874 585
R400 B.n872 B.n16 585
R401 B.n16 B.n15 585
R402 B.n871 B.n870 585
R403 B.n870 B.n869 585
R404 B.n18 B.n17 585
R405 B.n868 B.n18 585
R406 B.n866 B.n865 585
R407 B.n867 B.n866 585
R408 B.n864 B.n23 585
R409 B.n23 B.n22 585
R410 B.n863 B.n862 585
R411 B.n862 B.n861 585
R412 B.n25 B.n24 585
R413 B.n860 B.n25 585
R414 B.n858 B.n857 585
R415 B.n859 B.n858 585
R416 B.n856 B.n30 585
R417 B.n30 B.n29 585
R418 B.n855 B.n854 585
R419 B.n854 B.n853 585
R420 B.n32 B.n31 585
R421 B.n852 B.n32 585
R422 B.n850 B.n849 585
R423 B.n851 B.n850 585
R424 B.n887 B.n886 585
R425 B.n886 B.n885 585
R426 B.n187 B.t10 552.909
R427 B.n179 B.t2 552.909
R428 B.n70 B.t13 552.909
R429 B.n76 B.t6 552.909
R430 B.n495 B.n146 487.695
R431 B.n850 B.n37 487.695
R432 B.n497 B.n144 487.695
R433 B.n573 B.n35 487.695
R434 B.n187 B.t12 446.724
R435 B.n179 B.t5 446.724
R436 B.n70 B.t14 446.724
R437 B.n76 B.t8 446.724
R438 B.n188 B.t11 413.947
R439 B.n77 B.t9 413.947
R440 B.n180 B.t4 413.947
R441 B.n71 B.t15 413.947
R442 B.n574 B.n36 256.663
R443 B.n576 B.n36 256.663
R444 B.n582 B.n36 256.663
R445 B.n584 B.n36 256.663
R446 B.n590 B.n36 256.663
R447 B.n592 B.n36 256.663
R448 B.n598 B.n36 256.663
R449 B.n600 B.n36 256.663
R450 B.n606 B.n36 256.663
R451 B.n608 B.n36 256.663
R452 B.n614 B.n36 256.663
R453 B.n616 B.n36 256.663
R454 B.n622 B.n36 256.663
R455 B.n624 B.n36 256.663
R456 B.n630 B.n36 256.663
R457 B.n632 B.n36 256.663
R458 B.n638 B.n36 256.663
R459 B.n640 B.n36 256.663
R460 B.n646 B.n36 256.663
R461 B.n648 B.n36 256.663
R462 B.n654 B.n36 256.663
R463 B.n656 B.n36 256.663
R464 B.n662 B.n36 256.663
R465 B.n664 B.n36 256.663
R466 B.n670 B.n36 256.663
R467 B.n672 B.n36 256.663
R468 B.n678 B.n36 256.663
R469 B.n680 B.n36 256.663
R470 B.n686 B.n36 256.663
R471 B.n688 B.n36 256.663
R472 B.n694 B.n36 256.663
R473 B.n79 B.n36 256.663
R474 B.n700 B.n36 256.663
R475 B.n706 B.n36 256.663
R476 B.n708 B.n36 256.663
R477 B.n714 B.n36 256.663
R478 B.n716 B.n36 256.663
R479 B.n723 B.n36 256.663
R480 B.n725 B.n36 256.663
R481 B.n731 B.n36 256.663
R482 B.n733 B.n36 256.663
R483 B.n739 B.n36 256.663
R484 B.n741 B.n36 256.663
R485 B.n747 B.n36 256.663
R486 B.n749 B.n36 256.663
R487 B.n755 B.n36 256.663
R488 B.n757 B.n36 256.663
R489 B.n763 B.n36 256.663
R490 B.n765 B.n36 256.663
R491 B.n771 B.n36 256.663
R492 B.n773 B.n36 256.663
R493 B.n779 B.n36 256.663
R494 B.n781 B.n36 256.663
R495 B.n787 B.n36 256.663
R496 B.n789 B.n36 256.663
R497 B.n795 B.n36 256.663
R498 B.n797 B.n36 256.663
R499 B.n803 B.n36 256.663
R500 B.n805 B.n36 256.663
R501 B.n811 B.n36 256.663
R502 B.n813 B.n36 256.663
R503 B.n819 B.n36 256.663
R504 B.n821 B.n36 256.663
R505 B.n827 B.n36 256.663
R506 B.n829 B.n36 256.663
R507 B.n835 B.n36 256.663
R508 B.n837 B.n36 256.663
R509 B.n843 B.n36 256.663
R510 B.n845 B.n36 256.663
R511 B.n490 B.n145 256.663
R512 B.n148 B.n145 256.663
R513 B.n483 B.n145 256.663
R514 B.n477 B.n145 256.663
R515 B.n475 B.n145 256.663
R516 B.n469 B.n145 256.663
R517 B.n467 B.n145 256.663
R518 B.n461 B.n145 256.663
R519 B.n459 B.n145 256.663
R520 B.n453 B.n145 256.663
R521 B.n451 B.n145 256.663
R522 B.n445 B.n145 256.663
R523 B.n443 B.n145 256.663
R524 B.n437 B.n145 256.663
R525 B.n435 B.n145 256.663
R526 B.n429 B.n145 256.663
R527 B.n427 B.n145 256.663
R528 B.n421 B.n145 256.663
R529 B.n419 B.n145 256.663
R530 B.n413 B.n145 256.663
R531 B.n411 B.n145 256.663
R532 B.n405 B.n145 256.663
R533 B.n403 B.n145 256.663
R534 B.n397 B.n145 256.663
R535 B.n395 B.n145 256.663
R536 B.n389 B.n145 256.663
R537 B.n387 B.n145 256.663
R538 B.n381 B.n145 256.663
R539 B.n379 B.n145 256.663
R540 B.n373 B.n145 256.663
R541 B.n371 B.n145 256.663
R542 B.n364 B.n145 256.663
R543 B.n362 B.n145 256.663
R544 B.n356 B.n145 256.663
R545 B.n354 B.n145 256.663
R546 B.n348 B.n145 256.663
R547 B.n346 B.n145 256.663
R548 B.n340 B.n145 256.663
R549 B.n338 B.n145 256.663
R550 B.n332 B.n145 256.663
R551 B.n330 B.n145 256.663
R552 B.n324 B.n145 256.663
R553 B.n322 B.n145 256.663
R554 B.n316 B.n145 256.663
R555 B.n314 B.n145 256.663
R556 B.n308 B.n145 256.663
R557 B.n306 B.n145 256.663
R558 B.n300 B.n145 256.663
R559 B.n298 B.n145 256.663
R560 B.n292 B.n145 256.663
R561 B.n290 B.n145 256.663
R562 B.n284 B.n145 256.663
R563 B.n282 B.n145 256.663
R564 B.n276 B.n145 256.663
R565 B.n274 B.n145 256.663
R566 B.n268 B.n145 256.663
R567 B.n266 B.n145 256.663
R568 B.n260 B.n145 256.663
R569 B.n258 B.n145 256.663
R570 B.n252 B.n145 256.663
R571 B.n250 B.n145 256.663
R572 B.n244 B.n145 256.663
R573 B.n242 B.n145 256.663
R574 B.n236 B.n145 256.663
R575 B.n234 B.n145 256.663
R576 B.n228 B.n145 256.663
R577 B.n226 B.n145 256.663
R578 B.n220 B.n145 256.663
R579 B.n495 B.n140 163.367
R580 B.n503 B.n140 163.367
R581 B.n503 B.n138 163.367
R582 B.n507 B.n138 163.367
R583 B.n507 B.n132 163.367
R584 B.n515 B.n132 163.367
R585 B.n515 B.n130 163.367
R586 B.n519 B.n130 163.367
R587 B.n519 B.n124 163.367
R588 B.n527 B.n124 163.367
R589 B.n527 B.n122 163.367
R590 B.n531 B.n122 163.367
R591 B.n531 B.n116 163.367
R592 B.n540 B.n116 163.367
R593 B.n540 B.n114 163.367
R594 B.n544 B.n114 163.367
R595 B.n544 B.n2 163.367
R596 B.n886 B.n2 163.367
R597 B.n886 B.n3 163.367
R598 B.n882 B.n3 163.367
R599 B.n882 B.n9 163.367
R600 B.n878 B.n9 163.367
R601 B.n878 B.n11 163.367
R602 B.n874 B.n11 163.367
R603 B.n874 B.n16 163.367
R604 B.n870 B.n16 163.367
R605 B.n870 B.n18 163.367
R606 B.n866 B.n18 163.367
R607 B.n866 B.n23 163.367
R608 B.n862 B.n23 163.367
R609 B.n862 B.n25 163.367
R610 B.n858 B.n25 163.367
R611 B.n858 B.n30 163.367
R612 B.n854 B.n30 163.367
R613 B.n854 B.n32 163.367
R614 B.n850 B.n32 163.367
R615 B.n491 B.n489 163.367
R616 B.n489 B.n488 163.367
R617 B.n485 B.n484 163.367
R618 B.n482 B.n150 163.367
R619 B.n478 B.n476 163.367
R620 B.n474 B.n152 163.367
R621 B.n470 B.n468 163.367
R622 B.n466 B.n154 163.367
R623 B.n462 B.n460 163.367
R624 B.n458 B.n156 163.367
R625 B.n454 B.n452 163.367
R626 B.n450 B.n158 163.367
R627 B.n446 B.n444 163.367
R628 B.n442 B.n160 163.367
R629 B.n438 B.n436 163.367
R630 B.n434 B.n162 163.367
R631 B.n430 B.n428 163.367
R632 B.n426 B.n164 163.367
R633 B.n422 B.n420 163.367
R634 B.n418 B.n166 163.367
R635 B.n414 B.n412 163.367
R636 B.n410 B.n168 163.367
R637 B.n406 B.n404 163.367
R638 B.n402 B.n170 163.367
R639 B.n398 B.n396 163.367
R640 B.n394 B.n172 163.367
R641 B.n390 B.n388 163.367
R642 B.n386 B.n174 163.367
R643 B.n382 B.n380 163.367
R644 B.n378 B.n176 163.367
R645 B.n374 B.n372 163.367
R646 B.n370 B.n178 163.367
R647 B.n365 B.n363 163.367
R648 B.n361 B.n182 163.367
R649 B.n357 B.n355 163.367
R650 B.n353 B.n184 163.367
R651 B.n349 B.n347 163.367
R652 B.n345 B.n186 163.367
R653 B.n341 B.n339 163.367
R654 B.n337 B.n191 163.367
R655 B.n333 B.n331 163.367
R656 B.n329 B.n193 163.367
R657 B.n325 B.n323 163.367
R658 B.n321 B.n195 163.367
R659 B.n317 B.n315 163.367
R660 B.n313 B.n197 163.367
R661 B.n309 B.n307 163.367
R662 B.n305 B.n199 163.367
R663 B.n301 B.n299 163.367
R664 B.n297 B.n201 163.367
R665 B.n293 B.n291 163.367
R666 B.n289 B.n203 163.367
R667 B.n285 B.n283 163.367
R668 B.n281 B.n205 163.367
R669 B.n277 B.n275 163.367
R670 B.n273 B.n207 163.367
R671 B.n269 B.n267 163.367
R672 B.n265 B.n209 163.367
R673 B.n261 B.n259 163.367
R674 B.n257 B.n211 163.367
R675 B.n253 B.n251 163.367
R676 B.n249 B.n213 163.367
R677 B.n245 B.n243 163.367
R678 B.n241 B.n215 163.367
R679 B.n237 B.n235 163.367
R680 B.n233 B.n217 163.367
R681 B.n229 B.n227 163.367
R682 B.n225 B.n219 163.367
R683 B.n221 B.n144 163.367
R684 B.n497 B.n142 163.367
R685 B.n501 B.n142 163.367
R686 B.n501 B.n135 163.367
R687 B.n509 B.n135 163.367
R688 B.n509 B.n133 163.367
R689 B.n513 B.n133 163.367
R690 B.n513 B.n128 163.367
R691 B.n521 B.n128 163.367
R692 B.n521 B.n126 163.367
R693 B.n525 B.n126 163.367
R694 B.n525 B.n119 163.367
R695 B.n533 B.n119 163.367
R696 B.n533 B.n117 163.367
R697 B.n538 B.n117 163.367
R698 B.n538 B.n112 163.367
R699 B.n546 B.n112 163.367
R700 B.n547 B.n546 163.367
R701 B.n547 B.n5 163.367
R702 B.n6 B.n5 163.367
R703 B.n7 B.n6 163.367
R704 B.n552 B.n7 163.367
R705 B.n552 B.n12 163.367
R706 B.n13 B.n12 163.367
R707 B.n14 B.n13 163.367
R708 B.n557 B.n14 163.367
R709 B.n557 B.n19 163.367
R710 B.n20 B.n19 163.367
R711 B.n21 B.n20 163.367
R712 B.n562 B.n21 163.367
R713 B.n562 B.n26 163.367
R714 B.n27 B.n26 163.367
R715 B.n28 B.n27 163.367
R716 B.n567 B.n28 163.367
R717 B.n567 B.n33 163.367
R718 B.n34 B.n33 163.367
R719 B.n35 B.n34 163.367
R720 B.n846 B.n844 163.367
R721 B.n842 B.n39 163.367
R722 B.n838 B.n836 163.367
R723 B.n834 B.n41 163.367
R724 B.n830 B.n828 163.367
R725 B.n826 B.n43 163.367
R726 B.n822 B.n820 163.367
R727 B.n818 B.n45 163.367
R728 B.n814 B.n812 163.367
R729 B.n810 B.n47 163.367
R730 B.n806 B.n804 163.367
R731 B.n802 B.n49 163.367
R732 B.n798 B.n796 163.367
R733 B.n794 B.n51 163.367
R734 B.n790 B.n788 163.367
R735 B.n786 B.n53 163.367
R736 B.n782 B.n780 163.367
R737 B.n778 B.n55 163.367
R738 B.n774 B.n772 163.367
R739 B.n770 B.n57 163.367
R740 B.n766 B.n764 163.367
R741 B.n762 B.n59 163.367
R742 B.n758 B.n756 163.367
R743 B.n754 B.n61 163.367
R744 B.n750 B.n748 163.367
R745 B.n746 B.n63 163.367
R746 B.n742 B.n740 163.367
R747 B.n738 B.n65 163.367
R748 B.n734 B.n732 163.367
R749 B.n730 B.n67 163.367
R750 B.n726 B.n724 163.367
R751 B.n722 B.n69 163.367
R752 B.n717 B.n715 163.367
R753 B.n713 B.n73 163.367
R754 B.n709 B.n707 163.367
R755 B.n705 B.n75 163.367
R756 B.n701 B.n699 163.367
R757 B.n696 B.n695 163.367
R758 B.n693 B.n81 163.367
R759 B.n689 B.n687 163.367
R760 B.n685 B.n83 163.367
R761 B.n681 B.n679 163.367
R762 B.n677 B.n85 163.367
R763 B.n673 B.n671 163.367
R764 B.n669 B.n87 163.367
R765 B.n665 B.n663 163.367
R766 B.n661 B.n89 163.367
R767 B.n657 B.n655 163.367
R768 B.n653 B.n91 163.367
R769 B.n649 B.n647 163.367
R770 B.n645 B.n93 163.367
R771 B.n641 B.n639 163.367
R772 B.n637 B.n95 163.367
R773 B.n633 B.n631 163.367
R774 B.n629 B.n97 163.367
R775 B.n625 B.n623 163.367
R776 B.n621 B.n99 163.367
R777 B.n617 B.n615 163.367
R778 B.n613 B.n101 163.367
R779 B.n609 B.n607 163.367
R780 B.n605 B.n103 163.367
R781 B.n601 B.n599 163.367
R782 B.n597 B.n105 163.367
R783 B.n593 B.n591 163.367
R784 B.n589 B.n107 163.367
R785 B.n585 B.n583 163.367
R786 B.n581 B.n109 163.367
R787 B.n577 B.n575 163.367
R788 B.n490 B.n146 71.676
R789 B.n488 B.n148 71.676
R790 B.n484 B.n483 71.676
R791 B.n477 B.n150 71.676
R792 B.n476 B.n475 71.676
R793 B.n469 B.n152 71.676
R794 B.n468 B.n467 71.676
R795 B.n461 B.n154 71.676
R796 B.n460 B.n459 71.676
R797 B.n453 B.n156 71.676
R798 B.n452 B.n451 71.676
R799 B.n445 B.n158 71.676
R800 B.n444 B.n443 71.676
R801 B.n437 B.n160 71.676
R802 B.n436 B.n435 71.676
R803 B.n429 B.n162 71.676
R804 B.n428 B.n427 71.676
R805 B.n421 B.n164 71.676
R806 B.n420 B.n419 71.676
R807 B.n413 B.n166 71.676
R808 B.n412 B.n411 71.676
R809 B.n405 B.n168 71.676
R810 B.n404 B.n403 71.676
R811 B.n397 B.n170 71.676
R812 B.n396 B.n395 71.676
R813 B.n389 B.n172 71.676
R814 B.n388 B.n387 71.676
R815 B.n381 B.n174 71.676
R816 B.n380 B.n379 71.676
R817 B.n373 B.n176 71.676
R818 B.n372 B.n371 71.676
R819 B.n364 B.n178 71.676
R820 B.n363 B.n362 71.676
R821 B.n356 B.n182 71.676
R822 B.n355 B.n354 71.676
R823 B.n348 B.n184 71.676
R824 B.n347 B.n346 71.676
R825 B.n340 B.n186 71.676
R826 B.n339 B.n338 71.676
R827 B.n332 B.n191 71.676
R828 B.n331 B.n330 71.676
R829 B.n324 B.n193 71.676
R830 B.n323 B.n322 71.676
R831 B.n316 B.n195 71.676
R832 B.n315 B.n314 71.676
R833 B.n308 B.n197 71.676
R834 B.n307 B.n306 71.676
R835 B.n300 B.n199 71.676
R836 B.n299 B.n298 71.676
R837 B.n292 B.n201 71.676
R838 B.n291 B.n290 71.676
R839 B.n284 B.n203 71.676
R840 B.n283 B.n282 71.676
R841 B.n276 B.n205 71.676
R842 B.n275 B.n274 71.676
R843 B.n268 B.n207 71.676
R844 B.n267 B.n266 71.676
R845 B.n260 B.n209 71.676
R846 B.n259 B.n258 71.676
R847 B.n252 B.n211 71.676
R848 B.n251 B.n250 71.676
R849 B.n244 B.n213 71.676
R850 B.n243 B.n242 71.676
R851 B.n236 B.n215 71.676
R852 B.n235 B.n234 71.676
R853 B.n228 B.n217 71.676
R854 B.n227 B.n226 71.676
R855 B.n220 B.n219 71.676
R856 B.n845 B.n37 71.676
R857 B.n844 B.n843 71.676
R858 B.n837 B.n39 71.676
R859 B.n836 B.n835 71.676
R860 B.n829 B.n41 71.676
R861 B.n828 B.n827 71.676
R862 B.n821 B.n43 71.676
R863 B.n820 B.n819 71.676
R864 B.n813 B.n45 71.676
R865 B.n812 B.n811 71.676
R866 B.n805 B.n47 71.676
R867 B.n804 B.n803 71.676
R868 B.n797 B.n49 71.676
R869 B.n796 B.n795 71.676
R870 B.n789 B.n51 71.676
R871 B.n788 B.n787 71.676
R872 B.n781 B.n53 71.676
R873 B.n780 B.n779 71.676
R874 B.n773 B.n55 71.676
R875 B.n772 B.n771 71.676
R876 B.n765 B.n57 71.676
R877 B.n764 B.n763 71.676
R878 B.n757 B.n59 71.676
R879 B.n756 B.n755 71.676
R880 B.n749 B.n61 71.676
R881 B.n748 B.n747 71.676
R882 B.n741 B.n63 71.676
R883 B.n740 B.n739 71.676
R884 B.n733 B.n65 71.676
R885 B.n732 B.n731 71.676
R886 B.n725 B.n67 71.676
R887 B.n724 B.n723 71.676
R888 B.n716 B.n69 71.676
R889 B.n715 B.n714 71.676
R890 B.n708 B.n73 71.676
R891 B.n707 B.n706 71.676
R892 B.n700 B.n75 71.676
R893 B.n699 B.n79 71.676
R894 B.n695 B.n694 71.676
R895 B.n688 B.n81 71.676
R896 B.n687 B.n686 71.676
R897 B.n680 B.n83 71.676
R898 B.n679 B.n678 71.676
R899 B.n672 B.n85 71.676
R900 B.n671 B.n670 71.676
R901 B.n664 B.n87 71.676
R902 B.n663 B.n662 71.676
R903 B.n656 B.n89 71.676
R904 B.n655 B.n654 71.676
R905 B.n648 B.n91 71.676
R906 B.n647 B.n646 71.676
R907 B.n640 B.n93 71.676
R908 B.n639 B.n638 71.676
R909 B.n632 B.n95 71.676
R910 B.n631 B.n630 71.676
R911 B.n624 B.n97 71.676
R912 B.n623 B.n622 71.676
R913 B.n616 B.n99 71.676
R914 B.n615 B.n614 71.676
R915 B.n608 B.n101 71.676
R916 B.n607 B.n606 71.676
R917 B.n600 B.n103 71.676
R918 B.n599 B.n598 71.676
R919 B.n592 B.n105 71.676
R920 B.n591 B.n590 71.676
R921 B.n584 B.n107 71.676
R922 B.n583 B.n582 71.676
R923 B.n576 B.n109 71.676
R924 B.n575 B.n574 71.676
R925 B.n574 B.n573 71.676
R926 B.n577 B.n576 71.676
R927 B.n582 B.n581 71.676
R928 B.n585 B.n584 71.676
R929 B.n590 B.n589 71.676
R930 B.n593 B.n592 71.676
R931 B.n598 B.n597 71.676
R932 B.n601 B.n600 71.676
R933 B.n606 B.n605 71.676
R934 B.n609 B.n608 71.676
R935 B.n614 B.n613 71.676
R936 B.n617 B.n616 71.676
R937 B.n622 B.n621 71.676
R938 B.n625 B.n624 71.676
R939 B.n630 B.n629 71.676
R940 B.n633 B.n632 71.676
R941 B.n638 B.n637 71.676
R942 B.n641 B.n640 71.676
R943 B.n646 B.n645 71.676
R944 B.n649 B.n648 71.676
R945 B.n654 B.n653 71.676
R946 B.n657 B.n656 71.676
R947 B.n662 B.n661 71.676
R948 B.n665 B.n664 71.676
R949 B.n670 B.n669 71.676
R950 B.n673 B.n672 71.676
R951 B.n678 B.n677 71.676
R952 B.n681 B.n680 71.676
R953 B.n686 B.n685 71.676
R954 B.n689 B.n688 71.676
R955 B.n694 B.n693 71.676
R956 B.n696 B.n79 71.676
R957 B.n701 B.n700 71.676
R958 B.n706 B.n705 71.676
R959 B.n709 B.n708 71.676
R960 B.n714 B.n713 71.676
R961 B.n717 B.n716 71.676
R962 B.n723 B.n722 71.676
R963 B.n726 B.n725 71.676
R964 B.n731 B.n730 71.676
R965 B.n734 B.n733 71.676
R966 B.n739 B.n738 71.676
R967 B.n742 B.n741 71.676
R968 B.n747 B.n746 71.676
R969 B.n750 B.n749 71.676
R970 B.n755 B.n754 71.676
R971 B.n758 B.n757 71.676
R972 B.n763 B.n762 71.676
R973 B.n766 B.n765 71.676
R974 B.n771 B.n770 71.676
R975 B.n774 B.n773 71.676
R976 B.n779 B.n778 71.676
R977 B.n782 B.n781 71.676
R978 B.n787 B.n786 71.676
R979 B.n790 B.n789 71.676
R980 B.n795 B.n794 71.676
R981 B.n798 B.n797 71.676
R982 B.n803 B.n802 71.676
R983 B.n806 B.n805 71.676
R984 B.n811 B.n810 71.676
R985 B.n814 B.n813 71.676
R986 B.n819 B.n818 71.676
R987 B.n822 B.n821 71.676
R988 B.n827 B.n826 71.676
R989 B.n830 B.n829 71.676
R990 B.n835 B.n834 71.676
R991 B.n838 B.n837 71.676
R992 B.n843 B.n842 71.676
R993 B.n846 B.n845 71.676
R994 B.n491 B.n490 71.676
R995 B.n485 B.n148 71.676
R996 B.n483 B.n482 71.676
R997 B.n478 B.n477 71.676
R998 B.n475 B.n474 71.676
R999 B.n470 B.n469 71.676
R1000 B.n467 B.n466 71.676
R1001 B.n462 B.n461 71.676
R1002 B.n459 B.n458 71.676
R1003 B.n454 B.n453 71.676
R1004 B.n451 B.n450 71.676
R1005 B.n446 B.n445 71.676
R1006 B.n443 B.n442 71.676
R1007 B.n438 B.n437 71.676
R1008 B.n435 B.n434 71.676
R1009 B.n430 B.n429 71.676
R1010 B.n427 B.n426 71.676
R1011 B.n422 B.n421 71.676
R1012 B.n419 B.n418 71.676
R1013 B.n414 B.n413 71.676
R1014 B.n411 B.n410 71.676
R1015 B.n406 B.n405 71.676
R1016 B.n403 B.n402 71.676
R1017 B.n398 B.n397 71.676
R1018 B.n395 B.n394 71.676
R1019 B.n390 B.n389 71.676
R1020 B.n387 B.n386 71.676
R1021 B.n382 B.n381 71.676
R1022 B.n379 B.n378 71.676
R1023 B.n374 B.n373 71.676
R1024 B.n371 B.n370 71.676
R1025 B.n365 B.n364 71.676
R1026 B.n362 B.n361 71.676
R1027 B.n357 B.n356 71.676
R1028 B.n354 B.n353 71.676
R1029 B.n349 B.n348 71.676
R1030 B.n346 B.n345 71.676
R1031 B.n341 B.n340 71.676
R1032 B.n338 B.n337 71.676
R1033 B.n333 B.n332 71.676
R1034 B.n330 B.n329 71.676
R1035 B.n325 B.n324 71.676
R1036 B.n322 B.n321 71.676
R1037 B.n317 B.n316 71.676
R1038 B.n314 B.n313 71.676
R1039 B.n309 B.n308 71.676
R1040 B.n306 B.n305 71.676
R1041 B.n301 B.n300 71.676
R1042 B.n298 B.n297 71.676
R1043 B.n293 B.n292 71.676
R1044 B.n290 B.n289 71.676
R1045 B.n285 B.n284 71.676
R1046 B.n282 B.n281 71.676
R1047 B.n277 B.n276 71.676
R1048 B.n274 B.n273 71.676
R1049 B.n269 B.n268 71.676
R1050 B.n266 B.n265 71.676
R1051 B.n261 B.n260 71.676
R1052 B.n258 B.n257 71.676
R1053 B.n253 B.n252 71.676
R1054 B.n250 B.n249 71.676
R1055 B.n245 B.n244 71.676
R1056 B.n242 B.n241 71.676
R1057 B.n237 B.n236 71.676
R1058 B.n234 B.n233 71.676
R1059 B.n229 B.n228 71.676
R1060 B.n226 B.n225 71.676
R1061 B.n221 B.n220 71.676
R1062 B.n189 B.n188 59.5399
R1063 B.n367 B.n180 59.5399
R1064 B.n720 B.n71 59.5399
R1065 B.n78 B.n77 59.5399
R1066 B.n496 B.n145 56.0711
R1067 B.n851 B.n36 56.0711
R1068 B.n188 B.n187 32.7763
R1069 B.n180 B.n179 32.7763
R1070 B.n71 B.n70 32.7763
R1071 B.n77 B.n76 32.7763
R1072 B.n849 B.n848 31.6883
R1073 B.n572 B.n571 31.6883
R1074 B.n498 B.n143 31.6883
R1075 B.n494 B.n493 31.6883
R1076 B.n496 B.n141 30.0226
R1077 B.n502 B.n141 30.0226
R1078 B.n502 B.n136 30.0226
R1079 B.n508 B.n136 30.0226
R1080 B.n508 B.n137 30.0226
R1081 B.n514 B.n129 30.0226
R1082 B.n520 B.n129 30.0226
R1083 B.n520 B.n125 30.0226
R1084 B.n526 B.n125 30.0226
R1085 B.n526 B.n120 30.0226
R1086 B.n532 B.n120 30.0226
R1087 B.n532 B.n121 30.0226
R1088 B.n539 B.n113 30.0226
R1089 B.n545 B.n113 30.0226
R1090 B.n545 B.n4 30.0226
R1091 B.n885 B.n4 30.0226
R1092 B.n885 B.n884 30.0226
R1093 B.n884 B.n883 30.0226
R1094 B.n883 B.n8 30.0226
R1095 B.n877 B.n8 30.0226
R1096 B.n876 B.n875 30.0226
R1097 B.n875 B.n15 30.0226
R1098 B.n869 B.n15 30.0226
R1099 B.n869 B.n868 30.0226
R1100 B.n868 B.n867 30.0226
R1101 B.n867 B.n22 30.0226
R1102 B.n861 B.n22 30.0226
R1103 B.n860 B.n859 30.0226
R1104 B.n859 B.n29 30.0226
R1105 B.n853 B.n29 30.0226
R1106 B.n853 B.n852 30.0226
R1107 B.n852 B.n851 30.0226
R1108 B.n121 B.t0 27.3736
R1109 B.t1 B.n876 27.3736
R1110 B.n137 B.t3 22.0756
R1111 B.t7 B.n860 22.0756
R1112 B B.n887 18.0485
R1113 B.n848 B.n847 10.6151
R1114 B.n847 B.n38 10.6151
R1115 B.n841 B.n38 10.6151
R1116 B.n841 B.n840 10.6151
R1117 B.n840 B.n839 10.6151
R1118 B.n839 B.n40 10.6151
R1119 B.n833 B.n40 10.6151
R1120 B.n833 B.n832 10.6151
R1121 B.n832 B.n831 10.6151
R1122 B.n831 B.n42 10.6151
R1123 B.n825 B.n42 10.6151
R1124 B.n825 B.n824 10.6151
R1125 B.n824 B.n823 10.6151
R1126 B.n823 B.n44 10.6151
R1127 B.n817 B.n44 10.6151
R1128 B.n817 B.n816 10.6151
R1129 B.n816 B.n815 10.6151
R1130 B.n815 B.n46 10.6151
R1131 B.n809 B.n46 10.6151
R1132 B.n809 B.n808 10.6151
R1133 B.n808 B.n807 10.6151
R1134 B.n807 B.n48 10.6151
R1135 B.n801 B.n48 10.6151
R1136 B.n801 B.n800 10.6151
R1137 B.n800 B.n799 10.6151
R1138 B.n799 B.n50 10.6151
R1139 B.n793 B.n50 10.6151
R1140 B.n793 B.n792 10.6151
R1141 B.n792 B.n791 10.6151
R1142 B.n791 B.n52 10.6151
R1143 B.n785 B.n52 10.6151
R1144 B.n785 B.n784 10.6151
R1145 B.n784 B.n783 10.6151
R1146 B.n783 B.n54 10.6151
R1147 B.n777 B.n54 10.6151
R1148 B.n777 B.n776 10.6151
R1149 B.n776 B.n775 10.6151
R1150 B.n775 B.n56 10.6151
R1151 B.n769 B.n56 10.6151
R1152 B.n769 B.n768 10.6151
R1153 B.n768 B.n767 10.6151
R1154 B.n767 B.n58 10.6151
R1155 B.n761 B.n58 10.6151
R1156 B.n761 B.n760 10.6151
R1157 B.n760 B.n759 10.6151
R1158 B.n759 B.n60 10.6151
R1159 B.n753 B.n60 10.6151
R1160 B.n753 B.n752 10.6151
R1161 B.n752 B.n751 10.6151
R1162 B.n751 B.n62 10.6151
R1163 B.n745 B.n62 10.6151
R1164 B.n745 B.n744 10.6151
R1165 B.n744 B.n743 10.6151
R1166 B.n743 B.n64 10.6151
R1167 B.n737 B.n64 10.6151
R1168 B.n737 B.n736 10.6151
R1169 B.n736 B.n735 10.6151
R1170 B.n735 B.n66 10.6151
R1171 B.n729 B.n66 10.6151
R1172 B.n729 B.n728 10.6151
R1173 B.n728 B.n727 10.6151
R1174 B.n727 B.n68 10.6151
R1175 B.n721 B.n68 10.6151
R1176 B.n719 B.n718 10.6151
R1177 B.n718 B.n72 10.6151
R1178 B.n712 B.n72 10.6151
R1179 B.n712 B.n711 10.6151
R1180 B.n711 B.n710 10.6151
R1181 B.n710 B.n74 10.6151
R1182 B.n704 B.n74 10.6151
R1183 B.n704 B.n703 10.6151
R1184 B.n703 B.n702 10.6151
R1185 B.n698 B.n697 10.6151
R1186 B.n697 B.n80 10.6151
R1187 B.n692 B.n80 10.6151
R1188 B.n692 B.n691 10.6151
R1189 B.n691 B.n690 10.6151
R1190 B.n690 B.n82 10.6151
R1191 B.n684 B.n82 10.6151
R1192 B.n684 B.n683 10.6151
R1193 B.n683 B.n682 10.6151
R1194 B.n682 B.n84 10.6151
R1195 B.n676 B.n84 10.6151
R1196 B.n676 B.n675 10.6151
R1197 B.n675 B.n674 10.6151
R1198 B.n674 B.n86 10.6151
R1199 B.n668 B.n86 10.6151
R1200 B.n668 B.n667 10.6151
R1201 B.n667 B.n666 10.6151
R1202 B.n666 B.n88 10.6151
R1203 B.n660 B.n88 10.6151
R1204 B.n660 B.n659 10.6151
R1205 B.n659 B.n658 10.6151
R1206 B.n658 B.n90 10.6151
R1207 B.n652 B.n90 10.6151
R1208 B.n652 B.n651 10.6151
R1209 B.n651 B.n650 10.6151
R1210 B.n650 B.n92 10.6151
R1211 B.n644 B.n92 10.6151
R1212 B.n644 B.n643 10.6151
R1213 B.n643 B.n642 10.6151
R1214 B.n642 B.n94 10.6151
R1215 B.n636 B.n94 10.6151
R1216 B.n636 B.n635 10.6151
R1217 B.n635 B.n634 10.6151
R1218 B.n634 B.n96 10.6151
R1219 B.n628 B.n96 10.6151
R1220 B.n628 B.n627 10.6151
R1221 B.n627 B.n626 10.6151
R1222 B.n626 B.n98 10.6151
R1223 B.n620 B.n98 10.6151
R1224 B.n620 B.n619 10.6151
R1225 B.n619 B.n618 10.6151
R1226 B.n618 B.n100 10.6151
R1227 B.n612 B.n100 10.6151
R1228 B.n612 B.n611 10.6151
R1229 B.n611 B.n610 10.6151
R1230 B.n610 B.n102 10.6151
R1231 B.n604 B.n102 10.6151
R1232 B.n604 B.n603 10.6151
R1233 B.n603 B.n602 10.6151
R1234 B.n602 B.n104 10.6151
R1235 B.n596 B.n104 10.6151
R1236 B.n596 B.n595 10.6151
R1237 B.n595 B.n594 10.6151
R1238 B.n594 B.n106 10.6151
R1239 B.n588 B.n106 10.6151
R1240 B.n588 B.n587 10.6151
R1241 B.n587 B.n586 10.6151
R1242 B.n586 B.n108 10.6151
R1243 B.n580 B.n108 10.6151
R1244 B.n580 B.n579 10.6151
R1245 B.n579 B.n578 10.6151
R1246 B.n578 B.n110 10.6151
R1247 B.n572 B.n110 10.6151
R1248 B.n499 B.n498 10.6151
R1249 B.n500 B.n499 10.6151
R1250 B.n500 B.n134 10.6151
R1251 B.n510 B.n134 10.6151
R1252 B.n511 B.n510 10.6151
R1253 B.n512 B.n511 10.6151
R1254 B.n512 B.n127 10.6151
R1255 B.n522 B.n127 10.6151
R1256 B.n523 B.n522 10.6151
R1257 B.n524 B.n523 10.6151
R1258 B.n524 B.n118 10.6151
R1259 B.n534 B.n118 10.6151
R1260 B.n535 B.n534 10.6151
R1261 B.n537 B.n535 10.6151
R1262 B.n537 B.n536 10.6151
R1263 B.n536 B.n111 10.6151
R1264 B.n548 B.n111 10.6151
R1265 B.n549 B.n548 10.6151
R1266 B.n550 B.n549 10.6151
R1267 B.n551 B.n550 10.6151
R1268 B.n553 B.n551 10.6151
R1269 B.n554 B.n553 10.6151
R1270 B.n555 B.n554 10.6151
R1271 B.n556 B.n555 10.6151
R1272 B.n558 B.n556 10.6151
R1273 B.n559 B.n558 10.6151
R1274 B.n560 B.n559 10.6151
R1275 B.n561 B.n560 10.6151
R1276 B.n563 B.n561 10.6151
R1277 B.n564 B.n563 10.6151
R1278 B.n565 B.n564 10.6151
R1279 B.n566 B.n565 10.6151
R1280 B.n568 B.n566 10.6151
R1281 B.n569 B.n568 10.6151
R1282 B.n570 B.n569 10.6151
R1283 B.n571 B.n570 10.6151
R1284 B.n493 B.n492 10.6151
R1285 B.n492 B.n147 10.6151
R1286 B.n487 B.n147 10.6151
R1287 B.n487 B.n486 10.6151
R1288 B.n486 B.n149 10.6151
R1289 B.n481 B.n149 10.6151
R1290 B.n481 B.n480 10.6151
R1291 B.n480 B.n479 10.6151
R1292 B.n479 B.n151 10.6151
R1293 B.n473 B.n151 10.6151
R1294 B.n473 B.n472 10.6151
R1295 B.n472 B.n471 10.6151
R1296 B.n471 B.n153 10.6151
R1297 B.n465 B.n153 10.6151
R1298 B.n465 B.n464 10.6151
R1299 B.n464 B.n463 10.6151
R1300 B.n463 B.n155 10.6151
R1301 B.n457 B.n155 10.6151
R1302 B.n457 B.n456 10.6151
R1303 B.n456 B.n455 10.6151
R1304 B.n455 B.n157 10.6151
R1305 B.n449 B.n157 10.6151
R1306 B.n449 B.n448 10.6151
R1307 B.n448 B.n447 10.6151
R1308 B.n447 B.n159 10.6151
R1309 B.n441 B.n159 10.6151
R1310 B.n441 B.n440 10.6151
R1311 B.n440 B.n439 10.6151
R1312 B.n439 B.n161 10.6151
R1313 B.n433 B.n161 10.6151
R1314 B.n433 B.n432 10.6151
R1315 B.n432 B.n431 10.6151
R1316 B.n431 B.n163 10.6151
R1317 B.n425 B.n163 10.6151
R1318 B.n425 B.n424 10.6151
R1319 B.n424 B.n423 10.6151
R1320 B.n423 B.n165 10.6151
R1321 B.n417 B.n165 10.6151
R1322 B.n417 B.n416 10.6151
R1323 B.n416 B.n415 10.6151
R1324 B.n415 B.n167 10.6151
R1325 B.n409 B.n167 10.6151
R1326 B.n409 B.n408 10.6151
R1327 B.n408 B.n407 10.6151
R1328 B.n407 B.n169 10.6151
R1329 B.n401 B.n169 10.6151
R1330 B.n401 B.n400 10.6151
R1331 B.n400 B.n399 10.6151
R1332 B.n399 B.n171 10.6151
R1333 B.n393 B.n171 10.6151
R1334 B.n393 B.n392 10.6151
R1335 B.n392 B.n391 10.6151
R1336 B.n391 B.n173 10.6151
R1337 B.n385 B.n173 10.6151
R1338 B.n385 B.n384 10.6151
R1339 B.n384 B.n383 10.6151
R1340 B.n383 B.n175 10.6151
R1341 B.n377 B.n175 10.6151
R1342 B.n377 B.n376 10.6151
R1343 B.n376 B.n375 10.6151
R1344 B.n375 B.n177 10.6151
R1345 B.n369 B.n177 10.6151
R1346 B.n369 B.n368 10.6151
R1347 B.n366 B.n181 10.6151
R1348 B.n360 B.n181 10.6151
R1349 B.n360 B.n359 10.6151
R1350 B.n359 B.n358 10.6151
R1351 B.n358 B.n183 10.6151
R1352 B.n352 B.n183 10.6151
R1353 B.n352 B.n351 10.6151
R1354 B.n351 B.n350 10.6151
R1355 B.n350 B.n185 10.6151
R1356 B.n344 B.n343 10.6151
R1357 B.n343 B.n342 10.6151
R1358 B.n342 B.n190 10.6151
R1359 B.n336 B.n190 10.6151
R1360 B.n336 B.n335 10.6151
R1361 B.n335 B.n334 10.6151
R1362 B.n334 B.n192 10.6151
R1363 B.n328 B.n192 10.6151
R1364 B.n328 B.n327 10.6151
R1365 B.n327 B.n326 10.6151
R1366 B.n326 B.n194 10.6151
R1367 B.n320 B.n194 10.6151
R1368 B.n320 B.n319 10.6151
R1369 B.n319 B.n318 10.6151
R1370 B.n318 B.n196 10.6151
R1371 B.n312 B.n196 10.6151
R1372 B.n312 B.n311 10.6151
R1373 B.n311 B.n310 10.6151
R1374 B.n310 B.n198 10.6151
R1375 B.n304 B.n198 10.6151
R1376 B.n304 B.n303 10.6151
R1377 B.n303 B.n302 10.6151
R1378 B.n302 B.n200 10.6151
R1379 B.n296 B.n200 10.6151
R1380 B.n296 B.n295 10.6151
R1381 B.n295 B.n294 10.6151
R1382 B.n294 B.n202 10.6151
R1383 B.n288 B.n202 10.6151
R1384 B.n288 B.n287 10.6151
R1385 B.n287 B.n286 10.6151
R1386 B.n286 B.n204 10.6151
R1387 B.n280 B.n204 10.6151
R1388 B.n280 B.n279 10.6151
R1389 B.n279 B.n278 10.6151
R1390 B.n278 B.n206 10.6151
R1391 B.n272 B.n206 10.6151
R1392 B.n272 B.n271 10.6151
R1393 B.n271 B.n270 10.6151
R1394 B.n270 B.n208 10.6151
R1395 B.n264 B.n208 10.6151
R1396 B.n264 B.n263 10.6151
R1397 B.n263 B.n262 10.6151
R1398 B.n262 B.n210 10.6151
R1399 B.n256 B.n210 10.6151
R1400 B.n256 B.n255 10.6151
R1401 B.n255 B.n254 10.6151
R1402 B.n254 B.n212 10.6151
R1403 B.n248 B.n212 10.6151
R1404 B.n248 B.n247 10.6151
R1405 B.n247 B.n246 10.6151
R1406 B.n246 B.n214 10.6151
R1407 B.n240 B.n214 10.6151
R1408 B.n240 B.n239 10.6151
R1409 B.n239 B.n238 10.6151
R1410 B.n238 B.n216 10.6151
R1411 B.n232 B.n216 10.6151
R1412 B.n232 B.n231 10.6151
R1413 B.n231 B.n230 10.6151
R1414 B.n230 B.n218 10.6151
R1415 B.n224 B.n218 10.6151
R1416 B.n224 B.n223 10.6151
R1417 B.n223 B.n222 10.6151
R1418 B.n222 B.n143 10.6151
R1419 B.n494 B.n139 10.6151
R1420 B.n504 B.n139 10.6151
R1421 B.n505 B.n504 10.6151
R1422 B.n506 B.n505 10.6151
R1423 B.n506 B.n131 10.6151
R1424 B.n516 B.n131 10.6151
R1425 B.n517 B.n516 10.6151
R1426 B.n518 B.n517 10.6151
R1427 B.n518 B.n123 10.6151
R1428 B.n528 B.n123 10.6151
R1429 B.n529 B.n528 10.6151
R1430 B.n530 B.n529 10.6151
R1431 B.n530 B.n115 10.6151
R1432 B.n541 B.n115 10.6151
R1433 B.n542 B.n541 10.6151
R1434 B.n543 B.n542 10.6151
R1435 B.n543 B.n0 10.6151
R1436 B.n881 B.n1 10.6151
R1437 B.n881 B.n880 10.6151
R1438 B.n880 B.n879 10.6151
R1439 B.n879 B.n10 10.6151
R1440 B.n873 B.n10 10.6151
R1441 B.n873 B.n872 10.6151
R1442 B.n872 B.n871 10.6151
R1443 B.n871 B.n17 10.6151
R1444 B.n865 B.n17 10.6151
R1445 B.n865 B.n864 10.6151
R1446 B.n864 B.n863 10.6151
R1447 B.n863 B.n24 10.6151
R1448 B.n857 B.n24 10.6151
R1449 B.n857 B.n856 10.6151
R1450 B.n856 B.n855 10.6151
R1451 B.n855 B.n31 10.6151
R1452 B.n849 B.n31 10.6151
R1453 B.n721 B.n720 9.36635
R1454 B.n698 B.n78 9.36635
R1455 B.n368 B.n367 9.36635
R1456 B.n344 B.n189 9.36635
R1457 B.n514 B.t3 7.94752
R1458 B.n861 B.t7 7.94752
R1459 B.n887 B.n0 2.81026
R1460 B.n887 B.n1 2.81026
R1461 B.n539 B.t0 2.64951
R1462 B.n877 B.t1 2.64951
R1463 B.n720 B.n719 1.24928
R1464 B.n702 B.n78 1.24928
R1465 B.n367 B.n366 1.24928
R1466 B.n189 B.n185 1.24928
R1467 VP.n0 VP.t1 504.676
R1468 VP.n0 VP.t0 457.521
R1469 VP VP.n0 0.146778
R1470 VTAIL.n434 VTAIL.n330 289.615
R1471 VTAIL.n104 VTAIL.n0 289.615
R1472 VTAIL.n324 VTAIL.n220 289.615
R1473 VTAIL.n214 VTAIL.n110 289.615
R1474 VTAIL.n367 VTAIL.n366 185
R1475 VTAIL.n369 VTAIL.n368 185
R1476 VTAIL.n362 VTAIL.n361 185
R1477 VTAIL.n375 VTAIL.n374 185
R1478 VTAIL.n377 VTAIL.n376 185
R1479 VTAIL.n358 VTAIL.n357 185
R1480 VTAIL.n383 VTAIL.n382 185
R1481 VTAIL.n385 VTAIL.n384 185
R1482 VTAIL.n354 VTAIL.n353 185
R1483 VTAIL.n391 VTAIL.n390 185
R1484 VTAIL.n393 VTAIL.n392 185
R1485 VTAIL.n350 VTAIL.n349 185
R1486 VTAIL.n399 VTAIL.n398 185
R1487 VTAIL.n401 VTAIL.n400 185
R1488 VTAIL.n346 VTAIL.n345 185
R1489 VTAIL.n408 VTAIL.n407 185
R1490 VTAIL.n409 VTAIL.n344 185
R1491 VTAIL.n411 VTAIL.n410 185
R1492 VTAIL.n342 VTAIL.n341 185
R1493 VTAIL.n417 VTAIL.n416 185
R1494 VTAIL.n419 VTAIL.n418 185
R1495 VTAIL.n338 VTAIL.n337 185
R1496 VTAIL.n425 VTAIL.n424 185
R1497 VTAIL.n427 VTAIL.n426 185
R1498 VTAIL.n334 VTAIL.n333 185
R1499 VTAIL.n433 VTAIL.n432 185
R1500 VTAIL.n435 VTAIL.n434 185
R1501 VTAIL.n37 VTAIL.n36 185
R1502 VTAIL.n39 VTAIL.n38 185
R1503 VTAIL.n32 VTAIL.n31 185
R1504 VTAIL.n45 VTAIL.n44 185
R1505 VTAIL.n47 VTAIL.n46 185
R1506 VTAIL.n28 VTAIL.n27 185
R1507 VTAIL.n53 VTAIL.n52 185
R1508 VTAIL.n55 VTAIL.n54 185
R1509 VTAIL.n24 VTAIL.n23 185
R1510 VTAIL.n61 VTAIL.n60 185
R1511 VTAIL.n63 VTAIL.n62 185
R1512 VTAIL.n20 VTAIL.n19 185
R1513 VTAIL.n69 VTAIL.n68 185
R1514 VTAIL.n71 VTAIL.n70 185
R1515 VTAIL.n16 VTAIL.n15 185
R1516 VTAIL.n78 VTAIL.n77 185
R1517 VTAIL.n79 VTAIL.n14 185
R1518 VTAIL.n81 VTAIL.n80 185
R1519 VTAIL.n12 VTAIL.n11 185
R1520 VTAIL.n87 VTAIL.n86 185
R1521 VTAIL.n89 VTAIL.n88 185
R1522 VTAIL.n8 VTAIL.n7 185
R1523 VTAIL.n95 VTAIL.n94 185
R1524 VTAIL.n97 VTAIL.n96 185
R1525 VTAIL.n4 VTAIL.n3 185
R1526 VTAIL.n103 VTAIL.n102 185
R1527 VTAIL.n105 VTAIL.n104 185
R1528 VTAIL.n325 VTAIL.n324 185
R1529 VTAIL.n323 VTAIL.n322 185
R1530 VTAIL.n224 VTAIL.n223 185
R1531 VTAIL.n317 VTAIL.n316 185
R1532 VTAIL.n315 VTAIL.n314 185
R1533 VTAIL.n228 VTAIL.n227 185
R1534 VTAIL.n309 VTAIL.n308 185
R1535 VTAIL.n307 VTAIL.n306 185
R1536 VTAIL.n232 VTAIL.n231 185
R1537 VTAIL.n236 VTAIL.n234 185
R1538 VTAIL.n301 VTAIL.n300 185
R1539 VTAIL.n299 VTAIL.n298 185
R1540 VTAIL.n238 VTAIL.n237 185
R1541 VTAIL.n293 VTAIL.n292 185
R1542 VTAIL.n291 VTAIL.n290 185
R1543 VTAIL.n242 VTAIL.n241 185
R1544 VTAIL.n285 VTAIL.n284 185
R1545 VTAIL.n283 VTAIL.n282 185
R1546 VTAIL.n246 VTAIL.n245 185
R1547 VTAIL.n277 VTAIL.n276 185
R1548 VTAIL.n275 VTAIL.n274 185
R1549 VTAIL.n250 VTAIL.n249 185
R1550 VTAIL.n269 VTAIL.n268 185
R1551 VTAIL.n267 VTAIL.n266 185
R1552 VTAIL.n254 VTAIL.n253 185
R1553 VTAIL.n261 VTAIL.n260 185
R1554 VTAIL.n259 VTAIL.n258 185
R1555 VTAIL.n215 VTAIL.n214 185
R1556 VTAIL.n213 VTAIL.n212 185
R1557 VTAIL.n114 VTAIL.n113 185
R1558 VTAIL.n207 VTAIL.n206 185
R1559 VTAIL.n205 VTAIL.n204 185
R1560 VTAIL.n118 VTAIL.n117 185
R1561 VTAIL.n199 VTAIL.n198 185
R1562 VTAIL.n197 VTAIL.n196 185
R1563 VTAIL.n122 VTAIL.n121 185
R1564 VTAIL.n126 VTAIL.n124 185
R1565 VTAIL.n191 VTAIL.n190 185
R1566 VTAIL.n189 VTAIL.n188 185
R1567 VTAIL.n128 VTAIL.n127 185
R1568 VTAIL.n183 VTAIL.n182 185
R1569 VTAIL.n181 VTAIL.n180 185
R1570 VTAIL.n132 VTAIL.n131 185
R1571 VTAIL.n175 VTAIL.n174 185
R1572 VTAIL.n173 VTAIL.n172 185
R1573 VTAIL.n136 VTAIL.n135 185
R1574 VTAIL.n167 VTAIL.n166 185
R1575 VTAIL.n165 VTAIL.n164 185
R1576 VTAIL.n140 VTAIL.n139 185
R1577 VTAIL.n159 VTAIL.n158 185
R1578 VTAIL.n157 VTAIL.n156 185
R1579 VTAIL.n144 VTAIL.n143 185
R1580 VTAIL.n151 VTAIL.n150 185
R1581 VTAIL.n149 VTAIL.n148 185
R1582 VTAIL.n365 VTAIL.t1 147.659
R1583 VTAIL.n35 VTAIL.t3 147.659
R1584 VTAIL.n257 VTAIL.t2 147.659
R1585 VTAIL.n147 VTAIL.t0 147.659
R1586 VTAIL.n368 VTAIL.n367 104.615
R1587 VTAIL.n368 VTAIL.n361 104.615
R1588 VTAIL.n375 VTAIL.n361 104.615
R1589 VTAIL.n376 VTAIL.n375 104.615
R1590 VTAIL.n376 VTAIL.n357 104.615
R1591 VTAIL.n383 VTAIL.n357 104.615
R1592 VTAIL.n384 VTAIL.n383 104.615
R1593 VTAIL.n384 VTAIL.n353 104.615
R1594 VTAIL.n391 VTAIL.n353 104.615
R1595 VTAIL.n392 VTAIL.n391 104.615
R1596 VTAIL.n392 VTAIL.n349 104.615
R1597 VTAIL.n399 VTAIL.n349 104.615
R1598 VTAIL.n400 VTAIL.n399 104.615
R1599 VTAIL.n400 VTAIL.n345 104.615
R1600 VTAIL.n408 VTAIL.n345 104.615
R1601 VTAIL.n409 VTAIL.n408 104.615
R1602 VTAIL.n410 VTAIL.n409 104.615
R1603 VTAIL.n410 VTAIL.n341 104.615
R1604 VTAIL.n417 VTAIL.n341 104.615
R1605 VTAIL.n418 VTAIL.n417 104.615
R1606 VTAIL.n418 VTAIL.n337 104.615
R1607 VTAIL.n425 VTAIL.n337 104.615
R1608 VTAIL.n426 VTAIL.n425 104.615
R1609 VTAIL.n426 VTAIL.n333 104.615
R1610 VTAIL.n433 VTAIL.n333 104.615
R1611 VTAIL.n434 VTAIL.n433 104.615
R1612 VTAIL.n38 VTAIL.n37 104.615
R1613 VTAIL.n38 VTAIL.n31 104.615
R1614 VTAIL.n45 VTAIL.n31 104.615
R1615 VTAIL.n46 VTAIL.n45 104.615
R1616 VTAIL.n46 VTAIL.n27 104.615
R1617 VTAIL.n53 VTAIL.n27 104.615
R1618 VTAIL.n54 VTAIL.n53 104.615
R1619 VTAIL.n54 VTAIL.n23 104.615
R1620 VTAIL.n61 VTAIL.n23 104.615
R1621 VTAIL.n62 VTAIL.n61 104.615
R1622 VTAIL.n62 VTAIL.n19 104.615
R1623 VTAIL.n69 VTAIL.n19 104.615
R1624 VTAIL.n70 VTAIL.n69 104.615
R1625 VTAIL.n70 VTAIL.n15 104.615
R1626 VTAIL.n78 VTAIL.n15 104.615
R1627 VTAIL.n79 VTAIL.n78 104.615
R1628 VTAIL.n80 VTAIL.n79 104.615
R1629 VTAIL.n80 VTAIL.n11 104.615
R1630 VTAIL.n87 VTAIL.n11 104.615
R1631 VTAIL.n88 VTAIL.n87 104.615
R1632 VTAIL.n88 VTAIL.n7 104.615
R1633 VTAIL.n95 VTAIL.n7 104.615
R1634 VTAIL.n96 VTAIL.n95 104.615
R1635 VTAIL.n96 VTAIL.n3 104.615
R1636 VTAIL.n103 VTAIL.n3 104.615
R1637 VTAIL.n104 VTAIL.n103 104.615
R1638 VTAIL.n324 VTAIL.n323 104.615
R1639 VTAIL.n323 VTAIL.n223 104.615
R1640 VTAIL.n316 VTAIL.n223 104.615
R1641 VTAIL.n316 VTAIL.n315 104.615
R1642 VTAIL.n315 VTAIL.n227 104.615
R1643 VTAIL.n308 VTAIL.n227 104.615
R1644 VTAIL.n308 VTAIL.n307 104.615
R1645 VTAIL.n307 VTAIL.n231 104.615
R1646 VTAIL.n236 VTAIL.n231 104.615
R1647 VTAIL.n300 VTAIL.n236 104.615
R1648 VTAIL.n300 VTAIL.n299 104.615
R1649 VTAIL.n299 VTAIL.n237 104.615
R1650 VTAIL.n292 VTAIL.n237 104.615
R1651 VTAIL.n292 VTAIL.n291 104.615
R1652 VTAIL.n291 VTAIL.n241 104.615
R1653 VTAIL.n284 VTAIL.n241 104.615
R1654 VTAIL.n284 VTAIL.n283 104.615
R1655 VTAIL.n283 VTAIL.n245 104.615
R1656 VTAIL.n276 VTAIL.n245 104.615
R1657 VTAIL.n276 VTAIL.n275 104.615
R1658 VTAIL.n275 VTAIL.n249 104.615
R1659 VTAIL.n268 VTAIL.n249 104.615
R1660 VTAIL.n268 VTAIL.n267 104.615
R1661 VTAIL.n267 VTAIL.n253 104.615
R1662 VTAIL.n260 VTAIL.n253 104.615
R1663 VTAIL.n260 VTAIL.n259 104.615
R1664 VTAIL.n214 VTAIL.n213 104.615
R1665 VTAIL.n213 VTAIL.n113 104.615
R1666 VTAIL.n206 VTAIL.n113 104.615
R1667 VTAIL.n206 VTAIL.n205 104.615
R1668 VTAIL.n205 VTAIL.n117 104.615
R1669 VTAIL.n198 VTAIL.n117 104.615
R1670 VTAIL.n198 VTAIL.n197 104.615
R1671 VTAIL.n197 VTAIL.n121 104.615
R1672 VTAIL.n126 VTAIL.n121 104.615
R1673 VTAIL.n190 VTAIL.n126 104.615
R1674 VTAIL.n190 VTAIL.n189 104.615
R1675 VTAIL.n189 VTAIL.n127 104.615
R1676 VTAIL.n182 VTAIL.n127 104.615
R1677 VTAIL.n182 VTAIL.n181 104.615
R1678 VTAIL.n181 VTAIL.n131 104.615
R1679 VTAIL.n174 VTAIL.n131 104.615
R1680 VTAIL.n174 VTAIL.n173 104.615
R1681 VTAIL.n173 VTAIL.n135 104.615
R1682 VTAIL.n166 VTAIL.n135 104.615
R1683 VTAIL.n166 VTAIL.n165 104.615
R1684 VTAIL.n165 VTAIL.n139 104.615
R1685 VTAIL.n158 VTAIL.n139 104.615
R1686 VTAIL.n158 VTAIL.n157 104.615
R1687 VTAIL.n157 VTAIL.n143 104.615
R1688 VTAIL.n150 VTAIL.n143 104.615
R1689 VTAIL.n150 VTAIL.n149 104.615
R1690 VTAIL.n367 VTAIL.t1 52.3082
R1691 VTAIL.n37 VTAIL.t3 52.3082
R1692 VTAIL.n259 VTAIL.t2 52.3082
R1693 VTAIL.n149 VTAIL.t0 52.3082
R1694 VTAIL.n219 VTAIL.n109 32.2117
R1695 VTAIL.n439 VTAIL.n438 31.4096
R1696 VTAIL.n109 VTAIL.n108 31.4096
R1697 VTAIL.n329 VTAIL.n328 31.4096
R1698 VTAIL.n219 VTAIL.n218 31.4096
R1699 VTAIL.n439 VTAIL.n329 30.7548
R1700 VTAIL.n366 VTAIL.n365 15.6677
R1701 VTAIL.n36 VTAIL.n35 15.6677
R1702 VTAIL.n258 VTAIL.n257 15.6677
R1703 VTAIL.n148 VTAIL.n147 15.6677
R1704 VTAIL.n411 VTAIL.n342 13.1884
R1705 VTAIL.n81 VTAIL.n12 13.1884
R1706 VTAIL.n234 VTAIL.n232 13.1884
R1707 VTAIL.n124 VTAIL.n122 13.1884
R1708 VTAIL.n369 VTAIL.n364 12.8005
R1709 VTAIL.n412 VTAIL.n344 12.8005
R1710 VTAIL.n416 VTAIL.n415 12.8005
R1711 VTAIL.n39 VTAIL.n34 12.8005
R1712 VTAIL.n82 VTAIL.n14 12.8005
R1713 VTAIL.n86 VTAIL.n85 12.8005
R1714 VTAIL.n306 VTAIL.n305 12.8005
R1715 VTAIL.n302 VTAIL.n301 12.8005
R1716 VTAIL.n261 VTAIL.n256 12.8005
R1717 VTAIL.n196 VTAIL.n195 12.8005
R1718 VTAIL.n192 VTAIL.n191 12.8005
R1719 VTAIL.n151 VTAIL.n146 12.8005
R1720 VTAIL.n370 VTAIL.n362 12.0247
R1721 VTAIL.n407 VTAIL.n406 12.0247
R1722 VTAIL.n419 VTAIL.n340 12.0247
R1723 VTAIL.n40 VTAIL.n32 12.0247
R1724 VTAIL.n77 VTAIL.n76 12.0247
R1725 VTAIL.n89 VTAIL.n10 12.0247
R1726 VTAIL.n309 VTAIL.n230 12.0247
R1727 VTAIL.n298 VTAIL.n235 12.0247
R1728 VTAIL.n262 VTAIL.n254 12.0247
R1729 VTAIL.n199 VTAIL.n120 12.0247
R1730 VTAIL.n188 VTAIL.n125 12.0247
R1731 VTAIL.n152 VTAIL.n144 12.0247
R1732 VTAIL.n374 VTAIL.n373 11.249
R1733 VTAIL.n405 VTAIL.n346 11.249
R1734 VTAIL.n420 VTAIL.n338 11.249
R1735 VTAIL.n44 VTAIL.n43 11.249
R1736 VTAIL.n75 VTAIL.n16 11.249
R1737 VTAIL.n90 VTAIL.n8 11.249
R1738 VTAIL.n310 VTAIL.n228 11.249
R1739 VTAIL.n297 VTAIL.n238 11.249
R1740 VTAIL.n266 VTAIL.n265 11.249
R1741 VTAIL.n200 VTAIL.n118 11.249
R1742 VTAIL.n187 VTAIL.n128 11.249
R1743 VTAIL.n156 VTAIL.n155 11.249
R1744 VTAIL.n377 VTAIL.n360 10.4732
R1745 VTAIL.n402 VTAIL.n401 10.4732
R1746 VTAIL.n424 VTAIL.n423 10.4732
R1747 VTAIL.n47 VTAIL.n30 10.4732
R1748 VTAIL.n72 VTAIL.n71 10.4732
R1749 VTAIL.n94 VTAIL.n93 10.4732
R1750 VTAIL.n314 VTAIL.n313 10.4732
R1751 VTAIL.n294 VTAIL.n293 10.4732
R1752 VTAIL.n269 VTAIL.n252 10.4732
R1753 VTAIL.n204 VTAIL.n203 10.4732
R1754 VTAIL.n184 VTAIL.n183 10.4732
R1755 VTAIL.n159 VTAIL.n142 10.4732
R1756 VTAIL.n378 VTAIL.n358 9.69747
R1757 VTAIL.n398 VTAIL.n348 9.69747
R1758 VTAIL.n427 VTAIL.n336 9.69747
R1759 VTAIL.n48 VTAIL.n28 9.69747
R1760 VTAIL.n68 VTAIL.n18 9.69747
R1761 VTAIL.n97 VTAIL.n6 9.69747
R1762 VTAIL.n317 VTAIL.n226 9.69747
R1763 VTAIL.n290 VTAIL.n240 9.69747
R1764 VTAIL.n270 VTAIL.n250 9.69747
R1765 VTAIL.n207 VTAIL.n116 9.69747
R1766 VTAIL.n180 VTAIL.n130 9.69747
R1767 VTAIL.n160 VTAIL.n140 9.69747
R1768 VTAIL.n438 VTAIL.n437 9.45567
R1769 VTAIL.n108 VTAIL.n107 9.45567
R1770 VTAIL.n328 VTAIL.n327 9.45567
R1771 VTAIL.n218 VTAIL.n217 9.45567
R1772 VTAIL.n437 VTAIL.n436 9.3005
R1773 VTAIL.n431 VTAIL.n430 9.3005
R1774 VTAIL.n429 VTAIL.n428 9.3005
R1775 VTAIL.n336 VTAIL.n335 9.3005
R1776 VTAIL.n423 VTAIL.n422 9.3005
R1777 VTAIL.n421 VTAIL.n420 9.3005
R1778 VTAIL.n340 VTAIL.n339 9.3005
R1779 VTAIL.n415 VTAIL.n414 9.3005
R1780 VTAIL.n387 VTAIL.n386 9.3005
R1781 VTAIL.n356 VTAIL.n355 9.3005
R1782 VTAIL.n381 VTAIL.n380 9.3005
R1783 VTAIL.n379 VTAIL.n378 9.3005
R1784 VTAIL.n360 VTAIL.n359 9.3005
R1785 VTAIL.n373 VTAIL.n372 9.3005
R1786 VTAIL.n371 VTAIL.n370 9.3005
R1787 VTAIL.n364 VTAIL.n363 9.3005
R1788 VTAIL.n389 VTAIL.n388 9.3005
R1789 VTAIL.n352 VTAIL.n351 9.3005
R1790 VTAIL.n395 VTAIL.n394 9.3005
R1791 VTAIL.n397 VTAIL.n396 9.3005
R1792 VTAIL.n348 VTAIL.n347 9.3005
R1793 VTAIL.n403 VTAIL.n402 9.3005
R1794 VTAIL.n405 VTAIL.n404 9.3005
R1795 VTAIL.n406 VTAIL.n343 9.3005
R1796 VTAIL.n413 VTAIL.n412 9.3005
R1797 VTAIL.n332 VTAIL.n331 9.3005
R1798 VTAIL.n107 VTAIL.n106 9.3005
R1799 VTAIL.n101 VTAIL.n100 9.3005
R1800 VTAIL.n99 VTAIL.n98 9.3005
R1801 VTAIL.n6 VTAIL.n5 9.3005
R1802 VTAIL.n93 VTAIL.n92 9.3005
R1803 VTAIL.n91 VTAIL.n90 9.3005
R1804 VTAIL.n10 VTAIL.n9 9.3005
R1805 VTAIL.n85 VTAIL.n84 9.3005
R1806 VTAIL.n57 VTAIL.n56 9.3005
R1807 VTAIL.n26 VTAIL.n25 9.3005
R1808 VTAIL.n51 VTAIL.n50 9.3005
R1809 VTAIL.n49 VTAIL.n48 9.3005
R1810 VTAIL.n30 VTAIL.n29 9.3005
R1811 VTAIL.n43 VTAIL.n42 9.3005
R1812 VTAIL.n41 VTAIL.n40 9.3005
R1813 VTAIL.n34 VTAIL.n33 9.3005
R1814 VTAIL.n59 VTAIL.n58 9.3005
R1815 VTAIL.n22 VTAIL.n21 9.3005
R1816 VTAIL.n65 VTAIL.n64 9.3005
R1817 VTAIL.n67 VTAIL.n66 9.3005
R1818 VTAIL.n18 VTAIL.n17 9.3005
R1819 VTAIL.n73 VTAIL.n72 9.3005
R1820 VTAIL.n75 VTAIL.n74 9.3005
R1821 VTAIL.n76 VTAIL.n13 9.3005
R1822 VTAIL.n83 VTAIL.n82 9.3005
R1823 VTAIL.n2 VTAIL.n1 9.3005
R1824 VTAIL.n244 VTAIL.n243 9.3005
R1825 VTAIL.n287 VTAIL.n286 9.3005
R1826 VTAIL.n289 VTAIL.n288 9.3005
R1827 VTAIL.n240 VTAIL.n239 9.3005
R1828 VTAIL.n295 VTAIL.n294 9.3005
R1829 VTAIL.n297 VTAIL.n296 9.3005
R1830 VTAIL.n235 VTAIL.n233 9.3005
R1831 VTAIL.n303 VTAIL.n302 9.3005
R1832 VTAIL.n327 VTAIL.n326 9.3005
R1833 VTAIL.n222 VTAIL.n221 9.3005
R1834 VTAIL.n321 VTAIL.n320 9.3005
R1835 VTAIL.n319 VTAIL.n318 9.3005
R1836 VTAIL.n226 VTAIL.n225 9.3005
R1837 VTAIL.n313 VTAIL.n312 9.3005
R1838 VTAIL.n311 VTAIL.n310 9.3005
R1839 VTAIL.n230 VTAIL.n229 9.3005
R1840 VTAIL.n305 VTAIL.n304 9.3005
R1841 VTAIL.n281 VTAIL.n280 9.3005
R1842 VTAIL.n279 VTAIL.n278 9.3005
R1843 VTAIL.n248 VTAIL.n247 9.3005
R1844 VTAIL.n273 VTAIL.n272 9.3005
R1845 VTAIL.n271 VTAIL.n270 9.3005
R1846 VTAIL.n252 VTAIL.n251 9.3005
R1847 VTAIL.n265 VTAIL.n264 9.3005
R1848 VTAIL.n263 VTAIL.n262 9.3005
R1849 VTAIL.n256 VTAIL.n255 9.3005
R1850 VTAIL.n134 VTAIL.n133 9.3005
R1851 VTAIL.n177 VTAIL.n176 9.3005
R1852 VTAIL.n179 VTAIL.n178 9.3005
R1853 VTAIL.n130 VTAIL.n129 9.3005
R1854 VTAIL.n185 VTAIL.n184 9.3005
R1855 VTAIL.n187 VTAIL.n186 9.3005
R1856 VTAIL.n125 VTAIL.n123 9.3005
R1857 VTAIL.n193 VTAIL.n192 9.3005
R1858 VTAIL.n217 VTAIL.n216 9.3005
R1859 VTAIL.n112 VTAIL.n111 9.3005
R1860 VTAIL.n211 VTAIL.n210 9.3005
R1861 VTAIL.n209 VTAIL.n208 9.3005
R1862 VTAIL.n116 VTAIL.n115 9.3005
R1863 VTAIL.n203 VTAIL.n202 9.3005
R1864 VTAIL.n201 VTAIL.n200 9.3005
R1865 VTAIL.n120 VTAIL.n119 9.3005
R1866 VTAIL.n195 VTAIL.n194 9.3005
R1867 VTAIL.n171 VTAIL.n170 9.3005
R1868 VTAIL.n169 VTAIL.n168 9.3005
R1869 VTAIL.n138 VTAIL.n137 9.3005
R1870 VTAIL.n163 VTAIL.n162 9.3005
R1871 VTAIL.n161 VTAIL.n160 9.3005
R1872 VTAIL.n142 VTAIL.n141 9.3005
R1873 VTAIL.n155 VTAIL.n154 9.3005
R1874 VTAIL.n153 VTAIL.n152 9.3005
R1875 VTAIL.n146 VTAIL.n145 9.3005
R1876 VTAIL.n382 VTAIL.n381 8.92171
R1877 VTAIL.n397 VTAIL.n350 8.92171
R1878 VTAIL.n428 VTAIL.n334 8.92171
R1879 VTAIL.n52 VTAIL.n51 8.92171
R1880 VTAIL.n67 VTAIL.n20 8.92171
R1881 VTAIL.n98 VTAIL.n4 8.92171
R1882 VTAIL.n318 VTAIL.n224 8.92171
R1883 VTAIL.n289 VTAIL.n242 8.92171
R1884 VTAIL.n274 VTAIL.n273 8.92171
R1885 VTAIL.n208 VTAIL.n114 8.92171
R1886 VTAIL.n179 VTAIL.n132 8.92171
R1887 VTAIL.n164 VTAIL.n163 8.92171
R1888 VTAIL.n385 VTAIL.n356 8.14595
R1889 VTAIL.n394 VTAIL.n393 8.14595
R1890 VTAIL.n432 VTAIL.n431 8.14595
R1891 VTAIL.n55 VTAIL.n26 8.14595
R1892 VTAIL.n64 VTAIL.n63 8.14595
R1893 VTAIL.n102 VTAIL.n101 8.14595
R1894 VTAIL.n322 VTAIL.n321 8.14595
R1895 VTAIL.n286 VTAIL.n285 8.14595
R1896 VTAIL.n277 VTAIL.n248 8.14595
R1897 VTAIL.n212 VTAIL.n211 8.14595
R1898 VTAIL.n176 VTAIL.n175 8.14595
R1899 VTAIL.n167 VTAIL.n138 8.14595
R1900 VTAIL.n386 VTAIL.n354 7.3702
R1901 VTAIL.n390 VTAIL.n352 7.3702
R1902 VTAIL.n435 VTAIL.n332 7.3702
R1903 VTAIL.n438 VTAIL.n330 7.3702
R1904 VTAIL.n56 VTAIL.n24 7.3702
R1905 VTAIL.n60 VTAIL.n22 7.3702
R1906 VTAIL.n105 VTAIL.n2 7.3702
R1907 VTAIL.n108 VTAIL.n0 7.3702
R1908 VTAIL.n328 VTAIL.n220 7.3702
R1909 VTAIL.n325 VTAIL.n222 7.3702
R1910 VTAIL.n282 VTAIL.n244 7.3702
R1911 VTAIL.n278 VTAIL.n246 7.3702
R1912 VTAIL.n218 VTAIL.n110 7.3702
R1913 VTAIL.n215 VTAIL.n112 7.3702
R1914 VTAIL.n172 VTAIL.n134 7.3702
R1915 VTAIL.n168 VTAIL.n136 7.3702
R1916 VTAIL.n389 VTAIL.n354 6.59444
R1917 VTAIL.n390 VTAIL.n389 6.59444
R1918 VTAIL.n436 VTAIL.n435 6.59444
R1919 VTAIL.n436 VTAIL.n330 6.59444
R1920 VTAIL.n59 VTAIL.n24 6.59444
R1921 VTAIL.n60 VTAIL.n59 6.59444
R1922 VTAIL.n106 VTAIL.n105 6.59444
R1923 VTAIL.n106 VTAIL.n0 6.59444
R1924 VTAIL.n326 VTAIL.n220 6.59444
R1925 VTAIL.n326 VTAIL.n325 6.59444
R1926 VTAIL.n282 VTAIL.n281 6.59444
R1927 VTAIL.n281 VTAIL.n246 6.59444
R1928 VTAIL.n216 VTAIL.n110 6.59444
R1929 VTAIL.n216 VTAIL.n215 6.59444
R1930 VTAIL.n172 VTAIL.n171 6.59444
R1931 VTAIL.n171 VTAIL.n136 6.59444
R1932 VTAIL.n386 VTAIL.n385 5.81868
R1933 VTAIL.n393 VTAIL.n352 5.81868
R1934 VTAIL.n432 VTAIL.n332 5.81868
R1935 VTAIL.n56 VTAIL.n55 5.81868
R1936 VTAIL.n63 VTAIL.n22 5.81868
R1937 VTAIL.n102 VTAIL.n2 5.81868
R1938 VTAIL.n322 VTAIL.n222 5.81868
R1939 VTAIL.n285 VTAIL.n244 5.81868
R1940 VTAIL.n278 VTAIL.n277 5.81868
R1941 VTAIL.n212 VTAIL.n112 5.81868
R1942 VTAIL.n175 VTAIL.n134 5.81868
R1943 VTAIL.n168 VTAIL.n167 5.81868
R1944 VTAIL.n382 VTAIL.n356 5.04292
R1945 VTAIL.n394 VTAIL.n350 5.04292
R1946 VTAIL.n431 VTAIL.n334 5.04292
R1947 VTAIL.n52 VTAIL.n26 5.04292
R1948 VTAIL.n64 VTAIL.n20 5.04292
R1949 VTAIL.n101 VTAIL.n4 5.04292
R1950 VTAIL.n321 VTAIL.n224 5.04292
R1951 VTAIL.n286 VTAIL.n242 5.04292
R1952 VTAIL.n274 VTAIL.n248 5.04292
R1953 VTAIL.n211 VTAIL.n114 5.04292
R1954 VTAIL.n176 VTAIL.n132 5.04292
R1955 VTAIL.n164 VTAIL.n138 5.04292
R1956 VTAIL.n365 VTAIL.n363 4.38563
R1957 VTAIL.n35 VTAIL.n33 4.38563
R1958 VTAIL.n257 VTAIL.n255 4.38563
R1959 VTAIL.n147 VTAIL.n145 4.38563
R1960 VTAIL.n381 VTAIL.n358 4.26717
R1961 VTAIL.n398 VTAIL.n397 4.26717
R1962 VTAIL.n428 VTAIL.n427 4.26717
R1963 VTAIL.n51 VTAIL.n28 4.26717
R1964 VTAIL.n68 VTAIL.n67 4.26717
R1965 VTAIL.n98 VTAIL.n97 4.26717
R1966 VTAIL.n318 VTAIL.n317 4.26717
R1967 VTAIL.n290 VTAIL.n289 4.26717
R1968 VTAIL.n273 VTAIL.n250 4.26717
R1969 VTAIL.n208 VTAIL.n207 4.26717
R1970 VTAIL.n180 VTAIL.n179 4.26717
R1971 VTAIL.n163 VTAIL.n140 4.26717
R1972 VTAIL.n378 VTAIL.n377 3.49141
R1973 VTAIL.n401 VTAIL.n348 3.49141
R1974 VTAIL.n424 VTAIL.n336 3.49141
R1975 VTAIL.n48 VTAIL.n47 3.49141
R1976 VTAIL.n71 VTAIL.n18 3.49141
R1977 VTAIL.n94 VTAIL.n6 3.49141
R1978 VTAIL.n314 VTAIL.n226 3.49141
R1979 VTAIL.n293 VTAIL.n240 3.49141
R1980 VTAIL.n270 VTAIL.n269 3.49141
R1981 VTAIL.n204 VTAIL.n116 3.49141
R1982 VTAIL.n183 VTAIL.n130 3.49141
R1983 VTAIL.n160 VTAIL.n159 3.49141
R1984 VTAIL.n374 VTAIL.n360 2.71565
R1985 VTAIL.n402 VTAIL.n346 2.71565
R1986 VTAIL.n423 VTAIL.n338 2.71565
R1987 VTAIL.n44 VTAIL.n30 2.71565
R1988 VTAIL.n72 VTAIL.n16 2.71565
R1989 VTAIL.n93 VTAIL.n8 2.71565
R1990 VTAIL.n313 VTAIL.n228 2.71565
R1991 VTAIL.n294 VTAIL.n238 2.71565
R1992 VTAIL.n266 VTAIL.n252 2.71565
R1993 VTAIL.n203 VTAIL.n118 2.71565
R1994 VTAIL.n184 VTAIL.n128 2.71565
R1995 VTAIL.n156 VTAIL.n142 2.71565
R1996 VTAIL.n373 VTAIL.n362 1.93989
R1997 VTAIL.n407 VTAIL.n405 1.93989
R1998 VTAIL.n420 VTAIL.n419 1.93989
R1999 VTAIL.n43 VTAIL.n32 1.93989
R2000 VTAIL.n77 VTAIL.n75 1.93989
R2001 VTAIL.n90 VTAIL.n89 1.93989
R2002 VTAIL.n310 VTAIL.n309 1.93989
R2003 VTAIL.n298 VTAIL.n297 1.93989
R2004 VTAIL.n265 VTAIL.n254 1.93989
R2005 VTAIL.n200 VTAIL.n199 1.93989
R2006 VTAIL.n188 VTAIL.n187 1.93989
R2007 VTAIL.n155 VTAIL.n144 1.93989
R2008 VTAIL.n329 VTAIL.n219 1.19878
R2009 VTAIL.n370 VTAIL.n369 1.16414
R2010 VTAIL.n406 VTAIL.n344 1.16414
R2011 VTAIL.n416 VTAIL.n340 1.16414
R2012 VTAIL.n40 VTAIL.n39 1.16414
R2013 VTAIL.n76 VTAIL.n14 1.16414
R2014 VTAIL.n86 VTAIL.n10 1.16414
R2015 VTAIL.n306 VTAIL.n230 1.16414
R2016 VTAIL.n301 VTAIL.n235 1.16414
R2017 VTAIL.n262 VTAIL.n261 1.16414
R2018 VTAIL.n196 VTAIL.n120 1.16414
R2019 VTAIL.n191 VTAIL.n125 1.16414
R2020 VTAIL.n152 VTAIL.n151 1.16414
R2021 VTAIL VTAIL.n109 0.892741
R2022 VTAIL.n366 VTAIL.n364 0.388379
R2023 VTAIL.n412 VTAIL.n411 0.388379
R2024 VTAIL.n415 VTAIL.n342 0.388379
R2025 VTAIL.n36 VTAIL.n34 0.388379
R2026 VTAIL.n82 VTAIL.n81 0.388379
R2027 VTAIL.n85 VTAIL.n12 0.388379
R2028 VTAIL.n305 VTAIL.n232 0.388379
R2029 VTAIL.n302 VTAIL.n234 0.388379
R2030 VTAIL.n258 VTAIL.n256 0.388379
R2031 VTAIL.n195 VTAIL.n122 0.388379
R2032 VTAIL.n192 VTAIL.n124 0.388379
R2033 VTAIL.n148 VTAIL.n146 0.388379
R2034 VTAIL VTAIL.n439 0.306534
R2035 VTAIL.n371 VTAIL.n363 0.155672
R2036 VTAIL.n372 VTAIL.n371 0.155672
R2037 VTAIL.n372 VTAIL.n359 0.155672
R2038 VTAIL.n379 VTAIL.n359 0.155672
R2039 VTAIL.n380 VTAIL.n379 0.155672
R2040 VTAIL.n380 VTAIL.n355 0.155672
R2041 VTAIL.n387 VTAIL.n355 0.155672
R2042 VTAIL.n388 VTAIL.n387 0.155672
R2043 VTAIL.n388 VTAIL.n351 0.155672
R2044 VTAIL.n395 VTAIL.n351 0.155672
R2045 VTAIL.n396 VTAIL.n395 0.155672
R2046 VTAIL.n396 VTAIL.n347 0.155672
R2047 VTAIL.n403 VTAIL.n347 0.155672
R2048 VTAIL.n404 VTAIL.n403 0.155672
R2049 VTAIL.n404 VTAIL.n343 0.155672
R2050 VTAIL.n413 VTAIL.n343 0.155672
R2051 VTAIL.n414 VTAIL.n413 0.155672
R2052 VTAIL.n414 VTAIL.n339 0.155672
R2053 VTAIL.n421 VTAIL.n339 0.155672
R2054 VTAIL.n422 VTAIL.n421 0.155672
R2055 VTAIL.n422 VTAIL.n335 0.155672
R2056 VTAIL.n429 VTAIL.n335 0.155672
R2057 VTAIL.n430 VTAIL.n429 0.155672
R2058 VTAIL.n430 VTAIL.n331 0.155672
R2059 VTAIL.n437 VTAIL.n331 0.155672
R2060 VTAIL.n41 VTAIL.n33 0.155672
R2061 VTAIL.n42 VTAIL.n41 0.155672
R2062 VTAIL.n42 VTAIL.n29 0.155672
R2063 VTAIL.n49 VTAIL.n29 0.155672
R2064 VTAIL.n50 VTAIL.n49 0.155672
R2065 VTAIL.n50 VTAIL.n25 0.155672
R2066 VTAIL.n57 VTAIL.n25 0.155672
R2067 VTAIL.n58 VTAIL.n57 0.155672
R2068 VTAIL.n58 VTAIL.n21 0.155672
R2069 VTAIL.n65 VTAIL.n21 0.155672
R2070 VTAIL.n66 VTAIL.n65 0.155672
R2071 VTAIL.n66 VTAIL.n17 0.155672
R2072 VTAIL.n73 VTAIL.n17 0.155672
R2073 VTAIL.n74 VTAIL.n73 0.155672
R2074 VTAIL.n74 VTAIL.n13 0.155672
R2075 VTAIL.n83 VTAIL.n13 0.155672
R2076 VTAIL.n84 VTAIL.n83 0.155672
R2077 VTAIL.n84 VTAIL.n9 0.155672
R2078 VTAIL.n91 VTAIL.n9 0.155672
R2079 VTAIL.n92 VTAIL.n91 0.155672
R2080 VTAIL.n92 VTAIL.n5 0.155672
R2081 VTAIL.n99 VTAIL.n5 0.155672
R2082 VTAIL.n100 VTAIL.n99 0.155672
R2083 VTAIL.n100 VTAIL.n1 0.155672
R2084 VTAIL.n107 VTAIL.n1 0.155672
R2085 VTAIL.n327 VTAIL.n221 0.155672
R2086 VTAIL.n320 VTAIL.n221 0.155672
R2087 VTAIL.n320 VTAIL.n319 0.155672
R2088 VTAIL.n319 VTAIL.n225 0.155672
R2089 VTAIL.n312 VTAIL.n225 0.155672
R2090 VTAIL.n312 VTAIL.n311 0.155672
R2091 VTAIL.n311 VTAIL.n229 0.155672
R2092 VTAIL.n304 VTAIL.n229 0.155672
R2093 VTAIL.n304 VTAIL.n303 0.155672
R2094 VTAIL.n303 VTAIL.n233 0.155672
R2095 VTAIL.n296 VTAIL.n233 0.155672
R2096 VTAIL.n296 VTAIL.n295 0.155672
R2097 VTAIL.n295 VTAIL.n239 0.155672
R2098 VTAIL.n288 VTAIL.n239 0.155672
R2099 VTAIL.n288 VTAIL.n287 0.155672
R2100 VTAIL.n287 VTAIL.n243 0.155672
R2101 VTAIL.n280 VTAIL.n243 0.155672
R2102 VTAIL.n280 VTAIL.n279 0.155672
R2103 VTAIL.n279 VTAIL.n247 0.155672
R2104 VTAIL.n272 VTAIL.n247 0.155672
R2105 VTAIL.n272 VTAIL.n271 0.155672
R2106 VTAIL.n271 VTAIL.n251 0.155672
R2107 VTAIL.n264 VTAIL.n251 0.155672
R2108 VTAIL.n264 VTAIL.n263 0.155672
R2109 VTAIL.n263 VTAIL.n255 0.155672
R2110 VTAIL.n217 VTAIL.n111 0.155672
R2111 VTAIL.n210 VTAIL.n111 0.155672
R2112 VTAIL.n210 VTAIL.n209 0.155672
R2113 VTAIL.n209 VTAIL.n115 0.155672
R2114 VTAIL.n202 VTAIL.n115 0.155672
R2115 VTAIL.n202 VTAIL.n201 0.155672
R2116 VTAIL.n201 VTAIL.n119 0.155672
R2117 VTAIL.n194 VTAIL.n119 0.155672
R2118 VTAIL.n194 VTAIL.n193 0.155672
R2119 VTAIL.n193 VTAIL.n123 0.155672
R2120 VTAIL.n186 VTAIL.n123 0.155672
R2121 VTAIL.n186 VTAIL.n185 0.155672
R2122 VTAIL.n185 VTAIL.n129 0.155672
R2123 VTAIL.n178 VTAIL.n129 0.155672
R2124 VTAIL.n178 VTAIL.n177 0.155672
R2125 VTAIL.n177 VTAIL.n133 0.155672
R2126 VTAIL.n170 VTAIL.n133 0.155672
R2127 VTAIL.n170 VTAIL.n169 0.155672
R2128 VTAIL.n169 VTAIL.n137 0.155672
R2129 VTAIL.n162 VTAIL.n137 0.155672
R2130 VTAIL.n162 VTAIL.n161 0.155672
R2131 VTAIL.n161 VTAIL.n141 0.155672
R2132 VTAIL.n154 VTAIL.n141 0.155672
R2133 VTAIL.n154 VTAIL.n153 0.155672
R2134 VTAIL.n153 VTAIL.n145 0.155672
R2135 VDD1.n104 VDD1.n0 289.615
R2136 VDD1.n213 VDD1.n109 289.615
R2137 VDD1.n105 VDD1.n104 185
R2138 VDD1.n103 VDD1.n102 185
R2139 VDD1.n4 VDD1.n3 185
R2140 VDD1.n97 VDD1.n96 185
R2141 VDD1.n95 VDD1.n94 185
R2142 VDD1.n8 VDD1.n7 185
R2143 VDD1.n89 VDD1.n88 185
R2144 VDD1.n87 VDD1.n86 185
R2145 VDD1.n12 VDD1.n11 185
R2146 VDD1.n16 VDD1.n14 185
R2147 VDD1.n81 VDD1.n80 185
R2148 VDD1.n79 VDD1.n78 185
R2149 VDD1.n18 VDD1.n17 185
R2150 VDD1.n73 VDD1.n72 185
R2151 VDD1.n71 VDD1.n70 185
R2152 VDD1.n22 VDD1.n21 185
R2153 VDD1.n65 VDD1.n64 185
R2154 VDD1.n63 VDD1.n62 185
R2155 VDD1.n26 VDD1.n25 185
R2156 VDD1.n57 VDD1.n56 185
R2157 VDD1.n55 VDD1.n54 185
R2158 VDD1.n30 VDD1.n29 185
R2159 VDD1.n49 VDD1.n48 185
R2160 VDD1.n47 VDD1.n46 185
R2161 VDD1.n34 VDD1.n33 185
R2162 VDD1.n41 VDD1.n40 185
R2163 VDD1.n39 VDD1.n38 185
R2164 VDD1.n146 VDD1.n145 185
R2165 VDD1.n148 VDD1.n147 185
R2166 VDD1.n141 VDD1.n140 185
R2167 VDD1.n154 VDD1.n153 185
R2168 VDD1.n156 VDD1.n155 185
R2169 VDD1.n137 VDD1.n136 185
R2170 VDD1.n162 VDD1.n161 185
R2171 VDD1.n164 VDD1.n163 185
R2172 VDD1.n133 VDD1.n132 185
R2173 VDD1.n170 VDD1.n169 185
R2174 VDD1.n172 VDD1.n171 185
R2175 VDD1.n129 VDD1.n128 185
R2176 VDD1.n178 VDD1.n177 185
R2177 VDD1.n180 VDD1.n179 185
R2178 VDD1.n125 VDD1.n124 185
R2179 VDD1.n187 VDD1.n186 185
R2180 VDD1.n188 VDD1.n123 185
R2181 VDD1.n190 VDD1.n189 185
R2182 VDD1.n121 VDD1.n120 185
R2183 VDD1.n196 VDD1.n195 185
R2184 VDD1.n198 VDD1.n197 185
R2185 VDD1.n117 VDD1.n116 185
R2186 VDD1.n204 VDD1.n203 185
R2187 VDD1.n206 VDD1.n205 185
R2188 VDD1.n113 VDD1.n112 185
R2189 VDD1.n212 VDD1.n211 185
R2190 VDD1.n214 VDD1.n213 185
R2191 VDD1.n37 VDD1.t0 147.659
R2192 VDD1.n144 VDD1.t1 147.659
R2193 VDD1.n104 VDD1.n103 104.615
R2194 VDD1.n103 VDD1.n3 104.615
R2195 VDD1.n96 VDD1.n3 104.615
R2196 VDD1.n96 VDD1.n95 104.615
R2197 VDD1.n95 VDD1.n7 104.615
R2198 VDD1.n88 VDD1.n7 104.615
R2199 VDD1.n88 VDD1.n87 104.615
R2200 VDD1.n87 VDD1.n11 104.615
R2201 VDD1.n16 VDD1.n11 104.615
R2202 VDD1.n80 VDD1.n16 104.615
R2203 VDD1.n80 VDD1.n79 104.615
R2204 VDD1.n79 VDD1.n17 104.615
R2205 VDD1.n72 VDD1.n17 104.615
R2206 VDD1.n72 VDD1.n71 104.615
R2207 VDD1.n71 VDD1.n21 104.615
R2208 VDD1.n64 VDD1.n21 104.615
R2209 VDD1.n64 VDD1.n63 104.615
R2210 VDD1.n63 VDD1.n25 104.615
R2211 VDD1.n56 VDD1.n25 104.615
R2212 VDD1.n56 VDD1.n55 104.615
R2213 VDD1.n55 VDD1.n29 104.615
R2214 VDD1.n48 VDD1.n29 104.615
R2215 VDD1.n48 VDD1.n47 104.615
R2216 VDD1.n47 VDD1.n33 104.615
R2217 VDD1.n40 VDD1.n33 104.615
R2218 VDD1.n40 VDD1.n39 104.615
R2219 VDD1.n147 VDD1.n146 104.615
R2220 VDD1.n147 VDD1.n140 104.615
R2221 VDD1.n154 VDD1.n140 104.615
R2222 VDD1.n155 VDD1.n154 104.615
R2223 VDD1.n155 VDD1.n136 104.615
R2224 VDD1.n162 VDD1.n136 104.615
R2225 VDD1.n163 VDD1.n162 104.615
R2226 VDD1.n163 VDD1.n132 104.615
R2227 VDD1.n170 VDD1.n132 104.615
R2228 VDD1.n171 VDD1.n170 104.615
R2229 VDD1.n171 VDD1.n128 104.615
R2230 VDD1.n178 VDD1.n128 104.615
R2231 VDD1.n179 VDD1.n178 104.615
R2232 VDD1.n179 VDD1.n124 104.615
R2233 VDD1.n187 VDD1.n124 104.615
R2234 VDD1.n188 VDD1.n187 104.615
R2235 VDD1.n189 VDD1.n188 104.615
R2236 VDD1.n189 VDD1.n120 104.615
R2237 VDD1.n196 VDD1.n120 104.615
R2238 VDD1.n197 VDD1.n196 104.615
R2239 VDD1.n197 VDD1.n116 104.615
R2240 VDD1.n204 VDD1.n116 104.615
R2241 VDD1.n205 VDD1.n204 104.615
R2242 VDD1.n205 VDD1.n112 104.615
R2243 VDD1.n212 VDD1.n112 104.615
R2244 VDD1.n213 VDD1.n212 104.615
R2245 VDD1 VDD1.n217 92.4817
R2246 VDD1.n39 VDD1.t0 52.3082
R2247 VDD1.n146 VDD1.t1 52.3082
R2248 VDD1 VDD1.n108 48.5108
R2249 VDD1.n38 VDD1.n37 15.6677
R2250 VDD1.n145 VDD1.n144 15.6677
R2251 VDD1.n14 VDD1.n12 13.1884
R2252 VDD1.n190 VDD1.n121 13.1884
R2253 VDD1.n86 VDD1.n85 12.8005
R2254 VDD1.n82 VDD1.n81 12.8005
R2255 VDD1.n41 VDD1.n36 12.8005
R2256 VDD1.n148 VDD1.n143 12.8005
R2257 VDD1.n191 VDD1.n123 12.8005
R2258 VDD1.n195 VDD1.n194 12.8005
R2259 VDD1.n89 VDD1.n10 12.0247
R2260 VDD1.n78 VDD1.n15 12.0247
R2261 VDD1.n42 VDD1.n34 12.0247
R2262 VDD1.n149 VDD1.n141 12.0247
R2263 VDD1.n186 VDD1.n185 12.0247
R2264 VDD1.n198 VDD1.n119 12.0247
R2265 VDD1.n90 VDD1.n8 11.249
R2266 VDD1.n77 VDD1.n18 11.249
R2267 VDD1.n46 VDD1.n45 11.249
R2268 VDD1.n153 VDD1.n152 11.249
R2269 VDD1.n184 VDD1.n125 11.249
R2270 VDD1.n199 VDD1.n117 11.249
R2271 VDD1.n94 VDD1.n93 10.4732
R2272 VDD1.n74 VDD1.n73 10.4732
R2273 VDD1.n49 VDD1.n32 10.4732
R2274 VDD1.n156 VDD1.n139 10.4732
R2275 VDD1.n181 VDD1.n180 10.4732
R2276 VDD1.n203 VDD1.n202 10.4732
R2277 VDD1.n97 VDD1.n6 9.69747
R2278 VDD1.n70 VDD1.n20 9.69747
R2279 VDD1.n50 VDD1.n30 9.69747
R2280 VDD1.n157 VDD1.n137 9.69747
R2281 VDD1.n177 VDD1.n127 9.69747
R2282 VDD1.n206 VDD1.n115 9.69747
R2283 VDD1.n108 VDD1.n107 9.45567
R2284 VDD1.n217 VDD1.n216 9.45567
R2285 VDD1.n24 VDD1.n23 9.3005
R2286 VDD1.n67 VDD1.n66 9.3005
R2287 VDD1.n69 VDD1.n68 9.3005
R2288 VDD1.n20 VDD1.n19 9.3005
R2289 VDD1.n75 VDD1.n74 9.3005
R2290 VDD1.n77 VDD1.n76 9.3005
R2291 VDD1.n15 VDD1.n13 9.3005
R2292 VDD1.n83 VDD1.n82 9.3005
R2293 VDD1.n107 VDD1.n106 9.3005
R2294 VDD1.n2 VDD1.n1 9.3005
R2295 VDD1.n101 VDD1.n100 9.3005
R2296 VDD1.n99 VDD1.n98 9.3005
R2297 VDD1.n6 VDD1.n5 9.3005
R2298 VDD1.n93 VDD1.n92 9.3005
R2299 VDD1.n91 VDD1.n90 9.3005
R2300 VDD1.n10 VDD1.n9 9.3005
R2301 VDD1.n85 VDD1.n84 9.3005
R2302 VDD1.n61 VDD1.n60 9.3005
R2303 VDD1.n59 VDD1.n58 9.3005
R2304 VDD1.n28 VDD1.n27 9.3005
R2305 VDD1.n53 VDD1.n52 9.3005
R2306 VDD1.n51 VDD1.n50 9.3005
R2307 VDD1.n32 VDD1.n31 9.3005
R2308 VDD1.n45 VDD1.n44 9.3005
R2309 VDD1.n43 VDD1.n42 9.3005
R2310 VDD1.n36 VDD1.n35 9.3005
R2311 VDD1.n216 VDD1.n215 9.3005
R2312 VDD1.n210 VDD1.n209 9.3005
R2313 VDD1.n208 VDD1.n207 9.3005
R2314 VDD1.n115 VDD1.n114 9.3005
R2315 VDD1.n202 VDD1.n201 9.3005
R2316 VDD1.n200 VDD1.n199 9.3005
R2317 VDD1.n119 VDD1.n118 9.3005
R2318 VDD1.n194 VDD1.n193 9.3005
R2319 VDD1.n166 VDD1.n165 9.3005
R2320 VDD1.n135 VDD1.n134 9.3005
R2321 VDD1.n160 VDD1.n159 9.3005
R2322 VDD1.n158 VDD1.n157 9.3005
R2323 VDD1.n139 VDD1.n138 9.3005
R2324 VDD1.n152 VDD1.n151 9.3005
R2325 VDD1.n150 VDD1.n149 9.3005
R2326 VDD1.n143 VDD1.n142 9.3005
R2327 VDD1.n168 VDD1.n167 9.3005
R2328 VDD1.n131 VDD1.n130 9.3005
R2329 VDD1.n174 VDD1.n173 9.3005
R2330 VDD1.n176 VDD1.n175 9.3005
R2331 VDD1.n127 VDD1.n126 9.3005
R2332 VDD1.n182 VDD1.n181 9.3005
R2333 VDD1.n184 VDD1.n183 9.3005
R2334 VDD1.n185 VDD1.n122 9.3005
R2335 VDD1.n192 VDD1.n191 9.3005
R2336 VDD1.n111 VDD1.n110 9.3005
R2337 VDD1.n98 VDD1.n4 8.92171
R2338 VDD1.n69 VDD1.n22 8.92171
R2339 VDD1.n54 VDD1.n53 8.92171
R2340 VDD1.n161 VDD1.n160 8.92171
R2341 VDD1.n176 VDD1.n129 8.92171
R2342 VDD1.n207 VDD1.n113 8.92171
R2343 VDD1.n102 VDD1.n101 8.14595
R2344 VDD1.n66 VDD1.n65 8.14595
R2345 VDD1.n57 VDD1.n28 8.14595
R2346 VDD1.n164 VDD1.n135 8.14595
R2347 VDD1.n173 VDD1.n172 8.14595
R2348 VDD1.n211 VDD1.n210 8.14595
R2349 VDD1.n108 VDD1.n0 7.3702
R2350 VDD1.n105 VDD1.n2 7.3702
R2351 VDD1.n62 VDD1.n24 7.3702
R2352 VDD1.n58 VDD1.n26 7.3702
R2353 VDD1.n165 VDD1.n133 7.3702
R2354 VDD1.n169 VDD1.n131 7.3702
R2355 VDD1.n214 VDD1.n111 7.3702
R2356 VDD1.n217 VDD1.n109 7.3702
R2357 VDD1.n106 VDD1.n0 6.59444
R2358 VDD1.n106 VDD1.n105 6.59444
R2359 VDD1.n62 VDD1.n61 6.59444
R2360 VDD1.n61 VDD1.n26 6.59444
R2361 VDD1.n168 VDD1.n133 6.59444
R2362 VDD1.n169 VDD1.n168 6.59444
R2363 VDD1.n215 VDD1.n214 6.59444
R2364 VDD1.n215 VDD1.n109 6.59444
R2365 VDD1.n102 VDD1.n2 5.81868
R2366 VDD1.n65 VDD1.n24 5.81868
R2367 VDD1.n58 VDD1.n57 5.81868
R2368 VDD1.n165 VDD1.n164 5.81868
R2369 VDD1.n172 VDD1.n131 5.81868
R2370 VDD1.n211 VDD1.n111 5.81868
R2371 VDD1.n101 VDD1.n4 5.04292
R2372 VDD1.n66 VDD1.n22 5.04292
R2373 VDD1.n54 VDD1.n28 5.04292
R2374 VDD1.n161 VDD1.n135 5.04292
R2375 VDD1.n173 VDD1.n129 5.04292
R2376 VDD1.n210 VDD1.n113 5.04292
R2377 VDD1.n37 VDD1.n35 4.38563
R2378 VDD1.n144 VDD1.n142 4.38563
R2379 VDD1.n98 VDD1.n97 4.26717
R2380 VDD1.n70 VDD1.n69 4.26717
R2381 VDD1.n53 VDD1.n30 4.26717
R2382 VDD1.n160 VDD1.n137 4.26717
R2383 VDD1.n177 VDD1.n176 4.26717
R2384 VDD1.n207 VDD1.n206 4.26717
R2385 VDD1.n94 VDD1.n6 3.49141
R2386 VDD1.n73 VDD1.n20 3.49141
R2387 VDD1.n50 VDD1.n49 3.49141
R2388 VDD1.n157 VDD1.n156 3.49141
R2389 VDD1.n180 VDD1.n127 3.49141
R2390 VDD1.n203 VDD1.n115 3.49141
R2391 VDD1.n93 VDD1.n8 2.71565
R2392 VDD1.n74 VDD1.n18 2.71565
R2393 VDD1.n46 VDD1.n32 2.71565
R2394 VDD1.n153 VDD1.n139 2.71565
R2395 VDD1.n181 VDD1.n125 2.71565
R2396 VDD1.n202 VDD1.n117 2.71565
R2397 VDD1.n90 VDD1.n89 1.93989
R2398 VDD1.n78 VDD1.n77 1.93989
R2399 VDD1.n45 VDD1.n34 1.93989
R2400 VDD1.n152 VDD1.n141 1.93989
R2401 VDD1.n186 VDD1.n184 1.93989
R2402 VDD1.n199 VDD1.n198 1.93989
R2403 VDD1.n86 VDD1.n10 1.16414
R2404 VDD1.n81 VDD1.n15 1.16414
R2405 VDD1.n42 VDD1.n41 1.16414
R2406 VDD1.n149 VDD1.n148 1.16414
R2407 VDD1.n185 VDD1.n123 1.16414
R2408 VDD1.n195 VDD1.n119 1.16414
R2409 VDD1.n85 VDD1.n12 0.388379
R2410 VDD1.n82 VDD1.n14 0.388379
R2411 VDD1.n38 VDD1.n36 0.388379
R2412 VDD1.n145 VDD1.n143 0.388379
R2413 VDD1.n191 VDD1.n190 0.388379
R2414 VDD1.n194 VDD1.n121 0.388379
R2415 VDD1.n107 VDD1.n1 0.155672
R2416 VDD1.n100 VDD1.n1 0.155672
R2417 VDD1.n100 VDD1.n99 0.155672
R2418 VDD1.n99 VDD1.n5 0.155672
R2419 VDD1.n92 VDD1.n5 0.155672
R2420 VDD1.n92 VDD1.n91 0.155672
R2421 VDD1.n91 VDD1.n9 0.155672
R2422 VDD1.n84 VDD1.n9 0.155672
R2423 VDD1.n84 VDD1.n83 0.155672
R2424 VDD1.n83 VDD1.n13 0.155672
R2425 VDD1.n76 VDD1.n13 0.155672
R2426 VDD1.n76 VDD1.n75 0.155672
R2427 VDD1.n75 VDD1.n19 0.155672
R2428 VDD1.n68 VDD1.n19 0.155672
R2429 VDD1.n68 VDD1.n67 0.155672
R2430 VDD1.n67 VDD1.n23 0.155672
R2431 VDD1.n60 VDD1.n23 0.155672
R2432 VDD1.n60 VDD1.n59 0.155672
R2433 VDD1.n59 VDD1.n27 0.155672
R2434 VDD1.n52 VDD1.n27 0.155672
R2435 VDD1.n52 VDD1.n51 0.155672
R2436 VDD1.n51 VDD1.n31 0.155672
R2437 VDD1.n44 VDD1.n31 0.155672
R2438 VDD1.n44 VDD1.n43 0.155672
R2439 VDD1.n43 VDD1.n35 0.155672
R2440 VDD1.n150 VDD1.n142 0.155672
R2441 VDD1.n151 VDD1.n150 0.155672
R2442 VDD1.n151 VDD1.n138 0.155672
R2443 VDD1.n158 VDD1.n138 0.155672
R2444 VDD1.n159 VDD1.n158 0.155672
R2445 VDD1.n159 VDD1.n134 0.155672
R2446 VDD1.n166 VDD1.n134 0.155672
R2447 VDD1.n167 VDD1.n166 0.155672
R2448 VDD1.n167 VDD1.n130 0.155672
R2449 VDD1.n174 VDD1.n130 0.155672
R2450 VDD1.n175 VDD1.n174 0.155672
R2451 VDD1.n175 VDD1.n126 0.155672
R2452 VDD1.n182 VDD1.n126 0.155672
R2453 VDD1.n183 VDD1.n182 0.155672
R2454 VDD1.n183 VDD1.n122 0.155672
R2455 VDD1.n192 VDD1.n122 0.155672
R2456 VDD1.n193 VDD1.n192 0.155672
R2457 VDD1.n193 VDD1.n118 0.155672
R2458 VDD1.n200 VDD1.n118 0.155672
R2459 VDD1.n201 VDD1.n200 0.155672
R2460 VDD1.n201 VDD1.n114 0.155672
R2461 VDD1.n208 VDD1.n114 0.155672
R2462 VDD1.n209 VDD1.n208 0.155672
R2463 VDD1.n209 VDD1.n110 0.155672
R2464 VDD1.n216 VDD1.n110 0.155672
R2465 VN VN.t0 504.962
R2466 VN VN.t1 457.666
R2467 VDD2.n213 VDD2.n109 289.615
R2468 VDD2.n104 VDD2.n0 289.615
R2469 VDD2.n214 VDD2.n213 185
R2470 VDD2.n212 VDD2.n211 185
R2471 VDD2.n113 VDD2.n112 185
R2472 VDD2.n206 VDD2.n205 185
R2473 VDD2.n204 VDD2.n203 185
R2474 VDD2.n117 VDD2.n116 185
R2475 VDD2.n198 VDD2.n197 185
R2476 VDD2.n196 VDD2.n195 185
R2477 VDD2.n121 VDD2.n120 185
R2478 VDD2.n125 VDD2.n123 185
R2479 VDD2.n190 VDD2.n189 185
R2480 VDD2.n188 VDD2.n187 185
R2481 VDD2.n127 VDD2.n126 185
R2482 VDD2.n182 VDD2.n181 185
R2483 VDD2.n180 VDD2.n179 185
R2484 VDD2.n131 VDD2.n130 185
R2485 VDD2.n174 VDD2.n173 185
R2486 VDD2.n172 VDD2.n171 185
R2487 VDD2.n135 VDD2.n134 185
R2488 VDD2.n166 VDD2.n165 185
R2489 VDD2.n164 VDD2.n163 185
R2490 VDD2.n139 VDD2.n138 185
R2491 VDD2.n158 VDD2.n157 185
R2492 VDD2.n156 VDD2.n155 185
R2493 VDD2.n143 VDD2.n142 185
R2494 VDD2.n150 VDD2.n149 185
R2495 VDD2.n148 VDD2.n147 185
R2496 VDD2.n37 VDD2.n36 185
R2497 VDD2.n39 VDD2.n38 185
R2498 VDD2.n32 VDD2.n31 185
R2499 VDD2.n45 VDD2.n44 185
R2500 VDD2.n47 VDD2.n46 185
R2501 VDD2.n28 VDD2.n27 185
R2502 VDD2.n53 VDD2.n52 185
R2503 VDD2.n55 VDD2.n54 185
R2504 VDD2.n24 VDD2.n23 185
R2505 VDD2.n61 VDD2.n60 185
R2506 VDD2.n63 VDD2.n62 185
R2507 VDD2.n20 VDD2.n19 185
R2508 VDD2.n69 VDD2.n68 185
R2509 VDD2.n71 VDD2.n70 185
R2510 VDD2.n16 VDD2.n15 185
R2511 VDD2.n78 VDD2.n77 185
R2512 VDD2.n79 VDD2.n14 185
R2513 VDD2.n81 VDD2.n80 185
R2514 VDD2.n12 VDD2.n11 185
R2515 VDD2.n87 VDD2.n86 185
R2516 VDD2.n89 VDD2.n88 185
R2517 VDD2.n8 VDD2.n7 185
R2518 VDD2.n95 VDD2.n94 185
R2519 VDD2.n97 VDD2.n96 185
R2520 VDD2.n4 VDD2.n3 185
R2521 VDD2.n103 VDD2.n102 185
R2522 VDD2.n105 VDD2.n104 185
R2523 VDD2.n146 VDD2.t1 147.659
R2524 VDD2.n35 VDD2.t0 147.659
R2525 VDD2.n213 VDD2.n212 104.615
R2526 VDD2.n212 VDD2.n112 104.615
R2527 VDD2.n205 VDD2.n112 104.615
R2528 VDD2.n205 VDD2.n204 104.615
R2529 VDD2.n204 VDD2.n116 104.615
R2530 VDD2.n197 VDD2.n116 104.615
R2531 VDD2.n197 VDD2.n196 104.615
R2532 VDD2.n196 VDD2.n120 104.615
R2533 VDD2.n125 VDD2.n120 104.615
R2534 VDD2.n189 VDD2.n125 104.615
R2535 VDD2.n189 VDD2.n188 104.615
R2536 VDD2.n188 VDD2.n126 104.615
R2537 VDD2.n181 VDD2.n126 104.615
R2538 VDD2.n181 VDD2.n180 104.615
R2539 VDD2.n180 VDD2.n130 104.615
R2540 VDD2.n173 VDD2.n130 104.615
R2541 VDD2.n173 VDD2.n172 104.615
R2542 VDD2.n172 VDD2.n134 104.615
R2543 VDD2.n165 VDD2.n134 104.615
R2544 VDD2.n165 VDD2.n164 104.615
R2545 VDD2.n164 VDD2.n138 104.615
R2546 VDD2.n157 VDD2.n138 104.615
R2547 VDD2.n157 VDD2.n156 104.615
R2548 VDD2.n156 VDD2.n142 104.615
R2549 VDD2.n149 VDD2.n142 104.615
R2550 VDD2.n149 VDD2.n148 104.615
R2551 VDD2.n38 VDD2.n37 104.615
R2552 VDD2.n38 VDD2.n31 104.615
R2553 VDD2.n45 VDD2.n31 104.615
R2554 VDD2.n46 VDD2.n45 104.615
R2555 VDD2.n46 VDD2.n27 104.615
R2556 VDD2.n53 VDD2.n27 104.615
R2557 VDD2.n54 VDD2.n53 104.615
R2558 VDD2.n54 VDD2.n23 104.615
R2559 VDD2.n61 VDD2.n23 104.615
R2560 VDD2.n62 VDD2.n61 104.615
R2561 VDD2.n62 VDD2.n19 104.615
R2562 VDD2.n69 VDD2.n19 104.615
R2563 VDD2.n70 VDD2.n69 104.615
R2564 VDD2.n70 VDD2.n15 104.615
R2565 VDD2.n78 VDD2.n15 104.615
R2566 VDD2.n79 VDD2.n78 104.615
R2567 VDD2.n80 VDD2.n79 104.615
R2568 VDD2.n80 VDD2.n11 104.615
R2569 VDD2.n87 VDD2.n11 104.615
R2570 VDD2.n88 VDD2.n87 104.615
R2571 VDD2.n88 VDD2.n7 104.615
R2572 VDD2.n95 VDD2.n7 104.615
R2573 VDD2.n96 VDD2.n95 104.615
R2574 VDD2.n96 VDD2.n3 104.615
R2575 VDD2.n103 VDD2.n3 104.615
R2576 VDD2.n104 VDD2.n103 104.615
R2577 VDD2.n218 VDD2.n108 91.5927
R2578 VDD2.n148 VDD2.t1 52.3082
R2579 VDD2.n37 VDD2.t0 52.3082
R2580 VDD2.n218 VDD2.n217 48.0884
R2581 VDD2.n147 VDD2.n146 15.6677
R2582 VDD2.n36 VDD2.n35 15.6677
R2583 VDD2.n123 VDD2.n121 13.1884
R2584 VDD2.n81 VDD2.n12 13.1884
R2585 VDD2.n195 VDD2.n194 12.8005
R2586 VDD2.n191 VDD2.n190 12.8005
R2587 VDD2.n150 VDD2.n145 12.8005
R2588 VDD2.n39 VDD2.n34 12.8005
R2589 VDD2.n82 VDD2.n14 12.8005
R2590 VDD2.n86 VDD2.n85 12.8005
R2591 VDD2.n198 VDD2.n119 12.0247
R2592 VDD2.n187 VDD2.n124 12.0247
R2593 VDD2.n151 VDD2.n143 12.0247
R2594 VDD2.n40 VDD2.n32 12.0247
R2595 VDD2.n77 VDD2.n76 12.0247
R2596 VDD2.n89 VDD2.n10 12.0247
R2597 VDD2.n199 VDD2.n117 11.249
R2598 VDD2.n186 VDD2.n127 11.249
R2599 VDD2.n155 VDD2.n154 11.249
R2600 VDD2.n44 VDD2.n43 11.249
R2601 VDD2.n75 VDD2.n16 11.249
R2602 VDD2.n90 VDD2.n8 11.249
R2603 VDD2.n203 VDD2.n202 10.4732
R2604 VDD2.n183 VDD2.n182 10.4732
R2605 VDD2.n158 VDD2.n141 10.4732
R2606 VDD2.n47 VDD2.n30 10.4732
R2607 VDD2.n72 VDD2.n71 10.4732
R2608 VDD2.n94 VDD2.n93 10.4732
R2609 VDD2.n206 VDD2.n115 9.69747
R2610 VDD2.n179 VDD2.n129 9.69747
R2611 VDD2.n159 VDD2.n139 9.69747
R2612 VDD2.n48 VDD2.n28 9.69747
R2613 VDD2.n68 VDD2.n18 9.69747
R2614 VDD2.n97 VDD2.n6 9.69747
R2615 VDD2.n217 VDD2.n216 9.45567
R2616 VDD2.n108 VDD2.n107 9.45567
R2617 VDD2.n133 VDD2.n132 9.3005
R2618 VDD2.n176 VDD2.n175 9.3005
R2619 VDD2.n178 VDD2.n177 9.3005
R2620 VDD2.n129 VDD2.n128 9.3005
R2621 VDD2.n184 VDD2.n183 9.3005
R2622 VDD2.n186 VDD2.n185 9.3005
R2623 VDD2.n124 VDD2.n122 9.3005
R2624 VDD2.n192 VDD2.n191 9.3005
R2625 VDD2.n216 VDD2.n215 9.3005
R2626 VDD2.n111 VDD2.n110 9.3005
R2627 VDD2.n210 VDD2.n209 9.3005
R2628 VDD2.n208 VDD2.n207 9.3005
R2629 VDD2.n115 VDD2.n114 9.3005
R2630 VDD2.n202 VDD2.n201 9.3005
R2631 VDD2.n200 VDD2.n199 9.3005
R2632 VDD2.n119 VDD2.n118 9.3005
R2633 VDD2.n194 VDD2.n193 9.3005
R2634 VDD2.n170 VDD2.n169 9.3005
R2635 VDD2.n168 VDD2.n167 9.3005
R2636 VDD2.n137 VDD2.n136 9.3005
R2637 VDD2.n162 VDD2.n161 9.3005
R2638 VDD2.n160 VDD2.n159 9.3005
R2639 VDD2.n141 VDD2.n140 9.3005
R2640 VDD2.n154 VDD2.n153 9.3005
R2641 VDD2.n152 VDD2.n151 9.3005
R2642 VDD2.n145 VDD2.n144 9.3005
R2643 VDD2.n107 VDD2.n106 9.3005
R2644 VDD2.n101 VDD2.n100 9.3005
R2645 VDD2.n99 VDD2.n98 9.3005
R2646 VDD2.n6 VDD2.n5 9.3005
R2647 VDD2.n93 VDD2.n92 9.3005
R2648 VDD2.n91 VDD2.n90 9.3005
R2649 VDD2.n10 VDD2.n9 9.3005
R2650 VDD2.n85 VDD2.n84 9.3005
R2651 VDD2.n57 VDD2.n56 9.3005
R2652 VDD2.n26 VDD2.n25 9.3005
R2653 VDD2.n51 VDD2.n50 9.3005
R2654 VDD2.n49 VDD2.n48 9.3005
R2655 VDD2.n30 VDD2.n29 9.3005
R2656 VDD2.n43 VDD2.n42 9.3005
R2657 VDD2.n41 VDD2.n40 9.3005
R2658 VDD2.n34 VDD2.n33 9.3005
R2659 VDD2.n59 VDD2.n58 9.3005
R2660 VDD2.n22 VDD2.n21 9.3005
R2661 VDD2.n65 VDD2.n64 9.3005
R2662 VDD2.n67 VDD2.n66 9.3005
R2663 VDD2.n18 VDD2.n17 9.3005
R2664 VDD2.n73 VDD2.n72 9.3005
R2665 VDD2.n75 VDD2.n74 9.3005
R2666 VDD2.n76 VDD2.n13 9.3005
R2667 VDD2.n83 VDD2.n82 9.3005
R2668 VDD2.n2 VDD2.n1 9.3005
R2669 VDD2.n207 VDD2.n113 8.92171
R2670 VDD2.n178 VDD2.n131 8.92171
R2671 VDD2.n163 VDD2.n162 8.92171
R2672 VDD2.n52 VDD2.n51 8.92171
R2673 VDD2.n67 VDD2.n20 8.92171
R2674 VDD2.n98 VDD2.n4 8.92171
R2675 VDD2.n211 VDD2.n210 8.14595
R2676 VDD2.n175 VDD2.n174 8.14595
R2677 VDD2.n166 VDD2.n137 8.14595
R2678 VDD2.n55 VDD2.n26 8.14595
R2679 VDD2.n64 VDD2.n63 8.14595
R2680 VDD2.n102 VDD2.n101 8.14595
R2681 VDD2.n217 VDD2.n109 7.3702
R2682 VDD2.n214 VDD2.n111 7.3702
R2683 VDD2.n171 VDD2.n133 7.3702
R2684 VDD2.n167 VDD2.n135 7.3702
R2685 VDD2.n56 VDD2.n24 7.3702
R2686 VDD2.n60 VDD2.n22 7.3702
R2687 VDD2.n105 VDD2.n2 7.3702
R2688 VDD2.n108 VDD2.n0 7.3702
R2689 VDD2.n215 VDD2.n109 6.59444
R2690 VDD2.n215 VDD2.n214 6.59444
R2691 VDD2.n171 VDD2.n170 6.59444
R2692 VDD2.n170 VDD2.n135 6.59444
R2693 VDD2.n59 VDD2.n24 6.59444
R2694 VDD2.n60 VDD2.n59 6.59444
R2695 VDD2.n106 VDD2.n105 6.59444
R2696 VDD2.n106 VDD2.n0 6.59444
R2697 VDD2.n211 VDD2.n111 5.81868
R2698 VDD2.n174 VDD2.n133 5.81868
R2699 VDD2.n167 VDD2.n166 5.81868
R2700 VDD2.n56 VDD2.n55 5.81868
R2701 VDD2.n63 VDD2.n22 5.81868
R2702 VDD2.n102 VDD2.n2 5.81868
R2703 VDD2.n210 VDD2.n113 5.04292
R2704 VDD2.n175 VDD2.n131 5.04292
R2705 VDD2.n163 VDD2.n137 5.04292
R2706 VDD2.n52 VDD2.n26 5.04292
R2707 VDD2.n64 VDD2.n20 5.04292
R2708 VDD2.n101 VDD2.n4 5.04292
R2709 VDD2.n146 VDD2.n144 4.38563
R2710 VDD2.n35 VDD2.n33 4.38563
R2711 VDD2.n207 VDD2.n206 4.26717
R2712 VDD2.n179 VDD2.n178 4.26717
R2713 VDD2.n162 VDD2.n139 4.26717
R2714 VDD2.n51 VDD2.n28 4.26717
R2715 VDD2.n68 VDD2.n67 4.26717
R2716 VDD2.n98 VDD2.n97 4.26717
R2717 VDD2.n203 VDD2.n115 3.49141
R2718 VDD2.n182 VDD2.n129 3.49141
R2719 VDD2.n159 VDD2.n158 3.49141
R2720 VDD2.n48 VDD2.n47 3.49141
R2721 VDD2.n71 VDD2.n18 3.49141
R2722 VDD2.n94 VDD2.n6 3.49141
R2723 VDD2.n202 VDD2.n117 2.71565
R2724 VDD2.n183 VDD2.n127 2.71565
R2725 VDD2.n155 VDD2.n141 2.71565
R2726 VDD2.n44 VDD2.n30 2.71565
R2727 VDD2.n72 VDD2.n16 2.71565
R2728 VDD2.n93 VDD2.n8 2.71565
R2729 VDD2.n199 VDD2.n198 1.93989
R2730 VDD2.n187 VDD2.n186 1.93989
R2731 VDD2.n154 VDD2.n143 1.93989
R2732 VDD2.n43 VDD2.n32 1.93989
R2733 VDD2.n77 VDD2.n75 1.93989
R2734 VDD2.n90 VDD2.n89 1.93989
R2735 VDD2.n195 VDD2.n119 1.16414
R2736 VDD2.n190 VDD2.n124 1.16414
R2737 VDD2.n151 VDD2.n150 1.16414
R2738 VDD2.n40 VDD2.n39 1.16414
R2739 VDD2.n76 VDD2.n14 1.16414
R2740 VDD2.n86 VDD2.n10 1.16414
R2741 VDD2 VDD2.n218 0.422914
R2742 VDD2.n194 VDD2.n121 0.388379
R2743 VDD2.n191 VDD2.n123 0.388379
R2744 VDD2.n147 VDD2.n145 0.388379
R2745 VDD2.n36 VDD2.n34 0.388379
R2746 VDD2.n82 VDD2.n81 0.388379
R2747 VDD2.n85 VDD2.n12 0.388379
R2748 VDD2.n216 VDD2.n110 0.155672
R2749 VDD2.n209 VDD2.n110 0.155672
R2750 VDD2.n209 VDD2.n208 0.155672
R2751 VDD2.n208 VDD2.n114 0.155672
R2752 VDD2.n201 VDD2.n114 0.155672
R2753 VDD2.n201 VDD2.n200 0.155672
R2754 VDD2.n200 VDD2.n118 0.155672
R2755 VDD2.n193 VDD2.n118 0.155672
R2756 VDD2.n193 VDD2.n192 0.155672
R2757 VDD2.n192 VDD2.n122 0.155672
R2758 VDD2.n185 VDD2.n122 0.155672
R2759 VDD2.n185 VDD2.n184 0.155672
R2760 VDD2.n184 VDD2.n128 0.155672
R2761 VDD2.n177 VDD2.n128 0.155672
R2762 VDD2.n177 VDD2.n176 0.155672
R2763 VDD2.n176 VDD2.n132 0.155672
R2764 VDD2.n169 VDD2.n132 0.155672
R2765 VDD2.n169 VDD2.n168 0.155672
R2766 VDD2.n168 VDD2.n136 0.155672
R2767 VDD2.n161 VDD2.n136 0.155672
R2768 VDD2.n161 VDD2.n160 0.155672
R2769 VDD2.n160 VDD2.n140 0.155672
R2770 VDD2.n153 VDD2.n140 0.155672
R2771 VDD2.n153 VDD2.n152 0.155672
R2772 VDD2.n152 VDD2.n144 0.155672
R2773 VDD2.n41 VDD2.n33 0.155672
R2774 VDD2.n42 VDD2.n41 0.155672
R2775 VDD2.n42 VDD2.n29 0.155672
R2776 VDD2.n49 VDD2.n29 0.155672
R2777 VDD2.n50 VDD2.n49 0.155672
R2778 VDD2.n50 VDD2.n25 0.155672
R2779 VDD2.n57 VDD2.n25 0.155672
R2780 VDD2.n58 VDD2.n57 0.155672
R2781 VDD2.n58 VDD2.n21 0.155672
R2782 VDD2.n65 VDD2.n21 0.155672
R2783 VDD2.n66 VDD2.n65 0.155672
R2784 VDD2.n66 VDD2.n17 0.155672
R2785 VDD2.n73 VDD2.n17 0.155672
R2786 VDD2.n74 VDD2.n73 0.155672
R2787 VDD2.n74 VDD2.n13 0.155672
R2788 VDD2.n83 VDD2.n13 0.155672
R2789 VDD2.n84 VDD2.n83 0.155672
R2790 VDD2.n84 VDD2.n9 0.155672
R2791 VDD2.n91 VDD2.n9 0.155672
R2792 VDD2.n92 VDD2.n91 0.155672
R2793 VDD2.n92 VDD2.n5 0.155672
R2794 VDD2.n99 VDD2.n5 0.155672
R2795 VDD2.n100 VDD2.n99 0.155672
R2796 VDD2.n100 VDD2.n1 0.155672
R2797 VDD2.n107 VDD2.n1 0.155672
C0 VN VP 6.28586f
C1 VN VTAIL 3.09441f
C2 VDD1 VN 0.147888f
C3 VTAIL VP 3.10907f
C4 VDD2 VN 3.83843f
C5 VDD1 VP 3.96743f
C6 VDD1 VTAIL 7.42804f
C7 VDD2 VP 0.282384f
C8 VDD2 VTAIL 7.46534f
C9 VDD1 VDD2 0.532165f
C10 VDD2 B 5.368645f
C11 VDD1 B 8.43401f
C12 VTAIL B 9.66584f
C13 VN B 11.48697f
C14 VP B 5.368913f
C15 VDD2.n0 B 0.028672f
C16 VDD2.n1 B 0.020014f
C17 VDD2.n2 B 0.010755f
C18 VDD2.n3 B 0.02542f
C19 VDD2.n4 B 0.011387f
C20 VDD2.n5 B 0.020014f
C21 VDD2.n6 B 0.010755f
C22 VDD2.n7 B 0.02542f
C23 VDD2.n8 B 0.011387f
C24 VDD2.n9 B 0.020014f
C25 VDD2.n10 B 0.010755f
C26 VDD2.n11 B 0.02542f
C27 VDD2.n12 B 0.011071f
C28 VDD2.n13 B 0.020014f
C29 VDD2.n14 B 0.011387f
C30 VDD2.n15 B 0.02542f
C31 VDD2.n16 B 0.011387f
C32 VDD2.n17 B 0.020014f
C33 VDD2.n18 B 0.010755f
C34 VDD2.n19 B 0.02542f
C35 VDD2.n20 B 0.011387f
C36 VDD2.n21 B 0.020014f
C37 VDD2.n22 B 0.010755f
C38 VDD2.n23 B 0.02542f
C39 VDD2.n24 B 0.011387f
C40 VDD2.n25 B 0.020014f
C41 VDD2.n26 B 0.010755f
C42 VDD2.n27 B 0.02542f
C43 VDD2.n28 B 0.011387f
C44 VDD2.n29 B 0.020014f
C45 VDD2.n30 B 0.010755f
C46 VDD2.n31 B 0.02542f
C47 VDD2.n32 B 0.011387f
C48 VDD2.n33 B 1.72775f
C49 VDD2.n34 B 0.010755f
C50 VDD2.t0 B 0.042234f
C51 VDD2.n35 B 0.15382f
C52 VDD2.n36 B 0.015017f
C53 VDD2.n37 B 0.019065f
C54 VDD2.n38 B 0.02542f
C55 VDD2.n39 B 0.011387f
C56 VDD2.n40 B 0.010755f
C57 VDD2.n41 B 0.020014f
C58 VDD2.n42 B 0.020014f
C59 VDD2.n43 B 0.010755f
C60 VDD2.n44 B 0.011387f
C61 VDD2.n45 B 0.02542f
C62 VDD2.n46 B 0.02542f
C63 VDD2.n47 B 0.011387f
C64 VDD2.n48 B 0.010755f
C65 VDD2.n49 B 0.020014f
C66 VDD2.n50 B 0.020014f
C67 VDD2.n51 B 0.010755f
C68 VDD2.n52 B 0.011387f
C69 VDD2.n53 B 0.02542f
C70 VDD2.n54 B 0.02542f
C71 VDD2.n55 B 0.011387f
C72 VDD2.n56 B 0.010755f
C73 VDD2.n57 B 0.020014f
C74 VDD2.n58 B 0.020014f
C75 VDD2.n59 B 0.010755f
C76 VDD2.n60 B 0.011387f
C77 VDD2.n61 B 0.02542f
C78 VDD2.n62 B 0.02542f
C79 VDD2.n63 B 0.011387f
C80 VDD2.n64 B 0.010755f
C81 VDD2.n65 B 0.020014f
C82 VDD2.n66 B 0.020014f
C83 VDD2.n67 B 0.010755f
C84 VDD2.n68 B 0.011387f
C85 VDD2.n69 B 0.02542f
C86 VDD2.n70 B 0.02542f
C87 VDD2.n71 B 0.011387f
C88 VDD2.n72 B 0.010755f
C89 VDD2.n73 B 0.020014f
C90 VDD2.n74 B 0.020014f
C91 VDD2.n75 B 0.010755f
C92 VDD2.n76 B 0.010755f
C93 VDD2.n77 B 0.011387f
C94 VDD2.n78 B 0.02542f
C95 VDD2.n79 B 0.02542f
C96 VDD2.n80 B 0.02542f
C97 VDD2.n81 B 0.011071f
C98 VDD2.n82 B 0.010755f
C99 VDD2.n83 B 0.020014f
C100 VDD2.n84 B 0.020014f
C101 VDD2.n85 B 0.010755f
C102 VDD2.n86 B 0.011387f
C103 VDD2.n87 B 0.02542f
C104 VDD2.n88 B 0.02542f
C105 VDD2.n89 B 0.011387f
C106 VDD2.n90 B 0.010755f
C107 VDD2.n91 B 0.020014f
C108 VDD2.n92 B 0.020014f
C109 VDD2.n93 B 0.010755f
C110 VDD2.n94 B 0.011387f
C111 VDD2.n95 B 0.02542f
C112 VDD2.n96 B 0.02542f
C113 VDD2.n97 B 0.011387f
C114 VDD2.n98 B 0.010755f
C115 VDD2.n99 B 0.020014f
C116 VDD2.n100 B 0.020014f
C117 VDD2.n101 B 0.010755f
C118 VDD2.n102 B 0.011387f
C119 VDD2.n103 B 0.02542f
C120 VDD2.n104 B 0.055986f
C121 VDD2.n105 B 0.011387f
C122 VDD2.n106 B 0.010755f
C123 VDD2.n107 B 0.045168f
C124 VDD2.n108 B 0.754761f
C125 VDD2.n109 B 0.028672f
C126 VDD2.n110 B 0.020014f
C127 VDD2.n111 B 0.010755f
C128 VDD2.n112 B 0.02542f
C129 VDD2.n113 B 0.011387f
C130 VDD2.n114 B 0.020014f
C131 VDD2.n115 B 0.010755f
C132 VDD2.n116 B 0.02542f
C133 VDD2.n117 B 0.011387f
C134 VDD2.n118 B 0.020014f
C135 VDD2.n119 B 0.010755f
C136 VDD2.n120 B 0.02542f
C137 VDD2.n121 B 0.011071f
C138 VDD2.n122 B 0.020014f
C139 VDD2.n123 B 0.011071f
C140 VDD2.n124 B 0.010755f
C141 VDD2.n125 B 0.02542f
C142 VDD2.n126 B 0.02542f
C143 VDD2.n127 B 0.011387f
C144 VDD2.n128 B 0.020014f
C145 VDD2.n129 B 0.010755f
C146 VDD2.n130 B 0.02542f
C147 VDD2.n131 B 0.011387f
C148 VDD2.n132 B 0.020014f
C149 VDD2.n133 B 0.010755f
C150 VDD2.n134 B 0.02542f
C151 VDD2.n135 B 0.011387f
C152 VDD2.n136 B 0.020014f
C153 VDD2.n137 B 0.010755f
C154 VDD2.n138 B 0.02542f
C155 VDD2.n139 B 0.011387f
C156 VDD2.n140 B 0.020014f
C157 VDD2.n141 B 0.010755f
C158 VDD2.n142 B 0.02542f
C159 VDD2.n143 B 0.011387f
C160 VDD2.n144 B 1.72775f
C161 VDD2.n145 B 0.010755f
C162 VDD2.t1 B 0.042234f
C163 VDD2.n146 B 0.15382f
C164 VDD2.n147 B 0.015017f
C165 VDD2.n148 B 0.019065f
C166 VDD2.n149 B 0.02542f
C167 VDD2.n150 B 0.011387f
C168 VDD2.n151 B 0.010755f
C169 VDD2.n152 B 0.020014f
C170 VDD2.n153 B 0.020014f
C171 VDD2.n154 B 0.010755f
C172 VDD2.n155 B 0.011387f
C173 VDD2.n156 B 0.02542f
C174 VDD2.n157 B 0.02542f
C175 VDD2.n158 B 0.011387f
C176 VDD2.n159 B 0.010755f
C177 VDD2.n160 B 0.020014f
C178 VDD2.n161 B 0.020014f
C179 VDD2.n162 B 0.010755f
C180 VDD2.n163 B 0.011387f
C181 VDD2.n164 B 0.02542f
C182 VDD2.n165 B 0.02542f
C183 VDD2.n166 B 0.011387f
C184 VDD2.n167 B 0.010755f
C185 VDD2.n168 B 0.020014f
C186 VDD2.n169 B 0.020014f
C187 VDD2.n170 B 0.010755f
C188 VDD2.n171 B 0.011387f
C189 VDD2.n172 B 0.02542f
C190 VDD2.n173 B 0.02542f
C191 VDD2.n174 B 0.011387f
C192 VDD2.n175 B 0.010755f
C193 VDD2.n176 B 0.020014f
C194 VDD2.n177 B 0.020014f
C195 VDD2.n178 B 0.010755f
C196 VDD2.n179 B 0.011387f
C197 VDD2.n180 B 0.02542f
C198 VDD2.n181 B 0.02542f
C199 VDD2.n182 B 0.011387f
C200 VDD2.n183 B 0.010755f
C201 VDD2.n184 B 0.020014f
C202 VDD2.n185 B 0.020014f
C203 VDD2.n186 B 0.010755f
C204 VDD2.n187 B 0.011387f
C205 VDD2.n188 B 0.02542f
C206 VDD2.n189 B 0.02542f
C207 VDD2.n190 B 0.011387f
C208 VDD2.n191 B 0.010755f
C209 VDD2.n192 B 0.020014f
C210 VDD2.n193 B 0.020014f
C211 VDD2.n194 B 0.010755f
C212 VDD2.n195 B 0.011387f
C213 VDD2.n196 B 0.02542f
C214 VDD2.n197 B 0.02542f
C215 VDD2.n198 B 0.011387f
C216 VDD2.n199 B 0.010755f
C217 VDD2.n200 B 0.020014f
C218 VDD2.n201 B 0.020014f
C219 VDD2.n202 B 0.010755f
C220 VDD2.n203 B 0.011387f
C221 VDD2.n204 B 0.02542f
C222 VDD2.n205 B 0.02542f
C223 VDD2.n206 B 0.011387f
C224 VDD2.n207 B 0.010755f
C225 VDD2.n208 B 0.020014f
C226 VDD2.n209 B 0.020014f
C227 VDD2.n210 B 0.010755f
C228 VDD2.n211 B 0.011387f
C229 VDD2.n212 B 0.02542f
C230 VDD2.n213 B 0.055986f
C231 VDD2.n214 B 0.011387f
C232 VDD2.n215 B 0.010755f
C233 VDD2.n216 B 0.045168f
C234 VDD2.n217 B 0.045219f
C235 VDD2.n218 B 2.86801f
C236 VN.t1 B 3.42503f
C237 VN.t0 B 3.72089f
C238 VDD1.n0 B 0.028737f
C239 VDD1.n1 B 0.02006f
C240 VDD1.n2 B 0.010779f
C241 VDD1.n3 B 0.025478f
C242 VDD1.n4 B 0.011413f
C243 VDD1.n5 B 0.02006f
C244 VDD1.n6 B 0.010779f
C245 VDD1.n7 B 0.025478f
C246 VDD1.n8 B 0.011413f
C247 VDD1.n9 B 0.02006f
C248 VDD1.n10 B 0.010779f
C249 VDD1.n11 B 0.025478f
C250 VDD1.n12 B 0.011096f
C251 VDD1.n13 B 0.02006f
C252 VDD1.n14 B 0.011096f
C253 VDD1.n15 B 0.010779f
C254 VDD1.n16 B 0.025478f
C255 VDD1.n17 B 0.025478f
C256 VDD1.n18 B 0.011413f
C257 VDD1.n19 B 0.02006f
C258 VDD1.n20 B 0.010779f
C259 VDD1.n21 B 0.025478f
C260 VDD1.n22 B 0.011413f
C261 VDD1.n23 B 0.02006f
C262 VDD1.n24 B 0.010779f
C263 VDD1.n25 B 0.025478f
C264 VDD1.n26 B 0.011413f
C265 VDD1.n27 B 0.02006f
C266 VDD1.n28 B 0.010779f
C267 VDD1.n29 B 0.025478f
C268 VDD1.n30 B 0.011413f
C269 VDD1.n31 B 0.02006f
C270 VDD1.n32 B 0.010779f
C271 VDD1.n33 B 0.025478f
C272 VDD1.n34 B 0.011413f
C273 VDD1.n35 B 1.73171f
C274 VDD1.n36 B 0.010779f
C275 VDD1.t0 B 0.04233f
C276 VDD1.n37 B 0.154173f
C277 VDD1.n38 B 0.015051f
C278 VDD1.n39 B 0.019109f
C279 VDD1.n40 B 0.025478f
C280 VDD1.n41 B 0.011413f
C281 VDD1.n42 B 0.010779f
C282 VDD1.n43 B 0.02006f
C283 VDD1.n44 B 0.02006f
C284 VDD1.n45 B 0.010779f
C285 VDD1.n46 B 0.011413f
C286 VDD1.n47 B 0.025478f
C287 VDD1.n48 B 0.025478f
C288 VDD1.n49 B 0.011413f
C289 VDD1.n50 B 0.010779f
C290 VDD1.n51 B 0.02006f
C291 VDD1.n52 B 0.02006f
C292 VDD1.n53 B 0.010779f
C293 VDD1.n54 B 0.011413f
C294 VDD1.n55 B 0.025478f
C295 VDD1.n56 B 0.025478f
C296 VDD1.n57 B 0.011413f
C297 VDD1.n58 B 0.010779f
C298 VDD1.n59 B 0.02006f
C299 VDD1.n60 B 0.02006f
C300 VDD1.n61 B 0.010779f
C301 VDD1.n62 B 0.011413f
C302 VDD1.n63 B 0.025478f
C303 VDD1.n64 B 0.025478f
C304 VDD1.n65 B 0.011413f
C305 VDD1.n66 B 0.010779f
C306 VDD1.n67 B 0.02006f
C307 VDD1.n68 B 0.02006f
C308 VDD1.n69 B 0.010779f
C309 VDD1.n70 B 0.011413f
C310 VDD1.n71 B 0.025478f
C311 VDD1.n72 B 0.025478f
C312 VDD1.n73 B 0.011413f
C313 VDD1.n74 B 0.010779f
C314 VDD1.n75 B 0.02006f
C315 VDD1.n76 B 0.02006f
C316 VDD1.n77 B 0.010779f
C317 VDD1.n78 B 0.011413f
C318 VDD1.n79 B 0.025478f
C319 VDD1.n80 B 0.025478f
C320 VDD1.n81 B 0.011413f
C321 VDD1.n82 B 0.010779f
C322 VDD1.n83 B 0.02006f
C323 VDD1.n84 B 0.02006f
C324 VDD1.n85 B 0.010779f
C325 VDD1.n86 B 0.011413f
C326 VDD1.n87 B 0.025478f
C327 VDD1.n88 B 0.025478f
C328 VDD1.n89 B 0.011413f
C329 VDD1.n90 B 0.010779f
C330 VDD1.n91 B 0.02006f
C331 VDD1.n92 B 0.02006f
C332 VDD1.n93 B 0.010779f
C333 VDD1.n94 B 0.011413f
C334 VDD1.n95 B 0.025478f
C335 VDD1.n96 B 0.025478f
C336 VDD1.n97 B 0.011413f
C337 VDD1.n98 B 0.010779f
C338 VDD1.n99 B 0.02006f
C339 VDD1.n100 B 0.02006f
C340 VDD1.n101 B 0.010779f
C341 VDD1.n102 B 0.011413f
C342 VDD1.n103 B 0.025478f
C343 VDD1.n104 B 0.056114f
C344 VDD1.n105 B 0.011413f
C345 VDD1.n106 B 0.010779f
C346 VDD1.n107 B 0.045272f
C347 VDD1.n108 B 0.045891f
C348 VDD1.n109 B 0.028737f
C349 VDD1.n110 B 0.02006f
C350 VDD1.n111 B 0.010779f
C351 VDD1.n112 B 0.025478f
C352 VDD1.n113 B 0.011413f
C353 VDD1.n114 B 0.02006f
C354 VDD1.n115 B 0.010779f
C355 VDD1.n116 B 0.025478f
C356 VDD1.n117 B 0.011413f
C357 VDD1.n118 B 0.02006f
C358 VDD1.n119 B 0.010779f
C359 VDD1.n120 B 0.025478f
C360 VDD1.n121 B 0.011096f
C361 VDD1.n122 B 0.02006f
C362 VDD1.n123 B 0.011413f
C363 VDD1.n124 B 0.025478f
C364 VDD1.n125 B 0.011413f
C365 VDD1.n126 B 0.02006f
C366 VDD1.n127 B 0.010779f
C367 VDD1.n128 B 0.025478f
C368 VDD1.n129 B 0.011413f
C369 VDD1.n130 B 0.02006f
C370 VDD1.n131 B 0.010779f
C371 VDD1.n132 B 0.025478f
C372 VDD1.n133 B 0.011413f
C373 VDD1.n134 B 0.02006f
C374 VDD1.n135 B 0.010779f
C375 VDD1.n136 B 0.025478f
C376 VDD1.n137 B 0.011413f
C377 VDD1.n138 B 0.02006f
C378 VDD1.n139 B 0.010779f
C379 VDD1.n140 B 0.025478f
C380 VDD1.n141 B 0.011413f
C381 VDD1.n142 B 1.73171f
C382 VDD1.n143 B 0.010779f
C383 VDD1.t1 B 0.04233f
C384 VDD1.n144 B 0.154173f
C385 VDD1.n145 B 0.015051f
C386 VDD1.n146 B 0.019109f
C387 VDD1.n147 B 0.025478f
C388 VDD1.n148 B 0.011413f
C389 VDD1.n149 B 0.010779f
C390 VDD1.n150 B 0.02006f
C391 VDD1.n151 B 0.02006f
C392 VDD1.n152 B 0.010779f
C393 VDD1.n153 B 0.011413f
C394 VDD1.n154 B 0.025478f
C395 VDD1.n155 B 0.025478f
C396 VDD1.n156 B 0.011413f
C397 VDD1.n157 B 0.010779f
C398 VDD1.n158 B 0.02006f
C399 VDD1.n159 B 0.02006f
C400 VDD1.n160 B 0.010779f
C401 VDD1.n161 B 0.011413f
C402 VDD1.n162 B 0.025478f
C403 VDD1.n163 B 0.025478f
C404 VDD1.n164 B 0.011413f
C405 VDD1.n165 B 0.010779f
C406 VDD1.n166 B 0.02006f
C407 VDD1.n167 B 0.02006f
C408 VDD1.n168 B 0.010779f
C409 VDD1.n169 B 0.011413f
C410 VDD1.n170 B 0.025478f
C411 VDD1.n171 B 0.025478f
C412 VDD1.n172 B 0.011413f
C413 VDD1.n173 B 0.010779f
C414 VDD1.n174 B 0.02006f
C415 VDD1.n175 B 0.02006f
C416 VDD1.n176 B 0.010779f
C417 VDD1.n177 B 0.011413f
C418 VDD1.n178 B 0.025478f
C419 VDD1.n179 B 0.025478f
C420 VDD1.n180 B 0.011413f
C421 VDD1.n181 B 0.010779f
C422 VDD1.n182 B 0.02006f
C423 VDD1.n183 B 0.02006f
C424 VDD1.n184 B 0.010779f
C425 VDD1.n185 B 0.010779f
C426 VDD1.n186 B 0.011413f
C427 VDD1.n187 B 0.025478f
C428 VDD1.n188 B 0.025478f
C429 VDD1.n189 B 0.025478f
C430 VDD1.n190 B 0.011096f
C431 VDD1.n191 B 0.010779f
C432 VDD1.n192 B 0.02006f
C433 VDD1.n193 B 0.02006f
C434 VDD1.n194 B 0.010779f
C435 VDD1.n195 B 0.011413f
C436 VDD1.n196 B 0.025478f
C437 VDD1.n197 B 0.025478f
C438 VDD1.n198 B 0.011413f
C439 VDD1.n199 B 0.010779f
C440 VDD1.n200 B 0.02006f
C441 VDD1.n201 B 0.02006f
C442 VDD1.n202 B 0.010779f
C443 VDD1.n203 B 0.011413f
C444 VDD1.n204 B 0.025478f
C445 VDD1.n205 B 0.025478f
C446 VDD1.n206 B 0.011413f
C447 VDD1.n207 B 0.010779f
C448 VDD1.n208 B 0.02006f
C449 VDD1.n209 B 0.02006f
C450 VDD1.n210 B 0.010779f
C451 VDD1.n211 B 0.011413f
C452 VDD1.n212 B 0.025478f
C453 VDD1.n213 B 0.056114f
C454 VDD1.n214 B 0.011413f
C455 VDD1.n215 B 0.010779f
C456 VDD1.n216 B 0.045272f
C457 VDD1.n217 B 0.79136f
C458 VTAIL.n0 B 0.027964f
C459 VTAIL.n1 B 0.01952f
C460 VTAIL.n2 B 0.010489f
C461 VTAIL.n3 B 0.024793f
C462 VTAIL.n4 B 0.011106f
C463 VTAIL.n5 B 0.01952f
C464 VTAIL.n6 B 0.010489f
C465 VTAIL.n7 B 0.024793f
C466 VTAIL.n8 B 0.011106f
C467 VTAIL.n9 B 0.01952f
C468 VTAIL.n10 B 0.010489f
C469 VTAIL.n11 B 0.024793f
C470 VTAIL.n12 B 0.010798f
C471 VTAIL.n13 B 0.01952f
C472 VTAIL.n14 B 0.011106f
C473 VTAIL.n15 B 0.024793f
C474 VTAIL.n16 B 0.011106f
C475 VTAIL.n17 B 0.01952f
C476 VTAIL.n18 B 0.010489f
C477 VTAIL.n19 B 0.024793f
C478 VTAIL.n20 B 0.011106f
C479 VTAIL.n21 B 0.01952f
C480 VTAIL.n22 B 0.010489f
C481 VTAIL.n23 B 0.024793f
C482 VTAIL.n24 B 0.011106f
C483 VTAIL.n25 B 0.01952f
C484 VTAIL.n26 B 0.010489f
C485 VTAIL.n27 B 0.024793f
C486 VTAIL.n28 B 0.011106f
C487 VTAIL.n29 B 0.01952f
C488 VTAIL.n30 B 0.010489f
C489 VTAIL.n31 B 0.024793f
C490 VTAIL.n32 B 0.011106f
C491 VTAIL.n33 B 1.68512f
C492 VTAIL.n34 B 0.010489f
C493 VTAIL.t3 B 0.041191f
C494 VTAIL.n35 B 0.150025f
C495 VTAIL.n36 B 0.014646f
C496 VTAIL.n37 B 0.018595f
C497 VTAIL.n38 B 0.024793f
C498 VTAIL.n39 B 0.011106f
C499 VTAIL.n40 B 0.010489f
C500 VTAIL.n41 B 0.01952f
C501 VTAIL.n42 B 0.01952f
C502 VTAIL.n43 B 0.010489f
C503 VTAIL.n44 B 0.011106f
C504 VTAIL.n45 B 0.024793f
C505 VTAIL.n46 B 0.024793f
C506 VTAIL.n47 B 0.011106f
C507 VTAIL.n48 B 0.010489f
C508 VTAIL.n49 B 0.01952f
C509 VTAIL.n50 B 0.01952f
C510 VTAIL.n51 B 0.010489f
C511 VTAIL.n52 B 0.011106f
C512 VTAIL.n53 B 0.024793f
C513 VTAIL.n54 B 0.024793f
C514 VTAIL.n55 B 0.011106f
C515 VTAIL.n56 B 0.010489f
C516 VTAIL.n57 B 0.01952f
C517 VTAIL.n58 B 0.01952f
C518 VTAIL.n59 B 0.010489f
C519 VTAIL.n60 B 0.011106f
C520 VTAIL.n61 B 0.024793f
C521 VTAIL.n62 B 0.024793f
C522 VTAIL.n63 B 0.011106f
C523 VTAIL.n64 B 0.010489f
C524 VTAIL.n65 B 0.01952f
C525 VTAIL.n66 B 0.01952f
C526 VTAIL.n67 B 0.010489f
C527 VTAIL.n68 B 0.011106f
C528 VTAIL.n69 B 0.024793f
C529 VTAIL.n70 B 0.024793f
C530 VTAIL.n71 B 0.011106f
C531 VTAIL.n72 B 0.010489f
C532 VTAIL.n73 B 0.01952f
C533 VTAIL.n74 B 0.01952f
C534 VTAIL.n75 B 0.010489f
C535 VTAIL.n76 B 0.010489f
C536 VTAIL.n77 B 0.011106f
C537 VTAIL.n78 B 0.024793f
C538 VTAIL.n79 B 0.024793f
C539 VTAIL.n80 B 0.024793f
C540 VTAIL.n81 B 0.010798f
C541 VTAIL.n82 B 0.010489f
C542 VTAIL.n83 B 0.01952f
C543 VTAIL.n84 B 0.01952f
C544 VTAIL.n85 B 0.010489f
C545 VTAIL.n86 B 0.011106f
C546 VTAIL.n87 B 0.024793f
C547 VTAIL.n88 B 0.024793f
C548 VTAIL.n89 B 0.011106f
C549 VTAIL.n90 B 0.010489f
C550 VTAIL.n91 B 0.01952f
C551 VTAIL.n92 B 0.01952f
C552 VTAIL.n93 B 0.010489f
C553 VTAIL.n94 B 0.011106f
C554 VTAIL.n95 B 0.024793f
C555 VTAIL.n96 B 0.024793f
C556 VTAIL.n97 B 0.011106f
C557 VTAIL.n98 B 0.010489f
C558 VTAIL.n99 B 0.01952f
C559 VTAIL.n100 B 0.01952f
C560 VTAIL.n101 B 0.010489f
C561 VTAIL.n102 B 0.011106f
C562 VTAIL.n103 B 0.024793f
C563 VTAIL.n104 B 0.054604f
C564 VTAIL.n105 B 0.011106f
C565 VTAIL.n106 B 0.010489f
C566 VTAIL.n107 B 0.044054f
C567 VTAIL.n108 B 0.030616f
C568 VTAIL.n109 B 1.58557f
C569 VTAIL.n110 B 0.027964f
C570 VTAIL.n111 B 0.01952f
C571 VTAIL.n112 B 0.010489f
C572 VTAIL.n113 B 0.024793f
C573 VTAIL.n114 B 0.011106f
C574 VTAIL.n115 B 0.01952f
C575 VTAIL.n116 B 0.010489f
C576 VTAIL.n117 B 0.024793f
C577 VTAIL.n118 B 0.011106f
C578 VTAIL.n119 B 0.01952f
C579 VTAIL.n120 B 0.010489f
C580 VTAIL.n121 B 0.024793f
C581 VTAIL.n122 B 0.010798f
C582 VTAIL.n123 B 0.01952f
C583 VTAIL.n124 B 0.010798f
C584 VTAIL.n125 B 0.010489f
C585 VTAIL.n126 B 0.024793f
C586 VTAIL.n127 B 0.024793f
C587 VTAIL.n128 B 0.011106f
C588 VTAIL.n129 B 0.01952f
C589 VTAIL.n130 B 0.010489f
C590 VTAIL.n131 B 0.024793f
C591 VTAIL.n132 B 0.011106f
C592 VTAIL.n133 B 0.01952f
C593 VTAIL.n134 B 0.010489f
C594 VTAIL.n135 B 0.024793f
C595 VTAIL.n136 B 0.011106f
C596 VTAIL.n137 B 0.01952f
C597 VTAIL.n138 B 0.010489f
C598 VTAIL.n139 B 0.024793f
C599 VTAIL.n140 B 0.011106f
C600 VTAIL.n141 B 0.01952f
C601 VTAIL.n142 B 0.010489f
C602 VTAIL.n143 B 0.024793f
C603 VTAIL.n144 B 0.011106f
C604 VTAIL.n145 B 1.68512f
C605 VTAIL.n146 B 0.010489f
C606 VTAIL.t0 B 0.041191f
C607 VTAIL.n147 B 0.150025f
C608 VTAIL.n148 B 0.014646f
C609 VTAIL.n149 B 0.018595f
C610 VTAIL.n150 B 0.024793f
C611 VTAIL.n151 B 0.011106f
C612 VTAIL.n152 B 0.010489f
C613 VTAIL.n153 B 0.01952f
C614 VTAIL.n154 B 0.01952f
C615 VTAIL.n155 B 0.010489f
C616 VTAIL.n156 B 0.011106f
C617 VTAIL.n157 B 0.024793f
C618 VTAIL.n158 B 0.024793f
C619 VTAIL.n159 B 0.011106f
C620 VTAIL.n160 B 0.010489f
C621 VTAIL.n161 B 0.01952f
C622 VTAIL.n162 B 0.01952f
C623 VTAIL.n163 B 0.010489f
C624 VTAIL.n164 B 0.011106f
C625 VTAIL.n165 B 0.024793f
C626 VTAIL.n166 B 0.024793f
C627 VTAIL.n167 B 0.011106f
C628 VTAIL.n168 B 0.010489f
C629 VTAIL.n169 B 0.01952f
C630 VTAIL.n170 B 0.01952f
C631 VTAIL.n171 B 0.010489f
C632 VTAIL.n172 B 0.011106f
C633 VTAIL.n173 B 0.024793f
C634 VTAIL.n174 B 0.024793f
C635 VTAIL.n175 B 0.011106f
C636 VTAIL.n176 B 0.010489f
C637 VTAIL.n177 B 0.01952f
C638 VTAIL.n178 B 0.01952f
C639 VTAIL.n179 B 0.010489f
C640 VTAIL.n180 B 0.011106f
C641 VTAIL.n181 B 0.024793f
C642 VTAIL.n182 B 0.024793f
C643 VTAIL.n183 B 0.011106f
C644 VTAIL.n184 B 0.010489f
C645 VTAIL.n185 B 0.01952f
C646 VTAIL.n186 B 0.01952f
C647 VTAIL.n187 B 0.010489f
C648 VTAIL.n188 B 0.011106f
C649 VTAIL.n189 B 0.024793f
C650 VTAIL.n190 B 0.024793f
C651 VTAIL.n191 B 0.011106f
C652 VTAIL.n192 B 0.010489f
C653 VTAIL.n193 B 0.01952f
C654 VTAIL.n194 B 0.01952f
C655 VTAIL.n195 B 0.010489f
C656 VTAIL.n196 B 0.011106f
C657 VTAIL.n197 B 0.024793f
C658 VTAIL.n198 B 0.024793f
C659 VTAIL.n199 B 0.011106f
C660 VTAIL.n200 B 0.010489f
C661 VTAIL.n201 B 0.01952f
C662 VTAIL.n202 B 0.01952f
C663 VTAIL.n203 B 0.010489f
C664 VTAIL.n204 B 0.011106f
C665 VTAIL.n205 B 0.024793f
C666 VTAIL.n206 B 0.024793f
C667 VTAIL.n207 B 0.011106f
C668 VTAIL.n208 B 0.010489f
C669 VTAIL.n209 B 0.01952f
C670 VTAIL.n210 B 0.01952f
C671 VTAIL.n211 B 0.010489f
C672 VTAIL.n212 B 0.011106f
C673 VTAIL.n213 B 0.024793f
C674 VTAIL.n214 B 0.054604f
C675 VTAIL.n215 B 0.011106f
C676 VTAIL.n216 B 0.010489f
C677 VTAIL.n217 B 0.044054f
C678 VTAIL.n218 B 0.030616f
C679 VTAIL.n219 B 1.60482f
C680 VTAIL.n220 B 0.027964f
C681 VTAIL.n221 B 0.01952f
C682 VTAIL.n222 B 0.010489f
C683 VTAIL.n223 B 0.024793f
C684 VTAIL.n224 B 0.011106f
C685 VTAIL.n225 B 0.01952f
C686 VTAIL.n226 B 0.010489f
C687 VTAIL.n227 B 0.024793f
C688 VTAIL.n228 B 0.011106f
C689 VTAIL.n229 B 0.01952f
C690 VTAIL.n230 B 0.010489f
C691 VTAIL.n231 B 0.024793f
C692 VTAIL.n232 B 0.010798f
C693 VTAIL.n233 B 0.01952f
C694 VTAIL.n234 B 0.010798f
C695 VTAIL.n235 B 0.010489f
C696 VTAIL.n236 B 0.024793f
C697 VTAIL.n237 B 0.024793f
C698 VTAIL.n238 B 0.011106f
C699 VTAIL.n239 B 0.01952f
C700 VTAIL.n240 B 0.010489f
C701 VTAIL.n241 B 0.024793f
C702 VTAIL.n242 B 0.011106f
C703 VTAIL.n243 B 0.01952f
C704 VTAIL.n244 B 0.010489f
C705 VTAIL.n245 B 0.024793f
C706 VTAIL.n246 B 0.011106f
C707 VTAIL.n247 B 0.01952f
C708 VTAIL.n248 B 0.010489f
C709 VTAIL.n249 B 0.024793f
C710 VTAIL.n250 B 0.011106f
C711 VTAIL.n251 B 0.01952f
C712 VTAIL.n252 B 0.010489f
C713 VTAIL.n253 B 0.024793f
C714 VTAIL.n254 B 0.011106f
C715 VTAIL.n255 B 1.68512f
C716 VTAIL.n256 B 0.010489f
C717 VTAIL.t2 B 0.041191f
C718 VTAIL.n257 B 0.150025f
C719 VTAIL.n258 B 0.014646f
C720 VTAIL.n259 B 0.018595f
C721 VTAIL.n260 B 0.024793f
C722 VTAIL.n261 B 0.011106f
C723 VTAIL.n262 B 0.010489f
C724 VTAIL.n263 B 0.01952f
C725 VTAIL.n264 B 0.01952f
C726 VTAIL.n265 B 0.010489f
C727 VTAIL.n266 B 0.011106f
C728 VTAIL.n267 B 0.024793f
C729 VTAIL.n268 B 0.024793f
C730 VTAIL.n269 B 0.011106f
C731 VTAIL.n270 B 0.010489f
C732 VTAIL.n271 B 0.01952f
C733 VTAIL.n272 B 0.01952f
C734 VTAIL.n273 B 0.010489f
C735 VTAIL.n274 B 0.011106f
C736 VTAIL.n275 B 0.024793f
C737 VTAIL.n276 B 0.024793f
C738 VTAIL.n277 B 0.011106f
C739 VTAIL.n278 B 0.010489f
C740 VTAIL.n279 B 0.01952f
C741 VTAIL.n280 B 0.01952f
C742 VTAIL.n281 B 0.010489f
C743 VTAIL.n282 B 0.011106f
C744 VTAIL.n283 B 0.024793f
C745 VTAIL.n284 B 0.024793f
C746 VTAIL.n285 B 0.011106f
C747 VTAIL.n286 B 0.010489f
C748 VTAIL.n287 B 0.01952f
C749 VTAIL.n288 B 0.01952f
C750 VTAIL.n289 B 0.010489f
C751 VTAIL.n290 B 0.011106f
C752 VTAIL.n291 B 0.024793f
C753 VTAIL.n292 B 0.024793f
C754 VTAIL.n293 B 0.011106f
C755 VTAIL.n294 B 0.010489f
C756 VTAIL.n295 B 0.01952f
C757 VTAIL.n296 B 0.01952f
C758 VTAIL.n297 B 0.010489f
C759 VTAIL.n298 B 0.011106f
C760 VTAIL.n299 B 0.024793f
C761 VTAIL.n300 B 0.024793f
C762 VTAIL.n301 B 0.011106f
C763 VTAIL.n302 B 0.010489f
C764 VTAIL.n303 B 0.01952f
C765 VTAIL.n304 B 0.01952f
C766 VTAIL.n305 B 0.010489f
C767 VTAIL.n306 B 0.011106f
C768 VTAIL.n307 B 0.024793f
C769 VTAIL.n308 B 0.024793f
C770 VTAIL.n309 B 0.011106f
C771 VTAIL.n310 B 0.010489f
C772 VTAIL.n311 B 0.01952f
C773 VTAIL.n312 B 0.01952f
C774 VTAIL.n313 B 0.010489f
C775 VTAIL.n314 B 0.011106f
C776 VTAIL.n315 B 0.024793f
C777 VTAIL.n316 B 0.024793f
C778 VTAIL.n317 B 0.011106f
C779 VTAIL.n318 B 0.010489f
C780 VTAIL.n319 B 0.01952f
C781 VTAIL.n320 B 0.01952f
C782 VTAIL.n321 B 0.010489f
C783 VTAIL.n322 B 0.011106f
C784 VTAIL.n323 B 0.024793f
C785 VTAIL.n324 B 0.054604f
C786 VTAIL.n325 B 0.011106f
C787 VTAIL.n326 B 0.010489f
C788 VTAIL.n327 B 0.044054f
C789 VTAIL.n328 B 0.030616f
C790 VTAIL.n329 B 1.51318f
C791 VTAIL.n330 B 0.027964f
C792 VTAIL.n331 B 0.01952f
C793 VTAIL.n332 B 0.010489f
C794 VTAIL.n333 B 0.024793f
C795 VTAIL.n334 B 0.011106f
C796 VTAIL.n335 B 0.01952f
C797 VTAIL.n336 B 0.010489f
C798 VTAIL.n337 B 0.024793f
C799 VTAIL.n338 B 0.011106f
C800 VTAIL.n339 B 0.01952f
C801 VTAIL.n340 B 0.010489f
C802 VTAIL.n341 B 0.024793f
C803 VTAIL.n342 B 0.010798f
C804 VTAIL.n343 B 0.01952f
C805 VTAIL.n344 B 0.011106f
C806 VTAIL.n345 B 0.024793f
C807 VTAIL.n346 B 0.011106f
C808 VTAIL.n347 B 0.01952f
C809 VTAIL.n348 B 0.010489f
C810 VTAIL.n349 B 0.024793f
C811 VTAIL.n350 B 0.011106f
C812 VTAIL.n351 B 0.01952f
C813 VTAIL.n352 B 0.010489f
C814 VTAIL.n353 B 0.024793f
C815 VTAIL.n354 B 0.011106f
C816 VTAIL.n355 B 0.01952f
C817 VTAIL.n356 B 0.010489f
C818 VTAIL.n357 B 0.024793f
C819 VTAIL.n358 B 0.011106f
C820 VTAIL.n359 B 0.01952f
C821 VTAIL.n360 B 0.010489f
C822 VTAIL.n361 B 0.024793f
C823 VTAIL.n362 B 0.011106f
C824 VTAIL.n363 B 1.68512f
C825 VTAIL.n364 B 0.010489f
C826 VTAIL.t1 B 0.041191f
C827 VTAIL.n365 B 0.150025f
C828 VTAIL.n366 B 0.014646f
C829 VTAIL.n367 B 0.018595f
C830 VTAIL.n368 B 0.024793f
C831 VTAIL.n369 B 0.011106f
C832 VTAIL.n370 B 0.010489f
C833 VTAIL.n371 B 0.01952f
C834 VTAIL.n372 B 0.01952f
C835 VTAIL.n373 B 0.010489f
C836 VTAIL.n374 B 0.011106f
C837 VTAIL.n375 B 0.024793f
C838 VTAIL.n376 B 0.024793f
C839 VTAIL.n377 B 0.011106f
C840 VTAIL.n378 B 0.010489f
C841 VTAIL.n379 B 0.01952f
C842 VTAIL.n380 B 0.01952f
C843 VTAIL.n381 B 0.010489f
C844 VTAIL.n382 B 0.011106f
C845 VTAIL.n383 B 0.024793f
C846 VTAIL.n384 B 0.024793f
C847 VTAIL.n385 B 0.011106f
C848 VTAIL.n386 B 0.010489f
C849 VTAIL.n387 B 0.01952f
C850 VTAIL.n388 B 0.01952f
C851 VTAIL.n389 B 0.010489f
C852 VTAIL.n390 B 0.011106f
C853 VTAIL.n391 B 0.024793f
C854 VTAIL.n392 B 0.024793f
C855 VTAIL.n393 B 0.011106f
C856 VTAIL.n394 B 0.010489f
C857 VTAIL.n395 B 0.01952f
C858 VTAIL.n396 B 0.01952f
C859 VTAIL.n397 B 0.010489f
C860 VTAIL.n398 B 0.011106f
C861 VTAIL.n399 B 0.024793f
C862 VTAIL.n400 B 0.024793f
C863 VTAIL.n401 B 0.011106f
C864 VTAIL.n402 B 0.010489f
C865 VTAIL.n403 B 0.01952f
C866 VTAIL.n404 B 0.01952f
C867 VTAIL.n405 B 0.010489f
C868 VTAIL.n406 B 0.010489f
C869 VTAIL.n407 B 0.011106f
C870 VTAIL.n408 B 0.024793f
C871 VTAIL.n409 B 0.024793f
C872 VTAIL.n410 B 0.024793f
C873 VTAIL.n411 B 0.010798f
C874 VTAIL.n412 B 0.010489f
C875 VTAIL.n413 B 0.01952f
C876 VTAIL.n414 B 0.01952f
C877 VTAIL.n415 B 0.010489f
C878 VTAIL.n416 B 0.011106f
C879 VTAIL.n417 B 0.024793f
C880 VTAIL.n418 B 0.024793f
C881 VTAIL.n419 B 0.011106f
C882 VTAIL.n420 B 0.010489f
C883 VTAIL.n421 B 0.01952f
C884 VTAIL.n422 B 0.01952f
C885 VTAIL.n423 B 0.010489f
C886 VTAIL.n424 B 0.011106f
C887 VTAIL.n425 B 0.024793f
C888 VTAIL.n426 B 0.024793f
C889 VTAIL.n427 B 0.011106f
C890 VTAIL.n428 B 0.010489f
C891 VTAIL.n429 B 0.01952f
C892 VTAIL.n430 B 0.01952f
C893 VTAIL.n431 B 0.010489f
C894 VTAIL.n432 B 0.011106f
C895 VTAIL.n433 B 0.024793f
C896 VTAIL.n434 B 0.054604f
C897 VTAIL.n435 B 0.011106f
C898 VTAIL.n436 B 0.010489f
C899 VTAIL.n437 B 0.044054f
C900 VTAIL.n438 B 0.030616f
C901 VTAIL.n439 B 1.45706f
C902 VP.t1 B 3.79056f
C903 VP.t0 B 3.49239f
C904 VP.n0 B 6.07582f
.ends

