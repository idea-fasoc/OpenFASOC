* NGSPICE file created from diff_pair_sample_1288.ext - technology: sky130A

.subckt diff_pair_sample_1288 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t9 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
X1 B.t11 B.t9 B.t10 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=4.8321 pd=25.56 as=0 ps=0 w=12.39 l=1.85
X2 VTAIL.t17 VN.t1 VDD2.t6 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
X3 VDD2.t8 VN.t2 VTAIL.t16 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=4.8321 ps=25.56 w=12.39 l=1.85
X4 VDD2.t1 VN.t3 VTAIL.t15 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=4.8321 pd=25.56 as=2.04435 ps=12.72 w=12.39 l=1.85
X5 VDD1.t9 VP.t0 VTAIL.t4 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=4.8321 ps=25.56 w=12.39 l=1.85
X6 VDD1.t8 VP.t1 VTAIL.t2 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=4.8321 ps=25.56 w=12.39 l=1.85
X7 VTAIL.t8 VP.t2 VDD1.t7 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
X8 VTAIL.t1 VP.t3 VDD1.t6 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
X9 VTAIL.t14 VN.t4 VDD2.t5 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
X10 VDD1.t5 VP.t4 VTAIL.t7 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=4.8321 pd=25.56 as=2.04435 ps=12.72 w=12.39 l=1.85
X11 VDD2.t3 VN.t5 VTAIL.t13 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=4.8321 ps=25.56 w=12.39 l=1.85
X12 VTAIL.t19 VP.t5 VDD1.t4 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
X13 VDD1.t3 VP.t6 VTAIL.t5 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
X14 B.t8 B.t6 B.t7 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=4.8321 pd=25.56 as=0 ps=0 w=12.39 l=1.85
X15 B.t5 B.t3 B.t4 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=4.8321 pd=25.56 as=0 ps=0 w=12.39 l=1.85
X16 VTAIL.t12 VN.t6 VDD2.t0 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
X17 B.t2 B.t0 B.t1 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=4.8321 pd=25.56 as=0 ps=0 w=12.39 l=1.85
X18 VDD1.t2 VP.t7 VTAIL.t0 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=4.8321 pd=25.56 as=2.04435 ps=12.72 w=12.39 l=1.85
X19 VDD2.t2 VN.t7 VTAIL.t11 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
X20 VDD2.t7 VN.t8 VTAIL.t10 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
X21 VDD2.t4 VN.t9 VTAIL.t9 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=4.8321 pd=25.56 as=2.04435 ps=12.72 w=12.39 l=1.85
X22 VDD1.t1 VP.t8 VTAIL.t3 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
X23 VTAIL.t6 VP.t9 VDD1.t0 w_n3586_n3446# sky130_fd_pr__pfet_01v8 ad=2.04435 pd=12.72 as=2.04435 ps=12.72 w=12.39 l=1.85
R0 VN.n7 VN.t9 196.847
R1 VN.n39 VN.t5 196.847
R2 VN.n31 VN.n30 180.385
R3 VN.n63 VN.n62 180.385
R4 VN.n8 VN.t1 161.405
R5 VN.n15 VN.t7 161.405
R6 VN.n22 VN.t4 161.405
R7 VN.n30 VN.t2 161.405
R8 VN.n40 VN.t6 161.405
R9 VN.n47 VN.t8 161.405
R10 VN.n54 VN.t0 161.405
R11 VN.n62 VN.t3 161.405
R12 VN.n61 VN.n32 161.3
R13 VN.n60 VN.n59 161.3
R14 VN.n58 VN.n33 161.3
R15 VN.n57 VN.n56 161.3
R16 VN.n55 VN.n34 161.3
R17 VN.n53 VN.n52 161.3
R18 VN.n51 VN.n35 161.3
R19 VN.n50 VN.n49 161.3
R20 VN.n48 VN.n36 161.3
R21 VN.n46 VN.n45 161.3
R22 VN.n44 VN.n37 161.3
R23 VN.n43 VN.n42 161.3
R24 VN.n41 VN.n38 161.3
R25 VN.n29 VN.n0 161.3
R26 VN.n28 VN.n27 161.3
R27 VN.n26 VN.n1 161.3
R28 VN.n25 VN.n24 161.3
R29 VN.n23 VN.n2 161.3
R30 VN.n21 VN.n20 161.3
R31 VN.n19 VN.n3 161.3
R32 VN.n18 VN.n17 161.3
R33 VN.n16 VN.n4 161.3
R34 VN.n14 VN.n13 161.3
R35 VN.n12 VN.n5 161.3
R36 VN.n11 VN.n10 161.3
R37 VN.n9 VN.n6 161.3
R38 VN.n10 VN.n5 56.0336
R39 VN.n17 VN.n3 56.0336
R40 VN.n42 VN.n37 56.0336
R41 VN.n49 VN.n35 56.0336
R42 VN VN.n63 49.6539
R43 VN.n8 VN.n7 48.2603
R44 VN.n40 VN.n39 48.2603
R45 VN.n28 VN.n1 42.4359
R46 VN.n60 VN.n33 42.4359
R47 VN.n24 VN.n1 38.5509
R48 VN.n56 VN.n33 38.5509
R49 VN.n10 VN.n9 24.9531
R50 VN.n21 VN.n3 24.9531
R51 VN.n42 VN.n41 24.9531
R52 VN.n53 VN.n35 24.9531
R53 VN.n14 VN.n5 24.4675
R54 VN.n17 VN.n16 24.4675
R55 VN.n24 VN.n23 24.4675
R56 VN.n29 VN.n28 24.4675
R57 VN.n49 VN.n48 24.4675
R58 VN.n46 VN.n37 24.4675
R59 VN.n56 VN.n55 24.4675
R60 VN.n61 VN.n60 24.4675
R61 VN.n9 VN.n8 21.0421
R62 VN.n22 VN.n21 21.0421
R63 VN.n41 VN.n40 21.0421
R64 VN.n54 VN.n53 21.0421
R65 VN.n15 VN.n14 12.234
R66 VN.n16 VN.n15 12.234
R67 VN.n48 VN.n47 12.234
R68 VN.n47 VN.n46 12.234
R69 VN.n39 VN.n38 12.1797
R70 VN.n7 VN.n6 12.1797
R71 VN.n30 VN.n29 5.38324
R72 VN.n62 VN.n61 5.38324
R73 VN.n23 VN.n22 3.42588
R74 VN.n55 VN.n54 3.42588
R75 VN.n63 VN.n32 0.189894
R76 VN.n59 VN.n32 0.189894
R77 VN.n59 VN.n58 0.189894
R78 VN.n58 VN.n57 0.189894
R79 VN.n57 VN.n34 0.189894
R80 VN.n52 VN.n34 0.189894
R81 VN.n52 VN.n51 0.189894
R82 VN.n51 VN.n50 0.189894
R83 VN.n50 VN.n36 0.189894
R84 VN.n45 VN.n36 0.189894
R85 VN.n45 VN.n44 0.189894
R86 VN.n44 VN.n43 0.189894
R87 VN.n43 VN.n38 0.189894
R88 VN.n11 VN.n6 0.189894
R89 VN.n12 VN.n11 0.189894
R90 VN.n13 VN.n12 0.189894
R91 VN.n13 VN.n4 0.189894
R92 VN.n18 VN.n4 0.189894
R93 VN.n19 VN.n18 0.189894
R94 VN.n20 VN.n19 0.189894
R95 VN.n20 VN.n2 0.189894
R96 VN.n25 VN.n2 0.189894
R97 VN.n26 VN.n25 0.189894
R98 VN.n27 VN.n26 0.189894
R99 VN.n27 VN.n0 0.189894
R100 VN.n31 VN.n0 0.189894
R101 VN VN.n31 0.0516364
R102 VDD2.n1 VDD2.t4 76.1689
R103 VDD2.n4 VDD2.t1 74.2897
R104 VDD2.n3 VDD2.n2 73.0202
R105 VDD2 VDD2.n7 73.0174
R106 VDD2.n6 VDD2.n5 71.6663
R107 VDD2.n1 VDD2.n0 71.6661
R108 VDD2.n4 VDD2.n3 43.3231
R109 VDD2.n7 VDD2.t0 2.62399
R110 VDD2.n7 VDD2.t3 2.62399
R111 VDD2.n5 VDD2.t9 2.62399
R112 VDD2.n5 VDD2.t7 2.62399
R113 VDD2.n2 VDD2.t5 2.62399
R114 VDD2.n2 VDD2.t8 2.62399
R115 VDD2.n0 VDD2.t6 2.62399
R116 VDD2.n0 VDD2.t2 2.62399
R117 VDD2.n6 VDD2.n4 1.87981
R118 VDD2 VDD2.n6 0.528517
R119 VDD2.n3 VDD2.n1 0.414982
R120 VTAIL.n11 VTAIL.t13 57.6109
R121 VTAIL.n17 VTAIL.t16 57.6108
R122 VTAIL.n2 VTAIL.t2 57.6108
R123 VTAIL.n16 VTAIL.t4 57.6108
R124 VTAIL.n15 VTAIL.n14 54.9875
R125 VTAIL.n13 VTAIL.n12 54.9875
R126 VTAIL.n10 VTAIL.n9 54.9875
R127 VTAIL.n8 VTAIL.n7 54.9875
R128 VTAIL.n19 VTAIL.n18 54.9873
R129 VTAIL.n1 VTAIL.n0 54.9873
R130 VTAIL.n4 VTAIL.n3 54.9873
R131 VTAIL.n6 VTAIL.n5 54.9873
R132 VTAIL.n8 VTAIL.n6 26.8065
R133 VTAIL.n17 VTAIL.n16 24.9272
R134 VTAIL.n18 VTAIL.t11 2.62399
R135 VTAIL.n18 VTAIL.t14 2.62399
R136 VTAIL.n0 VTAIL.t9 2.62399
R137 VTAIL.n0 VTAIL.t17 2.62399
R138 VTAIL.n3 VTAIL.t5 2.62399
R139 VTAIL.n3 VTAIL.t19 2.62399
R140 VTAIL.n5 VTAIL.t7 2.62399
R141 VTAIL.n5 VTAIL.t8 2.62399
R142 VTAIL.n14 VTAIL.t3 2.62399
R143 VTAIL.n14 VTAIL.t1 2.62399
R144 VTAIL.n12 VTAIL.t0 2.62399
R145 VTAIL.n12 VTAIL.t6 2.62399
R146 VTAIL.n9 VTAIL.t10 2.62399
R147 VTAIL.n9 VTAIL.t12 2.62399
R148 VTAIL.n7 VTAIL.t15 2.62399
R149 VTAIL.n7 VTAIL.t18 2.62399
R150 VTAIL.n10 VTAIL.n8 1.87981
R151 VTAIL.n11 VTAIL.n10 1.87981
R152 VTAIL.n15 VTAIL.n13 1.87981
R153 VTAIL.n16 VTAIL.n15 1.87981
R154 VTAIL.n6 VTAIL.n4 1.87981
R155 VTAIL.n4 VTAIL.n2 1.87981
R156 VTAIL.n19 VTAIL.n17 1.87981
R157 VTAIL VTAIL.n1 1.46817
R158 VTAIL.n13 VTAIL.n11 1.40998
R159 VTAIL.n2 VTAIL.n1 1.40998
R160 VTAIL VTAIL.n19 0.412138
R161 B.n410 B.n409 585
R162 B.n408 B.n125 585
R163 B.n407 B.n406 585
R164 B.n405 B.n126 585
R165 B.n404 B.n403 585
R166 B.n402 B.n127 585
R167 B.n401 B.n400 585
R168 B.n399 B.n128 585
R169 B.n398 B.n397 585
R170 B.n396 B.n129 585
R171 B.n395 B.n394 585
R172 B.n393 B.n130 585
R173 B.n392 B.n391 585
R174 B.n390 B.n131 585
R175 B.n389 B.n388 585
R176 B.n387 B.n132 585
R177 B.n386 B.n385 585
R178 B.n384 B.n133 585
R179 B.n383 B.n382 585
R180 B.n381 B.n134 585
R181 B.n380 B.n379 585
R182 B.n378 B.n135 585
R183 B.n377 B.n376 585
R184 B.n375 B.n136 585
R185 B.n374 B.n373 585
R186 B.n372 B.n137 585
R187 B.n371 B.n370 585
R188 B.n369 B.n138 585
R189 B.n368 B.n367 585
R190 B.n366 B.n139 585
R191 B.n365 B.n364 585
R192 B.n363 B.n140 585
R193 B.n362 B.n361 585
R194 B.n360 B.n141 585
R195 B.n359 B.n358 585
R196 B.n357 B.n142 585
R197 B.n356 B.n355 585
R198 B.n354 B.n143 585
R199 B.n353 B.n352 585
R200 B.n351 B.n144 585
R201 B.n350 B.n349 585
R202 B.n348 B.n145 585
R203 B.n347 B.n346 585
R204 B.n344 B.n146 585
R205 B.n343 B.n342 585
R206 B.n341 B.n149 585
R207 B.n340 B.n339 585
R208 B.n338 B.n150 585
R209 B.n337 B.n336 585
R210 B.n335 B.n151 585
R211 B.n334 B.n333 585
R212 B.n332 B.n152 585
R213 B.n330 B.n329 585
R214 B.n328 B.n155 585
R215 B.n327 B.n326 585
R216 B.n325 B.n156 585
R217 B.n324 B.n323 585
R218 B.n322 B.n157 585
R219 B.n321 B.n320 585
R220 B.n319 B.n158 585
R221 B.n318 B.n317 585
R222 B.n316 B.n159 585
R223 B.n315 B.n314 585
R224 B.n313 B.n160 585
R225 B.n312 B.n311 585
R226 B.n310 B.n161 585
R227 B.n309 B.n308 585
R228 B.n307 B.n162 585
R229 B.n306 B.n305 585
R230 B.n304 B.n163 585
R231 B.n303 B.n302 585
R232 B.n301 B.n164 585
R233 B.n300 B.n299 585
R234 B.n298 B.n165 585
R235 B.n297 B.n296 585
R236 B.n295 B.n166 585
R237 B.n294 B.n293 585
R238 B.n292 B.n167 585
R239 B.n291 B.n290 585
R240 B.n289 B.n168 585
R241 B.n288 B.n287 585
R242 B.n286 B.n169 585
R243 B.n285 B.n284 585
R244 B.n283 B.n170 585
R245 B.n282 B.n281 585
R246 B.n280 B.n171 585
R247 B.n279 B.n278 585
R248 B.n277 B.n172 585
R249 B.n276 B.n275 585
R250 B.n274 B.n173 585
R251 B.n273 B.n272 585
R252 B.n271 B.n174 585
R253 B.n270 B.n269 585
R254 B.n268 B.n175 585
R255 B.n267 B.n266 585
R256 B.n411 B.n124 585
R257 B.n413 B.n412 585
R258 B.n414 B.n123 585
R259 B.n416 B.n415 585
R260 B.n417 B.n122 585
R261 B.n419 B.n418 585
R262 B.n420 B.n121 585
R263 B.n422 B.n421 585
R264 B.n423 B.n120 585
R265 B.n425 B.n424 585
R266 B.n426 B.n119 585
R267 B.n428 B.n427 585
R268 B.n429 B.n118 585
R269 B.n431 B.n430 585
R270 B.n432 B.n117 585
R271 B.n434 B.n433 585
R272 B.n435 B.n116 585
R273 B.n437 B.n436 585
R274 B.n438 B.n115 585
R275 B.n440 B.n439 585
R276 B.n441 B.n114 585
R277 B.n443 B.n442 585
R278 B.n444 B.n113 585
R279 B.n446 B.n445 585
R280 B.n447 B.n112 585
R281 B.n449 B.n448 585
R282 B.n450 B.n111 585
R283 B.n452 B.n451 585
R284 B.n453 B.n110 585
R285 B.n455 B.n454 585
R286 B.n456 B.n109 585
R287 B.n458 B.n457 585
R288 B.n459 B.n108 585
R289 B.n461 B.n460 585
R290 B.n462 B.n107 585
R291 B.n464 B.n463 585
R292 B.n465 B.n106 585
R293 B.n467 B.n466 585
R294 B.n468 B.n105 585
R295 B.n470 B.n469 585
R296 B.n471 B.n104 585
R297 B.n473 B.n472 585
R298 B.n474 B.n103 585
R299 B.n476 B.n475 585
R300 B.n477 B.n102 585
R301 B.n479 B.n478 585
R302 B.n480 B.n101 585
R303 B.n482 B.n481 585
R304 B.n483 B.n100 585
R305 B.n485 B.n484 585
R306 B.n486 B.n99 585
R307 B.n488 B.n487 585
R308 B.n489 B.n98 585
R309 B.n491 B.n490 585
R310 B.n492 B.n97 585
R311 B.n494 B.n493 585
R312 B.n495 B.n96 585
R313 B.n497 B.n496 585
R314 B.n498 B.n95 585
R315 B.n500 B.n499 585
R316 B.n501 B.n94 585
R317 B.n503 B.n502 585
R318 B.n504 B.n93 585
R319 B.n506 B.n505 585
R320 B.n507 B.n92 585
R321 B.n509 B.n508 585
R322 B.n510 B.n91 585
R323 B.n512 B.n511 585
R324 B.n513 B.n90 585
R325 B.n515 B.n514 585
R326 B.n516 B.n89 585
R327 B.n518 B.n517 585
R328 B.n519 B.n88 585
R329 B.n521 B.n520 585
R330 B.n522 B.n87 585
R331 B.n524 B.n523 585
R332 B.n525 B.n86 585
R333 B.n527 B.n526 585
R334 B.n528 B.n85 585
R335 B.n530 B.n529 585
R336 B.n531 B.n84 585
R337 B.n533 B.n532 585
R338 B.n534 B.n83 585
R339 B.n536 B.n535 585
R340 B.n537 B.n82 585
R341 B.n539 B.n538 585
R342 B.n540 B.n81 585
R343 B.n542 B.n541 585
R344 B.n543 B.n80 585
R345 B.n545 B.n544 585
R346 B.n546 B.n79 585
R347 B.n548 B.n547 585
R348 B.n549 B.n78 585
R349 B.n551 B.n550 585
R350 B.n694 B.n25 585
R351 B.n693 B.n692 585
R352 B.n691 B.n26 585
R353 B.n690 B.n689 585
R354 B.n688 B.n27 585
R355 B.n687 B.n686 585
R356 B.n685 B.n28 585
R357 B.n684 B.n683 585
R358 B.n682 B.n29 585
R359 B.n681 B.n680 585
R360 B.n679 B.n30 585
R361 B.n678 B.n677 585
R362 B.n676 B.n31 585
R363 B.n675 B.n674 585
R364 B.n673 B.n32 585
R365 B.n672 B.n671 585
R366 B.n670 B.n33 585
R367 B.n669 B.n668 585
R368 B.n667 B.n34 585
R369 B.n666 B.n665 585
R370 B.n664 B.n35 585
R371 B.n663 B.n662 585
R372 B.n661 B.n36 585
R373 B.n660 B.n659 585
R374 B.n658 B.n37 585
R375 B.n657 B.n656 585
R376 B.n655 B.n38 585
R377 B.n654 B.n653 585
R378 B.n652 B.n39 585
R379 B.n651 B.n650 585
R380 B.n649 B.n40 585
R381 B.n648 B.n647 585
R382 B.n646 B.n41 585
R383 B.n645 B.n644 585
R384 B.n643 B.n42 585
R385 B.n642 B.n641 585
R386 B.n640 B.n43 585
R387 B.n639 B.n638 585
R388 B.n637 B.n44 585
R389 B.n636 B.n635 585
R390 B.n634 B.n45 585
R391 B.n633 B.n632 585
R392 B.n631 B.n46 585
R393 B.n630 B.n629 585
R394 B.n628 B.n47 585
R395 B.n627 B.n626 585
R396 B.n625 B.n51 585
R397 B.n624 B.n623 585
R398 B.n622 B.n52 585
R399 B.n621 B.n620 585
R400 B.n619 B.n53 585
R401 B.n618 B.n617 585
R402 B.n615 B.n54 585
R403 B.n614 B.n613 585
R404 B.n612 B.n57 585
R405 B.n611 B.n610 585
R406 B.n609 B.n58 585
R407 B.n608 B.n607 585
R408 B.n606 B.n59 585
R409 B.n605 B.n604 585
R410 B.n603 B.n60 585
R411 B.n602 B.n601 585
R412 B.n600 B.n61 585
R413 B.n599 B.n598 585
R414 B.n597 B.n62 585
R415 B.n596 B.n595 585
R416 B.n594 B.n63 585
R417 B.n593 B.n592 585
R418 B.n591 B.n64 585
R419 B.n590 B.n589 585
R420 B.n588 B.n65 585
R421 B.n587 B.n586 585
R422 B.n585 B.n66 585
R423 B.n584 B.n583 585
R424 B.n582 B.n67 585
R425 B.n581 B.n580 585
R426 B.n579 B.n68 585
R427 B.n578 B.n577 585
R428 B.n576 B.n69 585
R429 B.n575 B.n574 585
R430 B.n573 B.n70 585
R431 B.n572 B.n571 585
R432 B.n570 B.n71 585
R433 B.n569 B.n568 585
R434 B.n567 B.n72 585
R435 B.n566 B.n565 585
R436 B.n564 B.n73 585
R437 B.n563 B.n562 585
R438 B.n561 B.n74 585
R439 B.n560 B.n559 585
R440 B.n558 B.n75 585
R441 B.n557 B.n556 585
R442 B.n555 B.n76 585
R443 B.n554 B.n553 585
R444 B.n552 B.n77 585
R445 B.n696 B.n695 585
R446 B.n697 B.n24 585
R447 B.n699 B.n698 585
R448 B.n700 B.n23 585
R449 B.n702 B.n701 585
R450 B.n703 B.n22 585
R451 B.n705 B.n704 585
R452 B.n706 B.n21 585
R453 B.n708 B.n707 585
R454 B.n709 B.n20 585
R455 B.n711 B.n710 585
R456 B.n712 B.n19 585
R457 B.n714 B.n713 585
R458 B.n715 B.n18 585
R459 B.n717 B.n716 585
R460 B.n718 B.n17 585
R461 B.n720 B.n719 585
R462 B.n721 B.n16 585
R463 B.n723 B.n722 585
R464 B.n724 B.n15 585
R465 B.n726 B.n725 585
R466 B.n727 B.n14 585
R467 B.n729 B.n728 585
R468 B.n730 B.n13 585
R469 B.n732 B.n731 585
R470 B.n733 B.n12 585
R471 B.n735 B.n734 585
R472 B.n736 B.n11 585
R473 B.n738 B.n737 585
R474 B.n739 B.n10 585
R475 B.n741 B.n740 585
R476 B.n742 B.n9 585
R477 B.n744 B.n743 585
R478 B.n745 B.n8 585
R479 B.n747 B.n746 585
R480 B.n748 B.n7 585
R481 B.n750 B.n749 585
R482 B.n751 B.n6 585
R483 B.n753 B.n752 585
R484 B.n754 B.n5 585
R485 B.n756 B.n755 585
R486 B.n757 B.n4 585
R487 B.n759 B.n758 585
R488 B.n760 B.n3 585
R489 B.n762 B.n761 585
R490 B.n763 B.n0 585
R491 B.n2 B.n1 585
R492 B.n199 B.n198 585
R493 B.n201 B.n200 585
R494 B.n202 B.n197 585
R495 B.n204 B.n203 585
R496 B.n205 B.n196 585
R497 B.n207 B.n206 585
R498 B.n208 B.n195 585
R499 B.n210 B.n209 585
R500 B.n211 B.n194 585
R501 B.n213 B.n212 585
R502 B.n214 B.n193 585
R503 B.n216 B.n215 585
R504 B.n217 B.n192 585
R505 B.n219 B.n218 585
R506 B.n220 B.n191 585
R507 B.n222 B.n221 585
R508 B.n223 B.n190 585
R509 B.n225 B.n224 585
R510 B.n226 B.n189 585
R511 B.n228 B.n227 585
R512 B.n229 B.n188 585
R513 B.n231 B.n230 585
R514 B.n232 B.n187 585
R515 B.n234 B.n233 585
R516 B.n235 B.n186 585
R517 B.n237 B.n236 585
R518 B.n238 B.n185 585
R519 B.n240 B.n239 585
R520 B.n241 B.n184 585
R521 B.n243 B.n242 585
R522 B.n244 B.n183 585
R523 B.n246 B.n245 585
R524 B.n247 B.n182 585
R525 B.n249 B.n248 585
R526 B.n250 B.n181 585
R527 B.n252 B.n251 585
R528 B.n253 B.n180 585
R529 B.n255 B.n254 585
R530 B.n256 B.n179 585
R531 B.n258 B.n257 585
R532 B.n259 B.n178 585
R533 B.n261 B.n260 585
R534 B.n262 B.n177 585
R535 B.n264 B.n263 585
R536 B.n265 B.n176 585
R537 B.n267 B.n176 521.33
R538 B.n409 B.n124 521.33
R539 B.n552 B.n551 521.33
R540 B.n696 B.n25 521.33
R541 B.n153 B.t9 367.947
R542 B.n147 B.t3 367.947
R543 B.n55 B.t6 367.947
R544 B.n48 B.t0 367.947
R545 B.n765 B.n764 256.663
R546 B.n764 B.n763 235.042
R547 B.n764 B.n2 235.042
R548 B.n268 B.n267 163.367
R549 B.n269 B.n268 163.367
R550 B.n269 B.n174 163.367
R551 B.n273 B.n174 163.367
R552 B.n274 B.n273 163.367
R553 B.n275 B.n274 163.367
R554 B.n275 B.n172 163.367
R555 B.n279 B.n172 163.367
R556 B.n280 B.n279 163.367
R557 B.n281 B.n280 163.367
R558 B.n281 B.n170 163.367
R559 B.n285 B.n170 163.367
R560 B.n286 B.n285 163.367
R561 B.n287 B.n286 163.367
R562 B.n287 B.n168 163.367
R563 B.n291 B.n168 163.367
R564 B.n292 B.n291 163.367
R565 B.n293 B.n292 163.367
R566 B.n293 B.n166 163.367
R567 B.n297 B.n166 163.367
R568 B.n298 B.n297 163.367
R569 B.n299 B.n298 163.367
R570 B.n299 B.n164 163.367
R571 B.n303 B.n164 163.367
R572 B.n304 B.n303 163.367
R573 B.n305 B.n304 163.367
R574 B.n305 B.n162 163.367
R575 B.n309 B.n162 163.367
R576 B.n310 B.n309 163.367
R577 B.n311 B.n310 163.367
R578 B.n311 B.n160 163.367
R579 B.n315 B.n160 163.367
R580 B.n316 B.n315 163.367
R581 B.n317 B.n316 163.367
R582 B.n317 B.n158 163.367
R583 B.n321 B.n158 163.367
R584 B.n322 B.n321 163.367
R585 B.n323 B.n322 163.367
R586 B.n323 B.n156 163.367
R587 B.n327 B.n156 163.367
R588 B.n328 B.n327 163.367
R589 B.n329 B.n328 163.367
R590 B.n329 B.n152 163.367
R591 B.n334 B.n152 163.367
R592 B.n335 B.n334 163.367
R593 B.n336 B.n335 163.367
R594 B.n336 B.n150 163.367
R595 B.n340 B.n150 163.367
R596 B.n341 B.n340 163.367
R597 B.n342 B.n341 163.367
R598 B.n342 B.n146 163.367
R599 B.n347 B.n146 163.367
R600 B.n348 B.n347 163.367
R601 B.n349 B.n348 163.367
R602 B.n349 B.n144 163.367
R603 B.n353 B.n144 163.367
R604 B.n354 B.n353 163.367
R605 B.n355 B.n354 163.367
R606 B.n355 B.n142 163.367
R607 B.n359 B.n142 163.367
R608 B.n360 B.n359 163.367
R609 B.n361 B.n360 163.367
R610 B.n361 B.n140 163.367
R611 B.n365 B.n140 163.367
R612 B.n366 B.n365 163.367
R613 B.n367 B.n366 163.367
R614 B.n367 B.n138 163.367
R615 B.n371 B.n138 163.367
R616 B.n372 B.n371 163.367
R617 B.n373 B.n372 163.367
R618 B.n373 B.n136 163.367
R619 B.n377 B.n136 163.367
R620 B.n378 B.n377 163.367
R621 B.n379 B.n378 163.367
R622 B.n379 B.n134 163.367
R623 B.n383 B.n134 163.367
R624 B.n384 B.n383 163.367
R625 B.n385 B.n384 163.367
R626 B.n385 B.n132 163.367
R627 B.n389 B.n132 163.367
R628 B.n390 B.n389 163.367
R629 B.n391 B.n390 163.367
R630 B.n391 B.n130 163.367
R631 B.n395 B.n130 163.367
R632 B.n396 B.n395 163.367
R633 B.n397 B.n396 163.367
R634 B.n397 B.n128 163.367
R635 B.n401 B.n128 163.367
R636 B.n402 B.n401 163.367
R637 B.n403 B.n402 163.367
R638 B.n403 B.n126 163.367
R639 B.n407 B.n126 163.367
R640 B.n408 B.n407 163.367
R641 B.n409 B.n408 163.367
R642 B.n551 B.n78 163.367
R643 B.n547 B.n78 163.367
R644 B.n547 B.n546 163.367
R645 B.n546 B.n545 163.367
R646 B.n545 B.n80 163.367
R647 B.n541 B.n80 163.367
R648 B.n541 B.n540 163.367
R649 B.n540 B.n539 163.367
R650 B.n539 B.n82 163.367
R651 B.n535 B.n82 163.367
R652 B.n535 B.n534 163.367
R653 B.n534 B.n533 163.367
R654 B.n533 B.n84 163.367
R655 B.n529 B.n84 163.367
R656 B.n529 B.n528 163.367
R657 B.n528 B.n527 163.367
R658 B.n527 B.n86 163.367
R659 B.n523 B.n86 163.367
R660 B.n523 B.n522 163.367
R661 B.n522 B.n521 163.367
R662 B.n521 B.n88 163.367
R663 B.n517 B.n88 163.367
R664 B.n517 B.n516 163.367
R665 B.n516 B.n515 163.367
R666 B.n515 B.n90 163.367
R667 B.n511 B.n90 163.367
R668 B.n511 B.n510 163.367
R669 B.n510 B.n509 163.367
R670 B.n509 B.n92 163.367
R671 B.n505 B.n92 163.367
R672 B.n505 B.n504 163.367
R673 B.n504 B.n503 163.367
R674 B.n503 B.n94 163.367
R675 B.n499 B.n94 163.367
R676 B.n499 B.n498 163.367
R677 B.n498 B.n497 163.367
R678 B.n497 B.n96 163.367
R679 B.n493 B.n96 163.367
R680 B.n493 B.n492 163.367
R681 B.n492 B.n491 163.367
R682 B.n491 B.n98 163.367
R683 B.n487 B.n98 163.367
R684 B.n487 B.n486 163.367
R685 B.n486 B.n485 163.367
R686 B.n485 B.n100 163.367
R687 B.n481 B.n100 163.367
R688 B.n481 B.n480 163.367
R689 B.n480 B.n479 163.367
R690 B.n479 B.n102 163.367
R691 B.n475 B.n102 163.367
R692 B.n475 B.n474 163.367
R693 B.n474 B.n473 163.367
R694 B.n473 B.n104 163.367
R695 B.n469 B.n104 163.367
R696 B.n469 B.n468 163.367
R697 B.n468 B.n467 163.367
R698 B.n467 B.n106 163.367
R699 B.n463 B.n106 163.367
R700 B.n463 B.n462 163.367
R701 B.n462 B.n461 163.367
R702 B.n461 B.n108 163.367
R703 B.n457 B.n108 163.367
R704 B.n457 B.n456 163.367
R705 B.n456 B.n455 163.367
R706 B.n455 B.n110 163.367
R707 B.n451 B.n110 163.367
R708 B.n451 B.n450 163.367
R709 B.n450 B.n449 163.367
R710 B.n449 B.n112 163.367
R711 B.n445 B.n112 163.367
R712 B.n445 B.n444 163.367
R713 B.n444 B.n443 163.367
R714 B.n443 B.n114 163.367
R715 B.n439 B.n114 163.367
R716 B.n439 B.n438 163.367
R717 B.n438 B.n437 163.367
R718 B.n437 B.n116 163.367
R719 B.n433 B.n116 163.367
R720 B.n433 B.n432 163.367
R721 B.n432 B.n431 163.367
R722 B.n431 B.n118 163.367
R723 B.n427 B.n118 163.367
R724 B.n427 B.n426 163.367
R725 B.n426 B.n425 163.367
R726 B.n425 B.n120 163.367
R727 B.n421 B.n120 163.367
R728 B.n421 B.n420 163.367
R729 B.n420 B.n419 163.367
R730 B.n419 B.n122 163.367
R731 B.n415 B.n122 163.367
R732 B.n415 B.n414 163.367
R733 B.n414 B.n413 163.367
R734 B.n413 B.n124 163.367
R735 B.n692 B.n25 163.367
R736 B.n692 B.n691 163.367
R737 B.n691 B.n690 163.367
R738 B.n690 B.n27 163.367
R739 B.n686 B.n27 163.367
R740 B.n686 B.n685 163.367
R741 B.n685 B.n684 163.367
R742 B.n684 B.n29 163.367
R743 B.n680 B.n29 163.367
R744 B.n680 B.n679 163.367
R745 B.n679 B.n678 163.367
R746 B.n678 B.n31 163.367
R747 B.n674 B.n31 163.367
R748 B.n674 B.n673 163.367
R749 B.n673 B.n672 163.367
R750 B.n672 B.n33 163.367
R751 B.n668 B.n33 163.367
R752 B.n668 B.n667 163.367
R753 B.n667 B.n666 163.367
R754 B.n666 B.n35 163.367
R755 B.n662 B.n35 163.367
R756 B.n662 B.n661 163.367
R757 B.n661 B.n660 163.367
R758 B.n660 B.n37 163.367
R759 B.n656 B.n37 163.367
R760 B.n656 B.n655 163.367
R761 B.n655 B.n654 163.367
R762 B.n654 B.n39 163.367
R763 B.n650 B.n39 163.367
R764 B.n650 B.n649 163.367
R765 B.n649 B.n648 163.367
R766 B.n648 B.n41 163.367
R767 B.n644 B.n41 163.367
R768 B.n644 B.n643 163.367
R769 B.n643 B.n642 163.367
R770 B.n642 B.n43 163.367
R771 B.n638 B.n43 163.367
R772 B.n638 B.n637 163.367
R773 B.n637 B.n636 163.367
R774 B.n636 B.n45 163.367
R775 B.n632 B.n45 163.367
R776 B.n632 B.n631 163.367
R777 B.n631 B.n630 163.367
R778 B.n630 B.n47 163.367
R779 B.n626 B.n47 163.367
R780 B.n626 B.n625 163.367
R781 B.n625 B.n624 163.367
R782 B.n624 B.n52 163.367
R783 B.n620 B.n52 163.367
R784 B.n620 B.n619 163.367
R785 B.n619 B.n618 163.367
R786 B.n618 B.n54 163.367
R787 B.n613 B.n54 163.367
R788 B.n613 B.n612 163.367
R789 B.n612 B.n611 163.367
R790 B.n611 B.n58 163.367
R791 B.n607 B.n58 163.367
R792 B.n607 B.n606 163.367
R793 B.n606 B.n605 163.367
R794 B.n605 B.n60 163.367
R795 B.n601 B.n60 163.367
R796 B.n601 B.n600 163.367
R797 B.n600 B.n599 163.367
R798 B.n599 B.n62 163.367
R799 B.n595 B.n62 163.367
R800 B.n595 B.n594 163.367
R801 B.n594 B.n593 163.367
R802 B.n593 B.n64 163.367
R803 B.n589 B.n64 163.367
R804 B.n589 B.n588 163.367
R805 B.n588 B.n587 163.367
R806 B.n587 B.n66 163.367
R807 B.n583 B.n66 163.367
R808 B.n583 B.n582 163.367
R809 B.n582 B.n581 163.367
R810 B.n581 B.n68 163.367
R811 B.n577 B.n68 163.367
R812 B.n577 B.n576 163.367
R813 B.n576 B.n575 163.367
R814 B.n575 B.n70 163.367
R815 B.n571 B.n70 163.367
R816 B.n571 B.n570 163.367
R817 B.n570 B.n569 163.367
R818 B.n569 B.n72 163.367
R819 B.n565 B.n72 163.367
R820 B.n565 B.n564 163.367
R821 B.n564 B.n563 163.367
R822 B.n563 B.n74 163.367
R823 B.n559 B.n74 163.367
R824 B.n559 B.n558 163.367
R825 B.n558 B.n557 163.367
R826 B.n557 B.n76 163.367
R827 B.n553 B.n76 163.367
R828 B.n553 B.n552 163.367
R829 B.n697 B.n696 163.367
R830 B.n698 B.n697 163.367
R831 B.n698 B.n23 163.367
R832 B.n702 B.n23 163.367
R833 B.n703 B.n702 163.367
R834 B.n704 B.n703 163.367
R835 B.n704 B.n21 163.367
R836 B.n708 B.n21 163.367
R837 B.n709 B.n708 163.367
R838 B.n710 B.n709 163.367
R839 B.n710 B.n19 163.367
R840 B.n714 B.n19 163.367
R841 B.n715 B.n714 163.367
R842 B.n716 B.n715 163.367
R843 B.n716 B.n17 163.367
R844 B.n720 B.n17 163.367
R845 B.n721 B.n720 163.367
R846 B.n722 B.n721 163.367
R847 B.n722 B.n15 163.367
R848 B.n726 B.n15 163.367
R849 B.n727 B.n726 163.367
R850 B.n728 B.n727 163.367
R851 B.n728 B.n13 163.367
R852 B.n732 B.n13 163.367
R853 B.n733 B.n732 163.367
R854 B.n734 B.n733 163.367
R855 B.n734 B.n11 163.367
R856 B.n738 B.n11 163.367
R857 B.n739 B.n738 163.367
R858 B.n740 B.n739 163.367
R859 B.n740 B.n9 163.367
R860 B.n744 B.n9 163.367
R861 B.n745 B.n744 163.367
R862 B.n746 B.n745 163.367
R863 B.n746 B.n7 163.367
R864 B.n750 B.n7 163.367
R865 B.n751 B.n750 163.367
R866 B.n752 B.n751 163.367
R867 B.n752 B.n5 163.367
R868 B.n756 B.n5 163.367
R869 B.n757 B.n756 163.367
R870 B.n758 B.n757 163.367
R871 B.n758 B.n3 163.367
R872 B.n762 B.n3 163.367
R873 B.n763 B.n762 163.367
R874 B.n198 B.n2 163.367
R875 B.n201 B.n198 163.367
R876 B.n202 B.n201 163.367
R877 B.n203 B.n202 163.367
R878 B.n203 B.n196 163.367
R879 B.n207 B.n196 163.367
R880 B.n208 B.n207 163.367
R881 B.n209 B.n208 163.367
R882 B.n209 B.n194 163.367
R883 B.n213 B.n194 163.367
R884 B.n214 B.n213 163.367
R885 B.n215 B.n214 163.367
R886 B.n215 B.n192 163.367
R887 B.n219 B.n192 163.367
R888 B.n220 B.n219 163.367
R889 B.n221 B.n220 163.367
R890 B.n221 B.n190 163.367
R891 B.n225 B.n190 163.367
R892 B.n226 B.n225 163.367
R893 B.n227 B.n226 163.367
R894 B.n227 B.n188 163.367
R895 B.n231 B.n188 163.367
R896 B.n232 B.n231 163.367
R897 B.n233 B.n232 163.367
R898 B.n233 B.n186 163.367
R899 B.n237 B.n186 163.367
R900 B.n238 B.n237 163.367
R901 B.n239 B.n238 163.367
R902 B.n239 B.n184 163.367
R903 B.n243 B.n184 163.367
R904 B.n244 B.n243 163.367
R905 B.n245 B.n244 163.367
R906 B.n245 B.n182 163.367
R907 B.n249 B.n182 163.367
R908 B.n250 B.n249 163.367
R909 B.n251 B.n250 163.367
R910 B.n251 B.n180 163.367
R911 B.n255 B.n180 163.367
R912 B.n256 B.n255 163.367
R913 B.n257 B.n256 163.367
R914 B.n257 B.n178 163.367
R915 B.n261 B.n178 163.367
R916 B.n262 B.n261 163.367
R917 B.n263 B.n262 163.367
R918 B.n263 B.n176 163.367
R919 B.n147 B.t4 152.207
R920 B.n55 B.t8 152.207
R921 B.n153 B.t10 152.191
R922 B.n48 B.t2 152.191
R923 B.n148 B.t5 109.927
R924 B.n56 B.t7 109.927
R925 B.n154 B.t11 109.912
R926 B.n49 B.t1 109.912
R927 B.n331 B.n154 59.5399
R928 B.n345 B.n148 59.5399
R929 B.n616 B.n56 59.5399
R930 B.n50 B.n49 59.5399
R931 B.n154 B.n153 42.2793
R932 B.n148 B.n147 42.2793
R933 B.n56 B.n55 42.2793
R934 B.n49 B.n48 42.2793
R935 B.n695 B.n694 33.8737
R936 B.n550 B.n77 33.8737
R937 B.n411 B.n410 33.8737
R938 B.n266 B.n265 33.8737
R939 B B.n765 18.0485
R940 B.n695 B.n24 10.6151
R941 B.n699 B.n24 10.6151
R942 B.n700 B.n699 10.6151
R943 B.n701 B.n700 10.6151
R944 B.n701 B.n22 10.6151
R945 B.n705 B.n22 10.6151
R946 B.n706 B.n705 10.6151
R947 B.n707 B.n706 10.6151
R948 B.n707 B.n20 10.6151
R949 B.n711 B.n20 10.6151
R950 B.n712 B.n711 10.6151
R951 B.n713 B.n712 10.6151
R952 B.n713 B.n18 10.6151
R953 B.n717 B.n18 10.6151
R954 B.n718 B.n717 10.6151
R955 B.n719 B.n718 10.6151
R956 B.n719 B.n16 10.6151
R957 B.n723 B.n16 10.6151
R958 B.n724 B.n723 10.6151
R959 B.n725 B.n724 10.6151
R960 B.n725 B.n14 10.6151
R961 B.n729 B.n14 10.6151
R962 B.n730 B.n729 10.6151
R963 B.n731 B.n730 10.6151
R964 B.n731 B.n12 10.6151
R965 B.n735 B.n12 10.6151
R966 B.n736 B.n735 10.6151
R967 B.n737 B.n736 10.6151
R968 B.n737 B.n10 10.6151
R969 B.n741 B.n10 10.6151
R970 B.n742 B.n741 10.6151
R971 B.n743 B.n742 10.6151
R972 B.n743 B.n8 10.6151
R973 B.n747 B.n8 10.6151
R974 B.n748 B.n747 10.6151
R975 B.n749 B.n748 10.6151
R976 B.n749 B.n6 10.6151
R977 B.n753 B.n6 10.6151
R978 B.n754 B.n753 10.6151
R979 B.n755 B.n754 10.6151
R980 B.n755 B.n4 10.6151
R981 B.n759 B.n4 10.6151
R982 B.n760 B.n759 10.6151
R983 B.n761 B.n760 10.6151
R984 B.n761 B.n0 10.6151
R985 B.n694 B.n693 10.6151
R986 B.n693 B.n26 10.6151
R987 B.n689 B.n26 10.6151
R988 B.n689 B.n688 10.6151
R989 B.n688 B.n687 10.6151
R990 B.n687 B.n28 10.6151
R991 B.n683 B.n28 10.6151
R992 B.n683 B.n682 10.6151
R993 B.n682 B.n681 10.6151
R994 B.n681 B.n30 10.6151
R995 B.n677 B.n30 10.6151
R996 B.n677 B.n676 10.6151
R997 B.n676 B.n675 10.6151
R998 B.n675 B.n32 10.6151
R999 B.n671 B.n32 10.6151
R1000 B.n671 B.n670 10.6151
R1001 B.n670 B.n669 10.6151
R1002 B.n669 B.n34 10.6151
R1003 B.n665 B.n34 10.6151
R1004 B.n665 B.n664 10.6151
R1005 B.n664 B.n663 10.6151
R1006 B.n663 B.n36 10.6151
R1007 B.n659 B.n36 10.6151
R1008 B.n659 B.n658 10.6151
R1009 B.n658 B.n657 10.6151
R1010 B.n657 B.n38 10.6151
R1011 B.n653 B.n38 10.6151
R1012 B.n653 B.n652 10.6151
R1013 B.n652 B.n651 10.6151
R1014 B.n651 B.n40 10.6151
R1015 B.n647 B.n40 10.6151
R1016 B.n647 B.n646 10.6151
R1017 B.n646 B.n645 10.6151
R1018 B.n645 B.n42 10.6151
R1019 B.n641 B.n42 10.6151
R1020 B.n641 B.n640 10.6151
R1021 B.n640 B.n639 10.6151
R1022 B.n639 B.n44 10.6151
R1023 B.n635 B.n44 10.6151
R1024 B.n635 B.n634 10.6151
R1025 B.n634 B.n633 10.6151
R1026 B.n633 B.n46 10.6151
R1027 B.n629 B.n628 10.6151
R1028 B.n628 B.n627 10.6151
R1029 B.n627 B.n51 10.6151
R1030 B.n623 B.n51 10.6151
R1031 B.n623 B.n622 10.6151
R1032 B.n622 B.n621 10.6151
R1033 B.n621 B.n53 10.6151
R1034 B.n617 B.n53 10.6151
R1035 B.n615 B.n614 10.6151
R1036 B.n614 B.n57 10.6151
R1037 B.n610 B.n57 10.6151
R1038 B.n610 B.n609 10.6151
R1039 B.n609 B.n608 10.6151
R1040 B.n608 B.n59 10.6151
R1041 B.n604 B.n59 10.6151
R1042 B.n604 B.n603 10.6151
R1043 B.n603 B.n602 10.6151
R1044 B.n602 B.n61 10.6151
R1045 B.n598 B.n61 10.6151
R1046 B.n598 B.n597 10.6151
R1047 B.n597 B.n596 10.6151
R1048 B.n596 B.n63 10.6151
R1049 B.n592 B.n63 10.6151
R1050 B.n592 B.n591 10.6151
R1051 B.n591 B.n590 10.6151
R1052 B.n590 B.n65 10.6151
R1053 B.n586 B.n65 10.6151
R1054 B.n586 B.n585 10.6151
R1055 B.n585 B.n584 10.6151
R1056 B.n584 B.n67 10.6151
R1057 B.n580 B.n67 10.6151
R1058 B.n580 B.n579 10.6151
R1059 B.n579 B.n578 10.6151
R1060 B.n578 B.n69 10.6151
R1061 B.n574 B.n69 10.6151
R1062 B.n574 B.n573 10.6151
R1063 B.n573 B.n572 10.6151
R1064 B.n572 B.n71 10.6151
R1065 B.n568 B.n71 10.6151
R1066 B.n568 B.n567 10.6151
R1067 B.n567 B.n566 10.6151
R1068 B.n566 B.n73 10.6151
R1069 B.n562 B.n73 10.6151
R1070 B.n562 B.n561 10.6151
R1071 B.n561 B.n560 10.6151
R1072 B.n560 B.n75 10.6151
R1073 B.n556 B.n75 10.6151
R1074 B.n556 B.n555 10.6151
R1075 B.n555 B.n554 10.6151
R1076 B.n554 B.n77 10.6151
R1077 B.n550 B.n549 10.6151
R1078 B.n549 B.n548 10.6151
R1079 B.n548 B.n79 10.6151
R1080 B.n544 B.n79 10.6151
R1081 B.n544 B.n543 10.6151
R1082 B.n543 B.n542 10.6151
R1083 B.n542 B.n81 10.6151
R1084 B.n538 B.n81 10.6151
R1085 B.n538 B.n537 10.6151
R1086 B.n537 B.n536 10.6151
R1087 B.n536 B.n83 10.6151
R1088 B.n532 B.n83 10.6151
R1089 B.n532 B.n531 10.6151
R1090 B.n531 B.n530 10.6151
R1091 B.n530 B.n85 10.6151
R1092 B.n526 B.n85 10.6151
R1093 B.n526 B.n525 10.6151
R1094 B.n525 B.n524 10.6151
R1095 B.n524 B.n87 10.6151
R1096 B.n520 B.n87 10.6151
R1097 B.n520 B.n519 10.6151
R1098 B.n519 B.n518 10.6151
R1099 B.n518 B.n89 10.6151
R1100 B.n514 B.n89 10.6151
R1101 B.n514 B.n513 10.6151
R1102 B.n513 B.n512 10.6151
R1103 B.n512 B.n91 10.6151
R1104 B.n508 B.n91 10.6151
R1105 B.n508 B.n507 10.6151
R1106 B.n507 B.n506 10.6151
R1107 B.n506 B.n93 10.6151
R1108 B.n502 B.n93 10.6151
R1109 B.n502 B.n501 10.6151
R1110 B.n501 B.n500 10.6151
R1111 B.n500 B.n95 10.6151
R1112 B.n496 B.n95 10.6151
R1113 B.n496 B.n495 10.6151
R1114 B.n495 B.n494 10.6151
R1115 B.n494 B.n97 10.6151
R1116 B.n490 B.n97 10.6151
R1117 B.n490 B.n489 10.6151
R1118 B.n489 B.n488 10.6151
R1119 B.n488 B.n99 10.6151
R1120 B.n484 B.n99 10.6151
R1121 B.n484 B.n483 10.6151
R1122 B.n483 B.n482 10.6151
R1123 B.n482 B.n101 10.6151
R1124 B.n478 B.n101 10.6151
R1125 B.n478 B.n477 10.6151
R1126 B.n477 B.n476 10.6151
R1127 B.n476 B.n103 10.6151
R1128 B.n472 B.n103 10.6151
R1129 B.n472 B.n471 10.6151
R1130 B.n471 B.n470 10.6151
R1131 B.n470 B.n105 10.6151
R1132 B.n466 B.n105 10.6151
R1133 B.n466 B.n465 10.6151
R1134 B.n465 B.n464 10.6151
R1135 B.n464 B.n107 10.6151
R1136 B.n460 B.n107 10.6151
R1137 B.n460 B.n459 10.6151
R1138 B.n459 B.n458 10.6151
R1139 B.n458 B.n109 10.6151
R1140 B.n454 B.n109 10.6151
R1141 B.n454 B.n453 10.6151
R1142 B.n453 B.n452 10.6151
R1143 B.n452 B.n111 10.6151
R1144 B.n448 B.n111 10.6151
R1145 B.n448 B.n447 10.6151
R1146 B.n447 B.n446 10.6151
R1147 B.n446 B.n113 10.6151
R1148 B.n442 B.n113 10.6151
R1149 B.n442 B.n441 10.6151
R1150 B.n441 B.n440 10.6151
R1151 B.n440 B.n115 10.6151
R1152 B.n436 B.n115 10.6151
R1153 B.n436 B.n435 10.6151
R1154 B.n435 B.n434 10.6151
R1155 B.n434 B.n117 10.6151
R1156 B.n430 B.n117 10.6151
R1157 B.n430 B.n429 10.6151
R1158 B.n429 B.n428 10.6151
R1159 B.n428 B.n119 10.6151
R1160 B.n424 B.n119 10.6151
R1161 B.n424 B.n423 10.6151
R1162 B.n423 B.n422 10.6151
R1163 B.n422 B.n121 10.6151
R1164 B.n418 B.n121 10.6151
R1165 B.n418 B.n417 10.6151
R1166 B.n417 B.n416 10.6151
R1167 B.n416 B.n123 10.6151
R1168 B.n412 B.n123 10.6151
R1169 B.n412 B.n411 10.6151
R1170 B.n199 B.n1 10.6151
R1171 B.n200 B.n199 10.6151
R1172 B.n200 B.n197 10.6151
R1173 B.n204 B.n197 10.6151
R1174 B.n205 B.n204 10.6151
R1175 B.n206 B.n205 10.6151
R1176 B.n206 B.n195 10.6151
R1177 B.n210 B.n195 10.6151
R1178 B.n211 B.n210 10.6151
R1179 B.n212 B.n211 10.6151
R1180 B.n212 B.n193 10.6151
R1181 B.n216 B.n193 10.6151
R1182 B.n217 B.n216 10.6151
R1183 B.n218 B.n217 10.6151
R1184 B.n218 B.n191 10.6151
R1185 B.n222 B.n191 10.6151
R1186 B.n223 B.n222 10.6151
R1187 B.n224 B.n223 10.6151
R1188 B.n224 B.n189 10.6151
R1189 B.n228 B.n189 10.6151
R1190 B.n229 B.n228 10.6151
R1191 B.n230 B.n229 10.6151
R1192 B.n230 B.n187 10.6151
R1193 B.n234 B.n187 10.6151
R1194 B.n235 B.n234 10.6151
R1195 B.n236 B.n235 10.6151
R1196 B.n236 B.n185 10.6151
R1197 B.n240 B.n185 10.6151
R1198 B.n241 B.n240 10.6151
R1199 B.n242 B.n241 10.6151
R1200 B.n242 B.n183 10.6151
R1201 B.n246 B.n183 10.6151
R1202 B.n247 B.n246 10.6151
R1203 B.n248 B.n247 10.6151
R1204 B.n248 B.n181 10.6151
R1205 B.n252 B.n181 10.6151
R1206 B.n253 B.n252 10.6151
R1207 B.n254 B.n253 10.6151
R1208 B.n254 B.n179 10.6151
R1209 B.n258 B.n179 10.6151
R1210 B.n259 B.n258 10.6151
R1211 B.n260 B.n259 10.6151
R1212 B.n260 B.n177 10.6151
R1213 B.n264 B.n177 10.6151
R1214 B.n265 B.n264 10.6151
R1215 B.n266 B.n175 10.6151
R1216 B.n270 B.n175 10.6151
R1217 B.n271 B.n270 10.6151
R1218 B.n272 B.n271 10.6151
R1219 B.n272 B.n173 10.6151
R1220 B.n276 B.n173 10.6151
R1221 B.n277 B.n276 10.6151
R1222 B.n278 B.n277 10.6151
R1223 B.n278 B.n171 10.6151
R1224 B.n282 B.n171 10.6151
R1225 B.n283 B.n282 10.6151
R1226 B.n284 B.n283 10.6151
R1227 B.n284 B.n169 10.6151
R1228 B.n288 B.n169 10.6151
R1229 B.n289 B.n288 10.6151
R1230 B.n290 B.n289 10.6151
R1231 B.n290 B.n167 10.6151
R1232 B.n294 B.n167 10.6151
R1233 B.n295 B.n294 10.6151
R1234 B.n296 B.n295 10.6151
R1235 B.n296 B.n165 10.6151
R1236 B.n300 B.n165 10.6151
R1237 B.n301 B.n300 10.6151
R1238 B.n302 B.n301 10.6151
R1239 B.n302 B.n163 10.6151
R1240 B.n306 B.n163 10.6151
R1241 B.n307 B.n306 10.6151
R1242 B.n308 B.n307 10.6151
R1243 B.n308 B.n161 10.6151
R1244 B.n312 B.n161 10.6151
R1245 B.n313 B.n312 10.6151
R1246 B.n314 B.n313 10.6151
R1247 B.n314 B.n159 10.6151
R1248 B.n318 B.n159 10.6151
R1249 B.n319 B.n318 10.6151
R1250 B.n320 B.n319 10.6151
R1251 B.n320 B.n157 10.6151
R1252 B.n324 B.n157 10.6151
R1253 B.n325 B.n324 10.6151
R1254 B.n326 B.n325 10.6151
R1255 B.n326 B.n155 10.6151
R1256 B.n330 B.n155 10.6151
R1257 B.n333 B.n332 10.6151
R1258 B.n333 B.n151 10.6151
R1259 B.n337 B.n151 10.6151
R1260 B.n338 B.n337 10.6151
R1261 B.n339 B.n338 10.6151
R1262 B.n339 B.n149 10.6151
R1263 B.n343 B.n149 10.6151
R1264 B.n344 B.n343 10.6151
R1265 B.n346 B.n145 10.6151
R1266 B.n350 B.n145 10.6151
R1267 B.n351 B.n350 10.6151
R1268 B.n352 B.n351 10.6151
R1269 B.n352 B.n143 10.6151
R1270 B.n356 B.n143 10.6151
R1271 B.n357 B.n356 10.6151
R1272 B.n358 B.n357 10.6151
R1273 B.n358 B.n141 10.6151
R1274 B.n362 B.n141 10.6151
R1275 B.n363 B.n362 10.6151
R1276 B.n364 B.n363 10.6151
R1277 B.n364 B.n139 10.6151
R1278 B.n368 B.n139 10.6151
R1279 B.n369 B.n368 10.6151
R1280 B.n370 B.n369 10.6151
R1281 B.n370 B.n137 10.6151
R1282 B.n374 B.n137 10.6151
R1283 B.n375 B.n374 10.6151
R1284 B.n376 B.n375 10.6151
R1285 B.n376 B.n135 10.6151
R1286 B.n380 B.n135 10.6151
R1287 B.n381 B.n380 10.6151
R1288 B.n382 B.n381 10.6151
R1289 B.n382 B.n133 10.6151
R1290 B.n386 B.n133 10.6151
R1291 B.n387 B.n386 10.6151
R1292 B.n388 B.n387 10.6151
R1293 B.n388 B.n131 10.6151
R1294 B.n392 B.n131 10.6151
R1295 B.n393 B.n392 10.6151
R1296 B.n394 B.n393 10.6151
R1297 B.n394 B.n129 10.6151
R1298 B.n398 B.n129 10.6151
R1299 B.n399 B.n398 10.6151
R1300 B.n400 B.n399 10.6151
R1301 B.n400 B.n127 10.6151
R1302 B.n404 B.n127 10.6151
R1303 B.n405 B.n404 10.6151
R1304 B.n406 B.n405 10.6151
R1305 B.n406 B.n125 10.6151
R1306 B.n410 B.n125 10.6151
R1307 B.n765 B.n0 8.11757
R1308 B.n765 B.n1 8.11757
R1309 B.n629 B.n50 6.5566
R1310 B.n617 B.n616 6.5566
R1311 B.n332 B.n331 6.5566
R1312 B.n345 B.n344 6.5566
R1313 B.n50 B.n46 4.05904
R1314 B.n616 B.n615 4.05904
R1315 B.n331 B.n330 4.05904
R1316 B.n346 B.n345 4.05904
R1317 VP.n17 VP.t7 196.847
R1318 VP.n42 VP.n9 180.385
R1319 VP.n74 VP.n73 180.385
R1320 VP.n41 VP.n40 180.385
R1321 VP.n9 VP.t4 161.405
R1322 VP.n51 VP.t2 161.405
R1323 VP.n58 VP.t6 161.405
R1324 VP.n65 VP.t5 161.405
R1325 VP.n73 VP.t1 161.405
R1326 VP.n40 VP.t0 161.405
R1327 VP.n32 VP.t3 161.405
R1328 VP.n25 VP.t8 161.405
R1329 VP.n18 VP.t9 161.405
R1330 VP.n19 VP.n16 161.3
R1331 VP.n21 VP.n20 161.3
R1332 VP.n22 VP.n15 161.3
R1333 VP.n24 VP.n23 161.3
R1334 VP.n26 VP.n14 161.3
R1335 VP.n28 VP.n27 161.3
R1336 VP.n29 VP.n13 161.3
R1337 VP.n31 VP.n30 161.3
R1338 VP.n33 VP.n12 161.3
R1339 VP.n35 VP.n34 161.3
R1340 VP.n36 VP.n11 161.3
R1341 VP.n38 VP.n37 161.3
R1342 VP.n39 VP.n10 161.3
R1343 VP.n72 VP.n0 161.3
R1344 VP.n71 VP.n70 161.3
R1345 VP.n69 VP.n1 161.3
R1346 VP.n68 VP.n67 161.3
R1347 VP.n66 VP.n2 161.3
R1348 VP.n64 VP.n63 161.3
R1349 VP.n62 VP.n3 161.3
R1350 VP.n61 VP.n60 161.3
R1351 VP.n59 VP.n4 161.3
R1352 VP.n57 VP.n56 161.3
R1353 VP.n55 VP.n5 161.3
R1354 VP.n54 VP.n53 161.3
R1355 VP.n52 VP.n6 161.3
R1356 VP.n50 VP.n49 161.3
R1357 VP.n48 VP.n7 161.3
R1358 VP.n47 VP.n46 161.3
R1359 VP.n45 VP.n8 161.3
R1360 VP.n44 VP.n43 161.3
R1361 VP.n53 VP.n5 56.0336
R1362 VP.n60 VP.n3 56.0336
R1363 VP.n27 VP.n13 56.0336
R1364 VP.n20 VP.n15 56.0336
R1365 VP.n42 VP.n41 49.2732
R1366 VP.n18 VP.n17 48.2603
R1367 VP.n46 VP.n45 42.4359
R1368 VP.n71 VP.n1 42.4359
R1369 VP.n38 VP.n11 42.4359
R1370 VP.n46 VP.n7 38.5509
R1371 VP.n67 VP.n1 38.5509
R1372 VP.n34 VP.n11 38.5509
R1373 VP.n53 VP.n52 24.9531
R1374 VP.n64 VP.n3 24.9531
R1375 VP.n31 VP.n13 24.9531
R1376 VP.n20 VP.n19 24.9531
R1377 VP.n45 VP.n44 24.4675
R1378 VP.n50 VP.n7 24.4675
R1379 VP.n57 VP.n5 24.4675
R1380 VP.n60 VP.n59 24.4675
R1381 VP.n67 VP.n66 24.4675
R1382 VP.n72 VP.n71 24.4675
R1383 VP.n39 VP.n38 24.4675
R1384 VP.n34 VP.n33 24.4675
R1385 VP.n24 VP.n15 24.4675
R1386 VP.n27 VP.n26 24.4675
R1387 VP.n52 VP.n51 21.0421
R1388 VP.n65 VP.n64 21.0421
R1389 VP.n32 VP.n31 21.0421
R1390 VP.n19 VP.n18 21.0421
R1391 VP.n58 VP.n57 12.234
R1392 VP.n59 VP.n58 12.234
R1393 VP.n25 VP.n24 12.234
R1394 VP.n26 VP.n25 12.234
R1395 VP.n17 VP.n16 12.1797
R1396 VP.n44 VP.n9 5.38324
R1397 VP.n73 VP.n72 5.38324
R1398 VP.n40 VP.n39 5.38324
R1399 VP.n51 VP.n50 3.42588
R1400 VP.n66 VP.n65 3.42588
R1401 VP.n33 VP.n32 3.42588
R1402 VP.n21 VP.n16 0.189894
R1403 VP.n22 VP.n21 0.189894
R1404 VP.n23 VP.n22 0.189894
R1405 VP.n23 VP.n14 0.189894
R1406 VP.n28 VP.n14 0.189894
R1407 VP.n29 VP.n28 0.189894
R1408 VP.n30 VP.n29 0.189894
R1409 VP.n30 VP.n12 0.189894
R1410 VP.n35 VP.n12 0.189894
R1411 VP.n36 VP.n35 0.189894
R1412 VP.n37 VP.n36 0.189894
R1413 VP.n37 VP.n10 0.189894
R1414 VP.n41 VP.n10 0.189894
R1415 VP.n43 VP.n42 0.189894
R1416 VP.n43 VP.n8 0.189894
R1417 VP.n47 VP.n8 0.189894
R1418 VP.n48 VP.n47 0.189894
R1419 VP.n49 VP.n48 0.189894
R1420 VP.n49 VP.n6 0.189894
R1421 VP.n54 VP.n6 0.189894
R1422 VP.n55 VP.n54 0.189894
R1423 VP.n56 VP.n55 0.189894
R1424 VP.n56 VP.n4 0.189894
R1425 VP.n61 VP.n4 0.189894
R1426 VP.n62 VP.n61 0.189894
R1427 VP.n63 VP.n62 0.189894
R1428 VP.n63 VP.n2 0.189894
R1429 VP.n68 VP.n2 0.189894
R1430 VP.n69 VP.n68 0.189894
R1431 VP.n70 VP.n69 0.189894
R1432 VP.n70 VP.n0 0.189894
R1433 VP.n74 VP.n0 0.189894
R1434 VP VP.n74 0.0516364
R1435 VDD1.n1 VDD1.t2 76.169
R1436 VDD1.n3 VDD1.t5 76.1689
R1437 VDD1.n5 VDD1.n4 73.0202
R1438 VDD1.n1 VDD1.n0 71.6663
R1439 VDD1.n7 VDD1.n6 71.6661
R1440 VDD1.n3 VDD1.n2 71.6661
R1441 VDD1.n7 VDD1.n5 44.8457
R1442 VDD1.n6 VDD1.t6 2.62399
R1443 VDD1.n6 VDD1.t9 2.62399
R1444 VDD1.n0 VDD1.t0 2.62399
R1445 VDD1.n0 VDD1.t1 2.62399
R1446 VDD1.n4 VDD1.t4 2.62399
R1447 VDD1.n4 VDD1.t8 2.62399
R1448 VDD1.n2 VDD1.t7 2.62399
R1449 VDD1.n2 VDD1.t3 2.62399
R1450 VDD1 VDD1.n7 1.35179
R1451 VDD1 VDD1.n1 0.528517
R1452 VDD1.n5 VDD1.n3 0.414982
C0 VDD1 VP 10.489599f
C1 VP VN 7.36228f
C2 VDD2 VTAIL 10.7923f
C3 VDD2 w_n3586_n3446# 2.63319f
C4 w_n3586_n3446# VTAIL 3.16824f
C5 VDD2 B 2.30231f
C6 VDD2 VDD1 1.68566f
C7 VDD2 VN 10.1572f
C8 VTAIL B 3.47566f
C9 w_n3586_n3446# B 9.39498f
C10 VDD2 VP 0.487861f
C11 VDD1 VTAIL 10.7476f
C12 VDD1 w_n3586_n3446# 2.52852f
C13 VTAIL VN 10.4727f
C14 w_n3586_n3446# VN 7.44433f
C15 VTAIL VP 10.4871f
C16 w_n3586_n3446# VP 7.9089f
C17 VDD1 B 2.2136f
C18 B VN 1.09709f
C19 B VP 1.87414f
C20 VDD1 VN 0.151509f
C21 VDD2 VSUBS 1.873185f
C22 VDD1 VSUBS 1.653886f
C23 VTAIL VSUBS 1.13801f
C24 VN VSUBS 6.47797f
C25 VP VSUBS 3.282002f
C26 B VSUBS 4.468581f
C27 w_n3586_n3446# VSUBS 0.152032p
C28 VDD1.t2 VSUBS 2.75711f
C29 VDD1.t0 VSUBS 0.268213f
C30 VDD1.t1 VSUBS 0.268213f
C31 VDD1.n0 VSUBS 2.09645f
C32 VDD1.n1 VSUBS 1.51092f
C33 VDD1.t5 VSUBS 2.7571f
C34 VDD1.t7 VSUBS 0.268213f
C35 VDD1.t3 VSUBS 0.268213f
C36 VDD1.n2 VSUBS 2.09645f
C37 VDD1.n3 VSUBS 1.50245f
C38 VDD1.t4 VSUBS 0.268213f
C39 VDD1.t8 VSUBS 0.268213f
C40 VDD1.n4 VSUBS 2.1117f
C41 VDD1.n5 VSUBS 3.1906f
C42 VDD1.t6 VSUBS 0.268213f
C43 VDD1.t9 VSUBS 0.268213f
C44 VDD1.n6 VSUBS 2.09644f
C45 VDD1.n7 VSUBS 3.46919f
C46 VP.n0 VSUBS 0.034333f
C47 VP.t1 VSUBS 2.14613f
C48 VP.n1 VSUBS 0.027932f
C49 VP.n2 VSUBS 0.034333f
C50 VP.t5 VSUBS 2.14613f
C51 VP.n3 VSUBS 0.040994f
C52 VP.n4 VSUBS 0.034333f
C53 VP.t6 VSUBS 2.14613f
C54 VP.n5 VSUBS 0.058647f
C55 VP.n6 VSUBS 0.034333f
C56 VP.t2 VSUBS 2.14613f
C57 VP.n7 VSUBS 0.068834f
C58 VP.n8 VSUBS 0.034333f
C59 VP.t4 VSUBS 2.14613f
C60 VP.n9 VSUBS 0.849955f
C61 VP.n10 VSUBS 0.034333f
C62 VP.t0 VSUBS 2.14613f
C63 VP.n11 VSUBS 0.027932f
C64 VP.n12 VSUBS 0.034333f
C65 VP.t3 VSUBS 2.14613f
C66 VP.n13 VSUBS 0.040994f
C67 VP.n14 VSUBS 0.034333f
C68 VP.t8 VSUBS 2.14613f
C69 VP.n15 VSUBS 0.058647f
C70 VP.n16 VSUBS 0.255061f
C71 VP.t9 VSUBS 2.14613f
C72 VP.t7 VSUBS 2.31424f
C73 VP.n17 VSUBS 0.840349f
C74 VP.n18 VSUBS 0.855826f
C75 VP.n19 VSUBS 0.060167f
C76 VP.n20 VSUBS 0.040994f
C77 VP.n21 VSUBS 0.034333f
C78 VP.n22 VSUBS 0.034333f
C79 VP.n23 VSUBS 0.034333f
C80 VP.n24 VSUBS 0.048193f
C81 VP.n25 VSUBS 0.766746f
C82 VP.n26 VSUBS 0.048193f
C83 VP.n27 VSUBS 0.058647f
C84 VP.n28 VSUBS 0.034333f
C85 VP.n29 VSUBS 0.034333f
C86 VP.n30 VSUBS 0.034333f
C87 VP.n31 VSUBS 0.060167f
C88 VP.n32 VSUBS 0.766746f
C89 VP.n33 VSUBS 0.03682f
C90 VP.n34 VSUBS 0.068834f
C91 VP.n35 VSUBS 0.034333f
C92 VP.n36 VSUBS 0.034333f
C93 VP.n37 VSUBS 0.034333f
C94 VP.n38 VSUBS 0.067464f
C95 VP.n39 VSUBS 0.039347f
C96 VP.n40 VSUBS 0.849955f
C97 VP.n41 VSUBS 1.83564f
C98 VP.n42 VSUBS 1.86069f
C99 VP.n43 VSUBS 0.034333f
C100 VP.n44 VSUBS 0.039347f
C101 VP.n45 VSUBS 0.067464f
C102 VP.n46 VSUBS 0.027932f
C103 VP.n47 VSUBS 0.034333f
C104 VP.n48 VSUBS 0.034333f
C105 VP.n49 VSUBS 0.034333f
C106 VP.n50 VSUBS 0.03682f
C107 VP.n51 VSUBS 0.766746f
C108 VP.n52 VSUBS 0.060167f
C109 VP.n53 VSUBS 0.040994f
C110 VP.n54 VSUBS 0.034333f
C111 VP.n55 VSUBS 0.034333f
C112 VP.n56 VSUBS 0.034333f
C113 VP.n57 VSUBS 0.048193f
C114 VP.n58 VSUBS 0.766746f
C115 VP.n59 VSUBS 0.048193f
C116 VP.n60 VSUBS 0.058647f
C117 VP.n61 VSUBS 0.034333f
C118 VP.n62 VSUBS 0.034333f
C119 VP.n63 VSUBS 0.034333f
C120 VP.n64 VSUBS 0.060167f
C121 VP.n65 VSUBS 0.766746f
C122 VP.n66 VSUBS 0.03682f
C123 VP.n67 VSUBS 0.068834f
C124 VP.n68 VSUBS 0.034333f
C125 VP.n69 VSUBS 0.034333f
C126 VP.n70 VSUBS 0.034333f
C127 VP.n71 VSUBS 0.067464f
C128 VP.n72 VSUBS 0.039347f
C129 VP.n73 VSUBS 0.849955f
C130 VP.n74 VSUBS 0.036452f
C131 B.n0 VSUBS 0.007698f
C132 B.n1 VSUBS 0.007698f
C133 B.n2 VSUBS 0.011385f
C134 B.n3 VSUBS 0.008724f
C135 B.n4 VSUBS 0.008724f
C136 B.n5 VSUBS 0.008724f
C137 B.n6 VSUBS 0.008724f
C138 B.n7 VSUBS 0.008724f
C139 B.n8 VSUBS 0.008724f
C140 B.n9 VSUBS 0.008724f
C141 B.n10 VSUBS 0.008724f
C142 B.n11 VSUBS 0.008724f
C143 B.n12 VSUBS 0.008724f
C144 B.n13 VSUBS 0.008724f
C145 B.n14 VSUBS 0.008724f
C146 B.n15 VSUBS 0.008724f
C147 B.n16 VSUBS 0.008724f
C148 B.n17 VSUBS 0.008724f
C149 B.n18 VSUBS 0.008724f
C150 B.n19 VSUBS 0.008724f
C151 B.n20 VSUBS 0.008724f
C152 B.n21 VSUBS 0.008724f
C153 B.n22 VSUBS 0.008724f
C154 B.n23 VSUBS 0.008724f
C155 B.n24 VSUBS 0.008724f
C156 B.n25 VSUBS 0.02141f
C157 B.n26 VSUBS 0.008724f
C158 B.n27 VSUBS 0.008724f
C159 B.n28 VSUBS 0.008724f
C160 B.n29 VSUBS 0.008724f
C161 B.n30 VSUBS 0.008724f
C162 B.n31 VSUBS 0.008724f
C163 B.n32 VSUBS 0.008724f
C164 B.n33 VSUBS 0.008724f
C165 B.n34 VSUBS 0.008724f
C166 B.n35 VSUBS 0.008724f
C167 B.n36 VSUBS 0.008724f
C168 B.n37 VSUBS 0.008724f
C169 B.n38 VSUBS 0.008724f
C170 B.n39 VSUBS 0.008724f
C171 B.n40 VSUBS 0.008724f
C172 B.n41 VSUBS 0.008724f
C173 B.n42 VSUBS 0.008724f
C174 B.n43 VSUBS 0.008724f
C175 B.n44 VSUBS 0.008724f
C176 B.n45 VSUBS 0.008724f
C177 B.n46 VSUBS 0.00603f
C178 B.n47 VSUBS 0.008724f
C179 B.t1 VSUBS 0.50494f
C180 B.t2 VSUBS 0.525274f
C181 B.t0 VSUBS 1.26706f
C182 B.n48 VSUBS 0.249668f
C183 B.n49 VSUBS 0.085638f
C184 B.n50 VSUBS 0.020213f
C185 B.n51 VSUBS 0.008724f
C186 B.n52 VSUBS 0.008724f
C187 B.n53 VSUBS 0.008724f
C188 B.n54 VSUBS 0.008724f
C189 B.t7 VSUBS 0.50493f
C190 B.t8 VSUBS 0.525264f
C191 B.t6 VSUBS 1.26706f
C192 B.n55 VSUBS 0.249678f
C193 B.n56 VSUBS 0.085649f
C194 B.n57 VSUBS 0.008724f
C195 B.n58 VSUBS 0.008724f
C196 B.n59 VSUBS 0.008724f
C197 B.n60 VSUBS 0.008724f
C198 B.n61 VSUBS 0.008724f
C199 B.n62 VSUBS 0.008724f
C200 B.n63 VSUBS 0.008724f
C201 B.n64 VSUBS 0.008724f
C202 B.n65 VSUBS 0.008724f
C203 B.n66 VSUBS 0.008724f
C204 B.n67 VSUBS 0.008724f
C205 B.n68 VSUBS 0.008724f
C206 B.n69 VSUBS 0.008724f
C207 B.n70 VSUBS 0.008724f
C208 B.n71 VSUBS 0.008724f
C209 B.n72 VSUBS 0.008724f
C210 B.n73 VSUBS 0.008724f
C211 B.n74 VSUBS 0.008724f
C212 B.n75 VSUBS 0.008724f
C213 B.n76 VSUBS 0.008724f
C214 B.n77 VSUBS 0.02141f
C215 B.n78 VSUBS 0.008724f
C216 B.n79 VSUBS 0.008724f
C217 B.n80 VSUBS 0.008724f
C218 B.n81 VSUBS 0.008724f
C219 B.n82 VSUBS 0.008724f
C220 B.n83 VSUBS 0.008724f
C221 B.n84 VSUBS 0.008724f
C222 B.n85 VSUBS 0.008724f
C223 B.n86 VSUBS 0.008724f
C224 B.n87 VSUBS 0.008724f
C225 B.n88 VSUBS 0.008724f
C226 B.n89 VSUBS 0.008724f
C227 B.n90 VSUBS 0.008724f
C228 B.n91 VSUBS 0.008724f
C229 B.n92 VSUBS 0.008724f
C230 B.n93 VSUBS 0.008724f
C231 B.n94 VSUBS 0.008724f
C232 B.n95 VSUBS 0.008724f
C233 B.n96 VSUBS 0.008724f
C234 B.n97 VSUBS 0.008724f
C235 B.n98 VSUBS 0.008724f
C236 B.n99 VSUBS 0.008724f
C237 B.n100 VSUBS 0.008724f
C238 B.n101 VSUBS 0.008724f
C239 B.n102 VSUBS 0.008724f
C240 B.n103 VSUBS 0.008724f
C241 B.n104 VSUBS 0.008724f
C242 B.n105 VSUBS 0.008724f
C243 B.n106 VSUBS 0.008724f
C244 B.n107 VSUBS 0.008724f
C245 B.n108 VSUBS 0.008724f
C246 B.n109 VSUBS 0.008724f
C247 B.n110 VSUBS 0.008724f
C248 B.n111 VSUBS 0.008724f
C249 B.n112 VSUBS 0.008724f
C250 B.n113 VSUBS 0.008724f
C251 B.n114 VSUBS 0.008724f
C252 B.n115 VSUBS 0.008724f
C253 B.n116 VSUBS 0.008724f
C254 B.n117 VSUBS 0.008724f
C255 B.n118 VSUBS 0.008724f
C256 B.n119 VSUBS 0.008724f
C257 B.n120 VSUBS 0.008724f
C258 B.n121 VSUBS 0.008724f
C259 B.n122 VSUBS 0.008724f
C260 B.n123 VSUBS 0.008724f
C261 B.n124 VSUBS 0.020416f
C262 B.n125 VSUBS 0.008724f
C263 B.n126 VSUBS 0.008724f
C264 B.n127 VSUBS 0.008724f
C265 B.n128 VSUBS 0.008724f
C266 B.n129 VSUBS 0.008724f
C267 B.n130 VSUBS 0.008724f
C268 B.n131 VSUBS 0.008724f
C269 B.n132 VSUBS 0.008724f
C270 B.n133 VSUBS 0.008724f
C271 B.n134 VSUBS 0.008724f
C272 B.n135 VSUBS 0.008724f
C273 B.n136 VSUBS 0.008724f
C274 B.n137 VSUBS 0.008724f
C275 B.n138 VSUBS 0.008724f
C276 B.n139 VSUBS 0.008724f
C277 B.n140 VSUBS 0.008724f
C278 B.n141 VSUBS 0.008724f
C279 B.n142 VSUBS 0.008724f
C280 B.n143 VSUBS 0.008724f
C281 B.n144 VSUBS 0.008724f
C282 B.n145 VSUBS 0.008724f
C283 B.n146 VSUBS 0.008724f
C284 B.t5 VSUBS 0.50493f
C285 B.t4 VSUBS 0.525264f
C286 B.t3 VSUBS 1.26706f
C287 B.n147 VSUBS 0.249678f
C288 B.n148 VSUBS 0.085649f
C289 B.n149 VSUBS 0.008724f
C290 B.n150 VSUBS 0.008724f
C291 B.n151 VSUBS 0.008724f
C292 B.n152 VSUBS 0.008724f
C293 B.t11 VSUBS 0.50494f
C294 B.t10 VSUBS 0.525274f
C295 B.t9 VSUBS 1.26706f
C296 B.n153 VSUBS 0.249668f
C297 B.n154 VSUBS 0.085638f
C298 B.n155 VSUBS 0.008724f
C299 B.n156 VSUBS 0.008724f
C300 B.n157 VSUBS 0.008724f
C301 B.n158 VSUBS 0.008724f
C302 B.n159 VSUBS 0.008724f
C303 B.n160 VSUBS 0.008724f
C304 B.n161 VSUBS 0.008724f
C305 B.n162 VSUBS 0.008724f
C306 B.n163 VSUBS 0.008724f
C307 B.n164 VSUBS 0.008724f
C308 B.n165 VSUBS 0.008724f
C309 B.n166 VSUBS 0.008724f
C310 B.n167 VSUBS 0.008724f
C311 B.n168 VSUBS 0.008724f
C312 B.n169 VSUBS 0.008724f
C313 B.n170 VSUBS 0.008724f
C314 B.n171 VSUBS 0.008724f
C315 B.n172 VSUBS 0.008724f
C316 B.n173 VSUBS 0.008724f
C317 B.n174 VSUBS 0.008724f
C318 B.n175 VSUBS 0.008724f
C319 B.n176 VSUBS 0.020416f
C320 B.n177 VSUBS 0.008724f
C321 B.n178 VSUBS 0.008724f
C322 B.n179 VSUBS 0.008724f
C323 B.n180 VSUBS 0.008724f
C324 B.n181 VSUBS 0.008724f
C325 B.n182 VSUBS 0.008724f
C326 B.n183 VSUBS 0.008724f
C327 B.n184 VSUBS 0.008724f
C328 B.n185 VSUBS 0.008724f
C329 B.n186 VSUBS 0.008724f
C330 B.n187 VSUBS 0.008724f
C331 B.n188 VSUBS 0.008724f
C332 B.n189 VSUBS 0.008724f
C333 B.n190 VSUBS 0.008724f
C334 B.n191 VSUBS 0.008724f
C335 B.n192 VSUBS 0.008724f
C336 B.n193 VSUBS 0.008724f
C337 B.n194 VSUBS 0.008724f
C338 B.n195 VSUBS 0.008724f
C339 B.n196 VSUBS 0.008724f
C340 B.n197 VSUBS 0.008724f
C341 B.n198 VSUBS 0.008724f
C342 B.n199 VSUBS 0.008724f
C343 B.n200 VSUBS 0.008724f
C344 B.n201 VSUBS 0.008724f
C345 B.n202 VSUBS 0.008724f
C346 B.n203 VSUBS 0.008724f
C347 B.n204 VSUBS 0.008724f
C348 B.n205 VSUBS 0.008724f
C349 B.n206 VSUBS 0.008724f
C350 B.n207 VSUBS 0.008724f
C351 B.n208 VSUBS 0.008724f
C352 B.n209 VSUBS 0.008724f
C353 B.n210 VSUBS 0.008724f
C354 B.n211 VSUBS 0.008724f
C355 B.n212 VSUBS 0.008724f
C356 B.n213 VSUBS 0.008724f
C357 B.n214 VSUBS 0.008724f
C358 B.n215 VSUBS 0.008724f
C359 B.n216 VSUBS 0.008724f
C360 B.n217 VSUBS 0.008724f
C361 B.n218 VSUBS 0.008724f
C362 B.n219 VSUBS 0.008724f
C363 B.n220 VSUBS 0.008724f
C364 B.n221 VSUBS 0.008724f
C365 B.n222 VSUBS 0.008724f
C366 B.n223 VSUBS 0.008724f
C367 B.n224 VSUBS 0.008724f
C368 B.n225 VSUBS 0.008724f
C369 B.n226 VSUBS 0.008724f
C370 B.n227 VSUBS 0.008724f
C371 B.n228 VSUBS 0.008724f
C372 B.n229 VSUBS 0.008724f
C373 B.n230 VSUBS 0.008724f
C374 B.n231 VSUBS 0.008724f
C375 B.n232 VSUBS 0.008724f
C376 B.n233 VSUBS 0.008724f
C377 B.n234 VSUBS 0.008724f
C378 B.n235 VSUBS 0.008724f
C379 B.n236 VSUBS 0.008724f
C380 B.n237 VSUBS 0.008724f
C381 B.n238 VSUBS 0.008724f
C382 B.n239 VSUBS 0.008724f
C383 B.n240 VSUBS 0.008724f
C384 B.n241 VSUBS 0.008724f
C385 B.n242 VSUBS 0.008724f
C386 B.n243 VSUBS 0.008724f
C387 B.n244 VSUBS 0.008724f
C388 B.n245 VSUBS 0.008724f
C389 B.n246 VSUBS 0.008724f
C390 B.n247 VSUBS 0.008724f
C391 B.n248 VSUBS 0.008724f
C392 B.n249 VSUBS 0.008724f
C393 B.n250 VSUBS 0.008724f
C394 B.n251 VSUBS 0.008724f
C395 B.n252 VSUBS 0.008724f
C396 B.n253 VSUBS 0.008724f
C397 B.n254 VSUBS 0.008724f
C398 B.n255 VSUBS 0.008724f
C399 B.n256 VSUBS 0.008724f
C400 B.n257 VSUBS 0.008724f
C401 B.n258 VSUBS 0.008724f
C402 B.n259 VSUBS 0.008724f
C403 B.n260 VSUBS 0.008724f
C404 B.n261 VSUBS 0.008724f
C405 B.n262 VSUBS 0.008724f
C406 B.n263 VSUBS 0.008724f
C407 B.n264 VSUBS 0.008724f
C408 B.n265 VSUBS 0.020416f
C409 B.n266 VSUBS 0.02141f
C410 B.n267 VSUBS 0.02141f
C411 B.n268 VSUBS 0.008724f
C412 B.n269 VSUBS 0.008724f
C413 B.n270 VSUBS 0.008724f
C414 B.n271 VSUBS 0.008724f
C415 B.n272 VSUBS 0.008724f
C416 B.n273 VSUBS 0.008724f
C417 B.n274 VSUBS 0.008724f
C418 B.n275 VSUBS 0.008724f
C419 B.n276 VSUBS 0.008724f
C420 B.n277 VSUBS 0.008724f
C421 B.n278 VSUBS 0.008724f
C422 B.n279 VSUBS 0.008724f
C423 B.n280 VSUBS 0.008724f
C424 B.n281 VSUBS 0.008724f
C425 B.n282 VSUBS 0.008724f
C426 B.n283 VSUBS 0.008724f
C427 B.n284 VSUBS 0.008724f
C428 B.n285 VSUBS 0.008724f
C429 B.n286 VSUBS 0.008724f
C430 B.n287 VSUBS 0.008724f
C431 B.n288 VSUBS 0.008724f
C432 B.n289 VSUBS 0.008724f
C433 B.n290 VSUBS 0.008724f
C434 B.n291 VSUBS 0.008724f
C435 B.n292 VSUBS 0.008724f
C436 B.n293 VSUBS 0.008724f
C437 B.n294 VSUBS 0.008724f
C438 B.n295 VSUBS 0.008724f
C439 B.n296 VSUBS 0.008724f
C440 B.n297 VSUBS 0.008724f
C441 B.n298 VSUBS 0.008724f
C442 B.n299 VSUBS 0.008724f
C443 B.n300 VSUBS 0.008724f
C444 B.n301 VSUBS 0.008724f
C445 B.n302 VSUBS 0.008724f
C446 B.n303 VSUBS 0.008724f
C447 B.n304 VSUBS 0.008724f
C448 B.n305 VSUBS 0.008724f
C449 B.n306 VSUBS 0.008724f
C450 B.n307 VSUBS 0.008724f
C451 B.n308 VSUBS 0.008724f
C452 B.n309 VSUBS 0.008724f
C453 B.n310 VSUBS 0.008724f
C454 B.n311 VSUBS 0.008724f
C455 B.n312 VSUBS 0.008724f
C456 B.n313 VSUBS 0.008724f
C457 B.n314 VSUBS 0.008724f
C458 B.n315 VSUBS 0.008724f
C459 B.n316 VSUBS 0.008724f
C460 B.n317 VSUBS 0.008724f
C461 B.n318 VSUBS 0.008724f
C462 B.n319 VSUBS 0.008724f
C463 B.n320 VSUBS 0.008724f
C464 B.n321 VSUBS 0.008724f
C465 B.n322 VSUBS 0.008724f
C466 B.n323 VSUBS 0.008724f
C467 B.n324 VSUBS 0.008724f
C468 B.n325 VSUBS 0.008724f
C469 B.n326 VSUBS 0.008724f
C470 B.n327 VSUBS 0.008724f
C471 B.n328 VSUBS 0.008724f
C472 B.n329 VSUBS 0.008724f
C473 B.n330 VSUBS 0.00603f
C474 B.n331 VSUBS 0.020213f
C475 B.n332 VSUBS 0.007056f
C476 B.n333 VSUBS 0.008724f
C477 B.n334 VSUBS 0.008724f
C478 B.n335 VSUBS 0.008724f
C479 B.n336 VSUBS 0.008724f
C480 B.n337 VSUBS 0.008724f
C481 B.n338 VSUBS 0.008724f
C482 B.n339 VSUBS 0.008724f
C483 B.n340 VSUBS 0.008724f
C484 B.n341 VSUBS 0.008724f
C485 B.n342 VSUBS 0.008724f
C486 B.n343 VSUBS 0.008724f
C487 B.n344 VSUBS 0.007056f
C488 B.n345 VSUBS 0.020213f
C489 B.n346 VSUBS 0.00603f
C490 B.n347 VSUBS 0.008724f
C491 B.n348 VSUBS 0.008724f
C492 B.n349 VSUBS 0.008724f
C493 B.n350 VSUBS 0.008724f
C494 B.n351 VSUBS 0.008724f
C495 B.n352 VSUBS 0.008724f
C496 B.n353 VSUBS 0.008724f
C497 B.n354 VSUBS 0.008724f
C498 B.n355 VSUBS 0.008724f
C499 B.n356 VSUBS 0.008724f
C500 B.n357 VSUBS 0.008724f
C501 B.n358 VSUBS 0.008724f
C502 B.n359 VSUBS 0.008724f
C503 B.n360 VSUBS 0.008724f
C504 B.n361 VSUBS 0.008724f
C505 B.n362 VSUBS 0.008724f
C506 B.n363 VSUBS 0.008724f
C507 B.n364 VSUBS 0.008724f
C508 B.n365 VSUBS 0.008724f
C509 B.n366 VSUBS 0.008724f
C510 B.n367 VSUBS 0.008724f
C511 B.n368 VSUBS 0.008724f
C512 B.n369 VSUBS 0.008724f
C513 B.n370 VSUBS 0.008724f
C514 B.n371 VSUBS 0.008724f
C515 B.n372 VSUBS 0.008724f
C516 B.n373 VSUBS 0.008724f
C517 B.n374 VSUBS 0.008724f
C518 B.n375 VSUBS 0.008724f
C519 B.n376 VSUBS 0.008724f
C520 B.n377 VSUBS 0.008724f
C521 B.n378 VSUBS 0.008724f
C522 B.n379 VSUBS 0.008724f
C523 B.n380 VSUBS 0.008724f
C524 B.n381 VSUBS 0.008724f
C525 B.n382 VSUBS 0.008724f
C526 B.n383 VSUBS 0.008724f
C527 B.n384 VSUBS 0.008724f
C528 B.n385 VSUBS 0.008724f
C529 B.n386 VSUBS 0.008724f
C530 B.n387 VSUBS 0.008724f
C531 B.n388 VSUBS 0.008724f
C532 B.n389 VSUBS 0.008724f
C533 B.n390 VSUBS 0.008724f
C534 B.n391 VSUBS 0.008724f
C535 B.n392 VSUBS 0.008724f
C536 B.n393 VSUBS 0.008724f
C537 B.n394 VSUBS 0.008724f
C538 B.n395 VSUBS 0.008724f
C539 B.n396 VSUBS 0.008724f
C540 B.n397 VSUBS 0.008724f
C541 B.n398 VSUBS 0.008724f
C542 B.n399 VSUBS 0.008724f
C543 B.n400 VSUBS 0.008724f
C544 B.n401 VSUBS 0.008724f
C545 B.n402 VSUBS 0.008724f
C546 B.n403 VSUBS 0.008724f
C547 B.n404 VSUBS 0.008724f
C548 B.n405 VSUBS 0.008724f
C549 B.n406 VSUBS 0.008724f
C550 B.n407 VSUBS 0.008724f
C551 B.n408 VSUBS 0.008724f
C552 B.n409 VSUBS 0.02141f
C553 B.n410 VSUBS 0.020416f
C554 B.n411 VSUBS 0.02141f
C555 B.n412 VSUBS 0.008724f
C556 B.n413 VSUBS 0.008724f
C557 B.n414 VSUBS 0.008724f
C558 B.n415 VSUBS 0.008724f
C559 B.n416 VSUBS 0.008724f
C560 B.n417 VSUBS 0.008724f
C561 B.n418 VSUBS 0.008724f
C562 B.n419 VSUBS 0.008724f
C563 B.n420 VSUBS 0.008724f
C564 B.n421 VSUBS 0.008724f
C565 B.n422 VSUBS 0.008724f
C566 B.n423 VSUBS 0.008724f
C567 B.n424 VSUBS 0.008724f
C568 B.n425 VSUBS 0.008724f
C569 B.n426 VSUBS 0.008724f
C570 B.n427 VSUBS 0.008724f
C571 B.n428 VSUBS 0.008724f
C572 B.n429 VSUBS 0.008724f
C573 B.n430 VSUBS 0.008724f
C574 B.n431 VSUBS 0.008724f
C575 B.n432 VSUBS 0.008724f
C576 B.n433 VSUBS 0.008724f
C577 B.n434 VSUBS 0.008724f
C578 B.n435 VSUBS 0.008724f
C579 B.n436 VSUBS 0.008724f
C580 B.n437 VSUBS 0.008724f
C581 B.n438 VSUBS 0.008724f
C582 B.n439 VSUBS 0.008724f
C583 B.n440 VSUBS 0.008724f
C584 B.n441 VSUBS 0.008724f
C585 B.n442 VSUBS 0.008724f
C586 B.n443 VSUBS 0.008724f
C587 B.n444 VSUBS 0.008724f
C588 B.n445 VSUBS 0.008724f
C589 B.n446 VSUBS 0.008724f
C590 B.n447 VSUBS 0.008724f
C591 B.n448 VSUBS 0.008724f
C592 B.n449 VSUBS 0.008724f
C593 B.n450 VSUBS 0.008724f
C594 B.n451 VSUBS 0.008724f
C595 B.n452 VSUBS 0.008724f
C596 B.n453 VSUBS 0.008724f
C597 B.n454 VSUBS 0.008724f
C598 B.n455 VSUBS 0.008724f
C599 B.n456 VSUBS 0.008724f
C600 B.n457 VSUBS 0.008724f
C601 B.n458 VSUBS 0.008724f
C602 B.n459 VSUBS 0.008724f
C603 B.n460 VSUBS 0.008724f
C604 B.n461 VSUBS 0.008724f
C605 B.n462 VSUBS 0.008724f
C606 B.n463 VSUBS 0.008724f
C607 B.n464 VSUBS 0.008724f
C608 B.n465 VSUBS 0.008724f
C609 B.n466 VSUBS 0.008724f
C610 B.n467 VSUBS 0.008724f
C611 B.n468 VSUBS 0.008724f
C612 B.n469 VSUBS 0.008724f
C613 B.n470 VSUBS 0.008724f
C614 B.n471 VSUBS 0.008724f
C615 B.n472 VSUBS 0.008724f
C616 B.n473 VSUBS 0.008724f
C617 B.n474 VSUBS 0.008724f
C618 B.n475 VSUBS 0.008724f
C619 B.n476 VSUBS 0.008724f
C620 B.n477 VSUBS 0.008724f
C621 B.n478 VSUBS 0.008724f
C622 B.n479 VSUBS 0.008724f
C623 B.n480 VSUBS 0.008724f
C624 B.n481 VSUBS 0.008724f
C625 B.n482 VSUBS 0.008724f
C626 B.n483 VSUBS 0.008724f
C627 B.n484 VSUBS 0.008724f
C628 B.n485 VSUBS 0.008724f
C629 B.n486 VSUBS 0.008724f
C630 B.n487 VSUBS 0.008724f
C631 B.n488 VSUBS 0.008724f
C632 B.n489 VSUBS 0.008724f
C633 B.n490 VSUBS 0.008724f
C634 B.n491 VSUBS 0.008724f
C635 B.n492 VSUBS 0.008724f
C636 B.n493 VSUBS 0.008724f
C637 B.n494 VSUBS 0.008724f
C638 B.n495 VSUBS 0.008724f
C639 B.n496 VSUBS 0.008724f
C640 B.n497 VSUBS 0.008724f
C641 B.n498 VSUBS 0.008724f
C642 B.n499 VSUBS 0.008724f
C643 B.n500 VSUBS 0.008724f
C644 B.n501 VSUBS 0.008724f
C645 B.n502 VSUBS 0.008724f
C646 B.n503 VSUBS 0.008724f
C647 B.n504 VSUBS 0.008724f
C648 B.n505 VSUBS 0.008724f
C649 B.n506 VSUBS 0.008724f
C650 B.n507 VSUBS 0.008724f
C651 B.n508 VSUBS 0.008724f
C652 B.n509 VSUBS 0.008724f
C653 B.n510 VSUBS 0.008724f
C654 B.n511 VSUBS 0.008724f
C655 B.n512 VSUBS 0.008724f
C656 B.n513 VSUBS 0.008724f
C657 B.n514 VSUBS 0.008724f
C658 B.n515 VSUBS 0.008724f
C659 B.n516 VSUBS 0.008724f
C660 B.n517 VSUBS 0.008724f
C661 B.n518 VSUBS 0.008724f
C662 B.n519 VSUBS 0.008724f
C663 B.n520 VSUBS 0.008724f
C664 B.n521 VSUBS 0.008724f
C665 B.n522 VSUBS 0.008724f
C666 B.n523 VSUBS 0.008724f
C667 B.n524 VSUBS 0.008724f
C668 B.n525 VSUBS 0.008724f
C669 B.n526 VSUBS 0.008724f
C670 B.n527 VSUBS 0.008724f
C671 B.n528 VSUBS 0.008724f
C672 B.n529 VSUBS 0.008724f
C673 B.n530 VSUBS 0.008724f
C674 B.n531 VSUBS 0.008724f
C675 B.n532 VSUBS 0.008724f
C676 B.n533 VSUBS 0.008724f
C677 B.n534 VSUBS 0.008724f
C678 B.n535 VSUBS 0.008724f
C679 B.n536 VSUBS 0.008724f
C680 B.n537 VSUBS 0.008724f
C681 B.n538 VSUBS 0.008724f
C682 B.n539 VSUBS 0.008724f
C683 B.n540 VSUBS 0.008724f
C684 B.n541 VSUBS 0.008724f
C685 B.n542 VSUBS 0.008724f
C686 B.n543 VSUBS 0.008724f
C687 B.n544 VSUBS 0.008724f
C688 B.n545 VSUBS 0.008724f
C689 B.n546 VSUBS 0.008724f
C690 B.n547 VSUBS 0.008724f
C691 B.n548 VSUBS 0.008724f
C692 B.n549 VSUBS 0.008724f
C693 B.n550 VSUBS 0.020416f
C694 B.n551 VSUBS 0.020416f
C695 B.n552 VSUBS 0.02141f
C696 B.n553 VSUBS 0.008724f
C697 B.n554 VSUBS 0.008724f
C698 B.n555 VSUBS 0.008724f
C699 B.n556 VSUBS 0.008724f
C700 B.n557 VSUBS 0.008724f
C701 B.n558 VSUBS 0.008724f
C702 B.n559 VSUBS 0.008724f
C703 B.n560 VSUBS 0.008724f
C704 B.n561 VSUBS 0.008724f
C705 B.n562 VSUBS 0.008724f
C706 B.n563 VSUBS 0.008724f
C707 B.n564 VSUBS 0.008724f
C708 B.n565 VSUBS 0.008724f
C709 B.n566 VSUBS 0.008724f
C710 B.n567 VSUBS 0.008724f
C711 B.n568 VSUBS 0.008724f
C712 B.n569 VSUBS 0.008724f
C713 B.n570 VSUBS 0.008724f
C714 B.n571 VSUBS 0.008724f
C715 B.n572 VSUBS 0.008724f
C716 B.n573 VSUBS 0.008724f
C717 B.n574 VSUBS 0.008724f
C718 B.n575 VSUBS 0.008724f
C719 B.n576 VSUBS 0.008724f
C720 B.n577 VSUBS 0.008724f
C721 B.n578 VSUBS 0.008724f
C722 B.n579 VSUBS 0.008724f
C723 B.n580 VSUBS 0.008724f
C724 B.n581 VSUBS 0.008724f
C725 B.n582 VSUBS 0.008724f
C726 B.n583 VSUBS 0.008724f
C727 B.n584 VSUBS 0.008724f
C728 B.n585 VSUBS 0.008724f
C729 B.n586 VSUBS 0.008724f
C730 B.n587 VSUBS 0.008724f
C731 B.n588 VSUBS 0.008724f
C732 B.n589 VSUBS 0.008724f
C733 B.n590 VSUBS 0.008724f
C734 B.n591 VSUBS 0.008724f
C735 B.n592 VSUBS 0.008724f
C736 B.n593 VSUBS 0.008724f
C737 B.n594 VSUBS 0.008724f
C738 B.n595 VSUBS 0.008724f
C739 B.n596 VSUBS 0.008724f
C740 B.n597 VSUBS 0.008724f
C741 B.n598 VSUBS 0.008724f
C742 B.n599 VSUBS 0.008724f
C743 B.n600 VSUBS 0.008724f
C744 B.n601 VSUBS 0.008724f
C745 B.n602 VSUBS 0.008724f
C746 B.n603 VSUBS 0.008724f
C747 B.n604 VSUBS 0.008724f
C748 B.n605 VSUBS 0.008724f
C749 B.n606 VSUBS 0.008724f
C750 B.n607 VSUBS 0.008724f
C751 B.n608 VSUBS 0.008724f
C752 B.n609 VSUBS 0.008724f
C753 B.n610 VSUBS 0.008724f
C754 B.n611 VSUBS 0.008724f
C755 B.n612 VSUBS 0.008724f
C756 B.n613 VSUBS 0.008724f
C757 B.n614 VSUBS 0.008724f
C758 B.n615 VSUBS 0.00603f
C759 B.n616 VSUBS 0.020213f
C760 B.n617 VSUBS 0.007056f
C761 B.n618 VSUBS 0.008724f
C762 B.n619 VSUBS 0.008724f
C763 B.n620 VSUBS 0.008724f
C764 B.n621 VSUBS 0.008724f
C765 B.n622 VSUBS 0.008724f
C766 B.n623 VSUBS 0.008724f
C767 B.n624 VSUBS 0.008724f
C768 B.n625 VSUBS 0.008724f
C769 B.n626 VSUBS 0.008724f
C770 B.n627 VSUBS 0.008724f
C771 B.n628 VSUBS 0.008724f
C772 B.n629 VSUBS 0.007056f
C773 B.n630 VSUBS 0.008724f
C774 B.n631 VSUBS 0.008724f
C775 B.n632 VSUBS 0.008724f
C776 B.n633 VSUBS 0.008724f
C777 B.n634 VSUBS 0.008724f
C778 B.n635 VSUBS 0.008724f
C779 B.n636 VSUBS 0.008724f
C780 B.n637 VSUBS 0.008724f
C781 B.n638 VSUBS 0.008724f
C782 B.n639 VSUBS 0.008724f
C783 B.n640 VSUBS 0.008724f
C784 B.n641 VSUBS 0.008724f
C785 B.n642 VSUBS 0.008724f
C786 B.n643 VSUBS 0.008724f
C787 B.n644 VSUBS 0.008724f
C788 B.n645 VSUBS 0.008724f
C789 B.n646 VSUBS 0.008724f
C790 B.n647 VSUBS 0.008724f
C791 B.n648 VSUBS 0.008724f
C792 B.n649 VSUBS 0.008724f
C793 B.n650 VSUBS 0.008724f
C794 B.n651 VSUBS 0.008724f
C795 B.n652 VSUBS 0.008724f
C796 B.n653 VSUBS 0.008724f
C797 B.n654 VSUBS 0.008724f
C798 B.n655 VSUBS 0.008724f
C799 B.n656 VSUBS 0.008724f
C800 B.n657 VSUBS 0.008724f
C801 B.n658 VSUBS 0.008724f
C802 B.n659 VSUBS 0.008724f
C803 B.n660 VSUBS 0.008724f
C804 B.n661 VSUBS 0.008724f
C805 B.n662 VSUBS 0.008724f
C806 B.n663 VSUBS 0.008724f
C807 B.n664 VSUBS 0.008724f
C808 B.n665 VSUBS 0.008724f
C809 B.n666 VSUBS 0.008724f
C810 B.n667 VSUBS 0.008724f
C811 B.n668 VSUBS 0.008724f
C812 B.n669 VSUBS 0.008724f
C813 B.n670 VSUBS 0.008724f
C814 B.n671 VSUBS 0.008724f
C815 B.n672 VSUBS 0.008724f
C816 B.n673 VSUBS 0.008724f
C817 B.n674 VSUBS 0.008724f
C818 B.n675 VSUBS 0.008724f
C819 B.n676 VSUBS 0.008724f
C820 B.n677 VSUBS 0.008724f
C821 B.n678 VSUBS 0.008724f
C822 B.n679 VSUBS 0.008724f
C823 B.n680 VSUBS 0.008724f
C824 B.n681 VSUBS 0.008724f
C825 B.n682 VSUBS 0.008724f
C826 B.n683 VSUBS 0.008724f
C827 B.n684 VSUBS 0.008724f
C828 B.n685 VSUBS 0.008724f
C829 B.n686 VSUBS 0.008724f
C830 B.n687 VSUBS 0.008724f
C831 B.n688 VSUBS 0.008724f
C832 B.n689 VSUBS 0.008724f
C833 B.n690 VSUBS 0.008724f
C834 B.n691 VSUBS 0.008724f
C835 B.n692 VSUBS 0.008724f
C836 B.n693 VSUBS 0.008724f
C837 B.n694 VSUBS 0.02141f
C838 B.n695 VSUBS 0.020416f
C839 B.n696 VSUBS 0.020416f
C840 B.n697 VSUBS 0.008724f
C841 B.n698 VSUBS 0.008724f
C842 B.n699 VSUBS 0.008724f
C843 B.n700 VSUBS 0.008724f
C844 B.n701 VSUBS 0.008724f
C845 B.n702 VSUBS 0.008724f
C846 B.n703 VSUBS 0.008724f
C847 B.n704 VSUBS 0.008724f
C848 B.n705 VSUBS 0.008724f
C849 B.n706 VSUBS 0.008724f
C850 B.n707 VSUBS 0.008724f
C851 B.n708 VSUBS 0.008724f
C852 B.n709 VSUBS 0.008724f
C853 B.n710 VSUBS 0.008724f
C854 B.n711 VSUBS 0.008724f
C855 B.n712 VSUBS 0.008724f
C856 B.n713 VSUBS 0.008724f
C857 B.n714 VSUBS 0.008724f
C858 B.n715 VSUBS 0.008724f
C859 B.n716 VSUBS 0.008724f
C860 B.n717 VSUBS 0.008724f
C861 B.n718 VSUBS 0.008724f
C862 B.n719 VSUBS 0.008724f
C863 B.n720 VSUBS 0.008724f
C864 B.n721 VSUBS 0.008724f
C865 B.n722 VSUBS 0.008724f
C866 B.n723 VSUBS 0.008724f
C867 B.n724 VSUBS 0.008724f
C868 B.n725 VSUBS 0.008724f
C869 B.n726 VSUBS 0.008724f
C870 B.n727 VSUBS 0.008724f
C871 B.n728 VSUBS 0.008724f
C872 B.n729 VSUBS 0.008724f
C873 B.n730 VSUBS 0.008724f
C874 B.n731 VSUBS 0.008724f
C875 B.n732 VSUBS 0.008724f
C876 B.n733 VSUBS 0.008724f
C877 B.n734 VSUBS 0.008724f
C878 B.n735 VSUBS 0.008724f
C879 B.n736 VSUBS 0.008724f
C880 B.n737 VSUBS 0.008724f
C881 B.n738 VSUBS 0.008724f
C882 B.n739 VSUBS 0.008724f
C883 B.n740 VSUBS 0.008724f
C884 B.n741 VSUBS 0.008724f
C885 B.n742 VSUBS 0.008724f
C886 B.n743 VSUBS 0.008724f
C887 B.n744 VSUBS 0.008724f
C888 B.n745 VSUBS 0.008724f
C889 B.n746 VSUBS 0.008724f
C890 B.n747 VSUBS 0.008724f
C891 B.n748 VSUBS 0.008724f
C892 B.n749 VSUBS 0.008724f
C893 B.n750 VSUBS 0.008724f
C894 B.n751 VSUBS 0.008724f
C895 B.n752 VSUBS 0.008724f
C896 B.n753 VSUBS 0.008724f
C897 B.n754 VSUBS 0.008724f
C898 B.n755 VSUBS 0.008724f
C899 B.n756 VSUBS 0.008724f
C900 B.n757 VSUBS 0.008724f
C901 B.n758 VSUBS 0.008724f
C902 B.n759 VSUBS 0.008724f
C903 B.n760 VSUBS 0.008724f
C904 B.n761 VSUBS 0.008724f
C905 B.n762 VSUBS 0.008724f
C906 B.n763 VSUBS 0.011385f
C907 B.n764 VSUBS 0.012128f
C908 B.n765 VSUBS 0.024117f
C909 VTAIL.t9 VSUBS 0.277002f
C910 VTAIL.t17 VSUBS 0.277002f
C911 VTAIL.n0 VSUBS 2.00221f
C912 VTAIL.n1 VSUBS 0.92933f
C913 VTAIL.t2 VSUBS 2.6447f
C914 VTAIL.n2 VSUBS 1.07983f
C915 VTAIL.t5 VSUBS 0.277002f
C916 VTAIL.t19 VSUBS 0.277002f
C917 VTAIL.n3 VSUBS 2.00221f
C918 VTAIL.n4 VSUBS 1.00969f
C919 VTAIL.t7 VSUBS 0.277002f
C920 VTAIL.t8 VSUBS 0.277002f
C921 VTAIL.n5 VSUBS 2.00221f
C922 VTAIL.n6 VSUBS 2.53902f
C923 VTAIL.t15 VSUBS 0.277002f
C924 VTAIL.t18 VSUBS 0.277002f
C925 VTAIL.n7 VSUBS 2.00222f
C926 VTAIL.n8 VSUBS 2.53901f
C927 VTAIL.t10 VSUBS 0.277002f
C928 VTAIL.t12 VSUBS 0.277002f
C929 VTAIL.n9 VSUBS 2.00222f
C930 VTAIL.n10 VSUBS 1.00968f
C931 VTAIL.t13 VSUBS 2.64472f
C932 VTAIL.n11 VSUBS 1.07981f
C933 VTAIL.t0 VSUBS 0.277002f
C934 VTAIL.t6 VSUBS 0.277002f
C935 VTAIL.n12 VSUBS 2.00222f
C936 VTAIL.n13 VSUBS 0.966847f
C937 VTAIL.t3 VSUBS 0.277002f
C938 VTAIL.t1 VSUBS 0.277002f
C939 VTAIL.n14 VSUBS 2.00222f
C940 VTAIL.n15 VSUBS 1.00968f
C941 VTAIL.t4 VSUBS 2.6447f
C942 VTAIL.n16 VSUBS 2.48067f
C943 VTAIL.t16 VSUBS 2.6447f
C944 VTAIL.n17 VSUBS 2.48067f
C945 VTAIL.t11 VSUBS 0.277002f
C946 VTAIL.t14 VSUBS 0.277002f
C947 VTAIL.n18 VSUBS 2.00221f
C948 VTAIL.n19 VSUBS 0.87589f
C949 VDD2.t4 VSUBS 2.76791f
C950 VDD2.t6 VSUBS 0.269265f
C951 VDD2.t2 VSUBS 0.269265f
C952 VDD2.n0 VSUBS 2.10467f
C953 VDD2.n1 VSUBS 1.50835f
C954 VDD2.t5 VSUBS 0.269265f
C955 VDD2.t8 VSUBS 0.269265f
C956 VDD2.n2 VSUBS 2.11998f
C957 VDD2.n3 VSUBS 3.08699f
C958 VDD2.t1 VSUBS 2.74829f
C959 VDD2.n4 VSUBS 3.46833f
C960 VDD2.t9 VSUBS 0.269265f
C961 VDD2.t7 VSUBS 0.269265f
C962 VDD2.n5 VSUBS 2.10468f
C963 VDD2.n6 VSUBS 0.740725f
C964 VDD2.t0 VSUBS 0.269265f
C965 VDD2.t3 VSUBS 0.269265f
C966 VDD2.n7 VSUBS 2.11993f
C967 VN.n0 VSUBS 0.033532f
C968 VN.t2 VSUBS 2.09604f
C969 VN.n1 VSUBS 0.02728f
C970 VN.n2 VSUBS 0.033532f
C971 VN.t4 VSUBS 2.09604f
C972 VN.n3 VSUBS 0.040037f
C973 VN.n4 VSUBS 0.033532f
C974 VN.t7 VSUBS 2.09604f
C975 VN.n5 VSUBS 0.057278f
C976 VN.n6 VSUBS 0.249109f
C977 VN.t1 VSUBS 2.09604f
C978 VN.t9 VSUBS 2.26023f
C979 VN.n7 VSUBS 0.820738f
C980 VN.n8 VSUBS 0.835853f
C981 VN.n9 VSUBS 0.058763f
C982 VN.n10 VSUBS 0.040037f
C983 VN.n11 VSUBS 0.033532f
C984 VN.n12 VSUBS 0.033532f
C985 VN.n13 VSUBS 0.033532f
C986 VN.n14 VSUBS 0.047068f
C987 VN.n15 VSUBS 0.748853f
C988 VN.n16 VSUBS 0.047068f
C989 VN.n17 VSUBS 0.057278f
C990 VN.n18 VSUBS 0.033532f
C991 VN.n19 VSUBS 0.033532f
C992 VN.n20 VSUBS 0.033532f
C993 VN.n21 VSUBS 0.058763f
C994 VN.n22 VSUBS 0.748853f
C995 VN.n23 VSUBS 0.035961f
C996 VN.n24 VSUBS 0.067227f
C997 VN.n25 VSUBS 0.033532f
C998 VN.n26 VSUBS 0.033532f
C999 VN.n27 VSUBS 0.033532f
C1000 VN.n28 VSUBS 0.06589f
C1001 VN.n29 VSUBS 0.038429f
C1002 VN.n30 VSUBS 0.830119f
C1003 VN.n31 VSUBS 0.035601f
C1004 VN.n32 VSUBS 0.033532f
C1005 VN.t3 VSUBS 2.09604f
C1006 VN.n33 VSUBS 0.02728f
C1007 VN.n34 VSUBS 0.033532f
C1008 VN.t0 VSUBS 2.09604f
C1009 VN.n35 VSUBS 0.040037f
C1010 VN.n36 VSUBS 0.033532f
C1011 VN.t8 VSUBS 2.09604f
C1012 VN.n37 VSUBS 0.057278f
C1013 VN.n38 VSUBS 0.249109f
C1014 VN.t6 VSUBS 2.09604f
C1015 VN.t5 VSUBS 2.26023f
C1016 VN.n39 VSUBS 0.820738f
C1017 VN.n40 VSUBS 0.835853f
C1018 VN.n41 VSUBS 0.058763f
C1019 VN.n42 VSUBS 0.040037f
C1020 VN.n43 VSUBS 0.033532f
C1021 VN.n44 VSUBS 0.033532f
C1022 VN.n45 VSUBS 0.033532f
C1023 VN.n46 VSUBS 0.047068f
C1024 VN.n47 VSUBS 0.748853f
C1025 VN.n48 VSUBS 0.047068f
C1026 VN.n49 VSUBS 0.057278f
C1027 VN.n50 VSUBS 0.033532f
C1028 VN.n51 VSUBS 0.033532f
C1029 VN.n52 VSUBS 0.033532f
C1030 VN.n53 VSUBS 0.058763f
C1031 VN.n54 VSUBS 0.748853f
C1032 VN.n55 VSUBS 0.035961f
C1033 VN.n56 VSUBS 0.067227f
C1034 VN.n57 VSUBS 0.033532f
C1035 VN.n58 VSUBS 0.033532f
C1036 VN.n59 VSUBS 0.033532f
C1037 VN.n60 VSUBS 0.06589f
C1038 VN.n61 VSUBS 0.038429f
C1039 VN.n62 VSUBS 0.830119f
C1040 VN.n63 VSUBS 1.81462f
.ends

