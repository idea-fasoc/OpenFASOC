* NGSPICE file created from diff_pair_sample_1751.ext - technology: sky130A

.subckt diff_pair_sample_1751 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4524 pd=3.1 as=0.4524 ps=3.1 w=1.16 l=1.97
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4524 pd=3.1 as=0 ps=0 w=1.16 l=1.97
X2 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4524 pd=3.1 as=0.4524 ps=3.1 w=1.16 l=1.97
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.4524 pd=3.1 as=0 ps=0 w=1.16 l=1.97
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.4524 pd=3.1 as=0.4524 ps=3.1 w=1.16 l=1.97
X5 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4524 pd=3.1 as=0.4524 ps=3.1 w=1.16 l=1.97
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.4524 pd=3.1 as=0 ps=0 w=1.16 l=1.97
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4524 pd=3.1 as=0 ps=0 w=1.16 l=1.97
R0 VP.n0 VP.t1 107.85
R1 VP.n0 VP.t0 73.0773
R2 VP VP.n0 0.241678
R3 VTAIL.n3 VTAIL.t0 156.886
R4 VTAIL.n0 VTAIL.t2 156.886
R5 VTAIL.n2 VTAIL.t3 156.886
R6 VTAIL.n1 VTAIL.t1 156.886
R7 VTAIL.n1 VTAIL.n0 17.3324
R8 VTAIL.n3 VTAIL.n2 15.3496
R9 VTAIL.n2 VTAIL.n1 1.46171
R10 VTAIL VTAIL.n0 1.02421
R11 VTAIL VTAIL.n3 0.438
R12 VDD1 VDD1.t1 203.209
R13 VDD1 VDD1.t0 174.118
R14 B.n330 B.n329 585
R15 B.n331 B.n330 585
R16 B.n118 B.n57 585
R17 B.n117 B.n116 585
R18 B.n115 B.n114 585
R19 B.n113 B.n112 585
R20 B.n111 B.n110 585
R21 B.n109 B.n108 585
R22 B.n107 B.n106 585
R23 B.n105 B.n104 585
R24 B.n103 B.n102 585
R25 B.n100 B.n99 585
R26 B.n98 B.n97 585
R27 B.n96 B.n95 585
R28 B.n94 B.n93 585
R29 B.n92 B.n91 585
R30 B.n90 B.n89 585
R31 B.n88 B.n87 585
R32 B.n86 B.n85 585
R33 B.n84 B.n83 585
R34 B.n82 B.n81 585
R35 B.n80 B.n79 585
R36 B.n78 B.n77 585
R37 B.n76 B.n75 585
R38 B.n74 B.n73 585
R39 B.n72 B.n71 585
R40 B.n70 B.n69 585
R41 B.n68 B.n67 585
R42 B.n66 B.n65 585
R43 B.n64 B.n63 585
R44 B.n328 B.n42 585
R45 B.n332 B.n42 585
R46 B.n327 B.n41 585
R47 B.n333 B.n41 585
R48 B.n326 B.n325 585
R49 B.n325 B.n37 585
R50 B.n324 B.n36 585
R51 B.n339 B.n36 585
R52 B.n323 B.n35 585
R53 B.n340 B.n35 585
R54 B.n322 B.n34 585
R55 B.n341 B.n34 585
R56 B.n321 B.n320 585
R57 B.n320 B.n33 585
R58 B.n319 B.n29 585
R59 B.n347 B.n29 585
R60 B.n318 B.n28 585
R61 B.n348 B.n28 585
R62 B.n317 B.n27 585
R63 B.n349 B.n27 585
R64 B.n316 B.n315 585
R65 B.n315 B.n23 585
R66 B.n314 B.n22 585
R67 B.n355 B.n22 585
R68 B.n313 B.n21 585
R69 B.n356 B.n21 585
R70 B.n312 B.n20 585
R71 B.n357 B.n20 585
R72 B.n311 B.n310 585
R73 B.n310 B.n16 585
R74 B.n309 B.n15 585
R75 B.n363 B.n15 585
R76 B.n308 B.n14 585
R77 B.n364 B.n14 585
R78 B.n307 B.n13 585
R79 B.n365 B.n13 585
R80 B.n306 B.n305 585
R81 B.n305 B.n12 585
R82 B.n304 B.n303 585
R83 B.n304 B.n8 585
R84 B.n302 B.n7 585
R85 B.n372 B.n7 585
R86 B.n301 B.n6 585
R87 B.n373 B.n6 585
R88 B.n300 B.n5 585
R89 B.n374 B.n5 585
R90 B.n299 B.n298 585
R91 B.n298 B.n4 585
R92 B.n297 B.n119 585
R93 B.n297 B.n296 585
R94 B.n287 B.n120 585
R95 B.n121 B.n120 585
R96 B.n289 B.n288 585
R97 B.n290 B.n289 585
R98 B.n286 B.n125 585
R99 B.n129 B.n125 585
R100 B.n285 B.n284 585
R101 B.n284 B.n283 585
R102 B.n127 B.n126 585
R103 B.n128 B.n127 585
R104 B.n276 B.n275 585
R105 B.n277 B.n276 585
R106 B.n274 B.n134 585
R107 B.n134 B.n133 585
R108 B.n273 B.n272 585
R109 B.n272 B.n271 585
R110 B.n136 B.n135 585
R111 B.n137 B.n136 585
R112 B.n264 B.n263 585
R113 B.n265 B.n264 585
R114 B.n262 B.n142 585
R115 B.n142 B.n141 585
R116 B.n261 B.n260 585
R117 B.n260 B.n259 585
R118 B.n144 B.n143 585
R119 B.n252 B.n144 585
R120 B.n251 B.n250 585
R121 B.n253 B.n251 585
R122 B.n249 B.n149 585
R123 B.n149 B.n148 585
R124 B.n248 B.n247 585
R125 B.n247 B.n246 585
R126 B.n151 B.n150 585
R127 B.n152 B.n151 585
R128 B.n239 B.n238 585
R129 B.n240 B.n239 585
R130 B.n237 B.n157 585
R131 B.n157 B.n156 585
R132 B.n231 B.n230 585
R133 B.n229 B.n173 585
R134 B.n228 B.n172 585
R135 B.n233 B.n172 585
R136 B.n227 B.n226 585
R137 B.n225 B.n224 585
R138 B.n223 B.n222 585
R139 B.n221 B.n220 585
R140 B.n219 B.n218 585
R141 B.n217 B.n216 585
R142 B.n215 B.n214 585
R143 B.n212 B.n211 585
R144 B.n210 B.n209 585
R145 B.n208 B.n207 585
R146 B.n206 B.n205 585
R147 B.n204 B.n203 585
R148 B.n202 B.n201 585
R149 B.n200 B.n199 585
R150 B.n198 B.n197 585
R151 B.n196 B.n195 585
R152 B.n194 B.n193 585
R153 B.n192 B.n191 585
R154 B.n190 B.n189 585
R155 B.n188 B.n187 585
R156 B.n186 B.n185 585
R157 B.n184 B.n183 585
R158 B.n182 B.n181 585
R159 B.n180 B.n179 585
R160 B.n159 B.n158 585
R161 B.n236 B.n235 585
R162 B.n155 B.n154 585
R163 B.n156 B.n155 585
R164 B.n242 B.n241 585
R165 B.n241 B.n240 585
R166 B.n243 B.n153 585
R167 B.n153 B.n152 585
R168 B.n245 B.n244 585
R169 B.n246 B.n245 585
R170 B.n147 B.n146 585
R171 B.n148 B.n147 585
R172 B.n255 B.n254 585
R173 B.n254 B.n253 585
R174 B.n256 B.n145 585
R175 B.n252 B.n145 585
R176 B.n258 B.n257 585
R177 B.n259 B.n258 585
R178 B.n140 B.n139 585
R179 B.n141 B.n140 585
R180 B.n267 B.n266 585
R181 B.n266 B.n265 585
R182 B.n268 B.n138 585
R183 B.n138 B.n137 585
R184 B.n270 B.n269 585
R185 B.n271 B.n270 585
R186 B.n132 B.n131 585
R187 B.n133 B.n132 585
R188 B.n279 B.n278 585
R189 B.n278 B.n277 585
R190 B.n280 B.n130 585
R191 B.n130 B.n128 585
R192 B.n282 B.n281 585
R193 B.n283 B.n282 585
R194 B.n124 B.n123 585
R195 B.n129 B.n124 585
R196 B.n292 B.n291 585
R197 B.n291 B.n290 585
R198 B.n293 B.n122 585
R199 B.n122 B.n121 585
R200 B.n295 B.n294 585
R201 B.n296 B.n295 585
R202 B.n3 B.n0 585
R203 B.n4 B.n3 585
R204 B.n371 B.n1 585
R205 B.n372 B.n371 585
R206 B.n370 B.n369 585
R207 B.n370 B.n8 585
R208 B.n368 B.n9 585
R209 B.n12 B.n9 585
R210 B.n367 B.n366 585
R211 B.n366 B.n365 585
R212 B.n11 B.n10 585
R213 B.n364 B.n11 585
R214 B.n362 B.n361 585
R215 B.n363 B.n362 585
R216 B.n360 B.n17 585
R217 B.n17 B.n16 585
R218 B.n359 B.n358 585
R219 B.n358 B.n357 585
R220 B.n19 B.n18 585
R221 B.n356 B.n19 585
R222 B.n354 B.n353 585
R223 B.n355 B.n354 585
R224 B.n352 B.n24 585
R225 B.n24 B.n23 585
R226 B.n351 B.n350 585
R227 B.n350 B.n349 585
R228 B.n26 B.n25 585
R229 B.n348 B.n26 585
R230 B.n346 B.n345 585
R231 B.n347 B.n346 585
R232 B.n344 B.n30 585
R233 B.n33 B.n30 585
R234 B.n343 B.n342 585
R235 B.n342 B.n341 585
R236 B.n32 B.n31 585
R237 B.n340 B.n32 585
R238 B.n338 B.n337 585
R239 B.n339 B.n338 585
R240 B.n336 B.n38 585
R241 B.n38 B.n37 585
R242 B.n335 B.n334 585
R243 B.n334 B.n333 585
R244 B.n40 B.n39 585
R245 B.n332 B.n40 585
R246 B.n375 B.n374 585
R247 B.n373 B.n2 585
R248 B.n63 B.n40 526.135
R249 B.n330 B.n42 526.135
R250 B.n235 B.n157 526.135
R251 B.n231 B.n155 526.135
R252 B.n331 B.n56 256.663
R253 B.n331 B.n55 256.663
R254 B.n331 B.n54 256.663
R255 B.n331 B.n53 256.663
R256 B.n331 B.n52 256.663
R257 B.n331 B.n51 256.663
R258 B.n331 B.n50 256.663
R259 B.n331 B.n49 256.663
R260 B.n331 B.n48 256.663
R261 B.n331 B.n47 256.663
R262 B.n331 B.n46 256.663
R263 B.n331 B.n45 256.663
R264 B.n331 B.n44 256.663
R265 B.n331 B.n43 256.663
R266 B.n233 B.n232 256.663
R267 B.n233 B.n160 256.663
R268 B.n233 B.n161 256.663
R269 B.n233 B.n162 256.663
R270 B.n233 B.n163 256.663
R271 B.n233 B.n164 256.663
R272 B.n233 B.n165 256.663
R273 B.n233 B.n166 256.663
R274 B.n233 B.n167 256.663
R275 B.n233 B.n168 256.663
R276 B.n233 B.n169 256.663
R277 B.n233 B.n170 256.663
R278 B.n233 B.n171 256.663
R279 B.n234 B.n233 256.663
R280 B.n377 B.n376 256.663
R281 B.n233 B.n156 227.351
R282 B.n332 B.n331 227.351
R283 B.n60 B.t13 221.037
R284 B.n58 B.t2 221.037
R285 B.n176 B.t10 221.037
R286 B.n174 B.t6 221.037
R287 B.n60 B.t14 192.07
R288 B.n58 B.t4 192.07
R289 B.n176 B.t12 192.07
R290 B.n174 B.t9 192.07
R291 B.n67 B.n66 163.367
R292 B.n71 B.n70 163.367
R293 B.n75 B.n74 163.367
R294 B.n79 B.n78 163.367
R295 B.n83 B.n82 163.367
R296 B.n87 B.n86 163.367
R297 B.n91 B.n90 163.367
R298 B.n95 B.n94 163.367
R299 B.n99 B.n98 163.367
R300 B.n104 B.n103 163.367
R301 B.n108 B.n107 163.367
R302 B.n112 B.n111 163.367
R303 B.n116 B.n115 163.367
R304 B.n330 B.n57 163.367
R305 B.n239 B.n157 163.367
R306 B.n239 B.n151 163.367
R307 B.n247 B.n151 163.367
R308 B.n247 B.n149 163.367
R309 B.n251 B.n149 163.367
R310 B.n251 B.n144 163.367
R311 B.n260 B.n144 163.367
R312 B.n260 B.n142 163.367
R313 B.n264 B.n142 163.367
R314 B.n264 B.n136 163.367
R315 B.n272 B.n136 163.367
R316 B.n272 B.n134 163.367
R317 B.n276 B.n134 163.367
R318 B.n276 B.n127 163.367
R319 B.n284 B.n127 163.367
R320 B.n284 B.n125 163.367
R321 B.n289 B.n125 163.367
R322 B.n289 B.n120 163.367
R323 B.n297 B.n120 163.367
R324 B.n298 B.n297 163.367
R325 B.n298 B.n5 163.367
R326 B.n6 B.n5 163.367
R327 B.n7 B.n6 163.367
R328 B.n304 B.n7 163.367
R329 B.n305 B.n304 163.367
R330 B.n305 B.n13 163.367
R331 B.n14 B.n13 163.367
R332 B.n15 B.n14 163.367
R333 B.n310 B.n15 163.367
R334 B.n310 B.n20 163.367
R335 B.n21 B.n20 163.367
R336 B.n22 B.n21 163.367
R337 B.n315 B.n22 163.367
R338 B.n315 B.n27 163.367
R339 B.n28 B.n27 163.367
R340 B.n29 B.n28 163.367
R341 B.n320 B.n29 163.367
R342 B.n320 B.n34 163.367
R343 B.n35 B.n34 163.367
R344 B.n36 B.n35 163.367
R345 B.n325 B.n36 163.367
R346 B.n325 B.n41 163.367
R347 B.n42 B.n41 163.367
R348 B.n173 B.n172 163.367
R349 B.n226 B.n172 163.367
R350 B.n224 B.n223 163.367
R351 B.n220 B.n219 163.367
R352 B.n216 B.n215 163.367
R353 B.n211 B.n210 163.367
R354 B.n207 B.n206 163.367
R355 B.n203 B.n202 163.367
R356 B.n199 B.n198 163.367
R357 B.n195 B.n194 163.367
R358 B.n191 B.n190 163.367
R359 B.n187 B.n186 163.367
R360 B.n183 B.n182 163.367
R361 B.n179 B.n159 163.367
R362 B.n241 B.n155 163.367
R363 B.n241 B.n153 163.367
R364 B.n245 B.n153 163.367
R365 B.n245 B.n147 163.367
R366 B.n254 B.n147 163.367
R367 B.n254 B.n145 163.367
R368 B.n258 B.n145 163.367
R369 B.n258 B.n140 163.367
R370 B.n266 B.n140 163.367
R371 B.n266 B.n138 163.367
R372 B.n270 B.n138 163.367
R373 B.n270 B.n132 163.367
R374 B.n278 B.n132 163.367
R375 B.n278 B.n130 163.367
R376 B.n282 B.n130 163.367
R377 B.n282 B.n124 163.367
R378 B.n291 B.n124 163.367
R379 B.n291 B.n122 163.367
R380 B.n295 B.n122 163.367
R381 B.n295 B.n3 163.367
R382 B.n375 B.n3 163.367
R383 B.n371 B.n2 163.367
R384 B.n371 B.n370 163.367
R385 B.n370 B.n9 163.367
R386 B.n366 B.n9 163.367
R387 B.n366 B.n11 163.367
R388 B.n362 B.n11 163.367
R389 B.n362 B.n17 163.367
R390 B.n358 B.n17 163.367
R391 B.n358 B.n19 163.367
R392 B.n354 B.n19 163.367
R393 B.n354 B.n24 163.367
R394 B.n350 B.n24 163.367
R395 B.n350 B.n26 163.367
R396 B.n346 B.n26 163.367
R397 B.n346 B.n30 163.367
R398 B.n342 B.n30 163.367
R399 B.n342 B.n32 163.367
R400 B.n338 B.n32 163.367
R401 B.n338 B.n38 163.367
R402 B.n334 B.n38 163.367
R403 B.n334 B.n40 163.367
R404 B.n61 B.t15 147.464
R405 B.n59 B.t5 147.464
R406 B.n177 B.t11 147.464
R407 B.n175 B.t8 147.464
R408 B.n240 B.n156 116.24
R409 B.n240 B.n152 116.24
R410 B.n246 B.n152 116.24
R411 B.n246 B.n148 116.24
R412 B.n253 B.n148 116.24
R413 B.n253 B.n252 116.24
R414 B.n259 B.n141 116.24
R415 B.n265 B.n141 116.24
R416 B.n265 B.n137 116.24
R417 B.n271 B.n137 116.24
R418 B.n271 B.n133 116.24
R419 B.n277 B.n133 116.24
R420 B.n277 B.n128 116.24
R421 B.n283 B.n128 116.24
R422 B.n283 B.n129 116.24
R423 B.n290 B.n121 116.24
R424 B.n296 B.n121 116.24
R425 B.n296 B.n4 116.24
R426 B.n374 B.n4 116.24
R427 B.n374 B.n373 116.24
R428 B.n373 B.n372 116.24
R429 B.n372 B.n8 116.24
R430 B.n12 B.n8 116.24
R431 B.n365 B.n12 116.24
R432 B.n364 B.n363 116.24
R433 B.n363 B.n16 116.24
R434 B.n357 B.n16 116.24
R435 B.n357 B.n356 116.24
R436 B.n356 B.n355 116.24
R437 B.n355 B.n23 116.24
R438 B.n349 B.n23 116.24
R439 B.n349 B.n348 116.24
R440 B.n348 B.n347 116.24
R441 B.n341 B.n33 116.24
R442 B.n341 B.n340 116.24
R443 B.n340 B.n339 116.24
R444 B.n339 B.n37 116.24
R445 B.n333 B.n37 116.24
R446 B.n333 B.n332 116.24
R447 B.n63 B.n43 71.676
R448 B.n67 B.n44 71.676
R449 B.n71 B.n45 71.676
R450 B.n75 B.n46 71.676
R451 B.n79 B.n47 71.676
R452 B.n83 B.n48 71.676
R453 B.n87 B.n49 71.676
R454 B.n91 B.n50 71.676
R455 B.n95 B.n51 71.676
R456 B.n99 B.n52 71.676
R457 B.n104 B.n53 71.676
R458 B.n108 B.n54 71.676
R459 B.n112 B.n55 71.676
R460 B.n116 B.n56 71.676
R461 B.n57 B.n56 71.676
R462 B.n115 B.n55 71.676
R463 B.n111 B.n54 71.676
R464 B.n107 B.n53 71.676
R465 B.n103 B.n52 71.676
R466 B.n98 B.n51 71.676
R467 B.n94 B.n50 71.676
R468 B.n90 B.n49 71.676
R469 B.n86 B.n48 71.676
R470 B.n82 B.n47 71.676
R471 B.n78 B.n46 71.676
R472 B.n74 B.n45 71.676
R473 B.n70 B.n44 71.676
R474 B.n66 B.n43 71.676
R475 B.n232 B.n231 71.676
R476 B.n226 B.n160 71.676
R477 B.n223 B.n161 71.676
R478 B.n219 B.n162 71.676
R479 B.n215 B.n163 71.676
R480 B.n210 B.n164 71.676
R481 B.n206 B.n165 71.676
R482 B.n202 B.n166 71.676
R483 B.n198 B.n167 71.676
R484 B.n194 B.n168 71.676
R485 B.n190 B.n169 71.676
R486 B.n186 B.n170 71.676
R487 B.n182 B.n171 71.676
R488 B.n234 B.n159 71.676
R489 B.n232 B.n173 71.676
R490 B.n224 B.n160 71.676
R491 B.n220 B.n161 71.676
R492 B.n216 B.n162 71.676
R493 B.n211 B.n163 71.676
R494 B.n207 B.n164 71.676
R495 B.n203 B.n165 71.676
R496 B.n199 B.n166 71.676
R497 B.n195 B.n167 71.676
R498 B.n191 B.n168 71.676
R499 B.n187 B.n169 71.676
R500 B.n183 B.n170 71.676
R501 B.n179 B.n171 71.676
R502 B.n235 B.n234 71.676
R503 B.n376 B.n375 71.676
R504 B.n376 B.n2 71.676
R505 B.n252 B.t7 63.2484
R506 B.n33 B.t3 63.2484
R507 B.n129 B.t1 59.8296
R508 B.t0 B.n364 59.8296
R509 B.n62 B.n61 59.5399
R510 B.n101 B.n59 59.5399
R511 B.n178 B.n177 59.5399
R512 B.n213 B.n175 59.5399
R513 B.n290 B.t1 56.4108
R514 B.n365 B.t0 56.4108
R515 B.n259 B.t7 52.992
R516 B.n347 B.t3 52.992
R517 B.n61 B.n60 44.6066
R518 B.n59 B.n58 44.6066
R519 B.n177 B.n176 44.6066
R520 B.n175 B.n174 44.6066
R521 B.n230 B.n154 34.1859
R522 B.n237 B.n236 34.1859
R523 B.n329 B.n328 34.1859
R524 B.n64 B.n39 34.1859
R525 B B.n377 18.0485
R526 B.n242 B.n154 10.6151
R527 B.n243 B.n242 10.6151
R528 B.n244 B.n243 10.6151
R529 B.n244 B.n146 10.6151
R530 B.n255 B.n146 10.6151
R531 B.n256 B.n255 10.6151
R532 B.n257 B.n256 10.6151
R533 B.n257 B.n139 10.6151
R534 B.n267 B.n139 10.6151
R535 B.n268 B.n267 10.6151
R536 B.n269 B.n268 10.6151
R537 B.n269 B.n131 10.6151
R538 B.n279 B.n131 10.6151
R539 B.n280 B.n279 10.6151
R540 B.n281 B.n280 10.6151
R541 B.n281 B.n123 10.6151
R542 B.n292 B.n123 10.6151
R543 B.n293 B.n292 10.6151
R544 B.n294 B.n293 10.6151
R545 B.n294 B.n0 10.6151
R546 B.n230 B.n229 10.6151
R547 B.n229 B.n228 10.6151
R548 B.n228 B.n227 10.6151
R549 B.n227 B.n225 10.6151
R550 B.n225 B.n222 10.6151
R551 B.n222 B.n221 10.6151
R552 B.n221 B.n218 10.6151
R553 B.n218 B.n217 10.6151
R554 B.n217 B.n214 10.6151
R555 B.n212 B.n209 10.6151
R556 B.n209 B.n208 10.6151
R557 B.n208 B.n205 10.6151
R558 B.n205 B.n204 10.6151
R559 B.n204 B.n201 10.6151
R560 B.n201 B.n200 10.6151
R561 B.n200 B.n197 10.6151
R562 B.n197 B.n196 10.6151
R563 B.n193 B.n192 10.6151
R564 B.n192 B.n189 10.6151
R565 B.n189 B.n188 10.6151
R566 B.n188 B.n185 10.6151
R567 B.n185 B.n184 10.6151
R568 B.n184 B.n181 10.6151
R569 B.n181 B.n180 10.6151
R570 B.n180 B.n158 10.6151
R571 B.n236 B.n158 10.6151
R572 B.n238 B.n237 10.6151
R573 B.n238 B.n150 10.6151
R574 B.n248 B.n150 10.6151
R575 B.n249 B.n248 10.6151
R576 B.n250 B.n249 10.6151
R577 B.n250 B.n143 10.6151
R578 B.n261 B.n143 10.6151
R579 B.n262 B.n261 10.6151
R580 B.n263 B.n262 10.6151
R581 B.n263 B.n135 10.6151
R582 B.n273 B.n135 10.6151
R583 B.n274 B.n273 10.6151
R584 B.n275 B.n274 10.6151
R585 B.n275 B.n126 10.6151
R586 B.n285 B.n126 10.6151
R587 B.n286 B.n285 10.6151
R588 B.n288 B.n286 10.6151
R589 B.n288 B.n287 10.6151
R590 B.n287 B.n119 10.6151
R591 B.n299 B.n119 10.6151
R592 B.n300 B.n299 10.6151
R593 B.n301 B.n300 10.6151
R594 B.n302 B.n301 10.6151
R595 B.n303 B.n302 10.6151
R596 B.n306 B.n303 10.6151
R597 B.n307 B.n306 10.6151
R598 B.n308 B.n307 10.6151
R599 B.n309 B.n308 10.6151
R600 B.n311 B.n309 10.6151
R601 B.n312 B.n311 10.6151
R602 B.n313 B.n312 10.6151
R603 B.n314 B.n313 10.6151
R604 B.n316 B.n314 10.6151
R605 B.n317 B.n316 10.6151
R606 B.n318 B.n317 10.6151
R607 B.n319 B.n318 10.6151
R608 B.n321 B.n319 10.6151
R609 B.n322 B.n321 10.6151
R610 B.n323 B.n322 10.6151
R611 B.n324 B.n323 10.6151
R612 B.n326 B.n324 10.6151
R613 B.n327 B.n326 10.6151
R614 B.n328 B.n327 10.6151
R615 B.n369 B.n1 10.6151
R616 B.n369 B.n368 10.6151
R617 B.n368 B.n367 10.6151
R618 B.n367 B.n10 10.6151
R619 B.n361 B.n10 10.6151
R620 B.n361 B.n360 10.6151
R621 B.n360 B.n359 10.6151
R622 B.n359 B.n18 10.6151
R623 B.n353 B.n18 10.6151
R624 B.n353 B.n352 10.6151
R625 B.n352 B.n351 10.6151
R626 B.n351 B.n25 10.6151
R627 B.n345 B.n25 10.6151
R628 B.n345 B.n344 10.6151
R629 B.n344 B.n343 10.6151
R630 B.n343 B.n31 10.6151
R631 B.n337 B.n31 10.6151
R632 B.n337 B.n336 10.6151
R633 B.n336 B.n335 10.6151
R634 B.n335 B.n39 10.6151
R635 B.n65 B.n64 10.6151
R636 B.n68 B.n65 10.6151
R637 B.n69 B.n68 10.6151
R638 B.n72 B.n69 10.6151
R639 B.n73 B.n72 10.6151
R640 B.n76 B.n73 10.6151
R641 B.n77 B.n76 10.6151
R642 B.n80 B.n77 10.6151
R643 B.n81 B.n80 10.6151
R644 B.n85 B.n84 10.6151
R645 B.n88 B.n85 10.6151
R646 B.n89 B.n88 10.6151
R647 B.n92 B.n89 10.6151
R648 B.n93 B.n92 10.6151
R649 B.n96 B.n93 10.6151
R650 B.n97 B.n96 10.6151
R651 B.n100 B.n97 10.6151
R652 B.n105 B.n102 10.6151
R653 B.n106 B.n105 10.6151
R654 B.n109 B.n106 10.6151
R655 B.n110 B.n109 10.6151
R656 B.n113 B.n110 10.6151
R657 B.n114 B.n113 10.6151
R658 B.n117 B.n114 10.6151
R659 B.n118 B.n117 10.6151
R660 B.n329 B.n118 10.6151
R661 B.n377 B.n0 8.11757
R662 B.n377 B.n1 8.11757
R663 B.n213 B.n212 6.5566
R664 B.n196 B.n178 6.5566
R665 B.n84 B.n62 6.5566
R666 B.n101 B.n100 6.5566
R667 B.n214 B.n213 4.05904
R668 B.n193 B.n178 4.05904
R669 B.n81 B.n62 4.05904
R670 B.n102 B.n101 4.05904
R671 VN VN.t1 108.041
R672 VN VN.t0 73.3184
R673 VDD2.n0 VDD2.t1 202.189
R674 VDD2.n0 VDD2.t0 173.564
R675 VDD2 VDD2.n0 0.554379
C0 VDD2 VTAIL 2.04194f
C1 VDD2 VN 0.484267f
C2 VDD1 VDD2 0.598277f
C3 VDD2 VP 0.314486f
C4 VN VTAIL 0.775817f
C5 VDD1 VTAIL 1.99313f
C6 VP VTAIL 0.789948f
C7 VDD1 VN 0.155683f
C8 VN VP 3.15675f
C9 VDD1 VP 0.641394f
C10 VDD2 B 2.227313f
C11 VDD1 B 2.32364f
C12 VTAIL B 2.329312f
C13 VN B 6.7471f
C14 VP B 4.652924f
C15 VDD2.t1 B 0.210121f
C16 VDD2.t0 B 0.11093f
C17 VDD2.n0 B 1.58954f
C18 VN.t0 B 0.400484f
C19 VN.t1 B 0.780232f
C20 VTAIL.t2 B 0.062394f
C21 VTAIL.n0 B 0.458118f
C22 VTAIL.t1 B 0.062394f
C23 VTAIL.n1 B 0.474319f
C24 VTAIL.t3 B 0.062394f
C25 VTAIL.n2 B 0.400893f
C26 VTAIL.t0 B 0.062394f
C27 VTAIL.n3 B 0.362982f
C28 VP.t1 B 0.785228f
C29 VP.t0 B 0.406157f
C30 VP.n0 B 1.95039f
.ends

