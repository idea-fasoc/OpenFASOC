* NGSPICE file created from diff_pair_sample_0773.ext - technology: sky130A

.subckt diff_pair_sample_0773 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t3 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=1.5249 pd=8.6 as=0.64515 ps=4.24 w=3.91 l=0.85
X1 VTAIL.t3 VP.t0 VDD1.t3 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=1.5249 pd=8.6 as=0.64515 ps=4.24 w=3.91 l=0.85
X2 VDD1.t2 VP.t1 VTAIL.t2 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=0.64515 pd=4.24 as=1.5249 ps=8.6 w=3.91 l=0.85
X3 B.t11 B.t9 B.t10 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=1.5249 pd=8.6 as=0 ps=0 w=3.91 l=0.85
X4 VDD2.t2 VN.t1 VTAIL.t6 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=0.64515 pd=4.24 as=1.5249 ps=8.6 w=3.91 l=0.85
X5 B.t8 B.t6 B.t7 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=1.5249 pd=8.6 as=0 ps=0 w=3.91 l=0.85
X6 VTAIL.t0 VP.t2 VDD1.t1 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=1.5249 pd=8.6 as=0.64515 ps=4.24 w=3.91 l=0.85
X7 B.t5 B.t3 B.t4 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=1.5249 pd=8.6 as=0 ps=0 w=3.91 l=0.85
X8 B.t2 B.t0 B.t1 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=1.5249 pd=8.6 as=0 ps=0 w=3.91 l=0.85
X9 VTAIL.t5 VN.t2 VDD2.t1 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=1.5249 pd=8.6 as=0.64515 ps=4.24 w=3.91 l=0.85
X10 VDD1.t0 VP.t3 VTAIL.t1 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=0.64515 pd=4.24 as=1.5249 ps=8.6 w=3.91 l=0.85
X11 VDD2.t0 VN.t3 VTAIL.t4 w_n1678_n1750# sky130_fd_pr__pfet_01v8 ad=0.64515 pd=4.24 as=1.5249 ps=8.6 w=3.91 l=0.85
R0 VN.n0 VN.t2 178.356
R1 VN.n1 VN.t1 178.356
R2 VN.n0 VN.t3 178.305
R3 VN.n1 VN.t0 178.305
R4 VN VN.n1 79.8912
R5 VN VN.n0 44.7132
R6 VDD2.n2 VDD2.n0 145.062
R7 VDD2.n2 VDD2.n1 114.925
R8 VDD2.n1 VDD2.t3 8.3138
R9 VDD2.n1 VDD2.t2 8.3138
R10 VDD2.n0 VDD2.t1 8.3138
R11 VDD2.n0 VDD2.t0 8.3138
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n154 VTAIL.n140 756.745
R14 VTAIL.n14 VTAIL.n0 756.745
R15 VTAIL.n34 VTAIL.n20 756.745
R16 VTAIL.n54 VTAIL.n40 756.745
R17 VTAIL.n134 VTAIL.n120 756.745
R18 VTAIL.n114 VTAIL.n100 756.745
R19 VTAIL.n94 VTAIL.n80 756.745
R20 VTAIL.n74 VTAIL.n60 756.745
R21 VTAIL.n147 VTAIL.n146 585
R22 VTAIL.n144 VTAIL.n143 585
R23 VTAIL.n153 VTAIL.n152 585
R24 VTAIL.n155 VTAIL.n154 585
R25 VTAIL.n7 VTAIL.n6 585
R26 VTAIL.n4 VTAIL.n3 585
R27 VTAIL.n13 VTAIL.n12 585
R28 VTAIL.n15 VTAIL.n14 585
R29 VTAIL.n27 VTAIL.n26 585
R30 VTAIL.n24 VTAIL.n23 585
R31 VTAIL.n33 VTAIL.n32 585
R32 VTAIL.n35 VTAIL.n34 585
R33 VTAIL.n47 VTAIL.n46 585
R34 VTAIL.n44 VTAIL.n43 585
R35 VTAIL.n53 VTAIL.n52 585
R36 VTAIL.n55 VTAIL.n54 585
R37 VTAIL.n135 VTAIL.n134 585
R38 VTAIL.n133 VTAIL.n132 585
R39 VTAIL.n124 VTAIL.n123 585
R40 VTAIL.n127 VTAIL.n126 585
R41 VTAIL.n115 VTAIL.n114 585
R42 VTAIL.n113 VTAIL.n112 585
R43 VTAIL.n104 VTAIL.n103 585
R44 VTAIL.n107 VTAIL.n106 585
R45 VTAIL.n95 VTAIL.n94 585
R46 VTAIL.n93 VTAIL.n92 585
R47 VTAIL.n84 VTAIL.n83 585
R48 VTAIL.n87 VTAIL.n86 585
R49 VTAIL.n75 VTAIL.n74 585
R50 VTAIL.n73 VTAIL.n72 585
R51 VTAIL.n64 VTAIL.n63 585
R52 VTAIL.n67 VTAIL.n66 585
R53 VTAIL.t4 VTAIL.n145 330.707
R54 VTAIL.t5 VTAIL.n5 330.707
R55 VTAIL.t1 VTAIL.n25 330.707
R56 VTAIL.t3 VTAIL.n45 330.707
R57 VTAIL.t2 VTAIL.n125 330.707
R58 VTAIL.t0 VTAIL.n105 330.707
R59 VTAIL.t6 VTAIL.n85 330.707
R60 VTAIL.t7 VTAIL.n65 330.707
R61 VTAIL.n146 VTAIL.n143 171.744
R62 VTAIL.n153 VTAIL.n143 171.744
R63 VTAIL.n154 VTAIL.n153 171.744
R64 VTAIL.n6 VTAIL.n3 171.744
R65 VTAIL.n13 VTAIL.n3 171.744
R66 VTAIL.n14 VTAIL.n13 171.744
R67 VTAIL.n26 VTAIL.n23 171.744
R68 VTAIL.n33 VTAIL.n23 171.744
R69 VTAIL.n34 VTAIL.n33 171.744
R70 VTAIL.n46 VTAIL.n43 171.744
R71 VTAIL.n53 VTAIL.n43 171.744
R72 VTAIL.n54 VTAIL.n53 171.744
R73 VTAIL.n134 VTAIL.n133 171.744
R74 VTAIL.n133 VTAIL.n123 171.744
R75 VTAIL.n126 VTAIL.n123 171.744
R76 VTAIL.n114 VTAIL.n113 171.744
R77 VTAIL.n113 VTAIL.n103 171.744
R78 VTAIL.n106 VTAIL.n103 171.744
R79 VTAIL.n94 VTAIL.n93 171.744
R80 VTAIL.n93 VTAIL.n83 171.744
R81 VTAIL.n86 VTAIL.n83 171.744
R82 VTAIL.n74 VTAIL.n73 171.744
R83 VTAIL.n73 VTAIL.n63 171.744
R84 VTAIL.n66 VTAIL.n63 171.744
R85 VTAIL.n146 VTAIL.t4 85.8723
R86 VTAIL.n6 VTAIL.t5 85.8723
R87 VTAIL.n26 VTAIL.t1 85.8723
R88 VTAIL.n46 VTAIL.t3 85.8723
R89 VTAIL.n126 VTAIL.t2 85.8723
R90 VTAIL.n106 VTAIL.t0 85.8723
R91 VTAIL.n86 VTAIL.t6 85.8723
R92 VTAIL.n66 VTAIL.t7 85.8723
R93 VTAIL.n159 VTAIL.n158 33.5429
R94 VTAIL.n19 VTAIL.n18 33.5429
R95 VTAIL.n39 VTAIL.n38 33.5429
R96 VTAIL.n59 VTAIL.n58 33.5429
R97 VTAIL.n139 VTAIL.n138 33.5429
R98 VTAIL.n119 VTAIL.n118 33.5429
R99 VTAIL.n99 VTAIL.n98 33.5429
R100 VTAIL.n79 VTAIL.n78 33.5429
R101 VTAIL.n159 VTAIL.n139 16.7548
R102 VTAIL.n79 VTAIL.n59 16.7548
R103 VTAIL.n147 VTAIL.n145 16.3201
R104 VTAIL.n7 VTAIL.n5 16.3201
R105 VTAIL.n27 VTAIL.n25 16.3201
R106 VTAIL.n47 VTAIL.n45 16.3201
R107 VTAIL.n127 VTAIL.n125 16.3201
R108 VTAIL.n107 VTAIL.n105 16.3201
R109 VTAIL.n87 VTAIL.n85 16.3201
R110 VTAIL.n67 VTAIL.n65 16.3201
R111 VTAIL.n148 VTAIL.n144 12.8005
R112 VTAIL.n8 VTAIL.n4 12.8005
R113 VTAIL.n28 VTAIL.n24 12.8005
R114 VTAIL.n48 VTAIL.n44 12.8005
R115 VTAIL.n128 VTAIL.n124 12.8005
R116 VTAIL.n108 VTAIL.n104 12.8005
R117 VTAIL.n88 VTAIL.n84 12.8005
R118 VTAIL.n68 VTAIL.n64 12.8005
R119 VTAIL.n152 VTAIL.n151 12.0247
R120 VTAIL.n12 VTAIL.n11 12.0247
R121 VTAIL.n32 VTAIL.n31 12.0247
R122 VTAIL.n52 VTAIL.n51 12.0247
R123 VTAIL.n132 VTAIL.n131 12.0247
R124 VTAIL.n112 VTAIL.n111 12.0247
R125 VTAIL.n92 VTAIL.n91 12.0247
R126 VTAIL.n72 VTAIL.n71 12.0247
R127 VTAIL.n155 VTAIL.n142 11.249
R128 VTAIL.n15 VTAIL.n2 11.249
R129 VTAIL.n35 VTAIL.n22 11.249
R130 VTAIL.n55 VTAIL.n42 11.249
R131 VTAIL.n135 VTAIL.n122 11.249
R132 VTAIL.n115 VTAIL.n102 11.249
R133 VTAIL.n95 VTAIL.n82 11.249
R134 VTAIL.n75 VTAIL.n62 11.249
R135 VTAIL.n156 VTAIL.n140 10.4732
R136 VTAIL.n16 VTAIL.n0 10.4732
R137 VTAIL.n36 VTAIL.n20 10.4732
R138 VTAIL.n56 VTAIL.n40 10.4732
R139 VTAIL.n136 VTAIL.n120 10.4732
R140 VTAIL.n116 VTAIL.n100 10.4732
R141 VTAIL.n96 VTAIL.n80 10.4732
R142 VTAIL.n76 VTAIL.n60 10.4732
R143 VTAIL.n158 VTAIL.n157 9.45567
R144 VTAIL.n18 VTAIL.n17 9.45567
R145 VTAIL.n38 VTAIL.n37 9.45567
R146 VTAIL.n58 VTAIL.n57 9.45567
R147 VTAIL.n138 VTAIL.n137 9.45567
R148 VTAIL.n118 VTAIL.n117 9.45567
R149 VTAIL.n98 VTAIL.n97 9.45567
R150 VTAIL.n78 VTAIL.n77 9.45567
R151 VTAIL.n157 VTAIL.n156 9.3005
R152 VTAIL.n142 VTAIL.n141 9.3005
R153 VTAIL.n151 VTAIL.n150 9.3005
R154 VTAIL.n149 VTAIL.n148 9.3005
R155 VTAIL.n17 VTAIL.n16 9.3005
R156 VTAIL.n2 VTAIL.n1 9.3005
R157 VTAIL.n11 VTAIL.n10 9.3005
R158 VTAIL.n9 VTAIL.n8 9.3005
R159 VTAIL.n37 VTAIL.n36 9.3005
R160 VTAIL.n22 VTAIL.n21 9.3005
R161 VTAIL.n31 VTAIL.n30 9.3005
R162 VTAIL.n29 VTAIL.n28 9.3005
R163 VTAIL.n57 VTAIL.n56 9.3005
R164 VTAIL.n42 VTAIL.n41 9.3005
R165 VTAIL.n51 VTAIL.n50 9.3005
R166 VTAIL.n49 VTAIL.n48 9.3005
R167 VTAIL.n137 VTAIL.n136 9.3005
R168 VTAIL.n122 VTAIL.n121 9.3005
R169 VTAIL.n131 VTAIL.n130 9.3005
R170 VTAIL.n129 VTAIL.n128 9.3005
R171 VTAIL.n117 VTAIL.n116 9.3005
R172 VTAIL.n102 VTAIL.n101 9.3005
R173 VTAIL.n111 VTAIL.n110 9.3005
R174 VTAIL.n109 VTAIL.n108 9.3005
R175 VTAIL.n97 VTAIL.n96 9.3005
R176 VTAIL.n82 VTAIL.n81 9.3005
R177 VTAIL.n91 VTAIL.n90 9.3005
R178 VTAIL.n89 VTAIL.n88 9.3005
R179 VTAIL.n77 VTAIL.n76 9.3005
R180 VTAIL.n62 VTAIL.n61 9.3005
R181 VTAIL.n71 VTAIL.n70 9.3005
R182 VTAIL.n69 VTAIL.n68 9.3005
R183 VTAIL.n149 VTAIL.n145 3.78097
R184 VTAIL.n9 VTAIL.n5 3.78097
R185 VTAIL.n29 VTAIL.n25 3.78097
R186 VTAIL.n49 VTAIL.n45 3.78097
R187 VTAIL.n129 VTAIL.n125 3.78097
R188 VTAIL.n109 VTAIL.n105 3.78097
R189 VTAIL.n89 VTAIL.n85 3.78097
R190 VTAIL.n69 VTAIL.n65 3.78097
R191 VTAIL.n158 VTAIL.n140 3.49141
R192 VTAIL.n18 VTAIL.n0 3.49141
R193 VTAIL.n38 VTAIL.n20 3.49141
R194 VTAIL.n58 VTAIL.n40 3.49141
R195 VTAIL.n138 VTAIL.n120 3.49141
R196 VTAIL.n118 VTAIL.n100 3.49141
R197 VTAIL.n98 VTAIL.n80 3.49141
R198 VTAIL.n78 VTAIL.n60 3.49141
R199 VTAIL.n156 VTAIL.n155 2.71565
R200 VTAIL.n16 VTAIL.n15 2.71565
R201 VTAIL.n36 VTAIL.n35 2.71565
R202 VTAIL.n56 VTAIL.n55 2.71565
R203 VTAIL.n136 VTAIL.n135 2.71565
R204 VTAIL.n116 VTAIL.n115 2.71565
R205 VTAIL.n96 VTAIL.n95 2.71565
R206 VTAIL.n76 VTAIL.n75 2.71565
R207 VTAIL.n152 VTAIL.n142 1.93989
R208 VTAIL.n12 VTAIL.n2 1.93989
R209 VTAIL.n32 VTAIL.n22 1.93989
R210 VTAIL.n52 VTAIL.n42 1.93989
R211 VTAIL.n132 VTAIL.n122 1.93989
R212 VTAIL.n112 VTAIL.n102 1.93989
R213 VTAIL.n92 VTAIL.n82 1.93989
R214 VTAIL.n72 VTAIL.n62 1.93989
R215 VTAIL.n151 VTAIL.n144 1.16414
R216 VTAIL.n11 VTAIL.n4 1.16414
R217 VTAIL.n31 VTAIL.n24 1.16414
R218 VTAIL.n51 VTAIL.n44 1.16414
R219 VTAIL.n131 VTAIL.n124 1.16414
R220 VTAIL.n111 VTAIL.n104 1.16414
R221 VTAIL.n91 VTAIL.n84 1.16414
R222 VTAIL.n71 VTAIL.n64 1.16414
R223 VTAIL.n99 VTAIL.n79 1.01774
R224 VTAIL.n139 VTAIL.n119 1.01774
R225 VTAIL.n59 VTAIL.n39 1.01774
R226 VTAIL VTAIL.n19 0.56731
R227 VTAIL.n119 VTAIL.n99 0.470328
R228 VTAIL.n39 VTAIL.n19 0.470328
R229 VTAIL VTAIL.n159 0.450931
R230 VTAIL.n148 VTAIL.n147 0.388379
R231 VTAIL.n8 VTAIL.n7 0.388379
R232 VTAIL.n28 VTAIL.n27 0.388379
R233 VTAIL.n48 VTAIL.n47 0.388379
R234 VTAIL.n128 VTAIL.n127 0.388379
R235 VTAIL.n108 VTAIL.n107 0.388379
R236 VTAIL.n88 VTAIL.n87 0.388379
R237 VTAIL.n68 VTAIL.n67 0.388379
R238 VTAIL.n150 VTAIL.n149 0.155672
R239 VTAIL.n150 VTAIL.n141 0.155672
R240 VTAIL.n157 VTAIL.n141 0.155672
R241 VTAIL.n10 VTAIL.n9 0.155672
R242 VTAIL.n10 VTAIL.n1 0.155672
R243 VTAIL.n17 VTAIL.n1 0.155672
R244 VTAIL.n30 VTAIL.n29 0.155672
R245 VTAIL.n30 VTAIL.n21 0.155672
R246 VTAIL.n37 VTAIL.n21 0.155672
R247 VTAIL.n50 VTAIL.n49 0.155672
R248 VTAIL.n50 VTAIL.n41 0.155672
R249 VTAIL.n57 VTAIL.n41 0.155672
R250 VTAIL.n137 VTAIL.n121 0.155672
R251 VTAIL.n130 VTAIL.n121 0.155672
R252 VTAIL.n130 VTAIL.n129 0.155672
R253 VTAIL.n117 VTAIL.n101 0.155672
R254 VTAIL.n110 VTAIL.n101 0.155672
R255 VTAIL.n110 VTAIL.n109 0.155672
R256 VTAIL.n97 VTAIL.n81 0.155672
R257 VTAIL.n90 VTAIL.n81 0.155672
R258 VTAIL.n90 VTAIL.n89 0.155672
R259 VTAIL.n77 VTAIL.n61 0.155672
R260 VTAIL.n70 VTAIL.n61 0.155672
R261 VTAIL.n70 VTAIL.n69 0.155672
R262 VP.n1 VP.t2 178.356
R263 VP.n1 VP.t1 178.305
R264 VP.n6 VP.n5 161.3
R265 VP.n4 VP.n0 161.3
R266 VP.n3 VP.n2 161.3
R267 VP.n3 VP.t0 157.359
R268 VP.n5 VP.t3 157.359
R269 VP.n2 VP.n1 79.5106
R270 VP.n4 VP.n3 24.1005
R271 VP.n5 VP.n4 24.1005
R272 VP.n2 VP.n0 0.189894
R273 VP.n6 VP.n0 0.189894
R274 VP VP.n6 0.0516364
R275 VDD1 VDD1.n1 145.588
R276 VDD1 VDD1.n0 114.984
R277 VDD1.n0 VDD1.t1 8.3138
R278 VDD1.n0 VDD1.t2 8.3138
R279 VDD1.n1 VDD1.t3 8.3138
R280 VDD1.n1 VDD1.t0 8.3138
R281 B.n186 B.n57 585
R282 B.n185 B.n184 585
R283 B.n183 B.n58 585
R284 B.n182 B.n181 585
R285 B.n180 B.n59 585
R286 B.n179 B.n178 585
R287 B.n177 B.n60 585
R288 B.n176 B.n175 585
R289 B.n174 B.n61 585
R290 B.n173 B.n172 585
R291 B.n171 B.n62 585
R292 B.n170 B.n169 585
R293 B.n168 B.n63 585
R294 B.n167 B.n166 585
R295 B.n165 B.n64 585
R296 B.n164 B.n163 585
R297 B.n162 B.n65 585
R298 B.n161 B.n160 585
R299 B.n159 B.n158 585
R300 B.n157 B.n69 585
R301 B.n156 B.n155 585
R302 B.n154 B.n70 585
R303 B.n153 B.n152 585
R304 B.n151 B.n71 585
R305 B.n150 B.n149 585
R306 B.n148 B.n72 585
R307 B.n147 B.n146 585
R308 B.n144 B.n73 585
R309 B.n143 B.n142 585
R310 B.n141 B.n76 585
R311 B.n140 B.n139 585
R312 B.n138 B.n77 585
R313 B.n137 B.n136 585
R314 B.n135 B.n78 585
R315 B.n134 B.n133 585
R316 B.n132 B.n79 585
R317 B.n131 B.n130 585
R318 B.n129 B.n80 585
R319 B.n128 B.n127 585
R320 B.n126 B.n81 585
R321 B.n125 B.n124 585
R322 B.n123 B.n82 585
R323 B.n122 B.n121 585
R324 B.n120 B.n83 585
R325 B.n119 B.n118 585
R326 B.n188 B.n187 585
R327 B.n189 B.n56 585
R328 B.n191 B.n190 585
R329 B.n192 B.n55 585
R330 B.n194 B.n193 585
R331 B.n195 B.n54 585
R332 B.n197 B.n196 585
R333 B.n198 B.n53 585
R334 B.n200 B.n199 585
R335 B.n201 B.n52 585
R336 B.n203 B.n202 585
R337 B.n204 B.n51 585
R338 B.n206 B.n205 585
R339 B.n207 B.n50 585
R340 B.n209 B.n208 585
R341 B.n210 B.n49 585
R342 B.n212 B.n211 585
R343 B.n213 B.n48 585
R344 B.n215 B.n214 585
R345 B.n216 B.n47 585
R346 B.n218 B.n217 585
R347 B.n219 B.n46 585
R348 B.n221 B.n220 585
R349 B.n222 B.n45 585
R350 B.n224 B.n223 585
R351 B.n225 B.n44 585
R352 B.n227 B.n226 585
R353 B.n228 B.n43 585
R354 B.n230 B.n229 585
R355 B.n231 B.n42 585
R356 B.n233 B.n232 585
R357 B.n234 B.n41 585
R358 B.n236 B.n235 585
R359 B.n237 B.n40 585
R360 B.n239 B.n238 585
R361 B.n240 B.n39 585
R362 B.n242 B.n241 585
R363 B.n243 B.n38 585
R364 B.n312 B.n11 585
R365 B.n311 B.n310 585
R366 B.n309 B.n12 585
R367 B.n308 B.n307 585
R368 B.n306 B.n13 585
R369 B.n305 B.n304 585
R370 B.n303 B.n14 585
R371 B.n302 B.n301 585
R372 B.n300 B.n15 585
R373 B.n299 B.n298 585
R374 B.n297 B.n16 585
R375 B.n296 B.n295 585
R376 B.n294 B.n17 585
R377 B.n293 B.n292 585
R378 B.n291 B.n18 585
R379 B.n290 B.n289 585
R380 B.n288 B.n19 585
R381 B.n287 B.n286 585
R382 B.n285 B.n284 585
R383 B.n283 B.n23 585
R384 B.n282 B.n281 585
R385 B.n280 B.n24 585
R386 B.n279 B.n278 585
R387 B.n277 B.n25 585
R388 B.n276 B.n275 585
R389 B.n274 B.n26 585
R390 B.n273 B.n272 585
R391 B.n270 B.n27 585
R392 B.n269 B.n268 585
R393 B.n267 B.n30 585
R394 B.n266 B.n265 585
R395 B.n264 B.n31 585
R396 B.n263 B.n262 585
R397 B.n261 B.n32 585
R398 B.n260 B.n259 585
R399 B.n258 B.n33 585
R400 B.n257 B.n256 585
R401 B.n255 B.n34 585
R402 B.n254 B.n253 585
R403 B.n252 B.n35 585
R404 B.n251 B.n250 585
R405 B.n249 B.n36 585
R406 B.n248 B.n247 585
R407 B.n246 B.n37 585
R408 B.n245 B.n244 585
R409 B.n314 B.n313 585
R410 B.n315 B.n10 585
R411 B.n317 B.n316 585
R412 B.n318 B.n9 585
R413 B.n320 B.n319 585
R414 B.n321 B.n8 585
R415 B.n323 B.n322 585
R416 B.n324 B.n7 585
R417 B.n326 B.n325 585
R418 B.n327 B.n6 585
R419 B.n329 B.n328 585
R420 B.n330 B.n5 585
R421 B.n332 B.n331 585
R422 B.n333 B.n4 585
R423 B.n335 B.n334 585
R424 B.n336 B.n3 585
R425 B.n338 B.n337 585
R426 B.n339 B.n0 585
R427 B.n2 B.n1 585
R428 B.n93 B.n92 585
R429 B.n95 B.n94 585
R430 B.n96 B.n91 585
R431 B.n98 B.n97 585
R432 B.n99 B.n90 585
R433 B.n101 B.n100 585
R434 B.n102 B.n89 585
R435 B.n104 B.n103 585
R436 B.n105 B.n88 585
R437 B.n107 B.n106 585
R438 B.n108 B.n87 585
R439 B.n110 B.n109 585
R440 B.n111 B.n86 585
R441 B.n113 B.n112 585
R442 B.n114 B.n85 585
R443 B.n116 B.n115 585
R444 B.n117 B.n84 585
R445 B.n118 B.n117 521.33
R446 B.n188 B.n57 521.33
R447 B.n244 B.n243 521.33
R448 B.n314 B.n11 521.33
R449 B.n74 B.t3 312.649
R450 B.n66 B.t9 312.649
R451 B.n28 B.t6 312.649
R452 B.n20 B.t0 312.649
R453 B.n66 B.t10 256.769
R454 B.n28 B.t8 256.769
R455 B.n74 B.t4 256.769
R456 B.n20 B.t2 256.769
R457 B.n341 B.n340 256.663
R458 B.n340 B.n339 235.042
R459 B.n340 B.n2 235.042
R460 B.n67 B.t11 233.885
R461 B.n29 B.t7 233.885
R462 B.n75 B.t5 233.883
R463 B.n21 B.t1 233.883
R464 B.n118 B.n83 163.367
R465 B.n122 B.n83 163.367
R466 B.n123 B.n122 163.367
R467 B.n124 B.n123 163.367
R468 B.n124 B.n81 163.367
R469 B.n128 B.n81 163.367
R470 B.n129 B.n128 163.367
R471 B.n130 B.n129 163.367
R472 B.n130 B.n79 163.367
R473 B.n134 B.n79 163.367
R474 B.n135 B.n134 163.367
R475 B.n136 B.n135 163.367
R476 B.n136 B.n77 163.367
R477 B.n140 B.n77 163.367
R478 B.n141 B.n140 163.367
R479 B.n142 B.n141 163.367
R480 B.n142 B.n73 163.367
R481 B.n147 B.n73 163.367
R482 B.n148 B.n147 163.367
R483 B.n149 B.n148 163.367
R484 B.n149 B.n71 163.367
R485 B.n153 B.n71 163.367
R486 B.n154 B.n153 163.367
R487 B.n155 B.n154 163.367
R488 B.n155 B.n69 163.367
R489 B.n159 B.n69 163.367
R490 B.n160 B.n159 163.367
R491 B.n160 B.n65 163.367
R492 B.n164 B.n65 163.367
R493 B.n165 B.n164 163.367
R494 B.n166 B.n165 163.367
R495 B.n166 B.n63 163.367
R496 B.n170 B.n63 163.367
R497 B.n171 B.n170 163.367
R498 B.n172 B.n171 163.367
R499 B.n172 B.n61 163.367
R500 B.n176 B.n61 163.367
R501 B.n177 B.n176 163.367
R502 B.n178 B.n177 163.367
R503 B.n178 B.n59 163.367
R504 B.n182 B.n59 163.367
R505 B.n183 B.n182 163.367
R506 B.n184 B.n183 163.367
R507 B.n184 B.n57 163.367
R508 B.n243 B.n242 163.367
R509 B.n242 B.n39 163.367
R510 B.n238 B.n39 163.367
R511 B.n238 B.n237 163.367
R512 B.n237 B.n236 163.367
R513 B.n236 B.n41 163.367
R514 B.n232 B.n41 163.367
R515 B.n232 B.n231 163.367
R516 B.n231 B.n230 163.367
R517 B.n230 B.n43 163.367
R518 B.n226 B.n43 163.367
R519 B.n226 B.n225 163.367
R520 B.n225 B.n224 163.367
R521 B.n224 B.n45 163.367
R522 B.n220 B.n45 163.367
R523 B.n220 B.n219 163.367
R524 B.n219 B.n218 163.367
R525 B.n218 B.n47 163.367
R526 B.n214 B.n47 163.367
R527 B.n214 B.n213 163.367
R528 B.n213 B.n212 163.367
R529 B.n212 B.n49 163.367
R530 B.n208 B.n49 163.367
R531 B.n208 B.n207 163.367
R532 B.n207 B.n206 163.367
R533 B.n206 B.n51 163.367
R534 B.n202 B.n51 163.367
R535 B.n202 B.n201 163.367
R536 B.n201 B.n200 163.367
R537 B.n200 B.n53 163.367
R538 B.n196 B.n53 163.367
R539 B.n196 B.n195 163.367
R540 B.n195 B.n194 163.367
R541 B.n194 B.n55 163.367
R542 B.n190 B.n55 163.367
R543 B.n190 B.n189 163.367
R544 B.n189 B.n188 163.367
R545 B.n310 B.n11 163.367
R546 B.n310 B.n309 163.367
R547 B.n309 B.n308 163.367
R548 B.n308 B.n13 163.367
R549 B.n304 B.n13 163.367
R550 B.n304 B.n303 163.367
R551 B.n303 B.n302 163.367
R552 B.n302 B.n15 163.367
R553 B.n298 B.n15 163.367
R554 B.n298 B.n297 163.367
R555 B.n297 B.n296 163.367
R556 B.n296 B.n17 163.367
R557 B.n292 B.n17 163.367
R558 B.n292 B.n291 163.367
R559 B.n291 B.n290 163.367
R560 B.n290 B.n19 163.367
R561 B.n286 B.n19 163.367
R562 B.n286 B.n285 163.367
R563 B.n285 B.n23 163.367
R564 B.n281 B.n23 163.367
R565 B.n281 B.n280 163.367
R566 B.n280 B.n279 163.367
R567 B.n279 B.n25 163.367
R568 B.n275 B.n25 163.367
R569 B.n275 B.n274 163.367
R570 B.n274 B.n273 163.367
R571 B.n273 B.n27 163.367
R572 B.n268 B.n27 163.367
R573 B.n268 B.n267 163.367
R574 B.n267 B.n266 163.367
R575 B.n266 B.n31 163.367
R576 B.n262 B.n31 163.367
R577 B.n262 B.n261 163.367
R578 B.n261 B.n260 163.367
R579 B.n260 B.n33 163.367
R580 B.n256 B.n33 163.367
R581 B.n256 B.n255 163.367
R582 B.n255 B.n254 163.367
R583 B.n254 B.n35 163.367
R584 B.n250 B.n35 163.367
R585 B.n250 B.n249 163.367
R586 B.n249 B.n248 163.367
R587 B.n248 B.n37 163.367
R588 B.n244 B.n37 163.367
R589 B.n315 B.n314 163.367
R590 B.n316 B.n315 163.367
R591 B.n316 B.n9 163.367
R592 B.n320 B.n9 163.367
R593 B.n321 B.n320 163.367
R594 B.n322 B.n321 163.367
R595 B.n322 B.n7 163.367
R596 B.n326 B.n7 163.367
R597 B.n327 B.n326 163.367
R598 B.n328 B.n327 163.367
R599 B.n328 B.n5 163.367
R600 B.n332 B.n5 163.367
R601 B.n333 B.n332 163.367
R602 B.n334 B.n333 163.367
R603 B.n334 B.n3 163.367
R604 B.n338 B.n3 163.367
R605 B.n339 B.n338 163.367
R606 B.n93 B.n2 163.367
R607 B.n94 B.n93 163.367
R608 B.n94 B.n91 163.367
R609 B.n98 B.n91 163.367
R610 B.n99 B.n98 163.367
R611 B.n100 B.n99 163.367
R612 B.n100 B.n89 163.367
R613 B.n104 B.n89 163.367
R614 B.n105 B.n104 163.367
R615 B.n106 B.n105 163.367
R616 B.n106 B.n87 163.367
R617 B.n110 B.n87 163.367
R618 B.n111 B.n110 163.367
R619 B.n112 B.n111 163.367
R620 B.n112 B.n85 163.367
R621 B.n116 B.n85 163.367
R622 B.n117 B.n116 163.367
R623 B.n145 B.n75 59.5399
R624 B.n68 B.n67 59.5399
R625 B.n271 B.n29 59.5399
R626 B.n22 B.n21 59.5399
R627 B.n313 B.n312 33.8737
R628 B.n245 B.n38 33.8737
R629 B.n187 B.n186 33.8737
R630 B.n119 B.n84 33.8737
R631 B.n75 B.n74 22.8853
R632 B.n67 B.n66 22.8853
R633 B.n29 B.n28 22.8853
R634 B.n21 B.n20 22.8853
R635 B B.n341 18.0485
R636 B.n313 B.n10 10.6151
R637 B.n317 B.n10 10.6151
R638 B.n318 B.n317 10.6151
R639 B.n319 B.n318 10.6151
R640 B.n319 B.n8 10.6151
R641 B.n323 B.n8 10.6151
R642 B.n324 B.n323 10.6151
R643 B.n325 B.n324 10.6151
R644 B.n325 B.n6 10.6151
R645 B.n329 B.n6 10.6151
R646 B.n330 B.n329 10.6151
R647 B.n331 B.n330 10.6151
R648 B.n331 B.n4 10.6151
R649 B.n335 B.n4 10.6151
R650 B.n336 B.n335 10.6151
R651 B.n337 B.n336 10.6151
R652 B.n337 B.n0 10.6151
R653 B.n312 B.n311 10.6151
R654 B.n311 B.n12 10.6151
R655 B.n307 B.n12 10.6151
R656 B.n307 B.n306 10.6151
R657 B.n306 B.n305 10.6151
R658 B.n305 B.n14 10.6151
R659 B.n301 B.n14 10.6151
R660 B.n301 B.n300 10.6151
R661 B.n300 B.n299 10.6151
R662 B.n299 B.n16 10.6151
R663 B.n295 B.n16 10.6151
R664 B.n295 B.n294 10.6151
R665 B.n294 B.n293 10.6151
R666 B.n293 B.n18 10.6151
R667 B.n289 B.n18 10.6151
R668 B.n289 B.n288 10.6151
R669 B.n288 B.n287 10.6151
R670 B.n284 B.n283 10.6151
R671 B.n283 B.n282 10.6151
R672 B.n282 B.n24 10.6151
R673 B.n278 B.n24 10.6151
R674 B.n278 B.n277 10.6151
R675 B.n277 B.n276 10.6151
R676 B.n276 B.n26 10.6151
R677 B.n272 B.n26 10.6151
R678 B.n270 B.n269 10.6151
R679 B.n269 B.n30 10.6151
R680 B.n265 B.n30 10.6151
R681 B.n265 B.n264 10.6151
R682 B.n264 B.n263 10.6151
R683 B.n263 B.n32 10.6151
R684 B.n259 B.n32 10.6151
R685 B.n259 B.n258 10.6151
R686 B.n258 B.n257 10.6151
R687 B.n257 B.n34 10.6151
R688 B.n253 B.n34 10.6151
R689 B.n253 B.n252 10.6151
R690 B.n252 B.n251 10.6151
R691 B.n251 B.n36 10.6151
R692 B.n247 B.n36 10.6151
R693 B.n247 B.n246 10.6151
R694 B.n246 B.n245 10.6151
R695 B.n241 B.n38 10.6151
R696 B.n241 B.n240 10.6151
R697 B.n240 B.n239 10.6151
R698 B.n239 B.n40 10.6151
R699 B.n235 B.n40 10.6151
R700 B.n235 B.n234 10.6151
R701 B.n234 B.n233 10.6151
R702 B.n233 B.n42 10.6151
R703 B.n229 B.n42 10.6151
R704 B.n229 B.n228 10.6151
R705 B.n228 B.n227 10.6151
R706 B.n227 B.n44 10.6151
R707 B.n223 B.n44 10.6151
R708 B.n223 B.n222 10.6151
R709 B.n222 B.n221 10.6151
R710 B.n221 B.n46 10.6151
R711 B.n217 B.n46 10.6151
R712 B.n217 B.n216 10.6151
R713 B.n216 B.n215 10.6151
R714 B.n215 B.n48 10.6151
R715 B.n211 B.n48 10.6151
R716 B.n211 B.n210 10.6151
R717 B.n210 B.n209 10.6151
R718 B.n209 B.n50 10.6151
R719 B.n205 B.n50 10.6151
R720 B.n205 B.n204 10.6151
R721 B.n204 B.n203 10.6151
R722 B.n203 B.n52 10.6151
R723 B.n199 B.n52 10.6151
R724 B.n199 B.n198 10.6151
R725 B.n198 B.n197 10.6151
R726 B.n197 B.n54 10.6151
R727 B.n193 B.n54 10.6151
R728 B.n193 B.n192 10.6151
R729 B.n192 B.n191 10.6151
R730 B.n191 B.n56 10.6151
R731 B.n187 B.n56 10.6151
R732 B.n92 B.n1 10.6151
R733 B.n95 B.n92 10.6151
R734 B.n96 B.n95 10.6151
R735 B.n97 B.n96 10.6151
R736 B.n97 B.n90 10.6151
R737 B.n101 B.n90 10.6151
R738 B.n102 B.n101 10.6151
R739 B.n103 B.n102 10.6151
R740 B.n103 B.n88 10.6151
R741 B.n107 B.n88 10.6151
R742 B.n108 B.n107 10.6151
R743 B.n109 B.n108 10.6151
R744 B.n109 B.n86 10.6151
R745 B.n113 B.n86 10.6151
R746 B.n114 B.n113 10.6151
R747 B.n115 B.n114 10.6151
R748 B.n115 B.n84 10.6151
R749 B.n120 B.n119 10.6151
R750 B.n121 B.n120 10.6151
R751 B.n121 B.n82 10.6151
R752 B.n125 B.n82 10.6151
R753 B.n126 B.n125 10.6151
R754 B.n127 B.n126 10.6151
R755 B.n127 B.n80 10.6151
R756 B.n131 B.n80 10.6151
R757 B.n132 B.n131 10.6151
R758 B.n133 B.n132 10.6151
R759 B.n133 B.n78 10.6151
R760 B.n137 B.n78 10.6151
R761 B.n138 B.n137 10.6151
R762 B.n139 B.n138 10.6151
R763 B.n139 B.n76 10.6151
R764 B.n143 B.n76 10.6151
R765 B.n144 B.n143 10.6151
R766 B.n146 B.n72 10.6151
R767 B.n150 B.n72 10.6151
R768 B.n151 B.n150 10.6151
R769 B.n152 B.n151 10.6151
R770 B.n152 B.n70 10.6151
R771 B.n156 B.n70 10.6151
R772 B.n157 B.n156 10.6151
R773 B.n158 B.n157 10.6151
R774 B.n162 B.n161 10.6151
R775 B.n163 B.n162 10.6151
R776 B.n163 B.n64 10.6151
R777 B.n167 B.n64 10.6151
R778 B.n168 B.n167 10.6151
R779 B.n169 B.n168 10.6151
R780 B.n169 B.n62 10.6151
R781 B.n173 B.n62 10.6151
R782 B.n174 B.n173 10.6151
R783 B.n175 B.n174 10.6151
R784 B.n175 B.n60 10.6151
R785 B.n179 B.n60 10.6151
R786 B.n180 B.n179 10.6151
R787 B.n181 B.n180 10.6151
R788 B.n181 B.n58 10.6151
R789 B.n185 B.n58 10.6151
R790 B.n186 B.n185 10.6151
R791 B.n341 B.n0 8.11757
R792 B.n341 B.n1 8.11757
R793 B.n284 B.n22 6.5566
R794 B.n272 B.n271 6.5566
R795 B.n146 B.n145 6.5566
R796 B.n158 B.n68 6.5566
R797 B.n287 B.n22 4.05904
R798 B.n271 B.n270 4.05904
R799 B.n145 B.n144 4.05904
R800 B.n161 B.n68 4.05904
C0 VN w_n1678_n1750# 2.35063f
C1 VTAIL VN 1.34856f
C2 VDD2 VP 0.287431f
C3 VP B 1.01878f
C4 VP VDD1 1.45537f
C5 VDD2 B 0.758106f
C6 VDD2 VDD1 0.601115f
C7 VP w_n1678_n1750# 2.56092f
C8 VTAIL VP 1.36266f
C9 VDD1 B 0.734336f
C10 VDD2 w_n1678_n1750# 0.893236f
C11 VDD2 VTAIL 3.15857f
C12 w_n1678_n1750# B 4.82304f
C13 VDD1 w_n1678_n1750# 0.876091f
C14 VTAIL VDD1 3.1161f
C15 VTAIL B 1.6773f
C16 VP VN 3.43471f
C17 VTAIL w_n1678_n1750# 2.0521f
C18 VDD2 VN 1.32013f
C19 VDD1 VN 0.151544f
C20 VN B 0.676522f
C21 VDD2 VSUBS 0.463743f
C22 VDD1 VSUBS 2.637449f
C23 VTAIL VSUBS 0.413518f
C24 VN VSUBS 4.00173f
C25 VP VSUBS 0.973639f
C26 B VSUBS 1.974743f
C27 w_n1678_n1750# VSUBS 36.9898f
C28 B.n0 VSUBS 0.006534f
C29 B.n1 VSUBS 0.006534f
C30 B.n2 VSUBS 0.009663f
C31 B.n3 VSUBS 0.007405f
C32 B.n4 VSUBS 0.007405f
C33 B.n5 VSUBS 0.007405f
C34 B.n6 VSUBS 0.007405f
C35 B.n7 VSUBS 0.007405f
C36 B.n8 VSUBS 0.007405f
C37 B.n9 VSUBS 0.007405f
C38 B.n10 VSUBS 0.007405f
C39 B.n11 VSUBS 0.01809f
C40 B.n12 VSUBS 0.007405f
C41 B.n13 VSUBS 0.007405f
C42 B.n14 VSUBS 0.007405f
C43 B.n15 VSUBS 0.007405f
C44 B.n16 VSUBS 0.007405f
C45 B.n17 VSUBS 0.007405f
C46 B.n18 VSUBS 0.007405f
C47 B.n19 VSUBS 0.007405f
C48 B.t1 VSUBS 0.059792f
C49 B.t2 VSUBS 0.0689f
C50 B.t0 VSUBS 0.159636f
C51 B.n20 VSUBS 0.126132f
C52 B.n21 VSUBS 0.112763f
C53 B.n22 VSUBS 0.017157f
C54 B.n23 VSUBS 0.007405f
C55 B.n24 VSUBS 0.007405f
C56 B.n25 VSUBS 0.007405f
C57 B.n26 VSUBS 0.007405f
C58 B.n27 VSUBS 0.007405f
C59 B.t7 VSUBS 0.059793f
C60 B.t8 VSUBS 0.068901f
C61 B.t6 VSUBS 0.159636f
C62 B.n28 VSUBS 0.126131f
C63 B.n29 VSUBS 0.112762f
C64 B.n30 VSUBS 0.007405f
C65 B.n31 VSUBS 0.007405f
C66 B.n32 VSUBS 0.007405f
C67 B.n33 VSUBS 0.007405f
C68 B.n34 VSUBS 0.007405f
C69 B.n35 VSUBS 0.007405f
C70 B.n36 VSUBS 0.007405f
C71 B.n37 VSUBS 0.007405f
C72 B.n38 VSUBS 0.017411f
C73 B.n39 VSUBS 0.007405f
C74 B.n40 VSUBS 0.007405f
C75 B.n41 VSUBS 0.007405f
C76 B.n42 VSUBS 0.007405f
C77 B.n43 VSUBS 0.007405f
C78 B.n44 VSUBS 0.007405f
C79 B.n45 VSUBS 0.007405f
C80 B.n46 VSUBS 0.007405f
C81 B.n47 VSUBS 0.007405f
C82 B.n48 VSUBS 0.007405f
C83 B.n49 VSUBS 0.007405f
C84 B.n50 VSUBS 0.007405f
C85 B.n51 VSUBS 0.007405f
C86 B.n52 VSUBS 0.007405f
C87 B.n53 VSUBS 0.007405f
C88 B.n54 VSUBS 0.007405f
C89 B.n55 VSUBS 0.007405f
C90 B.n56 VSUBS 0.007405f
C91 B.n57 VSUBS 0.01809f
C92 B.n58 VSUBS 0.007405f
C93 B.n59 VSUBS 0.007405f
C94 B.n60 VSUBS 0.007405f
C95 B.n61 VSUBS 0.007405f
C96 B.n62 VSUBS 0.007405f
C97 B.n63 VSUBS 0.007405f
C98 B.n64 VSUBS 0.007405f
C99 B.n65 VSUBS 0.007405f
C100 B.t11 VSUBS 0.059793f
C101 B.t10 VSUBS 0.068901f
C102 B.t9 VSUBS 0.159636f
C103 B.n66 VSUBS 0.126131f
C104 B.n67 VSUBS 0.112762f
C105 B.n68 VSUBS 0.017157f
C106 B.n69 VSUBS 0.007405f
C107 B.n70 VSUBS 0.007405f
C108 B.n71 VSUBS 0.007405f
C109 B.n72 VSUBS 0.007405f
C110 B.n73 VSUBS 0.007405f
C111 B.t5 VSUBS 0.059792f
C112 B.t4 VSUBS 0.0689f
C113 B.t3 VSUBS 0.159636f
C114 B.n74 VSUBS 0.126132f
C115 B.n75 VSUBS 0.112763f
C116 B.n76 VSUBS 0.007405f
C117 B.n77 VSUBS 0.007405f
C118 B.n78 VSUBS 0.007405f
C119 B.n79 VSUBS 0.007405f
C120 B.n80 VSUBS 0.007405f
C121 B.n81 VSUBS 0.007405f
C122 B.n82 VSUBS 0.007405f
C123 B.n83 VSUBS 0.007405f
C124 B.n84 VSUBS 0.017411f
C125 B.n85 VSUBS 0.007405f
C126 B.n86 VSUBS 0.007405f
C127 B.n87 VSUBS 0.007405f
C128 B.n88 VSUBS 0.007405f
C129 B.n89 VSUBS 0.007405f
C130 B.n90 VSUBS 0.007405f
C131 B.n91 VSUBS 0.007405f
C132 B.n92 VSUBS 0.007405f
C133 B.n93 VSUBS 0.007405f
C134 B.n94 VSUBS 0.007405f
C135 B.n95 VSUBS 0.007405f
C136 B.n96 VSUBS 0.007405f
C137 B.n97 VSUBS 0.007405f
C138 B.n98 VSUBS 0.007405f
C139 B.n99 VSUBS 0.007405f
C140 B.n100 VSUBS 0.007405f
C141 B.n101 VSUBS 0.007405f
C142 B.n102 VSUBS 0.007405f
C143 B.n103 VSUBS 0.007405f
C144 B.n104 VSUBS 0.007405f
C145 B.n105 VSUBS 0.007405f
C146 B.n106 VSUBS 0.007405f
C147 B.n107 VSUBS 0.007405f
C148 B.n108 VSUBS 0.007405f
C149 B.n109 VSUBS 0.007405f
C150 B.n110 VSUBS 0.007405f
C151 B.n111 VSUBS 0.007405f
C152 B.n112 VSUBS 0.007405f
C153 B.n113 VSUBS 0.007405f
C154 B.n114 VSUBS 0.007405f
C155 B.n115 VSUBS 0.007405f
C156 B.n116 VSUBS 0.007405f
C157 B.n117 VSUBS 0.017411f
C158 B.n118 VSUBS 0.01809f
C159 B.n119 VSUBS 0.01809f
C160 B.n120 VSUBS 0.007405f
C161 B.n121 VSUBS 0.007405f
C162 B.n122 VSUBS 0.007405f
C163 B.n123 VSUBS 0.007405f
C164 B.n124 VSUBS 0.007405f
C165 B.n125 VSUBS 0.007405f
C166 B.n126 VSUBS 0.007405f
C167 B.n127 VSUBS 0.007405f
C168 B.n128 VSUBS 0.007405f
C169 B.n129 VSUBS 0.007405f
C170 B.n130 VSUBS 0.007405f
C171 B.n131 VSUBS 0.007405f
C172 B.n132 VSUBS 0.007405f
C173 B.n133 VSUBS 0.007405f
C174 B.n134 VSUBS 0.007405f
C175 B.n135 VSUBS 0.007405f
C176 B.n136 VSUBS 0.007405f
C177 B.n137 VSUBS 0.007405f
C178 B.n138 VSUBS 0.007405f
C179 B.n139 VSUBS 0.007405f
C180 B.n140 VSUBS 0.007405f
C181 B.n141 VSUBS 0.007405f
C182 B.n142 VSUBS 0.007405f
C183 B.n143 VSUBS 0.007405f
C184 B.n144 VSUBS 0.005118f
C185 B.n145 VSUBS 0.017157f
C186 B.n146 VSUBS 0.005989f
C187 B.n147 VSUBS 0.007405f
C188 B.n148 VSUBS 0.007405f
C189 B.n149 VSUBS 0.007405f
C190 B.n150 VSUBS 0.007405f
C191 B.n151 VSUBS 0.007405f
C192 B.n152 VSUBS 0.007405f
C193 B.n153 VSUBS 0.007405f
C194 B.n154 VSUBS 0.007405f
C195 B.n155 VSUBS 0.007405f
C196 B.n156 VSUBS 0.007405f
C197 B.n157 VSUBS 0.007405f
C198 B.n158 VSUBS 0.005989f
C199 B.n159 VSUBS 0.007405f
C200 B.n160 VSUBS 0.007405f
C201 B.n161 VSUBS 0.005118f
C202 B.n162 VSUBS 0.007405f
C203 B.n163 VSUBS 0.007405f
C204 B.n164 VSUBS 0.007405f
C205 B.n165 VSUBS 0.007405f
C206 B.n166 VSUBS 0.007405f
C207 B.n167 VSUBS 0.007405f
C208 B.n168 VSUBS 0.007405f
C209 B.n169 VSUBS 0.007405f
C210 B.n170 VSUBS 0.007405f
C211 B.n171 VSUBS 0.007405f
C212 B.n172 VSUBS 0.007405f
C213 B.n173 VSUBS 0.007405f
C214 B.n174 VSUBS 0.007405f
C215 B.n175 VSUBS 0.007405f
C216 B.n176 VSUBS 0.007405f
C217 B.n177 VSUBS 0.007405f
C218 B.n178 VSUBS 0.007405f
C219 B.n179 VSUBS 0.007405f
C220 B.n180 VSUBS 0.007405f
C221 B.n181 VSUBS 0.007405f
C222 B.n182 VSUBS 0.007405f
C223 B.n183 VSUBS 0.007405f
C224 B.n184 VSUBS 0.007405f
C225 B.n185 VSUBS 0.007405f
C226 B.n186 VSUBS 0.017246f
C227 B.n187 VSUBS 0.018254f
C228 B.n188 VSUBS 0.017411f
C229 B.n189 VSUBS 0.007405f
C230 B.n190 VSUBS 0.007405f
C231 B.n191 VSUBS 0.007405f
C232 B.n192 VSUBS 0.007405f
C233 B.n193 VSUBS 0.007405f
C234 B.n194 VSUBS 0.007405f
C235 B.n195 VSUBS 0.007405f
C236 B.n196 VSUBS 0.007405f
C237 B.n197 VSUBS 0.007405f
C238 B.n198 VSUBS 0.007405f
C239 B.n199 VSUBS 0.007405f
C240 B.n200 VSUBS 0.007405f
C241 B.n201 VSUBS 0.007405f
C242 B.n202 VSUBS 0.007405f
C243 B.n203 VSUBS 0.007405f
C244 B.n204 VSUBS 0.007405f
C245 B.n205 VSUBS 0.007405f
C246 B.n206 VSUBS 0.007405f
C247 B.n207 VSUBS 0.007405f
C248 B.n208 VSUBS 0.007405f
C249 B.n209 VSUBS 0.007405f
C250 B.n210 VSUBS 0.007405f
C251 B.n211 VSUBS 0.007405f
C252 B.n212 VSUBS 0.007405f
C253 B.n213 VSUBS 0.007405f
C254 B.n214 VSUBS 0.007405f
C255 B.n215 VSUBS 0.007405f
C256 B.n216 VSUBS 0.007405f
C257 B.n217 VSUBS 0.007405f
C258 B.n218 VSUBS 0.007405f
C259 B.n219 VSUBS 0.007405f
C260 B.n220 VSUBS 0.007405f
C261 B.n221 VSUBS 0.007405f
C262 B.n222 VSUBS 0.007405f
C263 B.n223 VSUBS 0.007405f
C264 B.n224 VSUBS 0.007405f
C265 B.n225 VSUBS 0.007405f
C266 B.n226 VSUBS 0.007405f
C267 B.n227 VSUBS 0.007405f
C268 B.n228 VSUBS 0.007405f
C269 B.n229 VSUBS 0.007405f
C270 B.n230 VSUBS 0.007405f
C271 B.n231 VSUBS 0.007405f
C272 B.n232 VSUBS 0.007405f
C273 B.n233 VSUBS 0.007405f
C274 B.n234 VSUBS 0.007405f
C275 B.n235 VSUBS 0.007405f
C276 B.n236 VSUBS 0.007405f
C277 B.n237 VSUBS 0.007405f
C278 B.n238 VSUBS 0.007405f
C279 B.n239 VSUBS 0.007405f
C280 B.n240 VSUBS 0.007405f
C281 B.n241 VSUBS 0.007405f
C282 B.n242 VSUBS 0.007405f
C283 B.n243 VSUBS 0.017411f
C284 B.n244 VSUBS 0.01809f
C285 B.n245 VSUBS 0.01809f
C286 B.n246 VSUBS 0.007405f
C287 B.n247 VSUBS 0.007405f
C288 B.n248 VSUBS 0.007405f
C289 B.n249 VSUBS 0.007405f
C290 B.n250 VSUBS 0.007405f
C291 B.n251 VSUBS 0.007405f
C292 B.n252 VSUBS 0.007405f
C293 B.n253 VSUBS 0.007405f
C294 B.n254 VSUBS 0.007405f
C295 B.n255 VSUBS 0.007405f
C296 B.n256 VSUBS 0.007405f
C297 B.n257 VSUBS 0.007405f
C298 B.n258 VSUBS 0.007405f
C299 B.n259 VSUBS 0.007405f
C300 B.n260 VSUBS 0.007405f
C301 B.n261 VSUBS 0.007405f
C302 B.n262 VSUBS 0.007405f
C303 B.n263 VSUBS 0.007405f
C304 B.n264 VSUBS 0.007405f
C305 B.n265 VSUBS 0.007405f
C306 B.n266 VSUBS 0.007405f
C307 B.n267 VSUBS 0.007405f
C308 B.n268 VSUBS 0.007405f
C309 B.n269 VSUBS 0.007405f
C310 B.n270 VSUBS 0.005118f
C311 B.n271 VSUBS 0.017157f
C312 B.n272 VSUBS 0.005989f
C313 B.n273 VSUBS 0.007405f
C314 B.n274 VSUBS 0.007405f
C315 B.n275 VSUBS 0.007405f
C316 B.n276 VSUBS 0.007405f
C317 B.n277 VSUBS 0.007405f
C318 B.n278 VSUBS 0.007405f
C319 B.n279 VSUBS 0.007405f
C320 B.n280 VSUBS 0.007405f
C321 B.n281 VSUBS 0.007405f
C322 B.n282 VSUBS 0.007405f
C323 B.n283 VSUBS 0.007405f
C324 B.n284 VSUBS 0.005989f
C325 B.n285 VSUBS 0.007405f
C326 B.n286 VSUBS 0.007405f
C327 B.n287 VSUBS 0.005118f
C328 B.n288 VSUBS 0.007405f
C329 B.n289 VSUBS 0.007405f
C330 B.n290 VSUBS 0.007405f
C331 B.n291 VSUBS 0.007405f
C332 B.n292 VSUBS 0.007405f
C333 B.n293 VSUBS 0.007405f
C334 B.n294 VSUBS 0.007405f
C335 B.n295 VSUBS 0.007405f
C336 B.n296 VSUBS 0.007405f
C337 B.n297 VSUBS 0.007405f
C338 B.n298 VSUBS 0.007405f
C339 B.n299 VSUBS 0.007405f
C340 B.n300 VSUBS 0.007405f
C341 B.n301 VSUBS 0.007405f
C342 B.n302 VSUBS 0.007405f
C343 B.n303 VSUBS 0.007405f
C344 B.n304 VSUBS 0.007405f
C345 B.n305 VSUBS 0.007405f
C346 B.n306 VSUBS 0.007405f
C347 B.n307 VSUBS 0.007405f
C348 B.n308 VSUBS 0.007405f
C349 B.n309 VSUBS 0.007405f
C350 B.n310 VSUBS 0.007405f
C351 B.n311 VSUBS 0.007405f
C352 B.n312 VSUBS 0.01809f
C353 B.n313 VSUBS 0.017411f
C354 B.n314 VSUBS 0.017411f
C355 B.n315 VSUBS 0.007405f
C356 B.n316 VSUBS 0.007405f
C357 B.n317 VSUBS 0.007405f
C358 B.n318 VSUBS 0.007405f
C359 B.n319 VSUBS 0.007405f
C360 B.n320 VSUBS 0.007405f
C361 B.n321 VSUBS 0.007405f
C362 B.n322 VSUBS 0.007405f
C363 B.n323 VSUBS 0.007405f
C364 B.n324 VSUBS 0.007405f
C365 B.n325 VSUBS 0.007405f
C366 B.n326 VSUBS 0.007405f
C367 B.n327 VSUBS 0.007405f
C368 B.n328 VSUBS 0.007405f
C369 B.n329 VSUBS 0.007405f
C370 B.n330 VSUBS 0.007405f
C371 B.n331 VSUBS 0.007405f
C372 B.n332 VSUBS 0.007405f
C373 B.n333 VSUBS 0.007405f
C374 B.n334 VSUBS 0.007405f
C375 B.n335 VSUBS 0.007405f
C376 B.n336 VSUBS 0.007405f
C377 B.n337 VSUBS 0.007405f
C378 B.n338 VSUBS 0.007405f
C379 B.n339 VSUBS 0.009663f
C380 B.n340 VSUBS 0.010294f
C381 B.n341 VSUBS 0.02047f
C382 VDD1.t1 VSUBS 0.057113f
C383 VDD1.t2 VSUBS 0.057113f
C384 VDD1.n0 VSUBS 0.331492f
C385 VDD1.t3 VSUBS 0.057113f
C386 VDD1.t0 VSUBS 0.057113f
C387 VDD1.n1 VSUBS 0.51315f
C388 VP.n0 VSUBS 0.048096f
C389 VP.t1 VSUBS 0.501379f
C390 VP.t2 VSUBS 0.501465f
C391 VP.n1 VSUBS 1.11139f
C392 VP.n2 VSUBS 2.33178f
C393 VP.t0 VSUBS 0.472405f
C394 VP.n3 VSUBS 0.243178f
C395 VP.n4 VSUBS 0.010914f
C396 VP.t3 VSUBS 0.472405f
C397 VP.n5 VSUBS 0.243178f
C398 VP.n6 VSUBS 0.037272f
C399 VTAIL.n0 VSUBS 0.019805f
C400 VTAIL.n1 VSUBS 0.018451f
C401 VTAIL.n2 VSUBS 0.009915f
C402 VTAIL.n3 VSUBS 0.023435f
C403 VTAIL.n4 VSUBS 0.010498f
C404 VTAIL.n5 VSUBS 0.071148f
C405 VTAIL.t5 VSUBS 0.051658f
C406 VTAIL.n6 VSUBS 0.017576f
C407 VTAIL.n7 VSUBS 0.01474f
C408 VTAIL.n8 VSUBS 0.009915f
C409 VTAIL.n9 VSUBS 0.245936f
C410 VTAIL.n10 VSUBS 0.018451f
C411 VTAIL.n11 VSUBS 0.009915f
C412 VTAIL.n12 VSUBS 0.010498f
C413 VTAIL.n13 VSUBS 0.023435f
C414 VTAIL.n14 VSUBS 0.055138f
C415 VTAIL.n15 VSUBS 0.010498f
C416 VTAIL.n16 VSUBS 0.009915f
C417 VTAIL.n17 VSUBS 0.044413f
C418 VTAIL.n18 VSUBS 0.027711f
C419 VTAIL.n19 VSUBS 0.078386f
C420 VTAIL.n20 VSUBS 0.019805f
C421 VTAIL.n21 VSUBS 0.018451f
C422 VTAIL.n22 VSUBS 0.009915f
C423 VTAIL.n23 VSUBS 0.023435f
C424 VTAIL.n24 VSUBS 0.010498f
C425 VTAIL.n25 VSUBS 0.071148f
C426 VTAIL.t1 VSUBS 0.051658f
C427 VTAIL.n26 VSUBS 0.017576f
C428 VTAIL.n27 VSUBS 0.01474f
C429 VTAIL.n28 VSUBS 0.009915f
C430 VTAIL.n29 VSUBS 0.245936f
C431 VTAIL.n30 VSUBS 0.018451f
C432 VTAIL.n31 VSUBS 0.009915f
C433 VTAIL.n32 VSUBS 0.010498f
C434 VTAIL.n33 VSUBS 0.023435f
C435 VTAIL.n34 VSUBS 0.055138f
C436 VTAIL.n35 VSUBS 0.010498f
C437 VTAIL.n36 VSUBS 0.009915f
C438 VTAIL.n37 VSUBS 0.044413f
C439 VTAIL.n38 VSUBS 0.027711f
C440 VTAIL.n39 VSUBS 0.105165f
C441 VTAIL.n40 VSUBS 0.019805f
C442 VTAIL.n41 VSUBS 0.018451f
C443 VTAIL.n42 VSUBS 0.009915f
C444 VTAIL.n43 VSUBS 0.023435f
C445 VTAIL.n44 VSUBS 0.010498f
C446 VTAIL.n45 VSUBS 0.071148f
C447 VTAIL.t3 VSUBS 0.051658f
C448 VTAIL.n46 VSUBS 0.017576f
C449 VTAIL.n47 VSUBS 0.01474f
C450 VTAIL.n48 VSUBS 0.009915f
C451 VTAIL.n49 VSUBS 0.245936f
C452 VTAIL.n50 VSUBS 0.018451f
C453 VTAIL.n51 VSUBS 0.009915f
C454 VTAIL.n52 VSUBS 0.010498f
C455 VTAIL.n53 VSUBS 0.023435f
C456 VTAIL.n54 VSUBS 0.055138f
C457 VTAIL.n55 VSUBS 0.010498f
C458 VTAIL.n56 VSUBS 0.009915f
C459 VTAIL.n57 VSUBS 0.044413f
C460 VTAIL.n58 VSUBS 0.027711f
C461 VTAIL.n59 VSUBS 0.588739f
C462 VTAIL.n60 VSUBS 0.019805f
C463 VTAIL.n61 VSUBS 0.018451f
C464 VTAIL.n62 VSUBS 0.009915f
C465 VTAIL.n63 VSUBS 0.023435f
C466 VTAIL.n64 VSUBS 0.010498f
C467 VTAIL.n65 VSUBS 0.071148f
C468 VTAIL.t7 VSUBS 0.051658f
C469 VTAIL.n66 VSUBS 0.017576f
C470 VTAIL.n67 VSUBS 0.01474f
C471 VTAIL.n68 VSUBS 0.009915f
C472 VTAIL.n69 VSUBS 0.245936f
C473 VTAIL.n70 VSUBS 0.018451f
C474 VTAIL.n71 VSUBS 0.009915f
C475 VTAIL.n72 VSUBS 0.010498f
C476 VTAIL.n73 VSUBS 0.023435f
C477 VTAIL.n74 VSUBS 0.055138f
C478 VTAIL.n75 VSUBS 0.010498f
C479 VTAIL.n76 VSUBS 0.009915f
C480 VTAIL.n77 VSUBS 0.044413f
C481 VTAIL.n78 VSUBS 0.027711f
C482 VTAIL.n79 VSUBS 0.588739f
C483 VTAIL.n80 VSUBS 0.019805f
C484 VTAIL.n81 VSUBS 0.018451f
C485 VTAIL.n82 VSUBS 0.009915f
C486 VTAIL.n83 VSUBS 0.023435f
C487 VTAIL.n84 VSUBS 0.010498f
C488 VTAIL.n85 VSUBS 0.071148f
C489 VTAIL.t6 VSUBS 0.051658f
C490 VTAIL.n86 VSUBS 0.017576f
C491 VTAIL.n87 VSUBS 0.01474f
C492 VTAIL.n88 VSUBS 0.009915f
C493 VTAIL.n89 VSUBS 0.245936f
C494 VTAIL.n90 VSUBS 0.018451f
C495 VTAIL.n91 VSUBS 0.009915f
C496 VTAIL.n92 VSUBS 0.010498f
C497 VTAIL.n93 VSUBS 0.023435f
C498 VTAIL.n94 VSUBS 0.055138f
C499 VTAIL.n95 VSUBS 0.010498f
C500 VTAIL.n96 VSUBS 0.009915f
C501 VTAIL.n97 VSUBS 0.044413f
C502 VTAIL.n98 VSUBS 0.027711f
C503 VTAIL.n99 VSUBS 0.105165f
C504 VTAIL.n100 VSUBS 0.019805f
C505 VTAIL.n101 VSUBS 0.018451f
C506 VTAIL.n102 VSUBS 0.009915f
C507 VTAIL.n103 VSUBS 0.023435f
C508 VTAIL.n104 VSUBS 0.010498f
C509 VTAIL.n105 VSUBS 0.071148f
C510 VTAIL.t0 VSUBS 0.051658f
C511 VTAIL.n106 VSUBS 0.017576f
C512 VTAIL.n107 VSUBS 0.01474f
C513 VTAIL.n108 VSUBS 0.009915f
C514 VTAIL.n109 VSUBS 0.245936f
C515 VTAIL.n110 VSUBS 0.018451f
C516 VTAIL.n111 VSUBS 0.009915f
C517 VTAIL.n112 VSUBS 0.010498f
C518 VTAIL.n113 VSUBS 0.023435f
C519 VTAIL.n114 VSUBS 0.055138f
C520 VTAIL.n115 VSUBS 0.010498f
C521 VTAIL.n116 VSUBS 0.009915f
C522 VTAIL.n117 VSUBS 0.044413f
C523 VTAIL.n118 VSUBS 0.027711f
C524 VTAIL.n119 VSUBS 0.105165f
C525 VTAIL.n120 VSUBS 0.019805f
C526 VTAIL.n121 VSUBS 0.018451f
C527 VTAIL.n122 VSUBS 0.009915f
C528 VTAIL.n123 VSUBS 0.023435f
C529 VTAIL.n124 VSUBS 0.010498f
C530 VTAIL.n125 VSUBS 0.071148f
C531 VTAIL.t2 VSUBS 0.051658f
C532 VTAIL.n126 VSUBS 0.017576f
C533 VTAIL.n127 VSUBS 0.01474f
C534 VTAIL.n128 VSUBS 0.009915f
C535 VTAIL.n129 VSUBS 0.245936f
C536 VTAIL.n130 VSUBS 0.018451f
C537 VTAIL.n131 VSUBS 0.009915f
C538 VTAIL.n132 VSUBS 0.010498f
C539 VTAIL.n133 VSUBS 0.023435f
C540 VTAIL.n134 VSUBS 0.055138f
C541 VTAIL.n135 VSUBS 0.010498f
C542 VTAIL.n136 VSUBS 0.009915f
C543 VTAIL.n137 VSUBS 0.044413f
C544 VTAIL.n138 VSUBS 0.027711f
C545 VTAIL.n139 VSUBS 0.588739f
C546 VTAIL.n140 VSUBS 0.019805f
C547 VTAIL.n141 VSUBS 0.018451f
C548 VTAIL.n142 VSUBS 0.009915f
C549 VTAIL.n143 VSUBS 0.023435f
C550 VTAIL.n144 VSUBS 0.010498f
C551 VTAIL.n145 VSUBS 0.071148f
C552 VTAIL.t4 VSUBS 0.051658f
C553 VTAIL.n146 VSUBS 0.017576f
C554 VTAIL.n147 VSUBS 0.01474f
C555 VTAIL.n148 VSUBS 0.009915f
C556 VTAIL.n149 VSUBS 0.245936f
C557 VTAIL.n150 VSUBS 0.018451f
C558 VTAIL.n151 VSUBS 0.009915f
C559 VTAIL.n152 VSUBS 0.010498f
C560 VTAIL.n153 VSUBS 0.023435f
C561 VTAIL.n154 VSUBS 0.055138f
C562 VTAIL.n155 VSUBS 0.010498f
C563 VTAIL.n156 VSUBS 0.009915f
C564 VTAIL.n157 VSUBS 0.044413f
C565 VTAIL.n158 VSUBS 0.027711f
C566 VTAIL.n159 VSUBS 0.555041f
C567 VDD2.t1 VSUBS 0.060283f
C568 VDD2.t0 VSUBS 0.060283f
C569 VDD2.n0 VSUBS 0.530682f
C570 VDD2.t3 VSUBS 0.060283f
C571 VDD2.t2 VSUBS 0.060283f
C572 VDD2.n1 VSUBS 0.349715f
C573 VDD2.n2 VSUBS 2.01032f
C574 VN.t2 VSUBS 0.479348f
C575 VN.t3 VSUBS 0.479266f
C576 VN.n0 VSUBS 0.420367f
C577 VN.t1 VSUBS 0.479348f
C578 VN.t0 VSUBS 0.479266f
C579 VN.n1 VSUBS 1.07977f
.ends

