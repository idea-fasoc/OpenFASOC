* NGSPICE file created from opamp_sample_0005.ext - technology: sky130A

.subckt opamp_sample_0005 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 GND.t201 GND.t199 GND.t200 GND.t121 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X1 GND.t76 CS_BIAS.t20 VOUT.t29 GND.t62 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X2 GND.t198 GND.t196 GND.t197 GND.t99 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X3 VOUT.t37 GND.t214 VDD.t141 VDD.t98 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=1.5561 ps=8.76 w=3.99 l=3.26
X4 VN.t3 GND.t193 GND.t195 GND.t194 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X5 VDD.t93 VDD.t91 VDD.t92 VDD.t28 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X6 GND.t67 CS_BIAS.t21 VOUT.t28 GND.t45 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X7 VOUT.t27 CS_BIAS.t22 GND.t213 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=2.37
X8 GND.t29 CS_BIAS.t23 VOUT.t26 GND.t28 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X9 VOUT.t25 CS_BIAS.t24 GND.t47 GND.t10 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=2.37
X10 VOUT.t24 CS_BIAS.t25 GND.t27 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X11 GND.t192 GND.t189 GND.t191 GND.t190 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=0 ps=0 w=4.14 l=4.06
X12 GND.t188 GND.t186 GND.t187 GND.t121 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X13 a_n12854_10929# a_n12854_10929# a_n12854_10929# VDD.t1 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=1.7706 ps=10.64 w=2.27 l=5.93
X14 VOUT.t23 CS_BIAS.t26 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X15 GND.t75 CS_BIAS.t18 CS_BIAS.t19 GND.t62 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X16 a_n4580_9541.t12 GND.t178 GND.t179 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=5.93
X17 a_n7464_n776.t9 DIFFPAIR_BIAS.t10 GND.t83 GND.t82 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=4.06
X18 VOUT.t40 a_n4580_9541.t0 sky130_fd_pr__cap_mim_m3_1 l=10.72 w=5.27
X19 VDD.t140 GND.t215 a_n4580_9541.t8 VDD.t139 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=5.93
X20 VOUT.t41 a_n4580_9541.t0 sky130_fd_pr__cap_mim_m3_1 l=10.72 w=5.27
X21 GND.t66 CS_BIAS.t27 VOUT.t22 GND.t62 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X22 GND.t32 VN.t4 a_n7464_n776.t24 GND.t22 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=2.7963 ps=15.12 w=7.17 l=6.98
X23 VOUT.t21 CS_BIAS.t28 GND.t204 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=2.37
X24 VOUT.t31 GND.t216 VDD.t137 VDD.t126 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=1.5561 ps=8.76 w=3.99 l=3.26
X25 VOUT.t32 GND.t217 VDD.t138 VDD.t126 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=1.5561 ps=8.76 w=3.99 l=3.26
X26 VDD.t136 GND.t218 a_n11384_10929.t7 VDD.t135 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=5.93
X27 VDD.t90 VDD.t88 VDD.t89 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=5.93
X28 a_n7464_n776.t23 VN.t5 GND.t56 GND.t33 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X29 VOUT.t30 GND.t219 VDD.t134 VDD.t126 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=1.5561 ps=8.76 w=3.99 l=3.26
X30 GND.t42 VN.t6 a_n7464_n776.t22 GND.t4 sky130_fd_pr__nfet_01v8 ad=2.7963 pd=15.12 as=1.18305 ps=7.5 w=7.17 l=6.98
X31 GND.t185 GND.t183 GND.t184 GND.t125 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X32 GND.t211 VN.t7 a_n7464_n776.t21 GND.t84 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X33 GND.t44 VN.t8 a_n7464_n776.t20 GND.t43 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=2.7963 ps=15.12 w=7.17 l=6.98
X34 a_n7464_n776.t19 VN.t9 GND.t55 GND.t54 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X35 GND.t182 GND.t180 GND.t181 GND.t121 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X36 VN.t2 GND.t175 GND.t177 GND.t176 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X37 CS_BIAS.t17 CS_BIAS.t16 GND.t57 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=2.37
X38 VOUT.t20 CS_BIAS.t29 GND.t11 GND.t10 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=2.37
X39 VOUT.t35 GND.t220 VDD.t133 VDD.t98 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=1.5561 ps=8.76 w=3.99 l=3.26
X40 VP.t3 GND.t172 GND.t174 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X41 VDD.t87 VDD.t85 VDD.t86 VDD.t28 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X42 GND.t171 GND.t169 GND.t170 GND.t103 sky130_fd_pr__nfet_01v8 ad=2.7963 pd=15.12 as=0 ps=0 w=7.17 l=6.98
X43 VOUT.t42 a_n4580_9541.t0 sky130_fd_pr__cap_mim_m3_1 l=10.72 w=5.27
X44 CS_BIAS.t15 CS_BIAS.t14 GND.t53 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=2.37
X45 VDD.t84 VDD.t82 VDD.t83 VDD.t48 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X46 VOUT.t43 a_n4580_9541.t0 sky130_fd_pr__cap_mim_m3_1 l=10.72 w=5.27
X47 GND.t168 GND.t166 GND.t167 GND.t99 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X48 VDD.t81 VDD.t79 VDD.t80 VDD.t48 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X49 VDD.t78 VDD.t76 VDD.t77 VDD.t48 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X50 DIFFPAIR_BIAS.t9 DIFFPAIR_BIAS.t8 GND.t59 GND.t58 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=4.06
X51 VOUT.t34 GND.t221 VDD.t132 VDD.t126 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=1.5561 ps=8.76 w=3.99 l=3.26
X52 VDD.t75 VDD.t73 VDD.t74 VDD.t48 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X53 a_n7464_n776.t8 DIFFPAIR_BIAS.t11 GND.t81 GND.t80 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=4.06
X54 GND.t165 GND.t163 GND.t164 GND.t111 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X55 VOUT.t19 CS_BIAS.t30 GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=2.37
X56 VDD.t72 VDD.t70 VDD.t71 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=5.93
X57 a_n11384_10929.t11 GND.t161 GND.t162 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=5.93
X58 VDD.t69 VDD.t67 VDD.t68 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X59 VDD.t66 VDD.t64 VDD.t65 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=5.93
X60 VOUT.t18 CS_BIAS.t31 GND.t69 GND.t14 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=2.37
X61 VOUT.t17 CS_BIAS.t32 GND.t25 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X62 GND.t160 GND.t158 GND.t159 GND.t111 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X63 GND.t68 CS_BIAS.t33 VOUT.t16 GND.t45 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X64 VP.t2 GND.t155 GND.t157 GND.t156 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X65 a_n7464_n776.t7 DIFFPAIR_BIAS.t12 GND.t3 GND.t2 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=4.06
X66 GND.t154 GND.t152 GND.t153 GND.t125 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X67 GND.t87 VP.t4 a_n7464_n776.t14 GND.t37 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X68 a_n7464_n776.t13 VP.t5 GND.t86 GND.t35 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X69 VDD.t63 VDD.t60 VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=5.93
X70 VOUT.t15 CS_BIAS.t34 GND.t40 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=2.37
X71 GND.t73 CS_BIAS.t35 VOUT.t14 GND.t64 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X72 GND.t70 CS_BIAS.t12 CS_BIAS.t13 GND.t64 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X73 GND.t206 VN.t10 a_n7464_n776.t18 GND.t8 sky130_fd_pr__nfet_01v8 ad=2.7963 pd=15.12 as=1.18305 ps=7.5 w=7.17 l=6.98
X74 VDD.t59 VDD.t57 VDD.t58 VDD.t3 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X75 a_n11384_10929.t6 GND.t222 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=5.93
X76 VDD.t56 VDD.t54 VDD.t55 VDD.t3 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X77 CS_BIAS.t11 CS_BIAS.t10 GND.t212 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X78 GND.t151 GND.t149 GND.t150 GND.t99 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X79 GND.t97 GND.t96 a_n4580_9541.t11 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=5.93
X80 VDD.t53 VDD.t51 VDD.t52 VDD.t3 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X81 GND.t95 GND.t94 a_n11384_10929.t10 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=5.93
X82 GND.t148 GND.t146 GND.t147 GND.t111 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X83 VDD.t50 VDD.t47 VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X84 VDD.t129 GND.t223 a_n4580_9541.t7 VDD.t128 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=5.93
X85 VOUT.t38 GND.t224 VDD.t127 VDD.t126 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=1.5561 ps=8.76 w=3.99 l=3.26
X86 CS_BIAS.t9 CS_BIAS.t8 GND.t207 GND.t10 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=2.37
X87 VOUT.t13 CS_BIAS.t36 GND.t13 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X88 VOUT.t12 CS_BIAS.t37 GND.t74 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X89 GND.t41 CS_BIAS.t38 VOUT.t11 GND.t28 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X90 GND.t145 GND.t143 GND.t144 GND.t125 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X91 VDD.t46 VDD.t43 VDD.t45 VDD.t44 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=5.93
X92 VDD.t125 GND.t225 a_n11384_10929.t5 VDD.t124 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=5.93
X93 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.t6 GND.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=4.06
X94 VDD.t42 VDD.t40 VDD.t41 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X95 GND.t72 CS_BIAS.t39 VOUT.t10 GND.t28 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X96 GND.t142 GND.t141 a_n11384_10929.t9 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=5.93
X97 VDD.t39 VDD.t37 VDD.t38 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=5.93
X98 VOUT.t9 CS_BIAS.t40 GND.t24 GND.t10 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=2.37
X99 a_n7464_n776.t17 VN.t11 GND.t31 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X100 GND.t85 VP.t6 a_n7464_n776.t12 GND.t84 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X101 VOUT.t44 a_n4580_9541.t0 sky130_fd_pr__cap_mim_m3_1 l=10.72 w=5.27
X102 GND.t79 VP.t7 a_n7464_n776.t11 GND.t43 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=2.7963 ps=15.12 w=7.17 l=6.98
X103 VDD.t122 GND.t226 a_n11384_10929.t4 VDD.t121 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=5.93
X104 VOUT.t45 a_n4580_9541.t0 sky130_fd_pr__cap_mim_m3_1 l=10.72 w=5.27
X105 GND.t140 GND.t138 GND.t139 GND.t89 sky130_fd_pr__nfet_01v8 ad=2.7963 pd=15.12 as=0 ps=0 w=7.17 l=6.98
X106 a_n7464_n776.t10 VP.t8 GND.t78 GND.t54 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X107 GND.t137 GND.t135 VN.t1 GND.t136 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X108 GND.t132 GND.t131 a_n4580_9541.t10 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=5.93
X109 a_n11384_10929.t8 GND.t133 GND.t134 VDD.t119 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=5.93
X110 VOUT.t8 CS_BIAS.t41 GND.t71 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=2.37
X111 GND.t63 CS_BIAS.t42 VOUT.t7 GND.t62 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X112 VDD.t118 GND.t227 a_n11384_10929.t3 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.8853 ps=5.32 w=2.27 l=5.93
X113 VDD.t36 VDD.t34 VDD.t35 VDD.t28 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X114 VDD.t33 VDD.t31 VDD.t32 VDD.t28 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X115 GND.t130 GND.t128 VP.t1 GND.t129 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X116 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 GND.t61 GND.t60 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=4.06
X117 GND.t127 GND.t124 GND.t126 GND.t125 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X118 GND.t77 CS_BIAS.t6 CS_BIAS.t7 GND.t45 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X119 VDD.t30 VDD.t27 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X120 GND.t30 CS_BIAS.t4 CS_BIAS.t5 GND.t28 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X121 a_n11384_10929.t2 GND.t228 VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=5.93
X122 GND.t123 GND.t120 GND.t122 GND.t121 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X123 GND.t23 VP.t9 a_n7464_n776.t3 GND.t22 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=2.7963 ps=15.12 w=7.17 l=6.98
X124 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t7 GND.t6 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=4.06
X125 VDD.t26 VDD.t24 VDD.t25 VDD.t3 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X126 a_n4580_9541.t6 GND.t229 VDD.t114 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=5.93
X127 a_n7464_n776.t4 VP.t10 GND.t34 GND.t33 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X128 GND.t38 VN.t12 a_n7464_n776.t16 GND.t37 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X129 VDD.t23 VDD.t20 VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=5.93
X130 GND.t5 VP.t11 a_n7464_n776.t0 GND.t4 sky130_fd_pr__nfet_01v8 ad=2.7963 pd=15.12 as=1.18305 ps=7.5 w=7.17 l=6.98
X131 a_n7464_n776.t15 VN.t13 GND.t36 GND.t35 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X132 GND.t119 GND.t117 VP.t0 GND.t118 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X133 GND.t116 GND.t114 VN.t0 GND.t115 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X134 GND.t113 GND.t110 GND.t112 GND.t111 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X135 VOUT.t6 CS_BIAS.t43 GND.t51 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=2.37
X136 a_n11384_10929.t1 GND.t230 VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=5.93
X137 GND.t109 GND.t106 GND.t108 GND.t107 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=0 ps=0 w=4.14 l=4.06
X138 GND.t9 VP.t12 a_n7464_n776.t1 GND.t8 sky130_fd_pr__nfet_01v8 ad=2.7963 pd=15.12 as=1.18305 ps=7.5 w=7.17 l=6.98
X139 VDD.t19 VDD.t17 VDD.t18 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X140 VDD.t110 GND.t231 a_n4580_9541.t5 VDD.t109 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=5.93
X141 GND.t65 CS_BIAS.t44 VOUT.t5 GND.t64 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X142 VDD.t16 VDD.t14 VDD.t15 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X143 a_n4580_9541.t4 GND.t232 VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=5.93
X144 GND.t46 CS_BIAS.t45 VOUT.t4 GND.t45 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X145 VOUT.t3 CS_BIAS.t46 GND.t26 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X146 VOUT.t2 CS_BIAS.t47 GND.t203 GND.t14 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=2.37
X147 VDD.t13 VDD.t10 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0 ps=0 w=2.27 l=5.93
X148 VDD.t9 VDD.t6 VDD.t8 VDD.t7 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X149 CS_BIAS.t3 CS_BIAS.t2 GND.t205 GND.t14 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0.44715 ps=3.04 w=2.71 l=2.37
X150 GND.t105 GND.t102 GND.t104 GND.t103 sky130_fd_pr__nfet_01v8 ad=2.7963 pd=15.12 as=0 ps=0 w=7.17 l=6.98
X151 GND.t101 GND.t98 GND.t100 GND.t99 sky130_fd_pr__nfet_01v8 ad=1.0569 pd=6.2 as=0 ps=0 w=2.71 l=2.37
X152 VOUT.t46 a_n4580_9541.t0 sky130_fd_pr__cap_mim_m3_1 l=10.72 w=5.27
X153 a_n11384_10929.t0 GND.t233 VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=5.93
X154 a_11512_10929# a_11512_10929# a_11512_10929# VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=1.7706 ps=10.64 w=2.27 l=5.93
X155 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t209 GND.t208 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=4.06
X156 CS_BIAS.t1 CS_BIAS.t0 GND.t210 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X157 VOUT.t47 a_n4580_9541.t0 sky130_fd_pr__cap_mim_m3_1 l=10.72 w=5.27
X158 VOUT.t1 CS_BIAS.t48 GND.t50 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=1.0569 ps=6.2 w=2.71 l=2.37
X159 GND.t202 CS_BIAS.t49 VOUT.t0 GND.t64 sky130_fd_pr__nfet_01v8 ad=0.44715 pd=3.04 as=0.44715 ps=3.04 w=2.71 l=2.37
X160 VOUT.t33 GND.t234 VDD.t104 VDD.t98 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=1.5561 ps=8.76 w=3.99 l=3.26
X161 VOUT.t36 GND.t235 VDD.t103 VDD.t98 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=1.5561 ps=8.76 w=3.99 l=3.26
X162 a_n7464_n776.t2 VP.t13 GND.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=1.18305 pd=7.5 as=1.18305 ps=7.5 w=7.17 l=6.98
X163 a_n4580_9541.t9 GND.t92 GND.t93 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=5.93
X164 a_n4580_9541.t3 GND.t236 VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=5.93
X165 VOUT.t39 GND.t237 VDD.t99 VDD.t98 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=1.5561 ps=8.76 w=3.99 l=3.26
X166 VDD.t97 GND.t238 a_n4580_9541.t2 VDD.t96 sky130_fd_pr__pfet_01v8 ad=0.37455 pd=2.6 as=0.37455 ps=2.6 w=2.27 l=5.93
X167 VDD.t5 VDD.t2 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=1.5561 pd=8.76 as=0 ps=0 w=3.99 l=3.26
X168 a_n7464_n776.t6 DIFFPAIR_BIAS.t13 GND.t49 GND.t48 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=4.06
X169 a_n7464_n776.t5 DIFFPAIR_BIAS.t14 GND.t19 GND.t18 sky130_fd_pr__nfet_01v8 ad=1.6146 pd=9.06 as=1.6146 ps=9.06 w=4.14 l=4.06
X170 GND.t91 GND.t88 GND.t90 GND.t89 sky130_fd_pr__nfet_01v8 ad=2.7963 pd=15.12 as=0 ps=0 w=7.17 l=6.98
X171 a_n4580_9541.t1 GND.t239 VDD.t95 VDD.t94 sky130_fd_pr__pfet_01v8 ad=0.8853 pd=5.32 as=0.37455 ps=2.6 w=2.27 l=5.93
R0 GND.n8216 GND.n532 1529.15
R1 GND.n7375 GND.n1035 1031.54
R2 GND.n7221 GND.n1176 939.619
R3 GND.n382 GND.n242 763.976
R4 GND.n8447 GND.n251 763.976
R5 GND.n6450 GND.n6449 763.976
R6 GND.n6510 GND.n3070 763.976
R7 GND.n7043 GND.n1385 763.976
R8 GND.n7045 GND.n1379 763.976
R9 GND.n7115 GND.n7114 763.976
R10 GND.n7177 GND.n1246 763.976
R11 GND.n2829 GND.n2827 761.573
R12 GND.n6627 GND.n2903 761.573
R13 GND.n4319 GND.n2663 761.573
R14 GND.n6859 GND.n2665 761.573
R15 GND.n7374 GND.n1036 732.745
R16 GND.n8215 GND.n533 732.745
R17 GND.n8396 GND.n423 732.745
R18 GND.n7222 GND.n1177 732.745
R19 GND.n6271 GND.n247 718.33
R20 GND.n6294 GND.n252 718.33
R21 GND.n5820 GND.n3066 718.33
R22 GND.n6447 GND.n5822 718.33
R23 GND.n1935 GND.n1383 718.33
R24 GND.n6989 GND.n1381 718.33
R25 GND.n1291 GND.n1242 718.33
R26 GND.n7112 GND.n1293 718.33
R27 GND.n1935 GND.n1436 589.749
R28 GND.n6111 GND.n3066 588.893
R29 GND.n7370 GND.n1036 585
R30 GND.n1036 GND.n1035 585
R31 GND.n7369 GND.n7368 585
R32 GND.n7368 GND.n7367 585
R33 GND.n1039 GND.n1038 585
R34 GND.n7366 GND.n1039 585
R35 GND.n7364 GND.n7363 585
R36 GND.n7365 GND.n7364 585
R37 GND.n7362 GND.n1041 585
R38 GND.n1041 GND.n1040 585
R39 GND.n7361 GND.n7360 585
R40 GND.n7360 GND.n7359 585
R41 GND.n1047 GND.n1046 585
R42 GND.n7358 GND.n1047 585
R43 GND.n7356 GND.n7355 585
R44 GND.n7357 GND.n7356 585
R45 GND.n7354 GND.n1049 585
R46 GND.n1049 GND.n1048 585
R47 GND.n7353 GND.n7352 585
R48 GND.n7352 GND.n7351 585
R49 GND.n1055 GND.n1054 585
R50 GND.n7350 GND.n1055 585
R51 GND.n7348 GND.n7347 585
R52 GND.n7349 GND.n7348 585
R53 GND.n7346 GND.n1057 585
R54 GND.n1057 GND.n1056 585
R55 GND.n7345 GND.n7344 585
R56 GND.n7344 GND.n7343 585
R57 GND.n1063 GND.n1062 585
R58 GND.n7342 GND.n1063 585
R59 GND.n7340 GND.n7339 585
R60 GND.n7341 GND.n7340 585
R61 GND.n7338 GND.n1065 585
R62 GND.n1065 GND.n1064 585
R63 GND.n7337 GND.n7336 585
R64 GND.n7336 GND.n7335 585
R65 GND.n1071 GND.n1070 585
R66 GND.n7334 GND.n1071 585
R67 GND.n7332 GND.n7331 585
R68 GND.n7333 GND.n7332 585
R69 GND.n7330 GND.n1073 585
R70 GND.n1073 GND.n1072 585
R71 GND.n7329 GND.n7328 585
R72 GND.n7328 GND.n7327 585
R73 GND.n1079 GND.n1078 585
R74 GND.n7326 GND.n1079 585
R75 GND.n7324 GND.n7323 585
R76 GND.n7325 GND.n7324 585
R77 GND.n7322 GND.n1081 585
R78 GND.n1081 GND.n1080 585
R79 GND.n7321 GND.n7320 585
R80 GND.n7320 GND.n7319 585
R81 GND.n1087 GND.n1086 585
R82 GND.n7318 GND.n1087 585
R83 GND.n7316 GND.n7315 585
R84 GND.n7317 GND.n7316 585
R85 GND.n7314 GND.n1089 585
R86 GND.n1089 GND.n1088 585
R87 GND.n7313 GND.n7312 585
R88 GND.n7312 GND.n7311 585
R89 GND.n1095 GND.n1094 585
R90 GND.n7310 GND.n1095 585
R91 GND.n7308 GND.n7307 585
R92 GND.n7309 GND.n7308 585
R93 GND.n7306 GND.n1097 585
R94 GND.n1097 GND.n1096 585
R95 GND.n7305 GND.n7304 585
R96 GND.n7304 GND.n7303 585
R97 GND.n1103 GND.n1102 585
R98 GND.n7302 GND.n1103 585
R99 GND.n7300 GND.n7299 585
R100 GND.n7301 GND.n7300 585
R101 GND.n7298 GND.n1105 585
R102 GND.n1105 GND.n1104 585
R103 GND.n7297 GND.n7296 585
R104 GND.n7296 GND.n7295 585
R105 GND.n1111 GND.n1110 585
R106 GND.n7294 GND.n1111 585
R107 GND.n7292 GND.n7291 585
R108 GND.n7293 GND.n7292 585
R109 GND.n7290 GND.n1113 585
R110 GND.n1113 GND.n1112 585
R111 GND.n7289 GND.n7288 585
R112 GND.n7288 GND.n7287 585
R113 GND.n1119 GND.n1118 585
R114 GND.n7286 GND.n1119 585
R115 GND.n7284 GND.n7283 585
R116 GND.n7285 GND.n7284 585
R117 GND.n7282 GND.n1121 585
R118 GND.n1121 GND.n1120 585
R119 GND.n7281 GND.n7280 585
R120 GND.n7280 GND.n7279 585
R121 GND.n1127 GND.n1126 585
R122 GND.n7278 GND.n1127 585
R123 GND.n7276 GND.n7275 585
R124 GND.n7277 GND.n7276 585
R125 GND.n7274 GND.n1129 585
R126 GND.n1129 GND.n1128 585
R127 GND.n7273 GND.n7272 585
R128 GND.n7272 GND.n7271 585
R129 GND.n1135 GND.n1134 585
R130 GND.n7270 GND.n1135 585
R131 GND.n7268 GND.n7267 585
R132 GND.n7269 GND.n7268 585
R133 GND.n7266 GND.n1137 585
R134 GND.n1137 GND.n1136 585
R135 GND.n7265 GND.n7264 585
R136 GND.n7264 GND.n7263 585
R137 GND.n1143 GND.n1142 585
R138 GND.n7262 GND.n1143 585
R139 GND.n7260 GND.n7259 585
R140 GND.n7261 GND.n7260 585
R141 GND.n7258 GND.n1145 585
R142 GND.n1145 GND.n1144 585
R143 GND.n7257 GND.n7256 585
R144 GND.n7256 GND.n7255 585
R145 GND.n1151 GND.n1150 585
R146 GND.n7254 GND.n1151 585
R147 GND.n7252 GND.n7251 585
R148 GND.n7253 GND.n7252 585
R149 GND.n7250 GND.n1153 585
R150 GND.n1153 GND.n1152 585
R151 GND.n7249 GND.n7248 585
R152 GND.n7248 GND.n7247 585
R153 GND.n1159 GND.n1158 585
R154 GND.n7246 GND.n1159 585
R155 GND.n7244 GND.n7243 585
R156 GND.n7245 GND.n7244 585
R157 GND.n7242 GND.n1161 585
R158 GND.n1161 GND.n1160 585
R159 GND.n7241 GND.n7240 585
R160 GND.n7240 GND.n7239 585
R161 GND.n1167 GND.n1166 585
R162 GND.n7238 GND.n1167 585
R163 GND.n7236 GND.n7235 585
R164 GND.n7237 GND.n7236 585
R165 GND.n7234 GND.n1169 585
R166 GND.n1169 GND.n1168 585
R167 GND.n7233 GND.n7232 585
R168 GND.n7232 GND.n7231 585
R169 GND.n1175 GND.n1174 585
R170 GND.n7230 GND.n1175 585
R171 GND.n7228 GND.n7227 585
R172 GND.n7229 GND.n7228 585
R173 GND.n7226 GND.n1177 585
R174 GND.n1177 GND.n1176 585
R175 GND.n7374 GND.n7373 585
R176 GND.n7375 GND.n7374 585
R177 GND.n1034 GND.n1033 585
R178 GND.n7376 GND.n1034 585
R179 GND.n7379 GND.n7378 585
R180 GND.n7378 GND.n7377 585
R181 GND.n1031 GND.n1030 585
R182 GND.n1030 GND.n1029 585
R183 GND.n7384 GND.n7383 585
R184 GND.n7385 GND.n7384 585
R185 GND.n1028 GND.n1027 585
R186 GND.n7386 GND.n1028 585
R187 GND.n7389 GND.n7388 585
R188 GND.n7388 GND.n7387 585
R189 GND.n1025 GND.n1024 585
R190 GND.n1024 GND.n1023 585
R191 GND.n7394 GND.n7393 585
R192 GND.n7395 GND.n7394 585
R193 GND.n1022 GND.n1021 585
R194 GND.n7396 GND.n1022 585
R195 GND.n7399 GND.n7398 585
R196 GND.n7398 GND.n7397 585
R197 GND.n1019 GND.n1018 585
R198 GND.n1018 GND.n1017 585
R199 GND.n7404 GND.n7403 585
R200 GND.n7405 GND.n7404 585
R201 GND.n1016 GND.n1015 585
R202 GND.n7406 GND.n1016 585
R203 GND.n7409 GND.n7408 585
R204 GND.n7408 GND.n7407 585
R205 GND.n1013 GND.n1012 585
R206 GND.n1012 GND.n1011 585
R207 GND.n7414 GND.n7413 585
R208 GND.n7415 GND.n7414 585
R209 GND.n1010 GND.n1009 585
R210 GND.n7416 GND.n1010 585
R211 GND.n7419 GND.n7418 585
R212 GND.n7418 GND.n7417 585
R213 GND.n1007 GND.n1006 585
R214 GND.n1006 GND.n1005 585
R215 GND.n7424 GND.n7423 585
R216 GND.n7425 GND.n7424 585
R217 GND.n1004 GND.n1003 585
R218 GND.n7426 GND.n1004 585
R219 GND.n7429 GND.n7428 585
R220 GND.n7428 GND.n7427 585
R221 GND.n1001 GND.n1000 585
R222 GND.n1000 GND.n999 585
R223 GND.n7434 GND.n7433 585
R224 GND.n7435 GND.n7434 585
R225 GND.n998 GND.n997 585
R226 GND.n7436 GND.n998 585
R227 GND.n7439 GND.n7438 585
R228 GND.n7438 GND.n7437 585
R229 GND.n995 GND.n994 585
R230 GND.n994 GND.n993 585
R231 GND.n7444 GND.n7443 585
R232 GND.n7445 GND.n7444 585
R233 GND.n992 GND.n991 585
R234 GND.n7446 GND.n992 585
R235 GND.n7449 GND.n7448 585
R236 GND.n7448 GND.n7447 585
R237 GND.n989 GND.n988 585
R238 GND.n988 GND.n987 585
R239 GND.n7454 GND.n7453 585
R240 GND.n7455 GND.n7454 585
R241 GND.n986 GND.n985 585
R242 GND.n7456 GND.n986 585
R243 GND.n7459 GND.n7458 585
R244 GND.n7458 GND.n7457 585
R245 GND.n983 GND.n982 585
R246 GND.n982 GND.n981 585
R247 GND.n7464 GND.n7463 585
R248 GND.n7465 GND.n7464 585
R249 GND.n980 GND.n979 585
R250 GND.n7466 GND.n980 585
R251 GND.n7469 GND.n7468 585
R252 GND.n7468 GND.n7467 585
R253 GND.n977 GND.n976 585
R254 GND.n976 GND.n975 585
R255 GND.n7474 GND.n7473 585
R256 GND.n7475 GND.n7474 585
R257 GND.n974 GND.n973 585
R258 GND.n7476 GND.n974 585
R259 GND.n7479 GND.n7478 585
R260 GND.n7478 GND.n7477 585
R261 GND.n971 GND.n970 585
R262 GND.n970 GND.n969 585
R263 GND.n7484 GND.n7483 585
R264 GND.n7485 GND.n7484 585
R265 GND.n968 GND.n967 585
R266 GND.n7486 GND.n968 585
R267 GND.n7489 GND.n7488 585
R268 GND.n7488 GND.n7487 585
R269 GND.n965 GND.n964 585
R270 GND.n964 GND.n963 585
R271 GND.n7494 GND.n7493 585
R272 GND.n7495 GND.n7494 585
R273 GND.n962 GND.n961 585
R274 GND.n7496 GND.n962 585
R275 GND.n7499 GND.n7498 585
R276 GND.n7498 GND.n7497 585
R277 GND.n959 GND.n958 585
R278 GND.n958 GND.n957 585
R279 GND.n7504 GND.n7503 585
R280 GND.n7505 GND.n7504 585
R281 GND.n956 GND.n955 585
R282 GND.n7506 GND.n956 585
R283 GND.n7509 GND.n7508 585
R284 GND.n7508 GND.n7507 585
R285 GND.n953 GND.n952 585
R286 GND.n952 GND.n951 585
R287 GND.n7514 GND.n7513 585
R288 GND.n7515 GND.n7514 585
R289 GND.n950 GND.n949 585
R290 GND.n7516 GND.n950 585
R291 GND.n7519 GND.n7518 585
R292 GND.n7518 GND.n7517 585
R293 GND.n947 GND.n946 585
R294 GND.n946 GND.n945 585
R295 GND.n7524 GND.n7523 585
R296 GND.n7525 GND.n7524 585
R297 GND.n944 GND.n943 585
R298 GND.n7526 GND.n944 585
R299 GND.n7529 GND.n7528 585
R300 GND.n7528 GND.n7527 585
R301 GND.n941 GND.n940 585
R302 GND.n940 GND.n939 585
R303 GND.n7534 GND.n7533 585
R304 GND.n7535 GND.n7534 585
R305 GND.n938 GND.n937 585
R306 GND.n7536 GND.n938 585
R307 GND.n7539 GND.n7538 585
R308 GND.n7538 GND.n7537 585
R309 GND.n935 GND.n934 585
R310 GND.n934 GND.n933 585
R311 GND.n7544 GND.n7543 585
R312 GND.n7545 GND.n7544 585
R313 GND.n932 GND.n931 585
R314 GND.n7546 GND.n932 585
R315 GND.n7549 GND.n7548 585
R316 GND.n7548 GND.n7547 585
R317 GND.n929 GND.n928 585
R318 GND.n928 GND.n927 585
R319 GND.n7554 GND.n7553 585
R320 GND.n7555 GND.n7554 585
R321 GND.n926 GND.n925 585
R322 GND.n7556 GND.n926 585
R323 GND.n7559 GND.n7558 585
R324 GND.n7558 GND.n7557 585
R325 GND.n923 GND.n922 585
R326 GND.n922 GND.n921 585
R327 GND.n7564 GND.n7563 585
R328 GND.n7565 GND.n7564 585
R329 GND.n920 GND.n919 585
R330 GND.n7566 GND.n920 585
R331 GND.n7569 GND.n7568 585
R332 GND.n7568 GND.n7567 585
R333 GND.n917 GND.n916 585
R334 GND.n916 GND.n915 585
R335 GND.n7574 GND.n7573 585
R336 GND.n7575 GND.n7574 585
R337 GND.n914 GND.n913 585
R338 GND.n7576 GND.n914 585
R339 GND.n7579 GND.n7578 585
R340 GND.n7578 GND.n7577 585
R341 GND.n911 GND.n910 585
R342 GND.n910 GND.n909 585
R343 GND.n7584 GND.n7583 585
R344 GND.n7585 GND.n7584 585
R345 GND.n908 GND.n907 585
R346 GND.n7586 GND.n908 585
R347 GND.n7589 GND.n7588 585
R348 GND.n7588 GND.n7587 585
R349 GND.n905 GND.n904 585
R350 GND.n904 GND.n903 585
R351 GND.n7594 GND.n7593 585
R352 GND.n7595 GND.n7594 585
R353 GND.n902 GND.n901 585
R354 GND.n7596 GND.n902 585
R355 GND.n7599 GND.n7598 585
R356 GND.n7598 GND.n7597 585
R357 GND.n899 GND.n898 585
R358 GND.n898 GND.n897 585
R359 GND.n7604 GND.n7603 585
R360 GND.n7605 GND.n7604 585
R361 GND.n896 GND.n895 585
R362 GND.n7606 GND.n896 585
R363 GND.n7609 GND.n7608 585
R364 GND.n7608 GND.n7607 585
R365 GND.n893 GND.n892 585
R366 GND.n892 GND.n891 585
R367 GND.n7614 GND.n7613 585
R368 GND.n7615 GND.n7614 585
R369 GND.n890 GND.n889 585
R370 GND.n7616 GND.n890 585
R371 GND.n7619 GND.n7618 585
R372 GND.n7618 GND.n7617 585
R373 GND.n887 GND.n886 585
R374 GND.n886 GND.n885 585
R375 GND.n7624 GND.n7623 585
R376 GND.n7625 GND.n7624 585
R377 GND.n884 GND.n883 585
R378 GND.n7626 GND.n884 585
R379 GND.n7629 GND.n7628 585
R380 GND.n7628 GND.n7627 585
R381 GND.n881 GND.n880 585
R382 GND.n880 GND.n879 585
R383 GND.n7634 GND.n7633 585
R384 GND.n7635 GND.n7634 585
R385 GND.n878 GND.n877 585
R386 GND.n7636 GND.n878 585
R387 GND.n7639 GND.n7638 585
R388 GND.n7638 GND.n7637 585
R389 GND.n875 GND.n874 585
R390 GND.n874 GND.n873 585
R391 GND.n7644 GND.n7643 585
R392 GND.n7645 GND.n7644 585
R393 GND.n872 GND.n871 585
R394 GND.n7646 GND.n872 585
R395 GND.n7649 GND.n7648 585
R396 GND.n7648 GND.n7647 585
R397 GND.n869 GND.n868 585
R398 GND.n868 GND.n867 585
R399 GND.n7654 GND.n7653 585
R400 GND.n7655 GND.n7654 585
R401 GND.n866 GND.n865 585
R402 GND.n7656 GND.n866 585
R403 GND.n7659 GND.n7658 585
R404 GND.n7658 GND.n7657 585
R405 GND.n863 GND.n862 585
R406 GND.n862 GND.n861 585
R407 GND.n7664 GND.n7663 585
R408 GND.n7665 GND.n7664 585
R409 GND.n860 GND.n859 585
R410 GND.n7666 GND.n860 585
R411 GND.n7669 GND.n7668 585
R412 GND.n7668 GND.n7667 585
R413 GND.n857 GND.n856 585
R414 GND.n856 GND.n855 585
R415 GND.n7674 GND.n7673 585
R416 GND.n7675 GND.n7674 585
R417 GND.n854 GND.n853 585
R418 GND.n7676 GND.n854 585
R419 GND.n7679 GND.n7678 585
R420 GND.n7678 GND.n7677 585
R421 GND.n851 GND.n850 585
R422 GND.n850 GND.n849 585
R423 GND.n7684 GND.n7683 585
R424 GND.n7685 GND.n7684 585
R425 GND.n848 GND.n847 585
R426 GND.n7686 GND.n848 585
R427 GND.n7689 GND.n7688 585
R428 GND.n7688 GND.n7687 585
R429 GND.n845 GND.n844 585
R430 GND.n844 GND.n843 585
R431 GND.n7694 GND.n7693 585
R432 GND.n7695 GND.n7694 585
R433 GND.n842 GND.n841 585
R434 GND.n7696 GND.n842 585
R435 GND.n7699 GND.n7698 585
R436 GND.n7698 GND.n7697 585
R437 GND.n839 GND.n838 585
R438 GND.n838 GND.n837 585
R439 GND.n7704 GND.n7703 585
R440 GND.n7705 GND.n7704 585
R441 GND.n836 GND.n835 585
R442 GND.n7706 GND.n836 585
R443 GND.n7709 GND.n7708 585
R444 GND.n7708 GND.n7707 585
R445 GND.n833 GND.n832 585
R446 GND.n832 GND.n831 585
R447 GND.n7714 GND.n7713 585
R448 GND.n7715 GND.n7714 585
R449 GND.n830 GND.n829 585
R450 GND.n7716 GND.n830 585
R451 GND.n7719 GND.n7718 585
R452 GND.n7718 GND.n7717 585
R453 GND.n827 GND.n826 585
R454 GND.n826 GND.n825 585
R455 GND.n7724 GND.n7723 585
R456 GND.n7725 GND.n7724 585
R457 GND.n824 GND.n823 585
R458 GND.n7726 GND.n824 585
R459 GND.n7729 GND.n7728 585
R460 GND.n7728 GND.n7727 585
R461 GND.n821 GND.n820 585
R462 GND.n820 GND.n819 585
R463 GND.n7734 GND.n7733 585
R464 GND.n7735 GND.n7734 585
R465 GND.n818 GND.n817 585
R466 GND.n7736 GND.n818 585
R467 GND.n7739 GND.n7738 585
R468 GND.n7738 GND.n7737 585
R469 GND.n815 GND.n814 585
R470 GND.n814 GND.n813 585
R471 GND.n7744 GND.n7743 585
R472 GND.n7745 GND.n7744 585
R473 GND.n812 GND.n811 585
R474 GND.n7746 GND.n812 585
R475 GND.n7749 GND.n7748 585
R476 GND.n7748 GND.n7747 585
R477 GND.n809 GND.n808 585
R478 GND.n808 GND.n807 585
R479 GND.n7754 GND.n7753 585
R480 GND.n7755 GND.n7754 585
R481 GND.n806 GND.n805 585
R482 GND.n7756 GND.n806 585
R483 GND.n7759 GND.n7758 585
R484 GND.n7758 GND.n7757 585
R485 GND.n803 GND.n802 585
R486 GND.n802 GND.n801 585
R487 GND.n7764 GND.n7763 585
R488 GND.n7765 GND.n7764 585
R489 GND.n800 GND.n799 585
R490 GND.n7766 GND.n800 585
R491 GND.n7769 GND.n7768 585
R492 GND.n7768 GND.n7767 585
R493 GND.n797 GND.n796 585
R494 GND.n796 GND.n795 585
R495 GND.n7774 GND.n7773 585
R496 GND.n7775 GND.n7774 585
R497 GND.n794 GND.n793 585
R498 GND.n7776 GND.n794 585
R499 GND.n7779 GND.n7778 585
R500 GND.n7778 GND.n7777 585
R501 GND.n791 GND.n790 585
R502 GND.n790 GND.n789 585
R503 GND.n7784 GND.n7783 585
R504 GND.n7785 GND.n7784 585
R505 GND.n788 GND.n787 585
R506 GND.n7786 GND.n788 585
R507 GND.n7789 GND.n7788 585
R508 GND.n7788 GND.n7787 585
R509 GND.n785 GND.n784 585
R510 GND.n784 GND.n783 585
R511 GND.n7794 GND.n7793 585
R512 GND.n7795 GND.n7794 585
R513 GND.n782 GND.n781 585
R514 GND.n7796 GND.n782 585
R515 GND.n7799 GND.n7798 585
R516 GND.n7798 GND.n7797 585
R517 GND.n779 GND.n778 585
R518 GND.n778 GND.n777 585
R519 GND.n7804 GND.n7803 585
R520 GND.n7805 GND.n7804 585
R521 GND.n776 GND.n775 585
R522 GND.n7806 GND.n776 585
R523 GND.n7809 GND.n7808 585
R524 GND.n7808 GND.n7807 585
R525 GND.n773 GND.n772 585
R526 GND.n772 GND.n771 585
R527 GND.n7814 GND.n7813 585
R528 GND.n7815 GND.n7814 585
R529 GND.n770 GND.n769 585
R530 GND.n7816 GND.n770 585
R531 GND.n7819 GND.n7818 585
R532 GND.n7818 GND.n7817 585
R533 GND.n767 GND.n766 585
R534 GND.n766 GND.n765 585
R535 GND.n7824 GND.n7823 585
R536 GND.n7825 GND.n7824 585
R537 GND.n764 GND.n763 585
R538 GND.n7826 GND.n764 585
R539 GND.n7829 GND.n7828 585
R540 GND.n7828 GND.n7827 585
R541 GND.n761 GND.n760 585
R542 GND.n760 GND.n759 585
R543 GND.n7834 GND.n7833 585
R544 GND.n7835 GND.n7834 585
R545 GND.n758 GND.n757 585
R546 GND.n7836 GND.n758 585
R547 GND.n7839 GND.n7838 585
R548 GND.n7838 GND.n7837 585
R549 GND.n755 GND.n754 585
R550 GND.n754 GND.n753 585
R551 GND.n7844 GND.n7843 585
R552 GND.n7845 GND.n7844 585
R553 GND.n752 GND.n751 585
R554 GND.n7846 GND.n752 585
R555 GND.n7849 GND.n7848 585
R556 GND.n7848 GND.n7847 585
R557 GND.n749 GND.n748 585
R558 GND.n748 GND.n747 585
R559 GND.n7854 GND.n7853 585
R560 GND.n7855 GND.n7854 585
R561 GND.n746 GND.n745 585
R562 GND.n7856 GND.n746 585
R563 GND.n7859 GND.n7858 585
R564 GND.n7858 GND.n7857 585
R565 GND.n743 GND.n742 585
R566 GND.n742 GND.n741 585
R567 GND.n7864 GND.n7863 585
R568 GND.n7865 GND.n7864 585
R569 GND.n740 GND.n739 585
R570 GND.n7866 GND.n740 585
R571 GND.n7869 GND.n7868 585
R572 GND.n7868 GND.n7867 585
R573 GND.n737 GND.n736 585
R574 GND.n736 GND.n735 585
R575 GND.n7874 GND.n7873 585
R576 GND.n7875 GND.n7874 585
R577 GND.n734 GND.n733 585
R578 GND.n7876 GND.n734 585
R579 GND.n7879 GND.n7878 585
R580 GND.n7878 GND.n7877 585
R581 GND.n731 GND.n730 585
R582 GND.n730 GND.n729 585
R583 GND.n7884 GND.n7883 585
R584 GND.n7885 GND.n7884 585
R585 GND.n728 GND.n727 585
R586 GND.n7886 GND.n728 585
R587 GND.n7889 GND.n7888 585
R588 GND.n7888 GND.n7887 585
R589 GND.n725 GND.n724 585
R590 GND.n724 GND.n723 585
R591 GND.n7894 GND.n7893 585
R592 GND.n7895 GND.n7894 585
R593 GND.n722 GND.n721 585
R594 GND.n7896 GND.n722 585
R595 GND.n7899 GND.n7898 585
R596 GND.n7898 GND.n7897 585
R597 GND.n719 GND.n718 585
R598 GND.n718 GND.n717 585
R599 GND.n7904 GND.n7903 585
R600 GND.n7905 GND.n7904 585
R601 GND.n716 GND.n715 585
R602 GND.n7906 GND.n716 585
R603 GND.n7909 GND.n7908 585
R604 GND.n7908 GND.n7907 585
R605 GND.n713 GND.n712 585
R606 GND.n712 GND.n711 585
R607 GND.n7914 GND.n7913 585
R608 GND.n7915 GND.n7914 585
R609 GND.n710 GND.n709 585
R610 GND.n7916 GND.n710 585
R611 GND.n7919 GND.n7918 585
R612 GND.n7918 GND.n7917 585
R613 GND.n707 GND.n706 585
R614 GND.n706 GND.n705 585
R615 GND.n7924 GND.n7923 585
R616 GND.n7925 GND.n7924 585
R617 GND.n704 GND.n703 585
R618 GND.n7926 GND.n704 585
R619 GND.n7929 GND.n7928 585
R620 GND.n7928 GND.n7927 585
R621 GND.n701 GND.n700 585
R622 GND.n700 GND.n699 585
R623 GND.n7934 GND.n7933 585
R624 GND.n7935 GND.n7934 585
R625 GND.n698 GND.n697 585
R626 GND.n7936 GND.n698 585
R627 GND.n7939 GND.n7938 585
R628 GND.n7938 GND.n7937 585
R629 GND.n695 GND.n694 585
R630 GND.n694 GND.n693 585
R631 GND.n7944 GND.n7943 585
R632 GND.n7945 GND.n7944 585
R633 GND.n692 GND.n691 585
R634 GND.n7946 GND.n692 585
R635 GND.n7949 GND.n7948 585
R636 GND.n7948 GND.n7947 585
R637 GND.n689 GND.n688 585
R638 GND.n688 GND.n687 585
R639 GND.n7954 GND.n7953 585
R640 GND.n7955 GND.n7954 585
R641 GND.n686 GND.n685 585
R642 GND.n7956 GND.n686 585
R643 GND.n7959 GND.n7958 585
R644 GND.n7958 GND.n7957 585
R645 GND.n683 GND.n682 585
R646 GND.n682 GND.n681 585
R647 GND.n7964 GND.n7963 585
R648 GND.n7965 GND.n7964 585
R649 GND.n680 GND.n679 585
R650 GND.n7966 GND.n680 585
R651 GND.n7969 GND.n7968 585
R652 GND.n7968 GND.n7967 585
R653 GND.n677 GND.n676 585
R654 GND.n676 GND.n675 585
R655 GND.n7974 GND.n7973 585
R656 GND.n7975 GND.n7974 585
R657 GND.n674 GND.n673 585
R658 GND.n7976 GND.n674 585
R659 GND.n7979 GND.n7978 585
R660 GND.n7978 GND.n7977 585
R661 GND.n671 GND.n670 585
R662 GND.n670 GND.n669 585
R663 GND.n7984 GND.n7983 585
R664 GND.n7985 GND.n7984 585
R665 GND.n668 GND.n667 585
R666 GND.n7986 GND.n668 585
R667 GND.n7989 GND.n7988 585
R668 GND.n7988 GND.n7987 585
R669 GND.n665 GND.n664 585
R670 GND.n664 GND.n663 585
R671 GND.n7994 GND.n7993 585
R672 GND.n7995 GND.n7994 585
R673 GND.n662 GND.n661 585
R674 GND.n7996 GND.n662 585
R675 GND.n7999 GND.n7998 585
R676 GND.n7998 GND.n7997 585
R677 GND.n659 GND.n658 585
R678 GND.n658 GND.n657 585
R679 GND.n8004 GND.n8003 585
R680 GND.n8005 GND.n8004 585
R681 GND.n656 GND.n655 585
R682 GND.n8006 GND.n656 585
R683 GND.n8009 GND.n8008 585
R684 GND.n8008 GND.n8007 585
R685 GND.n653 GND.n652 585
R686 GND.n652 GND.n651 585
R687 GND.n8014 GND.n8013 585
R688 GND.n8015 GND.n8014 585
R689 GND.n650 GND.n649 585
R690 GND.n8016 GND.n650 585
R691 GND.n8019 GND.n8018 585
R692 GND.n8018 GND.n8017 585
R693 GND.n647 GND.n646 585
R694 GND.n646 GND.n645 585
R695 GND.n8024 GND.n8023 585
R696 GND.n8025 GND.n8024 585
R697 GND.n644 GND.n643 585
R698 GND.n8026 GND.n644 585
R699 GND.n8029 GND.n8028 585
R700 GND.n8028 GND.n8027 585
R701 GND.n641 GND.n640 585
R702 GND.n640 GND.n639 585
R703 GND.n8034 GND.n8033 585
R704 GND.n8035 GND.n8034 585
R705 GND.n638 GND.n637 585
R706 GND.n8036 GND.n638 585
R707 GND.n8039 GND.n8038 585
R708 GND.n8038 GND.n8037 585
R709 GND.n635 GND.n634 585
R710 GND.n634 GND.n633 585
R711 GND.n8044 GND.n8043 585
R712 GND.n8045 GND.n8044 585
R713 GND.n632 GND.n631 585
R714 GND.n8046 GND.n632 585
R715 GND.n8049 GND.n8048 585
R716 GND.n8048 GND.n8047 585
R717 GND.n629 GND.n628 585
R718 GND.n628 GND.n627 585
R719 GND.n8054 GND.n8053 585
R720 GND.n8055 GND.n8054 585
R721 GND.n626 GND.n625 585
R722 GND.n8056 GND.n626 585
R723 GND.n8059 GND.n8058 585
R724 GND.n8058 GND.n8057 585
R725 GND.n623 GND.n622 585
R726 GND.n622 GND.n621 585
R727 GND.n8064 GND.n8063 585
R728 GND.n8065 GND.n8064 585
R729 GND.n620 GND.n619 585
R730 GND.n8066 GND.n620 585
R731 GND.n8069 GND.n8068 585
R732 GND.n8068 GND.n8067 585
R733 GND.n617 GND.n616 585
R734 GND.n616 GND.n615 585
R735 GND.n8074 GND.n8073 585
R736 GND.n8075 GND.n8074 585
R737 GND.n614 GND.n613 585
R738 GND.n8076 GND.n614 585
R739 GND.n8079 GND.n8078 585
R740 GND.n8078 GND.n8077 585
R741 GND.n611 GND.n610 585
R742 GND.n610 GND.n609 585
R743 GND.n8084 GND.n8083 585
R744 GND.n8085 GND.n8084 585
R745 GND.n608 GND.n607 585
R746 GND.n8086 GND.n608 585
R747 GND.n8089 GND.n8088 585
R748 GND.n8088 GND.n8087 585
R749 GND.n605 GND.n604 585
R750 GND.n604 GND.n603 585
R751 GND.n8094 GND.n8093 585
R752 GND.n8095 GND.n8094 585
R753 GND.n602 GND.n601 585
R754 GND.n8096 GND.n602 585
R755 GND.n8099 GND.n8098 585
R756 GND.n8098 GND.n8097 585
R757 GND.n599 GND.n598 585
R758 GND.n598 GND.n597 585
R759 GND.n8104 GND.n8103 585
R760 GND.n8105 GND.n8104 585
R761 GND.n596 GND.n595 585
R762 GND.n8106 GND.n596 585
R763 GND.n8109 GND.n8108 585
R764 GND.n8108 GND.n8107 585
R765 GND.n593 GND.n592 585
R766 GND.n592 GND.n591 585
R767 GND.n8114 GND.n8113 585
R768 GND.n8115 GND.n8114 585
R769 GND.n590 GND.n589 585
R770 GND.n8116 GND.n590 585
R771 GND.n8119 GND.n8118 585
R772 GND.n8118 GND.n8117 585
R773 GND.n587 GND.n586 585
R774 GND.n586 GND.n585 585
R775 GND.n8124 GND.n8123 585
R776 GND.n8125 GND.n8124 585
R777 GND.n584 GND.n583 585
R778 GND.n8126 GND.n584 585
R779 GND.n8129 GND.n8128 585
R780 GND.n8128 GND.n8127 585
R781 GND.n581 GND.n580 585
R782 GND.n580 GND.n579 585
R783 GND.n8134 GND.n8133 585
R784 GND.n8135 GND.n8134 585
R785 GND.n578 GND.n577 585
R786 GND.n8136 GND.n578 585
R787 GND.n8139 GND.n8138 585
R788 GND.n8138 GND.n8137 585
R789 GND.n575 GND.n574 585
R790 GND.n574 GND.n573 585
R791 GND.n8144 GND.n8143 585
R792 GND.n8145 GND.n8144 585
R793 GND.n572 GND.n571 585
R794 GND.n8146 GND.n572 585
R795 GND.n8149 GND.n8148 585
R796 GND.n8148 GND.n8147 585
R797 GND.n569 GND.n568 585
R798 GND.n568 GND.n567 585
R799 GND.n8154 GND.n8153 585
R800 GND.n8155 GND.n8154 585
R801 GND.n566 GND.n565 585
R802 GND.n8156 GND.n566 585
R803 GND.n8159 GND.n8158 585
R804 GND.n8158 GND.n8157 585
R805 GND.n563 GND.n562 585
R806 GND.n562 GND.n561 585
R807 GND.n8164 GND.n8163 585
R808 GND.n8165 GND.n8164 585
R809 GND.n560 GND.n559 585
R810 GND.n8166 GND.n560 585
R811 GND.n8169 GND.n8168 585
R812 GND.n8168 GND.n8167 585
R813 GND.n557 GND.n556 585
R814 GND.n556 GND.n555 585
R815 GND.n8174 GND.n8173 585
R816 GND.n8175 GND.n8174 585
R817 GND.n554 GND.n553 585
R818 GND.n8176 GND.n554 585
R819 GND.n8179 GND.n8178 585
R820 GND.n8178 GND.n8177 585
R821 GND.n551 GND.n550 585
R822 GND.n550 GND.n549 585
R823 GND.n8184 GND.n8183 585
R824 GND.n8185 GND.n8184 585
R825 GND.n548 GND.n547 585
R826 GND.n8186 GND.n548 585
R827 GND.n8189 GND.n8188 585
R828 GND.n8188 GND.n8187 585
R829 GND.n545 GND.n544 585
R830 GND.n544 GND.n543 585
R831 GND.n8194 GND.n8193 585
R832 GND.n8195 GND.n8194 585
R833 GND.n542 GND.n541 585
R834 GND.n8196 GND.n542 585
R835 GND.n8199 GND.n8198 585
R836 GND.n8198 GND.n8197 585
R837 GND.n539 GND.n538 585
R838 GND.n538 GND.n537 585
R839 GND.n8205 GND.n8204 585
R840 GND.n8206 GND.n8205 585
R841 GND.n536 GND.n535 585
R842 GND.n8207 GND.n536 585
R843 GND.n8210 GND.n8209 585
R844 GND.n8209 GND.n8208 585
R845 GND.n8211 GND.n533 585
R846 GND.n533 GND.n532 585
R847 GND.n8396 GND.n8395 585
R848 GND.n8397 GND.n8396 585
R849 GND.n426 GND.n425 585
R850 GND.n425 GND.n424 585
R851 GND.n8390 GND.n8389 585
R852 GND.n8389 GND.n8388 585
R853 GND.n429 GND.n428 585
R854 GND.n8387 GND.n429 585
R855 GND.n8385 GND.n8384 585
R856 GND.n8386 GND.n8385 585
R857 GND.n432 GND.n431 585
R858 GND.n431 GND.n430 585
R859 GND.n8380 GND.n8379 585
R860 GND.n8379 GND.n8378 585
R861 GND.n435 GND.n434 585
R862 GND.n8377 GND.n435 585
R863 GND.n8375 GND.n8374 585
R864 GND.n8376 GND.n8375 585
R865 GND.n438 GND.n437 585
R866 GND.n437 GND.n436 585
R867 GND.n8370 GND.n8369 585
R868 GND.n8369 GND.n8368 585
R869 GND.n441 GND.n440 585
R870 GND.n8367 GND.n441 585
R871 GND.n8365 GND.n8364 585
R872 GND.n8366 GND.n8365 585
R873 GND.n444 GND.n443 585
R874 GND.n443 GND.n442 585
R875 GND.n8360 GND.n8359 585
R876 GND.n8359 GND.n8358 585
R877 GND.n447 GND.n446 585
R878 GND.n8357 GND.n447 585
R879 GND.n8355 GND.n8354 585
R880 GND.n8356 GND.n8355 585
R881 GND.n450 GND.n449 585
R882 GND.n449 GND.n448 585
R883 GND.n8350 GND.n8349 585
R884 GND.n8349 GND.n8348 585
R885 GND.n453 GND.n452 585
R886 GND.n8347 GND.n453 585
R887 GND.n8345 GND.n8344 585
R888 GND.n8346 GND.n8345 585
R889 GND.n456 GND.n455 585
R890 GND.n455 GND.n454 585
R891 GND.n8340 GND.n8339 585
R892 GND.n8339 GND.n8338 585
R893 GND.n459 GND.n458 585
R894 GND.n8337 GND.n459 585
R895 GND.n8335 GND.n8334 585
R896 GND.n8336 GND.n8335 585
R897 GND.n462 GND.n461 585
R898 GND.n461 GND.n460 585
R899 GND.n8330 GND.n8329 585
R900 GND.n8329 GND.n8328 585
R901 GND.n465 GND.n464 585
R902 GND.n8327 GND.n465 585
R903 GND.n8325 GND.n8324 585
R904 GND.n8326 GND.n8325 585
R905 GND.n468 GND.n467 585
R906 GND.n467 GND.n466 585
R907 GND.n8320 GND.n8319 585
R908 GND.n8319 GND.n8318 585
R909 GND.n471 GND.n470 585
R910 GND.n8317 GND.n471 585
R911 GND.n8315 GND.n8314 585
R912 GND.n8316 GND.n8315 585
R913 GND.n474 GND.n473 585
R914 GND.n473 GND.n472 585
R915 GND.n8310 GND.n8309 585
R916 GND.n8309 GND.n8308 585
R917 GND.n477 GND.n476 585
R918 GND.n8307 GND.n477 585
R919 GND.n8305 GND.n8304 585
R920 GND.n8306 GND.n8305 585
R921 GND.n480 GND.n479 585
R922 GND.n479 GND.n478 585
R923 GND.n8300 GND.n8299 585
R924 GND.n8299 GND.n8298 585
R925 GND.n483 GND.n482 585
R926 GND.n8297 GND.n483 585
R927 GND.n8295 GND.n8294 585
R928 GND.n8296 GND.n8295 585
R929 GND.n486 GND.n485 585
R930 GND.n485 GND.n484 585
R931 GND.n8290 GND.n8289 585
R932 GND.n8289 GND.n8288 585
R933 GND.n489 GND.n488 585
R934 GND.n8287 GND.n489 585
R935 GND.n8285 GND.n8284 585
R936 GND.n8286 GND.n8285 585
R937 GND.n492 GND.n491 585
R938 GND.n491 GND.n490 585
R939 GND.n8280 GND.n8279 585
R940 GND.n8279 GND.n8278 585
R941 GND.n495 GND.n494 585
R942 GND.n8277 GND.n495 585
R943 GND.n8275 GND.n8274 585
R944 GND.n8276 GND.n8275 585
R945 GND.n498 GND.n497 585
R946 GND.n497 GND.n496 585
R947 GND.n8270 GND.n8269 585
R948 GND.n8269 GND.n8268 585
R949 GND.n501 GND.n500 585
R950 GND.n8267 GND.n501 585
R951 GND.n8265 GND.n8264 585
R952 GND.n8266 GND.n8265 585
R953 GND.n504 GND.n503 585
R954 GND.n503 GND.n502 585
R955 GND.n8260 GND.n8259 585
R956 GND.n8259 GND.n8258 585
R957 GND.n507 GND.n506 585
R958 GND.n8257 GND.n507 585
R959 GND.n8255 GND.n8254 585
R960 GND.n8256 GND.n8255 585
R961 GND.n510 GND.n509 585
R962 GND.n509 GND.n508 585
R963 GND.n8250 GND.n8249 585
R964 GND.n8249 GND.n8248 585
R965 GND.n513 GND.n512 585
R966 GND.n8247 GND.n513 585
R967 GND.n8245 GND.n8244 585
R968 GND.n8246 GND.n8245 585
R969 GND.n516 GND.n515 585
R970 GND.n515 GND.n514 585
R971 GND.n8240 GND.n8239 585
R972 GND.n8239 GND.n8238 585
R973 GND.n519 GND.n518 585
R974 GND.n8237 GND.n519 585
R975 GND.n8235 GND.n8234 585
R976 GND.n8236 GND.n8235 585
R977 GND.n522 GND.n521 585
R978 GND.n521 GND.n520 585
R979 GND.n8230 GND.n8229 585
R980 GND.n8229 GND.n8228 585
R981 GND.n525 GND.n524 585
R982 GND.n8227 GND.n525 585
R983 GND.n8225 GND.n8224 585
R984 GND.n8226 GND.n8225 585
R985 GND.n528 GND.n527 585
R986 GND.n527 GND.n526 585
R987 GND.n8220 GND.n8219 585
R988 GND.n8219 GND.n8218 585
R989 GND.n531 GND.n530 585
R990 GND.n8217 GND.n531 585
R991 GND.n8215 GND.n8214 585
R992 GND.n8216 GND.n8215 585
R993 GND.n2514 GND.n1383 585
R994 GND.n7044 GND.n1383 585
R995 GND.n2516 GND.n2515 585
R996 GND.n2517 GND.n2516 585
R997 GND.n2513 GND.n1374 585
R998 GND.n2513 GND.n1964 585
R999 GND.n2512 GND.n1373 585
R1000 GND.n2512 GND.n2511 585
R1001 GND.n1966 GND.n1372 585
R1002 GND.n2491 GND.n1966 585
R1003 GND.n2500 GND.n2499 585
R1004 GND.n2501 GND.n2500 585
R1005 GND.n2498 GND.n1366 585
R1006 GND.n2498 GND.n2497 585
R1007 GND.n1979 GND.n1365 585
R1008 GND.n2476 GND.n1979 585
R1009 GND.n2465 GND.n1364 585
R1010 GND.n2465 GND.n2000 585
R1011 GND.n2467 GND.n2466 585
R1012 GND.n2468 GND.n2467 585
R1013 GND.n2464 GND.n1358 585
R1014 GND.n2464 GND.n2463 585
R1015 GND.n2010 GND.n1357 585
R1016 GND.n2022 GND.n2010 585
R1017 GND.n2019 GND.n1356 585
R1018 GND.n2449 GND.n2019 585
R1019 GND.n2437 GND.n2435 585
R1020 GND.n2437 GND.n2436 585
R1021 GND.n2438 GND.n1350 585
R1022 GND.n2439 GND.n2438 585
R1023 GND.n2434 GND.n1349 585
R1024 GND.n2434 GND.n2433 585
R1025 GND.n2031 GND.n1348 585
R1026 GND.n2044 GND.n2031 585
R1027 GND.n2042 GND.n2041 585
R1028 GND.n2423 GND.n2042 585
R1029 GND.n2352 GND.n1342 585
R1030 GND.n2353 GND.n2352 585
R1031 GND.n2083 GND.n1341 585
R1032 GND.n2350 GND.n2083 585
R1033 GND.n2394 GND.n1340 585
R1034 GND.n2394 GND.n2393 585
R1035 GND.n2396 GND.n2395 585
R1036 GND.n2397 GND.n2396 585
R1037 GND.n2075 GND.n1334 585
R1038 GND.n2402 GND.n2075 585
R1039 GND.n2074 GND.n1333 585
R1040 GND.n2074 GND.n2072 585
R1041 GND.n2061 GND.n1332 585
R1042 GND.n2064 GND.n2061 585
R1043 GND.n2412 GND.n2062 585
R1044 GND.n2412 GND.n2411 585
R1045 GND.n2413 GND.n1326 585
R1046 GND.n2414 GND.n2413 585
R1047 GND.n2060 GND.n1325 585
R1048 GND.n2097 GND.n2060 585
R1049 GND.n2099 GND.n1324 585
R1050 GND.n2326 GND.n2099 585
R1051 GND.n2316 GND.n2314 585
R1052 GND.n2316 GND.n2315 585
R1053 GND.n2317 GND.n1318 585
R1054 GND.n2318 GND.n2317 585
R1055 GND.n2313 GND.n1317 585
R1056 GND.n2313 GND.n2312 585
R1057 GND.n2108 GND.n1316 585
R1058 GND.n2122 GND.n2108 585
R1059 GND.n2120 GND.n2119 585
R1060 GND.n2303 GND.n2120 585
R1061 GND.n2291 GND.n1310 585
R1062 GND.n2291 GND.n2290 585
R1063 GND.n2292 GND.n1309 585
R1064 GND.n2293 GND.n2292 585
R1065 GND.n2289 GND.n1308 585
R1066 GND.n2289 GND.n2288 585
R1067 GND.n2133 GND.n2132 585
R1068 GND.n2145 GND.n2133 585
R1069 GND.n2143 GND.n1302 585
R1070 GND.n2279 GND.n2143 585
R1071 GND.n2267 GND.n1301 585
R1072 GND.n2267 GND.n2266 585
R1073 GND.n2268 GND.n1300 585
R1074 GND.n2269 GND.n2268 585
R1075 GND.n2154 GND.n2153 585
R1076 GND.n2217 GND.n2154 585
R1077 GND.n1295 GND.n1294 585
R1078 GND.n2173 GND.n1294 585
R1079 GND.n7112 GND.n7111 585
R1080 GND.n7113 GND.n7112 585
R1081 GND.n2190 GND.n1293 585
R1082 GND.n2192 GND.n2191 585
R1083 GND.n2194 GND.n2193 585
R1084 GND.n2186 GND.n2185 585
R1085 GND.n2198 GND.n2187 585
R1086 GND.n2200 GND.n2199 585
R1087 GND.n2202 GND.n2201 585
R1088 GND.n2182 GND.n2181 585
R1089 GND.n2206 GND.n2183 585
R1090 GND.n2207 GND.n2178 585
R1091 GND.n2208 GND.n1242 585
R1092 GND.n7179 GND.n1242 585
R1093 GND.n6990 GND.n6989 585
R1094 GND.n1923 GND.n1922 585
R1095 GND.n1954 GND.n1953 585
R1096 GND.n1952 GND.n1951 585
R1097 GND.n1950 GND.n1949 585
R1098 GND.n1948 GND.n1947 585
R1099 GND.n1946 GND.n1945 585
R1100 GND.n1944 GND.n1943 585
R1101 GND.n1942 GND.n1941 585
R1102 GND.n1940 GND.n1939 585
R1103 GND.n6987 GND.n1935 585
R1104 GND.n1989 GND.n1381 585
R1105 GND.n7044 GND.n1381 585
R1106 GND.n1990 GND.n1965 585
R1107 GND.n2517 GND.n1965 585
R1108 GND.n1992 GND.n1991 585
R1109 GND.n1991 GND.n1964 585
R1110 GND.n1993 GND.n1968 585
R1111 GND.n2511 GND.n1968 585
R1112 GND.n2493 GND.n2492 585
R1113 GND.n2492 GND.n2491 585
R1114 GND.n2494 GND.n1977 585
R1115 GND.n2501 GND.n1977 585
R1116 GND.n2496 GND.n2495 585
R1117 GND.n2497 GND.n2496 585
R1118 GND.n1982 GND.n1981 585
R1119 GND.n2476 GND.n1981 585
R1120 GND.n2459 GND.n2458 585
R1121 GND.n2458 GND.n2000 585
R1122 GND.n2460 GND.n2008 585
R1123 GND.n2468 GND.n2008 585
R1124 GND.n2462 GND.n2461 585
R1125 GND.n2463 GND.n2462 585
R1126 GND.n2013 GND.n2012 585
R1127 GND.n2022 GND.n2012 585
R1128 GND.n2451 GND.n2450 585
R1129 GND.n2450 GND.n2449 585
R1130 GND.n2016 GND.n2015 585
R1131 GND.n2436 GND.n2016 585
R1132 GND.n2430 GND.n2029 585
R1133 GND.n2439 GND.n2029 585
R1134 GND.n2432 GND.n2431 585
R1135 GND.n2433 GND.n2432 585
R1136 GND.n2035 GND.n2034 585
R1137 GND.n2044 GND.n2034 585
R1138 GND.n2425 GND.n2424 585
R1139 GND.n2424 GND.n2423 585
R1140 GND.n2038 GND.n2037 585
R1141 GND.n2353 GND.n2038 585
R1142 GND.n2346 GND.n2345 585
R1143 GND.n2350 GND.n2346 585
R1144 GND.n2086 GND.n2084 585
R1145 GND.n2393 GND.n2084 585
R1146 GND.n2341 GND.n2081 585
R1147 GND.n2397 GND.n2081 585
R1148 GND.n2340 GND.n2073 585
R1149 GND.n2402 GND.n2073 585
R1150 GND.n2334 GND.n2088 585
R1151 GND.n2334 GND.n2072 585
R1152 GND.n2336 GND.n2335 585
R1153 GND.n2335 GND.n2064 585
R1154 GND.n2333 GND.n2063 585
R1155 GND.n2411 GND.n2063 585
R1156 GND.n2332 GND.n2058 585
R1157 GND.n2414 GND.n2058 585
R1158 GND.n2094 GND.n2090 585
R1159 GND.n2097 GND.n2094 585
R1160 GND.n2328 GND.n2327 585
R1161 GND.n2327 GND.n2326 585
R1162 GND.n2093 GND.n2092 585
R1163 GND.n2315 GND.n2093 585
R1164 GND.n2113 GND.n2106 585
R1165 GND.n2318 GND.n2106 585
R1166 GND.n2311 GND.n2310 585
R1167 GND.n2312 GND.n2311 585
R1168 GND.n2112 GND.n2111 585
R1169 GND.n2122 GND.n2111 585
R1170 GND.n2305 GND.n2304 585
R1171 GND.n2304 GND.n2303 585
R1172 GND.n2116 GND.n2115 585
R1173 GND.n2290 GND.n2116 585
R1174 GND.n2137 GND.n2130 585
R1175 GND.n2293 GND.n2130 585
R1176 GND.n2287 GND.n2286 585
R1177 GND.n2288 GND.n2287 585
R1178 GND.n2136 GND.n2135 585
R1179 GND.n2145 GND.n2135 585
R1180 GND.n2281 GND.n2280 585
R1181 GND.n2280 GND.n2279 585
R1182 GND.n2140 GND.n2139 585
R1183 GND.n2266 GND.n2140 585
R1184 GND.n2176 GND.n2152 585
R1185 GND.n2269 GND.n2152 585
R1186 GND.n2216 GND.n2215 585
R1187 GND.n2217 GND.n2216 585
R1188 GND.n2175 GND.n2174 585
R1189 GND.n2174 GND.n2173 585
R1190 GND.n2210 GND.n1291 585
R1191 GND.n7113 GND.n1291 585
R1192 GND.n7043 GND.n7042 585
R1193 GND.n7044 GND.n7043 585
R1194 GND.n1386 GND.n1384 585
R1195 GND.n2517 GND.n1384 585
R1196 GND.n2508 GND.n1971 585
R1197 GND.n1971 GND.n1964 585
R1198 GND.n2510 GND.n2509 585
R1199 GND.n2511 GND.n2510 585
R1200 GND.n1972 GND.n1970 585
R1201 GND.n2491 GND.n1970 585
R1202 GND.n2503 GND.n2502 585
R1203 GND.n2502 GND.n2501 585
R1204 GND.n1975 GND.n1974 585
R1205 GND.n2497 GND.n1975 585
R1206 GND.n2475 GND.n2474 585
R1207 GND.n2476 GND.n2475 585
R1208 GND.n2003 GND.n2002 585
R1209 GND.n2002 GND.n2000 585
R1210 GND.n2470 GND.n2469 585
R1211 GND.n2469 GND.n2468 585
R1212 GND.n2006 GND.n2005 585
R1213 GND.n2463 GND.n2006 585
R1214 GND.n2446 GND.n2023 585
R1215 GND.n2023 GND.n2022 585
R1216 GND.n2448 GND.n2447 585
R1217 GND.n2449 GND.n2448 585
R1218 GND.n2024 GND.n2020 585
R1219 GND.n2436 GND.n2020 585
R1220 GND.n2441 GND.n2440 585
R1221 GND.n2440 GND.n2439 585
R1222 GND.n2027 GND.n2026 585
R1223 GND.n2433 GND.n2027 585
R1224 GND.n2420 GND.n2045 585
R1225 GND.n2045 GND.n2044 585
R1226 GND.n2422 GND.n2421 585
R1227 GND.n2423 GND.n2422 585
R1228 GND.n2046 GND.n2043 585
R1229 GND.n2353 GND.n2043 585
R1230 GND.n2349 GND.n2348 585
R1231 GND.n2350 GND.n2349 585
R1232 GND.n2347 GND.n2079 585
R1233 GND.n2393 GND.n2079 585
R1234 GND.n2399 GND.n2398 585
R1235 GND.n2398 GND.n2397 585
R1236 GND.n2401 GND.n2400 585
R1237 GND.n2402 GND.n2401 585
R1238 GND.n2078 GND.n2077 585
R1239 GND.n2078 GND.n2072 585
R1240 GND.n2076 GND.n2052 585
R1241 GND.n2076 GND.n2064 585
R1242 GND.n2056 GND.n2053 585
R1243 GND.n2411 GND.n2056 585
R1244 GND.n2416 GND.n2415 585
R1245 GND.n2415 GND.n2414 585
R1246 GND.n2055 GND.n2054 585
R1247 GND.n2097 GND.n2055 585
R1248 GND.n2325 GND.n2324 585
R1249 GND.n2326 GND.n2325 585
R1250 GND.n2101 GND.n2100 585
R1251 GND.n2315 GND.n2100 585
R1252 GND.n2320 GND.n2319 585
R1253 GND.n2319 GND.n2318 585
R1254 GND.n2104 GND.n2103 585
R1255 GND.n2312 GND.n2104 585
R1256 GND.n2300 GND.n2123 585
R1257 GND.n2123 GND.n2122 585
R1258 GND.n2302 GND.n2301 585
R1259 GND.n2303 GND.n2302 585
R1260 GND.n2124 GND.n2121 585
R1261 GND.n2290 GND.n2121 585
R1262 GND.n2295 GND.n2294 585
R1263 GND.n2294 GND.n2293 585
R1264 GND.n2127 GND.n2126 585
R1265 GND.n2288 GND.n2127 585
R1266 GND.n2276 GND.n2146 585
R1267 GND.n2146 GND.n2145 585
R1268 GND.n2278 GND.n2277 585
R1269 GND.n2279 GND.n2278 585
R1270 GND.n2147 GND.n2144 585
R1271 GND.n2266 GND.n2144 585
R1272 GND.n2271 GND.n2270 585
R1273 GND.n2270 GND.n2269 585
R1274 GND.n2150 GND.n2149 585
R1275 GND.n2217 GND.n2150 585
R1276 GND.n2172 GND.n2171 585
R1277 GND.n2173 GND.n2172 585
R1278 GND.n2168 GND.n1246 585
R1279 GND.n7113 GND.n1246 585
R1280 GND.n7177 GND.n7176 585
R1281 GND.n7175 GND.n1245 585
R1282 GND.n7174 GND.n1244 585
R1283 GND.n7179 GND.n1244 585
R1284 GND.n7173 GND.n7172 585
R1285 GND.n7171 GND.n7170 585
R1286 GND.n7169 GND.n7168 585
R1287 GND.n7167 GND.n7166 585
R1288 GND.n7165 GND.n7164 585
R1289 GND.n7163 GND.n7162 585
R1290 GND.n7161 GND.n7160 585
R1291 GND.n7159 GND.n7158 585
R1292 GND.n7157 GND.n7156 585
R1293 GND.n7155 GND.n7154 585
R1294 GND.n7153 GND.n7152 585
R1295 GND.n7151 GND.n7150 585
R1296 GND.n7149 GND.n7148 585
R1297 GND.n7147 GND.n7146 585
R1298 GND.n7145 GND.n7144 585
R1299 GND.n7143 GND.n7142 585
R1300 GND.n7141 GND.n7140 585
R1301 GND.n7139 GND.n1269 585
R1302 GND.n7138 GND.n7137 585
R1303 GND.n7136 GND.n7135 585
R1304 GND.n7134 GND.n7133 585
R1305 GND.n7132 GND.n7131 585
R1306 GND.n7130 GND.n7129 585
R1307 GND.n7128 GND.n7127 585
R1308 GND.n7126 GND.n7125 585
R1309 GND.n7124 GND.n7123 585
R1310 GND.n7122 GND.n7121 585
R1311 GND.n7120 GND.n1282 585
R1312 GND.n1286 GND.n1283 585
R1313 GND.n7116 GND.n7115 585
R1314 GND.n6994 GND.n1379 585
R1315 GND.n6995 GND.n1433 585
R1316 GND.n6996 GND.n1429 585
R1317 GND.n6997 GND.n1428 585
R1318 GND.n6975 GND.n1426 585
R1319 GND.n7001 GND.n1425 585
R1320 GND.n7002 GND.n1424 585
R1321 GND.n7003 GND.n1423 585
R1322 GND.n6978 GND.n1421 585
R1323 GND.n7007 GND.n1420 585
R1324 GND.n7008 GND.n1419 585
R1325 GND.n7009 GND.n1418 585
R1326 GND.n6981 GND.n1416 585
R1327 GND.n7013 GND.n1413 585
R1328 GND.n7014 GND.n1412 585
R1329 GND.n7015 GND.n1411 585
R1330 GND.n6984 GND.n1409 585
R1331 GND.n7019 GND.n1408 585
R1332 GND.n6987 GND.n6986 585
R1333 GND.n7021 GND.n1405 585
R1334 GND.n1932 GND.n1403 585
R1335 GND.n7025 GND.n1402 585
R1336 GND.n7026 GND.n1401 585
R1337 GND.n7027 GND.n1398 585
R1338 GND.n1929 GND.n1396 585
R1339 GND.n7031 GND.n1395 585
R1340 GND.n7032 GND.n1394 585
R1341 GND.n7033 GND.n1393 585
R1342 GND.n1926 GND.n1391 585
R1343 GND.n7037 GND.n1390 585
R1344 GND.n7038 GND.n1389 585
R1345 GND.n7039 GND.n1385 585
R1346 GND.n7046 GND.n7045 585
R1347 GND.n7045 GND.n7044 585
R1348 GND.n7047 GND.n1377 585
R1349 GND.n2517 GND.n1377 585
R1350 GND.n7048 GND.n1376 585
R1351 GND.n1964 GND.n1376 585
R1352 GND.n1967 GND.n1371 585
R1353 GND.n2511 GND.n1967 585
R1354 GND.n7052 GND.n1370 585
R1355 GND.n2491 GND.n1370 585
R1356 GND.n7053 GND.n1369 585
R1357 GND.n2501 GND.n1369 585
R1358 GND.n7054 GND.n1368 585
R1359 GND.n2497 GND.n1368 585
R1360 GND.n2001 GND.n1363 585
R1361 GND.n2476 GND.n2001 585
R1362 GND.n7058 GND.n1362 585
R1363 GND.n2000 GND.n1362 585
R1364 GND.n7059 GND.n1361 585
R1365 GND.n2468 GND.n1361 585
R1366 GND.n7060 GND.n1360 585
R1367 GND.n2463 GND.n1360 585
R1368 GND.n2021 GND.n1355 585
R1369 GND.n2022 GND.n2021 585
R1370 GND.n7064 GND.n1354 585
R1371 GND.n2449 GND.n1354 585
R1372 GND.n7065 GND.n1353 585
R1373 GND.n2436 GND.n1353 585
R1374 GND.n7066 GND.n1352 585
R1375 GND.n2439 GND.n1352 585
R1376 GND.n2033 GND.n1347 585
R1377 GND.n2433 GND.n2033 585
R1378 GND.n7070 GND.n1346 585
R1379 GND.n2044 GND.n1346 585
R1380 GND.n7071 GND.n1345 585
R1381 GND.n2423 GND.n1345 585
R1382 GND.n7072 GND.n1344 585
R1383 GND.n2353 GND.n1344 585
R1384 GND.n2085 GND.n1339 585
R1385 GND.n2350 GND.n2085 585
R1386 GND.n7076 GND.n1338 585
R1387 GND.n2393 GND.n1338 585
R1388 GND.n7077 GND.n1337 585
R1389 GND.n2397 GND.n1337 585
R1390 GND.n7078 GND.n1336 585
R1391 GND.n2402 GND.n1336 585
R1392 GND.n2071 GND.n1331 585
R1393 GND.n2072 GND.n2071 585
R1394 GND.n7082 GND.n1330 585
R1395 GND.n2064 GND.n1330 585
R1396 GND.n7083 GND.n1329 585
R1397 GND.n2411 GND.n1329 585
R1398 GND.n7084 GND.n1328 585
R1399 GND.n2414 GND.n1328 585
R1400 GND.n2096 GND.n1323 585
R1401 GND.n2097 GND.n2096 585
R1402 GND.n7088 GND.n1322 585
R1403 GND.n2326 GND.n1322 585
R1404 GND.n7089 GND.n1321 585
R1405 GND.n2315 GND.n1321 585
R1406 GND.n7090 GND.n1320 585
R1407 GND.n2318 GND.n1320 585
R1408 GND.n2110 GND.n1315 585
R1409 GND.n2312 GND.n2110 585
R1410 GND.n7094 GND.n1314 585
R1411 GND.n2122 GND.n1314 585
R1412 GND.n7095 GND.n1313 585
R1413 GND.n2303 GND.n1313 585
R1414 GND.n7096 GND.n1312 585
R1415 GND.n2290 GND.n1312 585
R1416 GND.n2129 GND.n1307 585
R1417 GND.n2293 GND.n2129 585
R1418 GND.n7100 GND.n1306 585
R1419 GND.n2288 GND.n1306 585
R1420 GND.n7101 GND.n1305 585
R1421 GND.n2145 GND.n1305 585
R1422 GND.n7102 GND.n1304 585
R1423 GND.n2279 GND.n1304 585
R1424 GND.n2265 GND.n1299 585
R1425 GND.n2266 GND.n2265 585
R1426 GND.n7106 GND.n1298 585
R1427 GND.n2269 GND.n1298 585
R1428 GND.n7107 GND.n1297 585
R1429 GND.n2217 GND.n1297 585
R1430 GND.n7108 GND.n1288 585
R1431 GND.n2173 GND.n1288 585
R1432 GND.n7114 GND.n1289 585
R1433 GND.n7114 GND.n7113 585
R1434 GND.n8450 GND.n247 585
R1435 GND.n8446 GND.n247 585
R1436 GND.n8452 GND.n8451 585
R1437 GND.n8453 GND.n8452 585
R1438 GND.n232 GND.n231 585
R1439 GND.n6302 GND.n232 585
R1440 GND.n8461 GND.n8460 585
R1441 GND.n8460 GND.n8459 585
R1442 GND.n8462 GND.n227 585
R1443 GND.n6335 GND.n227 585
R1444 GND.n8464 GND.n8463 585
R1445 GND.n8465 GND.n8464 585
R1446 GND.n211 GND.n210 585
R1447 GND.n6341 GND.n211 585
R1448 GND.n8473 GND.n8472 585
R1449 GND.n8472 GND.n8471 585
R1450 GND.n8474 GND.n206 585
R1451 GND.n6347 GND.n206 585
R1452 GND.n8476 GND.n8475 585
R1453 GND.n8477 GND.n8476 585
R1454 GND.n191 GND.n190 585
R1455 GND.n6353 GND.n191 585
R1456 GND.n8485 GND.n8484 585
R1457 GND.n8484 GND.n8483 585
R1458 GND.n8486 GND.n186 585
R1459 GND.n6239 GND.n186 585
R1460 GND.n8488 GND.n8487 585
R1461 GND.n8489 GND.n8488 585
R1462 GND.n171 GND.n170 585
R1463 GND.n6230 GND.n171 585
R1464 GND.n8497 GND.n8496 585
R1465 GND.n8496 GND.n8495 585
R1466 GND.n8498 GND.n165 585
R1467 GND.n6223 GND.n165 585
R1468 GND.n8500 GND.n8499 585
R1469 GND.n8501 GND.n8500 585
R1470 GND.n166 GND.n164 585
R1471 GND.n6215 GND.n164 585
R1472 GND.n5940 GND.n5939 585
R1473 GND.n5944 GND.n5940 585
R1474 GND.n6375 GND.n6374 585
R1475 GND.n6374 GND.n6373 585
R1476 GND.n6376 GND.n144 585
R1477 GND.n8508 GND.n144 585
R1478 GND.n6378 GND.n6377 585
R1479 GND.n6379 GND.n6378 585
R1480 GND.n5935 GND.n5934 585
R1481 GND.n5934 GND.n5926 585
R1482 GND.n5917 GND.n5916 585
R1483 GND.n6388 GND.n5917 585
R1484 GND.n6394 GND.n6393 585
R1485 GND.n6393 GND.n6392 585
R1486 GND.n6395 GND.n5912 585
R1487 GND.n6198 GND.n5912 585
R1488 GND.n6397 GND.n6396 585
R1489 GND.n6398 GND.n6397 585
R1490 GND.n5898 GND.n5897 585
R1491 GND.n6183 GND.n5898 585
R1492 GND.n6406 GND.n6405 585
R1493 GND.n6405 GND.n6404 585
R1494 GND.n6407 GND.n5893 585
R1495 GND.n6176 GND.n5893 585
R1496 GND.n6409 GND.n6408 585
R1497 GND.n6410 GND.n6409 585
R1498 GND.n5877 GND.n5876 585
R1499 GND.n6168 GND.n5877 585
R1500 GND.n6418 GND.n6417 585
R1501 GND.n6417 GND.n6416 585
R1502 GND.n6419 GND.n5872 585
R1503 GND.n6161 GND.n5872 585
R1504 GND.n6421 GND.n6420 585
R1505 GND.n6422 GND.n6421 585
R1506 GND.n5856 GND.n5855 585
R1507 GND.n6153 GND.n5856 585
R1508 GND.n6430 GND.n6429 585
R1509 GND.n6429 GND.n6428 585
R1510 GND.n6431 GND.n5849 585
R1511 GND.n6146 GND.n5849 585
R1512 GND.n6433 GND.n6432 585
R1513 GND.n6434 GND.n6433 585
R1514 GND.n5850 GND.n5848 585
R1515 GND.n6138 GND.n5848 585
R1516 GND.n5832 GND.n5825 585
R1517 GND.n6440 GND.n5832 585
R1518 GND.n6445 GND.n5823 585
R1519 GND.n6051 GND.n5823 585
R1520 GND.n6447 GND.n6446 585
R1521 GND.n6448 GND.n6447 585
R1522 GND.n6132 GND.n5822 585
R1523 GND.n6131 GND.n6130 585
R1524 GND.n6129 GND.n6128 585
R1525 GND.n6127 GND.n6126 585
R1526 GND.n6125 GND.n6124 585
R1527 GND.n6123 GND.n6122 585
R1528 GND.n6121 GND.n6120 585
R1529 GND.n6119 GND.n6118 585
R1530 GND.n6117 GND.n6116 585
R1531 GND.n6115 GND.n6112 585
R1532 GND.n6512 GND.n3066 585
R1533 GND.n6295 GND.n6294 585
R1534 GND.n6292 GND.n6260 585
R1535 GND.n6291 GND.n6290 585
R1536 GND.n6284 GND.n6262 585
R1537 GND.n6286 GND.n6285 585
R1538 GND.n6282 GND.n6264 585
R1539 GND.n6281 GND.n6280 585
R1540 GND.n6274 GND.n6266 585
R1541 GND.n6276 GND.n6275 585
R1542 GND.n6272 GND.n6268 585
R1543 GND.n6271 GND.n6270 585
R1544 GND.n6271 GND.n383 585
R1545 GND.n6298 GND.n252 585
R1546 GND.n8446 GND.n252 585
R1547 GND.n6299 GND.n245 585
R1548 GND.n8453 GND.n245 585
R1549 GND.n6301 GND.n6300 585
R1550 GND.n6302 GND.n6301 585
R1551 GND.n6252 GND.n234 585
R1552 GND.n8459 GND.n234 585
R1553 GND.n6337 GND.n6336 585
R1554 GND.n6336 GND.n6335 585
R1555 GND.n6338 GND.n225 585
R1556 GND.n8465 GND.n225 585
R1557 GND.n6340 GND.n6339 585
R1558 GND.n6341 GND.n6340 585
R1559 GND.n5964 GND.n214 585
R1560 GND.n8471 GND.n214 585
R1561 GND.n6349 GND.n6348 585
R1562 GND.n6348 GND.n6347 585
R1563 GND.n6350 GND.n204 585
R1564 GND.n8477 GND.n204 585
R1565 GND.n6352 GND.n6351 585
R1566 GND.n6353 GND.n6352 585
R1567 GND.n5960 GND.n194 585
R1568 GND.n8483 GND.n194 585
R1569 GND.n6238 GND.n6237 585
R1570 GND.n6239 GND.n6238 585
R1571 GND.n5966 GND.n184 585
R1572 GND.n8489 GND.n184 585
R1573 GND.n6232 GND.n6231 585
R1574 GND.n6231 GND.n6230 585
R1575 GND.n5968 GND.n174 585
R1576 GND.n8495 GND.n174 585
R1577 GND.n6222 GND.n6221 585
R1578 GND.n6223 GND.n6222 585
R1579 GND.n5970 GND.n162 585
R1580 GND.n8501 GND.n162 585
R1581 GND.n6217 GND.n6216 585
R1582 GND.n6216 GND.n6215 585
R1583 GND.n5973 GND.n5972 585
R1584 GND.n5973 GND.n5944 585
R1585 GND.n141 GND.n139 585
R1586 GND.n6373 GND.n141 585
R1587 GND.n8510 GND.n8509 585
R1588 GND.n8509 GND.n8508 585
R1589 GND.n140 GND.n138 585
R1590 GND.n6379 GND.n140 585
R1591 GND.n6193 GND.n6192 585
R1592 GND.n6192 GND.n5926 585
R1593 GND.n6194 GND.n5925 585
R1594 GND.n6388 GND.n5925 585
R1595 GND.n6195 GND.n5920 585
R1596 GND.n6392 GND.n5920 585
R1597 GND.n6197 GND.n6196 585
R1598 GND.n6198 GND.n6197 585
R1599 GND.n6036 GND.n5911 585
R1600 GND.n6398 GND.n5911 585
R1601 GND.n6185 GND.n6184 585
R1602 GND.n6184 GND.n6183 585
R1603 GND.n6038 GND.n5901 585
R1604 GND.n6404 GND.n5901 585
R1605 GND.n6175 GND.n6174 585
R1606 GND.n6176 GND.n6175 585
R1607 GND.n6040 GND.n5891 585
R1608 GND.n6410 GND.n5891 585
R1609 GND.n6170 GND.n6169 585
R1610 GND.n6169 GND.n6168 585
R1611 GND.n6042 GND.n5880 585
R1612 GND.n6416 GND.n5880 585
R1613 GND.n6160 GND.n6159 585
R1614 GND.n6161 GND.n6160 585
R1615 GND.n6044 GND.n5870 585
R1616 GND.n6422 GND.n5870 585
R1617 GND.n6155 GND.n6154 585
R1618 GND.n6154 GND.n6153 585
R1619 GND.n6046 GND.n5859 585
R1620 GND.n6428 GND.n5859 585
R1621 GND.n6145 GND.n6144 585
R1622 GND.n6146 GND.n6145 585
R1623 GND.n6048 GND.n5846 585
R1624 GND.n6434 GND.n5846 585
R1625 GND.n6140 GND.n6139 585
R1626 GND.n6139 GND.n6138 585
R1627 GND.n6137 GND.n5830 585
R1628 GND.n6440 GND.n5830 585
R1629 GND.n6136 GND.n6052 585
R1630 GND.n6052 GND.n6051 585
R1631 GND.n6050 GND.n5820 585
R1632 GND.n6448 GND.n5820 585
R1633 GND.n242 GND.n241 585
R1634 GND.n8446 GND.n242 585
R1635 GND.n8455 GND.n8454 585
R1636 GND.n8454 GND.n8453 585
R1637 GND.n8456 GND.n236 585
R1638 GND.n6302 GND.n236 585
R1639 GND.n8458 GND.n8457 585
R1640 GND.n8459 GND.n8458 585
R1641 GND.n222 GND.n221 585
R1642 GND.n6335 GND.n222 585
R1643 GND.n8467 GND.n8466 585
R1644 GND.n8466 GND.n8465 585
R1645 GND.n8468 GND.n216 585
R1646 GND.n6341 GND.n216 585
R1647 GND.n8470 GND.n8469 585
R1648 GND.n8471 GND.n8470 585
R1649 GND.n201 GND.n200 585
R1650 GND.n6347 GND.n201 585
R1651 GND.n8479 GND.n8478 585
R1652 GND.n8478 GND.n8477 585
R1653 GND.n8480 GND.n195 585
R1654 GND.n6353 GND.n195 585
R1655 GND.n8482 GND.n8481 585
R1656 GND.n8483 GND.n8482 585
R1657 GND.n181 GND.n180 585
R1658 GND.n6239 GND.n181 585
R1659 GND.n8491 GND.n8490 585
R1660 GND.n8490 GND.n8489 585
R1661 GND.n8492 GND.n176 585
R1662 GND.n6230 GND.n176 585
R1663 GND.n8494 GND.n8493 585
R1664 GND.n8495 GND.n8494 585
R1665 GND.n159 GND.n157 585
R1666 GND.n6223 GND.n159 585
R1667 GND.n8503 GND.n8502 585
R1668 GND.n8502 GND.n8501 585
R1669 GND.n158 GND.n156 585
R1670 GND.n6215 GND.n158 585
R1671 GND.n5943 GND.n5942 585
R1672 GND.n5944 GND.n5943 585
R1673 GND.n148 GND.n146 585
R1674 GND.n6373 GND.n146 585
R1675 GND.n8507 GND.n8506 585
R1676 GND.n8508 GND.n8507 585
R1677 GND.n147 GND.n145 585
R1678 GND.n6379 GND.n145 585
R1679 GND.n5923 GND.n5922 585
R1680 GND.n5926 GND.n5923 585
R1681 GND.n6389 GND.n154 585
R1682 GND.n6389 GND.n6388 585
R1683 GND.n6391 GND.n6390 585
R1684 GND.n6392 GND.n6391 585
R1685 GND.n5908 GND.n5907 585
R1686 GND.n6198 GND.n5908 585
R1687 GND.n6400 GND.n6399 585
R1688 GND.n6399 GND.n6398 585
R1689 GND.n6401 GND.n5903 585
R1690 GND.n6183 GND.n5903 585
R1691 GND.n6403 GND.n6402 585
R1692 GND.n6404 GND.n6403 585
R1693 GND.n5888 GND.n5887 585
R1694 GND.n6176 GND.n5888 585
R1695 GND.n6412 GND.n6411 585
R1696 GND.n6411 GND.n6410 585
R1697 GND.n6413 GND.n5882 585
R1698 GND.n6168 GND.n5882 585
R1699 GND.n6415 GND.n6414 585
R1700 GND.n6416 GND.n6415 585
R1701 GND.n5867 GND.n5866 585
R1702 GND.n6161 GND.n5867 585
R1703 GND.n6424 GND.n6423 585
R1704 GND.n6423 GND.n6422 585
R1705 GND.n6425 GND.n5861 585
R1706 GND.n6153 GND.n5861 585
R1707 GND.n6427 GND.n6426 585
R1708 GND.n6428 GND.n6427 585
R1709 GND.n5843 GND.n5842 585
R1710 GND.n6146 GND.n5843 585
R1711 GND.n6436 GND.n6435 585
R1712 GND.n6435 GND.n6434 585
R1713 GND.n6437 GND.n5834 585
R1714 GND.n6138 GND.n5834 585
R1715 GND.n6439 GND.n6438 585
R1716 GND.n6440 GND.n6439 585
R1717 GND.n5835 GND.n5833 585
R1718 GND.n6051 GND.n5833 585
R1719 GND.n5836 GND.n3070 585
R1720 GND.n6448 GND.n3070 585
R1721 GND.n6510 GND.n6509 585
R1722 GND.n6508 GND.n3069 585
R1723 GND.n6507 GND.n3068 585
R1724 GND.n6512 GND.n3068 585
R1725 GND.n6506 GND.n6505 585
R1726 GND.n6504 GND.n6503 585
R1727 GND.n6502 GND.n6501 585
R1728 GND.n6500 GND.n6499 585
R1729 GND.n6498 GND.n6497 585
R1730 GND.n6496 GND.n6495 585
R1731 GND.n6494 GND.n6493 585
R1732 GND.n6492 GND.n6491 585
R1733 GND.n6490 GND.n6489 585
R1734 GND.n6488 GND.n6487 585
R1735 GND.n6486 GND.n6485 585
R1736 GND.n6485 GND.n5791 585
R1737 GND.n6484 GND.n6483 585
R1738 GND.n6482 GND.n6481 585
R1739 GND.n6480 GND.n6479 585
R1740 GND.n6478 GND.n6477 585
R1741 GND.n6476 GND.n6475 585
R1742 GND.n6474 GND.n5798 585
R1743 GND.n6473 GND.n6472 585
R1744 GND.n6471 GND.n6470 585
R1745 GND.n6469 GND.n6468 585
R1746 GND.n6467 GND.n6466 585
R1747 GND.n6465 GND.n6464 585
R1748 GND.n6463 GND.n6462 585
R1749 GND.n6461 GND.n6460 585
R1750 GND.n6459 GND.n6458 585
R1751 GND.n6457 GND.n6456 585
R1752 GND.n6455 GND.n5811 585
R1753 GND.n5815 GND.n5812 585
R1754 GND.n6451 GND.n6450 585
R1755 GND.n311 GND.n251 585
R1756 GND.n317 GND.n316 585
R1757 GND.n319 GND.n318 585
R1758 GND.n321 GND.n320 585
R1759 GND.n323 GND.n322 585
R1760 GND.n325 GND.n324 585
R1761 GND.n327 GND.n326 585
R1762 GND.n329 GND.n328 585
R1763 GND.n331 GND.n330 585
R1764 GND.n333 GND.n332 585
R1765 GND.n335 GND.n334 585
R1766 GND.n301 GND.n298 585
R1767 GND.n339 GND.n302 585
R1768 GND.n341 GND.n340 585
R1769 GND.n343 GND.n342 585
R1770 GND.n345 GND.n344 585
R1771 GND.n347 GND.n346 585
R1772 GND.n349 GND.n348 585
R1773 GND.n351 GND.n350 585
R1774 GND.n353 GND.n352 585
R1775 GND.n355 GND.n354 585
R1776 GND.n358 GND.n357 585
R1777 GND.n356 GND.n287 585
R1778 GND.n363 GND.n362 585
R1779 GND.n365 GND.n364 585
R1780 GND.n367 GND.n366 585
R1781 GND.n369 GND.n368 585
R1782 GND.n371 GND.n370 585
R1783 GND.n373 GND.n372 585
R1784 GND.n376 GND.n375 585
R1785 GND.n374 GND.n281 585
R1786 GND.n380 GND.n278 585
R1787 GND.n382 GND.n381 585
R1788 GND.n383 GND.n382 585
R1789 GND.n8448 GND.n8447 585
R1790 GND.n8447 GND.n8446 585
R1791 GND.n250 GND.n244 585
R1792 GND.n8453 GND.n244 585
R1793 GND.n6304 GND.n6303 585
R1794 GND.n6303 GND.n6302 585
R1795 GND.n6305 GND.n233 585
R1796 GND.n8459 GND.n233 585
R1797 GND.n6307 GND.n6306 585
R1798 GND.n6335 GND.n6307 585
R1799 GND.n6247 GND.n224 585
R1800 GND.n8465 GND.n224 585
R1801 GND.n6343 GND.n6342 585
R1802 GND.n6342 GND.n6341 585
R1803 GND.n6344 GND.n213 585
R1804 GND.n8471 GND.n213 585
R1805 GND.n6346 GND.n6345 585
R1806 GND.n6347 GND.n6346 585
R1807 GND.n6245 GND.n203 585
R1808 GND.n8477 GND.n203 585
R1809 GND.n6244 GND.n5959 585
R1810 GND.n6353 GND.n5959 585
R1811 GND.n6242 GND.n193 585
R1812 GND.n8483 GND.n193 585
R1813 GND.n6241 GND.n6240 585
R1814 GND.n6240 GND.n6239 585
R1815 GND.n5965 GND.n183 585
R1816 GND.n8489 GND.n183 585
R1817 GND.n6229 GND.n6228 585
R1818 GND.n6230 GND.n6229 585
R1819 GND.n6226 GND.n173 585
R1820 GND.n8495 GND.n173 585
R1821 GND.n6225 GND.n6224 585
R1822 GND.n6224 GND.n6223 585
R1823 GND.n5969 GND.n161 585
R1824 GND.n8501 GND.n161 585
R1825 GND.n6214 GND.n6213 585
R1826 GND.n6215 GND.n6214 585
R1827 GND.n6210 GND.n5975 585
R1828 GND.n5975 GND.n5944 585
R1829 GND.n6209 GND.n5941 585
R1830 GND.n6373 GND.n5941 585
R1831 GND.n6208 GND.n142 585
R1832 GND.n8508 GND.n142 585
R1833 GND.n6207 GND.n5933 585
R1834 GND.n6379 GND.n5933 585
R1835 GND.n6206 GND.n6205 585
R1836 GND.n6205 GND.n5926 585
R1837 GND.n6202 GND.n5924 585
R1838 GND.n6388 GND.n5924 585
R1839 GND.n6201 GND.n5919 585
R1840 GND.n6392 GND.n5919 585
R1841 GND.n6200 GND.n6199 585
R1842 GND.n6199 GND.n6198 585
R1843 GND.n5976 GND.n5910 585
R1844 GND.n6398 GND.n5910 585
R1845 GND.n6182 GND.n6181 585
R1846 GND.n6183 GND.n6182 585
R1847 GND.n6179 GND.n5900 585
R1848 GND.n6404 GND.n5900 585
R1849 GND.n6178 GND.n6177 585
R1850 GND.n6177 GND.n6176 585
R1851 GND.n6039 GND.n5890 585
R1852 GND.n6410 GND.n5890 585
R1853 GND.n6167 GND.n6166 585
R1854 GND.n6168 GND.n6167 585
R1855 GND.n6164 GND.n5879 585
R1856 GND.n6416 GND.n5879 585
R1857 GND.n6163 GND.n6162 585
R1858 GND.n6162 GND.n6161 585
R1859 GND.n6043 GND.n5869 585
R1860 GND.n6422 GND.n5869 585
R1861 GND.n6152 GND.n6151 585
R1862 GND.n6153 GND.n6152 585
R1863 GND.n6149 GND.n5858 585
R1864 GND.n6428 GND.n5858 585
R1865 GND.n6148 GND.n6147 585
R1866 GND.n6147 GND.n6146 585
R1867 GND.n6047 GND.n5845 585
R1868 GND.n6434 GND.n5845 585
R1869 GND.n5828 GND.n5827 585
R1870 GND.n6138 GND.n5828 585
R1871 GND.n6442 GND.n6441 585
R1872 GND.n6441 GND.n6440 585
R1873 GND.n6443 GND.n5817 585
R1874 GND.n6051 GND.n5817 585
R1875 GND.n6449 GND.n5818 585
R1876 GND.n6449 GND.n6448 585
R1877 GND.n3026 GND.n3025 585
R1878 GND.n5728 GND.n3026 585
R1879 GND.n6530 GND.n6529 585
R1880 GND.n6529 GND.n6528 585
R1881 GND.n6531 GND.n3023 585
R1882 GND.n3028 GND.n3023 585
R1883 GND.n6533 GND.n6532 585
R1884 GND.n6534 GND.n6533 585
R1885 GND.n3024 GND.n3022 585
R1886 GND.n3022 GND.n3020 585
R1887 GND.n5716 GND.n5715 585
R1888 GND.n5717 GND.n5716 585
R1889 GND.n3009 GND.n3008 585
R1890 GND.n3012 GND.n3009 585
R1891 GND.n6544 GND.n6543 585
R1892 GND.n6543 GND.n6542 585
R1893 GND.n6545 GND.n3006 585
R1894 GND.n3010 GND.n3006 585
R1895 GND.n6547 GND.n6546 585
R1896 GND.n6548 GND.n6547 585
R1897 GND.n3007 GND.n3005 585
R1898 GND.n3005 GND.n3002 585
R1899 GND.n5703 GND.n5702 585
R1900 GND.n5704 GND.n5703 585
R1901 GND.n2992 GND.n2991 585
R1902 GND.n2994 GND.n2992 585
R1903 GND.n6558 GND.n6557 585
R1904 GND.n6557 GND.n6556 585
R1905 GND.n6559 GND.n2989 585
R1906 GND.n5695 GND.n2989 585
R1907 GND.n6561 GND.n6560 585
R1908 GND.n6562 GND.n6561 585
R1909 GND.n2990 GND.n2988 585
R1910 GND.n2988 GND.n2985 585
R1911 GND.n5689 GND.n5688 585
R1912 GND.n5690 GND.n5689 585
R1913 GND.n2974 GND.n2973 585
R1914 GND.n2977 GND.n2974 585
R1915 GND.n6572 GND.n6571 585
R1916 GND.n6571 GND.n6570 585
R1917 GND.n6573 GND.n2971 585
R1918 GND.n2975 GND.n2971 585
R1919 GND.n6575 GND.n6574 585
R1920 GND.n6576 GND.n6575 585
R1921 GND.n2972 GND.n2970 585
R1922 GND.n2970 GND.n2967 585
R1923 GND.n5676 GND.n5675 585
R1924 GND.n5677 GND.n5676 585
R1925 GND.n2956 GND.n2955 585
R1926 GND.n2959 GND.n2956 585
R1927 GND.n6586 GND.n6585 585
R1928 GND.n6585 GND.n6584 585
R1929 GND.n6587 GND.n2953 585
R1930 GND.n2953 GND.n2951 585
R1931 GND.n6589 GND.n6588 585
R1932 GND.n6590 GND.n6589 585
R1933 GND.n2954 GND.n2952 585
R1934 GND.n2952 GND.n2949 585
R1935 GND.n5663 GND.n5662 585
R1936 GND.n5664 GND.n5663 585
R1937 GND.n2938 GND.n2937 585
R1938 GND.n2941 GND.n2938 585
R1939 GND.n6600 GND.n6599 585
R1940 GND.n6599 GND.n6598 585
R1941 GND.n6601 GND.n2935 585
R1942 GND.n2935 GND.n2933 585
R1943 GND.n6603 GND.n6602 585
R1944 GND.n6604 GND.n6603 585
R1945 GND.n2936 GND.n2934 585
R1946 GND.n2934 GND.n2931 585
R1947 GND.n5650 GND.n5649 585
R1948 GND.n5651 GND.n5650 585
R1949 GND.n2920 GND.n2919 585
R1950 GND.n2923 GND.n2920 585
R1951 GND.n6614 GND.n6613 585
R1952 GND.n6613 GND.n6612 585
R1953 GND.n6615 GND.n2917 585
R1954 GND.n5642 GND.n2917 585
R1955 GND.n6617 GND.n6616 585
R1956 GND.n6618 GND.n6617 585
R1957 GND.n2918 GND.n2916 585
R1958 GND.n2916 GND.n2914 585
R1959 GND.n5636 GND.n5635 585
R1960 GND.n5637 GND.n5636 585
R1961 GND.n5634 GND.n3236 585
R1962 GND.n3236 GND.n2905 585
R1963 GND.n5633 GND.n5632 585
R1964 GND.n5632 GND.n2904 585
R1965 GND.n5631 GND.n3237 585
R1966 GND.n5631 GND.n5630 585
R1967 GND.n5618 GND.n3238 585
R1968 GND.n5577 GND.n3238 585
R1969 GND.n5620 GND.n5619 585
R1970 GND.n5621 GND.n5620 585
R1971 GND.n5617 GND.n3246 585
R1972 GND.n5611 GND.n3246 585
R1973 GND.n5616 GND.n5615 585
R1974 GND.n5615 GND.n5614 585
R1975 GND.n3248 GND.n3247 585
R1976 GND.n5587 GND.n3248 585
R1977 GND.n5600 GND.n5599 585
R1978 GND.n5601 GND.n5600 585
R1979 GND.n5598 GND.n3260 585
R1980 GND.n5593 GND.n3260 585
R1981 GND.n5597 GND.n5596 585
R1982 GND.n5596 GND.n5595 585
R1983 GND.n3262 GND.n3261 585
R1984 GND.n5562 GND.n3262 585
R1985 GND.n5553 GND.n3281 585
R1986 GND.n3281 GND.n3273 585
R1987 GND.n5555 GND.n5554 585
R1988 GND.n5556 GND.n5555 585
R1989 GND.n5552 GND.n3280 585
R1990 GND.n3286 GND.n3280 585
R1991 GND.n5551 GND.n5550 585
R1992 GND.n5550 GND.n5549 585
R1993 GND.n3283 GND.n3282 585
R1994 GND.n5459 GND.n3283 585
R1995 GND.n5534 GND.n5533 585
R1996 GND.n5535 GND.n5534 585
R1997 GND.n5532 GND.n3297 585
R1998 GND.n3297 GND.n3293 585
R1999 GND.n5531 GND.n5530 585
R2000 GND.n5530 GND.n5529 585
R2001 GND.n3299 GND.n3298 585
R2002 GND.n5466 GND.n3299 585
R2003 GND.n5506 GND.n5505 585
R2004 GND.n5507 GND.n5506 585
R2005 GND.n5504 GND.n3311 585
R2006 GND.n3311 GND.n3308 585
R2007 GND.n5503 GND.n5502 585
R2008 GND.n5502 GND.n5501 585
R2009 GND.n3313 GND.n3312 585
R2010 GND.n5473 GND.n3313 585
R2011 GND.n5486 GND.n5485 585
R2012 GND.n5487 GND.n5486 585
R2013 GND.n5484 GND.n3325 585
R2014 GND.n5479 GND.n3325 585
R2015 GND.n5483 GND.n5482 585
R2016 GND.n5482 GND.n5481 585
R2017 GND.n3327 GND.n3326 585
R2018 GND.n5454 GND.n3327 585
R2019 GND.n5440 GND.n5439 585
R2020 GND.n5439 GND.n5438 585
R2021 GND.n5441 GND.n3343 585
R2022 GND.n5436 GND.n3343 585
R2023 GND.n5443 GND.n5442 585
R2024 GND.n5444 GND.n5443 585
R2025 GND.n3344 GND.n3342 585
R2026 GND.n5430 GND.n3342 585
R2027 GND.n5427 GND.n5426 585
R2028 GND.n5428 GND.n5427 585
R2029 GND.n5425 GND.n3348 585
R2030 GND.n5419 GND.n3348 585
R2031 GND.n5424 GND.n5423 585
R2032 GND.n5423 GND.n5422 585
R2033 GND.n3350 GND.n3349 585
R2034 GND.n5408 GND.n3350 585
R2035 GND.n5397 GND.n3368 585
R2036 GND.n3368 GND.n3360 585
R2037 GND.n5399 GND.n5398 585
R2038 GND.n5400 GND.n5399 585
R2039 GND.n5396 GND.n3367 585
R2040 GND.n5337 GND.n3367 585
R2041 GND.n5395 GND.n5394 585
R2042 GND.n5394 GND.n5393 585
R2043 GND.n3370 GND.n3369 585
R2044 GND.n5281 GND.n3370 585
R2045 GND.n5381 GND.n5380 585
R2046 GND.n5382 GND.n5381 585
R2047 GND.n5379 GND.n3383 585
R2048 GND.n3383 GND.n3379 585
R2049 GND.n5378 GND.n5377 585
R2050 GND.n5377 GND.n5376 585
R2051 GND.n3385 GND.n3384 585
R2052 GND.n5288 GND.n3385 585
R2053 GND.n5327 GND.n5326 585
R2054 GND.n5328 GND.n5327 585
R2055 GND.n5325 GND.n3397 585
R2056 GND.n3397 GND.n3394 585
R2057 GND.n5324 GND.n5323 585
R2058 GND.n5323 GND.n5322 585
R2059 GND.n3399 GND.n3398 585
R2060 GND.n5295 GND.n3399 585
R2061 GND.n5308 GND.n5307 585
R2062 GND.n5309 GND.n5308 585
R2063 GND.n5306 GND.n3411 585
R2064 GND.n5301 GND.n3411 585
R2065 GND.n5305 GND.n5304 585
R2066 GND.n5304 GND.n5303 585
R2067 GND.n3413 GND.n3412 585
R2068 GND.n5276 GND.n3413 585
R2069 GND.n5262 GND.n5261 585
R2070 GND.n5261 GND.n5260 585
R2071 GND.n5263 GND.n3428 585
R2072 GND.n5258 GND.n3428 585
R2073 GND.n5265 GND.n5264 585
R2074 GND.n5266 GND.n5265 585
R2075 GND.n3429 GND.n3427 585
R2076 GND.n5252 GND.n3427 585
R2077 GND.n5249 GND.n5248 585
R2078 GND.n5250 GND.n5249 585
R2079 GND.n5247 GND.n3435 585
R2080 GND.n5242 GND.n3435 585
R2081 GND.n5246 GND.n5245 585
R2082 GND.n5245 GND.n5244 585
R2083 GND.n3437 GND.n3436 585
R2084 GND.n5231 GND.n3437 585
R2085 GND.n5220 GND.n3455 585
R2086 GND.n3455 GND.n3447 585
R2087 GND.n5222 GND.n5221 585
R2088 GND.n5223 GND.n5222 585
R2089 GND.n5219 GND.n3454 585
R2090 GND.n3460 GND.n3454 585
R2091 GND.n5218 GND.n5217 585
R2092 GND.n5217 GND.n5216 585
R2093 GND.n3457 GND.n3456 585
R2094 GND.n5106 GND.n3457 585
R2095 GND.n5204 GND.n5203 585
R2096 GND.n5205 GND.n5204 585
R2097 GND.n5202 GND.n3472 585
R2098 GND.n3472 GND.n3468 585
R2099 GND.n5201 GND.n5200 585
R2100 GND.n5200 GND.n5199 585
R2101 GND.n3474 GND.n3473 585
R2102 GND.n5114 GND.n3474 585
R2103 GND.n5153 GND.n5152 585
R2104 GND.n5154 GND.n5153 585
R2105 GND.n5151 GND.n3486 585
R2106 GND.n3486 GND.n3483 585
R2107 GND.n5150 GND.n5149 585
R2108 GND.n5149 GND.n5148 585
R2109 GND.n3488 GND.n3487 585
R2110 GND.n5121 GND.n3488 585
R2111 GND.n5134 GND.n5133 585
R2112 GND.n5135 GND.n5134 585
R2113 GND.n5132 GND.n3501 585
R2114 GND.n5127 GND.n3501 585
R2115 GND.n5131 GND.n5130 585
R2116 GND.n5130 GND.n5129 585
R2117 GND.n3503 GND.n3502 585
R2118 GND.n5101 GND.n3503 585
R2119 GND.n5087 GND.n5086 585
R2120 GND.n5086 GND.n5085 585
R2121 GND.n5088 GND.n3519 585
R2122 GND.n5083 GND.n3519 585
R2123 GND.n5090 GND.n5089 585
R2124 GND.n5091 GND.n5090 585
R2125 GND.n3520 GND.n3518 585
R2126 GND.n5077 GND.n3518 585
R2127 GND.n5074 GND.n5073 585
R2128 GND.n5075 GND.n5074 585
R2129 GND.n5072 GND.n3524 585
R2130 GND.n5067 GND.n3524 585
R2131 GND.n5071 GND.n5070 585
R2132 GND.n5070 GND.n5069 585
R2133 GND.n3526 GND.n3525 585
R2134 GND.n5056 GND.n3526 585
R2135 GND.n5045 GND.n3545 585
R2136 GND.n3545 GND.n3536 585
R2137 GND.n5047 GND.n5046 585
R2138 GND.n5048 GND.n5047 585
R2139 GND.n5044 GND.n3544 585
R2140 GND.n3550 GND.n3544 585
R2141 GND.n5043 GND.n5042 585
R2142 GND.n5042 GND.n5041 585
R2143 GND.n3547 GND.n3546 585
R2144 GND.n4931 GND.n3547 585
R2145 GND.n5029 GND.n5028 585
R2146 GND.n5030 GND.n5029 585
R2147 GND.n5027 GND.n3561 585
R2148 GND.n3561 GND.n3557 585
R2149 GND.n5026 GND.n5025 585
R2150 GND.n5025 GND.n5024 585
R2151 GND.n3563 GND.n3562 585
R2152 GND.n4938 GND.n3563 585
R2153 GND.n4977 GND.n4976 585
R2154 GND.n4978 GND.n4977 585
R2155 GND.n4975 GND.n3575 585
R2156 GND.n3575 GND.n3572 585
R2157 GND.n4974 GND.n4973 585
R2158 GND.n4973 GND.n4972 585
R2159 GND.n3577 GND.n3576 585
R2160 GND.n4945 GND.n3577 585
R2161 GND.n4958 GND.n4957 585
R2162 GND.n4959 GND.n4958 585
R2163 GND.n4956 GND.n3590 585
R2164 GND.n4951 GND.n3590 585
R2165 GND.n4955 GND.n4954 585
R2166 GND.n4954 GND.n4953 585
R2167 GND.n3592 GND.n3591 585
R2168 GND.n4926 GND.n3592 585
R2169 GND.n4912 GND.n4911 585
R2170 GND.n4911 GND.n4910 585
R2171 GND.n4913 GND.n3608 585
R2172 GND.n4908 GND.n3608 585
R2173 GND.n4915 GND.n4914 585
R2174 GND.n4916 GND.n4915 585
R2175 GND.n3609 GND.n3607 585
R2176 GND.n4902 GND.n3607 585
R2177 GND.n4899 GND.n4898 585
R2178 GND.n4900 GND.n4899 585
R2179 GND.n4897 GND.n3613 585
R2180 GND.n4892 GND.n3613 585
R2181 GND.n4896 GND.n4895 585
R2182 GND.n4895 GND.n4894 585
R2183 GND.n3615 GND.n3614 585
R2184 GND.n4880 GND.n3615 585
R2185 GND.n4869 GND.n3633 585
R2186 GND.n3633 GND.n3625 585
R2187 GND.n4871 GND.n4870 585
R2188 GND.n4872 GND.n4871 585
R2189 GND.n4868 GND.n3632 585
R2190 GND.n3638 GND.n3632 585
R2191 GND.n4867 GND.n4866 585
R2192 GND.n4866 GND.n4865 585
R2193 GND.n3635 GND.n3634 585
R2194 GND.n4754 GND.n3635 585
R2195 GND.n4852 GND.n4851 585
R2196 GND.n4853 GND.n4852 585
R2197 GND.n4850 GND.n3649 585
R2198 GND.n3649 GND.n3645 585
R2199 GND.n4849 GND.n4848 585
R2200 GND.n4848 GND.n4847 585
R2201 GND.n3651 GND.n3650 585
R2202 GND.n4761 GND.n3651 585
R2203 GND.n4801 GND.n4800 585
R2204 GND.n4802 GND.n4801 585
R2205 GND.n4799 GND.n3663 585
R2206 GND.n3663 GND.n3660 585
R2207 GND.n4798 GND.n4797 585
R2208 GND.n4797 GND.n4796 585
R2209 GND.n3665 GND.n3664 585
R2210 GND.n4768 GND.n3665 585
R2211 GND.n4781 GND.n4780 585
R2212 GND.n4782 GND.n4781 585
R2213 GND.n4779 GND.n3677 585
R2214 GND.n4774 GND.n3677 585
R2215 GND.n4778 GND.n4777 585
R2216 GND.n4777 GND.n4776 585
R2217 GND.n3679 GND.n3678 585
R2218 GND.n4749 GND.n3679 585
R2219 GND.n4735 GND.n4734 585
R2220 GND.n4734 GND.n4733 585
R2221 GND.n4736 GND.n3695 585
R2222 GND.n4731 GND.n3695 585
R2223 GND.n4738 GND.n4737 585
R2224 GND.n4739 GND.n4738 585
R2225 GND.n3696 GND.n3694 585
R2226 GND.n4725 GND.n3694 585
R2227 GND.n4722 GND.n4721 585
R2228 GND.n4723 GND.n4722 585
R2229 GND.n4720 GND.n3700 585
R2230 GND.n4714 GND.n3700 585
R2231 GND.n4719 GND.n4718 585
R2232 GND.n4718 GND.n4717 585
R2233 GND.n3702 GND.n3701 585
R2234 GND.n4703 GND.n3702 585
R2235 GND.n4692 GND.n3720 585
R2236 GND.n3720 GND.n3712 585
R2237 GND.n4694 GND.n4693 585
R2238 GND.n4695 GND.n4694 585
R2239 GND.n4691 GND.n3719 585
R2240 GND.n3726 GND.n3719 585
R2241 GND.n4690 GND.n4689 585
R2242 GND.n4689 GND.n4688 585
R2243 GND.n3722 GND.n3721 585
R2244 GND.n4537 GND.n3722 585
R2245 GND.n4676 GND.n4675 585
R2246 GND.n4677 GND.n4676 585
R2247 GND.n4674 GND.n3737 585
R2248 GND.n3737 GND.n3733 585
R2249 GND.n4673 GND.n4672 585
R2250 GND.n4672 GND.n4671 585
R2251 GND.n3739 GND.n3738 585
R2252 GND.n4544 GND.n3739 585
R2253 GND.n4624 GND.n4623 585
R2254 GND.n4625 GND.n4624 585
R2255 GND.n4622 GND.n3751 585
R2256 GND.n3751 GND.n3748 585
R2257 GND.n4621 GND.n4620 585
R2258 GND.n4620 GND.n4619 585
R2259 GND.n3753 GND.n3752 585
R2260 GND.n4551 GND.n3753 585
R2261 GND.n4605 GND.n4604 585
R2262 GND.n4606 GND.n4605 585
R2263 GND.n4603 GND.n3764 585
R2264 GND.n4598 GND.n3764 585
R2265 GND.n4602 GND.n4601 585
R2266 GND.n4601 GND.n4600 585
R2267 GND.n3766 GND.n3765 585
R2268 GND.n3779 GND.n3766 585
R2269 GND.n4574 GND.n4573 585
R2270 GND.n4573 GND.n3778 585
R2271 GND.n4575 GND.n3789 585
R2272 GND.n4561 GND.n3789 585
R2273 GND.n4577 GND.n4576 585
R2274 GND.n4578 GND.n4577 585
R2275 GND.n4572 GND.n3788 585
R2276 GND.n4567 GND.n3788 585
R2277 GND.n4571 GND.n4570 585
R2278 GND.n4570 GND.n4569 585
R2279 GND.n3791 GND.n3790 585
R2280 GND.n4531 GND.n3791 585
R2281 GND.n4517 GND.n3809 585
R2282 GND.n3809 GND.n3808 585
R2283 GND.n4519 GND.n4518 585
R2284 GND.n4520 GND.n4519 585
R2285 GND.n4516 GND.n3807 585
R2286 GND.n3807 GND.n3803 585
R2287 GND.n4515 GND.n4514 585
R2288 GND.n4514 GND.n4513 585
R2289 GND.n3811 GND.n3810 585
R2290 GND.n4453 GND.n3811 585
R2291 GND.n4492 GND.n4491 585
R2292 GND.n4493 GND.n4492 585
R2293 GND.n4490 GND.n3823 585
R2294 GND.n3823 GND.n3820 585
R2295 GND.n4489 GND.n4488 585
R2296 GND.n4488 GND.n4487 585
R2297 GND.n3825 GND.n3824 585
R2298 GND.n4461 GND.n3825 585
R2299 GND.n4474 GND.n4473 585
R2300 GND.n4475 GND.n4474 585
R2301 GND.n4472 GND.n3838 585
R2302 GND.n3838 GND.n3835 585
R2303 GND.n4471 GND.n4470 585
R2304 GND.n4470 GND.n4469 585
R2305 GND.n3840 GND.n3839 585
R2306 GND.n4399 GND.n3840 585
R2307 GND.n4442 GND.n4441 585
R2308 GND.n4443 GND.n4442 585
R2309 GND.n4440 GND.n3848 585
R2310 GND.n4435 GND.n3848 585
R2311 GND.n4439 GND.n4438 585
R2312 GND.n4438 GND.n4437 585
R2313 GND.n3850 GND.n3849 585
R2314 GND.n4365 GND.n3850 585
R2315 GND.n4415 GND.n4414 585
R2316 GND.n4416 GND.n4415 585
R2317 GND.n4413 GND.n3863 585
R2318 GND.n3863 GND.n3860 585
R2319 GND.n4412 GND.n4411 585
R2320 GND.n4411 GND.n4410 585
R2321 GND.n3865 GND.n3864 585
R2322 GND.n4372 GND.n3865 585
R2323 GND.n4385 GND.n4384 585
R2324 GND.n4386 GND.n4385 585
R2325 GND.n4383 GND.n3878 585
R2326 GND.n4378 GND.n3878 585
R2327 GND.n4382 GND.n4381 585
R2328 GND.n4381 GND.n4380 585
R2329 GND.n3880 GND.n3879 585
R2330 GND.n4358 GND.n3880 585
R2331 GND.n4344 GND.n3895 585
R2332 GND.n3895 GND.n3894 585
R2333 GND.n4346 GND.n4345 585
R2334 GND.n4347 GND.n4346 585
R2335 GND.n4343 GND.n3893 585
R2336 GND.n3893 GND.n3889 585
R2337 GND.n4342 GND.n4341 585
R2338 GND.n4341 GND.n4340 585
R2339 GND.n3897 GND.n3896 585
R2340 GND.n3897 GND.n2664 585
R2341 GND.n4207 GND.n4206 585
R2342 GND.n4206 GND.n2662 585
R2343 GND.n4209 GND.n4208 585
R2344 GND.n4210 GND.n4209 585
R2345 GND.n2652 GND.n2651 585
R2346 GND.n2654 GND.n2652 585
R2347 GND.n6870 GND.n6869 585
R2348 GND.n6869 GND.n6868 585
R2349 GND.n6871 GND.n2649 585
R2350 GND.n4192 GND.n2649 585
R2351 GND.n6873 GND.n6872 585
R2352 GND.n6874 GND.n6873 585
R2353 GND.n2650 GND.n2648 585
R2354 GND.n2648 GND.n2645 585
R2355 GND.n4186 GND.n4185 585
R2356 GND.n4187 GND.n4186 585
R2357 GND.n2634 GND.n2633 585
R2358 GND.n2637 GND.n2634 585
R2359 GND.n6884 GND.n6883 585
R2360 GND.n6883 GND.n6882 585
R2361 GND.n6885 GND.n2631 585
R2362 GND.n2635 GND.n2631 585
R2363 GND.n6887 GND.n6886 585
R2364 GND.n6888 GND.n6887 585
R2365 GND.n2632 GND.n2630 585
R2366 GND.n2630 GND.n2627 585
R2367 GND.n4173 GND.n4172 585
R2368 GND.n4174 GND.n4173 585
R2369 GND.n2616 GND.n2615 585
R2370 GND.n2619 GND.n2616 585
R2371 GND.n6898 GND.n6897 585
R2372 GND.n6897 GND.n6896 585
R2373 GND.n6899 GND.n2613 585
R2374 GND.n2617 GND.n2613 585
R2375 GND.n6901 GND.n6900 585
R2376 GND.n6902 GND.n6901 585
R2377 GND.n2614 GND.n2612 585
R2378 GND.n2612 GND.n2609 585
R2379 GND.n4160 GND.n4159 585
R2380 GND.n4161 GND.n4160 585
R2381 GND.n2598 GND.n2597 585
R2382 GND.n2601 GND.n2598 585
R2383 GND.n6912 GND.n6911 585
R2384 GND.n6911 GND.n6910 585
R2385 GND.n6913 GND.n2595 585
R2386 GND.n2595 GND.n2593 585
R2387 GND.n6915 GND.n6914 585
R2388 GND.n6916 GND.n6915 585
R2389 GND.n2596 GND.n2594 585
R2390 GND.n2594 GND.n2591 585
R2391 GND.n4147 GND.n4146 585
R2392 GND.n4148 GND.n4147 585
R2393 GND.n2580 GND.n2579 585
R2394 GND.n2583 GND.n2580 585
R2395 GND.n6926 GND.n6925 585
R2396 GND.n6925 GND.n6924 585
R2397 GND.n6927 GND.n2577 585
R2398 GND.n4139 GND.n2577 585
R2399 GND.n6929 GND.n6928 585
R2400 GND.n6930 GND.n6929 585
R2401 GND.n2578 GND.n2576 585
R2402 GND.n2576 GND.n2574 585
R2403 GND.n4133 GND.n4132 585
R2404 GND.n4134 GND.n4133 585
R2405 GND.n2563 GND.n2562 585
R2406 GND.n2566 GND.n2563 585
R2407 GND.n6940 GND.n6939 585
R2408 GND.n6939 GND.n6938 585
R2409 GND.n6941 GND.n2560 585
R2410 GND.n2560 GND.n2558 585
R2411 GND.n6943 GND.n6942 585
R2412 GND.n6944 GND.n6943 585
R2413 GND.n2561 GND.n2559 585
R2414 GND.n2559 GND.n2556 585
R2415 GND.n4120 GND.n4119 585
R2416 GND.n4121 GND.n4120 585
R2417 GND.n2545 GND.n2544 585
R2418 GND.n2548 GND.n2545 585
R2419 GND.n6953 GND.n6952 585
R2420 GND.n6952 GND.n6951 585
R2421 GND.n6954 GND.n2542 585
R2422 GND.n4112 GND.n2542 585
R2423 GND.n6956 GND.n6955 585
R2424 GND.n6957 GND.n6956 585
R2425 GND.n2543 GND.n2541 585
R2426 GND.n2541 GND.n2539 585
R2427 GND.n3976 GND.n3975 585
R2428 GND.n3979 GND.n3978 585
R2429 GND.n3980 GND.n3960 585
R2430 GND.n3960 GND.n2530 585
R2431 GND.n3982 GND.n3981 585
R2432 GND.n3984 GND.n3959 585
R2433 GND.n3987 GND.n3986 585
R2434 GND.n3988 GND.n3958 585
R2435 GND.n3990 GND.n3989 585
R2436 GND.n3992 GND.n3957 585
R2437 GND.n3995 GND.n3994 585
R2438 GND.n3996 GND.n3956 585
R2439 GND.n3998 GND.n3997 585
R2440 GND.n4000 GND.n3955 585
R2441 GND.n4003 GND.n4002 585
R2442 GND.n4004 GND.n3954 585
R2443 GND.n4006 GND.n4005 585
R2444 GND.n4008 GND.n3953 585
R2445 GND.n4011 GND.n4010 585
R2446 GND.n4012 GND.n3952 585
R2447 GND.n4014 GND.n4013 585
R2448 GND.n4016 GND.n3951 585
R2449 GND.n4019 GND.n4018 585
R2450 GND.n4020 GND.n3950 585
R2451 GND.n4022 GND.n4021 585
R2452 GND.n4024 GND.n3949 585
R2453 GND.n4027 GND.n4026 585
R2454 GND.n4028 GND.n3948 585
R2455 GND.n4030 GND.n4029 585
R2456 GND.n4032 GND.n3947 585
R2457 GND.n4035 GND.n4034 585
R2458 GND.n4036 GND.n3943 585
R2459 GND.n4038 GND.n4037 585
R2460 GND.n4040 GND.n3942 585
R2461 GND.n4041 GND.n1407 585
R2462 GND.n4043 GND.n1407 585
R2463 GND.n4046 GND.n4045 585
R2464 GND.n4047 GND.n3941 585
R2465 GND.n4049 GND.n4048 585
R2466 GND.n4051 GND.n3940 585
R2467 GND.n4054 GND.n4053 585
R2468 GND.n4055 GND.n3936 585
R2469 GND.n4057 GND.n4056 585
R2470 GND.n4059 GND.n3935 585
R2471 GND.n4062 GND.n4061 585
R2472 GND.n4063 GND.n3934 585
R2473 GND.n4065 GND.n4064 585
R2474 GND.n4067 GND.n3933 585
R2475 GND.n4070 GND.n4069 585
R2476 GND.n4071 GND.n3932 585
R2477 GND.n4073 GND.n4072 585
R2478 GND.n4075 GND.n3931 585
R2479 GND.n4078 GND.n4077 585
R2480 GND.n4079 GND.n3930 585
R2481 GND.n4081 GND.n4080 585
R2482 GND.n4083 GND.n3929 585
R2483 GND.n4086 GND.n4085 585
R2484 GND.n4087 GND.n3928 585
R2485 GND.n4089 GND.n4088 585
R2486 GND.n4091 GND.n3927 585
R2487 GND.n4094 GND.n4093 585
R2488 GND.n4095 GND.n3926 585
R2489 GND.n4097 GND.n4096 585
R2490 GND.n4099 GND.n3925 585
R2491 GND.n4102 GND.n4101 585
R2492 GND.n4103 GND.n3924 585
R2493 GND.n4105 GND.n4104 585
R2494 GND.n4107 GND.n3923 585
R2495 GND.n4108 GND.n3922 585
R2496 GND.n4108 GND.n2530 585
R2497 GND.n5731 GND.n5730 585
R2498 GND.n5732 GND.n3210 585
R2499 GND.n5734 GND.n5733 585
R2500 GND.n5736 GND.n3208 585
R2501 GND.n5738 GND.n5737 585
R2502 GND.n5739 GND.n3207 585
R2503 GND.n5741 GND.n5740 585
R2504 GND.n5743 GND.n3205 585
R2505 GND.n5745 GND.n5744 585
R2506 GND.n5746 GND.n3204 585
R2507 GND.n5748 GND.n5747 585
R2508 GND.n5750 GND.n3202 585
R2509 GND.n5752 GND.n5751 585
R2510 GND.n5753 GND.n3201 585
R2511 GND.n5755 GND.n5754 585
R2512 GND.n5757 GND.n3199 585
R2513 GND.n5759 GND.n5758 585
R2514 GND.n5760 GND.n3198 585
R2515 GND.n5762 GND.n5761 585
R2516 GND.n5764 GND.n3196 585
R2517 GND.n5766 GND.n5765 585
R2518 GND.n5767 GND.n3195 585
R2519 GND.n5769 GND.n5768 585
R2520 GND.n5771 GND.n3193 585
R2521 GND.n5773 GND.n5772 585
R2522 GND.n5774 GND.n3192 585
R2523 GND.n5776 GND.n5775 585
R2524 GND.n5778 GND.n3190 585
R2525 GND.n5780 GND.n5779 585
R2526 GND.n5782 GND.n3187 585
R2527 GND.n5784 GND.n5783 585
R2528 GND.n5786 GND.n3186 585
R2529 GND.n5787 GND.n3086 585
R2530 GND.n3184 GND.n3087 585
R2531 GND.n3183 GND.n3182 585
R2532 GND.n3181 GND.n3180 585
R2533 GND.n3179 GND.n3089 585
R2534 GND.n3177 GND.n3176 585
R2535 GND.n3172 GND.n3090 585
R2536 GND.n3171 GND.n3170 585
R2537 GND.n3168 GND.n3091 585
R2538 GND.n3166 GND.n3165 585
R2539 GND.n3164 GND.n3092 585
R2540 GND.n3163 GND.n3162 585
R2541 GND.n3160 GND.n3093 585
R2542 GND.n3158 GND.n3157 585
R2543 GND.n3156 GND.n3094 585
R2544 GND.n3155 GND.n3154 585
R2545 GND.n3152 GND.n3095 585
R2546 GND.n3150 GND.n3149 585
R2547 GND.n3148 GND.n3096 585
R2548 GND.n3147 GND.n3146 585
R2549 GND.n3144 GND.n3097 585
R2550 GND.n3142 GND.n3141 585
R2551 GND.n3140 GND.n3098 585
R2552 GND.n3139 GND.n3138 585
R2553 GND.n3136 GND.n3099 585
R2554 GND.n3134 GND.n3133 585
R2555 GND.n3132 GND.n3100 585
R2556 GND.n3131 GND.n3130 585
R2557 GND.n3128 GND.n3101 585
R2558 GND.n3126 GND.n3125 585
R2559 GND.n3124 GND.n3102 585
R2560 GND.n3123 GND.n3122 585
R2561 GND.n3120 GND.n3103 585
R2562 GND.n3118 GND.n3117 585
R2563 GND.n5729 GND.n5725 585
R2564 GND.n5729 GND.n5728 585
R2565 GND.n5724 GND.n3029 585
R2566 GND.n6528 GND.n3029 585
R2567 GND.n5723 GND.n5722 585
R2568 GND.n5722 GND.n3028 585
R2569 GND.n5721 GND.n3021 585
R2570 GND.n6534 GND.n3021 585
R2571 GND.n5720 GND.n5719 585
R2572 GND.n5719 GND.n3020 585
R2573 GND.n5718 GND.n3211 585
R2574 GND.n5718 GND.n5717 585
R2575 GND.n5713 GND.n5712 585
R2576 GND.n5713 GND.n3012 585
R2577 GND.n5711 GND.n3011 585
R2578 GND.n6542 GND.n3011 585
R2579 GND.n5710 GND.n5709 585
R2580 GND.n5709 GND.n3010 585
R2581 GND.n5708 GND.n3003 585
R2582 GND.n6548 GND.n3003 585
R2583 GND.n5707 GND.n5706 585
R2584 GND.n5706 GND.n3002 585
R2585 GND.n5705 GND.n3212 585
R2586 GND.n5705 GND.n5704 585
R2587 GND.n5700 GND.n5699 585
R2588 GND.n5700 GND.n2994 585
R2589 GND.n5698 GND.n2993 585
R2590 GND.n6556 GND.n2993 585
R2591 GND.n5697 GND.n5696 585
R2592 GND.n5696 GND.n5695 585
R2593 GND.n5694 GND.n2986 585
R2594 GND.n6562 GND.n2986 585
R2595 GND.n5693 GND.n5692 585
R2596 GND.n5692 GND.n2985 585
R2597 GND.n5691 GND.n3213 585
R2598 GND.n5691 GND.n5690 585
R2599 GND.n5686 GND.n5685 585
R2600 GND.n5686 GND.n2977 585
R2601 GND.n5684 GND.n2976 585
R2602 GND.n6570 GND.n2976 585
R2603 GND.n5683 GND.n5682 585
R2604 GND.n5682 GND.n2975 585
R2605 GND.n5681 GND.n2968 585
R2606 GND.n6576 GND.n2968 585
R2607 GND.n5680 GND.n5679 585
R2608 GND.n5679 GND.n2967 585
R2609 GND.n5678 GND.n3214 585
R2610 GND.n5678 GND.n5677 585
R2611 GND.n5673 GND.n5672 585
R2612 GND.n5673 GND.n2959 585
R2613 GND.n5671 GND.n2958 585
R2614 GND.n6584 GND.n2958 585
R2615 GND.n5670 GND.n5669 585
R2616 GND.n5669 GND.n2951 585
R2617 GND.n5668 GND.n2950 585
R2618 GND.n6590 GND.n2950 585
R2619 GND.n5667 GND.n5666 585
R2620 GND.n5666 GND.n2949 585
R2621 GND.n5665 GND.n3215 585
R2622 GND.n5665 GND.n5664 585
R2623 GND.n5660 GND.n5659 585
R2624 GND.n5660 GND.n2941 585
R2625 GND.n5658 GND.n2940 585
R2626 GND.n6598 GND.n2940 585
R2627 GND.n5657 GND.n5656 585
R2628 GND.n5656 GND.n2933 585
R2629 GND.n5655 GND.n2932 585
R2630 GND.n6604 GND.n2932 585
R2631 GND.n5654 GND.n5653 585
R2632 GND.n5653 GND.n2931 585
R2633 GND.n5652 GND.n3216 585
R2634 GND.n5652 GND.n5651 585
R2635 GND.n5647 GND.n5646 585
R2636 GND.n5647 GND.n2923 585
R2637 GND.n5645 GND.n2922 585
R2638 GND.n6612 GND.n2922 585
R2639 GND.n5644 GND.n5643 585
R2640 GND.n5643 GND.n5642 585
R2641 GND.n5641 GND.n2915 585
R2642 GND.n6618 GND.n2915 585
R2643 GND.n5640 GND.n5639 585
R2644 GND.n5639 GND.n2914 585
R2645 GND.n5638 GND.n3217 585
R2646 GND.n5638 GND.n5637 585
R2647 GND.n5625 GND.n3218 585
R2648 GND.n3218 GND.n2905 585
R2649 GND.n5626 GND.n3241 585
R2650 GND.n3241 GND.n2904 585
R2651 GND.n5628 GND.n5627 585
R2652 GND.n5630 GND.n5628 585
R2653 GND.n5624 GND.n3240 585
R2654 GND.n5577 GND.n3240 585
R2655 GND.n5623 GND.n5622 585
R2656 GND.n5622 GND.n5621 585
R2657 GND.n3243 GND.n3242 585
R2658 GND.n5611 GND.n3243 585
R2659 GND.n3266 GND.n3250 585
R2660 GND.n5614 GND.n3250 585
R2661 GND.n5589 GND.n5588 585
R2662 GND.n5588 GND.n5587 585
R2663 GND.n5590 GND.n3259 585
R2664 GND.n5601 GND.n3259 585
R2665 GND.n5592 GND.n5591 585
R2666 GND.n5593 GND.n5592 585
R2667 GND.n3265 GND.n3264 585
R2668 GND.n5595 GND.n3264 585
R2669 GND.n5561 GND.n5560 585
R2670 GND.n5562 GND.n5561 585
R2671 GND.n5559 GND.n3275 585
R2672 GND.n3275 GND.n3273 585
R2673 GND.n5558 GND.n5557 585
R2674 GND.n5557 GND.n5556 585
R2675 GND.n3277 GND.n3276 585
R2676 GND.n3286 GND.n3277 585
R2677 GND.n5458 GND.n3285 585
R2678 GND.n5549 GND.n3285 585
R2679 GND.n5461 GND.n5460 585
R2680 GND.n5460 GND.n5459 585
R2681 GND.n5462 GND.n3295 585
R2682 GND.n5535 GND.n3295 585
R2683 GND.n5464 GND.n5463 585
R2684 GND.n5463 GND.n3293 585
R2685 GND.n5465 GND.n3301 585
R2686 GND.n5529 GND.n3301 585
R2687 GND.n5468 GND.n5467 585
R2688 GND.n5467 GND.n5466 585
R2689 GND.n5469 GND.n3309 585
R2690 GND.n5507 GND.n3309 585
R2691 GND.n5471 GND.n5470 585
R2692 GND.n5470 GND.n3308 585
R2693 GND.n5472 GND.n3315 585
R2694 GND.n5501 GND.n3315 585
R2695 GND.n5475 GND.n5474 585
R2696 GND.n5474 GND.n5473 585
R2697 GND.n5476 GND.n3323 585
R2698 GND.n5487 GND.n3323 585
R2699 GND.n5478 GND.n5477 585
R2700 GND.n5479 GND.n5478 585
R2701 GND.n5457 GND.n3329 585
R2702 GND.n5481 GND.n3329 585
R2703 GND.n5456 GND.n5455 585
R2704 GND.n5455 GND.n5454 585
R2705 GND.n3331 GND.n3330 585
R2706 GND.n5438 GND.n3331 585
R2707 GND.n5435 GND.n5434 585
R2708 GND.n5436 GND.n5435 585
R2709 GND.n5433 GND.n3340 585
R2710 GND.n5444 GND.n3340 585
R2711 GND.n5432 GND.n5431 585
R2712 GND.n5431 GND.n5430 585
R2713 GND.n3346 GND.n3345 585
R2714 GND.n5428 GND.n3346 585
R2715 GND.n5404 GND.n3354 585
R2716 GND.n5419 GND.n3354 585
R2717 GND.n5405 GND.n3352 585
R2718 GND.n5422 GND.n3352 585
R2719 GND.n5407 GND.n5406 585
R2720 GND.n5408 GND.n5407 585
R2721 GND.n5403 GND.n3362 585
R2722 GND.n3362 GND.n3360 585
R2723 GND.n5402 GND.n5401 585
R2724 GND.n5401 GND.n5400 585
R2725 GND.n3364 GND.n3363 585
R2726 GND.n5337 GND.n3364 585
R2727 GND.n5280 GND.n3373 585
R2728 GND.n5393 GND.n3373 585
R2729 GND.n5283 GND.n5282 585
R2730 GND.n5282 GND.n5281 585
R2731 GND.n5284 GND.n3381 585
R2732 GND.n5382 GND.n3381 585
R2733 GND.n5286 GND.n5285 585
R2734 GND.n5285 GND.n3379 585
R2735 GND.n5287 GND.n3387 585
R2736 GND.n5376 GND.n3387 585
R2737 GND.n5290 GND.n5289 585
R2738 GND.n5289 GND.n5288 585
R2739 GND.n5291 GND.n3395 585
R2740 GND.n5328 GND.n3395 585
R2741 GND.n5293 GND.n5292 585
R2742 GND.n5292 GND.n3394 585
R2743 GND.n5294 GND.n3401 585
R2744 GND.n5322 GND.n3401 585
R2745 GND.n5297 GND.n5296 585
R2746 GND.n5296 GND.n5295 585
R2747 GND.n5298 GND.n3409 585
R2748 GND.n5309 GND.n3409 585
R2749 GND.n5300 GND.n5299 585
R2750 GND.n5301 GND.n5300 585
R2751 GND.n5279 GND.n3416 585
R2752 GND.n5303 GND.n3416 585
R2753 GND.n5278 GND.n5277 585
R2754 GND.n5277 GND.n5276 585
R2755 GND.n3418 GND.n3417 585
R2756 GND.n5260 GND.n3418 585
R2757 GND.n5257 GND.n5256 585
R2758 GND.n5258 GND.n5257 585
R2759 GND.n5255 GND.n3426 585
R2760 GND.n5266 GND.n3426 585
R2761 GND.n5254 GND.n5253 585
R2762 GND.n5253 GND.n5252 585
R2763 GND.n3432 GND.n3431 585
R2764 GND.n5250 GND.n3432 585
R2765 GND.n5227 GND.n3441 585
R2766 GND.n5242 GND.n3441 585
R2767 GND.n5228 GND.n3439 585
R2768 GND.n5244 GND.n3439 585
R2769 GND.n5230 GND.n5229 585
R2770 GND.n5231 GND.n5230 585
R2771 GND.n5226 GND.n3449 585
R2772 GND.n3449 GND.n3447 585
R2773 GND.n5225 GND.n5224 585
R2774 GND.n5224 GND.n5223 585
R2775 GND.n3451 GND.n3450 585
R2776 GND.n3460 GND.n3451 585
R2777 GND.n5105 GND.n3459 585
R2778 GND.n5216 GND.n3459 585
R2779 GND.n5108 GND.n5107 585
R2780 GND.n5107 GND.n5106 585
R2781 GND.n5109 GND.n3470 585
R2782 GND.n5205 GND.n3470 585
R2783 GND.n5111 GND.n5110 585
R2784 GND.n5110 GND.n3468 585
R2785 GND.n5112 GND.n3476 585
R2786 GND.n5199 GND.n3476 585
R2787 GND.n5116 GND.n5115 585
R2788 GND.n5115 GND.n5114 585
R2789 GND.n5117 GND.n3484 585
R2790 GND.n5154 GND.n3484 585
R2791 GND.n5119 GND.n5118 585
R2792 GND.n5118 GND.n3483 585
R2793 GND.n5120 GND.n3490 585
R2794 GND.n5148 GND.n3490 585
R2795 GND.n5123 GND.n5122 585
R2796 GND.n5122 GND.n5121 585
R2797 GND.n5124 GND.n3499 585
R2798 GND.n5135 GND.n3499 585
R2799 GND.n5126 GND.n5125 585
R2800 GND.n5127 GND.n5126 585
R2801 GND.n5104 GND.n3505 585
R2802 GND.n5129 GND.n3505 585
R2803 GND.n5103 GND.n5102 585
R2804 GND.n5102 GND.n5101 585
R2805 GND.n3507 GND.n3506 585
R2806 GND.n5085 GND.n3507 585
R2807 GND.n5082 GND.n5081 585
R2808 GND.n5083 GND.n5082 585
R2809 GND.n5080 GND.n3516 585
R2810 GND.n5091 GND.n3516 585
R2811 GND.n5079 GND.n5078 585
R2812 GND.n5078 GND.n5077 585
R2813 GND.n3522 GND.n3521 585
R2814 GND.n5075 GND.n3522 585
R2815 GND.n5052 GND.n3530 585
R2816 GND.n5067 GND.n3530 585
R2817 GND.n5053 GND.n3528 585
R2818 GND.n5069 GND.n3528 585
R2819 GND.n5055 GND.n5054 585
R2820 GND.n5056 GND.n5055 585
R2821 GND.n5051 GND.n3538 585
R2822 GND.n3538 GND.n3536 585
R2823 GND.n5050 GND.n5049 585
R2824 GND.n5049 GND.n5048 585
R2825 GND.n3540 GND.n3539 585
R2826 GND.n3550 GND.n3540 585
R2827 GND.n4930 GND.n3549 585
R2828 GND.n5041 GND.n3549 585
R2829 GND.n4933 GND.n4932 585
R2830 GND.n4932 GND.n4931 585
R2831 GND.n4934 GND.n3559 585
R2832 GND.n5030 GND.n3559 585
R2833 GND.n4936 GND.n4935 585
R2834 GND.n4935 GND.n3557 585
R2835 GND.n4937 GND.n3565 585
R2836 GND.n5024 GND.n3565 585
R2837 GND.n4940 GND.n4939 585
R2838 GND.n4939 GND.n4938 585
R2839 GND.n4941 GND.n3573 585
R2840 GND.n4978 GND.n3573 585
R2841 GND.n4943 GND.n4942 585
R2842 GND.n4942 GND.n3572 585
R2843 GND.n4944 GND.n3579 585
R2844 GND.n4972 GND.n3579 585
R2845 GND.n4947 GND.n4946 585
R2846 GND.n4946 GND.n4945 585
R2847 GND.n4948 GND.n3587 585
R2848 GND.n4959 GND.n3587 585
R2849 GND.n4950 GND.n4949 585
R2850 GND.n4951 GND.n4950 585
R2851 GND.n4929 GND.n3594 585
R2852 GND.n4953 GND.n3594 585
R2853 GND.n4928 GND.n4927 585
R2854 GND.n4927 GND.n4926 585
R2855 GND.n3596 GND.n3595 585
R2856 GND.n4910 GND.n3596 585
R2857 GND.n4907 GND.n4906 585
R2858 GND.n4908 GND.n4907 585
R2859 GND.n4905 GND.n3604 585
R2860 GND.n4916 GND.n3604 585
R2861 GND.n4904 GND.n4903 585
R2862 GND.n4903 GND.n4902 585
R2863 GND.n3611 GND.n3610 585
R2864 GND.n4900 GND.n3611 585
R2865 GND.n4876 GND.n3619 585
R2866 GND.n4892 GND.n3619 585
R2867 GND.n4877 GND.n3617 585
R2868 GND.n4894 GND.n3617 585
R2869 GND.n4879 GND.n4878 585
R2870 GND.n4880 GND.n4879 585
R2871 GND.n4875 GND.n3627 585
R2872 GND.n3627 GND.n3625 585
R2873 GND.n4874 GND.n4873 585
R2874 GND.n4873 GND.n4872 585
R2875 GND.n3629 GND.n3628 585
R2876 GND.n3638 GND.n3629 585
R2877 GND.n4753 GND.n3637 585
R2878 GND.n4865 GND.n3637 585
R2879 GND.n4756 GND.n4755 585
R2880 GND.n4755 GND.n4754 585
R2881 GND.n4757 GND.n3647 585
R2882 GND.n4853 GND.n3647 585
R2883 GND.n4759 GND.n4758 585
R2884 GND.n4758 GND.n3645 585
R2885 GND.n4760 GND.n3653 585
R2886 GND.n4847 GND.n3653 585
R2887 GND.n4763 GND.n4762 585
R2888 GND.n4762 GND.n4761 585
R2889 GND.n4764 GND.n3661 585
R2890 GND.n4802 GND.n3661 585
R2891 GND.n4766 GND.n4765 585
R2892 GND.n4765 GND.n3660 585
R2893 GND.n4767 GND.n3667 585
R2894 GND.n4796 GND.n3667 585
R2895 GND.n4770 GND.n4769 585
R2896 GND.n4769 GND.n4768 585
R2897 GND.n4771 GND.n3675 585
R2898 GND.n4782 GND.n3675 585
R2899 GND.n4773 GND.n4772 585
R2900 GND.n4774 GND.n4773 585
R2901 GND.n4752 GND.n3681 585
R2902 GND.n4776 GND.n3681 585
R2903 GND.n4751 GND.n4750 585
R2904 GND.n4750 GND.n4749 585
R2905 GND.n3683 GND.n3682 585
R2906 GND.n4733 GND.n3683 585
R2907 GND.n4730 GND.n4729 585
R2908 GND.n4731 GND.n4730 585
R2909 GND.n4728 GND.n3692 585
R2910 GND.n4739 GND.n3692 585
R2911 GND.n4727 GND.n4726 585
R2912 GND.n4726 GND.n4725 585
R2913 GND.n3698 GND.n3697 585
R2914 GND.n4723 GND.n3698 585
R2915 GND.n4699 GND.n3706 585
R2916 GND.n4714 GND.n3706 585
R2917 GND.n4700 GND.n3704 585
R2918 GND.n4717 GND.n3704 585
R2919 GND.n4702 GND.n4701 585
R2920 GND.n4703 GND.n4702 585
R2921 GND.n4698 GND.n3714 585
R2922 GND.n3714 GND.n3712 585
R2923 GND.n4697 GND.n4696 585
R2924 GND.n4696 GND.n4695 585
R2925 GND.n3716 GND.n3715 585
R2926 GND.n3726 GND.n3716 585
R2927 GND.n4536 GND.n3725 585
R2928 GND.n4688 GND.n3725 585
R2929 GND.n4539 GND.n4538 585
R2930 GND.n4538 GND.n4537 585
R2931 GND.n4540 GND.n3735 585
R2932 GND.n4677 GND.n3735 585
R2933 GND.n4542 GND.n4541 585
R2934 GND.n4541 GND.n3733 585
R2935 GND.n4543 GND.n3741 585
R2936 GND.n4671 GND.n3741 585
R2937 GND.n4546 GND.n4545 585
R2938 GND.n4545 GND.n4544 585
R2939 GND.n4547 GND.n3749 585
R2940 GND.n4625 GND.n3749 585
R2941 GND.n4549 GND.n4548 585
R2942 GND.n4548 GND.n3748 585
R2943 GND.n4550 GND.n3755 585
R2944 GND.n4619 GND.n3755 585
R2945 GND.n4553 GND.n4552 585
R2946 GND.n4552 GND.n4551 585
R2947 GND.n4554 GND.n3762 585
R2948 GND.n4606 GND.n3762 585
R2949 GND.n4555 GND.n3770 585
R2950 GND.n4598 GND.n3770 585
R2951 GND.n4556 GND.n3769 585
R2952 GND.n4600 GND.n3769 585
R2953 GND.n4558 GND.n4557 585
R2954 GND.n4558 GND.n3779 585
R2955 GND.n4559 GND.n4535 585
R2956 GND.n4559 GND.n3778 585
R2957 GND.n4563 GND.n4562 585
R2958 GND.n4562 GND.n4561 585
R2959 GND.n4564 GND.n3786 585
R2960 GND.n4578 GND.n3786 585
R2961 GND.n4566 GND.n4565 585
R2962 GND.n4567 GND.n4566 585
R2963 GND.n4534 GND.n3794 585
R2964 GND.n4569 GND.n3794 585
R2965 GND.n4533 GND.n4532 585
R2966 GND.n4532 GND.n4531 585
R2967 GND.n3796 GND.n3795 585
R2968 GND.n3808 GND.n3796 585
R2969 GND.n4447 GND.n3805 585
R2970 GND.n4520 GND.n3805 585
R2971 GND.n4449 GND.n4448 585
R2972 GND.n4448 GND.n3803 585
R2973 GND.n4450 GND.n3813 585
R2974 GND.n4513 GND.n3813 585
R2975 GND.n4455 GND.n4454 585
R2976 GND.n4454 GND.n4453 585
R2977 GND.n4456 GND.n3821 585
R2978 GND.n4493 GND.n3821 585
R2979 GND.n4458 GND.n4457 585
R2980 GND.n4457 GND.n3820 585
R2981 GND.n4459 GND.n3827 585
R2982 GND.n4487 GND.n3827 585
R2983 GND.n4463 GND.n4462 585
R2984 GND.n4462 GND.n4461 585
R2985 GND.n4464 GND.n3836 585
R2986 GND.n4475 GND.n3836 585
R2987 GND.n4465 GND.n3843 585
R2988 GND.n3843 GND.n3835 585
R2989 GND.n4467 GND.n4466 585
R2990 GND.n4469 GND.n4467 585
R2991 GND.n4446 GND.n3842 585
R2992 GND.n4399 GND.n3842 585
R2993 GND.n4445 GND.n4444 585
R2994 GND.n4444 GND.n4443 585
R2995 GND.n3845 GND.n3844 585
R2996 GND.n4435 GND.n3845 585
R2997 GND.n4362 GND.n3852 585
R2998 GND.n4437 GND.n3852 585
R2999 GND.n4367 GND.n4366 585
R3000 GND.n4366 GND.n4365 585
R3001 GND.n4368 GND.n3861 585
R3002 GND.n4416 GND.n3861 585
R3003 GND.n4370 GND.n4369 585
R3004 GND.n4369 GND.n3860 585
R3005 GND.n4371 GND.n3867 585
R3006 GND.n4410 GND.n3867 585
R3007 GND.n4374 GND.n4373 585
R3008 GND.n4373 GND.n4372 585
R3009 GND.n4375 GND.n3876 585
R3010 GND.n4386 GND.n3876 585
R3011 GND.n4377 GND.n4376 585
R3012 GND.n4378 GND.n4377 585
R3013 GND.n4361 GND.n3882 585
R3014 GND.n4380 GND.n3882 585
R3015 GND.n4360 GND.n4359 585
R3016 GND.n4359 GND.n4358 585
R3017 GND.n3884 GND.n3883 585
R3018 GND.n3894 GND.n3884 585
R3019 GND.n4197 GND.n3891 585
R3020 GND.n4347 GND.n3891 585
R3021 GND.n4199 GND.n4198 585
R3022 GND.n4198 GND.n3889 585
R3023 GND.n4200 GND.n3899 585
R3024 GND.n4340 GND.n3899 585
R3025 GND.n4202 GND.n4201 585
R3026 GND.n4201 GND.n2664 585
R3027 GND.n4203 GND.n3915 585
R3028 GND.n3915 GND.n2662 585
R3029 GND.n4205 GND.n4204 585
R3030 GND.n4210 GND.n4205 585
R3031 GND.n4196 GND.n3914 585
R3032 GND.n3914 GND.n2654 585
R3033 GND.n4195 GND.n2653 585
R3034 GND.n6868 GND.n2653 585
R3035 GND.n4194 GND.n4193 585
R3036 GND.n4193 GND.n4192 585
R3037 GND.n4191 GND.n2646 585
R3038 GND.n6874 GND.n2646 585
R3039 GND.n4190 GND.n4189 585
R3040 GND.n4189 GND.n2645 585
R3041 GND.n4188 GND.n3916 585
R3042 GND.n4188 GND.n4187 585
R3043 GND.n4183 GND.n4182 585
R3044 GND.n4183 GND.n2637 585
R3045 GND.n4181 GND.n2636 585
R3046 GND.n6882 GND.n2636 585
R3047 GND.n4180 GND.n4179 585
R3048 GND.n4179 GND.n2635 585
R3049 GND.n4178 GND.n2628 585
R3050 GND.n6888 GND.n2628 585
R3051 GND.n4177 GND.n4176 585
R3052 GND.n4176 GND.n2627 585
R3053 GND.n4175 GND.n3917 585
R3054 GND.n4175 GND.n4174 585
R3055 GND.n4170 GND.n4169 585
R3056 GND.n4170 GND.n2619 585
R3057 GND.n4168 GND.n2618 585
R3058 GND.n6896 GND.n2618 585
R3059 GND.n4167 GND.n4166 585
R3060 GND.n4166 GND.n2617 585
R3061 GND.n4165 GND.n2610 585
R3062 GND.n6902 GND.n2610 585
R3063 GND.n4164 GND.n4163 585
R3064 GND.n4163 GND.n2609 585
R3065 GND.n4162 GND.n3918 585
R3066 GND.n4162 GND.n4161 585
R3067 GND.n4157 GND.n4156 585
R3068 GND.n4157 GND.n2601 585
R3069 GND.n4155 GND.n2600 585
R3070 GND.n6910 GND.n2600 585
R3071 GND.n4154 GND.n4153 585
R3072 GND.n4153 GND.n2593 585
R3073 GND.n4152 GND.n2592 585
R3074 GND.n6916 GND.n2592 585
R3075 GND.n4151 GND.n4150 585
R3076 GND.n4150 GND.n2591 585
R3077 GND.n4149 GND.n3919 585
R3078 GND.n4149 GND.n4148 585
R3079 GND.n4144 GND.n4143 585
R3080 GND.n4144 GND.n2583 585
R3081 GND.n4142 GND.n2582 585
R3082 GND.n6924 GND.n2582 585
R3083 GND.n4141 GND.n4140 585
R3084 GND.n4140 GND.n4139 585
R3085 GND.n4138 GND.n2575 585
R3086 GND.n6930 GND.n2575 585
R3087 GND.n4137 GND.n4136 585
R3088 GND.n4136 GND.n2574 585
R3089 GND.n4135 GND.n3920 585
R3090 GND.n4135 GND.n4134 585
R3091 GND.n4130 GND.n4129 585
R3092 GND.n4130 GND.n2566 585
R3093 GND.n4128 GND.n2565 585
R3094 GND.n6938 GND.n2565 585
R3095 GND.n4127 GND.n4126 585
R3096 GND.n4126 GND.n2558 585
R3097 GND.n4125 GND.n2557 585
R3098 GND.n6944 GND.n2557 585
R3099 GND.n4124 GND.n4123 585
R3100 GND.n4123 GND.n2556 585
R3101 GND.n4122 GND.n3921 585
R3102 GND.n4122 GND.n4121 585
R3103 GND.n4117 GND.n4116 585
R3104 GND.n4117 GND.n2548 585
R3105 GND.n4115 GND.n2547 585
R3106 GND.n6951 GND.n2547 585
R3107 GND.n4114 GND.n4113 585
R3108 GND.n4113 GND.n4112 585
R3109 GND.n4111 GND.n2540 585
R3110 GND.n6957 GND.n2540 585
R3111 GND.n4110 GND.n4109 585
R3112 GND.n4109 GND.n2539 585
R3113 GND.n423 GND.n422 585
R3114 GND.n8398 GND.n423 585
R3115 GND.n8401 GND.n8400 585
R3116 GND.n8400 GND.n8399 585
R3117 GND.n8402 GND.n417 585
R3118 GND.n417 GND.n416 585
R3119 GND.n8404 GND.n8403 585
R3120 GND.n8405 GND.n8404 585
R3121 GND.n415 GND.n414 585
R3122 GND.n8406 GND.n415 585
R3123 GND.n8409 GND.n8408 585
R3124 GND.n8408 GND.n8407 585
R3125 GND.n8410 GND.n409 585
R3126 GND.n409 GND.n408 585
R3127 GND.n8412 GND.n8411 585
R3128 GND.n8413 GND.n8412 585
R3129 GND.n407 GND.n406 585
R3130 GND.n8414 GND.n407 585
R3131 GND.n8417 GND.n8416 585
R3132 GND.n8416 GND.n8415 585
R3133 GND.n8418 GND.n401 585
R3134 GND.n401 GND.n400 585
R3135 GND.n8420 GND.n8419 585
R3136 GND.n8421 GND.n8420 585
R3137 GND.n399 GND.n398 585
R3138 GND.n8422 GND.n399 585
R3139 GND.n8425 GND.n8424 585
R3140 GND.n8424 GND.n8423 585
R3141 GND.n8426 GND.n393 585
R3142 GND.n393 GND.n392 585
R3143 GND.n8428 GND.n8427 585
R3144 GND.n8429 GND.n8428 585
R3145 GND.n391 GND.n390 585
R3146 GND.n8430 GND.n391 585
R3147 GND.n8433 GND.n8432 585
R3148 GND.n8432 GND.n8431 585
R3149 GND.n8434 GND.n385 585
R3150 GND.n385 GND.n384 585
R3151 GND.n8436 GND.n8435 585
R3152 GND.n8437 GND.n8436 585
R3153 GND.n261 GND.n260 585
R3154 GND.n8438 GND.n261 585
R3155 GND.n8441 GND.n8440 585
R3156 GND.n8440 GND.n8439 585
R3157 GND.n8442 GND.n255 585
R3158 GND.n255 GND.n253 585
R3159 GND.n8444 GND.n8443 585
R3160 GND.n8445 GND.n8444 585
R3161 GND.n256 GND.n254 585
R3162 GND.n254 GND.n246 585
R3163 GND.n6330 GND.n6329 585
R3164 GND.n6329 GND.n243 585
R3165 GND.n6331 GND.n6309 585
R3166 GND.n6309 GND.n235 585
R3167 GND.n6333 GND.n6332 585
R3168 GND.n6334 GND.n6333 585
R3169 GND.n6310 GND.n6308 585
R3170 GND.n6308 GND.n226 585
R3171 GND.n6322 GND.n6321 585
R3172 GND.n6321 GND.n223 585
R3173 GND.n6320 GND.n6312 585
R3174 GND.n6320 GND.n215 585
R3175 GND.n6319 GND.n6318 585
R3176 GND.n6319 GND.n212 585
R3177 GND.n6314 GND.n6313 585
R3178 GND.n6313 GND.n205 585
R3179 GND.n5958 GND.n5957 585
R3180 GND.n5958 GND.n202 585
R3181 GND.n6356 GND.n6355 585
R3182 GND.n6355 GND.n6354 585
R3183 GND.n6357 GND.n5952 585
R3184 GND.n5952 GND.n192 585
R3185 GND.n6359 GND.n6358 585
R3186 GND.n6359 GND.n185 585
R3187 GND.n6360 GND.n5951 585
R3188 GND.n6360 GND.n182 585
R3189 GND.n6362 GND.n6361 585
R3190 GND.n6361 GND.n175 585
R3191 GND.n6363 GND.n5948 585
R3192 GND.n5948 GND.n172 585
R3193 GND.n6365 GND.n6364 585
R3194 GND.n6365 GND.n163 585
R3195 GND.n6367 GND.n6366 585
R3196 GND.n6366 GND.n160 585
R3197 GND.n6368 GND.n5945 585
R3198 GND.n5974 GND.n5945 585
R3199 GND.n6371 GND.n6370 585
R3200 GND.n6372 GND.n6371 585
R3201 GND.n5946 GND.n5931 585
R3202 GND.n5931 GND.n143 585
R3203 GND.n6382 GND.n6381 585
R3204 GND.n6381 GND.n6380 585
R3205 GND.n6383 GND.n5928 585
R3206 GND.n5932 GND.n5928 585
R3207 GND.n6386 GND.n6385 585
R3208 GND.n6387 GND.n6386 585
R3209 GND.n5929 GND.n5927 585
R3210 GND.n5927 GND.n5921 585
R3211 GND.n6032 GND.n5978 585
R3212 GND.n5978 GND.n5918 585
R3213 GND.n6034 GND.n6033 585
R3214 GND.n6035 GND.n6034 585
R3215 GND.n5979 GND.n5977 585
R3216 GND.n5977 GND.n5909 585
R3217 GND.n6027 GND.n6026 585
R3218 GND.n6026 GND.n5902 585
R3219 GND.n6025 GND.n5981 585
R3220 GND.n6025 GND.n5899 585
R3221 GND.n6024 GND.n6023 585
R3222 GND.n6024 GND.n5892 585
R3223 GND.n5983 GND.n5982 585
R3224 GND.n5982 GND.n5889 585
R3225 GND.n6019 GND.n6018 585
R3226 GND.n6018 GND.n5881 585
R3227 GND.n6017 GND.n5985 585
R3228 GND.n6017 GND.n5878 585
R3229 GND.n6016 GND.n6015 585
R3230 GND.n6016 GND.n5871 585
R3231 GND.n5987 GND.n5986 585
R3232 GND.n5986 GND.n5868 585
R3233 GND.n6011 GND.n6010 585
R3234 GND.n6010 GND.n5860 585
R3235 GND.n6009 GND.n5989 585
R3236 GND.n6009 GND.n5857 585
R3237 GND.n6008 GND.n6007 585
R3238 GND.n6008 GND.n5847 585
R3239 GND.n5991 GND.n5990 585
R3240 GND.n5990 GND.n5844 585
R3241 GND.n6003 GND.n6002 585
R3242 GND.n6002 GND.n5831 585
R3243 GND.n6001 GND.n5993 585
R3244 GND.n6001 GND.n5829 585
R3245 GND.n6000 GND.n5999 585
R3246 GND.n6000 GND.n5821 585
R3247 GND.n5995 GND.n5994 585
R3248 GND.n5994 GND.n5819 585
R3249 GND.n3045 GND.n3044 585
R3250 GND.n3067 GND.n3045 585
R3251 GND.n6515 GND.n6514 585
R3252 GND.n6514 GND.n6513 585
R3253 GND.n6516 GND.n3039 585
R3254 GND.n3039 GND.n3038 585
R3255 GND.n6518 GND.n6517 585
R3256 GND.n6519 GND.n6518 585
R3257 GND.n3036 GND.n3035 585
R3258 GND.n6520 GND.n3036 585
R3259 GND.n6523 GND.n6522 585
R3260 GND.n6522 GND.n6521 585
R3261 GND.n6524 GND.n3030 585
R3262 GND.n5727 GND.n3030 585
R3263 GND.n6526 GND.n6525 585
R3264 GND.n6527 GND.n6526 585
R3265 GND.n3019 GND.n3018 585
R3266 GND.n3027 GND.n3019 585
R3267 GND.n6537 GND.n6536 585
R3268 GND.n6536 GND.n6535 585
R3269 GND.n6538 GND.n3013 585
R3270 GND.n5714 GND.n3013 585
R3271 GND.n6540 GND.n6539 585
R3272 GND.n6541 GND.n6540 585
R3273 GND.n3001 GND.n3000 585
R3274 GND.n3004 GND.n3001 585
R3275 GND.n6551 GND.n6550 585
R3276 GND.n6550 GND.n6549 585
R3277 GND.n6552 GND.n2995 585
R3278 GND.n5701 GND.n2995 585
R3279 GND.n6554 GND.n6553 585
R3280 GND.n6555 GND.n6554 585
R3281 GND.n2984 GND.n2983 585
R3282 GND.n2987 GND.n2984 585
R3283 GND.n6565 GND.n6564 585
R3284 GND.n6564 GND.n6563 585
R3285 GND.n6566 GND.n2978 585
R3286 GND.n5687 GND.n2978 585
R3287 GND.n6568 GND.n6567 585
R3288 GND.n6569 GND.n6568 585
R3289 GND.n2966 GND.n2965 585
R3290 GND.n2969 GND.n2966 585
R3291 GND.n6579 GND.n6578 585
R3292 GND.n6578 GND.n6577 585
R3293 GND.n6580 GND.n2960 585
R3294 GND.n5674 GND.n2960 585
R3295 GND.n6582 GND.n6581 585
R3296 GND.n6583 GND.n6582 585
R3297 GND.n2948 GND.n2947 585
R3298 GND.n2957 GND.n2948 585
R3299 GND.n6593 GND.n6592 585
R3300 GND.n6592 GND.n6591 585
R3301 GND.n6594 GND.n2942 585
R3302 GND.n5661 GND.n2942 585
R3303 GND.n6596 GND.n6595 585
R3304 GND.n6597 GND.n6596 585
R3305 GND.n2930 GND.n2929 585
R3306 GND.n2939 GND.n2930 585
R3307 GND.n6607 GND.n6606 585
R3308 GND.n6606 GND.n6605 585
R3309 GND.n6608 GND.n2924 585
R3310 GND.n5648 GND.n2924 585
R3311 GND.n6610 GND.n6609 585
R3312 GND.n6611 GND.n6610 585
R3313 GND.n2913 GND.n2912 585
R3314 GND.n2921 GND.n2913 585
R3315 GND.n6621 GND.n6620 585
R3316 GND.n6620 GND.n6619 585
R3317 GND.n6622 GND.n2907 585
R3318 GND.n3235 GND.n2907 585
R3319 GND.n6624 GND.n6623 585
R3320 GND.n6625 GND.n6624 585
R3321 GND.n2908 GND.n2906 585
R3322 GND.n5629 GND.n2906 585
R3323 GND.n5579 GND.n5576 585
R3324 GND.n5579 GND.n5578 585
R3325 GND.n5581 GND.n5580 585
R3326 GND.n5580 GND.n3244 585
R3327 GND.n5582 GND.n3268 585
R3328 GND.n3268 GND.n3249 585
R3329 GND.n5584 GND.n5583 585
R3330 GND.n5585 GND.n5584 585
R3331 GND.n3269 GND.n3267 585
R3332 GND.n3267 GND.n3258 585
R3333 GND.n5568 GND.n5567 585
R3334 GND.n5567 GND.n3263 585
R3335 GND.n5566 GND.n3271 585
R3336 GND.n5566 GND.n5565 585
R3337 GND.n5545 GND.n3272 585
R3338 GND.n3278 GND.n3272 585
R3339 GND.n5547 GND.n5546 585
R3340 GND.n5548 GND.n5547 585
R3341 GND.n3289 GND.n3288 585
R3342 GND.n3296 GND.n3288 585
R3343 GND.n5540 GND.n5539 585
R3344 GND.n5539 GND.n5538 585
R3345 GND.n3292 GND.n3291 585
R3346 GND.n3300 GND.n3292 585
R3347 GND.n5495 GND.n3317 585
R3348 GND.n3317 GND.n3310 585
R3349 GND.n5497 GND.n5496 585
R3350 GND.n5498 GND.n5497 585
R3351 GND.n3318 GND.n3316 585
R3352 GND.n3316 GND.n3314 585
R3353 GND.n5490 GND.n5489 585
R3354 GND.n5489 GND.n5488 585
R3355 GND.n3321 GND.n3320 585
R3356 GND.n5480 GND.n3321 585
R3357 GND.n5452 GND.n5451 585
R3358 GND.n5453 GND.n5452 585
R3359 GND.n3335 GND.n3334 585
R3360 GND.n5437 GND.n3334 585
R3361 GND.n5447 GND.n5446 585
R3362 GND.n5446 GND.n5445 585
R3363 GND.n3338 GND.n3337 585
R3364 GND.n5429 GND.n3338 585
R3365 GND.n5417 GND.n5416 585
R3366 GND.n5418 GND.n5417 585
R3367 GND.n3356 GND.n3355 585
R3368 GND.n3355 GND.n3351 585
R3369 GND.n5412 GND.n5411 585
R3370 GND.n5411 GND.n5410 585
R3371 GND.n3359 GND.n3358 585
R3372 GND.n3365 GND.n3359 585
R3373 GND.n5391 GND.n5390 585
R3374 GND.n5392 GND.n5391 585
R3375 GND.n3375 GND.n3374 585
R3376 GND.n3382 GND.n3374 585
R3377 GND.n5386 GND.n5385 585
R3378 GND.n5385 GND.n5384 585
R3379 GND.n3378 GND.n3377 585
R3380 GND.n3386 GND.n3378 585
R3381 GND.n5317 GND.n3403 585
R3382 GND.n3403 GND.n3396 585
R3383 GND.n5319 GND.n5318 585
R3384 GND.n5320 GND.n5319 585
R3385 GND.n3404 GND.n3402 585
R3386 GND.n3402 GND.n3400 585
R3387 GND.n5312 GND.n5311 585
R3388 GND.n5311 GND.n5310 585
R3389 GND.n3407 GND.n3406 585
R3390 GND.n5302 GND.n3407 585
R3391 GND.n5274 GND.n5273 585
R3392 GND.n5275 GND.n5274 585
R3393 GND.n3421 GND.n3420 585
R3394 GND.n5259 GND.n3420 585
R3395 GND.n5269 GND.n5268 585
R3396 GND.n5268 GND.n5267 585
R3397 GND.n3424 GND.n3423 585
R3398 GND.n5251 GND.n3424 585
R3399 GND.n5240 GND.n5239 585
R3400 GND.n5241 GND.n5240 585
R3401 GND.n3443 GND.n3442 585
R3402 GND.n3442 GND.n3438 585
R3403 GND.n5235 GND.n5234 585
R3404 GND.n5234 GND.n5233 585
R3405 GND.n3446 GND.n3445 585
R3406 GND.n3452 GND.n3446 585
R3407 GND.n5214 GND.n5213 585
R3408 GND.n5215 GND.n5214 585
R3409 GND.n3464 GND.n3463 585
R3410 GND.n3471 GND.n3463 585
R3411 GND.n5209 GND.n5208 585
R3412 GND.n5208 GND.n5207 585
R3413 GND.n3467 GND.n3466 585
R3414 GND.n3475 GND.n3467 585
R3415 GND.n5143 GND.n3492 585
R3416 GND.n3492 GND.n3485 585
R3417 GND.n5145 GND.n5144 585
R3418 GND.n5146 GND.n5145 585
R3419 GND.n3493 GND.n3491 585
R3420 GND.n3491 GND.n3489 585
R3421 GND.n5138 GND.n5137 585
R3422 GND.n5137 GND.n5136 585
R3423 GND.n3496 GND.n3495 585
R3424 GND.n5128 GND.n3496 585
R3425 GND.n5099 GND.n5098 585
R3426 GND.n5100 GND.n5099 585
R3427 GND.n3510 GND.n3509 585
R3428 GND.n5084 GND.n3509 585
R3429 GND.n5094 GND.n5093 585
R3430 GND.n5093 GND.n5092 585
R3431 GND.n3513 GND.n3512 585
R3432 GND.n5076 GND.n3513 585
R3433 GND.n5065 GND.n5064 585
R3434 GND.n5066 GND.n5065 585
R3435 GND.n3532 GND.n3531 585
R3436 GND.n3531 GND.n3527 585
R3437 GND.n5060 GND.n5059 585
R3438 GND.n5059 GND.n5058 585
R3439 GND.n3535 GND.n3534 585
R3440 GND.n3541 GND.n3535 585
R3441 GND.n5039 GND.n5038 585
R3442 GND.n5040 GND.n5039 585
R3443 GND.n3553 GND.n3552 585
R3444 GND.n3560 GND.n3552 585
R3445 GND.n5034 GND.n5033 585
R3446 GND.n5033 GND.n5032 585
R3447 GND.n3556 GND.n3555 585
R3448 GND.n3564 GND.n3556 585
R3449 GND.n4967 GND.n3581 585
R3450 GND.n3581 GND.n3574 585
R3451 GND.n4969 GND.n4968 585
R3452 GND.n4970 GND.n4969 585
R3453 GND.n3582 GND.n3580 585
R3454 GND.n3580 GND.n3578 585
R3455 GND.n4962 GND.n4961 585
R3456 GND.n4961 GND.n4960 585
R3457 GND.n3585 GND.n3584 585
R3458 GND.n4952 GND.n3585 585
R3459 GND.n4924 GND.n4923 585
R3460 GND.n4925 GND.n4924 585
R3461 GND.n3599 GND.n3598 585
R3462 GND.n4909 GND.n3598 585
R3463 GND.n4919 GND.n4918 585
R3464 GND.n4918 GND.n4917 585
R3465 GND.n3602 GND.n3601 585
R3466 GND.n4901 GND.n3602 585
R3467 GND.n4890 GND.n4889 585
R3468 GND.n4891 GND.n4890 585
R3469 GND.n3621 GND.n3620 585
R3470 GND.n3620 GND.n3616 585
R3471 GND.n4885 GND.n4884 585
R3472 GND.n4884 GND.n4883 585
R3473 GND.n3624 GND.n3623 585
R3474 GND.n3630 GND.n3624 585
R3475 GND.n4863 GND.n4862 585
R3476 GND.n4864 GND.n4863 585
R3477 GND.n3641 GND.n3640 585
R3478 GND.n3648 GND.n3640 585
R3479 GND.n4858 GND.n4857 585
R3480 GND.n4857 GND.n4856 585
R3481 GND.n3644 GND.n3643 585
R3482 GND.n3652 GND.n3644 585
R3483 GND.n4790 GND.n3669 585
R3484 GND.n3669 GND.n3662 585
R3485 GND.n4792 GND.n4791 585
R3486 GND.n4793 GND.n4792 585
R3487 GND.n3670 GND.n3668 585
R3488 GND.n3668 GND.n3666 585
R3489 GND.n4785 GND.n4784 585
R3490 GND.n4784 GND.n4783 585
R3491 GND.n3673 GND.n3672 585
R3492 GND.n4775 GND.n3673 585
R3493 GND.n4747 GND.n4746 585
R3494 GND.n4748 GND.n4747 585
R3495 GND.n3687 GND.n3686 585
R3496 GND.n4732 GND.n3686 585
R3497 GND.n4742 GND.n4741 585
R3498 GND.n4741 GND.n4740 585
R3499 GND.n3690 GND.n3689 585
R3500 GND.n4724 GND.n3690 585
R3501 GND.n4712 GND.n4711 585
R3502 GND.n4713 GND.n4712 585
R3503 GND.n3708 GND.n3707 585
R3504 GND.n3707 GND.n3703 585
R3505 GND.n4707 GND.n4706 585
R3506 GND.n4706 GND.n4705 585
R3507 GND.n3711 GND.n3710 585
R3508 GND.n3717 GND.n3711 585
R3509 GND.n4686 GND.n4685 585
R3510 GND.n4687 GND.n4686 585
R3511 GND.n3729 GND.n3728 585
R3512 GND.n3736 GND.n3728 585
R3513 GND.n4681 GND.n4680 585
R3514 GND.n4680 GND.n4679 585
R3515 GND.n3732 GND.n3731 585
R3516 GND.n3740 GND.n3732 585
R3517 GND.n4614 GND.n3757 585
R3518 GND.n3757 GND.n3750 585
R3519 GND.n4616 GND.n4615 585
R3520 GND.n4617 GND.n4616 585
R3521 GND.n3758 GND.n3756 585
R3522 GND.n3756 GND.n3754 585
R3523 GND.n4609 GND.n4608 585
R3524 GND.n4608 GND.n4607 585
R3525 GND.n3761 GND.n3760 585
R3526 GND.n4599 GND.n3761 585
R3527 GND.n4586 GND.n4585 585
R3528 GND.n4587 GND.n4586 585
R3529 GND.n3781 GND.n3780 585
R3530 GND.n4560 GND.n3780 585
R3531 GND.n4581 GND.n4580 585
R3532 GND.n4580 GND.n4579 585
R3533 GND.n3784 GND.n3783 585
R3534 GND.n4568 GND.n3784 585
R3535 GND.n4529 GND.n4528 585
R3536 GND.n4530 GND.n4529 585
R3537 GND.n3799 GND.n3798 585
R3538 GND.n3806 GND.n3798 585
R3539 GND.n4524 GND.n4523 585
R3540 GND.n4523 GND.n4522 585
R3541 GND.n3802 GND.n3801 585
R3542 GND.n3812 GND.n3802 585
R3543 GND.n4483 GND.n3829 585
R3544 GND.n3829 GND.n3822 585
R3545 GND.n4485 GND.n4484 585
R3546 GND.n4486 GND.n4485 585
R3547 GND.n3830 GND.n3828 585
R3548 GND.n4460 GND.n3828 585
R3549 GND.n4478 GND.n4477 585
R3550 GND.n4477 GND.n4476 585
R3551 GND.n3833 GND.n3832 585
R3552 GND.n4468 GND.n3833 585
R3553 GND.n4401 GND.n4398 585
R3554 GND.n4401 GND.n4400 585
R3555 GND.n4402 GND.n4395 585
R3556 GND.n4402 GND.n3846 585
R3557 GND.n4404 GND.n4403 585
R3558 GND.n4403 GND.n3851 585
R3559 GND.n4405 GND.n3869 585
R3560 GND.n3869 GND.n3862 585
R3561 GND.n4407 GND.n4406 585
R3562 GND.n4408 GND.n4407 585
R3563 GND.n3870 GND.n3868 585
R3564 GND.n3868 GND.n3866 585
R3565 GND.n4389 GND.n4388 585
R3566 GND.n4388 GND.n4387 585
R3567 GND.n3873 GND.n3872 585
R3568 GND.n4379 GND.n3873 585
R3569 GND.n4356 GND.n4355 585
R3570 GND.n4357 GND.n4356 585
R3571 GND.n3887 GND.n3886 585
R3572 GND.n3892 GND.n3886 585
R3573 GND.n4351 GND.n4350 585
R3574 GND.n4350 GND.n4349 585
R3575 GND.n2661 GND.n2660 585
R3576 GND.n3898 GND.n2661 585
R3577 GND.n6863 GND.n6862 585
R3578 GND.n6862 GND.n6861 585
R3579 GND.n6864 GND.n2655 585
R3580 GND.n4211 GND.n2655 585
R3581 GND.n6866 GND.n6865 585
R3582 GND.n6867 GND.n6866 585
R3583 GND.n2644 GND.n2643 585
R3584 GND.n2647 GND.n2644 585
R3585 GND.n6877 GND.n6876 585
R3586 GND.n6876 GND.n6875 585
R3587 GND.n6878 GND.n2638 585
R3588 GND.n4184 GND.n2638 585
R3589 GND.n6880 GND.n6879 585
R3590 GND.n6881 GND.n6880 585
R3591 GND.n2626 GND.n2625 585
R3592 GND.n2629 GND.n2626 585
R3593 GND.n6891 GND.n6890 585
R3594 GND.n6890 GND.n6889 585
R3595 GND.n6892 GND.n2620 585
R3596 GND.n4171 GND.n2620 585
R3597 GND.n6894 GND.n6893 585
R3598 GND.n6895 GND.n6894 585
R3599 GND.n2608 GND.n2607 585
R3600 GND.n2611 GND.n2608 585
R3601 GND.n6905 GND.n6904 585
R3602 GND.n6904 GND.n6903 585
R3603 GND.n6906 GND.n2602 585
R3604 GND.n4158 GND.n2602 585
R3605 GND.n6908 GND.n6907 585
R3606 GND.n6909 GND.n6908 585
R3607 GND.n2590 GND.n2589 585
R3608 GND.n2599 GND.n2590 585
R3609 GND.n6919 GND.n6918 585
R3610 GND.n6918 GND.n6917 585
R3611 GND.n6920 GND.n2584 585
R3612 GND.n4145 GND.n2584 585
R3613 GND.n6922 GND.n6921 585
R3614 GND.n6923 GND.n6922 585
R3615 GND.n2573 GND.n2572 585
R3616 GND.n2581 GND.n2573 585
R3617 GND.n6933 GND.n6932 585
R3618 GND.n6932 GND.n6931 585
R3619 GND.n6934 GND.n2567 585
R3620 GND.n4131 GND.n2567 585
R3621 GND.n6936 GND.n6935 585
R3622 GND.n6937 GND.n6936 585
R3623 GND.n2555 GND.n2554 585
R3624 GND.n2564 GND.n2555 585
R3625 GND.n6946 GND.n6945 585
R3626 GND.n6945 GND.t136 585
R3627 GND.n6947 GND.n2549 585
R3628 GND.n4118 GND.n2549 585
R3629 GND.n6949 GND.n6948 585
R3630 GND.n6950 GND.n6949 585
R3631 GND.n2537 GND.n2536 585
R3632 GND.n2546 GND.n2537 585
R3633 GND.n6960 GND.n6959 585
R3634 GND.n6959 GND.n6958 585
R3635 GND.n6961 GND.n2531 585
R3636 GND.n2538 GND.n2531 585
R3637 GND.n6963 GND.n6962 585
R3638 GND.n6964 GND.n6963 585
R3639 GND.n2529 GND.n2528 585
R3640 GND.n6965 GND.n2529 585
R3641 GND.n6968 GND.n6967 585
R3642 GND.n6967 GND.n6966 585
R3643 GND.n6969 GND.n1958 585
R3644 GND.n1958 GND.n1956 585
R3645 GND.n6971 GND.n6970 585
R3646 GND.n6972 GND.n6971 585
R3647 GND.n1959 GND.n1957 585
R3648 GND.n1957 GND.n1924 585
R3649 GND.n2522 GND.n2521 585
R3650 GND.n2521 GND.n1382 585
R3651 GND.n2520 GND.n1961 585
R3652 GND.n2520 GND.n1380 585
R3653 GND.n2519 GND.n1963 585
R3654 GND.n2519 GND.n2518 585
R3655 GND.n2487 GND.n1962 585
R3656 GND.n1969 GND.n1962 585
R3657 GND.n2489 GND.n2488 585
R3658 GND.n2490 GND.n2489 585
R3659 GND.n1995 GND.n1994 585
R3660 GND.n1994 GND.n1978 585
R3661 GND.n2481 GND.n2480 585
R3662 GND.n2480 GND.n1976 585
R3663 GND.n2479 GND.n1997 585
R3664 GND.n2479 GND.n1980 585
R3665 GND.n2478 GND.n1999 585
R3666 GND.n2478 GND.n2477 585
R3667 GND.n2373 GND.n1998 585
R3668 GND.n2009 GND.n1998 585
R3669 GND.n2375 GND.n2374 585
R3670 GND.n2374 GND.n2007 585
R3671 GND.n2376 GND.n2366 585
R3672 GND.n2366 GND.n2011 585
R3673 GND.n2378 GND.n2377 585
R3674 GND.n2378 GND.n2018 585
R3675 GND.n2379 GND.n2365 585
R3676 GND.n2379 GND.n2017 585
R3677 GND.n2381 GND.n2380 585
R3678 GND.n2380 GND.n2030 585
R3679 GND.n2382 GND.n2360 585
R3680 GND.n2360 GND.n2028 585
R3681 GND.n2384 GND.n2383 585
R3682 GND.n2384 GND.n2032 585
R3683 GND.n2385 GND.n2359 585
R3684 GND.n2385 GND.n2040 585
R3685 GND.n2387 GND.n2386 585
R3686 GND.n2386 GND.n2039 585
R3687 GND.n2389 GND.n2355 585
R3688 GND.n2355 GND.n2354 585
R3689 GND.n2391 GND.n2390 585
R3690 GND.n2392 GND.n2391 585
R3691 GND.n2357 GND.n2351 585
R3692 GND.n2351 GND.n2082 585
R3693 GND.n2356 GND.n2069 585
R3694 GND.n2080 GND.n2069 585
R3695 GND.n2405 GND.n2404 585
R3696 GND.n2404 GND.n2403 585
R3697 GND.n2406 GND.n2066 585
R3698 GND.n2070 GND.n2066 585
R3699 GND.n2409 GND.n2408 585
R3700 GND.n2410 GND.n2409 585
R3701 GND.n2067 GND.n2065 585
R3702 GND.n2065 GND.n2059 585
R3703 GND.n2243 GND.n2239 585
R3704 GND.n2239 GND.n2057 585
R3705 GND.n2245 GND.n2244 585
R3706 GND.n2245 GND.n2098 585
R3707 GND.n2246 GND.n2238 585
R3708 GND.n2246 GND.n2095 585
R3709 GND.n2248 GND.n2247 585
R3710 GND.n2247 GND.n2107 585
R3711 GND.n2249 GND.n2233 585
R3712 GND.n2233 GND.n2105 585
R3713 GND.n2251 GND.n2250 585
R3714 GND.n2251 GND.n2109 585
R3715 GND.n2252 GND.n2232 585
R3716 GND.n2252 GND.n2118 585
R3717 GND.n2254 GND.n2253 585
R3718 GND.n2253 GND.n2117 585
R3719 GND.n2255 GND.n2227 585
R3720 GND.n2227 GND.n2131 585
R3721 GND.n2257 GND.n2256 585
R3722 GND.n2257 GND.n2128 585
R3723 GND.n2258 GND.n2226 585
R3724 GND.n2258 GND.n2134 585
R3725 GND.n2260 GND.n2259 585
R3726 GND.n2259 GND.n2142 585
R3727 GND.n2261 GND.n2156 585
R3728 GND.n2156 GND.n2141 585
R3729 GND.n2263 GND.n2262 585
R3730 GND.n2264 GND.n2263 585
R3731 GND.n2157 GND.n2155 585
R3732 GND.n2155 GND.n2151 585
R3733 GND.n2220 GND.n2219 585
R3734 GND.n2219 GND.n2218 585
R3735 GND.n2167 GND.n2159 585
R3736 GND.n2167 GND.n1292 585
R3737 GND.n2166 GND.n2165 585
R3738 GND.n2166 GND.n1290 585
R3739 GND.n2161 GND.n2160 585
R3740 GND.n2160 GND.n1243 585
R3741 GND.n1221 GND.n1220 585
R3742 GND.n7180 GND.n1221 585
R3743 GND.n7183 GND.n7182 585
R3744 GND.n7182 GND.n7181 585
R3745 GND.n7184 GND.n1215 585
R3746 GND.n1215 GND.n1214 585
R3747 GND.n7186 GND.n7185 585
R3748 GND.n7187 GND.n7186 585
R3749 GND.n1213 GND.n1212 585
R3750 GND.n7188 GND.n1213 585
R3751 GND.n7191 GND.n7190 585
R3752 GND.n7190 GND.n7189 585
R3753 GND.n7192 GND.n1207 585
R3754 GND.n1207 GND.n1206 585
R3755 GND.n7194 GND.n7193 585
R3756 GND.n7195 GND.n7194 585
R3757 GND.n1205 GND.n1204 585
R3758 GND.n7196 GND.n1205 585
R3759 GND.n7199 GND.n7198 585
R3760 GND.n7198 GND.n7197 585
R3761 GND.n7200 GND.n1199 585
R3762 GND.n1199 GND.n1198 585
R3763 GND.n7202 GND.n7201 585
R3764 GND.n7203 GND.n7202 585
R3765 GND.n1197 GND.n1196 585
R3766 GND.n7204 GND.n1197 585
R3767 GND.n7207 GND.n7206 585
R3768 GND.n7206 GND.n7205 585
R3769 GND.n7208 GND.n1191 585
R3770 GND.n1191 GND.n1190 585
R3771 GND.n7210 GND.n7209 585
R3772 GND.n7211 GND.n7210 585
R3773 GND.n1189 GND.n1188 585
R3774 GND.n7212 GND.n1189 585
R3775 GND.n7215 GND.n7214 585
R3776 GND.n7214 GND.n7213 585
R3777 GND.n7216 GND.n1184 585
R3778 GND.n1184 GND.n1183 585
R3779 GND.n7218 GND.n7217 585
R3780 GND.n7219 GND.n7218 585
R3781 GND.n1182 GND.n1181 585
R3782 GND.n7220 GND.n1182 585
R3783 GND.n7223 GND.n7222 585
R3784 GND.n7222 GND.n7221 585
R3785 GND.n2903 GND.n2899 585
R3786 GND.n3234 GND.n2903 585
R3787 GND.n6632 GND.n2898 585
R3788 GND.n6633 GND.n2897 585
R3789 GND.n6634 GND.n2896 585
R3790 GND.n6637 GND.n2891 585
R3791 GND.n6638 GND.n2890 585
R3792 GND.n6639 GND.n2889 585
R3793 GND.n3229 GND.n2887 585
R3794 GND.n6643 GND.n2886 585
R3795 GND.n6644 GND.n2885 585
R3796 GND.n6645 GND.n2884 585
R3797 GND.n3226 GND.n2882 585
R3798 GND.n6649 GND.n2881 585
R3799 GND.n6650 GND.n2880 585
R3800 GND.n6651 GND.n2879 585
R3801 GND.n3223 GND.n2877 585
R3802 GND.n6655 GND.n2876 585
R3803 GND.n6656 GND.n2875 585
R3804 GND.n6657 GND.n2874 585
R3805 GND.n3220 GND.n2832 585
R3806 GND.n6661 GND.n2831 585
R3807 GND.n6662 GND.n2830 585
R3808 GND.n6663 GND.n2829 585
R3809 GND.n6628 GND.n6627 585
R3810 GND.n6627 GND.n6626 585
R3811 GND.n2902 GND.n2901 585
R3812 GND.n3239 GND.n2902 585
R3813 GND.n3254 GND.n3252 585
R3814 GND.n3252 GND.n3245 585
R3815 GND.n5610 GND.n5609 585
R3816 GND.n5613 GND.n5610 585
R3817 GND.n3253 GND.n3251 585
R3818 GND.n5586 GND.n3251 585
R3819 GND.n5604 GND.n5603 585
R3820 GND.n5603 GND.n5602 585
R3821 GND.n3257 GND.n3256 585
R3822 GND.n5594 GND.n3257 585
R3823 GND.n5517 GND.n3274 585
R3824 GND.n5564 GND.n3274 585
R3825 GND.n5520 GND.n5516 585
R3826 GND.n5516 GND.n3279 585
R3827 GND.n5521 GND.n5515 585
R3828 GND.n5515 GND.n3287 585
R3829 GND.n5522 GND.n5514 585
R3830 GND.n5514 GND.n3284 585
R3831 GND.n3304 GND.n3294 585
R3832 GND.n5537 GND.n3294 585
R3833 GND.n5527 GND.n5526 585
R3834 GND.n5528 GND.n5527 585
R3835 GND.n3303 GND.n3302 585
R3836 GND.n5466 GND.n3302 585
R3837 GND.n5510 GND.n5509 585
R3838 GND.n5509 GND.n5508 585
R3839 GND.n3307 GND.n3306 585
R3840 GND.n5500 GND.n3307 585
R3841 GND.n5352 GND.n5351 585
R3842 GND.n5351 GND.n3324 585
R3843 GND.n5355 GND.n5350 585
R3844 GND.n5350 GND.n3322 585
R3845 GND.n5356 GND.n5349 585
R3846 GND.n5349 GND.n3328 585
R3847 GND.n5357 GND.n5348 585
R3848 GND.n5348 GND.n3333 585
R3849 GND.n5347 GND.n5345 585
R3850 GND.n5347 GND.n3341 585
R3851 GND.n5361 GND.n5344 585
R3852 GND.n5344 GND.n3339 585
R3853 GND.n5362 GND.n5343 585
R3854 GND.n5343 GND.n3347 585
R3855 GND.n5363 GND.n3353 585
R3856 GND.n5421 GND.n3353 585
R3857 GND.n5341 GND.n3361 585
R3858 GND.n5409 GND.n3361 585
R3859 GND.n5367 GND.n5340 585
R3860 GND.n5340 GND.n3366 585
R3861 GND.n5368 GND.n5339 585
R3862 GND.n5339 GND.n5338 585
R3863 GND.n5369 GND.n5336 585
R3864 GND.n5336 GND.n3372 585
R3865 GND.n3390 GND.n3380 585
R3866 GND.n5383 GND.n3380 585
R3867 GND.n5374 GND.n5373 585
R3868 GND.n5375 GND.n5374 585
R3869 GND.n3389 GND.n3388 585
R3870 GND.n5288 GND.n3388 585
R3871 GND.n5332 GND.n5331 585
R3872 GND.n5331 GND.n5330 585
R3873 GND.n3393 GND.n3392 585
R3874 GND.n5321 GND.n3393 585
R3875 GND.n5175 GND.n5174 585
R3876 GND.n5174 GND.n3410 585
R3877 GND.n5178 GND.n5173 585
R3878 GND.n5173 GND.n3408 585
R3879 GND.n5179 GND.n5172 585
R3880 GND.n5172 GND.n3415 585
R3881 GND.n5180 GND.n5171 585
R3882 GND.n5171 GND.n3419 585
R3883 GND.n5170 GND.n5168 585
R3884 GND.n5170 GND.n3430 585
R3885 GND.n5184 GND.n5167 585
R3886 GND.n5167 GND.n3425 585
R3887 GND.n5185 GND.n5166 585
R3888 GND.n5166 GND.n3434 585
R3889 GND.n5186 GND.n3440 585
R3890 GND.n5243 GND.n3440 585
R3891 GND.n5164 GND.n3448 585
R3892 GND.n5232 GND.n3448 585
R3893 GND.n5190 GND.n5163 585
R3894 GND.n5163 GND.n3453 585
R3895 GND.n5191 GND.n5162 585
R3896 GND.n5162 GND.n3462 585
R3897 GND.n5192 GND.n5161 585
R3898 GND.n5161 GND.n3458 585
R3899 GND.n3479 GND.n3469 585
R3900 GND.n5206 GND.n3469 585
R3901 GND.n5197 GND.n5196 585
R3902 GND.n5198 GND.n5197 585
R3903 GND.n3478 GND.n3477 585
R3904 GND.n5114 GND.n3477 585
R3905 GND.n5157 GND.n5156 585
R3906 GND.n5156 GND.n5155 585
R3907 GND.n3482 GND.n3481 585
R3908 GND.n5147 GND.n3482 585
R3909 GND.n4999 GND.n4998 585
R3910 GND.n4998 GND.n3500 585
R3911 GND.n5002 GND.n4997 585
R3912 GND.n4997 GND.n3498 585
R3913 GND.n5003 GND.n4996 585
R3914 GND.n4996 GND.n3504 585
R3915 GND.n5004 GND.n4995 585
R3916 GND.n4995 GND.n3508 585
R3917 GND.n4994 GND.n4992 585
R3918 GND.n4994 GND.n3517 585
R3919 GND.n5008 GND.n4991 585
R3920 GND.n4991 GND.n3515 585
R3921 GND.n5009 GND.n4990 585
R3922 GND.n4990 GND.n3523 585
R3923 GND.n5010 GND.n3529 585
R3924 GND.n5068 GND.n3529 585
R3925 GND.n4988 GND.n3537 585
R3926 GND.n5057 GND.n3537 585
R3927 GND.n5014 GND.n4987 585
R3928 GND.n4987 GND.n3543 585
R3929 GND.n5015 GND.n4986 585
R3930 GND.n4986 GND.n3551 585
R3931 GND.n5016 GND.n4985 585
R3932 GND.n4985 GND.n3548 585
R3933 GND.n3568 GND.n3558 585
R3934 GND.n5031 GND.n3558 585
R3935 GND.n5021 GND.n5020 585
R3936 GND.n5023 GND.n5021 585
R3937 GND.n3567 GND.n3566 585
R3938 GND.n4938 GND.n3566 585
R3939 GND.n4981 GND.n4980 585
R3940 GND.n4980 GND.n4979 585
R3941 GND.n3571 GND.n3570 585
R3942 GND.n4971 GND.n3571 585
R3943 GND.n4823 GND.n4822 585
R3944 GND.n4822 GND.n3589 585
R3945 GND.n4826 GND.n4821 585
R3946 GND.n4821 GND.n3586 585
R3947 GND.n4827 GND.n4820 585
R3948 GND.n4820 GND.n3593 585
R3949 GND.n4828 GND.n4819 585
R3950 GND.n4819 GND.n3597 585
R3951 GND.n4818 GND.n4816 585
R3952 GND.n4818 GND.n3606 585
R3953 GND.n4832 GND.n4815 585
R3954 GND.n4815 GND.n3603 585
R3955 GND.n4833 GND.n4814 585
R3956 GND.n4814 GND.n3612 585
R3957 GND.n4834 GND.n3618 585
R3958 GND.n4893 GND.n3618 585
R3959 GND.n4812 GND.n3626 585
R3960 GND.n4882 GND.n3626 585
R3961 GND.n4838 GND.n4811 585
R3962 GND.n4811 GND.n3631 585
R3963 GND.n4839 GND.n4810 585
R3964 GND.n4810 GND.n3639 585
R3965 GND.n4840 GND.n4809 585
R3966 GND.n4809 GND.n3636 585
R3967 GND.n3656 GND.n3646 585
R3968 GND.n4855 GND.n3646 585
R3969 GND.n4845 GND.n4844 585
R3970 GND.n4846 GND.n4845 585
R3971 GND.n3655 GND.n3654 585
R3972 GND.n4761 GND.n3654 585
R3973 GND.n4805 GND.n4804 585
R3974 GND.n4804 GND.n4803 585
R3975 GND.n3659 GND.n3658 585
R3976 GND.n4795 GND.n3659 585
R3977 GND.n4647 GND.n4646 585
R3978 GND.n4646 GND.n3676 585
R3979 GND.n4650 GND.n4645 585
R3980 GND.n4645 GND.n3674 585
R3981 GND.n4651 GND.n4644 585
R3982 GND.n4644 GND.n3680 585
R3983 GND.n4652 GND.n4643 585
R3984 GND.n4643 GND.n3685 585
R3985 GND.n4642 GND.n4640 585
R3986 GND.n4642 GND.n3693 585
R3987 GND.n4656 GND.n4639 585
R3988 GND.n4639 GND.n3691 585
R3989 GND.n4657 GND.n4638 585
R3990 GND.n4638 GND.n3699 585
R3991 GND.n4658 GND.n3705 585
R3992 GND.n4716 GND.n3705 585
R3993 GND.n4636 GND.n3713 585
R3994 GND.n4704 GND.n3713 585
R3995 GND.n4662 GND.n4635 585
R3996 GND.n4635 GND.n3718 585
R3997 GND.n4663 GND.n4634 585
R3998 GND.n4634 GND.n3727 585
R3999 GND.n4664 GND.n4633 585
R4000 GND.n4633 GND.n3724 585
R4001 GND.n3744 GND.n3734 585
R4002 GND.n4678 GND.n3734 585
R4003 GND.n4669 GND.n4668 585
R4004 GND.n4670 GND.n4669 585
R4005 GND.n3743 GND.n3742 585
R4006 GND.n4544 GND.n3742 585
R4007 GND.n4629 GND.n4628 585
R4008 GND.n4628 GND.n4627 585
R4009 GND.n3747 GND.n3746 585
R4010 GND.n4618 GND.n3747 585
R4011 GND.n3774 GND.n3772 585
R4012 GND.n3772 GND.n3763 585
R4013 GND.n4596 GND.n4595 585
R4014 GND.n4597 GND.n4596 585
R4015 GND.n3773 GND.n3771 585
R4016 GND.n3771 GND.n3768 585
R4017 GND.n4590 GND.n4589 585
R4018 GND.n4589 GND.n4588 585
R4019 GND.n3777 GND.n3776 585
R4020 GND.n3787 GND.n3777 585
R4021 GND.n4504 GND.n4502 585
R4022 GND.n4502 GND.n3785 585
R4023 GND.n4505 GND.n4501 585
R4024 GND.n4501 GND.n3793 585
R4025 GND.n4506 GND.n4500 585
R4026 GND.n4500 GND.n3797 585
R4027 GND.n3816 GND.n3804 585
R4028 GND.n4521 GND.n3804 585
R4029 GND.n4511 GND.n4510 585
R4030 GND.n4512 GND.n4511 585
R4031 GND.n3815 GND.n3814 585
R4032 GND.n4452 GND.n3814 585
R4033 GND.n4496 GND.n4495 585
R4034 GND.n4495 GND.n4494 585
R4035 GND.n3819 GND.n3818 585
R4036 GND.n3826 GND.n3819 585
R4037 GND.n4427 GND.n4425 585
R4038 GND.n4425 GND.n3837 585
R4039 GND.n4428 GND.n4424 585
R4040 GND.n4424 GND.n3835 585
R4041 GND.n4429 GND.n4423 585
R4042 GND.n4423 GND.n3841 585
R4043 GND.n3856 GND.n3854 585
R4044 GND.n3854 GND.n3847 585
R4045 GND.n4434 GND.n4433 585
R4046 GND.n4436 GND.n4434 585
R4047 GND.n3855 GND.n3853 585
R4048 GND.n4364 GND.n3853 585
R4049 GND.n4419 GND.n4418 585
R4050 GND.n4418 GND.n4417 585
R4051 GND.n3859 GND.n3858 585
R4052 GND.n4409 GND.n3859 585
R4053 GND.n4328 GND.n4327 585
R4054 GND.n4327 GND.n3877 585
R4055 GND.n4331 GND.n4326 585
R4056 GND.n4326 GND.n3875 585
R4057 GND.n4332 GND.n4325 585
R4058 GND.n4325 GND.n3881 585
R4059 GND.n4333 GND.n4324 585
R4060 GND.n4324 GND.n3885 585
R4061 GND.n3901 GND.n3890 585
R4062 GND.n4348 GND.n3890 585
R4063 GND.n4338 GND.n4337 585
R4064 GND.n4339 GND.n4338 585
R4065 GND.n3900 GND.n2663 585
R4066 GND.n6860 GND.n2663 585
R4067 GND.n4213 GND.n2665 585
R4068 GND.n4315 GND.n4314 585
R4069 GND.n4214 GND.n4212 585
R4070 GND.n4317 GND.n4212 585
R4071 GND.n4270 GND.n4216 585
R4072 GND.n4269 GND.n4217 585
R4073 GND.n4268 GND.n4218 585
R4074 GND.n4221 GND.n4219 585
R4075 GND.n4264 GND.n4222 585
R4076 GND.n4263 GND.n4223 585
R4077 GND.n4262 GND.n4224 585
R4078 GND.n4227 GND.n4225 585
R4079 GND.n4258 GND.n4228 585
R4080 GND.n4257 GND.n4229 585
R4081 GND.n4256 GND.n4230 585
R4082 GND.n4233 GND.n4231 585
R4083 GND.n4252 GND.n4234 585
R4084 GND.n4251 GND.n4235 585
R4085 GND.n4250 GND.n4236 585
R4086 GND.n4242 GND.n4237 585
R4087 GND.n4246 GND.n4243 585
R4088 GND.n4245 GND.n4244 585
R4089 GND.n3904 GND.n3903 585
R4090 GND.n4320 GND.n4319 585
R4091 GND.n6666 GND.n2827 585
R4092 GND.n6626 GND.n2827 585
R4093 GND.n6667 GND.n2826 585
R4094 GND.n3239 GND.n2826 585
R4095 GND.n6668 GND.n2825 585
R4096 GND.n3245 GND.n2825 585
R4097 GND.n5612 GND.n2823 585
R4098 GND.n5613 GND.n5612 585
R4099 GND.n6672 GND.n2822 585
R4100 GND.n5586 GND.n2822 585
R4101 GND.n6673 GND.n2821 585
R4102 GND.n5602 GND.n2821 585
R4103 GND.n6674 GND.n2820 585
R4104 GND.n5594 GND.n2820 585
R4105 GND.n5563 GND.n2818 585
R4106 GND.n5564 GND.n5563 585
R4107 GND.n6678 GND.n2817 585
R4108 GND.n3279 GND.n2817 585
R4109 GND.n6679 GND.n2816 585
R4110 GND.n3287 GND.n2816 585
R4111 GND.n6680 GND.n2815 585
R4112 GND.n3284 GND.n2815 585
R4113 GND.n5536 GND.n2813 585
R4114 GND.n5537 GND.n5536 585
R4115 GND.n6684 GND.n2812 585
R4116 GND.n5528 GND.n2812 585
R4117 GND.n6685 GND.n2811 585
R4118 GND.n5466 GND.n2811 585
R4119 GND.n6686 GND.n2810 585
R4120 GND.n5508 GND.n2810 585
R4121 GND.n5499 GND.n2808 585
R4122 GND.n5500 GND.n5499 585
R4123 GND.n6690 GND.n2807 585
R4124 GND.n3324 GND.n2807 585
R4125 GND.n6691 GND.n2806 585
R4126 GND.n3322 GND.n2806 585
R4127 GND.n6692 GND.n2805 585
R4128 GND.n3328 GND.n2805 585
R4129 GND.n3332 GND.n2803 585
R4130 GND.n3333 GND.n3332 585
R4131 GND.n6696 GND.n2802 585
R4132 GND.n3341 GND.n2802 585
R4133 GND.n6697 GND.n2801 585
R4134 GND.n3339 GND.n2801 585
R4135 GND.n6698 GND.n2800 585
R4136 GND.n3347 GND.n2800 585
R4137 GND.n5420 GND.n2798 585
R4138 GND.n5421 GND.n5420 585
R4139 GND.n6702 GND.n2797 585
R4140 GND.n5409 GND.n2797 585
R4141 GND.n6703 GND.n2796 585
R4142 GND.n3366 GND.n2796 585
R4143 GND.n6704 GND.n2795 585
R4144 GND.n5338 GND.n2795 585
R4145 GND.n3371 GND.n2793 585
R4146 GND.n3372 GND.n3371 585
R4147 GND.n6708 GND.n2792 585
R4148 GND.n5383 GND.n2792 585
R4149 GND.n6709 GND.n2791 585
R4150 GND.n5375 GND.n2791 585
R4151 GND.n6710 GND.n2790 585
R4152 GND.n5288 GND.n2790 585
R4153 GND.n5329 GND.n2788 585
R4154 GND.n5330 GND.n5329 585
R4155 GND.n6714 GND.n2787 585
R4156 GND.n5321 GND.n2787 585
R4157 GND.n6715 GND.n2786 585
R4158 GND.n3410 GND.n2786 585
R4159 GND.n6716 GND.n2785 585
R4160 GND.n3408 GND.n2785 585
R4161 GND.n3414 GND.n2783 585
R4162 GND.n3415 GND.n3414 585
R4163 GND.n6720 GND.n2782 585
R4164 GND.n3419 GND.n2782 585
R4165 GND.n6721 GND.n2781 585
R4166 GND.n3430 GND.n2781 585
R4167 GND.n6722 GND.n2780 585
R4168 GND.n3425 GND.n2780 585
R4169 GND.n3433 GND.n2778 585
R4170 GND.n3434 GND.n3433 585
R4171 GND.n6726 GND.n2777 585
R4172 GND.n5243 GND.n2777 585
R4173 GND.n6727 GND.n2776 585
R4174 GND.n5232 GND.n2776 585
R4175 GND.n6728 GND.n2775 585
R4176 GND.n3453 GND.n2775 585
R4177 GND.n3461 GND.n2773 585
R4178 GND.n3462 GND.n3461 585
R4179 GND.n6732 GND.n2772 585
R4180 GND.n3458 GND.n2772 585
R4181 GND.n6733 GND.n2771 585
R4182 GND.n5206 GND.n2771 585
R4183 GND.n6734 GND.n2770 585
R4184 GND.n5198 GND.n2770 585
R4185 GND.n5113 GND.n2768 585
R4186 GND.n5114 GND.n5113 585
R4187 GND.n6738 GND.n2767 585
R4188 GND.n5155 GND.n2767 585
R4189 GND.n6739 GND.n2766 585
R4190 GND.n5147 GND.n2766 585
R4191 GND.n6740 GND.n2765 585
R4192 GND.n3500 GND.n2765 585
R4193 GND.n3497 GND.n2763 585
R4194 GND.n3498 GND.n3497 585
R4195 GND.n6744 GND.n2762 585
R4196 GND.n3504 GND.n2762 585
R4197 GND.n6745 GND.n2761 585
R4198 GND.n3508 GND.n2761 585
R4199 GND.n6746 GND.n2760 585
R4200 GND.n3517 GND.n2760 585
R4201 GND.n3514 GND.n2758 585
R4202 GND.n3515 GND.n3514 585
R4203 GND.n6750 GND.n2757 585
R4204 GND.n3523 GND.n2757 585
R4205 GND.n6751 GND.n2756 585
R4206 GND.n5068 GND.n2756 585
R4207 GND.n6752 GND.n2755 585
R4208 GND.n5057 GND.n2755 585
R4209 GND.n3542 GND.n2753 585
R4210 GND.n3543 GND.n3542 585
R4211 GND.n6756 GND.n2752 585
R4212 GND.n3551 GND.n2752 585
R4213 GND.n6757 GND.n2751 585
R4214 GND.n3548 GND.n2751 585
R4215 GND.n6758 GND.n2750 585
R4216 GND.n5031 GND.n2750 585
R4217 GND.n5022 GND.n2748 585
R4218 GND.n5023 GND.n5022 585
R4219 GND.n6762 GND.n2747 585
R4220 GND.n4938 GND.n2747 585
R4221 GND.n6763 GND.n2746 585
R4222 GND.n4979 GND.n2746 585
R4223 GND.n6764 GND.n2745 585
R4224 GND.n4971 GND.n2745 585
R4225 GND.n3588 GND.n2743 585
R4226 GND.n3589 GND.n3588 585
R4227 GND.n6768 GND.n2742 585
R4228 GND.n3586 GND.n2742 585
R4229 GND.n6769 GND.n2741 585
R4230 GND.n3593 GND.n2741 585
R4231 GND.n6770 GND.n2740 585
R4232 GND.n3597 GND.n2740 585
R4233 GND.n3605 GND.n2738 585
R4234 GND.n3606 GND.n3605 585
R4235 GND.n6774 GND.n2737 585
R4236 GND.n3603 GND.n2737 585
R4237 GND.n6775 GND.n2736 585
R4238 GND.n3612 GND.n2736 585
R4239 GND.n6776 GND.n2735 585
R4240 GND.n4893 GND.n2735 585
R4241 GND.n4881 GND.n2733 585
R4242 GND.n4882 GND.n4881 585
R4243 GND.n6780 GND.n2732 585
R4244 GND.n3631 GND.n2732 585
R4245 GND.n6781 GND.n2731 585
R4246 GND.n3639 GND.n2731 585
R4247 GND.n6782 GND.n2730 585
R4248 GND.n3636 GND.n2730 585
R4249 GND.n4854 GND.n2728 585
R4250 GND.n4855 GND.n4854 585
R4251 GND.n6786 GND.n2727 585
R4252 GND.n4846 GND.n2727 585
R4253 GND.n6787 GND.n2726 585
R4254 GND.n4761 GND.n2726 585
R4255 GND.n6788 GND.n2725 585
R4256 GND.n4803 GND.n2725 585
R4257 GND.n4794 GND.n2723 585
R4258 GND.n4795 GND.n4794 585
R4259 GND.n6792 GND.n2722 585
R4260 GND.n3676 GND.n2722 585
R4261 GND.n6793 GND.n2721 585
R4262 GND.n3674 GND.n2721 585
R4263 GND.n6794 GND.n2720 585
R4264 GND.n3680 GND.n2720 585
R4265 GND.n3684 GND.n2718 585
R4266 GND.n3685 GND.n3684 585
R4267 GND.n6798 GND.n2717 585
R4268 GND.n3693 GND.n2717 585
R4269 GND.n6799 GND.n2716 585
R4270 GND.n3691 GND.n2716 585
R4271 GND.n6800 GND.n2715 585
R4272 GND.n3699 GND.n2715 585
R4273 GND.n4715 GND.n2713 585
R4274 GND.n4716 GND.n4715 585
R4275 GND.n6804 GND.n2712 585
R4276 GND.n4704 GND.n2712 585
R4277 GND.n6805 GND.n2711 585
R4278 GND.n3718 GND.n2711 585
R4279 GND.n6806 GND.n2710 585
R4280 GND.n3727 GND.n2710 585
R4281 GND.n3723 GND.n2708 585
R4282 GND.n3724 GND.n3723 585
R4283 GND.n6810 GND.n2707 585
R4284 GND.n4678 GND.n2707 585
R4285 GND.n6811 GND.n2706 585
R4286 GND.n4670 GND.n2706 585
R4287 GND.n6812 GND.n2705 585
R4288 GND.n4544 GND.n2705 585
R4289 GND.n4626 GND.n2703 585
R4290 GND.n4627 GND.n4626 585
R4291 GND.n6816 GND.n2702 585
R4292 GND.n4618 GND.n2702 585
R4293 GND.n6817 GND.n2701 585
R4294 GND.n3763 GND.n2701 585
R4295 GND.n6818 GND.n2700 585
R4296 GND.n4597 GND.n2700 585
R4297 GND.n3767 GND.n2698 585
R4298 GND.n3768 GND.n3767 585
R4299 GND.n6822 GND.n2697 585
R4300 GND.n4588 GND.n2697 585
R4301 GND.n6823 GND.n2696 585
R4302 GND.n3787 GND.n2696 585
R4303 GND.n6824 GND.n2695 585
R4304 GND.n3785 GND.n2695 585
R4305 GND.n3792 GND.n2693 585
R4306 GND.n3793 GND.n3792 585
R4307 GND.n6828 GND.n2692 585
R4308 GND.n3797 GND.n2692 585
R4309 GND.n6829 GND.n2691 585
R4310 GND.n4521 GND.n2691 585
R4311 GND.n6830 GND.n2690 585
R4312 GND.n4512 GND.n2690 585
R4313 GND.n4451 GND.n2688 585
R4314 GND.n4452 GND.n4451 585
R4315 GND.n6834 GND.n2687 585
R4316 GND.n4494 GND.n2687 585
R4317 GND.n6835 GND.n2686 585
R4318 GND.n3826 GND.n2686 585
R4319 GND.n6836 GND.n2685 585
R4320 GND.n3837 GND.n2685 585
R4321 GND.n3834 GND.n2683 585
R4322 GND.n3835 GND.n3834 585
R4323 GND.n6840 GND.n2682 585
R4324 GND.n3841 GND.n2682 585
R4325 GND.n6841 GND.n2681 585
R4326 GND.n3847 GND.n2681 585
R4327 GND.n6842 GND.n2680 585
R4328 GND.n4436 GND.n2680 585
R4329 GND.n4363 GND.n2678 585
R4330 GND.n4364 GND.n4363 585
R4331 GND.n6846 GND.n2677 585
R4332 GND.n4417 GND.n2677 585
R4333 GND.n6847 GND.n2676 585
R4334 GND.n4409 GND.n2676 585
R4335 GND.n6848 GND.n2675 585
R4336 GND.n3877 GND.n2675 585
R4337 GND.n3874 GND.n2673 585
R4338 GND.n3875 GND.n3874 585
R4339 GND.n6852 GND.n2672 585
R4340 GND.n3881 GND.n2672 585
R4341 GND.n6853 GND.n2671 585
R4342 GND.n3885 GND.n2671 585
R4343 GND.n6854 GND.n2670 585
R4344 GND.n4348 GND.n2670 585
R4345 GND.n2667 GND.n2666 585
R4346 GND.n4339 GND.n2666 585
R4347 GND.n6859 GND.n6858 585
R4348 GND.n6860 GND.n6859 585
R4349 GND.n3118 GND.n3026 502.111
R4350 GND.n5730 GND.n5729 502.111
R4351 GND.n4109 GND.n4108 502.111
R4352 GND.n3976 GND.n2541 502.111
R4353 GND.n8398 GND.n8397 391.433
R4354 GND.n3937 GND.t140 340.447
R4355 GND.n3188 GND.t104 340.447
R4356 GND.n3944 GND.t91 340.447
R4357 GND.n3173 GND.t170 340.447
R4358 GND.n8217 GND.n8216 301.784
R4359 GND.n8218 GND.n8217 301.784
R4360 GND.n8218 GND.n526 301.784
R4361 GND.n8226 GND.n526 301.784
R4362 GND.n8227 GND.n8226 301.784
R4363 GND.n8228 GND.n8227 301.784
R4364 GND.n8228 GND.n520 301.784
R4365 GND.n8236 GND.n520 301.784
R4366 GND.n8237 GND.n8236 301.784
R4367 GND.n8238 GND.n8237 301.784
R4368 GND.n8238 GND.n514 301.784
R4369 GND.n8246 GND.n514 301.784
R4370 GND.n8247 GND.n8246 301.784
R4371 GND.n8248 GND.n8247 301.784
R4372 GND.n8248 GND.n508 301.784
R4373 GND.n8256 GND.n508 301.784
R4374 GND.n8257 GND.n8256 301.784
R4375 GND.n8258 GND.n8257 301.784
R4376 GND.n8258 GND.n502 301.784
R4377 GND.n8266 GND.n502 301.784
R4378 GND.n8267 GND.n8266 301.784
R4379 GND.n8268 GND.n8267 301.784
R4380 GND.n8268 GND.n496 301.784
R4381 GND.n8276 GND.n496 301.784
R4382 GND.n8277 GND.n8276 301.784
R4383 GND.n8278 GND.n8277 301.784
R4384 GND.n8278 GND.n490 301.784
R4385 GND.n8286 GND.n490 301.784
R4386 GND.n8287 GND.n8286 301.784
R4387 GND.n8288 GND.n8287 301.784
R4388 GND.n8288 GND.n484 301.784
R4389 GND.n8296 GND.n484 301.784
R4390 GND.n8297 GND.n8296 301.784
R4391 GND.n8298 GND.n8297 301.784
R4392 GND.n8298 GND.n478 301.784
R4393 GND.n8306 GND.n478 301.784
R4394 GND.n8307 GND.n8306 301.784
R4395 GND.n8308 GND.n8307 301.784
R4396 GND.n8308 GND.n472 301.784
R4397 GND.n8316 GND.n472 301.784
R4398 GND.n8317 GND.n8316 301.784
R4399 GND.n8318 GND.n8317 301.784
R4400 GND.n8318 GND.n466 301.784
R4401 GND.n8326 GND.n466 301.784
R4402 GND.n8327 GND.n8326 301.784
R4403 GND.n8328 GND.n8327 301.784
R4404 GND.n8328 GND.n460 301.784
R4405 GND.n8336 GND.n460 301.784
R4406 GND.n8337 GND.n8336 301.784
R4407 GND.n8338 GND.n8337 301.784
R4408 GND.n8338 GND.n454 301.784
R4409 GND.n8346 GND.n454 301.784
R4410 GND.n8347 GND.n8346 301.784
R4411 GND.n8348 GND.n8347 301.784
R4412 GND.n8348 GND.n448 301.784
R4413 GND.n8356 GND.n448 301.784
R4414 GND.n8357 GND.n8356 301.784
R4415 GND.n8358 GND.n8357 301.784
R4416 GND.n8358 GND.n442 301.784
R4417 GND.n8366 GND.n442 301.784
R4418 GND.n8367 GND.n8366 301.784
R4419 GND.n8368 GND.n8367 301.784
R4420 GND.n8368 GND.n436 301.784
R4421 GND.n8376 GND.n436 301.784
R4422 GND.n8377 GND.n8376 301.784
R4423 GND.n8378 GND.n8377 301.784
R4424 GND.n8378 GND.n430 301.784
R4425 GND.n8386 GND.n430 301.784
R4426 GND.n8387 GND.n8386 301.784
R4427 GND.n8388 GND.n8387 301.784
R4428 GND.n8388 GND.n424 301.784
R4429 GND.n8397 GND.n424 301.784
R4430 GND.n3966 GND.n3965 294.49
R4431 GND.n3109 GND.n3108 294.49
R4432 GND.n21 GND.n15 289.615
R4433 GND.n36 GND.n30 289.615
R4434 GND.n52 GND.n46 289.615
R4435 GND.n6 GND.n0 289.615
R4436 GND.n82 GND.n76 289.615
R4437 GND.n97 GND.n91 289.615
R4438 GND.n113 GND.n107 289.615
R4439 GND.n129 GND.n123 289.615
R4440 GND.n3977 GND.n2530 256.663
R4441 GND.n3983 GND.n2530 256.663
R4442 GND.n3985 GND.n2530 256.663
R4443 GND.n3991 GND.n2530 256.663
R4444 GND.n3993 GND.n2530 256.663
R4445 GND.n3999 GND.n2530 256.663
R4446 GND.n4001 GND.n2530 256.663
R4447 GND.n4007 GND.n2530 256.663
R4448 GND.n4009 GND.n2530 256.663
R4449 GND.n4015 GND.n2530 256.663
R4450 GND.n4017 GND.n2530 256.663
R4451 GND.n4023 GND.n2530 256.663
R4452 GND.n4025 GND.n2530 256.663
R4453 GND.n4031 GND.n2530 256.663
R4454 GND.n4033 GND.n2530 256.663
R4455 GND.n4039 GND.n2530 256.663
R4456 GND.n4042 GND.n2530 256.663
R4457 GND.n4044 GND.n2530 256.663
R4458 GND.n4050 GND.n2530 256.663
R4459 GND.n4052 GND.n2530 256.663
R4460 GND.n4058 GND.n2530 256.663
R4461 GND.n4060 GND.n2530 256.663
R4462 GND.n4066 GND.n2530 256.663
R4463 GND.n4068 GND.n2530 256.663
R4464 GND.n4074 GND.n2530 256.663
R4465 GND.n4076 GND.n2530 256.663
R4466 GND.n4082 GND.n2530 256.663
R4467 GND.n4084 GND.n2530 256.663
R4468 GND.n4090 GND.n2530 256.663
R4469 GND.n4092 GND.n2530 256.663
R4470 GND.n4098 GND.n2530 256.663
R4471 GND.n4100 GND.n2530 256.663
R4472 GND.n4106 GND.n2530 256.663
R4473 GND.n5726 GND.n3037 256.663
R4474 GND.n5735 GND.n3037 256.663
R4475 GND.n3209 GND.n3037 256.663
R4476 GND.n5742 GND.n3037 256.663
R4477 GND.n3206 GND.n3037 256.663
R4478 GND.n5749 GND.n3037 256.663
R4479 GND.n3203 GND.n3037 256.663
R4480 GND.n5756 GND.n3037 256.663
R4481 GND.n3200 GND.n3037 256.663
R4482 GND.n5763 GND.n3037 256.663
R4483 GND.n3197 GND.n3037 256.663
R4484 GND.n5770 GND.n3037 256.663
R4485 GND.n3194 GND.n3037 256.663
R4486 GND.n5777 GND.n3037 256.663
R4487 GND.n3191 GND.n3037 256.663
R4488 GND.n5785 GND.n3037 256.663
R4489 GND.n5788 GND.n3037 256.663
R4490 GND.n5790 GND.n5789 256.663
R4491 GND.n3185 GND.n3037 256.663
R4492 GND.n3088 GND.n3037 256.663
R4493 GND.n3178 GND.n3037 256.663
R4494 GND.n3169 GND.n3037 256.663
R4495 GND.n3167 GND.n3037 256.663
R4496 GND.n3161 GND.n3037 256.663
R4497 GND.n3159 GND.n3037 256.663
R4498 GND.n3153 GND.n3037 256.663
R4499 GND.n3151 GND.n3037 256.663
R4500 GND.n3145 GND.n3037 256.663
R4501 GND.n3143 GND.n3037 256.663
R4502 GND.n3137 GND.n3037 256.663
R4503 GND.n3135 GND.n3037 256.663
R4504 GND.n3129 GND.n3037 256.663
R4505 GND.n3127 GND.n3037 256.663
R4506 GND.n3121 GND.n3037 256.663
R4507 GND.n3119 GND.n3037 256.663
R4508 GND.n7179 GND.n1237 242.672
R4509 GND.n7179 GND.n1238 242.672
R4510 GND.n7179 GND.n1239 242.672
R4511 GND.n7179 GND.n1240 242.672
R4512 GND.n7179 GND.n1241 242.672
R4513 GND.n6988 GND.n6987 242.672
R4514 GND.n6987 GND.n1955 242.672
R4515 GND.n6987 GND.n1938 242.672
R4516 GND.n6987 GND.n1937 242.672
R4517 GND.n6987 GND.n1936 242.672
R4518 GND.n7179 GND.n7178 242.672
R4519 GND.n7179 GND.n1222 242.672
R4520 GND.n7179 GND.n1223 242.672
R4521 GND.n7179 GND.n1224 242.672
R4522 GND.n7179 GND.n1225 242.672
R4523 GND.n7179 GND.n1226 242.672
R4524 GND.n7179 GND.n1227 242.672
R4525 GND.n7179 GND.n1228 242.672
R4526 GND.n7179 GND.n1229 242.672
R4527 GND.n7179 GND.n1230 242.672
R4528 GND.n7179 GND.n1231 242.672
R4529 GND.n7179 GND.n1232 242.672
R4530 GND.n7179 GND.n1233 242.672
R4531 GND.n7179 GND.n1234 242.672
R4532 GND.n7179 GND.n1235 242.672
R4533 GND.n7179 GND.n1236 242.672
R4534 GND.n6987 GND.n6973 242.672
R4535 GND.n6987 GND.n6974 242.672
R4536 GND.n6987 GND.n6976 242.672
R4537 GND.n6987 GND.n6977 242.672
R4538 GND.n6987 GND.n6979 242.672
R4539 GND.n6987 GND.n6980 242.672
R4540 GND.n6987 GND.n6982 242.672
R4541 GND.n6987 GND.n6983 242.672
R4542 GND.n6987 GND.n6985 242.672
R4543 GND.n7020 GND.n1406 242.672
R4544 GND.n6987 GND.n1934 242.672
R4545 GND.n6987 GND.n1933 242.672
R4546 GND.n6987 GND.n1931 242.672
R4547 GND.n6987 GND.n1930 242.672
R4548 GND.n6987 GND.n1928 242.672
R4549 GND.n6987 GND.n1927 242.672
R4550 GND.n6987 GND.n1925 242.672
R4551 GND.n6512 GND.n3061 242.672
R4552 GND.n6512 GND.n3062 242.672
R4553 GND.n6512 GND.n3063 242.672
R4554 GND.n6512 GND.n3064 242.672
R4555 GND.n6512 GND.n3065 242.672
R4556 GND.n6293 GND.n383 242.672
R4557 GND.n6261 GND.n383 242.672
R4558 GND.n6283 GND.n383 242.672
R4559 GND.n6265 GND.n383 242.672
R4560 GND.n6273 GND.n383 242.672
R4561 GND.n6512 GND.n6511 242.672
R4562 GND.n6512 GND.n3046 242.672
R4563 GND.n6512 GND.n3047 242.672
R4564 GND.n6512 GND.n3048 242.672
R4565 GND.n6512 GND.n3049 242.672
R4566 GND.n6512 GND.n3050 242.672
R4567 GND.n6512 GND.n3051 242.672
R4568 GND.n6512 GND.n3052 242.672
R4569 GND.n6512 GND.n3053 242.672
R4570 GND.n6512 GND.n3054 242.672
R4571 GND.n6512 GND.n3055 242.672
R4572 GND.n6512 GND.n3056 242.672
R4573 GND.n6512 GND.n3057 242.672
R4574 GND.n6512 GND.n3058 242.672
R4575 GND.n6512 GND.n3059 242.672
R4576 GND.n6512 GND.n3060 242.672
R4577 GND.n383 GND.n262 242.672
R4578 GND.n383 GND.n263 242.672
R4579 GND.n383 GND.n264 242.672
R4580 GND.n383 GND.n265 242.672
R4581 GND.n383 GND.n266 242.672
R4582 GND.n383 GND.n267 242.672
R4583 GND.n383 GND.n268 242.672
R4584 GND.n383 GND.n269 242.672
R4585 GND.n383 GND.n270 242.672
R4586 GND.n383 GND.n271 242.672
R4587 GND.n383 GND.n272 242.672
R4588 GND.n383 GND.n273 242.672
R4589 GND.n383 GND.n274 242.672
R4590 GND.n383 GND.n275 242.672
R4591 GND.n383 GND.n276 242.672
R4592 GND.n383 GND.n277 242.672
R4593 GND.n3234 GND.n3233 242.672
R4594 GND.n3234 GND.n3232 242.672
R4595 GND.n3234 GND.n3231 242.672
R4596 GND.n3234 GND.n3230 242.672
R4597 GND.n3234 GND.n3228 242.672
R4598 GND.n3234 GND.n3227 242.672
R4599 GND.n3234 GND.n3225 242.672
R4600 GND.n3234 GND.n3224 242.672
R4601 GND.n3234 GND.n3222 242.672
R4602 GND.n3234 GND.n3221 242.672
R4603 GND.n3234 GND.n3219 242.672
R4604 GND.n4317 GND.n4316 242.672
R4605 GND.n4317 GND.n3905 242.672
R4606 GND.n4317 GND.n3906 242.672
R4607 GND.n4317 GND.n3907 242.672
R4608 GND.n4317 GND.n3908 242.672
R4609 GND.n4317 GND.n3909 242.672
R4610 GND.n4317 GND.n3910 242.672
R4611 GND.n4317 GND.n3911 242.672
R4612 GND.n4317 GND.n3912 242.672
R4613 GND.n4317 GND.n3913 242.672
R4614 GND.n4318 GND.n4317 242.672
R4615 GND.n382 GND.n278 240.244
R4616 GND.n375 GND.n374 240.244
R4617 GND.n372 GND.n371 240.244
R4618 GND.n368 GND.n367 240.244
R4619 GND.n364 GND.n363 240.244
R4620 GND.n357 GND.n356 240.244
R4621 GND.n354 GND.n353 240.244
R4622 GND.n350 GND.n349 240.244
R4623 GND.n346 GND.n345 240.244
R4624 GND.n342 GND.n341 240.244
R4625 GND.n302 GND.n301 240.244
R4626 GND.n334 GND.n333 240.244
R4627 GND.n330 GND.n329 240.244
R4628 GND.n326 GND.n325 240.244
R4629 GND.n322 GND.n321 240.244
R4630 GND.n318 GND.n317 240.244
R4631 GND.n6449 GND.n5817 240.244
R4632 GND.n6441 GND.n5817 240.244
R4633 GND.n6441 GND.n5828 240.244
R4634 GND.n5845 GND.n5828 240.244
R4635 GND.n6147 GND.n5845 240.244
R4636 GND.n6147 GND.n5858 240.244
R4637 GND.n6152 GND.n5858 240.244
R4638 GND.n6152 GND.n5869 240.244
R4639 GND.n6162 GND.n5869 240.244
R4640 GND.n6162 GND.n5879 240.244
R4641 GND.n6167 GND.n5879 240.244
R4642 GND.n6167 GND.n5890 240.244
R4643 GND.n6177 GND.n5890 240.244
R4644 GND.n6177 GND.n5900 240.244
R4645 GND.n6182 GND.n5900 240.244
R4646 GND.n6182 GND.n5910 240.244
R4647 GND.n6199 GND.n5910 240.244
R4648 GND.n6199 GND.n5919 240.244
R4649 GND.n5924 GND.n5919 240.244
R4650 GND.n6205 GND.n5924 240.244
R4651 GND.n6205 GND.n5933 240.244
R4652 GND.n5933 GND.n142 240.244
R4653 GND.n5941 GND.n142 240.244
R4654 GND.n5975 GND.n5941 240.244
R4655 GND.n6214 GND.n5975 240.244
R4656 GND.n6214 GND.n161 240.244
R4657 GND.n6224 GND.n161 240.244
R4658 GND.n6224 GND.n173 240.244
R4659 GND.n6229 GND.n173 240.244
R4660 GND.n6229 GND.n183 240.244
R4661 GND.n6240 GND.n183 240.244
R4662 GND.n6240 GND.n193 240.244
R4663 GND.n5959 GND.n193 240.244
R4664 GND.n5959 GND.n203 240.244
R4665 GND.n6346 GND.n203 240.244
R4666 GND.n6346 GND.n213 240.244
R4667 GND.n6342 GND.n213 240.244
R4668 GND.n6342 GND.n224 240.244
R4669 GND.n6307 GND.n224 240.244
R4670 GND.n6307 GND.n233 240.244
R4671 GND.n6303 GND.n233 240.244
R4672 GND.n6303 GND.n244 240.244
R4673 GND.n8447 GND.n244 240.244
R4674 GND.n3069 GND.n3068 240.244
R4675 GND.n6505 GND.n3068 240.244
R4676 GND.n6503 GND.n6502 240.244
R4677 GND.n6499 GND.n6498 240.244
R4678 GND.n6495 GND.n6494 240.244
R4679 GND.n6491 GND.n6490 240.244
R4680 GND.n6487 GND.n6486 240.244
R4681 GND.n6483 GND.n5791 240.244
R4682 GND.n6481 GND.n6480 240.244
R4683 GND.n6477 GND.n6476 240.244
R4684 GND.n6472 GND.n5798 240.244
R4685 GND.n6470 GND.n6469 240.244
R4686 GND.n6466 GND.n6465 240.244
R4687 GND.n6462 GND.n6461 240.244
R4688 GND.n6458 GND.n6457 240.244
R4689 GND.n5812 GND.n5811 240.244
R4690 GND.n5833 GND.n3070 240.244
R4691 GND.n6439 GND.n5833 240.244
R4692 GND.n6439 GND.n5834 240.244
R4693 GND.n6435 GND.n5834 240.244
R4694 GND.n6435 GND.n5843 240.244
R4695 GND.n6427 GND.n5843 240.244
R4696 GND.n6427 GND.n5861 240.244
R4697 GND.n6423 GND.n5861 240.244
R4698 GND.n6423 GND.n5867 240.244
R4699 GND.n6415 GND.n5867 240.244
R4700 GND.n6415 GND.n5882 240.244
R4701 GND.n6411 GND.n5882 240.244
R4702 GND.n6411 GND.n5888 240.244
R4703 GND.n6403 GND.n5888 240.244
R4704 GND.n6403 GND.n5903 240.244
R4705 GND.n6399 GND.n5903 240.244
R4706 GND.n6399 GND.n5908 240.244
R4707 GND.n6391 GND.n5908 240.244
R4708 GND.n6391 GND.n6389 240.244
R4709 GND.n6389 GND.n5923 240.244
R4710 GND.n5923 GND.n145 240.244
R4711 GND.n8507 GND.n145 240.244
R4712 GND.n8507 GND.n146 240.244
R4713 GND.n5943 GND.n146 240.244
R4714 GND.n5943 GND.n158 240.244
R4715 GND.n8502 GND.n158 240.244
R4716 GND.n8502 GND.n159 240.244
R4717 GND.n8494 GND.n159 240.244
R4718 GND.n8494 GND.n176 240.244
R4719 GND.n8490 GND.n176 240.244
R4720 GND.n8490 GND.n181 240.244
R4721 GND.n8482 GND.n181 240.244
R4722 GND.n8482 GND.n195 240.244
R4723 GND.n8478 GND.n195 240.244
R4724 GND.n8478 GND.n201 240.244
R4725 GND.n8470 GND.n201 240.244
R4726 GND.n8470 GND.n216 240.244
R4727 GND.n8466 GND.n216 240.244
R4728 GND.n8466 GND.n222 240.244
R4729 GND.n8458 GND.n222 240.244
R4730 GND.n8458 GND.n236 240.244
R4731 GND.n8454 GND.n236 240.244
R4732 GND.n8454 GND.n242 240.244
R4733 GND.n6272 GND.n6271 240.244
R4734 GND.n6275 GND.n6274 240.244
R4735 GND.n6282 GND.n6281 240.244
R4736 GND.n6285 GND.n6284 240.244
R4737 GND.n6292 GND.n6291 240.244
R4738 GND.n6052 GND.n5820 240.244
R4739 GND.n6052 GND.n5830 240.244
R4740 GND.n6139 GND.n5830 240.244
R4741 GND.n6139 GND.n5846 240.244
R4742 GND.n6145 GND.n5846 240.244
R4743 GND.n6145 GND.n5859 240.244
R4744 GND.n6154 GND.n5859 240.244
R4745 GND.n6154 GND.n5870 240.244
R4746 GND.n6160 GND.n5870 240.244
R4747 GND.n6160 GND.n5880 240.244
R4748 GND.n6169 GND.n5880 240.244
R4749 GND.n6169 GND.n5891 240.244
R4750 GND.n6175 GND.n5891 240.244
R4751 GND.n6175 GND.n5901 240.244
R4752 GND.n6184 GND.n5901 240.244
R4753 GND.n6184 GND.n5911 240.244
R4754 GND.n6197 GND.n5911 240.244
R4755 GND.n6197 GND.n5920 240.244
R4756 GND.n5925 GND.n5920 240.244
R4757 GND.n6192 GND.n5925 240.244
R4758 GND.n6192 GND.n140 240.244
R4759 GND.n8509 GND.n140 240.244
R4760 GND.n8509 GND.n141 240.244
R4761 GND.n5973 GND.n141 240.244
R4762 GND.n6216 GND.n5973 240.244
R4763 GND.n6216 GND.n162 240.244
R4764 GND.n6222 GND.n162 240.244
R4765 GND.n6222 GND.n174 240.244
R4766 GND.n6231 GND.n174 240.244
R4767 GND.n6231 GND.n184 240.244
R4768 GND.n6238 GND.n184 240.244
R4769 GND.n6238 GND.n194 240.244
R4770 GND.n6352 GND.n194 240.244
R4771 GND.n6352 GND.n204 240.244
R4772 GND.n6348 GND.n204 240.244
R4773 GND.n6348 GND.n214 240.244
R4774 GND.n6340 GND.n214 240.244
R4775 GND.n6340 GND.n225 240.244
R4776 GND.n6336 GND.n225 240.244
R4777 GND.n6336 GND.n234 240.244
R4778 GND.n6301 GND.n234 240.244
R4779 GND.n6301 GND.n245 240.244
R4780 GND.n252 GND.n245 240.244
R4781 GND.n6130 GND.n6129 240.244
R4782 GND.n6126 GND.n6125 240.244
R4783 GND.n6122 GND.n6121 240.244
R4784 GND.n6118 GND.n6117 240.244
R4785 GND.n6112 GND.n3066 240.244
R4786 GND.n6447 GND.n5823 240.244
R4787 GND.n5832 GND.n5823 240.244
R4788 GND.n5848 GND.n5832 240.244
R4789 GND.n6433 GND.n5848 240.244
R4790 GND.n6433 GND.n5849 240.244
R4791 GND.n6429 GND.n5849 240.244
R4792 GND.n6429 GND.n5856 240.244
R4793 GND.n6421 GND.n5856 240.244
R4794 GND.n6421 GND.n5872 240.244
R4795 GND.n6417 GND.n5872 240.244
R4796 GND.n6417 GND.n5877 240.244
R4797 GND.n6409 GND.n5877 240.244
R4798 GND.n6409 GND.n5893 240.244
R4799 GND.n6405 GND.n5893 240.244
R4800 GND.n6405 GND.n5898 240.244
R4801 GND.n6397 GND.n5898 240.244
R4802 GND.n6397 GND.n5912 240.244
R4803 GND.n6393 GND.n5912 240.244
R4804 GND.n6393 GND.n5917 240.244
R4805 GND.n5934 GND.n5917 240.244
R4806 GND.n6378 GND.n5934 240.244
R4807 GND.n6378 GND.n144 240.244
R4808 GND.n6374 GND.n144 240.244
R4809 GND.n6374 GND.n5940 240.244
R4810 GND.n5940 GND.n164 240.244
R4811 GND.n8500 GND.n164 240.244
R4812 GND.n8500 GND.n165 240.244
R4813 GND.n8496 GND.n165 240.244
R4814 GND.n8496 GND.n171 240.244
R4815 GND.n8488 GND.n171 240.244
R4816 GND.n8488 GND.n186 240.244
R4817 GND.n8484 GND.n186 240.244
R4818 GND.n8484 GND.n191 240.244
R4819 GND.n8476 GND.n191 240.244
R4820 GND.n8476 GND.n206 240.244
R4821 GND.n8472 GND.n206 240.244
R4822 GND.n8472 GND.n211 240.244
R4823 GND.n8464 GND.n211 240.244
R4824 GND.n8464 GND.n227 240.244
R4825 GND.n8460 GND.n227 240.244
R4826 GND.n8460 GND.n232 240.244
R4827 GND.n8452 GND.n232 240.244
R4828 GND.n8452 GND.n247 240.244
R4829 GND.n1390 GND.n1389 240.244
R4830 GND.n1926 GND.n1393 240.244
R4831 GND.n1395 GND.n1394 240.244
R4832 GND.n1929 GND.n1398 240.244
R4833 GND.n1402 GND.n1401 240.244
R4834 GND.n1932 GND.n1405 240.244
R4835 GND.n6986 GND.n1408 240.244
R4836 GND.n6984 GND.n1411 240.244
R4837 GND.n1413 GND.n1412 240.244
R4838 GND.n6981 GND.n1418 240.244
R4839 GND.n1420 GND.n1419 240.244
R4840 GND.n6978 GND.n1423 240.244
R4841 GND.n1425 GND.n1424 240.244
R4842 GND.n6975 GND.n1428 240.244
R4843 GND.n1433 GND.n1429 240.244
R4844 GND.n7114 GND.n1288 240.244
R4845 GND.n1297 GND.n1288 240.244
R4846 GND.n1298 GND.n1297 240.244
R4847 GND.n2265 GND.n1298 240.244
R4848 GND.n2265 GND.n1304 240.244
R4849 GND.n1305 GND.n1304 240.244
R4850 GND.n1306 GND.n1305 240.244
R4851 GND.n2129 GND.n1306 240.244
R4852 GND.n2129 GND.n1312 240.244
R4853 GND.n1313 GND.n1312 240.244
R4854 GND.n1314 GND.n1313 240.244
R4855 GND.n2110 GND.n1314 240.244
R4856 GND.n2110 GND.n1320 240.244
R4857 GND.n1321 GND.n1320 240.244
R4858 GND.n1322 GND.n1321 240.244
R4859 GND.n2096 GND.n1322 240.244
R4860 GND.n2096 GND.n1328 240.244
R4861 GND.n1329 GND.n1328 240.244
R4862 GND.n1330 GND.n1329 240.244
R4863 GND.n2071 GND.n1330 240.244
R4864 GND.n2071 GND.n1336 240.244
R4865 GND.n1337 GND.n1336 240.244
R4866 GND.n1338 GND.n1337 240.244
R4867 GND.n2085 GND.n1338 240.244
R4868 GND.n2085 GND.n1344 240.244
R4869 GND.n1345 GND.n1344 240.244
R4870 GND.n1346 GND.n1345 240.244
R4871 GND.n2033 GND.n1346 240.244
R4872 GND.n2033 GND.n1352 240.244
R4873 GND.n1353 GND.n1352 240.244
R4874 GND.n1354 GND.n1353 240.244
R4875 GND.n2021 GND.n1354 240.244
R4876 GND.n2021 GND.n1360 240.244
R4877 GND.n1361 GND.n1360 240.244
R4878 GND.n1362 GND.n1361 240.244
R4879 GND.n2001 GND.n1362 240.244
R4880 GND.n2001 GND.n1368 240.244
R4881 GND.n1369 GND.n1368 240.244
R4882 GND.n1370 GND.n1369 240.244
R4883 GND.n1967 GND.n1370 240.244
R4884 GND.n1967 GND.n1376 240.244
R4885 GND.n1377 GND.n1376 240.244
R4886 GND.n7045 GND.n1377 240.244
R4887 GND.n1245 GND.n1244 240.244
R4888 GND.n7172 GND.n1244 240.244
R4889 GND.n7170 GND.n7169 240.244
R4890 GND.n7166 GND.n7165 240.244
R4891 GND.n7162 GND.n7161 240.244
R4892 GND.n7158 GND.n7157 240.244
R4893 GND.n7154 GND.n7153 240.244
R4894 GND.n7150 GND.n7149 240.244
R4895 GND.n7146 GND.n7145 240.244
R4896 GND.n7142 GND.n7141 240.244
R4897 GND.n7137 GND.n1269 240.244
R4898 GND.n7135 GND.n7134 240.244
R4899 GND.n7131 GND.n7130 240.244
R4900 GND.n7127 GND.n7126 240.244
R4901 GND.n7123 GND.n7122 240.244
R4902 GND.n1283 GND.n1282 240.244
R4903 GND.n2172 GND.n1246 240.244
R4904 GND.n2172 GND.n2150 240.244
R4905 GND.n2270 GND.n2150 240.244
R4906 GND.n2270 GND.n2144 240.244
R4907 GND.n2278 GND.n2144 240.244
R4908 GND.n2278 GND.n2146 240.244
R4909 GND.n2146 GND.n2127 240.244
R4910 GND.n2294 GND.n2127 240.244
R4911 GND.n2294 GND.n2121 240.244
R4912 GND.n2302 GND.n2121 240.244
R4913 GND.n2302 GND.n2123 240.244
R4914 GND.n2123 GND.n2104 240.244
R4915 GND.n2319 GND.n2104 240.244
R4916 GND.n2319 GND.n2100 240.244
R4917 GND.n2325 GND.n2100 240.244
R4918 GND.n2325 GND.n2055 240.244
R4919 GND.n2415 GND.n2055 240.244
R4920 GND.n2415 GND.n2056 240.244
R4921 GND.n2076 GND.n2056 240.244
R4922 GND.n2078 GND.n2076 240.244
R4923 GND.n2401 GND.n2078 240.244
R4924 GND.n2401 GND.n2398 240.244
R4925 GND.n2398 GND.n2079 240.244
R4926 GND.n2349 GND.n2079 240.244
R4927 GND.n2349 GND.n2043 240.244
R4928 GND.n2422 GND.n2043 240.244
R4929 GND.n2422 GND.n2045 240.244
R4930 GND.n2045 GND.n2027 240.244
R4931 GND.n2440 GND.n2027 240.244
R4932 GND.n2440 GND.n2020 240.244
R4933 GND.n2448 GND.n2020 240.244
R4934 GND.n2448 GND.n2023 240.244
R4935 GND.n2023 GND.n2006 240.244
R4936 GND.n2469 GND.n2006 240.244
R4937 GND.n2469 GND.n2002 240.244
R4938 GND.n2475 GND.n2002 240.244
R4939 GND.n2475 GND.n1975 240.244
R4940 GND.n2502 GND.n1975 240.244
R4941 GND.n2502 GND.n1970 240.244
R4942 GND.n2510 GND.n1970 240.244
R4943 GND.n2510 GND.n1971 240.244
R4944 GND.n1971 GND.n1384 240.244
R4945 GND.n7043 GND.n1384 240.244
R4946 GND.n1939 GND.n1935 240.244
R4947 GND.n1943 GND.n1942 240.244
R4948 GND.n1947 GND.n1946 240.244
R4949 GND.n1951 GND.n1950 240.244
R4950 GND.n1954 GND.n1923 240.244
R4951 GND.n2174 GND.n1291 240.244
R4952 GND.n2216 GND.n2174 240.244
R4953 GND.n2216 GND.n2152 240.244
R4954 GND.n2152 GND.n2140 240.244
R4955 GND.n2280 GND.n2140 240.244
R4956 GND.n2280 GND.n2135 240.244
R4957 GND.n2287 GND.n2135 240.244
R4958 GND.n2287 GND.n2130 240.244
R4959 GND.n2130 GND.n2116 240.244
R4960 GND.n2304 GND.n2116 240.244
R4961 GND.n2304 GND.n2111 240.244
R4962 GND.n2311 GND.n2111 240.244
R4963 GND.n2311 GND.n2106 240.244
R4964 GND.n2106 GND.n2093 240.244
R4965 GND.n2327 GND.n2093 240.244
R4966 GND.n2327 GND.n2094 240.244
R4967 GND.n2094 GND.n2058 240.244
R4968 GND.n2063 GND.n2058 240.244
R4969 GND.n2335 GND.n2063 240.244
R4970 GND.n2335 GND.n2334 240.244
R4971 GND.n2334 GND.n2073 240.244
R4972 GND.n2081 GND.n2073 240.244
R4973 GND.n2084 GND.n2081 240.244
R4974 GND.n2346 GND.n2084 240.244
R4975 GND.n2346 GND.n2038 240.244
R4976 GND.n2424 GND.n2038 240.244
R4977 GND.n2424 GND.n2034 240.244
R4978 GND.n2432 GND.n2034 240.244
R4979 GND.n2432 GND.n2029 240.244
R4980 GND.n2029 GND.n2016 240.244
R4981 GND.n2450 GND.n2016 240.244
R4982 GND.n2450 GND.n2012 240.244
R4983 GND.n2462 GND.n2012 240.244
R4984 GND.n2462 GND.n2008 240.244
R4985 GND.n2458 GND.n2008 240.244
R4986 GND.n2458 GND.n1981 240.244
R4987 GND.n2496 GND.n1981 240.244
R4988 GND.n2496 GND.n1977 240.244
R4989 GND.n2492 GND.n1977 240.244
R4990 GND.n2492 GND.n1968 240.244
R4991 GND.n1991 GND.n1968 240.244
R4992 GND.n1991 GND.n1965 240.244
R4993 GND.n1965 GND.n1381 240.244
R4994 GND.n2193 GND.n2192 240.244
R4995 GND.n2187 GND.n2186 240.244
R4996 GND.n2201 GND.n2200 240.244
R4997 GND.n2183 GND.n2182 240.244
R4998 GND.n2178 GND.n1242 240.244
R4999 GND.n7112 GND.n1294 240.244
R5000 GND.n2154 GND.n1294 240.244
R5001 GND.n2268 GND.n2154 240.244
R5002 GND.n2268 GND.n2267 240.244
R5003 GND.n2267 GND.n2143 240.244
R5004 GND.n2143 GND.n2133 240.244
R5005 GND.n2289 GND.n2133 240.244
R5006 GND.n2292 GND.n2289 240.244
R5007 GND.n2292 GND.n2291 240.244
R5008 GND.n2291 GND.n2120 240.244
R5009 GND.n2120 GND.n2108 240.244
R5010 GND.n2313 GND.n2108 240.244
R5011 GND.n2317 GND.n2313 240.244
R5012 GND.n2317 GND.n2316 240.244
R5013 GND.n2316 GND.n2099 240.244
R5014 GND.n2099 GND.n2060 240.244
R5015 GND.n2413 GND.n2060 240.244
R5016 GND.n2413 GND.n2412 240.244
R5017 GND.n2412 GND.n2061 240.244
R5018 GND.n2074 GND.n2061 240.244
R5019 GND.n2075 GND.n2074 240.244
R5020 GND.n2396 GND.n2075 240.244
R5021 GND.n2396 GND.n2394 240.244
R5022 GND.n2394 GND.n2083 240.244
R5023 GND.n2352 GND.n2083 240.244
R5024 GND.n2352 GND.n2042 240.244
R5025 GND.n2042 GND.n2031 240.244
R5026 GND.n2434 GND.n2031 240.244
R5027 GND.n2438 GND.n2434 240.244
R5028 GND.n2438 GND.n2437 240.244
R5029 GND.n2437 GND.n2019 240.244
R5030 GND.n2019 GND.n2010 240.244
R5031 GND.n2464 GND.n2010 240.244
R5032 GND.n2467 GND.n2464 240.244
R5033 GND.n2467 GND.n2465 240.244
R5034 GND.n2465 GND.n1979 240.244
R5035 GND.n2498 GND.n1979 240.244
R5036 GND.n2500 GND.n2498 240.244
R5037 GND.n2500 GND.n1966 240.244
R5038 GND.n2512 GND.n1966 240.244
R5039 GND.n2513 GND.n2512 240.244
R5040 GND.n2516 GND.n2513 240.244
R5041 GND.n2516 GND.n1383 240.244
R5042 GND.n7374 GND.n1034 240.244
R5043 GND.n7378 GND.n1034 240.244
R5044 GND.n7378 GND.n1030 240.244
R5045 GND.n7384 GND.n1030 240.244
R5046 GND.n7384 GND.n1028 240.244
R5047 GND.n7388 GND.n1028 240.244
R5048 GND.n7388 GND.n1024 240.244
R5049 GND.n7394 GND.n1024 240.244
R5050 GND.n7394 GND.n1022 240.244
R5051 GND.n7398 GND.n1022 240.244
R5052 GND.n7398 GND.n1018 240.244
R5053 GND.n7404 GND.n1018 240.244
R5054 GND.n7404 GND.n1016 240.244
R5055 GND.n7408 GND.n1016 240.244
R5056 GND.n7408 GND.n1012 240.244
R5057 GND.n7414 GND.n1012 240.244
R5058 GND.n7414 GND.n1010 240.244
R5059 GND.n7418 GND.n1010 240.244
R5060 GND.n7418 GND.n1006 240.244
R5061 GND.n7424 GND.n1006 240.244
R5062 GND.n7424 GND.n1004 240.244
R5063 GND.n7428 GND.n1004 240.244
R5064 GND.n7428 GND.n1000 240.244
R5065 GND.n7434 GND.n1000 240.244
R5066 GND.n7434 GND.n998 240.244
R5067 GND.n7438 GND.n998 240.244
R5068 GND.n7438 GND.n994 240.244
R5069 GND.n7444 GND.n994 240.244
R5070 GND.n7444 GND.n992 240.244
R5071 GND.n7448 GND.n992 240.244
R5072 GND.n7448 GND.n988 240.244
R5073 GND.n7454 GND.n988 240.244
R5074 GND.n7454 GND.n986 240.244
R5075 GND.n7458 GND.n986 240.244
R5076 GND.n7458 GND.n982 240.244
R5077 GND.n7464 GND.n982 240.244
R5078 GND.n7464 GND.n980 240.244
R5079 GND.n7468 GND.n980 240.244
R5080 GND.n7468 GND.n976 240.244
R5081 GND.n7474 GND.n976 240.244
R5082 GND.n7474 GND.n974 240.244
R5083 GND.n7478 GND.n974 240.244
R5084 GND.n7478 GND.n970 240.244
R5085 GND.n7484 GND.n970 240.244
R5086 GND.n7484 GND.n968 240.244
R5087 GND.n7488 GND.n968 240.244
R5088 GND.n7488 GND.n964 240.244
R5089 GND.n7494 GND.n964 240.244
R5090 GND.n7494 GND.n962 240.244
R5091 GND.n7498 GND.n962 240.244
R5092 GND.n7498 GND.n958 240.244
R5093 GND.n7504 GND.n958 240.244
R5094 GND.n7504 GND.n956 240.244
R5095 GND.n7508 GND.n956 240.244
R5096 GND.n7508 GND.n952 240.244
R5097 GND.n7514 GND.n952 240.244
R5098 GND.n7514 GND.n950 240.244
R5099 GND.n7518 GND.n950 240.244
R5100 GND.n7518 GND.n946 240.244
R5101 GND.n7524 GND.n946 240.244
R5102 GND.n7524 GND.n944 240.244
R5103 GND.n7528 GND.n944 240.244
R5104 GND.n7528 GND.n940 240.244
R5105 GND.n7534 GND.n940 240.244
R5106 GND.n7534 GND.n938 240.244
R5107 GND.n7538 GND.n938 240.244
R5108 GND.n7538 GND.n934 240.244
R5109 GND.n7544 GND.n934 240.244
R5110 GND.n7544 GND.n932 240.244
R5111 GND.n7548 GND.n932 240.244
R5112 GND.n7548 GND.n928 240.244
R5113 GND.n7554 GND.n928 240.244
R5114 GND.n7554 GND.n926 240.244
R5115 GND.n7558 GND.n926 240.244
R5116 GND.n7558 GND.n922 240.244
R5117 GND.n7564 GND.n922 240.244
R5118 GND.n7564 GND.n920 240.244
R5119 GND.n7568 GND.n920 240.244
R5120 GND.n7568 GND.n916 240.244
R5121 GND.n7574 GND.n916 240.244
R5122 GND.n7574 GND.n914 240.244
R5123 GND.n7578 GND.n914 240.244
R5124 GND.n7578 GND.n910 240.244
R5125 GND.n7584 GND.n910 240.244
R5126 GND.n7584 GND.n908 240.244
R5127 GND.n7588 GND.n908 240.244
R5128 GND.n7588 GND.n904 240.244
R5129 GND.n7594 GND.n904 240.244
R5130 GND.n7594 GND.n902 240.244
R5131 GND.n7598 GND.n902 240.244
R5132 GND.n7598 GND.n898 240.244
R5133 GND.n7604 GND.n898 240.244
R5134 GND.n7604 GND.n896 240.244
R5135 GND.n7608 GND.n896 240.244
R5136 GND.n7608 GND.n892 240.244
R5137 GND.n7614 GND.n892 240.244
R5138 GND.n7614 GND.n890 240.244
R5139 GND.n7618 GND.n890 240.244
R5140 GND.n7618 GND.n886 240.244
R5141 GND.n7624 GND.n886 240.244
R5142 GND.n7624 GND.n884 240.244
R5143 GND.n7628 GND.n884 240.244
R5144 GND.n7628 GND.n880 240.244
R5145 GND.n7634 GND.n880 240.244
R5146 GND.n7634 GND.n878 240.244
R5147 GND.n7638 GND.n878 240.244
R5148 GND.n7638 GND.n874 240.244
R5149 GND.n7644 GND.n874 240.244
R5150 GND.n7644 GND.n872 240.244
R5151 GND.n7648 GND.n872 240.244
R5152 GND.n7648 GND.n868 240.244
R5153 GND.n7654 GND.n868 240.244
R5154 GND.n7654 GND.n866 240.244
R5155 GND.n7658 GND.n866 240.244
R5156 GND.n7658 GND.n862 240.244
R5157 GND.n7664 GND.n862 240.244
R5158 GND.n7664 GND.n860 240.244
R5159 GND.n7668 GND.n860 240.244
R5160 GND.n7668 GND.n856 240.244
R5161 GND.n7674 GND.n856 240.244
R5162 GND.n7674 GND.n854 240.244
R5163 GND.n7678 GND.n854 240.244
R5164 GND.n7678 GND.n850 240.244
R5165 GND.n7684 GND.n850 240.244
R5166 GND.n7684 GND.n848 240.244
R5167 GND.n7688 GND.n848 240.244
R5168 GND.n7688 GND.n844 240.244
R5169 GND.n7694 GND.n844 240.244
R5170 GND.n7694 GND.n842 240.244
R5171 GND.n7698 GND.n842 240.244
R5172 GND.n7698 GND.n838 240.244
R5173 GND.n7704 GND.n838 240.244
R5174 GND.n7704 GND.n836 240.244
R5175 GND.n7708 GND.n836 240.244
R5176 GND.n7708 GND.n832 240.244
R5177 GND.n7714 GND.n832 240.244
R5178 GND.n7714 GND.n830 240.244
R5179 GND.n7718 GND.n830 240.244
R5180 GND.n7718 GND.n826 240.244
R5181 GND.n7724 GND.n826 240.244
R5182 GND.n7724 GND.n824 240.244
R5183 GND.n7728 GND.n824 240.244
R5184 GND.n7728 GND.n820 240.244
R5185 GND.n7734 GND.n820 240.244
R5186 GND.n7734 GND.n818 240.244
R5187 GND.n7738 GND.n818 240.244
R5188 GND.n7738 GND.n814 240.244
R5189 GND.n7744 GND.n814 240.244
R5190 GND.n7744 GND.n812 240.244
R5191 GND.n7748 GND.n812 240.244
R5192 GND.n7748 GND.n808 240.244
R5193 GND.n7754 GND.n808 240.244
R5194 GND.n7754 GND.n806 240.244
R5195 GND.n7758 GND.n806 240.244
R5196 GND.n7758 GND.n802 240.244
R5197 GND.n7764 GND.n802 240.244
R5198 GND.n7764 GND.n800 240.244
R5199 GND.n7768 GND.n800 240.244
R5200 GND.n7768 GND.n796 240.244
R5201 GND.n7774 GND.n796 240.244
R5202 GND.n7774 GND.n794 240.244
R5203 GND.n7778 GND.n794 240.244
R5204 GND.n7778 GND.n790 240.244
R5205 GND.n7784 GND.n790 240.244
R5206 GND.n7784 GND.n788 240.244
R5207 GND.n7788 GND.n788 240.244
R5208 GND.n7788 GND.n784 240.244
R5209 GND.n7794 GND.n784 240.244
R5210 GND.n7794 GND.n782 240.244
R5211 GND.n7798 GND.n782 240.244
R5212 GND.n7798 GND.n778 240.244
R5213 GND.n7804 GND.n778 240.244
R5214 GND.n7804 GND.n776 240.244
R5215 GND.n7808 GND.n776 240.244
R5216 GND.n7808 GND.n772 240.244
R5217 GND.n7814 GND.n772 240.244
R5218 GND.n7814 GND.n770 240.244
R5219 GND.n7818 GND.n770 240.244
R5220 GND.n7818 GND.n766 240.244
R5221 GND.n7824 GND.n766 240.244
R5222 GND.n7824 GND.n764 240.244
R5223 GND.n7828 GND.n764 240.244
R5224 GND.n7828 GND.n760 240.244
R5225 GND.n7834 GND.n760 240.244
R5226 GND.n7834 GND.n758 240.244
R5227 GND.n7838 GND.n758 240.244
R5228 GND.n7838 GND.n754 240.244
R5229 GND.n7844 GND.n754 240.244
R5230 GND.n7844 GND.n752 240.244
R5231 GND.n7848 GND.n752 240.244
R5232 GND.n7848 GND.n748 240.244
R5233 GND.n7854 GND.n748 240.244
R5234 GND.n7854 GND.n746 240.244
R5235 GND.n7858 GND.n746 240.244
R5236 GND.n7858 GND.n742 240.244
R5237 GND.n7864 GND.n742 240.244
R5238 GND.n7864 GND.n740 240.244
R5239 GND.n7868 GND.n740 240.244
R5240 GND.n7868 GND.n736 240.244
R5241 GND.n7874 GND.n736 240.244
R5242 GND.n7874 GND.n734 240.244
R5243 GND.n7878 GND.n734 240.244
R5244 GND.n7878 GND.n730 240.244
R5245 GND.n7884 GND.n730 240.244
R5246 GND.n7884 GND.n728 240.244
R5247 GND.n7888 GND.n728 240.244
R5248 GND.n7888 GND.n724 240.244
R5249 GND.n7894 GND.n724 240.244
R5250 GND.n7894 GND.n722 240.244
R5251 GND.n7898 GND.n722 240.244
R5252 GND.n7898 GND.n718 240.244
R5253 GND.n7904 GND.n718 240.244
R5254 GND.n7904 GND.n716 240.244
R5255 GND.n7908 GND.n716 240.244
R5256 GND.n7908 GND.n712 240.244
R5257 GND.n7914 GND.n712 240.244
R5258 GND.n7914 GND.n710 240.244
R5259 GND.n7918 GND.n710 240.244
R5260 GND.n7918 GND.n706 240.244
R5261 GND.n7924 GND.n706 240.244
R5262 GND.n7924 GND.n704 240.244
R5263 GND.n7928 GND.n704 240.244
R5264 GND.n7928 GND.n700 240.244
R5265 GND.n7934 GND.n700 240.244
R5266 GND.n7934 GND.n698 240.244
R5267 GND.n7938 GND.n698 240.244
R5268 GND.n7938 GND.n694 240.244
R5269 GND.n7944 GND.n694 240.244
R5270 GND.n7944 GND.n692 240.244
R5271 GND.n7948 GND.n692 240.244
R5272 GND.n7948 GND.n688 240.244
R5273 GND.n7954 GND.n688 240.244
R5274 GND.n7954 GND.n686 240.244
R5275 GND.n7958 GND.n686 240.244
R5276 GND.n7958 GND.n682 240.244
R5277 GND.n7964 GND.n682 240.244
R5278 GND.n7964 GND.n680 240.244
R5279 GND.n7968 GND.n680 240.244
R5280 GND.n7968 GND.n676 240.244
R5281 GND.n7974 GND.n676 240.244
R5282 GND.n7974 GND.n674 240.244
R5283 GND.n7978 GND.n674 240.244
R5284 GND.n7978 GND.n670 240.244
R5285 GND.n7984 GND.n670 240.244
R5286 GND.n7984 GND.n668 240.244
R5287 GND.n7988 GND.n668 240.244
R5288 GND.n7988 GND.n664 240.244
R5289 GND.n7994 GND.n664 240.244
R5290 GND.n7994 GND.n662 240.244
R5291 GND.n7998 GND.n662 240.244
R5292 GND.n7998 GND.n658 240.244
R5293 GND.n8004 GND.n658 240.244
R5294 GND.n8004 GND.n656 240.244
R5295 GND.n8008 GND.n656 240.244
R5296 GND.n8008 GND.n652 240.244
R5297 GND.n8014 GND.n652 240.244
R5298 GND.n8014 GND.n650 240.244
R5299 GND.n8018 GND.n650 240.244
R5300 GND.n8018 GND.n646 240.244
R5301 GND.n8024 GND.n646 240.244
R5302 GND.n8024 GND.n644 240.244
R5303 GND.n8028 GND.n644 240.244
R5304 GND.n8028 GND.n640 240.244
R5305 GND.n8034 GND.n640 240.244
R5306 GND.n8034 GND.n638 240.244
R5307 GND.n8038 GND.n638 240.244
R5308 GND.n8038 GND.n634 240.244
R5309 GND.n8044 GND.n634 240.244
R5310 GND.n8044 GND.n632 240.244
R5311 GND.n8048 GND.n632 240.244
R5312 GND.n8048 GND.n628 240.244
R5313 GND.n8054 GND.n628 240.244
R5314 GND.n8054 GND.n626 240.244
R5315 GND.n8058 GND.n626 240.244
R5316 GND.n8058 GND.n622 240.244
R5317 GND.n8064 GND.n622 240.244
R5318 GND.n8064 GND.n620 240.244
R5319 GND.n8068 GND.n620 240.244
R5320 GND.n8068 GND.n616 240.244
R5321 GND.n8074 GND.n616 240.244
R5322 GND.n8074 GND.n614 240.244
R5323 GND.n8078 GND.n614 240.244
R5324 GND.n8078 GND.n610 240.244
R5325 GND.n8084 GND.n610 240.244
R5326 GND.n8084 GND.n608 240.244
R5327 GND.n8088 GND.n608 240.244
R5328 GND.n8088 GND.n604 240.244
R5329 GND.n8094 GND.n604 240.244
R5330 GND.n8094 GND.n602 240.244
R5331 GND.n8098 GND.n602 240.244
R5332 GND.n8098 GND.n598 240.244
R5333 GND.n8104 GND.n598 240.244
R5334 GND.n8104 GND.n596 240.244
R5335 GND.n8108 GND.n596 240.244
R5336 GND.n8108 GND.n592 240.244
R5337 GND.n8114 GND.n592 240.244
R5338 GND.n8114 GND.n590 240.244
R5339 GND.n8118 GND.n590 240.244
R5340 GND.n8118 GND.n586 240.244
R5341 GND.n8124 GND.n586 240.244
R5342 GND.n8124 GND.n584 240.244
R5343 GND.n8128 GND.n584 240.244
R5344 GND.n8128 GND.n580 240.244
R5345 GND.n8134 GND.n580 240.244
R5346 GND.n8134 GND.n578 240.244
R5347 GND.n8138 GND.n578 240.244
R5348 GND.n8138 GND.n574 240.244
R5349 GND.n8144 GND.n574 240.244
R5350 GND.n8144 GND.n572 240.244
R5351 GND.n8148 GND.n572 240.244
R5352 GND.n8148 GND.n568 240.244
R5353 GND.n8154 GND.n568 240.244
R5354 GND.n8154 GND.n566 240.244
R5355 GND.n8158 GND.n566 240.244
R5356 GND.n8158 GND.n562 240.244
R5357 GND.n8164 GND.n562 240.244
R5358 GND.n8164 GND.n560 240.244
R5359 GND.n8168 GND.n560 240.244
R5360 GND.n8168 GND.n556 240.244
R5361 GND.n8174 GND.n556 240.244
R5362 GND.n8174 GND.n554 240.244
R5363 GND.n8178 GND.n554 240.244
R5364 GND.n8178 GND.n550 240.244
R5365 GND.n8184 GND.n550 240.244
R5366 GND.n8184 GND.n548 240.244
R5367 GND.n8188 GND.n548 240.244
R5368 GND.n8188 GND.n544 240.244
R5369 GND.n8194 GND.n544 240.244
R5370 GND.n8194 GND.n542 240.244
R5371 GND.n8198 GND.n542 240.244
R5372 GND.n8198 GND.n538 240.244
R5373 GND.n8205 GND.n538 240.244
R5374 GND.n8205 GND.n536 240.244
R5375 GND.n8209 GND.n536 240.244
R5376 GND.n8209 GND.n533 240.244
R5377 GND.n8215 GND.n531 240.244
R5378 GND.n8219 GND.n531 240.244
R5379 GND.n8219 GND.n527 240.244
R5380 GND.n8225 GND.n527 240.244
R5381 GND.n8225 GND.n525 240.244
R5382 GND.n8229 GND.n525 240.244
R5383 GND.n8229 GND.n521 240.244
R5384 GND.n8235 GND.n521 240.244
R5385 GND.n8235 GND.n519 240.244
R5386 GND.n8239 GND.n519 240.244
R5387 GND.n8239 GND.n515 240.244
R5388 GND.n8245 GND.n515 240.244
R5389 GND.n8245 GND.n513 240.244
R5390 GND.n8249 GND.n513 240.244
R5391 GND.n8249 GND.n509 240.244
R5392 GND.n8255 GND.n509 240.244
R5393 GND.n8255 GND.n507 240.244
R5394 GND.n8259 GND.n507 240.244
R5395 GND.n8259 GND.n503 240.244
R5396 GND.n8265 GND.n503 240.244
R5397 GND.n8265 GND.n501 240.244
R5398 GND.n8269 GND.n501 240.244
R5399 GND.n8269 GND.n497 240.244
R5400 GND.n8275 GND.n497 240.244
R5401 GND.n8275 GND.n495 240.244
R5402 GND.n8279 GND.n495 240.244
R5403 GND.n8279 GND.n491 240.244
R5404 GND.n8285 GND.n491 240.244
R5405 GND.n8285 GND.n489 240.244
R5406 GND.n8289 GND.n489 240.244
R5407 GND.n8289 GND.n485 240.244
R5408 GND.n8295 GND.n485 240.244
R5409 GND.n8295 GND.n483 240.244
R5410 GND.n8299 GND.n483 240.244
R5411 GND.n8299 GND.n479 240.244
R5412 GND.n8305 GND.n479 240.244
R5413 GND.n8305 GND.n477 240.244
R5414 GND.n8309 GND.n477 240.244
R5415 GND.n8309 GND.n473 240.244
R5416 GND.n8315 GND.n473 240.244
R5417 GND.n8315 GND.n471 240.244
R5418 GND.n8319 GND.n471 240.244
R5419 GND.n8319 GND.n467 240.244
R5420 GND.n8325 GND.n467 240.244
R5421 GND.n8325 GND.n465 240.244
R5422 GND.n8329 GND.n465 240.244
R5423 GND.n8329 GND.n461 240.244
R5424 GND.n8335 GND.n461 240.244
R5425 GND.n8335 GND.n459 240.244
R5426 GND.n8339 GND.n459 240.244
R5427 GND.n8339 GND.n455 240.244
R5428 GND.n8345 GND.n455 240.244
R5429 GND.n8345 GND.n453 240.244
R5430 GND.n8349 GND.n453 240.244
R5431 GND.n8349 GND.n449 240.244
R5432 GND.n8355 GND.n449 240.244
R5433 GND.n8355 GND.n447 240.244
R5434 GND.n8359 GND.n447 240.244
R5435 GND.n8359 GND.n443 240.244
R5436 GND.n8365 GND.n443 240.244
R5437 GND.n8365 GND.n441 240.244
R5438 GND.n8369 GND.n441 240.244
R5439 GND.n8369 GND.n437 240.244
R5440 GND.n8375 GND.n437 240.244
R5441 GND.n8375 GND.n435 240.244
R5442 GND.n8379 GND.n435 240.244
R5443 GND.n8379 GND.n431 240.244
R5444 GND.n8385 GND.n431 240.244
R5445 GND.n8385 GND.n429 240.244
R5446 GND.n8389 GND.n429 240.244
R5447 GND.n8389 GND.n425 240.244
R5448 GND.n8396 GND.n425 240.244
R5449 GND.n7222 GND.n1182 240.244
R5450 GND.n7218 GND.n1182 240.244
R5451 GND.n7218 GND.n1184 240.244
R5452 GND.n7214 GND.n1184 240.244
R5453 GND.n7214 GND.n1189 240.244
R5454 GND.n7210 GND.n1189 240.244
R5455 GND.n7210 GND.n1191 240.244
R5456 GND.n7206 GND.n1191 240.244
R5457 GND.n7206 GND.n1197 240.244
R5458 GND.n7202 GND.n1197 240.244
R5459 GND.n7202 GND.n1199 240.244
R5460 GND.n7198 GND.n1199 240.244
R5461 GND.n7198 GND.n1205 240.244
R5462 GND.n7194 GND.n1205 240.244
R5463 GND.n7194 GND.n1207 240.244
R5464 GND.n7190 GND.n1207 240.244
R5465 GND.n7190 GND.n1213 240.244
R5466 GND.n7186 GND.n1213 240.244
R5467 GND.n7186 GND.n1215 240.244
R5468 GND.n7182 GND.n1215 240.244
R5469 GND.n7182 GND.n1221 240.244
R5470 GND.n2160 GND.n1221 240.244
R5471 GND.n2166 GND.n2160 240.244
R5472 GND.n2167 GND.n2166 240.244
R5473 GND.n2219 GND.n2167 240.244
R5474 GND.n2219 GND.n2155 240.244
R5475 GND.n2263 GND.n2155 240.244
R5476 GND.n2263 GND.n2156 240.244
R5477 GND.n2259 GND.n2156 240.244
R5478 GND.n2259 GND.n2258 240.244
R5479 GND.n2258 GND.n2257 240.244
R5480 GND.n2257 GND.n2227 240.244
R5481 GND.n2253 GND.n2227 240.244
R5482 GND.n2253 GND.n2252 240.244
R5483 GND.n2252 GND.n2251 240.244
R5484 GND.n2251 GND.n2233 240.244
R5485 GND.n2247 GND.n2233 240.244
R5486 GND.n2247 GND.n2246 240.244
R5487 GND.n2246 GND.n2245 240.244
R5488 GND.n2245 GND.n2239 240.244
R5489 GND.n2239 GND.n2065 240.244
R5490 GND.n2409 GND.n2065 240.244
R5491 GND.n2409 GND.n2066 240.244
R5492 GND.n2404 GND.n2066 240.244
R5493 GND.n2404 GND.n2069 240.244
R5494 GND.n2351 GND.n2069 240.244
R5495 GND.n2391 GND.n2351 240.244
R5496 GND.n2391 GND.n2355 240.244
R5497 GND.n2386 GND.n2355 240.244
R5498 GND.n2386 GND.n2385 240.244
R5499 GND.n2385 GND.n2384 240.244
R5500 GND.n2384 GND.n2360 240.244
R5501 GND.n2380 GND.n2360 240.244
R5502 GND.n2380 GND.n2379 240.244
R5503 GND.n2379 GND.n2378 240.244
R5504 GND.n2378 GND.n2366 240.244
R5505 GND.n2374 GND.n2366 240.244
R5506 GND.n2374 GND.n1998 240.244
R5507 GND.n2478 GND.n1998 240.244
R5508 GND.n2479 GND.n2478 240.244
R5509 GND.n2480 GND.n2479 240.244
R5510 GND.n2480 GND.n1994 240.244
R5511 GND.n2489 GND.n1994 240.244
R5512 GND.n2489 GND.n1962 240.244
R5513 GND.n2519 GND.n1962 240.244
R5514 GND.n2520 GND.n2519 240.244
R5515 GND.n2521 GND.n2520 240.244
R5516 GND.n2521 GND.n1957 240.244
R5517 GND.n6971 GND.n1957 240.244
R5518 GND.n6971 GND.n1958 240.244
R5519 GND.n6967 GND.n1958 240.244
R5520 GND.n6967 GND.n2529 240.244
R5521 GND.n6963 GND.n2529 240.244
R5522 GND.n6963 GND.n2531 240.244
R5523 GND.n6959 GND.n2531 240.244
R5524 GND.n6959 GND.n2537 240.244
R5525 GND.n6949 GND.n2537 240.244
R5526 GND.n6949 GND.n2549 240.244
R5527 GND.n6945 GND.n2549 240.244
R5528 GND.n6945 GND.n2555 240.244
R5529 GND.n6936 GND.n2555 240.244
R5530 GND.n6936 GND.n2567 240.244
R5531 GND.n6932 GND.n2567 240.244
R5532 GND.n6932 GND.n2573 240.244
R5533 GND.n6922 GND.n2573 240.244
R5534 GND.n6922 GND.n2584 240.244
R5535 GND.n6918 GND.n2584 240.244
R5536 GND.n6918 GND.n2590 240.244
R5537 GND.n6908 GND.n2590 240.244
R5538 GND.n6908 GND.n2602 240.244
R5539 GND.n6904 GND.n2602 240.244
R5540 GND.n6904 GND.n2608 240.244
R5541 GND.n6894 GND.n2608 240.244
R5542 GND.n6894 GND.n2620 240.244
R5543 GND.n6890 GND.n2620 240.244
R5544 GND.n6890 GND.n2626 240.244
R5545 GND.n6880 GND.n2626 240.244
R5546 GND.n6880 GND.n2638 240.244
R5547 GND.n6876 GND.n2638 240.244
R5548 GND.n6876 GND.n2644 240.244
R5549 GND.n6866 GND.n2644 240.244
R5550 GND.n6866 GND.n2655 240.244
R5551 GND.n6862 GND.n2655 240.244
R5552 GND.n6862 GND.n2661 240.244
R5553 GND.n4350 GND.n2661 240.244
R5554 GND.n4350 GND.n3886 240.244
R5555 GND.n4356 GND.n3886 240.244
R5556 GND.n4356 GND.n3873 240.244
R5557 GND.n4388 GND.n3873 240.244
R5558 GND.n4388 GND.n3868 240.244
R5559 GND.n4407 GND.n3868 240.244
R5560 GND.n4407 GND.n3869 240.244
R5561 GND.n4403 GND.n3869 240.244
R5562 GND.n4403 GND.n4402 240.244
R5563 GND.n4402 GND.n4401 240.244
R5564 GND.n4401 GND.n3833 240.244
R5565 GND.n4477 GND.n3833 240.244
R5566 GND.n4477 GND.n3828 240.244
R5567 GND.n4485 GND.n3828 240.244
R5568 GND.n4485 GND.n3829 240.244
R5569 GND.n3829 GND.n3802 240.244
R5570 GND.n4523 GND.n3802 240.244
R5571 GND.n4523 GND.n3798 240.244
R5572 GND.n4529 GND.n3798 240.244
R5573 GND.n4529 GND.n3784 240.244
R5574 GND.n4580 GND.n3784 240.244
R5575 GND.n4580 GND.n3780 240.244
R5576 GND.n4586 GND.n3780 240.244
R5577 GND.n4586 GND.n3761 240.244
R5578 GND.n4608 GND.n3761 240.244
R5579 GND.n4608 GND.n3756 240.244
R5580 GND.n4616 GND.n3756 240.244
R5581 GND.n4616 GND.n3757 240.244
R5582 GND.n3757 GND.n3732 240.244
R5583 GND.n4680 GND.n3732 240.244
R5584 GND.n4680 GND.n3728 240.244
R5585 GND.n4686 GND.n3728 240.244
R5586 GND.n4686 GND.n3711 240.244
R5587 GND.n4706 GND.n3711 240.244
R5588 GND.n4706 GND.n3707 240.244
R5589 GND.n4712 GND.n3707 240.244
R5590 GND.n4712 GND.n3690 240.244
R5591 GND.n4741 GND.n3690 240.244
R5592 GND.n4741 GND.n3686 240.244
R5593 GND.n4747 GND.n3686 240.244
R5594 GND.n4747 GND.n3673 240.244
R5595 GND.n4784 GND.n3673 240.244
R5596 GND.n4784 GND.n3668 240.244
R5597 GND.n4792 GND.n3668 240.244
R5598 GND.n4792 GND.n3669 240.244
R5599 GND.n3669 GND.n3644 240.244
R5600 GND.n4857 GND.n3644 240.244
R5601 GND.n4857 GND.n3640 240.244
R5602 GND.n4863 GND.n3640 240.244
R5603 GND.n4863 GND.n3624 240.244
R5604 GND.n4884 GND.n3624 240.244
R5605 GND.n4884 GND.n3620 240.244
R5606 GND.n4890 GND.n3620 240.244
R5607 GND.n4890 GND.n3602 240.244
R5608 GND.n4918 GND.n3602 240.244
R5609 GND.n4918 GND.n3598 240.244
R5610 GND.n4924 GND.n3598 240.244
R5611 GND.n4924 GND.n3585 240.244
R5612 GND.n4961 GND.n3585 240.244
R5613 GND.n4961 GND.n3580 240.244
R5614 GND.n4969 GND.n3580 240.244
R5615 GND.n4969 GND.n3581 240.244
R5616 GND.n3581 GND.n3556 240.244
R5617 GND.n5033 GND.n3556 240.244
R5618 GND.n5033 GND.n3552 240.244
R5619 GND.n5039 GND.n3552 240.244
R5620 GND.n5039 GND.n3535 240.244
R5621 GND.n5059 GND.n3535 240.244
R5622 GND.n5059 GND.n3531 240.244
R5623 GND.n5065 GND.n3531 240.244
R5624 GND.n5065 GND.n3513 240.244
R5625 GND.n5093 GND.n3513 240.244
R5626 GND.n5093 GND.n3509 240.244
R5627 GND.n5099 GND.n3509 240.244
R5628 GND.n5099 GND.n3496 240.244
R5629 GND.n5137 GND.n3496 240.244
R5630 GND.n5137 GND.n3491 240.244
R5631 GND.n5145 GND.n3491 240.244
R5632 GND.n5145 GND.n3492 240.244
R5633 GND.n3492 GND.n3467 240.244
R5634 GND.n5208 GND.n3467 240.244
R5635 GND.n5208 GND.n3463 240.244
R5636 GND.n5214 GND.n3463 240.244
R5637 GND.n5214 GND.n3446 240.244
R5638 GND.n5234 GND.n3446 240.244
R5639 GND.n5234 GND.n3442 240.244
R5640 GND.n5240 GND.n3442 240.244
R5641 GND.n5240 GND.n3424 240.244
R5642 GND.n5268 GND.n3424 240.244
R5643 GND.n5268 GND.n3420 240.244
R5644 GND.n5274 GND.n3420 240.244
R5645 GND.n5274 GND.n3407 240.244
R5646 GND.n5311 GND.n3407 240.244
R5647 GND.n5311 GND.n3402 240.244
R5648 GND.n5319 GND.n3402 240.244
R5649 GND.n5319 GND.n3403 240.244
R5650 GND.n3403 GND.n3378 240.244
R5651 GND.n5385 GND.n3378 240.244
R5652 GND.n5385 GND.n3374 240.244
R5653 GND.n5391 GND.n3374 240.244
R5654 GND.n5391 GND.n3359 240.244
R5655 GND.n5411 GND.n3359 240.244
R5656 GND.n5411 GND.n3355 240.244
R5657 GND.n5417 GND.n3355 240.244
R5658 GND.n5417 GND.n3338 240.244
R5659 GND.n5446 GND.n3338 240.244
R5660 GND.n5446 GND.n3334 240.244
R5661 GND.n5452 GND.n3334 240.244
R5662 GND.n5452 GND.n3321 240.244
R5663 GND.n5489 GND.n3321 240.244
R5664 GND.n5489 GND.n3316 240.244
R5665 GND.n5497 GND.n3316 240.244
R5666 GND.n5497 GND.n3317 240.244
R5667 GND.n3317 GND.n3292 240.244
R5668 GND.n5539 GND.n3292 240.244
R5669 GND.n5539 GND.n3288 240.244
R5670 GND.n5547 GND.n3288 240.244
R5671 GND.n5547 GND.n3272 240.244
R5672 GND.n5566 GND.n3272 240.244
R5673 GND.n5567 GND.n5566 240.244
R5674 GND.n5567 GND.n3267 240.244
R5675 GND.n5584 GND.n3267 240.244
R5676 GND.n5584 GND.n3268 240.244
R5677 GND.n5580 GND.n3268 240.244
R5678 GND.n5580 GND.n5579 240.244
R5679 GND.n5579 GND.n2906 240.244
R5680 GND.n6624 GND.n2906 240.244
R5681 GND.n6624 GND.n2907 240.244
R5682 GND.n6620 GND.n2907 240.244
R5683 GND.n6620 GND.n2913 240.244
R5684 GND.n6610 GND.n2913 240.244
R5685 GND.n6610 GND.n2924 240.244
R5686 GND.n6606 GND.n2924 240.244
R5687 GND.n6606 GND.n2930 240.244
R5688 GND.n6596 GND.n2930 240.244
R5689 GND.n6596 GND.n2942 240.244
R5690 GND.n6592 GND.n2942 240.244
R5691 GND.n6592 GND.n2948 240.244
R5692 GND.n6582 GND.n2948 240.244
R5693 GND.n6582 GND.n2960 240.244
R5694 GND.n6578 GND.n2960 240.244
R5695 GND.n6578 GND.n2966 240.244
R5696 GND.n6568 GND.n2966 240.244
R5697 GND.n6568 GND.n2978 240.244
R5698 GND.n6564 GND.n2978 240.244
R5699 GND.n6564 GND.n2984 240.244
R5700 GND.n6554 GND.n2984 240.244
R5701 GND.n6554 GND.n2995 240.244
R5702 GND.n6550 GND.n2995 240.244
R5703 GND.n6550 GND.n3001 240.244
R5704 GND.n6540 GND.n3001 240.244
R5705 GND.n6540 GND.n3013 240.244
R5706 GND.n6536 GND.n3013 240.244
R5707 GND.n6536 GND.n3019 240.244
R5708 GND.n6526 GND.n3019 240.244
R5709 GND.n6526 GND.n3030 240.244
R5710 GND.n6522 GND.n3030 240.244
R5711 GND.n6522 GND.n3036 240.244
R5712 GND.n6518 GND.n3036 240.244
R5713 GND.n6518 GND.n3039 240.244
R5714 GND.n6514 GND.n3039 240.244
R5715 GND.n6514 GND.n3045 240.244
R5716 GND.n5994 GND.n3045 240.244
R5717 GND.n6000 GND.n5994 240.244
R5718 GND.n6001 GND.n6000 240.244
R5719 GND.n6002 GND.n6001 240.244
R5720 GND.n6002 GND.n5990 240.244
R5721 GND.n6008 GND.n5990 240.244
R5722 GND.n6009 GND.n6008 240.244
R5723 GND.n6010 GND.n6009 240.244
R5724 GND.n6010 GND.n5986 240.244
R5725 GND.n6016 GND.n5986 240.244
R5726 GND.n6017 GND.n6016 240.244
R5727 GND.n6018 GND.n6017 240.244
R5728 GND.n6018 GND.n5982 240.244
R5729 GND.n6024 GND.n5982 240.244
R5730 GND.n6025 GND.n6024 240.244
R5731 GND.n6026 GND.n6025 240.244
R5732 GND.n6026 GND.n5977 240.244
R5733 GND.n6034 GND.n5977 240.244
R5734 GND.n6034 GND.n5978 240.244
R5735 GND.n5978 GND.n5927 240.244
R5736 GND.n6386 GND.n5927 240.244
R5737 GND.n6386 GND.n5928 240.244
R5738 GND.n6381 GND.n5928 240.244
R5739 GND.n6381 GND.n5931 240.244
R5740 GND.n6371 GND.n5931 240.244
R5741 GND.n6371 GND.n5945 240.244
R5742 GND.n6366 GND.n5945 240.244
R5743 GND.n6366 GND.n6365 240.244
R5744 GND.n6365 GND.n5948 240.244
R5745 GND.n6361 GND.n5948 240.244
R5746 GND.n6361 GND.n6360 240.244
R5747 GND.n6360 GND.n6359 240.244
R5748 GND.n6359 GND.n5952 240.244
R5749 GND.n6355 GND.n5952 240.244
R5750 GND.n6355 GND.n5958 240.244
R5751 GND.n6313 GND.n5958 240.244
R5752 GND.n6319 GND.n6313 240.244
R5753 GND.n6320 GND.n6319 240.244
R5754 GND.n6321 GND.n6320 240.244
R5755 GND.n6321 GND.n6308 240.244
R5756 GND.n6333 GND.n6308 240.244
R5757 GND.n6333 GND.n6309 240.244
R5758 GND.n6329 GND.n6309 240.244
R5759 GND.n6329 GND.n254 240.244
R5760 GND.n8444 GND.n254 240.244
R5761 GND.n8444 GND.n255 240.244
R5762 GND.n8440 GND.n255 240.244
R5763 GND.n8440 GND.n261 240.244
R5764 GND.n8436 GND.n261 240.244
R5765 GND.n8436 GND.n385 240.244
R5766 GND.n8432 GND.n385 240.244
R5767 GND.n8432 GND.n391 240.244
R5768 GND.n8428 GND.n391 240.244
R5769 GND.n8428 GND.n393 240.244
R5770 GND.n8424 GND.n393 240.244
R5771 GND.n8424 GND.n399 240.244
R5772 GND.n8420 GND.n399 240.244
R5773 GND.n8420 GND.n401 240.244
R5774 GND.n8416 GND.n401 240.244
R5775 GND.n8416 GND.n407 240.244
R5776 GND.n8412 GND.n407 240.244
R5777 GND.n8412 GND.n409 240.244
R5778 GND.n8408 GND.n409 240.244
R5779 GND.n8408 GND.n415 240.244
R5780 GND.n8404 GND.n415 240.244
R5781 GND.n8404 GND.n417 240.244
R5782 GND.n8400 GND.n417 240.244
R5783 GND.n8400 GND.n423 240.244
R5784 GND.n7368 GND.n1036 240.244
R5785 GND.n7368 GND.n1039 240.244
R5786 GND.n7364 GND.n1039 240.244
R5787 GND.n7364 GND.n1041 240.244
R5788 GND.n7360 GND.n1041 240.244
R5789 GND.n7360 GND.n1047 240.244
R5790 GND.n7356 GND.n1047 240.244
R5791 GND.n7356 GND.n1049 240.244
R5792 GND.n7352 GND.n1049 240.244
R5793 GND.n7352 GND.n1055 240.244
R5794 GND.n7348 GND.n1055 240.244
R5795 GND.n7348 GND.n1057 240.244
R5796 GND.n7344 GND.n1057 240.244
R5797 GND.n7344 GND.n1063 240.244
R5798 GND.n7340 GND.n1063 240.244
R5799 GND.n7340 GND.n1065 240.244
R5800 GND.n7336 GND.n1065 240.244
R5801 GND.n7336 GND.n1071 240.244
R5802 GND.n7332 GND.n1071 240.244
R5803 GND.n7332 GND.n1073 240.244
R5804 GND.n7328 GND.n1073 240.244
R5805 GND.n7328 GND.n1079 240.244
R5806 GND.n7324 GND.n1079 240.244
R5807 GND.n7324 GND.n1081 240.244
R5808 GND.n7320 GND.n1081 240.244
R5809 GND.n7320 GND.n1087 240.244
R5810 GND.n7316 GND.n1087 240.244
R5811 GND.n7316 GND.n1089 240.244
R5812 GND.n7312 GND.n1089 240.244
R5813 GND.n7312 GND.n1095 240.244
R5814 GND.n7308 GND.n1095 240.244
R5815 GND.n7308 GND.n1097 240.244
R5816 GND.n7304 GND.n1097 240.244
R5817 GND.n7304 GND.n1103 240.244
R5818 GND.n7300 GND.n1103 240.244
R5819 GND.n7300 GND.n1105 240.244
R5820 GND.n7296 GND.n1105 240.244
R5821 GND.n7296 GND.n1111 240.244
R5822 GND.n7292 GND.n1111 240.244
R5823 GND.n7292 GND.n1113 240.244
R5824 GND.n7288 GND.n1113 240.244
R5825 GND.n7288 GND.n1119 240.244
R5826 GND.n7284 GND.n1119 240.244
R5827 GND.n7284 GND.n1121 240.244
R5828 GND.n7280 GND.n1121 240.244
R5829 GND.n7280 GND.n1127 240.244
R5830 GND.n7276 GND.n1127 240.244
R5831 GND.n7276 GND.n1129 240.244
R5832 GND.n7272 GND.n1129 240.244
R5833 GND.n7272 GND.n1135 240.244
R5834 GND.n7268 GND.n1135 240.244
R5835 GND.n7268 GND.n1137 240.244
R5836 GND.n7264 GND.n1137 240.244
R5837 GND.n7264 GND.n1143 240.244
R5838 GND.n7260 GND.n1143 240.244
R5839 GND.n7260 GND.n1145 240.244
R5840 GND.n7256 GND.n1145 240.244
R5841 GND.n7256 GND.n1151 240.244
R5842 GND.n7252 GND.n1151 240.244
R5843 GND.n7252 GND.n1153 240.244
R5844 GND.n7248 GND.n1153 240.244
R5845 GND.n7248 GND.n1159 240.244
R5846 GND.n7244 GND.n1159 240.244
R5847 GND.n7244 GND.n1161 240.244
R5848 GND.n7240 GND.n1161 240.244
R5849 GND.n7240 GND.n1167 240.244
R5850 GND.n7236 GND.n1167 240.244
R5851 GND.n7236 GND.n1169 240.244
R5852 GND.n7232 GND.n1169 240.244
R5853 GND.n7232 GND.n1175 240.244
R5854 GND.n7228 GND.n1175 240.244
R5855 GND.n7228 GND.n1177 240.244
R5856 GND.n2831 GND.n2830 240.244
R5857 GND.n3220 GND.n2874 240.244
R5858 GND.n2876 GND.n2875 240.244
R5859 GND.n3223 GND.n2879 240.244
R5860 GND.n2881 GND.n2880 240.244
R5861 GND.n3226 GND.n2884 240.244
R5862 GND.n2886 GND.n2885 240.244
R5863 GND.n3229 GND.n2889 240.244
R5864 GND.n2891 GND.n2890 240.244
R5865 GND.n2897 GND.n2896 240.244
R5866 GND.n2903 GND.n2898 240.244
R5867 GND.n4338 GND.n2663 240.244
R5868 GND.n4338 GND.n3890 240.244
R5869 GND.n4324 GND.n3890 240.244
R5870 GND.n4325 GND.n4324 240.244
R5871 GND.n4326 GND.n4325 240.244
R5872 GND.n4327 GND.n4326 240.244
R5873 GND.n4327 GND.n3859 240.244
R5874 GND.n4418 GND.n3859 240.244
R5875 GND.n4418 GND.n3853 240.244
R5876 GND.n4434 GND.n3853 240.244
R5877 GND.n4434 GND.n3854 240.244
R5878 GND.n4423 GND.n3854 240.244
R5879 GND.n4424 GND.n4423 240.244
R5880 GND.n4425 GND.n4424 240.244
R5881 GND.n4425 GND.n3819 240.244
R5882 GND.n4495 GND.n3819 240.244
R5883 GND.n4495 GND.n3814 240.244
R5884 GND.n4511 GND.n3814 240.244
R5885 GND.n4511 GND.n3804 240.244
R5886 GND.n4500 GND.n3804 240.244
R5887 GND.n4501 GND.n4500 240.244
R5888 GND.n4502 GND.n4501 240.244
R5889 GND.n4502 GND.n3777 240.244
R5890 GND.n4589 GND.n3777 240.244
R5891 GND.n4589 GND.n3771 240.244
R5892 GND.n4596 GND.n3771 240.244
R5893 GND.n4596 GND.n3772 240.244
R5894 GND.n3772 GND.n3747 240.244
R5895 GND.n4628 GND.n3747 240.244
R5896 GND.n4628 GND.n3742 240.244
R5897 GND.n4669 GND.n3742 240.244
R5898 GND.n4669 GND.n3734 240.244
R5899 GND.n4633 GND.n3734 240.244
R5900 GND.n4634 GND.n4633 240.244
R5901 GND.n4635 GND.n4634 240.244
R5902 GND.n4635 GND.n3713 240.244
R5903 GND.n3713 GND.n3705 240.244
R5904 GND.n4638 GND.n3705 240.244
R5905 GND.n4639 GND.n4638 240.244
R5906 GND.n4642 GND.n4639 240.244
R5907 GND.n4643 GND.n4642 240.244
R5908 GND.n4644 GND.n4643 240.244
R5909 GND.n4645 GND.n4644 240.244
R5910 GND.n4646 GND.n4645 240.244
R5911 GND.n4646 GND.n3659 240.244
R5912 GND.n4804 GND.n3659 240.244
R5913 GND.n4804 GND.n3654 240.244
R5914 GND.n4845 GND.n3654 240.244
R5915 GND.n4845 GND.n3646 240.244
R5916 GND.n4809 GND.n3646 240.244
R5917 GND.n4810 GND.n4809 240.244
R5918 GND.n4811 GND.n4810 240.244
R5919 GND.n4811 GND.n3626 240.244
R5920 GND.n3626 GND.n3618 240.244
R5921 GND.n4814 GND.n3618 240.244
R5922 GND.n4815 GND.n4814 240.244
R5923 GND.n4818 GND.n4815 240.244
R5924 GND.n4819 GND.n4818 240.244
R5925 GND.n4820 GND.n4819 240.244
R5926 GND.n4821 GND.n4820 240.244
R5927 GND.n4822 GND.n4821 240.244
R5928 GND.n4822 GND.n3571 240.244
R5929 GND.n4980 GND.n3571 240.244
R5930 GND.n4980 GND.n3566 240.244
R5931 GND.n5021 GND.n3566 240.244
R5932 GND.n5021 GND.n3558 240.244
R5933 GND.n4985 GND.n3558 240.244
R5934 GND.n4986 GND.n4985 240.244
R5935 GND.n4987 GND.n4986 240.244
R5936 GND.n4987 GND.n3537 240.244
R5937 GND.n3537 GND.n3529 240.244
R5938 GND.n4990 GND.n3529 240.244
R5939 GND.n4991 GND.n4990 240.244
R5940 GND.n4994 GND.n4991 240.244
R5941 GND.n4995 GND.n4994 240.244
R5942 GND.n4996 GND.n4995 240.244
R5943 GND.n4997 GND.n4996 240.244
R5944 GND.n4998 GND.n4997 240.244
R5945 GND.n4998 GND.n3482 240.244
R5946 GND.n5156 GND.n3482 240.244
R5947 GND.n5156 GND.n3477 240.244
R5948 GND.n5197 GND.n3477 240.244
R5949 GND.n5197 GND.n3469 240.244
R5950 GND.n5161 GND.n3469 240.244
R5951 GND.n5162 GND.n5161 240.244
R5952 GND.n5163 GND.n5162 240.244
R5953 GND.n5163 GND.n3448 240.244
R5954 GND.n3448 GND.n3440 240.244
R5955 GND.n5166 GND.n3440 240.244
R5956 GND.n5167 GND.n5166 240.244
R5957 GND.n5170 GND.n5167 240.244
R5958 GND.n5171 GND.n5170 240.244
R5959 GND.n5172 GND.n5171 240.244
R5960 GND.n5173 GND.n5172 240.244
R5961 GND.n5174 GND.n5173 240.244
R5962 GND.n5174 GND.n3393 240.244
R5963 GND.n5331 GND.n3393 240.244
R5964 GND.n5331 GND.n3388 240.244
R5965 GND.n5374 GND.n3388 240.244
R5966 GND.n5374 GND.n3380 240.244
R5967 GND.n5336 GND.n3380 240.244
R5968 GND.n5339 GND.n5336 240.244
R5969 GND.n5340 GND.n5339 240.244
R5970 GND.n5340 GND.n3361 240.244
R5971 GND.n3361 GND.n3353 240.244
R5972 GND.n5343 GND.n3353 240.244
R5973 GND.n5344 GND.n5343 240.244
R5974 GND.n5347 GND.n5344 240.244
R5975 GND.n5348 GND.n5347 240.244
R5976 GND.n5349 GND.n5348 240.244
R5977 GND.n5350 GND.n5349 240.244
R5978 GND.n5351 GND.n5350 240.244
R5979 GND.n5351 GND.n3307 240.244
R5980 GND.n5509 GND.n3307 240.244
R5981 GND.n5509 GND.n3302 240.244
R5982 GND.n5527 GND.n3302 240.244
R5983 GND.n5527 GND.n3294 240.244
R5984 GND.n5514 GND.n3294 240.244
R5985 GND.n5515 GND.n5514 240.244
R5986 GND.n5516 GND.n5515 240.244
R5987 GND.n5516 GND.n3274 240.244
R5988 GND.n3274 GND.n3257 240.244
R5989 GND.n5603 GND.n3257 240.244
R5990 GND.n5603 GND.n3251 240.244
R5991 GND.n5610 GND.n3251 240.244
R5992 GND.n5610 GND.n3252 240.244
R5993 GND.n3252 GND.n2902 240.244
R5994 GND.n6627 GND.n2902 240.244
R5995 GND.n4315 GND.n4212 240.244
R5996 GND.n4216 GND.n4212 240.244
R5997 GND.n4218 GND.n4217 240.244
R5998 GND.n4222 GND.n4221 240.244
R5999 GND.n4224 GND.n4223 240.244
R6000 GND.n4228 GND.n4227 240.244
R6001 GND.n4230 GND.n4229 240.244
R6002 GND.n4234 GND.n4233 240.244
R6003 GND.n4236 GND.n4235 240.244
R6004 GND.n4243 GND.n4242 240.244
R6005 GND.n4244 GND.n3904 240.244
R6006 GND.n6859 GND.n2666 240.244
R6007 GND.n2670 GND.n2666 240.244
R6008 GND.n2671 GND.n2670 240.244
R6009 GND.n2672 GND.n2671 240.244
R6010 GND.n3874 GND.n2672 240.244
R6011 GND.n3874 GND.n2675 240.244
R6012 GND.n2676 GND.n2675 240.244
R6013 GND.n2677 GND.n2676 240.244
R6014 GND.n4363 GND.n2677 240.244
R6015 GND.n4363 GND.n2680 240.244
R6016 GND.n2681 GND.n2680 240.244
R6017 GND.n2682 GND.n2681 240.244
R6018 GND.n3834 GND.n2682 240.244
R6019 GND.n3834 GND.n2685 240.244
R6020 GND.n2686 GND.n2685 240.244
R6021 GND.n2687 GND.n2686 240.244
R6022 GND.n4451 GND.n2687 240.244
R6023 GND.n4451 GND.n2690 240.244
R6024 GND.n2691 GND.n2690 240.244
R6025 GND.n2692 GND.n2691 240.244
R6026 GND.n3792 GND.n2692 240.244
R6027 GND.n3792 GND.n2695 240.244
R6028 GND.n2696 GND.n2695 240.244
R6029 GND.n2697 GND.n2696 240.244
R6030 GND.n3767 GND.n2697 240.244
R6031 GND.n3767 GND.n2700 240.244
R6032 GND.n2701 GND.n2700 240.244
R6033 GND.n2702 GND.n2701 240.244
R6034 GND.n4626 GND.n2702 240.244
R6035 GND.n4626 GND.n2705 240.244
R6036 GND.n2706 GND.n2705 240.244
R6037 GND.n2707 GND.n2706 240.244
R6038 GND.n3723 GND.n2707 240.244
R6039 GND.n3723 GND.n2710 240.244
R6040 GND.n2711 GND.n2710 240.244
R6041 GND.n2712 GND.n2711 240.244
R6042 GND.n4715 GND.n2712 240.244
R6043 GND.n4715 GND.n2715 240.244
R6044 GND.n2716 GND.n2715 240.244
R6045 GND.n2717 GND.n2716 240.244
R6046 GND.n3684 GND.n2717 240.244
R6047 GND.n3684 GND.n2720 240.244
R6048 GND.n2721 GND.n2720 240.244
R6049 GND.n2722 GND.n2721 240.244
R6050 GND.n4794 GND.n2722 240.244
R6051 GND.n4794 GND.n2725 240.244
R6052 GND.n2726 GND.n2725 240.244
R6053 GND.n2727 GND.n2726 240.244
R6054 GND.n4854 GND.n2727 240.244
R6055 GND.n4854 GND.n2730 240.244
R6056 GND.n2731 GND.n2730 240.244
R6057 GND.n2732 GND.n2731 240.244
R6058 GND.n4881 GND.n2732 240.244
R6059 GND.n4881 GND.n2735 240.244
R6060 GND.n2736 GND.n2735 240.244
R6061 GND.n2737 GND.n2736 240.244
R6062 GND.n3605 GND.n2737 240.244
R6063 GND.n3605 GND.n2740 240.244
R6064 GND.n2741 GND.n2740 240.244
R6065 GND.n2742 GND.n2741 240.244
R6066 GND.n3588 GND.n2742 240.244
R6067 GND.n3588 GND.n2745 240.244
R6068 GND.n2746 GND.n2745 240.244
R6069 GND.n2747 GND.n2746 240.244
R6070 GND.n5022 GND.n2747 240.244
R6071 GND.n5022 GND.n2750 240.244
R6072 GND.n2751 GND.n2750 240.244
R6073 GND.n2752 GND.n2751 240.244
R6074 GND.n3542 GND.n2752 240.244
R6075 GND.n3542 GND.n2755 240.244
R6076 GND.n2756 GND.n2755 240.244
R6077 GND.n2757 GND.n2756 240.244
R6078 GND.n3514 GND.n2757 240.244
R6079 GND.n3514 GND.n2760 240.244
R6080 GND.n2761 GND.n2760 240.244
R6081 GND.n2762 GND.n2761 240.244
R6082 GND.n3497 GND.n2762 240.244
R6083 GND.n3497 GND.n2765 240.244
R6084 GND.n2766 GND.n2765 240.244
R6085 GND.n2767 GND.n2766 240.244
R6086 GND.n5113 GND.n2767 240.244
R6087 GND.n5113 GND.n2770 240.244
R6088 GND.n2771 GND.n2770 240.244
R6089 GND.n2772 GND.n2771 240.244
R6090 GND.n3461 GND.n2772 240.244
R6091 GND.n3461 GND.n2775 240.244
R6092 GND.n2776 GND.n2775 240.244
R6093 GND.n2777 GND.n2776 240.244
R6094 GND.n3433 GND.n2777 240.244
R6095 GND.n3433 GND.n2780 240.244
R6096 GND.n2781 GND.n2780 240.244
R6097 GND.n2782 GND.n2781 240.244
R6098 GND.n3414 GND.n2782 240.244
R6099 GND.n3414 GND.n2785 240.244
R6100 GND.n2786 GND.n2785 240.244
R6101 GND.n2787 GND.n2786 240.244
R6102 GND.n5329 GND.n2787 240.244
R6103 GND.n5329 GND.n2790 240.244
R6104 GND.n2791 GND.n2790 240.244
R6105 GND.n2792 GND.n2791 240.244
R6106 GND.n3371 GND.n2792 240.244
R6107 GND.n3371 GND.n2795 240.244
R6108 GND.n2796 GND.n2795 240.244
R6109 GND.n2797 GND.n2796 240.244
R6110 GND.n5420 GND.n2797 240.244
R6111 GND.n5420 GND.n2800 240.244
R6112 GND.n2801 GND.n2800 240.244
R6113 GND.n2802 GND.n2801 240.244
R6114 GND.n3332 GND.n2802 240.244
R6115 GND.n3332 GND.n2805 240.244
R6116 GND.n2806 GND.n2805 240.244
R6117 GND.n2807 GND.n2806 240.244
R6118 GND.n5499 GND.n2807 240.244
R6119 GND.n5499 GND.n2810 240.244
R6120 GND.n2811 GND.n2810 240.244
R6121 GND.n2812 GND.n2811 240.244
R6122 GND.n5536 GND.n2812 240.244
R6123 GND.n5536 GND.n2815 240.244
R6124 GND.n2816 GND.n2815 240.244
R6125 GND.n2817 GND.n2816 240.244
R6126 GND.n5563 GND.n2817 240.244
R6127 GND.n5563 GND.n2820 240.244
R6128 GND.n2821 GND.n2820 240.244
R6129 GND.n2822 GND.n2821 240.244
R6130 GND.n5612 GND.n2822 240.244
R6131 GND.n5612 GND.n2825 240.244
R6132 GND.n2826 GND.n2825 240.244
R6133 GND.n2827 GND.n2826 240.244
R6134 GND.n6055 GND.n6053 237.732
R6135 GND.n3937 GND.t138 235.505
R6136 GND.n3188 GND.t102 235.505
R6137 GND.n3944 GND.t88 235.505
R6138 GND.n3173 GND.t169 235.505
R6139 GND.n1399 GND.t124 235.228
R6140 GND.n1414 GND.t143 235.228
R6141 GND.n1430 GND.t183 235.228
R6142 GND.n1920 GND.t152 235.228
R6143 GND.n2179 GND.t158 235.228
R6144 GND.n3081 GND.t196 235.228
R6145 GND.n5800 GND.t166 235.228
R6146 GND.n5813 GND.t149 235.228
R6147 GND.n312 GND.t180 235.228
R6148 GND.n299 GND.t186 235.228
R6149 GND.n288 GND.t120 235.228
R6150 GND.n6258 GND.t199 235.228
R6151 GND.n6113 GND.t98 235.228
R6152 GND.n1257 GND.t163 235.228
R6153 GND.n1271 GND.t146 235.228
R6154 GND.n1284 GND.t110 235.228
R6155 GND.n4239 GND.t189 234.108
R6156 GND.n2892 GND.t106 234.108
R6157 GND.n6055 GND.n6054 224.196
R6158 GND.n1910 GND.n1880 214.453
R6159 GND.n4303 GND.n4273 214.453
R6160 GND.n2863 GND.n2833 214.453
R6161 GND.n6096 GND.n6066 214.453
R6162 GND.n1934 GND.n1406 199.319
R6163 GND.n3938 GND.t139 198.677
R6164 GND.n3189 GND.t105 198.677
R6165 GND.n3945 GND.t90 198.677
R6166 GND.n3174 GND.t171 198.677
R6167 GND.n3966 GND.n3964 186.49
R6168 GND.n3109 GND.n3107 186.49
R6169 GND.n7376 GND.n7375 185.811
R6170 GND.n7377 GND.n7376 185.811
R6171 GND.n7377 GND.n1029 185.811
R6172 GND.n7385 GND.n1029 185.811
R6173 GND.n7386 GND.n7385 185.811
R6174 GND.n7387 GND.n7386 185.811
R6175 GND.n7387 GND.n1023 185.811
R6176 GND.n7395 GND.n1023 185.811
R6177 GND.n7396 GND.n7395 185.811
R6178 GND.n7397 GND.n7396 185.811
R6179 GND.n7397 GND.n1017 185.811
R6180 GND.n7405 GND.n1017 185.811
R6181 GND.n7406 GND.n7405 185.811
R6182 GND.n7407 GND.n7406 185.811
R6183 GND.n7407 GND.n1011 185.811
R6184 GND.n7415 GND.n1011 185.811
R6185 GND.n7416 GND.n7415 185.811
R6186 GND.n7417 GND.n7416 185.811
R6187 GND.n7417 GND.n1005 185.811
R6188 GND.n7425 GND.n1005 185.811
R6189 GND.n7426 GND.n7425 185.811
R6190 GND.n7427 GND.n7426 185.811
R6191 GND.n7427 GND.n999 185.811
R6192 GND.n7435 GND.n999 185.811
R6193 GND.n7436 GND.n7435 185.811
R6194 GND.n7437 GND.n7436 185.811
R6195 GND.n7437 GND.n993 185.811
R6196 GND.n7445 GND.n993 185.811
R6197 GND.n7446 GND.n7445 185.811
R6198 GND.n7447 GND.n7446 185.811
R6199 GND.n7447 GND.n987 185.811
R6200 GND.n7455 GND.n987 185.811
R6201 GND.n7456 GND.n7455 185.811
R6202 GND.n7457 GND.n7456 185.811
R6203 GND.n7457 GND.n981 185.811
R6204 GND.n7465 GND.n981 185.811
R6205 GND.n7466 GND.n7465 185.811
R6206 GND.n7467 GND.n7466 185.811
R6207 GND.n7467 GND.n975 185.811
R6208 GND.n7475 GND.n975 185.811
R6209 GND.n7476 GND.n7475 185.811
R6210 GND.n7477 GND.n7476 185.811
R6211 GND.n7477 GND.n969 185.811
R6212 GND.n7485 GND.n969 185.811
R6213 GND.n7486 GND.n7485 185.811
R6214 GND.n7487 GND.n7486 185.811
R6215 GND.n7487 GND.n963 185.811
R6216 GND.n7495 GND.n963 185.811
R6217 GND.n7496 GND.n7495 185.811
R6218 GND.n7497 GND.n7496 185.811
R6219 GND.n7497 GND.n957 185.811
R6220 GND.n7505 GND.n957 185.811
R6221 GND.n7506 GND.n7505 185.811
R6222 GND.n7507 GND.n7506 185.811
R6223 GND.n7507 GND.n951 185.811
R6224 GND.n7515 GND.n951 185.811
R6225 GND.n7516 GND.n7515 185.811
R6226 GND.n7517 GND.n7516 185.811
R6227 GND.n7517 GND.n945 185.811
R6228 GND.n7525 GND.n945 185.811
R6229 GND.n7526 GND.n7525 185.811
R6230 GND.n7527 GND.n7526 185.811
R6231 GND.n7527 GND.n939 185.811
R6232 GND.n7535 GND.n939 185.811
R6233 GND.n7536 GND.n7535 185.811
R6234 GND.n7537 GND.n7536 185.811
R6235 GND.n7537 GND.n933 185.811
R6236 GND.n7545 GND.n933 185.811
R6237 GND.n7546 GND.n7545 185.811
R6238 GND.n7547 GND.n7546 185.811
R6239 GND.n7547 GND.n927 185.811
R6240 GND.n7555 GND.n927 185.811
R6241 GND.n7556 GND.n7555 185.811
R6242 GND.n7557 GND.n7556 185.811
R6243 GND.n7557 GND.n921 185.811
R6244 GND.n7565 GND.n921 185.811
R6245 GND.n7566 GND.n7565 185.811
R6246 GND.n7567 GND.n7566 185.811
R6247 GND.n7567 GND.n915 185.811
R6248 GND.n7575 GND.n915 185.811
R6249 GND.n7576 GND.n7575 185.811
R6250 GND.n7577 GND.n7576 185.811
R6251 GND.n7577 GND.n909 185.811
R6252 GND.n7585 GND.n909 185.811
R6253 GND.n7586 GND.n7585 185.811
R6254 GND.n7587 GND.n7586 185.811
R6255 GND.n7587 GND.n903 185.811
R6256 GND.n7595 GND.n903 185.811
R6257 GND.n7596 GND.n7595 185.811
R6258 GND.n7597 GND.n7596 185.811
R6259 GND.n7597 GND.n897 185.811
R6260 GND.n7605 GND.n897 185.811
R6261 GND.n7606 GND.n7605 185.811
R6262 GND.n7607 GND.n7606 185.811
R6263 GND.n7607 GND.n891 185.811
R6264 GND.n7615 GND.n891 185.811
R6265 GND.n7616 GND.n7615 185.811
R6266 GND.n7617 GND.n7616 185.811
R6267 GND.n7617 GND.n885 185.811
R6268 GND.n7625 GND.n885 185.811
R6269 GND.n7626 GND.n7625 185.811
R6270 GND.n7627 GND.n7626 185.811
R6271 GND.n7627 GND.n879 185.811
R6272 GND.n7635 GND.n879 185.811
R6273 GND.n7636 GND.n7635 185.811
R6274 GND.n7637 GND.n7636 185.811
R6275 GND.n7637 GND.n873 185.811
R6276 GND.n7645 GND.n873 185.811
R6277 GND.n7646 GND.n7645 185.811
R6278 GND.n7647 GND.n7646 185.811
R6279 GND.n7647 GND.n867 185.811
R6280 GND.n7655 GND.n867 185.811
R6281 GND.n7656 GND.n7655 185.811
R6282 GND.n7657 GND.n7656 185.811
R6283 GND.n7657 GND.n861 185.811
R6284 GND.n7665 GND.n861 185.811
R6285 GND.n7666 GND.n7665 185.811
R6286 GND.n7667 GND.n7666 185.811
R6287 GND.n7667 GND.n855 185.811
R6288 GND.n7675 GND.n855 185.811
R6289 GND.n7676 GND.n7675 185.811
R6290 GND.n7677 GND.n7676 185.811
R6291 GND.n7677 GND.n849 185.811
R6292 GND.n7685 GND.n849 185.811
R6293 GND.n7686 GND.n7685 185.811
R6294 GND.n7687 GND.n7686 185.811
R6295 GND.n7687 GND.n843 185.811
R6296 GND.n7695 GND.n843 185.811
R6297 GND.n7696 GND.n7695 185.811
R6298 GND.n7697 GND.n7696 185.811
R6299 GND.n7697 GND.n837 185.811
R6300 GND.n7705 GND.n837 185.811
R6301 GND.n7706 GND.n7705 185.811
R6302 GND.n7707 GND.n7706 185.811
R6303 GND.n7707 GND.n831 185.811
R6304 GND.n7715 GND.n831 185.811
R6305 GND.n7716 GND.n7715 185.811
R6306 GND.n7717 GND.n7716 185.811
R6307 GND.n7717 GND.n825 185.811
R6308 GND.n7725 GND.n825 185.811
R6309 GND.n7726 GND.n7725 185.811
R6310 GND.n7727 GND.n7726 185.811
R6311 GND.n7727 GND.n819 185.811
R6312 GND.n7735 GND.n819 185.811
R6313 GND.n7736 GND.n7735 185.811
R6314 GND.n7737 GND.n7736 185.811
R6315 GND.n7737 GND.n813 185.811
R6316 GND.n7745 GND.n813 185.811
R6317 GND.n7746 GND.n7745 185.811
R6318 GND.n7747 GND.n7746 185.811
R6319 GND.n7747 GND.n807 185.811
R6320 GND.n7755 GND.n807 185.811
R6321 GND.n7756 GND.n7755 185.811
R6322 GND.n7757 GND.n7756 185.811
R6323 GND.n7757 GND.n801 185.811
R6324 GND.n7765 GND.n801 185.811
R6325 GND.n7766 GND.n7765 185.811
R6326 GND.n7767 GND.n7766 185.811
R6327 GND.n7767 GND.n795 185.811
R6328 GND.n7775 GND.n795 185.811
R6329 GND.n7776 GND.n7775 185.811
R6330 GND.n7777 GND.n7776 185.811
R6331 GND.n7777 GND.n789 185.811
R6332 GND.n7785 GND.n789 185.811
R6333 GND.n7786 GND.n7785 185.811
R6334 GND.n7787 GND.n7786 185.811
R6335 GND.n7787 GND.n783 185.811
R6336 GND.n7795 GND.n783 185.811
R6337 GND.n7796 GND.n7795 185.811
R6338 GND.n7797 GND.n7796 185.811
R6339 GND.n7797 GND.n777 185.811
R6340 GND.n7805 GND.n777 185.811
R6341 GND.n7806 GND.n7805 185.811
R6342 GND.n7807 GND.n7806 185.811
R6343 GND.n7807 GND.n771 185.811
R6344 GND.n7815 GND.n771 185.811
R6345 GND.n7816 GND.n7815 185.811
R6346 GND.n7817 GND.n7816 185.811
R6347 GND.n7817 GND.n765 185.811
R6348 GND.n7825 GND.n765 185.811
R6349 GND.n7826 GND.n7825 185.811
R6350 GND.n7827 GND.n7826 185.811
R6351 GND.n7827 GND.n759 185.811
R6352 GND.n7835 GND.n759 185.811
R6353 GND.n7836 GND.n7835 185.811
R6354 GND.n7837 GND.n7836 185.811
R6355 GND.n7837 GND.n753 185.811
R6356 GND.n7845 GND.n753 185.811
R6357 GND.n7846 GND.n7845 185.811
R6358 GND.n7847 GND.n7846 185.811
R6359 GND.n7847 GND.n747 185.811
R6360 GND.n7855 GND.n747 185.811
R6361 GND.n7856 GND.n7855 185.811
R6362 GND.n7857 GND.n7856 185.811
R6363 GND.n7857 GND.n741 185.811
R6364 GND.n7865 GND.n741 185.811
R6365 GND.n7866 GND.n7865 185.811
R6366 GND.n7867 GND.n7866 185.811
R6367 GND.n7867 GND.n735 185.811
R6368 GND.n7875 GND.n735 185.811
R6369 GND.n7876 GND.n7875 185.811
R6370 GND.n7877 GND.n7876 185.811
R6371 GND.n7877 GND.n729 185.811
R6372 GND.n7885 GND.n729 185.811
R6373 GND.n7886 GND.n7885 185.811
R6374 GND.n7887 GND.n7886 185.811
R6375 GND.n7887 GND.n723 185.811
R6376 GND.n7895 GND.n723 185.811
R6377 GND.n7896 GND.n7895 185.811
R6378 GND.n7897 GND.n7896 185.811
R6379 GND.n7897 GND.n717 185.811
R6380 GND.n7905 GND.n717 185.811
R6381 GND.n7906 GND.n7905 185.811
R6382 GND.n7907 GND.n7906 185.811
R6383 GND.n7907 GND.n711 185.811
R6384 GND.n7915 GND.n711 185.811
R6385 GND.n7916 GND.n7915 185.811
R6386 GND.n7917 GND.n7916 185.811
R6387 GND.n7917 GND.n705 185.811
R6388 GND.n7925 GND.n705 185.811
R6389 GND.n7926 GND.n7925 185.811
R6390 GND.n7927 GND.n7926 185.811
R6391 GND.n7927 GND.n699 185.811
R6392 GND.n7935 GND.n699 185.811
R6393 GND.n7936 GND.n7935 185.811
R6394 GND.n7937 GND.n7936 185.811
R6395 GND.n7937 GND.n693 185.811
R6396 GND.n7945 GND.n693 185.811
R6397 GND.n7946 GND.n7945 185.811
R6398 GND.n7947 GND.n7946 185.811
R6399 GND.n7947 GND.n687 185.811
R6400 GND.n7955 GND.n687 185.811
R6401 GND.n7956 GND.n7955 185.811
R6402 GND.n7957 GND.n7956 185.811
R6403 GND.n7957 GND.n681 185.811
R6404 GND.n7965 GND.n681 185.811
R6405 GND.n7966 GND.n7965 185.811
R6406 GND.n7967 GND.n7966 185.811
R6407 GND.n7967 GND.n675 185.811
R6408 GND.n7975 GND.n675 185.811
R6409 GND.n7976 GND.n7975 185.811
R6410 GND.n7977 GND.n7976 185.811
R6411 GND.n7977 GND.n669 185.811
R6412 GND.n7985 GND.n669 185.811
R6413 GND.n7986 GND.n7985 185.811
R6414 GND.n7987 GND.n7986 185.811
R6415 GND.n7987 GND.n663 185.811
R6416 GND.n7995 GND.n663 185.811
R6417 GND.n7996 GND.n7995 185.811
R6418 GND.n7997 GND.n7996 185.811
R6419 GND.n7997 GND.n657 185.811
R6420 GND.n8005 GND.n657 185.811
R6421 GND.n8006 GND.n8005 185.811
R6422 GND.n8007 GND.n8006 185.811
R6423 GND.n8007 GND.n651 185.811
R6424 GND.n8015 GND.n651 185.811
R6425 GND.n8016 GND.n8015 185.811
R6426 GND.n8017 GND.n8016 185.811
R6427 GND.n8017 GND.n645 185.811
R6428 GND.n8025 GND.n645 185.811
R6429 GND.n8026 GND.n8025 185.811
R6430 GND.n8027 GND.n8026 185.811
R6431 GND.n8027 GND.n639 185.811
R6432 GND.n8035 GND.n639 185.811
R6433 GND.n8036 GND.n8035 185.811
R6434 GND.n8037 GND.n8036 185.811
R6435 GND.n8037 GND.n633 185.811
R6436 GND.n8045 GND.n633 185.811
R6437 GND.n8046 GND.n8045 185.811
R6438 GND.n8047 GND.n8046 185.811
R6439 GND.n8047 GND.n627 185.811
R6440 GND.n8055 GND.n627 185.811
R6441 GND.n8056 GND.n8055 185.811
R6442 GND.n8057 GND.n8056 185.811
R6443 GND.n8057 GND.n621 185.811
R6444 GND.n8065 GND.n621 185.811
R6445 GND.n8066 GND.n8065 185.811
R6446 GND.n8067 GND.n8066 185.811
R6447 GND.n8067 GND.n615 185.811
R6448 GND.n8075 GND.n615 185.811
R6449 GND.n8076 GND.n8075 185.811
R6450 GND.n8077 GND.n8076 185.811
R6451 GND.n8077 GND.n609 185.811
R6452 GND.n8085 GND.n609 185.811
R6453 GND.n8086 GND.n8085 185.811
R6454 GND.n8087 GND.n8086 185.811
R6455 GND.n8087 GND.n603 185.811
R6456 GND.n8095 GND.n603 185.811
R6457 GND.n8096 GND.n8095 185.811
R6458 GND.n8097 GND.n8096 185.811
R6459 GND.n8097 GND.n597 185.811
R6460 GND.n8105 GND.n597 185.811
R6461 GND.n8106 GND.n8105 185.811
R6462 GND.n8107 GND.n8106 185.811
R6463 GND.n8107 GND.n591 185.811
R6464 GND.n8115 GND.n591 185.811
R6465 GND.n8116 GND.n8115 185.811
R6466 GND.n8117 GND.n8116 185.811
R6467 GND.n8117 GND.n585 185.811
R6468 GND.n8125 GND.n585 185.811
R6469 GND.n8126 GND.n8125 185.811
R6470 GND.n8127 GND.n8126 185.811
R6471 GND.n8127 GND.n579 185.811
R6472 GND.n8135 GND.n579 185.811
R6473 GND.n8136 GND.n8135 185.811
R6474 GND.n8137 GND.n8136 185.811
R6475 GND.n8137 GND.n573 185.811
R6476 GND.n8145 GND.n573 185.811
R6477 GND.n8146 GND.n8145 185.811
R6478 GND.n8147 GND.n8146 185.811
R6479 GND.n8147 GND.n567 185.811
R6480 GND.n8155 GND.n567 185.811
R6481 GND.n8156 GND.n8155 185.811
R6482 GND.n8157 GND.n8156 185.811
R6483 GND.n8157 GND.n561 185.811
R6484 GND.n8165 GND.n561 185.811
R6485 GND.n8166 GND.n8165 185.811
R6486 GND.n8167 GND.n8166 185.811
R6487 GND.n8167 GND.n555 185.811
R6488 GND.n8175 GND.n555 185.811
R6489 GND.n8176 GND.n8175 185.811
R6490 GND.n8177 GND.n8176 185.811
R6491 GND.n8177 GND.n549 185.811
R6492 GND.n8185 GND.n549 185.811
R6493 GND.n8186 GND.n8185 185.811
R6494 GND.n8187 GND.n8186 185.811
R6495 GND.n8187 GND.n543 185.811
R6496 GND.n8195 GND.n543 185.811
R6497 GND.n8196 GND.n8195 185.811
R6498 GND.n8197 GND.n8196 185.811
R6499 GND.n8197 GND.n537 185.811
R6500 GND.n8206 GND.n537 185.811
R6501 GND.n8207 GND.n8206 185.811
R6502 GND.n8208 GND.n8207 185.811
R6503 GND.n8208 GND.n532 185.811
R6504 GND.n22 GND.n21 185
R6505 GND.n20 GND.n19 185
R6506 GND.n37 GND.n36 185
R6507 GND.n35 GND.n34 185
R6508 GND.n53 GND.n52 185
R6509 GND.n51 GND.n50 185
R6510 GND.n7 GND.n6 185
R6511 GND.n5 GND.n4 185
R6512 GND.n1911 GND.n1910 185
R6513 GND.n1909 GND.n1908 185
R6514 GND.n1884 GND.n1883 185
R6515 GND.n1903 GND.n1902 185
R6516 GND.n1901 GND.n1900 185
R6517 GND.n1888 GND.n1887 185
R6518 GND.n1895 GND.n1894 185
R6519 GND.n1893 GND.n1892 185
R6520 GND.n4286 GND.n4285 185
R6521 GND.n4288 GND.n4287 185
R6522 GND.n4281 GND.n4280 185
R6523 GND.n4294 GND.n4293 185
R6524 GND.n4296 GND.n4295 185
R6525 GND.n4277 GND.n4276 185
R6526 GND.n4302 GND.n4301 185
R6527 GND.n4304 GND.n4303 185
R6528 GND.n2846 GND.n2845 185
R6529 GND.n2848 GND.n2847 185
R6530 GND.n2841 GND.n2840 185
R6531 GND.n2854 GND.n2853 185
R6532 GND.n2856 GND.n2855 185
R6533 GND.n2837 GND.n2836 185
R6534 GND.n2862 GND.n2861 185
R6535 GND.n2864 GND.n2863 185
R6536 GND.n83 GND.n82 185
R6537 GND.n81 GND.n80 185
R6538 GND.n98 GND.n97 185
R6539 GND.n96 GND.n95 185
R6540 GND.n114 GND.n113 185
R6541 GND.n112 GND.n111 185
R6542 GND.n130 GND.n129 185
R6543 GND.n128 GND.n127 185
R6544 GND.n6097 GND.n6096 185
R6545 GND.n6095 GND.n6094 185
R6546 GND.n6070 GND.n6069 185
R6547 GND.n6089 GND.n6088 185
R6548 GND.n6087 GND.n6086 185
R6549 GND.n6074 GND.n6073 185
R6550 GND.n6081 GND.n6080 185
R6551 GND.n6079 GND.n6078 185
R6552 GND.n1451 GND.t142 181.262
R6553 GND.n1587 GND.t162 181.262
R6554 GND.n64 GND.t19 180.314
R6555 GND.n1399 GND.t126 179.136
R6556 GND.n1414 GND.t144 179.136
R6557 GND.n1430 GND.t184 179.136
R6558 GND.n1920 GND.t153 179.136
R6559 GND.n2179 GND.t160 179.136
R6560 GND.n3081 GND.t198 179.136
R6561 GND.n5800 GND.t168 179.136
R6562 GND.n5813 GND.t151 179.136
R6563 GND.n312 GND.t181 179.136
R6564 GND.n299 GND.t187 179.136
R6565 GND.n288 GND.t122 179.136
R6566 GND.n6258 GND.t200 179.136
R6567 GND.n6113 GND.t101 179.136
R6568 GND.n1257 GND.t165 179.136
R6569 GND.n1271 GND.t148 179.136
R6570 GND.n1284 GND.t113 179.136
R6571 GND.n67 GND.t81 178.752
R6572 GND.n66 GND.t83 178.752
R6573 GND.n65 GND.t49 178.752
R6574 GND.n64 GND.t3 178.752
R6575 GND.n1451 GND.t134 178.565
R6576 GND.n1587 GND.t95 178.565
R6577 GND.n3122 GND.n3120 163.367
R6578 GND.n3126 GND.n3102 163.367
R6579 GND.n3130 GND.n3128 163.367
R6580 GND.n3134 GND.n3100 163.367
R6581 GND.n3138 GND.n3136 163.367
R6582 GND.n3142 GND.n3098 163.367
R6583 GND.n3146 GND.n3144 163.367
R6584 GND.n3150 GND.n3096 163.367
R6585 GND.n3154 GND.n3152 163.367
R6586 GND.n3158 GND.n3094 163.367
R6587 GND.n3162 GND.n3160 163.367
R6588 GND.n3166 GND.n3092 163.367
R6589 GND.n3170 GND.n3168 163.367
R6590 GND.n3177 GND.n3090 163.367
R6591 GND.n3180 GND.n3179 163.367
R6592 GND.n3184 GND.n3183 163.367
R6593 GND.n5787 GND.n5786 163.367
R6594 GND.n5784 GND.n3187 163.367
R6595 GND.n5779 GND.n5778 163.367
R6596 GND.n5776 GND.n3192 163.367
R6597 GND.n5772 GND.n5771 163.367
R6598 GND.n5769 GND.n3195 163.367
R6599 GND.n5765 GND.n5764 163.367
R6600 GND.n5762 GND.n3198 163.367
R6601 GND.n5758 GND.n5757 163.367
R6602 GND.n5755 GND.n3201 163.367
R6603 GND.n5751 GND.n5750 163.367
R6604 GND.n5748 GND.n3204 163.367
R6605 GND.n5744 GND.n5743 163.367
R6606 GND.n5741 GND.n3207 163.367
R6607 GND.n5737 GND.n5736 163.367
R6608 GND.n5734 GND.n3210 163.367
R6609 GND.n4109 GND.n2540 163.367
R6610 GND.n4113 GND.n2540 163.367
R6611 GND.n4113 GND.n2547 163.367
R6612 GND.n4117 GND.n2547 163.367
R6613 GND.n4122 GND.n4117 163.367
R6614 GND.n4123 GND.n4122 163.367
R6615 GND.n4123 GND.n2557 163.367
R6616 GND.n4126 GND.n2557 163.367
R6617 GND.n4126 GND.n2565 163.367
R6618 GND.n4130 GND.n2565 163.367
R6619 GND.n4135 GND.n4130 163.367
R6620 GND.n4136 GND.n4135 163.367
R6621 GND.n4136 GND.n2575 163.367
R6622 GND.n4140 GND.n2575 163.367
R6623 GND.n4140 GND.n2582 163.367
R6624 GND.n4144 GND.n2582 163.367
R6625 GND.n4149 GND.n4144 163.367
R6626 GND.n4150 GND.n4149 163.367
R6627 GND.n4150 GND.n2592 163.367
R6628 GND.n4153 GND.n2592 163.367
R6629 GND.n4153 GND.n2600 163.367
R6630 GND.n4157 GND.n2600 163.367
R6631 GND.n4162 GND.n4157 163.367
R6632 GND.n4163 GND.n4162 163.367
R6633 GND.n4163 GND.n2610 163.367
R6634 GND.n4166 GND.n2610 163.367
R6635 GND.n4166 GND.n2618 163.367
R6636 GND.n4170 GND.n2618 163.367
R6637 GND.n4175 GND.n4170 163.367
R6638 GND.n4176 GND.n4175 163.367
R6639 GND.n4176 GND.n2628 163.367
R6640 GND.n4179 GND.n2628 163.367
R6641 GND.n4179 GND.n2636 163.367
R6642 GND.n4183 GND.n2636 163.367
R6643 GND.n4188 GND.n4183 163.367
R6644 GND.n4189 GND.n4188 163.367
R6645 GND.n4189 GND.n2646 163.367
R6646 GND.n4193 GND.n2646 163.367
R6647 GND.n4193 GND.n2653 163.367
R6648 GND.n3914 GND.n2653 163.367
R6649 GND.n4205 GND.n3914 163.367
R6650 GND.n4205 GND.n3915 163.367
R6651 GND.n4201 GND.n3915 163.367
R6652 GND.n4201 GND.n3899 163.367
R6653 GND.n4198 GND.n3899 163.367
R6654 GND.n4198 GND.n3891 163.367
R6655 GND.n3891 GND.n3884 163.367
R6656 GND.n4359 GND.n3884 163.367
R6657 GND.n4359 GND.n3882 163.367
R6658 GND.n4377 GND.n3882 163.367
R6659 GND.n4377 GND.n3876 163.367
R6660 GND.n4373 GND.n3876 163.367
R6661 GND.n4373 GND.n3867 163.367
R6662 GND.n4369 GND.n3867 163.367
R6663 GND.n4369 GND.n3861 163.367
R6664 GND.n4366 GND.n3861 163.367
R6665 GND.n4366 GND.n3852 163.367
R6666 GND.n3852 GND.n3845 163.367
R6667 GND.n4444 GND.n3845 163.367
R6668 GND.n4444 GND.n3842 163.367
R6669 GND.n4467 GND.n3842 163.367
R6670 GND.n4467 GND.n3843 163.367
R6671 GND.n3843 GND.n3836 163.367
R6672 GND.n4462 GND.n3836 163.367
R6673 GND.n4462 GND.n3827 163.367
R6674 GND.n4457 GND.n3827 163.367
R6675 GND.n4457 GND.n3821 163.367
R6676 GND.n4454 GND.n3821 163.367
R6677 GND.n4454 GND.n3813 163.367
R6678 GND.n4448 GND.n3813 163.367
R6679 GND.n4448 GND.n3805 163.367
R6680 GND.n3805 GND.n3796 163.367
R6681 GND.n4532 GND.n3796 163.367
R6682 GND.n4532 GND.n3794 163.367
R6683 GND.n4566 GND.n3794 163.367
R6684 GND.n4566 GND.n3786 163.367
R6685 GND.n4562 GND.n3786 163.367
R6686 GND.n4562 GND.n4559 163.367
R6687 GND.n4559 GND.n4558 163.367
R6688 GND.n4558 GND.n3769 163.367
R6689 GND.n3770 GND.n3769 163.367
R6690 GND.n3770 GND.n3762 163.367
R6691 GND.n4552 GND.n3762 163.367
R6692 GND.n4552 GND.n3755 163.367
R6693 GND.n4548 GND.n3755 163.367
R6694 GND.n4548 GND.n3749 163.367
R6695 GND.n4545 GND.n3749 163.367
R6696 GND.n4545 GND.n3741 163.367
R6697 GND.n4541 GND.n3741 163.367
R6698 GND.n4541 GND.n3735 163.367
R6699 GND.n4538 GND.n3735 163.367
R6700 GND.n4538 GND.n3725 163.367
R6701 GND.n3725 GND.n3716 163.367
R6702 GND.n4696 GND.n3716 163.367
R6703 GND.n4696 GND.n3714 163.367
R6704 GND.n4702 GND.n3714 163.367
R6705 GND.n4702 GND.n3704 163.367
R6706 GND.n3706 GND.n3704 163.367
R6707 GND.n3706 GND.n3698 163.367
R6708 GND.n4726 GND.n3698 163.367
R6709 GND.n4726 GND.n3692 163.367
R6710 GND.n4730 GND.n3692 163.367
R6711 GND.n4730 GND.n3683 163.367
R6712 GND.n4750 GND.n3683 163.367
R6713 GND.n4750 GND.n3681 163.367
R6714 GND.n4773 GND.n3681 163.367
R6715 GND.n4773 GND.n3675 163.367
R6716 GND.n4769 GND.n3675 163.367
R6717 GND.n4769 GND.n3667 163.367
R6718 GND.n4765 GND.n3667 163.367
R6719 GND.n4765 GND.n3661 163.367
R6720 GND.n4762 GND.n3661 163.367
R6721 GND.n4762 GND.n3653 163.367
R6722 GND.n4758 GND.n3653 163.367
R6723 GND.n4758 GND.n3647 163.367
R6724 GND.n4755 GND.n3647 163.367
R6725 GND.n4755 GND.n3637 163.367
R6726 GND.n3637 GND.n3629 163.367
R6727 GND.n4873 GND.n3629 163.367
R6728 GND.n4873 GND.n3627 163.367
R6729 GND.n4879 GND.n3627 163.367
R6730 GND.n4879 GND.n3617 163.367
R6731 GND.n3619 GND.n3617 163.367
R6732 GND.n3619 GND.n3611 163.367
R6733 GND.n4903 GND.n3611 163.367
R6734 GND.n4903 GND.n3604 163.367
R6735 GND.n4907 GND.n3604 163.367
R6736 GND.n4907 GND.n3596 163.367
R6737 GND.n4927 GND.n3596 163.367
R6738 GND.n4927 GND.n3594 163.367
R6739 GND.n4950 GND.n3594 163.367
R6740 GND.n4950 GND.n3587 163.367
R6741 GND.n4946 GND.n3587 163.367
R6742 GND.n4946 GND.n3579 163.367
R6743 GND.n4942 GND.n3579 163.367
R6744 GND.n4942 GND.n3573 163.367
R6745 GND.n4939 GND.n3573 163.367
R6746 GND.n4939 GND.n3565 163.367
R6747 GND.n4935 GND.n3565 163.367
R6748 GND.n4935 GND.n3559 163.367
R6749 GND.n4932 GND.n3559 163.367
R6750 GND.n4932 GND.n3549 163.367
R6751 GND.n3549 GND.n3540 163.367
R6752 GND.n5049 GND.n3540 163.367
R6753 GND.n5049 GND.n3538 163.367
R6754 GND.n5055 GND.n3538 163.367
R6755 GND.n5055 GND.n3528 163.367
R6756 GND.n3530 GND.n3528 163.367
R6757 GND.n3530 GND.n3522 163.367
R6758 GND.n5078 GND.n3522 163.367
R6759 GND.n5078 GND.n3516 163.367
R6760 GND.n5082 GND.n3516 163.367
R6761 GND.n5082 GND.n3507 163.367
R6762 GND.n5102 GND.n3507 163.367
R6763 GND.n5102 GND.n3505 163.367
R6764 GND.n5126 GND.n3505 163.367
R6765 GND.n5126 GND.n3499 163.367
R6766 GND.n5122 GND.n3499 163.367
R6767 GND.n5122 GND.n3490 163.367
R6768 GND.n5118 GND.n3490 163.367
R6769 GND.n5118 GND.n3484 163.367
R6770 GND.n5115 GND.n3484 163.367
R6771 GND.n5115 GND.n3476 163.367
R6772 GND.n5110 GND.n3476 163.367
R6773 GND.n5110 GND.n3470 163.367
R6774 GND.n5107 GND.n3470 163.367
R6775 GND.n5107 GND.n3459 163.367
R6776 GND.n3459 GND.n3451 163.367
R6777 GND.n5224 GND.n3451 163.367
R6778 GND.n5224 GND.n3449 163.367
R6779 GND.n5230 GND.n3449 163.367
R6780 GND.n5230 GND.n3439 163.367
R6781 GND.n3441 GND.n3439 163.367
R6782 GND.n3441 GND.n3432 163.367
R6783 GND.n5253 GND.n3432 163.367
R6784 GND.n5253 GND.n3426 163.367
R6785 GND.n5257 GND.n3426 163.367
R6786 GND.n5257 GND.n3418 163.367
R6787 GND.n5277 GND.n3418 163.367
R6788 GND.n5277 GND.n3416 163.367
R6789 GND.n5300 GND.n3416 163.367
R6790 GND.n5300 GND.n3409 163.367
R6791 GND.n5296 GND.n3409 163.367
R6792 GND.n5296 GND.n3401 163.367
R6793 GND.n5292 GND.n3401 163.367
R6794 GND.n5292 GND.n3395 163.367
R6795 GND.n5289 GND.n3395 163.367
R6796 GND.n5289 GND.n3387 163.367
R6797 GND.n5285 GND.n3387 163.367
R6798 GND.n5285 GND.n3381 163.367
R6799 GND.n5282 GND.n3381 163.367
R6800 GND.n5282 GND.n3373 163.367
R6801 GND.n3373 GND.n3364 163.367
R6802 GND.n5401 GND.n3364 163.367
R6803 GND.n5401 GND.n3362 163.367
R6804 GND.n5407 GND.n3362 163.367
R6805 GND.n5407 GND.n3352 163.367
R6806 GND.n3354 GND.n3352 163.367
R6807 GND.n3354 GND.n3346 163.367
R6808 GND.n5431 GND.n3346 163.367
R6809 GND.n5431 GND.n3340 163.367
R6810 GND.n5435 GND.n3340 163.367
R6811 GND.n5435 GND.n3331 163.367
R6812 GND.n5455 GND.n3331 163.367
R6813 GND.n5455 GND.n3329 163.367
R6814 GND.n5478 GND.n3329 163.367
R6815 GND.n5478 GND.n3323 163.367
R6816 GND.n5474 GND.n3323 163.367
R6817 GND.n5474 GND.n3315 163.367
R6818 GND.n5470 GND.n3315 163.367
R6819 GND.n5470 GND.n3309 163.367
R6820 GND.n5467 GND.n3309 163.367
R6821 GND.n5467 GND.n3301 163.367
R6822 GND.n5463 GND.n3301 163.367
R6823 GND.n5463 GND.n3295 163.367
R6824 GND.n5460 GND.n3295 163.367
R6825 GND.n5460 GND.n3285 163.367
R6826 GND.n3285 GND.n3277 163.367
R6827 GND.n5557 GND.n3277 163.367
R6828 GND.n5557 GND.n3275 163.367
R6829 GND.n5561 GND.n3275 163.367
R6830 GND.n5561 GND.n3264 163.367
R6831 GND.n5592 GND.n3264 163.367
R6832 GND.n5592 GND.n3259 163.367
R6833 GND.n5588 GND.n3259 163.367
R6834 GND.n5588 GND.n3250 163.367
R6835 GND.n3250 GND.n3243 163.367
R6836 GND.n5622 GND.n3243 163.367
R6837 GND.n5622 GND.n3240 163.367
R6838 GND.n5628 GND.n3240 163.367
R6839 GND.n5628 GND.n3241 163.367
R6840 GND.n3241 GND.n3218 163.367
R6841 GND.n5638 GND.n3218 163.367
R6842 GND.n5639 GND.n5638 163.367
R6843 GND.n5639 GND.n2915 163.367
R6844 GND.n5643 GND.n2915 163.367
R6845 GND.n5643 GND.n2922 163.367
R6846 GND.n5647 GND.n2922 163.367
R6847 GND.n5652 GND.n5647 163.367
R6848 GND.n5653 GND.n5652 163.367
R6849 GND.n5653 GND.n2932 163.367
R6850 GND.n5656 GND.n2932 163.367
R6851 GND.n5656 GND.n2940 163.367
R6852 GND.n5660 GND.n2940 163.367
R6853 GND.n5665 GND.n5660 163.367
R6854 GND.n5666 GND.n5665 163.367
R6855 GND.n5666 GND.n2950 163.367
R6856 GND.n5669 GND.n2950 163.367
R6857 GND.n5669 GND.n2958 163.367
R6858 GND.n5673 GND.n2958 163.367
R6859 GND.n5678 GND.n5673 163.367
R6860 GND.n5679 GND.n5678 163.367
R6861 GND.n5679 GND.n2968 163.367
R6862 GND.n5682 GND.n2968 163.367
R6863 GND.n5682 GND.n2976 163.367
R6864 GND.n5686 GND.n2976 163.367
R6865 GND.n5691 GND.n5686 163.367
R6866 GND.n5692 GND.n5691 163.367
R6867 GND.n5692 GND.n2986 163.367
R6868 GND.n5696 GND.n2986 163.367
R6869 GND.n5696 GND.n2993 163.367
R6870 GND.n5700 GND.n2993 163.367
R6871 GND.n5705 GND.n5700 163.367
R6872 GND.n5706 GND.n5705 163.367
R6873 GND.n5706 GND.n3003 163.367
R6874 GND.n5709 GND.n3003 163.367
R6875 GND.n5709 GND.n3011 163.367
R6876 GND.n5713 GND.n3011 163.367
R6877 GND.n5718 GND.n5713 163.367
R6878 GND.n5719 GND.n5718 163.367
R6879 GND.n5719 GND.n3021 163.367
R6880 GND.n5722 GND.n3021 163.367
R6881 GND.n5722 GND.n3029 163.367
R6882 GND.n5729 GND.n3029 163.367
R6883 GND.n3978 GND.n3960 163.367
R6884 GND.n3982 GND.n3960 163.367
R6885 GND.n3986 GND.n3984 163.367
R6886 GND.n3990 GND.n3958 163.367
R6887 GND.n3994 GND.n3992 163.367
R6888 GND.n3998 GND.n3956 163.367
R6889 GND.n4002 GND.n4000 163.367
R6890 GND.n4006 GND.n3954 163.367
R6891 GND.n4010 GND.n4008 163.367
R6892 GND.n4014 GND.n3952 163.367
R6893 GND.n4018 GND.n4016 163.367
R6894 GND.n4022 GND.n3950 163.367
R6895 GND.n4026 GND.n4024 163.367
R6896 GND.n4030 GND.n3948 163.367
R6897 GND.n4034 GND.n4032 163.367
R6898 GND.n4038 GND.n3943 163.367
R6899 GND.n4041 GND.n4040 163.367
R6900 GND.n4045 GND.n4043 163.367
R6901 GND.n4049 GND.n3941 163.367
R6902 GND.n4053 GND.n4051 163.367
R6903 GND.n4057 GND.n3936 163.367
R6904 GND.n4061 GND.n4059 163.367
R6905 GND.n4065 GND.n3934 163.367
R6906 GND.n4069 GND.n4067 163.367
R6907 GND.n4073 GND.n3932 163.367
R6908 GND.n4077 GND.n4075 163.367
R6909 GND.n4081 GND.n3930 163.367
R6910 GND.n4085 GND.n4083 163.367
R6911 GND.n4089 GND.n3928 163.367
R6912 GND.n4093 GND.n4091 163.367
R6913 GND.n4097 GND.n3926 163.367
R6914 GND.n4101 GND.n4099 163.367
R6915 GND.n4105 GND.n3924 163.367
R6916 GND.n4108 GND.n4107 163.367
R6917 GND.n6956 GND.n2541 163.367
R6918 GND.n6956 GND.n2542 163.367
R6919 GND.n6952 GND.n2542 163.367
R6920 GND.n6952 GND.n2545 163.367
R6921 GND.n4120 GND.n2545 163.367
R6922 GND.n4120 GND.n2559 163.367
R6923 GND.n6943 GND.n2559 163.367
R6924 GND.n6943 GND.n2560 163.367
R6925 GND.n6939 GND.n2560 163.367
R6926 GND.n6939 GND.n2563 163.367
R6927 GND.n4133 GND.n2563 163.367
R6928 GND.n4133 GND.n2576 163.367
R6929 GND.n6929 GND.n2576 163.367
R6930 GND.n6929 GND.n2577 163.367
R6931 GND.n6925 GND.n2577 163.367
R6932 GND.n6925 GND.n2580 163.367
R6933 GND.n4147 GND.n2580 163.367
R6934 GND.n4147 GND.n2594 163.367
R6935 GND.n6915 GND.n2594 163.367
R6936 GND.n6915 GND.n2595 163.367
R6937 GND.n6911 GND.n2595 163.367
R6938 GND.n6911 GND.n2598 163.367
R6939 GND.n4160 GND.n2598 163.367
R6940 GND.n4160 GND.n2612 163.367
R6941 GND.n6901 GND.n2612 163.367
R6942 GND.n6901 GND.n2613 163.367
R6943 GND.n6897 GND.n2613 163.367
R6944 GND.n6897 GND.n2616 163.367
R6945 GND.n4173 GND.n2616 163.367
R6946 GND.n4173 GND.n2630 163.367
R6947 GND.n6887 GND.n2630 163.367
R6948 GND.n6887 GND.n2631 163.367
R6949 GND.n6883 GND.n2631 163.367
R6950 GND.n6883 GND.n2634 163.367
R6951 GND.n4186 GND.n2634 163.367
R6952 GND.n4186 GND.n2648 163.367
R6953 GND.n6873 GND.n2648 163.367
R6954 GND.n6873 GND.n2649 163.367
R6955 GND.n6869 GND.n2649 163.367
R6956 GND.n6869 GND.n2652 163.367
R6957 GND.n4209 GND.n2652 163.367
R6958 GND.n4209 GND.n4206 163.367
R6959 GND.n4206 GND.n3897 163.367
R6960 GND.n4341 GND.n3897 163.367
R6961 GND.n4341 GND.n3893 163.367
R6962 GND.n4346 GND.n3893 163.367
R6963 GND.n4346 GND.n3895 163.367
R6964 GND.n3895 GND.n3880 163.367
R6965 GND.n4381 GND.n3880 163.367
R6966 GND.n4381 GND.n3878 163.367
R6967 GND.n4385 GND.n3878 163.367
R6968 GND.n4385 GND.n3865 163.367
R6969 GND.n4411 GND.n3865 163.367
R6970 GND.n4411 GND.n3863 163.367
R6971 GND.n4415 GND.n3863 163.367
R6972 GND.n4415 GND.n3850 163.367
R6973 GND.n4438 GND.n3850 163.367
R6974 GND.n4438 GND.n3848 163.367
R6975 GND.n4442 GND.n3848 163.367
R6976 GND.n4442 GND.n3840 163.367
R6977 GND.n4470 GND.n3840 163.367
R6978 GND.n4470 GND.n3838 163.367
R6979 GND.n4474 GND.n3838 163.367
R6980 GND.n4474 GND.n3825 163.367
R6981 GND.n4488 GND.n3825 163.367
R6982 GND.n4488 GND.n3823 163.367
R6983 GND.n4492 GND.n3823 163.367
R6984 GND.n4492 GND.n3811 163.367
R6985 GND.n4514 GND.n3811 163.367
R6986 GND.n4514 GND.n3807 163.367
R6987 GND.n4519 GND.n3807 163.367
R6988 GND.n4519 GND.n3809 163.367
R6989 GND.n3809 GND.n3791 163.367
R6990 GND.n4570 GND.n3791 163.367
R6991 GND.n4570 GND.n3788 163.367
R6992 GND.n4577 GND.n3788 163.367
R6993 GND.n4577 GND.n3789 163.367
R6994 GND.n4573 GND.n3789 163.367
R6995 GND.n4573 GND.n3766 163.367
R6996 GND.n4601 GND.n3766 163.367
R6997 GND.n4601 GND.n3764 163.367
R6998 GND.n4605 GND.n3764 163.367
R6999 GND.n4605 GND.n3753 163.367
R7000 GND.n4620 GND.n3753 163.367
R7001 GND.n4620 GND.n3751 163.367
R7002 GND.n4624 GND.n3751 163.367
R7003 GND.n4624 GND.n3739 163.367
R7004 GND.n4672 GND.n3739 163.367
R7005 GND.n4672 GND.n3737 163.367
R7006 GND.n4676 GND.n3737 163.367
R7007 GND.n4676 GND.n3722 163.367
R7008 GND.n4689 GND.n3722 163.367
R7009 GND.n4689 GND.n3719 163.367
R7010 GND.n4694 GND.n3719 163.367
R7011 GND.n4694 GND.n3720 163.367
R7012 GND.n3720 GND.n3702 163.367
R7013 GND.n4718 GND.n3702 163.367
R7014 GND.n4718 GND.n3700 163.367
R7015 GND.n4722 GND.n3700 163.367
R7016 GND.n4722 GND.n3694 163.367
R7017 GND.n4738 GND.n3694 163.367
R7018 GND.n4738 GND.n3695 163.367
R7019 GND.n4734 GND.n3695 163.367
R7020 GND.n4734 GND.n3679 163.367
R7021 GND.n4777 GND.n3679 163.367
R7022 GND.n4777 GND.n3677 163.367
R7023 GND.n4781 GND.n3677 163.367
R7024 GND.n4781 GND.n3665 163.367
R7025 GND.n4797 GND.n3665 163.367
R7026 GND.n4797 GND.n3663 163.367
R7027 GND.n4801 GND.n3663 163.367
R7028 GND.n4801 GND.n3651 163.367
R7029 GND.n4848 GND.n3651 163.367
R7030 GND.n4848 GND.n3649 163.367
R7031 GND.n4852 GND.n3649 163.367
R7032 GND.n4852 GND.n3635 163.367
R7033 GND.n4866 GND.n3635 163.367
R7034 GND.n4866 GND.n3632 163.367
R7035 GND.n4871 GND.n3632 163.367
R7036 GND.n4871 GND.n3633 163.367
R7037 GND.n3633 GND.n3615 163.367
R7038 GND.n4895 GND.n3615 163.367
R7039 GND.n4895 GND.n3613 163.367
R7040 GND.n4899 GND.n3613 163.367
R7041 GND.n4899 GND.n3607 163.367
R7042 GND.n4915 GND.n3607 163.367
R7043 GND.n4915 GND.n3608 163.367
R7044 GND.n4911 GND.n3608 163.367
R7045 GND.n4911 GND.n3592 163.367
R7046 GND.n4954 GND.n3592 163.367
R7047 GND.n4954 GND.n3590 163.367
R7048 GND.n4958 GND.n3590 163.367
R7049 GND.n4958 GND.n3577 163.367
R7050 GND.n4973 GND.n3577 163.367
R7051 GND.n4973 GND.n3575 163.367
R7052 GND.n4977 GND.n3575 163.367
R7053 GND.n4977 GND.n3563 163.367
R7054 GND.n5025 GND.n3563 163.367
R7055 GND.n5025 GND.n3561 163.367
R7056 GND.n5029 GND.n3561 163.367
R7057 GND.n5029 GND.n3547 163.367
R7058 GND.n5042 GND.n3547 163.367
R7059 GND.n5042 GND.n3544 163.367
R7060 GND.n5047 GND.n3544 163.367
R7061 GND.n5047 GND.n3545 163.367
R7062 GND.n3545 GND.n3526 163.367
R7063 GND.n5070 GND.n3526 163.367
R7064 GND.n5070 GND.n3524 163.367
R7065 GND.n5074 GND.n3524 163.367
R7066 GND.n5074 GND.n3518 163.367
R7067 GND.n5090 GND.n3518 163.367
R7068 GND.n5090 GND.n3519 163.367
R7069 GND.n5086 GND.n3519 163.367
R7070 GND.n5086 GND.n3503 163.367
R7071 GND.n5130 GND.n3503 163.367
R7072 GND.n5130 GND.n3501 163.367
R7073 GND.n5134 GND.n3501 163.367
R7074 GND.n5134 GND.n3488 163.367
R7075 GND.n5149 GND.n3488 163.367
R7076 GND.n5149 GND.n3486 163.367
R7077 GND.n5153 GND.n3486 163.367
R7078 GND.n5153 GND.n3474 163.367
R7079 GND.n5200 GND.n3474 163.367
R7080 GND.n5200 GND.n3472 163.367
R7081 GND.n5204 GND.n3472 163.367
R7082 GND.n5204 GND.n3457 163.367
R7083 GND.n5217 GND.n3457 163.367
R7084 GND.n5217 GND.n3454 163.367
R7085 GND.n5222 GND.n3454 163.367
R7086 GND.n5222 GND.n3455 163.367
R7087 GND.n3455 GND.n3437 163.367
R7088 GND.n5245 GND.n3437 163.367
R7089 GND.n5245 GND.n3435 163.367
R7090 GND.n5249 GND.n3435 163.367
R7091 GND.n5249 GND.n3427 163.367
R7092 GND.n5265 GND.n3427 163.367
R7093 GND.n5265 GND.n3428 163.367
R7094 GND.n5261 GND.n3428 163.367
R7095 GND.n5261 GND.n3413 163.367
R7096 GND.n5304 GND.n3413 163.367
R7097 GND.n5304 GND.n3411 163.367
R7098 GND.n5308 GND.n3411 163.367
R7099 GND.n5308 GND.n3399 163.367
R7100 GND.n5323 GND.n3399 163.367
R7101 GND.n5323 GND.n3397 163.367
R7102 GND.n5327 GND.n3397 163.367
R7103 GND.n5327 GND.n3385 163.367
R7104 GND.n5377 GND.n3385 163.367
R7105 GND.n5377 GND.n3383 163.367
R7106 GND.n5381 GND.n3383 163.367
R7107 GND.n5381 GND.n3370 163.367
R7108 GND.n5394 GND.n3370 163.367
R7109 GND.n5394 GND.n3367 163.367
R7110 GND.n5399 GND.n3367 163.367
R7111 GND.n5399 GND.n3368 163.367
R7112 GND.n3368 GND.n3350 163.367
R7113 GND.n5423 GND.n3350 163.367
R7114 GND.n5423 GND.n3348 163.367
R7115 GND.n5427 GND.n3348 163.367
R7116 GND.n5427 GND.n3342 163.367
R7117 GND.n5443 GND.n3342 163.367
R7118 GND.n5443 GND.n3343 163.367
R7119 GND.n5439 GND.n3343 163.367
R7120 GND.n5439 GND.n3327 163.367
R7121 GND.n5482 GND.n3327 163.367
R7122 GND.n5482 GND.n3325 163.367
R7123 GND.n5486 GND.n3325 163.367
R7124 GND.n5486 GND.n3313 163.367
R7125 GND.n5502 GND.n3313 163.367
R7126 GND.n5502 GND.n3311 163.367
R7127 GND.n5506 GND.n3311 163.367
R7128 GND.n5506 GND.n3299 163.367
R7129 GND.n5530 GND.n3299 163.367
R7130 GND.n5530 GND.n3297 163.367
R7131 GND.n5534 GND.n3297 163.367
R7132 GND.n5534 GND.n3283 163.367
R7133 GND.n5550 GND.n3283 163.367
R7134 GND.n5550 GND.n3280 163.367
R7135 GND.n5555 GND.n3280 163.367
R7136 GND.n5555 GND.n3281 163.367
R7137 GND.n3281 GND.n3262 163.367
R7138 GND.n5596 GND.n3262 163.367
R7139 GND.n5596 GND.n3260 163.367
R7140 GND.n5600 GND.n3260 163.367
R7141 GND.n5600 GND.n3248 163.367
R7142 GND.n5615 GND.n3248 163.367
R7143 GND.n5615 GND.n3246 163.367
R7144 GND.n5620 GND.n3246 163.367
R7145 GND.n5620 GND.n3238 163.367
R7146 GND.n5631 GND.n3238 163.367
R7147 GND.n5632 GND.n5631 163.367
R7148 GND.n5632 GND.n3236 163.367
R7149 GND.n5636 GND.n3236 163.367
R7150 GND.n5636 GND.n2916 163.367
R7151 GND.n6617 GND.n2916 163.367
R7152 GND.n6617 GND.n2917 163.367
R7153 GND.n6613 GND.n2917 163.367
R7154 GND.n6613 GND.n2920 163.367
R7155 GND.n5650 GND.n2920 163.367
R7156 GND.n5650 GND.n2934 163.367
R7157 GND.n6603 GND.n2934 163.367
R7158 GND.n6603 GND.n2935 163.367
R7159 GND.n6599 GND.n2935 163.367
R7160 GND.n6599 GND.n2938 163.367
R7161 GND.n5663 GND.n2938 163.367
R7162 GND.n5663 GND.n2952 163.367
R7163 GND.n6589 GND.n2952 163.367
R7164 GND.n6589 GND.n2953 163.367
R7165 GND.n6585 GND.n2953 163.367
R7166 GND.n6585 GND.n2956 163.367
R7167 GND.n5676 GND.n2956 163.367
R7168 GND.n5676 GND.n2970 163.367
R7169 GND.n6575 GND.n2970 163.367
R7170 GND.n6575 GND.n2971 163.367
R7171 GND.n6571 GND.n2971 163.367
R7172 GND.n6571 GND.n2974 163.367
R7173 GND.n5689 GND.n2974 163.367
R7174 GND.n5689 GND.n2988 163.367
R7175 GND.n6561 GND.n2988 163.367
R7176 GND.n6561 GND.n2989 163.367
R7177 GND.n6557 GND.n2989 163.367
R7178 GND.n6557 GND.n2992 163.367
R7179 GND.n5703 GND.n2992 163.367
R7180 GND.n5703 GND.n3005 163.367
R7181 GND.n6547 GND.n3005 163.367
R7182 GND.n6547 GND.n3006 163.367
R7183 GND.n6543 GND.n3006 163.367
R7184 GND.n6543 GND.n3009 163.367
R7185 GND.n5716 GND.n3009 163.367
R7186 GND.n5716 GND.n3022 163.367
R7187 GND.n6533 GND.n3022 163.367
R7188 GND.n6533 GND.n3023 163.367
R7189 GND.n6529 GND.n3023 163.367
R7190 GND.n6529 GND.n3026 163.367
R7191 GND.n1566 GND.n1565 161.3
R7192 GND.n1567 GND.n1534 161.3
R7193 GND.n1569 GND.n1568 161.3
R7194 GND.n1570 GND.n1533 161.3
R7195 GND.n1572 GND.n1571 161.3
R7196 GND.n1573 GND.n1532 161.3
R7197 GND.n1575 GND.n1574 161.3
R7198 GND.n1576 GND.n1531 161.3
R7199 GND.n1578 GND.n1577 161.3
R7200 GND.n1579 GND.n1530 161.3
R7201 GND.n1581 GND.n1580 161.3
R7202 GND.n1582 GND.n1529 161.3
R7203 GND.n1544 GND.n1543 161.3
R7204 GND.n1545 GND.n1540 161.3
R7205 GND.n1547 GND.n1546 161.3
R7206 GND.n1548 GND.n1539 161.3
R7207 GND.n1550 GND.n1549 161.3
R7208 GND.n1551 GND.n1538 161.3
R7209 GND.n1553 GND.n1552 161.3
R7210 GND.n1554 GND.n1537 161.3
R7211 GND.n1556 GND.n1555 161.3
R7212 GND.n1557 GND.n1536 161.3
R7213 GND.n1559 GND.n1558 161.3
R7214 GND.n1560 GND.n1535 161.3
R7215 GND.n1859 GND.n1858 161.3
R7216 GND.n1860 GND.n1443 161.3
R7217 GND.n1862 GND.n1861 161.3
R7218 GND.n1863 GND.n1442 161.3
R7219 GND.n1865 GND.n1864 161.3
R7220 GND.n1866 GND.n1441 161.3
R7221 GND.n1868 GND.n1867 161.3
R7222 GND.n1869 GND.n1440 161.3
R7223 GND.n1871 GND.n1870 161.3
R7224 GND.n1872 GND.n1438 161.3
R7225 GND.n1838 GND.n1837 161.3
R7226 GND.n1839 GND.n1450 161.3
R7227 GND.n1841 GND.n1840 161.3
R7228 GND.n1842 GND.n1449 161.3
R7229 GND.n1844 GND.n1843 161.3
R7230 GND.n1845 GND.n1448 161.3
R7231 GND.n1847 GND.n1846 161.3
R7232 GND.n1848 GND.n1447 161.3
R7233 GND.n1850 GND.n1849 161.3
R7234 GND.n1851 GND.n1446 161.3
R7235 GND.n1853 GND.n1852 161.3
R7236 GND.n1854 GND.n1445 161.3
R7237 GND.n1648 GND.n1510 161.3
R7238 GND.n1647 GND.n1646 161.3
R7239 GND.n1645 GND.n1511 161.3
R7240 GND.n1644 GND.n1643 161.3
R7241 GND.n1642 GND.n1512 161.3
R7242 GND.n1641 GND.n1640 161.3
R7243 GND.n1639 GND.n1513 161.3
R7244 GND.n1638 GND.n1637 161.3
R7245 GND.n1636 GND.n1514 161.3
R7246 GND.n1635 GND.n1634 161.3
R7247 GND.n1633 GND.n1515 161.3
R7248 GND.n1632 GND.n1631 161.3
R7249 GND.n1629 GND.n1516 161.3
R7250 GND.n1628 GND.n1627 161.3
R7251 GND.n1626 GND.n1517 161.3
R7252 GND.n1625 GND.n1624 161.3
R7253 GND.n1623 GND.n1518 161.3
R7254 GND.n1622 GND.n1621 161.3
R7255 GND.n1620 GND.n1519 161.3
R7256 GND.n1619 GND.n1618 161.3
R7257 GND.n1617 GND.n1520 161.3
R7258 GND.n1616 GND.n1615 161.3
R7259 GND.n1614 GND.n1521 161.3
R7260 GND.n1613 GND.n1612 161.3
R7261 GND.n1611 GND.n1522 161.3
R7262 GND.n1609 GND.n1608 161.3
R7263 GND.n1607 GND.n1523 161.3
R7264 GND.n1606 GND.n1605 161.3
R7265 GND.n1604 GND.n1524 161.3
R7266 GND.n1603 GND.n1602 161.3
R7267 GND.n1601 GND.n1525 161.3
R7268 GND.n1600 GND.n1599 161.3
R7269 GND.n1598 GND.n1526 161.3
R7270 GND.n1597 GND.n1596 161.3
R7271 GND.n1595 GND.n1527 161.3
R7272 GND.n1594 GND.n1593 161.3
R7273 GND.n1592 GND.n1528 161.3
R7274 GND.n1709 GND.n1491 161.3
R7275 GND.n1708 GND.n1707 161.3
R7276 GND.n1706 GND.n1492 161.3
R7277 GND.n1705 GND.n1704 161.3
R7278 GND.n1703 GND.n1493 161.3
R7279 GND.n1702 GND.n1701 161.3
R7280 GND.n1700 GND.n1494 161.3
R7281 GND.n1699 GND.n1698 161.3
R7282 GND.n1697 GND.n1495 161.3
R7283 GND.n1696 GND.n1695 161.3
R7284 GND.n1694 GND.n1496 161.3
R7285 GND.n1693 GND.n1692 161.3
R7286 GND.n1690 GND.n1497 161.3
R7287 GND.n1689 GND.n1688 161.3
R7288 GND.n1687 GND.n1498 161.3
R7289 GND.n1686 GND.n1685 161.3
R7290 GND.n1684 GND.n1499 161.3
R7291 GND.n1683 GND.n1682 161.3
R7292 GND.n1681 GND.n1500 161.3
R7293 GND.n1680 GND.n1679 161.3
R7294 GND.n1678 GND.n1501 161.3
R7295 GND.n1677 GND.n1676 161.3
R7296 GND.n1675 GND.n1502 161.3
R7297 GND.n1674 GND.n1673 161.3
R7298 GND.n1672 GND.n1503 161.3
R7299 GND.n1670 GND.n1669 161.3
R7300 GND.n1668 GND.n1504 161.3
R7301 GND.n1667 GND.n1666 161.3
R7302 GND.n1665 GND.n1505 161.3
R7303 GND.n1664 GND.n1663 161.3
R7304 GND.n1662 GND.n1506 161.3
R7305 GND.n1661 GND.n1660 161.3
R7306 GND.n1659 GND.n1507 161.3
R7307 GND.n1658 GND.n1657 161.3
R7308 GND.n1656 GND.n1508 161.3
R7309 GND.n1655 GND.n1654 161.3
R7310 GND.n1653 GND.n1509 161.3
R7311 GND.n1770 GND.n1472 161.3
R7312 GND.n1769 GND.n1768 161.3
R7313 GND.n1767 GND.n1473 161.3
R7314 GND.n1766 GND.n1765 161.3
R7315 GND.n1764 GND.n1474 161.3
R7316 GND.n1763 GND.n1762 161.3
R7317 GND.n1761 GND.n1475 161.3
R7318 GND.n1760 GND.n1759 161.3
R7319 GND.n1758 GND.n1476 161.3
R7320 GND.n1757 GND.n1756 161.3
R7321 GND.n1755 GND.n1477 161.3
R7322 GND.n1754 GND.n1753 161.3
R7323 GND.n1751 GND.n1478 161.3
R7324 GND.n1750 GND.n1749 161.3
R7325 GND.n1748 GND.n1479 161.3
R7326 GND.n1747 GND.n1746 161.3
R7327 GND.n1745 GND.n1480 161.3
R7328 GND.n1744 GND.n1743 161.3
R7329 GND.n1742 GND.n1481 161.3
R7330 GND.n1741 GND.n1740 161.3
R7331 GND.n1739 GND.n1482 161.3
R7332 GND.n1738 GND.n1737 161.3
R7333 GND.n1736 GND.n1483 161.3
R7334 GND.n1735 GND.n1734 161.3
R7335 GND.n1733 GND.n1484 161.3
R7336 GND.n1731 GND.n1730 161.3
R7337 GND.n1729 GND.n1485 161.3
R7338 GND.n1728 GND.n1727 161.3
R7339 GND.n1726 GND.n1486 161.3
R7340 GND.n1725 GND.n1724 161.3
R7341 GND.n1723 GND.n1487 161.3
R7342 GND.n1722 GND.n1721 161.3
R7343 GND.n1720 GND.n1488 161.3
R7344 GND.n1719 GND.n1718 161.3
R7345 GND.n1717 GND.n1489 161.3
R7346 GND.n1716 GND.n1715 161.3
R7347 GND.n1714 GND.n1490 161.3
R7348 GND.n1831 GND.n1453 161.3
R7349 GND.n1830 GND.n1829 161.3
R7350 GND.n1828 GND.n1454 161.3
R7351 GND.n1827 GND.n1826 161.3
R7352 GND.n1825 GND.n1455 161.3
R7353 GND.n1824 GND.n1823 161.3
R7354 GND.n1822 GND.n1456 161.3
R7355 GND.n1821 GND.n1820 161.3
R7356 GND.n1819 GND.n1457 161.3
R7357 GND.n1818 GND.n1817 161.3
R7358 GND.n1816 GND.n1458 161.3
R7359 GND.n1815 GND.n1814 161.3
R7360 GND.n1812 GND.n1459 161.3
R7361 GND.n1811 GND.n1810 161.3
R7362 GND.n1809 GND.n1460 161.3
R7363 GND.n1808 GND.n1807 161.3
R7364 GND.n1806 GND.n1461 161.3
R7365 GND.n1805 GND.n1804 161.3
R7366 GND.n1803 GND.n1462 161.3
R7367 GND.n1802 GND.n1801 161.3
R7368 GND.n1800 GND.n1463 161.3
R7369 GND.n1799 GND.n1798 161.3
R7370 GND.n1797 GND.n1464 161.3
R7371 GND.n1796 GND.n1795 161.3
R7372 GND.n1794 GND.n1465 161.3
R7373 GND.n1792 GND.n1791 161.3
R7374 GND.n1790 GND.n1466 161.3
R7375 GND.n1789 GND.n1788 161.3
R7376 GND.n1787 GND.n1467 161.3
R7377 GND.n1786 GND.n1785 161.3
R7378 GND.n1784 GND.n1468 161.3
R7379 GND.n1783 GND.n1782 161.3
R7380 GND.n1781 GND.n1469 161.3
R7381 GND.n1780 GND.n1779 161.3
R7382 GND.n1778 GND.n1470 161.3
R7383 GND.n1777 GND.n1776 161.3
R7384 GND.n1775 GND.n1471 161.3
R7385 GND.n1439 GND.n1437 161.3
R7386 GND.n1874 GND.n1873 161.3
R7387 GND.n4239 GND.t192 157.496
R7388 GND.n2892 GND.t108 157.496
R7389 GND.n3106 GND.t155 153.965
R7390 GND.n18 GND.t40 153.582
R7391 GND.n33 GND.t51 153.582
R7392 GND.n49 GND.t50 153.582
R7393 GND.n3 GND.t57 153.582
R7394 GND.n79 GND.t71 153.582
R7395 GND.n94 GND.t213 153.582
R7396 GND.n110 GND.t204 153.582
R7397 GND.n126 GND.t53 153.582
R7398 GND.n3115 GND.n3114 152.776
R7399 GND.n3971 GND.n3961 152
R7400 GND.n3973 GND.n3972 152
R7401 GND.n3113 GND.n3104 152
R7402 GND.n4284 GND.t5 149.524
R7403 GND.n2844 GND.t206 149.524
R7404 GND.n1891 GND.t9 149.524
R7405 GND.n6077 GND.t42 149.524
R7406 GND.n5789 GND.n3185 143.351
R7407 GND.n5789 GND.n5788 143.351
R7408 GND.n3938 GND.n3937 141.77
R7409 GND.n3189 GND.n3188 141.77
R7410 GND.n3945 GND.n3944 141.77
R7411 GND.n3174 GND.n3173 141.77
R7412 GND.n3968 GND.t135 137.107
R7413 GND.n1400 GND.t127 126.772
R7414 GND.n1415 GND.t145 126.772
R7415 GND.n1431 GND.t185 126.772
R7416 GND.n1921 GND.t154 126.772
R7417 GND.n2180 GND.t159 126.772
R7418 GND.n3082 GND.t197 126.772
R7419 GND.n5801 GND.t167 126.772
R7420 GND.n5814 GND.t150 126.772
R7421 GND.n313 GND.t182 126.772
R7422 GND.n300 GND.t188 126.772
R7423 GND.n289 GND.t123 126.772
R7424 GND.n6259 GND.t201 126.772
R7425 GND.n6114 GND.t100 126.772
R7426 GND.n1258 GND.t164 126.772
R7427 GND.n1272 GND.t147 126.772
R7428 GND.n1285 GND.t112 126.772
R7429 GND.n3972 GND.t175 126.766
R7430 GND.n3970 GND.t114 126.766
R7431 GND.n3969 GND.t193 126.766
R7432 GND.n3105 GND.t117 126.766
R7433 GND.n3112 GND.t172 126.766
R7434 GND.n3114 GND.t128 126.766
R7435 GND.n21 GND.n20 104.615
R7436 GND.n36 GND.n35 104.615
R7437 GND.n52 GND.n51 104.615
R7438 GND.n6 GND.n5 104.615
R7439 GND.n1910 GND.n1909 104.615
R7440 GND.n1909 GND.n1883 104.615
R7441 GND.n1902 GND.n1883 104.615
R7442 GND.n1902 GND.n1901 104.615
R7443 GND.n1901 GND.n1887 104.615
R7444 GND.n1894 GND.n1887 104.615
R7445 GND.n1894 GND.n1893 104.615
R7446 GND.n4287 GND.n4286 104.615
R7447 GND.n4287 GND.n4280 104.615
R7448 GND.n4294 GND.n4280 104.615
R7449 GND.n4295 GND.n4294 104.615
R7450 GND.n4295 GND.n4276 104.615
R7451 GND.n4302 GND.n4276 104.615
R7452 GND.n4303 GND.n4302 104.615
R7453 GND.n2847 GND.n2846 104.615
R7454 GND.n2847 GND.n2840 104.615
R7455 GND.n2854 GND.n2840 104.615
R7456 GND.n2855 GND.n2854 104.615
R7457 GND.n2855 GND.n2836 104.615
R7458 GND.n2862 GND.n2836 104.615
R7459 GND.n2863 GND.n2862 104.615
R7460 GND.n82 GND.n81 104.615
R7461 GND.n97 GND.n96 104.615
R7462 GND.n113 GND.n112 104.615
R7463 GND.n129 GND.n128 104.615
R7464 GND.n6096 GND.n6095 104.615
R7465 GND.n6095 GND.n6069 104.615
R7466 GND.n6088 GND.n6069 104.615
R7467 GND.n6088 GND.n6087 104.615
R7468 GND.n6087 GND.n6073 104.615
R7469 GND.n6080 GND.n6073 104.615
R7470 GND.n6080 GND.n6079 104.615
R7471 GND.n374 GND.n277 99.6594
R7472 GND.n372 GND.n276 99.6594
R7473 GND.n368 GND.n275 99.6594
R7474 GND.n364 GND.n274 99.6594
R7475 GND.n356 GND.n273 99.6594
R7476 GND.n354 GND.n272 99.6594
R7477 GND.n350 GND.n271 99.6594
R7478 GND.n346 GND.n270 99.6594
R7479 GND.n342 GND.n269 99.6594
R7480 GND.n302 GND.n268 99.6594
R7481 GND.n334 GND.n267 99.6594
R7482 GND.n330 GND.n266 99.6594
R7483 GND.n326 GND.n265 99.6594
R7484 GND.n322 GND.n264 99.6594
R7485 GND.n318 GND.n263 99.6594
R7486 GND.n262 GND.n251 99.6594
R7487 GND.n6511 GND.n6510 99.6594
R7488 GND.n6505 GND.n3046 99.6594
R7489 GND.n6502 GND.n3047 99.6594
R7490 GND.n6498 GND.n3048 99.6594
R7491 GND.n6494 GND.n3049 99.6594
R7492 GND.n6490 GND.n3050 99.6594
R7493 GND.n6486 GND.n3051 99.6594
R7494 GND.n6483 GND.n3052 99.6594
R7495 GND.n6480 GND.n3053 99.6594
R7496 GND.n6476 GND.n3054 99.6594
R7497 GND.n6472 GND.n3055 99.6594
R7498 GND.n6469 GND.n3056 99.6594
R7499 GND.n6465 GND.n3057 99.6594
R7500 GND.n6461 GND.n3058 99.6594
R7501 GND.n6457 GND.n3059 99.6594
R7502 GND.n5812 GND.n3060 99.6594
R7503 GND.n6275 GND.n6273 99.6594
R7504 GND.n6281 GND.n6265 99.6594
R7505 GND.n6285 GND.n6283 99.6594
R7506 GND.n6291 GND.n6261 99.6594
R7507 GND.n6294 GND.n6293 99.6594
R7508 GND.n5822 GND.n3061 99.6594
R7509 GND.n6129 GND.n3062 99.6594
R7510 GND.n6125 GND.n3063 99.6594
R7511 GND.n6121 GND.n3064 99.6594
R7512 GND.n6117 GND.n3065 99.6594
R7513 GND.n1925 GND.n1389 99.6594
R7514 GND.n1927 GND.n1926 99.6594
R7515 GND.n1928 GND.n1394 99.6594
R7516 GND.n1930 GND.n1929 99.6594
R7517 GND.n1931 GND.n1401 99.6594
R7518 GND.n1933 GND.n1932 99.6594
R7519 GND.n6985 GND.n6984 99.6594
R7520 GND.n6983 GND.n1412 99.6594
R7521 GND.n6982 GND.n6981 99.6594
R7522 GND.n6980 GND.n1419 99.6594
R7523 GND.n6979 GND.n6978 99.6594
R7524 GND.n6977 GND.n1424 99.6594
R7525 GND.n6976 GND.n6975 99.6594
R7526 GND.n6974 GND.n1429 99.6594
R7527 GND.n6973 GND.n1379 99.6594
R7528 GND.n7178 GND.n7177 99.6594
R7529 GND.n7172 GND.n1222 99.6594
R7530 GND.n7169 GND.n1223 99.6594
R7531 GND.n7165 GND.n1224 99.6594
R7532 GND.n7161 GND.n1225 99.6594
R7533 GND.n7157 GND.n1226 99.6594
R7534 GND.n7153 GND.n1227 99.6594
R7535 GND.n7149 GND.n1228 99.6594
R7536 GND.n7145 GND.n1229 99.6594
R7537 GND.n7141 GND.n1230 99.6594
R7538 GND.n7137 GND.n1231 99.6594
R7539 GND.n7134 GND.n1232 99.6594
R7540 GND.n7130 GND.n1233 99.6594
R7541 GND.n7126 GND.n1234 99.6594
R7542 GND.n7122 GND.n1235 99.6594
R7543 GND.n1283 GND.n1236 99.6594
R7544 GND.n1942 GND.n1936 99.6594
R7545 GND.n1946 GND.n1937 99.6594
R7546 GND.n1950 GND.n1938 99.6594
R7547 GND.n1955 GND.n1954 99.6594
R7548 GND.n6989 GND.n6988 99.6594
R7549 GND.n1293 GND.n1237 99.6594
R7550 GND.n2193 GND.n1238 99.6594
R7551 GND.n2187 GND.n1239 99.6594
R7552 GND.n2201 GND.n1240 99.6594
R7553 GND.n2183 GND.n1241 99.6594
R7554 GND.n2192 GND.n1237 99.6594
R7555 GND.n2186 GND.n1238 99.6594
R7556 GND.n2200 GND.n1239 99.6594
R7557 GND.n2182 GND.n1240 99.6594
R7558 GND.n2178 GND.n1241 99.6594
R7559 GND.n6988 GND.n1923 99.6594
R7560 GND.n1955 GND.n1951 99.6594
R7561 GND.n1947 GND.n1938 99.6594
R7562 GND.n1943 GND.n1937 99.6594
R7563 GND.n1939 GND.n1936 99.6594
R7564 GND.n7178 GND.n1245 99.6594
R7565 GND.n7170 GND.n1222 99.6594
R7566 GND.n7166 GND.n1223 99.6594
R7567 GND.n7162 GND.n1224 99.6594
R7568 GND.n7158 GND.n1225 99.6594
R7569 GND.n7154 GND.n1226 99.6594
R7570 GND.n7150 GND.n1227 99.6594
R7571 GND.n7146 GND.n1228 99.6594
R7572 GND.n7142 GND.n1229 99.6594
R7573 GND.n1269 GND.n1230 99.6594
R7574 GND.n7135 GND.n1231 99.6594
R7575 GND.n7131 GND.n1232 99.6594
R7576 GND.n7127 GND.n1233 99.6594
R7577 GND.n7123 GND.n1234 99.6594
R7578 GND.n1282 GND.n1235 99.6594
R7579 GND.n7115 GND.n1236 99.6594
R7580 GND.n6973 GND.n1433 99.6594
R7581 GND.n6974 GND.n1428 99.6594
R7582 GND.n6976 GND.n1425 99.6594
R7583 GND.n6977 GND.n1423 99.6594
R7584 GND.n6979 GND.n1420 99.6594
R7585 GND.n6980 GND.n1418 99.6594
R7586 GND.n6982 GND.n1413 99.6594
R7587 GND.n6983 GND.n1411 99.6594
R7588 GND.n6985 GND.n1408 99.6594
R7589 GND.n6986 GND.n1406 99.6594
R7590 GND.n1934 GND.n1405 99.6594
R7591 GND.n1933 GND.n1402 99.6594
R7592 GND.n1931 GND.n1398 99.6594
R7593 GND.n1930 GND.n1395 99.6594
R7594 GND.n1928 GND.n1393 99.6594
R7595 GND.n1927 GND.n1390 99.6594
R7596 GND.n1925 GND.n1385 99.6594
R7597 GND.n6130 GND.n3061 99.6594
R7598 GND.n6126 GND.n3062 99.6594
R7599 GND.n6122 GND.n3063 99.6594
R7600 GND.n6118 GND.n3064 99.6594
R7601 GND.n6112 GND.n3065 99.6594
R7602 GND.n6293 GND.n6292 99.6594
R7603 GND.n6284 GND.n6261 99.6594
R7604 GND.n6283 GND.n6282 99.6594
R7605 GND.n6274 GND.n6265 99.6594
R7606 GND.n6273 GND.n6272 99.6594
R7607 GND.n6511 GND.n3069 99.6594
R7608 GND.n6503 GND.n3046 99.6594
R7609 GND.n6499 GND.n3047 99.6594
R7610 GND.n6495 GND.n3048 99.6594
R7611 GND.n6491 GND.n3049 99.6594
R7612 GND.n6487 GND.n3050 99.6594
R7613 GND.n5791 GND.n3051 99.6594
R7614 GND.n6481 GND.n3052 99.6594
R7615 GND.n6477 GND.n3053 99.6594
R7616 GND.n5798 GND.n3054 99.6594
R7617 GND.n6470 GND.n3055 99.6594
R7618 GND.n6466 GND.n3056 99.6594
R7619 GND.n6462 GND.n3057 99.6594
R7620 GND.n6458 GND.n3058 99.6594
R7621 GND.n5811 GND.n3059 99.6594
R7622 GND.n6450 GND.n3060 99.6594
R7623 GND.n317 GND.n262 99.6594
R7624 GND.n321 GND.n263 99.6594
R7625 GND.n325 GND.n264 99.6594
R7626 GND.n329 GND.n265 99.6594
R7627 GND.n333 GND.n266 99.6594
R7628 GND.n301 GND.n267 99.6594
R7629 GND.n341 GND.n268 99.6594
R7630 GND.n345 GND.n269 99.6594
R7631 GND.n349 GND.n270 99.6594
R7632 GND.n353 GND.n271 99.6594
R7633 GND.n357 GND.n272 99.6594
R7634 GND.n363 GND.n273 99.6594
R7635 GND.n367 GND.n274 99.6594
R7636 GND.n371 GND.n275 99.6594
R7637 GND.n375 GND.n276 99.6594
R7638 GND.n278 GND.n277 99.6594
R7639 GND.n3219 GND.n2829 99.6594
R7640 GND.n3221 GND.n2831 99.6594
R7641 GND.n3222 GND.n2874 99.6594
R7642 GND.n3224 GND.n2876 99.6594
R7643 GND.n3225 GND.n2879 99.6594
R7644 GND.n3227 GND.n2881 99.6594
R7645 GND.n3228 GND.n2884 99.6594
R7646 GND.n3230 GND.n2886 99.6594
R7647 GND.n3231 GND.n2889 99.6594
R7648 GND.n3232 GND.n2891 99.6594
R7649 GND.n3233 GND.n2897 99.6594
R7650 GND.n3233 GND.n2898 99.6594
R7651 GND.n3232 GND.n2896 99.6594
R7652 GND.n3231 GND.n2890 99.6594
R7653 GND.n3230 GND.n3229 99.6594
R7654 GND.n3228 GND.n2885 99.6594
R7655 GND.n3227 GND.n3226 99.6594
R7656 GND.n3225 GND.n2880 99.6594
R7657 GND.n3224 GND.n3223 99.6594
R7658 GND.n3222 GND.n2875 99.6594
R7659 GND.n3221 GND.n3220 99.6594
R7660 GND.n3219 GND.n2830 99.6594
R7661 GND.n4316 GND.n2665 99.6594
R7662 GND.n4216 GND.n3905 99.6594
R7663 GND.n4218 GND.n3906 99.6594
R7664 GND.n4222 GND.n3907 99.6594
R7665 GND.n4224 GND.n3908 99.6594
R7666 GND.n4228 GND.n3909 99.6594
R7667 GND.n4230 GND.n3910 99.6594
R7668 GND.n4234 GND.n3911 99.6594
R7669 GND.n4236 GND.n3912 99.6594
R7670 GND.n4243 GND.n3913 99.6594
R7671 GND.n4318 GND.n3904 99.6594
R7672 GND.n4316 GND.n4315 99.6594
R7673 GND.n4217 GND.n3905 99.6594
R7674 GND.n4221 GND.n3906 99.6594
R7675 GND.n4223 GND.n3907 99.6594
R7676 GND.n4227 GND.n3908 99.6594
R7677 GND.n4229 GND.n3909 99.6594
R7678 GND.n4233 GND.n3910 99.6594
R7679 GND.n4235 GND.n3911 99.6594
R7680 GND.n4242 GND.n3912 99.6594
R7681 GND.n4244 GND.n3913 99.6594
R7682 GND.n4319 GND.n4318 99.6594
R7683 GND.n1877 GND.n1876 85.6162
R7684 GND.n4311 GND.n4310 85.6161
R7685 GND.n2871 GND.n2870 85.6161
R7686 GND.n4240 GND.n4239 85.1399
R7687 GND.n2893 GND.n2892 85.1399
R7688 GND.n1879 GND.n1878 83.2531
R7689 GND.n6105 GND.n6104 83.2531
R7690 GND.n6102 GND.n6101 83.2531
R7691 GND.n4309 GND.n4308 83.253
R7692 GND.n2869 GND.n2868 83.253
R7693 GND.n7367 GND.n1035 81.3163
R7694 GND.n7367 GND.n7366 81.3163
R7695 GND.n7366 GND.n7365 81.3163
R7696 GND.n7365 GND.n1040 81.3163
R7697 GND.n7359 GND.n1040 81.3163
R7698 GND.n7359 GND.n7358 81.3163
R7699 GND.n7358 GND.n7357 81.3163
R7700 GND.n7357 GND.n1048 81.3163
R7701 GND.n7351 GND.n1048 81.3163
R7702 GND.n7351 GND.n7350 81.3163
R7703 GND.n7350 GND.n7349 81.3163
R7704 GND.n7349 GND.n1056 81.3163
R7705 GND.n7343 GND.n1056 81.3163
R7706 GND.n7343 GND.n7342 81.3163
R7707 GND.n7342 GND.n7341 81.3163
R7708 GND.n7341 GND.n1064 81.3163
R7709 GND.n7335 GND.n1064 81.3163
R7710 GND.n7335 GND.n7334 81.3163
R7711 GND.n7334 GND.n7333 81.3163
R7712 GND.n7333 GND.n1072 81.3163
R7713 GND.n7327 GND.n1072 81.3163
R7714 GND.n7327 GND.n7326 81.3163
R7715 GND.n7326 GND.n7325 81.3163
R7716 GND.n7325 GND.n1080 81.3163
R7717 GND.n7319 GND.n1080 81.3163
R7718 GND.n7319 GND.n7318 81.3163
R7719 GND.n7318 GND.n7317 81.3163
R7720 GND.n7317 GND.n1088 81.3163
R7721 GND.n7311 GND.n1088 81.3163
R7722 GND.n7311 GND.n7310 81.3163
R7723 GND.n7310 GND.n7309 81.3163
R7724 GND.n7309 GND.n1096 81.3163
R7725 GND.n7303 GND.n1096 81.3163
R7726 GND.n7303 GND.n7302 81.3163
R7727 GND.n7302 GND.n7301 81.3163
R7728 GND.n7301 GND.n1104 81.3163
R7729 GND.n7295 GND.n1104 81.3163
R7730 GND.n7295 GND.n7294 81.3163
R7731 GND.n7294 GND.n7293 81.3163
R7732 GND.n7293 GND.n1112 81.3163
R7733 GND.n7287 GND.n1112 81.3163
R7734 GND.n7287 GND.n7286 81.3163
R7735 GND.n7286 GND.n7285 81.3163
R7736 GND.n7285 GND.n1120 81.3163
R7737 GND.n7279 GND.n1120 81.3163
R7738 GND.n7279 GND.n7278 81.3163
R7739 GND.n7278 GND.n7277 81.3163
R7740 GND.n7277 GND.n1128 81.3163
R7741 GND.n7271 GND.n1128 81.3163
R7742 GND.n7271 GND.n7270 81.3163
R7743 GND.n7270 GND.n7269 81.3163
R7744 GND.n7269 GND.n1136 81.3163
R7745 GND.n7263 GND.n1136 81.3163
R7746 GND.n7263 GND.n7262 81.3163
R7747 GND.n7262 GND.n7261 81.3163
R7748 GND.n7261 GND.n1144 81.3163
R7749 GND.n7255 GND.n1144 81.3163
R7750 GND.n7255 GND.n7254 81.3163
R7751 GND.n7254 GND.n7253 81.3163
R7752 GND.n7253 GND.n1152 81.3163
R7753 GND.n7247 GND.n1152 81.3163
R7754 GND.n7247 GND.n7246 81.3163
R7755 GND.n7246 GND.n7245 81.3163
R7756 GND.n7245 GND.n1160 81.3163
R7757 GND.n7239 GND.n1160 81.3163
R7758 GND.n7239 GND.n7238 81.3163
R7759 GND.n7238 GND.n7237 81.3163
R7760 GND.n7237 GND.n1168 81.3163
R7761 GND.n7231 GND.n1168 81.3163
R7762 GND.n7231 GND.n7230 81.3163
R7763 GND.n7230 GND.n7229 81.3163
R7764 GND.n7229 GND.n1176 81.3163
R7765 GND.n68 GND.t21 78.6894
R7766 GND.n71 GND.t7 77.1283
R7767 GND.n70 GND.t209 77.1283
R7768 GND.n69 GND.t61 77.1283
R7769 GND.n68 GND.t59 77.1283
R7770 GND.n6056 GND.t234 76.2463
R7771 GND.n6060 GND.t216 76.2451
R7772 GND.n75 GND.n73 75.5577
R7773 GND.n90 GND.n88 75.5577
R7774 GND.n106 GND.n104 75.5577
R7775 GND.n122 GND.n120 75.5577
R7776 GND.n3968 GND.n3967 74.9819
R7777 GND.n27 GND.n26 74.3939
R7778 GND.n29 GND.n28 74.3939
R7779 GND.n42 GND.n41 74.3939
R7780 GND.n44 GND.n43 74.3939
R7781 GND.n58 GND.n57 74.3939
R7782 GND.n60 GND.n59 74.3939
R7783 GND.n12 GND.n11 74.3939
R7784 GND.n14 GND.n13 74.3939
R7785 GND.n75 GND.n74 74.3939
R7786 GND.n90 GND.n89 74.3939
R7787 GND.n106 GND.n105 74.3939
R7788 GND.n122 GND.n121 74.3939
R7789 GND.n6059 GND.t214 73.6933
R7790 GND.n6058 GND.t220 73.6933
R7791 GND.n6057 GND.t235 73.6933
R7792 GND.n6056 GND.t237 73.6933
R7793 GND.n6063 GND.t221 73.6921
R7794 GND.n6062 GND.t224 73.6921
R7795 GND.n6061 GND.t217 73.6921
R7796 GND.n6060 GND.t219 73.6921
R7797 GND.n3969 GND.n3963 72.8411
R7798 GND.n3970 GND.n3962 72.8411
R7799 GND.n3112 GND.n3111 72.8411
R7800 GND.n4240 GND.t191 72.3569
R7801 GND.n2893 GND.t109 72.3569
R7802 GND.n3120 GND.n3119 71.676
R7803 GND.n3121 GND.n3102 71.676
R7804 GND.n3128 GND.n3127 71.676
R7805 GND.n3129 GND.n3100 71.676
R7806 GND.n3136 GND.n3135 71.676
R7807 GND.n3137 GND.n3098 71.676
R7808 GND.n3144 GND.n3143 71.676
R7809 GND.n3145 GND.n3096 71.676
R7810 GND.n3152 GND.n3151 71.676
R7811 GND.n3153 GND.n3094 71.676
R7812 GND.n3160 GND.n3159 71.676
R7813 GND.n3161 GND.n3092 71.676
R7814 GND.n3168 GND.n3167 71.676
R7815 GND.n3169 GND.n3090 71.676
R7816 GND.n3179 GND.n3178 71.676
R7817 GND.n3183 GND.n3088 71.676
R7818 GND.n5788 GND.n5787 71.676
R7819 GND.n5785 GND.n5784 71.676
R7820 GND.n5779 GND.n3191 71.676
R7821 GND.n5777 GND.n5776 71.676
R7822 GND.n5772 GND.n3194 71.676
R7823 GND.n5770 GND.n5769 71.676
R7824 GND.n5765 GND.n3197 71.676
R7825 GND.n5763 GND.n5762 71.676
R7826 GND.n5758 GND.n3200 71.676
R7827 GND.n5756 GND.n5755 71.676
R7828 GND.n5751 GND.n3203 71.676
R7829 GND.n5749 GND.n5748 71.676
R7830 GND.n5744 GND.n3206 71.676
R7831 GND.n5742 GND.n5741 71.676
R7832 GND.n5737 GND.n3209 71.676
R7833 GND.n5735 GND.n5734 71.676
R7834 GND.n5730 GND.n5726 71.676
R7835 GND.n3977 GND.n3976 71.676
R7836 GND.n3983 GND.n3982 71.676
R7837 GND.n3986 GND.n3985 71.676
R7838 GND.n3991 GND.n3990 71.676
R7839 GND.n3994 GND.n3993 71.676
R7840 GND.n3999 GND.n3998 71.676
R7841 GND.n4002 GND.n4001 71.676
R7842 GND.n4007 GND.n4006 71.676
R7843 GND.n4010 GND.n4009 71.676
R7844 GND.n4015 GND.n4014 71.676
R7845 GND.n4018 GND.n4017 71.676
R7846 GND.n4023 GND.n4022 71.676
R7847 GND.n4026 GND.n4025 71.676
R7848 GND.n4031 GND.n4030 71.676
R7849 GND.n4034 GND.n4033 71.676
R7850 GND.n4039 GND.n4038 71.676
R7851 GND.n4042 GND.n4041 71.676
R7852 GND.n4045 GND.n4044 71.676
R7853 GND.n4050 GND.n4049 71.676
R7854 GND.n4053 GND.n4052 71.676
R7855 GND.n4058 GND.n4057 71.676
R7856 GND.n4061 GND.n4060 71.676
R7857 GND.n4066 GND.n4065 71.676
R7858 GND.n4069 GND.n4068 71.676
R7859 GND.n4074 GND.n4073 71.676
R7860 GND.n4077 GND.n4076 71.676
R7861 GND.n4082 GND.n4081 71.676
R7862 GND.n4085 GND.n4084 71.676
R7863 GND.n4090 GND.n4089 71.676
R7864 GND.n4093 GND.n4092 71.676
R7865 GND.n4098 GND.n4097 71.676
R7866 GND.n4101 GND.n4100 71.676
R7867 GND.n4106 GND.n4105 71.676
R7868 GND.n3978 GND.n3977 71.676
R7869 GND.n3984 GND.n3983 71.676
R7870 GND.n3985 GND.n3958 71.676
R7871 GND.n3992 GND.n3991 71.676
R7872 GND.n3993 GND.n3956 71.676
R7873 GND.n4000 GND.n3999 71.676
R7874 GND.n4001 GND.n3954 71.676
R7875 GND.n4008 GND.n4007 71.676
R7876 GND.n4009 GND.n3952 71.676
R7877 GND.n4016 GND.n4015 71.676
R7878 GND.n4017 GND.n3950 71.676
R7879 GND.n4024 GND.n4023 71.676
R7880 GND.n4025 GND.n3948 71.676
R7881 GND.n4032 GND.n4031 71.676
R7882 GND.n4033 GND.n3943 71.676
R7883 GND.n4040 GND.n4039 71.676
R7884 GND.n4043 GND.n4042 71.676
R7885 GND.n4044 GND.n3941 71.676
R7886 GND.n4051 GND.n4050 71.676
R7887 GND.n4052 GND.n3936 71.676
R7888 GND.n4059 GND.n4058 71.676
R7889 GND.n4060 GND.n3934 71.676
R7890 GND.n4067 GND.n4066 71.676
R7891 GND.n4068 GND.n3932 71.676
R7892 GND.n4075 GND.n4074 71.676
R7893 GND.n4076 GND.n3930 71.676
R7894 GND.n4083 GND.n4082 71.676
R7895 GND.n4084 GND.n3928 71.676
R7896 GND.n4091 GND.n4090 71.676
R7897 GND.n4092 GND.n3926 71.676
R7898 GND.n4099 GND.n4098 71.676
R7899 GND.n4100 GND.n3924 71.676
R7900 GND.n4107 GND.n4106 71.676
R7901 GND.n5726 GND.n3210 71.676
R7902 GND.n5736 GND.n5735 71.676
R7903 GND.n3209 GND.n3207 71.676
R7904 GND.n5743 GND.n5742 71.676
R7905 GND.n3206 GND.n3204 71.676
R7906 GND.n5750 GND.n5749 71.676
R7907 GND.n3203 GND.n3201 71.676
R7908 GND.n5757 GND.n5756 71.676
R7909 GND.n3200 GND.n3198 71.676
R7910 GND.n5764 GND.n5763 71.676
R7911 GND.n3197 GND.n3195 71.676
R7912 GND.n5771 GND.n5770 71.676
R7913 GND.n3194 GND.n3192 71.676
R7914 GND.n5778 GND.n5777 71.676
R7915 GND.n3191 GND.n3187 71.676
R7916 GND.n5786 GND.n5785 71.676
R7917 GND.n3185 GND.n3184 71.676
R7918 GND.n3180 GND.n3088 71.676
R7919 GND.n3178 GND.n3177 71.676
R7920 GND.n3170 GND.n3169 71.676
R7921 GND.n3167 GND.n3166 71.676
R7922 GND.n3162 GND.n3161 71.676
R7923 GND.n3159 GND.n3158 71.676
R7924 GND.n3154 GND.n3153 71.676
R7925 GND.n3151 GND.n3150 71.676
R7926 GND.n3146 GND.n3145 71.676
R7927 GND.n3143 GND.n3142 71.676
R7928 GND.n3138 GND.n3137 71.676
R7929 GND.n3135 GND.n3134 71.676
R7930 GND.n3130 GND.n3129 71.676
R7931 GND.n3127 GND.n3126 71.676
R7932 GND.n3122 GND.n3121 71.676
R7933 GND.n3119 GND.n3118 71.676
R7934 GND.n4309 GND.n4307 70.6332
R7935 GND.n2869 GND.n2867 70.6332
R7936 GND.n6102 GND.n6100 70.6332
R7937 GND.n1915 GND.n1914 67.4823
R7938 GND.n3974 GND.n3973 62.8652
R7939 GND.n3939 GND.n3938 59.5399
R7940 GND.n5781 GND.n3189 59.5399
R7941 GND.n3946 GND.n3945 59.5399
R7942 GND.n3175 GND.n3174 59.5399
R7943 GND.n3111 GND.n3106 59.441
R7944 GND.n1562 GND.n1561 58.7165
R7945 GND.n1542 GND.n1541 58.7165
R7946 GND.n1584 GND.n1583 58.7165
R7947 GND.n1564 GND.n1563 58.7165
R7948 GND.n1856 GND.n1855 58.7165
R7949 GND.n1836 GND.n1835 58.7165
R7950 GND.n1586 GND.n1585 58.7165
R7951 GND.n1857 GND.n1444 58.7165
R7952 GND.n1774 GND.n1773 58.2272
R7953 GND.n1833 GND.n1832 58.2272
R7954 GND.n1713 GND.n1712 58.2272
R7955 GND.n1772 GND.n1771 58.2272
R7956 GND.n1652 GND.n1651 58.2272
R7957 GND.n1711 GND.n1710 58.2272
R7958 GND.n1591 GND.n1590 58.2272
R7959 GND.n1650 GND.n1649 58.2272
R7960 GND.n1782 GND.n1468 56.5193
R7961 GND.n1824 GND.n1456 56.5193
R7962 GND.n1721 GND.n1487 56.5193
R7963 GND.n1763 GND.n1475 56.5193
R7964 GND.n1660 GND.n1506 56.5193
R7965 GND.n1702 GND.n1494 56.5193
R7966 GND.n1599 GND.n1525 56.5193
R7967 GND.n1641 GND.n1513 56.5193
R7968 GND.n1553 GND.n1538 56.5193
R7969 GND.n1575 GND.n1532 56.5193
R7970 GND.n1847 GND.n1448 56.5193
R7971 GND.n1867 GND.n1866 56.5193
R7972 GND.n1400 GND.n1399 52.3641
R7973 GND.n1415 GND.n1414 52.3641
R7974 GND.n1431 GND.n1430 52.3641
R7975 GND.n1921 GND.n1920 52.3641
R7976 GND.n2180 GND.n2179 52.3641
R7977 GND.n3082 GND.n3081 52.3641
R7978 GND.n5801 GND.n5800 52.3641
R7979 GND.n5814 GND.n5813 52.3641
R7980 GND.n313 GND.n312 52.3641
R7981 GND.n300 GND.n299 52.3641
R7982 GND.n289 GND.n288 52.3641
R7983 GND.n6259 GND.n6258 52.3641
R7984 GND.n6114 GND.n6113 52.3641
R7985 GND.n1258 GND.n1257 52.3641
R7986 GND.n1272 GND.n1271 52.3641
R7987 GND.n1285 GND.n1284 52.3641
R7988 GND.n20 GND.t40 52.3082
R7989 GND.n35 GND.t51 52.3082
R7990 GND.n51 GND.t50 52.3082
R7991 GND.n5 GND.t57 52.3082
R7992 GND.n1893 GND.t9 52.3082
R7993 GND.n4286 GND.t5 52.3082
R7994 GND.n2846 GND.t206 52.3082
R7995 GND.n81 GND.t71 52.3082
R7996 GND.n96 GND.t213 52.3082
R7997 GND.n112 GND.t204 52.3082
R7998 GND.n128 GND.t53 52.3082
R7999 GND.n6079 GND.t42 52.3082
R8000 GND.n3970 GND.n3969 48.2005
R8001 GND.n3112 GND.n3105 48.2005
R8002 GND.n3116 GND.n3115 44.3322
R8003 GND.n4241 GND.n4240 42.2793
R8004 GND.n7026 GND.n1400 42.2793
R8005 GND.n1416 GND.n1415 42.2793
R8006 GND.n6995 GND.n1431 42.2793
R8007 GND.n1922 GND.n1921 42.2793
R8008 GND.n2207 GND.n2180 42.2793
R8009 GND.n6493 GND.n3082 42.2793
R8010 GND.n6474 GND.n5801 42.2793
R8011 GND.n5815 GND.n5814 42.2793
R8012 GND.n316 GND.n313 42.2793
R8013 GND.n339 GND.n300 42.2793
R8014 GND.n362 GND.n289 42.2793
R8015 GND.n6260 GND.n6259 42.2793
R8016 GND.n6115 GND.n6114 42.2793
R8017 GND.n7160 GND.n1258 42.2793
R8018 GND.n7139 GND.n1272 42.2793
R8019 GND.n1286 GND.n1285 42.2793
R8020 GND.n2894 GND.n2893 42.2793
R8021 GND.n3967 GND.n3966 41.6274
R8022 GND.n3110 GND.n3109 41.6274
R8023 GND.n1801 GND.n1462 40.4934
R8024 GND.n1805 GND.n1462 40.4934
R8025 GND.n1740 GND.n1481 40.4934
R8026 GND.n1744 GND.n1481 40.4934
R8027 GND.n1679 GND.n1500 40.4934
R8028 GND.n1683 GND.n1500 40.4934
R8029 GND.n1618 GND.n1519 40.4934
R8030 GND.n1622 GND.n1519 40.4934
R8031 GND.n27 GND.n25 38.0037
R8032 GND.n42 GND.n40 38.0037
R8033 GND.n58 GND.n56 38.0037
R8034 GND.n12 GND.n10 38.0037
R8035 GND.n87 GND.n86 36.8399
R8036 GND.n102 GND.n101 36.8399
R8037 GND.n118 GND.n117 36.8399
R8038 GND.n134 GND.n133 36.8399
R8039 GND.n3969 GND.n3968 36.5361
R8040 GND.n7221 GND.n7220 33.0981
R8041 GND.n7220 GND.n7219 33.0981
R8042 GND.n7219 GND.n1183 33.0981
R8043 GND.n7213 GND.n1183 33.0981
R8044 GND.n7213 GND.n7212 33.0981
R8045 GND.n7212 GND.n7211 33.0981
R8046 GND.n7211 GND.n1190 33.0981
R8047 GND.n7205 GND.n1190 33.0981
R8048 GND.n7205 GND.n7204 33.0981
R8049 GND.n7204 GND.n7203 33.0981
R8050 GND.n7203 GND.n1198 33.0981
R8051 GND.n7197 GND.n1198 33.0981
R8052 GND.n7197 GND.n7196 33.0981
R8053 GND.n7196 GND.n7195 33.0981
R8054 GND.n7195 GND.n1206 33.0981
R8055 GND.n7189 GND.n1206 33.0981
R8056 GND.n7189 GND.n7188 33.0981
R8057 GND.n7188 GND.n7187 33.0981
R8058 GND.n7187 GND.n1214 33.0981
R8059 GND.n7181 GND.n1214 33.0981
R8060 GND.n7181 GND.n7180 33.0981
R8061 GND.n1290 GND.n1243 33.0981
R8062 GND.n1924 GND.n1382 33.0981
R8063 GND.n6972 GND.n1956 33.0981
R8064 GND.n6966 GND.n1956 33.0981
R8065 GND.n6966 GND.n6965 33.0981
R8066 GND.n6965 GND.n6964 33.0981
R8067 GND.n6520 GND.n6519 33.0981
R8068 GND.n6519 GND.n3038 33.0981
R8069 GND.n6513 GND.n3038 33.0981
R8070 GND.n5819 GND.n3067 33.0981
R8071 GND.n8445 GND.n253 33.0981
R8072 GND.n8439 GND.n8438 33.0981
R8073 GND.n8438 GND.n8437 33.0981
R8074 GND.n8437 GND.n384 33.0981
R8075 GND.n8431 GND.n384 33.0981
R8076 GND.n8431 GND.n8430 33.0981
R8077 GND.n8430 GND.n8429 33.0981
R8078 GND.n8429 GND.n392 33.0981
R8079 GND.n8423 GND.n392 33.0981
R8080 GND.n8423 GND.n8422 33.0981
R8081 GND.n8422 GND.n8421 33.0981
R8082 GND.n8421 GND.n400 33.0981
R8083 GND.n8415 GND.n400 33.0981
R8084 GND.n8415 GND.n8414 33.0981
R8085 GND.n8414 GND.n8413 33.0981
R8086 GND.n8413 GND.n408 33.0981
R8087 GND.n8407 GND.n408 33.0981
R8088 GND.n8407 GND.n8406 33.0981
R8089 GND.n8406 GND.n8405 33.0981
R8090 GND.n8405 GND.n416 33.0981
R8091 GND.n8399 GND.n416 33.0981
R8092 GND.n8399 GND.n8398 33.0981
R8093 GND.n5731 GND.n5725 32.6249
R8094 GND.n4110 GND.n3922 32.6249
R8095 GND.n2538 GND.n2530 32.1052
R8096 GND.n5727 GND.n3037 32.1052
R8097 GND.n7020 GND.n1407 30.6565
R8098 GND.n6485 GND.n5790 30.6565
R8099 GND.t129 GND.n6520 29.1264
R8100 GND.n3971 GND.n3970 27.0217
R8101 GND.n3113 GND.n3112 27.0217
R8102 GND.n3963 GND.n3962 25.8289
R8103 GND.n6987 GND.n6972 25.1547
R8104 GND.n6513 GND.n6512 25.1547
R8105 GND.n1776 GND.n1775 24.4675
R8106 GND.n1776 GND.n1470 24.4675
R8107 GND.n1780 GND.n1470 24.4675
R8108 GND.n1781 GND.n1780 24.4675
R8109 GND.n1782 GND.n1781 24.4675
R8110 GND.n1786 GND.n1468 24.4675
R8111 GND.n1787 GND.n1786 24.4675
R8112 GND.n1788 GND.n1787 24.4675
R8113 GND.n1788 GND.n1466 24.4675
R8114 GND.n1792 GND.n1466 24.4675
R8115 GND.n1795 GND.n1794 24.4675
R8116 GND.n1795 GND.n1464 24.4675
R8117 GND.n1799 GND.n1464 24.4675
R8118 GND.n1800 GND.n1799 24.4675
R8119 GND.n1801 GND.n1800 24.4675
R8120 GND.n1806 GND.n1805 24.4675
R8121 GND.n1807 GND.n1806 24.4675
R8122 GND.n1807 GND.n1460 24.4675
R8123 GND.n1811 GND.n1460 24.4675
R8124 GND.n1812 GND.n1811 24.4675
R8125 GND.n1814 GND.n1458 24.4675
R8126 GND.n1818 GND.n1458 24.4675
R8127 GND.n1819 GND.n1818 24.4675
R8128 GND.n1820 GND.n1819 24.4675
R8129 GND.n1820 GND.n1456 24.4675
R8130 GND.n1825 GND.n1824 24.4675
R8131 GND.n1826 GND.n1825 24.4675
R8132 GND.n1826 GND.n1454 24.4675
R8133 GND.n1830 GND.n1454 24.4675
R8134 GND.n1831 GND.n1830 24.4675
R8135 GND.n1715 GND.n1714 24.4675
R8136 GND.n1715 GND.n1489 24.4675
R8137 GND.n1719 GND.n1489 24.4675
R8138 GND.n1720 GND.n1719 24.4675
R8139 GND.n1721 GND.n1720 24.4675
R8140 GND.n1725 GND.n1487 24.4675
R8141 GND.n1726 GND.n1725 24.4675
R8142 GND.n1727 GND.n1726 24.4675
R8143 GND.n1727 GND.n1485 24.4675
R8144 GND.n1731 GND.n1485 24.4675
R8145 GND.n1734 GND.n1733 24.4675
R8146 GND.n1734 GND.n1483 24.4675
R8147 GND.n1738 GND.n1483 24.4675
R8148 GND.n1739 GND.n1738 24.4675
R8149 GND.n1740 GND.n1739 24.4675
R8150 GND.n1745 GND.n1744 24.4675
R8151 GND.n1746 GND.n1745 24.4675
R8152 GND.n1746 GND.n1479 24.4675
R8153 GND.n1750 GND.n1479 24.4675
R8154 GND.n1751 GND.n1750 24.4675
R8155 GND.n1753 GND.n1477 24.4675
R8156 GND.n1757 GND.n1477 24.4675
R8157 GND.n1758 GND.n1757 24.4675
R8158 GND.n1759 GND.n1758 24.4675
R8159 GND.n1759 GND.n1475 24.4675
R8160 GND.n1764 GND.n1763 24.4675
R8161 GND.n1765 GND.n1764 24.4675
R8162 GND.n1765 GND.n1473 24.4675
R8163 GND.n1769 GND.n1473 24.4675
R8164 GND.n1770 GND.n1769 24.4675
R8165 GND.n1654 GND.n1653 24.4675
R8166 GND.n1654 GND.n1508 24.4675
R8167 GND.n1658 GND.n1508 24.4675
R8168 GND.n1659 GND.n1658 24.4675
R8169 GND.n1660 GND.n1659 24.4675
R8170 GND.n1664 GND.n1506 24.4675
R8171 GND.n1665 GND.n1664 24.4675
R8172 GND.n1666 GND.n1665 24.4675
R8173 GND.n1666 GND.n1504 24.4675
R8174 GND.n1670 GND.n1504 24.4675
R8175 GND.n1673 GND.n1672 24.4675
R8176 GND.n1673 GND.n1502 24.4675
R8177 GND.n1677 GND.n1502 24.4675
R8178 GND.n1678 GND.n1677 24.4675
R8179 GND.n1679 GND.n1678 24.4675
R8180 GND.n1684 GND.n1683 24.4675
R8181 GND.n1685 GND.n1684 24.4675
R8182 GND.n1685 GND.n1498 24.4675
R8183 GND.n1689 GND.n1498 24.4675
R8184 GND.n1690 GND.n1689 24.4675
R8185 GND.n1692 GND.n1496 24.4675
R8186 GND.n1696 GND.n1496 24.4675
R8187 GND.n1697 GND.n1696 24.4675
R8188 GND.n1698 GND.n1697 24.4675
R8189 GND.n1698 GND.n1494 24.4675
R8190 GND.n1703 GND.n1702 24.4675
R8191 GND.n1704 GND.n1703 24.4675
R8192 GND.n1704 GND.n1492 24.4675
R8193 GND.n1708 GND.n1492 24.4675
R8194 GND.n1709 GND.n1708 24.4675
R8195 GND.n1593 GND.n1592 24.4675
R8196 GND.n1593 GND.n1527 24.4675
R8197 GND.n1597 GND.n1527 24.4675
R8198 GND.n1598 GND.n1597 24.4675
R8199 GND.n1599 GND.n1598 24.4675
R8200 GND.n1603 GND.n1525 24.4675
R8201 GND.n1604 GND.n1603 24.4675
R8202 GND.n1605 GND.n1604 24.4675
R8203 GND.n1605 GND.n1523 24.4675
R8204 GND.n1609 GND.n1523 24.4675
R8205 GND.n1612 GND.n1611 24.4675
R8206 GND.n1612 GND.n1521 24.4675
R8207 GND.n1616 GND.n1521 24.4675
R8208 GND.n1617 GND.n1616 24.4675
R8209 GND.n1618 GND.n1617 24.4675
R8210 GND.n1623 GND.n1622 24.4675
R8211 GND.n1624 GND.n1623 24.4675
R8212 GND.n1624 GND.n1517 24.4675
R8213 GND.n1628 GND.n1517 24.4675
R8214 GND.n1629 GND.n1628 24.4675
R8215 GND.n1631 GND.n1515 24.4675
R8216 GND.n1635 GND.n1515 24.4675
R8217 GND.n1636 GND.n1635 24.4675
R8218 GND.n1637 GND.n1636 24.4675
R8219 GND.n1637 GND.n1513 24.4675
R8220 GND.n1642 GND.n1641 24.4675
R8221 GND.n1643 GND.n1642 24.4675
R8222 GND.n1643 GND.n1511 24.4675
R8223 GND.n1647 GND.n1511 24.4675
R8224 GND.n1648 GND.n1647 24.4675
R8225 GND.n1560 GND.n1559 24.4675
R8226 GND.n1559 GND.n1536 24.4675
R8227 GND.n1555 GND.n1536 24.4675
R8228 GND.n1555 GND.n1554 24.4675
R8229 GND.n1554 GND.n1553 24.4675
R8230 GND.n1549 GND.n1538 24.4675
R8231 GND.n1549 GND.n1548 24.4675
R8232 GND.n1548 GND.n1547 24.4675
R8233 GND.n1547 GND.n1540 24.4675
R8234 GND.n1543 GND.n1540 24.4675
R8235 GND.n1582 GND.n1581 24.4675
R8236 GND.n1581 GND.n1530 24.4675
R8237 GND.n1577 GND.n1530 24.4675
R8238 GND.n1577 GND.n1576 24.4675
R8239 GND.n1576 GND.n1575 24.4675
R8240 GND.n1571 GND.n1532 24.4675
R8241 GND.n1571 GND.n1570 24.4675
R8242 GND.n1570 GND.n1569 24.4675
R8243 GND.n1569 GND.n1534 24.4675
R8244 GND.n1565 GND.n1534 24.4675
R8245 GND.n1854 GND.n1853 24.4675
R8246 GND.n1853 GND.n1446 24.4675
R8247 GND.n1849 GND.n1446 24.4675
R8248 GND.n1849 GND.n1848 24.4675
R8249 GND.n1848 GND.n1847 24.4675
R8250 GND.n1843 GND.n1448 24.4675
R8251 GND.n1843 GND.n1842 24.4675
R8252 GND.n1842 GND.n1841 24.4675
R8253 GND.n1841 GND.n1450 24.4675
R8254 GND.n1837 GND.n1450 24.4675
R8255 GND.n1873 GND.n1439 24.4675
R8256 GND.n1873 GND.n1872 24.4675
R8257 GND.n1872 GND.n1871 24.4675
R8258 GND.n1871 GND.n1440 24.4675
R8259 GND.n1867 GND.n1440 24.4675
R8260 GND.n1866 GND.n1865 24.4675
R8261 GND.n1865 GND.n1442 24.4675
R8262 GND.n1861 GND.n1442 24.4675
R8263 GND.n1861 GND.n1860 24.4675
R8264 GND.n1860 GND.n1859 24.4675
R8265 GND.n1877 GND.n1875 24.2758
R8266 GND.n1589 GND.n1584 23.9365
R8267 GND.n7180 GND.n7179 23.8308
R8268 GND.n8439 GND.n383 23.8308
R8269 GND.n1835 GND.n1834 23.7319
R8270 GND.n6944 GND.n2558 22.5069
R8271 GND.n4134 GND.n2566 22.5069
R8272 GND.n4148 GND.n2583 22.5069
R8273 GND.n6916 GND.n2593 22.5069
R8274 GND.n4161 GND.n2601 22.5069
R8275 GND.n6896 GND.n2617 22.5069
R8276 GND.n4174 GND.n2627 22.5069
R8277 GND.n6882 GND.n2635 22.5069
R8278 GND.n4187 GND.n2645 22.5069
R8279 GND.n4210 GND.n2662 22.5069
R8280 GND.n5637 GND.n2905 22.5069
R8281 GND.n5651 GND.n2923 22.5069
R8282 GND.n6604 GND.n2933 22.5069
R8283 GND.n5664 GND.n2941 22.5069
R8284 GND.n6590 GND.n2951 22.5069
R8285 GND.n5677 GND.n2967 22.5069
R8286 GND.n6570 GND.n2975 22.5069
R8287 GND.n5690 GND.n2985 22.5069
R8288 GND.n5704 GND.n3002 22.5069
R8289 GND.n6542 GND.n3010 22.5069
R8290 GND.n5717 GND.n3020 22.5069
R8291 GND.n6528 GND.n3028 22.5069
R8292 GND.n1588 GND.n1586 22.4289
R8293 GND.n6958 GND.n2539 21.8449
R8294 GND.n6957 GND.t115 21.8449
R8295 GND.n4158 GND.n2609 21.8449
R8296 GND.n6902 GND.n2611 21.8449
R8297 GND.n6584 GND.n2957 21.8449
R8298 GND.n5674 GND.n2959 21.8449
R8299 GND.n6106 GND.n6105 21.4888
R8300 GND.n6930 GND.t89 21.183
R8301 GND.n6556 GND.t103 21.183
R8302 GND.n3972 GND.n3971 21.1793
R8303 GND.n3114 GND.n3113 21.1793
R8304 GND.n1541 GND.n1452 21.141
R8305 GND.n2872 GND.n2871 20.961
R8306 GND.n4312 GND.n4311 20.548
R8307 GND.n6951 GND.n6950 20.521
R8308 GND.n6910 GND.n2599 20.521
R8309 GND.n4171 GND.n2619 20.521
R8310 GND.n5661 GND.n2949 20.521
R8311 GND.n6576 GND.n2969 20.521
R8312 GND.n6535 GND.n6534 20.521
R8313 GND.n3974 GND.n2543 20.4493
R8314 GND.n3116 GND.n3025 20.4493
R8315 GND.n3964 GND.t195 19.8005
R8316 GND.n3964 GND.t137 19.8005
R8317 GND.n3965 GND.t177 19.8005
R8318 GND.n3965 GND.t116 19.8005
R8319 GND.n3107 GND.t174 19.8005
R8320 GND.n3107 GND.t130 19.8005
R8321 GND.n3108 GND.t157 19.8005
R8322 GND.n3108 GND.t119 19.8005
R8323 GND.n1916 GND.n1915 19.5876
R8324 GND.n3962 GND.n3961 19.5087
R8325 GND.n4246 GND.n4245 19.3944
R8326 GND.n4245 GND.n3903 19.3944
R8327 GND.n4320 GND.n3903 19.3944
R8328 GND.n4314 GND.n4213 19.3944
R8329 GND.n4314 GND.n4214 19.3944
R8330 GND.n4270 GND.n4214 19.3944
R8331 GND.n4270 GND.n4269 19.3944
R8332 GND.n4269 GND.n4268 19.3944
R8333 GND.n4268 GND.n4219 19.3944
R8334 GND.n4264 GND.n4219 19.3944
R8335 GND.n4264 GND.n4263 19.3944
R8336 GND.n4263 GND.n4262 19.3944
R8337 GND.n4262 GND.n4225 19.3944
R8338 GND.n4258 GND.n4225 19.3944
R8339 GND.n4258 GND.n4257 19.3944
R8340 GND.n4257 GND.n4256 19.3944
R8341 GND.n4256 GND.n4231 19.3944
R8342 GND.n4252 GND.n4231 19.3944
R8343 GND.n4252 GND.n4251 19.3944
R8344 GND.n4251 GND.n4250 19.3944
R8345 GND.n4250 GND.n4237 19.3944
R8346 GND.n4337 GND.n3900 19.3944
R8347 GND.n4337 GND.n3901 19.3944
R8348 GND.n4333 GND.n3901 19.3944
R8349 GND.n4333 GND.n4332 19.3944
R8350 GND.n4332 GND.n4331 19.3944
R8351 GND.n4331 GND.n4328 19.3944
R8352 GND.n4328 GND.n3858 19.3944
R8353 GND.n4419 GND.n3858 19.3944
R8354 GND.n4419 GND.n3855 19.3944
R8355 GND.n4433 GND.n3855 19.3944
R8356 GND.n4433 GND.n3856 19.3944
R8357 GND.n4429 GND.n3856 19.3944
R8358 GND.n4429 GND.n4428 19.3944
R8359 GND.n4428 GND.n4427 19.3944
R8360 GND.n4427 GND.n3818 19.3944
R8361 GND.n4496 GND.n3818 19.3944
R8362 GND.n4496 GND.n3815 19.3944
R8363 GND.n4510 GND.n3815 19.3944
R8364 GND.n4510 GND.n3816 19.3944
R8365 GND.n4506 GND.n3816 19.3944
R8366 GND.n4506 GND.n4505 19.3944
R8367 GND.n4505 GND.n4504 19.3944
R8368 GND.n4504 GND.n3776 19.3944
R8369 GND.n4590 GND.n3776 19.3944
R8370 GND.n4590 GND.n3773 19.3944
R8371 GND.n4595 GND.n3773 19.3944
R8372 GND.n4595 GND.n3774 19.3944
R8373 GND.n3774 GND.n3746 19.3944
R8374 GND.n4629 GND.n3746 19.3944
R8375 GND.n4629 GND.n3743 19.3944
R8376 GND.n4668 GND.n3743 19.3944
R8377 GND.n4668 GND.n3744 19.3944
R8378 GND.n4664 GND.n3744 19.3944
R8379 GND.n4664 GND.n4663 19.3944
R8380 GND.n4663 GND.n4662 19.3944
R8381 GND.n4662 GND.n4636 19.3944
R8382 GND.n4658 GND.n4636 19.3944
R8383 GND.n4658 GND.n4657 19.3944
R8384 GND.n4657 GND.n4656 19.3944
R8385 GND.n4656 GND.n4640 19.3944
R8386 GND.n4652 GND.n4640 19.3944
R8387 GND.n4652 GND.n4651 19.3944
R8388 GND.n4651 GND.n4650 19.3944
R8389 GND.n4650 GND.n4647 19.3944
R8390 GND.n4647 GND.n3658 19.3944
R8391 GND.n4805 GND.n3658 19.3944
R8392 GND.n4805 GND.n3655 19.3944
R8393 GND.n4844 GND.n3655 19.3944
R8394 GND.n4844 GND.n3656 19.3944
R8395 GND.n4840 GND.n3656 19.3944
R8396 GND.n4840 GND.n4839 19.3944
R8397 GND.n4839 GND.n4838 19.3944
R8398 GND.n4838 GND.n4812 19.3944
R8399 GND.n4834 GND.n4812 19.3944
R8400 GND.n4834 GND.n4833 19.3944
R8401 GND.n4833 GND.n4832 19.3944
R8402 GND.n4832 GND.n4816 19.3944
R8403 GND.n4828 GND.n4816 19.3944
R8404 GND.n4828 GND.n4827 19.3944
R8405 GND.n4827 GND.n4826 19.3944
R8406 GND.n4826 GND.n4823 19.3944
R8407 GND.n4823 GND.n3570 19.3944
R8408 GND.n4981 GND.n3570 19.3944
R8409 GND.n4981 GND.n3567 19.3944
R8410 GND.n5020 GND.n3567 19.3944
R8411 GND.n5020 GND.n3568 19.3944
R8412 GND.n5016 GND.n3568 19.3944
R8413 GND.n5016 GND.n5015 19.3944
R8414 GND.n5015 GND.n5014 19.3944
R8415 GND.n5014 GND.n4988 19.3944
R8416 GND.n5010 GND.n4988 19.3944
R8417 GND.n5010 GND.n5009 19.3944
R8418 GND.n5009 GND.n5008 19.3944
R8419 GND.n5008 GND.n4992 19.3944
R8420 GND.n5004 GND.n4992 19.3944
R8421 GND.n5004 GND.n5003 19.3944
R8422 GND.n5003 GND.n5002 19.3944
R8423 GND.n5002 GND.n4999 19.3944
R8424 GND.n4999 GND.n3481 19.3944
R8425 GND.n5157 GND.n3481 19.3944
R8426 GND.n5157 GND.n3478 19.3944
R8427 GND.n5196 GND.n3478 19.3944
R8428 GND.n5196 GND.n3479 19.3944
R8429 GND.n5192 GND.n3479 19.3944
R8430 GND.n5192 GND.n5191 19.3944
R8431 GND.n5191 GND.n5190 19.3944
R8432 GND.n5190 GND.n5164 19.3944
R8433 GND.n5186 GND.n5164 19.3944
R8434 GND.n5186 GND.n5185 19.3944
R8435 GND.n5185 GND.n5184 19.3944
R8436 GND.n5184 GND.n5168 19.3944
R8437 GND.n5180 GND.n5168 19.3944
R8438 GND.n5180 GND.n5179 19.3944
R8439 GND.n5179 GND.n5178 19.3944
R8440 GND.n5178 GND.n5175 19.3944
R8441 GND.n5175 GND.n3392 19.3944
R8442 GND.n5332 GND.n3392 19.3944
R8443 GND.n5332 GND.n3389 19.3944
R8444 GND.n5373 GND.n3389 19.3944
R8445 GND.n5373 GND.n3390 19.3944
R8446 GND.n5369 GND.n3390 19.3944
R8447 GND.n5369 GND.n5368 19.3944
R8448 GND.n5368 GND.n5367 19.3944
R8449 GND.n5367 GND.n5341 19.3944
R8450 GND.n5363 GND.n5341 19.3944
R8451 GND.n5363 GND.n5362 19.3944
R8452 GND.n5362 GND.n5361 19.3944
R8453 GND.n5361 GND.n5345 19.3944
R8454 GND.n5357 GND.n5345 19.3944
R8455 GND.n5357 GND.n5356 19.3944
R8456 GND.n5356 GND.n5355 19.3944
R8457 GND.n5355 GND.n5352 19.3944
R8458 GND.n5352 GND.n3306 19.3944
R8459 GND.n5510 GND.n3306 19.3944
R8460 GND.n5510 GND.n3303 19.3944
R8461 GND.n5526 GND.n3303 19.3944
R8462 GND.n5526 GND.n3304 19.3944
R8463 GND.n5522 GND.n3304 19.3944
R8464 GND.n5522 GND.n5521 19.3944
R8465 GND.n5521 GND.n5520 19.3944
R8466 GND.n5520 GND.n5517 19.3944
R8467 GND.n5517 GND.n3256 19.3944
R8468 GND.n5604 GND.n3256 19.3944
R8469 GND.n5604 GND.n3253 19.3944
R8470 GND.n5609 GND.n3253 19.3944
R8471 GND.n5609 GND.n3254 19.3944
R8472 GND.n3254 GND.n2901 19.3944
R8473 GND.n6628 GND.n2901 19.3944
R8474 GND.n7108 GND.n1289 19.3944
R8475 GND.n7108 GND.n7107 19.3944
R8476 GND.n7107 GND.n7106 19.3944
R8477 GND.n7106 GND.n1299 19.3944
R8478 GND.n7102 GND.n1299 19.3944
R8479 GND.n7102 GND.n7101 19.3944
R8480 GND.n7101 GND.n7100 19.3944
R8481 GND.n7100 GND.n1307 19.3944
R8482 GND.n7096 GND.n1307 19.3944
R8483 GND.n7096 GND.n7095 19.3944
R8484 GND.n7095 GND.n7094 19.3944
R8485 GND.n7094 GND.n1315 19.3944
R8486 GND.n7090 GND.n1315 19.3944
R8487 GND.n7090 GND.n7089 19.3944
R8488 GND.n7089 GND.n7088 19.3944
R8489 GND.n7088 GND.n1323 19.3944
R8490 GND.n7084 GND.n1323 19.3944
R8491 GND.n7084 GND.n7083 19.3944
R8492 GND.n7083 GND.n7082 19.3944
R8493 GND.n7082 GND.n1331 19.3944
R8494 GND.n7078 GND.n1331 19.3944
R8495 GND.n7078 GND.n7077 19.3944
R8496 GND.n7077 GND.n7076 19.3944
R8497 GND.n7076 GND.n1339 19.3944
R8498 GND.n7072 GND.n1339 19.3944
R8499 GND.n7072 GND.n7071 19.3944
R8500 GND.n7071 GND.n7070 19.3944
R8501 GND.n7070 GND.n1347 19.3944
R8502 GND.n7066 GND.n1347 19.3944
R8503 GND.n7066 GND.n7065 19.3944
R8504 GND.n7065 GND.n7064 19.3944
R8505 GND.n7064 GND.n1355 19.3944
R8506 GND.n7060 GND.n1355 19.3944
R8507 GND.n7060 GND.n7059 19.3944
R8508 GND.n7059 GND.n7058 19.3944
R8509 GND.n7058 GND.n1363 19.3944
R8510 GND.n7054 GND.n1363 19.3944
R8511 GND.n7054 GND.n7053 19.3944
R8512 GND.n7053 GND.n7052 19.3944
R8513 GND.n7052 GND.n1371 19.3944
R8514 GND.n7048 GND.n1371 19.3944
R8515 GND.n7048 GND.n7047 19.3944
R8516 GND.n7047 GND.n7046 19.3944
R8517 GND.n7039 GND.n7038 19.3944
R8518 GND.n7038 GND.n7037 19.3944
R8519 GND.n7037 GND.n1391 19.3944
R8520 GND.n7033 GND.n1391 19.3944
R8521 GND.n7033 GND.n7032 19.3944
R8522 GND.n7032 GND.n7031 19.3944
R8523 GND.n7031 GND.n1396 19.3944
R8524 GND.n7027 GND.n1396 19.3944
R8525 GND.n7025 GND.n1403 19.3944
R8526 GND.n7021 GND.n1403 19.3944
R8527 GND.n7019 GND.n1409 19.3944
R8528 GND.n7015 GND.n1409 19.3944
R8529 GND.n7015 GND.n7014 19.3944
R8530 GND.n7014 GND.n7013 19.3944
R8531 GND.n7009 GND.n7008 19.3944
R8532 GND.n7008 GND.n7007 19.3944
R8533 GND.n7007 GND.n1421 19.3944
R8534 GND.n7003 GND.n1421 19.3944
R8535 GND.n7003 GND.n7002 19.3944
R8536 GND.n7002 GND.n7001 19.3944
R8537 GND.n7001 GND.n1426 19.3944
R8538 GND.n6997 GND.n1426 19.3944
R8539 GND.n6997 GND.n6996 19.3944
R8540 GND.n2210 GND.n2175 19.3944
R8541 GND.n2215 GND.n2175 19.3944
R8542 GND.n2215 GND.n2176 19.3944
R8543 GND.n2176 GND.n2139 19.3944
R8544 GND.n2281 GND.n2139 19.3944
R8545 GND.n2281 GND.n2136 19.3944
R8546 GND.n2286 GND.n2136 19.3944
R8547 GND.n2286 GND.n2137 19.3944
R8548 GND.n2137 GND.n2115 19.3944
R8549 GND.n2305 GND.n2115 19.3944
R8550 GND.n2305 GND.n2112 19.3944
R8551 GND.n2310 GND.n2112 19.3944
R8552 GND.n2310 GND.n2113 19.3944
R8553 GND.n2113 GND.n2092 19.3944
R8554 GND.n2328 GND.n2092 19.3944
R8555 GND.n2328 GND.n2090 19.3944
R8556 GND.n2332 GND.n2090 19.3944
R8557 GND.n2333 GND.n2332 19.3944
R8558 GND.n2336 GND.n2333 19.3944
R8559 GND.n2336 GND.n2088 19.3944
R8560 GND.n2340 GND.n2088 19.3944
R8561 GND.n2341 GND.n2340 19.3944
R8562 GND.n2341 GND.n2086 19.3944
R8563 GND.n2345 GND.n2086 19.3944
R8564 GND.n2345 GND.n2037 19.3944
R8565 GND.n2425 GND.n2037 19.3944
R8566 GND.n2425 GND.n2035 19.3944
R8567 GND.n2431 GND.n2035 19.3944
R8568 GND.n2431 GND.n2430 19.3944
R8569 GND.n2430 GND.n2015 19.3944
R8570 GND.n2451 GND.n2015 19.3944
R8571 GND.n2451 GND.n2013 19.3944
R8572 GND.n2461 GND.n2013 19.3944
R8573 GND.n2461 GND.n2460 19.3944
R8574 GND.n2460 GND.n2459 19.3944
R8575 GND.n2459 GND.n1982 19.3944
R8576 GND.n2495 GND.n1982 19.3944
R8577 GND.n2495 GND.n2494 19.3944
R8578 GND.n2494 GND.n2493 19.3944
R8579 GND.n2493 GND.n1993 19.3944
R8580 GND.n1993 GND.n1992 19.3944
R8581 GND.n1992 GND.n1990 19.3944
R8582 GND.n1990 GND.n1989 19.3944
R8583 GND.n1941 GND.n1940 19.3944
R8584 GND.n1945 GND.n1944 19.3944
R8585 GND.n1949 GND.n1948 19.3944
R8586 GND.n1953 GND.n1952 19.3944
R8587 GND.n2191 GND.n2190 19.3944
R8588 GND.n2194 GND.n2191 19.3944
R8589 GND.n2194 GND.n2185 19.3944
R8590 GND.n2198 GND.n2185 19.3944
R8591 GND.n2199 GND.n2198 19.3944
R8592 GND.n2202 GND.n2199 19.3944
R8593 GND.n2202 GND.n2181 19.3944
R8594 GND.n2206 GND.n2181 19.3944
R8595 GND.n7111 GND.n1295 19.3944
R8596 GND.n2153 GND.n1295 19.3944
R8597 GND.n2153 GND.n1300 19.3944
R8598 GND.n1301 GND.n1300 19.3944
R8599 GND.n1302 GND.n1301 19.3944
R8600 GND.n2132 GND.n1302 19.3944
R8601 GND.n2132 GND.n1308 19.3944
R8602 GND.n1309 GND.n1308 19.3944
R8603 GND.n1310 GND.n1309 19.3944
R8604 GND.n2119 GND.n1310 19.3944
R8605 GND.n2119 GND.n1316 19.3944
R8606 GND.n1317 GND.n1316 19.3944
R8607 GND.n1318 GND.n1317 19.3944
R8608 GND.n2314 GND.n1318 19.3944
R8609 GND.n2314 GND.n1324 19.3944
R8610 GND.n1325 GND.n1324 19.3944
R8611 GND.n1326 GND.n1325 19.3944
R8612 GND.n2062 GND.n1326 19.3944
R8613 GND.n2062 GND.n1332 19.3944
R8614 GND.n1333 GND.n1332 19.3944
R8615 GND.n1334 GND.n1333 19.3944
R8616 GND.n2395 GND.n1334 19.3944
R8617 GND.n2395 GND.n1340 19.3944
R8618 GND.n1341 GND.n1340 19.3944
R8619 GND.n1342 GND.n1341 19.3944
R8620 GND.n2041 GND.n1342 19.3944
R8621 GND.n2041 GND.n1348 19.3944
R8622 GND.n1349 GND.n1348 19.3944
R8623 GND.n1350 GND.n1349 19.3944
R8624 GND.n2435 GND.n1350 19.3944
R8625 GND.n2435 GND.n1356 19.3944
R8626 GND.n1357 GND.n1356 19.3944
R8627 GND.n1358 GND.n1357 19.3944
R8628 GND.n2466 GND.n1358 19.3944
R8629 GND.n2466 GND.n1364 19.3944
R8630 GND.n1365 GND.n1364 19.3944
R8631 GND.n1366 GND.n1365 19.3944
R8632 GND.n2499 GND.n1366 19.3944
R8633 GND.n2499 GND.n1372 19.3944
R8634 GND.n1373 GND.n1372 19.3944
R8635 GND.n1374 GND.n1373 19.3944
R8636 GND.n2515 GND.n1374 19.3944
R8637 GND.n2515 GND.n2514 19.3944
R8638 GND.n8214 GND.n530 19.3944
R8639 GND.n8220 GND.n530 19.3944
R8640 GND.n8220 GND.n528 19.3944
R8641 GND.n8224 GND.n528 19.3944
R8642 GND.n8224 GND.n524 19.3944
R8643 GND.n8230 GND.n524 19.3944
R8644 GND.n8230 GND.n522 19.3944
R8645 GND.n8234 GND.n522 19.3944
R8646 GND.n8234 GND.n518 19.3944
R8647 GND.n8240 GND.n518 19.3944
R8648 GND.n8240 GND.n516 19.3944
R8649 GND.n8244 GND.n516 19.3944
R8650 GND.n8244 GND.n512 19.3944
R8651 GND.n8250 GND.n512 19.3944
R8652 GND.n8250 GND.n510 19.3944
R8653 GND.n8254 GND.n510 19.3944
R8654 GND.n8254 GND.n506 19.3944
R8655 GND.n8260 GND.n506 19.3944
R8656 GND.n8260 GND.n504 19.3944
R8657 GND.n8264 GND.n504 19.3944
R8658 GND.n8264 GND.n500 19.3944
R8659 GND.n8270 GND.n500 19.3944
R8660 GND.n8270 GND.n498 19.3944
R8661 GND.n8274 GND.n498 19.3944
R8662 GND.n8274 GND.n494 19.3944
R8663 GND.n8280 GND.n494 19.3944
R8664 GND.n8280 GND.n492 19.3944
R8665 GND.n8284 GND.n492 19.3944
R8666 GND.n8284 GND.n488 19.3944
R8667 GND.n8290 GND.n488 19.3944
R8668 GND.n8290 GND.n486 19.3944
R8669 GND.n8294 GND.n486 19.3944
R8670 GND.n8294 GND.n482 19.3944
R8671 GND.n8300 GND.n482 19.3944
R8672 GND.n8300 GND.n480 19.3944
R8673 GND.n8304 GND.n480 19.3944
R8674 GND.n8304 GND.n476 19.3944
R8675 GND.n8310 GND.n476 19.3944
R8676 GND.n8310 GND.n474 19.3944
R8677 GND.n8314 GND.n474 19.3944
R8678 GND.n8314 GND.n470 19.3944
R8679 GND.n8320 GND.n470 19.3944
R8680 GND.n8320 GND.n468 19.3944
R8681 GND.n8324 GND.n468 19.3944
R8682 GND.n8324 GND.n464 19.3944
R8683 GND.n8330 GND.n464 19.3944
R8684 GND.n8330 GND.n462 19.3944
R8685 GND.n8334 GND.n462 19.3944
R8686 GND.n8334 GND.n458 19.3944
R8687 GND.n8340 GND.n458 19.3944
R8688 GND.n8340 GND.n456 19.3944
R8689 GND.n8344 GND.n456 19.3944
R8690 GND.n8344 GND.n452 19.3944
R8691 GND.n8350 GND.n452 19.3944
R8692 GND.n8350 GND.n450 19.3944
R8693 GND.n8354 GND.n450 19.3944
R8694 GND.n8354 GND.n446 19.3944
R8695 GND.n8360 GND.n446 19.3944
R8696 GND.n8360 GND.n444 19.3944
R8697 GND.n8364 GND.n444 19.3944
R8698 GND.n8364 GND.n440 19.3944
R8699 GND.n8370 GND.n440 19.3944
R8700 GND.n8370 GND.n438 19.3944
R8701 GND.n8374 GND.n438 19.3944
R8702 GND.n8374 GND.n434 19.3944
R8703 GND.n8380 GND.n434 19.3944
R8704 GND.n8380 GND.n432 19.3944
R8705 GND.n8384 GND.n432 19.3944
R8706 GND.n8384 GND.n428 19.3944
R8707 GND.n8390 GND.n428 19.3944
R8708 GND.n8390 GND.n426 19.3944
R8709 GND.n8395 GND.n426 19.3944
R8710 GND.n7373 GND.n1033 19.3944
R8711 GND.n7379 GND.n1033 19.3944
R8712 GND.n7379 GND.n1031 19.3944
R8713 GND.n7383 GND.n1031 19.3944
R8714 GND.n7383 GND.n1027 19.3944
R8715 GND.n7389 GND.n1027 19.3944
R8716 GND.n7389 GND.n1025 19.3944
R8717 GND.n7393 GND.n1025 19.3944
R8718 GND.n7393 GND.n1021 19.3944
R8719 GND.n7399 GND.n1021 19.3944
R8720 GND.n7399 GND.n1019 19.3944
R8721 GND.n7403 GND.n1019 19.3944
R8722 GND.n7403 GND.n1015 19.3944
R8723 GND.n7409 GND.n1015 19.3944
R8724 GND.n7409 GND.n1013 19.3944
R8725 GND.n7413 GND.n1013 19.3944
R8726 GND.n7413 GND.n1009 19.3944
R8727 GND.n7419 GND.n1009 19.3944
R8728 GND.n7419 GND.n1007 19.3944
R8729 GND.n7423 GND.n1007 19.3944
R8730 GND.n7423 GND.n1003 19.3944
R8731 GND.n7429 GND.n1003 19.3944
R8732 GND.n7429 GND.n1001 19.3944
R8733 GND.n7433 GND.n1001 19.3944
R8734 GND.n7433 GND.n997 19.3944
R8735 GND.n7439 GND.n997 19.3944
R8736 GND.n7439 GND.n995 19.3944
R8737 GND.n7443 GND.n995 19.3944
R8738 GND.n7443 GND.n991 19.3944
R8739 GND.n7449 GND.n991 19.3944
R8740 GND.n7449 GND.n989 19.3944
R8741 GND.n7453 GND.n989 19.3944
R8742 GND.n7453 GND.n985 19.3944
R8743 GND.n7459 GND.n985 19.3944
R8744 GND.n7459 GND.n983 19.3944
R8745 GND.n7463 GND.n983 19.3944
R8746 GND.n7463 GND.n979 19.3944
R8747 GND.n7469 GND.n979 19.3944
R8748 GND.n7469 GND.n977 19.3944
R8749 GND.n7473 GND.n977 19.3944
R8750 GND.n7473 GND.n973 19.3944
R8751 GND.n7479 GND.n973 19.3944
R8752 GND.n7479 GND.n971 19.3944
R8753 GND.n7483 GND.n971 19.3944
R8754 GND.n7483 GND.n967 19.3944
R8755 GND.n7489 GND.n967 19.3944
R8756 GND.n7489 GND.n965 19.3944
R8757 GND.n7493 GND.n965 19.3944
R8758 GND.n7493 GND.n961 19.3944
R8759 GND.n7499 GND.n961 19.3944
R8760 GND.n7499 GND.n959 19.3944
R8761 GND.n7503 GND.n959 19.3944
R8762 GND.n7503 GND.n955 19.3944
R8763 GND.n7509 GND.n955 19.3944
R8764 GND.n7509 GND.n953 19.3944
R8765 GND.n7513 GND.n953 19.3944
R8766 GND.n7513 GND.n949 19.3944
R8767 GND.n7519 GND.n949 19.3944
R8768 GND.n7519 GND.n947 19.3944
R8769 GND.n7523 GND.n947 19.3944
R8770 GND.n7523 GND.n943 19.3944
R8771 GND.n7529 GND.n943 19.3944
R8772 GND.n7529 GND.n941 19.3944
R8773 GND.n7533 GND.n941 19.3944
R8774 GND.n7533 GND.n937 19.3944
R8775 GND.n7539 GND.n937 19.3944
R8776 GND.n7539 GND.n935 19.3944
R8777 GND.n7543 GND.n935 19.3944
R8778 GND.n7543 GND.n931 19.3944
R8779 GND.n7549 GND.n931 19.3944
R8780 GND.n7549 GND.n929 19.3944
R8781 GND.n7553 GND.n929 19.3944
R8782 GND.n7553 GND.n925 19.3944
R8783 GND.n7559 GND.n925 19.3944
R8784 GND.n7559 GND.n923 19.3944
R8785 GND.n7563 GND.n923 19.3944
R8786 GND.n7563 GND.n919 19.3944
R8787 GND.n7569 GND.n919 19.3944
R8788 GND.n7569 GND.n917 19.3944
R8789 GND.n7573 GND.n917 19.3944
R8790 GND.n7573 GND.n913 19.3944
R8791 GND.n7579 GND.n913 19.3944
R8792 GND.n7579 GND.n911 19.3944
R8793 GND.n7583 GND.n911 19.3944
R8794 GND.n7583 GND.n907 19.3944
R8795 GND.n7589 GND.n907 19.3944
R8796 GND.n7589 GND.n905 19.3944
R8797 GND.n7593 GND.n905 19.3944
R8798 GND.n7593 GND.n901 19.3944
R8799 GND.n7599 GND.n901 19.3944
R8800 GND.n7599 GND.n899 19.3944
R8801 GND.n7603 GND.n899 19.3944
R8802 GND.n7603 GND.n895 19.3944
R8803 GND.n7609 GND.n895 19.3944
R8804 GND.n7609 GND.n893 19.3944
R8805 GND.n7613 GND.n893 19.3944
R8806 GND.n7613 GND.n889 19.3944
R8807 GND.n7619 GND.n889 19.3944
R8808 GND.n7619 GND.n887 19.3944
R8809 GND.n7623 GND.n887 19.3944
R8810 GND.n7623 GND.n883 19.3944
R8811 GND.n7629 GND.n883 19.3944
R8812 GND.n7629 GND.n881 19.3944
R8813 GND.n7633 GND.n881 19.3944
R8814 GND.n7633 GND.n877 19.3944
R8815 GND.n7639 GND.n877 19.3944
R8816 GND.n7639 GND.n875 19.3944
R8817 GND.n7643 GND.n875 19.3944
R8818 GND.n7643 GND.n871 19.3944
R8819 GND.n7649 GND.n871 19.3944
R8820 GND.n7649 GND.n869 19.3944
R8821 GND.n7653 GND.n869 19.3944
R8822 GND.n7653 GND.n865 19.3944
R8823 GND.n7659 GND.n865 19.3944
R8824 GND.n7659 GND.n863 19.3944
R8825 GND.n7663 GND.n863 19.3944
R8826 GND.n7663 GND.n859 19.3944
R8827 GND.n7669 GND.n859 19.3944
R8828 GND.n7669 GND.n857 19.3944
R8829 GND.n7673 GND.n857 19.3944
R8830 GND.n7673 GND.n853 19.3944
R8831 GND.n7679 GND.n853 19.3944
R8832 GND.n7679 GND.n851 19.3944
R8833 GND.n7683 GND.n851 19.3944
R8834 GND.n7683 GND.n847 19.3944
R8835 GND.n7689 GND.n847 19.3944
R8836 GND.n7689 GND.n845 19.3944
R8837 GND.n7693 GND.n845 19.3944
R8838 GND.n7693 GND.n841 19.3944
R8839 GND.n7699 GND.n841 19.3944
R8840 GND.n7699 GND.n839 19.3944
R8841 GND.n7703 GND.n839 19.3944
R8842 GND.n7703 GND.n835 19.3944
R8843 GND.n7709 GND.n835 19.3944
R8844 GND.n7709 GND.n833 19.3944
R8845 GND.n7713 GND.n833 19.3944
R8846 GND.n7713 GND.n829 19.3944
R8847 GND.n7719 GND.n829 19.3944
R8848 GND.n7719 GND.n827 19.3944
R8849 GND.n7723 GND.n827 19.3944
R8850 GND.n7723 GND.n823 19.3944
R8851 GND.n7729 GND.n823 19.3944
R8852 GND.n7729 GND.n821 19.3944
R8853 GND.n7733 GND.n821 19.3944
R8854 GND.n7733 GND.n817 19.3944
R8855 GND.n7739 GND.n817 19.3944
R8856 GND.n7739 GND.n815 19.3944
R8857 GND.n7743 GND.n815 19.3944
R8858 GND.n7743 GND.n811 19.3944
R8859 GND.n7749 GND.n811 19.3944
R8860 GND.n7749 GND.n809 19.3944
R8861 GND.n7753 GND.n809 19.3944
R8862 GND.n7753 GND.n805 19.3944
R8863 GND.n7759 GND.n805 19.3944
R8864 GND.n7759 GND.n803 19.3944
R8865 GND.n7763 GND.n803 19.3944
R8866 GND.n7763 GND.n799 19.3944
R8867 GND.n7769 GND.n799 19.3944
R8868 GND.n7769 GND.n797 19.3944
R8869 GND.n7773 GND.n797 19.3944
R8870 GND.n7773 GND.n793 19.3944
R8871 GND.n7779 GND.n793 19.3944
R8872 GND.n7779 GND.n791 19.3944
R8873 GND.n7783 GND.n791 19.3944
R8874 GND.n7783 GND.n787 19.3944
R8875 GND.n7789 GND.n787 19.3944
R8876 GND.n7789 GND.n785 19.3944
R8877 GND.n7793 GND.n785 19.3944
R8878 GND.n7793 GND.n781 19.3944
R8879 GND.n7799 GND.n781 19.3944
R8880 GND.n7799 GND.n779 19.3944
R8881 GND.n7803 GND.n779 19.3944
R8882 GND.n7803 GND.n775 19.3944
R8883 GND.n7809 GND.n775 19.3944
R8884 GND.n7809 GND.n773 19.3944
R8885 GND.n7813 GND.n773 19.3944
R8886 GND.n7813 GND.n769 19.3944
R8887 GND.n7819 GND.n769 19.3944
R8888 GND.n7819 GND.n767 19.3944
R8889 GND.n7823 GND.n767 19.3944
R8890 GND.n7823 GND.n763 19.3944
R8891 GND.n7829 GND.n763 19.3944
R8892 GND.n7829 GND.n761 19.3944
R8893 GND.n7833 GND.n761 19.3944
R8894 GND.n7833 GND.n757 19.3944
R8895 GND.n7839 GND.n757 19.3944
R8896 GND.n7839 GND.n755 19.3944
R8897 GND.n7843 GND.n755 19.3944
R8898 GND.n7843 GND.n751 19.3944
R8899 GND.n7849 GND.n751 19.3944
R8900 GND.n7849 GND.n749 19.3944
R8901 GND.n7853 GND.n749 19.3944
R8902 GND.n7853 GND.n745 19.3944
R8903 GND.n7859 GND.n745 19.3944
R8904 GND.n7859 GND.n743 19.3944
R8905 GND.n7863 GND.n743 19.3944
R8906 GND.n7863 GND.n739 19.3944
R8907 GND.n7869 GND.n739 19.3944
R8908 GND.n7869 GND.n737 19.3944
R8909 GND.n7873 GND.n737 19.3944
R8910 GND.n7873 GND.n733 19.3944
R8911 GND.n7879 GND.n733 19.3944
R8912 GND.n7879 GND.n731 19.3944
R8913 GND.n7883 GND.n731 19.3944
R8914 GND.n7883 GND.n727 19.3944
R8915 GND.n7889 GND.n727 19.3944
R8916 GND.n7889 GND.n725 19.3944
R8917 GND.n7893 GND.n725 19.3944
R8918 GND.n7893 GND.n721 19.3944
R8919 GND.n7899 GND.n721 19.3944
R8920 GND.n7899 GND.n719 19.3944
R8921 GND.n7903 GND.n719 19.3944
R8922 GND.n7903 GND.n715 19.3944
R8923 GND.n7909 GND.n715 19.3944
R8924 GND.n7909 GND.n713 19.3944
R8925 GND.n7913 GND.n713 19.3944
R8926 GND.n7913 GND.n709 19.3944
R8927 GND.n7919 GND.n709 19.3944
R8928 GND.n7919 GND.n707 19.3944
R8929 GND.n7923 GND.n707 19.3944
R8930 GND.n7923 GND.n703 19.3944
R8931 GND.n7929 GND.n703 19.3944
R8932 GND.n7929 GND.n701 19.3944
R8933 GND.n7933 GND.n701 19.3944
R8934 GND.n7933 GND.n697 19.3944
R8935 GND.n7939 GND.n697 19.3944
R8936 GND.n7939 GND.n695 19.3944
R8937 GND.n7943 GND.n695 19.3944
R8938 GND.n7943 GND.n691 19.3944
R8939 GND.n7949 GND.n691 19.3944
R8940 GND.n7949 GND.n689 19.3944
R8941 GND.n7953 GND.n689 19.3944
R8942 GND.n7953 GND.n685 19.3944
R8943 GND.n7959 GND.n685 19.3944
R8944 GND.n7959 GND.n683 19.3944
R8945 GND.n7963 GND.n683 19.3944
R8946 GND.n7963 GND.n679 19.3944
R8947 GND.n7969 GND.n679 19.3944
R8948 GND.n7969 GND.n677 19.3944
R8949 GND.n7973 GND.n677 19.3944
R8950 GND.n7973 GND.n673 19.3944
R8951 GND.n7979 GND.n673 19.3944
R8952 GND.n7979 GND.n671 19.3944
R8953 GND.n7983 GND.n671 19.3944
R8954 GND.n7983 GND.n667 19.3944
R8955 GND.n7989 GND.n667 19.3944
R8956 GND.n7989 GND.n665 19.3944
R8957 GND.n7993 GND.n665 19.3944
R8958 GND.n7993 GND.n661 19.3944
R8959 GND.n7999 GND.n661 19.3944
R8960 GND.n7999 GND.n659 19.3944
R8961 GND.n8003 GND.n659 19.3944
R8962 GND.n8003 GND.n655 19.3944
R8963 GND.n8009 GND.n655 19.3944
R8964 GND.n8009 GND.n653 19.3944
R8965 GND.n8013 GND.n653 19.3944
R8966 GND.n8013 GND.n649 19.3944
R8967 GND.n8019 GND.n649 19.3944
R8968 GND.n8019 GND.n647 19.3944
R8969 GND.n8023 GND.n647 19.3944
R8970 GND.n8023 GND.n643 19.3944
R8971 GND.n8029 GND.n643 19.3944
R8972 GND.n8029 GND.n641 19.3944
R8973 GND.n8033 GND.n641 19.3944
R8974 GND.n8033 GND.n637 19.3944
R8975 GND.n8039 GND.n637 19.3944
R8976 GND.n8039 GND.n635 19.3944
R8977 GND.n8043 GND.n635 19.3944
R8978 GND.n8043 GND.n631 19.3944
R8979 GND.n8049 GND.n631 19.3944
R8980 GND.n8049 GND.n629 19.3944
R8981 GND.n8053 GND.n629 19.3944
R8982 GND.n8053 GND.n625 19.3944
R8983 GND.n8059 GND.n625 19.3944
R8984 GND.n8059 GND.n623 19.3944
R8985 GND.n8063 GND.n623 19.3944
R8986 GND.n8063 GND.n619 19.3944
R8987 GND.n8069 GND.n619 19.3944
R8988 GND.n8069 GND.n617 19.3944
R8989 GND.n8073 GND.n617 19.3944
R8990 GND.n8073 GND.n613 19.3944
R8991 GND.n8079 GND.n613 19.3944
R8992 GND.n8079 GND.n611 19.3944
R8993 GND.n8083 GND.n611 19.3944
R8994 GND.n8083 GND.n607 19.3944
R8995 GND.n8089 GND.n607 19.3944
R8996 GND.n8089 GND.n605 19.3944
R8997 GND.n8093 GND.n605 19.3944
R8998 GND.n8093 GND.n601 19.3944
R8999 GND.n8099 GND.n601 19.3944
R9000 GND.n8099 GND.n599 19.3944
R9001 GND.n8103 GND.n599 19.3944
R9002 GND.n8103 GND.n595 19.3944
R9003 GND.n8109 GND.n595 19.3944
R9004 GND.n8109 GND.n593 19.3944
R9005 GND.n8113 GND.n593 19.3944
R9006 GND.n8113 GND.n589 19.3944
R9007 GND.n8119 GND.n589 19.3944
R9008 GND.n8119 GND.n587 19.3944
R9009 GND.n8123 GND.n587 19.3944
R9010 GND.n8123 GND.n583 19.3944
R9011 GND.n8129 GND.n583 19.3944
R9012 GND.n8129 GND.n581 19.3944
R9013 GND.n8133 GND.n581 19.3944
R9014 GND.n8133 GND.n577 19.3944
R9015 GND.n8139 GND.n577 19.3944
R9016 GND.n8139 GND.n575 19.3944
R9017 GND.n8143 GND.n575 19.3944
R9018 GND.n8143 GND.n571 19.3944
R9019 GND.n8149 GND.n571 19.3944
R9020 GND.n8149 GND.n569 19.3944
R9021 GND.n8153 GND.n569 19.3944
R9022 GND.n8153 GND.n565 19.3944
R9023 GND.n8159 GND.n565 19.3944
R9024 GND.n8159 GND.n563 19.3944
R9025 GND.n8163 GND.n563 19.3944
R9026 GND.n8163 GND.n559 19.3944
R9027 GND.n8169 GND.n559 19.3944
R9028 GND.n8169 GND.n557 19.3944
R9029 GND.n8173 GND.n557 19.3944
R9030 GND.n8173 GND.n553 19.3944
R9031 GND.n8179 GND.n553 19.3944
R9032 GND.n8179 GND.n551 19.3944
R9033 GND.n8183 GND.n551 19.3944
R9034 GND.n8183 GND.n547 19.3944
R9035 GND.n8189 GND.n547 19.3944
R9036 GND.n8189 GND.n545 19.3944
R9037 GND.n8193 GND.n545 19.3944
R9038 GND.n8193 GND.n541 19.3944
R9039 GND.n8199 GND.n541 19.3944
R9040 GND.n8199 GND.n539 19.3944
R9041 GND.n8204 GND.n539 19.3944
R9042 GND.n8204 GND.n535 19.3944
R9043 GND.n8210 GND.n535 19.3944
R9044 GND.n8211 GND.n8210 19.3944
R9045 GND.n6509 GND.n6508 19.3944
R9046 GND.n6508 GND.n6507 19.3944
R9047 GND.n6507 GND.n6506 19.3944
R9048 GND.n6506 GND.n6504 19.3944
R9049 GND.n6504 GND.n6501 19.3944
R9050 GND.n6501 GND.n6500 19.3944
R9051 GND.n6500 GND.n6497 19.3944
R9052 GND.n6497 GND.n6496 19.3944
R9053 GND.n6492 GND.n6489 19.3944
R9054 GND.n6489 GND.n6488 19.3944
R9055 GND.n6484 GND.n6482 19.3944
R9056 GND.n6482 GND.n6479 19.3944
R9057 GND.n6479 GND.n6478 19.3944
R9058 GND.n6478 GND.n6475 19.3944
R9059 GND.n6473 GND.n6471 19.3944
R9060 GND.n6471 GND.n6468 19.3944
R9061 GND.n6468 GND.n6467 19.3944
R9062 GND.n6467 GND.n6464 19.3944
R9063 GND.n6464 GND.n6463 19.3944
R9064 GND.n6463 GND.n6460 19.3944
R9065 GND.n6460 GND.n6459 19.3944
R9066 GND.n6459 GND.n6456 19.3944
R9067 GND.n6456 GND.n6455 19.3944
R9068 GND.n6443 GND.n5818 19.3944
R9069 GND.n6443 GND.n6442 19.3944
R9070 GND.n6442 GND.n5827 19.3944
R9071 GND.n6047 GND.n5827 19.3944
R9072 GND.n6148 GND.n6047 19.3944
R9073 GND.n6149 GND.n6148 19.3944
R9074 GND.n6151 GND.n6149 19.3944
R9075 GND.n6151 GND.n6043 19.3944
R9076 GND.n6163 GND.n6043 19.3944
R9077 GND.n6164 GND.n6163 19.3944
R9078 GND.n6166 GND.n6164 19.3944
R9079 GND.n6166 GND.n6039 19.3944
R9080 GND.n6178 GND.n6039 19.3944
R9081 GND.n6179 GND.n6178 19.3944
R9082 GND.n6181 GND.n6179 19.3944
R9083 GND.n6181 GND.n5976 19.3944
R9084 GND.n6200 GND.n5976 19.3944
R9085 GND.n6201 GND.n6200 19.3944
R9086 GND.n6202 GND.n6201 19.3944
R9087 GND.n6206 GND.n6202 19.3944
R9088 GND.n6207 GND.n6206 19.3944
R9089 GND.n6208 GND.n6207 19.3944
R9090 GND.n6209 GND.n6208 19.3944
R9091 GND.n6210 GND.n6209 19.3944
R9092 GND.n6213 GND.n6210 19.3944
R9093 GND.n6213 GND.n5969 19.3944
R9094 GND.n6225 GND.n5969 19.3944
R9095 GND.n6226 GND.n6225 19.3944
R9096 GND.n6228 GND.n6226 19.3944
R9097 GND.n6228 GND.n5965 19.3944
R9098 GND.n6241 GND.n5965 19.3944
R9099 GND.n6242 GND.n6241 19.3944
R9100 GND.n6244 GND.n6242 19.3944
R9101 GND.n6245 GND.n6244 19.3944
R9102 GND.n6345 GND.n6245 19.3944
R9103 GND.n6345 GND.n6344 19.3944
R9104 GND.n6344 GND.n6343 19.3944
R9105 GND.n6343 GND.n6247 19.3944
R9106 GND.n6306 GND.n6247 19.3944
R9107 GND.n6306 GND.n6305 19.3944
R9108 GND.n6305 GND.n6304 19.3944
R9109 GND.n6304 GND.n250 19.3944
R9110 GND.n8448 GND.n250 19.3944
R9111 GND.n6446 GND.n6445 19.3944
R9112 GND.n6445 GND.n5825 19.3944
R9113 GND.n5850 GND.n5825 19.3944
R9114 GND.n6432 GND.n5850 19.3944
R9115 GND.n6432 GND.n6431 19.3944
R9116 GND.n6431 GND.n6430 19.3944
R9117 GND.n6430 GND.n5855 19.3944
R9118 GND.n6420 GND.n5855 19.3944
R9119 GND.n6420 GND.n6419 19.3944
R9120 GND.n6419 GND.n6418 19.3944
R9121 GND.n6418 GND.n5876 19.3944
R9122 GND.n6408 GND.n5876 19.3944
R9123 GND.n6408 GND.n6407 19.3944
R9124 GND.n6407 GND.n6406 19.3944
R9125 GND.n6406 GND.n5897 19.3944
R9126 GND.n6396 GND.n5897 19.3944
R9127 GND.n6396 GND.n6395 19.3944
R9128 GND.n6395 GND.n6394 19.3944
R9129 GND.n6394 GND.n5916 19.3944
R9130 GND.n5935 GND.n5916 19.3944
R9131 GND.n6377 GND.n5935 19.3944
R9132 GND.n6377 GND.n6376 19.3944
R9133 GND.n6376 GND.n6375 19.3944
R9134 GND.n6375 GND.n5939 19.3944
R9135 GND.n5939 GND.n166 19.3944
R9136 GND.n8499 GND.n166 19.3944
R9137 GND.n8499 GND.n8498 19.3944
R9138 GND.n8498 GND.n8497 19.3944
R9139 GND.n8497 GND.n170 19.3944
R9140 GND.n8487 GND.n170 19.3944
R9141 GND.n8487 GND.n8486 19.3944
R9142 GND.n8486 GND.n8485 19.3944
R9143 GND.n8485 GND.n190 19.3944
R9144 GND.n8475 GND.n190 19.3944
R9145 GND.n8475 GND.n8474 19.3944
R9146 GND.n8474 GND.n8473 19.3944
R9147 GND.n8473 GND.n210 19.3944
R9148 GND.n8463 GND.n210 19.3944
R9149 GND.n8463 GND.n8462 19.3944
R9150 GND.n8462 GND.n8461 19.3944
R9151 GND.n8461 GND.n231 19.3944
R9152 GND.n8451 GND.n231 19.3944
R9153 GND.n8451 GND.n8450 19.3944
R9154 GND.n335 GND.n298 19.3944
R9155 GND.n335 GND.n332 19.3944
R9156 GND.n332 GND.n331 19.3944
R9157 GND.n331 GND.n328 19.3944
R9158 GND.n328 GND.n327 19.3944
R9159 GND.n327 GND.n324 19.3944
R9160 GND.n324 GND.n323 19.3944
R9161 GND.n323 GND.n320 19.3944
R9162 GND.n320 GND.n319 19.3944
R9163 GND.n358 GND.n287 19.3944
R9164 GND.n358 GND.n355 19.3944
R9165 GND.n355 GND.n352 19.3944
R9166 GND.n352 GND.n351 19.3944
R9167 GND.n351 GND.n348 19.3944
R9168 GND.n348 GND.n347 19.3944
R9169 GND.n347 GND.n344 19.3944
R9170 GND.n344 GND.n343 19.3944
R9171 GND.n343 GND.n340 19.3944
R9172 GND.n381 GND.n380 19.3944
R9173 GND.n380 GND.n281 19.3944
R9174 GND.n376 GND.n281 19.3944
R9175 GND.n376 GND.n373 19.3944
R9176 GND.n373 GND.n370 19.3944
R9177 GND.n370 GND.n369 19.3944
R9178 GND.n369 GND.n366 19.3944
R9179 GND.n366 GND.n365 19.3944
R9180 GND.n6270 GND.n6268 19.3944
R9181 GND.n6276 GND.n6268 19.3944
R9182 GND.n6276 GND.n6266 19.3944
R9183 GND.n6280 GND.n6266 19.3944
R9184 GND.n6280 GND.n6264 19.3944
R9185 GND.n6286 GND.n6264 19.3944
R9186 GND.n6286 GND.n6262 19.3944
R9187 GND.n6290 GND.n6262 19.3944
R9188 GND.n6136 GND.n6050 19.3944
R9189 GND.n6137 GND.n6136 19.3944
R9190 GND.n6140 GND.n6137 19.3944
R9191 GND.n6140 GND.n6048 19.3944
R9192 GND.n6144 GND.n6048 19.3944
R9193 GND.n6144 GND.n6046 19.3944
R9194 GND.n6155 GND.n6046 19.3944
R9195 GND.n6155 GND.n6044 19.3944
R9196 GND.n6159 GND.n6044 19.3944
R9197 GND.n6159 GND.n6042 19.3944
R9198 GND.n6170 GND.n6042 19.3944
R9199 GND.n6170 GND.n6040 19.3944
R9200 GND.n6174 GND.n6040 19.3944
R9201 GND.n6174 GND.n6038 19.3944
R9202 GND.n6185 GND.n6038 19.3944
R9203 GND.n6185 GND.n6036 19.3944
R9204 GND.n6196 GND.n6036 19.3944
R9205 GND.n6196 GND.n6195 19.3944
R9206 GND.n6195 GND.n6194 19.3944
R9207 GND.n6194 GND.n6193 19.3944
R9208 GND.n6193 GND.n138 19.3944
R9209 GND.n8510 GND.n138 19.3944
R9210 GND.n8510 GND.n139 19.3944
R9211 GND.n5972 GND.n139 19.3944
R9212 GND.n6217 GND.n5972 19.3944
R9213 GND.n6217 GND.n5970 19.3944
R9214 GND.n6221 GND.n5970 19.3944
R9215 GND.n6221 GND.n5968 19.3944
R9216 GND.n6232 GND.n5968 19.3944
R9217 GND.n6232 GND.n5966 19.3944
R9218 GND.n6237 GND.n5966 19.3944
R9219 GND.n6237 GND.n5960 19.3944
R9220 GND.n6351 GND.n5960 19.3944
R9221 GND.n6351 GND.n6350 19.3944
R9222 GND.n6350 GND.n6349 19.3944
R9223 GND.n6349 GND.n5964 19.3944
R9224 GND.n6339 GND.n5964 19.3944
R9225 GND.n6339 GND.n6338 19.3944
R9226 GND.n6338 GND.n6337 19.3944
R9227 GND.n6337 GND.n6252 19.3944
R9228 GND.n6300 GND.n6252 19.3944
R9229 GND.n6300 GND.n6299 19.3944
R9230 GND.n6299 GND.n6298 19.3944
R9231 GND.n6132 GND.n6131 19.3944
R9232 GND.n6128 GND.n6127 19.3944
R9233 GND.n6124 GND.n6123 19.3944
R9234 GND.n6120 GND.n6119 19.3944
R9235 GND.n5836 GND.n5835 19.3944
R9236 GND.n6438 GND.n5835 19.3944
R9237 GND.n6438 GND.n6437 19.3944
R9238 GND.n6437 GND.n6436 19.3944
R9239 GND.n6436 GND.n5842 19.3944
R9240 GND.n6426 GND.n5842 19.3944
R9241 GND.n6426 GND.n6425 19.3944
R9242 GND.n6425 GND.n6424 19.3944
R9243 GND.n6424 GND.n5866 19.3944
R9244 GND.n6414 GND.n5866 19.3944
R9245 GND.n6414 GND.n6413 19.3944
R9246 GND.n6413 GND.n6412 19.3944
R9247 GND.n6412 GND.n5887 19.3944
R9248 GND.n6402 GND.n5887 19.3944
R9249 GND.n6402 GND.n6401 19.3944
R9250 GND.n6401 GND.n6400 19.3944
R9251 GND.n6400 GND.n5907 19.3944
R9252 GND.n6390 GND.n154 19.3944
R9253 GND.n5922 GND.n154 19.3944
R9254 GND.n8506 GND.n147 19.3944
R9255 GND.n5942 GND.n148 19.3944
R9256 GND.n8503 GND.n156 19.3944
R9257 GND.n8503 GND.n157 19.3944
R9258 GND.n8493 GND.n157 19.3944
R9259 GND.n8493 GND.n8492 19.3944
R9260 GND.n8492 GND.n8491 19.3944
R9261 GND.n8491 GND.n180 19.3944
R9262 GND.n8481 GND.n180 19.3944
R9263 GND.n8481 GND.n8480 19.3944
R9264 GND.n8480 GND.n8479 19.3944
R9265 GND.n8479 GND.n200 19.3944
R9266 GND.n8469 GND.n200 19.3944
R9267 GND.n8469 GND.n8468 19.3944
R9268 GND.n8468 GND.n8467 19.3944
R9269 GND.n8467 GND.n221 19.3944
R9270 GND.n8457 GND.n221 19.3944
R9271 GND.n8457 GND.n8456 19.3944
R9272 GND.n8456 GND.n8455 19.3944
R9273 GND.n8455 GND.n241 19.3944
R9274 GND.n7223 GND.n1181 19.3944
R9275 GND.n7217 GND.n1181 19.3944
R9276 GND.n7217 GND.n7216 19.3944
R9277 GND.n7216 GND.n7215 19.3944
R9278 GND.n7215 GND.n1188 19.3944
R9279 GND.n7209 GND.n1188 19.3944
R9280 GND.n7209 GND.n7208 19.3944
R9281 GND.n7208 GND.n7207 19.3944
R9282 GND.n7207 GND.n1196 19.3944
R9283 GND.n7201 GND.n1196 19.3944
R9284 GND.n7201 GND.n7200 19.3944
R9285 GND.n7200 GND.n7199 19.3944
R9286 GND.n7199 GND.n1204 19.3944
R9287 GND.n7193 GND.n1204 19.3944
R9288 GND.n7193 GND.n7192 19.3944
R9289 GND.n7192 GND.n7191 19.3944
R9290 GND.n7191 GND.n1212 19.3944
R9291 GND.n7185 GND.n1212 19.3944
R9292 GND.n7185 GND.n7184 19.3944
R9293 GND.n7184 GND.n7183 19.3944
R9294 GND.n7183 GND.n1220 19.3944
R9295 GND.n2161 GND.n1220 19.3944
R9296 GND.n2165 GND.n2161 19.3944
R9297 GND.n2165 GND.n2159 19.3944
R9298 GND.n2220 GND.n2159 19.3944
R9299 GND.n2220 GND.n2157 19.3944
R9300 GND.n2262 GND.n2157 19.3944
R9301 GND.n2262 GND.n2261 19.3944
R9302 GND.n2261 GND.n2260 19.3944
R9303 GND.n2260 GND.n2226 19.3944
R9304 GND.n2256 GND.n2226 19.3944
R9305 GND.n2256 GND.n2255 19.3944
R9306 GND.n2255 GND.n2254 19.3944
R9307 GND.n2254 GND.n2232 19.3944
R9308 GND.n2250 GND.n2232 19.3944
R9309 GND.n2250 GND.n2249 19.3944
R9310 GND.n2249 GND.n2248 19.3944
R9311 GND.n2248 GND.n2238 19.3944
R9312 GND.n2244 GND.n2238 19.3944
R9313 GND.n2244 GND.n2243 19.3944
R9314 GND.n2408 GND.n2067 19.3944
R9315 GND.n2406 GND.n2405 19.3944
R9316 GND.n2357 GND.n2356 19.3944
R9317 GND.n2390 GND.n2389 19.3944
R9318 GND.n2387 GND.n2359 19.3944
R9319 GND.n2383 GND.n2359 19.3944
R9320 GND.n2383 GND.n2382 19.3944
R9321 GND.n2382 GND.n2381 19.3944
R9322 GND.n2381 GND.n2365 19.3944
R9323 GND.n2377 GND.n2365 19.3944
R9324 GND.n2377 GND.n2376 19.3944
R9325 GND.n2376 GND.n2375 19.3944
R9326 GND.n2375 GND.n2373 19.3944
R9327 GND.n2373 GND.n1999 19.3944
R9328 GND.n1999 GND.n1997 19.3944
R9329 GND.n2481 GND.n1997 19.3944
R9330 GND.n2481 GND.n1995 19.3944
R9331 GND.n2488 GND.n1995 19.3944
R9332 GND.n2488 GND.n2487 19.3944
R9333 GND.n2487 GND.n1963 19.3944
R9334 GND.n1963 GND.n1961 19.3944
R9335 GND.n2522 GND.n1961 19.3944
R9336 GND.n2522 GND.n1959 19.3944
R9337 GND.n6970 GND.n1959 19.3944
R9338 GND.n6970 GND.n6969 19.3944
R9339 GND.n6969 GND.n6968 19.3944
R9340 GND.n6968 GND.n2528 19.3944
R9341 GND.n6962 GND.n2528 19.3944
R9342 GND.n6962 GND.n6961 19.3944
R9343 GND.n6961 GND.n6960 19.3944
R9344 GND.n6960 GND.n2536 19.3944
R9345 GND.n6948 GND.n2536 19.3944
R9346 GND.n6948 GND.n6947 19.3944
R9347 GND.n6947 GND.n6946 19.3944
R9348 GND.n6946 GND.n2554 19.3944
R9349 GND.n6935 GND.n2554 19.3944
R9350 GND.n6935 GND.n6934 19.3944
R9351 GND.n6934 GND.n6933 19.3944
R9352 GND.n6933 GND.n2572 19.3944
R9353 GND.n6921 GND.n2572 19.3944
R9354 GND.n6921 GND.n6920 19.3944
R9355 GND.n6920 GND.n6919 19.3944
R9356 GND.n6919 GND.n2589 19.3944
R9357 GND.n6907 GND.n2589 19.3944
R9358 GND.n6907 GND.n6906 19.3944
R9359 GND.n6906 GND.n6905 19.3944
R9360 GND.n6905 GND.n2607 19.3944
R9361 GND.n6893 GND.n2607 19.3944
R9362 GND.n6893 GND.n6892 19.3944
R9363 GND.n6892 GND.n6891 19.3944
R9364 GND.n6891 GND.n2625 19.3944
R9365 GND.n6879 GND.n2625 19.3944
R9366 GND.n6879 GND.n6878 19.3944
R9367 GND.n6878 GND.n6877 19.3944
R9368 GND.n6877 GND.n2643 19.3944
R9369 GND.n6865 GND.n2643 19.3944
R9370 GND.n6865 GND.n6864 19.3944
R9371 GND.n6864 GND.n6863 19.3944
R9372 GND.n6863 GND.n2660 19.3944
R9373 GND.n4351 GND.n2660 19.3944
R9374 GND.n4351 GND.n3887 19.3944
R9375 GND.n4355 GND.n3887 19.3944
R9376 GND.n4355 GND.n3872 19.3944
R9377 GND.n4389 GND.n3872 19.3944
R9378 GND.n4389 GND.n3870 19.3944
R9379 GND.n4406 GND.n3870 19.3944
R9380 GND.n4406 GND.n4405 19.3944
R9381 GND.n4405 GND.n4404 19.3944
R9382 GND.n4404 GND.n4395 19.3944
R9383 GND.n4398 GND.n4395 19.3944
R9384 GND.n4398 GND.n3832 19.3944
R9385 GND.n4478 GND.n3832 19.3944
R9386 GND.n4478 GND.n3830 19.3944
R9387 GND.n4484 GND.n3830 19.3944
R9388 GND.n4484 GND.n4483 19.3944
R9389 GND.n4483 GND.n3801 19.3944
R9390 GND.n4524 GND.n3801 19.3944
R9391 GND.n4524 GND.n3799 19.3944
R9392 GND.n4528 GND.n3799 19.3944
R9393 GND.n4528 GND.n3783 19.3944
R9394 GND.n4581 GND.n3783 19.3944
R9395 GND.n4581 GND.n3781 19.3944
R9396 GND.n4585 GND.n3781 19.3944
R9397 GND.n4585 GND.n3760 19.3944
R9398 GND.n4609 GND.n3760 19.3944
R9399 GND.n4609 GND.n3758 19.3944
R9400 GND.n4615 GND.n3758 19.3944
R9401 GND.n4615 GND.n4614 19.3944
R9402 GND.n4614 GND.n3731 19.3944
R9403 GND.n4681 GND.n3731 19.3944
R9404 GND.n4681 GND.n3729 19.3944
R9405 GND.n4685 GND.n3729 19.3944
R9406 GND.n4685 GND.n3710 19.3944
R9407 GND.n4707 GND.n3710 19.3944
R9408 GND.n4707 GND.n3708 19.3944
R9409 GND.n4711 GND.n3708 19.3944
R9410 GND.n4711 GND.n3689 19.3944
R9411 GND.n4742 GND.n3689 19.3944
R9412 GND.n4742 GND.n3687 19.3944
R9413 GND.n4746 GND.n3687 19.3944
R9414 GND.n4746 GND.n3672 19.3944
R9415 GND.n4785 GND.n3672 19.3944
R9416 GND.n4785 GND.n3670 19.3944
R9417 GND.n4791 GND.n3670 19.3944
R9418 GND.n4791 GND.n4790 19.3944
R9419 GND.n4790 GND.n3643 19.3944
R9420 GND.n4858 GND.n3643 19.3944
R9421 GND.n4858 GND.n3641 19.3944
R9422 GND.n4862 GND.n3641 19.3944
R9423 GND.n4862 GND.n3623 19.3944
R9424 GND.n4885 GND.n3623 19.3944
R9425 GND.n4885 GND.n3621 19.3944
R9426 GND.n4889 GND.n3621 19.3944
R9427 GND.n4889 GND.n3601 19.3944
R9428 GND.n4919 GND.n3601 19.3944
R9429 GND.n4919 GND.n3599 19.3944
R9430 GND.n4923 GND.n3599 19.3944
R9431 GND.n4923 GND.n3584 19.3944
R9432 GND.n4962 GND.n3584 19.3944
R9433 GND.n4962 GND.n3582 19.3944
R9434 GND.n4968 GND.n3582 19.3944
R9435 GND.n4968 GND.n4967 19.3944
R9436 GND.n4967 GND.n3555 19.3944
R9437 GND.n5034 GND.n3555 19.3944
R9438 GND.n5034 GND.n3553 19.3944
R9439 GND.n5038 GND.n3553 19.3944
R9440 GND.n5038 GND.n3534 19.3944
R9441 GND.n5060 GND.n3534 19.3944
R9442 GND.n5060 GND.n3532 19.3944
R9443 GND.n5064 GND.n3532 19.3944
R9444 GND.n5064 GND.n3512 19.3944
R9445 GND.n5094 GND.n3512 19.3944
R9446 GND.n5094 GND.n3510 19.3944
R9447 GND.n5098 GND.n3510 19.3944
R9448 GND.n5098 GND.n3495 19.3944
R9449 GND.n5138 GND.n3495 19.3944
R9450 GND.n5138 GND.n3493 19.3944
R9451 GND.n5144 GND.n3493 19.3944
R9452 GND.n5144 GND.n5143 19.3944
R9453 GND.n5143 GND.n3466 19.3944
R9454 GND.n5209 GND.n3466 19.3944
R9455 GND.n5209 GND.n3464 19.3944
R9456 GND.n5213 GND.n3464 19.3944
R9457 GND.n5213 GND.n3445 19.3944
R9458 GND.n5235 GND.n3445 19.3944
R9459 GND.n5235 GND.n3443 19.3944
R9460 GND.n5239 GND.n3443 19.3944
R9461 GND.n5239 GND.n3423 19.3944
R9462 GND.n5269 GND.n3423 19.3944
R9463 GND.n5269 GND.n3421 19.3944
R9464 GND.n5273 GND.n3421 19.3944
R9465 GND.n5273 GND.n3406 19.3944
R9466 GND.n5312 GND.n3406 19.3944
R9467 GND.n5312 GND.n3404 19.3944
R9468 GND.n5318 GND.n3404 19.3944
R9469 GND.n5318 GND.n5317 19.3944
R9470 GND.n5317 GND.n3377 19.3944
R9471 GND.n5386 GND.n3377 19.3944
R9472 GND.n5386 GND.n3375 19.3944
R9473 GND.n5390 GND.n3375 19.3944
R9474 GND.n5390 GND.n3358 19.3944
R9475 GND.n5412 GND.n3358 19.3944
R9476 GND.n5412 GND.n3356 19.3944
R9477 GND.n5416 GND.n3356 19.3944
R9478 GND.n5416 GND.n3337 19.3944
R9479 GND.n5447 GND.n3337 19.3944
R9480 GND.n5447 GND.n3335 19.3944
R9481 GND.n5451 GND.n3335 19.3944
R9482 GND.n5451 GND.n3320 19.3944
R9483 GND.n5490 GND.n3320 19.3944
R9484 GND.n5490 GND.n3318 19.3944
R9485 GND.n5496 GND.n3318 19.3944
R9486 GND.n5496 GND.n5495 19.3944
R9487 GND.n5495 GND.n3291 19.3944
R9488 GND.n5540 GND.n3291 19.3944
R9489 GND.n5540 GND.n3289 19.3944
R9490 GND.n5546 GND.n3289 19.3944
R9491 GND.n5546 GND.n5545 19.3944
R9492 GND.n5545 GND.n3271 19.3944
R9493 GND.n5568 GND.n3271 19.3944
R9494 GND.n5568 GND.n3269 19.3944
R9495 GND.n5583 GND.n3269 19.3944
R9496 GND.n5583 GND.n5582 19.3944
R9497 GND.n5582 GND.n5581 19.3944
R9498 GND.n5581 GND.n5576 19.3944
R9499 GND.n5576 GND.n2908 19.3944
R9500 GND.n6623 GND.n2908 19.3944
R9501 GND.n6623 GND.n6622 19.3944
R9502 GND.n6622 GND.n6621 19.3944
R9503 GND.n6621 GND.n2912 19.3944
R9504 GND.n6609 GND.n2912 19.3944
R9505 GND.n6609 GND.n6608 19.3944
R9506 GND.n6608 GND.n6607 19.3944
R9507 GND.n6607 GND.n2929 19.3944
R9508 GND.n6595 GND.n2929 19.3944
R9509 GND.n6595 GND.n6594 19.3944
R9510 GND.n6594 GND.n6593 19.3944
R9511 GND.n6593 GND.n2947 19.3944
R9512 GND.n6581 GND.n2947 19.3944
R9513 GND.n6581 GND.n6580 19.3944
R9514 GND.n6580 GND.n6579 19.3944
R9515 GND.n6579 GND.n2965 19.3944
R9516 GND.n6567 GND.n2965 19.3944
R9517 GND.n6567 GND.n6566 19.3944
R9518 GND.n6566 GND.n6565 19.3944
R9519 GND.n6565 GND.n2983 19.3944
R9520 GND.n6553 GND.n2983 19.3944
R9521 GND.n6553 GND.n6552 19.3944
R9522 GND.n6552 GND.n6551 19.3944
R9523 GND.n6551 GND.n3000 19.3944
R9524 GND.n6539 GND.n3000 19.3944
R9525 GND.n6539 GND.n6538 19.3944
R9526 GND.n6538 GND.n6537 19.3944
R9527 GND.n6537 GND.n3018 19.3944
R9528 GND.n6525 GND.n3018 19.3944
R9529 GND.n6525 GND.n6524 19.3944
R9530 GND.n6524 GND.n6523 19.3944
R9531 GND.n6523 GND.n3035 19.3944
R9532 GND.n6517 GND.n3035 19.3944
R9533 GND.n6517 GND.n6516 19.3944
R9534 GND.n6516 GND.n6515 19.3944
R9535 GND.n6515 GND.n3044 19.3944
R9536 GND.n5995 GND.n3044 19.3944
R9537 GND.n5999 GND.n5995 19.3944
R9538 GND.n5999 GND.n5993 19.3944
R9539 GND.n6003 GND.n5993 19.3944
R9540 GND.n6003 GND.n5991 19.3944
R9541 GND.n6007 GND.n5991 19.3944
R9542 GND.n6007 GND.n5989 19.3944
R9543 GND.n6011 GND.n5989 19.3944
R9544 GND.n6011 GND.n5987 19.3944
R9545 GND.n6015 GND.n5987 19.3944
R9546 GND.n6015 GND.n5985 19.3944
R9547 GND.n6019 GND.n5985 19.3944
R9548 GND.n6019 GND.n5983 19.3944
R9549 GND.n6023 GND.n5983 19.3944
R9550 GND.n6023 GND.n5981 19.3944
R9551 GND.n6027 GND.n5981 19.3944
R9552 GND.n6027 GND.n5979 19.3944
R9553 GND.n6033 GND.n5979 19.3944
R9554 GND.n6033 GND.n6032 19.3944
R9555 GND.n6385 GND.n5929 19.3944
R9556 GND.n6383 GND.n6382 19.3944
R9557 GND.n6370 GND.n5946 19.3944
R9558 GND.n6368 GND.n6367 19.3944
R9559 GND.n6364 GND.n6363 19.3944
R9560 GND.n6363 GND.n6362 19.3944
R9561 GND.n6362 GND.n5951 19.3944
R9562 GND.n6358 GND.n5951 19.3944
R9563 GND.n6358 GND.n6357 19.3944
R9564 GND.n6357 GND.n6356 19.3944
R9565 GND.n6356 GND.n5957 19.3944
R9566 GND.n6314 GND.n5957 19.3944
R9567 GND.n6318 GND.n6314 19.3944
R9568 GND.n6318 GND.n6312 19.3944
R9569 GND.n6322 GND.n6312 19.3944
R9570 GND.n6322 GND.n6310 19.3944
R9571 GND.n6332 GND.n6310 19.3944
R9572 GND.n6332 GND.n6331 19.3944
R9573 GND.n6331 GND.n6330 19.3944
R9574 GND.n6330 GND.n256 19.3944
R9575 GND.n8443 GND.n256 19.3944
R9576 GND.n8443 GND.n8442 19.3944
R9577 GND.n8442 GND.n8441 19.3944
R9578 GND.n8441 GND.n260 19.3944
R9579 GND.n8435 GND.n260 19.3944
R9580 GND.n8435 GND.n8434 19.3944
R9581 GND.n8434 GND.n8433 19.3944
R9582 GND.n8433 GND.n390 19.3944
R9583 GND.n8427 GND.n390 19.3944
R9584 GND.n8427 GND.n8426 19.3944
R9585 GND.n8426 GND.n8425 19.3944
R9586 GND.n8425 GND.n398 19.3944
R9587 GND.n8419 GND.n398 19.3944
R9588 GND.n8419 GND.n8418 19.3944
R9589 GND.n8418 GND.n8417 19.3944
R9590 GND.n8417 GND.n406 19.3944
R9591 GND.n8411 GND.n406 19.3944
R9592 GND.n8411 GND.n8410 19.3944
R9593 GND.n8410 GND.n8409 19.3944
R9594 GND.n8409 GND.n414 19.3944
R9595 GND.n8403 GND.n414 19.3944
R9596 GND.n8403 GND.n8402 19.3944
R9597 GND.n8402 GND.n8401 19.3944
R9598 GND.n8401 GND.n422 19.3944
R9599 GND.n7176 GND.n7175 19.3944
R9600 GND.n7175 GND.n7174 19.3944
R9601 GND.n7174 GND.n7173 19.3944
R9602 GND.n7173 GND.n7171 19.3944
R9603 GND.n7171 GND.n7168 19.3944
R9604 GND.n7168 GND.n7167 19.3944
R9605 GND.n7167 GND.n7164 19.3944
R9606 GND.n7164 GND.n7163 19.3944
R9607 GND.n7159 GND.n7156 19.3944
R9608 GND.n7156 GND.n7155 19.3944
R9609 GND.n7155 GND.n7152 19.3944
R9610 GND.n7152 GND.n7151 19.3944
R9611 GND.n7151 GND.n7148 19.3944
R9612 GND.n7148 GND.n7147 19.3944
R9613 GND.n7147 GND.n7144 19.3944
R9614 GND.n7144 GND.n7143 19.3944
R9615 GND.n7143 GND.n7140 19.3944
R9616 GND.n7138 GND.n7136 19.3944
R9617 GND.n7136 GND.n7133 19.3944
R9618 GND.n7133 GND.n7132 19.3944
R9619 GND.n7132 GND.n7129 19.3944
R9620 GND.n7129 GND.n7128 19.3944
R9621 GND.n7128 GND.n7125 19.3944
R9622 GND.n7125 GND.n7124 19.3944
R9623 GND.n7124 GND.n7121 19.3944
R9624 GND.n7121 GND.n7120 19.3944
R9625 GND.n2171 GND.n2168 19.3944
R9626 GND.n2171 GND.n2149 19.3944
R9627 GND.n2271 GND.n2149 19.3944
R9628 GND.n2271 GND.n2147 19.3944
R9629 GND.n2277 GND.n2147 19.3944
R9630 GND.n2277 GND.n2276 19.3944
R9631 GND.n2276 GND.n2126 19.3944
R9632 GND.n2295 GND.n2126 19.3944
R9633 GND.n2295 GND.n2124 19.3944
R9634 GND.n2301 GND.n2124 19.3944
R9635 GND.n2301 GND.n2300 19.3944
R9636 GND.n2300 GND.n2103 19.3944
R9637 GND.n2320 GND.n2103 19.3944
R9638 GND.n2320 GND.n2101 19.3944
R9639 GND.n2324 GND.n2101 19.3944
R9640 GND.n2324 GND.n2054 19.3944
R9641 GND.n2416 GND.n2054 19.3944
R9642 GND.n2053 GND.n2052 19.3944
R9643 GND.n2077 GND.n2052 19.3944
R9644 GND.n2400 GND.n2399 19.3944
R9645 GND.n2348 GND.n2347 19.3944
R9646 GND.n2421 GND.n2046 19.3944
R9647 GND.n2421 GND.n2420 19.3944
R9648 GND.n2420 GND.n2026 19.3944
R9649 GND.n2441 GND.n2026 19.3944
R9650 GND.n2441 GND.n2024 19.3944
R9651 GND.n2447 GND.n2024 19.3944
R9652 GND.n2447 GND.n2446 19.3944
R9653 GND.n2446 GND.n2005 19.3944
R9654 GND.n2470 GND.n2005 19.3944
R9655 GND.n2470 GND.n2003 19.3944
R9656 GND.n2474 GND.n2003 19.3944
R9657 GND.n2474 GND.n1974 19.3944
R9658 GND.n2503 GND.n1974 19.3944
R9659 GND.n2503 GND.n1972 19.3944
R9660 GND.n2509 GND.n1972 19.3944
R9661 GND.n2509 GND.n2508 19.3944
R9662 GND.n2508 GND.n1386 19.3944
R9663 GND.n7042 GND.n1386 19.3944
R9664 GND.n7370 GND.n7369 19.3944
R9665 GND.n7369 GND.n1038 19.3944
R9666 GND.n7363 GND.n1038 19.3944
R9667 GND.n7363 GND.n7362 19.3944
R9668 GND.n7362 GND.n7361 19.3944
R9669 GND.n7361 GND.n1046 19.3944
R9670 GND.n7355 GND.n1046 19.3944
R9671 GND.n7355 GND.n7354 19.3944
R9672 GND.n7354 GND.n7353 19.3944
R9673 GND.n7353 GND.n1054 19.3944
R9674 GND.n7347 GND.n1054 19.3944
R9675 GND.n7347 GND.n7346 19.3944
R9676 GND.n7346 GND.n7345 19.3944
R9677 GND.n7345 GND.n1062 19.3944
R9678 GND.n7339 GND.n1062 19.3944
R9679 GND.n7339 GND.n7338 19.3944
R9680 GND.n7338 GND.n7337 19.3944
R9681 GND.n7337 GND.n1070 19.3944
R9682 GND.n7331 GND.n1070 19.3944
R9683 GND.n7331 GND.n7330 19.3944
R9684 GND.n7330 GND.n7329 19.3944
R9685 GND.n7329 GND.n1078 19.3944
R9686 GND.n7323 GND.n1078 19.3944
R9687 GND.n7323 GND.n7322 19.3944
R9688 GND.n7322 GND.n7321 19.3944
R9689 GND.n7321 GND.n1086 19.3944
R9690 GND.n7315 GND.n1086 19.3944
R9691 GND.n7315 GND.n7314 19.3944
R9692 GND.n7314 GND.n7313 19.3944
R9693 GND.n7313 GND.n1094 19.3944
R9694 GND.n7307 GND.n1094 19.3944
R9695 GND.n7307 GND.n7306 19.3944
R9696 GND.n7306 GND.n7305 19.3944
R9697 GND.n7305 GND.n1102 19.3944
R9698 GND.n7299 GND.n1102 19.3944
R9699 GND.n7299 GND.n7298 19.3944
R9700 GND.n7298 GND.n7297 19.3944
R9701 GND.n7297 GND.n1110 19.3944
R9702 GND.n7291 GND.n1110 19.3944
R9703 GND.n7291 GND.n7290 19.3944
R9704 GND.n7290 GND.n7289 19.3944
R9705 GND.n7289 GND.n1118 19.3944
R9706 GND.n7283 GND.n1118 19.3944
R9707 GND.n7283 GND.n7282 19.3944
R9708 GND.n7282 GND.n7281 19.3944
R9709 GND.n7281 GND.n1126 19.3944
R9710 GND.n7275 GND.n1126 19.3944
R9711 GND.n7275 GND.n7274 19.3944
R9712 GND.n7274 GND.n7273 19.3944
R9713 GND.n7273 GND.n1134 19.3944
R9714 GND.n7267 GND.n1134 19.3944
R9715 GND.n7267 GND.n7266 19.3944
R9716 GND.n7266 GND.n7265 19.3944
R9717 GND.n7265 GND.n1142 19.3944
R9718 GND.n7259 GND.n1142 19.3944
R9719 GND.n7259 GND.n7258 19.3944
R9720 GND.n7258 GND.n7257 19.3944
R9721 GND.n7257 GND.n1150 19.3944
R9722 GND.n7251 GND.n1150 19.3944
R9723 GND.n7251 GND.n7250 19.3944
R9724 GND.n7250 GND.n7249 19.3944
R9725 GND.n7249 GND.n1158 19.3944
R9726 GND.n7243 GND.n1158 19.3944
R9727 GND.n7243 GND.n7242 19.3944
R9728 GND.n7242 GND.n7241 19.3944
R9729 GND.n7241 GND.n1166 19.3944
R9730 GND.n7235 GND.n1166 19.3944
R9731 GND.n7235 GND.n7234 19.3944
R9732 GND.n7234 GND.n7233 19.3944
R9733 GND.n7233 GND.n1174 19.3944
R9734 GND.n7227 GND.n1174 19.3944
R9735 GND.n7227 GND.n7226 19.3944
R9736 GND.n6663 GND.n6662 19.3944
R9737 GND.n6662 GND.n6661 19.3944
R9738 GND.n6661 GND.n2832 19.3944
R9739 GND.n6657 GND.n2832 19.3944
R9740 GND.n6657 GND.n6656 19.3944
R9741 GND.n6656 GND.n6655 19.3944
R9742 GND.n6655 GND.n2877 19.3944
R9743 GND.n6651 GND.n2877 19.3944
R9744 GND.n6651 GND.n6650 19.3944
R9745 GND.n6650 GND.n6649 19.3944
R9746 GND.n6649 GND.n2882 19.3944
R9747 GND.n6645 GND.n2882 19.3944
R9748 GND.n6645 GND.n6644 19.3944
R9749 GND.n6644 GND.n6643 19.3944
R9750 GND.n6643 GND.n2887 19.3944
R9751 GND.n6639 GND.n2887 19.3944
R9752 GND.n6639 GND.n6638 19.3944
R9753 GND.n6638 GND.n6637 19.3944
R9754 GND.n6634 GND.n6633 19.3944
R9755 GND.n6633 GND.n6632 19.3944
R9756 GND.n6632 GND.n2899 19.3944
R9757 GND.n6858 GND.n2667 19.3944
R9758 GND.n6854 GND.n2667 19.3944
R9759 GND.n6854 GND.n6853 19.3944
R9760 GND.n6853 GND.n6852 19.3944
R9761 GND.n6852 GND.n2673 19.3944
R9762 GND.n6848 GND.n2673 19.3944
R9763 GND.n6848 GND.n6847 19.3944
R9764 GND.n6847 GND.n6846 19.3944
R9765 GND.n6846 GND.n2678 19.3944
R9766 GND.n6842 GND.n2678 19.3944
R9767 GND.n6842 GND.n6841 19.3944
R9768 GND.n6841 GND.n6840 19.3944
R9769 GND.n6840 GND.n2683 19.3944
R9770 GND.n6836 GND.n2683 19.3944
R9771 GND.n6836 GND.n6835 19.3944
R9772 GND.n6835 GND.n6834 19.3944
R9773 GND.n6834 GND.n2688 19.3944
R9774 GND.n6830 GND.n2688 19.3944
R9775 GND.n6830 GND.n6829 19.3944
R9776 GND.n6829 GND.n6828 19.3944
R9777 GND.n6828 GND.n2693 19.3944
R9778 GND.n6824 GND.n2693 19.3944
R9779 GND.n6824 GND.n6823 19.3944
R9780 GND.n6823 GND.n6822 19.3944
R9781 GND.n6822 GND.n2698 19.3944
R9782 GND.n6818 GND.n2698 19.3944
R9783 GND.n6818 GND.n6817 19.3944
R9784 GND.n6817 GND.n6816 19.3944
R9785 GND.n6816 GND.n2703 19.3944
R9786 GND.n6812 GND.n2703 19.3944
R9787 GND.n6812 GND.n6811 19.3944
R9788 GND.n6811 GND.n6810 19.3944
R9789 GND.n6810 GND.n2708 19.3944
R9790 GND.n6806 GND.n2708 19.3944
R9791 GND.n6806 GND.n6805 19.3944
R9792 GND.n6805 GND.n6804 19.3944
R9793 GND.n6804 GND.n2713 19.3944
R9794 GND.n6800 GND.n2713 19.3944
R9795 GND.n6800 GND.n6799 19.3944
R9796 GND.n6799 GND.n6798 19.3944
R9797 GND.n6798 GND.n2718 19.3944
R9798 GND.n6794 GND.n2718 19.3944
R9799 GND.n6794 GND.n6793 19.3944
R9800 GND.n6793 GND.n6792 19.3944
R9801 GND.n6792 GND.n2723 19.3944
R9802 GND.n6788 GND.n2723 19.3944
R9803 GND.n6788 GND.n6787 19.3944
R9804 GND.n6787 GND.n6786 19.3944
R9805 GND.n6786 GND.n2728 19.3944
R9806 GND.n6782 GND.n2728 19.3944
R9807 GND.n6782 GND.n6781 19.3944
R9808 GND.n6781 GND.n6780 19.3944
R9809 GND.n6780 GND.n2733 19.3944
R9810 GND.n6776 GND.n2733 19.3944
R9811 GND.n6776 GND.n6775 19.3944
R9812 GND.n6775 GND.n6774 19.3944
R9813 GND.n6774 GND.n2738 19.3944
R9814 GND.n6770 GND.n2738 19.3944
R9815 GND.n6770 GND.n6769 19.3944
R9816 GND.n6769 GND.n6768 19.3944
R9817 GND.n6768 GND.n2743 19.3944
R9818 GND.n6764 GND.n2743 19.3944
R9819 GND.n6764 GND.n6763 19.3944
R9820 GND.n6763 GND.n6762 19.3944
R9821 GND.n6762 GND.n2748 19.3944
R9822 GND.n6758 GND.n2748 19.3944
R9823 GND.n6758 GND.n6757 19.3944
R9824 GND.n6757 GND.n6756 19.3944
R9825 GND.n6756 GND.n2753 19.3944
R9826 GND.n6752 GND.n2753 19.3944
R9827 GND.n6752 GND.n6751 19.3944
R9828 GND.n6751 GND.n6750 19.3944
R9829 GND.n6750 GND.n2758 19.3944
R9830 GND.n6746 GND.n2758 19.3944
R9831 GND.n6746 GND.n6745 19.3944
R9832 GND.n6745 GND.n6744 19.3944
R9833 GND.n6744 GND.n2763 19.3944
R9834 GND.n6740 GND.n2763 19.3944
R9835 GND.n6740 GND.n6739 19.3944
R9836 GND.n6739 GND.n6738 19.3944
R9837 GND.n6738 GND.n2768 19.3944
R9838 GND.n6734 GND.n2768 19.3944
R9839 GND.n6734 GND.n6733 19.3944
R9840 GND.n6733 GND.n6732 19.3944
R9841 GND.n6732 GND.n2773 19.3944
R9842 GND.n6728 GND.n2773 19.3944
R9843 GND.n6728 GND.n6727 19.3944
R9844 GND.n6727 GND.n6726 19.3944
R9845 GND.n6726 GND.n2778 19.3944
R9846 GND.n6722 GND.n2778 19.3944
R9847 GND.n6722 GND.n6721 19.3944
R9848 GND.n6721 GND.n6720 19.3944
R9849 GND.n6720 GND.n2783 19.3944
R9850 GND.n6716 GND.n2783 19.3944
R9851 GND.n6716 GND.n6715 19.3944
R9852 GND.n6715 GND.n6714 19.3944
R9853 GND.n6714 GND.n2788 19.3944
R9854 GND.n6710 GND.n2788 19.3944
R9855 GND.n6710 GND.n6709 19.3944
R9856 GND.n6709 GND.n6708 19.3944
R9857 GND.n6708 GND.n2793 19.3944
R9858 GND.n6704 GND.n2793 19.3944
R9859 GND.n6704 GND.n6703 19.3944
R9860 GND.n6703 GND.n6702 19.3944
R9861 GND.n6702 GND.n2798 19.3944
R9862 GND.n6698 GND.n2798 19.3944
R9863 GND.n6698 GND.n6697 19.3944
R9864 GND.n6697 GND.n6696 19.3944
R9865 GND.n6696 GND.n2803 19.3944
R9866 GND.n6692 GND.n2803 19.3944
R9867 GND.n6692 GND.n6691 19.3944
R9868 GND.n6691 GND.n6690 19.3944
R9869 GND.n6690 GND.n2808 19.3944
R9870 GND.n6686 GND.n2808 19.3944
R9871 GND.n6686 GND.n6685 19.3944
R9872 GND.n6685 GND.n6684 19.3944
R9873 GND.n6684 GND.n2813 19.3944
R9874 GND.n6680 GND.n2813 19.3944
R9875 GND.n6680 GND.n6679 19.3944
R9876 GND.n6679 GND.n6678 19.3944
R9877 GND.n6678 GND.n2818 19.3944
R9878 GND.n6674 GND.n2818 19.3944
R9879 GND.n6674 GND.n6673 19.3944
R9880 GND.n6673 GND.n6672 19.3944
R9881 GND.n6672 GND.n2823 19.3944
R9882 GND.n6668 GND.n2823 19.3944
R9883 GND.n6668 GND.n6667 19.3944
R9884 GND.n6667 GND.n6666 19.3944
R9885 GND.t136 GND.n2556 19.1971
R9886 GND.n4145 GND.n2591 19.1971
R9887 GND.n6888 GND.n2629 19.1971
R9888 GND.n6598 GND.n2939 19.1971
R9889 GND.n5687 GND.n2977 19.1971
R9890 GND.n6541 GND.n3012 19.1971
R9891 GND.n1775 GND.n1774 19.0848
R9892 GND.n1832 GND.n1831 19.0848
R9893 GND.n1714 GND.n1713 19.0848
R9894 GND.n1771 GND.n1770 19.0848
R9895 GND.n1653 GND.n1652 19.0848
R9896 GND.n1710 GND.n1709 19.0848
R9897 GND.n1592 GND.n1591 19.0848
R9898 GND.n1649 GND.n1648 19.0848
R9899 GND.n3967 GND.n3963 18.7329
R9900 GND.n3111 GND.n3110 18.7329
R9901 GND.n7021 GND.n7020 18.6187
R9902 GND.n6488 GND.n6485 18.6187
R9903 GND.n1561 GND.n1560 18.5954
R9904 GND.n1543 GND.n1542 18.5954
R9905 GND.n1583 GND.n1582 18.5954
R9906 GND.n1565 GND.n1564 18.5954
R9907 GND.n1855 GND.n1854 18.5954
R9908 GND.n1837 GND.n1836 18.5954
R9909 GND.n1585 GND.n1439 18.5954
R9910 GND.n1859 GND.n1444 18.5954
R9911 GND.n1793 GND.n1792 18.1061
R9912 GND.n1814 GND.n1813 18.1061
R9913 GND.n1732 GND.n1731 18.1061
R9914 GND.n1753 GND.n1752 18.1061
R9915 GND.n1671 GND.n1670 18.1061
R9916 GND.n1692 GND.n1691 18.1061
R9917 GND.n1610 GND.n1609 18.1061
R9918 GND.n1631 GND.n1630 18.1061
R9919 GND.n6938 GND.n6937 17.8732
R9920 GND.n6924 GND.n2581 17.8732
R9921 GND.n4184 GND.n2637 17.8732
R9922 GND.n6867 GND.n2654 17.8732
R9923 GND.n6619 GND.n2914 17.8732
R9924 GND.n5648 GND.n2931 17.8732
R9925 GND.n6562 GND.n2987 17.8732
R9926 GND.n6549 GND.n6548 17.8732
R9927 GND.n7026 GND.n7025 17.2611
R9928 GND.n6493 GND.n6492 17.2611
R9929 GND.n362 GND.n287 17.2611
R9930 GND.n7160 GND.n7159 17.2611
R9931 GND.n7113 GND.n1292 17.2113
R9932 GND.n2218 GND.n2173 17.2113
R9933 GND.n2217 GND.n2151 17.2113
R9934 GND.n2266 GND.n2141 17.2113
R9935 GND.n2279 GND.n2142 17.2113
R9936 GND.n2145 GND.n2134 17.2113
R9937 GND.n2288 GND.n2128 17.2113
R9938 GND.n2293 GND.n2131 17.2113
R9939 GND.n2290 GND.n2117 17.2113
R9940 GND.n2303 GND.n2118 17.2113
R9941 GND.n2122 GND.n2109 17.2113
R9942 GND.n2312 GND.n2105 17.2113
R9943 GND.n2318 GND.n2107 17.2113
R9944 GND.n2315 GND.n2095 17.2113
R9945 GND.n2326 GND.n2098 17.2113
R9946 GND.n2414 GND.n2059 17.2113
R9947 GND.n2411 GND.n2410 17.2113
R9948 GND.n2070 GND.n2064 17.2113
R9949 GND.n2403 GND.n2072 17.2113
R9950 GND.n2397 GND.n2082 17.2113
R9951 GND.n2393 GND.n2392 17.2113
R9952 GND.n2354 GND.n2350 17.2113
R9953 GND.n2353 GND.n2039 17.2113
R9954 GND.n2423 GND.n2040 17.2113
R9955 GND.n2044 GND.n2032 17.2113
R9956 GND.n2433 GND.n2028 17.2113
R9957 GND.n2439 GND.n2030 17.2113
R9958 GND.n2436 GND.n2017 17.2113
R9959 GND.n2449 GND.n2018 17.2113
R9960 GND.n2463 GND.n2007 17.2113
R9961 GND.n2468 GND.n2009 17.2113
R9962 GND.n2477 GND.n2000 17.2113
R9963 GND.n2476 GND.n1980 17.2113
R9964 GND.n2497 GND.n1976 17.2113
R9965 GND.n2501 GND.n1978 17.2113
R9966 GND.n2491 GND.n2490 17.2113
R9967 GND.n2511 GND.n1969 17.2113
R9968 GND.n2518 GND.n1964 17.2113
R9969 GND.n2517 GND.n1380 17.2113
R9970 GND.n7044 GND.n1382 17.2113
R9971 GND.n6448 GND.n5819 17.2113
R9972 GND.n6051 GND.n5821 17.2113
R9973 GND.n6440 GND.n5829 17.2113
R9974 GND.n6138 GND.n5831 17.2113
R9975 GND.n6434 GND.n5844 17.2113
R9976 GND.n6146 GND.n5847 17.2113
R9977 GND.n6428 GND.n5857 17.2113
R9978 GND.n6153 GND.n5860 17.2113
R9979 GND.n6422 GND.n5868 17.2113
R9980 GND.n6161 GND.n5871 17.2113
R9981 GND.n6416 GND.n5878 17.2113
R9982 GND.n6410 GND.n5889 17.2113
R9983 GND.n6176 GND.n5892 17.2113
R9984 GND.n6404 GND.n5899 17.2113
R9985 GND.n6183 GND.n5902 17.2113
R9986 GND.n6398 GND.n5909 17.2113
R9987 GND.n6198 GND.n6035 17.2113
R9988 GND.n6392 GND.n5918 17.2113
R9989 GND.n6388 GND.n5921 17.2113
R9990 GND.n6387 GND.n5926 17.2113
R9991 GND.n6379 GND.n5932 17.2113
R9992 GND.n6373 GND.n143 17.2113
R9993 GND.n6372 GND.n5944 17.2113
R9994 GND.n6215 GND.n5974 17.2113
R9995 GND.n8501 GND.n160 17.2113
R9996 GND.n8495 GND.n172 17.2113
R9997 GND.n6230 GND.n175 17.2113
R9998 GND.n8489 GND.n182 17.2113
R9999 GND.n6239 GND.n185 17.2113
R10000 GND.n8483 GND.n192 17.2113
R10001 GND.n6354 GND.n6353 17.2113
R10002 GND.n8477 GND.n202 17.2113
R10003 GND.n6347 GND.n205 17.2113
R10004 GND.n8471 GND.n212 17.2113
R10005 GND.n6341 GND.n215 17.2113
R10006 GND.n8465 GND.n223 17.2113
R10007 GND.n6335 GND.n226 17.2113
R10008 GND.n6302 GND.n235 17.2113
R10009 GND.n8453 GND.n243 17.2113
R10010 GND.n8446 GND.n246 17.2113
R10011 GND.n2402 GND.t12 16.5493
R10012 GND.n4131 GND.n2574 16.5493
R10013 GND.n6931 GND.n2574 16.5493
R10014 GND.n6875 GND.n6874 16.5493
R10015 GND.n6874 GND.n2647 16.5493
R10016 GND.n6861 GND.n6860 16.5493
R10017 GND.n4349 GND.n4348 16.5493
R10018 GND.n4357 GND.n3881 16.5493
R10019 GND.n4387 GND.n3875 16.5493
R10020 GND.n4409 GND.n4408 16.5493
R10021 GND.n4364 GND.n3851 16.5493
R10022 GND.n4400 GND.n3847 16.5493
R10023 GND.n4468 GND.n3835 16.5493
R10024 GND.n4476 GND.n3835 16.5493
R10025 GND.n4460 GND.n3826 16.5493
R10026 GND.n4452 GND.n3822 16.5493
R10027 GND.n4522 GND.n4521 16.5493
R10028 GND.n4530 GND.n3793 16.5493
R10029 GND.n4579 GND.n3785 16.5493
R10030 GND.n4588 GND.n4587 16.5493
R10031 GND.n4618 GND.n4617 16.5493
R10032 GND.n4544 GND.n3750 16.5493
R10033 GND.n4544 GND.n3740 16.5493
R10034 GND.n4679 GND.n4678 16.5493
R10035 GND.n4687 GND.n3727 16.5493
R10036 GND.n4705 GND.n4704 16.5493
R10037 GND.n4713 GND.n3699 16.5493
R10038 GND.n4740 GND.n3691 16.5493
R10039 GND.n4748 GND.n3685 16.5493
R10040 GND.n4783 GND.n3674 16.5493
R10041 GND.n4795 GND.n4793 16.5493
R10042 GND.n4761 GND.n3662 16.5493
R10043 GND.n4761 GND.n3652 16.5493
R10044 GND.n4856 GND.n4855 16.5493
R10045 GND.n4864 GND.n3639 16.5493
R10046 GND.n4883 GND.n4882 16.5493
R10047 GND.n4891 GND.n3612 16.5493
R10048 GND.n4917 GND.n3603 16.5493
R10049 GND.n4925 GND.n3597 16.5493
R10050 GND.n4960 GND.n3586 16.5493
R10051 GND.n4971 GND.n4970 16.5493
R10052 GND.n4938 GND.n3574 16.5493
R10053 GND.n4938 GND.n3564 16.5493
R10054 GND.n5032 GND.n5031 16.5493
R10055 GND.n5040 GND.n3551 16.5493
R10056 GND.n5058 GND.n5057 16.5493
R10057 GND.n5066 GND.n3523 16.5493
R10058 GND.n5092 GND.n3515 16.5493
R10059 GND.n5100 GND.n3508 16.5493
R10060 GND.n5136 GND.n3498 16.5493
R10061 GND.n5147 GND.n5146 16.5493
R10062 GND.n5114 GND.n3485 16.5493
R10063 GND.n5114 GND.n3475 16.5493
R10064 GND.n5207 GND.n5206 16.5493
R10065 GND.n5215 GND.n3462 16.5493
R10066 GND.n5233 GND.n5232 16.5493
R10067 GND.n5241 GND.n3434 16.5493
R10068 GND.n5267 GND.n3425 16.5493
R10069 GND.n5275 GND.n3419 16.5493
R10070 GND.n5310 GND.n3408 16.5493
R10071 GND.n5321 GND.n5320 16.5493
R10072 GND.n5288 GND.n3396 16.5493
R10073 GND.n5288 GND.n3386 16.5493
R10074 GND.n5384 GND.n5383 16.5493
R10075 GND.n5410 GND.n5409 16.5493
R10076 GND.n5418 GND.n3347 16.5493
R10077 GND.n5445 GND.n3339 16.5493
R10078 GND.n5453 GND.n3333 16.5493
R10079 GND.n5488 GND.n3322 16.5493
R10080 GND.n5500 GND.n5498 16.5493
R10081 GND.n5466 GND.n3310 16.5493
R10082 GND.n5466 GND.n3300 16.5493
R10083 GND.n5538 GND.n5537 16.5493
R10084 GND.n5548 GND.n3287 16.5493
R10085 GND.n5565 GND.n5564 16.5493
R10086 GND.n5602 GND.n3258 16.5493
R10087 GND.n5586 GND.n3249 16.5493
R10088 GND.n5578 GND.n3245 16.5493
R10089 GND.n6626 GND.n6625 16.5493
R10090 GND.n6612 GND.n2921 16.5493
R10091 GND.n6612 GND.n6611 16.5493
R10092 GND.n6555 GND.n2994 16.5493
R10093 GND.n5701 GND.n2994 16.5493
R10094 GND.n8508 GND.t0 16.5493
R10095 GND.n7113 GND.n1290 15.8874
R10096 GND.n2173 GND.n1292 15.8874
R10097 GND.n2218 GND.n2217 15.8874
R10098 GND.n2269 GND.n2151 15.8874
R10099 GND.n2266 GND.n2264 15.8874
R10100 GND.n2279 GND.n2141 15.8874
R10101 GND.n2145 GND.n2142 15.8874
R10102 GND.n2288 GND.n2134 15.8874
R10103 GND.n2293 GND.n2128 15.8874
R10104 GND.n2290 GND.n2131 15.8874
R10105 GND.n2303 GND.n2117 15.8874
R10106 GND.n2312 GND.n2109 15.8874
R10107 GND.n2318 GND.n2105 15.8874
R10108 GND.n2315 GND.n2107 15.8874
R10109 GND.n2326 GND.n2095 15.8874
R10110 GND.n2098 GND.n2097 15.8874
R10111 GND.n2414 GND.n2057 15.8874
R10112 GND.n2411 GND.n2059 15.8874
R10113 GND.n2410 GND.n2064 15.8874
R10114 GND.n2072 GND.n2070 15.8874
R10115 GND.n2403 GND.n2402 15.8874
R10116 GND.n2397 GND.n2080 15.8874
R10117 GND.n2393 GND.n2082 15.8874
R10118 GND.n2392 GND.n2350 15.8874
R10119 GND.n2354 GND.n2353 15.8874
R10120 GND.n2423 GND.n2039 15.8874
R10121 GND.n2433 GND.n2032 15.8874
R10122 GND.n2439 GND.n2028 15.8874
R10123 GND.n2436 GND.n2030 15.8874
R10124 GND.n2449 GND.n2017 15.8874
R10125 GND.n2022 GND.n2018 15.8874
R10126 GND.n2463 GND.n2011 15.8874
R10127 GND.n2468 GND.n2007 15.8874
R10128 GND.n2009 GND.n2000 15.8874
R10129 GND.n2477 GND.n2476 15.8874
R10130 GND.n2497 GND.n1980 15.8874
R10131 GND.n2501 GND.n1976 15.8874
R10132 GND.n2491 GND.n1978 15.8874
R10133 GND.n1969 GND.n1964 15.8874
R10134 GND.n2518 GND.n2517 15.8874
R10135 GND.n7044 GND.n1380 15.8874
R10136 GND.n4358 GND.n3885 15.8874
R10137 GND.n4386 GND.n3877 15.8874
R10138 GND.n4531 GND.n3797 15.8874
R10139 GND.n4578 GND.n3787 15.8874
R10140 GND.n4739 GND.n3693 15.8874
R10141 GND.n4893 GND.n4892 15.8874
R10142 GND.n4916 GND.n3606 15.8874
R10143 GND.n5068 GND.n5067 15.8874
R10144 GND.n5091 GND.n3517 15.8874
R10145 GND.n5243 GND.n5242 15.8874
R10146 GND.n5421 GND.n5419 15.8874
R10147 GND.n5444 GND.n3341 15.8874
R10148 GND.n5594 GND.n5593 15.8874
R10149 GND.n5614 GND.n5613 15.8874
R10150 GND.n6448 GND.n5821 15.8874
R10151 GND.n6051 GND.n5829 15.8874
R10152 GND.n6440 GND.n5831 15.8874
R10153 GND.n6434 GND.n5847 15.8874
R10154 GND.n6146 GND.n5857 15.8874
R10155 GND.n6428 GND.n5860 15.8874
R10156 GND.n6153 GND.n5868 15.8874
R10157 GND.n6422 GND.n5871 15.8874
R10158 GND.n6161 GND.n5878 15.8874
R10159 GND.n6416 GND.n5881 15.8874
R10160 GND.n6168 GND.n5889 15.8874
R10161 GND.n6410 GND.n5892 15.8874
R10162 GND.n6176 GND.n5899 15.8874
R10163 GND.n6404 GND.n5902 15.8874
R10164 GND.n6183 GND.n5909 15.8874
R10165 GND.n6198 GND.n5918 15.8874
R10166 GND.n6392 GND.n5921 15.8874
R10167 GND.n6388 GND.n6387 15.8874
R10168 GND.n5932 GND.n5926 15.8874
R10169 GND.n6380 GND.n6379 15.8874
R10170 GND.n8508 GND.n143 15.8874
R10171 GND.n6373 GND.n6372 15.8874
R10172 GND.n5974 GND.n5944 15.8874
R10173 GND.n6215 GND.n160 15.8874
R10174 GND.n8501 GND.n163 15.8874
R10175 GND.n6223 GND.n172 15.8874
R10176 GND.n8495 GND.n175 15.8874
R10177 GND.n6230 GND.n182 15.8874
R10178 GND.n8489 GND.n185 15.8874
R10179 GND.n6239 GND.n192 15.8874
R10180 GND.n6353 GND.n202 15.8874
R10181 GND.n8477 GND.n205 15.8874
R10182 GND.n6347 GND.n212 15.8874
R10183 GND.n8471 GND.n215 15.8874
R10184 GND.n6341 GND.n223 15.8874
R10185 GND.n8465 GND.n226 15.8874
R10186 GND.n6335 GND.n6334 15.8874
R10187 GND.n8459 GND.n235 15.8874
R10188 GND.n6302 GND.n243 15.8874
R10189 GND.n8453 GND.n246 15.8874
R10190 GND.n8446 GND.n8445 15.8874
R10191 GND.n6938 GND.n2564 15.2254
R10192 GND.n6924 GND.n6923 15.2254
R10193 GND.n6881 GND.n2637 15.2254
R10194 GND.n4443 GND.n3846 15.2254
R10195 GND.n4487 GND.n4486 15.2254
R10196 GND.n4619 GND.n3754 15.2254
R10197 GND.n4677 GND.n3736 15.2254
R10198 GND.n4796 GND.n3666 15.2254
R10199 GND.n4853 GND.n3648 15.2254
R10200 GND.n4972 GND.n3578 15.2254
R10201 GND.n5030 GND.n3560 15.2254
R10202 GND.n5148 GND.n3489 15.2254
R10203 GND.n5205 GND.n3471 15.2254
R10204 GND.n5322 GND.n3400 15.2254
R10205 GND.n5382 GND.n3382 15.2254
R10206 GND.n5501 GND.n3314 15.2254
R10207 GND.n5535 GND.n3296 15.2254
R10208 GND.n6605 GND.n2931 15.2254
R10209 GND.n6563 GND.n6562 15.2254
R10210 GND.n6548 GND.n3004 15.2254
R10211 GND.n6527 GND.t173 15.2254
R10212 GND.n7009 GND.n1416 14.9338
R10213 GND.n6474 GND.n6473 14.9338
R10214 GND.n339 GND.n298 14.9338
R10215 GND.n7139 GND.n7138 14.9338
R10216 GND.n1452 GND.n1451 14.803
R10217 GND.n4192 GND.t8 14.5635
R10218 GND.n4339 GND.n3889 14.5635
R10219 GND.n4417 GND.n3860 14.5635
R10220 GND.n4512 GND.n3803 14.5635
R10221 GND.n3779 GND.n3768 14.5635
R10222 GND.n3718 GND.n3712 14.5635
R10223 GND.n4749 GND.n3680 14.5635
R10224 GND.n3631 GND.n3625 14.5635
R10225 GND.n5101 GND.n3504 14.5635
R10226 GND.n3453 GND.n3447 14.5635
R10227 GND.n5276 GND.n3415 14.5635
R10228 GND.n3366 GND.n3360 14.5635
R10229 GND.n5454 GND.n3328 14.5635
R10230 GND.n3279 GND.n3273 14.5635
R10231 GND.n5577 GND.n3239 14.5635
R10232 GND.n5642 GND.t22 14.5635
R10233 GND.n6054 GND.t179 14.3199
R10234 GND.n6054 GND.t97 14.3199
R10235 GND.n6053 GND.t93 14.3199
R10236 GND.n6053 GND.t132 14.3199
R10237 GND.t62 GND.n2057 13.9015
R10238 GND.n4118 GND.n2556 13.9015
R10239 GND.n6917 GND.n2591 13.9015
R10240 GND.n6889 GND.n6888 13.9015
R10241 GND.n3898 GND.n2664 13.9015
R10242 GND.n4365 GND.n3862 13.9015
R10243 GND.n4453 GND.n3812 13.9015
R10244 GND.n4599 GND.n4598 13.9015
R10245 GND.n3726 GND.n3717 13.9015
R10246 GND.n4775 GND.n4774 13.9015
R10247 GND.n3638 GND.n3630 13.9015
R10248 GND.n4952 GND.n4951 13.9015
R10249 GND.n3550 GND.n3541 13.9015
R10250 GND.n5128 GND.n5127 13.9015
R10251 GND.n3460 GND.n3452 13.9015
R10252 GND.n5302 GND.n5301 13.9015
R10253 GND.n5337 GND.n3365 13.9015
R10254 GND.n5480 GND.n5479 13.9015
R10255 GND.n3286 GND.n3278 13.9015
R10256 GND.n5629 GND.n2904 13.9015
R10257 GND.n6598 GND.n6597 13.9015
R10258 GND.n6569 GND.n2977 13.9015
R10259 GND.n5714 GND.n3012 13.9015
R10260 GND.t28 GND.n163 13.9015
R10261 GND.n1588 GND.n1587 13.507
R10262 GND.n6996 GND.n6995 13.3823
R10263 GND.n6990 GND.n1922 13.3823
R10264 GND.n2208 GND.n2207 13.3823
R10265 GND.n6455 GND.n5815 13.3823
R10266 GND.n319 GND.n316 13.3823
R10267 GND.n6295 GND.n6260 13.3823
R10268 GND.n7120 GND.n1286 13.3823
R10269 GND.n2264 GND.t111 13.2396
R10270 GND.n4121 GND.t194 13.2396
R10271 GND.n4437 GND.n4436 13.2396
R10272 GND.n4494 GND.n4493 13.2396
R10273 GND.n4606 GND.n3763 13.2396
R10274 GND.n4688 GND.n3724 13.2396
R10275 GND.n4782 GND.n3676 13.2396
R10276 GND.n4865 GND.n3636 13.2396
R10277 GND.n4959 GND.n3589 13.2396
R10278 GND.n5041 GND.n3548 13.2396
R10279 GND.n5135 GND.n3500 13.2396
R10280 GND.n5216 GND.n3458 13.2396
R10281 GND.n5309 GND.n3410 13.2396
R10282 GND.n5393 GND.n3372 13.2396
R10283 GND.n5487 GND.n3324 13.2396
R10284 GND.n5549 GND.n3284 13.2396
R10285 GND.n6334 GND.t121 13.2396
R10286 GND.n3973 GND.n3961 13.1884
R10287 GND.n3106 GND.n3105 13.1049
R10288 GND.n1912 GND.n1911 12.8005
R10289 GND.n4305 GND.n4304 12.8005
R10290 GND.n2865 GND.n2864 12.8005
R10291 GND.n6098 GND.n6097 12.8005
R10292 GND.n6995 GND.n6994 12.6066
R10293 GND.n2207 GND.n2206 12.6066
R10294 GND.n6451 GND.n5815 12.6066
R10295 GND.n316 GND.n311 12.6066
R10296 GND.n6290 GND.n6260 12.6066
R10297 GND.n6116 GND.n6115 12.6066
R10298 GND.n7116 GND.n1286 12.6066
R10299 GND.t45 GND.n2040 12.5776
R10300 GND.n6951 GND.n2546 12.5776
R10301 GND.n6910 GND.n6909 12.5776
R10302 GND.n6895 GND.n2619 12.5776
R10303 GND.n4347 GND.n3892 12.5776
R10304 GND.n4410 GND.n3866 12.5776
R10305 GND.n4520 GND.n3806 12.5776
R10306 GND.n4560 GND.n3778 12.5776
R10307 GND.n4703 GND.n3703 12.5776
R10308 GND.n4733 GND.n4732 12.5776
R10309 GND.n4880 GND.n3616 12.5776
R10310 GND.n4910 GND.n4909 12.5776
R10311 GND.n5056 GND.n3527 12.5776
R10312 GND.n5085 GND.n5084 12.5776
R10313 GND.n5231 GND.n3438 12.5776
R10314 GND.n5260 GND.n5259 12.5776
R10315 GND.n5408 GND.n3351 12.5776
R10316 GND.n5438 GND.n5437 12.5776
R10317 GND.n5562 GND.n3263 12.5776
R10318 GND.n5621 GND.n3244 12.5776
R10319 GND.n6591 GND.n2949 12.5776
R10320 GND.n6577 GND.n6576 12.5776
R10321 GND.n6035 GND.t64 12.5776
R10322 GND.n3115 GND.n3104 12.4126
R10323 GND.n6103 GND.n6065 12.349
R10324 GND.t48 GND.n3593 12.2466
R10325 GND.n3543 GND.t60 12.2466
R10326 GND.n3975 GND.n3974 12.1761
R10327 GND.n3117 GND.n3116 12.1761
R10328 GND.n1908 GND.n1882 12.0247
R10329 GND.n4301 GND.n4275 12.0247
R10330 GND.n2861 GND.n2835 12.0247
R10331 GND.n6094 GND.n6068 12.0247
R10332 GND.n2490 GND.t125 11.9156
R10333 GND.n4317 GND.n4211 11.9156
R10334 GND.n4461 GND.n3837 11.9156
R10335 GND.n4597 GND.t84 11.9156
R10336 GND.n4627 GND.n3748 11.9156
R10337 GND.n4670 GND.n3733 11.9156
R10338 GND.n4803 GND.n3660 11.9156
R10339 GND.n4846 GND.n3645 11.9156
R10340 GND.n4979 GND.n3572 11.9156
R10341 GND.n5023 GND.n3557 11.9156
R10342 GND.n5155 GND.n3483 11.9156
R10343 GND.n5198 GND.n3468 11.9156
R10344 GND.n5330 GND.n3394 11.9156
R10345 GND.n5375 GND.n3379 11.9156
R10346 GND.n5338 GND.t37 11.9156
R10347 GND.n5508 GND.n3308 11.9156
R10348 GND.n3235 GND.n3234 11.9156
R10349 GND.t99 GND.n5844 11.9156
R10350 GND.n6065 GND.n6055 11.8584
R10351 GND.n6903 GND.n2609 11.2537
R10352 GND.n6903 GND.n6902 11.2537
R10353 GND.n4380 GND.n4379 11.2537
R10354 GND.n4569 GND.n4568 11.2537
R10355 GND.n4568 GND.n4567 11.2537
R10356 GND.n4724 GND.n4723 11.2537
R10357 GND.n4725 GND.n4724 11.2537
R10358 GND.n4901 GND.n4900 11.2537
R10359 GND.n5077 GND.n5076 11.2537
R10360 GND.n5251 GND.n5250 11.2537
R10361 GND.n5252 GND.n5251 11.2537
R10362 GND.n5429 GND.n5428 11.2537
R10363 GND.n5430 GND.n5429 11.2537
R10364 GND.n5587 GND.n5585 11.2537
R10365 GND.n6584 GND.n6583 11.2537
R10366 GND.n6583 GND.n2959 11.2537
R10367 GND.n5728 GND.n5727 11.2537
R10368 GND.n1907 GND.n1884 11.249
R10369 GND.n4300 GND.n4277 11.249
R10370 GND.n2860 GND.n2837 11.249
R10371 GND.n6093 GND.n6070 11.249
R10372 GND.n7013 GND.n1416 11.055
R10373 GND.n6475 GND.n6474 11.055
R10374 GND.n340 GND.n339 11.055
R10375 GND.n7140 GND.n7139 11.055
R10376 GND.t2 GND.n4714 10.9227
R10377 GND.n5266 GND.t208 10.9227
R10378 GND.n3186 GND.n3086 10.6151
R10379 GND.n5783 GND.n3186 10.6151
R10380 GND.n5783 GND.n5782 10.6151
R10381 GND.n5780 GND.n3190 10.6151
R10382 GND.n5775 GND.n3190 10.6151
R10383 GND.n5775 GND.n5774 10.6151
R10384 GND.n5774 GND.n5773 10.6151
R10385 GND.n5773 GND.n3193 10.6151
R10386 GND.n5768 GND.n3193 10.6151
R10387 GND.n5768 GND.n5767 10.6151
R10388 GND.n5767 GND.n5766 10.6151
R10389 GND.n5766 GND.n3196 10.6151
R10390 GND.n5761 GND.n3196 10.6151
R10391 GND.n5761 GND.n5760 10.6151
R10392 GND.n5760 GND.n5759 10.6151
R10393 GND.n5759 GND.n3199 10.6151
R10394 GND.n5754 GND.n3199 10.6151
R10395 GND.n5754 GND.n5753 10.6151
R10396 GND.n5753 GND.n5752 10.6151
R10397 GND.n5752 GND.n3202 10.6151
R10398 GND.n5747 GND.n3202 10.6151
R10399 GND.n5747 GND.n5746 10.6151
R10400 GND.n5746 GND.n5745 10.6151
R10401 GND.n5745 GND.n3205 10.6151
R10402 GND.n5740 GND.n3205 10.6151
R10403 GND.n5740 GND.n5739 10.6151
R10404 GND.n5739 GND.n5738 10.6151
R10405 GND.n5738 GND.n3208 10.6151
R10406 GND.n5733 GND.n3208 10.6151
R10407 GND.n5733 GND.n5732 10.6151
R10408 GND.n5732 GND.n5731 10.6151
R10409 GND.n4111 GND.n4110 10.6151
R10410 GND.n4114 GND.n4111 10.6151
R10411 GND.n4115 GND.n4114 10.6151
R10412 GND.n4116 GND.n4115 10.6151
R10413 GND.n4116 GND.n3921 10.6151
R10414 GND.n4124 GND.n3921 10.6151
R10415 GND.n4125 GND.n4124 10.6151
R10416 GND.n4127 GND.n4125 10.6151
R10417 GND.n4128 GND.n4127 10.6151
R10418 GND.n4129 GND.n4128 10.6151
R10419 GND.n4129 GND.n3920 10.6151
R10420 GND.n4137 GND.n3920 10.6151
R10421 GND.n4138 GND.n4137 10.6151
R10422 GND.n4141 GND.n4138 10.6151
R10423 GND.n4142 GND.n4141 10.6151
R10424 GND.n4143 GND.n4142 10.6151
R10425 GND.n4143 GND.n3919 10.6151
R10426 GND.n4151 GND.n3919 10.6151
R10427 GND.n4152 GND.n4151 10.6151
R10428 GND.n4154 GND.n4152 10.6151
R10429 GND.n4155 GND.n4154 10.6151
R10430 GND.n4156 GND.n4155 10.6151
R10431 GND.n4156 GND.n3918 10.6151
R10432 GND.n4164 GND.n3918 10.6151
R10433 GND.n4165 GND.n4164 10.6151
R10434 GND.n4167 GND.n4165 10.6151
R10435 GND.n4168 GND.n4167 10.6151
R10436 GND.n4169 GND.n4168 10.6151
R10437 GND.n4169 GND.n3917 10.6151
R10438 GND.n4177 GND.n3917 10.6151
R10439 GND.n4178 GND.n4177 10.6151
R10440 GND.n4180 GND.n4178 10.6151
R10441 GND.n4181 GND.n4180 10.6151
R10442 GND.n4182 GND.n4181 10.6151
R10443 GND.n4182 GND.n3916 10.6151
R10444 GND.n4190 GND.n3916 10.6151
R10445 GND.n4191 GND.n4190 10.6151
R10446 GND.n4194 GND.n4191 10.6151
R10447 GND.n4195 GND.n4194 10.6151
R10448 GND.n4196 GND.n4195 10.6151
R10449 GND.n4204 GND.n4196 10.6151
R10450 GND.n4204 GND.n4203 10.6151
R10451 GND.n4203 GND.n4202 10.6151
R10452 GND.n4202 GND.n4200 10.6151
R10453 GND.n4200 GND.n4199 10.6151
R10454 GND.n4199 GND.n4197 10.6151
R10455 GND.n4197 GND.n3883 10.6151
R10456 GND.n4360 GND.n3883 10.6151
R10457 GND.n4361 GND.n4360 10.6151
R10458 GND.n4376 GND.n4361 10.6151
R10459 GND.n4376 GND.n4375 10.6151
R10460 GND.n4375 GND.n4374 10.6151
R10461 GND.n4374 GND.n4371 10.6151
R10462 GND.n4371 GND.n4370 10.6151
R10463 GND.n4370 GND.n4368 10.6151
R10464 GND.n4368 GND.n4367 10.6151
R10465 GND.n4367 GND.n4362 10.6151
R10466 GND.n4362 GND.n3844 10.6151
R10467 GND.n4445 GND.n3844 10.6151
R10468 GND.n4446 GND.n4445 10.6151
R10469 GND.n4466 GND.n4446 10.6151
R10470 GND.n4466 GND.n4465 10.6151
R10471 GND.n4465 GND.n4464 10.6151
R10472 GND.n4464 GND.n4463 10.6151
R10473 GND.n4463 GND.n4459 10.6151
R10474 GND.n4459 GND.n4458 10.6151
R10475 GND.n4458 GND.n4456 10.6151
R10476 GND.n4456 GND.n4455 10.6151
R10477 GND.n4455 GND.n4450 10.6151
R10478 GND.n4450 GND.n4449 10.6151
R10479 GND.n4449 GND.n4447 10.6151
R10480 GND.n4447 GND.n3795 10.6151
R10481 GND.n4533 GND.n3795 10.6151
R10482 GND.n4534 GND.n4533 10.6151
R10483 GND.n4565 GND.n4534 10.6151
R10484 GND.n4565 GND.n4564 10.6151
R10485 GND.n4564 GND.n4563 10.6151
R10486 GND.n4563 GND.n4535 10.6151
R10487 GND.n4557 GND.n4535 10.6151
R10488 GND.n4557 GND.n4556 10.6151
R10489 GND.n4556 GND.n4555 10.6151
R10490 GND.n4555 GND.n4554 10.6151
R10491 GND.n4554 GND.n4553 10.6151
R10492 GND.n4553 GND.n4550 10.6151
R10493 GND.n4550 GND.n4549 10.6151
R10494 GND.n4549 GND.n4547 10.6151
R10495 GND.n4547 GND.n4546 10.6151
R10496 GND.n4546 GND.n4543 10.6151
R10497 GND.n4543 GND.n4542 10.6151
R10498 GND.n4542 GND.n4540 10.6151
R10499 GND.n4540 GND.n4539 10.6151
R10500 GND.n4539 GND.n4536 10.6151
R10501 GND.n4536 GND.n3715 10.6151
R10502 GND.n4697 GND.n3715 10.6151
R10503 GND.n4698 GND.n4697 10.6151
R10504 GND.n4701 GND.n4698 10.6151
R10505 GND.n4701 GND.n4700 10.6151
R10506 GND.n4700 GND.n4699 10.6151
R10507 GND.n4699 GND.n3697 10.6151
R10508 GND.n4727 GND.n3697 10.6151
R10509 GND.n4728 GND.n4727 10.6151
R10510 GND.n4729 GND.n4728 10.6151
R10511 GND.n4729 GND.n3682 10.6151
R10512 GND.n4751 GND.n3682 10.6151
R10513 GND.n4752 GND.n4751 10.6151
R10514 GND.n4772 GND.n4752 10.6151
R10515 GND.n4772 GND.n4771 10.6151
R10516 GND.n4771 GND.n4770 10.6151
R10517 GND.n4770 GND.n4767 10.6151
R10518 GND.n4767 GND.n4766 10.6151
R10519 GND.n4766 GND.n4764 10.6151
R10520 GND.n4764 GND.n4763 10.6151
R10521 GND.n4763 GND.n4760 10.6151
R10522 GND.n4760 GND.n4759 10.6151
R10523 GND.n4759 GND.n4757 10.6151
R10524 GND.n4757 GND.n4756 10.6151
R10525 GND.n4756 GND.n4753 10.6151
R10526 GND.n4753 GND.n3628 10.6151
R10527 GND.n4874 GND.n3628 10.6151
R10528 GND.n4875 GND.n4874 10.6151
R10529 GND.n4878 GND.n4875 10.6151
R10530 GND.n4878 GND.n4877 10.6151
R10531 GND.n4877 GND.n4876 10.6151
R10532 GND.n4876 GND.n3610 10.6151
R10533 GND.n4904 GND.n3610 10.6151
R10534 GND.n4905 GND.n4904 10.6151
R10535 GND.n4906 GND.n4905 10.6151
R10536 GND.n4906 GND.n3595 10.6151
R10537 GND.n4928 GND.n3595 10.6151
R10538 GND.n4929 GND.n4928 10.6151
R10539 GND.n4949 GND.n4929 10.6151
R10540 GND.n4949 GND.n4948 10.6151
R10541 GND.n4948 GND.n4947 10.6151
R10542 GND.n4947 GND.n4944 10.6151
R10543 GND.n4944 GND.n4943 10.6151
R10544 GND.n4943 GND.n4941 10.6151
R10545 GND.n4941 GND.n4940 10.6151
R10546 GND.n4940 GND.n4937 10.6151
R10547 GND.n4937 GND.n4936 10.6151
R10548 GND.n4936 GND.n4934 10.6151
R10549 GND.n4934 GND.n4933 10.6151
R10550 GND.n4933 GND.n4930 10.6151
R10551 GND.n4930 GND.n3539 10.6151
R10552 GND.n5050 GND.n3539 10.6151
R10553 GND.n5051 GND.n5050 10.6151
R10554 GND.n5054 GND.n5051 10.6151
R10555 GND.n5054 GND.n5053 10.6151
R10556 GND.n5053 GND.n5052 10.6151
R10557 GND.n5052 GND.n3521 10.6151
R10558 GND.n5079 GND.n3521 10.6151
R10559 GND.n5080 GND.n5079 10.6151
R10560 GND.n5081 GND.n5080 10.6151
R10561 GND.n5081 GND.n3506 10.6151
R10562 GND.n5103 GND.n3506 10.6151
R10563 GND.n5104 GND.n5103 10.6151
R10564 GND.n5125 GND.n5104 10.6151
R10565 GND.n5125 GND.n5124 10.6151
R10566 GND.n5124 GND.n5123 10.6151
R10567 GND.n5123 GND.n5120 10.6151
R10568 GND.n5120 GND.n5119 10.6151
R10569 GND.n5119 GND.n5117 10.6151
R10570 GND.n5117 GND.n5116 10.6151
R10571 GND.n5116 GND.n5112 10.6151
R10572 GND.n5112 GND.n5111 10.6151
R10573 GND.n5111 GND.n5109 10.6151
R10574 GND.n5109 GND.n5108 10.6151
R10575 GND.n5108 GND.n5105 10.6151
R10576 GND.n5105 GND.n3450 10.6151
R10577 GND.n5225 GND.n3450 10.6151
R10578 GND.n5226 GND.n5225 10.6151
R10579 GND.n5229 GND.n5226 10.6151
R10580 GND.n5229 GND.n5228 10.6151
R10581 GND.n5228 GND.n5227 10.6151
R10582 GND.n5227 GND.n3431 10.6151
R10583 GND.n5254 GND.n3431 10.6151
R10584 GND.n5255 GND.n5254 10.6151
R10585 GND.n5256 GND.n5255 10.6151
R10586 GND.n5256 GND.n3417 10.6151
R10587 GND.n5278 GND.n3417 10.6151
R10588 GND.n5279 GND.n5278 10.6151
R10589 GND.n5299 GND.n5279 10.6151
R10590 GND.n5299 GND.n5298 10.6151
R10591 GND.n5298 GND.n5297 10.6151
R10592 GND.n5297 GND.n5294 10.6151
R10593 GND.n5294 GND.n5293 10.6151
R10594 GND.n5293 GND.n5291 10.6151
R10595 GND.n5291 GND.n5290 10.6151
R10596 GND.n5290 GND.n5287 10.6151
R10597 GND.n5287 GND.n5286 10.6151
R10598 GND.n5286 GND.n5284 10.6151
R10599 GND.n5284 GND.n5283 10.6151
R10600 GND.n5283 GND.n5280 10.6151
R10601 GND.n5280 GND.n3363 10.6151
R10602 GND.n5402 GND.n3363 10.6151
R10603 GND.n5403 GND.n5402 10.6151
R10604 GND.n5406 GND.n5403 10.6151
R10605 GND.n5406 GND.n5405 10.6151
R10606 GND.n5405 GND.n5404 10.6151
R10607 GND.n5404 GND.n3345 10.6151
R10608 GND.n5432 GND.n3345 10.6151
R10609 GND.n5433 GND.n5432 10.6151
R10610 GND.n5434 GND.n5433 10.6151
R10611 GND.n5434 GND.n3330 10.6151
R10612 GND.n5456 GND.n3330 10.6151
R10613 GND.n5457 GND.n5456 10.6151
R10614 GND.n5477 GND.n5457 10.6151
R10615 GND.n5477 GND.n5476 10.6151
R10616 GND.n5476 GND.n5475 10.6151
R10617 GND.n5475 GND.n5472 10.6151
R10618 GND.n5472 GND.n5471 10.6151
R10619 GND.n5471 GND.n5469 10.6151
R10620 GND.n5469 GND.n5468 10.6151
R10621 GND.n5468 GND.n5465 10.6151
R10622 GND.n5465 GND.n5464 10.6151
R10623 GND.n5464 GND.n5462 10.6151
R10624 GND.n5462 GND.n5461 10.6151
R10625 GND.n5461 GND.n5458 10.6151
R10626 GND.n5458 GND.n3276 10.6151
R10627 GND.n5558 GND.n3276 10.6151
R10628 GND.n5559 GND.n5558 10.6151
R10629 GND.n5560 GND.n5559 10.6151
R10630 GND.n5560 GND.n3265 10.6151
R10631 GND.n5591 GND.n3265 10.6151
R10632 GND.n5591 GND.n5590 10.6151
R10633 GND.n5590 GND.n5589 10.6151
R10634 GND.n5589 GND.n3266 10.6151
R10635 GND.n3266 GND.n3242 10.6151
R10636 GND.n5623 GND.n3242 10.6151
R10637 GND.n5624 GND.n5623 10.6151
R10638 GND.n5627 GND.n5624 10.6151
R10639 GND.n5627 GND.n5626 10.6151
R10640 GND.n5626 GND.n5625 10.6151
R10641 GND.n5625 GND.n3217 10.6151
R10642 GND.n5640 GND.n3217 10.6151
R10643 GND.n5641 GND.n5640 10.6151
R10644 GND.n5644 GND.n5641 10.6151
R10645 GND.n5645 GND.n5644 10.6151
R10646 GND.n5646 GND.n5645 10.6151
R10647 GND.n5646 GND.n3216 10.6151
R10648 GND.n5654 GND.n3216 10.6151
R10649 GND.n5655 GND.n5654 10.6151
R10650 GND.n5657 GND.n5655 10.6151
R10651 GND.n5658 GND.n5657 10.6151
R10652 GND.n5659 GND.n5658 10.6151
R10653 GND.n5659 GND.n3215 10.6151
R10654 GND.n5667 GND.n3215 10.6151
R10655 GND.n5668 GND.n5667 10.6151
R10656 GND.n5670 GND.n5668 10.6151
R10657 GND.n5671 GND.n5670 10.6151
R10658 GND.n5672 GND.n5671 10.6151
R10659 GND.n5672 GND.n3214 10.6151
R10660 GND.n5680 GND.n3214 10.6151
R10661 GND.n5681 GND.n5680 10.6151
R10662 GND.n5683 GND.n5681 10.6151
R10663 GND.n5684 GND.n5683 10.6151
R10664 GND.n5685 GND.n5684 10.6151
R10665 GND.n5685 GND.n3213 10.6151
R10666 GND.n5693 GND.n3213 10.6151
R10667 GND.n5694 GND.n5693 10.6151
R10668 GND.n5697 GND.n5694 10.6151
R10669 GND.n5698 GND.n5697 10.6151
R10670 GND.n5699 GND.n5698 10.6151
R10671 GND.n5699 GND.n3212 10.6151
R10672 GND.n5707 GND.n3212 10.6151
R10673 GND.n5708 GND.n5707 10.6151
R10674 GND.n5710 GND.n5708 10.6151
R10675 GND.n5711 GND.n5710 10.6151
R10676 GND.n5712 GND.n5711 10.6151
R10677 GND.n5712 GND.n3211 10.6151
R10678 GND.n5720 GND.n3211 10.6151
R10679 GND.n5721 GND.n5720 10.6151
R10680 GND.n5723 GND.n5721 10.6151
R10681 GND.n5724 GND.n5723 10.6151
R10682 GND.n5725 GND.n5724 10.6151
R10683 GND.n4047 GND.n4046 10.6151
R10684 GND.n4048 GND.n4047 10.6151
R10685 GND.n4048 GND.n3940 10.6151
R10686 GND.n4055 GND.n4054 10.6151
R10687 GND.n4056 GND.n4055 10.6151
R10688 GND.n4056 GND.n3935 10.6151
R10689 GND.n4062 GND.n3935 10.6151
R10690 GND.n4063 GND.n4062 10.6151
R10691 GND.n4064 GND.n4063 10.6151
R10692 GND.n4064 GND.n3933 10.6151
R10693 GND.n4070 GND.n3933 10.6151
R10694 GND.n4071 GND.n4070 10.6151
R10695 GND.n4072 GND.n4071 10.6151
R10696 GND.n4072 GND.n3931 10.6151
R10697 GND.n4078 GND.n3931 10.6151
R10698 GND.n4079 GND.n4078 10.6151
R10699 GND.n4080 GND.n4079 10.6151
R10700 GND.n4080 GND.n3929 10.6151
R10701 GND.n4086 GND.n3929 10.6151
R10702 GND.n4087 GND.n4086 10.6151
R10703 GND.n4088 GND.n4087 10.6151
R10704 GND.n4088 GND.n3927 10.6151
R10705 GND.n4094 GND.n3927 10.6151
R10706 GND.n4095 GND.n4094 10.6151
R10707 GND.n4096 GND.n4095 10.6151
R10708 GND.n4096 GND.n3925 10.6151
R10709 GND.n4102 GND.n3925 10.6151
R10710 GND.n4103 GND.n4102 10.6151
R10711 GND.n4104 GND.n4103 10.6151
R10712 GND.n4104 GND.n3923 10.6151
R10713 GND.n3923 GND.n3922 10.6151
R10714 GND.n3979 GND.n3975 10.6151
R10715 GND.n3980 GND.n3979 10.6151
R10716 GND.n3981 GND.n3980 10.6151
R10717 GND.n3981 GND.n3959 10.6151
R10718 GND.n3987 GND.n3959 10.6151
R10719 GND.n3988 GND.n3987 10.6151
R10720 GND.n3989 GND.n3988 10.6151
R10721 GND.n3989 GND.n3957 10.6151
R10722 GND.n3995 GND.n3957 10.6151
R10723 GND.n3996 GND.n3995 10.6151
R10724 GND.n3997 GND.n3996 10.6151
R10725 GND.n3997 GND.n3955 10.6151
R10726 GND.n4003 GND.n3955 10.6151
R10727 GND.n4004 GND.n4003 10.6151
R10728 GND.n4005 GND.n4004 10.6151
R10729 GND.n4005 GND.n3953 10.6151
R10730 GND.n4011 GND.n3953 10.6151
R10731 GND.n4012 GND.n4011 10.6151
R10732 GND.n4013 GND.n4012 10.6151
R10733 GND.n4013 GND.n3951 10.6151
R10734 GND.n4019 GND.n3951 10.6151
R10735 GND.n4020 GND.n4019 10.6151
R10736 GND.n4021 GND.n4020 10.6151
R10737 GND.n4021 GND.n3949 10.6151
R10738 GND.n4027 GND.n3949 10.6151
R10739 GND.n4028 GND.n4027 10.6151
R10740 GND.n4029 GND.n4028 10.6151
R10741 GND.n4029 GND.n3947 10.6151
R10742 GND.n4036 GND.n4035 10.6151
R10743 GND.n4037 GND.n4036 10.6151
R10744 GND.n4037 GND.n3942 10.6151
R10745 GND.n3117 GND.n3103 10.6151
R10746 GND.n3123 GND.n3103 10.6151
R10747 GND.n3124 GND.n3123 10.6151
R10748 GND.n3125 GND.n3124 10.6151
R10749 GND.n3125 GND.n3101 10.6151
R10750 GND.n3131 GND.n3101 10.6151
R10751 GND.n3132 GND.n3131 10.6151
R10752 GND.n3133 GND.n3132 10.6151
R10753 GND.n3133 GND.n3099 10.6151
R10754 GND.n3139 GND.n3099 10.6151
R10755 GND.n3140 GND.n3139 10.6151
R10756 GND.n3141 GND.n3140 10.6151
R10757 GND.n3141 GND.n3097 10.6151
R10758 GND.n3147 GND.n3097 10.6151
R10759 GND.n3148 GND.n3147 10.6151
R10760 GND.n3149 GND.n3148 10.6151
R10761 GND.n3149 GND.n3095 10.6151
R10762 GND.n3155 GND.n3095 10.6151
R10763 GND.n3156 GND.n3155 10.6151
R10764 GND.n3157 GND.n3156 10.6151
R10765 GND.n3157 GND.n3093 10.6151
R10766 GND.n3163 GND.n3093 10.6151
R10767 GND.n3164 GND.n3163 10.6151
R10768 GND.n3165 GND.n3164 10.6151
R10769 GND.n3165 GND.n3091 10.6151
R10770 GND.n3171 GND.n3091 10.6151
R10771 GND.n3172 GND.n3171 10.6151
R10772 GND.n3176 GND.n3172 10.6151
R10773 GND.n3181 GND.n3089 10.6151
R10774 GND.n3182 GND.n3181 10.6151
R10775 GND.n3182 GND.n3087 10.6151
R10776 GND.n6955 GND.n2543 10.6151
R10777 GND.n6955 GND.n6954 10.6151
R10778 GND.n6954 GND.n6953 10.6151
R10779 GND.n6953 GND.n2544 10.6151
R10780 GND.n4119 GND.n2544 10.6151
R10781 GND.n4119 GND.n2561 10.6151
R10782 GND.n6942 GND.n2561 10.6151
R10783 GND.n6942 GND.n6941 10.6151
R10784 GND.n6941 GND.n6940 10.6151
R10785 GND.n6940 GND.n2562 10.6151
R10786 GND.n4132 GND.n2562 10.6151
R10787 GND.n4132 GND.n2578 10.6151
R10788 GND.n6928 GND.n2578 10.6151
R10789 GND.n6928 GND.n6927 10.6151
R10790 GND.n6927 GND.n6926 10.6151
R10791 GND.n6926 GND.n2579 10.6151
R10792 GND.n4146 GND.n2579 10.6151
R10793 GND.n4146 GND.n2596 10.6151
R10794 GND.n6914 GND.n2596 10.6151
R10795 GND.n6914 GND.n6913 10.6151
R10796 GND.n6913 GND.n6912 10.6151
R10797 GND.n6912 GND.n2597 10.6151
R10798 GND.n4159 GND.n2597 10.6151
R10799 GND.n4159 GND.n2614 10.6151
R10800 GND.n6900 GND.n2614 10.6151
R10801 GND.n6900 GND.n6899 10.6151
R10802 GND.n6899 GND.n6898 10.6151
R10803 GND.n6898 GND.n2615 10.6151
R10804 GND.n4172 GND.n2615 10.6151
R10805 GND.n4172 GND.n2632 10.6151
R10806 GND.n6886 GND.n2632 10.6151
R10807 GND.n6886 GND.n6885 10.6151
R10808 GND.n6885 GND.n6884 10.6151
R10809 GND.n6884 GND.n2633 10.6151
R10810 GND.n4185 GND.n2633 10.6151
R10811 GND.n4185 GND.n2650 10.6151
R10812 GND.n6872 GND.n2650 10.6151
R10813 GND.n6872 GND.n6871 10.6151
R10814 GND.n6871 GND.n6870 10.6151
R10815 GND.n6870 GND.n2651 10.6151
R10816 GND.n4208 GND.n2651 10.6151
R10817 GND.n4208 GND.n4207 10.6151
R10818 GND.n4207 GND.n3896 10.6151
R10819 GND.n4342 GND.n3896 10.6151
R10820 GND.n4343 GND.n4342 10.6151
R10821 GND.n4345 GND.n4343 10.6151
R10822 GND.n4345 GND.n4344 10.6151
R10823 GND.n4344 GND.n3879 10.6151
R10824 GND.n4382 GND.n3879 10.6151
R10825 GND.n4383 GND.n4382 10.6151
R10826 GND.n4384 GND.n4383 10.6151
R10827 GND.n4384 GND.n3864 10.6151
R10828 GND.n4412 GND.n3864 10.6151
R10829 GND.n4413 GND.n4412 10.6151
R10830 GND.n4414 GND.n4413 10.6151
R10831 GND.n4414 GND.n3849 10.6151
R10832 GND.n4439 GND.n3849 10.6151
R10833 GND.n4440 GND.n4439 10.6151
R10834 GND.n4441 GND.n4440 10.6151
R10835 GND.n4441 GND.n3839 10.6151
R10836 GND.n4471 GND.n3839 10.6151
R10837 GND.n4472 GND.n4471 10.6151
R10838 GND.n4473 GND.n4472 10.6151
R10839 GND.n4473 GND.n3824 10.6151
R10840 GND.n4489 GND.n3824 10.6151
R10841 GND.n4490 GND.n4489 10.6151
R10842 GND.n4491 GND.n4490 10.6151
R10843 GND.n4491 GND.n3810 10.6151
R10844 GND.n4515 GND.n3810 10.6151
R10845 GND.n4516 GND.n4515 10.6151
R10846 GND.n4518 GND.n4516 10.6151
R10847 GND.n4518 GND.n4517 10.6151
R10848 GND.n4517 GND.n3790 10.6151
R10849 GND.n4571 GND.n3790 10.6151
R10850 GND.n4572 GND.n4571 10.6151
R10851 GND.n4576 GND.n4572 10.6151
R10852 GND.n4576 GND.n4575 10.6151
R10853 GND.n4575 GND.n4574 10.6151
R10854 GND.n4574 GND.n3765 10.6151
R10855 GND.n4602 GND.n3765 10.6151
R10856 GND.n4603 GND.n4602 10.6151
R10857 GND.n4604 GND.n4603 10.6151
R10858 GND.n4604 GND.n3752 10.6151
R10859 GND.n4621 GND.n3752 10.6151
R10860 GND.n4622 GND.n4621 10.6151
R10861 GND.n4623 GND.n4622 10.6151
R10862 GND.n4623 GND.n3738 10.6151
R10863 GND.n4673 GND.n3738 10.6151
R10864 GND.n4674 GND.n4673 10.6151
R10865 GND.n4675 GND.n4674 10.6151
R10866 GND.n4675 GND.n3721 10.6151
R10867 GND.n4690 GND.n3721 10.6151
R10868 GND.n4691 GND.n4690 10.6151
R10869 GND.n4693 GND.n4691 10.6151
R10870 GND.n4693 GND.n4692 10.6151
R10871 GND.n4692 GND.n3701 10.6151
R10872 GND.n4719 GND.n3701 10.6151
R10873 GND.n4720 GND.n4719 10.6151
R10874 GND.n4721 GND.n4720 10.6151
R10875 GND.n4721 GND.n3696 10.6151
R10876 GND.n4737 GND.n3696 10.6151
R10877 GND.n4737 GND.n4736 10.6151
R10878 GND.n4736 GND.n4735 10.6151
R10879 GND.n4735 GND.n3678 10.6151
R10880 GND.n4778 GND.n3678 10.6151
R10881 GND.n4779 GND.n4778 10.6151
R10882 GND.n4780 GND.n4779 10.6151
R10883 GND.n4780 GND.n3664 10.6151
R10884 GND.n4798 GND.n3664 10.6151
R10885 GND.n4799 GND.n4798 10.6151
R10886 GND.n4800 GND.n4799 10.6151
R10887 GND.n4800 GND.n3650 10.6151
R10888 GND.n4849 GND.n3650 10.6151
R10889 GND.n4850 GND.n4849 10.6151
R10890 GND.n4851 GND.n4850 10.6151
R10891 GND.n4851 GND.n3634 10.6151
R10892 GND.n4867 GND.n3634 10.6151
R10893 GND.n4868 GND.n4867 10.6151
R10894 GND.n4870 GND.n4868 10.6151
R10895 GND.n4870 GND.n4869 10.6151
R10896 GND.n4869 GND.n3614 10.6151
R10897 GND.n4896 GND.n3614 10.6151
R10898 GND.n4897 GND.n4896 10.6151
R10899 GND.n4898 GND.n4897 10.6151
R10900 GND.n4898 GND.n3609 10.6151
R10901 GND.n4914 GND.n3609 10.6151
R10902 GND.n4914 GND.n4913 10.6151
R10903 GND.n4913 GND.n4912 10.6151
R10904 GND.n4912 GND.n3591 10.6151
R10905 GND.n4955 GND.n3591 10.6151
R10906 GND.n4956 GND.n4955 10.6151
R10907 GND.n4957 GND.n4956 10.6151
R10908 GND.n4957 GND.n3576 10.6151
R10909 GND.n4974 GND.n3576 10.6151
R10910 GND.n4975 GND.n4974 10.6151
R10911 GND.n4976 GND.n4975 10.6151
R10912 GND.n4976 GND.n3562 10.6151
R10913 GND.n5026 GND.n3562 10.6151
R10914 GND.n5027 GND.n5026 10.6151
R10915 GND.n5028 GND.n5027 10.6151
R10916 GND.n5028 GND.n3546 10.6151
R10917 GND.n5043 GND.n3546 10.6151
R10918 GND.n5044 GND.n5043 10.6151
R10919 GND.n5046 GND.n5044 10.6151
R10920 GND.n5046 GND.n5045 10.6151
R10921 GND.n5045 GND.n3525 10.6151
R10922 GND.n5071 GND.n3525 10.6151
R10923 GND.n5072 GND.n5071 10.6151
R10924 GND.n5073 GND.n5072 10.6151
R10925 GND.n5073 GND.n3520 10.6151
R10926 GND.n5089 GND.n3520 10.6151
R10927 GND.n5089 GND.n5088 10.6151
R10928 GND.n5088 GND.n5087 10.6151
R10929 GND.n5087 GND.n3502 10.6151
R10930 GND.n5131 GND.n3502 10.6151
R10931 GND.n5132 GND.n5131 10.6151
R10932 GND.n5133 GND.n5132 10.6151
R10933 GND.n5133 GND.n3487 10.6151
R10934 GND.n5150 GND.n3487 10.6151
R10935 GND.n5151 GND.n5150 10.6151
R10936 GND.n5152 GND.n5151 10.6151
R10937 GND.n5152 GND.n3473 10.6151
R10938 GND.n5201 GND.n3473 10.6151
R10939 GND.n5202 GND.n5201 10.6151
R10940 GND.n5203 GND.n5202 10.6151
R10941 GND.n5203 GND.n3456 10.6151
R10942 GND.n5218 GND.n3456 10.6151
R10943 GND.n5219 GND.n5218 10.6151
R10944 GND.n5221 GND.n5219 10.6151
R10945 GND.n5221 GND.n5220 10.6151
R10946 GND.n5220 GND.n3436 10.6151
R10947 GND.n5246 GND.n3436 10.6151
R10948 GND.n5247 GND.n5246 10.6151
R10949 GND.n5248 GND.n5247 10.6151
R10950 GND.n5248 GND.n3429 10.6151
R10951 GND.n5264 GND.n3429 10.6151
R10952 GND.n5264 GND.n5263 10.6151
R10953 GND.n5263 GND.n5262 10.6151
R10954 GND.n5262 GND.n3412 10.6151
R10955 GND.n5305 GND.n3412 10.6151
R10956 GND.n5306 GND.n5305 10.6151
R10957 GND.n5307 GND.n5306 10.6151
R10958 GND.n5307 GND.n3398 10.6151
R10959 GND.n5324 GND.n3398 10.6151
R10960 GND.n5325 GND.n5324 10.6151
R10961 GND.n5326 GND.n5325 10.6151
R10962 GND.n5326 GND.n3384 10.6151
R10963 GND.n5378 GND.n3384 10.6151
R10964 GND.n5379 GND.n5378 10.6151
R10965 GND.n5380 GND.n5379 10.6151
R10966 GND.n5380 GND.n3369 10.6151
R10967 GND.n5395 GND.n3369 10.6151
R10968 GND.n5396 GND.n5395 10.6151
R10969 GND.n5398 GND.n5396 10.6151
R10970 GND.n5398 GND.n5397 10.6151
R10971 GND.n5397 GND.n3349 10.6151
R10972 GND.n5424 GND.n3349 10.6151
R10973 GND.n5425 GND.n5424 10.6151
R10974 GND.n5426 GND.n5425 10.6151
R10975 GND.n5426 GND.n3344 10.6151
R10976 GND.n5442 GND.n3344 10.6151
R10977 GND.n5442 GND.n5441 10.6151
R10978 GND.n5441 GND.n5440 10.6151
R10979 GND.n5440 GND.n3326 10.6151
R10980 GND.n5483 GND.n3326 10.6151
R10981 GND.n5484 GND.n5483 10.6151
R10982 GND.n5485 GND.n5484 10.6151
R10983 GND.n5485 GND.n3312 10.6151
R10984 GND.n5503 GND.n3312 10.6151
R10985 GND.n5504 GND.n5503 10.6151
R10986 GND.n5505 GND.n5504 10.6151
R10987 GND.n5505 GND.n3298 10.6151
R10988 GND.n5531 GND.n3298 10.6151
R10989 GND.n5532 GND.n5531 10.6151
R10990 GND.n5533 GND.n5532 10.6151
R10991 GND.n5533 GND.n3282 10.6151
R10992 GND.n5551 GND.n3282 10.6151
R10993 GND.n5552 GND.n5551 10.6151
R10994 GND.n5554 GND.n5552 10.6151
R10995 GND.n5554 GND.n5553 10.6151
R10996 GND.n5553 GND.n3261 10.6151
R10997 GND.n5597 GND.n3261 10.6151
R10998 GND.n5598 GND.n5597 10.6151
R10999 GND.n5599 GND.n5598 10.6151
R11000 GND.n5599 GND.n3247 10.6151
R11001 GND.n5616 GND.n3247 10.6151
R11002 GND.n5617 GND.n5616 10.6151
R11003 GND.n5619 GND.n5617 10.6151
R11004 GND.n5619 GND.n5618 10.6151
R11005 GND.n5618 GND.n3237 10.6151
R11006 GND.n5633 GND.n3237 10.6151
R11007 GND.n5634 GND.n5633 10.6151
R11008 GND.n5635 GND.n5634 10.6151
R11009 GND.n5635 GND.n2918 10.6151
R11010 GND.n6616 GND.n2918 10.6151
R11011 GND.n6616 GND.n6615 10.6151
R11012 GND.n6615 GND.n6614 10.6151
R11013 GND.n6614 GND.n2919 10.6151
R11014 GND.n5649 GND.n2919 10.6151
R11015 GND.n5649 GND.n2936 10.6151
R11016 GND.n6602 GND.n2936 10.6151
R11017 GND.n6602 GND.n6601 10.6151
R11018 GND.n6601 GND.n6600 10.6151
R11019 GND.n6600 GND.n2937 10.6151
R11020 GND.n5662 GND.n2937 10.6151
R11021 GND.n5662 GND.n2954 10.6151
R11022 GND.n6588 GND.n2954 10.6151
R11023 GND.n6588 GND.n6587 10.6151
R11024 GND.n6587 GND.n6586 10.6151
R11025 GND.n6586 GND.n2955 10.6151
R11026 GND.n5675 GND.n2955 10.6151
R11027 GND.n5675 GND.n2972 10.6151
R11028 GND.n6574 GND.n2972 10.6151
R11029 GND.n6574 GND.n6573 10.6151
R11030 GND.n6573 GND.n6572 10.6151
R11031 GND.n6572 GND.n2973 10.6151
R11032 GND.n5688 GND.n2973 10.6151
R11033 GND.n5688 GND.n2990 10.6151
R11034 GND.n6560 GND.n2990 10.6151
R11035 GND.n6560 GND.n6559 10.6151
R11036 GND.n6559 GND.n6558 10.6151
R11037 GND.n6558 GND.n2991 10.6151
R11038 GND.n5702 GND.n2991 10.6151
R11039 GND.n5702 GND.n3007 10.6151
R11040 GND.n6546 GND.n3007 10.6151
R11041 GND.n6546 GND.n6545 10.6151
R11042 GND.n6545 GND.n6544 10.6151
R11043 GND.n6544 GND.n3008 10.6151
R11044 GND.n5715 GND.n3008 10.6151
R11045 GND.n5715 GND.n3024 10.6151
R11046 GND.n6532 GND.n3024 10.6151
R11047 GND.n6532 GND.n6531 10.6151
R11048 GND.n6531 GND.n6530 10.6151
R11049 GND.n6530 GND.n3025 10.6151
R11050 GND.n2539 GND.t176 10.5917
R11051 GND.n4469 GND.n3841 10.5917
R11052 GND.n4475 GND.n3837 10.5917
R11053 GND.n4627 GND.n4625 10.5917
R11054 GND.n4671 GND.n4670 10.5917
R11055 GND.n4803 GND.n4802 10.5917
R11056 GND.n4979 GND.n4978 10.5917
R11057 GND.n5024 GND.n5023 10.5917
R11058 GND.n5199 GND.n5198 10.5917
R11059 GND.n5330 GND.n5328 10.5917
R11060 GND.n5376 GND.n5375 10.5917
R11061 GND.n5508 GND.n5507 10.5917
R11062 GND.n5529 GND.n5528 10.5917
R11063 GND.n1904 GND.n1903 10.4732
R11064 GND.n4297 GND.n4296 10.4732
R11065 GND.n2857 GND.n2856 10.4732
R11066 GND.n6090 GND.n6089 10.4732
R11067 GND.n1892 GND.n1891 10.2747
R11068 GND.n4285 GND.n4284 10.2747
R11069 GND.n2845 GND.n2844 10.2747
R11070 GND.n6078 GND.n6077 10.2747
R11071 GND.n19 GND.n18 10.1164
R11072 GND.n34 GND.n33 10.1164
R11073 GND.n50 GND.n49 10.1164
R11074 GND.n4 GND.n3 10.1164
R11075 GND.n80 GND.n79 10.1164
R11076 GND.n95 GND.n94 10.1164
R11077 GND.n111 GND.n110 10.1164
R11078 GND.n127 GND.n126 10.1164
R11079 GND.n2122 GND.t10 9.92979
R11080 GND.n2022 GND.t39 9.92979
R11081 GND.n4112 GND.n2546 9.92979
R11082 GND.n6909 GND.n2601 9.92979
R11083 GND.n6896 GND.n6895 9.92979
R11084 GND.n3894 GND.n3892 9.92979
R11085 GND.n4372 GND.n3866 9.92979
R11086 GND.n3808 GND.n3806 9.92979
R11087 GND.n4561 GND.n4560 9.92979
R11088 GND.n4717 GND.n3703 9.92979
R11089 GND.n4732 GND.n4731 9.92979
R11090 GND.n4894 GND.n3616 9.92979
R11091 GND.n4909 GND.n4908 9.92979
R11092 GND.n5069 GND.n3527 9.92979
R11093 GND.n5084 GND.n5083 9.92979
R11094 GND.n5244 GND.n3438 9.92979
R11095 GND.n5259 GND.n5258 9.92979
R11096 GND.n5422 GND.n3351 9.92979
R11097 GND.n5437 GND.n5436 9.92979
R11098 GND.n5595 GND.n3263 9.92979
R11099 GND.n5611 GND.n3244 9.92979
R11100 GND.n6591 GND.n6590 9.92979
R11101 GND.n6577 GND.n2967 9.92979
R11102 GND.n3028 GND.n3027 9.92979
R11103 GND.n6168 GND.t14 9.92979
R11104 GND.n8483 GND.t52 9.92979
R11105 GND.n1900 GND.n1886 9.69747
R11106 GND.n4293 GND.n4279 9.69747
R11107 GND.n2853 GND.n2839 9.69747
R11108 GND.n6086 GND.n6072 9.69747
R11109 GND.n25 GND.n24 9.45567
R11110 GND.n40 GND.n39 9.45567
R11111 GND.n56 GND.n55 9.45567
R11112 GND.n10 GND.n9 9.45567
R11113 GND.n1914 GND.n1913 9.45567
R11114 GND.n4307 GND.n4306 9.45567
R11115 GND.n2867 GND.n2866 9.45567
R11116 GND.n86 GND.n85 9.45567
R11117 GND.n101 GND.n100 9.45567
R11118 GND.n117 GND.n116 9.45567
R11119 GND.n133 GND.n132 9.45567
R11120 GND.n6100 GND.n6099 9.45567
R11121 GND.n5781 GND.n5780 9.36635
R11122 GND.n4054 GND.n3939 9.36635
R11123 GND.n3947 GND.n3946 9.36635
R11124 GND.n3176 GND.n3175 9.36635
R11125 GND.n1563 GND.n1562 9.35353
R11126 GND.n1857 GND.n1856 9.35353
R11127 GND.n24 GND.n23 9.3005
R11128 GND.n17 GND.n16 9.3005
R11129 GND.n39 GND.n38 9.3005
R11130 GND.n32 GND.n31 9.3005
R11131 GND.n55 GND.n54 9.3005
R11132 GND.n48 GND.n47 9.3005
R11133 GND.n9 GND.n8 9.3005
R11134 GND.n2 GND.n1 9.3005
R11135 GND.n1890 GND.n1889 9.3005
R11136 GND.n1897 GND.n1896 9.3005
R11137 GND.n1899 GND.n1898 9.3005
R11138 GND.n1886 GND.n1885 9.3005
R11139 GND.n1905 GND.n1904 9.3005
R11140 GND.n1907 GND.n1906 9.3005
R11141 GND.n1882 GND.n1881 9.3005
R11142 GND.n1913 GND.n1912 9.3005
R11143 GND.n4283 GND.n4282 9.3005
R11144 GND.n4290 GND.n4289 9.3005
R11145 GND.n4292 GND.n4291 9.3005
R11146 GND.n4279 GND.n4278 9.3005
R11147 GND.n4298 GND.n4297 9.3005
R11148 GND.n4300 GND.n4299 9.3005
R11149 GND.n4275 GND.n4274 9.3005
R11150 GND.n4306 GND.n4305 9.3005
R11151 GND.n2843 GND.n2842 9.3005
R11152 GND.n2850 GND.n2849 9.3005
R11153 GND.n2852 GND.n2851 9.3005
R11154 GND.n2839 GND.n2838 9.3005
R11155 GND.n2858 GND.n2857 9.3005
R11156 GND.n2860 GND.n2859 9.3005
R11157 GND.n2835 GND.n2834 9.3005
R11158 GND.n2866 GND.n2865 9.3005
R11159 GND.n2342 GND.n2341 9.3005
R11160 GND.n2343 GND.n2086 9.3005
R11161 GND.n2345 GND.n2344 9.3005
R11162 GND.n2037 GND.n2036 9.3005
R11163 GND.n2426 GND.n2425 9.3005
R11164 GND.n2427 GND.n2035 9.3005
R11165 GND.n2431 GND.n2428 9.3005
R11166 GND.n2430 GND.n2429 9.3005
R11167 GND.n2015 GND.n2014 9.3005
R11168 GND.n2452 GND.n2451 9.3005
R11169 GND.n2453 GND.n2013 9.3005
R11170 GND.n2461 GND.n2454 9.3005
R11171 GND.n2460 GND.n2455 9.3005
R11172 GND.n2459 GND.n2457 9.3005
R11173 GND.n2456 GND.n1982 9.3005
R11174 GND.n2495 GND.n1983 9.3005
R11175 GND.n2494 GND.n1984 9.3005
R11176 GND.n2493 GND.n1985 9.3005
R11177 GND.n1993 GND.n1986 9.3005
R11178 GND.n1992 GND.n1987 9.3005
R11179 GND.n1990 GND.n1988 9.3005
R11180 GND.n1989 GND.n1434 9.3005
R11181 GND.n7373 GND.n7372 9.3005
R11182 GND.n1033 GND.n1032 9.3005
R11183 GND.n7380 GND.n7379 9.3005
R11184 GND.n7381 GND.n1031 9.3005
R11185 GND.n7383 GND.n7382 9.3005
R11186 GND.n1027 GND.n1026 9.3005
R11187 GND.n7390 GND.n7389 9.3005
R11188 GND.n7391 GND.n1025 9.3005
R11189 GND.n7393 GND.n7392 9.3005
R11190 GND.n1021 GND.n1020 9.3005
R11191 GND.n7400 GND.n7399 9.3005
R11192 GND.n7401 GND.n1019 9.3005
R11193 GND.n7403 GND.n7402 9.3005
R11194 GND.n1015 GND.n1014 9.3005
R11195 GND.n7410 GND.n7409 9.3005
R11196 GND.n7411 GND.n1013 9.3005
R11197 GND.n7413 GND.n7412 9.3005
R11198 GND.n1009 GND.n1008 9.3005
R11199 GND.n7420 GND.n7419 9.3005
R11200 GND.n7421 GND.n1007 9.3005
R11201 GND.n7423 GND.n7422 9.3005
R11202 GND.n1003 GND.n1002 9.3005
R11203 GND.n7430 GND.n7429 9.3005
R11204 GND.n7431 GND.n1001 9.3005
R11205 GND.n7433 GND.n7432 9.3005
R11206 GND.n997 GND.n996 9.3005
R11207 GND.n7440 GND.n7439 9.3005
R11208 GND.n7441 GND.n995 9.3005
R11209 GND.n7443 GND.n7442 9.3005
R11210 GND.n991 GND.n990 9.3005
R11211 GND.n7450 GND.n7449 9.3005
R11212 GND.n7451 GND.n989 9.3005
R11213 GND.n7453 GND.n7452 9.3005
R11214 GND.n985 GND.n984 9.3005
R11215 GND.n7460 GND.n7459 9.3005
R11216 GND.n7461 GND.n983 9.3005
R11217 GND.n7463 GND.n7462 9.3005
R11218 GND.n979 GND.n978 9.3005
R11219 GND.n7470 GND.n7469 9.3005
R11220 GND.n7471 GND.n977 9.3005
R11221 GND.n7473 GND.n7472 9.3005
R11222 GND.n973 GND.n972 9.3005
R11223 GND.n7480 GND.n7479 9.3005
R11224 GND.n7481 GND.n971 9.3005
R11225 GND.n7483 GND.n7482 9.3005
R11226 GND.n967 GND.n966 9.3005
R11227 GND.n7490 GND.n7489 9.3005
R11228 GND.n7491 GND.n965 9.3005
R11229 GND.n7493 GND.n7492 9.3005
R11230 GND.n961 GND.n960 9.3005
R11231 GND.n7500 GND.n7499 9.3005
R11232 GND.n7501 GND.n959 9.3005
R11233 GND.n7503 GND.n7502 9.3005
R11234 GND.n955 GND.n954 9.3005
R11235 GND.n7510 GND.n7509 9.3005
R11236 GND.n7511 GND.n953 9.3005
R11237 GND.n7513 GND.n7512 9.3005
R11238 GND.n949 GND.n948 9.3005
R11239 GND.n7520 GND.n7519 9.3005
R11240 GND.n7521 GND.n947 9.3005
R11241 GND.n7523 GND.n7522 9.3005
R11242 GND.n943 GND.n942 9.3005
R11243 GND.n7530 GND.n7529 9.3005
R11244 GND.n7531 GND.n941 9.3005
R11245 GND.n7533 GND.n7532 9.3005
R11246 GND.n937 GND.n936 9.3005
R11247 GND.n7540 GND.n7539 9.3005
R11248 GND.n7541 GND.n935 9.3005
R11249 GND.n7543 GND.n7542 9.3005
R11250 GND.n931 GND.n930 9.3005
R11251 GND.n7550 GND.n7549 9.3005
R11252 GND.n7551 GND.n929 9.3005
R11253 GND.n7553 GND.n7552 9.3005
R11254 GND.n925 GND.n924 9.3005
R11255 GND.n7560 GND.n7559 9.3005
R11256 GND.n7561 GND.n923 9.3005
R11257 GND.n7563 GND.n7562 9.3005
R11258 GND.n919 GND.n918 9.3005
R11259 GND.n7570 GND.n7569 9.3005
R11260 GND.n7571 GND.n917 9.3005
R11261 GND.n7573 GND.n7572 9.3005
R11262 GND.n913 GND.n912 9.3005
R11263 GND.n7580 GND.n7579 9.3005
R11264 GND.n7581 GND.n911 9.3005
R11265 GND.n7583 GND.n7582 9.3005
R11266 GND.n907 GND.n906 9.3005
R11267 GND.n7590 GND.n7589 9.3005
R11268 GND.n7591 GND.n905 9.3005
R11269 GND.n7593 GND.n7592 9.3005
R11270 GND.n901 GND.n900 9.3005
R11271 GND.n7600 GND.n7599 9.3005
R11272 GND.n7601 GND.n899 9.3005
R11273 GND.n7603 GND.n7602 9.3005
R11274 GND.n895 GND.n894 9.3005
R11275 GND.n7610 GND.n7609 9.3005
R11276 GND.n7611 GND.n893 9.3005
R11277 GND.n7613 GND.n7612 9.3005
R11278 GND.n889 GND.n888 9.3005
R11279 GND.n7620 GND.n7619 9.3005
R11280 GND.n7621 GND.n887 9.3005
R11281 GND.n7623 GND.n7622 9.3005
R11282 GND.n883 GND.n882 9.3005
R11283 GND.n7630 GND.n7629 9.3005
R11284 GND.n7631 GND.n881 9.3005
R11285 GND.n7633 GND.n7632 9.3005
R11286 GND.n877 GND.n876 9.3005
R11287 GND.n7640 GND.n7639 9.3005
R11288 GND.n7641 GND.n875 9.3005
R11289 GND.n7643 GND.n7642 9.3005
R11290 GND.n871 GND.n870 9.3005
R11291 GND.n7650 GND.n7649 9.3005
R11292 GND.n7651 GND.n869 9.3005
R11293 GND.n7653 GND.n7652 9.3005
R11294 GND.n865 GND.n864 9.3005
R11295 GND.n7660 GND.n7659 9.3005
R11296 GND.n7661 GND.n863 9.3005
R11297 GND.n7663 GND.n7662 9.3005
R11298 GND.n859 GND.n858 9.3005
R11299 GND.n7670 GND.n7669 9.3005
R11300 GND.n7671 GND.n857 9.3005
R11301 GND.n7673 GND.n7672 9.3005
R11302 GND.n853 GND.n852 9.3005
R11303 GND.n7680 GND.n7679 9.3005
R11304 GND.n7681 GND.n851 9.3005
R11305 GND.n7683 GND.n7682 9.3005
R11306 GND.n847 GND.n846 9.3005
R11307 GND.n7690 GND.n7689 9.3005
R11308 GND.n7691 GND.n845 9.3005
R11309 GND.n7693 GND.n7692 9.3005
R11310 GND.n841 GND.n840 9.3005
R11311 GND.n7700 GND.n7699 9.3005
R11312 GND.n7701 GND.n839 9.3005
R11313 GND.n7703 GND.n7702 9.3005
R11314 GND.n835 GND.n834 9.3005
R11315 GND.n7710 GND.n7709 9.3005
R11316 GND.n7711 GND.n833 9.3005
R11317 GND.n7713 GND.n7712 9.3005
R11318 GND.n829 GND.n828 9.3005
R11319 GND.n7720 GND.n7719 9.3005
R11320 GND.n7721 GND.n827 9.3005
R11321 GND.n7723 GND.n7722 9.3005
R11322 GND.n823 GND.n822 9.3005
R11323 GND.n7730 GND.n7729 9.3005
R11324 GND.n7731 GND.n821 9.3005
R11325 GND.n7733 GND.n7732 9.3005
R11326 GND.n817 GND.n816 9.3005
R11327 GND.n7740 GND.n7739 9.3005
R11328 GND.n7741 GND.n815 9.3005
R11329 GND.n7743 GND.n7742 9.3005
R11330 GND.n811 GND.n810 9.3005
R11331 GND.n7750 GND.n7749 9.3005
R11332 GND.n7751 GND.n809 9.3005
R11333 GND.n7753 GND.n7752 9.3005
R11334 GND.n805 GND.n804 9.3005
R11335 GND.n7760 GND.n7759 9.3005
R11336 GND.n7761 GND.n803 9.3005
R11337 GND.n7763 GND.n7762 9.3005
R11338 GND.n799 GND.n798 9.3005
R11339 GND.n7770 GND.n7769 9.3005
R11340 GND.n7771 GND.n797 9.3005
R11341 GND.n7773 GND.n7772 9.3005
R11342 GND.n793 GND.n792 9.3005
R11343 GND.n7780 GND.n7779 9.3005
R11344 GND.n7781 GND.n791 9.3005
R11345 GND.n7783 GND.n7782 9.3005
R11346 GND.n787 GND.n786 9.3005
R11347 GND.n7790 GND.n7789 9.3005
R11348 GND.n7791 GND.n785 9.3005
R11349 GND.n7793 GND.n7792 9.3005
R11350 GND.n781 GND.n780 9.3005
R11351 GND.n7800 GND.n7799 9.3005
R11352 GND.n7801 GND.n779 9.3005
R11353 GND.n7803 GND.n7802 9.3005
R11354 GND.n775 GND.n774 9.3005
R11355 GND.n7810 GND.n7809 9.3005
R11356 GND.n7811 GND.n773 9.3005
R11357 GND.n7813 GND.n7812 9.3005
R11358 GND.n769 GND.n768 9.3005
R11359 GND.n7820 GND.n7819 9.3005
R11360 GND.n7821 GND.n767 9.3005
R11361 GND.n7823 GND.n7822 9.3005
R11362 GND.n763 GND.n762 9.3005
R11363 GND.n7830 GND.n7829 9.3005
R11364 GND.n7831 GND.n761 9.3005
R11365 GND.n7833 GND.n7832 9.3005
R11366 GND.n757 GND.n756 9.3005
R11367 GND.n7840 GND.n7839 9.3005
R11368 GND.n7841 GND.n755 9.3005
R11369 GND.n7843 GND.n7842 9.3005
R11370 GND.n751 GND.n750 9.3005
R11371 GND.n7850 GND.n7849 9.3005
R11372 GND.n7851 GND.n749 9.3005
R11373 GND.n7853 GND.n7852 9.3005
R11374 GND.n745 GND.n744 9.3005
R11375 GND.n7860 GND.n7859 9.3005
R11376 GND.n7861 GND.n743 9.3005
R11377 GND.n7863 GND.n7862 9.3005
R11378 GND.n739 GND.n738 9.3005
R11379 GND.n7870 GND.n7869 9.3005
R11380 GND.n7871 GND.n737 9.3005
R11381 GND.n7873 GND.n7872 9.3005
R11382 GND.n733 GND.n732 9.3005
R11383 GND.n7880 GND.n7879 9.3005
R11384 GND.n7881 GND.n731 9.3005
R11385 GND.n7883 GND.n7882 9.3005
R11386 GND.n727 GND.n726 9.3005
R11387 GND.n7890 GND.n7889 9.3005
R11388 GND.n7891 GND.n725 9.3005
R11389 GND.n7893 GND.n7892 9.3005
R11390 GND.n721 GND.n720 9.3005
R11391 GND.n7900 GND.n7899 9.3005
R11392 GND.n7901 GND.n719 9.3005
R11393 GND.n7903 GND.n7902 9.3005
R11394 GND.n715 GND.n714 9.3005
R11395 GND.n7910 GND.n7909 9.3005
R11396 GND.n7911 GND.n713 9.3005
R11397 GND.n7913 GND.n7912 9.3005
R11398 GND.n709 GND.n708 9.3005
R11399 GND.n7920 GND.n7919 9.3005
R11400 GND.n7921 GND.n707 9.3005
R11401 GND.n7923 GND.n7922 9.3005
R11402 GND.n703 GND.n702 9.3005
R11403 GND.n7930 GND.n7929 9.3005
R11404 GND.n7931 GND.n701 9.3005
R11405 GND.n7933 GND.n7932 9.3005
R11406 GND.n697 GND.n696 9.3005
R11407 GND.n7940 GND.n7939 9.3005
R11408 GND.n7941 GND.n695 9.3005
R11409 GND.n7943 GND.n7942 9.3005
R11410 GND.n691 GND.n690 9.3005
R11411 GND.n7950 GND.n7949 9.3005
R11412 GND.n7951 GND.n689 9.3005
R11413 GND.n7953 GND.n7952 9.3005
R11414 GND.n685 GND.n684 9.3005
R11415 GND.n7960 GND.n7959 9.3005
R11416 GND.n7961 GND.n683 9.3005
R11417 GND.n7963 GND.n7962 9.3005
R11418 GND.n679 GND.n678 9.3005
R11419 GND.n7970 GND.n7969 9.3005
R11420 GND.n7971 GND.n677 9.3005
R11421 GND.n7973 GND.n7972 9.3005
R11422 GND.n673 GND.n672 9.3005
R11423 GND.n7980 GND.n7979 9.3005
R11424 GND.n7981 GND.n671 9.3005
R11425 GND.n7983 GND.n7982 9.3005
R11426 GND.n667 GND.n666 9.3005
R11427 GND.n7990 GND.n7989 9.3005
R11428 GND.n7991 GND.n665 9.3005
R11429 GND.n7993 GND.n7992 9.3005
R11430 GND.n661 GND.n660 9.3005
R11431 GND.n8000 GND.n7999 9.3005
R11432 GND.n8001 GND.n659 9.3005
R11433 GND.n8003 GND.n8002 9.3005
R11434 GND.n655 GND.n654 9.3005
R11435 GND.n8010 GND.n8009 9.3005
R11436 GND.n8011 GND.n653 9.3005
R11437 GND.n8013 GND.n8012 9.3005
R11438 GND.n649 GND.n648 9.3005
R11439 GND.n8020 GND.n8019 9.3005
R11440 GND.n8021 GND.n647 9.3005
R11441 GND.n8023 GND.n8022 9.3005
R11442 GND.n643 GND.n642 9.3005
R11443 GND.n8030 GND.n8029 9.3005
R11444 GND.n8031 GND.n641 9.3005
R11445 GND.n8033 GND.n8032 9.3005
R11446 GND.n637 GND.n636 9.3005
R11447 GND.n8040 GND.n8039 9.3005
R11448 GND.n8041 GND.n635 9.3005
R11449 GND.n8043 GND.n8042 9.3005
R11450 GND.n631 GND.n630 9.3005
R11451 GND.n8050 GND.n8049 9.3005
R11452 GND.n8051 GND.n629 9.3005
R11453 GND.n8053 GND.n8052 9.3005
R11454 GND.n625 GND.n624 9.3005
R11455 GND.n8060 GND.n8059 9.3005
R11456 GND.n8061 GND.n623 9.3005
R11457 GND.n8063 GND.n8062 9.3005
R11458 GND.n619 GND.n618 9.3005
R11459 GND.n8070 GND.n8069 9.3005
R11460 GND.n8071 GND.n617 9.3005
R11461 GND.n8073 GND.n8072 9.3005
R11462 GND.n613 GND.n612 9.3005
R11463 GND.n8080 GND.n8079 9.3005
R11464 GND.n8081 GND.n611 9.3005
R11465 GND.n8083 GND.n8082 9.3005
R11466 GND.n607 GND.n606 9.3005
R11467 GND.n8090 GND.n8089 9.3005
R11468 GND.n8091 GND.n605 9.3005
R11469 GND.n8093 GND.n8092 9.3005
R11470 GND.n601 GND.n600 9.3005
R11471 GND.n8100 GND.n8099 9.3005
R11472 GND.n8101 GND.n599 9.3005
R11473 GND.n8103 GND.n8102 9.3005
R11474 GND.n595 GND.n594 9.3005
R11475 GND.n8110 GND.n8109 9.3005
R11476 GND.n8111 GND.n593 9.3005
R11477 GND.n8113 GND.n8112 9.3005
R11478 GND.n589 GND.n588 9.3005
R11479 GND.n8120 GND.n8119 9.3005
R11480 GND.n8121 GND.n587 9.3005
R11481 GND.n8123 GND.n8122 9.3005
R11482 GND.n583 GND.n582 9.3005
R11483 GND.n8130 GND.n8129 9.3005
R11484 GND.n8131 GND.n581 9.3005
R11485 GND.n8133 GND.n8132 9.3005
R11486 GND.n577 GND.n576 9.3005
R11487 GND.n8140 GND.n8139 9.3005
R11488 GND.n8141 GND.n575 9.3005
R11489 GND.n8143 GND.n8142 9.3005
R11490 GND.n571 GND.n570 9.3005
R11491 GND.n8150 GND.n8149 9.3005
R11492 GND.n8151 GND.n569 9.3005
R11493 GND.n8153 GND.n8152 9.3005
R11494 GND.n565 GND.n564 9.3005
R11495 GND.n8160 GND.n8159 9.3005
R11496 GND.n8161 GND.n563 9.3005
R11497 GND.n8163 GND.n8162 9.3005
R11498 GND.n559 GND.n558 9.3005
R11499 GND.n8170 GND.n8169 9.3005
R11500 GND.n8171 GND.n557 9.3005
R11501 GND.n8173 GND.n8172 9.3005
R11502 GND.n553 GND.n552 9.3005
R11503 GND.n8180 GND.n8179 9.3005
R11504 GND.n8181 GND.n551 9.3005
R11505 GND.n8183 GND.n8182 9.3005
R11506 GND.n547 GND.n546 9.3005
R11507 GND.n8190 GND.n8189 9.3005
R11508 GND.n8191 GND.n545 9.3005
R11509 GND.n8193 GND.n8192 9.3005
R11510 GND.n541 GND.n540 9.3005
R11511 GND.n8200 GND.n8199 9.3005
R11512 GND.n8201 GND.n539 9.3005
R11513 GND.n8204 GND.n8203 9.3005
R11514 GND.n8202 GND.n535 9.3005
R11515 GND.n8210 GND.n534 9.3005
R11516 GND.n8212 GND.n8211 9.3005
R11517 GND.n530 GND.n529 9.3005
R11518 GND.n8221 GND.n8220 9.3005
R11519 GND.n8222 GND.n528 9.3005
R11520 GND.n8224 GND.n8223 9.3005
R11521 GND.n524 GND.n523 9.3005
R11522 GND.n8231 GND.n8230 9.3005
R11523 GND.n8232 GND.n522 9.3005
R11524 GND.n8234 GND.n8233 9.3005
R11525 GND.n518 GND.n517 9.3005
R11526 GND.n8241 GND.n8240 9.3005
R11527 GND.n8242 GND.n516 9.3005
R11528 GND.n8244 GND.n8243 9.3005
R11529 GND.n512 GND.n511 9.3005
R11530 GND.n8251 GND.n8250 9.3005
R11531 GND.n8252 GND.n510 9.3005
R11532 GND.n8254 GND.n8253 9.3005
R11533 GND.n506 GND.n505 9.3005
R11534 GND.n8261 GND.n8260 9.3005
R11535 GND.n8262 GND.n504 9.3005
R11536 GND.n8264 GND.n8263 9.3005
R11537 GND.n500 GND.n499 9.3005
R11538 GND.n8271 GND.n8270 9.3005
R11539 GND.n8272 GND.n498 9.3005
R11540 GND.n8274 GND.n8273 9.3005
R11541 GND.n494 GND.n493 9.3005
R11542 GND.n8281 GND.n8280 9.3005
R11543 GND.n8282 GND.n492 9.3005
R11544 GND.n8284 GND.n8283 9.3005
R11545 GND.n488 GND.n487 9.3005
R11546 GND.n8291 GND.n8290 9.3005
R11547 GND.n8292 GND.n486 9.3005
R11548 GND.n8294 GND.n8293 9.3005
R11549 GND.n482 GND.n481 9.3005
R11550 GND.n8301 GND.n8300 9.3005
R11551 GND.n8302 GND.n480 9.3005
R11552 GND.n8304 GND.n8303 9.3005
R11553 GND.n476 GND.n475 9.3005
R11554 GND.n8311 GND.n8310 9.3005
R11555 GND.n8312 GND.n474 9.3005
R11556 GND.n8314 GND.n8313 9.3005
R11557 GND.n470 GND.n469 9.3005
R11558 GND.n8321 GND.n8320 9.3005
R11559 GND.n8322 GND.n468 9.3005
R11560 GND.n8324 GND.n8323 9.3005
R11561 GND.n464 GND.n463 9.3005
R11562 GND.n8331 GND.n8330 9.3005
R11563 GND.n8332 GND.n462 9.3005
R11564 GND.n8334 GND.n8333 9.3005
R11565 GND.n458 GND.n457 9.3005
R11566 GND.n8341 GND.n8340 9.3005
R11567 GND.n8342 GND.n456 9.3005
R11568 GND.n8344 GND.n8343 9.3005
R11569 GND.n452 GND.n451 9.3005
R11570 GND.n8351 GND.n8350 9.3005
R11571 GND.n8352 GND.n450 9.3005
R11572 GND.n8354 GND.n8353 9.3005
R11573 GND.n446 GND.n445 9.3005
R11574 GND.n8361 GND.n8360 9.3005
R11575 GND.n8362 GND.n444 9.3005
R11576 GND.n8364 GND.n8363 9.3005
R11577 GND.n440 GND.n439 9.3005
R11578 GND.n8371 GND.n8370 9.3005
R11579 GND.n8372 GND.n438 9.3005
R11580 GND.n8374 GND.n8373 9.3005
R11581 GND.n434 GND.n433 9.3005
R11582 GND.n8381 GND.n8380 9.3005
R11583 GND.n8382 GND.n432 9.3005
R11584 GND.n8384 GND.n8383 9.3005
R11585 GND.n428 GND.n427 9.3005
R11586 GND.n8391 GND.n8390 9.3005
R11587 GND.n8392 GND.n426 9.3005
R11588 GND.n8395 GND.n8394 9.3005
R11589 GND.n8214 GND.n8213 9.3005
R11590 GND.n85 GND.n84 9.3005
R11591 GND.n78 GND.n77 9.3005
R11592 GND.n100 GND.n99 9.3005
R11593 GND.n93 GND.n92 9.3005
R11594 GND.n116 GND.n115 9.3005
R11595 GND.n109 GND.n108 9.3005
R11596 GND.n132 GND.n131 9.3005
R11597 GND.n125 GND.n124 9.3005
R11598 GND.n6076 GND.n6075 9.3005
R11599 GND.n6083 GND.n6082 9.3005
R11600 GND.n6085 GND.n6084 9.3005
R11601 GND.n6072 GND.n6071 9.3005
R11602 GND.n6091 GND.n6090 9.3005
R11603 GND.n6093 GND.n6092 9.3005
R11604 GND.n6068 GND.n6067 9.3005
R11605 GND.n6099 GND.n6098 9.3005
R11606 GND.n6133 GND.n6132 9.3005
R11607 GND.n6136 GND.n6135 9.3005
R11608 GND.n6137 GND.n6049 9.3005
R11609 GND.n6141 GND.n6140 9.3005
R11610 GND.n6142 GND.n6048 9.3005
R11611 GND.n6144 GND.n6143 9.3005
R11612 GND.n6046 GND.n6045 9.3005
R11613 GND.n6156 GND.n6155 9.3005
R11614 GND.n6157 GND.n6044 9.3005
R11615 GND.n6159 GND.n6158 9.3005
R11616 GND.n6042 GND.n6041 9.3005
R11617 GND.n6171 GND.n6170 9.3005
R11618 GND.n6172 GND.n6040 9.3005
R11619 GND.n6174 GND.n6173 9.3005
R11620 GND.n6038 GND.n6037 9.3005
R11621 GND.n6186 GND.n6185 9.3005
R11622 GND.n6187 GND.n6036 9.3005
R11623 GND.n6196 GND.n6188 9.3005
R11624 GND.n6195 GND.n6189 9.3005
R11625 GND.n6194 GND.n6190 9.3005
R11626 GND.n6193 GND.n6191 9.3005
R11627 GND.n138 GND.n136 9.3005
R11628 GND.n6134 GND.n6050 9.3005
R11629 GND.n8511 GND.n8510 9.3005
R11630 GND.n139 GND.n137 9.3005
R11631 GND.n5972 GND.n5971 9.3005
R11632 GND.n6218 GND.n6217 9.3005
R11633 GND.n6219 GND.n5970 9.3005
R11634 GND.n6221 GND.n6220 9.3005
R11635 GND.n5968 GND.n5967 9.3005
R11636 GND.n6233 GND.n6232 9.3005
R11637 GND.n6234 GND.n5966 9.3005
R11638 GND.n6237 GND.n6236 9.3005
R11639 GND.n6235 GND.n5960 9.3005
R11640 GND.n6351 GND.n5961 9.3005
R11641 GND.n6350 GND.n5962 9.3005
R11642 GND.n6349 GND.n5963 9.3005
R11643 GND.n6248 GND.n5964 9.3005
R11644 GND.n6339 GND.n6249 9.3005
R11645 GND.n6338 GND.n6250 9.3005
R11646 GND.n6337 GND.n6251 9.3005
R11647 GND.n6254 GND.n6252 9.3005
R11648 GND.n6300 GND.n6255 9.3005
R11649 GND.n6299 GND.n6256 9.3005
R11650 GND.n6298 GND.n6297 9.3005
R11651 GND.n6268 GND.n6267 9.3005
R11652 GND.n6277 GND.n6276 9.3005
R11653 GND.n6278 GND.n6266 9.3005
R11654 GND.n6280 GND.n6279 9.3005
R11655 GND.n6264 GND.n6263 9.3005
R11656 GND.n6287 GND.n6286 9.3005
R11657 GND.n6288 GND.n6262 9.3005
R11658 GND.n6290 GND.n6289 9.3005
R11659 GND.n6260 GND.n6257 9.3005
R11660 GND.n6296 GND.n6295 9.3005
R11661 GND.n6270 GND.n6269 9.3005
R11662 GND.n380 GND.n379 9.3005
R11663 GND.n378 GND.n281 9.3005
R11664 GND.n377 GND.n376 9.3005
R11665 GND.n373 GND.n282 9.3005
R11666 GND.n370 GND.n283 9.3005
R11667 GND.n369 GND.n284 9.3005
R11668 GND.n366 GND.n285 9.3005
R11669 GND.n365 GND.n286 9.3005
R11670 GND.n362 GND.n361 9.3005
R11671 GND.n360 GND.n287 9.3005
R11672 GND.n359 GND.n358 9.3005
R11673 GND.n355 GND.n290 9.3005
R11674 GND.n352 GND.n291 9.3005
R11675 GND.n351 GND.n292 9.3005
R11676 GND.n348 GND.n293 9.3005
R11677 GND.n347 GND.n294 9.3005
R11678 GND.n344 GND.n295 9.3005
R11679 GND.n343 GND.n296 9.3005
R11680 GND.n340 GND.n297 9.3005
R11681 GND.n339 GND.n338 9.3005
R11682 GND.n337 GND.n298 9.3005
R11683 GND.n336 GND.n335 9.3005
R11684 GND.n332 GND.n303 9.3005
R11685 GND.n331 GND.n304 9.3005
R11686 GND.n328 GND.n305 9.3005
R11687 GND.n327 GND.n306 9.3005
R11688 GND.n324 GND.n307 9.3005
R11689 GND.n323 GND.n308 9.3005
R11690 GND.n320 GND.n309 9.3005
R11691 GND.n319 GND.n310 9.3005
R11692 GND.n316 GND.n315 9.3005
R11693 GND.n314 GND.n311 9.3005
R11694 GND.n381 GND.n280 9.3005
R11695 GND.n6445 GND.n6444 9.3005
R11696 GND.n5826 GND.n5825 9.3005
R11697 GND.n5851 GND.n5850 9.3005
R11698 GND.n6432 GND.n5852 9.3005
R11699 GND.n6431 GND.n5853 9.3005
R11700 GND.n6430 GND.n5854 9.3005
R11701 GND.n6150 GND.n5855 9.3005
R11702 GND.n6420 GND.n5873 9.3005
R11703 GND.n6419 GND.n5874 9.3005
R11704 GND.n6418 GND.n5875 9.3005
R11705 GND.n6165 GND.n5876 9.3005
R11706 GND.n6408 GND.n5894 9.3005
R11707 GND.n6407 GND.n5895 9.3005
R11708 GND.n6406 GND.n5896 9.3005
R11709 GND.n6180 GND.n5897 9.3005
R11710 GND.n6396 GND.n5913 9.3005
R11711 GND.n6395 GND.n5914 9.3005
R11712 GND.n6394 GND.n5915 9.3005
R11713 GND.n6203 GND.n5916 9.3005
R11714 GND.n6204 GND.n5935 9.3005
R11715 GND.n6377 GND.n5936 9.3005
R11716 GND.n6376 GND.n5937 9.3005
R11717 GND.n6375 GND.n5938 9.3005
R11718 GND.n6211 GND.n5939 9.3005
R11719 GND.n6212 GND.n166 9.3005
R11720 GND.n8499 GND.n167 9.3005
R11721 GND.n8498 GND.n168 9.3005
R11722 GND.n8497 GND.n169 9.3005
R11723 GND.n6227 GND.n170 9.3005
R11724 GND.n8487 GND.n187 9.3005
R11725 GND.n8486 GND.n188 9.3005
R11726 GND.n8485 GND.n189 9.3005
R11727 GND.n6243 GND.n190 9.3005
R11728 GND.n8475 GND.n207 9.3005
R11729 GND.n8474 GND.n208 9.3005
R11730 GND.n8473 GND.n209 9.3005
R11731 GND.n6246 GND.n210 9.3005
R11732 GND.n8463 GND.n228 9.3005
R11733 GND.n8462 GND.n229 9.3005
R11734 GND.n8461 GND.n230 9.3005
R11735 GND.n6253 GND.n231 9.3005
R11736 GND.n8451 GND.n248 9.3005
R11737 GND.n8450 GND.n8449 9.3005
R11738 GND.n6446 GND.n5824 9.3005
R11739 GND.n6444 GND.n6443 9.3005
R11740 GND.n6442 GND.n5826 9.3005
R11741 GND.n5851 GND.n5827 9.3005
R11742 GND.n6047 GND.n5852 9.3005
R11743 GND.n6148 GND.n5853 9.3005
R11744 GND.n6149 GND.n5854 9.3005
R11745 GND.n6151 GND.n6150 9.3005
R11746 GND.n6043 GND.n5873 9.3005
R11747 GND.n6163 GND.n5874 9.3005
R11748 GND.n6164 GND.n5875 9.3005
R11749 GND.n6166 GND.n6165 9.3005
R11750 GND.n6039 GND.n5894 9.3005
R11751 GND.n6178 GND.n5895 9.3005
R11752 GND.n6179 GND.n5896 9.3005
R11753 GND.n6181 GND.n6180 9.3005
R11754 GND.n5976 GND.n5913 9.3005
R11755 GND.n6200 GND.n5914 9.3005
R11756 GND.n6201 GND.n5915 9.3005
R11757 GND.n6203 GND.n6202 9.3005
R11758 GND.n6206 GND.n6204 9.3005
R11759 GND.n6207 GND.n5936 9.3005
R11760 GND.n6208 GND.n5937 9.3005
R11761 GND.n6209 GND.n5938 9.3005
R11762 GND.n6211 GND.n6210 9.3005
R11763 GND.n6213 GND.n6212 9.3005
R11764 GND.n5969 GND.n167 9.3005
R11765 GND.n6225 GND.n168 9.3005
R11766 GND.n6226 GND.n169 9.3005
R11767 GND.n6228 GND.n6227 9.3005
R11768 GND.n5965 GND.n187 9.3005
R11769 GND.n6241 GND.n188 9.3005
R11770 GND.n6242 GND.n189 9.3005
R11771 GND.n6244 GND.n6243 9.3005
R11772 GND.n6245 GND.n207 9.3005
R11773 GND.n6345 GND.n208 9.3005
R11774 GND.n6344 GND.n209 9.3005
R11775 GND.n6343 GND.n6246 9.3005
R11776 GND.n6247 GND.n228 9.3005
R11777 GND.n6306 GND.n229 9.3005
R11778 GND.n6305 GND.n230 9.3005
R11779 GND.n6304 GND.n6253 9.3005
R11780 GND.n250 GND.n248 9.3005
R11781 GND.n8449 GND.n8448 9.3005
R11782 GND.n5824 GND.n5818 9.3005
R11783 GND.n6455 GND.n6454 9.3005
R11784 GND.n6456 GND.n5810 9.3005
R11785 GND.n6459 GND.n5809 9.3005
R11786 GND.n6460 GND.n5808 9.3005
R11787 GND.n6463 GND.n5807 9.3005
R11788 GND.n6464 GND.n5806 9.3005
R11789 GND.n6467 GND.n5805 9.3005
R11790 GND.n6468 GND.n5804 9.3005
R11791 GND.n6471 GND.n5803 9.3005
R11792 GND.n6473 GND.n5802 9.3005
R11793 GND.n6474 GND.n5799 9.3005
R11794 GND.n6475 GND.n5797 9.3005
R11795 GND.n6478 GND.n5796 9.3005
R11796 GND.n6479 GND.n5795 9.3005
R11797 GND.n6482 GND.n5794 9.3005
R11798 GND.n6484 GND.n5793 9.3005
R11799 GND.n6488 GND.n3085 9.3005
R11800 GND.n6489 GND.n3084 9.3005
R11801 GND.n6492 GND.n3083 9.3005
R11802 GND.n6493 GND.n3080 9.3005
R11803 GND.n6496 GND.n3079 9.3005
R11804 GND.n6497 GND.n3078 9.3005
R11805 GND.n6500 GND.n3077 9.3005
R11806 GND.n6501 GND.n3076 9.3005
R11807 GND.n6504 GND.n3075 9.3005
R11808 GND.n6506 GND.n3074 9.3005
R11809 GND.n6507 GND.n3073 9.3005
R11810 GND.n6508 GND.n3072 9.3005
R11811 GND.n6509 GND.n3071 9.3005
R11812 GND.n6453 GND.n5815 9.3005
R11813 GND.n6452 GND.n6451 9.3005
R11814 GND.n5838 GND.n5835 9.3005
R11815 GND.n6438 GND.n5839 9.3005
R11816 GND.n6437 GND.n5840 9.3005
R11817 GND.n6436 GND.n5841 9.3005
R11818 GND.n5862 GND.n5842 9.3005
R11819 GND.n6426 GND.n5863 9.3005
R11820 GND.n6425 GND.n5864 9.3005
R11821 GND.n6424 GND.n5865 9.3005
R11822 GND.n5883 GND.n5866 9.3005
R11823 GND.n6414 GND.n5884 9.3005
R11824 GND.n6413 GND.n5885 9.3005
R11825 GND.n6412 GND.n5886 9.3005
R11826 GND.n5904 GND.n5887 9.3005
R11827 GND.n6402 GND.n5905 9.3005
R11828 GND.n6401 GND.n5906 9.3005
R11829 GND.n6400 GND.n150 9.3005
R11830 GND.n157 GND.n149 9.3005
R11831 GND.n8493 GND.n177 9.3005
R11832 GND.n8492 GND.n178 9.3005
R11833 GND.n8491 GND.n179 9.3005
R11834 GND.n196 GND.n180 9.3005
R11835 GND.n8481 GND.n197 9.3005
R11836 GND.n8480 GND.n198 9.3005
R11837 GND.n8479 GND.n199 9.3005
R11838 GND.n217 GND.n200 9.3005
R11839 GND.n8469 GND.n218 9.3005
R11840 GND.n8468 GND.n219 9.3005
R11841 GND.n8467 GND.n220 9.3005
R11842 GND.n237 GND.n221 9.3005
R11843 GND.n8457 GND.n238 9.3005
R11844 GND.n8456 GND.n239 9.3005
R11845 GND.n8455 GND.n240 9.3005
R11846 GND.n279 GND.n241 9.3005
R11847 GND.n5837 GND.n5836 9.3005
R11848 GND.n8504 GND.n154 9.3005
R11849 GND.n8504 GND.n8503 9.3005
R11850 GND.n2361 GND.n2359 9.3005
R11851 GND.n2383 GND.n2362 9.3005
R11852 GND.n2382 GND.n2363 9.3005
R11853 GND.n2381 GND.n2364 9.3005
R11854 GND.n2367 GND.n2365 9.3005
R11855 GND.n2377 GND.n2368 9.3005
R11856 GND.n2376 GND.n2369 9.3005
R11857 GND.n2375 GND.n2370 9.3005
R11858 GND.n2373 GND.n2372 9.3005
R11859 GND.n2371 GND.n1999 9.3005
R11860 GND.n1997 GND.n1996 9.3005
R11861 GND.n2482 GND.n2481 9.3005
R11862 GND.n2483 GND.n1995 9.3005
R11863 GND.n2488 GND.n2484 9.3005
R11864 GND.n2487 GND.n2486 9.3005
R11865 GND.n2485 GND.n1963 9.3005
R11866 GND.n1961 GND.n1960 9.3005
R11867 GND.n2523 GND.n2522 9.3005
R11868 GND.n2524 GND.n1959 9.3005
R11869 GND.n6970 GND.n2525 9.3005
R11870 GND.n6969 GND.n2526 9.3005
R11871 GND.n6968 GND.n2527 9.3005
R11872 GND.n2532 GND.n2528 9.3005
R11873 GND.n6962 GND.n2533 9.3005
R11874 GND.n6961 GND.n2534 9.3005
R11875 GND.n6960 GND.n2535 9.3005
R11876 GND.n2550 GND.n2536 9.3005
R11877 GND.n6948 GND.n2551 9.3005
R11878 GND.n6947 GND.n2552 9.3005
R11879 GND.n6946 GND.n2553 9.3005
R11880 GND.n2568 GND.n2554 9.3005
R11881 GND.n6935 GND.n2569 9.3005
R11882 GND.n6934 GND.n2570 9.3005
R11883 GND.n6933 GND.n2571 9.3005
R11884 GND.n2585 GND.n2572 9.3005
R11885 GND.n6921 GND.n2586 9.3005
R11886 GND.n6920 GND.n2587 9.3005
R11887 GND.n6919 GND.n2588 9.3005
R11888 GND.n2603 GND.n2589 9.3005
R11889 GND.n6907 GND.n2604 9.3005
R11890 GND.n6906 GND.n2605 9.3005
R11891 GND.n6905 GND.n2606 9.3005
R11892 GND.n2621 GND.n2607 9.3005
R11893 GND.n6893 GND.n2622 9.3005
R11894 GND.n6892 GND.n2623 9.3005
R11895 GND.n6891 GND.n2624 9.3005
R11896 GND.n2639 GND.n2625 9.3005
R11897 GND.n6879 GND.n2640 9.3005
R11898 GND.n6878 GND.n2641 9.3005
R11899 GND.n6877 GND.n2642 9.3005
R11900 GND.n2656 GND.n2643 9.3005
R11901 GND.n6865 GND.n2657 9.3005
R11902 GND.n6864 GND.n2658 9.3005
R11903 GND.n6863 GND.n2659 9.3005
R11904 GND.n3888 GND.n2660 9.3005
R11905 GND.n4352 GND.n4351 9.3005
R11906 GND.n4353 GND.n3887 9.3005
R11907 GND.n4355 GND.n4354 9.3005
R11908 GND.n3872 GND.n3871 9.3005
R11909 GND.n4390 GND.n4389 9.3005
R11910 GND.n4391 GND.n3870 9.3005
R11911 GND.n4406 GND.n4392 9.3005
R11912 GND.n4405 GND.n4393 9.3005
R11913 GND.n4404 GND.n4394 9.3005
R11914 GND.n4396 GND.n4395 9.3005
R11915 GND.n4398 GND.n4397 9.3005
R11916 GND.n3832 GND.n3831 9.3005
R11917 GND.n4479 GND.n4478 9.3005
R11918 GND.n4480 GND.n3830 9.3005
R11919 GND.n4484 GND.n4481 9.3005
R11920 GND.n4483 GND.n4482 9.3005
R11921 GND.n3801 GND.n3800 9.3005
R11922 GND.n4525 GND.n4524 9.3005
R11923 GND.n4526 GND.n3799 9.3005
R11924 GND.n4528 GND.n4527 9.3005
R11925 GND.n3783 GND.n3782 9.3005
R11926 GND.n4582 GND.n4581 9.3005
R11927 GND.n4583 GND.n3781 9.3005
R11928 GND.n4585 GND.n4584 9.3005
R11929 GND.n3760 GND.n3759 9.3005
R11930 GND.n4610 GND.n4609 9.3005
R11931 GND.n4611 GND.n3758 9.3005
R11932 GND.n4615 GND.n4612 9.3005
R11933 GND.n4614 GND.n4613 9.3005
R11934 GND.n3731 GND.n3730 9.3005
R11935 GND.n4682 GND.n4681 9.3005
R11936 GND.n4683 GND.n3729 9.3005
R11937 GND.n4685 GND.n4684 9.3005
R11938 GND.n3710 GND.n3709 9.3005
R11939 GND.n4708 GND.n4707 9.3005
R11940 GND.n4709 GND.n3708 9.3005
R11941 GND.n4711 GND.n4710 9.3005
R11942 GND.n3689 GND.n3688 9.3005
R11943 GND.n4743 GND.n4742 9.3005
R11944 GND.n4744 GND.n3687 9.3005
R11945 GND.n4746 GND.n4745 9.3005
R11946 GND.n3672 GND.n3671 9.3005
R11947 GND.n4786 GND.n4785 9.3005
R11948 GND.n4787 GND.n3670 9.3005
R11949 GND.n4791 GND.n4788 9.3005
R11950 GND.n4790 GND.n4789 9.3005
R11951 GND.n3643 GND.n3642 9.3005
R11952 GND.n4859 GND.n4858 9.3005
R11953 GND.n4860 GND.n3641 9.3005
R11954 GND.n4862 GND.n4861 9.3005
R11955 GND.n3623 GND.n3622 9.3005
R11956 GND.n4886 GND.n4885 9.3005
R11957 GND.n4887 GND.n3621 9.3005
R11958 GND.n4889 GND.n4888 9.3005
R11959 GND.n3601 GND.n3600 9.3005
R11960 GND.n4920 GND.n4919 9.3005
R11961 GND.n4921 GND.n3599 9.3005
R11962 GND.n4923 GND.n4922 9.3005
R11963 GND.n3584 GND.n3583 9.3005
R11964 GND.n4963 GND.n4962 9.3005
R11965 GND.n4964 GND.n3582 9.3005
R11966 GND.n4968 GND.n4965 9.3005
R11967 GND.n4967 GND.n4966 9.3005
R11968 GND.n3555 GND.n3554 9.3005
R11969 GND.n5035 GND.n5034 9.3005
R11970 GND.n5036 GND.n3553 9.3005
R11971 GND.n5038 GND.n5037 9.3005
R11972 GND.n3534 GND.n3533 9.3005
R11973 GND.n5061 GND.n5060 9.3005
R11974 GND.n5062 GND.n3532 9.3005
R11975 GND.n5064 GND.n5063 9.3005
R11976 GND.n3512 GND.n3511 9.3005
R11977 GND.n5095 GND.n5094 9.3005
R11978 GND.n5096 GND.n3510 9.3005
R11979 GND.n5098 GND.n5097 9.3005
R11980 GND.n3495 GND.n3494 9.3005
R11981 GND.n5139 GND.n5138 9.3005
R11982 GND.n5140 GND.n3493 9.3005
R11983 GND.n5144 GND.n5141 9.3005
R11984 GND.n5143 GND.n5142 9.3005
R11985 GND.n3466 GND.n3465 9.3005
R11986 GND.n5210 GND.n5209 9.3005
R11987 GND.n5211 GND.n3464 9.3005
R11988 GND.n5213 GND.n5212 9.3005
R11989 GND.n3445 GND.n3444 9.3005
R11990 GND.n5236 GND.n5235 9.3005
R11991 GND.n5237 GND.n3443 9.3005
R11992 GND.n5239 GND.n5238 9.3005
R11993 GND.n3423 GND.n3422 9.3005
R11994 GND.n5270 GND.n5269 9.3005
R11995 GND.n5271 GND.n3421 9.3005
R11996 GND.n5273 GND.n5272 9.3005
R11997 GND.n3406 GND.n3405 9.3005
R11998 GND.n5313 GND.n5312 9.3005
R11999 GND.n5314 GND.n3404 9.3005
R12000 GND.n5318 GND.n5315 9.3005
R12001 GND.n5317 GND.n5316 9.3005
R12002 GND.n3377 GND.n3376 9.3005
R12003 GND.n5387 GND.n5386 9.3005
R12004 GND.n5388 GND.n3375 9.3005
R12005 GND.n5390 GND.n5389 9.3005
R12006 GND.n3358 GND.n3357 9.3005
R12007 GND.n5413 GND.n5412 9.3005
R12008 GND.n5414 GND.n3356 9.3005
R12009 GND.n5416 GND.n5415 9.3005
R12010 GND.n3337 GND.n3336 9.3005
R12011 GND.n5448 GND.n5447 9.3005
R12012 GND.n5449 GND.n3335 9.3005
R12013 GND.n5451 GND.n5450 9.3005
R12014 GND.n3320 GND.n3319 9.3005
R12015 GND.n5491 GND.n5490 9.3005
R12016 GND.n5492 GND.n3318 9.3005
R12017 GND.n5496 GND.n5493 9.3005
R12018 GND.n5495 GND.n5494 9.3005
R12019 GND.n3291 GND.n3290 9.3005
R12020 GND.n5541 GND.n5540 9.3005
R12021 GND.n5542 GND.n3289 9.3005
R12022 GND.n5546 GND.n5543 9.3005
R12023 GND.n5545 GND.n5544 9.3005
R12024 GND.n3271 GND.n3270 9.3005
R12025 GND.n5569 GND.n5568 9.3005
R12026 GND.n5570 GND.n3269 9.3005
R12027 GND.n5583 GND.n5571 9.3005
R12028 GND.n5582 GND.n5572 9.3005
R12029 GND.n5581 GND.n5573 9.3005
R12030 GND.n5576 GND.n5575 9.3005
R12031 GND.n5574 GND.n2908 9.3005
R12032 GND.n6623 GND.n2909 9.3005
R12033 GND.n6622 GND.n2910 9.3005
R12034 GND.n6621 GND.n2911 9.3005
R12035 GND.n2925 GND.n2912 9.3005
R12036 GND.n6609 GND.n2926 9.3005
R12037 GND.n6608 GND.n2927 9.3005
R12038 GND.n6607 GND.n2928 9.3005
R12039 GND.n2943 GND.n2929 9.3005
R12040 GND.n6595 GND.n2944 9.3005
R12041 GND.n6594 GND.n2945 9.3005
R12042 GND.n6593 GND.n2946 9.3005
R12043 GND.n2961 GND.n2947 9.3005
R12044 GND.n6581 GND.n2962 9.3005
R12045 GND.n6580 GND.n2963 9.3005
R12046 GND.n6579 GND.n2964 9.3005
R12047 GND.n2979 GND.n2965 9.3005
R12048 GND.n6567 GND.n2980 9.3005
R12049 GND.n6566 GND.n2981 9.3005
R12050 GND.n6565 GND.n2982 9.3005
R12051 GND.n2996 GND.n2983 9.3005
R12052 GND.n6553 GND.n2997 9.3005
R12053 GND.n6552 GND.n2998 9.3005
R12054 GND.n6551 GND.n2999 9.3005
R12055 GND.n3014 GND.n3000 9.3005
R12056 GND.n6539 GND.n3015 9.3005
R12057 GND.n6538 GND.n3016 9.3005
R12058 GND.n6537 GND.n3017 9.3005
R12059 GND.n3031 GND.n3018 9.3005
R12060 GND.n6525 GND.n3032 9.3005
R12061 GND.n6524 GND.n3033 9.3005
R12062 GND.n6523 GND.n3034 9.3005
R12063 GND.n3040 GND.n3035 9.3005
R12064 GND.n6517 GND.n3041 9.3005
R12065 GND.n6516 GND.n3042 9.3005
R12066 GND.n6515 GND.n3043 9.3005
R12067 GND.n5996 GND.n3044 9.3005
R12068 GND.n5997 GND.n5995 9.3005
R12069 GND.n5999 GND.n5998 9.3005
R12070 GND.n5993 GND.n5992 9.3005
R12071 GND.n6004 GND.n6003 9.3005
R12072 GND.n6005 GND.n5991 9.3005
R12073 GND.n6007 GND.n6006 9.3005
R12074 GND.n5989 GND.n5988 9.3005
R12075 GND.n6012 GND.n6011 9.3005
R12076 GND.n6013 GND.n5987 9.3005
R12077 GND.n6015 GND.n6014 9.3005
R12078 GND.n5985 GND.n5984 9.3005
R12079 GND.n6020 GND.n6019 9.3005
R12080 GND.n6021 GND.n5983 9.3005
R12081 GND.n6023 GND.n6022 9.3005
R12082 GND.n5981 GND.n5980 9.3005
R12083 GND.n6028 GND.n6027 9.3005
R12084 GND.n6029 GND.n5979 9.3005
R12085 GND.n6033 GND.n6030 9.3005
R12086 GND.n6363 GND.n5949 9.3005
R12087 GND.n6362 GND.n5950 9.3005
R12088 GND.n5953 GND.n5951 9.3005
R12089 GND.n6358 GND.n5954 9.3005
R12090 GND.n6357 GND.n5955 9.3005
R12091 GND.n6356 GND.n5956 9.3005
R12092 GND.n6315 GND.n5957 9.3005
R12093 GND.n6316 GND.n6314 9.3005
R12094 GND.n6318 GND.n6317 9.3005
R12095 GND.n6312 GND.n6311 9.3005
R12096 GND.n6323 GND.n6322 9.3005
R12097 GND.n6324 GND.n6310 9.3005
R12098 GND.n6332 GND.n6325 9.3005
R12099 GND.n6331 GND.n6326 9.3005
R12100 GND.n6330 GND.n6328 9.3005
R12101 GND.n6327 GND.n256 9.3005
R12102 GND.n8443 GND.n257 9.3005
R12103 GND.n8442 GND.n258 9.3005
R12104 GND.n8441 GND.n259 9.3005
R12105 GND.n386 GND.n260 9.3005
R12106 GND.n8435 GND.n387 9.3005
R12107 GND.n8434 GND.n388 9.3005
R12108 GND.n8433 GND.n389 9.3005
R12109 GND.n394 GND.n390 9.3005
R12110 GND.n8427 GND.n395 9.3005
R12111 GND.n8426 GND.n396 9.3005
R12112 GND.n8425 GND.n397 9.3005
R12113 GND.n402 GND.n398 9.3005
R12114 GND.n8419 GND.n403 9.3005
R12115 GND.n8418 GND.n404 9.3005
R12116 GND.n8417 GND.n405 9.3005
R12117 GND.n410 GND.n406 9.3005
R12118 GND.n8411 GND.n411 9.3005
R12119 GND.n8410 GND.n412 9.3005
R12120 GND.n8409 GND.n413 9.3005
R12121 GND.n418 GND.n414 9.3005
R12122 GND.n8403 GND.n419 9.3005
R12123 GND.n8402 GND.n420 9.3005
R12124 GND.n8401 GND.n421 9.3005
R12125 GND.n8393 GND.n422 9.3005
R12126 GND.n7120 GND.n7119 9.3005
R12127 GND.n7121 GND.n1281 9.3005
R12128 GND.n7124 GND.n1280 9.3005
R12129 GND.n7125 GND.n1279 9.3005
R12130 GND.n7128 GND.n1278 9.3005
R12131 GND.n7129 GND.n1277 9.3005
R12132 GND.n7132 GND.n1276 9.3005
R12133 GND.n7133 GND.n1275 9.3005
R12134 GND.n7136 GND.n1274 9.3005
R12135 GND.n7138 GND.n1273 9.3005
R12136 GND.n7139 GND.n1270 9.3005
R12137 GND.n7140 GND.n1268 9.3005
R12138 GND.n7143 GND.n1267 9.3005
R12139 GND.n7144 GND.n1266 9.3005
R12140 GND.n7147 GND.n1265 9.3005
R12141 GND.n7148 GND.n1264 9.3005
R12142 GND.n7151 GND.n1263 9.3005
R12143 GND.n7152 GND.n1262 9.3005
R12144 GND.n7155 GND.n1261 9.3005
R12145 GND.n7156 GND.n1260 9.3005
R12146 GND.n7159 GND.n1259 9.3005
R12147 GND.n7160 GND.n1256 9.3005
R12148 GND.n7163 GND.n1255 9.3005
R12149 GND.n7164 GND.n1254 9.3005
R12150 GND.n7167 GND.n1253 9.3005
R12151 GND.n7168 GND.n1252 9.3005
R12152 GND.n7171 GND.n1251 9.3005
R12153 GND.n7173 GND.n1250 9.3005
R12154 GND.n7174 GND.n1249 9.3005
R12155 GND.n7175 GND.n1248 9.3005
R12156 GND.n7176 GND.n1247 9.3005
R12157 GND.n7118 GND.n1286 9.3005
R12158 GND.n7117 GND.n7116 9.3005
R12159 GND.n2171 GND.n2170 9.3005
R12160 GND.n2149 GND.n2148 9.3005
R12161 GND.n2272 GND.n2271 9.3005
R12162 GND.n2273 GND.n2147 9.3005
R12163 GND.n2277 GND.n2274 9.3005
R12164 GND.n2276 GND.n2275 9.3005
R12165 GND.n2126 GND.n2125 9.3005
R12166 GND.n2296 GND.n2295 9.3005
R12167 GND.n2297 GND.n2124 9.3005
R12168 GND.n2301 GND.n2298 9.3005
R12169 GND.n2300 GND.n2299 9.3005
R12170 GND.n2103 GND.n2102 9.3005
R12171 GND.n2321 GND.n2320 9.3005
R12172 GND.n2322 GND.n2101 9.3005
R12173 GND.n2324 GND.n2323 9.3005
R12174 GND.n2054 GND.n2047 9.3005
R12175 GND.n2420 GND.n2419 9.3005
R12176 GND.n2026 GND.n2025 9.3005
R12177 GND.n2442 GND.n2441 9.3005
R12178 GND.n2443 GND.n2024 9.3005
R12179 GND.n2447 GND.n2444 9.3005
R12180 GND.n2446 GND.n2445 9.3005
R12181 GND.n2005 GND.n2004 9.3005
R12182 GND.n2471 GND.n2470 9.3005
R12183 GND.n2472 GND.n2003 9.3005
R12184 GND.n2474 GND.n2473 9.3005
R12185 GND.n1974 GND.n1973 9.3005
R12186 GND.n2504 GND.n2503 9.3005
R12187 GND.n2505 GND.n1972 9.3005
R12188 GND.n2509 GND.n2506 9.3005
R12189 GND.n2508 GND.n2507 9.3005
R12190 GND.n1387 GND.n1386 9.3005
R12191 GND.n7042 GND.n7041 9.3005
R12192 GND.n2169 GND.n2168 9.3005
R12193 GND.n2418 GND.n2052 9.3005
R12194 GND.n2421 GND.n2418 9.3005
R12195 GND.n1181 GND.n1180 9.3005
R12196 GND.n7217 GND.n1185 9.3005
R12197 GND.n7216 GND.n1186 9.3005
R12198 GND.n7215 GND.n1187 9.3005
R12199 GND.n1192 GND.n1188 9.3005
R12200 GND.n7209 GND.n1193 9.3005
R12201 GND.n7208 GND.n1194 9.3005
R12202 GND.n7207 GND.n1195 9.3005
R12203 GND.n1200 GND.n1196 9.3005
R12204 GND.n7201 GND.n1201 9.3005
R12205 GND.n7200 GND.n1202 9.3005
R12206 GND.n7199 GND.n1203 9.3005
R12207 GND.n1208 GND.n1204 9.3005
R12208 GND.n7193 GND.n1209 9.3005
R12209 GND.n7192 GND.n1210 9.3005
R12210 GND.n7191 GND.n1211 9.3005
R12211 GND.n1216 GND.n1212 9.3005
R12212 GND.n7185 GND.n1217 9.3005
R12213 GND.n7184 GND.n1218 9.3005
R12214 GND.n7183 GND.n1219 9.3005
R12215 GND.n2162 GND.n1220 9.3005
R12216 GND.n2163 GND.n2161 9.3005
R12217 GND.n2165 GND.n2164 9.3005
R12218 GND.n2159 GND.n2158 9.3005
R12219 GND.n2221 GND.n2220 9.3005
R12220 GND.n2222 GND.n2157 9.3005
R12221 GND.n2262 GND.n2223 9.3005
R12222 GND.n2261 GND.n2224 9.3005
R12223 GND.n2260 GND.n2225 9.3005
R12224 GND.n2228 GND.n2226 9.3005
R12225 GND.n2256 GND.n2229 9.3005
R12226 GND.n2255 GND.n2230 9.3005
R12227 GND.n2254 GND.n2231 9.3005
R12228 GND.n2234 GND.n2232 9.3005
R12229 GND.n2250 GND.n2235 9.3005
R12230 GND.n2249 GND.n2236 9.3005
R12231 GND.n2248 GND.n2237 9.3005
R12232 GND.n2240 GND.n2238 9.3005
R12233 GND.n2244 GND.n2241 9.3005
R12234 GND.n7224 GND.n7223 9.3005
R12235 GND.n7227 GND.n1179 9.3005
R12236 GND.n1178 GND.n1174 9.3005
R12237 GND.n7233 GND.n1173 9.3005
R12238 GND.n7234 GND.n1172 9.3005
R12239 GND.n7235 GND.n1171 9.3005
R12240 GND.n1170 GND.n1166 9.3005
R12241 GND.n7241 GND.n1165 9.3005
R12242 GND.n7242 GND.n1164 9.3005
R12243 GND.n7243 GND.n1163 9.3005
R12244 GND.n1162 GND.n1158 9.3005
R12245 GND.n7249 GND.n1157 9.3005
R12246 GND.n7250 GND.n1156 9.3005
R12247 GND.n7251 GND.n1155 9.3005
R12248 GND.n1154 GND.n1150 9.3005
R12249 GND.n7257 GND.n1149 9.3005
R12250 GND.n7258 GND.n1148 9.3005
R12251 GND.n7259 GND.n1147 9.3005
R12252 GND.n1146 GND.n1142 9.3005
R12253 GND.n7265 GND.n1141 9.3005
R12254 GND.n7266 GND.n1140 9.3005
R12255 GND.n7267 GND.n1139 9.3005
R12256 GND.n1138 GND.n1134 9.3005
R12257 GND.n7273 GND.n1133 9.3005
R12258 GND.n7274 GND.n1132 9.3005
R12259 GND.n7275 GND.n1131 9.3005
R12260 GND.n1130 GND.n1126 9.3005
R12261 GND.n7281 GND.n1125 9.3005
R12262 GND.n7282 GND.n1124 9.3005
R12263 GND.n7283 GND.n1123 9.3005
R12264 GND.n1122 GND.n1118 9.3005
R12265 GND.n7289 GND.n1117 9.3005
R12266 GND.n7290 GND.n1116 9.3005
R12267 GND.n7291 GND.n1115 9.3005
R12268 GND.n1114 GND.n1110 9.3005
R12269 GND.n7297 GND.n1109 9.3005
R12270 GND.n7298 GND.n1108 9.3005
R12271 GND.n7299 GND.n1107 9.3005
R12272 GND.n1106 GND.n1102 9.3005
R12273 GND.n7305 GND.n1101 9.3005
R12274 GND.n7306 GND.n1100 9.3005
R12275 GND.n7307 GND.n1099 9.3005
R12276 GND.n1098 GND.n1094 9.3005
R12277 GND.n7313 GND.n1093 9.3005
R12278 GND.n7314 GND.n1092 9.3005
R12279 GND.n7315 GND.n1091 9.3005
R12280 GND.n1090 GND.n1086 9.3005
R12281 GND.n7321 GND.n1085 9.3005
R12282 GND.n7322 GND.n1084 9.3005
R12283 GND.n7323 GND.n1083 9.3005
R12284 GND.n1082 GND.n1078 9.3005
R12285 GND.n7329 GND.n1077 9.3005
R12286 GND.n7330 GND.n1076 9.3005
R12287 GND.n7331 GND.n1075 9.3005
R12288 GND.n1074 GND.n1070 9.3005
R12289 GND.n7337 GND.n1069 9.3005
R12290 GND.n7338 GND.n1068 9.3005
R12291 GND.n7339 GND.n1067 9.3005
R12292 GND.n1066 GND.n1062 9.3005
R12293 GND.n7345 GND.n1061 9.3005
R12294 GND.n7346 GND.n1060 9.3005
R12295 GND.n7347 GND.n1059 9.3005
R12296 GND.n1058 GND.n1054 9.3005
R12297 GND.n7353 GND.n1053 9.3005
R12298 GND.n7354 GND.n1052 9.3005
R12299 GND.n7355 GND.n1051 9.3005
R12300 GND.n1050 GND.n1046 9.3005
R12301 GND.n7361 GND.n1045 9.3005
R12302 GND.n7362 GND.n1044 9.3005
R12303 GND.n7363 GND.n1043 9.3005
R12304 GND.n1042 GND.n1038 9.3005
R12305 GND.n7369 GND.n1037 9.3005
R12306 GND.n7371 GND.n7370 9.3005
R12307 GND.n7226 GND.n7225 9.3005
R12308 GND.n6856 GND.n2667 9.3005
R12309 GND.n6855 GND.n6854 9.3005
R12310 GND.n6853 GND.n2669 9.3005
R12311 GND.n6852 GND.n6851 9.3005
R12312 GND.n6850 GND.n2673 9.3005
R12313 GND.n6849 GND.n6848 9.3005
R12314 GND.n6847 GND.n2674 9.3005
R12315 GND.n6846 GND.n6845 9.3005
R12316 GND.n6844 GND.n2678 9.3005
R12317 GND.n6843 GND.n6842 9.3005
R12318 GND.n6841 GND.n2679 9.3005
R12319 GND.n6840 GND.n6839 9.3005
R12320 GND.n6838 GND.n2683 9.3005
R12321 GND.n6837 GND.n6836 9.3005
R12322 GND.n6835 GND.n2684 9.3005
R12323 GND.n6834 GND.n6833 9.3005
R12324 GND.n6832 GND.n2688 9.3005
R12325 GND.n6831 GND.n6830 9.3005
R12326 GND.n6829 GND.n2689 9.3005
R12327 GND.n6828 GND.n6827 9.3005
R12328 GND.n6826 GND.n2693 9.3005
R12329 GND.n6825 GND.n6824 9.3005
R12330 GND.n6823 GND.n2694 9.3005
R12331 GND.n6822 GND.n6821 9.3005
R12332 GND.n6820 GND.n2698 9.3005
R12333 GND.n6819 GND.n6818 9.3005
R12334 GND.n6817 GND.n2699 9.3005
R12335 GND.n6816 GND.n6815 9.3005
R12336 GND.n6814 GND.n2703 9.3005
R12337 GND.n6813 GND.n6812 9.3005
R12338 GND.n6811 GND.n2704 9.3005
R12339 GND.n6810 GND.n6809 9.3005
R12340 GND.n6808 GND.n2708 9.3005
R12341 GND.n6807 GND.n6806 9.3005
R12342 GND.n6805 GND.n2709 9.3005
R12343 GND.n6804 GND.n6803 9.3005
R12344 GND.n6802 GND.n2713 9.3005
R12345 GND.n6801 GND.n6800 9.3005
R12346 GND.n6799 GND.n2714 9.3005
R12347 GND.n6798 GND.n6797 9.3005
R12348 GND.n6796 GND.n2718 9.3005
R12349 GND.n6795 GND.n6794 9.3005
R12350 GND.n6793 GND.n2719 9.3005
R12351 GND.n6792 GND.n6791 9.3005
R12352 GND.n6790 GND.n2723 9.3005
R12353 GND.n6789 GND.n6788 9.3005
R12354 GND.n6787 GND.n2724 9.3005
R12355 GND.n6786 GND.n6785 9.3005
R12356 GND.n6784 GND.n2728 9.3005
R12357 GND.n6783 GND.n6782 9.3005
R12358 GND.n6781 GND.n2729 9.3005
R12359 GND.n6780 GND.n6779 9.3005
R12360 GND.n6778 GND.n2733 9.3005
R12361 GND.n6777 GND.n6776 9.3005
R12362 GND.n6775 GND.n2734 9.3005
R12363 GND.n6774 GND.n6773 9.3005
R12364 GND.n6772 GND.n2738 9.3005
R12365 GND.n6771 GND.n6770 9.3005
R12366 GND.n6769 GND.n2739 9.3005
R12367 GND.n6768 GND.n6767 9.3005
R12368 GND.n6766 GND.n2743 9.3005
R12369 GND.n6765 GND.n6764 9.3005
R12370 GND.n6763 GND.n2744 9.3005
R12371 GND.n6762 GND.n6761 9.3005
R12372 GND.n6760 GND.n2748 9.3005
R12373 GND.n6759 GND.n6758 9.3005
R12374 GND.n6757 GND.n2749 9.3005
R12375 GND.n6756 GND.n6755 9.3005
R12376 GND.n6754 GND.n2753 9.3005
R12377 GND.n6753 GND.n6752 9.3005
R12378 GND.n6751 GND.n2754 9.3005
R12379 GND.n6750 GND.n6749 9.3005
R12380 GND.n6748 GND.n2758 9.3005
R12381 GND.n6747 GND.n6746 9.3005
R12382 GND.n6745 GND.n2759 9.3005
R12383 GND.n6744 GND.n6743 9.3005
R12384 GND.n6742 GND.n2763 9.3005
R12385 GND.n6741 GND.n6740 9.3005
R12386 GND.n6739 GND.n2764 9.3005
R12387 GND.n6738 GND.n6737 9.3005
R12388 GND.n6736 GND.n2768 9.3005
R12389 GND.n6735 GND.n6734 9.3005
R12390 GND.n6733 GND.n2769 9.3005
R12391 GND.n6732 GND.n6731 9.3005
R12392 GND.n6730 GND.n2773 9.3005
R12393 GND.n6729 GND.n6728 9.3005
R12394 GND.n6727 GND.n2774 9.3005
R12395 GND.n6726 GND.n6725 9.3005
R12396 GND.n6724 GND.n2778 9.3005
R12397 GND.n6723 GND.n6722 9.3005
R12398 GND.n6721 GND.n2779 9.3005
R12399 GND.n6720 GND.n6719 9.3005
R12400 GND.n6718 GND.n2783 9.3005
R12401 GND.n6717 GND.n6716 9.3005
R12402 GND.n6715 GND.n2784 9.3005
R12403 GND.n6714 GND.n6713 9.3005
R12404 GND.n6712 GND.n2788 9.3005
R12405 GND.n6711 GND.n6710 9.3005
R12406 GND.n6709 GND.n2789 9.3005
R12407 GND.n6708 GND.n6707 9.3005
R12408 GND.n6706 GND.n2793 9.3005
R12409 GND.n6705 GND.n6704 9.3005
R12410 GND.n6703 GND.n2794 9.3005
R12411 GND.n6702 GND.n6701 9.3005
R12412 GND.n6700 GND.n2798 9.3005
R12413 GND.n6699 GND.n6698 9.3005
R12414 GND.n6697 GND.n2799 9.3005
R12415 GND.n6696 GND.n6695 9.3005
R12416 GND.n6694 GND.n2803 9.3005
R12417 GND.n6693 GND.n6692 9.3005
R12418 GND.n6691 GND.n2804 9.3005
R12419 GND.n6690 GND.n6689 9.3005
R12420 GND.n6688 GND.n2808 9.3005
R12421 GND.n6687 GND.n6686 9.3005
R12422 GND.n6685 GND.n2809 9.3005
R12423 GND.n6684 GND.n6683 9.3005
R12424 GND.n6682 GND.n2813 9.3005
R12425 GND.n6681 GND.n6680 9.3005
R12426 GND.n6679 GND.n2814 9.3005
R12427 GND.n6678 GND.n6677 9.3005
R12428 GND.n6676 GND.n2818 9.3005
R12429 GND.n6675 GND.n6674 9.3005
R12430 GND.n6673 GND.n2819 9.3005
R12431 GND.n6672 GND.n6671 9.3005
R12432 GND.n6670 GND.n2823 9.3005
R12433 GND.n6669 GND.n6668 9.3005
R12434 GND.n6667 GND.n2824 9.3005
R12435 GND.n6666 GND.n6665 9.3005
R12436 GND.n6858 GND.n6857 9.3005
R12437 GND.n6662 GND.n2828 9.3005
R12438 GND.n6661 GND.n6660 9.3005
R12439 GND.n6659 GND.n2832 9.3005
R12440 GND.n6658 GND.n6657 9.3005
R12441 GND.n6656 GND.n2873 9.3005
R12442 GND.n6655 GND.n6654 9.3005
R12443 GND.n6653 GND.n2877 9.3005
R12444 GND.n6652 GND.n6651 9.3005
R12445 GND.n6650 GND.n2878 9.3005
R12446 GND.n6649 GND.n6648 9.3005
R12447 GND.n6647 GND.n2882 9.3005
R12448 GND.n6646 GND.n6645 9.3005
R12449 GND.n6644 GND.n2883 9.3005
R12450 GND.n6643 GND.n6642 9.3005
R12451 GND.n6641 GND.n2887 9.3005
R12452 GND.n6640 GND.n6639 9.3005
R12453 GND.n6638 GND.n2888 9.3005
R12454 GND.n6637 GND.n6636 9.3005
R12455 GND.n6635 GND.n6634 9.3005
R12456 GND.n6633 GND.n2895 9.3005
R12457 GND.n6632 GND.n6631 9.3005
R12458 GND.n6630 GND.n2899 9.3005
R12459 GND.n6664 GND.n6663 9.3005
R12460 GND.n4337 GND.n4336 9.3005
R12461 GND.n4335 GND.n3901 9.3005
R12462 GND.n4334 GND.n4333 9.3005
R12463 GND.n4332 GND.n4323 9.3005
R12464 GND.n4331 GND.n4330 9.3005
R12465 GND.n4329 GND.n4328 9.3005
R12466 GND.n3858 GND.n3857 9.3005
R12467 GND.n4420 GND.n4419 9.3005
R12468 GND.n4421 GND.n3855 9.3005
R12469 GND.n4433 GND.n4432 9.3005
R12470 GND.n4431 GND.n3856 9.3005
R12471 GND.n4430 GND.n4429 9.3005
R12472 GND.n4428 GND.n4422 9.3005
R12473 GND.n4427 GND.n4426 9.3005
R12474 GND.n3818 GND.n3817 9.3005
R12475 GND.n4497 GND.n4496 9.3005
R12476 GND.n4498 GND.n3815 9.3005
R12477 GND.n4510 GND.n4509 9.3005
R12478 GND.n4508 GND.n3816 9.3005
R12479 GND.n4507 GND.n4506 9.3005
R12480 GND.n4505 GND.n4499 9.3005
R12481 GND.n4504 GND.n4503 9.3005
R12482 GND.n3776 GND.n3775 9.3005
R12483 GND.n4591 GND.n4590 9.3005
R12484 GND.n4592 GND.n3773 9.3005
R12485 GND.n4595 GND.n4594 9.3005
R12486 GND.n4593 GND.n3774 9.3005
R12487 GND.n3746 GND.n3745 9.3005
R12488 GND.n4630 GND.n4629 9.3005
R12489 GND.n4631 GND.n3743 9.3005
R12490 GND.n4668 GND.n4667 9.3005
R12491 GND.n4666 GND.n3744 9.3005
R12492 GND.n4665 GND.n4664 9.3005
R12493 GND.n4663 GND.n4632 9.3005
R12494 GND.n4662 GND.n4661 9.3005
R12495 GND.n4660 GND.n4636 9.3005
R12496 GND.n4659 GND.n4658 9.3005
R12497 GND.n4657 GND.n4637 9.3005
R12498 GND.n4656 GND.n4655 9.3005
R12499 GND.n4654 GND.n4640 9.3005
R12500 GND.n4653 GND.n4652 9.3005
R12501 GND.n4651 GND.n4641 9.3005
R12502 GND.n4650 GND.n4649 9.3005
R12503 GND.n4648 GND.n4647 9.3005
R12504 GND.n3658 GND.n3657 9.3005
R12505 GND.n4806 GND.n4805 9.3005
R12506 GND.n4807 GND.n3655 9.3005
R12507 GND.n4844 GND.n4843 9.3005
R12508 GND.n4842 GND.n3656 9.3005
R12509 GND.n4841 GND.n4840 9.3005
R12510 GND.n4839 GND.n4808 9.3005
R12511 GND.n4838 GND.n4837 9.3005
R12512 GND.n4836 GND.n4812 9.3005
R12513 GND.n4835 GND.n4834 9.3005
R12514 GND.n4833 GND.n4813 9.3005
R12515 GND.n4832 GND.n4831 9.3005
R12516 GND.n4830 GND.n4816 9.3005
R12517 GND.n4829 GND.n4828 9.3005
R12518 GND.n4827 GND.n4817 9.3005
R12519 GND.n4826 GND.n4825 9.3005
R12520 GND.n4824 GND.n4823 9.3005
R12521 GND.n3570 GND.n3569 9.3005
R12522 GND.n4982 GND.n4981 9.3005
R12523 GND.n4983 GND.n3567 9.3005
R12524 GND.n5020 GND.n5019 9.3005
R12525 GND.n5018 GND.n3568 9.3005
R12526 GND.n5017 GND.n5016 9.3005
R12527 GND.n5015 GND.n4984 9.3005
R12528 GND.n5014 GND.n5013 9.3005
R12529 GND.n5012 GND.n4988 9.3005
R12530 GND.n5011 GND.n5010 9.3005
R12531 GND.n5009 GND.n4989 9.3005
R12532 GND.n5008 GND.n5007 9.3005
R12533 GND.n5006 GND.n4992 9.3005
R12534 GND.n5005 GND.n5004 9.3005
R12535 GND.n5003 GND.n4993 9.3005
R12536 GND.n5002 GND.n5001 9.3005
R12537 GND.n5000 GND.n4999 9.3005
R12538 GND.n3481 GND.n3480 9.3005
R12539 GND.n5158 GND.n5157 9.3005
R12540 GND.n5159 GND.n3478 9.3005
R12541 GND.n5196 GND.n5195 9.3005
R12542 GND.n5194 GND.n3479 9.3005
R12543 GND.n5193 GND.n5192 9.3005
R12544 GND.n5191 GND.n5160 9.3005
R12545 GND.n5190 GND.n5189 9.3005
R12546 GND.n5188 GND.n5164 9.3005
R12547 GND.n5187 GND.n5186 9.3005
R12548 GND.n5185 GND.n5165 9.3005
R12549 GND.n5184 GND.n5183 9.3005
R12550 GND.n5182 GND.n5168 9.3005
R12551 GND.n5181 GND.n5180 9.3005
R12552 GND.n5179 GND.n5169 9.3005
R12553 GND.n5178 GND.n5177 9.3005
R12554 GND.n5176 GND.n5175 9.3005
R12555 GND.n3392 GND.n3391 9.3005
R12556 GND.n5333 GND.n5332 9.3005
R12557 GND.n5334 GND.n3389 9.3005
R12558 GND.n5373 GND.n5372 9.3005
R12559 GND.n5371 GND.n3390 9.3005
R12560 GND.n5370 GND.n5369 9.3005
R12561 GND.n5368 GND.n5335 9.3005
R12562 GND.n5367 GND.n5366 9.3005
R12563 GND.n5365 GND.n5341 9.3005
R12564 GND.n5364 GND.n5363 9.3005
R12565 GND.n5362 GND.n5342 9.3005
R12566 GND.n5361 GND.n5360 9.3005
R12567 GND.n5359 GND.n5345 9.3005
R12568 GND.n5358 GND.n5357 9.3005
R12569 GND.n5356 GND.n5346 9.3005
R12570 GND.n5355 GND.n5354 9.3005
R12571 GND.n5353 GND.n5352 9.3005
R12572 GND.n3306 GND.n3305 9.3005
R12573 GND.n5511 GND.n5510 9.3005
R12574 GND.n5512 GND.n3303 9.3005
R12575 GND.n5526 GND.n5525 9.3005
R12576 GND.n5524 GND.n3304 9.3005
R12577 GND.n5523 GND.n5522 9.3005
R12578 GND.n5521 GND.n5513 9.3005
R12579 GND.n5520 GND.n5519 9.3005
R12580 GND.n5518 GND.n5517 9.3005
R12581 GND.n3256 GND.n3255 9.3005
R12582 GND.n5605 GND.n5604 9.3005
R12583 GND.n5606 GND.n3253 9.3005
R12584 GND.n5609 GND.n5608 9.3005
R12585 GND.n5607 GND.n3254 9.3005
R12586 GND.n2901 GND.n2900 9.3005
R12587 GND.n6629 GND.n6628 9.3005
R12588 GND.n4322 GND.n3900 9.3005
R12589 GND.n3903 GND.n3902 9.3005
R12590 GND.n4245 GND.n4238 9.3005
R12591 GND.n4247 GND.n4246 9.3005
R12592 GND.n4248 GND.n4237 9.3005
R12593 GND.n4250 GND.n4249 9.3005
R12594 GND.n4251 GND.n4232 9.3005
R12595 GND.n4253 GND.n4252 9.3005
R12596 GND.n4254 GND.n4231 9.3005
R12597 GND.n4256 GND.n4255 9.3005
R12598 GND.n4257 GND.n4226 9.3005
R12599 GND.n4259 GND.n4258 9.3005
R12600 GND.n4260 GND.n4225 9.3005
R12601 GND.n4262 GND.n4261 9.3005
R12602 GND.n4263 GND.n4220 9.3005
R12603 GND.n4265 GND.n4264 9.3005
R12604 GND.n4266 GND.n4219 9.3005
R12605 GND.n4268 GND.n4267 9.3005
R12606 GND.n4269 GND.n4215 9.3005
R12607 GND.n4271 GND.n4270 9.3005
R12608 GND.n4272 GND.n4214 9.3005
R12609 GND.n4314 GND.n4313 9.3005
R12610 GND.n4213 GND.n2668 9.3005
R12611 GND.n4321 GND.n4320 9.3005
R12612 GND.n6991 GND.n6990 9.3005
R12613 GND.n7022 GND.n7021 9.3005
R12614 GND.n7023 GND.n1403 9.3005
R12615 GND.n7025 GND.n7024 9.3005
R12616 GND.n7026 GND.n1397 9.3005
R12617 GND.n7028 GND.n7027 9.3005
R12618 GND.n7029 GND.n1396 9.3005
R12619 GND.n7031 GND.n7030 9.3005
R12620 GND.n7032 GND.n1392 9.3005
R12621 GND.n7034 GND.n7033 9.3005
R12622 GND.n7035 GND.n1391 9.3005
R12623 GND.n7037 GND.n7036 9.3005
R12624 GND.n7038 GND.n1388 9.3005
R12625 GND.n7040 GND.n7039 9.3005
R12626 GND.n7019 GND.n7018 9.3005
R12627 GND.n7017 GND.n1409 9.3005
R12628 GND.n7016 GND.n7015 9.3005
R12629 GND.n7014 GND.n1410 9.3005
R12630 GND.n7013 GND.n7012 9.3005
R12631 GND.n7011 GND.n1416 9.3005
R12632 GND.n7010 GND.n7009 9.3005
R12633 GND.n7008 GND.n1417 9.3005
R12634 GND.n7007 GND.n7006 9.3005
R12635 GND.n7005 GND.n1421 9.3005
R12636 GND.n7004 GND.n7003 9.3005
R12637 GND.n7002 GND.n1422 9.3005
R12638 GND.n7001 GND.n7000 9.3005
R12639 GND.n6999 GND.n1426 9.3005
R12640 GND.n6998 GND.n6997 9.3005
R12641 GND.n6996 GND.n1427 9.3005
R12642 GND.n6995 GND.n1432 9.3005
R12643 GND.n6994 GND.n6993 9.3005
R12644 GND.n7109 GND.n1295 9.3005
R12645 GND.n2153 GND.n1296 9.3005
R12646 GND.n7105 GND.n1300 9.3005
R12647 GND.n7104 GND.n1301 9.3005
R12648 GND.n7103 GND.n1302 9.3005
R12649 GND.n2132 GND.n1303 9.3005
R12650 GND.n7099 GND.n1308 9.3005
R12651 GND.n7098 GND.n1309 9.3005
R12652 GND.n7097 GND.n1310 9.3005
R12653 GND.n2119 GND.n1311 9.3005
R12654 GND.n7093 GND.n1316 9.3005
R12655 GND.n7092 GND.n1317 9.3005
R12656 GND.n7091 GND.n1318 9.3005
R12657 GND.n2314 GND.n1319 9.3005
R12658 GND.n7087 GND.n1324 9.3005
R12659 GND.n7086 GND.n1325 9.3005
R12660 GND.n7085 GND.n1326 9.3005
R12661 GND.n2062 GND.n1327 9.3005
R12662 GND.n7081 GND.n1332 9.3005
R12663 GND.n7080 GND.n1333 9.3005
R12664 GND.n7079 GND.n1334 9.3005
R12665 GND.n2395 GND.n1335 9.3005
R12666 GND.n7075 GND.n1340 9.3005
R12667 GND.n7074 GND.n1341 9.3005
R12668 GND.n7073 GND.n1342 9.3005
R12669 GND.n2041 GND.n1343 9.3005
R12670 GND.n7069 GND.n1348 9.3005
R12671 GND.n7068 GND.n1349 9.3005
R12672 GND.n7067 GND.n1350 9.3005
R12673 GND.n2435 GND.n1351 9.3005
R12674 GND.n7063 GND.n1356 9.3005
R12675 GND.n7062 GND.n1357 9.3005
R12676 GND.n7061 GND.n1358 9.3005
R12677 GND.n2466 GND.n1359 9.3005
R12678 GND.n7057 GND.n1364 9.3005
R12679 GND.n7056 GND.n1365 9.3005
R12680 GND.n7055 GND.n1366 9.3005
R12681 GND.n2499 GND.n1367 9.3005
R12682 GND.n7051 GND.n1372 9.3005
R12683 GND.n7050 GND.n1373 9.3005
R12684 GND.n7049 GND.n1374 9.3005
R12685 GND.n2515 GND.n1375 9.3005
R12686 GND.n2514 GND.n1378 9.3005
R12687 GND.n7111 GND.n7110 9.3005
R12688 GND.n7109 GND.n7108 9.3005
R12689 GND.n7107 GND.n1296 9.3005
R12690 GND.n7106 GND.n7105 9.3005
R12691 GND.n7104 GND.n1299 9.3005
R12692 GND.n7103 GND.n7102 9.3005
R12693 GND.n7101 GND.n1303 9.3005
R12694 GND.n7100 GND.n7099 9.3005
R12695 GND.n7098 GND.n1307 9.3005
R12696 GND.n7097 GND.n7096 9.3005
R12697 GND.n7095 GND.n1311 9.3005
R12698 GND.n7094 GND.n7093 9.3005
R12699 GND.n7092 GND.n1315 9.3005
R12700 GND.n7091 GND.n7090 9.3005
R12701 GND.n7089 GND.n1319 9.3005
R12702 GND.n7088 GND.n7087 9.3005
R12703 GND.n7086 GND.n1323 9.3005
R12704 GND.n7085 GND.n7084 9.3005
R12705 GND.n7083 GND.n1327 9.3005
R12706 GND.n7082 GND.n7081 9.3005
R12707 GND.n7080 GND.n1331 9.3005
R12708 GND.n7079 GND.n7078 9.3005
R12709 GND.n7077 GND.n1335 9.3005
R12710 GND.n7076 GND.n7075 9.3005
R12711 GND.n7074 GND.n1339 9.3005
R12712 GND.n7073 GND.n7072 9.3005
R12713 GND.n7071 GND.n1343 9.3005
R12714 GND.n7070 GND.n7069 9.3005
R12715 GND.n7068 GND.n1347 9.3005
R12716 GND.n7067 GND.n7066 9.3005
R12717 GND.n7065 GND.n1351 9.3005
R12718 GND.n7064 GND.n7063 9.3005
R12719 GND.n7062 GND.n1355 9.3005
R12720 GND.n7061 GND.n7060 9.3005
R12721 GND.n7059 GND.n1359 9.3005
R12722 GND.n7058 GND.n7057 9.3005
R12723 GND.n7056 GND.n1363 9.3005
R12724 GND.n7055 GND.n7054 9.3005
R12725 GND.n7053 GND.n1367 9.3005
R12726 GND.n7052 GND.n7051 9.3005
R12727 GND.n7050 GND.n1371 9.3005
R12728 GND.n7049 GND.n7048 9.3005
R12729 GND.n7047 GND.n1375 9.3005
R12730 GND.n7046 GND.n1378 9.3005
R12731 GND.n7110 GND.n1289 9.3005
R12732 GND.n2207 GND.n2177 9.3005
R12733 GND.n2206 GND.n2205 9.3005
R12734 GND.n2204 GND.n2181 9.3005
R12735 GND.n2203 GND.n2202 9.3005
R12736 GND.n2199 GND.n2184 9.3005
R12737 GND.n2198 GND.n2197 9.3005
R12738 GND.n2196 GND.n2185 9.3005
R12739 GND.n2195 GND.n2194 9.3005
R12740 GND.n2191 GND.n2188 9.3005
R12741 GND.n2190 GND.n2189 9.3005
R12742 GND.n2209 GND.n2208 9.3005
R12743 GND.n2212 GND.n2175 9.3005
R12744 GND.n2215 GND.n2214 9.3005
R12745 GND.n2213 GND.n2176 9.3005
R12746 GND.n2139 GND.n2138 9.3005
R12747 GND.n2282 GND.n2281 9.3005
R12748 GND.n2283 GND.n2136 9.3005
R12749 GND.n2286 GND.n2285 9.3005
R12750 GND.n2284 GND.n2137 9.3005
R12751 GND.n2115 GND.n2114 9.3005
R12752 GND.n2306 GND.n2305 9.3005
R12753 GND.n2307 GND.n2112 9.3005
R12754 GND.n2310 GND.n2309 9.3005
R12755 GND.n2308 GND.n2113 9.3005
R12756 GND.n2092 GND.n2091 9.3005
R12757 GND.n2329 GND.n2328 9.3005
R12758 GND.n2330 GND.n2090 9.3005
R12759 GND.n2332 GND.n2331 9.3005
R12760 GND.n2333 GND.n2089 9.3005
R12761 GND.n2337 GND.n2336 9.3005
R12762 GND.n2338 GND.n2088 9.3005
R12763 GND.n2340 GND.n2339 9.3005
R12764 GND.n2211 GND.n2210 9.3005
R12765 GND.n7179 GND.n1243 9.26784
R12766 GND.t194 GND.n2548 9.26784
R12767 GND.n4436 GND.n4435 9.26784
R12768 GND.n4494 GND.n3820 9.26784
R12769 GND.n4551 GND.n3763 9.26784
R12770 GND.n4537 GND.n3724 9.26784
R12771 GND.n4768 GND.n3676 9.26784
R12772 GND.n4754 GND.n3636 9.26784
R12773 GND.n4945 GND.n3589 9.26784
R12774 GND.n4931 GND.n3548 9.26784
R12775 GND.n5121 GND.n3500 9.26784
R12776 GND.n5106 GND.n3458 9.26784
R12777 GND.n5295 GND.n3410 9.26784
R12778 GND.n5281 GND.n3372 9.26784
R12779 GND.n5473 GND.n3324 9.26784
R12780 GND.n5459 GND.n3284 9.26784
R12781 GND.n383 GND.n253 9.26784
R12782 GND.n1774 GND.t222 9.22596
R12783 GND.n1793 GND.t225 9.22596
R12784 GND.n1813 GND.t230 9.22596
R12785 GND.n1832 GND.t218 9.22596
R12786 GND.n1713 GND.t228 9.22596
R12787 GND.n1732 GND.t226 9.22596
R12788 GND.n1752 GND.t233 9.22596
R12789 GND.n1771 GND.t227 9.22596
R12790 GND.n1652 GND.t236 9.22596
R12791 GND.n1671 GND.t238 9.22596
R12792 GND.n1691 GND.t229 9.22596
R12793 GND.n1710 GND.t215 9.22596
R12794 GND.n1591 GND.t239 9.22596
R12795 GND.n1610 GND.t231 9.22596
R12796 GND.n1630 GND.t232 9.22596
R12797 GND.n1649 GND.t223 9.22596
R12798 GND.n1561 GND.t141 9.22596
R12799 GND.n1542 GND.t133 9.22596
R12800 GND.n1583 GND.t92 9.22596
R12801 GND.n1564 GND.t131 9.22596
R12802 GND.n1855 GND.t178 9.22596
R12803 GND.n1836 GND.t96 9.22596
R12804 GND.n1585 GND.t94 9.22596
R12805 GND.n1444 GND.t161 9.22596
R12806 GND.n25 GND.n15 8.92171
R12807 GND.n40 GND.n30 8.92171
R12808 GND.n56 GND.n46 8.92171
R12809 GND.n10 GND.n0 8.92171
R12810 GND.n1899 GND.n1888 8.92171
R12811 GND.n4292 GND.n4281 8.92171
R12812 GND.n2852 GND.n2841 8.92171
R12813 GND.n86 GND.n76 8.92171
R12814 GND.n101 GND.n91 8.92171
R12815 GND.n117 GND.n107 8.92171
R12816 GND.n133 GND.n123 8.92171
R12817 GND.n6085 GND.n6074 8.92171
R12818 GND.n7027 GND.n7026 8.72777
R12819 GND.n6496 GND.n6493 8.72777
R12820 GND.n365 GND.n362 8.72777
R12821 GND.n7163 GND.n7160 8.72777
R12822 GND.n4121 GND.n4118 8.60589
R12823 GND.n6917 GND.n6916 8.60589
R12824 GND.n6889 GND.n2627 8.60589
R12825 GND.n4340 GND.n3898 8.60589
R12826 GND.n4416 GND.n3862 8.60589
R12827 GND.t16 GND.n3841 8.60589
R12828 GND.n4513 GND.n3812 8.60589
R12829 GND.n4600 GND.n4599 8.60589
R12830 GND.n4695 GND.n3717 8.60589
R12831 GND.n4776 GND.n4775 8.60589
R12832 GND.n4872 GND.n3630 8.60589
R12833 GND.n4953 GND.n4952 8.60589
R12834 GND.n5048 GND.n3541 8.60589
R12835 GND.n5129 GND.n5128 8.60589
R12836 GND.n5223 GND.n3452 8.60589
R12837 GND.n5303 GND.n5302 8.60589
R12838 GND.n5400 GND.n3365 8.60589
R12839 GND.n5481 GND.n5480 8.60589
R12840 GND.n5528 GND.t33 8.60589
R12841 GND.n5556 GND.n3278 8.60589
R12842 GND.n5630 GND.n5629 8.60589
R12843 GND.n6597 GND.n2941 8.60589
R12844 GND.n6570 GND.n6569 8.60589
R12845 GND.n8513 GND.n8512 8.60581
R12846 GND.n2087 GND.n63 8.60581
R12847 GND.n1590 GND.n1589 8.25845
R12848 GND.n1834 GND.n1833 8.25845
R12849 GND.n1914 GND.n1880 8.2187
R12850 GND.n4307 GND.n4273 8.2187
R12851 GND.n2867 GND.n2833 8.2187
R12852 GND.n6100 GND.n6066 8.2187
R12853 GND.n23 GND.n22 8.14595
R12854 GND.n38 GND.n37 8.14595
R12855 GND.n54 GND.n53 8.14595
R12856 GND.n8 GND.n7 8.14595
R12857 GND.n1896 GND.n1895 8.14595
R12858 GND.n4289 GND.n4288 8.14595
R12859 GND.n2849 GND.n2848 8.14595
R12860 GND.n84 GND.n83 8.14595
R12861 GND.n99 GND.n98 8.14595
R12862 GND.n115 GND.n114 8.14595
R12863 GND.n131 GND.n130 8.14595
R12864 GND.n6082 GND.n6081 8.14595
R12865 GND.n6987 GND.n1924 7.94393
R12866 GND.n6868 GND.t8 7.94393
R12867 GND.n4340 GND.n4339 7.94393
R12868 GND.n4417 GND.n4416 7.94393
R12869 GND.n4513 GND.n4512 7.94393
R12870 GND.n4600 GND.n3768 7.94393
R12871 GND.n4695 GND.n3718 7.94393
R12872 GND.n4776 GND.n3680 7.94393
R12873 GND.n4872 GND.n3631 7.94393
R12874 GND.n4902 GND.t43 7.94393
R12875 GND.n4953 GND.n3593 7.94393
R12876 GND.n5048 GND.n3543 7.94393
R12877 GND.t4 GND.n5075 7.94393
R12878 GND.n5129 GND.n3504 7.94393
R12879 GND.n5223 GND.n3453 7.94393
R12880 GND.n5303 GND.n3415 7.94393
R12881 GND.n5400 GND.n3366 7.94393
R12882 GND.n5481 GND.n3328 7.94393
R12883 GND.n5556 GND.n3279 7.94393
R12884 GND.n5630 GND.n3239 7.94393
R12885 GND.n6618 GND.t22 7.94393
R12886 GND.n6512 GND.n3067 7.94393
R12887 GND.n6064 GND.n6059 7.43975
R12888 GND.n19 GND.n17 7.3702
R12889 GND.n34 GND.n32 7.3702
R12890 GND.n50 GND.n48 7.3702
R12891 GND.n4 GND.n2 7.3702
R12892 GND.n1892 GND.n1890 7.3702
R12893 GND.n4285 GND.n4283 7.3702
R12894 GND.n2845 GND.n2843 7.3702
R12895 GND.n80 GND.n78 7.3702
R12896 GND.n95 GND.n93 7.3702
R12897 GND.n111 GND.n109 7.3702
R12898 GND.n127 GND.n125 7.3702
R12899 GND.n6078 GND.n6076 7.3702
R12900 GND.n26 GND.t27 7.30677
R12901 GND.n26 GND.t68 7.30677
R12902 GND.n28 GND.t24 7.30677
R12903 GND.n28 GND.t63 7.30677
R12904 GND.n41 GND.t74 7.30677
R12905 GND.n41 GND.t67 7.30677
R12906 GND.n43 GND.t11 7.30677
R12907 GND.n43 GND.t76 7.30677
R12908 GND.n57 GND.t13 7.30677
R12909 GND.n57 GND.t46 7.30677
R12910 GND.n59 GND.t47 7.30677
R12911 GND.n59 GND.t66 7.30677
R12912 GND.n11 GND.t212 7.30677
R12913 GND.n11 GND.t77 7.30677
R12914 GND.n13 GND.t207 7.30677
R12915 GND.n13 GND.t75 7.30677
R12916 GND.n74 GND.t25 7.30677
R12917 GND.n74 GND.t29 7.30677
R12918 GND.n73 GND.t203 7.30677
R12919 GND.n73 GND.t73 7.30677
R12920 GND.n89 GND.t1 7.30677
R12921 GND.n89 GND.t72 7.30677
R12922 GND.n88 GND.t69 7.30677
R12923 GND.n88 GND.t65 7.30677
R12924 GND.n105 GND.t26 7.30677
R12925 GND.n105 GND.t41 7.30677
R12926 GND.n104 GND.t15 7.30677
R12927 GND.n104 GND.t202 7.30677
R12928 GND.n121 GND.t210 7.30677
R12929 GND.n121 GND.t30 7.30677
R12930 GND.n120 GND.t205 7.30677
R12931 GND.n120 GND.t70 7.30677
R12932 GND.t39 GND.n2011 7.28198
R12933 GND.n2564 GND.n2558 7.28198
R12934 GND.n6923 GND.n2583 7.28198
R12935 GND.n6882 GND.n6881 7.28198
R12936 GND.n4211 GND.n4210 7.28198
R12937 GND.n4435 GND.n3846 7.28198
R12938 GND.n4551 GND.n3754 7.28198
R12939 GND.n4537 GND.n3736 7.28198
R12940 GND.n4768 GND.n3666 7.28198
R12941 GND.n4754 GND.n3648 7.28198
R12942 GND.n4945 GND.n3578 7.28198
R12943 GND.n4931 GND.n3560 7.28198
R12944 GND.n5121 GND.n3489 7.28198
R12945 GND.n5106 GND.n3471 7.28198
R12946 GND.n5295 GND.n3400 7.28198
R12947 GND.n5281 GND.n3382 7.28198
R12948 GND.n5459 GND.n3296 7.28198
R12949 GND.n5637 GND.n3235 7.28198
R12950 GND.n6605 GND.n6604 7.28198
R12951 GND.n6563 GND.n2985 7.28198
R12952 GND.n3010 GND.n3004 7.28198
R12953 GND.t14 GND.n5881 7.28198
R12954 GND.n4379 GND.t190 6.951
R12955 GND.n4847 GND.t58 6.951
R12956 GND.t82 GND.n5154 6.951
R12957 GND.n5585 GND.t107 6.951
R12958 GND.n63 GND.n62 6.81087
R12959 GND.n8513 GND.n135 6.81087
R12960 GND.n3894 GND.n3885 6.62003
R12961 GND.n4372 GND.n3877 6.62003
R12962 GND.n3808 GND.n3797 6.62003
R12963 GND.n4561 GND.n3787 6.62003
R12964 GND.n4717 GND.n4716 6.62003
R12965 GND.n4731 GND.n3693 6.62003
R12966 GND.n4894 GND.n4893 6.62003
R12967 GND.n4908 GND.n3606 6.62003
R12968 GND.n5069 GND.n5068 6.62003
R12969 GND.n5083 GND.n3517 6.62003
R12970 GND.n5244 GND.n5243 6.62003
R12971 GND.n5258 GND.n3430 6.62003
R12972 GND.n5422 GND.n5421 6.62003
R12973 GND.n5436 GND.n3341 6.62003
R12974 GND.n5595 GND.n5594 6.62003
R12975 GND.n5613 GND.n5611 6.62003
R12976 GND.n3027 GND.t118 6.62003
R12977 GND.n5728 GND.t173 6.62003
R12978 GND.n45 GND.n29 6.48757
R12979 GND.n1794 GND.n1793 6.36192
R12980 GND.n1813 GND.n1812 6.36192
R12981 GND.n1733 GND.n1732 6.36192
R12982 GND.n1752 GND.n1751 6.36192
R12983 GND.n1672 GND.n1671 6.36192
R12984 GND.n1691 GND.n1690 6.36192
R12985 GND.n1611 GND.n1610 6.36192
R12986 GND.n1630 GND.n1629 6.36192
R12987 GND.n6064 GND.n6063 6.26037
R12988 GND.t10 GND.n2118 5.95807
R12989 GND.n4134 GND.n4131 5.95807
R12990 GND.n6931 GND.n6930 5.95807
R12991 GND.n6875 GND.n2645 5.95807
R12992 GND.n4192 GND.n2647 5.95807
R12993 GND.n4469 GND.n4468 5.95807
R12994 GND.n4476 GND.n4475 5.95807
R12995 GND.n4625 GND.n3750 5.95807
R12996 GND.n4671 GND.n3740 5.95807
R12997 GND.n4802 GND.n3662 5.95807
R12998 GND.n4847 GND.n3652 5.95807
R12999 GND.n4978 GND.n3574 5.95807
R13000 GND.n5024 GND.n3564 5.95807
R13001 GND.n5154 GND.n3485 5.95807
R13002 GND.n5199 GND.n3475 5.95807
R13003 GND.n5328 GND.n3396 5.95807
R13004 GND.n5376 GND.n3386 5.95807
R13005 GND.n5507 GND.n3310 5.95807
R13006 GND.n5529 GND.n3300 5.95807
R13007 GND.n5642 GND.n2921 5.95807
R13008 GND.n6611 GND.n2923 5.95807
R13009 GND.n6556 GND.n6555 5.95807
R13010 GND.n5704 GND.n5701 5.95807
R13011 GND.n6534 GND.t118 5.95807
R13012 GND.n6354 GND.t52 5.95807
R13013 GND.n103 GND.n87 5.90567
R13014 GND.n22 GND.n17 5.81868
R13015 GND.n37 GND.n32 5.81868
R13016 GND.n53 GND.n48 5.81868
R13017 GND.n7 GND.n2 5.81868
R13018 GND.n1895 GND.n1890 5.81868
R13019 GND.n4288 GND.n4283 5.81868
R13020 GND.n2848 GND.n2843 5.81868
R13021 GND.n83 GND.n78 5.81868
R13022 GND.n98 GND.n93 5.81868
R13023 GND.n114 GND.n109 5.81868
R13024 GND.n130 GND.n125 5.81868
R13025 GND.n6081 GND.n6076 5.81868
R13026 GND.n4486 GND.t18 5.6271
R13027 GND.t6 GND.n3314 5.6271
R13028 GND.n1912 GND.n1880 5.3904
R13029 GND.n4305 GND.n4273 5.3904
R13030 GND.n2865 GND.n2833 5.3904
R13031 GND.n6098 GND.n6066 5.3904
R13032 GND.n62 GND.n14 5.35179
R13033 GND.n4380 GND.n3881 5.29612
R13034 GND.n4378 GND.n3875 5.29612
R13035 GND.n4569 GND.n3793 5.29612
R13036 GND.n4567 GND.n3785 5.29612
R13037 GND.n4723 GND.n3699 5.29612
R13038 GND.n4725 GND.n3691 5.29612
R13039 GND.n4900 GND.n3612 5.29612
R13040 GND.n4902 GND.n3603 5.29612
R13041 GND.n5075 GND.n3523 5.29612
R13042 GND.n5077 GND.n3515 5.29612
R13043 GND.n5250 GND.n3434 5.29612
R13044 GND.n5252 GND.n3425 5.29612
R13045 GND.n5428 GND.n3347 5.29612
R13046 GND.n5430 GND.n3339 5.29612
R13047 GND.n5602 GND.n5601 5.29612
R13048 GND.n5587 GND.n5586 5.29612
R13049 GND.n45 GND.n44 5.28929
R13050 GND.n61 GND.n60 5.28929
R13051 GND.n23 GND.n15 5.04292
R13052 GND.n38 GND.n30 5.04292
R13053 GND.n54 GND.n46 5.04292
R13054 GND.n8 GND.n0 5.04292
R13055 GND.n1896 GND.n1888 5.04292
R13056 GND.n4289 GND.n4281 5.04292
R13057 GND.n2849 GND.n2841 5.04292
R13058 GND.n84 GND.n76 5.04292
R13059 GND.n99 GND.n91 5.04292
R13060 GND.n115 GND.n107 5.04292
R13061 GND.n131 GND.n123 5.04292
R13062 GND.n6082 GND.n6074 5.04292
R13063 GND.n4716 GND.t2 4.96515
R13064 GND.n3430 GND.t208 4.96515
R13065 GND.n135 GND.n134 4.7699
R13066 GND.n1940 GND.n1436 4.74817
R13067 GND.n1941 GND.n1917 4.74817
R13068 GND.n1945 GND.n1918 4.74817
R13069 GND.n1949 GND.n1919 4.74817
R13070 GND.n6131 GND.n6107 4.74817
R13071 GND.n6127 GND.n6108 4.74817
R13072 GND.n6123 GND.n6109 4.74817
R13073 GND.n6119 GND.n6110 4.74817
R13074 GND.n6116 GND.n6110 4.74817
R13075 GND.n6120 GND.n6109 4.74817
R13076 GND.n6124 GND.n6108 4.74817
R13077 GND.n6128 GND.n6107 4.74817
R13078 GND.n5907 GND.n155 4.74817
R13079 GND.n153 GND.n147 4.74817
R13080 GND.n8505 GND.n148 4.74817
R13081 GND.n156 GND.n152 4.74817
R13082 GND.n6390 GND.n155 4.74817
R13083 GND.n5922 GND.n153 4.74817
R13084 GND.n8506 GND.n8505 4.74817
R13085 GND.n5942 GND.n152 4.74817
R13086 GND.n2243 GND.n2242 4.74817
R13087 GND.n2407 GND.n2406 4.74817
R13088 GND.n2356 GND.n2068 4.74817
R13089 GND.n2390 GND.n2358 4.74817
R13090 GND.n2388 GND.n2387 4.74817
R13091 GND.n6031 GND.n5929 4.74817
R13092 GND.n6384 GND.n6383 4.74817
R13093 GND.n5946 GND.n5930 4.74817
R13094 GND.n6369 GND.n6368 4.74817
R13095 GND.n6364 GND.n5947 4.74817
R13096 GND.n6032 GND.n6031 4.74817
R13097 GND.n6385 GND.n6384 4.74817
R13098 GND.n6382 GND.n5930 4.74817
R13099 GND.n6370 GND.n6369 4.74817
R13100 GND.n6367 GND.n5947 4.74817
R13101 GND.n2417 GND.n2416 4.74817
R13102 GND.n2400 GND.n2051 4.74817
R13103 GND.n2347 GND.n2050 4.74817
R13104 GND.n2049 GND.n2046 4.74817
R13105 GND.n2417 GND.n2053 4.74817
R13106 GND.n2077 GND.n2051 4.74817
R13107 GND.n2399 GND.n2050 4.74817
R13108 GND.n2348 GND.n2049 4.74817
R13109 GND.n2242 GND.n2067 4.74817
R13110 GND.n2408 GND.n2407 4.74817
R13111 GND.n2405 GND.n2068 4.74817
R13112 GND.n2358 GND.n2357 4.74817
R13113 GND.n2389 GND.n2388 4.74817
R13114 GND.n1944 GND.n1917 4.74817
R13115 GND.n1948 GND.n1918 4.74817
R13116 GND.n1952 GND.n1919 4.74817
R13117 GND.n103 GND.n102 4.7074
R13118 GND.n119 GND.n118 4.7074
R13119 GND.n6937 GND.n2566 4.63417
R13120 GND.n4139 GND.n2581 4.63417
R13121 GND.n4187 GND.n4184 4.63417
R13122 GND.n6868 GND.n6867 4.63417
R13123 GND.n4400 GND.n4399 4.63417
R13124 GND.n4461 GND.n4460 4.63417
R13125 GND.n4617 GND.n3748 4.63417
R13126 GND.n4679 GND.n3733 4.63417
R13127 GND.n4793 GND.n3660 4.63417
R13128 GND.n4856 GND.n3645 4.63417
R13129 GND.n4970 GND.n3572 4.63417
R13130 GND.n5032 GND.n3557 4.63417
R13131 GND.n5146 GND.n3483 4.63417
R13132 GND.n5207 GND.n3468 4.63417
R13133 GND.n5320 GND.n3394 4.63417
R13134 GND.n5384 GND.n3379 4.63417
R13135 GND.n5498 GND.n3308 4.63417
R13136 GND.n5538 GND.n3293 4.63417
R13137 GND.n6619 GND.n6618 4.63417
R13138 GND.n5651 GND.n5648 4.63417
R13139 GND.n5695 GND.n2987 4.63417
R13140 GND.n6549 GND.n3002 4.63417
R13141 GND.t156 GND.n5714 4.63417
R13142 GND.n6485 GND.n5792 4.6132
R13143 GND.n7020 GND.n1404 4.6132
R13144 GND.n72 GND.n67 4.4442
R13145 GND.t190 GND.n4378 4.30319
R13146 GND.n5601 GND.t107 4.30319
R13147 GND.n1900 GND.n1899 4.26717
R13148 GND.n4293 GND.n4292 4.26717
R13149 GND.n2853 GND.n2852 4.26717
R13150 GND.n6086 GND.n6085 4.26717
R13151 GND.n1712 GND.n1711 4.26641
R13152 GND.n2269 GND.t111 3.97222
R13153 GND.n2511 GND.t125 3.97222
R13154 GND.n4348 GND.n4347 3.97222
R13155 GND.n4410 GND.n4409 3.97222
R13156 GND.n4521 GND.n4520 3.97222
R13157 GND.n4588 GND.n3778 3.97222
R13158 GND.n4704 GND.n4703 3.97222
R13159 GND.n4882 GND.n4880 3.97222
R13160 GND.n4910 GND.n3597 3.97222
R13161 GND.n5057 GND.n5056 3.97222
R13162 GND.n5085 GND.n3508 3.97222
R13163 GND.n5260 GND.n3419 3.97222
R13164 GND.n5409 GND.n5408 3.97222
R13165 GND.n5438 GND.n3333 3.97222
R13166 GND.n5564 GND.n5562 3.97222
R13167 GND.n5621 GND.n3245 3.97222
R13168 GND.n5717 GND.t156 3.97222
R13169 GND.n6521 GND.t129 3.97222
R13170 GND.n6138 GND.t99 3.97222
R13171 GND.n8459 GND.t121 3.97222
R13172 GND.n6115 GND.n6111 3.8923
R13173 GND.n4241 GND.n4237 3.87929
R13174 GND.n6637 GND.n2894 3.87929
R13175 GND.n1922 GND.n1435 3.75785
R13176 GND.n1953 GND.n1435 3.75785
R13177 GND.t58 GND.n4846 3.64124
R13178 GND.n5155 GND.t82 3.64124
R13179 GND.n72 GND.n71 3.60163
R13180 GND.n1903 GND.n1886 3.49141
R13181 GND.n4296 GND.n4279 3.49141
R13182 GND.n2856 GND.n2839 3.49141
R13183 GND.n6089 GND.n6072 3.49141
R13184 GND.n6065 GND.n6064 3.4105
R13185 GND.n2097 GND.t62 3.31026
R13186 GND.n2044 GND.t45 3.31026
R13187 GND.t136 GND.n6944 3.31026
R13188 GND.n4148 GND.n4145 3.31026
R13189 GND.n2635 GND.n2629 3.31026
R13190 GND.n4317 GND.n2654 3.31026
R13191 GND.n6861 GND.n2662 3.31026
R13192 GND.n4437 GND.n3851 3.31026
R13193 GND.n4399 GND.t16 3.31026
R13194 GND.n4493 GND.n3822 3.31026
R13195 GND.n4607 GND.n4606 3.31026
R13196 GND.n4688 GND.n4687 3.31026
R13197 GND.n4733 GND.t54 3.31026
R13198 GND.n4783 GND.n4782 3.31026
R13199 GND.n4865 GND.n4864 3.31026
R13200 GND.t43 GND.n4901 3.31026
R13201 GND.n4960 GND.n4959 3.31026
R13202 GND.n5041 GND.n5040 3.31026
R13203 GND.n5076 GND.t4 3.31026
R13204 GND.n5136 GND.n5135 3.31026
R13205 GND.n5216 GND.n5215 3.31026
R13206 GND.t35 GND.n5231 3.31026
R13207 GND.n5310 GND.n5309 3.31026
R13208 GND.n5393 GND.n5392 3.31026
R13209 GND.n5488 GND.n5487 3.31026
R13210 GND.t33 GND.n3293 3.31026
R13211 GND.n5549 GND.n5548 3.31026
R13212 GND.n6625 GND.n2905 3.31026
R13213 GND.n3234 GND.n2914 3.31026
R13214 GND.n2939 GND.n2933 3.31026
R13215 GND.n5690 GND.n5687 3.31026
R13216 GND.n6542 GND.n6541 3.31026
R13217 GND.n6398 GND.t64 3.31026
R13218 GND.n6223 GND.t28 3.31026
R13219 GND.n1915 GND.n1879 3.15136
R13220 GND.n18 GND.n16 3.00987
R13221 GND.n33 GND.n31 3.00987
R13222 GND.n49 GND.n47 3.00987
R13223 GND.n3 GND.n1 3.00987
R13224 GND.n79 GND.n77 3.00987
R13225 GND.n94 GND.n92 3.00987
R13226 GND.n110 GND.n108 3.00987
R13227 GND.n126 GND.n124 3.00987
R13228 GND.n4607 GND.t20 2.97929
R13229 GND.n5392 GND.t80 2.97929
R13230 GND.n1651 GND.n1650 2.87436
R13231 GND.n1773 GND.n1772 2.87436
R13232 GND.n1891 GND.n1889 2.84305
R13233 GND.n4284 GND.n4282 2.84305
R13234 GND.n2844 GND.n2842 2.84305
R13235 GND.n6077 GND.n6075 2.84305
R13236 GND.n1834 GND.n1452 2.79595
R13237 GND.n6991 GND.n1435 2.77258
R13238 GND.n1876 GND.t78 2.76201
R13239 GND.n1876 GND.t79 2.76201
R13240 GND.n1878 GND.t17 2.76201
R13241 GND.n1878 GND.t85 2.76201
R13242 GND.n4310 GND.t34 2.76201
R13243 GND.n4310 GND.t23 2.76201
R13244 GND.n4308 GND.t86 2.76201
R13245 GND.n4308 GND.t87 2.76201
R13246 GND.n2870 GND.t55 2.76201
R13247 GND.n2870 GND.t44 2.76201
R13248 GND.n2868 GND.t31 2.76201
R13249 GND.n2868 GND.t211 2.76201
R13250 GND.n6104 GND.t56 2.76201
R13251 GND.n6104 GND.t32 2.76201
R13252 GND.n6101 GND.t36 2.76201
R13253 GND.n6101 GND.t38 2.76201
R13254 GND.n1904 GND.n1884 2.71565
R13255 GND.n4297 GND.n4277 2.71565
R13256 GND.n2857 GND.n2837 2.71565
R13257 GND.n4246 GND.n4241 2.71565
R13258 GND.n6090 GND.n6070 2.71565
R13259 GND.n6634 GND.n2894 2.71565
R13260 GND.n6133 GND.n6111 2.70535
R13261 GND.n6860 GND.n2664 2.64831
R13262 GND.n4365 GND.n4364 2.64831
R13263 GND.n4453 GND.n4452 2.64831
R13264 GND.n4598 GND.n4597 2.64831
R13265 GND.n3727 GND.n3726 2.64831
R13266 GND.n4774 GND.n3674 2.64831
R13267 GND.n3639 GND.n3638 2.64831
R13268 GND.n4951 GND.n3586 2.64831
R13269 GND.n3551 GND.n3550 2.64831
R13270 GND.n5127 GND.n3498 2.64831
R13271 GND.n3462 GND.n3460 2.64831
R13272 GND.n5301 GND.n3408 2.64831
R13273 GND.n5338 GND.n5337 2.64831
R13274 GND.n5479 GND.n3322 2.64831
R13275 GND.n3287 GND.n3286 2.64831
R13276 GND.n6626 GND.n2904 2.64831
R13277 GND.n6061 GND.n6060 2.55353
R13278 GND.n6062 GND.n6061 2.55353
R13279 GND.n6063 GND.n6062 2.55353
R13280 GND.n6057 GND.n6056 2.55353
R13281 GND.n6058 GND.n6057 2.55353
R13282 GND.n6059 GND.n6058 2.55353
R13283 GND.n6105 GND.n6103 2.36365
R13284 GND.n4926 GND.t48 2.31733
R13285 GND.t60 GND.n3536 2.31733
R13286 GND.n6133 GND.n6110 2.27742
R13287 GND.n6133 GND.n6109 2.27742
R13288 GND.n6133 GND.n6108 2.27742
R13289 GND.n6133 GND.n6107 2.27742
R13290 GND.n8504 GND.n155 2.27742
R13291 GND.n8504 GND.n153 2.27742
R13292 GND.n8505 GND.n8504 2.27742
R13293 GND.n8504 GND.n152 2.27742
R13294 GND.n6031 GND.n151 2.27742
R13295 GND.n6384 GND.n151 2.27742
R13296 GND.n5930 GND.n151 2.27742
R13297 GND.n6369 GND.n151 2.27742
R13298 GND.n5947 GND.n151 2.27742
R13299 GND.n2418 GND.n2417 2.27742
R13300 GND.n2418 GND.n2051 2.27742
R13301 GND.n2418 GND.n2050 2.27742
R13302 GND.n2418 GND.n2049 2.27742
R13303 GND.n2242 GND.n2048 2.27742
R13304 GND.n2407 GND.n2048 2.27742
R13305 GND.n2068 GND.n2048 2.27742
R13306 GND.n2358 GND.n2048 2.27742
R13307 GND.n2388 GND.n2048 2.27742
R13308 GND.n6991 GND.n1436 2.27742
R13309 GND.n6991 GND.n1917 2.27742
R13310 GND.n6991 GND.n1918 2.27742
R13311 GND.n6991 GND.n1919 2.27742
R13312 GND.n6950 GND.n2548 1.98636
R13313 GND.n2599 GND.n2593 1.98636
R13314 GND.n4174 GND.n4171 1.98636
R13315 GND.n4349 GND.n3889 1.98636
R13316 GND.n4408 GND.n3860 1.98636
R13317 GND.n4522 GND.n3803 1.98636
R13318 GND.n4587 GND.n3779 1.98636
R13319 GND.n4705 GND.n3712 1.98636
R13320 GND.n4749 GND.n4748 1.98636
R13321 GND.n4883 GND.n3625 1.98636
R13322 GND.n4926 GND.n4925 1.98636
R13323 GND.n5058 GND.n3536 1.98636
R13324 GND.n5101 GND.n5100 1.98636
R13325 GND.n5233 GND.n3447 1.98636
R13326 GND.n5276 GND.n5275 1.98636
R13327 GND.n5410 GND.n3360 1.98636
R13328 GND.n5454 GND.n5453 1.98636
R13329 GND.n5565 GND.n3273 1.98636
R13330 GND.n5578 GND.n5577 1.98636
R13331 GND.n5664 GND.n5661 1.98636
R13332 GND.n2975 GND.n2969 1.98636
R13333 GND.n6535 GND.n3020 1.98636
R13334 GND.n1908 GND.n1907 1.93989
R13335 GND.n4301 GND.n4300 1.93989
R13336 GND.n2861 GND.n2860 1.93989
R13337 GND.n6094 GND.n6093 1.93989
R13338 GND GND.n63 1.89648
R13339 GND.n62 GND.n61 1.73972
R13340 GND.n135 GND.n119 1.73972
R13341 GND.t18 GND.n3820 1.65538
R13342 GND.t84 GND.t20 1.65538
R13343 GND.t37 GND.t80 1.65538
R13344 GND.n5473 GND.t6 1.65538
R13345 GND.n65 GND.n64 1.56155
R13346 GND.n66 GND.n65 1.56155
R13347 GND.n67 GND.n66 1.56155
R13348 GND.n69 GND.n68 1.56155
R13349 GND.n70 GND.n69 1.56155
R13350 GND.n71 GND.n70 1.56155
R13351 GND.n4139 GND.t89 1.32441
R13352 GND.n4443 GND.n3847 1.32441
R13353 GND.n4487 GND.n3826 1.32441
R13354 GND.n4619 GND.n4618 1.32441
R13355 GND.n4678 GND.n4677 1.32441
R13356 GND.n4796 GND.n4795 1.32441
R13357 GND.n4855 GND.n4853 1.32441
R13358 GND.n4972 GND.n4971 1.32441
R13359 GND.n5031 GND.n5030 1.32441
R13360 GND.n5148 GND.n5147 1.32441
R13361 GND.n5206 GND.n5205 1.32441
R13362 GND.n5322 GND.n5321 1.32441
R13363 GND.n5383 GND.n5382 1.32441
R13364 GND.n5501 GND.n5500 1.32441
R13365 GND.n5537 GND.n5535 1.32441
R13366 GND.n5695 GND.t103 1.32441
R13367 GND.n1589 GND.n1588 1.30353
R13368 GND.n5782 GND.n5781 1.24928
R13369 GND.n3940 GND.n3939 1.24928
R13370 GND.n4035 GND.n3946 1.24928
R13371 GND.n3175 GND.n3089 1.24928
R13372 GND.n61 GND.n45 1.19878
R13373 GND.n119 GND.n103 1.19878
R13374 GND.n29 GND.n27 1.16429
R13375 GND.n44 GND.n42 1.16429
R13376 GND.n60 GND.n58 1.16429
R13377 GND.n14 GND.n12 1.16429
R13378 GND.n87 GND.n75 1.16429
R13379 GND.n102 GND.n90 1.16429
R13380 GND.n118 GND.n106 1.16429
R13381 GND.n134 GND.n122 1.16429
R13382 GND.n1911 GND.n1882 1.16414
R13383 GND.n4304 GND.n4275 1.16414
R13384 GND.n2864 GND.n2835 1.16414
R13385 GND.n6097 GND.n6068 1.16414
R13386 GND.n8514 GND.n8513 1.04891
R13387 GND.n6964 GND.n2530 0.993429
R13388 GND.n6521 GND.n3037 0.993429
R13389 GND.n1879 GND.n1877 0.788215
R13390 GND.n4311 GND.n4309 0.788215
R13391 GND.n2871 GND.n2869 0.788215
R13392 GND.n6103 GND.n6102 0.788215
R13393 GND.n3110 GND.n3104 0.776258
R13394 GND.n7020 GND.n7019 0.776258
R13395 GND.n6485 GND.n6484 0.776258
R13396 GND.n2080 GND.t12 0.662453
R13397 GND.t176 GND.n2538 0.662453
R13398 GND.n6958 GND.n6957 0.662453
R13399 GND.n4112 GND.t115 0.662453
R13400 GND.n4161 GND.n4158 0.662453
R13401 GND.n2617 GND.n2611 0.662453
R13402 GND.n4358 GND.n4357 0.662453
R13403 GND.n4387 GND.n4386 0.662453
R13404 GND.n4531 GND.n4530 0.662453
R13405 GND.n4579 GND.n4578 0.662453
R13406 GND.n4714 GND.n4713 0.662453
R13407 GND.n4740 GND.n4739 0.662453
R13408 GND.t54 GND.n3685 0.662453
R13409 GND.n4892 GND.n4891 0.662453
R13410 GND.n4917 GND.n4916 0.662453
R13411 GND.n5067 GND.n5066 0.662453
R13412 GND.n5092 GND.n5091 0.662453
R13413 GND.n5232 GND.t35 0.662453
R13414 GND.n5242 GND.n5241 0.662453
R13415 GND.n5267 GND.n5266 0.662453
R13416 GND.n5419 GND.n5418 0.662453
R13417 GND.n5445 GND.n5444 0.662453
R13418 GND.n5593 GND.n3258 0.662453
R13419 GND.n5614 GND.n3249 0.662453
R13420 GND.n2957 GND.n2951 0.662453
R13421 GND.n5677 GND.n5674 0.662453
R13422 GND.n6528 GND.n6527 0.662453
R13423 GND.n6380 GND.t0 0.662453
R13424 GND.n8504 GND.n151 0.597625
R13425 GND.n2418 GND.n2048 0.597625
R13426 GND.n1584 GND.n1529 0.502622
R13427 GND.n1566 GND.n1563 0.502622
R13428 GND.n1562 GND.n1535 0.502622
R13429 GND.n1544 GND.n1541 0.502622
R13430 GND.n1858 GND.n1857 0.502622
R13431 GND.n1856 GND.n1445 0.502622
R13432 GND.n1838 GND.n1835 0.502622
R13433 GND.n1590 GND.n1528 0.502622
R13434 GND.n1650 GND.n1510 0.502622
R13435 GND.n1651 GND.n1509 0.502622
R13436 GND.n1711 GND.n1491 0.502622
R13437 GND.n1712 GND.n1490 0.502622
R13438 GND.n1772 GND.n1472 0.502622
R13439 GND.n1773 GND.n1471 0.502622
R13440 GND.n1833 GND.n1453 0.502622
R13441 GND.n1586 GND.n1437 0.502622
R13442 GND.n280 GND.n279 0.485256
R13443 GND.n5837 GND.n3071 0.485256
R13444 GND.n7041 GND.n7040 0.485256
R13445 GND.n2169 GND.n1247 0.485256
R13446 GND.n6857 GND.n2668 0.483732
R13447 GND.n6665 GND.n6664 0.483732
R13448 GND.n6630 GND.n6629 0.483732
R13449 GND.n4322 GND.n4321 0.483732
R13450 GND.n7372 GND.n7371 0.465439
R13451 GND.n8213 GND.n8212 0.465439
R13452 GND.n8394 GND.n8393 0.465439
R13453 GND.n7225 GND.n7224 0.465439
R13454 GND.n2211 GND.n2209 0.456293
R13455 GND.n6297 GND.n6296 0.456293
R13456 GND GND.n8514 0.426242
R13457 GND.n5790 GND.n3086 0.312695
R13458 GND.n4046 GND.n1407 0.312695
R13459 GND.n3942 GND.n1407 0.312695
R13460 GND.n5790 GND.n3087 0.312695
R13461 GND.n8514 GND.n72 0.283597
R13462 GND.n314 GND.n249 0.279463
R13463 GND.n6452 GND.n5816 0.279463
R13464 GND.n7117 GND.n1287 0.279463
R13465 GND.n6993 GND.n6992 0.279463
R13466 GND.n6106 GND.n2872 0.277787
R13467 GND.n4312 GND.n1916 0.277787
R13468 GND.n6991 GND.n1434 0.268793
R13469 GND.n6134 GND.n6133 0.268793
R13470 GND.n6269 GND.n249 0.2505
R13471 GND.n2189 GND.n1287 0.2505
R13472 GND.n5792 GND.n3085 0.229039
R13473 GND.n5793 GND.n5792 0.229039
R13474 GND.n7022 GND.n1404 0.229039
R13475 GND.n7018 GND.n1404 0.229039
R13476 GND.n1580 GND.n1529 0.189894
R13477 GND.n1580 GND.n1579 0.189894
R13478 GND.n1579 GND.n1578 0.189894
R13479 GND.n1578 GND.n1531 0.189894
R13480 GND.n1574 GND.n1531 0.189894
R13481 GND.n1574 GND.n1573 0.189894
R13482 GND.n1573 GND.n1572 0.189894
R13483 GND.n1572 GND.n1533 0.189894
R13484 GND.n1568 GND.n1533 0.189894
R13485 GND.n1568 GND.n1567 0.189894
R13486 GND.n1567 GND.n1566 0.189894
R13487 GND.n1558 GND.n1535 0.189894
R13488 GND.n1558 GND.n1557 0.189894
R13489 GND.n1557 GND.n1556 0.189894
R13490 GND.n1556 GND.n1537 0.189894
R13491 GND.n1552 GND.n1537 0.189894
R13492 GND.n1552 GND.n1551 0.189894
R13493 GND.n1551 GND.n1550 0.189894
R13494 GND.n1550 GND.n1539 0.189894
R13495 GND.n1546 GND.n1539 0.189894
R13496 GND.n1546 GND.n1545 0.189894
R13497 GND.n1545 GND.n1544 0.189894
R13498 GND.n1870 GND.n1438 0.189894
R13499 GND.n1870 GND.n1869 0.189894
R13500 GND.n1869 GND.n1868 0.189894
R13501 GND.n1868 GND.n1441 0.189894
R13502 GND.n1864 GND.n1441 0.189894
R13503 GND.n1864 GND.n1863 0.189894
R13504 GND.n1863 GND.n1862 0.189894
R13505 GND.n1862 GND.n1443 0.189894
R13506 GND.n1858 GND.n1443 0.189894
R13507 GND.n1852 GND.n1445 0.189894
R13508 GND.n1852 GND.n1851 0.189894
R13509 GND.n1851 GND.n1850 0.189894
R13510 GND.n1850 GND.n1447 0.189894
R13511 GND.n1846 GND.n1447 0.189894
R13512 GND.n1846 GND.n1845 0.189894
R13513 GND.n1845 GND.n1844 0.189894
R13514 GND.n1844 GND.n1449 0.189894
R13515 GND.n1840 GND.n1449 0.189894
R13516 GND.n1840 GND.n1839 0.189894
R13517 GND.n1839 GND.n1838 0.189894
R13518 GND.n1594 GND.n1528 0.189894
R13519 GND.n1595 GND.n1594 0.189894
R13520 GND.n1596 GND.n1595 0.189894
R13521 GND.n1596 GND.n1526 0.189894
R13522 GND.n1600 GND.n1526 0.189894
R13523 GND.n1601 GND.n1600 0.189894
R13524 GND.n1602 GND.n1601 0.189894
R13525 GND.n1602 GND.n1524 0.189894
R13526 GND.n1606 GND.n1524 0.189894
R13527 GND.n1607 GND.n1606 0.189894
R13528 GND.n1608 GND.n1607 0.189894
R13529 GND.n1608 GND.n1522 0.189894
R13530 GND.n1613 GND.n1522 0.189894
R13531 GND.n1614 GND.n1613 0.189894
R13532 GND.n1615 GND.n1614 0.189894
R13533 GND.n1615 GND.n1520 0.189894
R13534 GND.n1619 GND.n1520 0.189894
R13535 GND.n1620 GND.n1619 0.189894
R13536 GND.n1621 GND.n1620 0.189894
R13537 GND.n1621 GND.n1518 0.189894
R13538 GND.n1625 GND.n1518 0.189894
R13539 GND.n1626 GND.n1625 0.189894
R13540 GND.n1627 GND.n1626 0.189894
R13541 GND.n1627 GND.n1516 0.189894
R13542 GND.n1632 GND.n1516 0.189894
R13543 GND.n1633 GND.n1632 0.189894
R13544 GND.n1634 GND.n1633 0.189894
R13545 GND.n1634 GND.n1514 0.189894
R13546 GND.n1638 GND.n1514 0.189894
R13547 GND.n1639 GND.n1638 0.189894
R13548 GND.n1640 GND.n1639 0.189894
R13549 GND.n1640 GND.n1512 0.189894
R13550 GND.n1644 GND.n1512 0.189894
R13551 GND.n1645 GND.n1644 0.189894
R13552 GND.n1646 GND.n1645 0.189894
R13553 GND.n1646 GND.n1510 0.189894
R13554 GND.n1655 GND.n1509 0.189894
R13555 GND.n1656 GND.n1655 0.189894
R13556 GND.n1657 GND.n1656 0.189894
R13557 GND.n1657 GND.n1507 0.189894
R13558 GND.n1661 GND.n1507 0.189894
R13559 GND.n1662 GND.n1661 0.189894
R13560 GND.n1663 GND.n1662 0.189894
R13561 GND.n1663 GND.n1505 0.189894
R13562 GND.n1667 GND.n1505 0.189894
R13563 GND.n1668 GND.n1667 0.189894
R13564 GND.n1669 GND.n1668 0.189894
R13565 GND.n1669 GND.n1503 0.189894
R13566 GND.n1674 GND.n1503 0.189894
R13567 GND.n1675 GND.n1674 0.189894
R13568 GND.n1676 GND.n1675 0.189894
R13569 GND.n1676 GND.n1501 0.189894
R13570 GND.n1680 GND.n1501 0.189894
R13571 GND.n1681 GND.n1680 0.189894
R13572 GND.n1682 GND.n1681 0.189894
R13573 GND.n1682 GND.n1499 0.189894
R13574 GND.n1686 GND.n1499 0.189894
R13575 GND.n1687 GND.n1686 0.189894
R13576 GND.n1688 GND.n1687 0.189894
R13577 GND.n1688 GND.n1497 0.189894
R13578 GND.n1693 GND.n1497 0.189894
R13579 GND.n1694 GND.n1693 0.189894
R13580 GND.n1695 GND.n1694 0.189894
R13581 GND.n1695 GND.n1495 0.189894
R13582 GND.n1699 GND.n1495 0.189894
R13583 GND.n1700 GND.n1699 0.189894
R13584 GND.n1701 GND.n1700 0.189894
R13585 GND.n1701 GND.n1493 0.189894
R13586 GND.n1705 GND.n1493 0.189894
R13587 GND.n1706 GND.n1705 0.189894
R13588 GND.n1707 GND.n1706 0.189894
R13589 GND.n1707 GND.n1491 0.189894
R13590 GND.n1716 GND.n1490 0.189894
R13591 GND.n1717 GND.n1716 0.189894
R13592 GND.n1718 GND.n1717 0.189894
R13593 GND.n1718 GND.n1488 0.189894
R13594 GND.n1722 GND.n1488 0.189894
R13595 GND.n1723 GND.n1722 0.189894
R13596 GND.n1724 GND.n1723 0.189894
R13597 GND.n1724 GND.n1486 0.189894
R13598 GND.n1728 GND.n1486 0.189894
R13599 GND.n1729 GND.n1728 0.189894
R13600 GND.n1730 GND.n1729 0.189894
R13601 GND.n1730 GND.n1484 0.189894
R13602 GND.n1735 GND.n1484 0.189894
R13603 GND.n1736 GND.n1735 0.189894
R13604 GND.n1737 GND.n1736 0.189894
R13605 GND.n1737 GND.n1482 0.189894
R13606 GND.n1741 GND.n1482 0.189894
R13607 GND.n1742 GND.n1741 0.189894
R13608 GND.n1743 GND.n1742 0.189894
R13609 GND.n1743 GND.n1480 0.189894
R13610 GND.n1747 GND.n1480 0.189894
R13611 GND.n1748 GND.n1747 0.189894
R13612 GND.n1749 GND.n1748 0.189894
R13613 GND.n1749 GND.n1478 0.189894
R13614 GND.n1754 GND.n1478 0.189894
R13615 GND.n1755 GND.n1754 0.189894
R13616 GND.n1756 GND.n1755 0.189894
R13617 GND.n1756 GND.n1476 0.189894
R13618 GND.n1760 GND.n1476 0.189894
R13619 GND.n1761 GND.n1760 0.189894
R13620 GND.n1762 GND.n1761 0.189894
R13621 GND.n1762 GND.n1474 0.189894
R13622 GND.n1766 GND.n1474 0.189894
R13623 GND.n1767 GND.n1766 0.189894
R13624 GND.n1768 GND.n1767 0.189894
R13625 GND.n1768 GND.n1472 0.189894
R13626 GND.n1777 GND.n1471 0.189894
R13627 GND.n1778 GND.n1777 0.189894
R13628 GND.n1779 GND.n1778 0.189894
R13629 GND.n1779 GND.n1469 0.189894
R13630 GND.n1783 GND.n1469 0.189894
R13631 GND.n1784 GND.n1783 0.189894
R13632 GND.n1785 GND.n1784 0.189894
R13633 GND.n1785 GND.n1467 0.189894
R13634 GND.n1789 GND.n1467 0.189894
R13635 GND.n1790 GND.n1789 0.189894
R13636 GND.n1791 GND.n1790 0.189894
R13637 GND.n1791 GND.n1465 0.189894
R13638 GND.n1796 GND.n1465 0.189894
R13639 GND.n1797 GND.n1796 0.189894
R13640 GND.n1798 GND.n1797 0.189894
R13641 GND.n1798 GND.n1463 0.189894
R13642 GND.n1802 GND.n1463 0.189894
R13643 GND.n1803 GND.n1802 0.189894
R13644 GND.n1804 GND.n1803 0.189894
R13645 GND.n1804 GND.n1461 0.189894
R13646 GND.n1808 GND.n1461 0.189894
R13647 GND.n1809 GND.n1808 0.189894
R13648 GND.n1810 GND.n1809 0.189894
R13649 GND.n1810 GND.n1459 0.189894
R13650 GND.n1815 GND.n1459 0.189894
R13651 GND.n1816 GND.n1815 0.189894
R13652 GND.n1817 GND.n1816 0.189894
R13653 GND.n1817 GND.n1457 0.189894
R13654 GND.n1821 GND.n1457 0.189894
R13655 GND.n1822 GND.n1821 0.189894
R13656 GND.n1823 GND.n1822 0.189894
R13657 GND.n1823 GND.n1455 0.189894
R13658 GND.n1827 GND.n1455 0.189894
R13659 GND.n1828 GND.n1827 0.189894
R13660 GND.n1829 GND.n1828 0.189894
R13661 GND.n1829 GND.n1453 0.189894
R13662 GND.n1874 GND.n1438 0.184609
R13663 GND.n24 GND.n16 0.155672
R13664 GND.n39 GND.n31 0.155672
R13665 GND.n55 GND.n47 0.155672
R13666 GND.n9 GND.n1 0.155672
R13667 GND.n1913 GND.n1881 0.155672
R13668 GND.n1906 GND.n1881 0.155672
R13669 GND.n1906 GND.n1905 0.155672
R13670 GND.n1905 GND.n1885 0.155672
R13671 GND.n1898 GND.n1885 0.155672
R13672 GND.n1898 GND.n1897 0.155672
R13673 GND.n1897 GND.n1889 0.155672
R13674 GND.n4290 GND.n4282 0.155672
R13675 GND.n4291 GND.n4290 0.155672
R13676 GND.n4291 GND.n4278 0.155672
R13677 GND.n4298 GND.n4278 0.155672
R13678 GND.n4299 GND.n4298 0.155672
R13679 GND.n4299 GND.n4274 0.155672
R13680 GND.n4306 GND.n4274 0.155672
R13681 GND.n2850 GND.n2842 0.155672
R13682 GND.n2851 GND.n2850 0.155672
R13683 GND.n2851 GND.n2838 0.155672
R13684 GND.n2858 GND.n2838 0.155672
R13685 GND.n2859 GND.n2858 0.155672
R13686 GND.n2859 GND.n2834 0.155672
R13687 GND.n2866 GND.n2834 0.155672
R13688 GND.n85 GND.n77 0.155672
R13689 GND.n100 GND.n92 0.155672
R13690 GND.n116 GND.n108 0.155672
R13691 GND.n132 GND.n124 0.155672
R13692 GND.n6099 GND.n6067 0.155672
R13693 GND.n6092 GND.n6067 0.155672
R13694 GND.n6092 GND.n6091 0.155672
R13695 GND.n6091 GND.n6071 0.155672
R13696 GND.n6084 GND.n6071 0.155672
R13697 GND.n6084 GND.n6083 0.155672
R13698 GND.n6083 GND.n6075 0.155672
R13699 GND.n2343 GND.n2342 0.152939
R13700 GND.n2344 GND.n2343 0.152939
R13701 GND.n2344 GND.n2036 0.152939
R13702 GND.n2426 GND.n2036 0.152939
R13703 GND.n2427 GND.n2426 0.152939
R13704 GND.n2428 GND.n2427 0.152939
R13705 GND.n2429 GND.n2428 0.152939
R13706 GND.n2429 GND.n2014 0.152939
R13707 GND.n2452 GND.n2014 0.152939
R13708 GND.n2453 GND.n2452 0.152939
R13709 GND.n2454 GND.n2453 0.152939
R13710 GND.n2455 GND.n2454 0.152939
R13711 GND.n2457 GND.n2455 0.152939
R13712 GND.n2457 GND.n2456 0.152939
R13713 GND.n2456 GND.n1983 0.152939
R13714 GND.n1984 GND.n1983 0.152939
R13715 GND.n1985 GND.n1984 0.152939
R13716 GND.n1986 GND.n1985 0.152939
R13717 GND.n1987 GND.n1986 0.152939
R13718 GND.n1988 GND.n1987 0.152939
R13719 GND.n1988 GND.n1434 0.152939
R13720 GND.n7372 GND.n1032 0.152939
R13721 GND.n7380 GND.n1032 0.152939
R13722 GND.n7381 GND.n7380 0.152939
R13723 GND.n7382 GND.n7381 0.152939
R13724 GND.n7382 GND.n1026 0.152939
R13725 GND.n7390 GND.n1026 0.152939
R13726 GND.n7391 GND.n7390 0.152939
R13727 GND.n7392 GND.n7391 0.152939
R13728 GND.n7392 GND.n1020 0.152939
R13729 GND.n7400 GND.n1020 0.152939
R13730 GND.n7401 GND.n7400 0.152939
R13731 GND.n7402 GND.n7401 0.152939
R13732 GND.n7402 GND.n1014 0.152939
R13733 GND.n7410 GND.n1014 0.152939
R13734 GND.n7411 GND.n7410 0.152939
R13735 GND.n7412 GND.n7411 0.152939
R13736 GND.n7412 GND.n1008 0.152939
R13737 GND.n7420 GND.n1008 0.152939
R13738 GND.n7421 GND.n7420 0.152939
R13739 GND.n7422 GND.n7421 0.152939
R13740 GND.n7422 GND.n1002 0.152939
R13741 GND.n7430 GND.n1002 0.152939
R13742 GND.n7431 GND.n7430 0.152939
R13743 GND.n7432 GND.n7431 0.152939
R13744 GND.n7432 GND.n996 0.152939
R13745 GND.n7440 GND.n996 0.152939
R13746 GND.n7441 GND.n7440 0.152939
R13747 GND.n7442 GND.n7441 0.152939
R13748 GND.n7442 GND.n990 0.152939
R13749 GND.n7450 GND.n990 0.152939
R13750 GND.n7451 GND.n7450 0.152939
R13751 GND.n7452 GND.n7451 0.152939
R13752 GND.n7452 GND.n984 0.152939
R13753 GND.n7460 GND.n984 0.152939
R13754 GND.n7461 GND.n7460 0.152939
R13755 GND.n7462 GND.n7461 0.152939
R13756 GND.n7462 GND.n978 0.152939
R13757 GND.n7470 GND.n978 0.152939
R13758 GND.n7471 GND.n7470 0.152939
R13759 GND.n7472 GND.n7471 0.152939
R13760 GND.n7472 GND.n972 0.152939
R13761 GND.n7480 GND.n972 0.152939
R13762 GND.n7481 GND.n7480 0.152939
R13763 GND.n7482 GND.n7481 0.152939
R13764 GND.n7482 GND.n966 0.152939
R13765 GND.n7490 GND.n966 0.152939
R13766 GND.n7491 GND.n7490 0.152939
R13767 GND.n7492 GND.n7491 0.152939
R13768 GND.n7492 GND.n960 0.152939
R13769 GND.n7500 GND.n960 0.152939
R13770 GND.n7501 GND.n7500 0.152939
R13771 GND.n7502 GND.n7501 0.152939
R13772 GND.n7502 GND.n954 0.152939
R13773 GND.n7510 GND.n954 0.152939
R13774 GND.n7511 GND.n7510 0.152939
R13775 GND.n7512 GND.n7511 0.152939
R13776 GND.n7512 GND.n948 0.152939
R13777 GND.n7520 GND.n948 0.152939
R13778 GND.n7521 GND.n7520 0.152939
R13779 GND.n7522 GND.n7521 0.152939
R13780 GND.n7522 GND.n942 0.152939
R13781 GND.n7530 GND.n942 0.152939
R13782 GND.n7531 GND.n7530 0.152939
R13783 GND.n7532 GND.n7531 0.152939
R13784 GND.n7532 GND.n936 0.152939
R13785 GND.n7540 GND.n936 0.152939
R13786 GND.n7541 GND.n7540 0.152939
R13787 GND.n7542 GND.n7541 0.152939
R13788 GND.n7542 GND.n930 0.152939
R13789 GND.n7550 GND.n930 0.152939
R13790 GND.n7551 GND.n7550 0.152939
R13791 GND.n7552 GND.n7551 0.152939
R13792 GND.n7552 GND.n924 0.152939
R13793 GND.n7560 GND.n924 0.152939
R13794 GND.n7561 GND.n7560 0.152939
R13795 GND.n7562 GND.n7561 0.152939
R13796 GND.n7562 GND.n918 0.152939
R13797 GND.n7570 GND.n918 0.152939
R13798 GND.n7571 GND.n7570 0.152939
R13799 GND.n7572 GND.n7571 0.152939
R13800 GND.n7572 GND.n912 0.152939
R13801 GND.n7580 GND.n912 0.152939
R13802 GND.n7581 GND.n7580 0.152939
R13803 GND.n7582 GND.n7581 0.152939
R13804 GND.n7582 GND.n906 0.152939
R13805 GND.n7590 GND.n906 0.152939
R13806 GND.n7591 GND.n7590 0.152939
R13807 GND.n7592 GND.n7591 0.152939
R13808 GND.n7592 GND.n900 0.152939
R13809 GND.n7600 GND.n900 0.152939
R13810 GND.n7601 GND.n7600 0.152939
R13811 GND.n7602 GND.n7601 0.152939
R13812 GND.n7602 GND.n894 0.152939
R13813 GND.n7610 GND.n894 0.152939
R13814 GND.n7611 GND.n7610 0.152939
R13815 GND.n7612 GND.n7611 0.152939
R13816 GND.n7612 GND.n888 0.152939
R13817 GND.n7620 GND.n888 0.152939
R13818 GND.n7621 GND.n7620 0.152939
R13819 GND.n7622 GND.n7621 0.152939
R13820 GND.n7622 GND.n882 0.152939
R13821 GND.n7630 GND.n882 0.152939
R13822 GND.n7631 GND.n7630 0.152939
R13823 GND.n7632 GND.n7631 0.152939
R13824 GND.n7632 GND.n876 0.152939
R13825 GND.n7640 GND.n876 0.152939
R13826 GND.n7641 GND.n7640 0.152939
R13827 GND.n7642 GND.n7641 0.152939
R13828 GND.n7642 GND.n870 0.152939
R13829 GND.n7650 GND.n870 0.152939
R13830 GND.n7651 GND.n7650 0.152939
R13831 GND.n7652 GND.n7651 0.152939
R13832 GND.n7652 GND.n864 0.152939
R13833 GND.n7660 GND.n864 0.152939
R13834 GND.n7661 GND.n7660 0.152939
R13835 GND.n7662 GND.n7661 0.152939
R13836 GND.n7662 GND.n858 0.152939
R13837 GND.n7670 GND.n858 0.152939
R13838 GND.n7671 GND.n7670 0.152939
R13839 GND.n7672 GND.n7671 0.152939
R13840 GND.n7672 GND.n852 0.152939
R13841 GND.n7680 GND.n852 0.152939
R13842 GND.n7681 GND.n7680 0.152939
R13843 GND.n7682 GND.n7681 0.152939
R13844 GND.n7682 GND.n846 0.152939
R13845 GND.n7690 GND.n846 0.152939
R13846 GND.n7691 GND.n7690 0.152939
R13847 GND.n7692 GND.n7691 0.152939
R13848 GND.n7692 GND.n840 0.152939
R13849 GND.n7700 GND.n840 0.152939
R13850 GND.n7701 GND.n7700 0.152939
R13851 GND.n7702 GND.n7701 0.152939
R13852 GND.n7702 GND.n834 0.152939
R13853 GND.n7710 GND.n834 0.152939
R13854 GND.n7711 GND.n7710 0.152939
R13855 GND.n7712 GND.n7711 0.152939
R13856 GND.n7712 GND.n828 0.152939
R13857 GND.n7720 GND.n828 0.152939
R13858 GND.n7721 GND.n7720 0.152939
R13859 GND.n7722 GND.n7721 0.152939
R13860 GND.n7722 GND.n822 0.152939
R13861 GND.n7730 GND.n822 0.152939
R13862 GND.n7731 GND.n7730 0.152939
R13863 GND.n7732 GND.n7731 0.152939
R13864 GND.n7732 GND.n816 0.152939
R13865 GND.n7740 GND.n816 0.152939
R13866 GND.n7741 GND.n7740 0.152939
R13867 GND.n7742 GND.n7741 0.152939
R13868 GND.n7742 GND.n810 0.152939
R13869 GND.n7750 GND.n810 0.152939
R13870 GND.n7751 GND.n7750 0.152939
R13871 GND.n7752 GND.n7751 0.152939
R13872 GND.n7752 GND.n804 0.152939
R13873 GND.n7760 GND.n804 0.152939
R13874 GND.n7761 GND.n7760 0.152939
R13875 GND.n7762 GND.n7761 0.152939
R13876 GND.n7762 GND.n798 0.152939
R13877 GND.n7770 GND.n798 0.152939
R13878 GND.n7771 GND.n7770 0.152939
R13879 GND.n7772 GND.n7771 0.152939
R13880 GND.n7772 GND.n792 0.152939
R13881 GND.n7780 GND.n792 0.152939
R13882 GND.n7781 GND.n7780 0.152939
R13883 GND.n7782 GND.n7781 0.152939
R13884 GND.n7782 GND.n786 0.152939
R13885 GND.n7790 GND.n786 0.152939
R13886 GND.n7791 GND.n7790 0.152939
R13887 GND.n7792 GND.n7791 0.152939
R13888 GND.n7792 GND.n780 0.152939
R13889 GND.n7800 GND.n780 0.152939
R13890 GND.n7801 GND.n7800 0.152939
R13891 GND.n7802 GND.n7801 0.152939
R13892 GND.n7802 GND.n774 0.152939
R13893 GND.n7810 GND.n774 0.152939
R13894 GND.n7811 GND.n7810 0.152939
R13895 GND.n7812 GND.n7811 0.152939
R13896 GND.n7812 GND.n768 0.152939
R13897 GND.n7820 GND.n768 0.152939
R13898 GND.n7821 GND.n7820 0.152939
R13899 GND.n7822 GND.n7821 0.152939
R13900 GND.n7822 GND.n762 0.152939
R13901 GND.n7830 GND.n762 0.152939
R13902 GND.n7831 GND.n7830 0.152939
R13903 GND.n7832 GND.n7831 0.152939
R13904 GND.n7832 GND.n756 0.152939
R13905 GND.n7840 GND.n756 0.152939
R13906 GND.n7841 GND.n7840 0.152939
R13907 GND.n7842 GND.n7841 0.152939
R13908 GND.n7842 GND.n750 0.152939
R13909 GND.n7850 GND.n750 0.152939
R13910 GND.n7851 GND.n7850 0.152939
R13911 GND.n7852 GND.n7851 0.152939
R13912 GND.n7852 GND.n744 0.152939
R13913 GND.n7860 GND.n744 0.152939
R13914 GND.n7861 GND.n7860 0.152939
R13915 GND.n7862 GND.n7861 0.152939
R13916 GND.n7862 GND.n738 0.152939
R13917 GND.n7870 GND.n738 0.152939
R13918 GND.n7871 GND.n7870 0.152939
R13919 GND.n7872 GND.n7871 0.152939
R13920 GND.n7872 GND.n732 0.152939
R13921 GND.n7880 GND.n732 0.152939
R13922 GND.n7881 GND.n7880 0.152939
R13923 GND.n7882 GND.n7881 0.152939
R13924 GND.n7882 GND.n726 0.152939
R13925 GND.n7890 GND.n726 0.152939
R13926 GND.n7891 GND.n7890 0.152939
R13927 GND.n7892 GND.n7891 0.152939
R13928 GND.n7892 GND.n720 0.152939
R13929 GND.n7900 GND.n720 0.152939
R13930 GND.n7901 GND.n7900 0.152939
R13931 GND.n7902 GND.n7901 0.152939
R13932 GND.n7902 GND.n714 0.152939
R13933 GND.n7910 GND.n714 0.152939
R13934 GND.n7911 GND.n7910 0.152939
R13935 GND.n7912 GND.n7911 0.152939
R13936 GND.n7912 GND.n708 0.152939
R13937 GND.n7920 GND.n708 0.152939
R13938 GND.n7921 GND.n7920 0.152939
R13939 GND.n7922 GND.n7921 0.152939
R13940 GND.n7922 GND.n702 0.152939
R13941 GND.n7930 GND.n702 0.152939
R13942 GND.n7931 GND.n7930 0.152939
R13943 GND.n7932 GND.n7931 0.152939
R13944 GND.n7932 GND.n696 0.152939
R13945 GND.n7940 GND.n696 0.152939
R13946 GND.n7941 GND.n7940 0.152939
R13947 GND.n7942 GND.n7941 0.152939
R13948 GND.n7942 GND.n690 0.152939
R13949 GND.n7950 GND.n690 0.152939
R13950 GND.n7951 GND.n7950 0.152939
R13951 GND.n7952 GND.n7951 0.152939
R13952 GND.n7952 GND.n684 0.152939
R13953 GND.n7960 GND.n684 0.152939
R13954 GND.n7961 GND.n7960 0.152939
R13955 GND.n7962 GND.n7961 0.152939
R13956 GND.n7962 GND.n678 0.152939
R13957 GND.n7970 GND.n678 0.152939
R13958 GND.n7971 GND.n7970 0.152939
R13959 GND.n7972 GND.n7971 0.152939
R13960 GND.n7972 GND.n672 0.152939
R13961 GND.n7980 GND.n672 0.152939
R13962 GND.n7981 GND.n7980 0.152939
R13963 GND.n7982 GND.n7981 0.152939
R13964 GND.n7982 GND.n666 0.152939
R13965 GND.n7990 GND.n666 0.152939
R13966 GND.n7991 GND.n7990 0.152939
R13967 GND.n7992 GND.n7991 0.152939
R13968 GND.n7992 GND.n660 0.152939
R13969 GND.n8000 GND.n660 0.152939
R13970 GND.n8001 GND.n8000 0.152939
R13971 GND.n8002 GND.n8001 0.152939
R13972 GND.n8002 GND.n654 0.152939
R13973 GND.n8010 GND.n654 0.152939
R13974 GND.n8011 GND.n8010 0.152939
R13975 GND.n8012 GND.n8011 0.152939
R13976 GND.n8012 GND.n648 0.152939
R13977 GND.n8020 GND.n648 0.152939
R13978 GND.n8021 GND.n8020 0.152939
R13979 GND.n8022 GND.n8021 0.152939
R13980 GND.n8022 GND.n642 0.152939
R13981 GND.n8030 GND.n642 0.152939
R13982 GND.n8031 GND.n8030 0.152939
R13983 GND.n8032 GND.n8031 0.152939
R13984 GND.n8032 GND.n636 0.152939
R13985 GND.n8040 GND.n636 0.152939
R13986 GND.n8041 GND.n8040 0.152939
R13987 GND.n8042 GND.n8041 0.152939
R13988 GND.n8042 GND.n630 0.152939
R13989 GND.n8050 GND.n630 0.152939
R13990 GND.n8051 GND.n8050 0.152939
R13991 GND.n8052 GND.n8051 0.152939
R13992 GND.n8052 GND.n624 0.152939
R13993 GND.n8060 GND.n624 0.152939
R13994 GND.n8061 GND.n8060 0.152939
R13995 GND.n8062 GND.n8061 0.152939
R13996 GND.n8062 GND.n618 0.152939
R13997 GND.n8070 GND.n618 0.152939
R13998 GND.n8071 GND.n8070 0.152939
R13999 GND.n8072 GND.n8071 0.152939
R14000 GND.n8072 GND.n612 0.152939
R14001 GND.n8080 GND.n612 0.152939
R14002 GND.n8081 GND.n8080 0.152939
R14003 GND.n8082 GND.n8081 0.152939
R14004 GND.n8082 GND.n606 0.152939
R14005 GND.n8090 GND.n606 0.152939
R14006 GND.n8091 GND.n8090 0.152939
R14007 GND.n8092 GND.n8091 0.152939
R14008 GND.n8092 GND.n600 0.152939
R14009 GND.n8100 GND.n600 0.152939
R14010 GND.n8101 GND.n8100 0.152939
R14011 GND.n8102 GND.n8101 0.152939
R14012 GND.n8102 GND.n594 0.152939
R14013 GND.n8110 GND.n594 0.152939
R14014 GND.n8111 GND.n8110 0.152939
R14015 GND.n8112 GND.n8111 0.152939
R14016 GND.n8112 GND.n588 0.152939
R14017 GND.n8120 GND.n588 0.152939
R14018 GND.n8121 GND.n8120 0.152939
R14019 GND.n8122 GND.n8121 0.152939
R14020 GND.n8122 GND.n582 0.152939
R14021 GND.n8130 GND.n582 0.152939
R14022 GND.n8131 GND.n8130 0.152939
R14023 GND.n8132 GND.n8131 0.152939
R14024 GND.n8132 GND.n576 0.152939
R14025 GND.n8140 GND.n576 0.152939
R14026 GND.n8141 GND.n8140 0.152939
R14027 GND.n8142 GND.n8141 0.152939
R14028 GND.n8142 GND.n570 0.152939
R14029 GND.n8150 GND.n570 0.152939
R14030 GND.n8151 GND.n8150 0.152939
R14031 GND.n8152 GND.n8151 0.152939
R14032 GND.n8152 GND.n564 0.152939
R14033 GND.n8160 GND.n564 0.152939
R14034 GND.n8161 GND.n8160 0.152939
R14035 GND.n8162 GND.n8161 0.152939
R14036 GND.n8162 GND.n558 0.152939
R14037 GND.n8170 GND.n558 0.152939
R14038 GND.n8171 GND.n8170 0.152939
R14039 GND.n8172 GND.n8171 0.152939
R14040 GND.n8172 GND.n552 0.152939
R14041 GND.n8180 GND.n552 0.152939
R14042 GND.n8181 GND.n8180 0.152939
R14043 GND.n8182 GND.n8181 0.152939
R14044 GND.n8182 GND.n546 0.152939
R14045 GND.n8190 GND.n546 0.152939
R14046 GND.n8191 GND.n8190 0.152939
R14047 GND.n8192 GND.n8191 0.152939
R14048 GND.n8192 GND.n540 0.152939
R14049 GND.n8200 GND.n540 0.152939
R14050 GND.n8201 GND.n8200 0.152939
R14051 GND.n8203 GND.n8201 0.152939
R14052 GND.n8203 GND.n8202 0.152939
R14053 GND.n8202 GND.n534 0.152939
R14054 GND.n8212 GND.n534 0.152939
R14055 GND.n8213 GND.n529 0.152939
R14056 GND.n8221 GND.n529 0.152939
R14057 GND.n8222 GND.n8221 0.152939
R14058 GND.n8223 GND.n8222 0.152939
R14059 GND.n8223 GND.n523 0.152939
R14060 GND.n8231 GND.n523 0.152939
R14061 GND.n8232 GND.n8231 0.152939
R14062 GND.n8233 GND.n8232 0.152939
R14063 GND.n8233 GND.n517 0.152939
R14064 GND.n8241 GND.n517 0.152939
R14065 GND.n8242 GND.n8241 0.152939
R14066 GND.n8243 GND.n8242 0.152939
R14067 GND.n8243 GND.n511 0.152939
R14068 GND.n8251 GND.n511 0.152939
R14069 GND.n8252 GND.n8251 0.152939
R14070 GND.n8253 GND.n8252 0.152939
R14071 GND.n8253 GND.n505 0.152939
R14072 GND.n8261 GND.n505 0.152939
R14073 GND.n8262 GND.n8261 0.152939
R14074 GND.n8263 GND.n8262 0.152939
R14075 GND.n8263 GND.n499 0.152939
R14076 GND.n8271 GND.n499 0.152939
R14077 GND.n8272 GND.n8271 0.152939
R14078 GND.n8273 GND.n8272 0.152939
R14079 GND.n8273 GND.n493 0.152939
R14080 GND.n8281 GND.n493 0.152939
R14081 GND.n8282 GND.n8281 0.152939
R14082 GND.n8283 GND.n8282 0.152939
R14083 GND.n8283 GND.n487 0.152939
R14084 GND.n8291 GND.n487 0.152939
R14085 GND.n8292 GND.n8291 0.152939
R14086 GND.n8293 GND.n8292 0.152939
R14087 GND.n8293 GND.n481 0.152939
R14088 GND.n8301 GND.n481 0.152939
R14089 GND.n8302 GND.n8301 0.152939
R14090 GND.n8303 GND.n8302 0.152939
R14091 GND.n8303 GND.n475 0.152939
R14092 GND.n8311 GND.n475 0.152939
R14093 GND.n8312 GND.n8311 0.152939
R14094 GND.n8313 GND.n8312 0.152939
R14095 GND.n8313 GND.n469 0.152939
R14096 GND.n8321 GND.n469 0.152939
R14097 GND.n8322 GND.n8321 0.152939
R14098 GND.n8323 GND.n8322 0.152939
R14099 GND.n8323 GND.n463 0.152939
R14100 GND.n8331 GND.n463 0.152939
R14101 GND.n8332 GND.n8331 0.152939
R14102 GND.n8333 GND.n8332 0.152939
R14103 GND.n8333 GND.n457 0.152939
R14104 GND.n8341 GND.n457 0.152939
R14105 GND.n8342 GND.n8341 0.152939
R14106 GND.n8343 GND.n8342 0.152939
R14107 GND.n8343 GND.n451 0.152939
R14108 GND.n8351 GND.n451 0.152939
R14109 GND.n8352 GND.n8351 0.152939
R14110 GND.n8353 GND.n8352 0.152939
R14111 GND.n8353 GND.n445 0.152939
R14112 GND.n8361 GND.n445 0.152939
R14113 GND.n8362 GND.n8361 0.152939
R14114 GND.n8363 GND.n8362 0.152939
R14115 GND.n8363 GND.n439 0.152939
R14116 GND.n8371 GND.n439 0.152939
R14117 GND.n8372 GND.n8371 0.152939
R14118 GND.n8373 GND.n8372 0.152939
R14119 GND.n8373 GND.n433 0.152939
R14120 GND.n8381 GND.n433 0.152939
R14121 GND.n8382 GND.n8381 0.152939
R14122 GND.n8383 GND.n8382 0.152939
R14123 GND.n8383 GND.n427 0.152939
R14124 GND.n8391 GND.n427 0.152939
R14125 GND.n8392 GND.n8391 0.152939
R14126 GND.n8394 GND.n8392 0.152939
R14127 GND.n5950 GND.n5949 0.152939
R14128 GND.n5953 GND.n5950 0.152939
R14129 GND.n5954 GND.n5953 0.152939
R14130 GND.n5955 GND.n5954 0.152939
R14131 GND.n5956 GND.n5955 0.152939
R14132 GND.n6315 GND.n5956 0.152939
R14133 GND.n6316 GND.n6315 0.152939
R14134 GND.n6317 GND.n6316 0.152939
R14135 GND.n6317 GND.n6311 0.152939
R14136 GND.n6323 GND.n6311 0.152939
R14137 GND.n6324 GND.n6323 0.152939
R14138 GND.n6325 GND.n6324 0.152939
R14139 GND.n6326 GND.n6325 0.152939
R14140 GND.n6328 GND.n6326 0.152939
R14141 GND.n6328 GND.n6327 0.152939
R14142 GND.n6327 GND.n257 0.152939
R14143 GND.n258 GND.n257 0.152939
R14144 GND.n259 GND.n258 0.152939
R14145 GND.n386 GND.n259 0.152939
R14146 GND.n387 GND.n386 0.152939
R14147 GND.n388 GND.n387 0.152939
R14148 GND.n389 GND.n388 0.152939
R14149 GND.n394 GND.n389 0.152939
R14150 GND.n395 GND.n394 0.152939
R14151 GND.n396 GND.n395 0.152939
R14152 GND.n397 GND.n396 0.152939
R14153 GND.n402 GND.n397 0.152939
R14154 GND.n403 GND.n402 0.152939
R14155 GND.n404 GND.n403 0.152939
R14156 GND.n405 GND.n404 0.152939
R14157 GND.n410 GND.n405 0.152939
R14158 GND.n411 GND.n410 0.152939
R14159 GND.n412 GND.n411 0.152939
R14160 GND.n413 GND.n412 0.152939
R14161 GND.n418 GND.n413 0.152939
R14162 GND.n419 GND.n418 0.152939
R14163 GND.n420 GND.n419 0.152939
R14164 GND.n421 GND.n420 0.152939
R14165 GND.n8393 GND.n421 0.152939
R14166 GND.n177 GND.n149 0.152939
R14167 GND.n178 GND.n177 0.152939
R14168 GND.n179 GND.n178 0.152939
R14169 GND.n196 GND.n179 0.152939
R14170 GND.n197 GND.n196 0.152939
R14171 GND.n198 GND.n197 0.152939
R14172 GND.n199 GND.n198 0.152939
R14173 GND.n217 GND.n199 0.152939
R14174 GND.n218 GND.n217 0.152939
R14175 GND.n219 GND.n218 0.152939
R14176 GND.n220 GND.n219 0.152939
R14177 GND.n237 GND.n220 0.152939
R14178 GND.n238 GND.n237 0.152939
R14179 GND.n239 GND.n238 0.152939
R14180 GND.n240 GND.n239 0.152939
R14181 GND.n279 GND.n240 0.152939
R14182 GND.n6135 GND.n6134 0.152939
R14183 GND.n6135 GND.n6049 0.152939
R14184 GND.n6141 GND.n6049 0.152939
R14185 GND.n6142 GND.n6141 0.152939
R14186 GND.n6143 GND.n6142 0.152939
R14187 GND.n6143 GND.n6045 0.152939
R14188 GND.n6156 GND.n6045 0.152939
R14189 GND.n6157 GND.n6156 0.152939
R14190 GND.n6158 GND.n6157 0.152939
R14191 GND.n6158 GND.n6041 0.152939
R14192 GND.n6171 GND.n6041 0.152939
R14193 GND.n6172 GND.n6171 0.152939
R14194 GND.n6173 GND.n6172 0.152939
R14195 GND.n6173 GND.n6037 0.152939
R14196 GND.n6186 GND.n6037 0.152939
R14197 GND.n6187 GND.n6186 0.152939
R14198 GND.n6188 GND.n6187 0.152939
R14199 GND.n6189 GND.n6188 0.152939
R14200 GND.n6190 GND.n6189 0.152939
R14201 GND.n6191 GND.n6190 0.152939
R14202 GND.n6191 GND.n136 0.152939
R14203 GND.n8511 GND.n137 0.152939
R14204 GND.n5971 GND.n137 0.152939
R14205 GND.n6218 GND.n5971 0.152939
R14206 GND.n6219 GND.n6218 0.152939
R14207 GND.n6220 GND.n6219 0.152939
R14208 GND.n6220 GND.n5967 0.152939
R14209 GND.n6233 GND.n5967 0.152939
R14210 GND.n6234 GND.n6233 0.152939
R14211 GND.n6236 GND.n6234 0.152939
R14212 GND.n6236 GND.n6235 0.152939
R14213 GND.n6235 GND.n5961 0.152939
R14214 GND.n5962 GND.n5961 0.152939
R14215 GND.n5963 GND.n5962 0.152939
R14216 GND.n6248 GND.n5963 0.152939
R14217 GND.n6249 GND.n6248 0.152939
R14218 GND.n6250 GND.n6249 0.152939
R14219 GND.n6251 GND.n6250 0.152939
R14220 GND.n6254 GND.n6251 0.152939
R14221 GND.n6255 GND.n6254 0.152939
R14222 GND.n6256 GND.n6255 0.152939
R14223 GND.n6297 GND.n6256 0.152939
R14224 GND.n6269 GND.n6267 0.152939
R14225 GND.n6277 GND.n6267 0.152939
R14226 GND.n6278 GND.n6277 0.152939
R14227 GND.n6279 GND.n6278 0.152939
R14228 GND.n6279 GND.n6263 0.152939
R14229 GND.n6287 GND.n6263 0.152939
R14230 GND.n6288 GND.n6287 0.152939
R14231 GND.n6289 GND.n6288 0.152939
R14232 GND.n6289 GND.n6257 0.152939
R14233 GND.n6296 GND.n6257 0.152939
R14234 GND.n379 GND.n280 0.152939
R14235 GND.n379 GND.n378 0.152939
R14236 GND.n378 GND.n377 0.152939
R14237 GND.n377 GND.n282 0.152939
R14238 GND.n283 GND.n282 0.152939
R14239 GND.n284 GND.n283 0.152939
R14240 GND.n285 GND.n284 0.152939
R14241 GND.n286 GND.n285 0.152939
R14242 GND.n361 GND.n286 0.152939
R14243 GND.n361 GND.n360 0.152939
R14244 GND.n360 GND.n359 0.152939
R14245 GND.n359 GND.n290 0.152939
R14246 GND.n291 GND.n290 0.152939
R14247 GND.n292 GND.n291 0.152939
R14248 GND.n293 GND.n292 0.152939
R14249 GND.n294 GND.n293 0.152939
R14250 GND.n295 GND.n294 0.152939
R14251 GND.n296 GND.n295 0.152939
R14252 GND.n297 GND.n296 0.152939
R14253 GND.n338 GND.n297 0.152939
R14254 GND.n338 GND.n337 0.152939
R14255 GND.n337 GND.n336 0.152939
R14256 GND.n336 GND.n303 0.152939
R14257 GND.n304 GND.n303 0.152939
R14258 GND.n305 GND.n304 0.152939
R14259 GND.n306 GND.n305 0.152939
R14260 GND.n307 GND.n306 0.152939
R14261 GND.n308 GND.n307 0.152939
R14262 GND.n309 GND.n308 0.152939
R14263 GND.n310 GND.n309 0.152939
R14264 GND.n315 GND.n310 0.152939
R14265 GND.n315 GND.n314 0.152939
R14266 GND.n3072 GND.n3071 0.152939
R14267 GND.n3073 GND.n3072 0.152939
R14268 GND.n3074 GND.n3073 0.152939
R14269 GND.n3075 GND.n3074 0.152939
R14270 GND.n3076 GND.n3075 0.152939
R14271 GND.n3077 GND.n3076 0.152939
R14272 GND.n3078 GND.n3077 0.152939
R14273 GND.n3079 GND.n3078 0.152939
R14274 GND.n3080 GND.n3079 0.152939
R14275 GND.n3083 GND.n3080 0.152939
R14276 GND.n3084 GND.n3083 0.152939
R14277 GND.n3085 GND.n3084 0.152939
R14278 GND.n5794 GND.n5793 0.152939
R14279 GND.n5795 GND.n5794 0.152939
R14280 GND.n5796 GND.n5795 0.152939
R14281 GND.n5797 GND.n5796 0.152939
R14282 GND.n5799 GND.n5797 0.152939
R14283 GND.n5802 GND.n5799 0.152939
R14284 GND.n5803 GND.n5802 0.152939
R14285 GND.n5804 GND.n5803 0.152939
R14286 GND.n5805 GND.n5804 0.152939
R14287 GND.n5806 GND.n5805 0.152939
R14288 GND.n5807 GND.n5806 0.152939
R14289 GND.n5808 GND.n5807 0.152939
R14290 GND.n5809 GND.n5808 0.152939
R14291 GND.n5810 GND.n5809 0.152939
R14292 GND.n6454 GND.n5810 0.152939
R14293 GND.n6454 GND.n6453 0.152939
R14294 GND.n6453 GND.n6452 0.152939
R14295 GND.n5838 GND.n5837 0.152939
R14296 GND.n5839 GND.n5838 0.152939
R14297 GND.n5840 GND.n5839 0.152939
R14298 GND.n5841 GND.n5840 0.152939
R14299 GND.n5862 GND.n5841 0.152939
R14300 GND.n5863 GND.n5862 0.152939
R14301 GND.n5864 GND.n5863 0.152939
R14302 GND.n5865 GND.n5864 0.152939
R14303 GND.n5883 GND.n5865 0.152939
R14304 GND.n5884 GND.n5883 0.152939
R14305 GND.n5885 GND.n5884 0.152939
R14306 GND.n5886 GND.n5885 0.152939
R14307 GND.n5904 GND.n5886 0.152939
R14308 GND.n5905 GND.n5904 0.152939
R14309 GND.n5906 GND.n5905 0.152939
R14310 GND.n5906 GND.n150 0.152939
R14311 GND.n2362 GND.n2361 0.152939
R14312 GND.n2363 GND.n2362 0.152939
R14313 GND.n2364 GND.n2363 0.152939
R14314 GND.n2367 GND.n2364 0.152939
R14315 GND.n2368 GND.n2367 0.152939
R14316 GND.n2369 GND.n2368 0.152939
R14317 GND.n2370 GND.n2369 0.152939
R14318 GND.n2372 GND.n2370 0.152939
R14319 GND.n2372 GND.n2371 0.152939
R14320 GND.n2371 GND.n1996 0.152939
R14321 GND.n2482 GND.n1996 0.152939
R14322 GND.n2483 GND.n2482 0.152939
R14323 GND.n2484 GND.n2483 0.152939
R14324 GND.n2486 GND.n2484 0.152939
R14325 GND.n2486 GND.n2485 0.152939
R14326 GND.n2485 GND.n1960 0.152939
R14327 GND.n2523 GND.n1960 0.152939
R14328 GND.n2524 GND.n2523 0.152939
R14329 GND.n2525 GND.n2524 0.152939
R14330 GND.n2526 GND.n2525 0.152939
R14331 GND.n2527 GND.n2526 0.152939
R14332 GND.n2532 GND.n2527 0.152939
R14333 GND.n2533 GND.n2532 0.152939
R14334 GND.n2534 GND.n2533 0.152939
R14335 GND.n2535 GND.n2534 0.152939
R14336 GND.n2550 GND.n2535 0.152939
R14337 GND.n2551 GND.n2550 0.152939
R14338 GND.n2552 GND.n2551 0.152939
R14339 GND.n2553 GND.n2552 0.152939
R14340 GND.n2568 GND.n2553 0.152939
R14341 GND.n2569 GND.n2568 0.152939
R14342 GND.n2570 GND.n2569 0.152939
R14343 GND.n2571 GND.n2570 0.152939
R14344 GND.n2585 GND.n2571 0.152939
R14345 GND.n2586 GND.n2585 0.152939
R14346 GND.n2587 GND.n2586 0.152939
R14347 GND.n2588 GND.n2587 0.152939
R14348 GND.n2603 GND.n2588 0.152939
R14349 GND.n2604 GND.n2603 0.152939
R14350 GND.n2605 GND.n2604 0.152939
R14351 GND.n2606 GND.n2605 0.152939
R14352 GND.n2621 GND.n2606 0.152939
R14353 GND.n2622 GND.n2621 0.152939
R14354 GND.n2623 GND.n2622 0.152939
R14355 GND.n2624 GND.n2623 0.152939
R14356 GND.n2639 GND.n2624 0.152939
R14357 GND.n2640 GND.n2639 0.152939
R14358 GND.n2641 GND.n2640 0.152939
R14359 GND.n2642 GND.n2641 0.152939
R14360 GND.n2656 GND.n2642 0.152939
R14361 GND.n2657 GND.n2656 0.152939
R14362 GND.n2658 GND.n2657 0.152939
R14363 GND.n2659 GND.n2658 0.152939
R14364 GND.n3888 GND.n2659 0.152939
R14365 GND.n4352 GND.n3888 0.152939
R14366 GND.n4353 GND.n4352 0.152939
R14367 GND.n4354 GND.n4353 0.152939
R14368 GND.n4354 GND.n3871 0.152939
R14369 GND.n4390 GND.n3871 0.152939
R14370 GND.n4391 GND.n4390 0.152939
R14371 GND.n4392 GND.n4391 0.152939
R14372 GND.n4393 GND.n4392 0.152939
R14373 GND.n4394 GND.n4393 0.152939
R14374 GND.n4396 GND.n4394 0.152939
R14375 GND.n4397 GND.n4396 0.152939
R14376 GND.n4397 GND.n3831 0.152939
R14377 GND.n4479 GND.n3831 0.152939
R14378 GND.n4480 GND.n4479 0.152939
R14379 GND.n4481 GND.n4480 0.152939
R14380 GND.n4482 GND.n4481 0.152939
R14381 GND.n4482 GND.n3800 0.152939
R14382 GND.n4525 GND.n3800 0.152939
R14383 GND.n4526 GND.n4525 0.152939
R14384 GND.n4527 GND.n4526 0.152939
R14385 GND.n4527 GND.n3782 0.152939
R14386 GND.n4582 GND.n3782 0.152939
R14387 GND.n4583 GND.n4582 0.152939
R14388 GND.n4584 GND.n4583 0.152939
R14389 GND.n4584 GND.n3759 0.152939
R14390 GND.n4610 GND.n3759 0.152939
R14391 GND.n4611 GND.n4610 0.152939
R14392 GND.n4612 GND.n4611 0.152939
R14393 GND.n4613 GND.n4612 0.152939
R14394 GND.n4613 GND.n3730 0.152939
R14395 GND.n4682 GND.n3730 0.152939
R14396 GND.n4683 GND.n4682 0.152939
R14397 GND.n4684 GND.n4683 0.152939
R14398 GND.n4684 GND.n3709 0.152939
R14399 GND.n4708 GND.n3709 0.152939
R14400 GND.n4709 GND.n4708 0.152939
R14401 GND.n4710 GND.n4709 0.152939
R14402 GND.n4710 GND.n3688 0.152939
R14403 GND.n4743 GND.n3688 0.152939
R14404 GND.n4744 GND.n4743 0.152939
R14405 GND.n4745 GND.n4744 0.152939
R14406 GND.n4745 GND.n3671 0.152939
R14407 GND.n4786 GND.n3671 0.152939
R14408 GND.n4787 GND.n4786 0.152939
R14409 GND.n4788 GND.n4787 0.152939
R14410 GND.n4789 GND.n4788 0.152939
R14411 GND.n4789 GND.n3642 0.152939
R14412 GND.n4859 GND.n3642 0.152939
R14413 GND.n4860 GND.n4859 0.152939
R14414 GND.n4861 GND.n4860 0.152939
R14415 GND.n4861 GND.n3622 0.152939
R14416 GND.n4886 GND.n3622 0.152939
R14417 GND.n4887 GND.n4886 0.152939
R14418 GND.n4888 GND.n4887 0.152939
R14419 GND.n4888 GND.n3600 0.152939
R14420 GND.n4920 GND.n3600 0.152939
R14421 GND.n4921 GND.n4920 0.152939
R14422 GND.n4922 GND.n4921 0.152939
R14423 GND.n4922 GND.n3583 0.152939
R14424 GND.n4963 GND.n3583 0.152939
R14425 GND.n4964 GND.n4963 0.152939
R14426 GND.n4965 GND.n4964 0.152939
R14427 GND.n4966 GND.n4965 0.152939
R14428 GND.n4966 GND.n3554 0.152939
R14429 GND.n5035 GND.n3554 0.152939
R14430 GND.n5036 GND.n5035 0.152939
R14431 GND.n5037 GND.n5036 0.152939
R14432 GND.n5037 GND.n3533 0.152939
R14433 GND.n5061 GND.n3533 0.152939
R14434 GND.n5062 GND.n5061 0.152939
R14435 GND.n5063 GND.n5062 0.152939
R14436 GND.n5063 GND.n3511 0.152939
R14437 GND.n5095 GND.n3511 0.152939
R14438 GND.n5096 GND.n5095 0.152939
R14439 GND.n5097 GND.n5096 0.152939
R14440 GND.n5097 GND.n3494 0.152939
R14441 GND.n5139 GND.n3494 0.152939
R14442 GND.n5140 GND.n5139 0.152939
R14443 GND.n5141 GND.n5140 0.152939
R14444 GND.n5142 GND.n5141 0.152939
R14445 GND.n5142 GND.n3465 0.152939
R14446 GND.n5210 GND.n3465 0.152939
R14447 GND.n5211 GND.n5210 0.152939
R14448 GND.n5212 GND.n5211 0.152939
R14449 GND.n5212 GND.n3444 0.152939
R14450 GND.n5236 GND.n3444 0.152939
R14451 GND.n5237 GND.n5236 0.152939
R14452 GND.n5238 GND.n5237 0.152939
R14453 GND.n5238 GND.n3422 0.152939
R14454 GND.n5270 GND.n3422 0.152939
R14455 GND.n5271 GND.n5270 0.152939
R14456 GND.n5272 GND.n5271 0.152939
R14457 GND.n5272 GND.n3405 0.152939
R14458 GND.n5313 GND.n3405 0.152939
R14459 GND.n5314 GND.n5313 0.152939
R14460 GND.n5315 GND.n5314 0.152939
R14461 GND.n5316 GND.n5315 0.152939
R14462 GND.n5316 GND.n3376 0.152939
R14463 GND.n5387 GND.n3376 0.152939
R14464 GND.n5388 GND.n5387 0.152939
R14465 GND.n5389 GND.n5388 0.152939
R14466 GND.n5389 GND.n3357 0.152939
R14467 GND.n5413 GND.n3357 0.152939
R14468 GND.n5414 GND.n5413 0.152939
R14469 GND.n5415 GND.n5414 0.152939
R14470 GND.n5415 GND.n3336 0.152939
R14471 GND.n5448 GND.n3336 0.152939
R14472 GND.n5449 GND.n5448 0.152939
R14473 GND.n5450 GND.n5449 0.152939
R14474 GND.n5450 GND.n3319 0.152939
R14475 GND.n5491 GND.n3319 0.152939
R14476 GND.n5492 GND.n5491 0.152939
R14477 GND.n5493 GND.n5492 0.152939
R14478 GND.n5494 GND.n5493 0.152939
R14479 GND.n5494 GND.n3290 0.152939
R14480 GND.n5541 GND.n3290 0.152939
R14481 GND.n5542 GND.n5541 0.152939
R14482 GND.n5543 GND.n5542 0.152939
R14483 GND.n5544 GND.n5543 0.152939
R14484 GND.n5544 GND.n3270 0.152939
R14485 GND.n5569 GND.n3270 0.152939
R14486 GND.n5570 GND.n5569 0.152939
R14487 GND.n5571 GND.n5570 0.152939
R14488 GND.n5572 GND.n5571 0.152939
R14489 GND.n5573 GND.n5572 0.152939
R14490 GND.n5575 GND.n5573 0.152939
R14491 GND.n5575 GND.n5574 0.152939
R14492 GND.n5574 GND.n2909 0.152939
R14493 GND.n2910 GND.n2909 0.152939
R14494 GND.n2911 GND.n2910 0.152939
R14495 GND.n2925 GND.n2911 0.152939
R14496 GND.n2926 GND.n2925 0.152939
R14497 GND.n2927 GND.n2926 0.152939
R14498 GND.n2928 GND.n2927 0.152939
R14499 GND.n2943 GND.n2928 0.152939
R14500 GND.n2944 GND.n2943 0.152939
R14501 GND.n2945 GND.n2944 0.152939
R14502 GND.n2946 GND.n2945 0.152939
R14503 GND.n2961 GND.n2946 0.152939
R14504 GND.n2962 GND.n2961 0.152939
R14505 GND.n2963 GND.n2962 0.152939
R14506 GND.n2964 GND.n2963 0.152939
R14507 GND.n2979 GND.n2964 0.152939
R14508 GND.n2980 GND.n2979 0.152939
R14509 GND.n2981 GND.n2980 0.152939
R14510 GND.n2982 GND.n2981 0.152939
R14511 GND.n2996 GND.n2982 0.152939
R14512 GND.n2997 GND.n2996 0.152939
R14513 GND.n2998 GND.n2997 0.152939
R14514 GND.n2999 GND.n2998 0.152939
R14515 GND.n3014 GND.n2999 0.152939
R14516 GND.n3015 GND.n3014 0.152939
R14517 GND.n3016 GND.n3015 0.152939
R14518 GND.n3017 GND.n3016 0.152939
R14519 GND.n3031 GND.n3017 0.152939
R14520 GND.n3032 GND.n3031 0.152939
R14521 GND.n3033 GND.n3032 0.152939
R14522 GND.n3034 GND.n3033 0.152939
R14523 GND.n3040 GND.n3034 0.152939
R14524 GND.n3041 GND.n3040 0.152939
R14525 GND.n3042 GND.n3041 0.152939
R14526 GND.n3043 GND.n3042 0.152939
R14527 GND.n5996 GND.n3043 0.152939
R14528 GND.n5997 GND.n5996 0.152939
R14529 GND.n5998 GND.n5997 0.152939
R14530 GND.n5998 GND.n5992 0.152939
R14531 GND.n6004 GND.n5992 0.152939
R14532 GND.n6005 GND.n6004 0.152939
R14533 GND.n6006 GND.n6005 0.152939
R14534 GND.n6006 GND.n5988 0.152939
R14535 GND.n6012 GND.n5988 0.152939
R14536 GND.n6013 GND.n6012 0.152939
R14537 GND.n6014 GND.n6013 0.152939
R14538 GND.n6014 GND.n5984 0.152939
R14539 GND.n6020 GND.n5984 0.152939
R14540 GND.n6021 GND.n6020 0.152939
R14541 GND.n6022 GND.n6021 0.152939
R14542 GND.n6022 GND.n5980 0.152939
R14543 GND.n6028 GND.n5980 0.152939
R14544 GND.n6029 GND.n6028 0.152939
R14545 GND.n6030 GND.n6029 0.152939
R14546 GND.n2419 GND.n2025 0.152939
R14547 GND.n2442 GND.n2025 0.152939
R14548 GND.n2443 GND.n2442 0.152939
R14549 GND.n2444 GND.n2443 0.152939
R14550 GND.n2445 GND.n2444 0.152939
R14551 GND.n2445 GND.n2004 0.152939
R14552 GND.n2471 GND.n2004 0.152939
R14553 GND.n2472 GND.n2471 0.152939
R14554 GND.n2473 GND.n2472 0.152939
R14555 GND.n2473 GND.n1973 0.152939
R14556 GND.n2504 GND.n1973 0.152939
R14557 GND.n2505 GND.n2504 0.152939
R14558 GND.n2506 GND.n2505 0.152939
R14559 GND.n2507 GND.n2506 0.152939
R14560 GND.n2507 GND.n1387 0.152939
R14561 GND.n7041 GND.n1387 0.152939
R14562 GND.n1248 GND.n1247 0.152939
R14563 GND.n1249 GND.n1248 0.152939
R14564 GND.n1250 GND.n1249 0.152939
R14565 GND.n1251 GND.n1250 0.152939
R14566 GND.n1252 GND.n1251 0.152939
R14567 GND.n1253 GND.n1252 0.152939
R14568 GND.n1254 GND.n1253 0.152939
R14569 GND.n1255 GND.n1254 0.152939
R14570 GND.n1256 GND.n1255 0.152939
R14571 GND.n1259 GND.n1256 0.152939
R14572 GND.n1260 GND.n1259 0.152939
R14573 GND.n1261 GND.n1260 0.152939
R14574 GND.n1262 GND.n1261 0.152939
R14575 GND.n1263 GND.n1262 0.152939
R14576 GND.n1264 GND.n1263 0.152939
R14577 GND.n1265 GND.n1264 0.152939
R14578 GND.n1266 GND.n1265 0.152939
R14579 GND.n1267 GND.n1266 0.152939
R14580 GND.n1268 GND.n1267 0.152939
R14581 GND.n1270 GND.n1268 0.152939
R14582 GND.n1273 GND.n1270 0.152939
R14583 GND.n1274 GND.n1273 0.152939
R14584 GND.n1275 GND.n1274 0.152939
R14585 GND.n1276 GND.n1275 0.152939
R14586 GND.n1277 GND.n1276 0.152939
R14587 GND.n1278 GND.n1277 0.152939
R14588 GND.n1279 GND.n1278 0.152939
R14589 GND.n1280 GND.n1279 0.152939
R14590 GND.n1281 GND.n1280 0.152939
R14591 GND.n7119 GND.n1281 0.152939
R14592 GND.n7119 GND.n7118 0.152939
R14593 GND.n7118 GND.n7117 0.152939
R14594 GND.n2170 GND.n2169 0.152939
R14595 GND.n2170 GND.n2148 0.152939
R14596 GND.n2272 GND.n2148 0.152939
R14597 GND.n2273 GND.n2272 0.152939
R14598 GND.n2274 GND.n2273 0.152939
R14599 GND.n2275 GND.n2274 0.152939
R14600 GND.n2275 GND.n2125 0.152939
R14601 GND.n2296 GND.n2125 0.152939
R14602 GND.n2297 GND.n2296 0.152939
R14603 GND.n2298 GND.n2297 0.152939
R14604 GND.n2299 GND.n2298 0.152939
R14605 GND.n2299 GND.n2102 0.152939
R14606 GND.n2321 GND.n2102 0.152939
R14607 GND.n2322 GND.n2321 0.152939
R14608 GND.n2323 GND.n2322 0.152939
R14609 GND.n2323 GND.n2047 0.152939
R14610 GND.n7224 GND.n1180 0.152939
R14611 GND.n1185 GND.n1180 0.152939
R14612 GND.n1186 GND.n1185 0.152939
R14613 GND.n1187 GND.n1186 0.152939
R14614 GND.n1192 GND.n1187 0.152939
R14615 GND.n1193 GND.n1192 0.152939
R14616 GND.n1194 GND.n1193 0.152939
R14617 GND.n1195 GND.n1194 0.152939
R14618 GND.n1200 GND.n1195 0.152939
R14619 GND.n1201 GND.n1200 0.152939
R14620 GND.n1202 GND.n1201 0.152939
R14621 GND.n1203 GND.n1202 0.152939
R14622 GND.n1208 GND.n1203 0.152939
R14623 GND.n1209 GND.n1208 0.152939
R14624 GND.n1210 GND.n1209 0.152939
R14625 GND.n1211 GND.n1210 0.152939
R14626 GND.n1216 GND.n1211 0.152939
R14627 GND.n1217 GND.n1216 0.152939
R14628 GND.n1218 GND.n1217 0.152939
R14629 GND.n1219 GND.n1218 0.152939
R14630 GND.n2162 GND.n1219 0.152939
R14631 GND.n2163 GND.n2162 0.152939
R14632 GND.n2164 GND.n2163 0.152939
R14633 GND.n2164 GND.n2158 0.152939
R14634 GND.n2221 GND.n2158 0.152939
R14635 GND.n2222 GND.n2221 0.152939
R14636 GND.n2223 GND.n2222 0.152939
R14637 GND.n2224 GND.n2223 0.152939
R14638 GND.n2225 GND.n2224 0.152939
R14639 GND.n2228 GND.n2225 0.152939
R14640 GND.n2229 GND.n2228 0.152939
R14641 GND.n2230 GND.n2229 0.152939
R14642 GND.n2231 GND.n2230 0.152939
R14643 GND.n2234 GND.n2231 0.152939
R14644 GND.n2235 GND.n2234 0.152939
R14645 GND.n2236 GND.n2235 0.152939
R14646 GND.n2237 GND.n2236 0.152939
R14647 GND.n2240 GND.n2237 0.152939
R14648 GND.n2241 GND.n2240 0.152939
R14649 GND.n7371 GND.n1037 0.152939
R14650 GND.n1042 GND.n1037 0.152939
R14651 GND.n1043 GND.n1042 0.152939
R14652 GND.n1044 GND.n1043 0.152939
R14653 GND.n1045 GND.n1044 0.152939
R14654 GND.n1050 GND.n1045 0.152939
R14655 GND.n1051 GND.n1050 0.152939
R14656 GND.n1052 GND.n1051 0.152939
R14657 GND.n1053 GND.n1052 0.152939
R14658 GND.n1058 GND.n1053 0.152939
R14659 GND.n1059 GND.n1058 0.152939
R14660 GND.n1060 GND.n1059 0.152939
R14661 GND.n1061 GND.n1060 0.152939
R14662 GND.n1066 GND.n1061 0.152939
R14663 GND.n1067 GND.n1066 0.152939
R14664 GND.n1068 GND.n1067 0.152939
R14665 GND.n1069 GND.n1068 0.152939
R14666 GND.n1074 GND.n1069 0.152939
R14667 GND.n1075 GND.n1074 0.152939
R14668 GND.n1076 GND.n1075 0.152939
R14669 GND.n1077 GND.n1076 0.152939
R14670 GND.n1082 GND.n1077 0.152939
R14671 GND.n1083 GND.n1082 0.152939
R14672 GND.n1084 GND.n1083 0.152939
R14673 GND.n1085 GND.n1084 0.152939
R14674 GND.n1090 GND.n1085 0.152939
R14675 GND.n1091 GND.n1090 0.152939
R14676 GND.n1092 GND.n1091 0.152939
R14677 GND.n1093 GND.n1092 0.152939
R14678 GND.n1098 GND.n1093 0.152939
R14679 GND.n1099 GND.n1098 0.152939
R14680 GND.n1100 GND.n1099 0.152939
R14681 GND.n1101 GND.n1100 0.152939
R14682 GND.n1106 GND.n1101 0.152939
R14683 GND.n1107 GND.n1106 0.152939
R14684 GND.n1108 GND.n1107 0.152939
R14685 GND.n1109 GND.n1108 0.152939
R14686 GND.n1114 GND.n1109 0.152939
R14687 GND.n1115 GND.n1114 0.152939
R14688 GND.n1116 GND.n1115 0.152939
R14689 GND.n1117 GND.n1116 0.152939
R14690 GND.n1122 GND.n1117 0.152939
R14691 GND.n1123 GND.n1122 0.152939
R14692 GND.n1124 GND.n1123 0.152939
R14693 GND.n1125 GND.n1124 0.152939
R14694 GND.n1130 GND.n1125 0.152939
R14695 GND.n1131 GND.n1130 0.152939
R14696 GND.n1132 GND.n1131 0.152939
R14697 GND.n1133 GND.n1132 0.152939
R14698 GND.n1138 GND.n1133 0.152939
R14699 GND.n1139 GND.n1138 0.152939
R14700 GND.n1140 GND.n1139 0.152939
R14701 GND.n1141 GND.n1140 0.152939
R14702 GND.n1146 GND.n1141 0.152939
R14703 GND.n1147 GND.n1146 0.152939
R14704 GND.n1148 GND.n1147 0.152939
R14705 GND.n1149 GND.n1148 0.152939
R14706 GND.n1154 GND.n1149 0.152939
R14707 GND.n1155 GND.n1154 0.152939
R14708 GND.n1156 GND.n1155 0.152939
R14709 GND.n1157 GND.n1156 0.152939
R14710 GND.n1162 GND.n1157 0.152939
R14711 GND.n1163 GND.n1162 0.152939
R14712 GND.n1164 GND.n1163 0.152939
R14713 GND.n1165 GND.n1164 0.152939
R14714 GND.n1170 GND.n1165 0.152939
R14715 GND.n1171 GND.n1170 0.152939
R14716 GND.n1172 GND.n1171 0.152939
R14717 GND.n1173 GND.n1172 0.152939
R14718 GND.n1178 GND.n1173 0.152939
R14719 GND.n1179 GND.n1178 0.152939
R14720 GND.n7225 GND.n1179 0.152939
R14721 GND.n6857 GND.n6856 0.152939
R14722 GND.n6856 GND.n6855 0.152939
R14723 GND.n6855 GND.n2669 0.152939
R14724 GND.n6851 GND.n2669 0.152939
R14725 GND.n6851 GND.n6850 0.152939
R14726 GND.n6850 GND.n6849 0.152939
R14727 GND.n6849 GND.n2674 0.152939
R14728 GND.n6845 GND.n2674 0.152939
R14729 GND.n6845 GND.n6844 0.152939
R14730 GND.n6844 GND.n6843 0.152939
R14731 GND.n6843 GND.n2679 0.152939
R14732 GND.n6839 GND.n2679 0.152939
R14733 GND.n6839 GND.n6838 0.152939
R14734 GND.n6838 GND.n6837 0.152939
R14735 GND.n6837 GND.n2684 0.152939
R14736 GND.n6833 GND.n2684 0.152939
R14737 GND.n6833 GND.n6832 0.152939
R14738 GND.n6832 GND.n6831 0.152939
R14739 GND.n6831 GND.n2689 0.152939
R14740 GND.n6827 GND.n2689 0.152939
R14741 GND.n6827 GND.n6826 0.152939
R14742 GND.n6826 GND.n6825 0.152939
R14743 GND.n6825 GND.n2694 0.152939
R14744 GND.n6821 GND.n2694 0.152939
R14745 GND.n6821 GND.n6820 0.152939
R14746 GND.n6820 GND.n6819 0.152939
R14747 GND.n6819 GND.n2699 0.152939
R14748 GND.n6815 GND.n2699 0.152939
R14749 GND.n6815 GND.n6814 0.152939
R14750 GND.n6814 GND.n6813 0.152939
R14751 GND.n6813 GND.n2704 0.152939
R14752 GND.n6809 GND.n2704 0.152939
R14753 GND.n6809 GND.n6808 0.152939
R14754 GND.n6808 GND.n6807 0.152939
R14755 GND.n6807 GND.n2709 0.152939
R14756 GND.n6803 GND.n2709 0.152939
R14757 GND.n6803 GND.n6802 0.152939
R14758 GND.n6802 GND.n6801 0.152939
R14759 GND.n6801 GND.n2714 0.152939
R14760 GND.n6797 GND.n2714 0.152939
R14761 GND.n6797 GND.n6796 0.152939
R14762 GND.n6796 GND.n6795 0.152939
R14763 GND.n6795 GND.n2719 0.152939
R14764 GND.n6791 GND.n2719 0.152939
R14765 GND.n6791 GND.n6790 0.152939
R14766 GND.n6790 GND.n6789 0.152939
R14767 GND.n6789 GND.n2724 0.152939
R14768 GND.n6785 GND.n2724 0.152939
R14769 GND.n6785 GND.n6784 0.152939
R14770 GND.n6784 GND.n6783 0.152939
R14771 GND.n6783 GND.n2729 0.152939
R14772 GND.n6779 GND.n2729 0.152939
R14773 GND.n6779 GND.n6778 0.152939
R14774 GND.n6778 GND.n6777 0.152939
R14775 GND.n6777 GND.n2734 0.152939
R14776 GND.n6773 GND.n2734 0.152939
R14777 GND.n6773 GND.n6772 0.152939
R14778 GND.n6772 GND.n6771 0.152939
R14779 GND.n6771 GND.n2739 0.152939
R14780 GND.n6767 GND.n2739 0.152939
R14781 GND.n6767 GND.n6766 0.152939
R14782 GND.n6766 GND.n6765 0.152939
R14783 GND.n6765 GND.n2744 0.152939
R14784 GND.n6761 GND.n2744 0.152939
R14785 GND.n6761 GND.n6760 0.152939
R14786 GND.n6760 GND.n6759 0.152939
R14787 GND.n6759 GND.n2749 0.152939
R14788 GND.n6755 GND.n2749 0.152939
R14789 GND.n6755 GND.n6754 0.152939
R14790 GND.n6754 GND.n6753 0.152939
R14791 GND.n6753 GND.n2754 0.152939
R14792 GND.n6749 GND.n2754 0.152939
R14793 GND.n6749 GND.n6748 0.152939
R14794 GND.n6748 GND.n6747 0.152939
R14795 GND.n6747 GND.n2759 0.152939
R14796 GND.n6743 GND.n2759 0.152939
R14797 GND.n6743 GND.n6742 0.152939
R14798 GND.n6742 GND.n6741 0.152939
R14799 GND.n6741 GND.n2764 0.152939
R14800 GND.n6737 GND.n2764 0.152939
R14801 GND.n6737 GND.n6736 0.152939
R14802 GND.n6736 GND.n6735 0.152939
R14803 GND.n6735 GND.n2769 0.152939
R14804 GND.n6731 GND.n2769 0.152939
R14805 GND.n6731 GND.n6730 0.152939
R14806 GND.n6730 GND.n6729 0.152939
R14807 GND.n6729 GND.n2774 0.152939
R14808 GND.n6725 GND.n2774 0.152939
R14809 GND.n6725 GND.n6724 0.152939
R14810 GND.n6724 GND.n6723 0.152939
R14811 GND.n6723 GND.n2779 0.152939
R14812 GND.n6719 GND.n2779 0.152939
R14813 GND.n6719 GND.n6718 0.152939
R14814 GND.n6718 GND.n6717 0.152939
R14815 GND.n6717 GND.n2784 0.152939
R14816 GND.n6713 GND.n2784 0.152939
R14817 GND.n6713 GND.n6712 0.152939
R14818 GND.n6712 GND.n6711 0.152939
R14819 GND.n6711 GND.n2789 0.152939
R14820 GND.n6707 GND.n2789 0.152939
R14821 GND.n6707 GND.n6706 0.152939
R14822 GND.n6706 GND.n6705 0.152939
R14823 GND.n6705 GND.n2794 0.152939
R14824 GND.n6701 GND.n2794 0.152939
R14825 GND.n6701 GND.n6700 0.152939
R14826 GND.n6700 GND.n6699 0.152939
R14827 GND.n6699 GND.n2799 0.152939
R14828 GND.n6695 GND.n2799 0.152939
R14829 GND.n6695 GND.n6694 0.152939
R14830 GND.n6694 GND.n6693 0.152939
R14831 GND.n6693 GND.n2804 0.152939
R14832 GND.n6689 GND.n2804 0.152939
R14833 GND.n6689 GND.n6688 0.152939
R14834 GND.n6688 GND.n6687 0.152939
R14835 GND.n6687 GND.n2809 0.152939
R14836 GND.n6683 GND.n2809 0.152939
R14837 GND.n6683 GND.n6682 0.152939
R14838 GND.n6682 GND.n6681 0.152939
R14839 GND.n6681 GND.n2814 0.152939
R14840 GND.n6677 GND.n2814 0.152939
R14841 GND.n6677 GND.n6676 0.152939
R14842 GND.n6676 GND.n6675 0.152939
R14843 GND.n6675 GND.n2819 0.152939
R14844 GND.n6671 GND.n2819 0.152939
R14845 GND.n6671 GND.n6670 0.152939
R14846 GND.n6670 GND.n6669 0.152939
R14847 GND.n6669 GND.n2824 0.152939
R14848 GND.n6665 GND.n2824 0.152939
R14849 GND.n6664 GND.n2828 0.152939
R14850 GND.n6660 GND.n6659 0.152939
R14851 GND.n6659 GND.n6658 0.152939
R14852 GND.n6658 GND.n2873 0.152939
R14853 GND.n6654 GND.n2873 0.152939
R14854 GND.n6654 GND.n6653 0.152939
R14855 GND.n6653 GND.n6652 0.152939
R14856 GND.n6652 GND.n2878 0.152939
R14857 GND.n6648 GND.n2878 0.152939
R14858 GND.n6648 GND.n6647 0.152939
R14859 GND.n6647 GND.n6646 0.152939
R14860 GND.n6646 GND.n2883 0.152939
R14861 GND.n6642 GND.n2883 0.152939
R14862 GND.n6642 GND.n6641 0.152939
R14863 GND.n6641 GND.n6640 0.152939
R14864 GND.n6640 GND.n2888 0.152939
R14865 GND.n6636 GND.n2888 0.152939
R14866 GND.n6636 GND.n6635 0.152939
R14867 GND.n6635 GND.n2895 0.152939
R14868 GND.n6631 GND.n2895 0.152939
R14869 GND.n6631 GND.n6630 0.152939
R14870 GND.n4336 GND.n4322 0.152939
R14871 GND.n4336 GND.n4335 0.152939
R14872 GND.n4335 GND.n4334 0.152939
R14873 GND.n4334 GND.n4323 0.152939
R14874 GND.n4330 GND.n4323 0.152939
R14875 GND.n4330 GND.n4329 0.152939
R14876 GND.n4329 GND.n3857 0.152939
R14877 GND.n4420 GND.n3857 0.152939
R14878 GND.n4421 GND.n4420 0.152939
R14879 GND.n4432 GND.n4421 0.152939
R14880 GND.n4432 GND.n4431 0.152939
R14881 GND.n4431 GND.n4430 0.152939
R14882 GND.n4430 GND.n4422 0.152939
R14883 GND.n4426 GND.n4422 0.152939
R14884 GND.n4426 GND.n3817 0.152939
R14885 GND.n4497 GND.n3817 0.152939
R14886 GND.n4498 GND.n4497 0.152939
R14887 GND.n4509 GND.n4498 0.152939
R14888 GND.n4509 GND.n4508 0.152939
R14889 GND.n4508 GND.n4507 0.152939
R14890 GND.n4507 GND.n4499 0.152939
R14891 GND.n4503 GND.n4499 0.152939
R14892 GND.n4503 GND.n3775 0.152939
R14893 GND.n4591 GND.n3775 0.152939
R14894 GND.n4592 GND.n4591 0.152939
R14895 GND.n4594 GND.n4592 0.152939
R14896 GND.n4594 GND.n4593 0.152939
R14897 GND.n4593 GND.n3745 0.152939
R14898 GND.n4630 GND.n3745 0.152939
R14899 GND.n4631 GND.n4630 0.152939
R14900 GND.n4667 GND.n4631 0.152939
R14901 GND.n4667 GND.n4666 0.152939
R14902 GND.n4666 GND.n4665 0.152939
R14903 GND.n4665 GND.n4632 0.152939
R14904 GND.n4661 GND.n4632 0.152939
R14905 GND.n4661 GND.n4660 0.152939
R14906 GND.n4660 GND.n4659 0.152939
R14907 GND.n4659 GND.n4637 0.152939
R14908 GND.n4655 GND.n4637 0.152939
R14909 GND.n4655 GND.n4654 0.152939
R14910 GND.n4654 GND.n4653 0.152939
R14911 GND.n4653 GND.n4641 0.152939
R14912 GND.n4649 GND.n4641 0.152939
R14913 GND.n4649 GND.n4648 0.152939
R14914 GND.n4648 GND.n3657 0.152939
R14915 GND.n4806 GND.n3657 0.152939
R14916 GND.n4807 GND.n4806 0.152939
R14917 GND.n4843 GND.n4807 0.152939
R14918 GND.n4843 GND.n4842 0.152939
R14919 GND.n4842 GND.n4841 0.152939
R14920 GND.n4841 GND.n4808 0.152939
R14921 GND.n4837 GND.n4808 0.152939
R14922 GND.n4837 GND.n4836 0.152939
R14923 GND.n4836 GND.n4835 0.152939
R14924 GND.n4835 GND.n4813 0.152939
R14925 GND.n4831 GND.n4813 0.152939
R14926 GND.n4831 GND.n4830 0.152939
R14927 GND.n4830 GND.n4829 0.152939
R14928 GND.n4829 GND.n4817 0.152939
R14929 GND.n4825 GND.n4817 0.152939
R14930 GND.n4825 GND.n4824 0.152939
R14931 GND.n4824 GND.n3569 0.152939
R14932 GND.n4982 GND.n3569 0.152939
R14933 GND.n4983 GND.n4982 0.152939
R14934 GND.n5019 GND.n4983 0.152939
R14935 GND.n5019 GND.n5018 0.152939
R14936 GND.n5018 GND.n5017 0.152939
R14937 GND.n5017 GND.n4984 0.152939
R14938 GND.n5013 GND.n4984 0.152939
R14939 GND.n5013 GND.n5012 0.152939
R14940 GND.n5012 GND.n5011 0.152939
R14941 GND.n5011 GND.n4989 0.152939
R14942 GND.n5007 GND.n4989 0.152939
R14943 GND.n5007 GND.n5006 0.152939
R14944 GND.n5006 GND.n5005 0.152939
R14945 GND.n5005 GND.n4993 0.152939
R14946 GND.n5001 GND.n4993 0.152939
R14947 GND.n5001 GND.n5000 0.152939
R14948 GND.n5000 GND.n3480 0.152939
R14949 GND.n5158 GND.n3480 0.152939
R14950 GND.n5159 GND.n5158 0.152939
R14951 GND.n5195 GND.n5159 0.152939
R14952 GND.n5195 GND.n5194 0.152939
R14953 GND.n5194 GND.n5193 0.152939
R14954 GND.n5193 GND.n5160 0.152939
R14955 GND.n5189 GND.n5160 0.152939
R14956 GND.n5189 GND.n5188 0.152939
R14957 GND.n5188 GND.n5187 0.152939
R14958 GND.n5187 GND.n5165 0.152939
R14959 GND.n5183 GND.n5165 0.152939
R14960 GND.n5183 GND.n5182 0.152939
R14961 GND.n5182 GND.n5181 0.152939
R14962 GND.n5181 GND.n5169 0.152939
R14963 GND.n5177 GND.n5169 0.152939
R14964 GND.n5177 GND.n5176 0.152939
R14965 GND.n5176 GND.n3391 0.152939
R14966 GND.n5333 GND.n3391 0.152939
R14967 GND.n5334 GND.n5333 0.152939
R14968 GND.n5372 GND.n5334 0.152939
R14969 GND.n5372 GND.n5371 0.152939
R14970 GND.n5371 GND.n5370 0.152939
R14971 GND.n5370 GND.n5335 0.152939
R14972 GND.n5366 GND.n5335 0.152939
R14973 GND.n5366 GND.n5365 0.152939
R14974 GND.n5365 GND.n5364 0.152939
R14975 GND.n5364 GND.n5342 0.152939
R14976 GND.n5360 GND.n5342 0.152939
R14977 GND.n5360 GND.n5359 0.152939
R14978 GND.n5359 GND.n5358 0.152939
R14979 GND.n5358 GND.n5346 0.152939
R14980 GND.n5354 GND.n5346 0.152939
R14981 GND.n5354 GND.n5353 0.152939
R14982 GND.n5353 GND.n3305 0.152939
R14983 GND.n5511 GND.n3305 0.152939
R14984 GND.n5512 GND.n5511 0.152939
R14985 GND.n5525 GND.n5512 0.152939
R14986 GND.n5525 GND.n5524 0.152939
R14987 GND.n5524 GND.n5523 0.152939
R14988 GND.n5523 GND.n5513 0.152939
R14989 GND.n5519 GND.n5513 0.152939
R14990 GND.n5519 GND.n5518 0.152939
R14991 GND.n5518 GND.n3255 0.152939
R14992 GND.n5605 GND.n3255 0.152939
R14993 GND.n5606 GND.n5605 0.152939
R14994 GND.n5608 GND.n5606 0.152939
R14995 GND.n5608 GND.n5607 0.152939
R14996 GND.n5607 GND.n2900 0.152939
R14997 GND.n6629 GND.n2900 0.152939
R14998 GND.n4313 GND.n2668 0.152939
R14999 GND.n4272 GND.n4271 0.152939
R15000 GND.n4271 GND.n4215 0.152939
R15001 GND.n4267 GND.n4215 0.152939
R15002 GND.n4267 GND.n4266 0.152939
R15003 GND.n4266 GND.n4265 0.152939
R15004 GND.n4265 GND.n4220 0.152939
R15005 GND.n4261 GND.n4220 0.152939
R15006 GND.n4261 GND.n4260 0.152939
R15007 GND.n4260 GND.n4259 0.152939
R15008 GND.n4259 GND.n4226 0.152939
R15009 GND.n4255 GND.n4226 0.152939
R15010 GND.n4255 GND.n4254 0.152939
R15011 GND.n4254 GND.n4253 0.152939
R15012 GND.n4253 GND.n4232 0.152939
R15013 GND.n4249 GND.n4232 0.152939
R15014 GND.n4249 GND.n4248 0.152939
R15015 GND.n4248 GND.n4247 0.152939
R15016 GND.n4247 GND.n4238 0.152939
R15017 GND.n4238 GND.n3902 0.152939
R15018 GND.n4321 GND.n3902 0.152939
R15019 GND.n7040 GND.n1388 0.152939
R15020 GND.n7036 GND.n1388 0.152939
R15021 GND.n7036 GND.n7035 0.152939
R15022 GND.n7035 GND.n7034 0.152939
R15023 GND.n7034 GND.n1392 0.152939
R15024 GND.n7030 GND.n1392 0.152939
R15025 GND.n7030 GND.n7029 0.152939
R15026 GND.n7029 GND.n7028 0.152939
R15027 GND.n7028 GND.n1397 0.152939
R15028 GND.n7024 GND.n1397 0.152939
R15029 GND.n7024 GND.n7023 0.152939
R15030 GND.n7023 GND.n7022 0.152939
R15031 GND.n7018 GND.n7017 0.152939
R15032 GND.n7017 GND.n7016 0.152939
R15033 GND.n7016 GND.n1410 0.152939
R15034 GND.n7012 GND.n1410 0.152939
R15035 GND.n7012 GND.n7011 0.152939
R15036 GND.n7011 GND.n7010 0.152939
R15037 GND.n7010 GND.n1417 0.152939
R15038 GND.n7006 GND.n1417 0.152939
R15039 GND.n7006 GND.n7005 0.152939
R15040 GND.n7005 GND.n7004 0.152939
R15041 GND.n7004 GND.n1422 0.152939
R15042 GND.n7000 GND.n1422 0.152939
R15043 GND.n7000 GND.n6999 0.152939
R15044 GND.n6999 GND.n6998 0.152939
R15045 GND.n6998 GND.n1427 0.152939
R15046 GND.n1432 GND.n1427 0.152939
R15047 GND.n6993 GND.n1432 0.152939
R15048 GND.n2189 GND.n2188 0.152939
R15049 GND.n2195 GND.n2188 0.152939
R15050 GND.n2196 GND.n2195 0.152939
R15051 GND.n2197 GND.n2196 0.152939
R15052 GND.n2197 GND.n2184 0.152939
R15053 GND.n2203 GND.n2184 0.152939
R15054 GND.n2204 GND.n2203 0.152939
R15055 GND.n2205 GND.n2204 0.152939
R15056 GND.n2205 GND.n2177 0.152939
R15057 GND.n2209 GND.n2177 0.152939
R15058 GND.n2212 GND.n2211 0.152939
R15059 GND.n2214 GND.n2212 0.152939
R15060 GND.n2214 GND.n2213 0.152939
R15061 GND.n2213 GND.n2138 0.152939
R15062 GND.n2282 GND.n2138 0.152939
R15063 GND.n2283 GND.n2282 0.152939
R15064 GND.n2285 GND.n2283 0.152939
R15065 GND.n2285 GND.n2284 0.152939
R15066 GND.n2284 GND.n2114 0.152939
R15067 GND.n2306 GND.n2114 0.152939
R15068 GND.n2307 GND.n2306 0.152939
R15069 GND.n2309 GND.n2307 0.152939
R15070 GND.n2309 GND.n2308 0.152939
R15071 GND.n2308 GND.n2091 0.152939
R15072 GND.n2329 GND.n2091 0.152939
R15073 GND.n2330 GND.n2329 0.152939
R15074 GND.n2331 GND.n2330 0.152939
R15075 GND.n2331 GND.n2089 0.152939
R15076 GND.n2337 GND.n2089 0.152939
R15077 GND.n2338 GND.n2337 0.152939
R15078 GND.n2339 GND.n2338 0.152939
R15079 GND.n5949 GND.n151 0.14989
R15080 GND.n2241 GND.n2048 0.14989
R15081 GND.n2872 GND.n2828 0.142268
R15082 GND.n4313 GND.n4312 0.142268
R15083 GND.n1875 GND.n1437 0.112242
R15084 GND.n8504 GND.n149 0.0767195
R15085 GND.n8504 GND.n150 0.0767195
R15086 GND.n2419 GND.n2418 0.0767195
R15087 GND.n2418 GND.n2047 0.0767195
R15088 GND.n2342 GND.n2087 0.0695946
R15089 GND.n8512 GND.n136 0.0695946
R15090 GND.n8512 GND.n8511 0.0695946
R15091 GND.n2339 GND.n2087 0.0695946
R15092 GND.n6133 GND.n5816 0.063
R15093 GND.n6992 GND.n6991 0.063
R15094 GND.n6133 GND.n6106 0.0541717
R15095 GND.n6991 GND.n1916 0.0541717
R15096 GND.n5824 GND.n5816 0.046356
R15097 GND.n8449 GND.n249 0.046356
R15098 GND.n7110 GND.n1287 0.046356
R15099 GND.n6992 GND.n1378 0.046356
R15100 GND.n1875 GND.n1874 0.0455581
R15101 GND.n6444 GND.n5824 0.0344674
R15102 GND.n6444 GND.n5826 0.0344674
R15103 GND.n5851 GND.n5826 0.0344674
R15104 GND.n5852 GND.n5851 0.0344674
R15105 GND.n5853 GND.n5852 0.0344674
R15106 GND.n5854 GND.n5853 0.0344674
R15107 GND.n6150 GND.n5854 0.0344674
R15108 GND.n6150 GND.n5873 0.0344674
R15109 GND.n5874 GND.n5873 0.0344674
R15110 GND.n5875 GND.n5874 0.0344674
R15111 GND.n6165 GND.n5875 0.0344674
R15112 GND.n6165 GND.n5894 0.0344674
R15113 GND.n5895 GND.n5894 0.0344674
R15114 GND.n5896 GND.n5895 0.0344674
R15115 GND.n6180 GND.n5896 0.0344674
R15116 GND.n6180 GND.n5913 0.0344674
R15117 GND.n5914 GND.n5913 0.0344674
R15118 GND.n5915 GND.n5914 0.0344674
R15119 GND.n6203 GND.n5915 0.0344674
R15120 GND.n6204 GND.n6203 0.0344674
R15121 GND.n6204 GND.n5936 0.0344674
R15122 GND.n5937 GND.n5936 0.0344674
R15123 GND.n5938 GND.n5937 0.0344674
R15124 GND.n6211 GND.n5938 0.0344674
R15125 GND.n6212 GND.n6211 0.0344674
R15126 GND.n6212 GND.n167 0.0344674
R15127 GND.n168 GND.n167 0.0344674
R15128 GND.n169 GND.n168 0.0344674
R15129 GND.n6227 GND.n169 0.0344674
R15130 GND.n6227 GND.n187 0.0344674
R15131 GND.n188 GND.n187 0.0344674
R15132 GND.n189 GND.n188 0.0344674
R15133 GND.n6243 GND.n189 0.0344674
R15134 GND.n6243 GND.n207 0.0344674
R15135 GND.n208 GND.n207 0.0344674
R15136 GND.n209 GND.n208 0.0344674
R15137 GND.n6246 GND.n209 0.0344674
R15138 GND.n6246 GND.n228 0.0344674
R15139 GND.n229 GND.n228 0.0344674
R15140 GND.n230 GND.n229 0.0344674
R15141 GND.n6253 GND.n230 0.0344674
R15142 GND.n6253 GND.n248 0.0344674
R15143 GND.n8449 GND.n248 0.0344674
R15144 GND.n7110 GND.n7109 0.0344674
R15145 GND.n7109 GND.n1296 0.0344674
R15146 GND.n7105 GND.n1296 0.0344674
R15147 GND.n7105 GND.n7104 0.0344674
R15148 GND.n7104 GND.n7103 0.0344674
R15149 GND.n7103 GND.n1303 0.0344674
R15150 GND.n7099 GND.n1303 0.0344674
R15151 GND.n7099 GND.n7098 0.0344674
R15152 GND.n7098 GND.n7097 0.0344674
R15153 GND.n7097 GND.n1311 0.0344674
R15154 GND.n7093 GND.n1311 0.0344674
R15155 GND.n7093 GND.n7092 0.0344674
R15156 GND.n7092 GND.n7091 0.0344674
R15157 GND.n7091 GND.n1319 0.0344674
R15158 GND.n7087 GND.n1319 0.0344674
R15159 GND.n7087 GND.n7086 0.0344674
R15160 GND.n7086 GND.n7085 0.0344674
R15161 GND.n7085 GND.n1327 0.0344674
R15162 GND.n7081 GND.n1327 0.0344674
R15163 GND.n7081 GND.n7080 0.0344674
R15164 GND.n7080 GND.n7079 0.0344674
R15165 GND.n7079 GND.n1335 0.0344674
R15166 GND.n7075 GND.n1335 0.0344674
R15167 GND.n7075 GND.n7074 0.0344674
R15168 GND.n7074 GND.n7073 0.0344674
R15169 GND.n7073 GND.n1343 0.0344674
R15170 GND.n7069 GND.n1343 0.0344674
R15171 GND.n7069 GND.n7068 0.0344674
R15172 GND.n7068 GND.n7067 0.0344674
R15173 GND.n7067 GND.n1351 0.0344674
R15174 GND.n7063 GND.n1351 0.0344674
R15175 GND.n7063 GND.n7062 0.0344674
R15176 GND.n7062 GND.n7061 0.0344674
R15177 GND.n7061 GND.n1359 0.0344674
R15178 GND.n7057 GND.n1359 0.0344674
R15179 GND.n7057 GND.n7056 0.0344674
R15180 GND.n7056 GND.n7055 0.0344674
R15181 GND.n7055 GND.n1367 0.0344674
R15182 GND.n7051 GND.n1367 0.0344674
R15183 GND.n7051 GND.n7050 0.0344674
R15184 GND.n7050 GND.n7049 0.0344674
R15185 GND.n7049 GND.n1375 0.0344674
R15186 GND.n1378 GND.n1375 0.0344674
R15187 GND.n6660 GND.n2872 0.0111707
R15188 GND.n4312 GND.n4272 0.0111707
R15189 GND.n2361 GND.n2048 0.00354878
R15190 GND.n6030 GND.n151 0.00354878
R15191 CS_BIAS.n50 CS_BIAS.n44 289.615
R15192 CS_BIAS.n183 CS_BIAS.n177 289.615
R15193 CS_BIAS.n51 CS_BIAS.n50 185
R15194 CS_BIAS.n49 CS_BIAS.n48 185
R15195 CS_BIAS.n184 CS_BIAS.n183 185
R15196 CS_BIAS.n182 CS_BIAS.n181 185
R15197 CS_BIAS.n167 CS_BIAS.n132 161.3
R15198 CS_BIAS.n166 CS_BIAS.n165 161.3
R15199 CS_BIAS.n164 CS_BIAS.n133 161.3
R15200 CS_BIAS.n163 CS_BIAS.n162 161.3
R15201 CS_BIAS.n161 CS_BIAS.n134 161.3
R15202 CS_BIAS.n160 CS_BIAS.n159 161.3
R15203 CS_BIAS.n158 CS_BIAS.n157 161.3
R15204 CS_BIAS.n156 CS_BIAS.n136 161.3
R15205 CS_BIAS.n155 CS_BIAS.n154 161.3
R15206 CS_BIAS.n153 CS_BIAS.n137 161.3
R15207 CS_BIAS.n152 CS_BIAS.n151 161.3
R15208 CS_BIAS.n149 CS_BIAS.n138 161.3
R15209 CS_BIAS.n148 CS_BIAS.n147 161.3
R15210 CS_BIAS.n146 CS_BIAS.n139 161.3
R15211 CS_BIAS.n145 CS_BIAS.n144 161.3
R15212 CS_BIAS.n143 CS_BIAS.n140 161.3
R15213 CS_BIAS.n104 CS_BIAS.n101 161.3
R15214 CS_BIAS.n106 CS_BIAS.n105 161.3
R15215 CS_BIAS.n107 CS_BIAS.n100 161.3
R15216 CS_BIAS.n109 CS_BIAS.n108 161.3
R15217 CS_BIAS.n110 CS_BIAS.n99 161.3
R15218 CS_BIAS.n113 CS_BIAS.n112 161.3
R15219 CS_BIAS.n114 CS_BIAS.n98 161.3
R15220 CS_BIAS.n116 CS_BIAS.n115 161.3
R15221 CS_BIAS.n117 CS_BIAS.n97 161.3
R15222 CS_BIAS.n119 CS_BIAS.n118 161.3
R15223 CS_BIAS.n121 CS_BIAS.n120 161.3
R15224 CS_BIAS.n122 CS_BIAS.n95 161.3
R15225 CS_BIAS.n124 CS_BIAS.n123 161.3
R15226 CS_BIAS.n125 CS_BIAS.n94 161.3
R15227 CS_BIAS.n127 CS_BIAS.n126 161.3
R15228 CS_BIAS.n128 CS_BIAS.n93 161.3
R15229 CS_BIAS.n17 CS_BIAS.n14 161.3
R15230 CS_BIAS.n19 CS_BIAS.n18 161.3
R15231 CS_BIAS.n20 CS_BIAS.n13 161.3
R15232 CS_BIAS.n22 CS_BIAS.n21 161.3
R15233 CS_BIAS.n23 CS_BIAS.n12 161.3
R15234 CS_BIAS.n26 CS_BIAS.n25 161.3
R15235 CS_BIAS.n27 CS_BIAS.n11 161.3
R15236 CS_BIAS.n29 CS_BIAS.n28 161.3
R15237 CS_BIAS.n30 CS_BIAS.n10 161.3
R15238 CS_BIAS.n32 CS_BIAS.n31 161.3
R15239 CS_BIAS.n34 CS_BIAS.n33 161.3
R15240 CS_BIAS.n35 CS_BIAS.n8 161.3
R15241 CS_BIAS.n37 CS_BIAS.n36 161.3
R15242 CS_BIAS.n38 CS_BIAS.n7 161.3
R15243 CS_BIAS.n40 CS_BIAS.n39 161.3
R15244 CS_BIAS.n41 CS_BIAS.n6 161.3
R15245 CS_BIAS.n66 CS_BIAS.n65 161.3
R15246 CS_BIAS.n67 CS_BIAS.n62 161.3
R15247 CS_BIAS.n69 CS_BIAS.n68 161.3
R15248 CS_BIAS.n70 CS_BIAS.n61 161.3
R15249 CS_BIAS.n72 CS_BIAS.n71 161.3
R15250 CS_BIAS.n75 CS_BIAS.n74 161.3
R15251 CS_BIAS.n76 CS_BIAS.n5 161.3
R15252 CS_BIAS.n78 CS_BIAS.n77 161.3
R15253 CS_BIAS.n79 CS_BIAS.n4 161.3
R15254 CS_BIAS.n81 CS_BIAS.n80 161.3
R15255 CS_BIAS.n83 CS_BIAS.n82 161.3
R15256 CS_BIAS.n84 CS_BIAS.n2 161.3
R15257 CS_BIAS.n86 CS_BIAS.n85 161.3
R15258 CS_BIAS.n87 CS_BIAS.n1 161.3
R15259 CS_BIAS.n89 CS_BIAS.n88 161.3
R15260 CS_BIAS.n90 CS_BIAS.n0 161.3
R15261 CS_BIAS.n338 CS_BIAS.n303 161.3
R15262 CS_BIAS.n337 CS_BIAS.n336 161.3
R15263 CS_BIAS.n335 CS_BIAS.n304 161.3
R15264 CS_BIAS.n334 CS_BIAS.n333 161.3
R15265 CS_BIAS.n332 CS_BIAS.n305 161.3
R15266 CS_BIAS.n331 CS_BIAS.n330 161.3
R15267 CS_BIAS.n329 CS_BIAS.n328 161.3
R15268 CS_BIAS.n327 CS_BIAS.n307 161.3
R15269 CS_BIAS.n326 CS_BIAS.n325 161.3
R15270 CS_BIAS.n324 CS_BIAS.n308 161.3
R15271 CS_BIAS.n323 CS_BIAS.n322 161.3
R15272 CS_BIAS.n320 CS_BIAS.n309 161.3
R15273 CS_BIAS.n319 CS_BIAS.n318 161.3
R15274 CS_BIAS.n317 CS_BIAS.n310 161.3
R15275 CS_BIAS.n316 CS_BIAS.n315 161.3
R15276 CS_BIAS.n314 CS_BIAS.n311 161.3
R15277 CS_BIAS.n299 CS_BIAS.n264 161.3
R15278 CS_BIAS.n298 CS_BIAS.n297 161.3
R15279 CS_BIAS.n296 CS_BIAS.n265 161.3
R15280 CS_BIAS.n295 CS_BIAS.n294 161.3
R15281 CS_BIAS.n293 CS_BIAS.n266 161.3
R15282 CS_BIAS.n292 CS_BIAS.n291 161.3
R15283 CS_BIAS.n290 CS_BIAS.n289 161.3
R15284 CS_BIAS.n288 CS_BIAS.n268 161.3
R15285 CS_BIAS.n287 CS_BIAS.n286 161.3
R15286 CS_BIAS.n285 CS_BIAS.n269 161.3
R15287 CS_BIAS.n284 CS_BIAS.n283 161.3
R15288 CS_BIAS.n281 CS_BIAS.n270 161.3
R15289 CS_BIAS.n280 CS_BIAS.n279 161.3
R15290 CS_BIAS.n278 CS_BIAS.n271 161.3
R15291 CS_BIAS.n277 CS_BIAS.n276 161.3
R15292 CS_BIAS.n275 CS_BIAS.n272 161.3
R15293 CS_BIAS.n225 CS_BIAS.n190 161.3
R15294 CS_BIAS.n224 CS_BIAS.n223 161.3
R15295 CS_BIAS.n222 CS_BIAS.n191 161.3
R15296 CS_BIAS.n221 CS_BIAS.n220 161.3
R15297 CS_BIAS.n219 CS_BIAS.n192 161.3
R15298 CS_BIAS.n218 CS_BIAS.n217 161.3
R15299 CS_BIAS.n216 CS_BIAS.n215 161.3
R15300 CS_BIAS.n214 CS_BIAS.n194 161.3
R15301 CS_BIAS.n213 CS_BIAS.n212 161.3
R15302 CS_BIAS.n211 CS_BIAS.n195 161.3
R15303 CS_BIAS.n210 CS_BIAS.n209 161.3
R15304 CS_BIAS.n207 CS_BIAS.n196 161.3
R15305 CS_BIAS.n206 CS_BIAS.n205 161.3
R15306 CS_BIAS.n204 CS_BIAS.n197 161.3
R15307 CS_BIAS.n203 CS_BIAS.n202 161.3
R15308 CS_BIAS.n201 CS_BIAS.n198 161.3
R15309 CS_BIAS.n243 CS_BIAS.n242 161.3
R15310 CS_BIAS.n241 CS_BIAS.n232 161.3
R15311 CS_BIAS.n240 CS_BIAS.n239 161.3
R15312 CS_BIAS.n238 CS_BIAS.n233 161.3
R15313 CS_BIAS.n237 CS_BIAS.n236 161.3
R15314 CS_BIAS.n261 CS_BIAS.n171 161.3
R15315 CS_BIAS.n260 CS_BIAS.n259 161.3
R15316 CS_BIAS.n258 CS_BIAS.n172 161.3
R15317 CS_BIAS.n257 CS_BIAS.n256 161.3
R15318 CS_BIAS.n255 CS_BIAS.n173 161.3
R15319 CS_BIAS.n254 CS_BIAS.n253 161.3
R15320 CS_BIAS.n252 CS_BIAS.n251 161.3
R15321 CS_BIAS.n250 CS_BIAS.n175 161.3
R15322 CS_BIAS.n249 CS_BIAS.n248 161.3
R15323 CS_BIAS.n247 CS_BIAS.n176 161.3
R15324 CS_BIAS.n246 CS_BIAS.n245 161.3
R15325 CS_BIAS.n47 CS_BIAS.t3 153.582
R15326 CS_BIAS.n180 CS_BIAS.t9 153.582
R15327 CS_BIAS.n50 CS_BIAS.n49 104.615
R15328 CS_BIAS.n183 CS_BIAS.n182 104.615
R15329 CS_BIAS.n169 CS_BIAS.n168 103.416
R15330 CS_BIAS.n130 CS_BIAS.n129 103.416
R15331 CS_BIAS.n43 CS_BIAS.n42 103.416
R15332 CS_BIAS.n92 CS_BIAS.n91 103.416
R15333 CS_BIAS.n340 CS_BIAS.n339 103.416
R15334 CS_BIAS.n301 CS_BIAS.n300 103.416
R15335 CS_BIAS.n227 CS_BIAS.n226 103.416
R15336 CS_BIAS.n263 CS_BIAS.n262 103.416
R15337 CS_BIAS.n59 CS_BIAS.n58 103.194
R15338 CS_BIAS.n57 CS_BIAS.n56 102.322
R15339 CS_BIAS.n229 CS_BIAS.n228 102.322
R15340 CS_BIAS.n189 CS_BIAS.n188 102.322
R15341 CS_BIAS.n189 CS_BIAS.n187 65.931
R15342 CS_BIAS.n55 CS_BIAS.n54 64.7672
R15343 CS_BIAS.n141 CS_BIAS.t41 60.3741
R15344 CS_BIAS.n102 CS_BIAS.t22 60.3741
R15345 CS_BIAS.n15 CS_BIAS.t14 60.3741
R15346 CS_BIAS.n64 CS_BIAS.t28 60.3741
R15347 CS_BIAS.n312 CS_BIAS.t40 60.3741
R15348 CS_BIAS.n273 CS_BIAS.t29 60.3741
R15349 CS_BIAS.n199 CS_BIAS.t8 60.3741
R15350 CS_BIAS.n235 CS_BIAS.t24 60.3741
R15351 CS_BIAS.n162 CS_BIAS.n133 56.5193
R15352 CS_BIAS.n123 CS_BIAS.n94 56.5193
R15353 CS_BIAS.n36 CS_BIAS.n7 56.5193
R15354 CS_BIAS.n85 CS_BIAS.n1 56.5193
R15355 CS_BIAS.n333 CS_BIAS.n304 56.5193
R15356 CS_BIAS.n294 CS_BIAS.n265 56.5193
R15357 CS_BIAS.n220 CS_BIAS.n191 56.5193
R15358 CS_BIAS.n256 CS_BIAS.n172 56.5193
R15359 CS_BIAS.n49 CS_BIAS.t3 52.3082
R15360 CS_BIAS.n182 CS_BIAS.t9 52.3082
R15361 CS_BIAS.n142 CS_BIAS.n141 50.2654
R15362 CS_BIAS.n103 CS_BIAS.n102 50.2654
R15363 CS_BIAS.n16 CS_BIAS.n15 50.2654
R15364 CS_BIAS.n64 CS_BIAS.n63 50.2654
R15365 CS_BIAS.n313 CS_BIAS.n312 50.2654
R15366 CS_BIAS.n274 CS_BIAS.n273 50.2654
R15367 CS_BIAS.n200 CS_BIAS.n199 50.2654
R15368 CS_BIAS.n235 CS_BIAS.n234 50.2654
R15369 CS_BIAS.n144 CS_BIAS.n139 50.2061
R15370 CS_BIAS.n156 CS_BIAS.n155 50.2061
R15371 CS_BIAS.n117 CS_BIAS.n116 50.2061
R15372 CS_BIAS.n105 CS_BIAS.n100 50.2061
R15373 CS_BIAS.n30 CS_BIAS.n29 50.2061
R15374 CS_BIAS.n18 CS_BIAS.n13 50.2061
R15375 CS_BIAS.n79 CS_BIAS.n78 50.2061
R15376 CS_BIAS.n68 CS_BIAS.n67 50.2061
R15377 CS_BIAS.n315 CS_BIAS.n310 50.2061
R15378 CS_BIAS.n327 CS_BIAS.n326 50.2061
R15379 CS_BIAS.n276 CS_BIAS.n271 50.2061
R15380 CS_BIAS.n288 CS_BIAS.n287 50.2061
R15381 CS_BIAS.n202 CS_BIAS.n197 50.2061
R15382 CS_BIAS.n214 CS_BIAS.n213 50.2061
R15383 CS_BIAS.n250 CS_BIAS.n249 50.2061
R15384 CS_BIAS.n239 CS_BIAS.n238 50.2061
R15385 CS_BIAS.n148 CS_BIAS.n139 30.7807
R15386 CS_BIAS.n155 CS_BIAS.n137 30.7807
R15387 CS_BIAS.n116 CS_BIAS.n98 30.7807
R15388 CS_BIAS.n109 CS_BIAS.n100 30.7807
R15389 CS_BIAS.n29 CS_BIAS.n11 30.7807
R15390 CS_BIAS.n22 CS_BIAS.n13 30.7807
R15391 CS_BIAS.n78 CS_BIAS.n5 30.7807
R15392 CS_BIAS.n68 CS_BIAS.n61 30.7807
R15393 CS_BIAS.n319 CS_BIAS.n310 30.7807
R15394 CS_BIAS.n326 CS_BIAS.n308 30.7807
R15395 CS_BIAS.n280 CS_BIAS.n271 30.7807
R15396 CS_BIAS.n287 CS_BIAS.n269 30.7807
R15397 CS_BIAS.n206 CS_BIAS.n197 30.7807
R15398 CS_BIAS.n213 CS_BIAS.n195 30.7807
R15399 CS_BIAS.n249 CS_BIAS.n176 30.7807
R15400 CS_BIAS.n239 CS_BIAS.n232 30.7807
R15401 CS_BIAS.n142 CS_BIAS.t23 27.5579
R15402 CS_BIAS.n150 CS_BIAS.t32 27.5579
R15403 CS_BIAS.n135 CS_BIAS.t35 27.5579
R15404 CS_BIAS.n168 CS_BIAS.t47 27.5579
R15405 CS_BIAS.n129 CS_BIAS.t31 27.5579
R15406 CS_BIAS.n96 CS_BIAS.t44 27.5579
R15407 CS_BIAS.n111 CS_BIAS.t26 27.5579
R15408 CS_BIAS.n103 CS_BIAS.t39 27.5579
R15409 CS_BIAS.n42 CS_BIAS.t2 27.5579
R15410 CS_BIAS.n9 CS_BIAS.t12 27.5579
R15411 CS_BIAS.n24 CS_BIAS.t0 27.5579
R15412 CS_BIAS.n16 CS_BIAS.t4 27.5579
R15413 CS_BIAS.n91 CS_BIAS.t30 27.5579
R15414 CS_BIAS.n3 CS_BIAS.t49 27.5579
R15415 CS_BIAS.n73 CS_BIAS.t46 27.5579
R15416 CS_BIAS.n63 CS_BIAS.t38 27.5579
R15417 CS_BIAS.n313 CS_BIAS.t42 27.5579
R15418 CS_BIAS.n321 CS_BIAS.t25 27.5579
R15419 CS_BIAS.n306 CS_BIAS.t33 27.5579
R15420 CS_BIAS.n339 CS_BIAS.t34 27.5579
R15421 CS_BIAS.n274 CS_BIAS.t20 27.5579
R15422 CS_BIAS.n282 CS_BIAS.t37 27.5579
R15423 CS_BIAS.n267 CS_BIAS.t21 27.5579
R15424 CS_BIAS.n300 CS_BIAS.t43 27.5579
R15425 CS_BIAS.n200 CS_BIAS.t18 27.5579
R15426 CS_BIAS.n208 CS_BIAS.t10 27.5579
R15427 CS_BIAS.n193 CS_BIAS.t6 27.5579
R15428 CS_BIAS.n226 CS_BIAS.t16 27.5579
R15429 CS_BIAS.n262 CS_BIAS.t48 27.5579
R15430 CS_BIAS.n174 CS_BIAS.t45 27.5579
R15431 CS_BIAS.n234 CS_BIAS.t27 27.5579
R15432 CS_BIAS.n244 CS_BIAS.t36 27.5579
R15433 CS_BIAS.n144 CS_BIAS.n143 24.4675
R15434 CS_BIAS.n151 CS_BIAS.n137 24.4675
R15435 CS_BIAS.n149 CS_BIAS.n148 24.4675
R15436 CS_BIAS.n162 CS_BIAS.n161 24.4675
R15437 CS_BIAS.n161 CS_BIAS.n160 24.4675
R15438 CS_BIAS.n157 CS_BIAS.n156 24.4675
R15439 CS_BIAS.n167 CS_BIAS.n166 24.4675
R15440 CS_BIAS.n166 CS_BIAS.n133 24.4675
R15441 CS_BIAS.n128 CS_BIAS.n127 24.4675
R15442 CS_BIAS.n127 CS_BIAS.n94 24.4675
R15443 CS_BIAS.n123 CS_BIAS.n122 24.4675
R15444 CS_BIAS.n122 CS_BIAS.n121 24.4675
R15445 CS_BIAS.n118 CS_BIAS.n117 24.4675
R15446 CS_BIAS.n112 CS_BIAS.n98 24.4675
R15447 CS_BIAS.n110 CS_BIAS.n109 24.4675
R15448 CS_BIAS.n105 CS_BIAS.n104 24.4675
R15449 CS_BIAS.n41 CS_BIAS.n40 24.4675
R15450 CS_BIAS.n40 CS_BIAS.n7 24.4675
R15451 CS_BIAS.n36 CS_BIAS.n35 24.4675
R15452 CS_BIAS.n35 CS_BIAS.n34 24.4675
R15453 CS_BIAS.n31 CS_BIAS.n30 24.4675
R15454 CS_BIAS.n25 CS_BIAS.n11 24.4675
R15455 CS_BIAS.n23 CS_BIAS.n22 24.4675
R15456 CS_BIAS.n18 CS_BIAS.n17 24.4675
R15457 CS_BIAS.n90 CS_BIAS.n89 24.4675
R15458 CS_BIAS.n89 CS_BIAS.n1 24.4675
R15459 CS_BIAS.n85 CS_BIAS.n84 24.4675
R15460 CS_BIAS.n84 CS_BIAS.n83 24.4675
R15461 CS_BIAS.n80 CS_BIAS.n79 24.4675
R15462 CS_BIAS.n74 CS_BIAS.n5 24.4675
R15463 CS_BIAS.n72 CS_BIAS.n61 24.4675
R15464 CS_BIAS.n67 CS_BIAS.n66 24.4675
R15465 CS_BIAS.n315 CS_BIAS.n314 24.4675
R15466 CS_BIAS.n320 CS_BIAS.n319 24.4675
R15467 CS_BIAS.n322 CS_BIAS.n308 24.4675
R15468 CS_BIAS.n328 CS_BIAS.n327 24.4675
R15469 CS_BIAS.n332 CS_BIAS.n331 24.4675
R15470 CS_BIAS.n333 CS_BIAS.n332 24.4675
R15471 CS_BIAS.n337 CS_BIAS.n304 24.4675
R15472 CS_BIAS.n338 CS_BIAS.n337 24.4675
R15473 CS_BIAS.n276 CS_BIAS.n275 24.4675
R15474 CS_BIAS.n281 CS_BIAS.n280 24.4675
R15475 CS_BIAS.n283 CS_BIAS.n269 24.4675
R15476 CS_BIAS.n289 CS_BIAS.n288 24.4675
R15477 CS_BIAS.n293 CS_BIAS.n292 24.4675
R15478 CS_BIAS.n294 CS_BIAS.n293 24.4675
R15479 CS_BIAS.n298 CS_BIAS.n265 24.4675
R15480 CS_BIAS.n299 CS_BIAS.n298 24.4675
R15481 CS_BIAS.n202 CS_BIAS.n201 24.4675
R15482 CS_BIAS.n207 CS_BIAS.n206 24.4675
R15483 CS_BIAS.n209 CS_BIAS.n195 24.4675
R15484 CS_BIAS.n215 CS_BIAS.n214 24.4675
R15485 CS_BIAS.n219 CS_BIAS.n218 24.4675
R15486 CS_BIAS.n220 CS_BIAS.n219 24.4675
R15487 CS_BIAS.n224 CS_BIAS.n191 24.4675
R15488 CS_BIAS.n225 CS_BIAS.n224 24.4675
R15489 CS_BIAS.n260 CS_BIAS.n172 24.4675
R15490 CS_BIAS.n261 CS_BIAS.n260 24.4675
R15491 CS_BIAS.n251 CS_BIAS.n250 24.4675
R15492 CS_BIAS.n255 CS_BIAS.n254 24.4675
R15493 CS_BIAS.n256 CS_BIAS.n255 24.4675
R15494 CS_BIAS.n238 CS_BIAS.n237 24.4675
R15495 CS_BIAS.n243 CS_BIAS.n232 24.4675
R15496 CS_BIAS.n245 CS_BIAS.n176 24.4675
R15497 CS_BIAS.n143 CS_BIAS.n142 22.0208
R15498 CS_BIAS.n157 CS_BIAS.n135 22.0208
R15499 CS_BIAS.n118 CS_BIAS.n96 22.0208
R15500 CS_BIAS.n104 CS_BIAS.n103 22.0208
R15501 CS_BIAS.n31 CS_BIAS.n9 22.0208
R15502 CS_BIAS.n17 CS_BIAS.n16 22.0208
R15503 CS_BIAS.n80 CS_BIAS.n3 22.0208
R15504 CS_BIAS.n66 CS_BIAS.n63 22.0208
R15505 CS_BIAS.n314 CS_BIAS.n313 22.0208
R15506 CS_BIAS.n328 CS_BIAS.n306 22.0208
R15507 CS_BIAS.n275 CS_BIAS.n274 22.0208
R15508 CS_BIAS.n289 CS_BIAS.n267 22.0208
R15509 CS_BIAS.n201 CS_BIAS.n200 22.0208
R15510 CS_BIAS.n215 CS_BIAS.n193 22.0208
R15511 CS_BIAS.n251 CS_BIAS.n174 22.0208
R15512 CS_BIAS.n237 CS_BIAS.n234 22.0208
R15513 CS_BIAS.n342 CS_BIAS.n170 12.7372
R15514 CS_BIAS.n151 CS_BIAS.n150 12.234
R15515 CS_BIAS.n150 CS_BIAS.n149 12.234
R15516 CS_BIAS.n112 CS_BIAS.n111 12.234
R15517 CS_BIAS.n111 CS_BIAS.n110 12.234
R15518 CS_BIAS.n25 CS_BIAS.n24 12.234
R15519 CS_BIAS.n24 CS_BIAS.n23 12.234
R15520 CS_BIAS.n74 CS_BIAS.n73 12.234
R15521 CS_BIAS.n73 CS_BIAS.n72 12.234
R15522 CS_BIAS.n321 CS_BIAS.n320 12.234
R15523 CS_BIAS.n322 CS_BIAS.n321 12.234
R15524 CS_BIAS.n282 CS_BIAS.n281 12.234
R15525 CS_BIAS.n283 CS_BIAS.n282 12.234
R15526 CS_BIAS.n208 CS_BIAS.n207 12.234
R15527 CS_BIAS.n209 CS_BIAS.n208 12.234
R15528 CS_BIAS.n244 CS_BIAS.n243 12.234
R15529 CS_BIAS.n245 CS_BIAS.n244 12.234
R15530 CS_BIAS.n229 CS_BIAS.n227 11.8921
R15531 CS_BIAS.n55 CS_BIAS.n43 11.3102
R15532 CS_BIAS.n48 CS_BIAS.n47 10.1164
R15533 CS_BIAS.n181 CS_BIAS.n180 10.1164
R15534 CS_BIAS.n60 CS_BIAS.n59 9.50363
R15535 CS_BIAS.n231 CS_BIAS.n230 9.50363
R15536 CS_BIAS.n54 CS_BIAS.n53 9.45567
R15537 CS_BIAS.n187 CS_BIAS.n186 9.45567
R15538 CS_BIAS.n342 CS_BIAS.n341 9.32527
R15539 CS_BIAS.n53 CS_BIAS.n52 9.3005
R15540 CS_BIAS.n46 CS_BIAS.n45 9.3005
R15541 CS_BIAS.n186 CS_BIAS.n185 9.3005
R15542 CS_BIAS.n179 CS_BIAS.n178 9.3005
R15543 CS_BIAS.n54 CS_BIAS.n44 8.92171
R15544 CS_BIAS.n187 CS_BIAS.n177 8.92171
R15545 CS_BIAS.n52 CS_BIAS.n51 8.14595
R15546 CS_BIAS.n185 CS_BIAS.n184 8.14595
R15547 CS_BIAS.n48 CS_BIAS.n46 7.3702
R15548 CS_BIAS.n181 CS_BIAS.n179 7.3702
R15549 CS_BIAS.n168 CS_BIAS.n167 7.3406
R15550 CS_BIAS.n129 CS_BIAS.n128 7.3406
R15551 CS_BIAS.n42 CS_BIAS.n41 7.3406
R15552 CS_BIAS.n91 CS_BIAS.n90 7.3406
R15553 CS_BIAS.n339 CS_BIAS.n338 7.3406
R15554 CS_BIAS.n300 CS_BIAS.n299 7.3406
R15555 CS_BIAS.n226 CS_BIAS.n225 7.3406
R15556 CS_BIAS.n262 CS_BIAS.n261 7.3406
R15557 CS_BIAS.n58 CS_BIAS.t5 7.30677
R15558 CS_BIAS.n58 CS_BIAS.t15 7.30677
R15559 CS_BIAS.n56 CS_BIAS.t13 7.30677
R15560 CS_BIAS.n56 CS_BIAS.t1 7.30677
R15561 CS_BIAS.n228 CS_BIAS.t7 7.30677
R15562 CS_BIAS.n228 CS_BIAS.t17 7.30677
R15563 CS_BIAS.n188 CS_BIAS.t19 7.30677
R15564 CS_BIAS.n188 CS_BIAS.t11 7.30677
R15565 CS_BIAS.n131 CS_BIAS.n92 7.08717
R15566 CS_BIAS.n302 CS_BIAS.n263 7.08717
R15567 CS_BIAS.n141 CS_BIAS.n140 7.01727
R15568 CS_BIAS.n102 CS_BIAS.n101 7.01727
R15569 CS_BIAS.n15 CS_BIAS.n14 7.01727
R15570 CS_BIAS.n65 CS_BIAS.n64 7.01727
R15571 CS_BIAS.n312 CS_BIAS.n311 7.01727
R15572 CS_BIAS.n273 CS_BIAS.n272 7.01727
R15573 CS_BIAS.n199 CS_BIAS.n198 7.01727
R15574 CS_BIAS.n236 CS_BIAS.n235 7.01727
R15575 CS_BIAS.n51 CS_BIAS.n46 5.81868
R15576 CS_BIAS.n184 CS_BIAS.n179 5.81868
R15577 CS_BIAS.n52 CS_BIAS.n44 5.04292
R15578 CS_BIAS.n185 CS_BIAS.n177 5.04292
R15579 CS_BIAS.n170 CS_BIAS.n169 5.01898
R15580 CS_BIAS.n131 CS_BIAS.n130 5.01898
R15581 CS_BIAS.n341 CS_BIAS.n340 5.01898
R15582 CS_BIAS.n302 CS_BIAS.n301 5.01898
R15583 CS_BIAS CS_BIAS.n342 4.14131
R15584 CS_BIAS.n47 CS_BIAS.n45 3.00987
R15585 CS_BIAS.n180 CS_BIAS.n178 3.00987
R15586 CS_BIAS.n160 CS_BIAS.n135 2.4472
R15587 CS_BIAS.n121 CS_BIAS.n96 2.4472
R15588 CS_BIAS.n34 CS_BIAS.n9 2.4472
R15589 CS_BIAS.n83 CS_BIAS.n3 2.4472
R15590 CS_BIAS.n331 CS_BIAS.n306 2.4472
R15591 CS_BIAS.n292 CS_BIAS.n267 2.4472
R15592 CS_BIAS.n218 CS_BIAS.n193 2.4472
R15593 CS_BIAS.n254 CS_BIAS.n174 2.4472
R15594 CS_BIAS.n170 CS_BIAS.n131 2.06868
R15595 CS_BIAS.n341 CS_BIAS.n302 2.06868
R15596 CS_BIAS.n57 CS_BIAS.n55 1.16429
R15597 CS_BIAS.n230 CS_BIAS.n229 0.873345
R15598 CS_BIAS.n59 CS_BIAS.n57 0.291448
R15599 CS_BIAS.n230 CS_BIAS.n189 0.291448
R15600 CS_BIAS.n169 CS_BIAS.n132 0.278367
R15601 CS_BIAS.n130 CS_BIAS.n93 0.278367
R15602 CS_BIAS.n43 CS_BIAS.n6 0.278367
R15603 CS_BIAS.n92 CS_BIAS.n0 0.278367
R15604 CS_BIAS.n340 CS_BIAS.n303 0.278367
R15605 CS_BIAS.n301 CS_BIAS.n264 0.278367
R15606 CS_BIAS.n227 CS_BIAS.n190 0.278367
R15607 CS_BIAS.n263 CS_BIAS.n171 0.278367
R15608 CS_BIAS.n165 CS_BIAS.n132 0.189894
R15609 CS_BIAS.n165 CS_BIAS.n164 0.189894
R15610 CS_BIAS.n164 CS_BIAS.n163 0.189894
R15611 CS_BIAS.n163 CS_BIAS.n134 0.189894
R15612 CS_BIAS.n159 CS_BIAS.n134 0.189894
R15613 CS_BIAS.n159 CS_BIAS.n158 0.189894
R15614 CS_BIAS.n158 CS_BIAS.n136 0.189894
R15615 CS_BIAS.n154 CS_BIAS.n136 0.189894
R15616 CS_BIAS.n154 CS_BIAS.n153 0.189894
R15617 CS_BIAS.n153 CS_BIAS.n152 0.189894
R15618 CS_BIAS.n152 CS_BIAS.n138 0.189894
R15619 CS_BIAS.n147 CS_BIAS.n138 0.189894
R15620 CS_BIAS.n147 CS_BIAS.n146 0.189894
R15621 CS_BIAS.n146 CS_BIAS.n145 0.189894
R15622 CS_BIAS.n145 CS_BIAS.n140 0.189894
R15623 CS_BIAS.n126 CS_BIAS.n93 0.189894
R15624 CS_BIAS.n126 CS_BIAS.n125 0.189894
R15625 CS_BIAS.n125 CS_BIAS.n124 0.189894
R15626 CS_BIAS.n124 CS_BIAS.n95 0.189894
R15627 CS_BIAS.n120 CS_BIAS.n95 0.189894
R15628 CS_BIAS.n120 CS_BIAS.n119 0.189894
R15629 CS_BIAS.n119 CS_BIAS.n97 0.189894
R15630 CS_BIAS.n115 CS_BIAS.n97 0.189894
R15631 CS_BIAS.n115 CS_BIAS.n114 0.189894
R15632 CS_BIAS.n114 CS_BIAS.n113 0.189894
R15633 CS_BIAS.n113 CS_BIAS.n99 0.189894
R15634 CS_BIAS.n108 CS_BIAS.n99 0.189894
R15635 CS_BIAS.n108 CS_BIAS.n107 0.189894
R15636 CS_BIAS.n107 CS_BIAS.n106 0.189894
R15637 CS_BIAS.n106 CS_BIAS.n101 0.189894
R15638 CS_BIAS.n39 CS_BIAS.n6 0.189894
R15639 CS_BIAS.n39 CS_BIAS.n38 0.189894
R15640 CS_BIAS.n38 CS_BIAS.n37 0.189894
R15641 CS_BIAS.n37 CS_BIAS.n8 0.189894
R15642 CS_BIAS.n33 CS_BIAS.n8 0.189894
R15643 CS_BIAS.n33 CS_BIAS.n32 0.189894
R15644 CS_BIAS.n32 CS_BIAS.n10 0.189894
R15645 CS_BIAS.n28 CS_BIAS.n10 0.189894
R15646 CS_BIAS.n28 CS_BIAS.n27 0.189894
R15647 CS_BIAS.n27 CS_BIAS.n26 0.189894
R15648 CS_BIAS.n26 CS_BIAS.n12 0.189894
R15649 CS_BIAS.n21 CS_BIAS.n12 0.189894
R15650 CS_BIAS.n21 CS_BIAS.n20 0.189894
R15651 CS_BIAS.n20 CS_BIAS.n19 0.189894
R15652 CS_BIAS.n19 CS_BIAS.n14 0.189894
R15653 CS_BIAS.n71 CS_BIAS.n70 0.189894
R15654 CS_BIAS.n70 CS_BIAS.n69 0.189894
R15655 CS_BIAS.n69 CS_BIAS.n62 0.189894
R15656 CS_BIAS.n65 CS_BIAS.n62 0.189894
R15657 CS_BIAS.n88 CS_BIAS.n0 0.189894
R15658 CS_BIAS.n88 CS_BIAS.n87 0.189894
R15659 CS_BIAS.n87 CS_BIAS.n86 0.189894
R15660 CS_BIAS.n86 CS_BIAS.n2 0.189894
R15661 CS_BIAS.n82 CS_BIAS.n2 0.189894
R15662 CS_BIAS.n82 CS_BIAS.n81 0.189894
R15663 CS_BIAS.n81 CS_BIAS.n4 0.189894
R15664 CS_BIAS.n77 CS_BIAS.n4 0.189894
R15665 CS_BIAS.n77 CS_BIAS.n76 0.189894
R15666 CS_BIAS.n76 CS_BIAS.n75 0.189894
R15667 CS_BIAS.n316 CS_BIAS.n311 0.189894
R15668 CS_BIAS.n317 CS_BIAS.n316 0.189894
R15669 CS_BIAS.n318 CS_BIAS.n317 0.189894
R15670 CS_BIAS.n318 CS_BIAS.n309 0.189894
R15671 CS_BIAS.n323 CS_BIAS.n309 0.189894
R15672 CS_BIAS.n324 CS_BIAS.n323 0.189894
R15673 CS_BIAS.n325 CS_BIAS.n324 0.189894
R15674 CS_BIAS.n325 CS_BIAS.n307 0.189894
R15675 CS_BIAS.n329 CS_BIAS.n307 0.189894
R15676 CS_BIAS.n330 CS_BIAS.n329 0.189894
R15677 CS_BIAS.n330 CS_BIAS.n305 0.189894
R15678 CS_BIAS.n334 CS_BIAS.n305 0.189894
R15679 CS_BIAS.n335 CS_BIAS.n334 0.189894
R15680 CS_BIAS.n336 CS_BIAS.n335 0.189894
R15681 CS_BIAS.n336 CS_BIAS.n303 0.189894
R15682 CS_BIAS.n277 CS_BIAS.n272 0.189894
R15683 CS_BIAS.n278 CS_BIAS.n277 0.189894
R15684 CS_BIAS.n279 CS_BIAS.n278 0.189894
R15685 CS_BIAS.n279 CS_BIAS.n270 0.189894
R15686 CS_BIAS.n284 CS_BIAS.n270 0.189894
R15687 CS_BIAS.n285 CS_BIAS.n284 0.189894
R15688 CS_BIAS.n286 CS_BIAS.n285 0.189894
R15689 CS_BIAS.n286 CS_BIAS.n268 0.189894
R15690 CS_BIAS.n290 CS_BIAS.n268 0.189894
R15691 CS_BIAS.n291 CS_BIAS.n290 0.189894
R15692 CS_BIAS.n291 CS_BIAS.n266 0.189894
R15693 CS_BIAS.n295 CS_BIAS.n266 0.189894
R15694 CS_BIAS.n296 CS_BIAS.n295 0.189894
R15695 CS_BIAS.n297 CS_BIAS.n296 0.189894
R15696 CS_BIAS.n297 CS_BIAS.n264 0.189894
R15697 CS_BIAS.n203 CS_BIAS.n198 0.189894
R15698 CS_BIAS.n204 CS_BIAS.n203 0.189894
R15699 CS_BIAS.n205 CS_BIAS.n204 0.189894
R15700 CS_BIAS.n205 CS_BIAS.n196 0.189894
R15701 CS_BIAS.n210 CS_BIAS.n196 0.189894
R15702 CS_BIAS.n211 CS_BIAS.n210 0.189894
R15703 CS_BIAS.n212 CS_BIAS.n211 0.189894
R15704 CS_BIAS.n212 CS_BIAS.n194 0.189894
R15705 CS_BIAS.n216 CS_BIAS.n194 0.189894
R15706 CS_BIAS.n217 CS_BIAS.n216 0.189894
R15707 CS_BIAS.n217 CS_BIAS.n192 0.189894
R15708 CS_BIAS.n221 CS_BIAS.n192 0.189894
R15709 CS_BIAS.n222 CS_BIAS.n221 0.189894
R15710 CS_BIAS.n223 CS_BIAS.n222 0.189894
R15711 CS_BIAS.n223 CS_BIAS.n190 0.189894
R15712 CS_BIAS.n236 CS_BIAS.n233 0.189894
R15713 CS_BIAS.n240 CS_BIAS.n233 0.189894
R15714 CS_BIAS.n241 CS_BIAS.n240 0.189894
R15715 CS_BIAS.n242 CS_BIAS.n241 0.189894
R15716 CS_BIAS.n247 CS_BIAS.n246 0.189894
R15717 CS_BIAS.n248 CS_BIAS.n247 0.189894
R15718 CS_BIAS.n248 CS_BIAS.n175 0.189894
R15719 CS_BIAS.n252 CS_BIAS.n175 0.189894
R15720 CS_BIAS.n253 CS_BIAS.n252 0.189894
R15721 CS_BIAS.n253 CS_BIAS.n173 0.189894
R15722 CS_BIAS.n257 CS_BIAS.n173 0.189894
R15723 CS_BIAS.n258 CS_BIAS.n257 0.189894
R15724 CS_BIAS.n259 CS_BIAS.n258 0.189894
R15725 CS_BIAS.n259 CS_BIAS.n171 0.189894
R15726 CS_BIAS.n53 CS_BIAS.n45 0.155672
R15727 CS_BIAS.n186 CS_BIAS.n178 0.155672
R15728 CS_BIAS.n71 CS_BIAS.n60 0.0762576
R15729 CS_BIAS.n75 CS_BIAS.n60 0.0762576
R15730 CS_BIAS.n242 CS_BIAS.n231 0.0762576
R15731 CS_BIAS.n246 CS_BIAS.n231 0.0762576
R15732 VOUT.n212 VOUT.n198 756.745
R15733 VOUT.n192 VOUT.n178 756.745
R15734 VOUT.n172 VOUT.n158 756.745
R15735 VOUT.n152 VOUT.n138 756.745
R15736 VOUT.n133 VOUT.n119 756.745
R15737 VOUT.n93 VOUT.n79 756.745
R15738 VOUT.n73 VOUT.n59 756.745
R15739 VOUT.n53 VOUT.n39 756.745
R15740 VOUT.n33 VOUT.n19 756.745
R15741 VOUT.n14 VOUT.n0 756.745
R15742 VOUT.n213 VOUT.n212 585
R15743 VOUT.n211 VOUT.n210 585
R15744 VOUT.n202 VOUT.n201 585
R15745 VOUT.n205 VOUT.n204 585
R15746 VOUT.n193 VOUT.n192 585
R15747 VOUT.n191 VOUT.n190 585
R15748 VOUT.n182 VOUT.n181 585
R15749 VOUT.n185 VOUT.n184 585
R15750 VOUT.n173 VOUT.n172 585
R15751 VOUT.n171 VOUT.n170 585
R15752 VOUT.n162 VOUT.n161 585
R15753 VOUT.n165 VOUT.n164 585
R15754 VOUT.n153 VOUT.n152 585
R15755 VOUT.n151 VOUT.n150 585
R15756 VOUT.n142 VOUT.n141 585
R15757 VOUT.n145 VOUT.n144 585
R15758 VOUT.n134 VOUT.n133 585
R15759 VOUT.n132 VOUT.n131 585
R15760 VOUT.n123 VOUT.n122 585
R15761 VOUT.n126 VOUT.n125 585
R15762 VOUT.n94 VOUT.n93 585
R15763 VOUT.n92 VOUT.n91 585
R15764 VOUT.n83 VOUT.n82 585
R15765 VOUT.n86 VOUT.n85 585
R15766 VOUT.n74 VOUT.n73 585
R15767 VOUT.n72 VOUT.n71 585
R15768 VOUT.n63 VOUT.n62 585
R15769 VOUT.n66 VOUT.n65 585
R15770 VOUT.n54 VOUT.n53 585
R15771 VOUT.n52 VOUT.n51 585
R15772 VOUT.n43 VOUT.n42 585
R15773 VOUT.n46 VOUT.n45 585
R15774 VOUT.n34 VOUT.n33 585
R15775 VOUT.n32 VOUT.n31 585
R15776 VOUT.n23 VOUT.n22 585
R15777 VOUT.n26 VOUT.n25 585
R15778 VOUT.n15 VOUT.n14 585
R15779 VOUT.n13 VOUT.n12 585
R15780 VOUT.n4 VOUT.n3 585
R15781 VOUT.n7 VOUT.n6 585
R15782 VOUT.t31 VOUT.n203 330.707
R15783 VOUT.t30 VOUT.n183 330.707
R15784 VOUT.t32 VOUT.n163 330.707
R15785 VOUT.t38 VOUT.n143 330.707
R15786 VOUT.t34 VOUT.n124 330.707
R15787 VOUT.t33 VOUT.n84 330.707
R15788 VOUT.t39 VOUT.n64 330.707
R15789 VOUT.t36 VOUT.n44 330.707
R15790 VOUT.t35 VOUT.n24 330.707
R15791 VOUT.t37 VOUT.n5 330.707
R15792 VOUT.n256 VOUT.n250 289.615
R15793 VOUT.n240 VOUT.n234 289.615
R15794 VOUT.n225 VOUT.n219 289.615
R15795 VOUT.n307 VOUT.n301 289.615
R15796 VOUT.n291 VOUT.n285 289.615
R15797 VOUT.n276 VOUT.n270 289.615
R15798 VOUT.n257 VOUT.n256 185
R15799 VOUT.n255 VOUT.n254 185
R15800 VOUT.n241 VOUT.n240 185
R15801 VOUT.n239 VOUT.n238 185
R15802 VOUT.n226 VOUT.n225 185
R15803 VOUT.n224 VOUT.n223 185
R15804 VOUT.n308 VOUT.n307 185
R15805 VOUT.n306 VOUT.n305 185
R15806 VOUT.n292 VOUT.n291 185
R15807 VOUT.n290 VOUT.n289 185
R15808 VOUT.n277 VOUT.n276 185
R15809 VOUT.n275 VOUT.n274 185
R15810 VOUT.n212 VOUT.n211 171.744
R15811 VOUT.n211 VOUT.n201 171.744
R15812 VOUT.n204 VOUT.n201 171.744
R15813 VOUT.n192 VOUT.n191 171.744
R15814 VOUT.n191 VOUT.n181 171.744
R15815 VOUT.n184 VOUT.n181 171.744
R15816 VOUT.n172 VOUT.n171 171.744
R15817 VOUT.n171 VOUT.n161 171.744
R15818 VOUT.n164 VOUT.n161 171.744
R15819 VOUT.n152 VOUT.n151 171.744
R15820 VOUT.n151 VOUT.n141 171.744
R15821 VOUT.n144 VOUT.n141 171.744
R15822 VOUT.n133 VOUT.n132 171.744
R15823 VOUT.n132 VOUT.n122 171.744
R15824 VOUT.n125 VOUT.n122 171.744
R15825 VOUT.n93 VOUT.n92 171.744
R15826 VOUT.n92 VOUT.n82 171.744
R15827 VOUT.n85 VOUT.n82 171.744
R15828 VOUT.n73 VOUT.n72 171.744
R15829 VOUT.n72 VOUT.n62 171.744
R15830 VOUT.n65 VOUT.n62 171.744
R15831 VOUT.n53 VOUT.n52 171.744
R15832 VOUT.n52 VOUT.n42 171.744
R15833 VOUT.n45 VOUT.n42 171.744
R15834 VOUT.n33 VOUT.n32 171.744
R15835 VOUT.n32 VOUT.n22 171.744
R15836 VOUT.n25 VOUT.n22 171.744
R15837 VOUT.n14 VOUT.n13 171.744
R15838 VOUT.n13 VOUT.n3 171.744
R15839 VOUT.n6 VOUT.n3 171.744
R15840 VOUT.n253 VOUT.t2 153.582
R15841 VOUT.n237 VOUT.t18 153.582
R15842 VOUT.n222 VOUT.t19 153.582
R15843 VOUT.n304 VOUT.t9 153.582
R15844 VOUT.n288 VOUT.t20 153.582
R15845 VOUT.n273 VOUT.t25 153.582
R15846 VOUT.n256 VOUT.n255 104.615
R15847 VOUT.n240 VOUT.n239 104.615
R15848 VOUT.n225 VOUT.n224 104.615
R15849 VOUT.n307 VOUT.n306 104.615
R15850 VOUT.n291 VOUT.n290 104.615
R15851 VOUT.n276 VOUT.n275 104.615
R15852 VOUT.n300 VOUT.n298 103.484
R15853 VOUT.n284 VOUT.n282 103.484
R15854 VOUT.n269 VOUT.n267 103.484
R15855 VOUT.n264 VOUT.n263 102.322
R15856 VOUT.n262 VOUT.n261 102.322
R15857 VOUT.n248 VOUT.n247 102.322
R15858 VOUT.n246 VOUT.n245 102.322
R15859 VOUT.n233 VOUT.n232 102.322
R15860 VOUT.n231 VOUT.n230 102.322
R15861 VOUT.n300 VOUT.n299 102.322
R15862 VOUT.n284 VOUT.n283 102.322
R15863 VOUT.n269 VOUT.n268 102.322
R15864 VOUT.n204 VOUT.t31 85.8723
R15865 VOUT.n184 VOUT.t30 85.8723
R15866 VOUT.n164 VOUT.t32 85.8723
R15867 VOUT.n144 VOUT.t38 85.8723
R15868 VOUT.n125 VOUT.t34 85.8723
R15869 VOUT.n85 VOUT.t33 85.8723
R15870 VOUT.n65 VOUT.t39 85.8723
R15871 VOUT.n45 VOUT.t36 85.8723
R15872 VOUT.n25 VOUT.t35 85.8723
R15873 VOUT.n6 VOUT.t37 85.8723
R15874 VOUT.n157 VOUT.n137 75.8593
R15875 VOUT.n38 VOUT.n18 75.0856
R15876 VOUT.n217 VOUT.n216 74.3852
R15877 VOUT.n197 VOUT.n196 74.3852
R15878 VOUT.n177 VOUT.n176 74.3852
R15879 VOUT.n157 VOUT.n156 74.3852
R15880 VOUT.n98 VOUT.n97 73.6115
R15881 VOUT.n78 VOUT.n77 73.6115
R15882 VOUT.n58 VOUT.n57 73.6115
R15883 VOUT.n38 VOUT.n37 73.6115
R15884 VOUT.n262 VOUT.n260 65.931
R15885 VOUT.n246 VOUT.n244 65.931
R15886 VOUT.n231 VOUT.n229 65.931
R15887 VOUT.n312 VOUT.n311 64.7672
R15888 VOUT.n296 VOUT.n295 64.7672
R15889 VOUT.n281 VOUT.n280 64.7672
R15890 VOUT.n255 VOUT.t2 52.3082
R15891 VOUT.n239 VOUT.t18 52.3082
R15892 VOUT.n224 VOUT.t19 52.3082
R15893 VOUT.n306 VOUT.t9 52.3082
R15894 VOUT.n290 VOUT.t20 52.3082
R15895 VOUT.n275 VOUT.t25 52.3082
R15896 VOUT.n205 VOUT.n203 16.3201
R15897 VOUT.n185 VOUT.n183 16.3201
R15898 VOUT.n165 VOUT.n163 16.3201
R15899 VOUT.n145 VOUT.n143 16.3201
R15900 VOUT.n126 VOUT.n124 16.3201
R15901 VOUT.n86 VOUT.n84 16.3201
R15902 VOUT.n66 VOUT.n64 16.3201
R15903 VOUT.n46 VOUT.n44 16.3201
R15904 VOUT.n26 VOUT.n24 16.3201
R15905 VOUT.n7 VOUT.n5 16.3201
R15906 VOUT.n206 VOUT.n202 12.8005
R15907 VOUT.n186 VOUT.n182 12.8005
R15908 VOUT.n166 VOUT.n162 12.8005
R15909 VOUT.n146 VOUT.n142 12.8005
R15910 VOUT.n127 VOUT.n123 12.8005
R15911 VOUT.n87 VOUT.n83 12.8005
R15912 VOUT.n67 VOUT.n63 12.8005
R15913 VOUT.n47 VOUT.n43 12.8005
R15914 VOUT.n27 VOUT.n23 12.8005
R15915 VOUT.n8 VOUT.n4 12.8005
R15916 VOUT.n210 VOUT.n209 12.0247
R15917 VOUT.n190 VOUT.n189 12.0247
R15918 VOUT.n170 VOUT.n169 12.0247
R15919 VOUT.n150 VOUT.n149 12.0247
R15920 VOUT.n131 VOUT.n130 12.0247
R15921 VOUT.n91 VOUT.n90 12.0247
R15922 VOUT.n71 VOUT.n70 12.0247
R15923 VOUT.n51 VOUT.n50 12.0247
R15924 VOUT.n31 VOUT.n30 12.0247
R15925 VOUT.n12 VOUT.n11 12.0247
R15926 VOUT.n213 VOUT.n200 11.249
R15927 VOUT.n193 VOUT.n180 11.249
R15928 VOUT.n173 VOUT.n160 11.249
R15929 VOUT.n153 VOUT.n140 11.249
R15930 VOUT.n134 VOUT.n121 11.249
R15931 VOUT.n94 VOUT.n81 11.249
R15932 VOUT.n74 VOUT.n61 11.249
R15933 VOUT.n54 VOUT.n41 11.249
R15934 VOUT.n34 VOUT.n21 11.249
R15935 VOUT.n15 VOUT.n2 11.249
R15936 VOUT.n214 VOUT.n198 10.4732
R15937 VOUT.n194 VOUT.n178 10.4732
R15938 VOUT.n174 VOUT.n158 10.4732
R15939 VOUT.n154 VOUT.n138 10.4732
R15940 VOUT.n135 VOUT.n119 10.4732
R15941 VOUT.n95 VOUT.n79 10.4732
R15942 VOUT.n75 VOUT.n59 10.4732
R15943 VOUT.n55 VOUT.n39 10.4732
R15944 VOUT.n35 VOUT.n19 10.4732
R15945 VOUT.n16 VOUT.n0 10.4732
R15946 VOUT.n254 VOUT.n253 10.1164
R15947 VOUT.n238 VOUT.n237 10.1164
R15948 VOUT.n223 VOUT.n222 10.1164
R15949 VOUT.n305 VOUT.n304 10.1164
R15950 VOUT.n289 VOUT.n288 10.1164
R15951 VOUT.n274 VOUT.n273 10.1164
R15952 VOUT.n216 VOUT.n215 9.45567
R15953 VOUT.n196 VOUT.n195 9.45567
R15954 VOUT.n176 VOUT.n175 9.45567
R15955 VOUT.n156 VOUT.n155 9.45567
R15956 VOUT.n137 VOUT.n136 9.45567
R15957 VOUT.n97 VOUT.n96 9.45567
R15958 VOUT.n77 VOUT.n76 9.45567
R15959 VOUT.n57 VOUT.n56 9.45567
R15960 VOUT.n37 VOUT.n36 9.45567
R15961 VOUT.n18 VOUT.n17 9.45567
R15962 VOUT.n260 VOUT.n259 9.45567
R15963 VOUT.n244 VOUT.n243 9.45567
R15964 VOUT.n229 VOUT.n228 9.45567
R15965 VOUT.n311 VOUT.n310 9.45567
R15966 VOUT.n295 VOUT.n294 9.45567
R15967 VOUT.n280 VOUT.n279 9.45567
R15968 VOUT.n215 VOUT.n214 9.3005
R15969 VOUT.n200 VOUT.n199 9.3005
R15970 VOUT.n209 VOUT.n208 9.3005
R15971 VOUT.n207 VOUT.n206 9.3005
R15972 VOUT.n195 VOUT.n194 9.3005
R15973 VOUT.n180 VOUT.n179 9.3005
R15974 VOUT.n189 VOUT.n188 9.3005
R15975 VOUT.n187 VOUT.n186 9.3005
R15976 VOUT.n175 VOUT.n174 9.3005
R15977 VOUT.n160 VOUT.n159 9.3005
R15978 VOUT.n169 VOUT.n168 9.3005
R15979 VOUT.n167 VOUT.n166 9.3005
R15980 VOUT.n155 VOUT.n154 9.3005
R15981 VOUT.n140 VOUT.n139 9.3005
R15982 VOUT.n149 VOUT.n148 9.3005
R15983 VOUT.n147 VOUT.n146 9.3005
R15984 VOUT.n136 VOUT.n135 9.3005
R15985 VOUT.n121 VOUT.n120 9.3005
R15986 VOUT.n130 VOUT.n129 9.3005
R15987 VOUT.n128 VOUT.n127 9.3005
R15988 VOUT.n96 VOUT.n95 9.3005
R15989 VOUT.n81 VOUT.n80 9.3005
R15990 VOUT.n90 VOUT.n89 9.3005
R15991 VOUT.n88 VOUT.n87 9.3005
R15992 VOUT.n76 VOUT.n75 9.3005
R15993 VOUT.n61 VOUT.n60 9.3005
R15994 VOUT.n70 VOUT.n69 9.3005
R15995 VOUT.n68 VOUT.n67 9.3005
R15996 VOUT.n56 VOUT.n55 9.3005
R15997 VOUT.n41 VOUT.n40 9.3005
R15998 VOUT.n50 VOUT.n49 9.3005
R15999 VOUT.n48 VOUT.n47 9.3005
R16000 VOUT.n36 VOUT.n35 9.3005
R16001 VOUT.n21 VOUT.n20 9.3005
R16002 VOUT.n30 VOUT.n29 9.3005
R16003 VOUT.n28 VOUT.n27 9.3005
R16004 VOUT.n17 VOUT.n16 9.3005
R16005 VOUT.n2 VOUT.n1 9.3005
R16006 VOUT.n11 VOUT.n10 9.3005
R16007 VOUT.n9 VOUT.n8 9.3005
R16008 VOUT.n259 VOUT.n258 9.3005
R16009 VOUT.n252 VOUT.n251 9.3005
R16010 VOUT.n243 VOUT.n242 9.3005
R16011 VOUT.n236 VOUT.n235 9.3005
R16012 VOUT.n228 VOUT.n227 9.3005
R16013 VOUT.n221 VOUT.n220 9.3005
R16014 VOUT.n310 VOUT.n309 9.3005
R16015 VOUT.n303 VOUT.n302 9.3005
R16016 VOUT.n294 VOUT.n293 9.3005
R16017 VOUT.n287 VOUT.n286 9.3005
R16018 VOUT.n279 VOUT.n278 9.3005
R16019 VOUT.n272 VOUT.n271 9.3005
R16020 VOUT.n260 VOUT.n250 8.92171
R16021 VOUT.n244 VOUT.n234 8.92171
R16022 VOUT.n229 VOUT.n219 8.92171
R16023 VOUT.n311 VOUT.n301 8.92171
R16024 VOUT.n295 VOUT.n285 8.92171
R16025 VOUT.n280 VOUT.n270 8.92171
R16026 VOUT.n266 VOUT.n218 8.86899
R16027 VOUT.n258 VOUT.n257 8.14595
R16028 VOUT.n242 VOUT.n241 8.14595
R16029 VOUT.n227 VOUT.n226 8.14595
R16030 VOUT.n309 VOUT.n308 8.14595
R16031 VOUT.n293 VOUT.n292 8.14595
R16032 VOUT.n278 VOUT.n277 8.14595
R16033 VOUT.n254 VOUT.n252 7.3702
R16034 VOUT.n238 VOUT.n236 7.3702
R16035 VOUT.n223 VOUT.n221 7.3702
R16036 VOUT.n305 VOUT.n303 7.3702
R16037 VOUT.n289 VOUT.n287 7.3702
R16038 VOUT.n274 VOUT.n272 7.3702
R16039 VOUT.n263 VOUT.t26 7.30677
R16040 VOUT.n263 VOUT.t8 7.30677
R16041 VOUT.n261 VOUT.t14 7.30677
R16042 VOUT.n261 VOUT.t17 7.30677
R16043 VOUT.n247 VOUT.t10 7.30677
R16044 VOUT.n247 VOUT.t27 7.30677
R16045 VOUT.n245 VOUT.t5 7.30677
R16046 VOUT.n245 VOUT.t23 7.30677
R16047 VOUT.n232 VOUT.t11 7.30677
R16048 VOUT.n232 VOUT.t21 7.30677
R16049 VOUT.n230 VOUT.t0 7.30677
R16050 VOUT.n230 VOUT.t3 7.30677
R16051 VOUT.n298 VOUT.t16 7.30677
R16052 VOUT.n298 VOUT.t15 7.30677
R16053 VOUT.n299 VOUT.t7 7.30677
R16054 VOUT.n299 VOUT.t24 7.30677
R16055 VOUT.n282 VOUT.t28 7.30677
R16056 VOUT.n282 VOUT.t6 7.30677
R16057 VOUT.n283 VOUT.t29 7.30677
R16058 VOUT.n283 VOUT.t12 7.30677
R16059 VOUT.n267 VOUT.t4 7.30677
R16060 VOUT.n267 VOUT.t1 7.30677
R16061 VOUT.n268 VOUT.t22 7.30677
R16062 VOUT.n268 VOUT.t13 7.30677
R16063 VOUT.n249 VOUT.n233 6.74619
R16064 VOUT.n266 VOUT.n265 6.348
R16065 VOUT.n314 VOUT.n313 6.348
R16066 VOUT.n297 VOUT.n281 6.16429
R16067 VOUT.n257 VOUT.n252 5.81868
R16068 VOUT.n241 VOUT.n236 5.81868
R16069 VOUT.n226 VOUT.n221 5.81868
R16070 VOUT.n308 VOUT.n303 5.81868
R16071 VOUT.n292 VOUT.n287 5.81868
R16072 VOUT.n277 VOUT.n272 5.81868
R16073 VOUT.n265 VOUT.n264 5.54791
R16074 VOUT.n249 VOUT.n248 5.54791
R16075 VOUT.n258 VOUT.n250 5.04292
R16076 VOUT.n242 VOUT.n234 5.04292
R16077 VOUT.n227 VOUT.n219 5.04292
R16078 VOUT.n309 VOUT.n301 5.04292
R16079 VOUT.n293 VOUT.n285 5.04292
R16080 VOUT.n278 VOUT.n270 5.04292
R16081 VOUT.n218 VOUT.n99 5.02041
R16082 VOUT.n313 VOUT.n312 4.96602
R16083 VOUT.n297 VOUT.n296 4.96602
R16084 VOUT.n315 VOUT.n99 4.87831
R16085 VOUT.n218 VOUT.n217 4.78873
R16086 VOUT.n99 VOUT.n98 4.78873
R16087 VOUT.n314 VOUT.n266 4.36899
R16088 VOUT.n315 VOUT.n314 3.97168
R16089 VOUT.n207 VOUT.n203 3.78097
R16090 VOUT.n187 VOUT.n183 3.78097
R16091 VOUT.n167 VOUT.n163 3.78097
R16092 VOUT.n147 VOUT.n143 3.78097
R16093 VOUT.n128 VOUT.n124 3.78097
R16094 VOUT.n88 VOUT.n84 3.78097
R16095 VOUT.n68 VOUT.n64 3.78097
R16096 VOUT.n48 VOUT.n44 3.78097
R16097 VOUT.n28 VOUT.n24 3.78097
R16098 VOUT.n9 VOUT.n5 3.78097
R16099 VOUT.n216 VOUT.n198 3.49141
R16100 VOUT.n196 VOUT.n178 3.49141
R16101 VOUT.n176 VOUT.n158 3.49141
R16102 VOUT.n156 VOUT.n138 3.49141
R16103 VOUT.n137 VOUT.n119 3.49141
R16104 VOUT.n97 VOUT.n79 3.49141
R16105 VOUT.n77 VOUT.n59 3.49141
R16106 VOUT.n57 VOUT.n39 3.49141
R16107 VOUT.n37 VOUT.n19 3.49141
R16108 VOUT.n18 VOUT.n0 3.49141
R16109 VOUT.n253 VOUT.n251 3.00987
R16110 VOUT.n237 VOUT.n235 3.00987
R16111 VOUT.n222 VOUT.n220 3.00987
R16112 VOUT.n304 VOUT.n302 3.00987
R16113 VOUT.n288 VOUT.n286 3.00987
R16114 VOUT.n273 VOUT.n271 3.00987
R16115 VOUT.n118 VOUT 2.9239
R16116 VOUT.n214 VOUT.n213 2.71565
R16117 VOUT.n194 VOUT.n193 2.71565
R16118 VOUT.n174 VOUT.n173 2.71565
R16119 VOUT.n154 VOUT.n153 2.71565
R16120 VOUT.n135 VOUT.n134 2.71565
R16121 VOUT.n95 VOUT.n94 2.71565
R16122 VOUT.n75 VOUT.n74 2.71565
R16123 VOUT.n55 VOUT.n54 2.71565
R16124 VOUT.n35 VOUT.n34 2.71565
R16125 VOUT.n16 VOUT.n15 2.71565
R16126 VOUT.n210 VOUT.n200 1.93989
R16127 VOUT.n190 VOUT.n180 1.93989
R16128 VOUT.n170 VOUT.n160 1.93989
R16129 VOUT.n150 VOUT.n140 1.93989
R16130 VOUT.n131 VOUT.n121 1.93989
R16131 VOUT.n91 VOUT.n81 1.93989
R16132 VOUT.n71 VOUT.n61 1.93989
R16133 VOUT.n51 VOUT.n41 1.93989
R16134 VOUT.n31 VOUT.n21 1.93989
R16135 VOUT.n12 VOUT.n2 1.93989
R16136 VOUT.n217 VOUT.n197 1.47464
R16137 VOUT.n197 VOUT.n177 1.47464
R16138 VOUT.n177 VOUT.n157 1.47464
R16139 VOUT.n98 VOUT.n78 1.47464
R16140 VOUT.n78 VOUT.n58 1.47464
R16141 VOUT.n58 VOUT.n38 1.47464
R16142 VOUT.n265 VOUT.n249 1.19878
R16143 VOUT.n313 VOUT.n297 1.19878
R16144 VOUT.n264 VOUT.n262 1.16429
R16145 VOUT.n248 VOUT.n246 1.16429
R16146 VOUT.n233 VOUT.n231 1.16429
R16147 VOUT.n312 VOUT.n300 1.16429
R16148 VOUT.n296 VOUT.n284 1.16429
R16149 VOUT.n281 VOUT.n269 1.16429
R16150 VOUT.n209 VOUT.n202 1.16414
R16151 VOUT.n189 VOUT.n182 1.16414
R16152 VOUT.n169 VOUT.n162 1.16414
R16153 VOUT.n149 VOUT.n142 1.16414
R16154 VOUT.n130 VOUT.n123 1.16414
R16155 VOUT.n90 VOUT.n83 1.16414
R16156 VOUT.n70 VOUT.n63 1.16414
R16157 VOUT.n50 VOUT.n43 1.16414
R16158 VOUT.n30 VOUT.n23 1.16414
R16159 VOUT.n11 VOUT.n4 1.16414
R16160 VOUT.n206 VOUT.n205 0.388379
R16161 VOUT.n186 VOUT.n185 0.388379
R16162 VOUT.n166 VOUT.n165 0.388379
R16163 VOUT.n146 VOUT.n145 0.388379
R16164 VOUT.n127 VOUT.n126 0.388379
R16165 VOUT.n87 VOUT.n86 0.388379
R16166 VOUT.n67 VOUT.n66 0.388379
R16167 VOUT.n47 VOUT.n46 0.388379
R16168 VOUT.n27 VOUT.n26 0.388379
R16169 VOUT.n8 VOUT.n7 0.388379
R16170 VOUT.n118 VOUT.n117 0.349024
R16171 VOUT.n315 VOUT.n118 0.28344
R16172 VOUT.n215 VOUT.n199 0.155672
R16173 VOUT.n208 VOUT.n199 0.155672
R16174 VOUT.n208 VOUT.n207 0.155672
R16175 VOUT.n195 VOUT.n179 0.155672
R16176 VOUT.n188 VOUT.n179 0.155672
R16177 VOUT.n188 VOUT.n187 0.155672
R16178 VOUT.n175 VOUT.n159 0.155672
R16179 VOUT.n168 VOUT.n159 0.155672
R16180 VOUT.n168 VOUT.n167 0.155672
R16181 VOUT.n155 VOUT.n139 0.155672
R16182 VOUT.n148 VOUT.n139 0.155672
R16183 VOUT.n148 VOUT.n147 0.155672
R16184 VOUT.n136 VOUT.n120 0.155672
R16185 VOUT.n129 VOUT.n120 0.155672
R16186 VOUT.n129 VOUT.n128 0.155672
R16187 VOUT.n96 VOUT.n80 0.155672
R16188 VOUT.n89 VOUT.n80 0.155672
R16189 VOUT.n89 VOUT.n88 0.155672
R16190 VOUT.n76 VOUT.n60 0.155672
R16191 VOUT.n69 VOUT.n60 0.155672
R16192 VOUT.n69 VOUT.n68 0.155672
R16193 VOUT.n56 VOUT.n40 0.155672
R16194 VOUT.n49 VOUT.n40 0.155672
R16195 VOUT.n49 VOUT.n48 0.155672
R16196 VOUT.n36 VOUT.n20 0.155672
R16197 VOUT.n29 VOUT.n20 0.155672
R16198 VOUT.n29 VOUT.n28 0.155672
R16199 VOUT.n17 VOUT.n1 0.155672
R16200 VOUT.n10 VOUT.n1 0.155672
R16201 VOUT.n10 VOUT.n9 0.155672
R16202 VOUT.n259 VOUT.n251 0.155672
R16203 VOUT.n243 VOUT.n235 0.155672
R16204 VOUT.n228 VOUT.n220 0.155672
R16205 VOUT.n310 VOUT.n302 0.155672
R16206 VOUT.n294 VOUT.n286 0.155672
R16207 VOUT.n279 VOUT.n271 0.155672
R16208 VOUT.n104 VOUT.t46 0.144808
R16209 VOUT.n107 VOUT.t43 0.144808
R16210 VOUT.n113 VOUT.t45 0.144808
R16211 VOUT.n115 VOUT.t40 0.144808
R16212 VOUT.n117 VOUT.t41 0.144808
R16213 VOUT.n106 VOUT.t46 0.144753
R16214 VOUT.n109 VOUT.t43 0.144753
R16215 VOUT.t45 VOUT.n112 0.144753
R16216 VOUT.t40 VOUT.n114 0.144753
R16217 VOUT.t41 VOUT.n116 0.144753
R16218 VOUT.n104 VOUT.n103 0.107924
R16219 VOUT.n110 VOUT.n109 0.107284
R16220 VOUT.n112 VOUT.n111 0.107284
R16221 VOUT.n107 VOUT.n106 0.0978715
R16222 VOUT.n114 VOUT.n113 0.0978715
R16223 VOUT.n116 VOUT.n115 0.0978715
R16224 VOUT.n110 VOUT.t42 0.073695
R16225 VOUT.n111 VOUT.t44 0.073695
R16226 VOUT.n103 VOUT.t47 0.0732793
R16227 VOUT.n111 VOUT.n110 0.066909
R16228 VOUT.n103 VOUT.n100 0.0507055
R16229 VOUT.n108 VOUT.n102 0.0391444
R16230 VOUT.n105 VOUT.n101 0.0391444
R16231 VOUT.n105 VOUT.n104 0.0242263
R16232 VOUT.n108 VOUT.n107 0.0242263
R16233 VOUT.n113 VOUT.n102 0.0242263
R16234 VOUT.n115 VOUT.n101 0.0242263
R16235 VOUT.n117 VOUT.n100 0.0242263
R16236 VOUT.n106 VOUT.n105 0.0225754
R16237 VOUT.n109 VOUT.n108 0.0225754
R16238 VOUT.n112 VOUT.n102 0.0225754
R16239 VOUT.n114 VOUT.n101 0.0225754
R16240 VOUT.n116 VOUT.n100 0.0225754
R16241 VOUT VOUT.n315 0.0099
R16242 VDD.n3397 VDD.n3383 756.745
R16243 VDD.n3377 VDD.n3363 756.745
R16244 VDD.n3357 VDD.n3343 756.745
R16245 VDD.n3337 VDD.n3323 756.745
R16246 VDD.n3318 VDD.n3304 756.745
R16247 VDD.n1433 VDD.n1419 756.745
R16248 VDD.n1413 VDD.n1399 756.745
R16249 VDD.n1393 VDD.n1379 756.745
R16250 VDD.n1373 VDD.n1359 756.745
R16251 VDD.n1354 VDD.n1340 756.745
R16252 VDD.n3398 VDD.n3397 585
R16253 VDD.n3396 VDD.n3395 585
R16254 VDD.n3387 VDD.n3386 585
R16255 VDD.n3390 VDD.n3389 585
R16256 VDD.n3378 VDD.n3377 585
R16257 VDD.n3376 VDD.n3375 585
R16258 VDD.n3367 VDD.n3366 585
R16259 VDD.n3370 VDD.n3369 585
R16260 VDD.n3358 VDD.n3357 585
R16261 VDD.n3356 VDD.n3355 585
R16262 VDD.n3347 VDD.n3346 585
R16263 VDD.n3350 VDD.n3349 585
R16264 VDD.n3338 VDD.n3337 585
R16265 VDD.n3336 VDD.n3335 585
R16266 VDD.n3327 VDD.n3326 585
R16267 VDD.n3330 VDD.n3329 585
R16268 VDD.n3319 VDD.n3318 585
R16269 VDD.n3317 VDD.n3316 585
R16270 VDD.n3308 VDD.n3307 585
R16271 VDD.n3311 VDD.n3310 585
R16272 VDD.n1434 VDD.n1433 585
R16273 VDD.n1432 VDD.n1431 585
R16274 VDD.n1423 VDD.n1422 585
R16275 VDD.n1426 VDD.n1425 585
R16276 VDD.n1414 VDD.n1413 585
R16277 VDD.n1412 VDD.n1411 585
R16278 VDD.n1403 VDD.n1402 585
R16279 VDD.n1406 VDD.n1405 585
R16280 VDD.n1394 VDD.n1393 585
R16281 VDD.n1392 VDD.n1391 585
R16282 VDD.n1383 VDD.n1382 585
R16283 VDD.n1386 VDD.n1385 585
R16284 VDD.n1374 VDD.n1373 585
R16285 VDD.n1372 VDD.n1371 585
R16286 VDD.n1363 VDD.n1362 585
R16287 VDD.n1366 VDD.n1365 585
R16288 VDD.n1355 VDD.n1354 585
R16289 VDD.n1353 VDD.n1352 585
R16290 VDD.n1344 VDD.n1343 585
R16291 VDD.n1347 VDD.n1346 585
R16292 VDD.n2907 VDD.n59 446.341
R16293 VDD.n3077 VDD.n2995 446.341
R16294 VDD.n3269 VDD.n2997 446.341
R16295 VDD.n2910 VDD.n61 446.341
R16296 VDD.n1555 VDD.n962 446.341
R16297 VDD.n1558 VDD.n1557 446.341
R16298 VDD.n1287 VDD.n1039 446.341
R16299 VDD.n1289 VDD.n1037 446.341
R16300 VDD.t137 VDD.n3388 330.707
R16301 VDD.t134 VDD.n3368 330.707
R16302 VDD.t138 VDD.n3348 330.707
R16303 VDD.t127 VDD.n3328 330.707
R16304 VDD.t132 VDD.n3309 330.707
R16305 VDD.t104 VDD.n1424 330.707
R16306 VDD.t99 VDD.n1404 330.707
R16307 VDD.t103 VDD.n1384 330.707
R16308 VDD.t133 VDD.n1364 330.707
R16309 VDD.t141 VDD.n1345 330.707
R16310 VDD.n2727 VDD.n166 313.171
R16311 VDD.n2701 VDD.n180 313.171
R16312 VDD.n2401 VDD.n2400 313.171
R16313 VDD.n2429 VDD.n417 313.171
R16314 VDD.n2116 VDD.n440 313.171
R16315 VDD.n2087 VDD.n2086 313.171
R16316 VDD.n1770 VDD.n1769 313.171
R16317 VDD.n1798 VDD.n697 313.171
R16318 VDD.n2679 VDD.n2678 313.171
R16319 VDD.n2737 VDD.n158 313.171
R16320 VDD.n2278 VDD.n2131 313.171
R16321 VDD.n2433 VDD.n421 313.171
R16322 VDD.n2072 VDD.n2071 313.171
R16323 VDD.n2041 VDD.n432 313.171
R16324 VDD.n900 VDD.n713 313.171
R16325 VDD.n769 VDD.n693 313.171
R16326 VDD.n1042 VDD.t26 305.06
R16327 VDD.n1058 VDD.t5 305.06
R16328 VDD.n1076 VDD.t56 305.06
R16329 VDD.n1093 VDD.t53 305.06
R16330 VDD.n1110 VDD.t59 305.06
R16331 VDD.n1510 VDD.t83 305.06
R16332 VDD.n956 VDD.t77 305.06
R16333 VDD.n925 VDD.t49 305.06
R16334 VDD.n753 VDD.t80 305.06
R16335 VDD.n729 VDD.t74 305.06
R16336 VDD.n3032 VDD.t92 305.06
R16337 VDD.n3042 VDD.t86 305.06
R16338 VDD.n3050 VDD.t32 305.06
R16339 VDD.n3059 VDD.t29 305.06
R16340 VDD.n3069 VDD.t35 305.06
R16341 VDD.n114 VDD.t19 305.06
R16342 VDD.n140 VDD.t16 305.06
R16343 VDD.n2856 VDD.t9 305.06
R16344 VDD.n64 VDD.t69 305.06
R16345 VDD.n2756 VDD.t42 305.06
R16346 VDD.n784 VDD.t66 295.156
R16347 VDD.n460 VDD.t22 295.156
R16348 VDD.n1647 VDD.t13 295.156
R16349 VDD.n443 VDD.t38 295.156
R16350 VDD.n2132 VDD.t90 295.156
R16351 VDD.n176 VDD.t45 295.156
R16352 VDD.n2281 VDD.t63 295.156
R16353 VDD.n154 VDD.t71 295.156
R16354 VDD.n1042 VDD.t24 238.362
R16355 VDD.n1058 VDD.t2 238.362
R16356 VDD.n1076 VDD.t54 238.362
R16357 VDD.n1093 VDD.t51 238.362
R16358 VDD.n1110 VDD.t57 238.362
R16359 VDD.n1510 VDD.t82 238.362
R16360 VDD.n956 VDD.t76 238.362
R16361 VDD.n925 VDD.t47 238.362
R16362 VDD.n753 VDD.t79 238.362
R16363 VDD.n729 VDD.t73 238.362
R16364 VDD.n3032 VDD.t91 238.362
R16365 VDD.n3042 VDD.t85 238.362
R16366 VDD.n3050 VDD.t31 238.362
R16367 VDD.n3059 VDD.t27 238.362
R16368 VDD.n3069 VDD.t34 238.362
R16369 VDD.n114 VDD.t17 238.362
R16370 VDD.n140 VDD.t14 238.362
R16371 VDD.n2856 VDD.t6 238.362
R16372 VDD.n64 VDD.t67 238.362
R16373 VDD.n2756 VDD.t40 238.362
R16374 VDD.n1043 VDD.t25 235.435
R16375 VDD.n1059 VDD.t4 235.435
R16376 VDD.n1077 VDD.t55 235.435
R16377 VDD.n1094 VDD.t52 235.435
R16378 VDD.n1111 VDD.t58 235.435
R16379 VDD.n1511 VDD.t84 235.435
R16380 VDD.n957 VDD.t78 235.435
R16381 VDD.n926 VDD.t50 235.435
R16382 VDD.n754 VDD.t81 235.435
R16383 VDD.n730 VDD.t75 235.435
R16384 VDD.n3033 VDD.t93 235.435
R16385 VDD.n3043 VDD.t87 235.435
R16386 VDD.n3051 VDD.t33 235.435
R16387 VDD.n3060 VDD.t30 235.435
R16388 VDD.n3070 VDD.t36 235.435
R16389 VDD.n115 VDD.t18 235.435
R16390 VDD.n141 VDD.t15 235.435
R16391 VDD.n2857 VDD.t8 235.435
R16392 VDD.n65 VDD.t68 235.435
R16393 VDD.n2757 VDD.t41 235.435
R16394 VDD.n784 VDD.t64 210.653
R16395 VDD.n460 VDD.t20 210.653
R16396 VDD.n1647 VDD.t10 210.653
R16397 VDD.n443 VDD.t37 210.653
R16398 VDD.n2132 VDD.t88 210.653
R16399 VDD.n176 VDD.t43 210.653
R16400 VDD.n2281 VDD.t60 210.653
R16401 VDD.n154 VDD.t70 210.653
R16402 VDD.n9 VDD.n7 194.87
R16403 VDD.n2 VDD.n0 194.87
R16404 VDD.n9 VDD.n8 192.173
R16405 VDD.n11 VDD.n10 192.173
R16406 VDD.n13 VDD.n12 192.173
R16407 VDD.n6 VDD.n5 192.173
R16408 VDD.n4 VDD.n3 192.173
R16409 VDD.n2 VDD.n1 192.173
R16410 VDD.t0 VDD.t94 191.406
R16411 VDD.t135 VDD.t1 191.406
R16412 VDD.n721 VDD.t0 191.147
R16413 VDD.n2909 VDD.t1 191.147
R16414 VDD.n2680 VDD.n2679 185
R16415 VDD.n2679 VDD.n163 185
R16416 VDD.n2681 VDD.n164 185
R16417 VDD.n2732 VDD.n164 185
R16418 VDD.n2683 VDD.n2682 185
R16419 VDD.n2682 VDD.n161 185
R16420 VDD.n2684 VDD.n185 185
R16421 VDD.n2694 VDD.n185 185
R16422 VDD.n2685 VDD.n193 185
R16423 VDD.n193 VDD.n183 185
R16424 VDD.n2687 VDD.n2686 185
R16425 VDD.n2688 VDD.n2687 185
R16426 VDD.n2663 VDD.n192 185
R16427 VDD.n192 VDD.n189 185
R16428 VDD.n2662 VDD.n2661 185
R16429 VDD.n2661 VDD.n2660 185
R16430 VDD.n195 VDD.n194 185
R16431 VDD.n196 VDD.n195 185
R16432 VDD.n2653 VDD.n2652 185
R16433 VDD.n2654 VDD.n2653 185
R16434 VDD.n2651 VDD.n205 185
R16435 VDD.n205 VDD.n202 185
R16436 VDD.n2650 VDD.n2649 185
R16437 VDD.n2649 VDD.n2648 185
R16438 VDD.n207 VDD.n206 185
R16439 VDD.n208 VDD.n207 185
R16440 VDD.n2641 VDD.n2640 185
R16441 VDD.n2642 VDD.n2641 185
R16442 VDD.n2639 VDD.n217 185
R16443 VDD.n217 VDD.n214 185
R16444 VDD.n2638 VDD.n2637 185
R16445 VDD.n2637 VDD.n2636 185
R16446 VDD.n219 VDD.n218 185
R16447 VDD.n220 VDD.n219 185
R16448 VDD.n2629 VDD.n2628 185
R16449 VDD.n2630 VDD.n2629 185
R16450 VDD.n2627 VDD.n229 185
R16451 VDD.n229 VDD.n226 185
R16452 VDD.n2626 VDD.n2625 185
R16453 VDD.n2625 VDD.n2624 185
R16454 VDD.n231 VDD.n230 185
R16455 VDD.n232 VDD.n231 185
R16456 VDD.n2617 VDD.n2616 185
R16457 VDD.n2618 VDD.n2617 185
R16458 VDD.n2615 VDD.n241 185
R16459 VDD.n241 VDD.n238 185
R16460 VDD.n2614 VDD.n2613 185
R16461 VDD.n2613 VDD.n2612 185
R16462 VDD.n243 VDD.n242 185
R16463 VDD.n244 VDD.n243 185
R16464 VDD.n2605 VDD.n2604 185
R16465 VDD.n2606 VDD.n2605 185
R16466 VDD.n2603 VDD.n253 185
R16467 VDD.n253 VDD.n250 185
R16468 VDD.n2602 VDD.n2601 185
R16469 VDD.n2601 VDD.n2600 185
R16470 VDD.n255 VDD.n254 185
R16471 VDD.n256 VDD.n255 185
R16472 VDD.n2593 VDD.n2592 185
R16473 VDD.n2594 VDD.n2593 185
R16474 VDD.n2591 VDD.n265 185
R16475 VDD.n265 VDD.n262 185
R16476 VDD.n2590 VDD.n2589 185
R16477 VDD.n2589 VDD.n2588 185
R16478 VDD.n267 VDD.n266 185
R16479 VDD.n275 VDD.n267 185
R16480 VDD.n2581 VDD.n2580 185
R16481 VDD.n2582 VDD.n2581 185
R16482 VDD.n2579 VDD.n276 185
R16483 VDD.n282 VDD.n276 185
R16484 VDD.n2578 VDD.n2577 185
R16485 VDD.n2577 VDD.n2576 185
R16486 VDD.n278 VDD.n277 185
R16487 VDD.n279 VDD.n278 185
R16488 VDD.n2569 VDD.n2568 185
R16489 VDD.n2570 VDD.n2569 185
R16490 VDD.n2567 VDD.n289 185
R16491 VDD.n289 VDD.n286 185
R16492 VDD.n2566 VDD.n2565 185
R16493 VDD.n2565 VDD.n2564 185
R16494 VDD.n291 VDD.n290 185
R16495 VDD.n292 VDD.n291 185
R16496 VDD.n2557 VDD.n2556 185
R16497 VDD.n2558 VDD.n2557 185
R16498 VDD.n2555 VDD.n301 185
R16499 VDD.n301 VDD.n298 185
R16500 VDD.n2554 VDD.n2553 185
R16501 VDD.n2553 VDD.n2552 185
R16502 VDD.n303 VDD.n302 185
R16503 VDD.n304 VDD.n303 185
R16504 VDD.n2545 VDD.n2544 185
R16505 VDD.n2546 VDD.n2545 185
R16506 VDD.n2543 VDD.n313 185
R16507 VDD.n313 VDD.n310 185
R16508 VDD.n2542 VDD.n2541 185
R16509 VDD.n2541 VDD.n2540 185
R16510 VDD.n315 VDD.n314 185
R16511 VDD.n316 VDD.n315 185
R16512 VDD.n2533 VDD.n2532 185
R16513 VDD.n2534 VDD.n2533 185
R16514 VDD.n2531 VDD.n325 185
R16515 VDD.n325 VDD.n322 185
R16516 VDD.n2530 VDD.n2529 185
R16517 VDD.n2529 VDD.n2528 185
R16518 VDD.n327 VDD.n326 185
R16519 VDD.n336 VDD.n327 185
R16520 VDD.n2521 VDD.n2520 185
R16521 VDD.n2522 VDD.n2521 185
R16522 VDD.n2519 VDD.n337 185
R16523 VDD.n337 VDD.n333 185
R16524 VDD.n2518 VDD.n2517 185
R16525 VDD.n2517 VDD.n2516 185
R16526 VDD.n339 VDD.n338 185
R16527 VDD.n340 VDD.n339 185
R16528 VDD.n2509 VDD.n2508 185
R16529 VDD.n2510 VDD.n2509 185
R16530 VDD.n2507 VDD.n349 185
R16531 VDD.n349 VDD.n346 185
R16532 VDD.n2506 VDD.n2505 185
R16533 VDD.n2505 VDD.n2504 185
R16534 VDD.n351 VDD.n350 185
R16535 VDD.n352 VDD.n351 185
R16536 VDD.n2497 VDD.n2496 185
R16537 VDD.n2498 VDD.n2497 185
R16538 VDD.n2495 VDD.n361 185
R16539 VDD.n361 VDD.n358 185
R16540 VDD.n2494 VDD.n2493 185
R16541 VDD.n2493 VDD.n2492 185
R16542 VDD.n363 VDD.n362 185
R16543 VDD.n364 VDD.n363 185
R16544 VDD.n2485 VDD.n2484 185
R16545 VDD.n2486 VDD.n2485 185
R16546 VDD.n2483 VDD.n373 185
R16547 VDD.n373 VDD.n370 185
R16548 VDD.n2482 VDD.n2481 185
R16549 VDD.n2481 VDD.n2480 185
R16550 VDD.n375 VDD.n374 185
R16551 VDD.n376 VDD.n375 185
R16552 VDD.n2473 VDD.n2472 185
R16553 VDD.n2474 VDD.n2473 185
R16554 VDD.n2471 VDD.n384 185
R16555 VDD.n389 VDD.n384 185
R16556 VDD.n2470 VDD.n2469 185
R16557 VDD.n2469 VDD.n2468 185
R16558 VDD.n386 VDD.n385 185
R16559 VDD.n396 VDD.n386 185
R16560 VDD.n2461 VDD.n2460 185
R16561 VDD.n2462 VDD.n2461 185
R16562 VDD.n2459 VDD.n397 185
R16563 VDD.n397 VDD.n393 185
R16564 VDD.n2458 VDD.n2457 185
R16565 VDD.n2457 VDD.n2456 185
R16566 VDD.n399 VDD.n398 185
R16567 VDD.n400 VDD.n399 185
R16568 VDD.n2449 VDD.n2448 185
R16569 VDD.n2450 VDD.n2449 185
R16570 VDD.n2447 VDD.n409 185
R16571 VDD.n409 VDD.n406 185
R16572 VDD.n2446 VDD.n2445 185
R16573 VDD.n2445 VDD.n2444 185
R16574 VDD.n411 VDD.n410 185
R16575 VDD.n412 VDD.n411 185
R16576 VDD.n2437 VDD.n2436 185
R16577 VDD.n2438 VDD.n2437 185
R16578 VDD.n2435 VDD.n421 185
R16579 VDD.n421 VDD.n418 185
R16580 VDD.n2434 VDD.n2433 185
R16581 VDD.n423 VDD.n422 185
R16582 VDD.n2136 VDD.n2135 185
R16583 VDD.n2138 VDD.n2137 185
R16584 VDD.n2140 VDD.n2139 185
R16585 VDD.n2142 VDD.n2141 185
R16586 VDD.n2144 VDD.n2143 185
R16587 VDD.n2146 VDD.n2145 185
R16588 VDD.n2148 VDD.n2147 185
R16589 VDD.n2150 VDD.n2149 185
R16590 VDD.n2152 VDD.n2151 185
R16591 VDD.n2154 VDD.n2153 185
R16592 VDD.n2156 VDD.n2155 185
R16593 VDD.n2157 VDD.n2130 185
R16594 VDD.n2278 VDD.n2277 185
R16595 VDD.n2431 VDD.n2278 185
R16596 VDD.n2737 VDD.n2736 185
R16597 VDD.n2739 VDD.n156 185
R16598 VDD.n2741 VDD.n2740 185
R16599 VDD.n2743 VDD.n153 185
R16600 VDD.n2745 VDD.n2744 185
R16601 VDD.n2747 VDD.n152 185
R16602 VDD.n2748 VDD.n149 185
R16603 VDD.n2751 VDD.n2750 185
R16604 VDD.n150 VDD.n148 185
R16605 VDD.n2670 VDD.n2667 185
R16606 VDD.n2672 VDD.n2671 185
R16607 VDD.n2673 VDD.n2666 185
R16608 VDD.n2675 VDD.n2674 185
R16609 VDD.n2677 VDD.n2665 185
R16610 VDD.n2678 VDD.n2664 185
R16611 VDD.n2678 VDD.n151 185
R16612 VDD.n2735 VDD.n158 185
R16613 VDD.n163 VDD.n158 185
R16614 VDD.n2734 VDD.n2733 185
R16615 VDD.n2733 VDD.n2732 185
R16616 VDD.n160 VDD.n159 185
R16617 VDD.n161 VDD.n160 185
R16618 VDD.n2158 VDD.n184 185
R16619 VDD.n2694 VDD.n184 185
R16620 VDD.n2160 VDD.n2159 185
R16621 VDD.n2159 VDD.n183 185
R16622 VDD.n2161 VDD.n191 185
R16623 VDD.n2688 VDD.n191 185
R16624 VDD.n2163 VDD.n2162 185
R16625 VDD.n2162 VDD.n189 185
R16626 VDD.n2164 VDD.n198 185
R16627 VDD.n2660 VDD.n198 185
R16628 VDD.n2166 VDD.n2165 185
R16629 VDD.n2165 VDD.n196 185
R16630 VDD.n2167 VDD.n204 185
R16631 VDD.n2654 VDD.n204 185
R16632 VDD.n2169 VDD.n2168 185
R16633 VDD.n2168 VDD.n202 185
R16634 VDD.n2170 VDD.n210 185
R16635 VDD.n2648 VDD.n210 185
R16636 VDD.n2172 VDD.n2171 185
R16637 VDD.n2171 VDD.n208 185
R16638 VDD.n2173 VDD.n216 185
R16639 VDD.n2642 VDD.n216 185
R16640 VDD.n2175 VDD.n2174 185
R16641 VDD.n2174 VDD.n214 185
R16642 VDD.n2176 VDD.n222 185
R16643 VDD.n2636 VDD.n222 185
R16644 VDD.n2178 VDD.n2177 185
R16645 VDD.n2177 VDD.n220 185
R16646 VDD.n2179 VDD.n228 185
R16647 VDD.n2630 VDD.n228 185
R16648 VDD.n2181 VDD.n2180 185
R16649 VDD.n2180 VDD.n226 185
R16650 VDD.n2182 VDD.n234 185
R16651 VDD.n2624 VDD.n234 185
R16652 VDD.n2184 VDD.n2183 185
R16653 VDD.n2183 VDD.n232 185
R16654 VDD.n2185 VDD.n240 185
R16655 VDD.n2618 VDD.n240 185
R16656 VDD.n2187 VDD.n2186 185
R16657 VDD.n2186 VDD.n238 185
R16658 VDD.n2188 VDD.n246 185
R16659 VDD.n2612 VDD.n246 185
R16660 VDD.n2190 VDD.n2189 185
R16661 VDD.n2189 VDD.n244 185
R16662 VDD.n2191 VDD.n252 185
R16663 VDD.n2606 VDD.n252 185
R16664 VDD.n2193 VDD.n2192 185
R16665 VDD.n2192 VDD.n250 185
R16666 VDD.n2194 VDD.n258 185
R16667 VDD.n2600 VDD.n258 185
R16668 VDD.n2196 VDD.n2195 185
R16669 VDD.n2195 VDD.n256 185
R16670 VDD.n2197 VDD.n264 185
R16671 VDD.n2594 VDD.n264 185
R16672 VDD.n2199 VDD.n2198 185
R16673 VDD.n2198 VDD.n262 185
R16674 VDD.n2200 VDD.n269 185
R16675 VDD.n2588 VDD.n269 185
R16676 VDD.n2202 VDD.n2201 185
R16677 VDD.n2201 VDD.n275 185
R16678 VDD.n2203 VDD.n274 185
R16679 VDD.n2582 VDD.n274 185
R16680 VDD.n2205 VDD.n2204 185
R16681 VDD.n2204 VDD.n282 185
R16682 VDD.n2206 VDD.n281 185
R16683 VDD.n2576 VDD.n281 185
R16684 VDD.n2208 VDD.n2207 185
R16685 VDD.n2207 VDD.n279 185
R16686 VDD.n2209 VDD.n288 185
R16687 VDD.n2570 VDD.n288 185
R16688 VDD.n2211 VDD.n2210 185
R16689 VDD.n2210 VDD.n286 185
R16690 VDD.n2212 VDD.n294 185
R16691 VDD.n2564 VDD.n294 185
R16692 VDD.n2214 VDD.n2213 185
R16693 VDD.n2213 VDD.n292 185
R16694 VDD.n2215 VDD.n300 185
R16695 VDD.n2558 VDD.n300 185
R16696 VDD.n2217 VDD.n2216 185
R16697 VDD.n2216 VDD.n298 185
R16698 VDD.n2218 VDD.n306 185
R16699 VDD.n2552 VDD.n306 185
R16700 VDD.n2220 VDD.n2219 185
R16701 VDD.n2219 VDD.n304 185
R16702 VDD.n2221 VDD.n312 185
R16703 VDD.n2546 VDD.n312 185
R16704 VDD.n2223 VDD.n2222 185
R16705 VDD.n2222 VDD.n310 185
R16706 VDD.n2224 VDD.n318 185
R16707 VDD.n2540 VDD.n318 185
R16708 VDD.n2226 VDD.n2225 185
R16709 VDD.n2225 VDD.n316 185
R16710 VDD.n2227 VDD.n324 185
R16711 VDD.n2534 VDD.n324 185
R16712 VDD.n2229 VDD.n2228 185
R16713 VDD.n2228 VDD.n322 185
R16714 VDD.n2230 VDD.n329 185
R16715 VDD.n2528 VDD.n329 185
R16716 VDD.n2232 VDD.n2231 185
R16717 VDD.n2231 VDD.n336 185
R16718 VDD.n2233 VDD.n335 185
R16719 VDD.n2522 VDD.n335 185
R16720 VDD.n2235 VDD.n2234 185
R16721 VDD.n2234 VDD.n333 185
R16722 VDD.n2236 VDD.n342 185
R16723 VDD.n2516 VDD.n342 185
R16724 VDD.n2238 VDD.n2237 185
R16725 VDD.n2237 VDD.n340 185
R16726 VDD.n2239 VDD.n348 185
R16727 VDD.n2510 VDD.n348 185
R16728 VDD.n2241 VDD.n2240 185
R16729 VDD.n2240 VDD.n346 185
R16730 VDD.n2242 VDD.n354 185
R16731 VDD.n2504 VDD.n354 185
R16732 VDD.n2244 VDD.n2243 185
R16733 VDD.n2243 VDD.n352 185
R16734 VDD.n2245 VDD.n360 185
R16735 VDD.n2498 VDD.n360 185
R16736 VDD.n2247 VDD.n2246 185
R16737 VDD.n2246 VDD.n358 185
R16738 VDD.n2248 VDD.n366 185
R16739 VDD.n2492 VDD.n366 185
R16740 VDD.n2250 VDD.n2249 185
R16741 VDD.n2249 VDD.n364 185
R16742 VDD.n2251 VDD.n372 185
R16743 VDD.n2486 VDD.n372 185
R16744 VDD.n2253 VDD.n2252 185
R16745 VDD.n2252 VDD.n370 185
R16746 VDD.n2254 VDD.n378 185
R16747 VDD.n2480 VDD.n378 185
R16748 VDD.n2256 VDD.n2255 185
R16749 VDD.n2255 VDD.n376 185
R16750 VDD.n2257 VDD.n383 185
R16751 VDD.n2474 VDD.n383 185
R16752 VDD.n2259 VDD.n2258 185
R16753 VDD.n2258 VDD.n389 185
R16754 VDD.n2260 VDD.n388 185
R16755 VDD.n2468 VDD.n388 185
R16756 VDD.n2262 VDD.n2261 185
R16757 VDD.n2261 VDD.n396 185
R16758 VDD.n2263 VDD.n395 185
R16759 VDD.n2462 VDD.n395 185
R16760 VDD.n2265 VDD.n2264 185
R16761 VDD.n2264 VDD.n393 185
R16762 VDD.n2266 VDD.n402 185
R16763 VDD.n2456 VDD.n402 185
R16764 VDD.n2268 VDD.n2267 185
R16765 VDD.n2267 VDD.n400 185
R16766 VDD.n2269 VDD.n408 185
R16767 VDD.n2450 VDD.n408 185
R16768 VDD.n2271 VDD.n2270 185
R16769 VDD.n2270 VDD.n406 185
R16770 VDD.n2272 VDD.n414 185
R16771 VDD.n2444 VDD.n414 185
R16772 VDD.n2274 VDD.n2273 185
R16773 VDD.n2273 VDD.n412 185
R16774 VDD.n2275 VDD.n420 185
R16775 VDD.n2438 VDD.n420 185
R16776 VDD.n2276 VDD.n2131 185
R16777 VDD.n2131 VDD.n418 185
R16778 VDD.n442 VDD.n440 185
R16779 VDD.n440 VDD.n424 185
R16780 VDD.n2083 VDD.n2082 185
R16781 VDD.n2084 VDD.n2083 185
R16782 VDD.n2081 VDD.n451 185
R16783 VDD.n451 VDD.n448 185
R16784 VDD.n2080 VDD.n2079 185
R16785 VDD.n2079 VDD.n2078 185
R16786 VDD.n453 VDD.n452 185
R16787 VDD.n454 VDD.n453 185
R16788 VDD.n2032 VDD.n2031 185
R16789 VDD.n2033 VDD.n2032 185
R16790 VDD.n2030 VDD.n468 185
R16791 VDD.n468 VDD.n465 185
R16792 VDD.n2029 VDD.n2028 185
R16793 VDD.n2028 VDD.n2027 185
R16794 VDD.n470 VDD.n469 185
R16795 VDD.n471 VDD.n470 185
R16796 VDD.n2018 VDD.n2017 185
R16797 VDD.n2019 VDD.n2018 185
R16798 VDD.n2016 VDD.n481 185
R16799 VDD.n481 VDD.n478 185
R16800 VDD.n2015 VDD.n2014 185
R16801 VDD.n2014 VDD.n2013 185
R16802 VDD.n483 VDD.n482 185
R16803 VDD.n484 VDD.n483 185
R16804 VDD.n2006 VDD.n2005 185
R16805 VDD.n2007 VDD.n2006 185
R16806 VDD.n2004 VDD.n493 185
R16807 VDD.n493 VDD.n490 185
R16808 VDD.n2003 VDD.n2002 185
R16809 VDD.n2002 VDD.n2001 185
R16810 VDD.n495 VDD.n494 185
R16811 VDD.n496 VDD.n495 185
R16812 VDD.n1994 VDD.n1993 185
R16813 VDD.n1995 VDD.n1994 185
R16814 VDD.n1992 VDD.n505 185
R16815 VDD.n505 VDD.n502 185
R16816 VDD.n1991 VDD.n1990 185
R16817 VDD.n1990 VDD.n1989 185
R16818 VDD.n507 VDD.n506 185
R16819 VDD.n508 VDD.n507 185
R16820 VDD.n1982 VDD.n1981 185
R16821 VDD.n1983 VDD.n1982 185
R16822 VDD.n1980 VDD.n517 185
R16823 VDD.n517 VDD.n514 185
R16824 VDD.n1979 VDD.n1978 185
R16825 VDD.n1978 VDD.n1977 185
R16826 VDD.n519 VDD.n518 185
R16827 VDD.n520 VDD.n519 185
R16828 VDD.n1970 VDD.n1969 185
R16829 VDD.n1971 VDD.n1970 185
R16830 VDD.n1968 VDD.n529 185
R16831 VDD.n529 VDD.n526 185
R16832 VDD.n1967 VDD.n1966 185
R16833 VDD.n1966 VDD.n1965 185
R16834 VDD.n531 VDD.n530 185
R16835 VDD.n532 VDD.n531 185
R16836 VDD.n1958 VDD.n1957 185
R16837 VDD.n1959 VDD.n1958 185
R16838 VDD.n1956 VDD.n541 185
R16839 VDD.n541 VDD.n538 185
R16840 VDD.n1955 VDD.n1954 185
R16841 VDD.n1954 VDD.n1953 185
R16842 VDD.n543 VDD.n542 185
R16843 VDD.n552 VDD.n543 185
R16844 VDD.n1946 VDD.n1945 185
R16845 VDD.n1947 VDD.n1946 185
R16846 VDD.n1944 VDD.n553 185
R16847 VDD.n553 VDD.n549 185
R16848 VDD.n1943 VDD.n1942 185
R16849 VDD.n1942 VDD.n1941 185
R16850 VDD.n555 VDD.n554 185
R16851 VDD.n556 VDD.n555 185
R16852 VDD.n1934 VDD.n1933 185
R16853 VDD.n1935 VDD.n1934 185
R16854 VDD.n1932 VDD.n565 185
R16855 VDD.n565 VDD.n562 185
R16856 VDD.n1931 VDD.n1930 185
R16857 VDD.n1930 VDD.n1929 185
R16858 VDD.n567 VDD.n566 185
R16859 VDD.n568 VDD.n567 185
R16860 VDD.n1922 VDD.n1921 185
R16861 VDD.n1923 VDD.n1922 185
R16862 VDD.n1920 VDD.n577 185
R16863 VDD.n577 VDD.n574 185
R16864 VDD.n1919 VDD.n1918 185
R16865 VDD.n1918 VDD.n1917 185
R16866 VDD.n579 VDD.n578 185
R16867 VDD.n580 VDD.n579 185
R16868 VDD.n1910 VDD.n1909 185
R16869 VDD.n1911 VDD.n1910 185
R16870 VDD.n1908 VDD.n589 185
R16871 VDD.n589 VDD.n586 185
R16872 VDD.n1907 VDD.n1906 185
R16873 VDD.n1906 VDD.n1905 185
R16874 VDD.n591 VDD.n590 185
R16875 VDD.n592 VDD.n591 185
R16876 VDD.n1898 VDD.n1897 185
R16877 VDD.n1899 VDD.n1898 185
R16878 VDD.n1896 VDD.n601 185
R16879 VDD.n601 VDD.n598 185
R16880 VDD.n1895 VDD.n1894 185
R16881 VDD.n1894 VDD.n1893 185
R16882 VDD.n603 VDD.n602 185
R16883 VDD.n604 VDD.n603 185
R16884 VDD.n1886 VDD.n1885 185
R16885 VDD.n1887 VDD.n1886 185
R16886 VDD.n1884 VDD.n613 185
R16887 VDD.n613 VDD.n610 185
R16888 VDD.n1883 VDD.n1882 185
R16889 VDD.n1882 VDD.n1881 185
R16890 VDD.n615 VDD.n614 185
R16891 VDD.n616 VDD.n615 185
R16892 VDD.n1874 VDD.n1873 185
R16893 VDD.n1875 VDD.n1874 185
R16894 VDD.n1872 VDD.n625 185
R16895 VDD.n625 VDD.n622 185
R16896 VDD.n1871 VDD.n1870 185
R16897 VDD.n1870 VDD.n1869 185
R16898 VDD.n627 VDD.n626 185
R16899 VDD.n628 VDD.n627 185
R16900 VDD.n1862 VDD.n1861 185
R16901 VDD.n1863 VDD.n1862 185
R16902 VDD.n1860 VDD.n637 185
R16903 VDD.n637 VDD.n634 185
R16904 VDD.n1859 VDD.n1858 185
R16905 VDD.n1858 VDD.n1857 185
R16906 VDD.n639 VDD.n638 185
R16907 VDD.n640 VDD.n639 185
R16908 VDD.n1850 VDD.n1849 185
R16909 VDD.n1851 VDD.n1850 185
R16910 VDD.n1848 VDD.n649 185
R16911 VDD.n649 VDD.n646 185
R16912 VDD.n1847 VDD.n1846 185
R16913 VDD.n1846 VDD.n1845 185
R16914 VDD.n651 VDD.n650 185
R16915 VDD.n660 VDD.n651 185
R16916 VDD.n1838 VDD.n1837 185
R16917 VDD.n1839 VDD.n1838 185
R16918 VDD.n1836 VDD.n661 185
R16919 VDD.n661 VDD.n657 185
R16920 VDD.n1835 VDD.n1834 185
R16921 VDD.n1834 VDD.n1833 185
R16922 VDD.n663 VDD.n662 185
R16923 VDD.n672 VDD.n663 185
R16924 VDD.n1826 VDD.n1825 185
R16925 VDD.n1827 VDD.n1826 185
R16926 VDD.n1824 VDD.n673 185
R16927 VDD.n673 VDD.n669 185
R16928 VDD.n1823 VDD.n1822 185
R16929 VDD.n1822 VDD.n1821 185
R16930 VDD.n675 VDD.n674 185
R16931 VDD.n676 VDD.n675 185
R16932 VDD.n1814 VDD.n1813 185
R16933 VDD.n1815 VDD.n1814 185
R16934 VDD.n1812 VDD.n685 185
R16935 VDD.n685 VDD.n682 185
R16936 VDD.n1811 VDD.n1810 185
R16937 VDD.n1810 VDD.n1809 185
R16938 VDD.n687 VDD.n686 185
R16939 VDD.n688 VDD.n687 185
R16940 VDD.n1802 VDD.n1801 185
R16941 VDD.n1803 VDD.n1802 185
R16942 VDD.n1800 VDD.n697 185
R16943 VDD.n697 VDD.n694 185
R16944 VDD.n1799 VDD.n1798 185
R16945 VDD.n699 VDD.n698 185
R16946 VDD.n1795 VDD.n1794 185
R16947 VDD.n1796 VDD.n1795 185
R16948 VDD.n1793 VDD.n714 185
R16949 VDD.n1792 VDD.n1791 185
R16950 VDD.n1790 VDD.n1789 185
R16951 VDD.n1788 VDD.n1787 185
R16952 VDD.n1786 VDD.n1785 185
R16953 VDD.n1784 VDD.n1783 185
R16954 VDD.n1782 VDD.n1781 185
R16955 VDD.n1780 VDD.n1779 185
R16956 VDD.n1778 VDD.n1777 185
R16957 VDD.n1775 VDD.n1774 185
R16958 VDD.n1773 VDD.n1772 185
R16959 VDD.n1771 VDD.n1770 185
R16960 VDD.n2088 VDD.n2087 185
R16961 VDD.n2090 VDD.n2089 185
R16962 VDD.n2092 VDD.n2091 185
R16963 VDD.n2095 VDD.n2094 185
R16964 VDD.n2097 VDD.n2096 185
R16965 VDD.n2099 VDD.n2098 185
R16966 VDD.n2101 VDD.n2100 185
R16967 VDD.n2103 VDD.n2102 185
R16968 VDD.n2105 VDD.n2104 185
R16969 VDD.n2107 VDD.n2106 185
R16970 VDD.n2109 VDD.n2108 185
R16971 VDD.n2111 VDD.n2110 185
R16972 VDD.n2113 VDD.n2112 185
R16973 VDD.n2114 VDD.n441 185
R16974 VDD.n2116 VDD.n2115 185
R16975 VDD.n2117 VDD.n2116 185
R16976 VDD.n2086 VDD.n445 185
R16977 VDD.n2086 VDD.n424 185
R16978 VDD.n2085 VDD.n447 185
R16979 VDD.n2085 VDD.n2084 185
R16980 VDD.n1649 VDD.n446 185
R16981 VDD.n448 VDD.n446 185
R16982 VDD.n1650 VDD.n455 185
R16983 VDD.n2078 VDD.n455 185
R16984 VDD.n1652 VDD.n1651 185
R16985 VDD.n1651 VDD.n454 185
R16986 VDD.n1653 VDD.n466 185
R16987 VDD.n2033 VDD.n466 185
R16988 VDD.n1655 VDD.n1654 185
R16989 VDD.n1654 VDD.n465 185
R16990 VDD.n1656 VDD.n472 185
R16991 VDD.n2027 VDD.n472 185
R16992 VDD.n1658 VDD.n1657 185
R16993 VDD.n1657 VDD.n471 185
R16994 VDD.n1659 VDD.n479 185
R16995 VDD.n2019 VDD.n479 185
R16996 VDD.n1661 VDD.n1660 185
R16997 VDD.n1660 VDD.n478 185
R16998 VDD.n1662 VDD.n485 185
R16999 VDD.n2013 VDD.n485 185
R17000 VDD.n1664 VDD.n1663 185
R17001 VDD.n1663 VDD.n484 185
R17002 VDD.n1665 VDD.n491 185
R17003 VDD.n2007 VDD.n491 185
R17004 VDD.n1667 VDD.n1666 185
R17005 VDD.n1666 VDD.n490 185
R17006 VDD.n1668 VDD.n497 185
R17007 VDD.n2001 VDD.n497 185
R17008 VDD.n1670 VDD.n1669 185
R17009 VDD.n1669 VDD.n496 185
R17010 VDD.n1671 VDD.n503 185
R17011 VDD.n1995 VDD.n503 185
R17012 VDD.n1673 VDD.n1672 185
R17013 VDD.n1672 VDD.n502 185
R17014 VDD.n1674 VDD.n509 185
R17015 VDD.n1989 VDD.n509 185
R17016 VDD.n1676 VDD.n1675 185
R17017 VDD.n1675 VDD.n508 185
R17018 VDD.n1677 VDD.n515 185
R17019 VDD.n1983 VDD.n515 185
R17020 VDD.n1679 VDD.n1678 185
R17021 VDD.n1678 VDD.n514 185
R17022 VDD.n1680 VDD.n521 185
R17023 VDD.n1977 VDD.n521 185
R17024 VDD.n1682 VDD.n1681 185
R17025 VDD.n1681 VDD.n520 185
R17026 VDD.n1683 VDD.n527 185
R17027 VDD.n1971 VDD.n527 185
R17028 VDD.n1685 VDD.n1684 185
R17029 VDD.n1684 VDD.n526 185
R17030 VDD.n1686 VDD.n533 185
R17031 VDD.n1965 VDD.n533 185
R17032 VDD.n1688 VDD.n1687 185
R17033 VDD.n1687 VDD.n532 185
R17034 VDD.n1689 VDD.n539 185
R17035 VDD.n1959 VDD.n539 185
R17036 VDD.n1691 VDD.n1690 185
R17037 VDD.n1690 VDD.n538 185
R17038 VDD.n1692 VDD.n544 185
R17039 VDD.n1953 VDD.n544 185
R17040 VDD.n1694 VDD.n1693 185
R17041 VDD.n1693 VDD.n552 185
R17042 VDD.n1695 VDD.n550 185
R17043 VDD.n1947 VDD.n550 185
R17044 VDD.n1697 VDD.n1696 185
R17045 VDD.n1696 VDD.n549 185
R17046 VDD.n1698 VDD.n557 185
R17047 VDD.n1941 VDD.n557 185
R17048 VDD.n1700 VDD.n1699 185
R17049 VDD.n1699 VDD.n556 185
R17050 VDD.n1701 VDD.n563 185
R17051 VDD.n1935 VDD.n563 185
R17052 VDD.n1703 VDD.n1702 185
R17053 VDD.n1702 VDD.n562 185
R17054 VDD.n1704 VDD.n569 185
R17055 VDD.n1929 VDD.n569 185
R17056 VDD.n1706 VDD.n1705 185
R17057 VDD.n1705 VDD.n568 185
R17058 VDD.n1707 VDD.n575 185
R17059 VDD.n1923 VDD.n575 185
R17060 VDD.n1709 VDD.n1708 185
R17061 VDD.n1708 VDD.n574 185
R17062 VDD.n1710 VDD.n581 185
R17063 VDD.n1917 VDD.n581 185
R17064 VDD.n1712 VDD.n1711 185
R17065 VDD.n1711 VDD.n580 185
R17066 VDD.n1713 VDD.n587 185
R17067 VDD.n1911 VDD.n587 185
R17068 VDD.n1715 VDD.n1714 185
R17069 VDD.n1714 VDD.n586 185
R17070 VDD.n1716 VDD.n593 185
R17071 VDD.n1905 VDD.n593 185
R17072 VDD.n1718 VDD.n1717 185
R17073 VDD.n1717 VDD.n592 185
R17074 VDD.n1719 VDD.n599 185
R17075 VDD.n1899 VDD.n599 185
R17076 VDD.n1721 VDD.n1720 185
R17077 VDD.n1720 VDD.n598 185
R17078 VDD.n1722 VDD.n605 185
R17079 VDD.n1893 VDD.n605 185
R17080 VDD.n1724 VDD.n1723 185
R17081 VDD.n1723 VDD.n604 185
R17082 VDD.n1725 VDD.n611 185
R17083 VDD.n1887 VDD.n611 185
R17084 VDD.n1727 VDD.n1726 185
R17085 VDD.n1726 VDD.n610 185
R17086 VDD.n1728 VDD.n617 185
R17087 VDD.n1881 VDD.n617 185
R17088 VDD.n1730 VDD.n1729 185
R17089 VDD.n1729 VDD.n616 185
R17090 VDD.n1731 VDD.n623 185
R17091 VDD.n1875 VDD.n623 185
R17092 VDD.n1733 VDD.n1732 185
R17093 VDD.n1732 VDD.n622 185
R17094 VDD.n1734 VDD.n629 185
R17095 VDD.n1869 VDD.n629 185
R17096 VDD.n1736 VDD.n1735 185
R17097 VDD.n1735 VDD.n628 185
R17098 VDD.n1737 VDD.n635 185
R17099 VDD.n1863 VDD.n635 185
R17100 VDD.n1739 VDD.n1738 185
R17101 VDD.n1738 VDD.n634 185
R17102 VDD.n1740 VDD.n641 185
R17103 VDD.n1857 VDD.n641 185
R17104 VDD.n1742 VDD.n1741 185
R17105 VDD.n1741 VDD.n640 185
R17106 VDD.n1743 VDD.n647 185
R17107 VDD.n1851 VDD.n647 185
R17108 VDD.n1745 VDD.n1744 185
R17109 VDD.n1744 VDD.n646 185
R17110 VDD.n1746 VDD.n652 185
R17111 VDD.n1845 VDD.n652 185
R17112 VDD.n1748 VDD.n1747 185
R17113 VDD.n1747 VDD.n660 185
R17114 VDD.n1749 VDD.n658 185
R17115 VDD.n1839 VDD.n658 185
R17116 VDD.n1751 VDD.n1750 185
R17117 VDD.n1750 VDD.n657 185
R17118 VDD.n1752 VDD.n664 185
R17119 VDD.n1833 VDD.n664 185
R17120 VDD.n1754 VDD.n1753 185
R17121 VDD.n1753 VDD.n672 185
R17122 VDD.n1755 VDD.n670 185
R17123 VDD.n1827 VDD.n670 185
R17124 VDD.n1757 VDD.n1756 185
R17125 VDD.n1756 VDD.n669 185
R17126 VDD.n1758 VDD.n677 185
R17127 VDD.n1821 VDD.n677 185
R17128 VDD.n1760 VDD.n1759 185
R17129 VDD.n1759 VDD.n676 185
R17130 VDD.n1761 VDD.n683 185
R17131 VDD.n1815 VDD.n683 185
R17132 VDD.n1763 VDD.n1762 185
R17133 VDD.n1762 VDD.n682 185
R17134 VDD.n1764 VDD.n689 185
R17135 VDD.n1809 VDD.n689 185
R17136 VDD.n1766 VDD.n1765 185
R17137 VDD.n1765 VDD.n688 185
R17138 VDD.n1767 VDD.n695 185
R17139 VDD.n1803 VDD.n695 185
R17140 VDD.n1769 VDD.n1768 185
R17141 VDD.n1769 VDD.n694 185
R17142 VDD.n2729 VDD.n166 185
R17143 VDD.n166 VDD.n163 185
R17144 VDD.n2731 VDD.n2730 185
R17145 VDD.n2732 VDD.n2731 185
R17146 VDD.n167 VDD.n165 185
R17147 VDD.n165 VDD.n161 185
R17148 VDD.n2693 VDD.n2692 185
R17149 VDD.n2694 VDD.n2693 185
R17150 VDD.n2691 VDD.n186 185
R17151 VDD.n186 VDD.n183 185
R17152 VDD.n2690 VDD.n2689 185
R17153 VDD.n2689 VDD.n2688 185
R17154 VDD.n188 VDD.n187 185
R17155 VDD.n189 VDD.n188 185
R17156 VDD.n2659 VDD.n2658 185
R17157 VDD.n2660 VDD.n2659 185
R17158 VDD.n2657 VDD.n199 185
R17159 VDD.n199 VDD.n196 185
R17160 VDD.n2656 VDD.n2655 185
R17161 VDD.n2655 VDD.n2654 185
R17162 VDD.n201 VDD.n200 185
R17163 VDD.n202 VDD.n201 185
R17164 VDD.n2647 VDD.n2646 185
R17165 VDD.n2648 VDD.n2647 185
R17166 VDD.n2645 VDD.n211 185
R17167 VDD.n211 VDD.n208 185
R17168 VDD.n2644 VDD.n2643 185
R17169 VDD.n2643 VDD.n2642 185
R17170 VDD.n213 VDD.n212 185
R17171 VDD.n214 VDD.n213 185
R17172 VDD.n2635 VDD.n2634 185
R17173 VDD.n2636 VDD.n2635 185
R17174 VDD.n2633 VDD.n223 185
R17175 VDD.n223 VDD.n220 185
R17176 VDD.n2632 VDD.n2631 185
R17177 VDD.n2631 VDD.n2630 185
R17178 VDD.n225 VDD.n224 185
R17179 VDD.n226 VDD.n225 185
R17180 VDD.n2623 VDD.n2622 185
R17181 VDD.n2624 VDD.n2623 185
R17182 VDD.n2621 VDD.n235 185
R17183 VDD.n235 VDD.n232 185
R17184 VDD.n2620 VDD.n2619 185
R17185 VDD.n2619 VDD.n2618 185
R17186 VDD.n237 VDD.n236 185
R17187 VDD.n238 VDD.n237 185
R17188 VDD.n2611 VDD.n2610 185
R17189 VDD.n2612 VDD.n2611 185
R17190 VDD.n2609 VDD.n247 185
R17191 VDD.n247 VDD.n244 185
R17192 VDD.n2608 VDD.n2607 185
R17193 VDD.n2607 VDD.n2606 185
R17194 VDD.n249 VDD.n248 185
R17195 VDD.n250 VDD.n249 185
R17196 VDD.n2599 VDD.n2598 185
R17197 VDD.n2600 VDD.n2599 185
R17198 VDD.n2597 VDD.n259 185
R17199 VDD.n259 VDD.n256 185
R17200 VDD.n2596 VDD.n2595 185
R17201 VDD.n2595 VDD.n2594 185
R17202 VDD.n261 VDD.n260 185
R17203 VDD.n262 VDD.n261 185
R17204 VDD.n2587 VDD.n2586 185
R17205 VDD.n2588 VDD.n2587 185
R17206 VDD.n2585 VDD.n270 185
R17207 VDD.n275 VDD.n270 185
R17208 VDD.n2584 VDD.n2583 185
R17209 VDD.n2583 VDD.n2582 185
R17210 VDD.n272 VDD.n271 185
R17211 VDD.n282 VDD.n272 185
R17212 VDD.n2575 VDD.n2574 185
R17213 VDD.n2576 VDD.n2575 185
R17214 VDD.n2573 VDD.n283 185
R17215 VDD.n283 VDD.n279 185
R17216 VDD.n2572 VDD.n2571 185
R17217 VDD.n2571 VDD.n2570 185
R17218 VDD.n285 VDD.n284 185
R17219 VDD.n286 VDD.n285 185
R17220 VDD.n2563 VDD.n2562 185
R17221 VDD.n2564 VDD.n2563 185
R17222 VDD.n2561 VDD.n295 185
R17223 VDD.n295 VDD.n292 185
R17224 VDD.n2560 VDD.n2559 185
R17225 VDD.n2559 VDD.n2558 185
R17226 VDD.n297 VDD.n296 185
R17227 VDD.n298 VDD.n297 185
R17228 VDD.n2551 VDD.n2550 185
R17229 VDD.n2552 VDD.n2551 185
R17230 VDD.n2549 VDD.n307 185
R17231 VDD.n307 VDD.n304 185
R17232 VDD.n2548 VDD.n2547 185
R17233 VDD.n2547 VDD.n2546 185
R17234 VDD.n309 VDD.n308 185
R17235 VDD.n310 VDD.n309 185
R17236 VDD.n2539 VDD.n2538 185
R17237 VDD.n2540 VDD.n2539 185
R17238 VDD.n2537 VDD.n319 185
R17239 VDD.n319 VDD.n316 185
R17240 VDD.n2536 VDD.n2535 185
R17241 VDD.n2535 VDD.n2534 185
R17242 VDD.n321 VDD.n320 185
R17243 VDD.n322 VDD.n321 185
R17244 VDD.n2527 VDD.n2526 185
R17245 VDD.n2528 VDD.n2527 185
R17246 VDD.n2525 VDD.n330 185
R17247 VDD.n336 VDD.n330 185
R17248 VDD.n2524 VDD.n2523 185
R17249 VDD.n2523 VDD.n2522 185
R17250 VDD.n332 VDD.n331 185
R17251 VDD.n333 VDD.n332 185
R17252 VDD.n2515 VDD.n2514 185
R17253 VDD.n2516 VDD.n2515 185
R17254 VDD.n2513 VDD.n343 185
R17255 VDD.n343 VDD.n340 185
R17256 VDD.n2512 VDD.n2511 185
R17257 VDD.n2511 VDD.n2510 185
R17258 VDD.n345 VDD.n344 185
R17259 VDD.n346 VDD.n345 185
R17260 VDD.n2503 VDD.n2502 185
R17261 VDD.n2504 VDD.n2503 185
R17262 VDD.n2501 VDD.n355 185
R17263 VDD.n355 VDD.n352 185
R17264 VDD.n2500 VDD.n2499 185
R17265 VDD.n2499 VDD.n2498 185
R17266 VDD.n357 VDD.n356 185
R17267 VDD.n358 VDD.n357 185
R17268 VDD.n2491 VDD.n2490 185
R17269 VDD.n2492 VDD.n2491 185
R17270 VDD.n2489 VDD.n367 185
R17271 VDD.n367 VDD.n364 185
R17272 VDD.n2488 VDD.n2487 185
R17273 VDD.n2487 VDD.n2486 185
R17274 VDD.n369 VDD.n368 185
R17275 VDD.n370 VDD.n369 185
R17276 VDD.n2479 VDD.n2478 185
R17277 VDD.n2480 VDD.n2479 185
R17278 VDD.n2477 VDD.n379 185
R17279 VDD.n379 VDD.n376 185
R17280 VDD.n2476 VDD.n2475 185
R17281 VDD.n2475 VDD.n2474 185
R17282 VDD.n381 VDD.n380 185
R17283 VDD.n389 VDD.n381 185
R17284 VDD.n2467 VDD.n2466 185
R17285 VDD.n2468 VDD.n2467 185
R17286 VDD.n2465 VDD.n390 185
R17287 VDD.n396 VDD.n390 185
R17288 VDD.n2464 VDD.n2463 185
R17289 VDD.n2463 VDD.n2462 185
R17290 VDD.n392 VDD.n391 185
R17291 VDD.n393 VDD.n392 185
R17292 VDD.n2455 VDD.n2454 185
R17293 VDD.n2456 VDD.n2455 185
R17294 VDD.n2453 VDD.n403 185
R17295 VDD.n403 VDD.n400 185
R17296 VDD.n2452 VDD.n2451 185
R17297 VDD.n2451 VDD.n2450 185
R17298 VDD.n405 VDD.n404 185
R17299 VDD.n406 VDD.n405 185
R17300 VDD.n2443 VDD.n2442 185
R17301 VDD.n2444 VDD.n2443 185
R17302 VDD.n2441 VDD.n415 185
R17303 VDD.n415 VDD.n412 185
R17304 VDD.n2440 VDD.n2439 185
R17305 VDD.n2439 VDD.n2438 185
R17306 VDD.n417 VDD.n416 185
R17307 VDD.n418 VDD.n417 185
R17308 VDD.n2429 VDD.n2428 185
R17309 VDD.n2427 VDD.n2280 185
R17310 VDD.n2426 VDD.n2279 185
R17311 VDD.n2431 VDD.n2279 185
R17312 VDD.n2425 VDD.n2424 185
R17313 VDD.n2423 VDD.n2422 185
R17314 VDD.n2421 VDD.n2420 185
R17315 VDD.n2419 VDD.n2418 185
R17316 VDD.n2417 VDD.n2416 185
R17317 VDD.n2415 VDD.n2414 185
R17318 VDD.n2413 VDD.n2412 185
R17319 VDD.n2411 VDD.n2410 185
R17320 VDD.n2409 VDD.n2408 185
R17321 VDD.n2406 VDD.n2405 185
R17322 VDD.n2404 VDD.n2403 185
R17323 VDD.n2402 VDD.n2401 185
R17324 VDD.n2701 VDD.n2700 185
R17325 VDD.n2703 VDD.n178 185
R17326 VDD.n2705 VDD.n2704 185
R17327 VDD.n2707 VDD.n175 185
R17328 VDD.n2709 VDD.n2708 185
R17329 VDD.n2711 VDD.n173 185
R17330 VDD.n2713 VDD.n2712 185
R17331 VDD.n2715 VDD.n172 185
R17332 VDD.n2717 VDD.n2716 185
R17333 VDD.n2719 VDD.n170 185
R17334 VDD.n2721 VDD.n2720 185
R17335 VDD.n2722 VDD.n169 185
R17336 VDD.n2724 VDD.n2723 185
R17337 VDD.n2726 VDD.n168 185
R17338 VDD.n2728 VDD.n2727 185
R17339 VDD.n2727 VDD.n151 185
R17340 VDD.n2699 VDD.n180 185
R17341 VDD.n180 VDD.n163 185
R17342 VDD.n2698 VDD.n162 185
R17343 VDD.n2732 VDD.n162 185
R17344 VDD.n2697 VDD.n2696 185
R17345 VDD.n2696 VDD.n161 185
R17346 VDD.n2695 VDD.n181 185
R17347 VDD.n2695 VDD.n2694 185
R17348 VDD.n2283 VDD.n182 185
R17349 VDD.n183 VDD.n182 185
R17350 VDD.n2284 VDD.n190 185
R17351 VDD.n2688 VDD.n190 185
R17352 VDD.n2286 VDD.n2285 185
R17353 VDD.n2285 VDD.n189 185
R17354 VDD.n2287 VDD.n197 185
R17355 VDD.n2660 VDD.n197 185
R17356 VDD.n2289 VDD.n2288 185
R17357 VDD.n2288 VDD.n196 185
R17358 VDD.n2290 VDD.n203 185
R17359 VDD.n2654 VDD.n203 185
R17360 VDD.n2292 VDD.n2291 185
R17361 VDD.n2291 VDD.n202 185
R17362 VDD.n2293 VDD.n209 185
R17363 VDD.n2648 VDD.n209 185
R17364 VDD.n2295 VDD.n2294 185
R17365 VDD.n2294 VDD.n208 185
R17366 VDD.n2296 VDD.n215 185
R17367 VDD.n2642 VDD.n215 185
R17368 VDD.n2298 VDD.n2297 185
R17369 VDD.n2297 VDD.n214 185
R17370 VDD.n2299 VDD.n221 185
R17371 VDD.n2636 VDD.n221 185
R17372 VDD.n2301 VDD.n2300 185
R17373 VDD.n2300 VDD.n220 185
R17374 VDD.n2302 VDD.n227 185
R17375 VDD.n2630 VDD.n227 185
R17376 VDD.n2304 VDD.n2303 185
R17377 VDD.n2303 VDD.n226 185
R17378 VDD.n2305 VDD.n233 185
R17379 VDD.n2624 VDD.n233 185
R17380 VDD.n2307 VDD.n2306 185
R17381 VDD.n2306 VDD.n232 185
R17382 VDD.n2308 VDD.n239 185
R17383 VDD.n2618 VDD.n239 185
R17384 VDD.n2310 VDD.n2309 185
R17385 VDD.n2309 VDD.n238 185
R17386 VDD.n2311 VDD.n245 185
R17387 VDD.n2612 VDD.n245 185
R17388 VDD.n2313 VDD.n2312 185
R17389 VDD.n2312 VDD.n244 185
R17390 VDD.n2314 VDD.n251 185
R17391 VDD.n2606 VDD.n251 185
R17392 VDD.n2316 VDD.n2315 185
R17393 VDD.n2315 VDD.n250 185
R17394 VDD.n2317 VDD.n257 185
R17395 VDD.n2600 VDD.n257 185
R17396 VDD.n2319 VDD.n2318 185
R17397 VDD.n2318 VDD.n256 185
R17398 VDD.n2320 VDD.n263 185
R17399 VDD.n2594 VDD.n263 185
R17400 VDD.n2322 VDD.n2321 185
R17401 VDD.n2321 VDD.n262 185
R17402 VDD.n2323 VDD.n268 185
R17403 VDD.n2588 VDD.n268 185
R17404 VDD.n2325 VDD.n2324 185
R17405 VDD.n2324 VDD.n275 185
R17406 VDD.n2326 VDD.n273 185
R17407 VDD.n2582 VDD.n273 185
R17408 VDD.n2328 VDD.n2327 185
R17409 VDD.n2327 VDD.n282 185
R17410 VDD.n2329 VDD.n280 185
R17411 VDD.n2576 VDD.n280 185
R17412 VDD.n2331 VDD.n2330 185
R17413 VDD.n2330 VDD.n279 185
R17414 VDD.n2332 VDD.n287 185
R17415 VDD.n2570 VDD.n287 185
R17416 VDD.n2334 VDD.n2333 185
R17417 VDD.n2333 VDD.n286 185
R17418 VDD.n2335 VDD.n293 185
R17419 VDD.n2564 VDD.n293 185
R17420 VDD.n2337 VDD.n2336 185
R17421 VDD.n2336 VDD.n292 185
R17422 VDD.n2338 VDD.n299 185
R17423 VDD.n2558 VDD.n299 185
R17424 VDD.n2340 VDD.n2339 185
R17425 VDD.n2339 VDD.n298 185
R17426 VDD.n2341 VDD.n305 185
R17427 VDD.n2552 VDD.n305 185
R17428 VDD.n2343 VDD.n2342 185
R17429 VDD.n2342 VDD.n304 185
R17430 VDD.n2344 VDD.n311 185
R17431 VDD.n2546 VDD.n311 185
R17432 VDD.n2346 VDD.n2345 185
R17433 VDD.n2345 VDD.n310 185
R17434 VDD.n2347 VDD.n317 185
R17435 VDD.n2540 VDD.n317 185
R17436 VDD.n2349 VDD.n2348 185
R17437 VDD.n2348 VDD.n316 185
R17438 VDD.n2350 VDD.n323 185
R17439 VDD.n2534 VDD.n323 185
R17440 VDD.n2352 VDD.n2351 185
R17441 VDD.n2351 VDD.n322 185
R17442 VDD.n2353 VDD.n328 185
R17443 VDD.n2528 VDD.n328 185
R17444 VDD.n2355 VDD.n2354 185
R17445 VDD.n2354 VDD.n336 185
R17446 VDD.n2356 VDD.n334 185
R17447 VDD.n2522 VDD.n334 185
R17448 VDD.n2358 VDD.n2357 185
R17449 VDD.n2357 VDD.n333 185
R17450 VDD.n2359 VDD.n341 185
R17451 VDD.n2516 VDD.n341 185
R17452 VDD.n2361 VDD.n2360 185
R17453 VDD.n2360 VDD.n340 185
R17454 VDD.n2362 VDD.n347 185
R17455 VDD.n2510 VDD.n347 185
R17456 VDD.n2364 VDD.n2363 185
R17457 VDD.n2363 VDD.n346 185
R17458 VDD.n2365 VDD.n353 185
R17459 VDD.n2504 VDD.n353 185
R17460 VDD.n2367 VDD.n2366 185
R17461 VDD.n2366 VDD.n352 185
R17462 VDD.n2368 VDD.n359 185
R17463 VDD.n2498 VDD.n359 185
R17464 VDD.n2370 VDD.n2369 185
R17465 VDD.n2369 VDD.n358 185
R17466 VDD.n2371 VDD.n365 185
R17467 VDD.n2492 VDD.n365 185
R17468 VDD.n2373 VDD.n2372 185
R17469 VDD.n2372 VDD.n364 185
R17470 VDD.n2374 VDD.n371 185
R17471 VDD.n2486 VDD.n371 185
R17472 VDD.n2376 VDD.n2375 185
R17473 VDD.n2375 VDD.n370 185
R17474 VDD.n2377 VDD.n377 185
R17475 VDD.n2480 VDD.n377 185
R17476 VDD.n2379 VDD.n2378 185
R17477 VDD.n2378 VDD.n376 185
R17478 VDD.n2380 VDD.n382 185
R17479 VDD.n2474 VDD.n382 185
R17480 VDD.n2382 VDD.n2381 185
R17481 VDD.n2381 VDD.n389 185
R17482 VDD.n2383 VDD.n387 185
R17483 VDD.n2468 VDD.n387 185
R17484 VDD.n2385 VDD.n2384 185
R17485 VDD.n2384 VDD.n396 185
R17486 VDD.n2386 VDD.n394 185
R17487 VDD.n2462 VDD.n394 185
R17488 VDD.n2388 VDD.n2387 185
R17489 VDD.n2387 VDD.n393 185
R17490 VDD.n2389 VDD.n401 185
R17491 VDD.n2456 VDD.n401 185
R17492 VDD.n2391 VDD.n2390 185
R17493 VDD.n2390 VDD.n400 185
R17494 VDD.n2392 VDD.n407 185
R17495 VDD.n2450 VDD.n407 185
R17496 VDD.n2394 VDD.n2393 185
R17497 VDD.n2393 VDD.n406 185
R17498 VDD.n2395 VDD.n413 185
R17499 VDD.n2444 VDD.n413 185
R17500 VDD.n2397 VDD.n2396 185
R17501 VDD.n2396 VDD.n412 185
R17502 VDD.n2398 VDD.n419 185
R17503 VDD.n2438 VDD.n419 185
R17504 VDD.n2400 VDD.n2399 185
R17505 VDD.n2400 VDD.n418 185
R17506 VDD.n1555 VDD.n1554 185
R17507 VDD.n1556 VDD.n1555 185
R17508 VDD.n963 VDD.n961 185
R17509 VDD.n961 VDD.n960 185
R17510 VDD.n1489 VDD.n1488 185
R17511 VDD.n1488 VDD.n1487 185
R17512 VDD.n966 VDD.n965 185
R17513 VDD.n967 VDD.n966 185
R17514 VDD.n1475 VDD.n1474 185
R17515 VDD.n1476 VDD.n1475 185
R17516 VDD.n976 VDD.n975 185
R17517 VDD.n975 VDD.n974 185
R17518 VDD.n1470 VDD.n1469 185
R17519 VDD.n1469 VDD.n1468 185
R17520 VDD.n979 VDD.n978 185
R17521 VDD.n980 VDD.n979 185
R17522 VDD.n1459 VDD.n1458 185
R17523 VDD.n1460 VDD.n1459 185
R17524 VDD.n988 VDD.n987 185
R17525 VDD.n987 VDD.n986 185
R17526 VDD.n1454 VDD.n1453 185
R17527 VDD.n1453 VDD.n1452 185
R17528 VDD.n991 VDD.n990 185
R17529 VDD.n992 VDD.n991 185
R17530 VDD.n1443 VDD.n1442 185
R17531 VDD.n1444 VDD.n1443 185
R17532 VDD.n999 VDD.n998 185
R17533 VDD.n998 VDD.t98 185
R17534 VDD.n1338 VDD.n1337 185
R17535 VDD.n1337 VDD.n1336 185
R17536 VDD.n1002 VDD.n1001 185
R17537 VDD.n1003 VDD.n1002 185
R17538 VDD.n1327 VDD.n1326 185
R17539 VDD.n1328 VDD.n1327 185
R17540 VDD.n1011 VDD.n1010 185
R17541 VDD.n1010 VDD.n1009 185
R17542 VDD.n1322 VDD.n1321 185
R17543 VDD.n1321 VDD.n1320 185
R17544 VDD.n1014 VDD.n1013 185
R17545 VDD.n1015 VDD.n1014 185
R17546 VDD.n1311 VDD.n1310 185
R17547 VDD.n1312 VDD.n1311 185
R17548 VDD.n1023 VDD.n1022 185
R17549 VDD.n1022 VDD.n1021 185
R17550 VDD.n1306 VDD.n1305 185
R17551 VDD.n1305 VDD.n1304 185
R17552 VDD.n1026 VDD.n1025 185
R17553 VDD.n1033 VDD.n1026 185
R17554 VDD.n1295 VDD.n1294 185
R17555 VDD.n1296 VDD.n1295 185
R17556 VDD.n1035 VDD.n1034 185
R17557 VDD.n1034 VDD.n1032 185
R17558 VDD.n1290 VDD.n1289 185
R17559 VDD.n1289 VDD.n1288 185
R17560 VDD.n1120 VDD.n1037 185
R17561 VDD.n1123 VDD.n1122 185
R17562 VDD.n1119 VDD.n1118 185
R17563 VDD.n1118 VDD.n1038 185
R17564 VDD.n1128 VDD.n1127 185
R17565 VDD.n1130 VDD.n1117 185
R17566 VDD.n1133 VDD.n1132 185
R17567 VDD.n1115 VDD.n1114 185
R17568 VDD.n1140 VDD.n1139 185
R17569 VDD.n1142 VDD.n1113 185
R17570 VDD.n1143 VDD.n1112 185
R17571 VDD.n1146 VDD.n1145 185
R17572 VDD.n1147 VDD.n1109 185
R17573 VDD.n1106 VDD.n1105 185
R17574 VDD.n1152 VDD.n1151 185
R17575 VDD.n1154 VDD.n1104 185
R17576 VDD.n1157 VDD.n1156 185
R17577 VDD.n1102 VDD.n1101 185
R17578 VDD.n1162 VDD.n1161 185
R17579 VDD.n1164 VDD.n1100 185
R17580 VDD.n1167 VDD.n1166 185
R17581 VDD.n1098 VDD.n1097 185
R17582 VDD.n1174 VDD.n1173 185
R17583 VDD.n1176 VDD.n1096 185
R17584 VDD.n1177 VDD.n1095 185
R17585 VDD.n1180 VDD.n1179 185
R17586 VDD.n1181 VDD.n1092 185
R17587 VDD.n1089 VDD.n1088 185
R17588 VDD.n1186 VDD.n1185 185
R17589 VDD.n1188 VDD.n1087 185
R17590 VDD.n1191 VDD.n1190 185
R17591 VDD.n1085 VDD.n1084 185
R17592 VDD.n1196 VDD.n1195 185
R17593 VDD.n1198 VDD.n1083 185
R17594 VDD.n1201 VDD.n1200 185
R17595 VDD.n1081 VDD.n1080 185
R17596 VDD.n1208 VDD.n1207 185
R17597 VDD.n1210 VDD.n1079 185
R17598 VDD.n1211 VDD.n1078 185
R17599 VDD.n1214 VDD.n1213 185
R17600 VDD.n1215 VDD.n1075 185
R17601 VDD.n1072 VDD.n1071 185
R17602 VDD.n1220 VDD.n1219 185
R17603 VDD.n1222 VDD.n1070 185
R17604 VDD.n1225 VDD.n1224 185
R17605 VDD.n1068 VDD.n1067 185
R17606 VDD.n1230 VDD.n1229 185
R17607 VDD.n1232 VDD.n1066 185
R17608 VDD.n1235 VDD.n1234 185
R17609 VDD.n1064 VDD.n1063 185
R17610 VDD.n1241 VDD.n1240 185
R17611 VDD.n1243 VDD.n1062 185
R17612 VDD.n1246 VDD.n1245 185
R17613 VDD.n1247 VDD.n1057 185
R17614 VDD.n1251 VDD.n1250 185
R17615 VDD.n1253 VDD.n1056 185
R17616 VDD.n1256 VDD.n1255 185
R17617 VDD.n1054 VDD.n1053 185
R17618 VDD.n1261 VDD.n1260 185
R17619 VDD.n1263 VDD.n1052 185
R17620 VDD.n1266 VDD.n1265 185
R17621 VDD.n1050 VDD.n1049 185
R17622 VDD.n1271 VDD.n1270 185
R17623 VDD.n1273 VDD.n1048 185
R17624 VDD.n1277 VDD.n1276 185
R17625 VDD.n1274 VDD.n1044 185
R17626 VDD.n1281 VDD.n1046 185
R17627 VDD.n1282 VDD.n1041 185
R17628 VDD.n1283 VDD.n1039 185
R17629 VDD.n1039 VDD.n1038 185
R17630 VDD.n1558 VDD.n955 185
R17631 VDD.n1561 VDD.n1560 185
R17632 VDD.n1562 VDD.n954 185
R17633 VDD.n952 VDD.n950 185
R17634 VDD.n1566 VDD.n949 185
R17635 VDD.n1567 VDD.n947 185
R17636 VDD.n1568 VDD.n946 185
R17637 VDD.n944 VDD.n942 185
R17638 VDD.n1572 VDD.n941 185
R17639 VDD.n1573 VDD.n939 185
R17640 VDD.n1574 VDD.n938 185
R17641 VDD.n936 VDD.n934 185
R17642 VDD.n1578 VDD.n933 185
R17643 VDD.n1579 VDD.n931 185
R17644 VDD.n1580 VDD.n930 185
R17645 VDD.n1583 VDD.n924 185
R17646 VDD.n1584 VDD.n923 185
R17647 VDD.n1585 VDD.n921 185
R17648 VDD.n920 VDD.n918 185
R17649 VDD.n768 VDD.n767 185
R17650 VDD.n1590 VDD.n1589 185
R17651 VDD.n1592 VDD.n765 185
R17652 VDD.n1594 VDD.n1593 185
R17653 VDD.n1595 VDD.n761 185
R17654 VDD.n1597 VDD.n1596 185
R17655 VDD.n1599 VDD.n758 185
R17656 VDD.n1601 VDD.n1600 185
R17657 VDD.n759 VDD.n752 185
R17658 VDD.n1605 VDD.n756 185
R17659 VDD.n1606 VDD.n748 185
R17660 VDD.n1608 VDD.n1607 185
R17661 VDD.n1610 VDD.n746 185
R17662 VDD.n1612 VDD.n1611 185
R17663 VDD.n1613 VDD.n741 185
R17664 VDD.n1615 VDD.n1614 185
R17665 VDD.n1617 VDD.n739 185
R17666 VDD.n1619 VDD.n1618 185
R17667 VDD.n1620 VDD.n735 185
R17668 VDD.n1622 VDD.n1621 185
R17669 VDD.n1624 VDD.n733 185
R17670 VDD.n1626 VDD.n1625 185
R17671 VDD.n728 VDD.n727 185
R17672 VDD.n1631 VDD.n1630 185
R17673 VDD.n1633 VDD.n725 185
R17674 VDD.n1635 VDD.n1634 185
R17675 VDD.n1636 VDD.n723 185
R17676 VDD.n1638 VDD.n1637 185
R17677 VDD.n1640 VDD.n722 185
R17678 VDD.n1641 VDD.n718 185
R17679 VDD.n1644 VDD.n1643 185
R17680 VDD.n720 VDD.n719 185
R17681 VDD.n1524 VDD.n1519 185
R17682 VDD.n1526 VDD.n1525 185
R17683 VDD.n1528 VDD.n1517 185
R17684 VDD.n1529 VDD.n1516 185
R17685 VDD.n1532 VDD.n1531 185
R17686 VDD.n1533 VDD.n1513 185
R17687 VDD.n1534 VDD.n1506 185
R17688 VDD.n1536 VDD.n1535 185
R17689 VDD.n1538 VDD.n1504 185
R17690 VDD.n1540 VDD.n1539 185
R17691 VDD.n1541 VDD.n1498 185
R17692 VDD.n1543 VDD.n1542 185
R17693 VDD.n1545 VDD.n1497 185
R17694 VDD.n1546 VDD.n1496 185
R17695 VDD.n1549 VDD.n1548 185
R17696 VDD.n1550 VDD.n1494 185
R17697 VDD.n1551 VDD.n962 185
R17698 VDD.n1557 VDD.n959 185
R17699 VDD.n1557 VDD.n1556 185
R17700 VDD.n970 VDD.n958 185
R17701 VDD.n960 VDD.n958 185
R17702 VDD.n1486 VDD.n1485 185
R17703 VDD.n1487 VDD.n1486 185
R17704 VDD.n969 VDD.n968 185
R17705 VDD.n968 VDD.n967 185
R17706 VDD.n1478 VDD.n1477 185
R17707 VDD.n1477 VDD.n1476 185
R17708 VDD.n973 VDD.n972 185
R17709 VDD.n974 VDD.n973 185
R17710 VDD.n1467 VDD.n1466 185
R17711 VDD.n1468 VDD.n1467 185
R17712 VDD.n982 VDD.n981 185
R17713 VDD.n981 VDD.n980 185
R17714 VDD.n1462 VDD.n1461 185
R17715 VDD.n1461 VDD.n1460 185
R17716 VDD.n985 VDD.n984 185
R17717 VDD.n986 VDD.n985 185
R17718 VDD.n1451 VDD.n1450 185
R17719 VDD.n1452 VDD.n1451 185
R17720 VDD.n994 VDD.n993 185
R17721 VDD.n993 VDD.n992 185
R17722 VDD.n1446 VDD.n1445 185
R17723 VDD.n1445 VDD.n1444 185
R17724 VDD.n997 VDD.n996 185
R17725 VDD.t98 VDD.n997 185
R17726 VDD.n1335 VDD.n1334 185
R17727 VDD.n1336 VDD.n1335 185
R17728 VDD.n1005 VDD.n1004 185
R17729 VDD.n1004 VDD.n1003 185
R17730 VDD.n1330 VDD.n1329 185
R17731 VDD.n1329 VDD.n1328 185
R17732 VDD.n1008 VDD.n1007 185
R17733 VDD.n1009 VDD.n1008 185
R17734 VDD.n1319 VDD.n1318 185
R17735 VDD.n1320 VDD.n1319 185
R17736 VDD.n1017 VDD.n1016 185
R17737 VDD.n1016 VDD.n1015 185
R17738 VDD.n1314 VDD.n1313 185
R17739 VDD.n1313 VDD.n1312 185
R17740 VDD.n1020 VDD.n1019 185
R17741 VDD.n1021 VDD.n1020 185
R17742 VDD.n1303 VDD.n1302 185
R17743 VDD.n1304 VDD.n1303 185
R17744 VDD.n1028 VDD.n1027 185
R17745 VDD.n1033 VDD.n1027 185
R17746 VDD.n1298 VDD.n1297 185
R17747 VDD.n1297 VDD.n1296 185
R17748 VDD.n1031 VDD.n1030 185
R17749 VDD.n1032 VDD.n1031 185
R17750 VDD.n1287 VDD.n1286 185
R17751 VDD.n1288 VDD.n1287 185
R17752 VDD.n2907 VDD.n2906 185
R17753 VDD.n2905 VDD.n101 185
R17754 VDD.n2904 VDD.n100 185
R17755 VDD.n2909 VDD.n100 185
R17756 VDD.n2903 VDD.n2902 185
R17757 VDD.n2901 VDD.n2900 185
R17758 VDD.n2899 VDD.n2898 185
R17759 VDD.n2897 VDD.n2896 185
R17760 VDD.n2895 VDD.n2894 185
R17761 VDD.n2893 VDD.n2892 185
R17762 VDD.n2891 VDD.n2890 185
R17763 VDD.n2889 VDD.n2888 185
R17764 VDD.n2887 VDD.n2886 185
R17765 VDD.n2885 VDD.n2884 185
R17766 VDD.n2883 VDD.n2882 185
R17767 VDD.n2881 VDD.n2880 185
R17768 VDD.n2879 VDD.n2878 185
R17769 VDD.n2877 VDD.n2876 185
R17770 VDD.n2875 VDD.n2874 185
R17771 VDD.n2873 VDD.n2872 185
R17772 VDD.n2871 VDD.n2870 185
R17773 VDD.n2869 VDD.n2868 185
R17774 VDD.n2867 VDD.n2866 185
R17775 VDD.n2865 VDD.n2864 185
R17776 VDD.n2863 VDD.n2862 185
R17777 VDD.n2861 VDD.n2860 185
R17778 VDD.n2859 VDD.n2858 185
R17779 VDD.n2850 VDD.n127 185
R17780 VDD.n2852 VDD.n2851 185
R17781 VDD.n2849 VDD.n2848 185
R17782 VDD.n2847 VDD.n2846 185
R17783 VDD.n2845 VDD.n2844 185
R17784 VDD.n2843 VDD.n2842 185
R17785 VDD.n2841 VDD.n2840 185
R17786 VDD.n2839 VDD.n2838 185
R17787 VDD.n2837 VDD.n2836 185
R17788 VDD.n2835 VDD.n2834 185
R17789 VDD.n2833 VDD.n2832 185
R17790 VDD.n2831 VDD.n2830 185
R17791 VDD.n2829 VDD.n2828 185
R17792 VDD.n2827 VDD.n2826 185
R17793 VDD.n2820 VDD.n139 185
R17794 VDD.n2822 VDD.n2821 185
R17795 VDD.n2819 VDD.n2818 185
R17796 VDD.n2817 VDD.n2816 185
R17797 VDD.n2815 VDD.n2814 185
R17798 VDD.n2813 VDD.n2812 185
R17799 VDD.n2811 VDD.n2810 185
R17800 VDD.n2809 VDD.n2808 185
R17801 VDD.n2807 VDD.n2806 185
R17802 VDD.n2805 VDD.n2804 185
R17803 VDD.n2803 VDD.n2802 185
R17804 VDD.n2801 VDD.n2800 185
R17805 VDD.n2799 VDD.n2798 185
R17806 VDD.n2797 VDD.n2796 185
R17807 VDD.n2795 VDD.n2794 185
R17808 VDD.n2793 VDD.n2792 185
R17809 VDD.n2791 VDD.n2790 185
R17810 VDD.n2789 VDD.n2788 185
R17811 VDD.n2787 VDD.n2786 185
R17812 VDD.n2785 VDD.n2784 185
R17813 VDD.n2783 VDD.n2782 185
R17814 VDD.n2781 VDD.n2780 185
R17815 VDD.n2779 VDD.n2778 185
R17816 VDD.n2777 VDD.n2776 185
R17817 VDD.n2775 VDD.n2774 185
R17818 VDD.n2773 VDD.n2772 185
R17819 VDD.n67 VDD.n66 185
R17820 VDD.n2911 VDD.n2910 185
R17821 VDD.n2910 VDD.n2909 185
R17822 VDD.n3269 VDD.n3268 185
R17823 VDD.n3034 VDD.n3031 185
R17824 VDD.n3241 VDD.n3240 185
R17825 VDD.n3239 VDD.n3238 185
R17826 VDD.n3237 VDD.n3236 185
R17827 VDD.n3230 VDD.n3036 185
R17828 VDD.n3232 VDD.n3231 185
R17829 VDD.n3229 VDD.n3228 185
R17830 VDD.n3227 VDD.n3226 185
R17831 VDD.n3220 VDD.n3038 185
R17832 VDD.n3222 VDD.n3221 185
R17833 VDD.n3219 VDD.n3218 185
R17834 VDD.n3217 VDD.n3216 185
R17835 VDD.n3210 VDD.n3040 185
R17836 VDD.n3212 VDD.n3211 185
R17837 VDD.n3208 VDD.n3207 185
R17838 VDD.n3206 VDD.n3205 185
R17839 VDD.n3199 VDD.n3044 185
R17840 VDD.n3201 VDD.n3200 185
R17841 VDD.n3198 VDD.n3197 185
R17842 VDD.n3196 VDD.n3195 185
R17843 VDD.n3189 VDD.n3046 185
R17844 VDD.n3191 VDD.n3190 185
R17845 VDD.n3188 VDD.n3187 185
R17846 VDD.n3186 VDD.n3185 185
R17847 VDD.n3179 VDD.n3048 185
R17848 VDD.n3181 VDD.n3180 185
R17849 VDD.n3178 VDD.n3177 185
R17850 VDD.n3176 VDD.n3175 185
R17851 VDD.n3174 VDD.n3173 185
R17852 VDD.n3172 VDD.n3053 185
R17853 VDD.n3168 VDD.n3167 185
R17854 VDD.n3166 VDD.n3165 185
R17855 VDD.n3164 VDD.n3163 185
R17856 VDD.n3162 VDD.n3055 185
R17857 VDD.n3158 VDD.n3157 185
R17858 VDD.n3156 VDD.n3155 185
R17859 VDD.n3154 VDD.n3153 185
R17860 VDD.n3152 VDD.n3057 185
R17861 VDD.n3148 VDD.n3147 185
R17862 VDD.n3146 VDD.n3145 185
R17863 VDD.n3144 VDD.n3143 185
R17864 VDD.n3142 VDD.n3061 185
R17865 VDD.n3138 VDD.n3137 185
R17866 VDD.n3136 VDD.n3135 185
R17867 VDD.n3134 VDD.n3133 185
R17868 VDD.n3132 VDD.n3063 185
R17869 VDD.n3128 VDD.n3127 185
R17870 VDD.n3126 VDD.n3125 185
R17871 VDD.n3124 VDD.n3123 185
R17872 VDD.n3122 VDD.n3065 185
R17873 VDD.n3118 VDD.n3117 185
R17874 VDD.n3116 VDD.n3115 185
R17875 VDD.n3114 VDD.n3113 185
R17876 VDD.n3112 VDD.n3067 185
R17877 VDD.n3108 VDD.n3107 185
R17878 VDD.n3106 VDD.n3105 185
R17879 VDD.n3104 VDD.n3103 185
R17880 VDD.n3102 VDD.n3071 185
R17881 VDD.n3098 VDD.n3097 185
R17882 VDD.n3096 VDD.n3095 185
R17883 VDD.n3094 VDD.n3093 185
R17884 VDD.n3092 VDD.n3073 185
R17885 VDD.n3088 VDD.n3087 185
R17886 VDD.n3086 VDD.n3085 185
R17887 VDD.n3084 VDD.n3083 185
R17888 VDD.n3082 VDD.n3075 185
R17889 VDD.n3078 VDD.n3077 185
R17890 VDD.n3265 VDD.n2997 185
R17891 VDD.n3272 VDD.n2997 185
R17892 VDD.n3264 VDD.n2996 185
R17893 VDD.n3273 VDD.n2996 185
R17894 VDD.n3263 VDD.n3262 185
R17895 VDD.n3262 VDD.n2988 185
R17896 VDD.n3245 VDD.n2987 185
R17897 VDD.n3279 VDD.n2987 185
R17898 VDD.n3258 VDD.n2986 185
R17899 VDD.n3280 VDD.n2986 185
R17900 VDD.n3257 VDD.n2985 185
R17901 VDD.n3281 VDD.n2985 185
R17902 VDD.n3256 VDD.n3255 185
R17903 VDD.n3255 VDD.n2977 185
R17904 VDD.n3247 VDD.n2976 185
R17905 VDD.n3287 VDD.n2976 185
R17906 VDD.n3251 VDD.n2975 185
R17907 VDD.n3288 VDD.n2975 185
R17908 VDD.n3250 VDD.n2974 185
R17909 VDD.n3289 VDD.n2974 185
R17910 VDD.n2966 VDD.n2965 185
R17911 VDD.n2967 VDD.n2966 185
R17912 VDD.n3297 VDD.n3296 185
R17913 VDD.n3296 VDD.n3295 185
R17914 VDD.n3298 VDD.n25 185
R17915 VDD.n25 VDD.n23 185
R17916 VDD.n3300 VDD.n3299 185
R17917 VDD.t126 VDD.n3300 185
R17918 VDD.n26 VDD.n24 185
R17919 VDD.n24 VDD.n22 185
R17920 VDD.n2959 VDD.n2958 185
R17921 VDD.n2958 VDD.n2957 185
R17922 VDD.n29 VDD.n28 185
R17923 VDD.n30 VDD.n29 185
R17924 VDD.n2948 VDD.n2947 185
R17925 VDD.n2949 VDD.n2948 185
R17926 VDD.n38 VDD.n37 185
R17927 VDD.n37 VDD.n36 185
R17928 VDD.n2943 VDD.n2942 185
R17929 VDD.n2942 VDD.n2941 185
R17930 VDD.n41 VDD.n40 185
R17931 VDD.n42 VDD.n41 185
R17932 VDD.n2932 VDD.n2931 185
R17933 VDD.n2933 VDD.n2932 185
R17934 VDD.n50 VDD.n49 185
R17935 VDD.n49 VDD.n48 185
R17936 VDD.n2927 VDD.n2926 185
R17937 VDD.n2926 VDD.n2925 185
R17938 VDD.n53 VDD.n52 185
R17939 VDD.n54 VDD.n53 185
R17940 VDD.n2916 VDD.n2915 185
R17941 VDD.n2917 VDD.n2916 185
R17942 VDD.n62 VDD.n61 185
R17943 VDD.n61 VDD.n60 185
R17944 VDD.n59 VDD.n58 185
R17945 VDD.n60 VDD.n59 185
R17946 VDD.n2919 VDD.n2918 185
R17947 VDD.n2918 VDD.n2917 185
R17948 VDD.n56 VDD.n55 185
R17949 VDD.n55 VDD.n54 185
R17950 VDD.n2924 VDD.n2923 185
R17951 VDD.n2925 VDD.n2924 185
R17952 VDD.n47 VDD.n46 185
R17953 VDD.n48 VDD.n47 185
R17954 VDD.n2935 VDD.n2934 185
R17955 VDD.n2934 VDD.n2933 185
R17956 VDD.n44 VDD.n43 185
R17957 VDD.n43 VDD.n42 185
R17958 VDD.n2940 VDD.n2939 185
R17959 VDD.n2941 VDD.n2940 185
R17960 VDD.n35 VDD.n34 185
R17961 VDD.n36 VDD.n35 185
R17962 VDD.n2951 VDD.n2950 185
R17963 VDD.n2950 VDD.n2949 185
R17964 VDD.n32 VDD.n31 185
R17965 VDD.n31 VDD.n30 185
R17966 VDD.n2956 VDD.n2955 185
R17967 VDD.n2957 VDD.n2956 185
R17968 VDD.n20 VDD.n18 185
R17969 VDD.n22 VDD.n20 185
R17970 VDD.n3302 VDD.n3301 185
R17971 VDD.n3301 VDD.t126 185
R17972 VDD.n21 VDD.n19 185
R17973 VDD.n23 VDD.n21 185
R17974 VDD.n3294 VDD.n3293 185
R17975 VDD.n3295 VDD.n3294 185
R17976 VDD.n3292 VDD.n2968 185
R17977 VDD.n2968 VDD.n2967 185
R17978 VDD.n3291 VDD.n3290 185
R17979 VDD.n3290 VDD.n3289 185
R17980 VDD.n2973 VDD.n2972 185
R17981 VDD.n3288 VDD.n2973 185
R17982 VDD.n3286 VDD.n3285 185
R17983 VDD.n3287 VDD.n3286 185
R17984 VDD.n3284 VDD.n2978 185
R17985 VDD.n2978 VDD.n2977 185
R17986 VDD.n3283 VDD.n3282 185
R17987 VDD.n3282 VDD.n3281 185
R17988 VDD.n2984 VDD.n2983 185
R17989 VDD.n3280 VDD.n2984 185
R17990 VDD.n3278 VDD.n3277 185
R17991 VDD.n3279 VDD.n3278 185
R17992 VDD.n3276 VDD.n2989 185
R17993 VDD.n2989 VDD.n2988 185
R17994 VDD.n3275 VDD.n3274 185
R17995 VDD.n3274 VDD.n3273 185
R17996 VDD.n2995 VDD.n2994 185
R17997 VDD.n3272 VDD.n2995 185
R17998 VDD.n2073 VDD.n2072 185
R17999 VDD.n2072 VDD.n424 185
R18000 VDD.n2074 VDD.n450 185
R18001 VDD.n2084 VDD.n450 185
R18002 VDD.n2075 VDD.n458 185
R18003 VDD.n458 VDD.n448 185
R18004 VDD.n2077 VDD.n2076 185
R18005 VDD.n2078 VDD.n2077 185
R18006 VDD.n459 VDD.n457 185
R18007 VDD.n457 VDD.n454 185
R18008 VDD.n2023 VDD.n467 185
R18009 VDD.n2033 VDD.n467 185
R18010 VDD.n2024 VDD.n475 185
R18011 VDD.n475 VDD.n465 185
R18012 VDD.n2026 VDD.n2025 185
R18013 VDD.n2027 VDD.n2026 185
R18014 VDD.n2022 VDD.n474 185
R18015 VDD.n474 VDD.n471 185
R18016 VDD.n2021 VDD.n2020 185
R18017 VDD.n2020 VDD.n2019 185
R18018 VDD.n477 VDD.n476 185
R18019 VDD.n478 VDD.n477 185
R18020 VDD.n2012 VDD.n2011 185
R18021 VDD.n2013 VDD.n2012 185
R18022 VDD.n2010 VDD.n487 185
R18023 VDD.n487 VDD.n484 185
R18024 VDD.n2009 VDD.n2008 185
R18025 VDD.n2008 VDD.n2007 185
R18026 VDD.n489 VDD.n488 185
R18027 VDD.n490 VDD.n489 185
R18028 VDD.n2000 VDD.n1999 185
R18029 VDD.n2001 VDD.n2000 185
R18030 VDD.n1998 VDD.n499 185
R18031 VDD.n499 VDD.n496 185
R18032 VDD.n1997 VDD.n1996 185
R18033 VDD.n1996 VDD.n1995 185
R18034 VDD.n501 VDD.n500 185
R18035 VDD.n502 VDD.n501 185
R18036 VDD.n1988 VDD.n1987 185
R18037 VDD.n1989 VDD.n1988 185
R18038 VDD.n1986 VDD.n511 185
R18039 VDD.n511 VDD.n508 185
R18040 VDD.n1985 VDD.n1984 185
R18041 VDD.n1984 VDD.n1983 185
R18042 VDD.n513 VDD.n512 185
R18043 VDD.n514 VDD.n513 185
R18044 VDD.n1976 VDD.n1975 185
R18045 VDD.n1977 VDD.n1976 185
R18046 VDD.n1974 VDD.n523 185
R18047 VDD.n523 VDD.n520 185
R18048 VDD.n1973 VDD.n1972 185
R18049 VDD.n1972 VDD.n1971 185
R18050 VDD.n525 VDD.n524 185
R18051 VDD.n526 VDD.n525 185
R18052 VDD.n1964 VDD.n1963 185
R18053 VDD.n1965 VDD.n1964 185
R18054 VDD.n1962 VDD.n535 185
R18055 VDD.n535 VDD.n532 185
R18056 VDD.n1961 VDD.n1960 185
R18057 VDD.n1960 VDD.n1959 185
R18058 VDD.n537 VDD.n536 185
R18059 VDD.n538 VDD.n537 185
R18060 VDD.n1952 VDD.n1951 185
R18061 VDD.n1953 VDD.n1952 185
R18062 VDD.n1950 VDD.n546 185
R18063 VDD.n552 VDD.n546 185
R18064 VDD.n1949 VDD.n1948 185
R18065 VDD.n1948 VDD.n1947 185
R18066 VDD.n548 VDD.n547 185
R18067 VDD.n549 VDD.n548 185
R18068 VDD.n1940 VDD.n1939 185
R18069 VDD.n1941 VDD.n1940 185
R18070 VDD.n1938 VDD.n559 185
R18071 VDD.n559 VDD.n556 185
R18072 VDD.n1937 VDD.n1936 185
R18073 VDD.n1936 VDD.n1935 185
R18074 VDD.n561 VDD.n560 185
R18075 VDD.n562 VDD.n561 185
R18076 VDD.n1928 VDD.n1927 185
R18077 VDD.n1929 VDD.n1928 185
R18078 VDD.n1926 VDD.n571 185
R18079 VDD.n571 VDD.n568 185
R18080 VDD.n1925 VDD.n1924 185
R18081 VDD.n1924 VDD.n1923 185
R18082 VDD.n573 VDD.n572 185
R18083 VDD.n574 VDD.n573 185
R18084 VDD.n1916 VDD.n1915 185
R18085 VDD.n1917 VDD.n1916 185
R18086 VDD.n1914 VDD.n583 185
R18087 VDD.n583 VDD.n580 185
R18088 VDD.n1913 VDD.n1912 185
R18089 VDD.n1912 VDD.n1911 185
R18090 VDD.n585 VDD.n584 185
R18091 VDD.n586 VDD.n585 185
R18092 VDD.n1904 VDD.n1903 185
R18093 VDD.n1905 VDD.n1904 185
R18094 VDD.n1902 VDD.n595 185
R18095 VDD.n595 VDD.n592 185
R18096 VDD.n1901 VDD.n1900 185
R18097 VDD.n1900 VDD.n1899 185
R18098 VDD.n597 VDD.n596 185
R18099 VDD.n598 VDD.n597 185
R18100 VDD.n1892 VDD.n1891 185
R18101 VDD.n1893 VDD.n1892 185
R18102 VDD.n1890 VDD.n607 185
R18103 VDD.n607 VDD.n604 185
R18104 VDD.n1889 VDD.n1888 185
R18105 VDD.n1888 VDD.n1887 185
R18106 VDD.n609 VDD.n608 185
R18107 VDD.n610 VDD.n609 185
R18108 VDD.n1880 VDD.n1879 185
R18109 VDD.n1881 VDD.n1880 185
R18110 VDD.n1878 VDD.n619 185
R18111 VDD.n619 VDD.n616 185
R18112 VDD.n1877 VDD.n1876 185
R18113 VDD.n1876 VDD.n1875 185
R18114 VDD.n621 VDD.n620 185
R18115 VDD.n622 VDD.n621 185
R18116 VDD.n1868 VDD.n1867 185
R18117 VDD.n1869 VDD.n1868 185
R18118 VDD.n1866 VDD.n631 185
R18119 VDD.n631 VDD.n628 185
R18120 VDD.n1865 VDD.n1864 185
R18121 VDD.n1864 VDD.n1863 185
R18122 VDD.n633 VDD.n632 185
R18123 VDD.n634 VDD.n633 185
R18124 VDD.n1856 VDD.n1855 185
R18125 VDD.n1857 VDD.n1856 185
R18126 VDD.n1854 VDD.n643 185
R18127 VDD.n643 VDD.n640 185
R18128 VDD.n1853 VDD.n1852 185
R18129 VDD.n1852 VDD.n1851 185
R18130 VDD.n645 VDD.n644 185
R18131 VDD.n646 VDD.n645 185
R18132 VDD.n1844 VDD.n1843 185
R18133 VDD.n1845 VDD.n1844 185
R18134 VDD.n1842 VDD.n654 185
R18135 VDD.n660 VDD.n654 185
R18136 VDD.n1841 VDD.n1840 185
R18137 VDD.n1840 VDD.n1839 185
R18138 VDD.n656 VDD.n655 185
R18139 VDD.n657 VDD.n656 185
R18140 VDD.n1832 VDD.n1831 185
R18141 VDD.n1833 VDD.n1832 185
R18142 VDD.n1830 VDD.n666 185
R18143 VDD.n672 VDD.n666 185
R18144 VDD.n1829 VDD.n1828 185
R18145 VDD.n1828 VDD.n1827 185
R18146 VDD.n668 VDD.n667 185
R18147 VDD.n669 VDD.n668 185
R18148 VDD.n1820 VDD.n1819 185
R18149 VDD.n1821 VDD.n1820 185
R18150 VDD.n1818 VDD.n679 185
R18151 VDD.n679 VDD.n676 185
R18152 VDD.n1817 VDD.n1816 185
R18153 VDD.n1816 VDD.n1815 185
R18154 VDD.n681 VDD.n680 185
R18155 VDD.n682 VDD.n681 185
R18156 VDD.n1808 VDD.n1807 185
R18157 VDD.n1809 VDD.n1808 185
R18158 VDD.n1806 VDD.n691 185
R18159 VDD.n691 VDD.n688 185
R18160 VDD.n1805 VDD.n1804 185
R18161 VDD.n1804 VDD.n1803 185
R18162 VDD.n693 VDD.n692 185
R18163 VDD.n694 VDD.n693 185
R18164 VDD.n2043 VDD.n432 185
R18165 VDD.n2117 VDD.n432 185
R18166 VDD.n2045 VDD.n2044 185
R18167 VDD.n2047 VDD.n2046 185
R18168 VDD.n2049 VDD.n2048 185
R18169 VDD.n2051 VDD.n2050 185
R18170 VDD.n2053 VDD.n2052 185
R18171 VDD.n2055 VDD.n2054 185
R18172 VDD.n2057 VDD.n2056 185
R18173 VDD.n2059 VDD.n2058 185
R18174 VDD.n2061 VDD.n2060 185
R18175 VDD.n2063 VDD.n2062 185
R18176 VDD.n2065 VDD.n2064 185
R18177 VDD.n2067 VDD.n2066 185
R18178 VDD.n2069 VDD.n2068 185
R18179 VDD.n2071 VDD.n2070 185
R18180 VDD.n2042 VDD.n2041 185
R18181 VDD.n2041 VDD.n424 185
R18182 VDD.n2040 VDD.n449 185
R18183 VDD.n2084 VDD.n449 185
R18184 VDD.n2039 VDD.n2038 185
R18185 VDD.n2038 VDD.n448 185
R18186 VDD.n2037 VDD.n456 185
R18187 VDD.n2078 VDD.n456 185
R18188 VDD.n2036 VDD.n2035 185
R18189 VDD.n2035 VDD.n454 185
R18190 VDD.n2034 VDD.n463 185
R18191 VDD.n2034 VDD.n2033 185
R18192 VDD.n787 VDD.n464 185
R18193 VDD.n465 VDD.n464 185
R18194 VDD.n788 VDD.n473 185
R18195 VDD.n2027 VDD.n473 185
R18196 VDD.n790 VDD.n789 185
R18197 VDD.n789 VDD.n471 185
R18198 VDD.n791 VDD.n480 185
R18199 VDD.n2019 VDD.n480 185
R18200 VDD.n793 VDD.n792 185
R18201 VDD.n792 VDD.n478 185
R18202 VDD.n794 VDD.n486 185
R18203 VDD.n2013 VDD.n486 185
R18204 VDD.n796 VDD.n795 185
R18205 VDD.n795 VDD.n484 185
R18206 VDD.n797 VDD.n492 185
R18207 VDD.n2007 VDD.n492 185
R18208 VDD.n799 VDD.n798 185
R18209 VDD.n798 VDD.n490 185
R18210 VDD.n800 VDD.n498 185
R18211 VDD.n2001 VDD.n498 185
R18212 VDD.n802 VDD.n801 185
R18213 VDD.n801 VDD.n496 185
R18214 VDD.n803 VDD.n504 185
R18215 VDD.n1995 VDD.n504 185
R18216 VDD.n805 VDD.n804 185
R18217 VDD.n804 VDD.n502 185
R18218 VDD.n806 VDD.n510 185
R18219 VDD.n1989 VDD.n510 185
R18220 VDD.n808 VDD.n807 185
R18221 VDD.n807 VDD.n508 185
R18222 VDD.n809 VDD.n516 185
R18223 VDD.n1983 VDD.n516 185
R18224 VDD.n811 VDD.n810 185
R18225 VDD.n810 VDD.n514 185
R18226 VDD.n812 VDD.n522 185
R18227 VDD.n1977 VDD.n522 185
R18228 VDD.n814 VDD.n813 185
R18229 VDD.n813 VDD.n520 185
R18230 VDD.n815 VDD.n528 185
R18231 VDD.n1971 VDD.n528 185
R18232 VDD.n817 VDD.n816 185
R18233 VDD.n816 VDD.n526 185
R18234 VDD.n818 VDD.n534 185
R18235 VDD.n1965 VDD.n534 185
R18236 VDD.n820 VDD.n819 185
R18237 VDD.n819 VDD.n532 185
R18238 VDD.n821 VDD.n540 185
R18239 VDD.n1959 VDD.n540 185
R18240 VDD.n823 VDD.n822 185
R18241 VDD.n822 VDD.n538 185
R18242 VDD.n824 VDD.n545 185
R18243 VDD.n1953 VDD.n545 185
R18244 VDD.n826 VDD.n825 185
R18245 VDD.n825 VDD.n552 185
R18246 VDD.n827 VDD.n551 185
R18247 VDD.n1947 VDD.n551 185
R18248 VDD.n829 VDD.n828 185
R18249 VDD.n828 VDD.n549 185
R18250 VDD.n830 VDD.n558 185
R18251 VDD.n1941 VDD.n558 185
R18252 VDD.n832 VDD.n831 185
R18253 VDD.n831 VDD.n556 185
R18254 VDD.n833 VDD.n564 185
R18255 VDD.n1935 VDD.n564 185
R18256 VDD.n835 VDD.n834 185
R18257 VDD.n834 VDD.n562 185
R18258 VDD.n836 VDD.n570 185
R18259 VDD.n1929 VDD.n570 185
R18260 VDD.n838 VDD.n837 185
R18261 VDD.n837 VDD.n568 185
R18262 VDD.n839 VDD.n576 185
R18263 VDD.n1923 VDD.n576 185
R18264 VDD.n841 VDD.n840 185
R18265 VDD.n840 VDD.n574 185
R18266 VDD.n842 VDD.n582 185
R18267 VDD.n1917 VDD.n582 185
R18268 VDD.n844 VDD.n843 185
R18269 VDD.n843 VDD.n580 185
R18270 VDD.n845 VDD.n588 185
R18271 VDD.n1911 VDD.n588 185
R18272 VDD.n847 VDD.n846 185
R18273 VDD.n846 VDD.n586 185
R18274 VDD.n848 VDD.n594 185
R18275 VDD.n1905 VDD.n594 185
R18276 VDD.n850 VDD.n849 185
R18277 VDD.n849 VDD.n592 185
R18278 VDD.n851 VDD.n600 185
R18279 VDD.n1899 VDD.n600 185
R18280 VDD.n853 VDD.n852 185
R18281 VDD.n852 VDD.n598 185
R18282 VDD.n854 VDD.n606 185
R18283 VDD.n1893 VDD.n606 185
R18284 VDD.n856 VDD.n855 185
R18285 VDD.n855 VDD.n604 185
R18286 VDD.n857 VDD.n612 185
R18287 VDD.n1887 VDD.n612 185
R18288 VDD.n859 VDD.n858 185
R18289 VDD.n858 VDD.n610 185
R18290 VDD.n860 VDD.n618 185
R18291 VDD.n1881 VDD.n618 185
R18292 VDD.n862 VDD.n861 185
R18293 VDD.n861 VDD.n616 185
R18294 VDD.n863 VDD.n624 185
R18295 VDD.n1875 VDD.n624 185
R18296 VDD.n865 VDD.n864 185
R18297 VDD.n864 VDD.n622 185
R18298 VDD.n866 VDD.n630 185
R18299 VDD.n1869 VDD.n630 185
R18300 VDD.n868 VDD.n867 185
R18301 VDD.n867 VDD.n628 185
R18302 VDD.n869 VDD.n636 185
R18303 VDD.n1863 VDD.n636 185
R18304 VDD.n871 VDD.n870 185
R18305 VDD.n870 VDD.n634 185
R18306 VDD.n872 VDD.n642 185
R18307 VDD.n1857 VDD.n642 185
R18308 VDD.n874 VDD.n873 185
R18309 VDD.n873 VDD.n640 185
R18310 VDD.n875 VDD.n648 185
R18311 VDD.n1851 VDD.n648 185
R18312 VDD.n877 VDD.n876 185
R18313 VDD.n876 VDD.n646 185
R18314 VDD.n878 VDD.n653 185
R18315 VDD.n1845 VDD.n653 185
R18316 VDD.n880 VDD.n879 185
R18317 VDD.n879 VDD.n660 185
R18318 VDD.n881 VDD.n659 185
R18319 VDD.n1839 VDD.n659 185
R18320 VDD.n883 VDD.n882 185
R18321 VDD.n882 VDD.n657 185
R18322 VDD.n884 VDD.n665 185
R18323 VDD.n1833 VDD.n665 185
R18324 VDD.n886 VDD.n885 185
R18325 VDD.n885 VDD.n672 185
R18326 VDD.n887 VDD.n671 185
R18327 VDD.n1827 VDD.n671 185
R18328 VDD.n889 VDD.n888 185
R18329 VDD.n888 VDD.n669 185
R18330 VDD.n890 VDD.n678 185
R18331 VDD.n1821 VDD.n678 185
R18332 VDD.n892 VDD.n891 185
R18333 VDD.n891 VDD.n676 185
R18334 VDD.n893 VDD.n684 185
R18335 VDD.n1815 VDD.n684 185
R18336 VDD.n895 VDD.n894 185
R18337 VDD.n894 VDD.n682 185
R18338 VDD.n896 VDD.n690 185
R18339 VDD.n1809 VDD.n690 185
R18340 VDD.n898 VDD.n897 185
R18341 VDD.n897 VDD.n688 185
R18342 VDD.n899 VDD.n696 185
R18343 VDD.n1803 VDD.n696 185
R18344 VDD.n901 VDD.n900 185
R18345 VDD.n900 VDD.n694 185
R18346 VDD.n770 VDD.n769 185
R18347 VDD.n772 VDD.n771 185
R18348 VDD.n774 VDD.n773 185
R18349 VDD.n776 VDD.n775 185
R18350 VDD.n778 VDD.n777 185
R18351 VDD.n780 VDD.n779 185
R18352 VDD.n782 VDD.n781 185
R18353 VDD.n915 VDD.n783 185
R18354 VDD.n914 VDD.n913 185
R18355 VDD.n912 VDD.n911 185
R18356 VDD.n910 VDD.n909 185
R18357 VDD.n908 VDD.n907 185
R18358 VDD.n906 VDD.n905 185
R18359 VDD.n904 VDD.n903 185
R18360 VDD.n902 VDD.n713 185
R18361 VDD.n1796 VDD.n713 185
R18362 VDD.n785 VDD.t65 173.75
R18363 VDD.n461 VDD.t23 173.75
R18364 VDD.n1648 VDD.t12 173.75
R18365 VDD.n444 VDD.t39 173.75
R18366 VDD.n2133 VDD.t89 173.75
R18367 VDD.n177 VDD.t46 173.75
R18368 VDD.n2282 VDD.t62 173.75
R18369 VDD.n155 VDD.t72 173.75
R18370 VDD.n3397 VDD.n3396 171.744
R18371 VDD.n3396 VDD.n3386 171.744
R18372 VDD.n3389 VDD.n3386 171.744
R18373 VDD.n3377 VDD.n3376 171.744
R18374 VDD.n3376 VDD.n3366 171.744
R18375 VDD.n3369 VDD.n3366 171.744
R18376 VDD.n3357 VDD.n3356 171.744
R18377 VDD.n3356 VDD.n3346 171.744
R18378 VDD.n3349 VDD.n3346 171.744
R18379 VDD.n3337 VDD.n3336 171.744
R18380 VDD.n3336 VDD.n3326 171.744
R18381 VDD.n3329 VDD.n3326 171.744
R18382 VDD.n3318 VDD.n3317 171.744
R18383 VDD.n3317 VDD.n3307 171.744
R18384 VDD.n3310 VDD.n3307 171.744
R18385 VDD.n1433 VDD.n1432 171.744
R18386 VDD.n1432 VDD.n1422 171.744
R18387 VDD.n1425 VDD.n1422 171.744
R18388 VDD.n1413 VDD.n1412 171.744
R18389 VDD.n1412 VDD.n1402 171.744
R18390 VDD.n1405 VDD.n1402 171.744
R18391 VDD.n1393 VDD.n1392 171.744
R18392 VDD.n1392 VDD.n1382 171.744
R18393 VDD.n1385 VDD.n1382 171.744
R18394 VDD.n1373 VDD.n1372 171.744
R18395 VDD.n1372 VDD.n1362 171.744
R18396 VDD.n1365 VDD.n1362 171.744
R18397 VDD.n1354 VDD.n1353 171.744
R18398 VDD.n1353 VDD.n1343 171.744
R18399 VDD.n1346 VDD.n1343 171.744
R18400 VDD.t94 VDD.t109 163.022
R18401 VDD.t109 VDD.t107 163.022
R18402 VDD.t107 VDD.t128 163.022
R18403 VDD.t130 VDD.t124 163.022
R18404 VDD.t124 VDD.t111 163.022
R18405 VDD.t111 VDD.t135 163.022
R18406 VDD.n2918 VDD.n59 146.341
R18407 VDD.n2918 VDD.n55 146.341
R18408 VDD.n2924 VDD.n55 146.341
R18409 VDD.n2924 VDD.n47 146.341
R18410 VDD.n2934 VDD.n47 146.341
R18411 VDD.n2934 VDD.n43 146.341
R18412 VDD.n2940 VDD.n43 146.341
R18413 VDD.n2940 VDD.n35 146.341
R18414 VDD.n2950 VDD.n35 146.341
R18415 VDD.n2950 VDD.n31 146.341
R18416 VDD.n2956 VDD.n31 146.341
R18417 VDD.n2956 VDD.n20 146.341
R18418 VDD.n3301 VDD.n20 146.341
R18419 VDD.n3301 VDD.n21 146.341
R18420 VDD.n3294 VDD.n21 146.341
R18421 VDD.n3294 VDD.n2968 146.341
R18422 VDD.n3290 VDD.n2968 146.341
R18423 VDD.n3290 VDD.n2973 146.341
R18424 VDD.n3286 VDD.n2973 146.341
R18425 VDD.n3286 VDD.n2978 146.341
R18426 VDD.n3282 VDD.n2978 146.341
R18427 VDD.n3282 VDD.n2984 146.341
R18428 VDD.n3278 VDD.n2984 146.341
R18429 VDD.n3278 VDD.n2989 146.341
R18430 VDD.n3274 VDD.n2989 146.341
R18431 VDD.n3274 VDD.n2995 146.341
R18432 VDD.n3083 VDD.n3082 146.341
R18433 VDD.n3087 VDD.n3086 146.341
R18434 VDD.n3093 VDD.n3092 146.341
R18435 VDD.n3097 VDD.n3096 146.341
R18436 VDD.n3103 VDD.n3102 146.341
R18437 VDD.n3107 VDD.n3106 146.341
R18438 VDD.n3113 VDD.n3112 146.341
R18439 VDD.n3117 VDD.n3116 146.341
R18440 VDD.n3123 VDD.n3122 146.341
R18441 VDD.n3127 VDD.n3126 146.341
R18442 VDD.n3133 VDD.n3132 146.341
R18443 VDD.n3137 VDD.n3136 146.341
R18444 VDD.n3143 VDD.n3142 146.341
R18445 VDD.n3147 VDD.n3146 146.341
R18446 VDD.n3153 VDD.n3152 146.341
R18447 VDD.n3157 VDD.n3156 146.341
R18448 VDD.n3163 VDD.n3162 146.341
R18449 VDD.n3167 VDD.n3166 146.341
R18450 VDD.n3173 VDD.n3172 146.341
R18451 VDD.n3177 VDD.n3176 146.341
R18452 VDD.n3180 VDD.n3179 146.341
R18453 VDD.n3187 VDD.n3186 146.341
R18454 VDD.n3190 VDD.n3189 146.341
R18455 VDD.n3197 VDD.n3196 146.341
R18456 VDD.n3200 VDD.n3199 146.341
R18457 VDD.n3207 VDD.n3206 146.341
R18458 VDD.n3211 VDD.n3210 146.341
R18459 VDD.n3218 VDD.n3217 146.341
R18460 VDD.n3221 VDD.n3220 146.341
R18461 VDD.n3228 VDD.n3227 146.341
R18462 VDD.n3231 VDD.n3230 146.341
R18463 VDD.n3238 VDD.n3237 146.341
R18464 VDD.n3240 VDD.n3031 146.341
R18465 VDD.n2916 VDD.n61 146.341
R18466 VDD.n2916 VDD.n53 146.341
R18467 VDD.n2926 VDD.n53 146.341
R18468 VDD.n2926 VDD.n49 146.341
R18469 VDD.n2932 VDD.n49 146.341
R18470 VDD.n2932 VDD.n41 146.341
R18471 VDD.n2942 VDD.n41 146.341
R18472 VDD.n2942 VDD.n37 146.341
R18473 VDD.n2948 VDD.n37 146.341
R18474 VDD.n2948 VDD.n29 146.341
R18475 VDD.n2958 VDD.n29 146.341
R18476 VDD.n2958 VDD.n24 146.341
R18477 VDD.n3300 VDD.n24 146.341
R18478 VDD.n3300 VDD.n25 146.341
R18479 VDD.n3296 VDD.n25 146.341
R18480 VDD.n3296 VDD.n2966 146.341
R18481 VDD.n2974 VDD.n2966 146.341
R18482 VDD.n2975 VDD.n2974 146.341
R18483 VDD.n2976 VDD.n2975 146.341
R18484 VDD.n3255 VDD.n2976 146.341
R18485 VDD.n3255 VDD.n2985 146.341
R18486 VDD.n2986 VDD.n2985 146.341
R18487 VDD.n2987 VDD.n2986 146.341
R18488 VDD.n3262 VDD.n2987 146.341
R18489 VDD.n3262 VDD.n2996 146.341
R18490 VDD.n2997 VDD.n2996 146.341
R18491 VDD.n101 VDD.n100 146.341
R18492 VDD.n2902 VDD.n100 146.341
R18493 VDD.n2900 VDD.n2899 146.341
R18494 VDD.n2896 VDD.n2895 146.341
R18495 VDD.n2892 VDD.n2891 146.341
R18496 VDD.n2888 VDD.n2887 146.341
R18497 VDD.n2884 VDD.n2883 146.341
R18498 VDD.n2880 VDD.n2879 146.341
R18499 VDD.n2876 VDD.n2875 146.341
R18500 VDD.n2872 VDD.n2871 146.341
R18501 VDD.n2868 VDD.n2867 146.341
R18502 VDD.n2864 VDD.n2863 146.341
R18503 VDD.n2860 VDD.n2859 146.341
R18504 VDD.n2851 VDD.n2850 146.341
R18505 VDD.n2848 VDD.n2847 146.341
R18506 VDD.n2844 VDD.n2843 146.341
R18507 VDD.n2840 VDD.n2839 146.341
R18508 VDD.n2836 VDD.n2835 146.341
R18509 VDD.n2832 VDD.n2831 146.341
R18510 VDD.n2828 VDD.n2827 146.341
R18511 VDD.n2821 VDD.n2820 146.341
R18512 VDD.n2818 VDD.n2817 146.341
R18513 VDD.n2814 VDD.n2813 146.341
R18514 VDD.n2810 VDD.n2809 146.341
R18515 VDD.n2806 VDD.n2805 146.341
R18516 VDD.n2802 VDD.n2801 146.341
R18517 VDD.n2798 VDD.n2797 146.341
R18518 VDD.n2794 VDD.n2793 146.341
R18519 VDD.n2790 VDD.n2789 146.341
R18520 VDD.n2786 VDD.n2785 146.341
R18521 VDD.n2782 VDD.n2781 146.341
R18522 VDD.n2778 VDD.n2777 146.341
R18523 VDD.n2774 VDD.n2773 146.341
R18524 VDD.n2910 VDD.n67 146.341
R18525 VDD.n1548 VDD.n1494 146.341
R18526 VDD.n1546 VDD.n1545 146.341
R18527 VDD.n1543 VDD.n1498 146.341
R18528 VDD.n1539 VDD.n1538 146.341
R18529 VDD.n1536 VDD.n1506 146.341
R18530 VDD.n1531 VDD.n1513 146.341
R18531 VDD.n1529 VDD.n1528 146.341
R18532 VDD.n1526 VDD.n1519 146.341
R18533 VDD.n1643 VDD.n720 146.341
R18534 VDD.n1641 VDD.n1640 146.341
R18535 VDD.n1638 VDD.n723 146.341
R18536 VDD.n1634 VDD.n1633 146.341
R18537 VDD.n1631 VDD.n727 146.341
R18538 VDD.n1625 VDD.n1624 146.341
R18539 VDD.n1622 VDD.n735 146.341
R18540 VDD.n1618 VDD.n1617 146.341
R18541 VDD.n1615 VDD.n741 146.341
R18542 VDD.n1611 VDD.n1610 146.341
R18543 VDD.n1608 VDD.n748 146.341
R18544 VDD.n759 VDD.n756 146.341
R18545 VDD.n1600 VDD.n1599 146.341
R18546 VDD.n1597 VDD.n761 146.341
R18547 VDD.n1593 VDD.n1592 146.341
R18548 VDD.n1590 VDD.n767 146.341
R18549 VDD.n921 VDD.n920 146.341
R18550 VDD.n924 VDD.n923 146.341
R18551 VDD.n931 VDD.n930 146.341
R18552 VDD.n936 VDD.n933 146.341
R18553 VDD.n939 VDD.n938 146.341
R18554 VDD.n944 VDD.n941 146.341
R18555 VDD.n947 VDD.n946 146.341
R18556 VDD.n952 VDD.n949 146.341
R18557 VDD.n1560 VDD.n954 146.341
R18558 VDD.n1287 VDD.n1031 146.341
R18559 VDD.n1297 VDD.n1031 146.341
R18560 VDD.n1297 VDD.n1027 146.341
R18561 VDD.n1303 VDD.n1027 146.341
R18562 VDD.n1303 VDD.n1020 146.341
R18563 VDD.n1313 VDD.n1020 146.341
R18564 VDD.n1313 VDD.n1016 146.341
R18565 VDD.n1319 VDD.n1016 146.341
R18566 VDD.n1319 VDD.n1008 146.341
R18567 VDD.n1329 VDD.n1008 146.341
R18568 VDD.n1329 VDD.n1004 146.341
R18569 VDD.n1335 VDD.n1004 146.341
R18570 VDD.n1335 VDD.n997 146.341
R18571 VDD.n1445 VDD.n997 146.341
R18572 VDD.n1445 VDD.n993 146.341
R18573 VDD.n1451 VDD.n993 146.341
R18574 VDD.n1451 VDD.n985 146.341
R18575 VDD.n1461 VDD.n985 146.341
R18576 VDD.n1461 VDD.n981 146.341
R18577 VDD.n1467 VDD.n981 146.341
R18578 VDD.n1467 VDD.n973 146.341
R18579 VDD.n1477 VDD.n973 146.341
R18580 VDD.n1477 VDD.n968 146.341
R18581 VDD.n1486 VDD.n968 146.341
R18582 VDD.n1486 VDD.n958 146.341
R18583 VDD.n1557 VDD.n958 146.341
R18584 VDD.n1122 VDD.n1118 146.341
R18585 VDD.n1128 VDD.n1118 146.341
R18586 VDD.n1132 VDD.n1130 146.341
R18587 VDD.n1140 VDD.n1114 146.341
R18588 VDD.n1143 VDD.n1142 146.341
R18589 VDD.n1145 VDD.n1109 146.341
R18590 VDD.n1152 VDD.n1105 146.341
R18591 VDD.n1156 VDD.n1154 146.341
R18592 VDD.n1162 VDD.n1101 146.341
R18593 VDD.n1166 VDD.n1164 146.341
R18594 VDD.n1174 VDD.n1097 146.341
R18595 VDD.n1177 VDD.n1176 146.341
R18596 VDD.n1179 VDD.n1092 146.341
R18597 VDD.n1186 VDD.n1088 146.341
R18598 VDD.n1190 VDD.n1188 146.341
R18599 VDD.n1196 VDD.n1084 146.341
R18600 VDD.n1200 VDD.n1198 146.341
R18601 VDD.n1208 VDD.n1080 146.341
R18602 VDD.n1211 VDD.n1210 146.341
R18603 VDD.n1213 VDD.n1075 146.341
R18604 VDD.n1220 VDD.n1071 146.341
R18605 VDD.n1224 VDD.n1222 146.341
R18606 VDD.n1230 VDD.n1067 146.341
R18607 VDD.n1234 VDD.n1232 146.341
R18608 VDD.n1241 VDD.n1063 146.341
R18609 VDD.n1245 VDD.n1243 146.341
R18610 VDD.n1251 VDD.n1057 146.341
R18611 VDD.n1255 VDD.n1253 146.341
R18612 VDD.n1261 VDD.n1053 146.341
R18613 VDD.n1265 VDD.n1263 146.341
R18614 VDD.n1271 VDD.n1049 146.341
R18615 VDD.n1276 VDD.n1273 146.341
R18616 VDD.n1274 VDD.n1046 146.341
R18617 VDD.n1041 VDD.n1039 146.341
R18618 VDD.n1289 VDD.n1034 146.341
R18619 VDD.n1295 VDD.n1034 146.341
R18620 VDD.n1295 VDD.n1026 146.341
R18621 VDD.n1305 VDD.n1026 146.341
R18622 VDD.n1305 VDD.n1022 146.341
R18623 VDD.n1311 VDD.n1022 146.341
R18624 VDD.n1311 VDD.n1014 146.341
R18625 VDD.n1321 VDD.n1014 146.341
R18626 VDD.n1321 VDD.n1010 146.341
R18627 VDD.n1327 VDD.n1010 146.341
R18628 VDD.n1327 VDD.n1002 146.341
R18629 VDD.n1337 VDD.n1002 146.341
R18630 VDD.n1337 VDD.n998 146.341
R18631 VDD.n1443 VDD.n998 146.341
R18632 VDD.n1443 VDD.n991 146.341
R18633 VDD.n1453 VDD.n991 146.341
R18634 VDD.n1453 VDD.n987 146.341
R18635 VDD.n1459 VDD.n987 146.341
R18636 VDD.n1459 VDD.n979 146.341
R18637 VDD.n1469 VDD.n979 146.341
R18638 VDD.n1469 VDD.n975 146.341
R18639 VDD.n1475 VDD.n975 146.341
R18640 VDD.n1475 VDD.n966 146.341
R18641 VDD.n1488 VDD.n966 146.341
R18642 VDD.n1488 VDD.n961 146.341
R18643 VDD.n1555 VDD.n961 146.341
R18644 VDD.n785 VDD.n784 121.406
R18645 VDD.n461 VDD.n460 121.406
R18646 VDD.n1648 VDD.n1647 121.406
R18647 VDD.n444 VDD.n443 121.406
R18648 VDD.n2133 VDD.n2132 121.406
R18649 VDD.n177 VDD.n176 121.406
R18650 VDD.n2282 VDD.n2281 121.406
R18651 VDD.n155 VDD.n154 121.406
R18652 VDD.n2727 VDD.n2726 99.5127
R18653 VDD.n2724 VDD.n169 99.5127
R18654 VDD.n2720 VDD.n2719 99.5127
R18655 VDD.n2717 VDD.n172 99.5127
R18656 VDD.n2712 VDD.n2711 99.5127
R18657 VDD.n2709 VDD.n175 99.5127
R18658 VDD.n2704 VDD.n2703 99.5127
R18659 VDD.n2400 VDD.n419 99.5127
R18660 VDD.n2396 VDD.n419 99.5127
R18661 VDD.n2396 VDD.n413 99.5127
R18662 VDD.n2393 VDD.n413 99.5127
R18663 VDD.n2393 VDD.n407 99.5127
R18664 VDD.n2390 VDD.n407 99.5127
R18665 VDD.n2390 VDD.n401 99.5127
R18666 VDD.n2387 VDD.n401 99.5127
R18667 VDD.n2387 VDD.n394 99.5127
R18668 VDD.n2384 VDD.n394 99.5127
R18669 VDD.n2384 VDD.n387 99.5127
R18670 VDD.n2381 VDD.n387 99.5127
R18671 VDD.n2381 VDD.n382 99.5127
R18672 VDD.n2378 VDD.n382 99.5127
R18673 VDD.n2378 VDD.n377 99.5127
R18674 VDD.n2375 VDD.n377 99.5127
R18675 VDD.n2375 VDD.n371 99.5127
R18676 VDD.n2372 VDD.n371 99.5127
R18677 VDD.n2372 VDD.n365 99.5127
R18678 VDD.n2369 VDD.n365 99.5127
R18679 VDD.n2369 VDD.n359 99.5127
R18680 VDD.n2366 VDD.n359 99.5127
R18681 VDD.n2366 VDD.n353 99.5127
R18682 VDD.n2363 VDD.n353 99.5127
R18683 VDD.n2363 VDD.n347 99.5127
R18684 VDD.n2360 VDD.n347 99.5127
R18685 VDD.n2360 VDD.n341 99.5127
R18686 VDD.n2357 VDD.n341 99.5127
R18687 VDD.n2357 VDD.n334 99.5127
R18688 VDD.n2354 VDD.n334 99.5127
R18689 VDD.n2354 VDD.n328 99.5127
R18690 VDD.n2351 VDD.n328 99.5127
R18691 VDD.n2351 VDD.n323 99.5127
R18692 VDD.n2348 VDD.n323 99.5127
R18693 VDD.n2348 VDD.n317 99.5127
R18694 VDD.n2345 VDD.n317 99.5127
R18695 VDD.n2345 VDD.n311 99.5127
R18696 VDD.n2342 VDD.n311 99.5127
R18697 VDD.n2342 VDD.n305 99.5127
R18698 VDD.n2339 VDD.n305 99.5127
R18699 VDD.n2339 VDD.n299 99.5127
R18700 VDD.n2336 VDD.n299 99.5127
R18701 VDD.n2336 VDD.n293 99.5127
R18702 VDD.n2333 VDD.n293 99.5127
R18703 VDD.n2333 VDD.n287 99.5127
R18704 VDD.n2330 VDD.n287 99.5127
R18705 VDD.n2330 VDD.n280 99.5127
R18706 VDD.n2327 VDD.n280 99.5127
R18707 VDD.n2327 VDD.n273 99.5127
R18708 VDD.n2324 VDD.n273 99.5127
R18709 VDD.n2324 VDD.n268 99.5127
R18710 VDD.n2321 VDD.n268 99.5127
R18711 VDD.n2321 VDD.n263 99.5127
R18712 VDD.n2318 VDD.n263 99.5127
R18713 VDD.n2318 VDD.n257 99.5127
R18714 VDD.n2315 VDD.n257 99.5127
R18715 VDD.n2315 VDD.n251 99.5127
R18716 VDD.n2312 VDD.n251 99.5127
R18717 VDD.n2312 VDD.n245 99.5127
R18718 VDD.n2309 VDD.n245 99.5127
R18719 VDD.n2309 VDD.n239 99.5127
R18720 VDD.n2306 VDD.n239 99.5127
R18721 VDD.n2306 VDD.n233 99.5127
R18722 VDD.n2303 VDD.n233 99.5127
R18723 VDD.n2303 VDD.n227 99.5127
R18724 VDD.n2300 VDD.n227 99.5127
R18725 VDD.n2300 VDD.n221 99.5127
R18726 VDD.n2297 VDD.n221 99.5127
R18727 VDD.n2297 VDD.n215 99.5127
R18728 VDD.n2294 VDD.n215 99.5127
R18729 VDD.n2294 VDD.n209 99.5127
R18730 VDD.n2291 VDD.n209 99.5127
R18731 VDD.n2291 VDD.n203 99.5127
R18732 VDD.n2288 VDD.n203 99.5127
R18733 VDD.n2288 VDD.n197 99.5127
R18734 VDD.n2285 VDD.n197 99.5127
R18735 VDD.n2285 VDD.n190 99.5127
R18736 VDD.n190 VDD.n182 99.5127
R18737 VDD.n2695 VDD.n182 99.5127
R18738 VDD.n2696 VDD.n2695 99.5127
R18739 VDD.n2696 VDD.n162 99.5127
R18740 VDD.n180 VDD.n162 99.5127
R18741 VDD.n2280 VDD.n2279 99.5127
R18742 VDD.n2424 VDD.n2279 99.5127
R18743 VDD.n2422 VDD.n2421 99.5127
R18744 VDD.n2418 VDD.n2417 99.5127
R18745 VDD.n2414 VDD.n2413 99.5127
R18746 VDD.n2410 VDD.n2409 99.5127
R18747 VDD.n2405 VDD.n2404 99.5127
R18748 VDD.n2439 VDD.n417 99.5127
R18749 VDD.n2439 VDD.n415 99.5127
R18750 VDD.n2443 VDD.n415 99.5127
R18751 VDD.n2443 VDD.n405 99.5127
R18752 VDD.n2451 VDD.n405 99.5127
R18753 VDD.n2451 VDD.n403 99.5127
R18754 VDD.n2455 VDD.n403 99.5127
R18755 VDD.n2455 VDD.n392 99.5127
R18756 VDD.n2463 VDD.n392 99.5127
R18757 VDD.n2463 VDD.n390 99.5127
R18758 VDD.n2467 VDD.n390 99.5127
R18759 VDD.n2467 VDD.n381 99.5127
R18760 VDD.n2475 VDD.n381 99.5127
R18761 VDD.n2475 VDD.n379 99.5127
R18762 VDD.n2479 VDD.n379 99.5127
R18763 VDD.n2479 VDD.n369 99.5127
R18764 VDD.n2487 VDD.n369 99.5127
R18765 VDD.n2487 VDD.n367 99.5127
R18766 VDD.n2491 VDD.n367 99.5127
R18767 VDD.n2491 VDD.n357 99.5127
R18768 VDD.n2499 VDD.n357 99.5127
R18769 VDD.n2499 VDD.n355 99.5127
R18770 VDD.n2503 VDD.n355 99.5127
R18771 VDD.n2503 VDD.n345 99.5127
R18772 VDD.n2511 VDD.n345 99.5127
R18773 VDD.n2511 VDD.n343 99.5127
R18774 VDD.n2515 VDD.n343 99.5127
R18775 VDD.n2515 VDD.n332 99.5127
R18776 VDD.n2523 VDD.n332 99.5127
R18777 VDD.n2523 VDD.n330 99.5127
R18778 VDD.n2527 VDD.n330 99.5127
R18779 VDD.n2527 VDD.n321 99.5127
R18780 VDD.n2535 VDD.n321 99.5127
R18781 VDD.n2535 VDD.n319 99.5127
R18782 VDD.n2539 VDD.n319 99.5127
R18783 VDD.n2539 VDD.n309 99.5127
R18784 VDD.n2547 VDD.n309 99.5127
R18785 VDD.n2547 VDD.n307 99.5127
R18786 VDD.n2551 VDD.n307 99.5127
R18787 VDD.n2551 VDD.n297 99.5127
R18788 VDD.n2559 VDD.n297 99.5127
R18789 VDD.n2559 VDD.n295 99.5127
R18790 VDD.n2563 VDD.n295 99.5127
R18791 VDD.n2563 VDD.n285 99.5127
R18792 VDD.n2571 VDD.n285 99.5127
R18793 VDD.n2571 VDD.n283 99.5127
R18794 VDD.n2575 VDD.n283 99.5127
R18795 VDD.n2575 VDD.n272 99.5127
R18796 VDD.n2583 VDD.n272 99.5127
R18797 VDD.n2583 VDD.n270 99.5127
R18798 VDD.n2587 VDD.n270 99.5127
R18799 VDD.n2587 VDD.n261 99.5127
R18800 VDD.n2595 VDD.n261 99.5127
R18801 VDD.n2595 VDD.n259 99.5127
R18802 VDD.n2599 VDD.n259 99.5127
R18803 VDD.n2599 VDD.n249 99.5127
R18804 VDD.n2607 VDD.n249 99.5127
R18805 VDD.n2607 VDD.n247 99.5127
R18806 VDD.n2611 VDD.n247 99.5127
R18807 VDD.n2611 VDD.n237 99.5127
R18808 VDD.n2619 VDD.n237 99.5127
R18809 VDD.n2619 VDD.n235 99.5127
R18810 VDD.n2623 VDD.n235 99.5127
R18811 VDD.n2623 VDD.n225 99.5127
R18812 VDD.n2631 VDD.n225 99.5127
R18813 VDD.n2631 VDD.n223 99.5127
R18814 VDD.n2635 VDD.n223 99.5127
R18815 VDD.n2635 VDD.n213 99.5127
R18816 VDD.n2643 VDD.n213 99.5127
R18817 VDD.n2643 VDD.n211 99.5127
R18818 VDD.n2647 VDD.n211 99.5127
R18819 VDD.n2647 VDD.n201 99.5127
R18820 VDD.n2655 VDD.n201 99.5127
R18821 VDD.n2655 VDD.n199 99.5127
R18822 VDD.n2659 VDD.n199 99.5127
R18823 VDD.n2659 VDD.n188 99.5127
R18824 VDD.n2689 VDD.n188 99.5127
R18825 VDD.n2689 VDD.n186 99.5127
R18826 VDD.n2693 VDD.n186 99.5127
R18827 VDD.n2693 VDD.n165 99.5127
R18828 VDD.n2731 VDD.n165 99.5127
R18829 VDD.n2731 VDD.n166 99.5127
R18830 VDD.n2116 VDD.n441 99.5127
R18831 VDD.n2112 VDD.n2111 99.5127
R18832 VDD.n2108 VDD.n2107 99.5127
R18833 VDD.n2104 VDD.n2103 99.5127
R18834 VDD.n2100 VDD.n2099 99.5127
R18835 VDD.n2096 VDD.n2095 99.5127
R18836 VDD.n2091 VDD.n2090 99.5127
R18837 VDD.n1769 VDD.n695 99.5127
R18838 VDD.n1765 VDD.n695 99.5127
R18839 VDD.n1765 VDD.n689 99.5127
R18840 VDD.n1762 VDD.n689 99.5127
R18841 VDD.n1762 VDD.n683 99.5127
R18842 VDD.n1759 VDD.n683 99.5127
R18843 VDD.n1759 VDD.n677 99.5127
R18844 VDD.n1756 VDD.n677 99.5127
R18845 VDD.n1756 VDD.n670 99.5127
R18846 VDD.n1753 VDD.n670 99.5127
R18847 VDD.n1753 VDD.n664 99.5127
R18848 VDD.n1750 VDD.n664 99.5127
R18849 VDD.n1750 VDD.n658 99.5127
R18850 VDD.n1747 VDD.n658 99.5127
R18851 VDD.n1747 VDD.n652 99.5127
R18852 VDD.n1744 VDD.n652 99.5127
R18853 VDD.n1744 VDD.n647 99.5127
R18854 VDD.n1741 VDD.n647 99.5127
R18855 VDD.n1741 VDD.n641 99.5127
R18856 VDD.n1738 VDD.n641 99.5127
R18857 VDD.n1738 VDD.n635 99.5127
R18858 VDD.n1735 VDD.n635 99.5127
R18859 VDD.n1735 VDD.n629 99.5127
R18860 VDD.n1732 VDD.n629 99.5127
R18861 VDD.n1732 VDD.n623 99.5127
R18862 VDD.n1729 VDD.n623 99.5127
R18863 VDD.n1729 VDD.n617 99.5127
R18864 VDD.n1726 VDD.n617 99.5127
R18865 VDD.n1726 VDD.n611 99.5127
R18866 VDD.n1723 VDD.n611 99.5127
R18867 VDD.n1723 VDD.n605 99.5127
R18868 VDD.n1720 VDD.n605 99.5127
R18869 VDD.n1720 VDD.n599 99.5127
R18870 VDD.n1717 VDD.n599 99.5127
R18871 VDD.n1717 VDD.n593 99.5127
R18872 VDD.n1714 VDD.n593 99.5127
R18873 VDD.n1714 VDD.n587 99.5127
R18874 VDD.n1711 VDD.n587 99.5127
R18875 VDD.n1711 VDD.n581 99.5127
R18876 VDD.n1708 VDD.n581 99.5127
R18877 VDD.n1708 VDD.n575 99.5127
R18878 VDD.n1705 VDD.n575 99.5127
R18879 VDD.n1705 VDD.n569 99.5127
R18880 VDD.n1702 VDD.n569 99.5127
R18881 VDD.n1702 VDD.n563 99.5127
R18882 VDD.n1699 VDD.n563 99.5127
R18883 VDD.n1699 VDD.n557 99.5127
R18884 VDD.n1696 VDD.n557 99.5127
R18885 VDD.n1696 VDD.n550 99.5127
R18886 VDD.n1693 VDD.n550 99.5127
R18887 VDD.n1693 VDD.n544 99.5127
R18888 VDD.n1690 VDD.n544 99.5127
R18889 VDD.n1690 VDD.n539 99.5127
R18890 VDD.n1687 VDD.n539 99.5127
R18891 VDD.n1687 VDD.n533 99.5127
R18892 VDD.n1684 VDD.n533 99.5127
R18893 VDD.n1684 VDD.n527 99.5127
R18894 VDD.n1681 VDD.n527 99.5127
R18895 VDD.n1681 VDD.n521 99.5127
R18896 VDD.n1678 VDD.n521 99.5127
R18897 VDD.n1678 VDD.n515 99.5127
R18898 VDD.n1675 VDD.n515 99.5127
R18899 VDD.n1675 VDD.n509 99.5127
R18900 VDD.n1672 VDD.n509 99.5127
R18901 VDD.n1672 VDD.n503 99.5127
R18902 VDD.n1669 VDD.n503 99.5127
R18903 VDD.n1669 VDD.n497 99.5127
R18904 VDD.n1666 VDD.n497 99.5127
R18905 VDD.n1666 VDD.n491 99.5127
R18906 VDD.n1663 VDD.n491 99.5127
R18907 VDD.n1663 VDD.n485 99.5127
R18908 VDD.n1660 VDD.n485 99.5127
R18909 VDD.n1660 VDD.n479 99.5127
R18910 VDD.n1657 VDD.n479 99.5127
R18911 VDD.n1657 VDD.n472 99.5127
R18912 VDD.n1654 VDD.n472 99.5127
R18913 VDD.n1654 VDD.n466 99.5127
R18914 VDD.n1651 VDD.n466 99.5127
R18915 VDD.n1651 VDD.n455 99.5127
R18916 VDD.n455 VDD.n446 99.5127
R18917 VDD.n2085 VDD.n446 99.5127
R18918 VDD.n2086 VDD.n2085 99.5127
R18919 VDD.n1795 VDD.n699 99.5127
R18920 VDD.n1795 VDD.n714 99.5127
R18921 VDD.n1791 VDD.n1790 99.5127
R18922 VDD.n1787 VDD.n1786 99.5127
R18923 VDD.n1783 VDD.n1782 99.5127
R18924 VDD.n1779 VDD.n1778 99.5127
R18925 VDD.n1774 VDD.n1773 99.5127
R18926 VDD.n1802 VDD.n697 99.5127
R18927 VDD.n1802 VDD.n687 99.5127
R18928 VDD.n1810 VDD.n687 99.5127
R18929 VDD.n1810 VDD.n685 99.5127
R18930 VDD.n1814 VDD.n685 99.5127
R18931 VDD.n1814 VDD.n675 99.5127
R18932 VDD.n1822 VDD.n675 99.5127
R18933 VDD.n1822 VDD.n673 99.5127
R18934 VDD.n1826 VDD.n673 99.5127
R18935 VDD.n1826 VDD.n663 99.5127
R18936 VDD.n1834 VDD.n663 99.5127
R18937 VDD.n1834 VDD.n661 99.5127
R18938 VDD.n1838 VDD.n661 99.5127
R18939 VDD.n1838 VDD.n651 99.5127
R18940 VDD.n1846 VDD.n651 99.5127
R18941 VDD.n1846 VDD.n649 99.5127
R18942 VDD.n1850 VDD.n649 99.5127
R18943 VDD.n1850 VDD.n639 99.5127
R18944 VDD.n1858 VDD.n639 99.5127
R18945 VDD.n1858 VDD.n637 99.5127
R18946 VDD.n1862 VDD.n637 99.5127
R18947 VDD.n1862 VDD.n627 99.5127
R18948 VDD.n1870 VDD.n627 99.5127
R18949 VDD.n1870 VDD.n625 99.5127
R18950 VDD.n1874 VDD.n625 99.5127
R18951 VDD.n1874 VDD.n615 99.5127
R18952 VDD.n1882 VDD.n615 99.5127
R18953 VDD.n1882 VDD.n613 99.5127
R18954 VDD.n1886 VDD.n613 99.5127
R18955 VDD.n1886 VDD.n603 99.5127
R18956 VDD.n1894 VDD.n603 99.5127
R18957 VDD.n1894 VDD.n601 99.5127
R18958 VDD.n1898 VDD.n601 99.5127
R18959 VDD.n1898 VDD.n591 99.5127
R18960 VDD.n1906 VDD.n591 99.5127
R18961 VDD.n1906 VDD.n589 99.5127
R18962 VDD.n1910 VDD.n589 99.5127
R18963 VDD.n1910 VDD.n579 99.5127
R18964 VDD.n1918 VDD.n579 99.5127
R18965 VDD.n1918 VDD.n577 99.5127
R18966 VDD.n1922 VDD.n577 99.5127
R18967 VDD.n1922 VDD.n567 99.5127
R18968 VDD.n1930 VDD.n567 99.5127
R18969 VDD.n1930 VDD.n565 99.5127
R18970 VDD.n1934 VDD.n565 99.5127
R18971 VDD.n1934 VDD.n555 99.5127
R18972 VDD.n1942 VDD.n555 99.5127
R18973 VDD.n1942 VDD.n553 99.5127
R18974 VDD.n1946 VDD.n553 99.5127
R18975 VDD.n1946 VDD.n543 99.5127
R18976 VDD.n1954 VDD.n543 99.5127
R18977 VDD.n1954 VDD.n541 99.5127
R18978 VDD.n1958 VDD.n541 99.5127
R18979 VDD.n1958 VDD.n531 99.5127
R18980 VDD.n1966 VDD.n531 99.5127
R18981 VDD.n1966 VDD.n529 99.5127
R18982 VDD.n1970 VDD.n529 99.5127
R18983 VDD.n1970 VDD.n519 99.5127
R18984 VDD.n1978 VDD.n519 99.5127
R18985 VDD.n1978 VDD.n517 99.5127
R18986 VDD.n1982 VDD.n517 99.5127
R18987 VDD.n1982 VDD.n507 99.5127
R18988 VDD.n1990 VDD.n507 99.5127
R18989 VDD.n1990 VDD.n505 99.5127
R18990 VDD.n1994 VDD.n505 99.5127
R18991 VDD.n1994 VDD.n495 99.5127
R18992 VDD.n2002 VDD.n495 99.5127
R18993 VDD.n2002 VDD.n493 99.5127
R18994 VDD.n2006 VDD.n493 99.5127
R18995 VDD.n2006 VDD.n483 99.5127
R18996 VDD.n2014 VDD.n483 99.5127
R18997 VDD.n2014 VDD.n481 99.5127
R18998 VDD.n2018 VDD.n481 99.5127
R18999 VDD.n2018 VDD.n470 99.5127
R19000 VDD.n2028 VDD.n470 99.5127
R19001 VDD.n2028 VDD.n468 99.5127
R19002 VDD.n2032 VDD.n468 99.5127
R19003 VDD.n2032 VDD.n453 99.5127
R19004 VDD.n2079 VDD.n453 99.5127
R19005 VDD.n2079 VDD.n451 99.5127
R19006 VDD.n2083 VDD.n451 99.5127
R19007 VDD.n2083 VDD.n440 99.5127
R19008 VDD.n2678 VDD.n2677 99.5127
R19009 VDD.n2675 VDD.n2666 99.5127
R19010 VDD.n2671 VDD.n2670 99.5127
R19011 VDD.n2750 VDD.n150 99.5127
R19012 VDD.n2748 VDD.n2747 99.5127
R19013 VDD.n2745 VDD.n153 99.5127
R19014 VDD.n2740 VDD.n2739 99.5127
R19015 VDD.n2131 VDD.n420 99.5127
R19016 VDD.n2273 VDD.n420 99.5127
R19017 VDD.n2273 VDD.n414 99.5127
R19018 VDD.n2270 VDD.n414 99.5127
R19019 VDD.n2270 VDD.n408 99.5127
R19020 VDD.n2267 VDD.n408 99.5127
R19021 VDD.n2267 VDD.n402 99.5127
R19022 VDD.n2264 VDD.n402 99.5127
R19023 VDD.n2264 VDD.n395 99.5127
R19024 VDD.n2261 VDD.n395 99.5127
R19025 VDD.n2261 VDD.n388 99.5127
R19026 VDD.n2258 VDD.n388 99.5127
R19027 VDD.n2258 VDD.n383 99.5127
R19028 VDD.n2255 VDD.n383 99.5127
R19029 VDD.n2255 VDD.n378 99.5127
R19030 VDD.n2252 VDD.n378 99.5127
R19031 VDD.n2252 VDD.n372 99.5127
R19032 VDD.n2249 VDD.n372 99.5127
R19033 VDD.n2249 VDD.n366 99.5127
R19034 VDD.n2246 VDD.n366 99.5127
R19035 VDD.n2246 VDD.n360 99.5127
R19036 VDD.n2243 VDD.n360 99.5127
R19037 VDD.n2243 VDD.n354 99.5127
R19038 VDD.n2240 VDD.n354 99.5127
R19039 VDD.n2240 VDD.n348 99.5127
R19040 VDD.n2237 VDD.n348 99.5127
R19041 VDD.n2237 VDD.n342 99.5127
R19042 VDD.n2234 VDD.n342 99.5127
R19043 VDD.n2234 VDD.n335 99.5127
R19044 VDD.n2231 VDD.n335 99.5127
R19045 VDD.n2231 VDD.n329 99.5127
R19046 VDD.n2228 VDD.n329 99.5127
R19047 VDD.n2228 VDD.n324 99.5127
R19048 VDD.n2225 VDD.n324 99.5127
R19049 VDD.n2225 VDD.n318 99.5127
R19050 VDD.n2222 VDD.n318 99.5127
R19051 VDD.n2222 VDD.n312 99.5127
R19052 VDD.n2219 VDD.n312 99.5127
R19053 VDD.n2219 VDD.n306 99.5127
R19054 VDD.n2216 VDD.n306 99.5127
R19055 VDD.n2216 VDD.n300 99.5127
R19056 VDD.n2213 VDD.n300 99.5127
R19057 VDD.n2213 VDD.n294 99.5127
R19058 VDD.n2210 VDD.n294 99.5127
R19059 VDD.n2210 VDD.n288 99.5127
R19060 VDD.n2207 VDD.n288 99.5127
R19061 VDD.n2207 VDD.n281 99.5127
R19062 VDD.n2204 VDD.n281 99.5127
R19063 VDD.n2204 VDD.n274 99.5127
R19064 VDD.n2201 VDD.n274 99.5127
R19065 VDD.n2201 VDD.n269 99.5127
R19066 VDD.n2198 VDD.n269 99.5127
R19067 VDD.n2198 VDD.n264 99.5127
R19068 VDD.n2195 VDD.n264 99.5127
R19069 VDD.n2195 VDD.n258 99.5127
R19070 VDD.n2192 VDD.n258 99.5127
R19071 VDD.n2192 VDD.n252 99.5127
R19072 VDD.n2189 VDD.n252 99.5127
R19073 VDD.n2189 VDD.n246 99.5127
R19074 VDD.n2186 VDD.n246 99.5127
R19075 VDD.n2186 VDD.n240 99.5127
R19076 VDD.n2183 VDD.n240 99.5127
R19077 VDD.n2183 VDD.n234 99.5127
R19078 VDD.n2180 VDD.n234 99.5127
R19079 VDD.n2180 VDD.n228 99.5127
R19080 VDD.n2177 VDD.n228 99.5127
R19081 VDD.n2177 VDD.n222 99.5127
R19082 VDD.n2174 VDD.n222 99.5127
R19083 VDD.n2174 VDD.n216 99.5127
R19084 VDD.n2171 VDD.n216 99.5127
R19085 VDD.n2171 VDD.n210 99.5127
R19086 VDD.n2168 VDD.n210 99.5127
R19087 VDD.n2168 VDD.n204 99.5127
R19088 VDD.n2165 VDD.n204 99.5127
R19089 VDD.n2165 VDD.n198 99.5127
R19090 VDD.n2162 VDD.n198 99.5127
R19091 VDD.n2162 VDD.n191 99.5127
R19092 VDD.n2159 VDD.n191 99.5127
R19093 VDD.n2159 VDD.n184 99.5127
R19094 VDD.n184 VDD.n160 99.5127
R19095 VDD.n2733 VDD.n160 99.5127
R19096 VDD.n2733 VDD.n158 99.5127
R19097 VDD.n2135 VDD.n423 99.5127
R19098 VDD.n2139 VDD.n2138 99.5127
R19099 VDD.n2143 VDD.n2142 99.5127
R19100 VDD.n2147 VDD.n2146 99.5127
R19101 VDD.n2151 VDD.n2150 99.5127
R19102 VDD.n2155 VDD.n2154 99.5127
R19103 VDD.n2278 VDD.n2130 99.5127
R19104 VDD.n2437 VDD.n421 99.5127
R19105 VDD.n2437 VDD.n411 99.5127
R19106 VDD.n2445 VDD.n411 99.5127
R19107 VDD.n2445 VDD.n409 99.5127
R19108 VDD.n2449 VDD.n409 99.5127
R19109 VDD.n2449 VDD.n399 99.5127
R19110 VDD.n2457 VDD.n399 99.5127
R19111 VDD.n2457 VDD.n397 99.5127
R19112 VDD.n2461 VDD.n397 99.5127
R19113 VDD.n2461 VDD.n386 99.5127
R19114 VDD.n2469 VDD.n386 99.5127
R19115 VDD.n2469 VDD.n384 99.5127
R19116 VDD.n2473 VDD.n384 99.5127
R19117 VDD.n2473 VDD.n375 99.5127
R19118 VDD.n2481 VDD.n375 99.5127
R19119 VDD.n2481 VDD.n373 99.5127
R19120 VDD.n2485 VDD.n373 99.5127
R19121 VDD.n2485 VDD.n363 99.5127
R19122 VDD.n2493 VDD.n363 99.5127
R19123 VDD.n2493 VDD.n361 99.5127
R19124 VDD.n2497 VDD.n361 99.5127
R19125 VDD.n2497 VDD.n351 99.5127
R19126 VDD.n2505 VDD.n351 99.5127
R19127 VDD.n2505 VDD.n349 99.5127
R19128 VDD.n2509 VDD.n349 99.5127
R19129 VDD.n2509 VDD.n339 99.5127
R19130 VDD.n2517 VDD.n339 99.5127
R19131 VDD.n2517 VDD.n337 99.5127
R19132 VDD.n2521 VDD.n337 99.5127
R19133 VDD.n2521 VDD.n327 99.5127
R19134 VDD.n2529 VDD.n327 99.5127
R19135 VDD.n2529 VDD.n325 99.5127
R19136 VDD.n2533 VDD.n325 99.5127
R19137 VDD.n2533 VDD.n315 99.5127
R19138 VDD.n2541 VDD.n315 99.5127
R19139 VDD.n2541 VDD.n313 99.5127
R19140 VDD.n2545 VDD.n313 99.5127
R19141 VDD.n2545 VDD.n303 99.5127
R19142 VDD.n2553 VDD.n303 99.5127
R19143 VDD.n2553 VDD.n301 99.5127
R19144 VDD.n2557 VDD.n301 99.5127
R19145 VDD.n2557 VDD.n291 99.5127
R19146 VDD.n2565 VDD.n291 99.5127
R19147 VDD.n2565 VDD.n289 99.5127
R19148 VDD.n2569 VDD.n289 99.5127
R19149 VDD.n2569 VDD.n278 99.5127
R19150 VDD.n2577 VDD.n278 99.5127
R19151 VDD.n2577 VDD.n276 99.5127
R19152 VDD.n2581 VDD.n276 99.5127
R19153 VDD.n2581 VDD.n267 99.5127
R19154 VDD.n2589 VDD.n267 99.5127
R19155 VDD.n2589 VDD.n265 99.5127
R19156 VDD.n2593 VDD.n265 99.5127
R19157 VDD.n2593 VDD.n255 99.5127
R19158 VDD.n2601 VDD.n255 99.5127
R19159 VDD.n2601 VDD.n253 99.5127
R19160 VDD.n2605 VDD.n253 99.5127
R19161 VDD.n2605 VDD.n243 99.5127
R19162 VDD.n2613 VDD.n243 99.5127
R19163 VDD.n2613 VDD.n241 99.5127
R19164 VDD.n2617 VDD.n241 99.5127
R19165 VDD.n2617 VDD.n231 99.5127
R19166 VDD.n2625 VDD.n231 99.5127
R19167 VDD.n2625 VDD.n229 99.5127
R19168 VDD.n2629 VDD.n229 99.5127
R19169 VDD.n2629 VDD.n219 99.5127
R19170 VDD.n2637 VDD.n219 99.5127
R19171 VDD.n2637 VDD.n217 99.5127
R19172 VDD.n2641 VDD.n217 99.5127
R19173 VDD.n2641 VDD.n207 99.5127
R19174 VDD.n2649 VDD.n207 99.5127
R19175 VDD.n2649 VDD.n205 99.5127
R19176 VDD.n2653 VDD.n205 99.5127
R19177 VDD.n2653 VDD.n195 99.5127
R19178 VDD.n2661 VDD.n195 99.5127
R19179 VDD.n2661 VDD.n192 99.5127
R19180 VDD.n2687 VDD.n192 99.5127
R19181 VDD.n2687 VDD.n193 99.5127
R19182 VDD.n193 VDD.n185 99.5127
R19183 VDD.n2682 VDD.n185 99.5127
R19184 VDD.n2682 VDD.n164 99.5127
R19185 VDD.n2679 VDD.n164 99.5127
R19186 VDD.n2068 VDD.n2067 99.5127
R19187 VDD.n2064 VDD.n2063 99.5127
R19188 VDD.n2060 VDD.n2059 99.5127
R19189 VDD.n2056 VDD.n2055 99.5127
R19190 VDD.n2052 VDD.n2051 99.5127
R19191 VDD.n2048 VDD.n2047 99.5127
R19192 VDD.n2044 VDD.n432 99.5127
R19193 VDD.n900 VDD.n696 99.5127
R19194 VDD.n897 VDD.n696 99.5127
R19195 VDD.n897 VDD.n690 99.5127
R19196 VDD.n894 VDD.n690 99.5127
R19197 VDD.n894 VDD.n684 99.5127
R19198 VDD.n891 VDD.n684 99.5127
R19199 VDD.n891 VDD.n678 99.5127
R19200 VDD.n888 VDD.n678 99.5127
R19201 VDD.n888 VDD.n671 99.5127
R19202 VDD.n885 VDD.n671 99.5127
R19203 VDD.n885 VDD.n665 99.5127
R19204 VDD.n882 VDD.n665 99.5127
R19205 VDD.n882 VDD.n659 99.5127
R19206 VDD.n879 VDD.n659 99.5127
R19207 VDD.n879 VDD.n653 99.5127
R19208 VDD.n876 VDD.n653 99.5127
R19209 VDD.n876 VDD.n648 99.5127
R19210 VDD.n873 VDD.n648 99.5127
R19211 VDD.n873 VDD.n642 99.5127
R19212 VDD.n870 VDD.n642 99.5127
R19213 VDD.n870 VDD.n636 99.5127
R19214 VDD.n867 VDD.n636 99.5127
R19215 VDD.n867 VDD.n630 99.5127
R19216 VDD.n864 VDD.n630 99.5127
R19217 VDD.n864 VDD.n624 99.5127
R19218 VDD.n861 VDD.n624 99.5127
R19219 VDD.n861 VDD.n618 99.5127
R19220 VDD.n858 VDD.n618 99.5127
R19221 VDD.n858 VDD.n612 99.5127
R19222 VDD.n855 VDD.n612 99.5127
R19223 VDD.n855 VDD.n606 99.5127
R19224 VDD.n852 VDD.n606 99.5127
R19225 VDD.n852 VDD.n600 99.5127
R19226 VDD.n849 VDD.n600 99.5127
R19227 VDD.n849 VDD.n594 99.5127
R19228 VDD.n846 VDD.n594 99.5127
R19229 VDD.n846 VDD.n588 99.5127
R19230 VDD.n843 VDD.n588 99.5127
R19231 VDD.n843 VDD.n582 99.5127
R19232 VDD.n840 VDD.n582 99.5127
R19233 VDD.n840 VDD.n576 99.5127
R19234 VDD.n837 VDD.n576 99.5127
R19235 VDD.n837 VDD.n570 99.5127
R19236 VDD.n834 VDD.n570 99.5127
R19237 VDD.n834 VDD.n564 99.5127
R19238 VDD.n831 VDD.n564 99.5127
R19239 VDD.n831 VDD.n558 99.5127
R19240 VDD.n828 VDD.n558 99.5127
R19241 VDD.n828 VDD.n551 99.5127
R19242 VDD.n825 VDD.n551 99.5127
R19243 VDD.n825 VDD.n545 99.5127
R19244 VDD.n822 VDD.n545 99.5127
R19245 VDD.n822 VDD.n540 99.5127
R19246 VDD.n819 VDD.n540 99.5127
R19247 VDD.n819 VDD.n534 99.5127
R19248 VDD.n816 VDD.n534 99.5127
R19249 VDD.n816 VDD.n528 99.5127
R19250 VDD.n813 VDD.n528 99.5127
R19251 VDD.n813 VDD.n522 99.5127
R19252 VDD.n810 VDD.n522 99.5127
R19253 VDD.n810 VDD.n516 99.5127
R19254 VDD.n807 VDD.n516 99.5127
R19255 VDD.n807 VDD.n510 99.5127
R19256 VDD.n804 VDD.n510 99.5127
R19257 VDD.n804 VDD.n504 99.5127
R19258 VDD.n801 VDD.n504 99.5127
R19259 VDD.n801 VDD.n498 99.5127
R19260 VDD.n798 VDD.n498 99.5127
R19261 VDD.n798 VDD.n492 99.5127
R19262 VDD.n795 VDD.n492 99.5127
R19263 VDD.n795 VDD.n486 99.5127
R19264 VDD.n792 VDD.n486 99.5127
R19265 VDD.n792 VDD.n480 99.5127
R19266 VDD.n789 VDD.n480 99.5127
R19267 VDD.n789 VDD.n473 99.5127
R19268 VDD.n473 VDD.n464 99.5127
R19269 VDD.n2034 VDD.n464 99.5127
R19270 VDD.n2035 VDD.n2034 99.5127
R19271 VDD.n2035 VDD.n456 99.5127
R19272 VDD.n2038 VDD.n456 99.5127
R19273 VDD.n2038 VDD.n449 99.5127
R19274 VDD.n2041 VDD.n449 99.5127
R19275 VDD.n773 VDD.n772 99.5127
R19276 VDD.n777 VDD.n776 99.5127
R19277 VDD.n781 VDD.n780 99.5127
R19278 VDD.n913 VDD.n783 99.5127
R19279 VDD.n911 VDD.n910 99.5127
R19280 VDD.n907 VDD.n906 99.5127
R19281 VDD.n903 VDD.n713 99.5127
R19282 VDD.n1804 VDD.n693 99.5127
R19283 VDD.n1804 VDD.n691 99.5127
R19284 VDD.n1808 VDD.n691 99.5127
R19285 VDD.n1808 VDD.n681 99.5127
R19286 VDD.n1816 VDD.n681 99.5127
R19287 VDD.n1816 VDD.n679 99.5127
R19288 VDD.n1820 VDD.n679 99.5127
R19289 VDD.n1820 VDD.n668 99.5127
R19290 VDD.n1828 VDD.n668 99.5127
R19291 VDD.n1828 VDD.n666 99.5127
R19292 VDD.n1832 VDD.n666 99.5127
R19293 VDD.n1832 VDD.n656 99.5127
R19294 VDD.n1840 VDD.n656 99.5127
R19295 VDD.n1840 VDD.n654 99.5127
R19296 VDD.n1844 VDD.n654 99.5127
R19297 VDD.n1844 VDD.n645 99.5127
R19298 VDD.n1852 VDD.n645 99.5127
R19299 VDD.n1852 VDD.n643 99.5127
R19300 VDD.n1856 VDD.n643 99.5127
R19301 VDD.n1856 VDD.n633 99.5127
R19302 VDD.n1864 VDD.n633 99.5127
R19303 VDD.n1864 VDD.n631 99.5127
R19304 VDD.n1868 VDD.n631 99.5127
R19305 VDD.n1868 VDD.n621 99.5127
R19306 VDD.n1876 VDD.n621 99.5127
R19307 VDD.n1876 VDD.n619 99.5127
R19308 VDD.n1880 VDD.n619 99.5127
R19309 VDD.n1880 VDD.n609 99.5127
R19310 VDD.n1888 VDD.n609 99.5127
R19311 VDD.n1888 VDD.n607 99.5127
R19312 VDD.n1892 VDD.n607 99.5127
R19313 VDD.n1892 VDD.n597 99.5127
R19314 VDD.n1900 VDD.n597 99.5127
R19315 VDD.n1900 VDD.n595 99.5127
R19316 VDD.n1904 VDD.n595 99.5127
R19317 VDD.n1904 VDD.n585 99.5127
R19318 VDD.n1912 VDD.n585 99.5127
R19319 VDD.n1912 VDD.n583 99.5127
R19320 VDD.n1916 VDD.n583 99.5127
R19321 VDD.n1916 VDD.n573 99.5127
R19322 VDD.n1924 VDD.n573 99.5127
R19323 VDD.n1924 VDD.n571 99.5127
R19324 VDD.n1928 VDD.n571 99.5127
R19325 VDD.n1928 VDD.n561 99.5127
R19326 VDD.n1936 VDD.n561 99.5127
R19327 VDD.n1936 VDD.n559 99.5127
R19328 VDD.n1940 VDD.n559 99.5127
R19329 VDD.n1940 VDD.n548 99.5127
R19330 VDD.n1948 VDD.n548 99.5127
R19331 VDD.n1948 VDD.n546 99.5127
R19332 VDD.n1952 VDD.n546 99.5127
R19333 VDD.n1952 VDD.n537 99.5127
R19334 VDD.n1960 VDD.n537 99.5127
R19335 VDD.n1960 VDD.n535 99.5127
R19336 VDD.n1964 VDD.n535 99.5127
R19337 VDD.n1964 VDD.n525 99.5127
R19338 VDD.n1972 VDD.n525 99.5127
R19339 VDD.n1972 VDD.n523 99.5127
R19340 VDD.n1976 VDD.n523 99.5127
R19341 VDD.n1976 VDD.n513 99.5127
R19342 VDD.n1984 VDD.n513 99.5127
R19343 VDD.n1984 VDD.n511 99.5127
R19344 VDD.n1988 VDD.n511 99.5127
R19345 VDD.n1988 VDD.n501 99.5127
R19346 VDD.n1996 VDD.n501 99.5127
R19347 VDD.n1996 VDD.n499 99.5127
R19348 VDD.n2000 VDD.n499 99.5127
R19349 VDD.n2000 VDD.n489 99.5127
R19350 VDD.n2008 VDD.n489 99.5127
R19351 VDD.n2008 VDD.n487 99.5127
R19352 VDD.n2012 VDD.n487 99.5127
R19353 VDD.n2012 VDD.n477 99.5127
R19354 VDD.n2020 VDD.n477 99.5127
R19355 VDD.n2020 VDD.n474 99.5127
R19356 VDD.n2026 VDD.n474 99.5127
R19357 VDD.n2026 VDD.n475 99.5127
R19358 VDD.n475 VDD.n467 99.5127
R19359 VDD.n467 VDD.n457 99.5127
R19360 VDD.n2077 VDD.n457 99.5127
R19361 VDD.n2077 VDD.n458 99.5127
R19362 VDD.n458 VDD.n450 99.5127
R19363 VDD.n2072 VDD.n450 99.5127
R19364 VDD.n1796 VDD.t128 98.1776
R19365 VDD.n151 VDD.t130 98.1776
R19366 VDD.n2431 VDD.n2117 94.5317
R19367 VDD.n3389 VDD.t137 85.8723
R19368 VDD.n3369 VDD.t134 85.8723
R19369 VDD.n3349 VDD.t138 85.8723
R19370 VDD.n3329 VDD.t127 85.8723
R19371 VDD.n3310 VDD.t132 85.8723
R19372 VDD.n1425 VDD.t104 85.8723
R19373 VDD.n1405 VDD.t99 85.8723
R19374 VDD.n1385 VDD.t103 85.8723
R19375 VDD.n1365 VDD.t133 85.8723
R19376 VDD.n1346 VDD.t141 85.8723
R19377 VDD.n2432 VDD.n2431 72.8958
R19378 VDD.n2431 VDD.n2124 72.8958
R19379 VDD.n2431 VDD.n2125 72.8958
R19380 VDD.n2431 VDD.n2126 72.8958
R19381 VDD.n2431 VDD.n2127 72.8958
R19382 VDD.n2431 VDD.n2128 72.8958
R19383 VDD.n2431 VDD.n2129 72.8958
R19384 VDD.n2738 VDD.n151 72.8958
R19385 VDD.n157 VDD.n151 72.8958
R19386 VDD.n2746 VDD.n151 72.8958
R19387 VDD.n2749 VDD.n151 72.8958
R19388 VDD.n2669 VDD.n151 72.8958
R19389 VDD.n2668 VDD.n151 72.8958
R19390 VDD.n2676 VDD.n151 72.8958
R19391 VDD.n1797 VDD.n1796 72.8958
R19392 VDD.n1796 VDD.n700 72.8958
R19393 VDD.n1796 VDD.n701 72.8958
R19394 VDD.n1796 VDD.n702 72.8958
R19395 VDD.n1796 VDD.n703 72.8958
R19396 VDD.n1796 VDD.n704 72.8958
R19397 VDD.n1796 VDD.n705 72.8958
R19398 VDD.n2117 VDD.n433 72.8958
R19399 VDD.n2117 VDD.n434 72.8958
R19400 VDD.n2117 VDD.n435 72.8958
R19401 VDD.n2117 VDD.n436 72.8958
R19402 VDD.n2117 VDD.n437 72.8958
R19403 VDD.n2117 VDD.n438 72.8958
R19404 VDD.n2117 VDD.n439 72.8958
R19405 VDD.n2431 VDD.n2430 72.8958
R19406 VDD.n2431 VDD.n2118 72.8958
R19407 VDD.n2431 VDD.n2119 72.8958
R19408 VDD.n2431 VDD.n2120 72.8958
R19409 VDD.n2431 VDD.n2121 72.8958
R19410 VDD.n2431 VDD.n2122 72.8958
R19411 VDD.n2431 VDD.n2123 72.8958
R19412 VDD.n2702 VDD.n151 72.8958
R19413 VDD.n179 VDD.n151 72.8958
R19414 VDD.n2710 VDD.n151 72.8958
R19415 VDD.n174 VDD.n151 72.8958
R19416 VDD.n2718 VDD.n151 72.8958
R19417 VDD.n171 VDD.n151 72.8958
R19418 VDD.n2725 VDD.n151 72.8958
R19419 VDD.n2117 VDD.n431 72.8958
R19420 VDD.n2117 VDD.n430 72.8958
R19421 VDD.n2117 VDD.n429 72.8958
R19422 VDD.n2117 VDD.n428 72.8958
R19423 VDD.n2117 VDD.n427 72.8958
R19424 VDD.n2117 VDD.n426 72.8958
R19425 VDD.n2117 VDD.n425 72.8958
R19426 VDD.n1796 VDD.n706 72.8958
R19427 VDD.n1796 VDD.n707 72.8958
R19428 VDD.n1796 VDD.n708 72.8958
R19429 VDD.n1796 VDD.n709 72.8958
R19430 VDD.n1796 VDD.n710 72.8958
R19431 VDD.n1796 VDD.n711 72.8958
R19432 VDD.n1796 VDD.n712 72.8958
R19433 VDD.n1043 VDD.n1042 69.6247
R19434 VDD.n1059 VDD.n1058 69.6247
R19435 VDD.n1077 VDD.n1076 69.6247
R19436 VDD.n1094 VDD.n1093 69.6247
R19437 VDD.n1111 VDD.n1110 69.6247
R19438 VDD.n1511 VDD.n1510 69.6247
R19439 VDD.n957 VDD.n956 69.6247
R19440 VDD.n926 VDD.n925 69.6247
R19441 VDD.n754 VDD.n753 69.6247
R19442 VDD.n730 VDD.n729 69.6247
R19443 VDD.n3033 VDD.n3032 69.6247
R19444 VDD.n3043 VDD.n3042 69.6247
R19445 VDD.n3051 VDD.n3050 69.6247
R19446 VDD.n3060 VDD.n3059 69.6247
R19447 VDD.n3070 VDD.n3069 69.6247
R19448 VDD.n115 VDD.n114 69.6247
R19449 VDD.n141 VDD.n140 69.6247
R19450 VDD.n2857 VDD.n2856 69.6247
R19451 VDD.n65 VDD.n64 69.6247
R19452 VDD.n2757 VDD.n2756 69.6247
R19453 VDD.n1121 VDD.n1038 66.2847
R19454 VDD.n1129 VDD.n1038 66.2847
R19455 VDD.n1131 VDD.n1038 66.2847
R19456 VDD.n1141 VDD.n1038 66.2847
R19457 VDD.n1144 VDD.n1038 66.2847
R19458 VDD.n1108 VDD.n1038 66.2847
R19459 VDD.n1153 VDD.n1038 66.2847
R19460 VDD.n1155 VDD.n1038 66.2847
R19461 VDD.n1163 VDD.n1038 66.2847
R19462 VDD.n1165 VDD.n1038 66.2847
R19463 VDD.n1175 VDD.n1038 66.2847
R19464 VDD.n1178 VDD.n1038 66.2847
R19465 VDD.n1091 VDD.n1038 66.2847
R19466 VDD.n1187 VDD.n1038 66.2847
R19467 VDD.n1189 VDD.n1038 66.2847
R19468 VDD.n1197 VDD.n1038 66.2847
R19469 VDD.n1199 VDD.n1038 66.2847
R19470 VDD.n1209 VDD.n1038 66.2847
R19471 VDD.n1212 VDD.n1038 66.2847
R19472 VDD.n1074 VDD.n1038 66.2847
R19473 VDD.n1221 VDD.n1038 66.2847
R19474 VDD.n1223 VDD.n1038 66.2847
R19475 VDD.n1231 VDD.n1038 66.2847
R19476 VDD.n1233 VDD.n1038 66.2847
R19477 VDD.n1242 VDD.n1038 66.2847
R19478 VDD.n1244 VDD.n1038 66.2847
R19479 VDD.n1252 VDD.n1038 66.2847
R19480 VDD.n1254 VDD.n1038 66.2847
R19481 VDD.n1262 VDD.n1038 66.2847
R19482 VDD.n1264 VDD.n1038 66.2847
R19483 VDD.n1272 VDD.n1038 66.2847
R19484 VDD.n1275 VDD.n1038 66.2847
R19485 VDD.n1045 VDD.n1038 66.2847
R19486 VDD.n1559 VDD.n721 66.2847
R19487 VDD.n953 VDD.n721 66.2847
R19488 VDD.n948 VDD.n721 66.2847
R19489 VDD.n945 VDD.n721 66.2847
R19490 VDD.n940 VDD.n721 66.2847
R19491 VDD.n937 VDD.n721 66.2847
R19492 VDD.n932 VDD.n721 66.2847
R19493 VDD.n929 VDD.n721 66.2847
R19494 VDD.n922 VDD.n721 66.2847
R19495 VDD.n919 VDD.n721 66.2847
R19496 VDD.n1591 VDD.n721 66.2847
R19497 VDD.n766 VDD.n721 66.2847
R19498 VDD.n1598 VDD.n721 66.2847
R19499 VDD.n760 VDD.n721 66.2847
R19500 VDD.n755 VDD.n721 66.2847
R19501 VDD.n1609 VDD.n721 66.2847
R19502 VDD.n747 VDD.n721 66.2847
R19503 VDD.n1616 VDD.n721 66.2847
R19504 VDD.n740 VDD.n721 66.2847
R19505 VDD.n1623 VDD.n721 66.2847
R19506 VDD.n734 VDD.n721 66.2847
R19507 VDD.n1632 VDD.n721 66.2847
R19508 VDD.n726 VDD.n721 66.2847
R19509 VDD.n1639 VDD.n721 66.2847
R19510 VDD.n1642 VDD.n721 66.2847
R19511 VDD.n1518 VDD.n721 66.2847
R19512 VDD.n1527 VDD.n721 66.2847
R19513 VDD.n1530 VDD.n721 66.2847
R19514 VDD.n1512 VDD.n721 66.2847
R19515 VDD.n1537 VDD.n721 66.2847
R19516 VDD.n1505 VDD.n721 66.2847
R19517 VDD.n1544 VDD.n721 66.2847
R19518 VDD.n1547 VDD.n721 66.2847
R19519 VDD.n1493 VDD.n721 66.2847
R19520 VDD.n2909 VDD.n2908 66.2847
R19521 VDD.n2909 VDD.n68 66.2847
R19522 VDD.n2909 VDD.n69 66.2847
R19523 VDD.n2909 VDD.n70 66.2847
R19524 VDD.n2909 VDD.n71 66.2847
R19525 VDD.n2909 VDD.n72 66.2847
R19526 VDD.n2909 VDD.n73 66.2847
R19527 VDD.n2909 VDD.n74 66.2847
R19528 VDD.n2909 VDD.n75 66.2847
R19529 VDD.n2909 VDD.n76 66.2847
R19530 VDD.n2909 VDD.n77 66.2847
R19531 VDD.n2909 VDD.n78 66.2847
R19532 VDD.n2909 VDD.n79 66.2847
R19533 VDD.n2909 VDD.n80 66.2847
R19534 VDD.n2909 VDD.n81 66.2847
R19535 VDD.n2909 VDD.n82 66.2847
R19536 VDD.n2909 VDD.n83 66.2847
R19537 VDD.n2909 VDD.n84 66.2847
R19538 VDD.n2909 VDD.n85 66.2847
R19539 VDD.n2909 VDD.n86 66.2847
R19540 VDD.n2909 VDD.n87 66.2847
R19541 VDD.n2909 VDD.n88 66.2847
R19542 VDD.n2909 VDD.n89 66.2847
R19543 VDD.n2909 VDD.n90 66.2847
R19544 VDD.n2909 VDD.n91 66.2847
R19545 VDD.n2909 VDD.n92 66.2847
R19546 VDD.n2909 VDD.n93 66.2847
R19547 VDD.n2909 VDD.n94 66.2847
R19548 VDD.n2909 VDD.n95 66.2847
R19549 VDD.n2909 VDD.n96 66.2847
R19550 VDD.n2909 VDD.n97 66.2847
R19551 VDD.n2909 VDD.n98 66.2847
R19552 VDD.n2909 VDD.n99 66.2847
R19553 VDD.n3271 VDD.n3270 66.2847
R19554 VDD.n3271 VDD.n3030 66.2847
R19555 VDD.n3271 VDD.n3029 66.2847
R19556 VDD.n3271 VDD.n3028 66.2847
R19557 VDD.n3271 VDD.n3027 66.2847
R19558 VDD.n3271 VDD.n3026 66.2847
R19559 VDD.n3271 VDD.n3025 66.2847
R19560 VDD.n3271 VDD.n3024 66.2847
R19561 VDD.n3271 VDD.n3023 66.2847
R19562 VDD.n3271 VDD.n3022 66.2847
R19563 VDD.n3271 VDD.n3021 66.2847
R19564 VDD.n3271 VDD.n3020 66.2847
R19565 VDD.n3271 VDD.n3019 66.2847
R19566 VDD.n3271 VDD.n3018 66.2847
R19567 VDD.n3271 VDD.n3017 66.2847
R19568 VDD.n3271 VDD.n3016 66.2847
R19569 VDD.n3271 VDD.n3015 66.2847
R19570 VDD.n3271 VDD.n3014 66.2847
R19571 VDD.n3271 VDD.n3013 66.2847
R19572 VDD.n3271 VDD.n3012 66.2847
R19573 VDD.n3271 VDD.n3011 66.2847
R19574 VDD.n3271 VDD.n3010 66.2847
R19575 VDD.n3271 VDD.n3009 66.2847
R19576 VDD.n3271 VDD.n3008 66.2847
R19577 VDD.n3271 VDD.n3007 66.2847
R19578 VDD.n3271 VDD.n3006 66.2847
R19579 VDD.n3271 VDD.n3005 66.2847
R19580 VDD.n3271 VDD.n3004 66.2847
R19581 VDD.n3271 VDD.n3003 66.2847
R19582 VDD.n3271 VDD.n3002 66.2847
R19583 VDD.n3271 VDD.n3001 66.2847
R19584 VDD.n3271 VDD.n3000 66.2847
R19585 VDD.n3271 VDD.n2999 66.2847
R19586 VDD.n3271 VDD.n2998 66.2847
R19587 VDD.n3082 VDD.n2998 52.4337
R19588 VDD.n3086 VDD.n2999 52.4337
R19589 VDD.n3092 VDD.n3000 52.4337
R19590 VDD.n3096 VDD.n3001 52.4337
R19591 VDD.n3102 VDD.n3002 52.4337
R19592 VDD.n3106 VDD.n3003 52.4337
R19593 VDD.n3112 VDD.n3004 52.4337
R19594 VDD.n3116 VDD.n3005 52.4337
R19595 VDD.n3122 VDD.n3006 52.4337
R19596 VDD.n3126 VDD.n3007 52.4337
R19597 VDD.n3132 VDD.n3008 52.4337
R19598 VDD.n3136 VDD.n3009 52.4337
R19599 VDD.n3142 VDD.n3010 52.4337
R19600 VDD.n3146 VDD.n3011 52.4337
R19601 VDD.n3152 VDD.n3012 52.4337
R19602 VDD.n3156 VDD.n3013 52.4337
R19603 VDD.n3162 VDD.n3014 52.4337
R19604 VDD.n3166 VDD.n3015 52.4337
R19605 VDD.n3172 VDD.n3016 52.4337
R19606 VDD.n3176 VDD.n3017 52.4337
R19607 VDD.n3180 VDD.n3018 52.4337
R19608 VDD.n3186 VDD.n3019 52.4337
R19609 VDD.n3190 VDD.n3020 52.4337
R19610 VDD.n3196 VDD.n3021 52.4337
R19611 VDD.n3200 VDD.n3022 52.4337
R19612 VDD.n3206 VDD.n3023 52.4337
R19613 VDD.n3211 VDD.n3024 52.4337
R19614 VDD.n3217 VDD.n3025 52.4337
R19615 VDD.n3221 VDD.n3026 52.4337
R19616 VDD.n3227 VDD.n3027 52.4337
R19617 VDD.n3231 VDD.n3028 52.4337
R19618 VDD.n3237 VDD.n3029 52.4337
R19619 VDD.n3240 VDD.n3030 52.4337
R19620 VDD.n3270 VDD.n3269 52.4337
R19621 VDD.n2908 VDD.n2907 52.4337
R19622 VDD.n2902 VDD.n68 52.4337
R19623 VDD.n2899 VDD.n69 52.4337
R19624 VDD.n2895 VDD.n70 52.4337
R19625 VDD.n2891 VDD.n71 52.4337
R19626 VDD.n2887 VDD.n72 52.4337
R19627 VDD.n2883 VDD.n73 52.4337
R19628 VDD.n2879 VDD.n74 52.4337
R19629 VDD.n2875 VDD.n75 52.4337
R19630 VDD.n2871 VDD.n76 52.4337
R19631 VDD.n2867 VDD.n77 52.4337
R19632 VDD.n2863 VDD.n78 52.4337
R19633 VDD.n2859 VDD.n79 52.4337
R19634 VDD.n2851 VDD.n80 52.4337
R19635 VDD.n2847 VDD.n81 52.4337
R19636 VDD.n2843 VDD.n82 52.4337
R19637 VDD.n2839 VDD.n83 52.4337
R19638 VDD.n2835 VDD.n84 52.4337
R19639 VDD.n2831 VDD.n85 52.4337
R19640 VDD.n2827 VDD.n86 52.4337
R19641 VDD.n2821 VDD.n87 52.4337
R19642 VDD.n2817 VDD.n88 52.4337
R19643 VDD.n2813 VDD.n89 52.4337
R19644 VDD.n2809 VDD.n90 52.4337
R19645 VDD.n2805 VDD.n91 52.4337
R19646 VDD.n2801 VDD.n92 52.4337
R19647 VDD.n2797 VDD.n93 52.4337
R19648 VDD.n2793 VDD.n94 52.4337
R19649 VDD.n2789 VDD.n95 52.4337
R19650 VDD.n2785 VDD.n96 52.4337
R19651 VDD.n2781 VDD.n97 52.4337
R19652 VDD.n2777 VDD.n98 52.4337
R19653 VDD.n2773 VDD.n99 52.4337
R19654 VDD.n1494 VDD.n1493 52.4337
R19655 VDD.n1547 VDD.n1546 52.4337
R19656 VDD.n1544 VDD.n1543 52.4337
R19657 VDD.n1539 VDD.n1505 52.4337
R19658 VDD.n1537 VDD.n1536 52.4337
R19659 VDD.n1513 VDD.n1512 52.4337
R19660 VDD.n1530 VDD.n1529 52.4337
R19661 VDD.n1527 VDD.n1526 52.4337
R19662 VDD.n1518 VDD.n720 52.4337
R19663 VDD.n1642 VDD.n1641 52.4337
R19664 VDD.n1639 VDD.n1638 52.4337
R19665 VDD.n1634 VDD.n726 52.4337
R19666 VDD.n1632 VDD.n1631 52.4337
R19667 VDD.n1625 VDD.n734 52.4337
R19668 VDD.n1623 VDD.n1622 52.4337
R19669 VDD.n1618 VDD.n740 52.4337
R19670 VDD.n1616 VDD.n1615 52.4337
R19671 VDD.n1611 VDD.n747 52.4337
R19672 VDD.n1609 VDD.n1608 52.4337
R19673 VDD.n756 VDD.n755 52.4337
R19674 VDD.n1600 VDD.n760 52.4337
R19675 VDD.n1598 VDD.n1597 52.4337
R19676 VDD.n1593 VDD.n766 52.4337
R19677 VDD.n1591 VDD.n1590 52.4337
R19678 VDD.n920 VDD.n919 52.4337
R19679 VDD.n923 VDD.n922 52.4337
R19680 VDD.n930 VDD.n929 52.4337
R19681 VDD.n933 VDD.n932 52.4337
R19682 VDD.n938 VDD.n937 52.4337
R19683 VDD.n941 VDD.n940 52.4337
R19684 VDD.n946 VDD.n945 52.4337
R19685 VDD.n949 VDD.n948 52.4337
R19686 VDD.n954 VDD.n953 52.4337
R19687 VDD.n1559 VDD.n1558 52.4337
R19688 VDD.n1121 VDD.n1037 52.4337
R19689 VDD.n1129 VDD.n1128 52.4337
R19690 VDD.n1132 VDD.n1131 52.4337
R19691 VDD.n1141 VDD.n1140 52.4337
R19692 VDD.n1144 VDD.n1143 52.4337
R19693 VDD.n1109 VDD.n1108 52.4337
R19694 VDD.n1153 VDD.n1152 52.4337
R19695 VDD.n1156 VDD.n1155 52.4337
R19696 VDD.n1163 VDD.n1162 52.4337
R19697 VDD.n1166 VDD.n1165 52.4337
R19698 VDD.n1175 VDD.n1174 52.4337
R19699 VDD.n1178 VDD.n1177 52.4337
R19700 VDD.n1092 VDD.n1091 52.4337
R19701 VDD.n1187 VDD.n1186 52.4337
R19702 VDD.n1190 VDD.n1189 52.4337
R19703 VDD.n1197 VDD.n1196 52.4337
R19704 VDD.n1200 VDD.n1199 52.4337
R19705 VDD.n1209 VDD.n1208 52.4337
R19706 VDD.n1212 VDD.n1211 52.4337
R19707 VDD.n1075 VDD.n1074 52.4337
R19708 VDD.n1221 VDD.n1220 52.4337
R19709 VDD.n1224 VDD.n1223 52.4337
R19710 VDD.n1231 VDD.n1230 52.4337
R19711 VDD.n1234 VDD.n1233 52.4337
R19712 VDD.n1242 VDD.n1241 52.4337
R19713 VDD.n1245 VDD.n1244 52.4337
R19714 VDD.n1252 VDD.n1251 52.4337
R19715 VDD.n1255 VDD.n1254 52.4337
R19716 VDD.n1262 VDD.n1261 52.4337
R19717 VDD.n1265 VDD.n1264 52.4337
R19718 VDD.n1272 VDD.n1271 52.4337
R19719 VDD.n1276 VDD.n1275 52.4337
R19720 VDD.n1046 VDD.n1045 52.4337
R19721 VDD.n1122 VDD.n1121 52.4337
R19722 VDD.n1130 VDD.n1129 52.4337
R19723 VDD.n1131 VDD.n1114 52.4337
R19724 VDD.n1142 VDD.n1141 52.4337
R19725 VDD.n1145 VDD.n1144 52.4337
R19726 VDD.n1108 VDD.n1105 52.4337
R19727 VDD.n1154 VDD.n1153 52.4337
R19728 VDD.n1155 VDD.n1101 52.4337
R19729 VDD.n1164 VDD.n1163 52.4337
R19730 VDD.n1165 VDD.n1097 52.4337
R19731 VDD.n1176 VDD.n1175 52.4337
R19732 VDD.n1179 VDD.n1178 52.4337
R19733 VDD.n1091 VDD.n1088 52.4337
R19734 VDD.n1188 VDD.n1187 52.4337
R19735 VDD.n1189 VDD.n1084 52.4337
R19736 VDD.n1198 VDD.n1197 52.4337
R19737 VDD.n1199 VDD.n1080 52.4337
R19738 VDD.n1210 VDD.n1209 52.4337
R19739 VDD.n1213 VDD.n1212 52.4337
R19740 VDD.n1074 VDD.n1071 52.4337
R19741 VDD.n1222 VDD.n1221 52.4337
R19742 VDD.n1223 VDD.n1067 52.4337
R19743 VDD.n1232 VDD.n1231 52.4337
R19744 VDD.n1233 VDD.n1063 52.4337
R19745 VDD.n1243 VDD.n1242 52.4337
R19746 VDD.n1244 VDD.n1057 52.4337
R19747 VDD.n1253 VDD.n1252 52.4337
R19748 VDD.n1254 VDD.n1053 52.4337
R19749 VDD.n1263 VDD.n1262 52.4337
R19750 VDD.n1264 VDD.n1049 52.4337
R19751 VDD.n1273 VDD.n1272 52.4337
R19752 VDD.n1275 VDD.n1274 52.4337
R19753 VDD.n1045 VDD.n1041 52.4337
R19754 VDD.n1560 VDD.n1559 52.4337
R19755 VDD.n953 VDD.n952 52.4337
R19756 VDD.n948 VDD.n947 52.4337
R19757 VDD.n945 VDD.n944 52.4337
R19758 VDD.n940 VDD.n939 52.4337
R19759 VDD.n937 VDD.n936 52.4337
R19760 VDD.n932 VDD.n931 52.4337
R19761 VDD.n929 VDD.n924 52.4337
R19762 VDD.n922 VDD.n921 52.4337
R19763 VDD.n919 VDD.n767 52.4337
R19764 VDD.n1592 VDD.n1591 52.4337
R19765 VDD.n766 VDD.n761 52.4337
R19766 VDD.n1599 VDD.n1598 52.4337
R19767 VDD.n760 VDD.n759 52.4337
R19768 VDD.n755 VDD.n748 52.4337
R19769 VDD.n1610 VDD.n1609 52.4337
R19770 VDD.n747 VDD.n741 52.4337
R19771 VDD.n1617 VDD.n1616 52.4337
R19772 VDD.n740 VDD.n735 52.4337
R19773 VDD.n1624 VDD.n1623 52.4337
R19774 VDD.n734 VDD.n727 52.4337
R19775 VDD.n1633 VDD.n1632 52.4337
R19776 VDD.n726 VDD.n723 52.4337
R19777 VDD.n1640 VDD.n1639 52.4337
R19778 VDD.n1643 VDD.n1642 52.4337
R19779 VDD.n1519 VDD.n1518 52.4337
R19780 VDD.n1528 VDD.n1527 52.4337
R19781 VDD.n1531 VDD.n1530 52.4337
R19782 VDD.n1512 VDD.n1506 52.4337
R19783 VDD.n1538 VDD.n1537 52.4337
R19784 VDD.n1505 VDD.n1498 52.4337
R19785 VDD.n1545 VDD.n1544 52.4337
R19786 VDD.n1548 VDD.n1547 52.4337
R19787 VDD.n1493 VDD.n962 52.4337
R19788 VDD.n2908 VDD.n101 52.4337
R19789 VDD.n2900 VDD.n68 52.4337
R19790 VDD.n2896 VDD.n69 52.4337
R19791 VDD.n2892 VDD.n70 52.4337
R19792 VDD.n2888 VDD.n71 52.4337
R19793 VDD.n2884 VDD.n72 52.4337
R19794 VDD.n2880 VDD.n73 52.4337
R19795 VDD.n2876 VDD.n74 52.4337
R19796 VDD.n2872 VDD.n75 52.4337
R19797 VDD.n2868 VDD.n76 52.4337
R19798 VDD.n2864 VDD.n77 52.4337
R19799 VDD.n2860 VDD.n78 52.4337
R19800 VDD.n2850 VDD.n79 52.4337
R19801 VDD.n2848 VDD.n80 52.4337
R19802 VDD.n2844 VDD.n81 52.4337
R19803 VDD.n2840 VDD.n82 52.4337
R19804 VDD.n2836 VDD.n83 52.4337
R19805 VDD.n2832 VDD.n84 52.4337
R19806 VDD.n2828 VDD.n85 52.4337
R19807 VDD.n2820 VDD.n86 52.4337
R19808 VDD.n2818 VDD.n87 52.4337
R19809 VDD.n2814 VDD.n88 52.4337
R19810 VDD.n2810 VDD.n89 52.4337
R19811 VDD.n2806 VDD.n90 52.4337
R19812 VDD.n2802 VDD.n91 52.4337
R19813 VDD.n2798 VDD.n92 52.4337
R19814 VDD.n2794 VDD.n93 52.4337
R19815 VDD.n2790 VDD.n94 52.4337
R19816 VDD.n2786 VDD.n95 52.4337
R19817 VDD.n2782 VDD.n96 52.4337
R19818 VDD.n2778 VDD.n97 52.4337
R19819 VDD.n2774 VDD.n98 52.4337
R19820 VDD.n99 VDD.n67 52.4337
R19821 VDD.n3270 VDD.n3031 52.4337
R19822 VDD.n3238 VDD.n3030 52.4337
R19823 VDD.n3230 VDD.n3029 52.4337
R19824 VDD.n3228 VDD.n3028 52.4337
R19825 VDD.n3220 VDD.n3027 52.4337
R19826 VDD.n3218 VDD.n3026 52.4337
R19827 VDD.n3210 VDD.n3025 52.4337
R19828 VDD.n3207 VDD.n3024 52.4337
R19829 VDD.n3199 VDD.n3023 52.4337
R19830 VDD.n3197 VDD.n3022 52.4337
R19831 VDD.n3189 VDD.n3021 52.4337
R19832 VDD.n3187 VDD.n3020 52.4337
R19833 VDD.n3179 VDD.n3019 52.4337
R19834 VDD.n3177 VDD.n3018 52.4337
R19835 VDD.n3173 VDD.n3017 52.4337
R19836 VDD.n3167 VDD.n3016 52.4337
R19837 VDD.n3163 VDD.n3015 52.4337
R19838 VDD.n3157 VDD.n3014 52.4337
R19839 VDD.n3153 VDD.n3013 52.4337
R19840 VDD.n3147 VDD.n3012 52.4337
R19841 VDD.n3143 VDD.n3011 52.4337
R19842 VDD.n3137 VDD.n3010 52.4337
R19843 VDD.n3133 VDD.n3009 52.4337
R19844 VDD.n3127 VDD.n3008 52.4337
R19845 VDD.n3123 VDD.n3007 52.4337
R19846 VDD.n3117 VDD.n3006 52.4337
R19847 VDD.n3113 VDD.n3005 52.4337
R19848 VDD.n3107 VDD.n3004 52.4337
R19849 VDD.n3103 VDD.n3003 52.4337
R19850 VDD.n3097 VDD.n3002 52.4337
R19851 VDD.n3093 VDD.n3001 52.4337
R19852 VDD.n3087 VDD.n3000 52.4337
R19853 VDD.n3083 VDD.n2999 52.4337
R19854 VDD.n3077 VDD.n2998 52.4337
R19855 VDD.n1378 VDD.n1358 47.6734
R19856 VDD.n3342 VDD.n3322 46.8997
R19857 VDD.n1438 VDD.n1437 46.1993
R19858 VDD.n1418 VDD.n1417 46.1993
R19859 VDD.n1398 VDD.n1397 46.1993
R19860 VDD.n1378 VDD.n1377 46.1993
R19861 VDD.n3402 VDD.n3401 45.4256
R19862 VDD.n3382 VDD.n3381 45.4256
R19863 VDD.n3362 VDD.n3361 45.4256
R19864 VDD.n3342 VDD.n3341 45.4256
R19865 VDD.n2725 VDD.n2724 39.2114
R19866 VDD.n2720 VDD.n171 39.2114
R19867 VDD.n2718 VDD.n2717 39.2114
R19868 VDD.n2712 VDD.n174 39.2114
R19869 VDD.n2710 VDD.n2709 39.2114
R19870 VDD.n2704 VDD.n179 39.2114
R19871 VDD.n2702 VDD.n2701 39.2114
R19872 VDD.n2430 VDD.n2429 39.2114
R19873 VDD.n2424 VDD.n2118 39.2114
R19874 VDD.n2421 VDD.n2119 39.2114
R19875 VDD.n2417 VDD.n2120 39.2114
R19876 VDD.n2413 VDD.n2121 39.2114
R19877 VDD.n2409 VDD.n2122 39.2114
R19878 VDD.n2404 VDD.n2123 39.2114
R19879 VDD.n2112 VDD.n439 39.2114
R19880 VDD.n2108 VDD.n438 39.2114
R19881 VDD.n2104 VDD.n437 39.2114
R19882 VDD.n2100 VDD.n436 39.2114
R19883 VDD.n2096 VDD.n435 39.2114
R19884 VDD.n2091 VDD.n434 39.2114
R19885 VDD.n2087 VDD.n433 39.2114
R19886 VDD.n1798 VDD.n1797 39.2114
R19887 VDD.n714 VDD.n700 39.2114
R19888 VDD.n1790 VDD.n701 39.2114
R19889 VDD.n1786 VDD.n702 39.2114
R19890 VDD.n1782 VDD.n703 39.2114
R19891 VDD.n1778 VDD.n704 39.2114
R19892 VDD.n1773 VDD.n705 39.2114
R19893 VDD.n2676 VDD.n2675 39.2114
R19894 VDD.n2671 VDD.n2668 39.2114
R19895 VDD.n2669 VDD.n150 39.2114
R19896 VDD.n2749 VDD.n2748 39.2114
R19897 VDD.n2746 VDD.n2745 39.2114
R19898 VDD.n2740 VDD.n157 39.2114
R19899 VDD.n2738 VDD.n2737 39.2114
R19900 VDD.n2433 VDD.n2432 39.2114
R19901 VDD.n2135 VDD.n2124 39.2114
R19902 VDD.n2139 VDD.n2125 39.2114
R19903 VDD.n2143 VDD.n2126 39.2114
R19904 VDD.n2147 VDD.n2127 39.2114
R19905 VDD.n2151 VDD.n2128 39.2114
R19906 VDD.n2155 VDD.n2129 39.2114
R19907 VDD.n2432 VDD.n423 39.2114
R19908 VDD.n2138 VDD.n2124 39.2114
R19909 VDD.n2142 VDD.n2125 39.2114
R19910 VDD.n2146 VDD.n2126 39.2114
R19911 VDD.n2150 VDD.n2127 39.2114
R19912 VDD.n2154 VDD.n2128 39.2114
R19913 VDD.n2130 VDD.n2129 39.2114
R19914 VDD.n2739 VDD.n2738 39.2114
R19915 VDD.n157 VDD.n153 39.2114
R19916 VDD.n2747 VDD.n2746 39.2114
R19917 VDD.n2750 VDD.n2749 39.2114
R19918 VDD.n2670 VDD.n2669 39.2114
R19919 VDD.n2668 VDD.n2666 39.2114
R19920 VDD.n2677 VDD.n2676 39.2114
R19921 VDD.n1797 VDD.n699 39.2114
R19922 VDD.n1791 VDD.n700 39.2114
R19923 VDD.n1787 VDD.n701 39.2114
R19924 VDD.n1783 VDD.n702 39.2114
R19925 VDD.n1779 VDD.n703 39.2114
R19926 VDD.n1774 VDD.n704 39.2114
R19927 VDD.n1770 VDD.n705 39.2114
R19928 VDD.n2090 VDD.n433 39.2114
R19929 VDD.n2095 VDD.n434 39.2114
R19930 VDD.n2099 VDD.n435 39.2114
R19931 VDD.n2103 VDD.n436 39.2114
R19932 VDD.n2107 VDD.n437 39.2114
R19933 VDD.n2111 VDD.n438 39.2114
R19934 VDD.n441 VDD.n439 39.2114
R19935 VDD.n2430 VDD.n2280 39.2114
R19936 VDD.n2422 VDD.n2118 39.2114
R19937 VDD.n2418 VDD.n2119 39.2114
R19938 VDD.n2414 VDD.n2120 39.2114
R19939 VDD.n2410 VDD.n2121 39.2114
R19940 VDD.n2405 VDD.n2122 39.2114
R19941 VDD.n2401 VDD.n2123 39.2114
R19942 VDD.n2703 VDD.n2702 39.2114
R19943 VDD.n179 VDD.n175 39.2114
R19944 VDD.n2711 VDD.n2710 39.2114
R19945 VDD.n174 VDD.n172 39.2114
R19946 VDD.n2719 VDD.n2718 39.2114
R19947 VDD.n171 VDD.n169 39.2114
R19948 VDD.n2726 VDD.n2725 39.2114
R19949 VDD.n2071 VDD.n425 39.2114
R19950 VDD.n2067 VDD.n426 39.2114
R19951 VDD.n2063 VDD.n427 39.2114
R19952 VDD.n2059 VDD.n428 39.2114
R19953 VDD.n2055 VDD.n429 39.2114
R19954 VDD.n2051 VDD.n430 39.2114
R19955 VDD.n2047 VDD.n431 39.2114
R19956 VDD.n769 VDD.n706 39.2114
R19957 VDD.n773 VDD.n707 39.2114
R19958 VDD.n777 VDD.n708 39.2114
R19959 VDD.n781 VDD.n709 39.2114
R19960 VDD.n913 VDD.n710 39.2114
R19961 VDD.n910 VDD.n711 39.2114
R19962 VDD.n906 VDD.n712 39.2114
R19963 VDD.n2044 VDD.n431 39.2114
R19964 VDD.n2048 VDD.n430 39.2114
R19965 VDD.n2052 VDD.n429 39.2114
R19966 VDD.n2056 VDD.n428 39.2114
R19967 VDD.n2060 VDD.n427 39.2114
R19968 VDD.n2064 VDD.n426 39.2114
R19969 VDD.n2068 VDD.n425 39.2114
R19970 VDD.n772 VDD.n706 39.2114
R19971 VDD.n776 VDD.n707 39.2114
R19972 VDD.n780 VDD.n708 39.2114
R19973 VDD.n783 VDD.n709 39.2114
R19974 VDD.n911 VDD.n710 39.2114
R19975 VDD.n907 VDD.n711 39.2114
R19976 VDD.n903 VDD.n712 39.2114
R19977 VDD.n1282 VDD.n1043 37.2369
R19978 VDD.n1060 VDD.n1059 37.2369
R19979 VDD.n1215 VDD.n1077 37.2369
R19980 VDD.n1181 VDD.n1094 37.2369
R19981 VDD.n1147 VDD.n1111 37.2369
R19982 VDD.n1533 VDD.n1511 37.2369
R19983 VDD.n1561 VDD.n957 37.2369
R19984 VDD.n927 VDD.n926 37.2369
R19985 VDD.n1605 VDD.n754 37.2369
R19986 VDD.n1630 VDD.n730 37.2369
R19987 VDD.n3034 VDD.n3033 37.2369
R19988 VDD.n3209 VDD.n3043 37.2369
R19989 VDD.n3175 VDD.n3051 37.2369
R19990 VDD.n3061 VDD.n3060 37.2369
R19991 VDD.n3105 VDD.n3070 37.2369
R19992 VDD.n2886 VDD.n115 37.2369
R19993 VDD.n2826 VDD.n141 37.2369
R19994 VDD.n2858 VDD.n2857 37.2369
R19995 VDD.n66 VDD.n65 37.2369
R19996 VDD.n2758 VDD.n2757 37.2369
R19997 VDD.n2115 VDD.n442 33.4054
R19998 VDD.n2088 VDD.n445 33.4054
R19999 VDD.n1771 VDD.n1768 33.4054
R20000 VDD.n1800 VDD.n1799 33.4054
R20001 VDD.n2402 VDD.n2399 33.4054
R20002 VDD.n2700 VDD.n2699 33.4054
R20003 VDD.n2428 VDD.n416 33.4054
R20004 VDD.n2729 VDD.n2728 33.4054
R20005 VDD.n2680 VDD.n2664 33.4054
R20006 VDD.n2736 VDD.n2735 33.4054
R20007 VDD.n2277 VDD.n2276 33.4054
R20008 VDD.n2435 VDD.n2434 33.4054
R20009 VDD.n770 VDD.n692 33.4054
R20010 VDD.n2073 VDD.n2070 33.4054
R20011 VDD.n2043 VDD.n2042 33.4054
R20012 VDD.n902 VDD.n901 33.4054
R20013 VDD.n786 VDD.n785 30.449
R20014 VDD.n462 VDD.n461 30.449
R20015 VDD.n1776 VDD.n1648 30.449
R20016 VDD.n2093 VDD.n444 30.449
R20017 VDD.n2134 VDD.n2133 30.449
R20018 VDD.n2706 VDD.n177 30.449
R20019 VDD.n2407 VDD.n2282 30.449
R20020 VDD.n2742 VDD.n155 30.449
R20021 VDD.n1288 VDD.n1038 24.3495
R20022 VDD.n1556 VDD.n721 24.3495
R20023 VDD.n2909 VDD.n60 24.3495
R20024 VDD.n3272 VDD.n3271 24.3495
R20025 VDD.n1286 VDD.n1030 19.3944
R20026 VDD.n1298 VDD.n1030 19.3944
R20027 VDD.n1298 VDD.n1028 19.3944
R20028 VDD.n1302 VDD.n1028 19.3944
R20029 VDD.n1302 VDD.n1019 19.3944
R20030 VDD.n1314 VDD.n1019 19.3944
R20031 VDD.n1314 VDD.n1017 19.3944
R20032 VDD.n1318 VDD.n1017 19.3944
R20033 VDD.n1318 VDD.n1007 19.3944
R20034 VDD.n1330 VDD.n1007 19.3944
R20035 VDD.n1330 VDD.n1005 19.3944
R20036 VDD.n1334 VDD.n1005 19.3944
R20037 VDD.n1334 VDD.n996 19.3944
R20038 VDD.n1446 VDD.n996 19.3944
R20039 VDD.n1446 VDD.n994 19.3944
R20040 VDD.n1450 VDD.n994 19.3944
R20041 VDD.n1450 VDD.n984 19.3944
R20042 VDD.n1462 VDD.n984 19.3944
R20043 VDD.n1462 VDD.n982 19.3944
R20044 VDD.n1466 VDD.n982 19.3944
R20045 VDD.n1466 VDD.n972 19.3944
R20046 VDD.n1478 VDD.n972 19.3944
R20047 VDD.n1478 VDD.n969 19.3944
R20048 VDD.n1485 VDD.n969 19.3944
R20049 VDD.n1485 VDD.n970 19.3944
R20050 VDD.n970 VDD.n959 19.3944
R20051 VDD.n1250 VDD.n1056 19.3944
R20052 VDD.n1256 VDD.n1056 19.3944
R20053 VDD.n1256 VDD.n1054 19.3944
R20054 VDD.n1260 VDD.n1054 19.3944
R20055 VDD.n1260 VDD.n1052 19.3944
R20056 VDD.n1266 VDD.n1052 19.3944
R20057 VDD.n1266 VDD.n1050 19.3944
R20058 VDD.n1270 VDD.n1050 19.3944
R20059 VDD.n1270 VDD.n1048 19.3944
R20060 VDD.n1277 VDD.n1048 19.3944
R20061 VDD.n1277 VDD.n1044 19.3944
R20062 VDD.n1281 VDD.n1044 19.3944
R20063 VDD.n1219 VDD.n1072 19.3944
R20064 VDD.n1219 VDD.n1070 19.3944
R20065 VDD.n1225 VDD.n1070 19.3944
R20066 VDD.n1225 VDD.n1068 19.3944
R20067 VDD.n1229 VDD.n1068 19.3944
R20068 VDD.n1229 VDD.n1066 19.3944
R20069 VDD.n1235 VDD.n1066 19.3944
R20070 VDD.n1235 VDD.n1064 19.3944
R20071 VDD.n1240 VDD.n1064 19.3944
R20072 VDD.n1240 VDD.n1062 19.3944
R20073 VDD.n1246 VDD.n1062 19.3944
R20074 VDD.n1247 VDD.n1246 19.3944
R20075 VDD.n1185 VDD.n1089 19.3944
R20076 VDD.n1185 VDD.n1087 19.3944
R20077 VDD.n1191 VDD.n1087 19.3944
R20078 VDD.n1191 VDD.n1085 19.3944
R20079 VDD.n1195 VDD.n1085 19.3944
R20080 VDD.n1195 VDD.n1083 19.3944
R20081 VDD.n1201 VDD.n1083 19.3944
R20082 VDD.n1201 VDD.n1081 19.3944
R20083 VDD.n1207 VDD.n1081 19.3944
R20084 VDD.n1207 VDD.n1079 19.3944
R20085 VDD.n1079 VDD.n1078 19.3944
R20086 VDD.n1214 VDD.n1078 19.3944
R20087 VDD.n1151 VDD.n1106 19.3944
R20088 VDD.n1151 VDD.n1104 19.3944
R20089 VDD.n1157 VDD.n1104 19.3944
R20090 VDD.n1157 VDD.n1102 19.3944
R20091 VDD.n1161 VDD.n1102 19.3944
R20092 VDD.n1161 VDD.n1100 19.3944
R20093 VDD.n1167 VDD.n1100 19.3944
R20094 VDD.n1167 VDD.n1098 19.3944
R20095 VDD.n1173 VDD.n1098 19.3944
R20096 VDD.n1173 VDD.n1096 19.3944
R20097 VDD.n1096 VDD.n1095 19.3944
R20098 VDD.n1180 VDD.n1095 19.3944
R20099 VDD.n1123 VDD.n1120 19.3944
R20100 VDD.n1123 VDD.n1119 19.3944
R20101 VDD.n1127 VDD.n1119 19.3944
R20102 VDD.n1127 VDD.n1117 19.3944
R20103 VDD.n1133 VDD.n1117 19.3944
R20104 VDD.n1133 VDD.n1115 19.3944
R20105 VDD.n1139 VDD.n1115 19.3944
R20106 VDD.n1139 VDD.n1113 19.3944
R20107 VDD.n1113 VDD.n1112 19.3944
R20108 VDD.n1146 VDD.n1112 19.3944
R20109 VDD.n1551 VDD.n1550 19.3944
R20110 VDD.n1550 VDD.n1549 19.3944
R20111 VDD.n1549 VDD.n1496 19.3944
R20112 VDD.n1497 VDD.n1496 19.3944
R20113 VDD.n1542 VDD.n1497 19.3944
R20114 VDD.n1542 VDD.n1541 19.3944
R20115 VDD.n1541 VDD.n1540 19.3944
R20116 VDD.n1540 VDD.n1504 19.3944
R20117 VDD.n1535 VDD.n1504 19.3944
R20118 VDD.n1535 VDD.n1534 19.3944
R20119 VDD.n1290 VDD.n1035 19.3944
R20120 VDD.n1294 VDD.n1035 19.3944
R20121 VDD.n1294 VDD.n1025 19.3944
R20122 VDD.n1306 VDD.n1025 19.3944
R20123 VDD.n1306 VDD.n1023 19.3944
R20124 VDD.n1310 VDD.n1023 19.3944
R20125 VDD.n1310 VDD.n1013 19.3944
R20126 VDD.n1322 VDD.n1013 19.3944
R20127 VDD.n1322 VDD.n1011 19.3944
R20128 VDD.n1326 VDD.n1011 19.3944
R20129 VDD.n1326 VDD.n1001 19.3944
R20130 VDD.n1338 VDD.n1001 19.3944
R20131 VDD.n1338 VDD.n999 19.3944
R20132 VDD.n1442 VDD.n999 19.3944
R20133 VDD.n1442 VDD.n990 19.3944
R20134 VDD.n1454 VDD.n990 19.3944
R20135 VDD.n1454 VDD.n988 19.3944
R20136 VDD.n1458 VDD.n988 19.3944
R20137 VDD.n1458 VDD.n978 19.3944
R20138 VDD.n1470 VDD.n978 19.3944
R20139 VDD.n1470 VDD.n976 19.3944
R20140 VDD.n1474 VDD.n976 19.3944
R20141 VDD.n1474 VDD.n965 19.3944
R20142 VDD.n1489 VDD.n965 19.3944
R20143 VDD.n1489 VDD.n963 19.3944
R20144 VDD.n1554 VDD.n963 19.3944
R20145 VDD.n1580 VDD.n1579 19.3944
R20146 VDD.n1579 VDD.n1578 19.3944
R20147 VDD.n1578 VDD.n934 19.3944
R20148 VDD.n1574 VDD.n934 19.3944
R20149 VDD.n1574 VDD.n1573 19.3944
R20150 VDD.n1573 VDD.n1572 19.3944
R20151 VDD.n1572 VDD.n942 19.3944
R20152 VDD.n1568 VDD.n942 19.3944
R20153 VDD.n1568 VDD.n1567 19.3944
R20154 VDD.n1567 VDD.n1566 19.3944
R20155 VDD.n1566 VDD.n950 19.3944
R20156 VDD.n1562 VDD.n950 19.3944
R20157 VDD.n1601 VDD.n752 19.3944
R20158 VDD.n1601 VDD.n758 19.3944
R20159 VDD.n1596 VDD.n758 19.3944
R20160 VDD.n1596 VDD.n1595 19.3944
R20161 VDD.n1595 VDD.n1594 19.3944
R20162 VDD.n1594 VDD.n765 19.3944
R20163 VDD.n1589 VDD.n768 19.3944
R20164 VDD.n1585 VDD.n918 19.3944
R20165 VDD.n1585 VDD.n1584 19.3944
R20166 VDD.n1584 VDD.n1583 19.3944
R20167 VDD.n1626 VDD.n728 19.3944
R20168 VDD.n1626 VDD.n733 19.3944
R20169 VDD.n1621 VDD.n733 19.3944
R20170 VDD.n1621 VDD.n1620 19.3944
R20171 VDD.n1620 VDD.n1619 19.3944
R20172 VDD.n1619 VDD.n739 19.3944
R20173 VDD.n1614 VDD.n739 19.3944
R20174 VDD.n1614 VDD.n1613 19.3944
R20175 VDD.n1613 VDD.n1612 19.3944
R20176 VDD.n1612 VDD.n746 19.3944
R20177 VDD.n1607 VDD.n746 19.3944
R20178 VDD.n1607 VDD.n1606 19.3944
R20179 VDD.n1532 VDD.n1516 19.3944
R20180 VDD.n1517 VDD.n1516 19.3944
R20181 VDD.n1525 VDD.n1517 19.3944
R20182 VDD.n1525 VDD.n1524 19.3944
R20183 VDD.n1524 VDD.n719 19.3944
R20184 VDD.n1644 VDD.n719 19.3944
R20185 VDD.n722 VDD.n718 19.3944
R20186 VDD.n1637 VDD.n1636 19.3944
R20187 VDD.n1636 VDD.n1635 19.3944
R20188 VDD.n1635 VDD.n725 19.3944
R20189 VDD.n2915 VDD.n62 19.3944
R20190 VDD.n2915 VDD.n52 19.3944
R20191 VDD.n2927 VDD.n52 19.3944
R20192 VDD.n2927 VDD.n50 19.3944
R20193 VDD.n2931 VDD.n50 19.3944
R20194 VDD.n2931 VDD.n40 19.3944
R20195 VDD.n2943 VDD.n40 19.3944
R20196 VDD.n2943 VDD.n38 19.3944
R20197 VDD.n2947 VDD.n38 19.3944
R20198 VDD.n2947 VDD.n28 19.3944
R20199 VDD.n2959 VDD.n28 19.3944
R20200 VDD.n2959 VDD.n26 19.3944
R20201 VDD.n3299 VDD.n26 19.3944
R20202 VDD.n3299 VDD.n3298 19.3944
R20203 VDD.n3298 VDD.n3297 19.3944
R20204 VDD.n3297 VDD.n2965 19.3944
R20205 VDD.n3250 VDD.n2965 19.3944
R20206 VDD.n3251 VDD.n3250 19.3944
R20207 VDD.n3251 VDD.n3247 19.3944
R20208 VDD.n3256 VDD.n3247 19.3944
R20209 VDD.n3257 VDD.n3256 19.3944
R20210 VDD.n3258 VDD.n3257 19.3944
R20211 VDD.n3258 VDD.n3245 19.3944
R20212 VDD.n3263 VDD.n3245 19.3944
R20213 VDD.n3264 VDD.n3263 19.3944
R20214 VDD.n3265 VDD.n3264 19.3944
R20215 VDD.n3212 VDD.n3040 19.3944
R20216 VDD.n3216 VDD.n3040 19.3944
R20217 VDD.n3219 VDD.n3216 19.3944
R20218 VDD.n3222 VDD.n3219 19.3944
R20219 VDD.n3222 VDD.n3038 19.3944
R20220 VDD.n3226 VDD.n3038 19.3944
R20221 VDD.n3229 VDD.n3226 19.3944
R20222 VDD.n3232 VDD.n3229 19.3944
R20223 VDD.n3232 VDD.n3036 19.3944
R20224 VDD.n3236 VDD.n3036 19.3944
R20225 VDD.n3239 VDD.n3236 19.3944
R20226 VDD.n3241 VDD.n3239 19.3944
R20227 VDD.n3181 VDD.n3178 19.3944
R20228 VDD.n3181 VDD.n3048 19.3944
R20229 VDD.n3185 VDD.n3048 19.3944
R20230 VDD.n3188 VDD.n3185 19.3944
R20231 VDD.n3191 VDD.n3188 19.3944
R20232 VDD.n3191 VDD.n3046 19.3944
R20233 VDD.n3195 VDD.n3046 19.3944
R20234 VDD.n3198 VDD.n3195 19.3944
R20235 VDD.n3201 VDD.n3198 19.3944
R20236 VDD.n3201 VDD.n3044 19.3944
R20237 VDD.n3205 VDD.n3044 19.3944
R20238 VDD.n3208 VDD.n3205 19.3944
R20239 VDD.n3145 VDD.n3144 19.3944
R20240 VDD.n3148 VDD.n3145 19.3944
R20241 VDD.n3148 VDD.n3057 19.3944
R20242 VDD.n3154 VDD.n3057 19.3944
R20243 VDD.n3155 VDD.n3154 19.3944
R20244 VDD.n3158 VDD.n3155 19.3944
R20245 VDD.n3158 VDD.n3055 19.3944
R20246 VDD.n3164 VDD.n3055 19.3944
R20247 VDD.n3165 VDD.n3164 19.3944
R20248 VDD.n3168 VDD.n3165 19.3944
R20249 VDD.n3168 VDD.n3053 19.3944
R20250 VDD.n3174 VDD.n3053 19.3944
R20251 VDD.n3108 VDD.n3067 19.3944
R20252 VDD.n3114 VDD.n3067 19.3944
R20253 VDD.n3115 VDD.n3114 19.3944
R20254 VDD.n3118 VDD.n3115 19.3944
R20255 VDD.n3118 VDD.n3065 19.3944
R20256 VDD.n3124 VDD.n3065 19.3944
R20257 VDD.n3125 VDD.n3124 19.3944
R20258 VDD.n3128 VDD.n3125 19.3944
R20259 VDD.n3128 VDD.n3063 19.3944
R20260 VDD.n3134 VDD.n3063 19.3944
R20261 VDD.n3135 VDD.n3134 19.3944
R20262 VDD.n3138 VDD.n3135 19.3944
R20263 VDD.n3078 VDD.n3075 19.3944
R20264 VDD.n3084 VDD.n3075 19.3944
R20265 VDD.n3085 VDD.n3084 19.3944
R20266 VDD.n3088 VDD.n3085 19.3944
R20267 VDD.n3088 VDD.n3073 19.3944
R20268 VDD.n3094 VDD.n3073 19.3944
R20269 VDD.n3095 VDD.n3094 19.3944
R20270 VDD.n3098 VDD.n3095 19.3944
R20271 VDD.n3098 VDD.n3071 19.3944
R20272 VDD.n3104 VDD.n3071 19.3944
R20273 VDD.n2919 VDD.n58 19.3944
R20274 VDD.n2919 VDD.n56 19.3944
R20275 VDD.n2923 VDD.n56 19.3944
R20276 VDD.n2923 VDD.n46 19.3944
R20277 VDD.n2935 VDD.n46 19.3944
R20278 VDD.n2935 VDD.n44 19.3944
R20279 VDD.n2939 VDD.n44 19.3944
R20280 VDD.n2939 VDD.n34 19.3944
R20281 VDD.n2951 VDD.n34 19.3944
R20282 VDD.n2951 VDD.n32 19.3944
R20283 VDD.n2955 VDD.n32 19.3944
R20284 VDD.n2955 VDD.n18 19.3944
R20285 VDD.n3302 VDD.n18 19.3944
R20286 VDD.n3302 VDD.n19 19.3944
R20287 VDD.n3293 VDD.n19 19.3944
R20288 VDD.n3293 VDD.n3292 19.3944
R20289 VDD.n3292 VDD.n3291 19.3944
R20290 VDD.n3291 VDD.n2972 19.3944
R20291 VDD.n3285 VDD.n2972 19.3944
R20292 VDD.n3285 VDD.n3284 19.3944
R20293 VDD.n3284 VDD.n3283 19.3944
R20294 VDD.n3283 VDD.n2983 19.3944
R20295 VDD.n3277 VDD.n2983 19.3944
R20296 VDD.n3277 VDD.n3276 19.3944
R20297 VDD.n3276 VDD.n3275 19.3944
R20298 VDD.n3275 VDD.n2994 19.3944
R20299 VDD.n2906 VDD.n2905 19.3944
R20300 VDD.n2905 VDD.n2904 19.3944
R20301 VDD.n2904 VDD.n2903 19.3944
R20302 VDD.n2903 VDD.n2901 19.3944
R20303 VDD.n2901 VDD.n2898 19.3944
R20304 VDD.n2898 VDD.n2897 19.3944
R20305 VDD.n2897 VDD.n2894 19.3944
R20306 VDD.n2894 VDD.n2893 19.3944
R20307 VDD.n2893 VDD.n2890 19.3944
R20308 VDD.n2890 VDD.n2889 19.3944
R20309 VDD.n2852 VDD.n127 19.3944
R20310 VDD.n2852 VDD.n2849 19.3944
R20311 VDD.n2849 VDD.n2846 19.3944
R20312 VDD.n2846 VDD.n2845 19.3944
R20313 VDD.n2845 VDD.n2842 19.3944
R20314 VDD.n2842 VDD.n2841 19.3944
R20315 VDD.n2841 VDD.n2838 19.3944
R20316 VDD.n2838 VDD.n2837 19.3944
R20317 VDD.n2837 VDD.n2834 19.3944
R20318 VDD.n2834 VDD.n2833 19.3944
R20319 VDD.n2833 VDD.n2830 19.3944
R20320 VDD.n2830 VDD.n2829 19.3944
R20321 VDD.n2885 VDD.n2882 19.3944
R20322 VDD.n2882 VDD.n2881 19.3944
R20323 VDD.n2881 VDD.n2878 19.3944
R20324 VDD.n2878 VDD.n2877 19.3944
R20325 VDD.n2877 VDD.n2874 19.3944
R20326 VDD.n2874 VDD.n2873 19.3944
R20327 VDD.n2870 VDD.n2869 19.3944
R20328 VDD.n2866 VDD.n2865 19.3944
R20329 VDD.n2865 VDD.n2862 19.3944
R20330 VDD.n2862 VDD.n2861 19.3944
R20331 VDD.n2796 VDD.n2795 19.3944
R20332 VDD.n2795 VDD.n2792 19.3944
R20333 VDD.n2792 VDD.n2791 19.3944
R20334 VDD.n2791 VDD.n2788 19.3944
R20335 VDD.n2788 VDD.n2787 19.3944
R20336 VDD.n2787 VDD.n2784 19.3944
R20337 VDD.n2784 VDD.n2783 19.3944
R20338 VDD.n2783 VDD.n2780 19.3944
R20339 VDD.n2780 VDD.n2779 19.3944
R20340 VDD.n2779 VDD.n2776 19.3944
R20341 VDD.n2776 VDD.n2775 19.3944
R20342 VDD.n2775 VDD.n2772 19.3944
R20343 VDD.n2822 VDD.n139 19.3944
R20344 VDD.n2822 VDD.n2819 19.3944
R20345 VDD.n2819 VDD.n2816 19.3944
R20346 VDD.n2816 VDD.n2815 19.3944
R20347 VDD.n2815 VDD.n2812 19.3944
R20348 VDD.n2812 VDD.n2811 19.3944
R20349 VDD.n2808 VDD.n2807 19.3944
R20350 VDD.n2804 VDD.n2803 19.3944
R20351 VDD.n2803 VDD.n2800 19.3944
R20352 VDD.n2800 VDD.n2799 19.3944
R20353 VDD.n1215 VDD.n1072 19.2005
R20354 VDD.n1147 VDD.n1146 19.2005
R20355 VDD.n1534 VDD.n1533 19.2005
R20356 VDD.n1605 VDD.n752 19.2005
R20357 VDD.n3178 VDD.n3175 19.2005
R20358 VDD.n3105 VDD.n3104 19.2005
R20359 VDD.n2889 VDD.n2886 19.2005
R20360 VDD.n2826 VDD.n139 19.2005
R20361 VDD.n1796 VDD.n694 17.188
R20362 VDD.n2117 VDD.n424 17.188
R20363 VDD.n2431 VDD.n418 17.188
R20364 VDD.n163 VDD.n151 17.188
R20365 VDD.n3390 VDD.n3388 16.3201
R20366 VDD.n3370 VDD.n3368 16.3201
R20367 VDD.n3350 VDD.n3348 16.3201
R20368 VDD.n3330 VDD.n3328 16.3201
R20369 VDD.n3311 VDD.n3309 16.3201
R20370 VDD.n1426 VDD.n1424 16.3201
R20371 VDD.n1406 VDD.n1404 16.3201
R20372 VDD.n1386 VDD.n1384 16.3201
R20373 VDD.n1366 VDD.n1364 16.3201
R20374 VDD.n1347 VDD.n1345 16.3201
R20375 VDD.n7 VDD.t112 14.3199
R20376 VDD.n7 VDD.t136 14.3199
R20377 VDD.n8 VDD.t131 14.3199
R20378 VDD.n8 VDD.t125 14.3199
R20379 VDD.n10 VDD.t106 14.3199
R20380 VDD.n10 VDD.t118 14.3199
R20381 VDD.n12 VDD.t116 14.3199
R20382 VDD.n12 VDD.t122 14.3199
R20383 VDD.n5 VDD.t114 14.3199
R20384 VDD.n5 VDD.t140 14.3199
R20385 VDD.n3 VDD.t101 14.3199
R20386 VDD.n3 VDD.t97 14.3199
R20387 VDD.n1 VDD.t108 14.3199
R20388 VDD.n1 VDD.t129 14.3199
R20389 VDD.n0 VDD.t95 14.3199
R20390 VDD.n0 VDD.t110 14.3199
R20391 VDD.n1282 VDD.n1281 13.7702
R20392 VDD.n1562 VDD.n1561 13.7702
R20393 VDD.n3241 VDD.n3034 13.7702
R20394 VDD.n2772 VDD.n66 13.7702
R20395 VDD.n1288 VDD.n1032 13.0213
R20396 VDD.n1296 VDD.n1032 13.0213
R20397 VDD.n1296 VDD.n1033 13.0213
R20398 VDD.n1304 VDD.n1021 13.0213
R20399 VDD.n1312 VDD.n1021 13.0213
R20400 VDD.n1312 VDD.n1015 13.0213
R20401 VDD.n1320 VDD.n1015 13.0213
R20402 VDD.n1320 VDD.n1009 13.0213
R20403 VDD.n1328 VDD.n1009 13.0213
R20404 VDD.n1328 VDD.n1003 13.0213
R20405 VDD.n1336 VDD.n1003 13.0213
R20406 VDD.n1336 VDD.t98 13.0213
R20407 VDD.n1444 VDD.t98 13.0213
R20408 VDD.n1444 VDD.n992 13.0213
R20409 VDD.n1452 VDD.n992 13.0213
R20410 VDD.n1452 VDD.n986 13.0213
R20411 VDD.n1460 VDD.n986 13.0213
R20412 VDD.n1460 VDD.n980 13.0213
R20413 VDD.n1468 VDD.n980 13.0213
R20414 VDD.n1468 VDD.n974 13.0213
R20415 VDD.n1476 VDD.n974 13.0213
R20416 VDD.n1487 VDD.n967 13.0213
R20417 VDD.n1487 VDD.n960 13.0213
R20418 VDD.n1556 VDD.n960 13.0213
R20419 VDD.n2917 VDD.n60 13.0213
R20420 VDD.n2917 VDD.n54 13.0213
R20421 VDD.n2925 VDD.n54 13.0213
R20422 VDD.n2933 VDD.n48 13.0213
R20423 VDD.n2933 VDD.n42 13.0213
R20424 VDD.n2941 VDD.n42 13.0213
R20425 VDD.n2941 VDD.n36 13.0213
R20426 VDD.n2949 VDD.n36 13.0213
R20427 VDD.n2949 VDD.n30 13.0213
R20428 VDD.n2957 VDD.n30 13.0213
R20429 VDD.n2957 VDD.n22 13.0213
R20430 VDD.t126 VDD.n22 13.0213
R20431 VDD.t126 VDD.n23 13.0213
R20432 VDD.n3295 VDD.n23 13.0213
R20433 VDD.n3295 VDD.n2967 13.0213
R20434 VDD.n3289 VDD.n2967 13.0213
R20435 VDD.n3289 VDD.n3288 13.0213
R20436 VDD.n3288 VDD.n3287 13.0213
R20437 VDD.n3287 VDD.n2977 13.0213
R20438 VDD.n3281 VDD.n2977 13.0213
R20439 VDD.n3281 VDD.n3280 13.0213
R20440 VDD.n3279 VDD.n2988 13.0213
R20441 VDD.n3273 VDD.n2988 13.0213
R20442 VDD.n3273 VDD.n3272 13.0213
R20443 VDD.n1181 VDD.n1089 12.9944
R20444 VDD.n1181 VDD.n1180 12.9944
R20445 VDD.n1630 VDD.n728 12.9944
R20446 VDD.n1630 VDD.n725 12.9944
R20447 VDD.n3144 VDD.n3061 12.9944
R20448 VDD.n3138 VDD.n3061 12.9944
R20449 VDD.n2858 VDD.n127 12.9944
R20450 VDD.n2861 VDD.n2858 12.9944
R20451 VDD.n3391 VDD.n3387 12.8005
R20452 VDD.n3371 VDD.n3367 12.8005
R20453 VDD.n3351 VDD.n3347 12.8005
R20454 VDD.n3331 VDD.n3327 12.8005
R20455 VDD.n3312 VDD.n3308 12.8005
R20456 VDD.n1427 VDD.n1423 12.8005
R20457 VDD.n1407 VDD.n1403 12.8005
R20458 VDD.n1387 VDD.n1383 12.8005
R20459 VDD.n1367 VDD.n1363 12.8005
R20460 VDD.n1348 VDD.n1344 12.8005
R20461 VDD.n1283 VDD.n1282 12.2187
R20462 VDD.n1561 VDD.n955 12.2187
R20463 VDD.n2911 VDD.n66 12.2187
R20464 VDD.n3268 VDD.n3034 12.2187
R20465 VDD.n3395 VDD.n3394 12.0247
R20466 VDD.n3375 VDD.n3374 12.0247
R20467 VDD.n3355 VDD.n3354 12.0247
R20468 VDD.n3335 VDD.n3334 12.0247
R20469 VDD.n3316 VDD.n3315 12.0247
R20470 VDD.n1431 VDD.n1430 12.0247
R20471 VDD.n1411 VDD.n1410 12.0247
R20472 VDD.n1391 VDD.n1390 12.0247
R20473 VDD.n1371 VDD.n1370 12.0247
R20474 VDD.n1352 VDD.n1351 12.0247
R20475 VDD.n1785 VDD.n1646 11.6152
R20476 VDD.n2715 VDD.n2714 11.6152
R20477 VDD.n2752 VDD.n2751 11.6152
R20478 VDD.n1587 VDD.n915 11.6152
R20479 VDD.n3398 VDD.n3385 11.249
R20480 VDD.n3378 VDD.n3365 11.249
R20481 VDD.n3358 VDD.n3345 11.249
R20482 VDD.n3338 VDD.n3325 11.249
R20483 VDD.n3319 VDD.n3306 11.249
R20484 VDD.n1434 VDD.n1421 11.249
R20485 VDD.n1414 VDD.n1401 11.249
R20486 VDD.n1394 VDD.n1381 11.249
R20487 VDD.n1374 VDD.n1361 11.249
R20488 VDD.n1355 VDD.n1342 11.249
R20489 VDD.n2115 VDD.n2114 10.6151
R20490 VDD.n2114 VDD.n2113 10.6151
R20491 VDD.n2113 VDD.n2110 10.6151
R20492 VDD.n2110 VDD.n2109 10.6151
R20493 VDD.n2109 VDD.n2106 10.6151
R20494 VDD.n2106 VDD.n2105 10.6151
R20495 VDD.n2105 VDD.n2102 10.6151
R20496 VDD.n2102 VDD.n2101 10.6151
R20497 VDD.n2101 VDD.n2098 10.6151
R20498 VDD.n2098 VDD.n2097 10.6151
R20499 VDD.n2097 VDD.n2094 10.6151
R20500 VDD.n2092 VDD.n2089 10.6151
R20501 VDD.n2089 VDD.n2088 10.6151
R20502 VDD.n1768 VDD.n1767 10.6151
R20503 VDD.n1767 VDD.n1766 10.6151
R20504 VDD.n1766 VDD.n1764 10.6151
R20505 VDD.n1764 VDD.n1763 10.6151
R20506 VDD.n1763 VDD.n1761 10.6151
R20507 VDD.n1761 VDD.n1760 10.6151
R20508 VDD.n1760 VDD.n1758 10.6151
R20509 VDD.n1758 VDD.n1757 10.6151
R20510 VDD.n1757 VDD.n1755 10.6151
R20511 VDD.n1755 VDD.n1754 10.6151
R20512 VDD.n1754 VDD.n1752 10.6151
R20513 VDD.n1752 VDD.n1751 10.6151
R20514 VDD.n1751 VDD.n1749 10.6151
R20515 VDD.n1749 VDD.n1748 10.6151
R20516 VDD.n1748 VDD.n1746 10.6151
R20517 VDD.n1746 VDD.n1745 10.6151
R20518 VDD.n1745 VDD.n1743 10.6151
R20519 VDD.n1743 VDD.n1742 10.6151
R20520 VDD.n1742 VDD.n1740 10.6151
R20521 VDD.n1740 VDD.n1739 10.6151
R20522 VDD.n1739 VDD.n1737 10.6151
R20523 VDD.n1737 VDD.n1736 10.6151
R20524 VDD.n1736 VDD.n1734 10.6151
R20525 VDD.n1734 VDD.n1733 10.6151
R20526 VDD.n1733 VDD.n1731 10.6151
R20527 VDD.n1731 VDD.n1730 10.6151
R20528 VDD.n1730 VDD.n1728 10.6151
R20529 VDD.n1728 VDD.n1727 10.6151
R20530 VDD.n1727 VDD.n1725 10.6151
R20531 VDD.n1725 VDD.n1724 10.6151
R20532 VDD.n1724 VDD.n1722 10.6151
R20533 VDD.n1722 VDD.n1721 10.6151
R20534 VDD.n1721 VDD.n1719 10.6151
R20535 VDD.n1719 VDD.n1718 10.6151
R20536 VDD.n1718 VDD.n1716 10.6151
R20537 VDD.n1716 VDD.n1715 10.6151
R20538 VDD.n1715 VDD.n1713 10.6151
R20539 VDD.n1713 VDD.n1712 10.6151
R20540 VDD.n1712 VDD.n1710 10.6151
R20541 VDD.n1710 VDD.n1709 10.6151
R20542 VDD.n1709 VDD.n1707 10.6151
R20543 VDD.n1707 VDD.n1706 10.6151
R20544 VDD.n1706 VDD.n1704 10.6151
R20545 VDD.n1704 VDD.n1703 10.6151
R20546 VDD.n1703 VDD.n1701 10.6151
R20547 VDD.n1701 VDD.n1700 10.6151
R20548 VDD.n1700 VDD.n1698 10.6151
R20549 VDD.n1698 VDD.n1697 10.6151
R20550 VDD.n1697 VDD.n1695 10.6151
R20551 VDD.n1695 VDD.n1694 10.6151
R20552 VDD.n1694 VDD.n1692 10.6151
R20553 VDD.n1692 VDD.n1691 10.6151
R20554 VDD.n1691 VDD.n1689 10.6151
R20555 VDD.n1689 VDD.n1688 10.6151
R20556 VDD.n1688 VDD.n1686 10.6151
R20557 VDD.n1686 VDD.n1685 10.6151
R20558 VDD.n1685 VDD.n1683 10.6151
R20559 VDD.n1683 VDD.n1682 10.6151
R20560 VDD.n1682 VDD.n1680 10.6151
R20561 VDD.n1680 VDD.n1679 10.6151
R20562 VDD.n1679 VDD.n1677 10.6151
R20563 VDD.n1677 VDD.n1676 10.6151
R20564 VDD.n1676 VDD.n1674 10.6151
R20565 VDD.n1674 VDD.n1673 10.6151
R20566 VDD.n1673 VDD.n1671 10.6151
R20567 VDD.n1671 VDD.n1670 10.6151
R20568 VDD.n1670 VDD.n1668 10.6151
R20569 VDD.n1668 VDD.n1667 10.6151
R20570 VDD.n1667 VDD.n1665 10.6151
R20571 VDD.n1665 VDD.n1664 10.6151
R20572 VDD.n1664 VDD.n1662 10.6151
R20573 VDD.n1662 VDD.n1661 10.6151
R20574 VDD.n1661 VDD.n1659 10.6151
R20575 VDD.n1659 VDD.n1658 10.6151
R20576 VDD.n1658 VDD.n1656 10.6151
R20577 VDD.n1656 VDD.n1655 10.6151
R20578 VDD.n1655 VDD.n1653 10.6151
R20579 VDD.n1653 VDD.n1652 10.6151
R20580 VDD.n1652 VDD.n1650 10.6151
R20581 VDD.n1650 VDD.n1649 10.6151
R20582 VDD.n1649 VDD.n447 10.6151
R20583 VDD.n447 VDD.n445 10.6151
R20584 VDD.n1799 VDD.n698 10.6151
R20585 VDD.n1794 VDD.n698 10.6151
R20586 VDD.n1794 VDD.n1793 10.6151
R20587 VDD.n1793 VDD.n1792 10.6151
R20588 VDD.n1792 VDD.n1789 10.6151
R20589 VDD.n1789 VDD.n1788 10.6151
R20590 VDD.n1788 VDD.n1785 10.6151
R20591 VDD.n1785 VDD.n1784 10.6151
R20592 VDD.n1784 VDD.n1781 10.6151
R20593 VDD.n1781 VDD.n1780 10.6151
R20594 VDD.n1780 VDD.n1777 10.6151
R20595 VDD.n1775 VDD.n1772 10.6151
R20596 VDD.n1772 VDD.n1771 10.6151
R20597 VDD.n1801 VDD.n1800 10.6151
R20598 VDD.n1801 VDD.n686 10.6151
R20599 VDD.n1811 VDD.n686 10.6151
R20600 VDD.n1812 VDD.n1811 10.6151
R20601 VDD.n1813 VDD.n1812 10.6151
R20602 VDD.n1813 VDD.n674 10.6151
R20603 VDD.n1823 VDD.n674 10.6151
R20604 VDD.n1824 VDD.n1823 10.6151
R20605 VDD.n1825 VDD.n1824 10.6151
R20606 VDD.n1825 VDD.n662 10.6151
R20607 VDD.n1835 VDD.n662 10.6151
R20608 VDD.n1836 VDD.n1835 10.6151
R20609 VDD.n1837 VDD.n1836 10.6151
R20610 VDD.n1837 VDD.n650 10.6151
R20611 VDD.n1847 VDD.n650 10.6151
R20612 VDD.n1848 VDD.n1847 10.6151
R20613 VDD.n1849 VDD.n1848 10.6151
R20614 VDD.n1849 VDD.n638 10.6151
R20615 VDD.n1859 VDD.n638 10.6151
R20616 VDD.n1860 VDD.n1859 10.6151
R20617 VDD.n1861 VDD.n1860 10.6151
R20618 VDD.n1861 VDD.n626 10.6151
R20619 VDD.n1871 VDD.n626 10.6151
R20620 VDD.n1872 VDD.n1871 10.6151
R20621 VDD.n1873 VDD.n1872 10.6151
R20622 VDD.n1873 VDD.n614 10.6151
R20623 VDD.n1883 VDD.n614 10.6151
R20624 VDD.n1884 VDD.n1883 10.6151
R20625 VDD.n1885 VDD.n1884 10.6151
R20626 VDD.n1885 VDD.n602 10.6151
R20627 VDD.n1895 VDD.n602 10.6151
R20628 VDD.n1896 VDD.n1895 10.6151
R20629 VDD.n1897 VDD.n1896 10.6151
R20630 VDD.n1897 VDD.n590 10.6151
R20631 VDD.n1907 VDD.n590 10.6151
R20632 VDD.n1908 VDD.n1907 10.6151
R20633 VDD.n1909 VDD.n1908 10.6151
R20634 VDD.n1909 VDD.n578 10.6151
R20635 VDD.n1919 VDD.n578 10.6151
R20636 VDD.n1920 VDD.n1919 10.6151
R20637 VDD.n1921 VDD.n1920 10.6151
R20638 VDD.n1921 VDD.n566 10.6151
R20639 VDD.n1931 VDD.n566 10.6151
R20640 VDD.n1932 VDD.n1931 10.6151
R20641 VDD.n1933 VDD.n1932 10.6151
R20642 VDD.n1933 VDD.n554 10.6151
R20643 VDD.n1943 VDD.n554 10.6151
R20644 VDD.n1944 VDD.n1943 10.6151
R20645 VDD.n1945 VDD.n1944 10.6151
R20646 VDD.n1945 VDD.n542 10.6151
R20647 VDD.n1955 VDD.n542 10.6151
R20648 VDD.n1956 VDD.n1955 10.6151
R20649 VDD.n1957 VDD.n1956 10.6151
R20650 VDD.n1957 VDD.n530 10.6151
R20651 VDD.n1967 VDD.n530 10.6151
R20652 VDD.n1968 VDD.n1967 10.6151
R20653 VDD.n1969 VDD.n1968 10.6151
R20654 VDD.n1969 VDD.n518 10.6151
R20655 VDD.n1979 VDD.n518 10.6151
R20656 VDD.n1980 VDD.n1979 10.6151
R20657 VDD.n1981 VDD.n1980 10.6151
R20658 VDD.n1981 VDD.n506 10.6151
R20659 VDD.n1991 VDD.n506 10.6151
R20660 VDD.n1992 VDD.n1991 10.6151
R20661 VDD.n1993 VDD.n1992 10.6151
R20662 VDD.n1993 VDD.n494 10.6151
R20663 VDD.n2003 VDD.n494 10.6151
R20664 VDD.n2004 VDD.n2003 10.6151
R20665 VDD.n2005 VDD.n2004 10.6151
R20666 VDD.n2005 VDD.n482 10.6151
R20667 VDD.n2015 VDD.n482 10.6151
R20668 VDD.n2016 VDD.n2015 10.6151
R20669 VDD.n2017 VDD.n2016 10.6151
R20670 VDD.n2017 VDD.n469 10.6151
R20671 VDD.n2029 VDD.n469 10.6151
R20672 VDD.n2030 VDD.n2029 10.6151
R20673 VDD.n2031 VDD.n2030 10.6151
R20674 VDD.n2031 VDD.n452 10.6151
R20675 VDD.n2080 VDD.n452 10.6151
R20676 VDD.n2081 VDD.n2080 10.6151
R20677 VDD.n2082 VDD.n2081 10.6151
R20678 VDD.n2082 VDD.n442 10.6151
R20679 VDD.n2399 VDD.n2398 10.6151
R20680 VDD.n2398 VDD.n2397 10.6151
R20681 VDD.n2397 VDD.n2395 10.6151
R20682 VDD.n2395 VDD.n2394 10.6151
R20683 VDD.n2394 VDD.n2392 10.6151
R20684 VDD.n2392 VDD.n2391 10.6151
R20685 VDD.n2391 VDD.n2389 10.6151
R20686 VDD.n2389 VDD.n2388 10.6151
R20687 VDD.n2388 VDD.n2386 10.6151
R20688 VDD.n2386 VDD.n2385 10.6151
R20689 VDD.n2385 VDD.n2383 10.6151
R20690 VDD.n2383 VDD.n2382 10.6151
R20691 VDD.n2382 VDD.n2380 10.6151
R20692 VDD.n2380 VDD.n2379 10.6151
R20693 VDD.n2379 VDD.n2377 10.6151
R20694 VDD.n2377 VDD.n2376 10.6151
R20695 VDD.n2376 VDD.n2374 10.6151
R20696 VDD.n2374 VDD.n2373 10.6151
R20697 VDD.n2373 VDD.n2371 10.6151
R20698 VDD.n2371 VDD.n2370 10.6151
R20699 VDD.n2370 VDD.n2368 10.6151
R20700 VDD.n2368 VDD.n2367 10.6151
R20701 VDD.n2367 VDD.n2365 10.6151
R20702 VDD.n2365 VDD.n2364 10.6151
R20703 VDD.n2364 VDD.n2362 10.6151
R20704 VDD.n2362 VDD.n2361 10.6151
R20705 VDD.n2361 VDD.n2359 10.6151
R20706 VDD.n2359 VDD.n2358 10.6151
R20707 VDD.n2358 VDD.n2356 10.6151
R20708 VDD.n2356 VDD.n2355 10.6151
R20709 VDD.n2355 VDD.n2353 10.6151
R20710 VDD.n2353 VDD.n2352 10.6151
R20711 VDD.n2352 VDD.n2350 10.6151
R20712 VDD.n2350 VDD.n2349 10.6151
R20713 VDD.n2349 VDD.n2347 10.6151
R20714 VDD.n2347 VDD.n2346 10.6151
R20715 VDD.n2346 VDD.n2344 10.6151
R20716 VDD.n2344 VDD.n2343 10.6151
R20717 VDD.n2343 VDD.n2341 10.6151
R20718 VDD.n2341 VDD.n2340 10.6151
R20719 VDD.n2340 VDD.n2338 10.6151
R20720 VDD.n2338 VDD.n2337 10.6151
R20721 VDD.n2337 VDD.n2335 10.6151
R20722 VDD.n2335 VDD.n2334 10.6151
R20723 VDD.n2334 VDD.n2332 10.6151
R20724 VDD.n2332 VDD.n2331 10.6151
R20725 VDD.n2331 VDD.n2329 10.6151
R20726 VDD.n2329 VDD.n2328 10.6151
R20727 VDD.n2328 VDD.n2326 10.6151
R20728 VDD.n2326 VDD.n2325 10.6151
R20729 VDD.n2325 VDD.n2323 10.6151
R20730 VDD.n2323 VDD.n2322 10.6151
R20731 VDD.n2322 VDD.n2320 10.6151
R20732 VDD.n2320 VDD.n2319 10.6151
R20733 VDD.n2319 VDD.n2317 10.6151
R20734 VDD.n2317 VDD.n2316 10.6151
R20735 VDD.n2316 VDD.n2314 10.6151
R20736 VDD.n2314 VDD.n2313 10.6151
R20737 VDD.n2313 VDD.n2311 10.6151
R20738 VDD.n2311 VDD.n2310 10.6151
R20739 VDD.n2310 VDD.n2308 10.6151
R20740 VDD.n2308 VDD.n2307 10.6151
R20741 VDD.n2307 VDD.n2305 10.6151
R20742 VDD.n2305 VDD.n2304 10.6151
R20743 VDD.n2304 VDD.n2302 10.6151
R20744 VDD.n2302 VDD.n2301 10.6151
R20745 VDD.n2301 VDD.n2299 10.6151
R20746 VDD.n2299 VDD.n2298 10.6151
R20747 VDD.n2298 VDD.n2296 10.6151
R20748 VDD.n2296 VDD.n2295 10.6151
R20749 VDD.n2295 VDD.n2293 10.6151
R20750 VDD.n2293 VDD.n2292 10.6151
R20751 VDD.n2292 VDD.n2290 10.6151
R20752 VDD.n2290 VDD.n2289 10.6151
R20753 VDD.n2289 VDD.n2287 10.6151
R20754 VDD.n2287 VDD.n2286 10.6151
R20755 VDD.n2286 VDD.n2284 10.6151
R20756 VDD.n2284 VDD.n2283 10.6151
R20757 VDD.n2283 VDD.n181 10.6151
R20758 VDD.n2697 VDD.n181 10.6151
R20759 VDD.n2698 VDD.n2697 10.6151
R20760 VDD.n2699 VDD.n2698 10.6151
R20761 VDD.n2428 VDD.n2427 10.6151
R20762 VDD.n2427 VDD.n2426 10.6151
R20763 VDD.n2426 VDD.n2425 10.6151
R20764 VDD.n2425 VDD.n2423 10.6151
R20765 VDD.n2423 VDD.n2420 10.6151
R20766 VDD.n2420 VDD.n2419 10.6151
R20767 VDD.n2419 VDD.n2416 10.6151
R20768 VDD.n2416 VDD.n2415 10.6151
R20769 VDD.n2415 VDD.n2412 10.6151
R20770 VDD.n2412 VDD.n2411 10.6151
R20771 VDD.n2411 VDD.n2408 10.6151
R20772 VDD.n2406 VDD.n2403 10.6151
R20773 VDD.n2403 VDD.n2402 10.6151
R20774 VDD.n2440 VDD.n416 10.6151
R20775 VDD.n2441 VDD.n2440 10.6151
R20776 VDD.n2442 VDD.n2441 10.6151
R20777 VDD.n2442 VDD.n404 10.6151
R20778 VDD.n2452 VDD.n404 10.6151
R20779 VDD.n2453 VDD.n2452 10.6151
R20780 VDD.n2454 VDD.n2453 10.6151
R20781 VDD.n2454 VDD.n391 10.6151
R20782 VDD.n2464 VDD.n391 10.6151
R20783 VDD.n2465 VDD.n2464 10.6151
R20784 VDD.n2466 VDD.n2465 10.6151
R20785 VDD.n2466 VDD.n380 10.6151
R20786 VDD.n2476 VDD.n380 10.6151
R20787 VDD.n2477 VDD.n2476 10.6151
R20788 VDD.n2478 VDD.n2477 10.6151
R20789 VDD.n2478 VDD.n368 10.6151
R20790 VDD.n2488 VDD.n368 10.6151
R20791 VDD.n2489 VDD.n2488 10.6151
R20792 VDD.n2490 VDD.n2489 10.6151
R20793 VDD.n2490 VDD.n356 10.6151
R20794 VDD.n2500 VDD.n356 10.6151
R20795 VDD.n2501 VDD.n2500 10.6151
R20796 VDD.n2502 VDD.n2501 10.6151
R20797 VDD.n2502 VDD.n344 10.6151
R20798 VDD.n2512 VDD.n344 10.6151
R20799 VDD.n2513 VDD.n2512 10.6151
R20800 VDD.n2514 VDD.n2513 10.6151
R20801 VDD.n2514 VDD.n331 10.6151
R20802 VDD.n2524 VDD.n331 10.6151
R20803 VDD.n2525 VDD.n2524 10.6151
R20804 VDD.n2526 VDD.n2525 10.6151
R20805 VDD.n2526 VDD.n320 10.6151
R20806 VDD.n2536 VDD.n320 10.6151
R20807 VDD.n2537 VDD.n2536 10.6151
R20808 VDD.n2538 VDD.n2537 10.6151
R20809 VDD.n2538 VDD.n308 10.6151
R20810 VDD.n2548 VDD.n308 10.6151
R20811 VDD.n2549 VDD.n2548 10.6151
R20812 VDD.n2550 VDD.n2549 10.6151
R20813 VDD.n2550 VDD.n296 10.6151
R20814 VDD.n2560 VDD.n296 10.6151
R20815 VDD.n2561 VDD.n2560 10.6151
R20816 VDD.n2562 VDD.n2561 10.6151
R20817 VDD.n2562 VDD.n284 10.6151
R20818 VDD.n2572 VDD.n284 10.6151
R20819 VDD.n2573 VDD.n2572 10.6151
R20820 VDD.n2574 VDD.n2573 10.6151
R20821 VDD.n2574 VDD.n271 10.6151
R20822 VDD.n2584 VDD.n271 10.6151
R20823 VDD.n2585 VDD.n2584 10.6151
R20824 VDD.n2586 VDD.n2585 10.6151
R20825 VDD.n2586 VDD.n260 10.6151
R20826 VDD.n2596 VDD.n260 10.6151
R20827 VDD.n2597 VDD.n2596 10.6151
R20828 VDD.n2598 VDD.n2597 10.6151
R20829 VDD.n2598 VDD.n248 10.6151
R20830 VDD.n2608 VDD.n248 10.6151
R20831 VDD.n2609 VDD.n2608 10.6151
R20832 VDD.n2610 VDD.n2609 10.6151
R20833 VDD.n2610 VDD.n236 10.6151
R20834 VDD.n2620 VDD.n236 10.6151
R20835 VDD.n2621 VDD.n2620 10.6151
R20836 VDD.n2622 VDD.n2621 10.6151
R20837 VDD.n2622 VDD.n224 10.6151
R20838 VDD.n2632 VDD.n224 10.6151
R20839 VDD.n2633 VDD.n2632 10.6151
R20840 VDD.n2634 VDD.n2633 10.6151
R20841 VDD.n2634 VDD.n212 10.6151
R20842 VDD.n2644 VDD.n212 10.6151
R20843 VDD.n2645 VDD.n2644 10.6151
R20844 VDD.n2646 VDD.n2645 10.6151
R20845 VDD.n2646 VDD.n200 10.6151
R20846 VDD.n2656 VDD.n200 10.6151
R20847 VDD.n2657 VDD.n2656 10.6151
R20848 VDD.n2658 VDD.n2657 10.6151
R20849 VDD.n2658 VDD.n187 10.6151
R20850 VDD.n2690 VDD.n187 10.6151
R20851 VDD.n2691 VDD.n2690 10.6151
R20852 VDD.n2692 VDD.n2691 10.6151
R20853 VDD.n2692 VDD.n167 10.6151
R20854 VDD.n2730 VDD.n167 10.6151
R20855 VDD.n2730 VDD.n2729 10.6151
R20856 VDD.n2728 VDD.n168 10.6151
R20857 VDD.n2723 VDD.n168 10.6151
R20858 VDD.n2723 VDD.n2722 10.6151
R20859 VDD.n2722 VDD.n2721 10.6151
R20860 VDD.n2721 VDD.n170 10.6151
R20861 VDD.n2716 VDD.n170 10.6151
R20862 VDD.n2716 VDD.n2715 10.6151
R20863 VDD.n2715 VDD.n2713 10.6151
R20864 VDD.n2713 VDD.n173 10.6151
R20865 VDD.n2708 VDD.n173 10.6151
R20866 VDD.n2708 VDD.n2707 10.6151
R20867 VDD.n2705 VDD.n178 10.6151
R20868 VDD.n2700 VDD.n178 10.6151
R20869 VDD.n2665 VDD.n2664 10.6151
R20870 VDD.n2674 VDD.n2665 10.6151
R20871 VDD.n2674 VDD.n2673 10.6151
R20872 VDD.n2673 VDD.n2672 10.6151
R20873 VDD.n2672 VDD.n2667 10.6151
R20874 VDD.n2667 VDD.n148 10.6151
R20875 VDD.n2751 VDD.n148 10.6151
R20876 VDD.n2751 VDD.n149 10.6151
R20877 VDD.n152 VDD.n149 10.6151
R20878 VDD.n2744 VDD.n152 10.6151
R20879 VDD.n2744 VDD.n2743 10.6151
R20880 VDD.n2741 VDD.n156 10.6151
R20881 VDD.n2736 VDD.n156 10.6151
R20882 VDD.n2276 VDD.n2275 10.6151
R20883 VDD.n2275 VDD.n2274 10.6151
R20884 VDD.n2274 VDD.n2272 10.6151
R20885 VDD.n2272 VDD.n2271 10.6151
R20886 VDD.n2271 VDD.n2269 10.6151
R20887 VDD.n2269 VDD.n2268 10.6151
R20888 VDD.n2268 VDD.n2266 10.6151
R20889 VDD.n2266 VDD.n2265 10.6151
R20890 VDD.n2265 VDD.n2263 10.6151
R20891 VDD.n2263 VDD.n2262 10.6151
R20892 VDD.n2262 VDD.n2260 10.6151
R20893 VDD.n2260 VDD.n2259 10.6151
R20894 VDD.n2259 VDD.n2257 10.6151
R20895 VDD.n2257 VDD.n2256 10.6151
R20896 VDD.n2256 VDD.n2254 10.6151
R20897 VDD.n2254 VDD.n2253 10.6151
R20898 VDD.n2253 VDD.n2251 10.6151
R20899 VDD.n2251 VDD.n2250 10.6151
R20900 VDD.n2250 VDD.n2248 10.6151
R20901 VDD.n2248 VDD.n2247 10.6151
R20902 VDD.n2247 VDD.n2245 10.6151
R20903 VDD.n2245 VDD.n2244 10.6151
R20904 VDD.n2244 VDD.n2242 10.6151
R20905 VDD.n2242 VDD.n2241 10.6151
R20906 VDD.n2241 VDD.n2239 10.6151
R20907 VDD.n2239 VDD.n2238 10.6151
R20908 VDD.n2238 VDD.n2236 10.6151
R20909 VDD.n2236 VDD.n2235 10.6151
R20910 VDD.n2235 VDD.n2233 10.6151
R20911 VDD.n2233 VDD.n2232 10.6151
R20912 VDD.n2232 VDD.n2230 10.6151
R20913 VDD.n2230 VDD.n2229 10.6151
R20914 VDD.n2229 VDD.n2227 10.6151
R20915 VDD.n2227 VDD.n2226 10.6151
R20916 VDD.n2226 VDD.n2224 10.6151
R20917 VDD.n2224 VDD.n2223 10.6151
R20918 VDD.n2223 VDD.n2221 10.6151
R20919 VDD.n2221 VDD.n2220 10.6151
R20920 VDD.n2220 VDD.n2218 10.6151
R20921 VDD.n2218 VDD.n2217 10.6151
R20922 VDD.n2217 VDD.n2215 10.6151
R20923 VDD.n2215 VDD.n2214 10.6151
R20924 VDD.n2214 VDD.n2212 10.6151
R20925 VDD.n2212 VDD.n2211 10.6151
R20926 VDD.n2211 VDD.n2209 10.6151
R20927 VDD.n2209 VDD.n2208 10.6151
R20928 VDD.n2208 VDD.n2206 10.6151
R20929 VDD.n2206 VDD.n2205 10.6151
R20930 VDD.n2205 VDD.n2203 10.6151
R20931 VDD.n2203 VDD.n2202 10.6151
R20932 VDD.n2202 VDD.n2200 10.6151
R20933 VDD.n2200 VDD.n2199 10.6151
R20934 VDD.n2199 VDD.n2197 10.6151
R20935 VDD.n2197 VDD.n2196 10.6151
R20936 VDD.n2196 VDD.n2194 10.6151
R20937 VDD.n2194 VDD.n2193 10.6151
R20938 VDD.n2193 VDD.n2191 10.6151
R20939 VDD.n2191 VDD.n2190 10.6151
R20940 VDD.n2190 VDD.n2188 10.6151
R20941 VDD.n2188 VDD.n2187 10.6151
R20942 VDD.n2187 VDD.n2185 10.6151
R20943 VDD.n2185 VDD.n2184 10.6151
R20944 VDD.n2184 VDD.n2182 10.6151
R20945 VDD.n2182 VDD.n2181 10.6151
R20946 VDD.n2181 VDD.n2179 10.6151
R20947 VDD.n2179 VDD.n2178 10.6151
R20948 VDD.n2178 VDD.n2176 10.6151
R20949 VDD.n2176 VDD.n2175 10.6151
R20950 VDD.n2175 VDD.n2173 10.6151
R20951 VDD.n2173 VDD.n2172 10.6151
R20952 VDD.n2172 VDD.n2170 10.6151
R20953 VDD.n2170 VDD.n2169 10.6151
R20954 VDD.n2169 VDD.n2167 10.6151
R20955 VDD.n2167 VDD.n2166 10.6151
R20956 VDD.n2166 VDD.n2164 10.6151
R20957 VDD.n2164 VDD.n2163 10.6151
R20958 VDD.n2163 VDD.n2161 10.6151
R20959 VDD.n2161 VDD.n2160 10.6151
R20960 VDD.n2160 VDD.n2158 10.6151
R20961 VDD.n2158 VDD.n159 10.6151
R20962 VDD.n2734 VDD.n159 10.6151
R20963 VDD.n2735 VDD.n2734 10.6151
R20964 VDD.n2434 VDD.n422 10.6151
R20965 VDD.n2136 VDD.n422 10.6151
R20966 VDD.n2137 VDD.n2136 10.6151
R20967 VDD.n2140 VDD.n2137 10.6151
R20968 VDD.n2141 VDD.n2140 10.6151
R20969 VDD.n2144 VDD.n2141 10.6151
R20970 VDD.n2145 VDD.n2144 10.6151
R20971 VDD.n2148 VDD.n2145 10.6151
R20972 VDD.n2149 VDD.n2148 10.6151
R20973 VDD.n2152 VDD.n2149 10.6151
R20974 VDD.n2153 VDD.n2152 10.6151
R20975 VDD.n2157 VDD.n2156 10.6151
R20976 VDD.n2277 VDD.n2157 10.6151
R20977 VDD.n2436 VDD.n2435 10.6151
R20978 VDD.n2436 VDD.n410 10.6151
R20979 VDD.n2446 VDD.n410 10.6151
R20980 VDD.n2447 VDD.n2446 10.6151
R20981 VDD.n2448 VDD.n2447 10.6151
R20982 VDD.n2448 VDD.n398 10.6151
R20983 VDD.n2458 VDD.n398 10.6151
R20984 VDD.n2459 VDD.n2458 10.6151
R20985 VDD.n2460 VDD.n2459 10.6151
R20986 VDD.n2460 VDD.n385 10.6151
R20987 VDD.n2470 VDD.n385 10.6151
R20988 VDD.n2471 VDD.n2470 10.6151
R20989 VDD.n2472 VDD.n2471 10.6151
R20990 VDD.n2472 VDD.n374 10.6151
R20991 VDD.n2482 VDD.n374 10.6151
R20992 VDD.n2483 VDD.n2482 10.6151
R20993 VDD.n2484 VDD.n2483 10.6151
R20994 VDD.n2484 VDD.n362 10.6151
R20995 VDD.n2494 VDD.n362 10.6151
R20996 VDD.n2495 VDD.n2494 10.6151
R20997 VDD.n2496 VDD.n2495 10.6151
R20998 VDD.n2496 VDD.n350 10.6151
R20999 VDD.n2506 VDD.n350 10.6151
R21000 VDD.n2507 VDD.n2506 10.6151
R21001 VDD.n2508 VDD.n2507 10.6151
R21002 VDD.n2508 VDD.n338 10.6151
R21003 VDD.n2518 VDD.n338 10.6151
R21004 VDD.n2519 VDD.n2518 10.6151
R21005 VDD.n2520 VDD.n2519 10.6151
R21006 VDD.n2520 VDD.n326 10.6151
R21007 VDD.n2530 VDD.n326 10.6151
R21008 VDD.n2531 VDD.n2530 10.6151
R21009 VDD.n2532 VDD.n2531 10.6151
R21010 VDD.n2532 VDD.n314 10.6151
R21011 VDD.n2542 VDD.n314 10.6151
R21012 VDD.n2543 VDD.n2542 10.6151
R21013 VDD.n2544 VDD.n2543 10.6151
R21014 VDD.n2544 VDD.n302 10.6151
R21015 VDD.n2554 VDD.n302 10.6151
R21016 VDD.n2555 VDD.n2554 10.6151
R21017 VDD.n2556 VDD.n2555 10.6151
R21018 VDD.n2556 VDD.n290 10.6151
R21019 VDD.n2566 VDD.n290 10.6151
R21020 VDD.n2567 VDD.n2566 10.6151
R21021 VDD.n2568 VDD.n2567 10.6151
R21022 VDD.n2568 VDD.n277 10.6151
R21023 VDD.n2578 VDD.n277 10.6151
R21024 VDD.n2579 VDD.n2578 10.6151
R21025 VDD.n2580 VDD.n2579 10.6151
R21026 VDD.n2580 VDD.n266 10.6151
R21027 VDD.n2590 VDD.n266 10.6151
R21028 VDD.n2591 VDD.n2590 10.6151
R21029 VDD.n2592 VDD.n2591 10.6151
R21030 VDD.n2592 VDD.n254 10.6151
R21031 VDD.n2602 VDD.n254 10.6151
R21032 VDD.n2603 VDD.n2602 10.6151
R21033 VDD.n2604 VDD.n2603 10.6151
R21034 VDD.n2604 VDD.n242 10.6151
R21035 VDD.n2614 VDD.n242 10.6151
R21036 VDD.n2615 VDD.n2614 10.6151
R21037 VDD.n2616 VDD.n2615 10.6151
R21038 VDD.n2616 VDD.n230 10.6151
R21039 VDD.n2626 VDD.n230 10.6151
R21040 VDD.n2627 VDD.n2626 10.6151
R21041 VDD.n2628 VDD.n2627 10.6151
R21042 VDD.n2628 VDD.n218 10.6151
R21043 VDD.n2638 VDD.n218 10.6151
R21044 VDD.n2639 VDD.n2638 10.6151
R21045 VDD.n2640 VDD.n2639 10.6151
R21046 VDD.n2640 VDD.n206 10.6151
R21047 VDD.n2650 VDD.n206 10.6151
R21048 VDD.n2651 VDD.n2650 10.6151
R21049 VDD.n2652 VDD.n2651 10.6151
R21050 VDD.n2652 VDD.n194 10.6151
R21051 VDD.n2662 VDD.n194 10.6151
R21052 VDD.n2663 VDD.n2662 10.6151
R21053 VDD.n2686 VDD.n2663 10.6151
R21054 VDD.n2686 VDD.n2685 10.6151
R21055 VDD.n2685 VDD.n2684 10.6151
R21056 VDD.n2684 VDD.n2683 10.6151
R21057 VDD.n2683 VDD.n2681 10.6151
R21058 VDD.n2681 VDD.n2680 10.6151
R21059 VDD.n1805 VDD.n692 10.6151
R21060 VDD.n1806 VDD.n1805 10.6151
R21061 VDD.n1807 VDD.n1806 10.6151
R21062 VDD.n1807 VDD.n680 10.6151
R21063 VDD.n1817 VDD.n680 10.6151
R21064 VDD.n1818 VDD.n1817 10.6151
R21065 VDD.n1819 VDD.n1818 10.6151
R21066 VDD.n1819 VDD.n667 10.6151
R21067 VDD.n1829 VDD.n667 10.6151
R21068 VDD.n1830 VDD.n1829 10.6151
R21069 VDD.n1831 VDD.n1830 10.6151
R21070 VDD.n1831 VDD.n655 10.6151
R21071 VDD.n1841 VDD.n655 10.6151
R21072 VDD.n1842 VDD.n1841 10.6151
R21073 VDD.n1843 VDD.n1842 10.6151
R21074 VDD.n1843 VDD.n644 10.6151
R21075 VDD.n1853 VDD.n644 10.6151
R21076 VDD.n1854 VDD.n1853 10.6151
R21077 VDD.n1855 VDD.n1854 10.6151
R21078 VDD.n1855 VDD.n632 10.6151
R21079 VDD.n1865 VDD.n632 10.6151
R21080 VDD.n1866 VDD.n1865 10.6151
R21081 VDD.n1867 VDD.n1866 10.6151
R21082 VDD.n1867 VDD.n620 10.6151
R21083 VDD.n1877 VDD.n620 10.6151
R21084 VDD.n1878 VDD.n1877 10.6151
R21085 VDD.n1879 VDD.n1878 10.6151
R21086 VDD.n1879 VDD.n608 10.6151
R21087 VDD.n1889 VDD.n608 10.6151
R21088 VDD.n1890 VDD.n1889 10.6151
R21089 VDD.n1891 VDD.n1890 10.6151
R21090 VDD.n1891 VDD.n596 10.6151
R21091 VDD.n1901 VDD.n596 10.6151
R21092 VDD.n1902 VDD.n1901 10.6151
R21093 VDD.n1903 VDD.n1902 10.6151
R21094 VDD.n1903 VDD.n584 10.6151
R21095 VDD.n1913 VDD.n584 10.6151
R21096 VDD.n1914 VDD.n1913 10.6151
R21097 VDD.n1915 VDD.n1914 10.6151
R21098 VDD.n1915 VDD.n572 10.6151
R21099 VDD.n1925 VDD.n572 10.6151
R21100 VDD.n1926 VDD.n1925 10.6151
R21101 VDD.n1927 VDD.n1926 10.6151
R21102 VDD.n1927 VDD.n560 10.6151
R21103 VDD.n1937 VDD.n560 10.6151
R21104 VDD.n1938 VDD.n1937 10.6151
R21105 VDD.n1939 VDD.n1938 10.6151
R21106 VDD.n1939 VDD.n547 10.6151
R21107 VDD.n1949 VDD.n547 10.6151
R21108 VDD.n1950 VDD.n1949 10.6151
R21109 VDD.n1951 VDD.n1950 10.6151
R21110 VDD.n1951 VDD.n536 10.6151
R21111 VDD.n1961 VDD.n536 10.6151
R21112 VDD.n1962 VDD.n1961 10.6151
R21113 VDD.n1963 VDD.n1962 10.6151
R21114 VDD.n1963 VDD.n524 10.6151
R21115 VDD.n1973 VDD.n524 10.6151
R21116 VDD.n1974 VDD.n1973 10.6151
R21117 VDD.n1975 VDD.n1974 10.6151
R21118 VDD.n1975 VDD.n512 10.6151
R21119 VDD.n1985 VDD.n512 10.6151
R21120 VDD.n1986 VDD.n1985 10.6151
R21121 VDD.n1987 VDD.n1986 10.6151
R21122 VDD.n1987 VDD.n500 10.6151
R21123 VDD.n1997 VDD.n500 10.6151
R21124 VDD.n1998 VDD.n1997 10.6151
R21125 VDD.n1999 VDD.n1998 10.6151
R21126 VDD.n1999 VDD.n488 10.6151
R21127 VDD.n2009 VDD.n488 10.6151
R21128 VDD.n2010 VDD.n2009 10.6151
R21129 VDD.n2011 VDD.n2010 10.6151
R21130 VDD.n2011 VDD.n476 10.6151
R21131 VDD.n2021 VDD.n476 10.6151
R21132 VDD.n2022 VDD.n2021 10.6151
R21133 VDD.n2025 VDD.n2022 10.6151
R21134 VDD.n2025 VDD.n2024 10.6151
R21135 VDD.n2024 VDD.n2023 10.6151
R21136 VDD.n2023 VDD.n459 10.6151
R21137 VDD.n2076 VDD.n459 10.6151
R21138 VDD.n2076 VDD.n2075 10.6151
R21139 VDD.n2075 VDD.n2074 10.6151
R21140 VDD.n2074 VDD.n2073 10.6151
R21141 VDD.n2070 VDD.n2069 10.6151
R21142 VDD.n2069 VDD.n2066 10.6151
R21143 VDD.n2066 VDD.n2065 10.6151
R21144 VDD.n2065 VDD.n2062 10.6151
R21145 VDD.n2062 VDD.n2061 10.6151
R21146 VDD.n2061 VDD.n2058 10.6151
R21147 VDD.n2058 VDD.n2057 10.6151
R21148 VDD.n2057 VDD.n2054 10.6151
R21149 VDD.n2054 VDD.n2053 10.6151
R21150 VDD.n2053 VDD.n2050 10.6151
R21151 VDD.n2050 VDD.n2049 10.6151
R21152 VDD.n2046 VDD.n2045 10.6151
R21153 VDD.n2045 VDD.n2043 10.6151
R21154 VDD.n901 VDD.n899 10.6151
R21155 VDD.n899 VDD.n898 10.6151
R21156 VDD.n898 VDD.n896 10.6151
R21157 VDD.n896 VDD.n895 10.6151
R21158 VDD.n895 VDD.n893 10.6151
R21159 VDD.n893 VDD.n892 10.6151
R21160 VDD.n892 VDD.n890 10.6151
R21161 VDD.n890 VDD.n889 10.6151
R21162 VDD.n889 VDD.n887 10.6151
R21163 VDD.n887 VDD.n886 10.6151
R21164 VDD.n886 VDD.n884 10.6151
R21165 VDD.n884 VDD.n883 10.6151
R21166 VDD.n883 VDD.n881 10.6151
R21167 VDD.n881 VDD.n880 10.6151
R21168 VDD.n880 VDD.n878 10.6151
R21169 VDD.n878 VDD.n877 10.6151
R21170 VDD.n877 VDD.n875 10.6151
R21171 VDD.n875 VDD.n874 10.6151
R21172 VDD.n874 VDD.n872 10.6151
R21173 VDD.n872 VDD.n871 10.6151
R21174 VDD.n871 VDD.n869 10.6151
R21175 VDD.n869 VDD.n868 10.6151
R21176 VDD.n868 VDD.n866 10.6151
R21177 VDD.n866 VDD.n865 10.6151
R21178 VDD.n865 VDD.n863 10.6151
R21179 VDD.n863 VDD.n862 10.6151
R21180 VDD.n862 VDD.n860 10.6151
R21181 VDD.n860 VDD.n859 10.6151
R21182 VDD.n859 VDD.n857 10.6151
R21183 VDD.n857 VDD.n856 10.6151
R21184 VDD.n856 VDD.n854 10.6151
R21185 VDD.n854 VDD.n853 10.6151
R21186 VDD.n853 VDD.n851 10.6151
R21187 VDD.n851 VDD.n850 10.6151
R21188 VDD.n850 VDD.n848 10.6151
R21189 VDD.n848 VDD.n847 10.6151
R21190 VDD.n847 VDD.n845 10.6151
R21191 VDD.n845 VDD.n844 10.6151
R21192 VDD.n844 VDD.n842 10.6151
R21193 VDD.n842 VDD.n841 10.6151
R21194 VDD.n841 VDD.n839 10.6151
R21195 VDD.n839 VDD.n838 10.6151
R21196 VDD.n838 VDD.n836 10.6151
R21197 VDD.n836 VDD.n835 10.6151
R21198 VDD.n835 VDD.n833 10.6151
R21199 VDD.n833 VDD.n832 10.6151
R21200 VDD.n832 VDD.n830 10.6151
R21201 VDD.n830 VDD.n829 10.6151
R21202 VDD.n829 VDD.n827 10.6151
R21203 VDD.n827 VDD.n826 10.6151
R21204 VDD.n826 VDD.n824 10.6151
R21205 VDD.n824 VDD.n823 10.6151
R21206 VDD.n823 VDD.n821 10.6151
R21207 VDD.n821 VDD.n820 10.6151
R21208 VDD.n820 VDD.n818 10.6151
R21209 VDD.n818 VDD.n817 10.6151
R21210 VDD.n817 VDD.n815 10.6151
R21211 VDD.n815 VDD.n814 10.6151
R21212 VDD.n814 VDD.n812 10.6151
R21213 VDD.n812 VDD.n811 10.6151
R21214 VDD.n811 VDD.n809 10.6151
R21215 VDD.n809 VDD.n808 10.6151
R21216 VDD.n808 VDD.n806 10.6151
R21217 VDD.n806 VDD.n805 10.6151
R21218 VDD.n805 VDD.n803 10.6151
R21219 VDD.n803 VDD.n802 10.6151
R21220 VDD.n802 VDD.n800 10.6151
R21221 VDD.n800 VDD.n799 10.6151
R21222 VDD.n799 VDD.n797 10.6151
R21223 VDD.n797 VDD.n796 10.6151
R21224 VDD.n796 VDD.n794 10.6151
R21225 VDD.n794 VDD.n793 10.6151
R21226 VDD.n793 VDD.n791 10.6151
R21227 VDD.n791 VDD.n790 10.6151
R21228 VDD.n790 VDD.n788 10.6151
R21229 VDD.n788 VDD.n787 10.6151
R21230 VDD.n787 VDD.n463 10.6151
R21231 VDD.n2036 VDD.n463 10.6151
R21232 VDD.n2037 VDD.n2036 10.6151
R21233 VDD.n2039 VDD.n2037 10.6151
R21234 VDD.n2040 VDD.n2039 10.6151
R21235 VDD.n2042 VDD.n2040 10.6151
R21236 VDD.n771 VDD.n770 10.6151
R21237 VDD.n774 VDD.n771 10.6151
R21238 VDD.n775 VDD.n774 10.6151
R21239 VDD.n778 VDD.n775 10.6151
R21240 VDD.n779 VDD.n778 10.6151
R21241 VDD.n782 VDD.n779 10.6151
R21242 VDD.n915 VDD.n782 10.6151
R21243 VDD.n915 VDD.n914 10.6151
R21244 VDD.n914 VDD.n912 10.6151
R21245 VDD.n912 VDD.n909 10.6151
R21246 VDD.n909 VDD.n908 10.6151
R21247 VDD.n905 VDD.n904 10.6151
R21248 VDD.n904 VDD.n902 10.6151
R21249 VDD.n3399 VDD.n3383 10.4732
R21250 VDD.n3379 VDD.n3363 10.4732
R21251 VDD.n3359 VDD.n3343 10.4732
R21252 VDD.n3339 VDD.n3323 10.4732
R21253 VDD.n3320 VDD.n3304 10.4732
R21254 VDD.n1435 VDD.n1419 10.4732
R21255 VDD.n1415 VDD.n1399 10.4732
R21256 VDD.n1395 VDD.n1379 10.4732
R21257 VDD.n1375 VDD.n1359 10.4732
R21258 VDD.n1356 VDD.n1340 10.4732
R21259 VDD.n3401 VDD.n3400 9.45567
R21260 VDD.n3381 VDD.n3380 9.45567
R21261 VDD.n3361 VDD.n3360 9.45567
R21262 VDD.n3341 VDD.n3340 9.45567
R21263 VDD.n3322 VDD.n3321 9.45567
R21264 VDD.n1437 VDD.n1436 9.45567
R21265 VDD.n1417 VDD.n1416 9.45567
R21266 VDD.n1397 VDD.n1396 9.45567
R21267 VDD.n1377 VDD.n1376 9.45567
R21268 VDD.n1358 VDD.n1357 9.45567
R21269 VDD.n1442 VDD.n1441 9.3005
R21270 VDD.n990 VDD.n989 9.3005
R21271 VDD.n1455 VDD.n1454 9.3005
R21272 VDD.n1456 VDD.n988 9.3005
R21273 VDD.n1458 VDD.n1457 9.3005
R21274 VDD.n978 VDD.n977 9.3005
R21275 VDD.n1471 VDD.n1470 9.3005
R21276 VDD.n1472 VDD.n976 9.3005
R21277 VDD.n1474 VDD.n1473 9.3005
R21278 VDD.n965 VDD.n964 9.3005
R21279 VDD.n1490 VDD.n1489 9.3005
R21280 VDD.n1491 VDD.n963 9.3005
R21281 VDD.n1554 VDD.n1553 9.3005
R21282 VDD.n1550 VDD.n1492 9.3005
R21283 VDD.n1549 VDD.n1495 9.3005
R21284 VDD.n1499 VDD.n1496 9.3005
R21285 VDD.n1500 VDD.n1497 9.3005
R21286 VDD.n1542 VDD.n1501 9.3005
R21287 VDD.n1541 VDD.n1502 9.3005
R21288 VDD.n1540 VDD.n1503 9.3005
R21289 VDD.n1507 VDD.n1504 9.3005
R21290 VDD.n1535 VDD.n1508 9.3005
R21291 VDD.n1534 VDD.n1509 9.3005
R21292 VDD.n1552 VDD.n1551 9.3005
R21293 VDD.n1533 VDD.n1514 9.3005
R21294 VDD.n1628 VDD.n728 9.3005
R21295 VDD.n1627 VDD.n1626 9.3005
R21296 VDD.n733 VDD.n732 9.3005
R21297 VDD.n1621 VDD.n736 9.3005
R21298 VDD.n1620 VDD.n737 9.3005
R21299 VDD.n1619 VDD.n738 9.3005
R21300 VDD.n742 VDD.n739 9.3005
R21301 VDD.n1614 VDD.n743 9.3005
R21302 VDD.n1613 VDD.n744 9.3005
R21303 VDD.n1612 VDD.n745 9.3005
R21304 VDD.n749 VDD.n746 9.3005
R21305 VDD.n1607 VDD.n750 9.3005
R21306 VDD.n1606 VDD.n751 9.3005
R21307 VDD.n1605 VDD.n1604 9.3005
R21308 VDD.n1603 VDD.n752 9.3005
R21309 VDD.n1602 VDD.n1601 9.3005
R21310 VDD.n758 VDD.n757 9.3005
R21311 VDD.n1596 VDD.n762 9.3005
R21312 VDD.n1595 VDD.n763 9.3005
R21313 VDD.n1594 VDD.n764 9.3005
R21314 VDD.n1630 VDD.n1629 9.3005
R21315 VDD.n1532 VDD.n1515 9.3005
R21316 VDD.n1520 VDD.n1516 9.3005
R21317 VDD.n1521 VDD.n1517 9.3005
R21318 VDD.n1525 VDD.n1522 9.3005
R21319 VDD.n1524 VDD.n1523 9.3005
R21320 VDD.n719 VDD.n715 9.3005
R21321 VDD.n1636 VDD.n716 9.3005
R21322 VDD.n1635 VDD.n724 9.3005
R21323 VDD.n731 VDD.n725 9.3005
R21324 VDD.n3400 VDD.n3399 9.3005
R21325 VDD.n3385 VDD.n3384 9.3005
R21326 VDD.n3394 VDD.n3393 9.3005
R21327 VDD.n3392 VDD.n3391 9.3005
R21328 VDD.n3380 VDD.n3379 9.3005
R21329 VDD.n3365 VDD.n3364 9.3005
R21330 VDD.n3374 VDD.n3373 9.3005
R21331 VDD.n3372 VDD.n3371 9.3005
R21332 VDD.n3360 VDD.n3359 9.3005
R21333 VDD.n3345 VDD.n3344 9.3005
R21334 VDD.n3354 VDD.n3353 9.3005
R21335 VDD.n3352 VDD.n3351 9.3005
R21336 VDD.n3340 VDD.n3339 9.3005
R21337 VDD.n3325 VDD.n3324 9.3005
R21338 VDD.n3334 VDD.n3333 9.3005
R21339 VDD.n3332 VDD.n3331 9.3005
R21340 VDD.n3321 VDD.n3320 9.3005
R21341 VDD.n3306 VDD.n3305 9.3005
R21342 VDD.n3315 VDD.n3314 9.3005
R21343 VDD.n3313 VDD.n3312 9.3005
R21344 VDD.n2826 VDD.n2825 9.3005
R21345 VDD.n2829 VDD.n138 9.3005
R21346 VDD.n2830 VDD.n137 9.3005
R21347 VDD.n2833 VDD.n136 9.3005
R21348 VDD.n2834 VDD.n135 9.3005
R21349 VDD.n2837 VDD.n134 9.3005
R21350 VDD.n2838 VDD.n133 9.3005
R21351 VDD.n2841 VDD.n132 9.3005
R21352 VDD.n2842 VDD.n131 9.3005
R21353 VDD.n2845 VDD.n130 9.3005
R21354 VDD.n2846 VDD.n129 9.3005
R21355 VDD.n2849 VDD.n128 9.3005
R21356 VDD.n2853 VDD.n2852 9.3005
R21357 VDD.n2854 VDD.n127 9.3005
R21358 VDD.n2858 VDD.n2855 9.3005
R21359 VDD.n2861 VDD.n126 9.3005
R21360 VDD.n2862 VDD.n125 9.3005
R21361 VDD.n2865 VDD.n124 9.3005
R21362 VDD.n2874 VDD.n121 9.3005
R21363 VDD.n2877 VDD.n120 9.3005
R21364 VDD.n2878 VDD.n119 9.3005
R21365 VDD.n2881 VDD.n118 9.3005
R21366 VDD.n2882 VDD.n117 9.3005
R21367 VDD.n2885 VDD.n116 9.3005
R21368 VDD.n2889 VDD.n112 9.3005
R21369 VDD.n2890 VDD.n111 9.3005
R21370 VDD.n2893 VDD.n110 9.3005
R21371 VDD.n2894 VDD.n109 9.3005
R21372 VDD.n2897 VDD.n108 9.3005
R21373 VDD.n2898 VDD.n107 9.3005
R21374 VDD.n2901 VDD.n106 9.3005
R21375 VDD.n2903 VDD.n105 9.3005
R21376 VDD.n2904 VDD.n104 9.3005
R21377 VDD.n2905 VDD.n103 9.3005
R21378 VDD.n2906 VDD.n102 9.3005
R21379 VDD.n2886 VDD.n113 9.3005
R21380 VDD.n58 VDD.n57 9.3005
R21381 VDD.n2920 VDD.n2919 9.3005
R21382 VDD.n2921 VDD.n56 9.3005
R21383 VDD.n2923 VDD.n2922 9.3005
R21384 VDD.n46 VDD.n45 9.3005
R21385 VDD.n2936 VDD.n2935 9.3005
R21386 VDD.n2937 VDD.n44 9.3005
R21387 VDD.n2939 VDD.n2938 9.3005
R21388 VDD.n34 VDD.n33 9.3005
R21389 VDD.n2952 VDD.n2951 9.3005
R21390 VDD.n2953 VDD.n32 9.3005
R21391 VDD.n2955 VDD.n2954 9.3005
R21392 VDD.n18 VDD.n16 9.3005
R21393 VDD.n3303 VDD.n3302 9.3005
R21394 VDD.n19 VDD.n17 9.3005
R21395 VDD.n3293 VDD.n2969 9.3005
R21396 VDD.n3292 VDD.n2970 9.3005
R21397 VDD.n3291 VDD.n2971 9.3005
R21398 VDD.n2979 VDD.n2972 9.3005
R21399 VDD.n3285 VDD.n2980 9.3005
R21400 VDD.n3284 VDD.n2981 9.3005
R21401 VDD.n3283 VDD.n2982 9.3005
R21402 VDD.n2990 VDD.n2983 9.3005
R21403 VDD.n3277 VDD.n2991 9.3005
R21404 VDD.n3276 VDD.n2992 9.3005
R21405 VDD.n3275 VDD.n2993 9.3005
R21406 VDD.n3076 VDD.n2994 9.3005
R21407 VDD.n3080 VDD.n3075 9.3005
R21408 VDD.n3084 VDD.n3081 9.3005
R21409 VDD.n3085 VDD.n3074 9.3005
R21410 VDD.n3089 VDD.n3088 9.3005
R21411 VDD.n3090 VDD.n3073 9.3005
R21412 VDD.n3094 VDD.n3091 9.3005
R21413 VDD.n3095 VDD.n3072 9.3005
R21414 VDD.n3099 VDD.n3098 9.3005
R21415 VDD.n3100 VDD.n3071 9.3005
R21416 VDD.n3104 VDD.n3101 9.3005
R21417 VDD.n3105 VDD.n3068 9.3005
R21418 VDD.n3109 VDD.n3108 9.3005
R21419 VDD.n3110 VDD.n3067 9.3005
R21420 VDD.n3114 VDD.n3111 9.3005
R21421 VDD.n3115 VDD.n3066 9.3005
R21422 VDD.n3119 VDD.n3118 9.3005
R21423 VDD.n3120 VDD.n3065 9.3005
R21424 VDD.n3124 VDD.n3121 9.3005
R21425 VDD.n3125 VDD.n3064 9.3005
R21426 VDD.n3129 VDD.n3128 9.3005
R21427 VDD.n3130 VDD.n3063 9.3005
R21428 VDD.n3134 VDD.n3131 9.3005
R21429 VDD.n3135 VDD.n3062 9.3005
R21430 VDD.n3139 VDD.n3138 9.3005
R21431 VDD.n3140 VDD.n3061 9.3005
R21432 VDD.n3144 VDD.n3141 9.3005
R21433 VDD.n3145 VDD.n3058 9.3005
R21434 VDD.n3149 VDD.n3148 9.3005
R21435 VDD.n3150 VDD.n3057 9.3005
R21436 VDD.n3154 VDD.n3151 9.3005
R21437 VDD.n3155 VDD.n3056 9.3005
R21438 VDD.n3159 VDD.n3158 9.3005
R21439 VDD.n3160 VDD.n3055 9.3005
R21440 VDD.n3164 VDD.n3161 9.3005
R21441 VDD.n3165 VDD.n3054 9.3005
R21442 VDD.n3169 VDD.n3168 9.3005
R21443 VDD.n3170 VDD.n3053 9.3005
R21444 VDD.n3174 VDD.n3171 9.3005
R21445 VDD.n3175 VDD.n3052 9.3005
R21446 VDD.n3178 VDD.n3049 9.3005
R21447 VDD.n3182 VDD.n3181 9.3005
R21448 VDD.n3183 VDD.n3048 9.3005
R21449 VDD.n3185 VDD.n3184 9.3005
R21450 VDD.n3188 VDD.n3047 9.3005
R21451 VDD.n3192 VDD.n3191 9.3005
R21452 VDD.n3193 VDD.n3046 9.3005
R21453 VDD.n3195 VDD.n3194 9.3005
R21454 VDD.n3198 VDD.n3045 9.3005
R21455 VDD.n3202 VDD.n3201 9.3005
R21456 VDD.n3203 VDD.n3044 9.3005
R21457 VDD.n3205 VDD.n3204 9.3005
R21458 VDD.n3208 VDD.n3041 9.3005
R21459 VDD.n3213 VDD.n3212 9.3005
R21460 VDD.n3214 VDD.n3040 9.3005
R21461 VDD.n3216 VDD.n3215 9.3005
R21462 VDD.n3219 VDD.n3039 9.3005
R21463 VDD.n3223 VDD.n3222 9.3005
R21464 VDD.n3224 VDD.n3038 9.3005
R21465 VDD.n3226 VDD.n3225 9.3005
R21466 VDD.n3229 VDD.n3037 9.3005
R21467 VDD.n3233 VDD.n3232 9.3005
R21468 VDD.n3234 VDD.n3036 9.3005
R21469 VDD.n3236 VDD.n3235 9.3005
R21470 VDD.n3239 VDD.n3035 9.3005
R21471 VDD.n3242 VDD.n3241 9.3005
R21472 VDD.n3243 VDD.n3034 9.3005
R21473 VDD.n3268 VDD.n3267 9.3005
R21474 VDD.n3079 VDD.n3078 9.3005
R21475 VDD.n2915 VDD.n2914 9.3005
R21476 VDD.n52 VDD.n51 9.3005
R21477 VDD.n2928 VDD.n2927 9.3005
R21478 VDD.n2929 VDD.n50 9.3005
R21479 VDD.n2931 VDD.n2930 9.3005
R21480 VDD.n40 VDD.n39 9.3005
R21481 VDD.n2944 VDD.n2943 9.3005
R21482 VDD.n2945 VDD.n38 9.3005
R21483 VDD.n2947 VDD.n2946 9.3005
R21484 VDD.n28 VDD.n27 9.3005
R21485 VDD.n2960 VDD.n2959 9.3005
R21486 VDD.n2961 VDD.n26 9.3005
R21487 VDD.n3299 VDD.n2962 9.3005
R21488 VDD.n3298 VDD.n2963 9.3005
R21489 VDD.n3297 VDD.n2964 9.3005
R21490 VDD.n3248 VDD.n2965 9.3005
R21491 VDD.n3250 VDD.n3249 9.3005
R21492 VDD.n3252 VDD.n3251 9.3005
R21493 VDD.n3253 VDD.n3247 9.3005
R21494 VDD.n3256 VDD.n3254 9.3005
R21495 VDD.n3257 VDD.n3246 9.3005
R21496 VDD.n3259 VDD.n3258 9.3005
R21497 VDD.n3260 VDD.n3245 9.3005
R21498 VDD.n3263 VDD.n3261 9.3005
R21499 VDD.n3264 VDD.n3244 9.3005
R21500 VDD.n3266 VDD.n3265 9.3005
R21501 VDD.n2913 VDD.n62 9.3005
R21502 VDD.n2912 VDD.n2911 9.3005
R21503 VDD.n66 VDD.n63 9.3005
R21504 VDD.n2772 VDD.n2771 9.3005
R21505 VDD.n2775 VDD.n2770 9.3005
R21506 VDD.n2776 VDD.n2769 9.3005
R21507 VDD.n2779 VDD.n2768 9.3005
R21508 VDD.n2780 VDD.n2767 9.3005
R21509 VDD.n2783 VDD.n2766 9.3005
R21510 VDD.n2784 VDD.n2765 9.3005
R21511 VDD.n2787 VDD.n2764 9.3005
R21512 VDD.n2788 VDD.n2763 9.3005
R21513 VDD.n2791 VDD.n2762 9.3005
R21514 VDD.n2792 VDD.n2761 9.3005
R21515 VDD.n2795 VDD.n2760 9.3005
R21516 VDD.n2796 VDD.n2759 9.3005
R21517 VDD.n2799 VDD.n2755 9.3005
R21518 VDD.n2800 VDD.n2754 9.3005
R21519 VDD.n2803 VDD.n2753 9.3005
R21520 VDD.n2812 VDD.n145 9.3005
R21521 VDD.n2815 VDD.n144 9.3005
R21522 VDD.n2816 VDD.n143 9.3005
R21523 VDD.n2819 VDD.n142 9.3005
R21524 VDD.n2823 VDD.n2822 9.3005
R21525 VDD.n2824 VDD.n139 9.3005
R21526 VDD.n1586 VDD.n1585 9.3005
R21527 VDD.n1584 VDD.n917 9.3005
R21528 VDD.n1583 VDD.n1582 9.3005
R21529 VDD.n1581 VDD.n1580 9.3005
R21530 VDD.n1579 VDD.n928 9.3005
R21531 VDD.n1578 VDD.n1577 9.3005
R21532 VDD.n1576 VDD.n934 9.3005
R21533 VDD.n1575 VDD.n1574 9.3005
R21534 VDD.n1573 VDD.n935 9.3005
R21535 VDD.n1572 VDD.n1571 9.3005
R21536 VDD.n1570 VDD.n942 9.3005
R21537 VDD.n1569 VDD.n1568 9.3005
R21538 VDD.n1567 VDD.n943 9.3005
R21539 VDD.n1566 VDD.n1565 9.3005
R21540 VDD.n1564 VDD.n950 9.3005
R21541 VDD.n1563 VDD.n1562 9.3005
R21542 VDD.n1561 VDD.n951 9.3005
R21543 VDD.n1481 VDD.n955 9.3005
R21544 VDD.n1030 VDD.n1029 9.3005
R21545 VDD.n1299 VDD.n1298 9.3005
R21546 VDD.n1300 VDD.n1028 9.3005
R21547 VDD.n1302 VDD.n1301 9.3005
R21548 VDD.n1019 VDD.n1018 9.3005
R21549 VDD.n1315 VDD.n1314 9.3005
R21550 VDD.n1316 VDD.n1017 9.3005
R21551 VDD.n1318 VDD.n1317 9.3005
R21552 VDD.n1007 VDD.n1006 9.3005
R21553 VDD.n1331 VDD.n1330 9.3005
R21554 VDD.n1332 VDD.n1005 9.3005
R21555 VDD.n1334 VDD.n1333 9.3005
R21556 VDD.n996 VDD.n995 9.3005
R21557 VDD.n1447 VDD.n1446 9.3005
R21558 VDD.n1448 VDD.n994 9.3005
R21559 VDD.n1450 VDD.n1449 9.3005
R21560 VDD.n984 VDD.n983 9.3005
R21561 VDD.n1463 VDD.n1462 9.3005
R21562 VDD.n1464 VDD.n982 9.3005
R21563 VDD.n1466 VDD.n1465 9.3005
R21564 VDD.n972 VDD.n971 9.3005
R21565 VDD.n1479 VDD.n1478 9.3005
R21566 VDD.n1480 VDD.n969 9.3005
R21567 VDD.n1485 VDD.n1484 9.3005
R21568 VDD.n1483 VDD.n970 9.3005
R21569 VDD.n1482 VDD.n959 9.3005
R21570 VDD.n1286 VDD.n1285 9.3005
R21571 VDD.n1281 VDD.n1280 9.3005
R21572 VDD.n1279 VDD.n1044 9.3005
R21573 VDD.n1278 VDD.n1277 9.3005
R21574 VDD.n1048 VDD.n1047 9.3005
R21575 VDD.n1270 VDD.n1269 9.3005
R21576 VDD.n1268 VDD.n1050 9.3005
R21577 VDD.n1267 VDD.n1266 9.3005
R21578 VDD.n1052 VDD.n1051 9.3005
R21579 VDD.n1260 VDD.n1259 9.3005
R21580 VDD.n1258 VDD.n1054 9.3005
R21581 VDD.n1257 VDD.n1256 9.3005
R21582 VDD.n1056 VDD.n1055 9.3005
R21583 VDD.n1250 VDD.n1249 9.3005
R21584 VDD.n1248 VDD.n1247 9.3005
R21585 VDD.n1246 VDD.n1061 9.3005
R21586 VDD.n1238 VDD.n1062 9.3005
R21587 VDD.n1240 VDD.n1239 9.3005
R21588 VDD.n1237 VDD.n1064 9.3005
R21589 VDD.n1236 VDD.n1235 9.3005
R21590 VDD.n1066 VDD.n1065 9.3005
R21591 VDD.n1229 VDD.n1228 9.3005
R21592 VDD.n1227 VDD.n1068 9.3005
R21593 VDD.n1226 VDD.n1225 9.3005
R21594 VDD.n1070 VDD.n1069 9.3005
R21595 VDD.n1219 VDD.n1218 9.3005
R21596 VDD.n1217 VDD.n1072 9.3005
R21597 VDD.n1216 VDD.n1215 9.3005
R21598 VDD.n1214 VDD.n1073 9.3005
R21599 VDD.n1204 VDD.n1078 9.3005
R21600 VDD.n1205 VDD.n1079 9.3005
R21601 VDD.n1207 VDD.n1206 9.3005
R21602 VDD.n1203 VDD.n1081 9.3005
R21603 VDD.n1202 VDD.n1201 9.3005
R21604 VDD.n1083 VDD.n1082 9.3005
R21605 VDD.n1195 VDD.n1194 9.3005
R21606 VDD.n1193 VDD.n1085 9.3005
R21607 VDD.n1192 VDD.n1191 9.3005
R21608 VDD.n1087 VDD.n1086 9.3005
R21609 VDD.n1185 VDD.n1184 9.3005
R21610 VDD.n1183 VDD.n1089 9.3005
R21611 VDD.n1182 VDD.n1181 9.3005
R21612 VDD.n1180 VDD.n1090 9.3005
R21613 VDD.n1170 VDD.n1095 9.3005
R21614 VDD.n1171 VDD.n1096 9.3005
R21615 VDD.n1173 VDD.n1172 9.3005
R21616 VDD.n1169 VDD.n1098 9.3005
R21617 VDD.n1168 VDD.n1167 9.3005
R21618 VDD.n1100 VDD.n1099 9.3005
R21619 VDD.n1161 VDD.n1160 9.3005
R21620 VDD.n1159 VDD.n1102 9.3005
R21621 VDD.n1158 VDD.n1157 9.3005
R21622 VDD.n1104 VDD.n1103 9.3005
R21623 VDD.n1151 VDD.n1150 9.3005
R21624 VDD.n1149 VDD.n1106 9.3005
R21625 VDD.n1146 VDD.n1107 9.3005
R21626 VDD.n1136 VDD.n1112 9.3005
R21627 VDD.n1137 VDD.n1113 9.3005
R21628 VDD.n1139 VDD.n1138 9.3005
R21629 VDD.n1135 VDD.n1115 9.3005
R21630 VDD.n1134 VDD.n1133 9.3005
R21631 VDD.n1117 VDD.n1116 9.3005
R21632 VDD.n1127 VDD.n1126 9.3005
R21633 VDD.n1125 VDD.n1119 9.3005
R21634 VDD.n1124 VDD.n1123 9.3005
R21635 VDD.n1120 VDD.n1036 9.3005
R21636 VDD.n1148 VDD.n1147 9.3005
R21637 VDD.n1282 VDD.n1040 9.3005
R21638 VDD.n1284 VDD.n1283 9.3005
R21639 VDD.n1292 VDD.n1035 9.3005
R21640 VDD.n1294 VDD.n1293 9.3005
R21641 VDD.n1025 VDD.n1024 9.3005
R21642 VDD.n1307 VDD.n1306 9.3005
R21643 VDD.n1308 VDD.n1023 9.3005
R21644 VDD.n1310 VDD.n1309 9.3005
R21645 VDD.n1013 VDD.n1012 9.3005
R21646 VDD.n1323 VDD.n1322 9.3005
R21647 VDD.n1324 VDD.n1011 9.3005
R21648 VDD.n1326 VDD.n1325 9.3005
R21649 VDD.n1001 VDD.n1000 9.3005
R21650 VDD.n1339 VDD.n1338 9.3005
R21651 VDD.n1291 VDD.n1290 9.3005
R21652 VDD.n1440 VDD.n999 9.3005
R21653 VDD.n1436 VDD.n1435 9.3005
R21654 VDD.n1421 VDD.n1420 9.3005
R21655 VDD.n1430 VDD.n1429 9.3005
R21656 VDD.n1428 VDD.n1427 9.3005
R21657 VDD.n1416 VDD.n1415 9.3005
R21658 VDD.n1401 VDD.n1400 9.3005
R21659 VDD.n1410 VDD.n1409 9.3005
R21660 VDD.n1408 VDD.n1407 9.3005
R21661 VDD.n1396 VDD.n1395 9.3005
R21662 VDD.n1381 VDD.n1380 9.3005
R21663 VDD.n1390 VDD.n1389 9.3005
R21664 VDD.n1388 VDD.n1387 9.3005
R21665 VDD.n1376 VDD.n1375 9.3005
R21666 VDD.n1361 VDD.n1360 9.3005
R21667 VDD.n1370 VDD.n1369 9.3005
R21668 VDD.n1368 VDD.n1367 9.3005
R21669 VDD.n1357 VDD.n1356 9.3005
R21670 VDD.n1342 VDD.n1341 9.3005
R21671 VDD.n1351 VDD.n1350 9.3005
R21672 VDD.n1349 VDD.n1348 9.3005
R21673 VDD.n1803 VDD.n694 8.85467
R21674 VDD.n1803 VDD.n688 8.85467
R21675 VDD.n1809 VDD.n688 8.85467
R21676 VDD.n1809 VDD.n682 8.85467
R21677 VDD.n1815 VDD.n682 8.85467
R21678 VDD.n1815 VDD.n676 8.85467
R21679 VDD.n1821 VDD.n676 8.85467
R21680 VDD.n1821 VDD.n669 8.85467
R21681 VDD.n1827 VDD.n669 8.85467
R21682 VDD.n1827 VDD.n672 8.85467
R21683 VDD.n1833 VDD.n657 8.85467
R21684 VDD.n1839 VDD.n657 8.85467
R21685 VDD.n1839 VDD.n660 8.85467
R21686 VDD.n1845 VDD.n646 8.85467
R21687 VDD.n1851 VDD.n646 8.85467
R21688 VDD.n1851 VDD.n640 8.85467
R21689 VDD.n1857 VDD.n640 8.85467
R21690 VDD.n1857 VDD.n634 8.85467
R21691 VDD.n1863 VDD.n634 8.85467
R21692 VDD.n1863 VDD.n628 8.85467
R21693 VDD.n1869 VDD.n628 8.85467
R21694 VDD.n1869 VDD.n622 8.85467
R21695 VDD.n1875 VDD.n622 8.85467
R21696 VDD.n1875 VDD.n616 8.85467
R21697 VDD.n1881 VDD.n616 8.85467
R21698 VDD.n1881 VDD.n610 8.85467
R21699 VDD.n1887 VDD.n610 8.85467
R21700 VDD.n1887 VDD.n604 8.85467
R21701 VDD.n1893 VDD.n604 8.85467
R21702 VDD.n1899 VDD.n598 8.85467
R21703 VDD.n1905 VDD.n592 8.85467
R21704 VDD.n1905 VDD.n586 8.85467
R21705 VDD.n1911 VDD.n586 8.85467
R21706 VDD.n1911 VDD.n580 8.85467
R21707 VDD.n1917 VDD.n580 8.85467
R21708 VDD.n1917 VDD.n574 8.85467
R21709 VDD.n1923 VDD.n574 8.85467
R21710 VDD.n1923 VDD.n568 8.85467
R21711 VDD.n1929 VDD.n568 8.85467
R21712 VDD.n1929 VDD.n562 8.85467
R21713 VDD.n1935 VDD.n562 8.85467
R21714 VDD.n1935 VDD.n556 8.85467
R21715 VDD.n1941 VDD.n556 8.85467
R21716 VDD.n1941 VDD.n549 8.85467
R21717 VDD.n1947 VDD.n549 8.85467
R21718 VDD.n1947 VDD.n552 8.85467
R21719 VDD.n1959 VDD.n538 8.85467
R21720 VDD.n1959 VDD.n532 8.85467
R21721 VDD.n1965 VDD.n532 8.85467
R21722 VDD.n1965 VDD.n526 8.85467
R21723 VDD.n1971 VDD.n526 8.85467
R21724 VDD.n1971 VDD.n520 8.85467
R21725 VDD.n1977 VDD.n520 8.85467
R21726 VDD.n1977 VDD.n514 8.85467
R21727 VDD.n1983 VDD.n514 8.85467
R21728 VDD.n1983 VDD.n508 8.85467
R21729 VDD.n1989 VDD.n508 8.85467
R21730 VDD.n1989 VDD.n502 8.85467
R21731 VDD.n1995 VDD.n502 8.85467
R21732 VDD.n1995 VDD.n496 8.85467
R21733 VDD.n2001 VDD.n496 8.85467
R21734 VDD.n2001 VDD.n490 8.85467
R21735 VDD.n2007 VDD.n490 8.85467
R21736 VDD.n2013 VDD.n484 8.85467
R21737 VDD.n2019 VDD.n478 8.85467
R21738 VDD.n2019 VDD.n471 8.85467
R21739 VDD.n2027 VDD.n471 8.85467
R21740 VDD.n2027 VDD.n465 8.85467
R21741 VDD.n2033 VDD.n465 8.85467
R21742 VDD.n2033 VDD.n454 8.85467
R21743 VDD.n2078 VDD.n454 8.85467
R21744 VDD.n2078 VDD.n448 8.85467
R21745 VDD.n2084 VDD.n448 8.85467
R21746 VDD.n2084 VDD.n424 8.85467
R21747 VDD.n2438 VDD.n418 8.85467
R21748 VDD.n2438 VDD.n412 8.85467
R21749 VDD.n2444 VDD.n412 8.85467
R21750 VDD.n2444 VDD.n406 8.85467
R21751 VDD.n2450 VDD.n406 8.85467
R21752 VDD.n2450 VDD.n400 8.85467
R21753 VDD.n2456 VDD.n400 8.85467
R21754 VDD.n2456 VDD.n393 8.85467
R21755 VDD.n2462 VDD.n393 8.85467
R21756 VDD.n2462 VDD.n396 8.85467
R21757 VDD.n2468 VDD.n389 8.85467
R21758 VDD.n2474 VDD.n376 8.85467
R21759 VDD.n2480 VDD.n376 8.85467
R21760 VDD.n2480 VDD.n370 8.85467
R21761 VDD.n2486 VDD.n370 8.85467
R21762 VDD.n2486 VDD.n364 8.85467
R21763 VDD.n2492 VDD.n364 8.85467
R21764 VDD.n2492 VDD.n358 8.85467
R21765 VDD.n2498 VDD.n358 8.85467
R21766 VDD.n2498 VDD.n352 8.85467
R21767 VDD.n2504 VDD.n352 8.85467
R21768 VDD.n2504 VDD.n346 8.85467
R21769 VDD.n2510 VDD.n346 8.85467
R21770 VDD.n2510 VDD.n340 8.85467
R21771 VDD.n2516 VDD.n340 8.85467
R21772 VDD.n2516 VDD.n333 8.85467
R21773 VDD.n2522 VDD.n333 8.85467
R21774 VDD.n2522 VDD.n336 8.85467
R21775 VDD.n2534 VDD.n322 8.85467
R21776 VDD.n2534 VDD.n316 8.85467
R21777 VDD.n2540 VDD.n316 8.85467
R21778 VDD.n2540 VDD.n310 8.85467
R21779 VDD.n2546 VDD.n310 8.85467
R21780 VDD.n2546 VDD.n304 8.85467
R21781 VDD.n2552 VDD.n304 8.85467
R21782 VDD.n2552 VDD.n298 8.85467
R21783 VDD.n2558 VDD.n298 8.85467
R21784 VDD.n2558 VDD.n292 8.85467
R21785 VDD.n2564 VDD.n292 8.85467
R21786 VDD.n2564 VDD.n286 8.85467
R21787 VDD.n2570 VDD.n286 8.85467
R21788 VDD.n2570 VDD.n279 8.85467
R21789 VDD.n2576 VDD.n279 8.85467
R21790 VDD.n2576 VDD.n282 8.85467
R21791 VDD.n2582 VDD.n275 8.85467
R21792 VDD.n2588 VDD.n262 8.85467
R21793 VDD.n2594 VDD.n262 8.85467
R21794 VDD.n2594 VDD.n256 8.85467
R21795 VDD.n2600 VDD.n256 8.85467
R21796 VDD.n2600 VDD.n250 8.85467
R21797 VDD.n2606 VDD.n250 8.85467
R21798 VDD.n2606 VDD.n244 8.85467
R21799 VDD.n2612 VDD.n244 8.85467
R21800 VDD.n2612 VDD.n238 8.85467
R21801 VDD.n2618 VDD.n238 8.85467
R21802 VDD.n2618 VDD.n232 8.85467
R21803 VDD.n2624 VDD.n232 8.85467
R21804 VDD.n2624 VDD.n226 8.85467
R21805 VDD.n2630 VDD.n226 8.85467
R21806 VDD.n2630 VDD.n220 8.85467
R21807 VDD.n2636 VDD.n220 8.85467
R21808 VDD.n2642 VDD.n214 8.85467
R21809 VDD.n2642 VDD.n208 8.85467
R21810 VDD.n2648 VDD.n208 8.85467
R21811 VDD.n2654 VDD.n202 8.85467
R21812 VDD.n2654 VDD.n196 8.85467
R21813 VDD.n2660 VDD.n196 8.85467
R21814 VDD.n2660 VDD.n189 8.85467
R21815 VDD.n2688 VDD.n189 8.85467
R21816 VDD.n2688 VDD.n183 8.85467
R21817 VDD.n2694 VDD.n183 8.85467
R21818 VDD.n2694 VDD.n161 8.85467
R21819 VDD.n2732 VDD.n161 8.85467
R21820 VDD.n2732 VDD.n163 8.85467
R21821 VDD.n2007 VDD.t139 8.72446
R21822 VDD.n2474 VDD.t115 8.72446
R21823 VDD.n15 VDD.n14 8.44301
R21824 VDD.n1033 VDD.t3 8.33383
R21825 VDD.t48 VDD.n967 8.33383
R21826 VDD.n2925 VDD.t7 8.33383
R21827 VDD.t28 VDD.n3279 8.33383
R21828 VDD.t96 VDD.n592 7.42238
R21829 VDD.n282 VDD.t105 7.42238
R21830 VDD.n1833 VDD.t11 7.29217
R21831 VDD.n2013 VDD.t21 7.29217
R21832 VDD.n2468 VDD.t61 7.29217
R21833 VDD.n2648 VDD.t44 7.29217
R21834 VDD.n1893 VDD.t102 7.03175
R21835 VDD.n1953 VDD.t120 7.03175
R21836 VDD.n2528 VDD.t123 7.03175
R21837 VDD.n2588 VDD.t119 7.03175
R21838 VDD.n1215 VDD.n1214 6.78838
R21839 VDD.n1147 VDD.n1106 6.78838
R21840 VDD.n1606 VDD.n1605 6.78838
R21841 VDD.n1533 VDD.n1532 6.78838
R21842 VDD.n3175 VDD.n3174 6.78838
R21843 VDD.n3108 VDD.n3105 6.78838
R21844 VDD.n2829 VDD.n2826 6.78838
R21845 VDD.n2886 VDD.n2885 6.78838
R21846 VDD.n660 VDD.t100 6.64112
R21847 VDD.t117 VDD.n214 6.64112
R21848 VDD.n1250 VDD.n1060 6.01262
R21849 VDD.n1580 VDD.n927 6.01262
R21850 VDD.n3212 VDD.n3209 6.01262
R21851 VDD.n2796 VDD.n2758 6.01262
R21852 VDD.n2094 VDD.n2093 5.93221
R21853 VDD.n1777 VDD.n1776 5.93221
R21854 VDD.n2408 VDD.n2407 5.93221
R21855 VDD.n2707 VDD.n2706 5.93221
R21856 VDD.n2743 VDD.n2742 5.93221
R21857 VDD.n2153 VDD.n2134 5.93221
R21858 VDD.n2049 VDD.n462 5.93221
R21859 VDD.n908 VDD.n786 5.93221
R21860 VDD.n1953 VDD.t113 5.07862
R21861 VDD.n2528 VDD.t121 5.07862
R21862 VDD.n1588 VDD.n765 4.74817
R21863 VDD.n916 VDD.n768 4.74817
R21864 VDD.n1645 VDD.n1644 4.74817
R21865 VDD.n722 VDD.n717 4.74817
R21866 VDD.n1645 VDD.n718 4.74817
R21867 VDD.n1637 VDD.n717 4.74817
R21868 VDD.n2873 VDD.n122 4.74817
R21869 VDD.n2866 VDD.n123 4.74817
R21870 VDD.n2869 VDD.n123 4.74817
R21871 VDD.n2870 VDD.n122 4.74817
R21872 VDD.n2808 VDD.n146 4.74817
R21873 VDD.n2804 VDD.n147 4.74817
R21874 VDD.n2807 VDD.n147 4.74817
R21875 VDD.n2811 VDD.n146 4.74817
R21876 VDD.n1589 VDD.n1588 4.74817
R21877 VDD.n918 VDD.n916 4.74817
R21878 VDD.n1304 VDD.t3 4.688
R21879 VDD.n1476 VDD.t48 4.688
R21880 VDD.t7 VDD.n48 4.688
R21881 VDD.n3280 VDD.t28 4.688
R21882 VDD.n2093 VDD.n2092 4.68343
R21883 VDD.n1776 VDD.n1775 4.68343
R21884 VDD.n2407 VDD.n2406 4.68343
R21885 VDD.n2706 VDD.n2705 4.68343
R21886 VDD.n2742 VDD.n2741 4.68343
R21887 VDD.n2156 VDD.n2134 4.68343
R21888 VDD.n2046 VDD.n462 4.68343
R21889 VDD.n905 VDD.n786 4.68343
R21890 VDD.n3403 VDD.n3303 4.65387
R21891 VDD.n1440 VDD.n1439 4.65387
R21892 VDD.n1439 VDD.n15 4.04185
R21893 VDD VDD.n3403 4.03401
R21894 VDD.n3392 VDD.n3388 3.78097
R21895 VDD.n3372 VDD.n3368 3.78097
R21896 VDD.n3352 VDD.n3348 3.78097
R21897 VDD.n3332 VDD.n3328 3.78097
R21898 VDD.n3313 VDD.n3309 3.78097
R21899 VDD.n1428 VDD.n1424 3.78097
R21900 VDD.n1408 VDD.n1404 3.78097
R21901 VDD.n1388 VDD.n1384 3.78097
R21902 VDD.n1368 VDD.n1364 3.78097
R21903 VDD.n1349 VDD.n1345 3.78097
R21904 VDD.t113 VDD.n538 3.77654
R21905 VDD.n336 VDD.t121 3.77654
R21906 VDD.n3401 VDD.n3383 3.49141
R21907 VDD.n3381 VDD.n3363 3.49141
R21908 VDD.n3361 VDD.n3343 3.49141
R21909 VDD.n3341 VDD.n3323 3.49141
R21910 VDD.n3322 VDD.n3304 3.49141
R21911 VDD.n1437 VDD.n1419 3.49141
R21912 VDD.n1417 VDD.n1399 3.49141
R21913 VDD.n1397 VDD.n1379 3.49141
R21914 VDD.n1377 VDD.n1359 3.49141
R21915 VDD.n1358 VDD.n1340 3.49141
R21916 VDD.n4 VDD.n2 3.3852
R21917 VDD.n11 VDD.n9 3.3852
R21918 VDD.n3399 VDD.n3398 2.71565
R21919 VDD.n3379 VDD.n3378 2.71565
R21920 VDD.n3359 VDD.n3358 2.71565
R21921 VDD.n3339 VDD.n3338 2.71565
R21922 VDD.n3320 VDD.n3319 2.71565
R21923 VDD.n1435 VDD.n1434 2.71565
R21924 VDD.n1415 VDD.n1414 2.71565
R21925 VDD.n1395 VDD.n1394 2.71565
R21926 VDD.n1375 VDD.n1374 2.71565
R21927 VDD.n1356 VDD.n1355 2.71565
R21928 VDD.n6 VDD.n4 2.69878
R21929 VDD.n13 VDD.n11 2.69878
R21930 VDD.n1646 VDD.n1645 2.27742
R21931 VDD.n1646 VDD.n717 2.27742
R21932 VDD.n2714 VDD.n123 2.27742
R21933 VDD.n2714 VDD.n122 2.27742
R21934 VDD.n2752 VDD.n147 2.27742
R21935 VDD.n2752 VDD.n146 2.27742
R21936 VDD.n1588 VDD.n1587 2.27742
R21937 VDD.n1587 VDD.n916 2.27742
R21938 VDD.n1845 VDD.t100 2.21404
R21939 VDD.n2636 VDD.t117 2.21404
R21940 VDD.n14 VDD.n6 2.08886
R21941 VDD.n14 VDD.n13 2.08886
R21942 VDD.n3395 VDD.n3385 1.93989
R21943 VDD.n3375 VDD.n3365 1.93989
R21944 VDD.n3355 VDD.n3345 1.93989
R21945 VDD.n3335 VDD.n3325 1.93989
R21946 VDD.n3316 VDD.n3306 1.93989
R21947 VDD.n1431 VDD.n1421 1.93989
R21948 VDD.n1411 VDD.n1401 1.93989
R21949 VDD.n1391 VDD.n1381 1.93989
R21950 VDD.n1371 VDD.n1361 1.93989
R21951 VDD.n1352 VDD.n1342 1.93989
R21952 VDD.t102 VDD.n598 1.82342
R21953 VDD.n552 VDD.t120 1.82342
R21954 VDD.t123 VDD.n322 1.82342
R21955 VDD.n275 VDD.t119 1.82342
R21956 VDD.n672 VDD.t11 1.563
R21957 VDD.t21 VDD.n478 1.563
R21958 VDD.n396 VDD.t61 1.563
R21959 VDD.t44 VDD.n202 1.563
R21960 VDD.n3402 VDD.n3382 1.47464
R21961 VDD.n3382 VDD.n3362 1.47464
R21962 VDD.n3362 VDD.n3342 1.47464
R21963 VDD.n1438 VDD.n1418 1.47464
R21964 VDD.n1418 VDD.n1398 1.47464
R21965 VDD.n1398 VDD.n1378 1.47464
R21966 VDD.n1899 VDD.t96 1.43279
R21967 VDD.n2582 VDD.t105 1.43279
R21968 VDD.n3394 VDD.n3387 1.16414
R21969 VDD.n3374 VDD.n3367 1.16414
R21970 VDD.n3354 VDD.n3347 1.16414
R21971 VDD.n3334 VDD.n3327 1.16414
R21972 VDD.n3315 VDD.n3308 1.16414
R21973 VDD.n1430 VDD.n1423 1.16414
R21974 VDD.n1410 VDD.n1403 1.16414
R21975 VDD.n1390 VDD.n1383 1.16414
R21976 VDD.n1370 VDD.n1363 1.16414
R21977 VDD.n1351 VDD.n1344 1.16414
R21978 VDD.n1247 VDD.n1060 0.582318
R21979 VDD.n1583 VDD.n927 0.582318
R21980 VDD.n3209 VDD.n3208 0.582318
R21981 VDD.n2799 VDD.n2758 0.582318
R21982 VDD.n3403 VDD.n3402 0.539233
R21983 VDD.n1439 VDD.n1438 0.539233
R21984 VDD.n1553 VDD.n1552 0.465439
R21985 VDD.n102 VDD.n57 0.465439
R21986 VDD.n3079 VDD.n3076 0.465439
R21987 VDD.n3267 VDD.n3266 0.465439
R21988 VDD.n2913 VDD.n2912 0.465439
R21989 VDD.n1482 VDD.n1481 0.465439
R21990 VDD.n1285 VDD.n1284 0.465439
R21991 VDD.n1291 VDD.n1036 0.465439
R21992 VDD.n3391 VDD.n3390 0.388379
R21993 VDD.n3371 VDD.n3370 0.388379
R21994 VDD.n3351 VDD.n3350 0.388379
R21995 VDD.n3331 VDD.n3330 0.388379
R21996 VDD.n3312 VDD.n3311 0.388379
R21997 VDD.n1427 VDD.n1426 0.388379
R21998 VDD.n1407 VDD.n1406 0.388379
R21999 VDD.n1387 VDD.n1386 0.388379
R22000 VDD.n1367 VDD.n1366 0.388379
R22001 VDD.n1348 VDD.n1347 0.388379
R22002 VDD.n3400 VDD.n3384 0.155672
R22003 VDD.n3393 VDD.n3384 0.155672
R22004 VDD.n3393 VDD.n3392 0.155672
R22005 VDD.n3380 VDD.n3364 0.155672
R22006 VDD.n3373 VDD.n3364 0.155672
R22007 VDD.n3373 VDD.n3372 0.155672
R22008 VDD.n3360 VDD.n3344 0.155672
R22009 VDD.n3353 VDD.n3344 0.155672
R22010 VDD.n3353 VDD.n3352 0.155672
R22011 VDD.n3340 VDD.n3324 0.155672
R22012 VDD.n3333 VDD.n3324 0.155672
R22013 VDD.n3333 VDD.n3332 0.155672
R22014 VDD.n3321 VDD.n3305 0.155672
R22015 VDD.n3314 VDD.n3305 0.155672
R22016 VDD.n3314 VDD.n3313 0.155672
R22017 VDD.n1436 VDD.n1420 0.155672
R22018 VDD.n1429 VDD.n1420 0.155672
R22019 VDD.n1429 VDD.n1428 0.155672
R22020 VDD.n1416 VDD.n1400 0.155672
R22021 VDD.n1409 VDD.n1400 0.155672
R22022 VDD.n1409 VDD.n1408 0.155672
R22023 VDD.n1396 VDD.n1380 0.155672
R22024 VDD.n1389 VDD.n1380 0.155672
R22025 VDD.n1389 VDD.n1388 0.155672
R22026 VDD.n1376 VDD.n1360 0.155672
R22027 VDD.n1369 VDD.n1360 0.155672
R22028 VDD.n1369 VDD.n1368 0.155672
R22029 VDD.n1357 VDD.n1341 0.155672
R22030 VDD.n1350 VDD.n1341 0.155672
R22031 VDD.n1350 VDD.n1349 0.155672
R22032 VDD.n1441 VDD.n989 0.152939
R22033 VDD.n1455 VDD.n989 0.152939
R22034 VDD.n1456 VDD.n1455 0.152939
R22035 VDD.n1457 VDD.n1456 0.152939
R22036 VDD.n1457 VDD.n977 0.152939
R22037 VDD.n1471 VDD.n977 0.152939
R22038 VDD.n1472 VDD.n1471 0.152939
R22039 VDD.n1473 VDD.n1472 0.152939
R22040 VDD.n1473 VDD.n964 0.152939
R22041 VDD.n1490 VDD.n964 0.152939
R22042 VDD.n1491 VDD.n1490 0.152939
R22043 VDD.n1553 VDD.n1491 0.152939
R22044 VDD.n1552 VDD.n1492 0.152939
R22045 VDD.n1495 VDD.n1492 0.152939
R22046 VDD.n1499 VDD.n1495 0.152939
R22047 VDD.n1500 VDD.n1499 0.152939
R22048 VDD.n1501 VDD.n1500 0.152939
R22049 VDD.n1502 VDD.n1501 0.152939
R22050 VDD.n1503 VDD.n1502 0.152939
R22051 VDD.n1507 VDD.n1503 0.152939
R22052 VDD.n1508 VDD.n1507 0.152939
R22053 VDD.n1509 VDD.n1508 0.152939
R22054 VDD.n1514 VDD.n1509 0.152939
R22055 VDD.n1515 VDD.n1514 0.152939
R22056 VDD.n1520 VDD.n1515 0.152939
R22057 VDD.n1521 VDD.n1520 0.152939
R22058 VDD.n1522 VDD.n1521 0.152939
R22059 VDD.n1523 VDD.n1522 0.152939
R22060 VDD.n1523 VDD.n715 0.152939
R22061 VDD.n724 VDD.n716 0.152939
R22062 VDD.n731 VDD.n724 0.152939
R22063 VDD.n1629 VDD.n731 0.152939
R22064 VDD.n1629 VDD.n1628 0.152939
R22065 VDD.n1628 VDD.n1627 0.152939
R22066 VDD.n1627 VDD.n732 0.152939
R22067 VDD.n736 VDD.n732 0.152939
R22068 VDD.n737 VDD.n736 0.152939
R22069 VDD.n738 VDD.n737 0.152939
R22070 VDD.n742 VDD.n738 0.152939
R22071 VDD.n743 VDD.n742 0.152939
R22072 VDD.n744 VDD.n743 0.152939
R22073 VDD.n745 VDD.n744 0.152939
R22074 VDD.n749 VDD.n745 0.152939
R22075 VDD.n750 VDD.n749 0.152939
R22076 VDD.n751 VDD.n750 0.152939
R22077 VDD.n1604 VDD.n751 0.152939
R22078 VDD.n1604 VDD.n1603 0.152939
R22079 VDD.n1603 VDD.n1602 0.152939
R22080 VDD.n1602 VDD.n757 0.152939
R22081 VDD.n762 VDD.n757 0.152939
R22082 VDD.n763 VDD.n762 0.152939
R22083 VDD.n764 VDD.n763 0.152939
R22084 VDD.n125 VDD.n124 0.152939
R22085 VDD.n126 VDD.n125 0.152939
R22086 VDD.n2855 VDD.n126 0.152939
R22087 VDD.n2855 VDD.n2854 0.152939
R22088 VDD.n2854 VDD.n2853 0.152939
R22089 VDD.n2853 VDD.n128 0.152939
R22090 VDD.n129 VDD.n128 0.152939
R22091 VDD.n130 VDD.n129 0.152939
R22092 VDD.n131 VDD.n130 0.152939
R22093 VDD.n132 VDD.n131 0.152939
R22094 VDD.n133 VDD.n132 0.152939
R22095 VDD.n134 VDD.n133 0.152939
R22096 VDD.n135 VDD.n134 0.152939
R22097 VDD.n136 VDD.n135 0.152939
R22098 VDD.n137 VDD.n136 0.152939
R22099 VDD.n138 VDD.n137 0.152939
R22100 VDD.n2825 VDD.n138 0.152939
R22101 VDD.n2825 VDD.n2824 0.152939
R22102 VDD.n2824 VDD.n2823 0.152939
R22103 VDD.n2823 VDD.n142 0.152939
R22104 VDD.n143 VDD.n142 0.152939
R22105 VDD.n144 VDD.n143 0.152939
R22106 VDD.n145 VDD.n144 0.152939
R22107 VDD.n103 VDD.n102 0.152939
R22108 VDD.n104 VDD.n103 0.152939
R22109 VDD.n105 VDD.n104 0.152939
R22110 VDD.n106 VDD.n105 0.152939
R22111 VDD.n107 VDD.n106 0.152939
R22112 VDD.n108 VDD.n107 0.152939
R22113 VDD.n109 VDD.n108 0.152939
R22114 VDD.n110 VDD.n109 0.152939
R22115 VDD.n111 VDD.n110 0.152939
R22116 VDD.n112 VDD.n111 0.152939
R22117 VDD.n113 VDD.n112 0.152939
R22118 VDD.n116 VDD.n113 0.152939
R22119 VDD.n117 VDD.n116 0.152939
R22120 VDD.n118 VDD.n117 0.152939
R22121 VDD.n119 VDD.n118 0.152939
R22122 VDD.n120 VDD.n119 0.152939
R22123 VDD.n121 VDD.n120 0.152939
R22124 VDD.n2920 VDD.n57 0.152939
R22125 VDD.n2921 VDD.n2920 0.152939
R22126 VDD.n2922 VDD.n2921 0.152939
R22127 VDD.n2922 VDD.n45 0.152939
R22128 VDD.n2936 VDD.n45 0.152939
R22129 VDD.n2937 VDD.n2936 0.152939
R22130 VDD.n2938 VDD.n2937 0.152939
R22131 VDD.n2938 VDD.n33 0.152939
R22132 VDD.n2952 VDD.n33 0.152939
R22133 VDD.n2953 VDD.n2952 0.152939
R22134 VDD.n2954 VDD.n2953 0.152939
R22135 VDD.n2954 VDD.n16 0.152939
R22136 VDD.n2969 VDD.n17 0.152939
R22137 VDD.n2970 VDD.n2969 0.152939
R22138 VDD.n2971 VDD.n2970 0.152939
R22139 VDD.n2979 VDD.n2971 0.152939
R22140 VDD.n2980 VDD.n2979 0.152939
R22141 VDD.n2981 VDD.n2980 0.152939
R22142 VDD.n2982 VDD.n2981 0.152939
R22143 VDD.n2990 VDD.n2982 0.152939
R22144 VDD.n2991 VDD.n2990 0.152939
R22145 VDD.n2992 VDD.n2991 0.152939
R22146 VDD.n2993 VDD.n2992 0.152939
R22147 VDD.n3076 VDD.n2993 0.152939
R22148 VDD.n3080 VDD.n3079 0.152939
R22149 VDD.n3081 VDD.n3080 0.152939
R22150 VDD.n3081 VDD.n3074 0.152939
R22151 VDD.n3089 VDD.n3074 0.152939
R22152 VDD.n3090 VDD.n3089 0.152939
R22153 VDD.n3091 VDD.n3090 0.152939
R22154 VDD.n3091 VDD.n3072 0.152939
R22155 VDD.n3099 VDD.n3072 0.152939
R22156 VDD.n3100 VDD.n3099 0.152939
R22157 VDD.n3101 VDD.n3100 0.152939
R22158 VDD.n3101 VDD.n3068 0.152939
R22159 VDD.n3109 VDD.n3068 0.152939
R22160 VDD.n3110 VDD.n3109 0.152939
R22161 VDD.n3111 VDD.n3110 0.152939
R22162 VDD.n3111 VDD.n3066 0.152939
R22163 VDD.n3119 VDD.n3066 0.152939
R22164 VDD.n3120 VDD.n3119 0.152939
R22165 VDD.n3121 VDD.n3120 0.152939
R22166 VDD.n3121 VDD.n3064 0.152939
R22167 VDD.n3129 VDD.n3064 0.152939
R22168 VDD.n3130 VDD.n3129 0.152939
R22169 VDD.n3131 VDD.n3130 0.152939
R22170 VDD.n3131 VDD.n3062 0.152939
R22171 VDD.n3139 VDD.n3062 0.152939
R22172 VDD.n3140 VDD.n3139 0.152939
R22173 VDD.n3141 VDD.n3140 0.152939
R22174 VDD.n3141 VDD.n3058 0.152939
R22175 VDD.n3149 VDD.n3058 0.152939
R22176 VDD.n3150 VDD.n3149 0.152939
R22177 VDD.n3151 VDD.n3150 0.152939
R22178 VDD.n3151 VDD.n3056 0.152939
R22179 VDD.n3159 VDD.n3056 0.152939
R22180 VDD.n3160 VDD.n3159 0.152939
R22181 VDD.n3161 VDD.n3160 0.152939
R22182 VDD.n3161 VDD.n3054 0.152939
R22183 VDD.n3169 VDD.n3054 0.152939
R22184 VDD.n3170 VDD.n3169 0.152939
R22185 VDD.n3171 VDD.n3170 0.152939
R22186 VDD.n3171 VDD.n3052 0.152939
R22187 VDD.n3052 VDD.n3049 0.152939
R22188 VDD.n3182 VDD.n3049 0.152939
R22189 VDD.n3183 VDD.n3182 0.152939
R22190 VDD.n3184 VDD.n3183 0.152939
R22191 VDD.n3184 VDD.n3047 0.152939
R22192 VDD.n3192 VDD.n3047 0.152939
R22193 VDD.n3193 VDD.n3192 0.152939
R22194 VDD.n3194 VDD.n3193 0.152939
R22195 VDD.n3194 VDD.n3045 0.152939
R22196 VDD.n3202 VDD.n3045 0.152939
R22197 VDD.n3203 VDD.n3202 0.152939
R22198 VDD.n3204 VDD.n3203 0.152939
R22199 VDD.n3204 VDD.n3041 0.152939
R22200 VDD.n3213 VDD.n3041 0.152939
R22201 VDD.n3214 VDD.n3213 0.152939
R22202 VDD.n3215 VDD.n3214 0.152939
R22203 VDD.n3215 VDD.n3039 0.152939
R22204 VDD.n3223 VDD.n3039 0.152939
R22205 VDD.n3224 VDD.n3223 0.152939
R22206 VDD.n3225 VDD.n3224 0.152939
R22207 VDD.n3225 VDD.n3037 0.152939
R22208 VDD.n3233 VDD.n3037 0.152939
R22209 VDD.n3234 VDD.n3233 0.152939
R22210 VDD.n3235 VDD.n3234 0.152939
R22211 VDD.n3235 VDD.n3035 0.152939
R22212 VDD.n3242 VDD.n3035 0.152939
R22213 VDD.n3243 VDD.n3242 0.152939
R22214 VDD.n3267 VDD.n3243 0.152939
R22215 VDD.n2914 VDD.n2913 0.152939
R22216 VDD.n2914 VDD.n51 0.152939
R22217 VDD.n2928 VDD.n51 0.152939
R22218 VDD.n2929 VDD.n2928 0.152939
R22219 VDD.n2930 VDD.n2929 0.152939
R22220 VDD.n2930 VDD.n39 0.152939
R22221 VDD.n2944 VDD.n39 0.152939
R22222 VDD.n2945 VDD.n2944 0.152939
R22223 VDD.n2946 VDD.n2945 0.152939
R22224 VDD.n2946 VDD.n27 0.152939
R22225 VDD.n2960 VDD.n27 0.152939
R22226 VDD.n2961 VDD.n2960 0.152939
R22227 VDD.n2962 VDD.n2961 0.152939
R22228 VDD.n2963 VDD.n2962 0.152939
R22229 VDD.n2964 VDD.n2963 0.152939
R22230 VDD.n3248 VDD.n2964 0.152939
R22231 VDD.n3249 VDD.n3248 0.152939
R22232 VDD.n3252 VDD.n3249 0.152939
R22233 VDD.n3253 VDD.n3252 0.152939
R22234 VDD.n3254 VDD.n3253 0.152939
R22235 VDD.n3254 VDD.n3246 0.152939
R22236 VDD.n3259 VDD.n3246 0.152939
R22237 VDD.n3260 VDD.n3259 0.152939
R22238 VDD.n3261 VDD.n3260 0.152939
R22239 VDD.n3261 VDD.n3244 0.152939
R22240 VDD.n3266 VDD.n3244 0.152939
R22241 VDD.n2754 VDD.n2753 0.152939
R22242 VDD.n2755 VDD.n2754 0.152939
R22243 VDD.n2759 VDD.n2755 0.152939
R22244 VDD.n2760 VDD.n2759 0.152939
R22245 VDD.n2761 VDD.n2760 0.152939
R22246 VDD.n2762 VDD.n2761 0.152939
R22247 VDD.n2763 VDD.n2762 0.152939
R22248 VDD.n2764 VDD.n2763 0.152939
R22249 VDD.n2765 VDD.n2764 0.152939
R22250 VDD.n2766 VDD.n2765 0.152939
R22251 VDD.n2767 VDD.n2766 0.152939
R22252 VDD.n2768 VDD.n2767 0.152939
R22253 VDD.n2769 VDD.n2768 0.152939
R22254 VDD.n2770 VDD.n2769 0.152939
R22255 VDD.n2771 VDD.n2770 0.152939
R22256 VDD.n2771 VDD.n63 0.152939
R22257 VDD.n2912 VDD.n63 0.152939
R22258 VDD.n1586 VDD.n917 0.152939
R22259 VDD.n1582 VDD.n917 0.152939
R22260 VDD.n1582 VDD.n1581 0.152939
R22261 VDD.n1581 VDD.n928 0.152939
R22262 VDD.n1577 VDD.n928 0.152939
R22263 VDD.n1577 VDD.n1576 0.152939
R22264 VDD.n1576 VDD.n1575 0.152939
R22265 VDD.n1575 VDD.n935 0.152939
R22266 VDD.n1571 VDD.n935 0.152939
R22267 VDD.n1571 VDD.n1570 0.152939
R22268 VDD.n1570 VDD.n1569 0.152939
R22269 VDD.n1569 VDD.n943 0.152939
R22270 VDD.n1565 VDD.n943 0.152939
R22271 VDD.n1565 VDD.n1564 0.152939
R22272 VDD.n1564 VDD.n1563 0.152939
R22273 VDD.n1563 VDD.n951 0.152939
R22274 VDD.n1481 VDD.n951 0.152939
R22275 VDD.n1285 VDD.n1029 0.152939
R22276 VDD.n1299 VDD.n1029 0.152939
R22277 VDD.n1300 VDD.n1299 0.152939
R22278 VDD.n1301 VDD.n1300 0.152939
R22279 VDD.n1301 VDD.n1018 0.152939
R22280 VDD.n1315 VDD.n1018 0.152939
R22281 VDD.n1316 VDD.n1315 0.152939
R22282 VDD.n1317 VDD.n1316 0.152939
R22283 VDD.n1317 VDD.n1006 0.152939
R22284 VDD.n1331 VDD.n1006 0.152939
R22285 VDD.n1332 VDD.n1331 0.152939
R22286 VDD.n1333 VDD.n1332 0.152939
R22287 VDD.n1333 VDD.n995 0.152939
R22288 VDD.n1447 VDD.n995 0.152939
R22289 VDD.n1448 VDD.n1447 0.152939
R22290 VDD.n1449 VDD.n1448 0.152939
R22291 VDD.n1449 VDD.n983 0.152939
R22292 VDD.n1463 VDD.n983 0.152939
R22293 VDD.n1464 VDD.n1463 0.152939
R22294 VDD.n1465 VDD.n1464 0.152939
R22295 VDD.n1465 VDD.n971 0.152939
R22296 VDD.n1479 VDD.n971 0.152939
R22297 VDD.n1480 VDD.n1479 0.152939
R22298 VDD.n1484 VDD.n1480 0.152939
R22299 VDD.n1484 VDD.n1483 0.152939
R22300 VDD.n1483 VDD.n1482 0.152939
R22301 VDD.n1124 VDD.n1036 0.152939
R22302 VDD.n1125 VDD.n1124 0.152939
R22303 VDD.n1126 VDD.n1125 0.152939
R22304 VDD.n1126 VDD.n1116 0.152939
R22305 VDD.n1134 VDD.n1116 0.152939
R22306 VDD.n1135 VDD.n1134 0.152939
R22307 VDD.n1138 VDD.n1135 0.152939
R22308 VDD.n1138 VDD.n1137 0.152939
R22309 VDD.n1137 VDD.n1136 0.152939
R22310 VDD.n1136 VDD.n1107 0.152939
R22311 VDD.n1148 VDD.n1107 0.152939
R22312 VDD.n1149 VDD.n1148 0.152939
R22313 VDD.n1150 VDD.n1149 0.152939
R22314 VDD.n1150 VDD.n1103 0.152939
R22315 VDD.n1158 VDD.n1103 0.152939
R22316 VDD.n1159 VDD.n1158 0.152939
R22317 VDD.n1160 VDD.n1159 0.152939
R22318 VDD.n1160 VDD.n1099 0.152939
R22319 VDD.n1168 VDD.n1099 0.152939
R22320 VDD.n1169 VDD.n1168 0.152939
R22321 VDD.n1172 VDD.n1169 0.152939
R22322 VDD.n1172 VDD.n1171 0.152939
R22323 VDD.n1171 VDD.n1170 0.152939
R22324 VDD.n1170 VDD.n1090 0.152939
R22325 VDD.n1182 VDD.n1090 0.152939
R22326 VDD.n1183 VDD.n1182 0.152939
R22327 VDD.n1184 VDD.n1183 0.152939
R22328 VDD.n1184 VDD.n1086 0.152939
R22329 VDD.n1192 VDD.n1086 0.152939
R22330 VDD.n1193 VDD.n1192 0.152939
R22331 VDD.n1194 VDD.n1193 0.152939
R22332 VDD.n1194 VDD.n1082 0.152939
R22333 VDD.n1202 VDD.n1082 0.152939
R22334 VDD.n1203 VDD.n1202 0.152939
R22335 VDD.n1206 VDD.n1203 0.152939
R22336 VDD.n1206 VDD.n1205 0.152939
R22337 VDD.n1205 VDD.n1204 0.152939
R22338 VDD.n1204 VDD.n1073 0.152939
R22339 VDD.n1216 VDD.n1073 0.152939
R22340 VDD.n1217 VDD.n1216 0.152939
R22341 VDD.n1218 VDD.n1217 0.152939
R22342 VDD.n1218 VDD.n1069 0.152939
R22343 VDD.n1226 VDD.n1069 0.152939
R22344 VDD.n1227 VDD.n1226 0.152939
R22345 VDD.n1228 VDD.n1227 0.152939
R22346 VDD.n1228 VDD.n1065 0.152939
R22347 VDD.n1236 VDD.n1065 0.152939
R22348 VDD.n1237 VDD.n1236 0.152939
R22349 VDD.n1239 VDD.n1237 0.152939
R22350 VDD.n1239 VDD.n1238 0.152939
R22351 VDD.n1238 VDD.n1061 0.152939
R22352 VDD.n1248 VDD.n1061 0.152939
R22353 VDD.n1249 VDD.n1248 0.152939
R22354 VDD.n1249 VDD.n1055 0.152939
R22355 VDD.n1257 VDD.n1055 0.152939
R22356 VDD.n1258 VDD.n1257 0.152939
R22357 VDD.n1259 VDD.n1258 0.152939
R22358 VDD.n1259 VDD.n1051 0.152939
R22359 VDD.n1267 VDD.n1051 0.152939
R22360 VDD.n1268 VDD.n1267 0.152939
R22361 VDD.n1269 VDD.n1268 0.152939
R22362 VDD.n1269 VDD.n1047 0.152939
R22363 VDD.n1278 VDD.n1047 0.152939
R22364 VDD.n1279 VDD.n1278 0.152939
R22365 VDD.n1280 VDD.n1279 0.152939
R22366 VDD.n1280 VDD.n1040 0.152939
R22367 VDD.n1284 VDD.n1040 0.152939
R22368 VDD.n1292 VDD.n1291 0.152939
R22369 VDD.n1293 VDD.n1292 0.152939
R22370 VDD.n1293 VDD.n1024 0.152939
R22371 VDD.n1307 VDD.n1024 0.152939
R22372 VDD.n1308 VDD.n1307 0.152939
R22373 VDD.n1309 VDD.n1308 0.152939
R22374 VDD.n1309 VDD.n1012 0.152939
R22375 VDD.n1323 VDD.n1012 0.152939
R22376 VDD.n1324 VDD.n1323 0.152939
R22377 VDD.n1325 VDD.n1324 0.152939
R22378 VDD.n1325 VDD.n1000 0.152939
R22379 VDD.n1339 VDD.n1000 0.152939
R22380 VDD.n1441 VDD.n1440 0.145814
R22381 VDD.n3303 VDD.n16 0.145814
R22382 VDD.n3303 VDD.n17 0.145814
R22383 VDD.n1440 VDD.n1339 0.145814
R22384 VDD.t139 VDD.n484 0.130708
R22385 VDD.n389 VDD.t115 0.130708
R22386 VDD.n1646 VDD.n716 0.1255
R22387 VDD.n1587 VDD.n764 0.1255
R22388 VDD.n2714 VDD.n124 0.1255
R22389 VDD.n2752 VDD.n145 0.1255
R22390 VDD.n1646 VDD.n715 0.027939
R22391 VDD.n2714 VDD.n121 0.027939
R22392 VDD.n2753 VDD.n2752 0.027939
R22393 VDD.n1587 VDD.n1586 0.027939
R22394 VDD VDD.n15 0.00833333
R22395 VN.n190 VN.t1 243.97
R22396 VN.n191 VN.t2 243.255
R22397 VN.n190 VN.n189 223.454
R22398 VN.n186 VN.n185 161.3
R22399 VN.n184 VN.n95 161.3
R22400 VN.n183 VN.n182 161.3
R22401 VN.n181 VN.n96 161.3
R22402 VN.n180 VN.n179 161.3
R22403 VN.n178 VN.n97 161.3
R22404 VN.n177 VN.n176 161.3
R22405 VN.n175 VN.n98 161.3
R22406 VN.n174 VN.n173 161.3
R22407 VN.n172 VN.n99 161.3
R22408 VN.n171 VN.n170 161.3
R22409 VN.n169 VN.n100 161.3
R22410 VN.n168 VN.n167 161.3
R22411 VN.n166 VN.n101 161.3
R22412 VN.n164 VN.n163 161.3
R22413 VN.n162 VN.n102 161.3
R22414 VN.n161 VN.n160 161.3
R22415 VN.n159 VN.n103 161.3
R22416 VN.n158 VN.n157 161.3
R22417 VN.n156 VN.n104 161.3
R22418 VN.n155 VN.n154 161.3
R22419 VN.n153 VN.n105 161.3
R22420 VN.n152 VN.n151 161.3
R22421 VN.n150 VN.n106 161.3
R22422 VN.n149 VN.n148 161.3
R22423 VN.n147 VN.n107 161.3
R22424 VN.n146 VN.n145 161.3
R22425 VN.n144 VN.n108 161.3
R22426 VN.n143 VN.n142 161.3
R22427 VN.n140 VN.n109 161.3
R22428 VN.n139 VN.n138 161.3
R22429 VN.n137 VN.n110 161.3
R22430 VN.n136 VN.n135 161.3
R22431 VN.n134 VN.n111 161.3
R22432 VN.n133 VN.n132 161.3
R22433 VN.n131 VN.n112 161.3
R22434 VN.n130 VN.n129 161.3
R22435 VN.n128 VN.n113 161.3
R22436 VN.n127 VN.n126 161.3
R22437 VN.n125 VN.n114 161.3
R22438 VN.n124 VN.n123 161.3
R22439 VN.n122 VN.n115 161.3
R22440 VN.n121 VN.n120 161.3
R22441 VN.n119 VN.n116 161.3
R22442 VN.n25 VN.n22 161.3
R22443 VN.n27 VN.n26 161.3
R22444 VN.n28 VN.n21 161.3
R22445 VN.n30 VN.n29 161.3
R22446 VN.n31 VN.n20 161.3
R22447 VN.n33 VN.n32 161.3
R22448 VN.n34 VN.n19 161.3
R22449 VN.n36 VN.n35 161.3
R22450 VN.n37 VN.n18 161.3
R22451 VN.n39 VN.n38 161.3
R22452 VN.n40 VN.n17 161.3
R22453 VN.n42 VN.n41 161.3
R22454 VN.n43 VN.n16 161.3
R22455 VN.n45 VN.n44 161.3
R22456 VN.n46 VN.n15 161.3
R22457 VN.n49 VN.n48 161.3
R22458 VN.n50 VN.n14 161.3
R22459 VN.n52 VN.n51 161.3
R22460 VN.n53 VN.n13 161.3
R22461 VN.n55 VN.n54 161.3
R22462 VN.n56 VN.n12 161.3
R22463 VN.n58 VN.n57 161.3
R22464 VN.n59 VN.n11 161.3
R22465 VN.n61 VN.n60 161.3
R22466 VN.n62 VN.n10 161.3
R22467 VN.n64 VN.n63 161.3
R22468 VN.n65 VN.n9 161.3
R22469 VN.n67 VN.n66 161.3
R22470 VN.n68 VN.n8 161.3
R22471 VN.n70 VN.n69 161.3
R22472 VN.n72 VN.n7 161.3
R22473 VN.n74 VN.n73 161.3
R22474 VN.n75 VN.n6 161.3
R22475 VN.n77 VN.n76 161.3
R22476 VN.n78 VN.n5 161.3
R22477 VN.n80 VN.n79 161.3
R22478 VN.n81 VN.n4 161.3
R22479 VN.n83 VN.n82 161.3
R22480 VN.n84 VN.n3 161.3
R22481 VN.n86 VN.n85 161.3
R22482 VN.n87 VN.n2 161.3
R22483 VN.n89 VN.n88 161.3
R22484 VN.n90 VN.n1 161.3
R22485 VN.n92 VN.n91 161.3
R22486 VN.n118 VN.n117 72.9837
R22487 VN.n24 VN.n23 72.9837
R22488 VN.n188 VN.n187 59.4459
R22489 VN.n187 VN.n94 58.5146
R22490 VN.n93 VN.n0 58.5146
R22491 VN.n118 VN.t6 58.337
R22492 VN.n24 VN.t8 58.3365
R22493 VN.n177 VN.n98 56.5193
R22494 VN.n83 VN.n4 56.5193
R22495 VN.n129 VN.n112 49.7204
R22496 VN.n153 VN.n152 49.7204
R22497 VN.n59 VN.n58 49.7204
R22498 VN.n35 VN.n18 49.7204
R22499 VN.n129 VN.n128 31.2664
R22500 VN.n154 VN.n153 31.2664
R22501 VN.n60 VN.n59 31.2664
R22502 VN.n35 VN.n34 31.2664
R22503 VN.n117 VN.t13 24.7565
R22504 VN.n141 VN.t12 24.7565
R22505 VN.n165 VN.t5 24.7565
R22506 VN.n94 VN.t4 24.7565
R22507 VN.n0 VN.t10 24.7565
R22508 VN.n71 VN.t11 24.7565
R22509 VN.n47 VN.t7 24.7565
R22510 VN.n23 VN.t9 24.7565
R22511 VN.n121 VN.n116 24.4675
R22512 VN.n122 VN.n121 24.4675
R22513 VN.n123 VN.n122 24.4675
R22514 VN.n123 VN.n114 24.4675
R22515 VN.n127 VN.n114 24.4675
R22516 VN.n128 VN.n127 24.4675
R22517 VN.n133 VN.n112 24.4675
R22518 VN.n134 VN.n133 24.4675
R22519 VN.n135 VN.n134 24.4675
R22520 VN.n135 VN.n110 24.4675
R22521 VN.n139 VN.n110 24.4675
R22522 VN.n140 VN.n139 24.4675
R22523 VN.n142 VN.n108 24.4675
R22524 VN.n146 VN.n108 24.4675
R22525 VN.n147 VN.n146 24.4675
R22526 VN.n148 VN.n147 24.4675
R22527 VN.n148 VN.n106 24.4675
R22528 VN.n152 VN.n106 24.4675
R22529 VN.n154 VN.n104 24.4675
R22530 VN.n158 VN.n104 24.4675
R22531 VN.n159 VN.n158 24.4675
R22532 VN.n160 VN.n159 24.4675
R22533 VN.n160 VN.n102 24.4675
R22534 VN.n164 VN.n102 24.4675
R22535 VN.n167 VN.n166 24.4675
R22536 VN.n167 VN.n100 24.4675
R22537 VN.n171 VN.n100 24.4675
R22538 VN.n172 VN.n171 24.4675
R22539 VN.n173 VN.n172 24.4675
R22540 VN.n173 VN.n98 24.4675
R22541 VN.n178 VN.n177 24.4675
R22542 VN.n179 VN.n178 24.4675
R22543 VN.n179 VN.n96 24.4675
R22544 VN.n183 VN.n96 24.4675
R22545 VN.n184 VN.n183 24.4675
R22546 VN.n185 VN.n184 24.4675
R22547 VN.n91 VN.n90 24.4675
R22548 VN.n90 VN.n89 24.4675
R22549 VN.n89 VN.n2 24.4675
R22550 VN.n85 VN.n2 24.4675
R22551 VN.n85 VN.n84 24.4675
R22552 VN.n84 VN.n83 24.4675
R22553 VN.n79 VN.n4 24.4675
R22554 VN.n79 VN.n78 24.4675
R22555 VN.n78 VN.n77 24.4675
R22556 VN.n77 VN.n6 24.4675
R22557 VN.n73 VN.n6 24.4675
R22558 VN.n73 VN.n72 24.4675
R22559 VN.n70 VN.n8 24.4675
R22560 VN.n66 VN.n8 24.4675
R22561 VN.n66 VN.n65 24.4675
R22562 VN.n65 VN.n64 24.4675
R22563 VN.n64 VN.n10 24.4675
R22564 VN.n60 VN.n10 24.4675
R22565 VN.n58 VN.n12 24.4675
R22566 VN.n54 VN.n12 24.4675
R22567 VN.n54 VN.n53 24.4675
R22568 VN.n53 VN.n52 24.4675
R22569 VN.n52 VN.n14 24.4675
R22570 VN.n48 VN.n14 24.4675
R22571 VN.n46 VN.n45 24.4675
R22572 VN.n45 VN.n16 24.4675
R22573 VN.n41 VN.n16 24.4675
R22574 VN.n41 VN.n40 24.4675
R22575 VN.n40 VN.n39 24.4675
R22576 VN.n39 VN.n18 24.4675
R22577 VN.n34 VN.n33 24.4675
R22578 VN.n33 VN.n20 24.4675
R22579 VN.n29 VN.n20 24.4675
R22580 VN.n29 VN.n28 24.4675
R22581 VN.n28 VN.n27 24.4675
R22582 VN.n27 VN.n22 24.4675
R22583 VN.n166 VN.n165 21.5315
R22584 VN.n72 VN.n71 21.5315
R22585 VN.n189 VN.t0 19.8005
R22586 VN.n189 VN.t3 19.8005
R22587 VN VN.n192 18.5481
R22588 VN.n185 VN.n94 18.1061
R22589 VN.n91 VN.n0 18.1061
R22590 VN.n188 VN.n93 15.0596
R22591 VN.n141 VN.n140 12.234
R22592 VN.n142 VN.n141 12.234
R22593 VN.n48 VN.n47 12.234
R22594 VN.n47 VN.n46 12.234
R22595 VN.n192 VN.n191 5.04791
R22596 VN.n117 VN.n116 2.93654
R22597 VN.n165 VN.n164 2.93654
R22598 VN.n71 VN.n70 2.93654
R22599 VN.n23 VN.n22 2.93654
R22600 VN.n192 VN.n188 1.188
R22601 VN.n119 VN.n118 0.780565
R22602 VN.n25 VN.n24 0.780562
R22603 VN.n191 VN.n190 0.716017
R22604 VN.n187 VN.n186 0.529113
R22605 VN.n93 VN.n92 0.529113
R22606 VN.n120 VN.n119 0.189894
R22607 VN.n120 VN.n115 0.189894
R22608 VN.n124 VN.n115 0.189894
R22609 VN.n125 VN.n124 0.189894
R22610 VN.n126 VN.n125 0.189894
R22611 VN.n126 VN.n113 0.189894
R22612 VN.n130 VN.n113 0.189894
R22613 VN.n131 VN.n130 0.189894
R22614 VN.n132 VN.n131 0.189894
R22615 VN.n132 VN.n111 0.189894
R22616 VN.n136 VN.n111 0.189894
R22617 VN.n137 VN.n136 0.189894
R22618 VN.n138 VN.n137 0.189894
R22619 VN.n138 VN.n109 0.189894
R22620 VN.n143 VN.n109 0.189894
R22621 VN.n144 VN.n143 0.189894
R22622 VN.n145 VN.n144 0.189894
R22623 VN.n145 VN.n107 0.189894
R22624 VN.n149 VN.n107 0.189894
R22625 VN.n150 VN.n149 0.189894
R22626 VN.n151 VN.n150 0.189894
R22627 VN.n151 VN.n105 0.189894
R22628 VN.n155 VN.n105 0.189894
R22629 VN.n156 VN.n155 0.189894
R22630 VN.n157 VN.n156 0.189894
R22631 VN.n157 VN.n103 0.189894
R22632 VN.n161 VN.n103 0.189894
R22633 VN.n162 VN.n161 0.189894
R22634 VN.n163 VN.n162 0.189894
R22635 VN.n163 VN.n101 0.189894
R22636 VN.n168 VN.n101 0.189894
R22637 VN.n169 VN.n168 0.189894
R22638 VN.n170 VN.n169 0.189894
R22639 VN.n170 VN.n99 0.189894
R22640 VN.n174 VN.n99 0.189894
R22641 VN.n175 VN.n174 0.189894
R22642 VN.n176 VN.n175 0.189894
R22643 VN.n176 VN.n97 0.189894
R22644 VN.n180 VN.n97 0.189894
R22645 VN.n181 VN.n180 0.189894
R22646 VN.n182 VN.n181 0.189894
R22647 VN.n182 VN.n95 0.189894
R22648 VN.n186 VN.n95 0.189894
R22649 VN.n92 VN.n1 0.189894
R22650 VN.n88 VN.n1 0.189894
R22651 VN.n88 VN.n87 0.189894
R22652 VN.n87 VN.n86 0.189894
R22653 VN.n86 VN.n3 0.189894
R22654 VN.n82 VN.n3 0.189894
R22655 VN.n82 VN.n81 0.189894
R22656 VN.n81 VN.n80 0.189894
R22657 VN.n80 VN.n5 0.189894
R22658 VN.n76 VN.n5 0.189894
R22659 VN.n76 VN.n75 0.189894
R22660 VN.n75 VN.n74 0.189894
R22661 VN.n74 VN.n7 0.189894
R22662 VN.n69 VN.n7 0.189894
R22663 VN.n69 VN.n68 0.189894
R22664 VN.n68 VN.n67 0.189894
R22665 VN.n67 VN.n9 0.189894
R22666 VN.n63 VN.n9 0.189894
R22667 VN.n63 VN.n62 0.189894
R22668 VN.n62 VN.n61 0.189894
R22669 VN.n61 VN.n11 0.189894
R22670 VN.n57 VN.n11 0.189894
R22671 VN.n57 VN.n56 0.189894
R22672 VN.n56 VN.n55 0.189894
R22673 VN.n55 VN.n13 0.189894
R22674 VN.n51 VN.n13 0.189894
R22675 VN.n51 VN.n50 0.189894
R22676 VN.n50 VN.n49 0.189894
R22677 VN.n49 VN.n15 0.189894
R22678 VN.n44 VN.n15 0.189894
R22679 VN.n44 VN.n43 0.189894
R22680 VN.n43 VN.n42 0.189894
R22681 VN.n42 VN.n17 0.189894
R22682 VN.n38 VN.n17 0.189894
R22683 VN.n38 VN.n37 0.189894
R22684 VN.n37 VN.n36 0.189894
R22685 VN.n36 VN.n19 0.189894
R22686 VN.n32 VN.n19 0.189894
R22687 VN.n32 VN.n31 0.189894
R22688 VN.n31 VN.n30 0.189894
R22689 VN.n30 VN.n21 0.189894
R22690 VN.n26 VN.n21 0.189894
R22691 VN.n26 VN.n25 0.189894
R22692 a_n4580_9541.n8 a_n4580_9541.t10 181.263
R22693 a_n4580_9541.n3 a_n4580_9541.t8 181.262
R22694 a_n4580_9541.n1 a_n4580_9541.t11 181.262
R22695 a_n4580_9541.n8 a_n4580_9541.t9 178.565
R22696 a_n4580_9541.n0 a_n4580_9541.t3 178.565
R22697 a_n4580_9541.n0 a_n4580_9541.t7 178.565
R22698 a_n4580_9541.n6 a_n4580_9541.t1 178.565
R22699 a_n4580_9541.n1 a_n4580_9541.t12 178.565
R22700 a_n4580_9541.n3 a_n4580_9541.n2 164.245
R22701 a_n4580_9541.n5 a_n4580_9541.n4 164.245
R22702 a_n4580_9541.n7 a_n4580_9541.n1 32.021
R22703 a_n4580_9541.n2 a_n4580_9541.t2 14.3199
R22704 a_n4580_9541.n2 a_n4580_9541.t6 14.3199
R22705 a_n4580_9541.n4 a_n4580_9541.t5 14.3199
R22706 a_n4580_9541.n4 a_n4580_9541.t4 14.3199
R22707 a_n4580_9541.n9 a_n4580_9541.n8 13.6858
R22708 a_n4580_9541.t0 a_n4580_9541.n9 12.2257
R22709 a_n4580_9541.n7 a_n4580_9541.n6 6.35395
R22710 a_n4580_9541.n5 a_n4580_9541.n0 3.3852
R22711 a_n4580_9541.n9 a_n4580_9541.n7 2.79595
R22712 a_n4580_9541.n6 a_n4580_9541.n5 2.69878
R22713 a_n4580_9541.n0 a_n4580_9541.n3 2.69878
R22714 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t3 122.907
R22715 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t1 121.347
R22716 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.t5 121.347
R22717 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.t9 121.347
R22718 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t7 121.347
R22719 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.t2 62.0876
R22720 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t11 61.4537
R22721 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.t0 58.964
R22722 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.t4 58.964
R22723 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.t8 58.964
R22724 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.t6 58.964
R22725 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.t13 58.3302
R22726 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.t12 58.3302
R22727 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.t14 58.3302
R22728 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t10 58.3302
R22729 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 6.10807
R22730 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n4 4.66322
R22731 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n9 4.58428
R22732 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 3.12528
R22733 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 3.12528
R22734 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n5 3.12528
R22735 DIFFPAIR_BIAS.n11 DIFFPAIR_BIAS.n10 3.12523
R22736 DIFFPAIR_BIAS.n12 DIFFPAIR_BIAS.n11 3.12523
R22737 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n0 2.19804
R22738 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.n3 1.56155
R22739 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 1.56155
R22740 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 1.56155
R22741 DIFFPAIR_BIAS DIFFPAIR_BIAS.n13 0.684875
R22742 DIFFPAIR_BIAS.n13 DIFFPAIR_BIAS.n12 0.636994
R22743 a_n7464_n776.n10 a_n7464_n776.t8 222.97
R22744 a_n7464_n776.n43 a_n7464_n776.t9 222.97
R22745 a_n7464_n776.n44 a_n7464_n776.t6 222.97
R22746 a_n7464_n776.n45 a_n7464_n776.t7 222.97
R22747 a_n7464_n776.n46 a_n7464_n776.t5 222.97
R22748 a_n7464_n776.n136 a_n7464_n776.n113 214.453
R22749 a_n7464_n776.n34 a_n7464_n776.n11 214.453
R22750 a_n7464_n776.n107 a_n7464_n776.n84 214.453
R22751 a_n7464_n776.n75 a_n7464_n776.n52 214.453
R22752 a_n7464_n776.n137 a_n7464_n776.n136 185
R22753 a_n7464_n776.n135 a_n7464_n776.n134 185
R22754 a_n7464_n776.n116 a_n7464_n776.n115 185
R22755 a_n7464_n776.n131 a_n7464_n776.n130 185
R22756 a_n7464_n776.n129 a_n7464_n776.n128 185
R22757 a_n7464_n776.n119 a_n7464_n776.n118 185
R22758 a_n7464_n776.n125 a_n7464_n776.n124 185
R22759 a_n7464_n776.n123 a_n7464_n776.n122 185
R22760 a_n7464_n776.n35 a_n7464_n776.n34 185
R22761 a_n7464_n776.n33 a_n7464_n776.n32 185
R22762 a_n7464_n776.n14 a_n7464_n776.n13 185
R22763 a_n7464_n776.n29 a_n7464_n776.n28 185
R22764 a_n7464_n776.n27 a_n7464_n776.n26 185
R22765 a_n7464_n776.n17 a_n7464_n776.n16 185
R22766 a_n7464_n776.n23 a_n7464_n776.n22 185
R22767 a_n7464_n776.n21 a_n7464_n776.n20 185
R22768 a_n7464_n776.n94 a_n7464_n776.n93 185
R22769 a_n7464_n776.n96 a_n7464_n776.n95 185
R22770 a_n7464_n776.n90 a_n7464_n776.n89 185
R22771 a_n7464_n776.n100 a_n7464_n776.n99 185
R22772 a_n7464_n776.n102 a_n7464_n776.n101 185
R22773 a_n7464_n776.n87 a_n7464_n776.n86 185
R22774 a_n7464_n776.n106 a_n7464_n776.n105 185
R22775 a_n7464_n776.n108 a_n7464_n776.n107 185
R22776 a_n7464_n776.n62 a_n7464_n776.n61 185
R22777 a_n7464_n776.n64 a_n7464_n776.n63 185
R22778 a_n7464_n776.n58 a_n7464_n776.n57 185
R22779 a_n7464_n776.n68 a_n7464_n776.n67 185
R22780 a_n7464_n776.n70 a_n7464_n776.n69 185
R22781 a_n7464_n776.n55 a_n7464_n776.n54 185
R22782 a_n7464_n776.n74 a_n7464_n776.n73 185
R22783 a_n7464_n776.n76 a_n7464_n776.n75 185
R22784 a_n7464_n776.n92 a_n7464_n776.t3 149.524
R22785 a_n7464_n776.n60 a_n7464_n776.t20 149.524
R22786 a_n7464_n776.n121 a_n7464_n776.t24 149.524
R22787 a_n7464_n776.n19 a_n7464_n776.t11 149.524
R22788 a_n7464_n776.n136 a_n7464_n776.n135 104.615
R22789 a_n7464_n776.n135 a_n7464_n776.n115 104.615
R22790 a_n7464_n776.n130 a_n7464_n776.n115 104.615
R22791 a_n7464_n776.n130 a_n7464_n776.n129 104.615
R22792 a_n7464_n776.n129 a_n7464_n776.n118 104.615
R22793 a_n7464_n776.n124 a_n7464_n776.n118 104.615
R22794 a_n7464_n776.n124 a_n7464_n776.n123 104.615
R22795 a_n7464_n776.n34 a_n7464_n776.n33 104.615
R22796 a_n7464_n776.n33 a_n7464_n776.n13 104.615
R22797 a_n7464_n776.n28 a_n7464_n776.n13 104.615
R22798 a_n7464_n776.n28 a_n7464_n776.n27 104.615
R22799 a_n7464_n776.n27 a_n7464_n776.n16 104.615
R22800 a_n7464_n776.n22 a_n7464_n776.n16 104.615
R22801 a_n7464_n776.n22 a_n7464_n776.n21 104.615
R22802 a_n7464_n776.n95 a_n7464_n776.n94 104.615
R22803 a_n7464_n776.n95 a_n7464_n776.n89 104.615
R22804 a_n7464_n776.n100 a_n7464_n776.n89 104.615
R22805 a_n7464_n776.n101 a_n7464_n776.n100 104.615
R22806 a_n7464_n776.n101 a_n7464_n776.n86 104.615
R22807 a_n7464_n776.n106 a_n7464_n776.n86 104.615
R22808 a_n7464_n776.n107 a_n7464_n776.n106 104.615
R22809 a_n7464_n776.n63 a_n7464_n776.n62 104.615
R22810 a_n7464_n776.n63 a_n7464_n776.n57 104.615
R22811 a_n7464_n776.n68 a_n7464_n776.n57 104.615
R22812 a_n7464_n776.n69 a_n7464_n776.n68 104.615
R22813 a_n7464_n776.n69 a_n7464_n776.n54 104.615
R22814 a_n7464_n776.n74 a_n7464_n776.n54 104.615
R22815 a_n7464_n776.n75 a_n7464_n776.n74 104.615
R22816 a_n7464_n776.n9 a_n7464_n776.n8 55.3258
R22817 a_n7464_n776.n40 a_n7464_n776.n39 55.3258
R22818 a_n7464_n776.n42 a_n7464_n776.n41 55.3258
R22819 a_n7464_n776.n83 a_n7464_n776.n82 55.3257
R22820 a_n7464_n776.n81 a_n7464_n776.n80 55.3257
R22821 a_n7464_n776.n51 a_n7464_n776.n50 55.3257
R22822 a_n7464_n776.n49 a_n7464_n776.n48 55.3257
R22823 a_n7464_n776.n142 a_n7464_n776.n141 55.3257
R22824 a_n7464_n776.n123 a_n7464_n776.t24 52.3082
R22825 a_n7464_n776.n21 a_n7464_n776.t11 52.3082
R22826 a_n7464_n776.n94 a_n7464_n776.t3 52.3082
R22827 a_n7464_n776.n62 a_n7464_n776.t20 52.3082
R22828 a_n7464_n776.n140 a_n7464_n776.n139 39.555
R22829 a_n7464_n776.n38 a_n7464_n776.n37 39.555
R22830 a_n7464_n776.n111 a_n7464_n776.n110 39.555
R22831 a_n7464_n776.n79 a_n7464_n776.n78 39.555
R22832 a_n7464_n776.n47 a_n7464_n776.n42 15.2562
R22833 a_n7464_n776.n140 a_n7464_n776.n112 13.6808
R22834 a_n7464_n776.n138 a_n7464_n776.n137 12.8005
R22835 a_n7464_n776.n36 a_n7464_n776.n35 12.8005
R22836 a_n7464_n776.n109 a_n7464_n776.n108 12.8005
R22837 a_n7464_n776.n77 a_n7464_n776.n76 12.8005
R22838 a_n7464_n776.n134 a_n7464_n776.n114 12.0247
R22839 a_n7464_n776.n32 a_n7464_n776.n12 12.0247
R22840 a_n7464_n776.n105 a_n7464_n776.n85 12.0247
R22841 a_n7464_n776.n73 a_n7464_n776.n53 12.0247
R22842 a_n7464_n776.n133 a_n7464_n776.n116 11.249
R22843 a_n7464_n776.n31 a_n7464_n776.n14 11.249
R22844 a_n7464_n776.n104 a_n7464_n776.n87 11.249
R22845 a_n7464_n776.n72 a_n7464_n776.n55 11.249
R22846 a_n7464_n776.n132 a_n7464_n776.n131 10.4732
R22847 a_n7464_n776.n30 a_n7464_n776.n29 10.4732
R22848 a_n7464_n776.n103 a_n7464_n776.n102 10.4732
R22849 a_n7464_n776.n71 a_n7464_n776.n70 10.4732
R22850 a_n7464_n776.n122 a_n7464_n776.n121 10.2747
R22851 a_n7464_n776.n20 a_n7464_n776.n19 10.2747
R22852 a_n7464_n776.n93 a_n7464_n776.n92 10.2747
R22853 a_n7464_n776.n61 a_n7464_n776.n60 10.2747
R22854 a_n7464_n776.n128 a_n7464_n776.n117 9.69747
R22855 a_n7464_n776.n26 a_n7464_n776.n15 9.69747
R22856 a_n7464_n776.n99 a_n7464_n776.n88 9.69747
R22857 a_n7464_n776.n67 a_n7464_n776.n56 9.69747
R22858 a_n7464_n776.n139 a_n7464_n776.n7 9.45567
R22859 a_n7464_n776.n37 a_n7464_n776.n5 9.45567
R22860 a_n7464_n776.n110 a_n7464_n776.n2 9.45567
R22861 a_n7464_n776.n78 a_n7464_n776.n0 9.45567
R22862 a_n7464_n776.n120 a_n7464_n776.n6 9.3005
R22863 a_n7464_n776.n6 a_n7464_n776.n126 9.3005
R22864 a_n7464_n776.n127 a_n7464_n776.n7 9.3005
R22865 a_n7464_n776.n117 a_n7464_n776.n7 9.3005
R22866 a_n7464_n776.n7 a_n7464_n776.n132 9.3005
R22867 a_n7464_n776.n133 a_n7464_n776.n7 9.3005
R22868 a_n7464_n776.n114 a_n7464_n776.n7 9.3005
R22869 a_n7464_n776.n7 a_n7464_n776.n138 9.3005
R22870 a_n7464_n776.n18 a_n7464_n776.n4 9.3005
R22871 a_n7464_n776.n4 a_n7464_n776.n24 9.3005
R22872 a_n7464_n776.n25 a_n7464_n776.n5 9.3005
R22873 a_n7464_n776.n15 a_n7464_n776.n5 9.3005
R22874 a_n7464_n776.n5 a_n7464_n776.n30 9.3005
R22875 a_n7464_n776.n31 a_n7464_n776.n5 9.3005
R22876 a_n7464_n776.n12 a_n7464_n776.n5 9.3005
R22877 a_n7464_n776.n5 a_n7464_n776.n36 9.3005
R22878 a_n7464_n776.n91 a_n7464_n776.n3 9.3005
R22879 a_n7464_n776.n3 a_n7464_n776.n97 9.3005
R22880 a_n7464_n776.n98 a_n7464_n776.n3 9.3005
R22881 a_n7464_n776.n88 a_n7464_n776.n3 9.3005
R22882 a_n7464_n776.n3 a_n7464_n776.n103 9.3005
R22883 a_n7464_n776.n104 a_n7464_n776.n3 9.3005
R22884 a_n7464_n776.n85 a_n7464_n776.n2 9.3005
R22885 a_n7464_n776.n2 a_n7464_n776.n109 9.3005
R22886 a_n7464_n776.n59 a_n7464_n776.n1 9.3005
R22887 a_n7464_n776.n1 a_n7464_n776.n65 9.3005
R22888 a_n7464_n776.n66 a_n7464_n776.n1 9.3005
R22889 a_n7464_n776.n56 a_n7464_n776.n1 9.3005
R22890 a_n7464_n776.n1 a_n7464_n776.n71 9.3005
R22891 a_n7464_n776.n72 a_n7464_n776.n1 9.3005
R22892 a_n7464_n776.n53 a_n7464_n776.n0 9.3005
R22893 a_n7464_n776.n0 a_n7464_n776.n77 9.3005
R22894 a_n7464_n776.n127 a_n7464_n776.n119 8.92171
R22895 a_n7464_n776.n25 a_n7464_n776.n17 8.92171
R22896 a_n7464_n776.n98 a_n7464_n776.n90 8.92171
R22897 a_n7464_n776.n66 a_n7464_n776.n58 8.92171
R22898 a_n7464_n776.n139 a_n7464_n776.n113 8.2187
R22899 a_n7464_n776.n37 a_n7464_n776.n11 8.2187
R22900 a_n7464_n776.n110 a_n7464_n776.n84 8.2187
R22901 a_n7464_n776.n78 a_n7464_n776.n52 8.2187
R22902 a_n7464_n776.n126 a_n7464_n776.n125 8.14595
R22903 a_n7464_n776.n24 a_n7464_n776.n23 8.14595
R22904 a_n7464_n776.n97 a_n7464_n776.n96 8.14595
R22905 a_n7464_n776.n65 a_n7464_n776.n64 8.14595
R22906 a_n7464_n776.n49 a_n7464_n776.n47 8.04791
R22907 a_n7464_n776.n122 a_n7464_n776.n120 7.3702
R22908 a_n7464_n776.n20 a_n7464_n776.n18 7.3702
R22909 a_n7464_n776.n93 a_n7464_n776.n91 7.3702
R22910 a_n7464_n776.n61 a_n7464_n776.n59 7.3702
R22911 a_n7464_n776.n112 a_n7464_n776.n111 6.47248
R22912 a_n7464_n776.n112 a_n7464_n776.n10 6.26581
R22913 a_n7464_n776.n125 a_n7464_n776.n120 5.81868
R22914 a_n7464_n776.n23 a_n7464_n776.n18 5.81868
R22915 a_n7464_n776.n96 a_n7464_n776.n91 5.81868
R22916 a_n7464_n776.n64 a_n7464_n776.n59 5.81868
R22917 a_n7464_n776.n138 a_n7464_n776.n113 5.3904
R22918 a_n7464_n776.n36 a_n7464_n776.n11 5.3904
R22919 a_n7464_n776.n109 a_n7464_n776.n84 5.3904
R22920 a_n7464_n776.n77 a_n7464_n776.n52 5.3904
R22921 a_n7464_n776.n126 a_n7464_n776.n119 5.04292
R22922 a_n7464_n776.n24 a_n7464_n776.n17 5.04292
R22923 a_n7464_n776.n97 a_n7464_n776.n90 5.04292
R22924 a_n7464_n776.n65 a_n7464_n776.n58 5.04292
R22925 a_n7464_n776.n47 a_n7464_n776.n46 4.8472
R22926 a_n7464_n776.n128 a_n7464_n776.n127 4.26717
R22927 a_n7464_n776.n26 a_n7464_n776.n25 4.26717
R22928 a_n7464_n776.n99 a_n7464_n776.n98 4.26717
R22929 a_n7464_n776.n67 a_n7464_n776.n66 4.26717
R22930 a_n7464_n776.n131 a_n7464_n776.n117 3.49141
R22931 a_n7464_n776.n29 a_n7464_n776.n15 3.49141
R22932 a_n7464_n776.n102 a_n7464_n776.n88 3.49141
R22933 a_n7464_n776.n70 a_n7464_n776.n56 3.49141
R22934 a_n7464_n776.n51 a_n7464_n776.n49 3.15136
R22935 a_n7464_n776.n79 a_n7464_n776.n51 3.15136
R22936 a_n7464_n776.n83 a_n7464_n776.n81 3.15136
R22937 a_n7464_n776.n111 a_n7464_n776.n83 3.15136
R22938 a_n7464_n776.n42 a_n7464_n776.n40 3.15136
R22939 a_n7464_n776.n40 a_n7464_n776.n38 3.15136
R22940 a_n7464_n776.n141 a_n7464_n776.n9 3.15136
R22941 a_n7464_n776.n141 a_n7464_n776.n140 3.15136
R22942 a_n7464_n776.n121 a_n7464_n776.n6 2.84305
R22943 a_n7464_n776.n19 a_n7464_n776.n4 2.84305
R22944 a_n7464_n776.n92 a_n7464_n776.n3 2.84305
R22945 a_n7464_n776.n60 a_n7464_n776.n1 2.84305
R22946 a_n7464_n776.n8 a_n7464_n776.t22 2.76201
R22947 a_n7464_n776.n8 a_n7464_n776.t15 2.76201
R22948 a_n7464_n776.n39 a_n7464_n776.t12 2.76201
R22949 a_n7464_n776.n39 a_n7464_n776.t10 2.76201
R22950 a_n7464_n776.n41 a_n7464_n776.t1 2.76201
R22951 a_n7464_n776.n41 a_n7464_n776.t2 2.76201
R22952 a_n7464_n776.n82 a_n7464_n776.t14 2.76201
R22953 a_n7464_n776.n82 a_n7464_n776.t4 2.76201
R22954 a_n7464_n776.n80 a_n7464_n776.t0 2.76201
R22955 a_n7464_n776.n80 a_n7464_n776.t13 2.76201
R22956 a_n7464_n776.n50 a_n7464_n776.t21 2.76201
R22957 a_n7464_n776.n50 a_n7464_n776.t19 2.76201
R22958 a_n7464_n776.n48 a_n7464_n776.t18 2.76201
R22959 a_n7464_n776.n48 a_n7464_n776.t17 2.76201
R22960 a_n7464_n776.n142 a_n7464_n776.t16 2.76201
R22961 a_n7464_n776.t23 a_n7464_n776.n142 2.76201
R22962 a_n7464_n776.n132 a_n7464_n776.n116 2.71565
R22963 a_n7464_n776.n30 a_n7464_n776.n14 2.71565
R22964 a_n7464_n776.n103 a_n7464_n776.n87 2.71565
R22965 a_n7464_n776.n71 a_n7464_n776.n55 2.71565
R22966 a_n7464_n776.n134 a_n7464_n776.n133 1.93989
R22967 a_n7464_n776.n32 a_n7464_n776.n31 1.93989
R22968 a_n7464_n776.n105 a_n7464_n776.n104 1.93989
R22969 a_n7464_n776.n73 a_n7464_n776.n72 1.93989
R22970 a_n7464_n776.n81 a_n7464_n776.n79 1.81084
R22971 a_n7464_n776.n38 a_n7464_n776.n9 1.81084
R22972 a_n7464_n776.n46 a_n7464_n776.n45 1.56155
R22973 a_n7464_n776.n45 a_n7464_n776.n44 1.56155
R22974 a_n7464_n776.n44 a_n7464_n776.n43 1.56155
R22975 a_n7464_n776.n43 a_n7464_n776.n10 1.56155
R22976 a_n7464_n776.n137 a_n7464_n776.n114 1.16414
R22977 a_n7464_n776.n35 a_n7464_n776.n12 1.16414
R22978 a_n7464_n776.n108 a_n7464_n776.n85 1.16414
R22979 a_n7464_n776.n76 a_n7464_n776.n53 1.16414
R22980 a_n7464_n776.n7 a_n7464_n776.n6 1.08671
R22981 a_n7464_n776.n5 a_n7464_n776.n4 1.08671
R22982 a_n7464_n776.n3 a_n7464_n776.n2 1.08671
R22983 a_n7464_n776.n1 a_n7464_n776.n0 1.08671
R22984 a_n11384_10929.n6 a_n11384_10929.n5 215.486
R22985 a_n11384_10929.n6 a_n11384_10929.n4 210.219
R22986 a_n11384_10929.n0 a_n11384_10929.t2 181.262
R22987 a_n11384_10929.n0 a_n11384_10929.t6 178.565
R22988 a_n11384_10929.n0 a_n11384_10929.t3 178.565
R22989 a_n11384_10929.t7 a_n11384_10929.n1 178.565
R22990 a_n11384_10929.n1 a_n11384_10929.n3 164.245
R22991 a_n11384_10929.n0 a_n11384_10929.n2 164.245
R22992 a_n11384_10929.n3 a_n11384_10929.t5 14.3199
R22993 a_n11384_10929.n3 a_n11384_10929.t1 14.3199
R22994 a_n11384_10929.n2 a_n11384_10929.t4 14.3199
R22995 a_n11384_10929.n2 a_n11384_10929.t0 14.3199
R22996 a_n11384_10929.n4 a_n11384_10929.t9 14.3199
R22997 a_n11384_10929.n4 a_n11384_10929.t8 14.3199
R22998 a_n11384_10929.n5 a_n11384_10929.t10 14.3199
R22999 a_n11384_10929.n5 a_n11384_10929.t11 14.3199
R23000 a_n11384_10929.n1 a_n11384_10929.n0 8.78175
R23001 a_n11384_10929.n1 a_n11384_10929.n6 6.35395
R23002 VP.n190 VP.t2 243.97
R23003 VP.n191 VP.t1 243.255
R23004 VP.n190 VP.n189 223.454
R23005 VP.n119 VP.n116 161.3
R23006 VP.n121 VP.n120 161.3
R23007 VP.n122 VP.n115 161.3
R23008 VP.n124 VP.n123 161.3
R23009 VP.n125 VP.n114 161.3
R23010 VP.n127 VP.n126 161.3
R23011 VP.n128 VP.n113 161.3
R23012 VP.n130 VP.n129 161.3
R23013 VP.n131 VP.n112 161.3
R23014 VP.n133 VP.n132 161.3
R23015 VP.n134 VP.n111 161.3
R23016 VP.n136 VP.n135 161.3
R23017 VP.n137 VP.n110 161.3
R23018 VP.n139 VP.n138 161.3
R23019 VP.n140 VP.n109 161.3
R23020 VP.n143 VP.n142 161.3
R23021 VP.n144 VP.n108 161.3
R23022 VP.n146 VP.n145 161.3
R23023 VP.n147 VP.n107 161.3
R23024 VP.n149 VP.n148 161.3
R23025 VP.n150 VP.n106 161.3
R23026 VP.n152 VP.n151 161.3
R23027 VP.n153 VP.n105 161.3
R23028 VP.n155 VP.n154 161.3
R23029 VP.n156 VP.n104 161.3
R23030 VP.n158 VP.n157 161.3
R23031 VP.n159 VP.n103 161.3
R23032 VP.n161 VP.n160 161.3
R23033 VP.n162 VP.n102 161.3
R23034 VP.n164 VP.n163 161.3
R23035 VP.n166 VP.n101 161.3
R23036 VP.n168 VP.n167 161.3
R23037 VP.n169 VP.n100 161.3
R23038 VP.n171 VP.n170 161.3
R23039 VP.n172 VP.n99 161.3
R23040 VP.n174 VP.n173 161.3
R23041 VP.n175 VP.n98 161.3
R23042 VP.n177 VP.n176 161.3
R23043 VP.n178 VP.n97 161.3
R23044 VP.n180 VP.n179 161.3
R23045 VP.n181 VP.n96 161.3
R23046 VP.n183 VP.n182 161.3
R23047 VP.n184 VP.n95 161.3
R23048 VP.n186 VP.n185 161.3
R23049 VP.n92 VP.n91 161.3
R23050 VP.n90 VP.n1 161.3
R23051 VP.n89 VP.n88 161.3
R23052 VP.n87 VP.n2 161.3
R23053 VP.n86 VP.n85 161.3
R23054 VP.n84 VP.n3 161.3
R23055 VP.n83 VP.n82 161.3
R23056 VP.n81 VP.n4 161.3
R23057 VP.n80 VP.n79 161.3
R23058 VP.n78 VP.n5 161.3
R23059 VP.n77 VP.n76 161.3
R23060 VP.n75 VP.n6 161.3
R23061 VP.n74 VP.n73 161.3
R23062 VP.n72 VP.n7 161.3
R23063 VP.n70 VP.n69 161.3
R23064 VP.n68 VP.n8 161.3
R23065 VP.n67 VP.n66 161.3
R23066 VP.n65 VP.n9 161.3
R23067 VP.n64 VP.n63 161.3
R23068 VP.n62 VP.n10 161.3
R23069 VP.n61 VP.n60 161.3
R23070 VP.n59 VP.n11 161.3
R23071 VP.n58 VP.n57 161.3
R23072 VP.n56 VP.n12 161.3
R23073 VP.n55 VP.n54 161.3
R23074 VP.n53 VP.n13 161.3
R23075 VP.n52 VP.n51 161.3
R23076 VP.n50 VP.n14 161.3
R23077 VP.n49 VP.n48 161.3
R23078 VP.n46 VP.n15 161.3
R23079 VP.n45 VP.n44 161.3
R23080 VP.n43 VP.n16 161.3
R23081 VP.n42 VP.n41 161.3
R23082 VP.n40 VP.n17 161.3
R23083 VP.n39 VP.n38 161.3
R23084 VP.n37 VP.n18 161.3
R23085 VP.n36 VP.n35 161.3
R23086 VP.n34 VP.n19 161.3
R23087 VP.n33 VP.n32 161.3
R23088 VP.n31 VP.n20 161.3
R23089 VP.n30 VP.n29 161.3
R23090 VP.n28 VP.n21 161.3
R23091 VP.n27 VP.n26 161.3
R23092 VP.n25 VP.n22 161.3
R23093 VP.n118 VP.n117 72.9837
R23094 VP.n24 VP.n23 72.9837
R23095 VP.n188 VP.n187 59.6618
R23096 VP.n187 VP.n94 58.5146
R23097 VP.n93 VP.n0 58.5146
R23098 VP.n24 VP.t11 58.337
R23099 VP.n118 VP.t7 58.3365
R23100 VP.n177 VP.n98 56.5193
R23101 VP.n83 VP.n4 56.5193
R23102 VP.n153 VP.n152 49.7204
R23103 VP.n129 VP.n112 49.7204
R23104 VP.n35 VP.n18 49.7204
R23105 VP.n59 VP.n58 49.7204
R23106 VP.n154 VP.n153 31.2664
R23107 VP.n129 VP.n128 31.2664
R23108 VP.n35 VP.n34 31.2664
R23109 VP.n60 VP.n59 31.2664
R23110 VP.n94 VP.t12 24.7565
R23111 VP.n165 VP.t13 24.7565
R23112 VP.n141 VP.t6 24.7565
R23113 VP.n117 VP.t8 24.7565
R23114 VP.n23 VP.t5 24.7565
R23115 VP.n47 VP.t4 24.7565
R23116 VP.n71 VP.t10 24.7565
R23117 VP.n0 VP.t9 24.7565
R23118 VP.n185 VP.n184 24.4675
R23119 VP.n184 VP.n183 24.4675
R23120 VP.n183 VP.n96 24.4675
R23121 VP.n179 VP.n96 24.4675
R23122 VP.n179 VP.n178 24.4675
R23123 VP.n178 VP.n177 24.4675
R23124 VP.n173 VP.n98 24.4675
R23125 VP.n173 VP.n172 24.4675
R23126 VP.n172 VP.n171 24.4675
R23127 VP.n171 VP.n100 24.4675
R23128 VP.n167 VP.n100 24.4675
R23129 VP.n167 VP.n166 24.4675
R23130 VP.n164 VP.n102 24.4675
R23131 VP.n160 VP.n102 24.4675
R23132 VP.n160 VP.n159 24.4675
R23133 VP.n159 VP.n158 24.4675
R23134 VP.n158 VP.n104 24.4675
R23135 VP.n154 VP.n104 24.4675
R23136 VP.n152 VP.n106 24.4675
R23137 VP.n148 VP.n106 24.4675
R23138 VP.n148 VP.n147 24.4675
R23139 VP.n147 VP.n146 24.4675
R23140 VP.n146 VP.n108 24.4675
R23141 VP.n142 VP.n108 24.4675
R23142 VP.n140 VP.n139 24.4675
R23143 VP.n139 VP.n110 24.4675
R23144 VP.n135 VP.n110 24.4675
R23145 VP.n135 VP.n134 24.4675
R23146 VP.n134 VP.n133 24.4675
R23147 VP.n133 VP.n112 24.4675
R23148 VP.n128 VP.n127 24.4675
R23149 VP.n127 VP.n114 24.4675
R23150 VP.n123 VP.n114 24.4675
R23151 VP.n123 VP.n122 24.4675
R23152 VP.n122 VP.n121 24.4675
R23153 VP.n121 VP.n116 24.4675
R23154 VP.n27 VP.n22 24.4675
R23155 VP.n28 VP.n27 24.4675
R23156 VP.n29 VP.n28 24.4675
R23157 VP.n29 VP.n20 24.4675
R23158 VP.n33 VP.n20 24.4675
R23159 VP.n34 VP.n33 24.4675
R23160 VP.n39 VP.n18 24.4675
R23161 VP.n40 VP.n39 24.4675
R23162 VP.n41 VP.n40 24.4675
R23163 VP.n41 VP.n16 24.4675
R23164 VP.n45 VP.n16 24.4675
R23165 VP.n46 VP.n45 24.4675
R23166 VP.n48 VP.n14 24.4675
R23167 VP.n52 VP.n14 24.4675
R23168 VP.n53 VP.n52 24.4675
R23169 VP.n54 VP.n53 24.4675
R23170 VP.n54 VP.n12 24.4675
R23171 VP.n58 VP.n12 24.4675
R23172 VP.n60 VP.n10 24.4675
R23173 VP.n64 VP.n10 24.4675
R23174 VP.n65 VP.n64 24.4675
R23175 VP.n66 VP.n65 24.4675
R23176 VP.n66 VP.n8 24.4675
R23177 VP.n70 VP.n8 24.4675
R23178 VP.n73 VP.n72 24.4675
R23179 VP.n73 VP.n6 24.4675
R23180 VP.n77 VP.n6 24.4675
R23181 VP.n78 VP.n77 24.4675
R23182 VP.n79 VP.n78 24.4675
R23183 VP.n79 VP.n4 24.4675
R23184 VP.n84 VP.n83 24.4675
R23185 VP.n85 VP.n84 24.4675
R23186 VP.n85 VP.n2 24.4675
R23187 VP.n89 VP.n2 24.4675
R23188 VP.n90 VP.n89 24.4675
R23189 VP.n91 VP.n90 24.4675
R23190 VP.n166 VP.n165 21.5315
R23191 VP.n72 VP.n71 21.5315
R23192 VP.n189 VP.t0 19.8005
R23193 VP.n189 VP.t3 19.8005
R23194 VP.n185 VP.n94 18.1061
R23195 VP.n91 VP.n0 18.1061
R23196 VP.n188 VP.n93 15.2755
R23197 VP.n142 VP.n141 12.234
R23198 VP.n141 VP.n140 12.234
R23199 VP.n47 VP.n46 12.234
R23200 VP.n48 VP.n47 12.234
R23201 VP VP.n192 11.5771
R23202 VP.n192 VP.n191 4.80222
R23203 VP.n165 VP.n164 2.93654
R23204 VP.n117 VP.n116 2.93654
R23205 VP.n23 VP.n22 2.93654
R23206 VP.n71 VP.n70 2.93654
R23207 VP.n192 VP.n188 0.972091
R23208 VP.n25 VP.n24 0.780565
R23209 VP.n119 VP.n118 0.780562
R23210 VP.n191 VP.n190 0.716017
R23211 VP.n187 VP.n186 0.529113
R23212 VP.n93 VP.n92 0.529113
R23213 VP.n186 VP.n95 0.189894
R23214 VP.n182 VP.n95 0.189894
R23215 VP.n182 VP.n181 0.189894
R23216 VP.n181 VP.n180 0.189894
R23217 VP.n180 VP.n97 0.189894
R23218 VP.n176 VP.n97 0.189894
R23219 VP.n176 VP.n175 0.189894
R23220 VP.n175 VP.n174 0.189894
R23221 VP.n174 VP.n99 0.189894
R23222 VP.n170 VP.n99 0.189894
R23223 VP.n170 VP.n169 0.189894
R23224 VP.n169 VP.n168 0.189894
R23225 VP.n168 VP.n101 0.189894
R23226 VP.n163 VP.n101 0.189894
R23227 VP.n163 VP.n162 0.189894
R23228 VP.n162 VP.n161 0.189894
R23229 VP.n161 VP.n103 0.189894
R23230 VP.n157 VP.n103 0.189894
R23231 VP.n157 VP.n156 0.189894
R23232 VP.n156 VP.n155 0.189894
R23233 VP.n155 VP.n105 0.189894
R23234 VP.n151 VP.n105 0.189894
R23235 VP.n151 VP.n150 0.189894
R23236 VP.n150 VP.n149 0.189894
R23237 VP.n149 VP.n107 0.189894
R23238 VP.n145 VP.n107 0.189894
R23239 VP.n145 VP.n144 0.189894
R23240 VP.n144 VP.n143 0.189894
R23241 VP.n143 VP.n109 0.189894
R23242 VP.n138 VP.n109 0.189894
R23243 VP.n138 VP.n137 0.189894
R23244 VP.n137 VP.n136 0.189894
R23245 VP.n136 VP.n111 0.189894
R23246 VP.n132 VP.n111 0.189894
R23247 VP.n132 VP.n131 0.189894
R23248 VP.n131 VP.n130 0.189894
R23249 VP.n130 VP.n113 0.189894
R23250 VP.n126 VP.n113 0.189894
R23251 VP.n126 VP.n125 0.189894
R23252 VP.n125 VP.n124 0.189894
R23253 VP.n124 VP.n115 0.189894
R23254 VP.n120 VP.n115 0.189894
R23255 VP.n120 VP.n119 0.189894
R23256 VP.n26 VP.n25 0.189894
R23257 VP.n26 VP.n21 0.189894
R23258 VP.n30 VP.n21 0.189894
R23259 VP.n31 VP.n30 0.189894
R23260 VP.n32 VP.n31 0.189894
R23261 VP.n32 VP.n19 0.189894
R23262 VP.n36 VP.n19 0.189894
R23263 VP.n37 VP.n36 0.189894
R23264 VP.n38 VP.n37 0.189894
R23265 VP.n38 VP.n17 0.189894
R23266 VP.n42 VP.n17 0.189894
R23267 VP.n43 VP.n42 0.189894
R23268 VP.n44 VP.n43 0.189894
R23269 VP.n44 VP.n15 0.189894
R23270 VP.n49 VP.n15 0.189894
R23271 VP.n50 VP.n49 0.189894
R23272 VP.n51 VP.n50 0.189894
R23273 VP.n51 VP.n13 0.189894
R23274 VP.n55 VP.n13 0.189894
R23275 VP.n56 VP.n55 0.189894
R23276 VP.n57 VP.n56 0.189894
R23277 VP.n57 VP.n11 0.189894
R23278 VP.n61 VP.n11 0.189894
R23279 VP.n62 VP.n61 0.189894
R23280 VP.n63 VP.n62 0.189894
R23281 VP.n63 VP.n9 0.189894
R23282 VP.n67 VP.n9 0.189894
R23283 VP.n68 VP.n67 0.189894
R23284 VP.n69 VP.n68 0.189894
R23285 VP.n69 VP.n7 0.189894
R23286 VP.n74 VP.n7 0.189894
R23287 VP.n75 VP.n74 0.189894
R23288 VP.n76 VP.n75 0.189894
R23289 VP.n76 VP.n5 0.189894
R23290 VP.n80 VP.n5 0.189894
R23291 VP.n81 VP.n80 0.189894
R23292 VP.n82 VP.n81 0.189894
R23293 VP.n82 VP.n3 0.189894
R23294 VP.n86 VP.n3 0.189894
R23295 VP.n87 VP.n86 0.189894
R23296 VP.n88 VP.n87 0.189894
R23297 VP.n88 VP.n1 0.189894
R23298 VP.n92 VP.n1 0.189894
C0 VDD VOUT 30.5405f
C1 VOUT VP 2.82844f
C2 VDD VN 0.295246f
C3 a_n12854_10929# VDD 1.81267f
C4 VOUT VN 1.23337f
C5 VOUT CS_BIAS 20.1905f
C6 VP VN 17.263401f
C7 VP CS_BIAS 0.631755f
C8 VN CS_BIAS 0.561641f
C9 VP DIFFPAIR_BIAS 7.75e-19
C10 VN DIFFPAIR_BIAS 0.001896f
C11 a_11512_10929# VDD 1.81267f
C12 DIFFPAIR_BIAS GND 54.876038f
C13 CS_BIAS GND 94.5312f
C14 VN GND 72.70878f
C15 VP GND 55.67877f
C16 VOUT GND 79.35675f
C17 VDD GND 0.889864p
C18 a_11512_10929# GND 1.35906f
C19 a_n12854_10929# GND 1.36714f
C20 VP.t9 GND 1.5212f
C21 VP.n0 GND 0.594179f
C22 VP.n1 GND 0.011375f
C23 VP.n2 GND 0.0212f
C24 VP.n3 GND 0.011375f
C25 VP.n4 GND 0.015497f
C26 VP.n5 GND 0.011375f
C27 VP.n6 GND 0.0212f
C28 VP.n7 GND 0.011375f
C29 VP.t10 GND 1.5212f
C30 VP.n8 GND 0.0212f
C31 VP.n9 GND 0.011375f
C32 VP.n10 GND 0.0212f
C33 VP.n11 GND 0.011375f
C34 VP.n12 GND 0.0212f
C35 VP.n13 GND 0.011375f
C36 VP.n14 GND 0.0212f
C37 VP.n15 GND 0.011375f
C38 VP.t4 GND 1.5212f
C39 VP.n16 GND 0.0212f
C40 VP.n17 GND 0.011375f
C41 VP.n18 GND 0.020987f
C42 VP.n19 GND 0.011375f
C43 VP.n20 GND 0.0212f
C44 VP.n21 GND 0.011375f
C45 VP.n22 GND 0.011989f
C46 VP.t5 GND 1.5212f
C47 VP.n23 GND 0.586354f
C48 VP.t11 GND 1.90055f
C49 VP.n24 GND 0.684358f
C50 VP.n25 GND 0.115124f
C51 VP.n26 GND 0.011375f
C52 VP.n27 GND 0.0212f
C53 VP.n28 GND 0.0212f
C54 VP.n29 GND 0.0212f
C55 VP.n30 GND 0.011375f
C56 VP.n31 GND 0.011375f
C57 VP.n32 GND 0.011375f
C58 VP.n33 GND 0.0212f
C59 VP.n34 GND 0.022839f
C60 VP.n35 GND 0.010587f
C61 VP.n36 GND 0.011375f
C62 VP.n37 GND 0.011375f
C63 VP.n38 GND 0.011375f
C64 VP.n39 GND 0.0212f
C65 VP.n40 GND 0.0212f
C66 VP.n41 GND 0.0212f
C67 VP.n42 GND 0.011375f
C68 VP.n43 GND 0.011375f
C69 VP.n44 GND 0.011375f
C70 VP.n45 GND 0.0212f
C71 VP.n46 GND 0.015967f
C72 VP.n47 GND 0.542256f
C73 VP.n48 GND 0.015967f
C74 VP.n49 GND 0.011375f
C75 VP.n50 GND 0.011375f
C76 VP.n51 GND 0.011375f
C77 VP.n52 GND 0.0212f
C78 VP.n53 GND 0.0212f
C79 VP.n54 GND 0.0212f
C80 VP.n55 GND 0.011375f
C81 VP.n56 GND 0.011375f
C82 VP.n57 GND 0.011375f
C83 VP.n58 GND 0.020987f
C84 VP.n59 GND 0.010587f
C85 VP.n60 GND 0.022839f
C86 VP.n61 GND 0.011375f
C87 VP.n62 GND 0.011375f
C88 VP.n63 GND 0.011375f
C89 VP.n64 GND 0.0212f
C90 VP.n65 GND 0.0212f
C91 VP.n66 GND 0.0212f
C92 VP.n67 GND 0.011375f
C93 VP.n68 GND 0.011375f
C94 VP.n69 GND 0.011375f
C95 VP.n70 GND 0.011989f
C96 VP.n71 GND 0.542256f
C97 VP.n72 GND 0.019944f
C98 VP.n73 GND 0.0212f
C99 VP.n74 GND 0.011375f
C100 VP.n75 GND 0.011375f
C101 VP.n76 GND 0.011375f
C102 VP.n77 GND 0.0212f
C103 VP.n78 GND 0.0212f
C104 VP.n79 GND 0.0212f
C105 VP.n80 GND 0.011375f
C106 VP.n81 GND 0.011375f
C107 VP.n82 GND 0.011375f
C108 VP.n83 GND 0.017716f
C109 VP.n84 GND 0.0212f
C110 VP.n85 GND 0.0212f
C111 VP.n86 GND 0.011375f
C112 VP.n87 GND 0.011375f
C113 VP.n88 GND 0.011375f
C114 VP.n89 GND 0.0212f
C115 VP.n90 GND 0.0212f
C116 VP.n91 GND 0.018479f
C117 VP.n92 GND 0.028294f
C118 VP.n93 GND 0.322699f
C119 VP.t12 GND 1.5212f
C120 VP.n94 GND 0.594179f
C121 VP.n95 GND 0.011375f
C122 VP.n96 GND 0.0212f
C123 VP.n97 GND 0.011375f
C124 VP.n98 GND 0.015497f
C125 VP.n99 GND 0.011375f
C126 VP.n100 GND 0.0212f
C127 VP.n101 GND 0.011375f
C128 VP.t13 GND 1.5212f
C129 VP.n102 GND 0.0212f
C130 VP.n103 GND 0.011375f
C131 VP.n104 GND 0.0212f
C132 VP.n105 GND 0.011375f
C133 VP.n106 GND 0.0212f
C134 VP.n107 GND 0.011375f
C135 VP.n108 GND 0.0212f
C136 VP.n109 GND 0.011375f
C137 VP.t6 GND 1.5212f
C138 VP.n110 GND 0.0212f
C139 VP.n111 GND 0.011375f
C140 VP.n112 GND 0.020987f
C141 VP.n113 GND 0.011375f
C142 VP.n114 GND 0.0212f
C143 VP.n115 GND 0.011375f
C144 VP.n116 GND 0.011989f
C145 VP.t7 GND 1.90055f
C146 VP.t8 GND 1.5212f
C147 VP.n117 GND 0.586354f
C148 VP.n118 GND 0.684362f
C149 VP.n119 GND 0.115124f
C150 VP.n120 GND 0.011375f
C151 VP.n121 GND 0.0212f
C152 VP.n122 GND 0.0212f
C153 VP.n123 GND 0.0212f
C154 VP.n124 GND 0.011375f
C155 VP.n125 GND 0.011375f
C156 VP.n126 GND 0.011375f
C157 VP.n127 GND 0.0212f
C158 VP.n128 GND 0.022839f
C159 VP.n129 GND 0.010587f
C160 VP.n130 GND 0.011375f
C161 VP.n131 GND 0.011375f
C162 VP.n132 GND 0.011375f
C163 VP.n133 GND 0.0212f
C164 VP.n134 GND 0.0212f
C165 VP.n135 GND 0.0212f
C166 VP.n136 GND 0.011375f
C167 VP.n137 GND 0.011375f
C168 VP.n138 GND 0.011375f
C169 VP.n139 GND 0.0212f
C170 VP.n140 GND 0.015967f
C171 VP.n141 GND 0.542256f
C172 VP.n142 GND 0.015967f
C173 VP.n143 GND 0.011375f
C174 VP.n144 GND 0.011375f
C175 VP.n145 GND 0.011375f
C176 VP.n146 GND 0.0212f
C177 VP.n147 GND 0.0212f
C178 VP.n148 GND 0.0212f
C179 VP.n149 GND 0.011375f
C180 VP.n150 GND 0.011375f
C181 VP.n151 GND 0.011375f
C182 VP.n152 GND 0.020987f
C183 VP.n153 GND 0.010587f
C184 VP.n154 GND 0.022839f
C185 VP.n155 GND 0.011375f
C186 VP.n156 GND 0.011375f
C187 VP.n157 GND 0.011375f
C188 VP.n158 GND 0.0212f
C189 VP.n159 GND 0.0212f
C190 VP.n160 GND 0.0212f
C191 VP.n161 GND 0.011375f
C192 VP.n162 GND 0.011375f
C193 VP.n163 GND 0.011375f
C194 VP.n164 GND 0.011989f
C195 VP.n165 GND 0.542256f
C196 VP.n166 GND 0.019944f
C197 VP.n167 GND 0.0212f
C198 VP.n168 GND 0.011375f
C199 VP.n169 GND 0.011375f
C200 VP.n170 GND 0.011375f
C201 VP.n171 GND 0.0212f
C202 VP.n172 GND 0.0212f
C203 VP.n173 GND 0.0212f
C204 VP.n174 GND 0.011375f
C205 VP.n175 GND 0.011375f
C206 VP.n176 GND 0.011375f
C207 VP.n177 GND 0.017716f
C208 VP.n178 GND 0.0212f
C209 VP.n179 GND 0.0212f
C210 VP.n180 GND 0.011375f
C211 VP.n181 GND 0.011375f
C212 VP.n182 GND 0.011375f
C213 VP.n183 GND 0.0212f
C214 VP.n184 GND 0.0212f
C215 VP.n185 GND 0.018479f
C216 VP.n186 GND 0.028294f
C217 VP.n187 GND 0.966526f
C218 VP.n188 GND 1.11203f
C219 VP.t2 GND 0.019636f
C220 VP.t0 GND 0.003507f
C221 VP.t3 GND 0.003507f
C222 VP.n189 GND 0.011372f
C223 VP.n190 GND 0.088284f
C224 VP.t1 GND 0.019517f
C225 VP.n191 GND 0.052963f
C226 VP.n192 GND 0.723621f
C227 a_n11384_10929.n0 GND 3.55508f
C228 a_n11384_10929.n1 GND 2.51726f
C229 a_n11384_10929.t2 GND 0.182684f
C230 a_n11384_10929.t4 GND 0.026687f
C231 a_n11384_10929.t0 GND 0.026687f
C232 a_n11384_10929.n2 GND 0.112037f
C233 a_n11384_10929.t3 GND 0.172139f
C234 a_n11384_10929.t6 GND 0.172139f
C235 a_n11384_10929.t5 GND 0.026687f
C236 a_n11384_10929.t1 GND 0.026687f
C237 a_n11384_10929.n3 GND 0.112037f
C238 a_n11384_10929.t9 GND 0.026687f
C239 a_n11384_10929.t8 GND 0.026687f
C240 a_n11384_10929.n4 GND 0.448985f
C241 a_n11384_10929.t10 GND 0.026687f
C242 a_n11384_10929.t11 GND 0.026687f
C243 a_n11384_10929.n5 GND 0.861407f
C244 a_n11384_10929.n6 GND 13.480599f
C245 a_n11384_10929.t7 GND 0.172138f
C246 a_n7464_n776.n0 GND 0.027698f
C247 a_n7464_n776.n1 GND 0.273898f
C248 a_n7464_n776.n2 GND 0.027698f
C249 a_n7464_n776.n3 GND 0.273898f
C250 a_n7464_n776.n4 GND 0.241639f
C251 a_n7464_n776.n5 GND 0.059957f
C252 a_n7464_n776.n6 GND 0.241639f
C253 a_n7464_n776.n7 GND 0.059957f
C254 a_n7464_n776.t16 GND 0.045695f
C255 a_n7464_n776.t22 GND 0.045695f
C256 a_n7464_n776.t15 GND 0.045695f
C257 a_n7464_n776.n8 GND 0.379192f
C258 a_n7464_n776.n9 GND 0.584563f
C259 a_n7464_n776.t8 GND 0.351628f
C260 a_n7464_n776.n10 GND 1.77309f
C261 a_n7464_n776.n11 GND 0.010727f
C262 a_n7464_n776.n12 GND 0.004334f
C263 a_n7464_n776.n13 GND 0.010243f
C264 a_n7464_n776.n14 GND 0.004589f
C265 a_n7464_n776.n15 GND 0.004334f
C266 a_n7464_n776.n16 GND 0.010243f
C267 a_n7464_n776.n17 GND 0.004589f
C268 a_n7464_n776.n18 GND 0.004334f
C269 a_n7464_n776.t11 GND 0.0171f
C270 a_n7464_n776.n19 GND 0.043208f
C271 a_n7464_n776.n20 GND 0.007241f
C272 a_n7464_n776.n21 GND 0.007682f
C273 a_n7464_n776.n22 GND 0.010243f
C274 a_n7464_n776.n23 GND 0.004589f
C275 a_n7464_n776.n24 GND 0.004334f
C276 a_n7464_n776.n25 GND 0.004334f
C277 a_n7464_n776.n26 GND 0.004589f
C278 a_n7464_n776.n27 GND 0.010243f
C279 a_n7464_n776.n28 GND 0.010243f
C280 a_n7464_n776.n29 GND 0.004589f
C281 a_n7464_n776.n30 GND 0.004334f
C282 a_n7464_n776.n31 GND 0.004334f
C283 a_n7464_n776.n32 GND 0.004589f
C284 a_n7464_n776.n33 GND 0.010243f
C285 a_n7464_n776.n34 GND 0.020664f
C286 a_n7464_n776.n35 GND 0.004589f
C287 a_n7464_n776.n36 GND 0.008474f
C288 a_n7464_n776.n37 GND 0.022804f
C289 a_n7464_n776.n38 GND 0.524965f
C290 a_n7464_n776.t12 GND 0.045695f
C291 a_n7464_n776.t10 GND 0.045695f
C292 a_n7464_n776.n39 GND 0.379192f
C293 a_n7464_n776.n40 GND 0.723906f
C294 a_n7464_n776.t1 GND 0.045695f
C295 a_n7464_n776.t2 GND 0.045695f
C296 a_n7464_n776.n41 GND 0.379192f
C297 a_n7464_n776.n42 GND 1.17212f
C298 a_n7464_n776.t9 GND 0.351628f
C299 a_n7464_n776.n43 GND 0.813636f
C300 a_n7464_n776.t6 GND 0.351628f
C301 a_n7464_n776.n44 GND 0.813636f
C302 a_n7464_n776.t7 GND 0.351628f
C303 a_n7464_n776.n45 GND 0.813636f
C304 a_n7464_n776.t5 GND 0.351628f
C305 a_n7464_n776.n46 GND 1.41504f
C306 a_n7464_n776.n47 GND 1.13303f
C307 a_n7464_n776.t18 GND 0.045695f
C308 a_n7464_n776.t17 GND 0.045695f
C309 a_n7464_n776.n48 GND 0.379189f
C310 a_n7464_n776.n49 GND 0.976712f
C311 a_n7464_n776.t21 GND 0.045695f
C312 a_n7464_n776.t19 GND 0.045695f
C313 a_n7464_n776.n50 GND 0.379189f
C314 a_n7464_n776.n51 GND 0.723909f
C315 a_n7464_n776.n52 GND 0.010727f
C316 a_n7464_n776.n53 GND 0.004334f
C317 a_n7464_n776.n54 GND 0.010243f
C318 a_n7464_n776.n55 GND 0.004589f
C319 a_n7464_n776.n56 GND 0.004334f
C320 a_n7464_n776.n57 GND 0.010243f
C321 a_n7464_n776.n58 GND 0.004589f
C322 a_n7464_n776.n59 GND 0.004334f
C323 a_n7464_n776.t20 GND 0.0171f
C324 a_n7464_n776.n60 GND 0.043208f
C325 a_n7464_n776.n61 GND 0.007241f
C326 a_n7464_n776.n62 GND 0.007682f
C327 a_n7464_n776.n63 GND 0.010243f
C328 a_n7464_n776.n64 GND 0.004589f
C329 a_n7464_n776.n65 GND 0.004334f
C330 a_n7464_n776.n66 GND 0.004334f
C331 a_n7464_n776.n67 GND 0.004589f
C332 a_n7464_n776.n68 GND 0.010243f
C333 a_n7464_n776.n69 GND 0.010243f
C334 a_n7464_n776.n70 GND 0.004589f
C335 a_n7464_n776.n71 GND 0.004334f
C336 a_n7464_n776.n72 GND 0.004334f
C337 a_n7464_n776.n73 GND 0.004589f
C338 a_n7464_n776.n74 GND 0.010243f
C339 a_n7464_n776.n75 GND 0.020664f
C340 a_n7464_n776.n76 GND 0.004589f
C341 a_n7464_n776.n77 GND 0.008474f
C342 a_n7464_n776.n78 GND 0.022804f
C343 a_n7464_n776.n79 GND 0.524965f
C344 a_n7464_n776.t0 GND 0.045695f
C345 a_n7464_n776.t13 GND 0.045695f
C346 a_n7464_n776.n80 GND 0.379189f
C347 a_n7464_n776.n81 GND 0.584566f
C348 a_n7464_n776.t14 GND 0.045695f
C349 a_n7464_n776.t4 GND 0.045695f
C350 a_n7464_n776.n82 GND 0.379189f
C351 a_n7464_n776.n83 GND 0.723909f
C352 a_n7464_n776.n84 GND 0.010727f
C353 a_n7464_n776.n85 GND 0.004334f
C354 a_n7464_n776.n86 GND 0.010243f
C355 a_n7464_n776.n87 GND 0.004589f
C356 a_n7464_n776.n88 GND 0.004334f
C357 a_n7464_n776.n89 GND 0.010243f
C358 a_n7464_n776.n90 GND 0.004589f
C359 a_n7464_n776.n91 GND 0.004334f
C360 a_n7464_n776.t3 GND 0.0171f
C361 a_n7464_n776.n92 GND 0.043208f
C362 a_n7464_n776.n93 GND 0.007241f
C363 a_n7464_n776.n94 GND 0.007682f
C364 a_n7464_n776.n95 GND 0.010243f
C365 a_n7464_n776.n96 GND 0.004589f
C366 a_n7464_n776.n97 GND 0.004334f
C367 a_n7464_n776.n98 GND 0.004334f
C368 a_n7464_n776.n99 GND 0.004589f
C369 a_n7464_n776.n100 GND 0.010243f
C370 a_n7464_n776.n101 GND 0.010243f
C371 a_n7464_n776.n102 GND 0.004589f
C372 a_n7464_n776.n103 GND 0.004334f
C373 a_n7464_n776.n104 GND 0.004334f
C374 a_n7464_n776.n105 GND 0.004589f
C375 a_n7464_n776.n106 GND 0.010243f
C376 a_n7464_n776.n107 GND 0.020664f
C377 a_n7464_n776.n108 GND 0.004589f
C378 a_n7464_n776.n109 GND 0.008474f
C379 a_n7464_n776.n110 GND 0.022804f
C380 a_n7464_n776.n111 GND 0.69099f
C381 a_n7464_n776.n112 GND 1.25151f
C382 a_n7464_n776.n113 GND 0.010727f
C383 a_n7464_n776.n114 GND 0.004334f
C384 a_n7464_n776.n115 GND 0.010243f
C385 a_n7464_n776.n116 GND 0.004589f
C386 a_n7464_n776.n117 GND 0.004334f
C387 a_n7464_n776.n118 GND 0.010243f
C388 a_n7464_n776.n119 GND 0.004589f
C389 a_n7464_n776.n120 GND 0.004334f
C390 a_n7464_n776.t24 GND 0.0171f
C391 a_n7464_n776.n121 GND 0.043208f
C392 a_n7464_n776.n122 GND 0.007241f
C393 a_n7464_n776.n123 GND 0.007682f
C394 a_n7464_n776.n124 GND 0.010243f
C395 a_n7464_n776.n125 GND 0.004589f
C396 a_n7464_n776.n126 GND 0.004334f
C397 a_n7464_n776.n127 GND 0.004334f
C398 a_n7464_n776.n128 GND 0.004589f
C399 a_n7464_n776.n129 GND 0.010243f
C400 a_n7464_n776.n130 GND 0.010243f
C401 a_n7464_n776.n131 GND 0.004589f
C402 a_n7464_n776.n132 GND 0.004334f
C403 a_n7464_n776.n133 GND 0.004334f
C404 a_n7464_n776.n134 GND 0.004589f
C405 a_n7464_n776.n135 GND 0.010243f
C406 a_n7464_n776.n136 GND 0.020664f
C407 a_n7464_n776.n137 GND 0.004589f
C408 a_n7464_n776.n138 GND 0.008474f
C409 a_n7464_n776.n139 GND 0.022804f
C410 a_n7464_n776.n140 GND 0.85547f
C411 a_n7464_n776.n141 GND 0.723911f
C412 a_n7464_n776.n142 GND 0.379187f
C413 a_n7464_n776.t23 GND 0.045695f
C414 DIFFPAIR_BIAS.t11 GND 0.108792f
C415 DIFFPAIR_BIAS.t10 GND 0.104772f
C416 DIFFPAIR_BIAS.n0 GND 0.1437f
C417 DIFFPAIR_BIAS.t3 GND 0.023563f
C418 DIFFPAIR_BIAS.t1 GND 0.022814f
C419 DIFFPAIR_BIAS.n1 GND 0.121226f
C420 DIFFPAIR_BIAS.t5 GND 0.022814f
C421 DIFFPAIR_BIAS.n2 GND 0.062985f
C422 DIFFPAIR_BIAS.t9 GND 0.022814f
C423 DIFFPAIR_BIAS.n3 GND 0.062985f
C424 DIFFPAIR_BIAS.t7 GND 0.022814f
C425 DIFFPAIR_BIAS.n4 GND 0.072295f
C426 DIFFPAIR_BIAS.t2 GND 0.105489f
C427 DIFFPAIR_BIAS.t0 GND 0.102298f
C428 DIFFPAIR_BIAS.n5 GND 0.131841f
C429 DIFFPAIR_BIAS.t4 GND 0.102298f
C430 DIFFPAIR_BIAS.n6 GND 0.071608f
C431 DIFFPAIR_BIAS.t8 GND 0.102298f
C432 DIFFPAIR_BIAS.n7 GND 0.071608f
C433 DIFFPAIR_BIAS.t6 GND 0.102298f
C434 DIFFPAIR_BIAS.n8 GND 0.075748f
C435 DIFFPAIR_BIAS.n9 GND 0.091744f
C436 DIFFPAIR_BIAS.t14 GND 0.104772f
C437 DIFFPAIR_BIAS.n10 GND 0.068876f
C438 DIFFPAIR_BIAS.t12 GND 0.104772f
C439 DIFFPAIR_BIAS.n11 GND 0.074108f
C440 DIFFPAIR_BIAS.t13 GND 0.104772f
C441 DIFFPAIR_BIAS.n12 GND 0.058225f
C442 DIFFPAIR_BIAS.n13 GND 0.036228f
C443 a_n4580_9541.n0 GND 1.04069f
C444 a_n4580_9541.t0 GND 50.9266f
C445 a_n4580_9541.t11 GND 0.1148f
C446 a_n4580_9541.t12 GND 0.108173f
C447 a_n4580_9541.n1 GND 2.82283f
C448 a_n4580_9541.t8 GND 0.1148f
C449 a_n4580_9541.t2 GND 0.01677f
C450 a_n4580_9541.t6 GND 0.01677f
C451 a_n4580_9541.n2 GND 0.070405f
C452 a_n4580_9541.n3 GND 1.19334f
C453 a_n4580_9541.t3 GND 0.108173f
C454 a_n4580_9541.t7 GND 0.108173f
C455 a_n4580_9541.t5 GND 0.01677f
C456 a_n4580_9541.t4 GND 0.01677f
C457 a_n4580_9541.n4 GND 0.070405f
C458 a_n4580_9541.n5 GND 0.754799f
C459 a_n4580_9541.t1 GND 0.108173f
C460 a_n4580_9541.n6 GND 0.827061f
C461 a_n4580_9541.n7 GND 2.48323f
C462 a_n4580_9541.t10 GND 0.114799f
C463 a_n4580_9541.t9 GND 0.108173f
C464 a_n4580_9541.n8 GND 2.35059f
C465 a_n4580_9541.n9 GND 1.60773f
C466 VN.t10 GND 1.09435f
C467 VN.n0 GND 0.42745f
C468 VN.n1 GND 0.008183f
C469 VN.n2 GND 0.015251f
C470 VN.n3 GND 0.008183f
C471 VN.n4 GND 0.011148f
C472 VN.n5 GND 0.008183f
C473 VN.n6 GND 0.015251f
C474 VN.n7 GND 0.008183f
C475 VN.t11 GND 1.09435f
C476 VN.n8 GND 0.015251f
C477 VN.n9 GND 0.008183f
C478 VN.n10 GND 0.015251f
C479 VN.n11 GND 0.008183f
C480 VN.n12 GND 0.015251f
C481 VN.n13 GND 0.008183f
C482 VN.n14 GND 0.015251f
C483 VN.n15 GND 0.008183f
C484 VN.t7 GND 1.09435f
C485 VN.n16 GND 0.015251f
C486 VN.n17 GND 0.008183f
C487 VN.n18 GND 0.015098f
C488 VN.n19 GND 0.008183f
C489 VN.n20 GND 0.015251f
C490 VN.n21 GND 0.008183f
C491 VN.n22 GND 0.008625f
C492 VN.t8 GND 1.36725f
C493 VN.t9 GND 1.09435f
C494 VN.n23 GND 0.421821f
C495 VN.n24 GND 0.492328f
C496 VN.n25 GND 0.08282f
C497 VN.n26 GND 0.008183f
C498 VN.n27 GND 0.015251f
C499 VN.n28 GND 0.015251f
C500 VN.n29 GND 0.015251f
C501 VN.n30 GND 0.008183f
C502 VN.n31 GND 0.008183f
C503 VN.n32 GND 0.008183f
C504 VN.n33 GND 0.015251f
C505 VN.n34 GND 0.01643f
C506 VN.n35 GND 0.007616f
C507 VN.n36 GND 0.008183f
C508 VN.n37 GND 0.008183f
C509 VN.n38 GND 0.008183f
C510 VN.n39 GND 0.015251f
C511 VN.n40 GND 0.015251f
C512 VN.n41 GND 0.015251f
C513 VN.n42 GND 0.008183f
C514 VN.n43 GND 0.008183f
C515 VN.n44 GND 0.008183f
C516 VN.n45 GND 0.015251f
C517 VN.n46 GND 0.011486f
C518 VN.n47 GND 0.390097f
C519 VN.n48 GND 0.011486f
C520 VN.n49 GND 0.008183f
C521 VN.n50 GND 0.008183f
C522 VN.n51 GND 0.008183f
C523 VN.n52 GND 0.015251f
C524 VN.n53 GND 0.015251f
C525 VN.n54 GND 0.015251f
C526 VN.n55 GND 0.008183f
C527 VN.n56 GND 0.008183f
C528 VN.n57 GND 0.008183f
C529 VN.n58 GND 0.015098f
C530 VN.n59 GND 0.007616f
C531 VN.n60 GND 0.01643f
C532 VN.n61 GND 0.008183f
C533 VN.n62 GND 0.008183f
C534 VN.n63 GND 0.008183f
C535 VN.n64 GND 0.015251f
C536 VN.n65 GND 0.015251f
C537 VN.n66 GND 0.015251f
C538 VN.n67 GND 0.008183f
C539 VN.n68 GND 0.008183f
C540 VN.n69 GND 0.008183f
C541 VN.n70 GND 0.008625f
C542 VN.n71 GND 0.390097f
C543 VN.n72 GND 0.014348f
C544 VN.n73 GND 0.015251f
C545 VN.n74 GND 0.008183f
C546 VN.n75 GND 0.008183f
C547 VN.n76 GND 0.008183f
C548 VN.n77 GND 0.015251f
C549 VN.n78 GND 0.015251f
C550 VN.n79 GND 0.015251f
C551 VN.n80 GND 0.008183f
C552 VN.n81 GND 0.008183f
C553 VN.n82 GND 0.008183f
C554 VN.n83 GND 0.012745f
C555 VN.n84 GND 0.015251f
C556 VN.n85 GND 0.015251f
C557 VN.n86 GND 0.008183f
C558 VN.n87 GND 0.008183f
C559 VN.n88 GND 0.008183f
C560 VN.n89 GND 0.015251f
C561 VN.n90 GND 0.015251f
C562 VN.n91 GND 0.013293f
C563 VN.n92 GND 0.020355f
C564 VN.n93 GND 0.230054f
C565 VN.t4 GND 1.09435f
C566 VN.n94 GND 0.42745f
C567 VN.n95 GND 0.008183f
C568 VN.n96 GND 0.015251f
C569 VN.n97 GND 0.008183f
C570 VN.n98 GND 0.011148f
C571 VN.n99 GND 0.008183f
C572 VN.n100 GND 0.015251f
C573 VN.n101 GND 0.008183f
C574 VN.t5 GND 1.09435f
C575 VN.n102 GND 0.015251f
C576 VN.n103 GND 0.008183f
C577 VN.n104 GND 0.015251f
C578 VN.n105 GND 0.008183f
C579 VN.n106 GND 0.015251f
C580 VN.n107 GND 0.008183f
C581 VN.n108 GND 0.015251f
C582 VN.n109 GND 0.008183f
C583 VN.t12 GND 1.09435f
C584 VN.n110 GND 0.015251f
C585 VN.n111 GND 0.008183f
C586 VN.n112 GND 0.015098f
C587 VN.n113 GND 0.008183f
C588 VN.n114 GND 0.015251f
C589 VN.n115 GND 0.008183f
C590 VN.n116 GND 0.008625f
C591 VN.t13 GND 1.09435f
C592 VN.n117 GND 0.421821f
C593 VN.t6 GND 1.36725f
C594 VN.n118 GND 0.492325f
C595 VN.n119 GND 0.08282f
C596 VN.n120 GND 0.008183f
C597 VN.n121 GND 0.015251f
C598 VN.n122 GND 0.015251f
C599 VN.n123 GND 0.015251f
C600 VN.n124 GND 0.008183f
C601 VN.n125 GND 0.008183f
C602 VN.n126 GND 0.008183f
C603 VN.n127 GND 0.015251f
C604 VN.n128 GND 0.01643f
C605 VN.n129 GND 0.007616f
C606 VN.n130 GND 0.008183f
C607 VN.n131 GND 0.008183f
C608 VN.n132 GND 0.008183f
C609 VN.n133 GND 0.015251f
C610 VN.n134 GND 0.015251f
C611 VN.n135 GND 0.015251f
C612 VN.n136 GND 0.008183f
C613 VN.n137 GND 0.008183f
C614 VN.n138 GND 0.008183f
C615 VN.n139 GND 0.015251f
C616 VN.n140 GND 0.011486f
C617 VN.n141 GND 0.390097f
C618 VN.n142 GND 0.011486f
C619 VN.n143 GND 0.008183f
C620 VN.n144 GND 0.008183f
C621 VN.n145 GND 0.008183f
C622 VN.n146 GND 0.015251f
C623 VN.n147 GND 0.015251f
C624 VN.n148 GND 0.015251f
C625 VN.n149 GND 0.008183f
C626 VN.n150 GND 0.008183f
C627 VN.n151 GND 0.008183f
C628 VN.n152 GND 0.015098f
C629 VN.n153 GND 0.007616f
C630 VN.n154 GND 0.01643f
C631 VN.n155 GND 0.008183f
C632 VN.n156 GND 0.008183f
C633 VN.n157 GND 0.008183f
C634 VN.n158 GND 0.015251f
C635 VN.n159 GND 0.015251f
C636 VN.n160 GND 0.015251f
C637 VN.n161 GND 0.008183f
C638 VN.n162 GND 0.008183f
C639 VN.n163 GND 0.008183f
C640 VN.n164 GND 0.008625f
C641 VN.n165 GND 0.390097f
C642 VN.n166 GND 0.014348f
C643 VN.n167 GND 0.015251f
C644 VN.n168 GND 0.008183f
C645 VN.n169 GND 0.008183f
C646 VN.n170 GND 0.008183f
C647 VN.n171 GND 0.015251f
C648 VN.n172 GND 0.015251f
C649 VN.n173 GND 0.015251f
C650 VN.n174 GND 0.008183f
C651 VN.n175 GND 0.008183f
C652 VN.n176 GND 0.008183f
C653 VN.n177 GND 0.012745f
C654 VN.n178 GND 0.015251f
C655 VN.n179 GND 0.015251f
C656 VN.n180 GND 0.008183f
C657 VN.n181 GND 0.008183f
C658 VN.n182 GND 0.008183f
C659 VN.n183 GND 0.015251f
C660 VN.n184 GND 0.015251f
C661 VN.n185 GND 0.013293f
C662 VN.n186 GND 0.020355f
C663 VN.n187 GND 0.692173f
C664 VN.n188 GND 0.796604f
C665 VN.t1 GND 0.014126f
C666 VN.t0 GND 0.002523f
C667 VN.t3 GND 0.002523f
C668 VN.n189 GND 0.008181f
C669 VN.n190 GND 0.063511f
C670 VN.t2 GND 0.01404f
C671 VN.n191 GND 0.04254f
C672 VN.n192 GND 2.16212f
C673 VDD.t95 GND 0.001629f
C674 VDD.t110 GND 0.001629f
C675 VDD.n0 GND 0.009559f
C676 VDD.t108 GND 0.001629f
C677 VDD.t129 GND 0.001629f
C678 VDD.n1 GND 0.008529f
C679 VDD.n2 GND 0.155114f
C680 VDD.t101 GND 0.001629f
C681 VDD.t97 GND 0.001629f
C682 VDD.n3 GND 0.008529f
C683 VDD.n4 GND 0.081723f
C684 VDD.t114 GND 0.001629f
C685 VDD.t140 GND 0.001629f
C686 VDD.n5 GND 0.008529f
C687 VDD.n6 GND 0.066551f
C688 VDD.t112 GND 0.001629f
C689 VDD.t136 GND 0.001629f
C690 VDD.n7 GND 0.009559f
C691 VDD.t131 GND 0.001629f
C692 VDD.t125 GND 0.001629f
C693 VDD.n8 GND 0.008529f
C694 VDD.n9 GND 0.155114f
C695 VDD.t106 GND 0.001629f
C696 VDD.t118 GND 0.001629f
C697 VDD.n10 GND 0.008529f
C698 VDD.n11 GND 0.081723f
C699 VDD.t116 GND 0.001629f
C700 VDD.t122 GND 0.001629f
C701 VDD.n12 GND 0.008529f
C702 VDD.n13 GND 0.066551f
C703 VDD.n14 GND 0.057336f
C704 VDD.n15 GND 0.988416f
C705 VDD.n16 GND 0.001777f
C706 VDD.n17 GND 0.001777f
C707 VDD.n18 GND 0.001435f
C708 VDD.n19 GND 0.001435f
C709 VDD.n20 GND 0.001783f
C710 VDD.n21 GND 0.001783f
C711 VDD.n22 GND 0.158648f
C712 VDD.n23 GND 0.158648f
C713 VDD.n24 GND 0.001783f
C714 VDD.n25 GND 0.001783f
C715 VDD.n26 GND 0.001435f
C716 VDD.n27 GND 0.001783f
C717 VDD.n28 GND 0.001435f
C718 VDD.n29 GND 0.001783f
C719 VDD.n30 GND 0.158648f
C720 VDD.n31 GND 0.001783f
C721 VDD.n32 GND 0.001435f
C722 VDD.n33 GND 0.001783f
C723 VDD.n34 GND 0.001435f
C724 VDD.n35 GND 0.001783f
C725 VDD.n36 GND 0.158648f
C726 VDD.n37 GND 0.001783f
C727 VDD.n38 GND 0.001435f
C728 VDD.n39 GND 0.001783f
C729 VDD.n40 GND 0.001435f
C730 VDD.n41 GND 0.001783f
C731 VDD.n42 GND 0.158648f
C732 VDD.n43 GND 0.001783f
C733 VDD.n44 GND 0.001435f
C734 VDD.n45 GND 0.001783f
C735 VDD.n46 GND 0.001435f
C736 VDD.n47 GND 0.001783f
C737 VDD.n48 GND 0.107881f
C738 VDD.n49 GND 0.001783f
C739 VDD.n50 GND 0.001435f
C740 VDD.n51 GND 0.001783f
C741 VDD.n52 GND 0.001435f
C742 VDD.n53 GND 0.001783f
C743 VDD.n54 GND 0.158648f
C744 VDD.t7 GND 0.079324f
C745 VDD.n55 GND 0.001783f
C746 VDD.n56 GND 0.001435f
C747 VDD.n57 GND 0.003894f
C748 VDD.n58 GND 0.001191f
C749 VDD.n59 GND 0.003894f
C750 VDD.n60 GND 0.22766f
C751 VDD.n61 GND 0.003894f
C752 VDD.n62 GND 0.001191f
C753 VDD.n63 GND 0.001783f
C754 VDD.t68 GND 0.010031f
C755 VDD.t69 GND 0.014304f
C756 VDD.t67 GND 0.109243f
C757 VDD.n64 GND 0.024442f
C758 VDD.n65 GND 0.019628f
C759 VDD.n66 GND 0.002928f
C760 VDD.n67 GND 0.001783f
C761 VDD.t1 GND 2.33054f
C762 VDD.n100 GND 0.001783f
C763 VDD.n101 GND 0.001783f
C764 VDD.n102 GND 0.004059f
C765 VDD.n103 GND 0.001783f
C766 VDD.n104 GND 0.001783f
C767 VDD.n105 GND 0.001783f
C768 VDD.n106 GND 0.001783f
C769 VDD.n107 GND 0.001783f
C770 VDD.n108 GND 0.001783f
C771 VDD.n109 GND 0.001783f
C772 VDD.n110 GND 0.001783f
C773 VDD.n111 GND 0.001783f
C774 VDD.n112 GND 0.001783f
C775 VDD.n113 GND 0.001783f
C776 VDD.t18 GND 0.010031f
C777 VDD.t19 GND 0.014304f
C778 VDD.t17 GND 0.109243f
C779 VDD.n114 GND 0.024442f
C780 VDD.n115 GND 0.019628f
C781 VDD.n116 GND 0.001783f
C782 VDD.n117 GND 0.001783f
C783 VDD.n118 GND 0.001783f
C784 VDD.n119 GND 0.001783f
C785 VDD.n120 GND 0.001783f
C786 VDD.n121 GND 0.001052f
C787 VDD.n124 GND 0.001623f
C788 VDD.n125 GND 0.001783f
C789 VDD.n126 GND 0.001783f
C790 VDD.n127 GND 0.001198f
C791 VDD.n128 GND 0.001783f
C792 VDD.n129 GND 0.001783f
C793 VDD.n130 GND 0.001783f
C794 VDD.n131 GND 0.001783f
C795 VDD.n132 GND 0.001783f
C796 VDD.n133 GND 0.001783f
C797 VDD.n134 GND 0.001783f
C798 VDD.n135 GND 0.001783f
C799 VDD.n136 GND 0.001783f
C800 VDD.n137 GND 0.001783f
C801 VDD.n138 GND 0.001783f
C802 VDD.n139 GND 0.001428f
C803 VDD.t15 GND 0.010031f
C804 VDD.t16 GND 0.014304f
C805 VDD.t14 GND 0.109243f
C806 VDD.n140 GND 0.024442f
C807 VDD.n141 GND 0.019628f
C808 VDD.n142 GND 0.001783f
C809 VDD.n143 GND 0.001783f
C810 VDD.n144 GND 0.001783f
C811 VDD.n145 GND 0.001623f
C812 VDD.n148 GND 0.001212f
C813 VDD.n149 GND 0.001212f
C814 VDD.n150 GND 0.001212f
C815 VDD.t135 GND 2.1592f
C816 VDD.t111 GND 1.98627f
C817 VDD.t124 GND 1.98627f
C818 VDD.t130 GND 1.59124f
C819 VDD.n151 GND 0.70281f
C820 VDD.n152 GND 0.001212f
C821 VDD.n153 GND 0.001212f
C822 VDD.t72 GND 0.00872f
C823 VDD.t71 GND 0.013318f
C824 VDD.t70 GND 0.116692f
C825 VDD.n154 GND 0.016902f
C826 VDD.n155 GND 0.011832f
C827 VDD.n156 GND 0.001212f
C828 VDD.n158 GND 0.002794f
C829 VDD.n159 GND 0.001212f
C830 VDD.n160 GND 0.001212f
C831 VDD.n161 GND 0.107881f
C832 VDD.n162 GND 0.001212f
C833 VDD.n163 GND 0.158648f
C834 VDD.n164 GND 0.001212f
C835 VDD.n165 GND 0.001212f
C836 VDD.n166 GND 0.002794f
C837 VDD.n167 GND 0.001212f
C838 VDD.n168 GND 0.001212f
C839 VDD.n169 GND 0.001212f
C840 VDD.n170 GND 0.001212f
C841 VDD.n172 GND 0.001212f
C842 VDD.n173 GND 0.001212f
C843 VDD.n175 GND 0.001212f
C844 VDD.t46 GND 0.00872f
C845 VDD.t45 GND 0.013318f
C846 VDD.t43 GND 0.116692f
C847 VDD.n176 GND 0.016902f
C848 VDD.n177 GND 0.011832f
C849 VDD.n178 GND 0.001212f
C850 VDD.n180 GND 0.002794f
C851 VDD.n181 GND 0.001212f
C852 VDD.n182 GND 0.001212f
C853 VDD.n183 GND 0.107881f
C854 VDD.n184 GND 0.001212f
C855 VDD.n185 GND 0.001212f
C856 VDD.n186 GND 0.001212f
C857 VDD.n187 GND 0.001212f
C858 VDD.n188 GND 0.001212f
C859 VDD.n189 GND 0.107881f
C860 VDD.n190 GND 0.001212f
C861 VDD.n191 GND 0.001212f
C862 VDD.n192 GND 0.001212f
C863 VDD.n193 GND 0.001212f
C864 VDD.n194 GND 0.001212f
C865 VDD.n195 GND 0.001212f
C866 VDD.n196 GND 0.107881f
C867 VDD.n197 GND 0.001212f
C868 VDD.n198 GND 0.001212f
C869 VDD.n199 GND 0.001212f
C870 VDD.n200 GND 0.001212f
C871 VDD.n201 GND 0.001212f
C872 VDD.n202 GND 0.063459f
C873 VDD.n203 GND 0.001212f
C874 VDD.n204 GND 0.001212f
C875 VDD.n205 GND 0.001212f
C876 VDD.n206 GND 0.001212f
C877 VDD.n207 GND 0.001212f
C878 VDD.n208 GND 0.107881f
C879 VDD.n209 GND 0.001212f
C880 VDD.n210 GND 0.001212f
C881 VDD.t44 GND 0.05394f
C882 VDD.n211 GND 0.001212f
C883 VDD.n212 GND 0.001212f
C884 VDD.n213 GND 0.001212f
C885 VDD.n214 GND 0.094396f
C886 VDD.n215 GND 0.001212f
C887 VDD.n216 GND 0.001212f
C888 VDD.n217 GND 0.001212f
C889 VDD.n218 GND 0.001212f
C890 VDD.n219 GND 0.001212f
C891 VDD.n220 GND 0.107881f
C892 VDD.n221 GND 0.001212f
C893 VDD.n222 GND 0.001212f
C894 VDD.t117 GND 0.05394f
C895 VDD.n223 GND 0.001212f
C896 VDD.n224 GND 0.001212f
C897 VDD.n225 GND 0.001212f
C898 VDD.n226 GND 0.107881f
C899 VDD.n227 GND 0.001212f
C900 VDD.n228 GND 0.001212f
C901 VDD.n229 GND 0.001212f
C902 VDD.n230 GND 0.001212f
C903 VDD.n231 GND 0.001212f
C904 VDD.n232 GND 0.107881f
C905 VDD.n233 GND 0.001212f
C906 VDD.n234 GND 0.001212f
C907 VDD.n235 GND 0.001212f
C908 VDD.n236 GND 0.001212f
C909 VDD.n237 GND 0.001212f
C910 VDD.n238 GND 0.107881f
C911 VDD.n239 GND 0.001212f
C912 VDD.n240 GND 0.001212f
C913 VDD.n241 GND 0.001212f
C914 VDD.n242 GND 0.001212f
C915 VDD.n243 GND 0.001212f
C916 VDD.n244 GND 0.107881f
C917 VDD.n245 GND 0.001212f
C918 VDD.n246 GND 0.001212f
C919 VDD.n247 GND 0.001212f
C920 VDD.n248 GND 0.001212f
C921 VDD.n249 GND 0.001212f
C922 VDD.n250 GND 0.107881f
C923 VDD.n251 GND 0.001212f
C924 VDD.n252 GND 0.001212f
C925 VDD.n253 GND 0.001212f
C926 VDD.n254 GND 0.001212f
C927 VDD.n255 GND 0.001212f
C928 VDD.n256 GND 0.107881f
C929 VDD.n257 GND 0.001212f
C930 VDD.n258 GND 0.001212f
C931 VDD.n259 GND 0.001212f
C932 VDD.n260 GND 0.001212f
C933 VDD.n261 GND 0.001212f
C934 VDD.n262 GND 0.107881f
C935 VDD.n263 GND 0.001212f
C936 VDD.n264 GND 0.001212f
C937 VDD.n265 GND 0.001212f
C938 VDD.n266 GND 0.001212f
C939 VDD.n267 GND 0.001212f
C940 VDD.t119 GND 0.05394f
C941 VDD.n268 GND 0.001212f
C942 VDD.n269 GND 0.001212f
C943 VDD.n270 GND 0.001212f
C944 VDD.n271 GND 0.001212f
C945 VDD.n272 GND 0.001212f
C946 VDD.t105 GND 0.05394f
C947 VDD.n273 GND 0.001212f
C948 VDD.n274 GND 0.001212f
C949 VDD.n275 GND 0.065046f
C950 VDD.n276 GND 0.001212f
C951 VDD.n277 GND 0.001212f
C952 VDD.n278 GND 0.001212f
C953 VDD.n279 GND 0.107881f
C954 VDD.n280 GND 0.001212f
C955 VDD.n281 GND 0.001212f
C956 VDD.n282 GND 0.099155f
C957 VDD.n283 GND 0.001212f
C958 VDD.n284 GND 0.001212f
C959 VDD.n285 GND 0.001212f
C960 VDD.n286 GND 0.107881f
C961 VDD.n287 GND 0.001212f
C962 VDD.n288 GND 0.001212f
C963 VDD.n289 GND 0.001212f
C964 VDD.n290 GND 0.001212f
C965 VDD.n291 GND 0.001212f
C966 VDD.n292 GND 0.107881f
C967 VDD.n293 GND 0.001212f
C968 VDD.n294 GND 0.001212f
C969 VDD.n295 GND 0.001212f
C970 VDD.n296 GND 0.001212f
C971 VDD.n297 GND 0.001212f
C972 VDD.n298 GND 0.107881f
C973 VDD.n299 GND 0.001212f
C974 VDD.n300 GND 0.001212f
C975 VDD.n301 GND 0.001212f
C976 VDD.n302 GND 0.001212f
C977 VDD.n303 GND 0.001212f
C978 VDD.n304 GND 0.107881f
C979 VDD.n305 GND 0.001212f
C980 VDD.n306 GND 0.001212f
C981 VDD.n307 GND 0.001212f
C982 VDD.n308 GND 0.001212f
C983 VDD.n309 GND 0.001212f
C984 VDD.n310 GND 0.107881f
C985 VDD.n311 GND 0.001212f
C986 VDD.n312 GND 0.001212f
C987 VDD.n313 GND 0.001212f
C988 VDD.n314 GND 0.001212f
C989 VDD.n315 GND 0.001212f
C990 VDD.n316 GND 0.107881f
C991 VDD.n317 GND 0.001212f
C992 VDD.n318 GND 0.001212f
C993 VDD.n319 GND 0.001212f
C994 VDD.n320 GND 0.001212f
C995 VDD.n321 GND 0.001212f
C996 VDD.n322 GND 0.065046f
C997 VDD.n323 GND 0.001212f
C998 VDD.n324 GND 0.001212f
C999 VDD.n325 GND 0.001212f
C1000 VDD.n326 GND 0.001212f
C1001 VDD.n327 GND 0.001212f
C1002 VDD.t121 GND 0.05394f
C1003 VDD.n328 GND 0.001212f
C1004 VDD.n329 GND 0.001212f
C1005 VDD.t123 GND 0.05394f
C1006 VDD.n330 GND 0.001212f
C1007 VDD.n331 GND 0.001212f
C1008 VDD.n332 GND 0.001212f
C1009 VDD.n333 GND 0.107881f
C1010 VDD.n334 GND 0.001212f
C1011 VDD.n335 GND 0.001212f
C1012 VDD.n336 GND 0.076944f
C1013 VDD.n337 GND 0.001212f
C1014 VDD.n338 GND 0.001212f
C1015 VDD.n339 GND 0.001212f
C1016 VDD.n340 GND 0.107881f
C1017 VDD.n341 GND 0.001212f
C1018 VDD.n342 GND 0.001212f
C1019 VDD.n343 GND 0.001212f
C1020 VDD.n344 GND 0.001212f
C1021 VDD.n345 GND 0.001212f
C1022 VDD.n346 GND 0.107881f
C1023 VDD.n347 GND 0.001212f
C1024 VDD.n348 GND 0.001212f
C1025 VDD.n349 GND 0.001212f
C1026 VDD.n350 GND 0.001212f
C1027 VDD.n351 GND 0.001212f
C1028 VDD.n352 GND 0.107881f
C1029 VDD.n353 GND 0.001212f
C1030 VDD.n354 GND 0.001212f
C1031 VDD.n355 GND 0.001212f
C1032 VDD.n356 GND 0.001212f
C1033 VDD.n357 GND 0.001212f
C1034 VDD.n358 GND 0.107881f
C1035 VDD.n359 GND 0.001212f
C1036 VDD.n360 GND 0.001212f
C1037 VDD.n361 GND 0.001212f
C1038 VDD.n362 GND 0.001212f
C1039 VDD.n363 GND 0.001212f
C1040 VDD.n364 GND 0.107881f
C1041 VDD.n365 GND 0.001212f
C1042 VDD.n366 GND 0.001212f
C1043 VDD.n367 GND 0.001212f
C1044 VDD.n368 GND 0.001212f
C1045 VDD.n369 GND 0.001212f
C1046 VDD.n370 GND 0.107881f
C1047 VDD.n371 GND 0.001212f
C1048 VDD.n372 GND 0.001212f
C1049 VDD.n373 GND 0.001212f
C1050 VDD.n374 GND 0.001212f
C1051 VDD.n375 GND 0.001212f
C1052 VDD.n376 GND 0.107881f
C1053 VDD.n377 GND 0.001212f
C1054 VDD.n378 GND 0.001212f
C1055 VDD.n379 GND 0.001212f
C1056 VDD.n380 GND 0.001212f
C1057 VDD.n381 GND 0.001212f
C1058 VDD.t115 GND 0.05394f
C1059 VDD.n382 GND 0.001212f
C1060 VDD.n383 GND 0.001212f
C1061 VDD.n384 GND 0.001212f
C1062 VDD.n385 GND 0.001212f
C1063 VDD.n386 GND 0.001212f
C1064 VDD.t61 GND 0.05394f
C1065 VDD.n387 GND 0.001212f
C1066 VDD.n388 GND 0.001212f
C1067 VDD.n389 GND 0.054734f
C1068 VDD.n390 GND 0.001212f
C1069 VDD.n391 GND 0.001212f
C1070 VDD.n392 GND 0.001212f
C1071 VDD.n393 GND 0.107881f
C1072 VDD.n394 GND 0.001212f
C1073 VDD.n395 GND 0.001212f
C1074 VDD.n396 GND 0.063459f
C1075 VDD.n397 GND 0.001212f
C1076 VDD.n398 GND 0.001212f
C1077 VDD.n399 GND 0.001212f
C1078 VDD.n400 GND 0.107881f
C1079 VDD.n401 GND 0.001212f
C1080 VDD.n402 GND 0.001212f
C1081 VDD.n403 GND 0.001212f
C1082 VDD.n404 GND 0.001212f
C1083 VDD.n405 GND 0.001212f
C1084 VDD.n406 GND 0.107881f
C1085 VDD.n407 GND 0.001212f
C1086 VDD.n408 GND 0.001212f
C1087 VDD.n409 GND 0.001212f
C1088 VDD.n410 GND 0.001212f
C1089 VDD.n411 GND 0.001212f
C1090 VDD.n412 GND 0.107881f
C1091 VDD.n413 GND 0.001212f
C1092 VDD.n414 GND 0.001212f
C1093 VDD.n415 GND 0.001212f
C1094 VDD.n416 GND 0.002794f
C1095 VDD.n417 GND 0.002794f
C1096 VDD.n418 GND 0.158648f
C1097 VDD.n419 GND 0.001212f
C1098 VDD.n420 GND 0.001212f
C1099 VDD.n421 GND 0.002794f
C1100 VDD.n422 GND 0.001212f
C1101 VDD.n423 GND 0.001212f
C1102 VDD.n424 GND 0.158648f
C1103 VDD.n432 GND 0.002965f
C1104 VDD.n440 GND 0.002794f
C1105 VDD.n441 GND 0.001212f
C1106 VDD.n442 GND 0.002794f
C1107 VDD.t39 GND 0.00872f
C1108 VDD.t38 GND 0.013318f
C1109 VDD.t37 GND 0.116692f
C1110 VDD.n443 GND 0.016902f
C1111 VDD.n444 GND 0.011832f
C1112 VDD.n445 GND 0.002934f
C1113 VDD.n446 GND 0.001212f
C1114 VDD.n447 GND 0.001212f
C1115 VDD.n448 GND 0.107881f
C1116 VDD.n449 GND 0.001212f
C1117 VDD.n450 GND 0.001212f
C1118 VDD.n451 GND 0.001212f
C1119 VDD.n452 GND 0.001212f
C1120 VDD.n453 GND 0.001212f
C1121 VDD.n454 GND 0.107881f
C1122 VDD.n455 GND 0.001212f
C1123 VDD.n456 GND 0.001212f
C1124 VDD.n457 GND 0.001212f
C1125 VDD.n458 GND 0.001212f
C1126 VDD.n459 GND 0.001212f
C1127 VDD.t23 GND 0.00872f
C1128 VDD.t22 GND 0.013318f
C1129 VDD.t20 GND 0.116692f
C1130 VDD.n460 GND 0.016902f
C1131 VDD.n461 GND 0.011832f
C1132 VDD.n462 GND 0.001733f
C1133 VDD.n463 GND 0.001212f
C1134 VDD.n464 GND 0.001212f
C1135 VDD.n465 GND 0.107881f
C1136 VDD.n466 GND 0.001212f
C1137 VDD.n467 GND 0.001212f
C1138 VDD.n468 GND 0.001212f
C1139 VDD.n469 GND 0.001212f
C1140 VDD.n470 GND 0.001212f
C1141 VDD.n471 GND 0.107881f
C1142 VDD.n472 GND 0.001212f
C1143 VDD.n473 GND 0.001212f
C1144 VDD.n474 GND 0.001212f
C1145 VDD.n475 GND 0.001212f
C1146 VDD.n476 GND 0.001212f
C1147 VDD.n477 GND 0.001212f
C1148 VDD.n478 GND 0.063459f
C1149 VDD.n479 GND 0.001212f
C1150 VDD.n480 GND 0.001212f
C1151 VDD.n481 GND 0.001212f
C1152 VDD.n482 GND 0.001212f
C1153 VDD.n483 GND 0.001212f
C1154 VDD.n484 GND 0.054734f
C1155 VDD.n485 GND 0.001212f
C1156 VDD.n486 GND 0.001212f
C1157 VDD.t21 GND 0.05394f
C1158 VDD.n487 GND 0.001212f
C1159 VDD.n488 GND 0.001212f
C1160 VDD.n489 GND 0.001212f
C1161 VDD.n490 GND 0.107881f
C1162 VDD.n491 GND 0.001212f
C1163 VDD.n492 GND 0.001212f
C1164 VDD.t139 GND 0.05394f
C1165 VDD.n493 GND 0.001212f
C1166 VDD.n494 GND 0.001212f
C1167 VDD.n495 GND 0.001212f
C1168 VDD.n496 GND 0.107881f
C1169 VDD.n497 GND 0.001212f
C1170 VDD.n498 GND 0.001212f
C1171 VDD.n499 GND 0.001212f
C1172 VDD.n500 GND 0.001212f
C1173 VDD.n501 GND 0.001212f
C1174 VDD.n502 GND 0.107881f
C1175 VDD.n503 GND 0.001212f
C1176 VDD.n504 GND 0.001212f
C1177 VDD.n505 GND 0.001212f
C1178 VDD.n506 GND 0.001212f
C1179 VDD.n507 GND 0.001212f
C1180 VDD.n508 GND 0.107881f
C1181 VDD.n509 GND 0.001212f
C1182 VDD.n510 GND 0.001212f
C1183 VDD.n511 GND 0.001212f
C1184 VDD.n512 GND 0.001212f
C1185 VDD.n513 GND 0.001212f
C1186 VDD.n514 GND 0.107881f
C1187 VDD.n515 GND 0.001212f
C1188 VDD.n516 GND 0.001212f
C1189 VDD.n517 GND 0.001212f
C1190 VDD.n518 GND 0.001212f
C1191 VDD.n519 GND 0.001212f
C1192 VDD.n520 GND 0.107881f
C1193 VDD.n521 GND 0.001212f
C1194 VDD.n522 GND 0.001212f
C1195 VDD.n523 GND 0.001212f
C1196 VDD.n524 GND 0.001212f
C1197 VDD.n525 GND 0.001212f
C1198 VDD.n526 GND 0.107881f
C1199 VDD.n527 GND 0.001212f
C1200 VDD.n528 GND 0.001212f
C1201 VDD.n529 GND 0.001212f
C1202 VDD.n530 GND 0.001212f
C1203 VDD.n531 GND 0.001212f
C1204 VDD.n532 GND 0.107881f
C1205 VDD.n533 GND 0.001212f
C1206 VDD.n534 GND 0.001212f
C1207 VDD.n535 GND 0.001212f
C1208 VDD.n536 GND 0.001212f
C1209 VDD.n537 GND 0.001212f
C1210 VDD.n538 GND 0.076944f
C1211 VDD.n539 GND 0.001212f
C1212 VDD.n540 GND 0.001212f
C1213 VDD.n541 GND 0.001212f
C1214 VDD.n542 GND 0.001212f
C1215 VDD.n543 GND 0.001212f
C1216 VDD.t120 GND 0.05394f
C1217 VDD.n544 GND 0.001212f
C1218 VDD.n545 GND 0.001212f
C1219 VDD.t113 GND 0.05394f
C1220 VDD.n546 GND 0.001212f
C1221 VDD.n547 GND 0.001212f
C1222 VDD.n548 GND 0.001212f
C1223 VDD.n549 GND 0.107881f
C1224 VDD.n550 GND 0.001212f
C1225 VDD.n551 GND 0.001212f
C1226 VDD.n552 GND 0.065046f
C1227 VDD.n553 GND 0.001212f
C1228 VDD.n554 GND 0.001212f
C1229 VDD.n555 GND 0.001212f
C1230 VDD.n556 GND 0.107881f
C1231 VDD.n557 GND 0.001212f
C1232 VDD.n558 GND 0.001212f
C1233 VDD.n559 GND 0.001212f
C1234 VDD.n560 GND 0.001212f
C1235 VDD.n561 GND 0.001212f
C1236 VDD.n562 GND 0.107881f
C1237 VDD.n563 GND 0.001212f
C1238 VDD.n564 GND 0.001212f
C1239 VDD.n565 GND 0.001212f
C1240 VDD.n566 GND 0.001212f
C1241 VDD.n567 GND 0.001212f
C1242 VDD.n568 GND 0.107881f
C1243 VDD.n569 GND 0.001212f
C1244 VDD.n570 GND 0.001212f
C1245 VDD.n571 GND 0.001212f
C1246 VDD.n572 GND 0.001212f
C1247 VDD.n573 GND 0.001212f
C1248 VDD.n574 GND 0.107881f
C1249 VDD.n575 GND 0.001212f
C1250 VDD.n576 GND 0.001212f
C1251 VDD.n577 GND 0.001212f
C1252 VDD.n578 GND 0.001212f
C1253 VDD.n579 GND 0.001212f
C1254 VDD.n580 GND 0.107881f
C1255 VDD.n581 GND 0.001212f
C1256 VDD.n582 GND 0.001212f
C1257 VDD.n583 GND 0.001212f
C1258 VDD.n584 GND 0.001212f
C1259 VDD.n585 GND 0.001212f
C1260 VDD.n586 GND 0.107881f
C1261 VDD.n587 GND 0.001212f
C1262 VDD.n588 GND 0.001212f
C1263 VDD.n589 GND 0.001212f
C1264 VDD.n590 GND 0.001212f
C1265 VDD.n591 GND 0.001212f
C1266 VDD.n592 GND 0.099155f
C1267 VDD.n593 GND 0.001212f
C1268 VDD.n594 GND 0.001212f
C1269 VDD.n595 GND 0.001212f
C1270 VDD.n596 GND 0.001212f
C1271 VDD.n597 GND 0.001212f
C1272 VDD.n598 GND 0.065046f
C1273 VDD.n599 GND 0.001212f
C1274 VDD.n600 GND 0.001212f
C1275 VDD.t96 GND 0.05394f
C1276 VDD.n601 GND 0.001212f
C1277 VDD.n602 GND 0.001212f
C1278 VDD.n603 GND 0.001212f
C1279 VDD.n604 GND 0.107881f
C1280 VDD.n605 GND 0.001212f
C1281 VDD.n606 GND 0.001212f
C1282 VDD.t102 GND 0.05394f
C1283 VDD.n607 GND 0.001212f
C1284 VDD.n608 GND 0.001212f
C1285 VDD.n609 GND 0.001212f
C1286 VDD.n610 GND 0.107881f
C1287 VDD.n611 GND 0.001212f
C1288 VDD.n612 GND 0.001212f
C1289 VDD.n613 GND 0.001212f
C1290 VDD.n614 GND 0.001212f
C1291 VDD.n615 GND 0.001212f
C1292 VDD.n616 GND 0.107881f
C1293 VDD.n617 GND 0.001212f
C1294 VDD.n618 GND 0.001212f
C1295 VDD.n619 GND 0.001212f
C1296 VDD.n620 GND 0.001212f
C1297 VDD.n621 GND 0.001212f
C1298 VDD.n622 GND 0.107881f
C1299 VDD.n623 GND 0.001212f
C1300 VDD.n624 GND 0.001212f
C1301 VDD.n625 GND 0.001212f
C1302 VDD.n626 GND 0.001212f
C1303 VDD.n627 GND 0.001212f
C1304 VDD.n628 GND 0.107881f
C1305 VDD.n629 GND 0.001212f
C1306 VDD.n630 GND 0.001212f
C1307 VDD.n631 GND 0.001212f
C1308 VDD.n632 GND 0.001212f
C1309 VDD.n633 GND 0.001212f
C1310 VDD.n634 GND 0.107881f
C1311 VDD.n635 GND 0.001212f
C1312 VDD.n636 GND 0.001212f
C1313 VDD.n637 GND 0.001212f
C1314 VDD.n638 GND 0.001212f
C1315 VDD.n639 GND 0.001212f
C1316 VDD.n640 GND 0.107881f
C1317 VDD.n641 GND 0.001212f
C1318 VDD.n642 GND 0.001212f
C1319 VDD.n643 GND 0.001212f
C1320 VDD.n644 GND 0.001212f
C1321 VDD.n645 GND 0.001212f
C1322 VDD.n646 GND 0.107881f
C1323 VDD.n647 GND 0.001212f
C1324 VDD.n648 GND 0.001212f
C1325 VDD.n649 GND 0.001212f
C1326 VDD.n650 GND 0.001212f
C1327 VDD.n651 GND 0.001212f
C1328 VDD.t100 GND 0.05394f
C1329 VDD.n652 GND 0.001212f
C1330 VDD.n653 GND 0.001212f
C1331 VDD.n654 GND 0.001212f
C1332 VDD.n655 GND 0.001212f
C1333 VDD.n656 GND 0.001212f
C1334 VDD.n657 GND 0.107881f
C1335 VDD.n658 GND 0.001212f
C1336 VDD.n659 GND 0.001212f
C1337 VDD.n660 GND 0.094396f
C1338 VDD.n661 GND 0.001212f
C1339 VDD.n662 GND 0.001212f
C1340 VDD.n663 GND 0.001212f
C1341 VDD.t11 GND 0.05394f
C1342 VDD.n664 GND 0.001212f
C1343 VDD.n665 GND 0.001212f
C1344 VDD.n666 GND 0.001212f
C1345 VDD.n667 GND 0.001212f
C1346 VDD.n668 GND 0.001212f
C1347 VDD.n669 GND 0.107881f
C1348 VDD.n670 GND 0.001212f
C1349 VDD.n671 GND 0.001212f
C1350 VDD.n672 GND 0.063459f
C1351 VDD.n673 GND 0.001212f
C1352 VDD.n674 GND 0.001212f
C1353 VDD.n675 GND 0.001212f
C1354 VDD.n676 GND 0.107881f
C1355 VDD.n677 GND 0.001212f
C1356 VDD.n678 GND 0.001212f
C1357 VDD.n679 GND 0.001212f
C1358 VDD.n680 GND 0.001212f
C1359 VDD.n681 GND 0.001212f
C1360 VDD.n682 GND 0.107881f
C1361 VDD.n683 GND 0.001212f
C1362 VDD.n684 GND 0.001212f
C1363 VDD.n685 GND 0.001212f
C1364 VDD.n686 GND 0.001212f
C1365 VDD.n687 GND 0.001212f
C1366 VDD.n688 GND 0.107881f
C1367 VDD.n689 GND 0.001212f
C1368 VDD.n690 GND 0.001212f
C1369 VDD.n691 GND 0.001212f
C1370 VDD.n692 GND 0.002794f
C1371 VDD.n693 GND 0.002794f
C1372 VDD.n694 GND 0.158648f
C1373 VDD.n695 GND 0.001212f
C1374 VDD.n696 GND 0.001212f
C1375 VDD.n697 GND 0.002794f
C1376 VDD.n698 GND 0.001212f
C1377 VDD.n699 GND 0.001212f
C1378 VDD.t128 GND 1.59124f
C1379 VDD.n713 GND 0.002965f
C1380 VDD.n714 GND 0.001212f
C1381 VDD.n715 GND 0.001052f
C1382 VDD.n716 GND 0.001623f
C1383 VDD.n718 GND 0.001435f
C1384 VDD.n719 GND 0.001435f
C1385 VDD.n720 GND 0.001783f
C1386 VDD.t107 GND 1.98627f
C1387 VDD.t109 GND 1.98627f
C1388 VDD.t94 GND 2.1592f
C1389 VDD.t0 GND 2.33054f
C1390 VDD.n721 GND 1.31281f
C1391 VDD.n722 GND 0.001435f
C1392 VDD.n723 GND 0.001783f
C1393 VDD.n724 GND 0.001783f
C1394 VDD.n725 GND 0.001198f
C1395 VDD.n727 GND 0.001783f
C1396 VDD.n728 GND 0.001198f
C1397 VDD.t75 GND 0.010031f
C1398 VDD.t74 GND 0.014304f
C1399 VDD.t73 GND 0.109243f
C1400 VDD.n729 GND 0.024442f
C1401 VDD.n730 GND 0.019628f
C1402 VDD.n731 GND 0.001783f
C1403 VDD.n732 GND 0.001783f
C1404 VDD.n733 GND 0.001435f
C1405 VDD.n735 GND 0.001783f
C1406 VDD.n736 GND 0.001783f
C1407 VDD.n737 GND 0.001783f
C1408 VDD.n738 GND 0.001783f
C1409 VDD.n739 GND 0.001435f
C1410 VDD.n741 GND 0.001783f
C1411 VDD.n742 GND 0.001783f
C1412 VDD.n743 GND 0.001783f
C1413 VDD.n744 GND 0.001783f
C1414 VDD.n745 GND 0.001783f
C1415 VDD.n746 GND 0.001435f
C1416 VDD.n748 GND 0.001783f
C1417 VDD.n749 GND 0.001783f
C1418 VDD.n750 GND 0.001783f
C1419 VDD.n751 GND 0.001783f
C1420 VDD.n752 GND 0.001428f
C1421 VDD.t81 GND 0.010031f
C1422 VDD.t80 GND 0.014304f
C1423 VDD.t79 GND 0.109243f
C1424 VDD.n753 GND 0.024442f
C1425 VDD.n754 GND 0.019628f
C1426 VDD.n756 GND 0.001783f
C1427 VDD.n757 GND 0.001783f
C1428 VDD.n758 GND 0.001435f
C1429 VDD.n759 GND 0.001783f
C1430 VDD.n761 GND 0.001783f
C1431 VDD.n762 GND 0.001783f
C1432 VDD.n763 GND 0.001783f
C1433 VDD.n764 GND 0.001623f
C1434 VDD.n765 GND 0.001435f
C1435 VDD.n767 GND 0.001783f
C1436 VDD.n768 GND 0.001435f
C1437 VDD.n769 GND 0.002965f
C1438 VDD.n770 GND 0.002965f
C1439 VDD.n771 GND 0.001212f
C1440 VDD.n772 GND 0.001212f
C1441 VDD.n773 GND 0.001212f
C1442 VDD.n774 GND 0.001212f
C1443 VDD.n775 GND 0.001212f
C1444 VDD.n776 GND 0.001212f
C1445 VDD.n777 GND 0.001212f
C1446 VDD.n778 GND 0.001212f
C1447 VDD.n779 GND 0.001212f
C1448 VDD.n780 GND 0.001212f
C1449 VDD.n781 GND 0.001212f
C1450 VDD.n782 GND 0.001212f
C1451 VDD.n783 GND 0.001212f
C1452 VDD.t65 GND 0.00872f
C1453 VDD.t66 GND 0.013318f
C1454 VDD.t64 GND 0.116692f
C1455 VDD.n784 GND 0.016902f
C1456 VDD.n785 GND 0.011832f
C1457 VDD.n786 GND 0.001733f
C1458 VDD.n787 GND 0.001212f
C1459 VDD.n788 GND 0.001212f
C1460 VDD.n789 GND 0.001212f
C1461 VDD.n790 GND 0.001212f
C1462 VDD.n791 GND 0.001212f
C1463 VDD.n792 GND 0.001212f
C1464 VDD.n793 GND 0.001212f
C1465 VDD.n794 GND 0.001212f
C1466 VDD.n795 GND 0.001212f
C1467 VDD.n796 GND 0.001212f
C1468 VDD.n797 GND 0.001212f
C1469 VDD.n798 GND 0.001212f
C1470 VDD.n799 GND 0.001212f
C1471 VDD.n800 GND 0.001212f
C1472 VDD.n801 GND 0.001212f
C1473 VDD.n802 GND 0.001212f
C1474 VDD.n803 GND 0.001212f
C1475 VDD.n804 GND 0.001212f
C1476 VDD.n805 GND 0.001212f
C1477 VDD.n806 GND 0.001212f
C1478 VDD.n807 GND 0.001212f
C1479 VDD.n808 GND 0.001212f
C1480 VDD.n809 GND 0.001212f
C1481 VDD.n810 GND 0.001212f
C1482 VDD.n811 GND 0.001212f
C1483 VDD.n812 GND 0.001212f
C1484 VDD.n813 GND 0.001212f
C1485 VDD.n814 GND 0.001212f
C1486 VDD.n815 GND 0.001212f
C1487 VDD.n816 GND 0.001212f
C1488 VDD.n817 GND 0.001212f
C1489 VDD.n818 GND 0.001212f
C1490 VDD.n819 GND 0.001212f
C1491 VDD.n820 GND 0.001212f
C1492 VDD.n821 GND 0.001212f
C1493 VDD.n822 GND 0.001212f
C1494 VDD.n823 GND 0.001212f
C1495 VDD.n824 GND 0.001212f
C1496 VDD.n825 GND 0.001212f
C1497 VDD.n826 GND 0.001212f
C1498 VDD.n827 GND 0.001212f
C1499 VDD.n828 GND 0.001212f
C1500 VDD.n829 GND 0.001212f
C1501 VDD.n830 GND 0.001212f
C1502 VDD.n831 GND 0.001212f
C1503 VDD.n832 GND 0.001212f
C1504 VDD.n833 GND 0.001212f
C1505 VDD.n834 GND 0.001212f
C1506 VDD.n835 GND 0.001212f
C1507 VDD.n836 GND 0.001212f
C1508 VDD.n837 GND 0.001212f
C1509 VDD.n838 GND 0.001212f
C1510 VDD.n839 GND 0.001212f
C1511 VDD.n840 GND 0.001212f
C1512 VDD.n841 GND 0.001212f
C1513 VDD.n842 GND 0.001212f
C1514 VDD.n843 GND 0.001212f
C1515 VDD.n844 GND 0.001212f
C1516 VDD.n845 GND 0.001212f
C1517 VDD.n846 GND 0.001212f
C1518 VDD.n847 GND 0.001212f
C1519 VDD.n848 GND 0.001212f
C1520 VDD.n849 GND 0.001212f
C1521 VDD.n850 GND 0.001212f
C1522 VDD.n851 GND 0.001212f
C1523 VDD.n852 GND 0.001212f
C1524 VDD.n853 GND 0.001212f
C1525 VDD.n854 GND 0.001212f
C1526 VDD.n855 GND 0.001212f
C1527 VDD.n856 GND 0.001212f
C1528 VDD.n857 GND 0.001212f
C1529 VDD.n858 GND 0.001212f
C1530 VDD.n859 GND 0.001212f
C1531 VDD.n860 GND 0.001212f
C1532 VDD.n861 GND 0.001212f
C1533 VDD.n862 GND 0.001212f
C1534 VDD.n863 GND 0.001212f
C1535 VDD.n864 GND 0.001212f
C1536 VDD.n865 GND 0.001212f
C1537 VDD.n866 GND 0.001212f
C1538 VDD.n867 GND 0.001212f
C1539 VDD.n868 GND 0.001212f
C1540 VDD.n869 GND 0.001212f
C1541 VDD.n870 GND 0.001212f
C1542 VDD.n871 GND 0.001212f
C1543 VDD.n872 GND 0.001212f
C1544 VDD.n873 GND 0.001212f
C1545 VDD.n874 GND 0.001212f
C1546 VDD.n875 GND 0.001212f
C1547 VDD.n876 GND 0.001212f
C1548 VDD.n877 GND 0.001212f
C1549 VDD.n878 GND 0.001212f
C1550 VDD.n879 GND 0.001212f
C1551 VDD.n880 GND 0.001212f
C1552 VDD.n881 GND 0.001212f
C1553 VDD.n882 GND 0.001212f
C1554 VDD.n883 GND 0.001212f
C1555 VDD.n884 GND 0.001212f
C1556 VDD.n885 GND 0.001212f
C1557 VDD.n886 GND 0.001212f
C1558 VDD.n887 GND 0.001212f
C1559 VDD.n888 GND 0.001212f
C1560 VDD.n889 GND 0.001212f
C1561 VDD.n890 GND 0.001212f
C1562 VDD.n891 GND 0.001212f
C1563 VDD.n892 GND 0.001212f
C1564 VDD.n893 GND 0.001212f
C1565 VDD.n894 GND 0.001212f
C1566 VDD.n895 GND 0.001212f
C1567 VDD.n896 GND 0.001212f
C1568 VDD.n897 GND 0.001212f
C1569 VDD.n898 GND 0.001212f
C1570 VDD.n899 GND 0.001212f
C1571 VDD.n900 GND 0.002794f
C1572 VDD.n901 GND 0.002794f
C1573 VDD.n902 GND 0.002965f
C1574 VDD.n903 GND 0.001212f
C1575 VDD.n904 GND 0.001212f
C1576 VDD.n905 GND 8.74e-19
C1577 VDD.n906 GND 0.001212f
C1578 VDD.n907 GND 0.001212f
C1579 VDD.n908 GND 9.45e-19
C1580 VDD.n909 GND 0.001212f
C1581 VDD.n910 GND 0.001212f
C1582 VDD.n911 GND 0.001212f
C1583 VDD.n912 GND 0.001212f
C1584 VDD.n913 GND 0.001212f
C1585 VDD.n914 GND 0.001212f
C1586 VDD.n915 GND 0.065701f
C1587 VDD.n917 GND 0.001783f
C1588 VDD.n918 GND 0.001435f
C1589 VDD.n920 GND 0.001783f
C1590 VDD.n921 GND 0.001783f
C1591 VDD.n923 GND 0.001783f
C1592 VDD.n924 GND 0.001783f
C1593 VDD.t50 GND 0.010031f
C1594 VDD.t49 GND 0.014304f
C1595 VDD.t47 GND 0.109243f
C1596 VDD.n925 GND 0.024442f
C1597 VDD.n926 GND 0.019628f
C1598 VDD.n927 GND 0.00221f
C1599 VDD.n928 GND 0.001783f
C1600 VDD.n930 GND 0.001783f
C1601 VDD.n931 GND 0.001783f
C1602 VDD.n933 GND 0.001783f
C1603 VDD.n934 GND 0.001435f
C1604 VDD.n935 GND 0.001783f
C1605 VDD.n936 GND 0.001783f
C1606 VDD.n938 GND 0.001783f
C1607 VDD.n939 GND 0.001783f
C1608 VDD.n941 GND 0.001783f
C1609 VDD.n942 GND 0.001435f
C1610 VDD.n943 GND 0.001783f
C1611 VDD.n944 GND 0.001783f
C1612 VDD.n946 GND 0.001783f
C1613 VDD.n947 GND 0.001783f
C1614 VDD.n949 GND 0.001783f
C1615 VDD.n950 GND 0.001435f
C1616 VDD.n951 GND 0.001783f
C1617 VDD.n952 GND 0.001783f
C1618 VDD.n954 GND 0.001783f
C1619 VDD.n955 GND 9.26e-19
C1620 VDD.t78 GND 0.010031f
C1621 VDD.t77 GND 0.014304f
C1622 VDD.t76 GND 0.109243f
C1623 VDD.n956 GND 0.024442f
C1624 VDD.n957 GND 0.019628f
C1625 VDD.n958 GND 0.001783f
C1626 VDD.n959 GND 0.001191f
C1627 VDD.n960 GND 0.158648f
C1628 VDD.n961 GND 0.001783f
C1629 VDD.n962 GND 0.004059f
C1630 VDD.n963 GND 0.001435f
C1631 VDD.n964 GND 0.001783f
C1632 VDD.n965 GND 0.001435f
C1633 VDD.n966 GND 0.001783f
C1634 VDD.n967 GND 0.130091f
C1635 VDD.n968 GND 0.001783f
C1636 VDD.n969 GND 0.001435f
C1637 VDD.n970 GND 0.001435f
C1638 VDD.n971 GND 0.001783f
C1639 VDD.n972 GND 0.001435f
C1640 VDD.n973 GND 0.001783f
C1641 VDD.n974 GND 0.158648f
C1642 VDD.t48 GND 0.079324f
C1643 VDD.n975 GND 0.001783f
C1644 VDD.n976 GND 0.001435f
C1645 VDD.n977 GND 0.001783f
C1646 VDD.n978 GND 0.001435f
C1647 VDD.n979 GND 0.001783f
C1648 VDD.n980 GND 0.158648f
C1649 VDD.n981 GND 0.001783f
C1650 VDD.n982 GND 0.001435f
C1651 VDD.n983 GND 0.001783f
C1652 VDD.n984 GND 0.001435f
C1653 VDD.n985 GND 0.001783f
C1654 VDD.n986 GND 0.158648f
C1655 VDD.n987 GND 0.001783f
C1656 VDD.n988 GND 0.001435f
C1657 VDD.n989 GND 0.001783f
C1658 VDD.n990 GND 0.001435f
C1659 VDD.n991 GND 0.001783f
C1660 VDD.n992 GND 0.158648f
C1661 VDD.n993 GND 0.001783f
C1662 VDD.n994 GND 0.001435f
C1663 VDD.n995 GND 0.001783f
C1664 VDD.n996 GND 0.001435f
C1665 VDD.n997 GND 0.001783f
C1666 VDD.t98 GND 0.158648f
C1667 VDD.n998 GND 0.001783f
C1668 VDD.n999 GND 0.001435f
C1669 VDD.n1000 GND 0.001783f
C1670 VDD.n1001 GND 0.001435f
C1671 VDD.n1002 GND 0.001783f
C1672 VDD.n1003 GND 0.158648f
C1673 VDD.n1004 GND 0.001783f
C1674 VDD.n1005 GND 0.001435f
C1675 VDD.n1006 GND 0.001783f
C1676 VDD.n1007 GND 0.001435f
C1677 VDD.n1008 GND 0.001783f
C1678 VDD.n1009 GND 0.158648f
C1679 VDD.n1010 GND 0.001783f
C1680 VDD.n1011 GND 0.001435f
C1681 VDD.n1012 GND 0.001783f
C1682 VDD.n1013 GND 0.001435f
C1683 VDD.n1014 GND 0.001783f
C1684 VDD.n1015 GND 0.158648f
C1685 VDD.n1016 GND 0.001783f
C1686 VDD.n1017 GND 0.001435f
C1687 VDD.n1018 GND 0.001783f
C1688 VDD.n1019 GND 0.001435f
C1689 VDD.n1020 GND 0.001783f
C1690 VDD.n1021 GND 0.158648f
C1691 VDD.n1022 GND 0.001783f
C1692 VDD.n1023 GND 0.001435f
C1693 VDD.n1024 GND 0.001783f
C1694 VDD.n1025 GND 0.001435f
C1695 VDD.n1026 GND 0.001783f
C1696 VDD.t3 GND 0.079324f
C1697 VDD.n1027 GND 0.001783f
C1698 VDD.n1028 GND 0.001435f
C1699 VDD.n1029 GND 0.001783f
C1700 VDD.n1030 GND 0.001435f
C1701 VDD.n1031 GND 0.001783f
C1702 VDD.n1032 GND 0.158648f
C1703 VDD.n1033 GND 0.130091f
C1704 VDD.n1034 GND 0.001783f
C1705 VDD.n1035 GND 0.001435f
C1706 VDD.n1036 GND 0.004059f
C1707 VDD.n1037 GND 0.004059f
C1708 VDD.n1038 GND 0.372029f
C1709 VDD.n1039 GND 0.004059f
C1710 VDD.n1040 GND 0.001783f
C1711 VDD.n1041 GND 0.001783f
C1712 VDD.t25 GND 0.010031f
C1713 VDD.t26 GND 0.014304f
C1714 VDD.t24 GND 0.109243f
C1715 VDD.n1042 GND 0.024442f
C1716 VDD.n1043 GND 0.019628f
C1717 VDD.n1044 GND 0.001435f
C1718 VDD.n1046 GND 0.001783f
C1719 VDD.n1047 GND 0.001783f
C1720 VDD.n1048 GND 0.001435f
C1721 VDD.n1049 GND 0.001783f
C1722 VDD.n1050 GND 0.001435f
C1723 VDD.n1051 GND 0.001783f
C1724 VDD.n1052 GND 0.001435f
C1725 VDD.n1053 GND 0.001783f
C1726 VDD.n1054 GND 0.001435f
C1727 VDD.n1055 GND 0.001783f
C1728 VDD.n1056 GND 0.001435f
C1729 VDD.n1057 GND 0.001783f
C1730 VDD.t4 GND 0.010031f
C1731 VDD.t5 GND 0.014304f
C1732 VDD.t2 GND 0.109243f
C1733 VDD.n1058 GND 0.024442f
C1734 VDD.n1059 GND 0.019628f
C1735 VDD.n1060 GND 0.00221f
C1736 VDD.n1061 GND 0.001783f
C1737 VDD.n1062 GND 0.001435f
C1738 VDD.n1063 GND 0.001783f
C1739 VDD.n1064 GND 0.001435f
C1740 VDD.n1065 GND 0.001783f
C1741 VDD.n1066 GND 0.001435f
C1742 VDD.n1067 GND 0.001783f
C1743 VDD.n1068 GND 0.001435f
C1744 VDD.n1069 GND 0.001783f
C1745 VDD.n1070 GND 0.001435f
C1746 VDD.n1071 GND 0.001783f
C1747 VDD.n1072 GND 0.001428f
C1748 VDD.n1073 GND 0.001783f
C1749 VDD.n1075 GND 0.001783f
C1750 VDD.t55 GND 0.010031f
C1751 VDD.t56 GND 0.014304f
C1752 VDD.t54 GND 0.109243f
C1753 VDD.n1076 GND 0.024442f
C1754 VDD.n1077 GND 0.019628f
C1755 VDD.n1078 GND 0.001435f
C1756 VDD.n1079 GND 0.001435f
C1757 VDD.n1080 GND 0.001783f
C1758 VDD.n1081 GND 0.001435f
C1759 VDD.n1082 GND 0.001783f
C1760 VDD.n1083 GND 0.001435f
C1761 VDD.n1084 GND 0.001783f
C1762 VDD.n1085 GND 0.001435f
C1763 VDD.n1086 GND 0.001783f
C1764 VDD.n1087 GND 0.001435f
C1765 VDD.n1088 GND 0.001783f
C1766 VDD.n1089 GND 0.001198f
C1767 VDD.n1090 GND 0.001783f
C1768 VDD.n1092 GND 0.001783f
C1769 VDD.t52 GND 0.010031f
C1770 VDD.t53 GND 0.014304f
C1771 VDD.t51 GND 0.109243f
C1772 VDD.n1093 GND 0.024442f
C1773 VDD.n1094 GND 0.019628f
C1774 VDD.n1095 GND 0.001435f
C1775 VDD.n1096 GND 0.001435f
C1776 VDD.n1097 GND 0.001783f
C1777 VDD.n1098 GND 0.001435f
C1778 VDD.n1099 GND 0.001783f
C1779 VDD.n1100 GND 0.001435f
C1780 VDD.n1101 GND 0.001783f
C1781 VDD.n1102 GND 0.001435f
C1782 VDD.n1103 GND 0.001783f
C1783 VDD.n1104 GND 0.001435f
C1784 VDD.n1105 GND 0.001783f
C1785 VDD.n1106 GND 9.69e-19
C1786 VDD.n1107 GND 0.001783f
C1787 VDD.n1109 GND 0.001783f
C1788 VDD.t58 GND 0.010031f
C1789 VDD.t59 GND 0.014304f
C1790 VDD.t57 GND 0.109243f
C1791 VDD.n1110 GND 0.024442f
C1792 VDD.n1111 GND 0.019628f
C1793 VDD.n1112 GND 0.001435f
C1794 VDD.n1113 GND 0.001435f
C1795 VDD.n1114 GND 0.001783f
C1796 VDD.n1115 GND 0.001435f
C1797 VDD.n1116 GND 0.001783f
C1798 VDD.n1117 GND 0.001435f
C1799 VDD.n1118 GND 0.001783f
C1800 VDD.n1119 GND 0.001435f
C1801 VDD.n1120 GND 0.001191f
C1802 VDD.n1122 GND 0.001783f
C1803 VDD.n1123 GND 0.001435f
C1804 VDD.n1124 GND 0.001783f
C1805 VDD.n1125 GND 0.001783f
C1806 VDD.n1126 GND 0.001783f
C1807 VDD.n1127 GND 0.001435f
C1808 VDD.n1128 GND 0.001783f
C1809 VDD.n1130 GND 0.001783f
C1810 VDD.n1132 GND 0.001783f
C1811 VDD.n1133 GND 0.001435f
C1812 VDD.n1134 GND 0.001783f
C1813 VDD.n1135 GND 0.001783f
C1814 VDD.n1136 GND 0.001783f
C1815 VDD.n1137 GND 0.001783f
C1816 VDD.n1138 GND 0.001783f
C1817 VDD.n1139 GND 0.001435f
C1818 VDD.n1140 GND 0.001783f
C1819 VDD.n1142 GND 0.001783f
C1820 VDD.n1143 GND 0.001783f
C1821 VDD.n1145 GND 0.001783f
C1822 VDD.n1146 GND 0.001428f
C1823 VDD.n1147 GND 0.002928f
C1824 VDD.n1148 GND 0.001783f
C1825 VDD.n1149 GND 0.001783f
C1826 VDD.n1150 GND 0.001783f
C1827 VDD.n1151 GND 0.001435f
C1828 VDD.n1152 GND 0.001783f
C1829 VDD.n1154 GND 0.001783f
C1830 VDD.n1156 GND 0.001783f
C1831 VDD.n1157 GND 0.001435f
C1832 VDD.n1158 GND 0.001783f
C1833 VDD.n1159 GND 0.001783f
C1834 VDD.n1160 GND 0.001783f
C1835 VDD.n1161 GND 0.001435f
C1836 VDD.n1162 GND 0.001783f
C1837 VDD.n1164 GND 0.001783f
C1838 VDD.n1166 GND 0.001783f
C1839 VDD.n1167 GND 0.001435f
C1840 VDD.n1168 GND 0.001783f
C1841 VDD.n1169 GND 0.001783f
C1842 VDD.n1170 GND 0.001783f
C1843 VDD.n1171 GND 0.001783f
C1844 VDD.n1172 GND 0.001783f
C1845 VDD.n1173 GND 0.001435f
C1846 VDD.n1174 GND 0.001783f
C1847 VDD.n1176 GND 0.001783f
C1848 VDD.n1177 GND 0.001783f
C1849 VDD.n1179 GND 0.001783f
C1850 VDD.n1180 GND 0.001198f
C1851 VDD.n1181 GND 0.002928f
C1852 VDD.n1182 GND 0.001783f
C1853 VDD.n1183 GND 0.001783f
C1854 VDD.n1184 GND 0.001783f
C1855 VDD.n1185 GND 0.001435f
C1856 VDD.n1186 GND 0.001783f
C1857 VDD.n1188 GND 0.001783f
C1858 VDD.n1190 GND 0.001783f
C1859 VDD.n1191 GND 0.001435f
C1860 VDD.n1192 GND 0.001783f
C1861 VDD.n1193 GND 0.001783f
C1862 VDD.n1194 GND 0.001783f
C1863 VDD.n1195 GND 0.001435f
C1864 VDD.n1196 GND 0.001783f
C1865 VDD.n1198 GND 0.001783f
C1866 VDD.n1200 GND 0.001783f
C1867 VDD.n1201 GND 0.001435f
C1868 VDD.n1202 GND 0.001783f
C1869 VDD.n1203 GND 0.001783f
C1870 VDD.n1204 GND 0.001783f
C1871 VDD.n1205 GND 0.001783f
C1872 VDD.n1206 GND 0.001783f
C1873 VDD.n1207 GND 0.001435f
C1874 VDD.n1208 GND 0.001783f
C1875 VDD.n1210 GND 0.001783f
C1876 VDD.n1211 GND 0.001783f
C1877 VDD.n1213 GND 0.001783f
C1878 VDD.n1214 GND 9.69e-19
C1879 VDD.n1215 GND 0.002928f
C1880 VDD.n1216 GND 0.001783f
C1881 VDD.n1217 GND 0.001783f
C1882 VDD.n1218 GND 0.001783f
C1883 VDD.n1219 GND 0.001435f
C1884 VDD.n1220 GND 0.001783f
C1885 VDD.n1222 GND 0.001783f
C1886 VDD.n1224 GND 0.001783f
C1887 VDD.n1225 GND 0.001435f
C1888 VDD.n1226 GND 0.001783f
C1889 VDD.n1227 GND 0.001783f
C1890 VDD.n1228 GND 0.001783f
C1891 VDD.n1229 GND 0.001435f
C1892 VDD.n1230 GND 0.001783f
C1893 VDD.n1232 GND 0.001783f
C1894 VDD.n1234 GND 0.001783f
C1895 VDD.n1235 GND 0.001435f
C1896 VDD.n1236 GND 0.001783f
C1897 VDD.n1237 GND 0.001783f
C1898 VDD.n1238 GND 0.001783f
C1899 VDD.n1239 GND 0.001783f
C1900 VDD.n1240 GND 0.001435f
C1901 VDD.n1241 GND 0.001783f
C1902 VDD.n1243 GND 0.001783f
C1903 VDD.n1245 GND 0.001783f
C1904 VDD.n1246 GND 0.001435f
C1905 VDD.n1247 GND 7.39e-19
C1906 VDD.n1248 GND 0.001783f
C1907 VDD.n1249 GND 0.001783f
C1908 VDD.n1250 GND 9.4e-19
C1909 VDD.n1251 GND 0.001783f
C1910 VDD.n1253 GND 0.001783f
C1911 VDD.n1255 GND 0.001783f
C1912 VDD.n1256 GND 0.001435f
C1913 VDD.n1257 GND 0.001783f
C1914 VDD.n1258 GND 0.001783f
C1915 VDD.n1259 GND 0.001783f
C1916 VDD.n1260 GND 0.001435f
C1917 VDD.n1261 GND 0.001783f
C1918 VDD.n1263 GND 0.001783f
C1919 VDD.n1265 GND 0.001783f
C1920 VDD.n1266 GND 0.001435f
C1921 VDD.n1267 GND 0.001783f
C1922 VDD.n1268 GND 0.001783f
C1923 VDD.n1269 GND 0.001783f
C1924 VDD.n1270 GND 0.001435f
C1925 VDD.n1271 GND 0.001783f
C1926 VDD.n1273 GND 0.001783f
C1927 VDD.n1274 GND 0.001783f
C1928 VDD.n1276 GND 0.001783f
C1929 VDD.n1277 GND 0.001435f
C1930 VDD.n1278 GND 0.001783f
C1931 VDD.n1279 GND 0.001783f
C1932 VDD.n1280 GND 0.001783f
C1933 VDD.n1281 GND 0.001227f
C1934 VDD.n1282 GND 0.002928f
C1935 VDD.n1283 GND 9.26e-19
C1936 VDD.n1284 GND 0.004059f
C1937 VDD.n1285 GND 0.003894f
C1938 VDD.n1286 GND 0.001191f
C1939 VDD.n1287 GND 0.003894f
C1940 VDD.n1288 GND 0.22766f
C1941 VDD.n1289 GND 0.003894f
C1942 VDD.n1290 GND 0.001191f
C1943 VDD.n1291 GND 0.003894f
C1944 VDD.n1292 GND 0.001783f
C1945 VDD.n1293 GND 0.001783f
C1946 VDD.n1294 GND 0.001435f
C1947 VDD.n1295 GND 0.001783f
C1948 VDD.n1296 GND 0.158648f
C1949 VDD.n1297 GND 0.001783f
C1950 VDD.n1298 GND 0.001435f
C1951 VDD.n1299 GND 0.001783f
C1952 VDD.n1300 GND 0.001783f
C1953 VDD.n1301 GND 0.001783f
C1954 VDD.n1302 GND 0.001435f
C1955 VDD.n1303 GND 0.001783f
C1956 VDD.n1304 GND 0.107881f
C1957 VDD.n1305 GND 0.001783f
C1958 VDD.n1306 GND 0.001435f
C1959 VDD.n1307 GND 0.001783f
C1960 VDD.n1308 GND 0.001783f
C1961 VDD.n1309 GND 0.001783f
C1962 VDD.n1310 GND 0.001435f
C1963 VDD.n1311 GND 0.001783f
C1964 VDD.n1312 GND 0.158648f
C1965 VDD.n1313 GND 0.001783f
C1966 VDD.n1314 GND 0.001435f
C1967 VDD.n1315 GND 0.001783f
C1968 VDD.n1316 GND 0.001783f
C1969 VDD.n1317 GND 0.001783f
C1970 VDD.n1318 GND 0.001435f
C1971 VDD.n1319 GND 0.001783f
C1972 VDD.n1320 GND 0.158648f
C1973 VDD.n1321 GND 0.001783f
C1974 VDD.n1322 GND 0.001435f
C1975 VDD.n1323 GND 0.001783f
C1976 VDD.n1324 GND 0.001783f
C1977 VDD.n1325 GND 0.001783f
C1978 VDD.n1326 GND 0.001435f
C1979 VDD.n1327 GND 0.001783f
C1980 VDD.n1328 GND 0.158648f
C1981 VDD.n1329 GND 0.001783f
C1982 VDD.n1330 GND 0.001435f
C1983 VDD.n1331 GND 0.001783f
C1984 VDD.n1332 GND 0.001783f
C1985 VDD.n1333 GND 0.001783f
C1986 VDD.n1334 GND 0.001435f
C1987 VDD.n1335 GND 0.001783f
C1988 VDD.n1336 GND 0.158648f
C1989 VDD.n1337 GND 0.001783f
C1990 VDD.n1338 GND 0.001435f
C1991 VDD.n1339 GND 0.001777f
C1992 VDD.n1340 GND 0.001005f
C1993 VDD.n1341 GND 9.08e-19
C1994 VDD.n1342 GND 4.88e-19
C1995 VDD.n1343 GND 0.001153f
C1996 VDD.n1344 GND 5.17e-19
C1997 VDD.n1345 GND 0.003542f
C1998 VDD.t141 GND 0.002562f
C1999 VDD.n1346 GND 8.65e-19
C2000 VDD.n1347 GND 7.25e-19
C2001 VDD.n1348 GND 4.88e-19
C2002 VDD.n1349 GND 0.012395f
C2003 VDD.n1350 GND 9.08e-19
C2004 VDD.n1351 GND 4.88e-19
C2005 VDD.n1352 GND 5.17e-19
C2006 VDD.n1353 GND 0.001153f
C2007 VDD.n1354 GND 0.002818f
C2008 VDD.n1355 GND 5.17e-19
C2009 VDD.n1356 GND 4.88e-19
C2010 VDD.n1357 GND 0.002285f
C2011 VDD.n1358 GND 0.005716f
C2012 VDD.n1359 GND 0.001005f
C2013 VDD.n1360 GND 9.08e-19
C2014 VDD.n1361 GND 4.88e-19
C2015 VDD.n1362 GND 0.001153f
C2016 VDD.n1363 GND 5.17e-19
C2017 VDD.n1364 GND 0.003542f
C2018 VDD.t133 GND 0.002562f
C2019 VDD.n1365 GND 8.65e-19
C2020 VDD.n1366 GND 7.25e-19
C2021 VDD.n1367 GND 4.88e-19
C2022 VDD.n1368 GND 0.012395f
C2023 VDD.n1369 GND 9.08e-19
C2024 VDD.n1370 GND 4.88e-19
C2025 VDD.n1371 GND 5.17e-19
C2026 VDD.n1372 GND 0.001153f
C2027 VDD.n1373 GND 0.002818f
C2028 VDD.n1374 GND 5.17e-19
C2029 VDD.n1375 GND 4.88e-19
C2030 VDD.n1376 GND 0.002285f
C2031 VDD.n1377 GND 0.004436f
C2032 VDD.n1378 GND 0.097672f
C2033 VDD.n1379 GND 0.001005f
C2034 VDD.n1380 GND 9.08e-19
C2035 VDD.n1381 GND 4.88e-19
C2036 VDD.n1382 GND 0.001153f
C2037 VDD.n1383 GND 5.17e-19
C2038 VDD.n1384 GND 0.003542f
C2039 VDD.t103 GND 0.002562f
C2040 VDD.n1385 GND 8.65e-19
C2041 VDD.n1386 GND 7.25e-19
C2042 VDD.n1387 GND 4.88e-19
C2043 VDD.n1388 GND 0.012395f
C2044 VDD.n1389 GND 9.08e-19
C2045 VDD.n1390 GND 4.88e-19
C2046 VDD.n1391 GND 5.17e-19
C2047 VDD.n1392 GND 0.001153f
C2048 VDD.n1393 GND 0.002818f
C2049 VDD.n1394 GND 5.17e-19
C2050 VDD.n1395 GND 4.88e-19
C2051 VDD.n1396 GND 0.002285f
C2052 VDD.n1397 GND 0.004436f
C2053 VDD.n1398 GND 0.05756f
C2054 VDD.n1399 GND 0.001005f
C2055 VDD.n1400 GND 9.08e-19
C2056 VDD.n1401 GND 4.88e-19
C2057 VDD.n1402 GND 0.001153f
C2058 VDD.n1403 GND 5.17e-19
C2059 VDD.n1404 GND 0.003542f
C2060 VDD.t99 GND 0.002562f
C2061 VDD.n1405 GND 8.65e-19
C2062 VDD.n1406 GND 7.25e-19
C2063 VDD.n1407 GND 4.88e-19
C2064 VDD.n1408 GND 0.012395f
C2065 VDD.n1409 GND 9.08e-19
C2066 VDD.n1410 GND 4.88e-19
C2067 VDD.n1411 GND 5.17e-19
C2068 VDD.n1412 GND 0.001153f
C2069 VDD.n1413 GND 0.002818f
C2070 VDD.n1414 GND 5.17e-19
C2071 VDD.n1415 GND 4.88e-19
C2072 VDD.n1416 GND 0.002285f
C2073 VDD.n1417 GND 0.004436f
C2074 VDD.n1418 GND 0.05756f
C2075 VDD.n1419 GND 0.001005f
C2076 VDD.n1420 GND 9.08e-19
C2077 VDD.n1421 GND 4.88e-19
C2078 VDD.n1422 GND 0.001153f
C2079 VDD.n1423 GND 5.17e-19
C2080 VDD.n1424 GND 0.003542f
C2081 VDD.t104 GND 0.002562f
C2082 VDD.n1425 GND 8.65e-19
C2083 VDD.n1426 GND 7.25e-19
C2084 VDD.n1427 GND 4.88e-19
C2085 VDD.n1428 GND 0.012395f
C2086 VDD.n1429 GND 9.08e-19
C2087 VDD.n1430 GND 4.88e-19
C2088 VDD.n1431 GND 5.17e-19
C2089 VDD.n1432 GND 0.001153f
C2090 VDD.n1433 GND 0.002818f
C2091 VDD.n1434 GND 5.17e-19
C2092 VDD.n1435 GND 4.88e-19
C2093 VDD.n1436 GND 0.002285f
C2094 VDD.n1437 GND 0.004436f
C2095 VDD.n1438 GND 0.054484f
C2096 VDD.n1439 GND 0.411326f
C2097 VDD.n1440 GND 0.003335f
C2098 VDD.n1441 GND 0.001777f
C2099 VDD.n1442 GND 0.001435f
C2100 VDD.n1443 GND 0.001783f
C2101 VDD.n1444 GND 0.158648f
C2102 VDD.n1445 GND 0.001783f
C2103 VDD.n1446 GND 0.001435f
C2104 VDD.n1447 GND 0.001783f
C2105 VDD.n1448 GND 0.001783f
C2106 VDD.n1449 GND 0.001783f
C2107 VDD.n1450 GND 0.001435f
C2108 VDD.n1451 GND 0.001783f
C2109 VDD.n1452 GND 0.158648f
C2110 VDD.n1453 GND 0.001783f
C2111 VDD.n1454 GND 0.001435f
C2112 VDD.n1455 GND 0.001783f
C2113 VDD.n1456 GND 0.001783f
C2114 VDD.n1457 GND 0.001783f
C2115 VDD.n1458 GND 0.001435f
C2116 VDD.n1459 GND 0.001783f
C2117 VDD.n1460 GND 0.158648f
C2118 VDD.n1461 GND 0.001783f
C2119 VDD.n1462 GND 0.001435f
C2120 VDD.n1463 GND 0.001783f
C2121 VDD.n1464 GND 0.001783f
C2122 VDD.n1465 GND 0.001783f
C2123 VDD.n1466 GND 0.001435f
C2124 VDD.n1467 GND 0.001783f
C2125 VDD.n1468 GND 0.158648f
C2126 VDD.n1469 GND 0.001783f
C2127 VDD.n1470 GND 0.001435f
C2128 VDD.n1471 GND 0.001783f
C2129 VDD.n1472 GND 0.001783f
C2130 VDD.n1473 GND 0.001783f
C2131 VDD.n1474 GND 0.001435f
C2132 VDD.n1475 GND 0.001783f
C2133 VDD.n1476 GND 0.107881f
C2134 VDD.n1477 GND 0.001783f
C2135 VDD.n1478 GND 0.001435f
C2136 VDD.n1479 GND 0.001783f
C2137 VDD.n1480 GND 0.001783f
C2138 VDD.n1481 GND 0.004059f
C2139 VDD.n1482 GND 0.003894f
C2140 VDD.n1483 GND 0.001783f
C2141 VDD.n1484 GND 0.001783f
C2142 VDD.n1485 GND 0.001435f
C2143 VDD.n1486 GND 0.001783f
C2144 VDD.n1487 GND 0.158648f
C2145 VDD.n1488 GND 0.001783f
C2146 VDD.n1489 GND 0.001435f
C2147 VDD.n1490 GND 0.001783f
C2148 VDD.n1491 GND 0.001783f
C2149 VDD.n1492 GND 0.001783f
C2150 VDD.n1494 GND 0.001783f
C2151 VDD.n1495 GND 0.001783f
C2152 VDD.n1496 GND 0.001435f
C2153 VDD.n1497 GND 0.001435f
C2154 VDD.n1498 GND 0.001783f
C2155 VDD.n1499 GND 0.001783f
C2156 VDD.n1500 GND 0.001783f
C2157 VDD.n1501 GND 0.001783f
C2158 VDD.n1502 GND 0.001783f
C2159 VDD.n1503 GND 0.001783f
C2160 VDD.n1504 GND 0.001435f
C2161 VDD.n1506 GND 0.001783f
C2162 VDD.n1507 GND 0.001783f
C2163 VDD.n1508 GND 0.001783f
C2164 VDD.n1509 GND 0.001783f
C2165 VDD.t84 GND 0.010031f
C2166 VDD.t83 GND 0.014304f
C2167 VDD.t82 GND 0.109243f
C2168 VDD.n1510 GND 0.024442f
C2169 VDD.n1511 GND 0.019628f
C2170 VDD.n1513 GND 0.001783f
C2171 VDD.n1514 GND 0.001783f
C2172 VDD.n1515 GND 0.001783f
C2173 VDD.n1516 GND 0.001435f
C2174 VDD.n1517 GND 0.001435f
C2175 VDD.n1519 GND 0.001783f
C2176 VDD.n1520 GND 0.001783f
C2177 VDD.n1521 GND 0.001783f
C2178 VDD.n1522 GND 0.001783f
C2179 VDD.n1523 GND 0.001783f
C2180 VDD.n1524 GND 0.001435f
C2181 VDD.n1525 GND 0.001435f
C2182 VDD.n1526 GND 0.001783f
C2183 VDD.n1528 GND 0.001783f
C2184 VDD.n1529 GND 0.001783f
C2185 VDD.n1531 GND 0.001783f
C2186 VDD.n1532 GND 9.69e-19
C2187 VDD.n1533 GND 0.002928f
C2188 VDD.n1534 GND 0.001428f
C2189 VDD.n1535 GND 0.001435f
C2190 VDD.n1536 GND 0.001783f
C2191 VDD.n1538 GND 0.001783f
C2192 VDD.n1539 GND 0.001783f
C2193 VDD.n1540 GND 0.001435f
C2194 VDD.n1541 GND 0.001435f
C2195 VDD.n1542 GND 0.001435f
C2196 VDD.n1543 GND 0.001783f
C2197 VDD.n1545 GND 0.001783f
C2198 VDD.n1546 GND 0.001783f
C2199 VDD.n1548 GND 0.001783f
C2200 VDD.n1549 GND 0.001435f
C2201 VDD.n1550 GND 0.001435f
C2202 VDD.n1551 GND 0.001191f
C2203 VDD.n1552 GND 0.004059f
C2204 VDD.n1553 GND 0.003894f
C2205 VDD.n1554 GND 0.001191f
C2206 VDD.n1555 GND 0.003894f
C2207 VDD.n1556 GND 0.22766f
C2208 VDD.n1557 GND 0.003894f
C2209 VDD.n1558 GND 0.004059f
C2210 VDD.n1560 GND 0.001783f
C2211 VDD.n1561 GND 0.002928f
C2212 VDD.n1562 GND 0.001227f
C2213 VDD.n1563 GND 0.001783f
C2214 VDD.n1564 GND 0.001783f
C2215 VDD.n1565 GND 0.001783f
C2216 VDD.n1566 GND 0.001435f
C2217 VDD.n1567 GND 0.001435f
C2218 VDD.n1568 GND 0.001435f
C2219 VDD.n1569 GND 0.001783f
C2220 VDD.n1570 GND 0.001783f
C2221 VDD.n1571 GND 0.001783f
C2222 VDD.n1572 GND 0.001435f
C2223 VDD.n1573 GND 0.001435f
C2224 VDD.n1574 GND 0.001435f
C2225 VDD.n1575 GND 0.001783f
C2226 VDD.n1576 GND 0.001783f
C2227 VDD.n1577 GND 0.001783f
C2228 VDD.n1578 GND 0.001435f
C2229 VDD.n1579 GND 0.001435f
C2230 VDD.n1580 GND 9.4e-19
C2231 VDD.n1581 GND 0.001783f
C2232 VDD.n1582 GND 0.001783f
C2233 VDD.n1583 GND 7.39e-19
C2234 VDD.n1584 GND 0.001435f
C2235 VDD.n1585 GND 0.001435f
C2236 VDD.n1586 GND 0.001052f
C2237 VDD.n1587 GND 0.584215f
C2238 VDD.n1589 GND 0.001435f
C2239 VDD.n1590 GND 0.001783f
C2240 VDD.n1592 GND 0.001783f
C2241 VDD.n1593 GND 0.001783f
C2242 VDD.n1594 GND 0.001435f
C2243 VDD.n1595 GND 0.001435f
C2244 VDD.n1596 GND 0.001435f
C2245 VDD.n1597 GND 0.001783f
C2246 VDD.n1599 GND 0.001783f
C2247 VDD.n1600 GND 0.001783f
C2248 VDD.n1601 GND 0.001435f
C2249 VDD.n1602 GND 0.001783f
C2250 VDD.n1603 GND 0.001783f
C2251 VDD.n1604 GND 0.001783f
C2252 VDD.n1605 GND 0.002928f
C2253 VDD.n1606 GND 9.69e-19
C2254 VDD.n1607 GND 0.001435f
C2255 VDD.n1608 GND 0.001783f
C2256 VDD.n1610 GND 0.001783f
C2257 VDD.n1611 GND 0.001783f
C2258 VDD.n1612 GND 0.001435f
C2259 VDD.n1613 GND 0.001435f
C2260 VDD.n1614 GND 0.001435f
C2261 VDD.n1615 GND 0.001783f
C2262 VDD.n1617 GND 0.001783f
C2263 VDD.n1618 GND 0.001783f
C2264 VDD.n1619 GND 0.001435f
C2265 VDD.n1620 GND 0.001435f
C2266 VDD.n1621 GND 0.001435f
C2267 VDD.n1622 GND 0.001783f
C2268 VDD.n1624 GND 0.001783f
C2269 VDD.n1625 GND 0.001783f
C2270 VDD.n1626 GND 0.001435f
C2271 VDD.n1627 GND 0.001783f
C2272 VDD.n1628 GND 0.001783f
C2273 VDD.n1629 GND 0.001783f
C2274 VDD.n1630 GND 0.002928f
C2275 VDD.n1631 GND 0.001783f
C2276 VDD.n1633 GND 0.001783f
C2277 VDD.n1634 GND 0.001783f
C2278 VDD.n1635 GND 0.001435f
C2279 VDD.n1636 GND 0.001435f
C2280 VDD.n1637 GND 0.001435f
C2281 VDD.n1638 GND 0.001783f
C2282 VDD.n1640 GND 0.001783f
C2283 VDD.n1641 GND 0.001783f
C2284 VDD.n1643 GND 0.001783f
C2285 VDD.n1644 GND 0.001435f
C2286 VDD.n1646 GND 0.584215f
C2287 VDD.t12 GND 0.00872f
C2288 VDD.t13 GND 0.013318f
C2289 VDD.t10 GND 0.116692f
C2290 VDD.n1647 GND 0.016902f
C2291 VDD.n1648 GND 0.011832f
C2292 VDD.n1649 GND 0.001212f
C2293 VDD.n1650 GND 0.001212f
C2294 VDD.n1651 GND 0.001212f
C2295 VDD.n1652 GND 0.001212f
C2296 VDD.n1653 GND 0.001212f
C2297 VDD.n1654 GND 0.001212f
C2298 VDD.n1655 GND 0.001212f
C2299 VDD.n1656 GND 0.001212f
C2300 VDD.n1657 GND 0.001212f
C2301 VDD.n1658 GND 0.001212f
C2302 VDD.n1659 GND 0.001212f
C2303 VDD.n1660 GND 0.001212f
C2304 VDD.n1661 GND 0.001212f
C2305 VDD.n1662 GND 0.001212f
C2306 VDD.n1663 GND 0.001212f
C2307 VDD.n1664 GND 0.001212f
C2308 VDD.n1665 GND 0.001212f
C2309 VDD.n1666 GND 0.001212f
C2310 VDD.n1667 GND 0.001212f
C2311 VDD.n1668 GND 0.001212f
C2312 VDD.n1669 GND 0.001212f
C2313 VDD.n1670 GND 0.001212f
C2314 VDD.n1671 GND 0.001212f
C2315 VDD.n1672 GND 0.001212f
C2316 VDD.n1673 GND 0.001212f
C2317 VDD.n1674 GND 0.001212f
C2318 VDD.n1675 GND 0.001212f
C2319 VDD.n1676 GND 0.001212f
C2320 VDD.n1677 GND 0.001212f
C2321 VDD.n1678 GND 0.001212f
C2322 VDD.n1679 GND 0.001212f
C2323 VDD.n1680 GND 0.001212f
C2324 VDD.n1681 GND 0.001212f
C2325 VDD.n1682 GND 0.001212f
C2326 VDD.n1683 GND 0.001212f
C2327 VDD.n1684 GND 0.001212f
C2328 VDD.n1685 GND 0.001212f
C2329 VDD.n1686 GND 0.001212f
C2330 VDD.n1687 GND 0.001212f
C2331 VDD.n1688 GND 0.001212f
C2332 VDD.n1689 GND 0.001212f
C2333 VDD.n1690 GND 0.001212f
C2334 VDD.n1691 GND 0.001212f
C2335 VDD.n1692 GND 0.001212f
C2336 VDD.n1693 GND 0.001212f
C2337 VDD.n1694 GND 0.001212f
C2338 VDD.n1695 GND 0.001212f
C2339 VDD.n1696 GND 0.001212f
C2340 VDD.n1697 GND 0.001212f
C2341 VDD.n1698 GND 0.001212f
C2342 VDD.n1699 GND 0.001212f
C2343 VDD.n1700 GND 0.001212f
C2344 VDD.n1701 GND 0.001212f
C2345 VDD.n1702 GND 0.001212f
C2346 VDD.n1703 GND 0.001212f
C2347 VDD.n1704 GND 0.001212f
C2348 VDD.n1705 GND 0.001212f
C2349 VDD.n1706 GND 0.001212f
C2350 VDD.n1707 GND 0.001212f
C2351 VDD.n1708 GND 0.001212f
C2352 VDD.n1709 GND 0.001212f
C2353 VDD.n1710 GND 0.001212f
C2354 VDD.n1711 GND 0.001212f
C2355 VDD.n1712 GND 0.001212f
C2356 VDD.n1713 GND 0.001212f
C2357 VDD.n1714 GND 0.001212f
C2358 VDD.n1715 GND 0.001212f
C2359 VDD.n1716 GND 0.001212f
C2360 VDD.n1717 GND 0.001212f
C2361 VDD.n1718 GND 0.001212f
C2362 VDD.n1719 GND 0.001212f
C2363 VDD.n1720 GND 0.001212f
C2364 VDD.n1721 GND 0.001212f
C2365 VDD.n1722 GND 0.001212f
C2366 VDD.n1723 GND 0.001212f
C2367 VDD.n1724 GND 0.001212f
C2368 VDD.n1725 GND 0.001212f
C2369 VDD.n1726 GND 0.001212f
C2370 VDD.n1727 GND 0.001212f
C2371 VDD.n1728 GND 0.001212f
C2372 VDD.n1729 GND 0.001212f
C2373 VDD.n1730 GND 0.001212f
C2374 VDD.n1731 GND 0.001212f
C2375 VDD.n1732 GND 0.001212f
C2376 VDD.n1733 GND 0.001212f
C2377 VDD.n1734 GND 0.001212f
C2378 VDD.n1735 GND 0.001212f
C2379 VDD.n1736 GND 0.001212f
C2380 VDD.n1737 GND 0.001212f
C2381 VDD.n1738 GND 0.001212f
C2382 VDD.n1739 GND 0.001212f
C2383 VDD.n1740 GND 0.001212f
C2384 VDD.n1741 GND 0.001212f
C2385 VDD.n1742 GND 0.001212f
C2386 VDD.n1743 GND 0.001212f
C2387 VDD.n1744 GND 0.001212f
C2388 VDD.n1745 GND 0.001212f
C2389 VDD.n1746 GND 0.001212f
C2390 VDD.n1747 GND 0.001212f
C2391 VDD.n1748 GND 0.001212f
C2392 VDD.n1749 GND 0.001212f
C2393 VDD.n1750 GND 0.001212f
C2394 VDD.n1751 GND 0.001212f
C2395 VDD.n1752 GND 0.001212f
C2396 VDD.n1753 GND 0.001212f
C2397 VDD.n1754 GND 0.001212f
C2398 VDD.n1755 GND 0.001212f
C2399 VDD.n1756 GND 0.001212f
C2400 VDD.n1757 GND 0.001212f
C2401 VDD.n1758 GND 0.001212f
C2402 VDD.n1759 GND 0.001212f
C2403 VDD.n1760 GND 0.001212f
C2404 VDD.n1761 GND 0.001212f
C2405 VDD.n1762 GND 0.001212f
C2406 VDD.n1763 GND 0.001212f
C2407 VDD.n1764 GND 0.001212f
C2408 VDD.n1765 GND 0.001212f
C2409 VDD.n1766 GND 0.001212f
C2410 VDD.n1767 GND 0.001212f
C2411 VDD.n1768 GND 0.002794f
C2412 VDD.n1769 GND 0.002794f
C2413 VDD.n1770 GND 0.002965f
C2414 VDD.n1771 GND 0.002965f
C2415 VDD.n1772 GND 0.001212f
C2416 VDD.n1773 GND 0.001212f
C2417 VDD.n1774 GND 0.001212f
C2418 VDD.n1775 GND 8.74e-19
C2419 VDD.n1776 GND 0.001733f
C2420 VDD.n1777 GND 9.45e-19
C2421 VDD.n1778 GND 0.001212f
C2422 VDD.n1779 GND 0.001212f
C2423 VDD.n1780 GND 0.001212f
C2424 VDD.n1781 GND 0.001212f
C2425 VDD.n1782 GND 0.001212f
C2426 VDD.n1783 GND 0.001212f
C2427 VDD.n1784 GND 0.001212f
C2428 VDD.n1785 GND 0.065701f
C2429 VDD.n1786 GND 0.001212f
C2430 VDD.n1787 GND 0.001212f
C2431 VDD.n1788 GND 0.001212f
C2432 VDD.n1789 GND 0.001212f
C2433 VDD.n1790 GND 0.001212f
C2434 VDD.n1791 GND 0.001212f
C2435 VDD.n1792 GND 0.001212f
C2436 VDD.n1793 GND 0.001212f
C2437 VDD.n1794 GND 0.001212f
C2438 VDD.n1795 GND 0.001212f
C2439 VDD.n1796 GND 0.70281f
C2440 VDD.n1798 GND 0.002965f
C2441 VDD.n1799 GND 0.002965f
C2442 VDD.n1800 GND 0.002794f
C2443 VDD.n1801 GND 0.001212f
C2444 VDD.n1802 GND 0.001212f
C2445 VDD.n1803 GND 0.107881f
C2446 VDD.n1804 GND 0.001212f
C2447 VDD.n1805 GND 0.001212f
C2448 VDD.n1806 GND 0.001212f
C2449 VDD.n1807 GND 0.001212f
C2450 VDD.n1808 GND 0.001212f
C2451 VDD.n1809 GND 0.107881f
C2452 VDD.n1810 GND 0.001212f
C2453 VDD.n1811 GND 0.001212f
C2454 VDD.n1812 GND 0.001212f
C2455 VDD.n1813 GND 0.001212f
C2456 VDD.n1814 GND 0.001212f
C2457 VDD.n1815 GND 0.107881f
C2458 VDD.n1816 GND 0.001212f
C2459 VDD.n1817 GND 0.001212f
C2460 VDD.n1818 GND 0.001212f
C2461 VDD.n1819 GND 0.001212f
C2462 VDD.n1820 GND 0.001212f
C2463 VDD.n1821 GND 0.107881f
C2464 VDD.n1822 GND 0.001212f
C2465 VDD.n1823 GND 0.001212f
C2466 VDD.n1824 GND 0.001212f
C2467 VDD.n1825 GND 0.001212f
C2468 VDD.n1826 GND 0.001212f
C2469 VDD.n1827 GND 0.107881f
C2470 VDD.n1828 GND 0.001212f
C2471 VDD.n1829 GND 0.001212f
C2472 VDD.n1830 GND 0.001212f
C2473 VDD.n1831 GND 0.001212f
C2474 VDD.n1832 GND 0.001212f
C2475 VDD.n1833 GND 0.098362f
C2476 VDD.n1834 GND 0.001212f
C2477 VDD.n1835 GND 0.001212f
C2478 VDD.n1836 GND 0.001212f
C2479 VDD.n1837 GND 0.001212f
C2480 VDD.n1838 GND 0.001212f
C2481 VDD.n1839 GND 0.107881f
C2482 VDD.n1840 GND 0.001212f
C2483 VDD.n1841 GND 0.001212f
C2484 VDD.n1842 GND 0.001212f
C2485 VDD.n1843 GND 0.001212f
C2486 VDD.n1844 GND 0.001212f
C2487 VDD.n1845 GND 0.067425f
C2488 VDD.n1846 GND 0.001212f
C2489 VDD.n1847 GND 0.001212f
C2490 VDD.n1848 GND 0.001212f
C2491 VDD.n1849 GND 0.001212f
C2492 VDD.n1850 GND 0.001212f
C2493 VDD.n1851 GND 0.107881f
C2494 VDD.n1852 GND 0.001212f
C2495 VDD.n1853 GND 0.001212f
C2496 VDD.n1854 GND 0.001212f
C2497 VDD.n1855 GND 0.001212f
C2498 VDD.n1856 GND 0.001212f
C2499 VDD.n1857 GND 0.107881f
C2500 VDD.n1858 GND 0.001212f
C2501 VDD.n1859 GND 0.001212f
C2502 VDD.n1860 GND 0.001212f
C2503 VDD.n1861 GND 0.001212f
C2504 VDD.n1862 GND 0.001212f
C2505 VDD.n1863 GND 0.107881f
C2506 VDD.n1864 GND 0.001212f
C2507 VDD.n1865 GND 0.001212f
C2508 VDD.n1866 GND 0.001212f
C2509 VDD.n1867 GND 0.001212f
C2510 VDD.n1868 GND 0.001212f
C2511 VDD.n1869 GND 0.107881f
C2512 VDD.n1870 GND 0.001212f
C2513 VDD.n1871 GND 0.001212f
C2514 VDD.n1872 GND 0.001212f
C2515 VDD.n1873 GND 0.001212f
C2516 VDD.n1874 GND 0.001212f
C2517 VDD.n1875 GND 0.107881f
C2518 VDD.n1876 GND 0.001212f
C2519 VDD.n1877 GND 0.001212f
C2520 VDD.n1878 GND 0.001212f
C2521 VDD.n1879 GND 0.001212f
C2522 VDD.n1880 GND 0.001212f
C2523 VDD.n1881 GND 0.107881f
C2524 VDD.n1882 GND 0.001212f
C2525 VDD.n1883 GND 0.001212f
C2526 VDD.n1884 GND 0.001212f
C2527 VDD.n1885 GND 0.001212f
C2528 VDD.n1886 GND 0.001212f
C2529 VDD.n1887 GND 0.107881f
C2530 VDD.n1888 GND 0.001212f
C2531 VDD.n1889 GND 0.001212f
C2532 VDD.n1890 GND 0.001212f
C2533 VDD.n1891 GND 0.001212f
C2534 VDD.n1892 GND 0.001212f
C2535 VDD.n1893 GND 0.096775f
C2536 VDD.n1894 GND 0.001212f
C2537 VDD.n1895 GND 0.001212f
C2538 VDD.n1896 GND 0.001212f
C2539 VDD.n1897 GND 0.001212f
C2540 VDD.n1898 GND 0.001212f
C2541 VDD.n1899 GND 0.062666f
C2542 VDD.n1900 GND 0.001212f
C2543 VDD.n1901 GND 0.001212f
C2544 VDD.n1902 GND 0.001212f
C2545 VDD.n1903 GND 0.001212f
C2546 VDD.n1904 GND 0.001212f
C2547 VDD.n1905 GND 0.107881f
C2548 VDD.n1906 GND 0.001212f
C2549 VDD.n1907 GND 0.001212f
C2550 VDD.n1908 GND 0.001212f
C2551 VDD.n1909 GND 0.001212f
C2552 VDD.n1910 GND 0.001212f
C2553 VDD.n1911 GND 0.107881f
C2554 VDD.n1912 GND 0.001212f
C2555 VDD.n1913 GND 0.001212f
C2556 VDD.n1914 GND 0.001212f
C2557 VDD.n1915 GND 0.001212f
C2558 VDD.n1916 GND 0.001212f
C2559 VDD.n1917 GND 0.107881f
C2560 VDD.n1918 GND 0.001212f
C2561 VDD.n1919 GND 0.001212f
C2562 VDD.n1920 GND 0.001212f
C2563 VDD.n1921 GND 0.001212f
C2564 VDD.n1922 GND 0.001212f
C2565 VDD.n1923 GND 0.107881f
C2566 VDD.n1924 GND 0.001212f
C2567 VDD.n1925 GND 0.001212f
C2568 VDD.n1926 GND 0.001212f
C2569 VDD.n1927 GND 0.001212f
C2570 VDD.n1928 GND 0.001212f
C2571 VDD.n1929 GND 0.107881f
C2572 VDD.n1930 GND 0.001212f
C2573 VDD.n1931 GND 0.001212f
C2574 VDD.n1932 GND 0.001212f
C2575 VDD.n1933 GND 0.001212f
C2576 VDD.n1934 GND 0.001212f
C2577 VDD.n1935 GND 0.107881f
C2578 VDD.n1936 GND 0.001212f
C2579 VDD.n1937 GND 0.001212f
C2580 VDD.n1938 GND 0.001212f
C2581 VDD.n1939 GND 0.001212f
C2582 VDD.n1940 GND 0.001212f
C2583 VDD.n1941 GND 0.107881f
C2584 VDD.n1942 GND 0.001212f
C2585 VDD.n1943 GND 0.001212f
C2586 VDD.n1944 GND 0.001212f
C2587 VDD.n1945 GND 0.001212f
C2588 VDD.n1946 GND 0.001212f
C2589 VDD.n1947 GND 0.107881f
C2590 VDD.n1948 GND 0.001212f
C2591 VDD.n1949 GND 0.001212f
C2592 VDD.n1950 GND 0.001212f
C2593 VDD.n1951 GND 0.001212f
C2594 VDD.n1952 GND 0.001212f
C2595 VDD.n1953 GND 0.073771f
C2596 VDD.n1954 GND 0.001212f
C2597 VDD.n1955 GND 0.001212f
C2598 VDD.n1956 GND 0.001212f
C2599 VDD.n1957 GND 0.001212f
C2600 VDD.n1958 GND 0.001212f
C2601 VDD.n1959 GND 0.107881f
C2602 VDD.n1960 GND 0.001212f
C2603 VDD.n1961 GND 0.001212f
C2604 VDD.n1962 GND 0.001212f
C2605 VDD.n1963 GND 0.001212f
C2606 VDD.n1964 GND 0.001212f
C2607 VDD.n1965 GND 0.107881f
C2608 VDD.n1966 GND 0.001212f
C2609 VDD.n1967 GND 0.001212f
C2610 VDD.n1968 GND 0.001212f
C2611 VDD.n1969 GND 0.001212f
C2612 VDD.n1970 GND 0.001212f
C2613 VDD.n1971 GND 0.107881f
C2614 VDD.n1972 GND 0.001212f
C2615 VDD.n1973 GND 0.001212f
C2616 VDD.n1974 GND 0.001212f
C2617 VDD.n1975 GND 0.001212f
C2618 VDD.n1976 GND 0.001212f
C2619 VDD.n1977 GND 0.107881f
C2620 VDD.n1978 GND 0.001212f
C2621 VDD.n1979 GND 0.001212f
C2622 VDD.n1980 GND 0.001212f
C2623 VDD.n1981 GND 0.001212f
C2624 VDD.n1982 GND 0.001212f
C2625 VDD.n1983 GND 0.107881f
C2626 VDD.n1984 GND 0.001212f
C2627 VDD.n1985 GND 0.001212f
C2628 VDD.n1986 GND 0.001212f
C2629 VDD.n1987 GND 0.001212f
C2630 VDD.n1988 GND 0.001212f
C2631 VDD.n1989 GND 0.107881f
C2632 VDD.n1990 GND 0.001212f
C2633 VDD.n1991 GND 0.001212f
C2634 VDD.n1992 GND 0.001212f
C2635 VDD.n1993 GND 0.001212f
C2636 VDD.n1994 GND 0.001212f
C2637 VDD.n1995 GND 0.107881f
C2638 VDD.n1996 GND 0.001212f
C2639 VDD.n1997 GND 0.001212f
C2640 VDD.n1998 GND 0.001212f
C2641 VDD.n1999 GND 0.001212f
C2642 VDD.n2000 GND 0.001212f
C2643 VDD.n2001 GND 0.107881f
C2644 VDD.n2002 GND 0.001212f
C2645 VDD.n2003 GND 0.001212f
C2646 VDD.n2004 GND 0.001212f
C2647 VDD.n2005 GND 0.001212f
C2648 VDD.n2006 GND 0.001212f
C2649 VDD.n2007 GND 0.107087f
C2650 VDD.n2008 GND 0.001212f
C2651 VDD.n2009 GND 0.001212f
C2652 VDD.n2010 GND 0.001212f
C2653 VDD.n2011 GND 0.001212f
C2654 VDD.n2012 GND 0.001212f
C2655 VDD.n2013 GND 0.098362f
C2656 VDD.n2014 GND 0.001212f
C2657 VDD.n2015 GND 0.001212f
C2658 VDD.n2016 GND 0.001212f
C2659 VDD.n2017 GND 0.001212f
C2660 VDD.n2018 GND 0.001212f
C2661 VDD.n2019 GND 0.107881f
C2662 VDD.n2020 GND 0.001212f
C2663 VDD.n2021 GND 0.001212f
C2664 VDD.n2022 GND 0.001212f
C2665 VDD.n2023 GND 0.001212f
C2666 VDD.n2024 GND 0.001212f
C2667 VDD.n2025 GND 0.001212f
C2668 VDD.n2026 GND 0.001212f
C2669 VDD.n2027 GND 0.107881f
C2670 VDD.n2028 GND 0.001212f
C2671 VDD.n2029 GND 0.001212f
C2672 VDD.n2030 GND 0.001212f
C2673 VDD.n2031 GND 0.001212f
C2674 VDD.n2032 GND 0.001212f
C2675 VDD.n2033 GND 0.107881f
C2676 VDD.n2034 GND 0.001212f
C2677 VDD.n2035 GND 0.001212f
C2678 VDD.n2036 GND 0.001212f
C2679 VDD.n2037 GND 0.001212f
C2680 VDD.n2038 GND 0.001212f
C2681 VDD.n2039 GND 0.001212f
C2682 VDD.n2040 GND 0.001212f
C2683 VDD.n2041 GND 0.002794f
C2684 VDD.n2042 GND 0.002934f
C2685 VDD.n2043 GND 0.002825f
C2686 VDD.n2044 GND 0.001212f
C2687 VDD.n2045 GND 0.001212f
C2688 VDD.n2046 GND 8.74e-19
C2689 VDD.n2047 GND 0.001212f
C2690 VDD.n2048 GND 0.001212f
C2691 VDD.n2049 GND 9.45e-19
C2692 VDD.n2050 GND 0.001212f
C2693 VDD.n2051 GND 0.001212f
C2694 VDD.n2052 GND 0.001212f
C2695 VDD.n2053 GND 0.001212f
C2696 VDD.n2054 GND 0.001212f
C2697 VDD.n2055 GND 0.001212f
C2698 VDD.n2056 GND 0.001212f
C2699 VDD.n2057 GND 0.001212f
C2700 VDD.n2058 GND 0.001212f
C2701 VDD.n2059 GND 0.001212f
C2702 VDD.n2060 GND 0.001212f
C2703 VDD.n2061 GND 0.001212f
C2704 VDD.n2062 GND 0.001212f
C2705 VDD.n2063 GND 0.001212f
C2706 VDD.n2064 GND 0.001212f
C2707 VDD.n2065 GND 0.001212f
C2708 VDD.n2066 GND 0.001212f
C2709 VDD.n2067 GND 0.001212f
C2710 VDD.n2068 GND 0.001212f
C2711 VDD.n2069 GND 0.001212f
C2712 VDD.n2070 GND 0.002965f
C2713 VDD.n2071 GND 0.002965f
C2714 VDD.n2072 GND 0.002794f
C2715 VDD.n2073 GND 0.002794f
C2716 VDD.n2074 GND 0.001212f
C2717 VDD.n2075 GND 0.001212f
C2718 VDD.n2076 GND 0.001212f
C2719 VDD.n2077 GND 0.001212f
C2720 VDD.n2078 GND 0.107881f
C2721 VDD.n2079 GND 0.001212f
C2722 VDD.n2080 GND 0.001212f
C2723 VDD.n2081 GND 0.001212f
C2724 VDD.n2082 GND 0.001212f
C2725 VDD.n2083 GND 0.001212f
C2726 VDD.n2084 GND 0.107881f
C2727 VDD.n2085 GND 0.001212f
C2728 VDD.n2086 GND 0.002794f
C2729 VDD.n2087 GND 0.002965f
C2730 VDD.n2088 GND 0.002825f
C2731 VDD.n2089 GND 0.001212f
C2732 VDD.n2090 GND 0.001212f
C2733 VDD.n2091 GND 0.001212f
C2734 VDD.n2092 GND 8.74e-19
C2735 VDD.n2093 GND 0.001733f
C2736 VDD.n2094 GND 9.45e-19
C2737 VDD.n2095 GND 0.001212f
C2738 VDD.n2096 GND 0.001212f
C2739 VDD.n2097 GND 0.001212f
C2740 VDD.n2098 GND 0.001212f
C2741 VDD.n2099 GND 0.001212f
C2742 VDD.n2100 GND 0.001212f
C2743 VDD.n2101 GND 0.001212f
C2744 VDD.n2102 GND 0.001212f
C2745 VDD.n2103 GND 0.001212f
C2746 VDD.n2104 GND 0.001212f
C2747 VDD.n2105 GND 0.001212f
C2748 VDD.n2106 GND 0.001212f
C2749 VDD.n2107 GND 0.001212f
C2750 VDD.n2108 GND 0.001212f
C2751 VDD.n2109 GND 0.001212f
C2752 VDD.n2110 GND 0.001212f
C2753 VDD.n2111 GND 0.001212f
C2754 VDD.n2112 GND 0.001212f
C2755 VDD.n2113 GND 0.001212f
C2756 VDD.n2114 GND 0.001212f
C2757 VDD.n2115 GND 0.002965f
C2758 VDD.n2116 GND 0.002965f
C2759 VDD.n2117 GND 0.680599f
C2760 VDD.n2130 GND 0.001212f
C2761 VDD.n2131 GND 0.002794f
C2762 VDD.t89 GND 0.00872f
C2763 VDD.t90 GND 0.013318f
C2764 VDD.t88 GND 0.116692f
C2765 VDD.n2132 GND 0.016902f
C2766 VDD.n2133 GND 0.011832f
C2767 VDD.n2134 GND 0.001733f
C2768 VDD.n2135 GND 0.001212f
C2769 VDD.n2136 GND 0.001212f
C2770 VDD.n2137 GND 0.001212f
C2771 VDD.n2138 GND 0.001212f
C2772 VDD.n2139 GND 0.001212f
C2773 VDD.n2140 GND 0.001212f
C2774 VDD.n2141 GND 0.001212f
C2775 VDD.n2142 GND 0.001212f
C2776 VDD.n2143 GND 0.001212f
C2777 VDD.n2144 GND 0.001212f
C2778 VDD.n2145 GND 0.001212f
C2779 VDD.n2146 GND 0.001212f
C2780 VDD.n2147 GND 0.001212f
C2781 VDD.n2148 GND 0.001212f
C2782 VDD.n2149 GND 0.001212f
C2783 VDD.n2150 GND 0.001212f
C2784 VDD.n2151 GND 0.001212f
C2785 VDD.n2152 GND 0.001212f
C2786 VDD.n2153 GND 9.45e-19
C2787 VDD.n2154 GND 0.001212f
C2788 VDD.n2155 GND 0.001212f
C2789 VDD.n2156 GND 8.74e-19
C2790 VDD.n2157 GND 0.001212f
C2791 VDD.n2158 GND 0.001212f
C2792 VDD.n2159 GND 0.001212f
C2793 VDD.n2160 GND 0.001212f
C2794 VDD.n2161 GND 0.001212f
C2795 VDD.n2162 GND 0.001212f
C2796 VDD.n2163 GND 0.001212f
C2797 VDD.n2164 GND 0.001212f
C2798 VDD.n2165 GND 0.001212f
C2799 VDD.n2166 GND 0.001212f
C2800 VDD.n2167 GND 0.001212f
C2801 VDD.n2168 GND 0.001212f
C2802 VDD.n2169 GND 0.001212f
C2803 VDD.n2170 GND 0.001212f
C2804 VDD.n2171 GND 0.001212f
C2805 VDD.n2172 GND 0.001212f
C2806 VDD.n2173 GND 0.001212f
C2807 VDD.n2174 GND 0.001212f
C2808 VDD.n2175 GND 0.001212f
C2809 VDD.n2176 GND 0.001212f
C2810 VDD.n2177 GND 0.001212f
C2811 VDD.n2178 GND 0.001212f
C2812 VDD.n2179 GND 0.001212f
C2813 VDD.n2180 GND 0.001212f
C2814 VDD.n2181 GND 0.001212f
C2815 VDD.n2182 GND 0.001212f
C2816 VDD.n2183 GND 0.001212f
C2817 VDD.n2184 GND 0.001212f
C2818 VDD.n2185 GND 0.001212f
C2819 VDD.n2186 GND 0.001212f
C2820 VDD.n2187 GND 0.001212f
C2821 VDD.n2188 GND 0.001212f
C2822 VDD.n2189 GND 0.001212f
C2823 VDD.n2190 GND 0.001212f
C2824 VDD.n2191 GND 0.001212f
C2825 VDD.n2192 GND 0.001212f
C2826 VDD.n2193 GND 0.001212f
C2827 VDD.n2194 GND 0.001212f
C2828 VDD.n2195 GND 0.001212f
C2829 VDD.n2196 GND 0.001212f
C2830 VDD.n2197 GND 0.001212f
C2831 VDD.n2198 GND 0.001212f
C2832 VDD.n2199 GND 0.001212f
C2833 VDD.n2200 GND 0.001212f
C2834 VDD.n2201 GND 0.001212f
C2835 VDD.n2202 GND 0.001212f
C2836 VDD.n2203 GND 0.001212f
C2837 VDD.n2204 GND 0.001212f
C2838 VDD.n2205 GND 0.001212f
C2839 VDD.n2206 GND 0.001212f
C2840 VDD.n2207 GND 0.001212f
C2841 VDD.n2208 GND 0.001212f
C2842 VDD.n2209 GND 0.001212f
C2843 VDD.n2210 GND 0.001212f
C2844 VDD.n2211 GND 0.001212f
C2845 VDD.n2212 GND 0.001212f
C2846 VDD.n2213 GND 0.001212f
C2847 VDD.n2214 GND 0.001212f
C2848 VDD.n2215 GND 0.001212f
C2849 VDD.n2216 GND 0.001212f
C2850 VDD.n2217 GND 0.001212f
C2851 VDD.n2218 GND 0.001212f
C2852 VDD.n2219 GND 0.001212f
C2853 VDD.n2220 GND 0.001212f
C2854 VDD.n2221 GND 0.001212f
C2855 VDD.n2222 GND 0.001212f
C2856 VDD.n2223 GND 0.001212f
C2857 VDD.n2224 GND 0.001212f
C2858 VDD.n2225 GND 0.001212f
C2859 VDD.n2226 GND 0.001212f
C2860 VDD.n2227 GND 0.001212f
C2861 VDD.n2228 GND 0.001212f
C2862 VDD.n2229 GND 0.001212f
C2863 VDD.n2230 GND 0.001212f
C2864 VDD.n2231 GND 0.001212f
C2865 VDD.n2232 GND 0.001212f
C2866 VDD.n2233 GND 0.001212f
C2867 VDD.n2234 GND 0.001212f
C2868 VDD.n2235 GND 0.001212f
C2869 VDD.n2236 GND 0.001212f
C2870 VDD.n2237 GND 0.001212f
C2871 VDD.n2238 GND 0.001212f
C2872 VDD.n2239 GND 0.001212f
C2873 VDD.n2240 GND 0.001212f
C2874 VDD.n2241 GND 0.001212f
C2875 VDD.n2242 GND 0.001212f
C2876 VDD.n2243 GND 0.001212f
C2877 VDD.n2244 GND 0.001212f
C2878 VDD.n2245 GND 0.001212f
C2879 VDD.n2246 GND 0.001212f
C2880 VDD.n2247 GND 0.001212f
C2881 VDD.n2248 GND 0.001212f
C2882 VDD.n2249 GND 0.001212f
C2883 VDD.n2250 GND 0.001212f
C2884 VDD.n2251 GND 0.001212f
C2885 VDD.n2252 GND 0.001212f
C2886 VDD.n2253 GND 0.001212f
C2887 VDD.n2254 GND 0.001212f
C2888 VDD.n2255 GND 0.001212f
C2889 VDD.n2256 GND 0.001212f
C2890 VDD.n2257 GND 0.001212f
C2891 VDD.n2258 GND 0.001212f
C2892 VDD.n2259 GND 0.001212f
C2893 VDD.n2260 GND 0.001212f
C2894 VDD.n2261 GND 0.001212f
C2895 VDD.n2262 GND 0.001212f
C2896 VDD.n2263 GND 0.001212f
C2897 VDD.n2264 GND 0.001212f
C2898 VDD.n2265 GND 0.001212f
C2899 VDD.n2266 GND 0.001212f
C2900 VDD.n2267 GND 0.001212f
C2901 VDD.n2268 GND 0.001212f
C2902 VDD.n2269 GND 0.001212f
C2903 VDD.n2270 GND 0.001212f
C2904 VDD.n2271 GND 0.001212f
C2905 VDD.n2272 GND 0.001212f
C2906 VDD.n2273 GND 0.001212f
C2907 VDD.n2274 GND 0.001212f
C2908 VDD.n2275 GND 0.001212f
C2909 VDD.n2276 GND 0.002794f
C2910 VDD.n2277 GND 0.002965f
C2911 VDD.n2278 GND 0.002965f
C2912 VDD.n2279 GND 0.001212f
C2913 VDD.n2280 GND 0.001212f
C2914 VDD.t62 GND 0.00872f
C2915 VDD.t63 GND 0.013318f
C2916 VDD.t60 GND 0.116692f
C2917 VDD.n2281 GND 0.016902f
C2918 VDD.n2282 GND 0.011832f
C2919 VDD.n2283 GND 0.001212f
C2920 VDD.n2284 GND 0.001212f
C2921 VDD.n2285 GND 0.001212f
C2922 VDD.n2286 GND 0.001212f
C2923 VDD.n2287 GND 0.001212f
C2924 VDD.n2288 GND 0.001212f
C2925 VDD.n2289 GND 0.001212f
C2926 VDD.n2290 GND 0.001212f
C2927 VDD.n2291 GND 0.001212f
C2928 VDD.n2292 GND 0.001212f
C2929 VDD.n2293 GND 0.001212f
C2930 VDD.n2294 GND 0.001212f
C2931 VDD.n2295 GND 0.001212f
C2932 VDD.n2296 GND 0.001212f
C2933 VDD.n2297 GND 0.001212f
C2934 VDD.n2298 GND 0.001212f
C2935 VDD.n2299 GND 0.001212f
C2936 VDD.n2300 GND 0.001212f
C2937 VDD.n2301 GND 0.001212f
C2938 VDD.n2302 GND 0.001212f
C2939 VDD.n2303 GND 0.001212f
C2940 VDD.n2304 GND 0.001212f
C2941 VDD.n2305 GND 0.001212f
C2942 VDD.n2306 GND 0.001212f
C2943 VDD.n2307 GND 0.001212f
C2944 VDD.n2308 GND 0.001212f
C2945 VDD.n2309 GND 0.001212f
C2946 VDD.n2310 GND 0.001212f
C2947 VDD.n2311 GND 0.001212f
C2948 VDD.n2312 GND 0.001212f
C2949 VDD.n2313 GND 0.001212f
C2950 VDD.n2314 GND 0.001212f
C2951 VDD.n2315 GND 0.001212f
C2952 VDD.n2316 GND 0.001212f
C2953 VDD.n2317 GND 0.001212f
C2954 VDD.n2318 GND 0.001212f
C2955 VDD.n2319 GND 0.001212f
C2956 VDD.n2320 GND 0.001212f
C2957 VDD.n2321 GND 0.001212f
C2958 VDD.n2322 GND 0.001212f
C2959 VDD.n2323 GND 0.001212f
C2960 VDD.n2324 GND 0.001212f
C2961 VDD.n2325 GND 0.001212f
C2962 VDD.n2326 GND 0.001212f
C2963 VDD.n2327 GND 0.001212f
C2964 VDD.n2328 GND 0.001212f
C2965 VDD.n2329 GND 0.001212f
C2966 VDD.n2330 GND 0.001212f
C2967 VDD.n2331 GND 0.001212f
C2968 VDD.n2332 GND 0.001212f
C2969 VDD.n2333 GND 0.001212f
C2970 VDD.n2334 GND 0.001212f
C2971 VDD.n2335 GND 0.001212f
C2972 VDD.n2336 GND 0.001212f
C2973 VDD.n2337 GND 0.001212f
C2974 VDD.n2338 GND 0.001212f
C2975 VDD.n2339 GND 0.001212f
C2976 VDD.n2340 GND 0.001212f
C2977 VDD.n2341 GND 0.001212f
C2978 VDD.n2342 GND 0.001212f
C2979 VDD.n2343 GND 0.001212f
C2980 VDD.n2344 GND 0.001212f
C2981 VDD.n2345 GND 0.001212f
C2982 VDD.n2346 GND 0.001212f
C2983 VDD.n2347 GND 0.001212f
C2984 VDD.n2348 GND 0.001212f
C2985 VDD.n2349 GND 0.001212f
C2986 VDD.n2350 GND 0.001212f
C2987 VDD.n2351 GND 0.001212f
C2988 VDD.n2352 GND 0.001212f
C2989 VDD.n2353 GND 0.001212f
C2990 VDD.n2354 GND 0.001212f
C2991 VDD.n2355 GND 0.001212f
C2992 VDD.n2356 GND 0.001212f
C2993 VDD.n2357 GND 0.001212f
C2994 VDD.n2358 GND 0.001212f
C2995 VDD.n2359 GND 0.001212f
C2996 VDD.n2360 GND 0.001212f
C2997 VDD.n2361 GND 0.001212f
C2998 VDD.n2362 GND 0.001212f
C2999 VDD.n2363 GND 0.001212f
C3000 VDD.n2364 GND 0.001212f
C3001 VDD.n2365 GND 0.001212f
C3002 VDD.n2366 GND 0.001212f
C3003 VDD.n2367 GND 0.001212f
C3004 VDD.n2368 GND 0.001212f
C3005 VDD.n2369 GND 0.001212f
C3006 VDD.n2370 GND 0.001212f
C3007 VDD.n2371 GND 0.001212f
C3008 VDD.n2372 GND 0.001212f
C3009 VDD.n2373 GND 0.001212f
C3010 VDD.n2374 GND 0.001212f
C3011 VDD.n2375 GND 0.001212f
C3012 VDD.n2376 GND 0.001212f
C3013 VDD.n2377 GND 0.001212f
C3014 VDD.n2378 GND 0.001212f
C3015 VDD.n2379 GND 0.001212f
C3016 VDD.n2380 GND 0.001212f
C3017 VDD.n2381 GND 0.001212f
C3018 VDD.n2382 GND 0.001212f
C3019 VDD.n2383 GND 0.001212f
C3020 VDD.n2384 GND 0.001212f
C3021 VDD.n2385 GND 0.001212f
C3022 VDD.n2386 GND 0.001212f
C3023 VDD.n2387 GND 0.001212f
C3024 VDD.n2388 GND 0.001212f
C3025 VDD.n2389 GND 0.001212f
C3026 VDD.n2390 GND 0.001212f
C3027 VDD.n2391 GND 0.001212f
C3028 VDD.n2392 GND 0.001212f
C3029 VDD.n2393 GND 0.001212f
C3030 VDD.n2394 GND 0.001212f
C3031 VDD.n2395 GND 0.001212f
C3032 VDD.n2396 GND 0.001212f
C3033 VDD.n2397 GND 0.001212f
C3034 VDD.n2398 GND 0.001212f
C3035 VDD.n2399 GND 0.002794f
C3036 VDD.n2400 GND 0.002794f
C3037 VDD.n2401 GND 0.002965f
C3038 VDD.n2402 GND 0.002965f
C3039 VDD.n2403 GND 0.001212f
C3040 VDD.n2404 GND 0.001212f
C3041 VDD.n2405 GND 0.001212f
C3042 VDD.n2406 GND 8.74e-19
C3043 VDD.n2407 GND 0.001733f
C3044 VDD.n2408 GND 9.45e-19
C3045 VDD.n2409 GND 0.001212f
C3046 VDD.n2410 GND 0.001212f
C3047 VDD.n2411 GND 0.001212f
C3048 VDD.n2412 GND 0.001212f
C3049 VDD.n2413 GND 0.001212f
C3050 VDD.n2414 GND 0.001212f
C3051 VDD.n2415 GND 0.001212f
C3052 VDD.n2416 GND 0.001212f
C3053 VDD.n2417 GND 0.001212f
C3054 VDD.n2418 GND 0.001212f
C3055 VDD.n2419 GND 0.001212f
C3056 VDD.n2420 GND 0.001212f
C3057 VDD.n2421 GND 0.001212f
C3058 VDD.n2422 GND 0.001212f
C3059 VDD.n2423 GND 0.001212f
C3060 VDD.n2424 GND 0.001212f
C3061 VDD.n2425 GND 0.001212f
C3062 VDD.n2426 GND 0.001212f
C3063 VDD.n2427 GND 0.001212f
C3064 VDD.n2428 GND 0.002965f
C3065 VDD.n2429 GND 0.002965f
C3066 VDD.n2431 GND 0.680599f
C3067 VDD.n2433 GND 0.002965f
C3068 VDD.n2434 GND 0.002965f
C3069 VDD.n2435 GND 0.002794f
C3070 VDD.n2436 GND 0.001212f
C3071 VDD.n2437 GND 0.001212f
C3072 VDD.n2438 GND 0.107881f
C3073 VDD.n2439 GND 0.001212f
C3074 VDD.n2440 GND 0.001212f
C3075 VDD.n2441 GND 0.001212f
C3076 VDD.n2442 GND 0.001212f
C3077 VDD.n2443 GND 0.001212f
C3078 VDD.n2444 GND 0.107881f
C3079 VDD.n2445 GND 0.001212f
C3080 VDD.n2446 GND 0.001212f
C3081 VDD.n2447 GND 0.001212f
C3082 VDD.n2448 GND 0.001212f
C3083 VDD.n2449 GND 0.001212f
C3084 VDD.n2450 GND 0.107881f
C3085 VDD.n2451 GND 0.001212f
C3086 VDD.n2452 GND 0.001212f
C3087 VDD.n2453 GND 0.001212f
C3088 VDD.n2454 GND 0.001212f
C3089 VDD.n2455 GND 0.001212f
C3090 VDD.n2456 GND 0.107881f
C3091 VDD.n2457 GND 0.001212f
C3092 VDD.n2458 GND 0.001212f
C3093 VDD.n2459 GND 0.001212f
C3094 VDD.n2460 GND 0.001212f
C3095 VDD.n2461 GND 0.001212f
C3096 VDD.n2462 GND 0.107881f
C3097 VDD.n2463 GND 0.001212f
C3098 VDD.n2464 GND 0.001212f
C3099 VDD.n2465 GND 0.001212f
C3100 VDD.n2466 GND 0.001212f
C3101 VDD.n2467 GND 0.001212f
C3102 VDD.n2468 GND 0.098362f
C3103 VDD.n2469 GND 0.001212f
C3104 VDD.n2470 GND 0.001212f
C3105 VDD.n2471 GND 0.001212f
C3106 VDD.n2472 GND 0.001212f
C3107 VDD.n2473 GND 0.001212f
C3108 VDD.n2474 GND 0.107087f
C3109 VDD.n2475 GND 0.001212f
C3110 VDD.n2476 GND 0.001212f
C3111 VDD.n2477 GND 0.001212f
C3112 VDD.n2478 GND 0.001212f
C3113 VDD.n2479 GND 0.001212f
C3114 VDD.n2480 GND 0.107881f
C3115 VDD.n2481 GND 0.001212f
C3116 VDD.n2482 GND 0.001212f
C3117 VDD.n2483 GND 0.001212f
C3118 VDD.n2484 GND 0.001212f
C3119 VDD.n2485 GND 0.001212f
C3120 VDD.n2486 GND 0.107881f
C3121 VDD.n2487 GND 0.001212f
C3122 VDD.n2488 GND 0.001212f
C3123 VDD.n2489 GND 0.001212f
C3124 VDD.n2490 GND 0.001212f
C3125 VDD.n2491 GND 0.001212f
C3126 VDD.n2492 GND 0.107881f
C3127 VDD.n2493 GND 0.001212f
C3128 VDD.n2494 GND 0.001212f
C3129 VDD.n2495 GND 0.001212f
C3130 VDD.n2496 GND 0.001212f
C3131 VDD.n2497 GND 0.001212f
C3132 VDD.n2498 GND 0.107881f
C3133 VDD.n2499 GND 0.001212f
C3134 VDD.n2500 GND 0.001212f
C3135 VDD.n2501 GND 0.001212f
C3136 VDD.n2502 GND 0.001212f
C3137 VDD.n2503 GND 0.001212f
C3138 VDD.n2504 GND 0.107881f
C3139 VDD.n2505 GND 0.001212f
C3140 VDD.n2506 GND 0.001212f
C3141 VDD.n2507 GND 0.001212f
C3142 VDD.n2508 GND 0.001212f
C3143 VDD.n2509 GND 0.001212f
C3144 VDD.n2510 GND 0.107881f
C3145 VDD.n2511 GND 0.001212f
C3146 VDD.n2512 GND 0.001212f
C3147 VDD.n2513 GND 0.001212f
C3148 VDD.n2514 GND 0.001212f
C3149 VDD.n2515 GND 0.001212f
C3150 VDD.n2516 GND 0.107881f
C3151 VDD.n2517 GND 0.001212f
C3152 VDD.n2518 GND 0.001212f
C3153 VDD.n2519 GND 0.001212f
C3154 VDD.n2520 GND 0.001212f
C3155 VDD.n2521 GND 0.001212f
C3156 VDD.n2522 GND 0.107881f
C3157 VDD.n2523 GND 0.001212f
C3158 VDD.n2524 GND 0.001212f
C3159 VDD.n2525 GND 0.001212f
C3160 VDD.n2526 GND 0.001212f
C3161 VDD.n2527 GND 0.001212f
C3162 VDD.n2528 GND 0.073771f
C3163 VDD.n2529 GND 0.001212f
C3164 VDD.n2530 GND 0.001212f
C3165 VDD.n2531 GND 0.001212f
C3166 VDD.n2532 GND 0.001212f
C3167 VDD.n2533 GND 0.001212f
C3168 VDD.n2534 GND 0.107881f
C3169 VDD.n2535 GND 0.001212f
C3170 VDD.n2536 GND 0.001212f
C3171 VDD.n2537 GND 0.001212f
C3172 VDD.n2538 GND 0.001212f
C3173 VDD.n2539 GND 0.001212f
C3174 VDD.n2540 GND 0.107881f
C3175 VDD.n2541 GND 0.001212f
C3176 VDD.n2542 GND 0.001212f
C3177 VDD.n2543 GND 0.001212f
C3178 VDD.n2544 GND 0.001212f
C3179 VDD.n2545 GND 0.001212f
C3180 VDD.n2546 GND 0.107881f
C3181 VDD.n2547 GND 0.001212f
C3182 VDD.n2548 GND 0.001212f
C3183 VDD.n2549 GND 0.001212f
C3184 VDD.n2550 GND 0.001212f
C3185 VDD.n2551 GND 0.001212f
C3186 VDD.n2552 GND 0.107881f
C3187 VDD.n2553 GND 0.001212f
C3188 VDD.n2554 GND 0.001212f
C3189 VDD.n2555 GND 0.001212f
C3190 VDD.n2556 GND 0.001212f
C3191 VDD.n2557 GND 0.001212f
C3192 VDD.n2558 GND 0.107881f
C3193 VDD.n2559 GND 0.001212f
C3194 VDD.n2560 GND 0.001212f
C3195 VDD.n2561 GND 0.001212f
C3196 VDD.n2562 GND 0.001212f
C3197 VDD.n2563 GND 0.001212f
C3198 VDD.n2564 GND 0.107881f
C3199 VDD.n2565 GND 0.001212f
C3200 VDD.n2566 GND 0.001212f
C3201 VDD.n2567 GND 0.001212f
C3202 VDD.n2568 GND 0.001212f
C3203 VDD.n2569 GND 0.001212f
C3204 VDD.n2570 GND 0.107881f
C3205 VDD.n2571 GND 0.001212f
C3206 VDD.n2572 GND 0.001212f
C3207 VDD.n2573 GND 0.001212f
C3208 VDD.n2574 GND 0.001212f
C3209 VDD.n2575 GND 0.001212f
C3210 VDD.n2576 GND 0.107881f
C3211 VDD.n2577 GND 0.001212f
C3212 VDD.n2578 GND 0.001212f
C3213 VDD.n2579 GND 0.001212f
C3214 VDD.n2580 GND 0.001212f
C3215 VDD.n2581 GND 0.001212f
C3216 VDD.n2582 GND 0.062666f
C3217 VDD.n2583 GND 0.001212f
C3218 VDD.n2584 GND 0.001212f
C3219 VDD.n2585 GND 0.001212f
C3220 VDD.n2586 GND 0.001212f
C3221 VDD.n2587 GND 0.001212f
C3222 VDD.n2588 GND 0.096775f
C3223 VDD.n2589 GND 0.001212f
C3224 VDD.n2590 GND 0.001212f
C3225 VDD.n2591 GND 0.001212f
C3226 VDD.n2592 GND 0.001212f
C3227 VDD.n2593 GND 0.001212f
C3228 VDD.n2594 GND 0.107881f
C3229 VDD.n2595 GND 0.001212f
C3230 VDD.n2596 GND 0.001212f
C3231 VDD.n2597 GND 0.001212f
C3232 VDD.n2598 GND 0.001212f
C3233 VDD.n2599 GND 0.001212f
C3234 VDD.n2600 GND 0.107881f
C3235 VDD.n2601 GND 0.001212f
C3236 VDD.n2602 GND 0.001212f
C3237 VDD.n2603 GND 0.001212f
C3238 VDD.n2604 GND 0.001212f
C3239 VDD.n2605 GND 0.001212f
C3240 VDD.n2606 GND 0.107881f
C3241 VDD.n2607 GND 0.001212f
C3242 VDD.n2608 GND 0.001212f
C3243 VDD.n2609 GND 0.001212f
C3244 VDD.n2610 GND 0.001212f
C3245 VDD.n2611 GND 0.001212f
C3246 VDD.n2612 GND 0.107881f
C3247 VDD.n2613 GND 0.001212f
C3248 VDD.n2614 GND 0.001212f
C3249 VDD.n2615 GND 0.001212f
C3250 VDD.n2616 GND 0.001212f
C3251 VDD.n2617 GND 0.001212f
C3252 VDD.n2618 GND 0.107881f
C3253 VDD.n2619 GND 0.001212f
C3254 VDD.n2620 GND 0.001212f
C3255 VDD.n2621 GND 0.001212f
C3256 VDD.n2622 GND 0.001212f
C3257 VDD.n2623 GND 0.001212f
C3258 VDD.n2624 GND 0.107881f
C3259 VDD.n2625 GND 0.001212f
C3260 VDD.n2626 GND 0.001212f
C3261 VDD.n2627 GND 0.001212f
C3262 VDD.n2628 GND 0.001212f
C3263 VDD.n2629 GND 0.001212f
C3264 VDD.n2630 GND 0.107881f
C3265 VDD.n2631 GND 0.001212f
C3266 VDD.n2632 GND 0.001212f
C3267 VDD.n2633 GND 0.001212f
C3268 VDD.n2634 GND 0.001212f
C3269 VDD.n2635 GND 0.001212f
C3270 VDD.n2636 GND 0.067425f
C3271 VDD.n2637 GND 0.001212f
C3272 VDD.n2638 GND 0.001212f
C3273 VDD.n2639 GND 0.001212f
C3274 VDD.n2640 GND 0.001212f
C3275 VDD.n2641 GND 0.001212f
C3276 VDD.n2642 GND 0.107881f
C3277 VDD.n2643 GND 0.001212f
C3278 VDD.n2644 GND 0.001212f
C3279 VDD.n2645 GND 0.001212f
C3280 VDD.n2646 GND 0.001212f
C3281 VDD.n2647 GND 0.001212f
C3282 VDD.n2648 GND 0.098362f
C3283 VDD.n2649 GND 0.001212f
C3284 VDD.n2650 GND 0.001212f
C3285 VDD.n2651 GND 0.001212f
C3286 VDD.n2652 GND 0.001212f
C3287 VDD.n2653 GND 0.001212f
C3288 VDD.n2654 GND 0.107881f
C3289 VDD.n2655 GND 0.001212f
C3290 VDD.n2656 GND 0.001212f
C3291 VDD.n2657 GND 0.001212f
C3292 VDD.n2658 GND 0.001212f
C3293 VDD.n2659 GND 0.001212f
C3294 VDD.n2660 GND 0.107881f
C3295 VDD.n2661 GND 0.001212f
C3296 VDD.n2662 GND 0.001212f
C3297 VDD.n2663 GND 0.001212f
C3298 VDD.n2664 GND 0.002965f
C3299 VDD.n2665 GND 0.001212f
C3300 VDD.n2666 GND 0.001212f
C3301 VDD.n2667 GND 0.001212f
C3302 VDD.n2670 GND 0.001212f
C3303 VDD.n2671 GND 0.001212f
C3304 VDD.n2672 GND 0.001212f
C3305 VDD.n2673 GND 0.001212f
C3306 VDD.n2674 GND 0.001212f
C3307 VDD.n2675 GND 0.001212f
C3308 VDD.n2677 GND 0.001212f
C3309 VDD.n2678 GND 0.002965f
C3310 VDD.n2679 GND 0.002794f
C3311 VDD.n2680 GND 0.002794f
C3312 VDD.n2681 GND 0.001212f
C3313 VDD.n2682 GND 0.001212f
C3314 VDD.n2683 GND 0.001212f
C3315 VDD.n2684 GND 0.001212f
C3316 VDD.n2685 GND 0.001212f
C3317 VDD.n2686 GND 0.001212f
C3318 VDD.n2687 GND 0.001212f
C3319 VDD.n2688 GND 0.107881f
C3320 VDD.n2689 GND 0.001212f
C3321 VDD.n2690 GND 0.001212f
C3322 VDD.n2691 GND 0.001212f
C3323 VDD.n2692 GND 0.001212f
C3324 VDD.n2693 GND 0.001212f
C3325 VDD.n2694 GND 0.107881f
C3326 VDD.n2695 GND 0.001212f
C3327 VDD.n2696 GND 0.001212f
C3328 VDD.n2697 GND 0.001212f
C3329 VDD.n2698 GND 0.001212f
C3330 VDD.n2699 GND 0.002934f
C3331 VDD.n2700 GND 0.002825f
C3332 VDD.n2701 GND 0.002965f
C3333 VDD.n2703 GND 0.001212f
C3334 VDD.n2704 GND 0.001212f
C3335 VDD.n2705 GND 8.74e-19
C3336 VDD.n2706 GND 0.001733f
C3337 VDD.n2707 GND 9.45e-19
C3338 VDD.n2708 GND 0.001212f
C3339 VDD.n2709 GND 0.001212f
C3340 VDD.n2711 GND 0.001212f
C3341 VDD.n2712 GND 0.001212f
C3342 VDD.n2713 GND 0.001212f
C3343 VDD.n2714 GND 0.584801f
C3344 VDD.n2715 GND 0.065115f
C3345 VDD.n2716 GND 0.001212f
C3346 VDD.n2717 GND 0.001212f
C3347 VDD.n2719 GND 0.001212f
C3348 VDD.n2720 GND 0.001212f
C3349 VDD.n2721 GND 0.001212f
C3350 VDD.n2722 GND 0.001212f
C3351 VDD.n2723 GND 0.001212f
C3352 VDD.n2724 GND 0.001212f
C3353 VDD.n2726 GND 0.001212f
C3354 VDD.n2727 GND 0.002965f
C3355 VDD.n2728 GND 0.002965f
C3356 VDD.n2729 GND 0.002794f
C3357 VDD.n2730 GND 0.001212f
C3358 VDD.n2731 GND 0.001212f
C3359 VDD.n2732 GND 0.107881f
C3360 VDD.n2733 GND 0.001212f
C3361 VDD.n2734 GND 0.001212f
C3362 VDD.n2735 GND 0.002934f
C3363 VDD.n2736 GND 0.002825f
C3364 VDD.n2737 GND 0.002965f
C3365 VDD.n2739 GND 0.001212f
C3366 VDD.n2740 GND 0.001212f
C3367 VDD.n2741 GND 8.74e-19
C3368 VDD.n2742 GND 0.001733f
C3369 VDD.n2743 GND 9.45e-19
C3370 VDD.n2744 GND 0.001212f
C3371 VDD.n2745 GND 0.001212f
C3372 VDD.n2747 GND 0.001212f
C3373 VDD.n2748 GND 0.001212f
C3374 VDD.n2750 GND 0.001212f
C3375 VDD.n2751 GND 0.065115f
C3376 VDD.n2752 GND 0.584801f
C3377 VDD.n2753 GND 0.001052f
C3378 VDD.n2754 GND 0.001783f
C3379 VDD.n2755 GND 0.001783f
C3380 VDD.t41 GND 0.010031f
C3381 VDD.t42 GND 0.014304f
C3382 VDD.t40 GND 0.109243f
C3383 VDD.n2756 GND 0.024442f
C3384 VDD.n2757 GND 0.019628f
C3385 VDD.n2758 GND 0.00221f
C3386 VDD.n2759 GND 0.001783f
C3387 VDD.n2760 GND 0.001783f
C3388 VDD.n2761 GND 0.001783f
C3389 VDD.n2762 GND 0.001783f
C3390 VDD.n2763 GND 0.001783f
C3391 VDD.n2764 GND 0.001783f
C3392 VDD.n2765 GND 0.001783f
C3393 VDD.n2766 GND 0.001783f
C3394 VDD.n2767 GND 0.001783f
C3395 VDD.n2768 GND 0.001783f
C3396 VDD.n2769 GND 0.001783f
C3397 VDD.n2770 GND 0.001783f
C3398 VDD.n2771 GND 0.001783f
C3399 VDD.n2772 GND 0.001227f
C3400 VDD.n2773 GND 0.001783f
C3401 VDD.n2774 GND 0.001783f
C3402 VDD.n2775 GND 0.001435f
C3403 VDD.n2776 GND 0.001435f
C3404 VDD.n2777 GND 0.001783f
C3405 VDD.n2778 GND 0.001783f
C3406 VDD.n2779 GND 0.001435f
C3407 VDD.n2780 GND 0.001435f
C3408 VDD.n2781 GND 0.001783f
C3409 VDD.n2782 GND 0.001783f
C3410 VDD.n2783 GND 0.001435f
C3411 VDD.n2784 GND 0.001435f
C3412 VDD.n2785 GND 0.001783f
C3413 VDD.n2786 GND 0.001783f
C3414 VDD.n2787 GND 0.001435f
C3415 VDD.n2788 GND 0.001435f
C3416 VDD.n2789 GND 0.001783f
C3417 VDD.n2790 GND 0.001783f
C3418 VDD.n2791 GND 0.001435f
C3419 VDD.n2792 GND 0.001435f
C3420 VDD.n2793 GND 0.001783f
C3421 VDD.n2794 GND 0.001783f
C3422 VDD.n2795 GND 0.001435f
C3423 VDD.n2796 GND 9.4e-19
C3424 VDD.n2797 GND 0.001783f
C3425 VDD.n2798 GND 0.001783f
C3426 VDD.n2799 GND 7.39e-19
C3427 VDD.n2800 GND 0.001435f
C3428 VDD.n2801 GND 0.001783f
C3429 VDD.n2802 GND 0.001783f
C3430 VDD.n2803 GND 0.001435f
C3431 VDD.n2804 GND 0.001435f
C3432 VDD.n2805 GND 0.001783f
C3433 VDD.n2806 GND 0.001783f
C3434 VDD.n2807 GND 0.001435f
C3435 VDD.n2808 GND 0.001435f
C3436 VDD.n2809 GND 0.001783f
C3437 VDD.n2810 GND 0.001783f
C3438 VDD.n2811 GND 0.001435f
C3439 VDD.n2812 GND 0.001435f
C3440 VDD.n2813 GND 0.001783f
C3441 VDD.n2814 GND 0.001783f
C3442 VDD.n2815 GND 0.001435f
C3443 VDD.n2816 GND 0.001435f
C3444 VDD.n2817 GND 0.001783f
C3445 VDD.n2818 GND 0.001783f
C3446 VDD.n2819 GND 0.001435f
C3447 VDD.n2820 GND 0.001783f
C3448 VDD.n2821 GND 0.001783f
C3449 VDD.n2822 GND 0.001435f
C3450 VDD.n2823 GND 0.001783f
C3451 VDD.n2824 GND 0.001783f
C3452 VDD.n2825 GND 0.001783f
C3453 VDD.n2826 GND 0.002928f
C3454 VDD.n2827 GND 0.001783f
C3455 VDD.n2828 GND 0.001783f
C3456 VDD.n2829 GND 9.69e-19
C3457 VDD.n2830 GND 0.001435f
C3458 VDD.n2831 GND 0.001783f
C3459 VDD.n2832 GND 0.001783f
C3460 VDD.n2833 GND 0.001435f
C3461 VDD.n2834 GND 0.001435f
C3462 VDD.n2835 GND 0.001783f
C3463 VDD.n2836 GND 0.001783f
C3464 VDD.n2837 GND 0.001435f
C3465 VDD.n2838 GND 0.001435f
C3466 VDD.n2839 GND 0.001783f
C3467 VDD.n2840 GND 0.001783f
C3468 VDD.n2841 GND 0.001435f
C3469 VDD.n2842 GND 0.001435f
C3470 VDD.n2843 GND 0.001783f
C3471 VDD.n2844 GND 0.001783f
C3472 VDD.n2845 GND 0.001435f
C3473 VDD.n2846 GND 0.001435f
C3474 VDD.n2847 GND 0.001783f
C3475 VDD.n2848 GND 0.001783f
C3476 VDD.n2849 GND 0.001435f
C3477 VDD.n2850 GND 0.001783f
C3478 VDD.n2851 GND 0.001783f
C3479 VDD.n2852 GND 0.001435f
C3480 VDD.n2853 GND 0.001783f
C3481 VDD.n2854 GND 0.001783f
C3482 VDD.n2855 GND 0.001783f
C3483 VDD.t8 GND 0.010031f
C3484 VDD.t9 GND 0.014304f
C3485 VDD.t6 GND 0.109243f
C3486 VDD.n2856 GND 0.024442f
C3487 VDD.n2857 GND 0.019628f
C3488 VDD.n2858 GND 0.002928f
C3489 VDD.n2859 GND 0.001783f
C3490 VDD.n2860 GND 0.001783f
C3491 VDD.n2861 GND 0.001198f
C3492 VDD.n2862 GND 0.001435f
C3493 VDD.n2863 GND 0.001783f
C3494 VDD.n2864 GND 0.001783f
C3495 VDD.n2865 GND 0.001435f
C3496 VDD.n2866 GND 0.001435f
C3497 VDD.n2867 GND 0.001783f
C3498 VDD.n2868 GND 0.001783f
C3499 VDD.n2869 GND 0.001435f
C3500 VDD.n2870 GND 0.001435f
C3501 VDD.n2871 GND 0.001783f
C3502 VDD.n2872 GND 0.001783f
C3503 VDD.n2873 GND 0.001435f
C3504 VDD.n2874 GND 0.001435f
C3505 VDD.n2875 GND 0.001783f
C3506 VDD.n2876 GND 0.001783f
C3507 VDD.n2877 GND 0.001435f
C3508 VDD.n2878 GND 0.001435f
C3509 VDD.n2879 GND 0.001783f
C3510 VDD.n2880 GND 0.001783f
C3511 VDD.n2881 GND 0.001435f
C3512 VDD.n2882 GND 0.001435f
C3513 VDD.n2883 GND 0.001783f
C3514 VDD.n2884 GND 0.001783f
C3515 VDD.n2885 GND 9.69e-19
C3516 VDD.n2886 GND 0.002928f
C3517 VDD.n2887 GND 0.001783f
C3518 VDD.n2888 GND 0.001783f
C3519 VDD.n2889 GND 0.001428f
C3520 VDD.n2890 GND 0.001435f
C3521 VDD.n2891 GND 0.001783f
C3522 VDD.n2892 GND 0.001783f
C3523 VDD.n2893 GND 0.001435f
C3524 VDD.n2894 GND 0.001435f
C3525 VDD.n2895 GND 0.001783f
C3526 VDD.n2896 GND 0.001783f
C3527 VDD.n2897 GND 0.001435f
C3528 VDD.n2898 GND 0.001435f
C3529 VDD.n2899 GND 0.001783f
C3530 VDD.n2900 GND 0.001783f
C3531 VDD.n2901 GND 0.001435f
C3532 VDD.n2902 GND 0.001783f
C3533 VDD.n2903 GND 0.001435f
C3534 VDD.n2904 GND 0.001435f
C3535 VDD.n2905 GND 0.001435f
C3536 VDD.n2906 GND 0.001191f
C3537 VDD.n2907 GND 0.004059f
C3538 VDD.n2909 GND 1.31281f
C3539 VDD.n2910 GND 0.004059f
C3540 VDD.n2911 GND 9.26e-19
C3541 VDD.n2912 GND 0.004059f
C3542 VDD.n2913 GND 0.003894f
C3543 VDD.n2914 GND 0.001783f
C3544 VDD.n2915 GND 0.001435f
C3545 VDD.n2916 GND 0.001783f
C3546 VDD.n2917 GND 0.158648f
C3547 VDD.n2918 GND 0.001783f
C3548 VDD.n2919 GND 0.001435f
C3549 VDD.n2920 GND 0.001783f
C3550 VDD.n2921 GND 0.001783f
C3551 VDD.n2922 GND 0.001783f
C3552 VDD.n2923 GND 0.001435f
C3553 VDD.n2924 GND 0.001783f
C3554 VDD.n2925 GND 0.130091f
C3555 VDD.n2926 GND 0.001783f
C3556 VDD.n2927 GND 0.001435f
C3557 VDD.n2928 GND 0.001783f
C3558 VDD.n2929 GND 0.001783f
C3559 VDD.n2930 GND 0.001783f
C3560 VDD.n2931 GND 0.001435f
C3561 VDD.n2932 GND 0.001783f
C3562 VDD.n2933 GND 0.158648f
C3563 VDD.n2934 GND 0.001783f
C3564 VDD.n2935 GND 0.001435f
C3565 VDD.n2936 GND 0.001783f
C3566 VDD.n2937 GND 0.001783f
C3567 VDD.n2938 GND 0.001783f
C3568 VDD.n2939 GND 0.001435f
C3569 VDD.n2940 GND 0.001783f
C3570 VDD.n2941 GND 0.158648f
C3571 VDD.n2942 GND 0.001783f
C3572 VDD.n2943 GND 0.001435f
C3573 VDD.n2944 GND 0.001783f
C3574 VDD.n2945 GND 0.001783f
C3575 VDD.n2946 GND 0.001783f
C3576 VDD.n2947 GND 0.001435f
C3577 VDD.n2948 GND 0.001783f
C3578 VDD.n2949 GND 0.158648f
C3579 VDD.n2950 GND 0.001783f
C3580 VDD.n2951 GND 0.001435f
C3581 VDD.n2952 GND 0.001783f
C3582 VDD.n2953 GND 0.001783f
C3583 VDD.n2954 GND 0.001783f
C3584 VDD.n2955 GND 0.001435f
C3585 VDD.n2956 GND 0.001783f
C3586 VDD.n2957 GND 0.158648f
C3587 VDD.n2958 GND 0.001783f
C3588 VDD.n2959 GND 0.001435f
C3589 VDD.n2960 GND 0.001783f
C3590 VDD.n2961 GND 0.001783f
C3591 VDD.n2962 GND 0.001783f
C3592 VDD.n2963 GND 0.001783f
C3593 VDD.n2964 GND 0.001783f
C3594 VDD.n2965 GND 0.001435f
C3595 VDD.n2966 GND 0.001783f
C3596 VDD.n2967 GND 0.158648f
C3597 VDD.n2968 GND 0.001783f
C3598 VDD.n2969 GND 0.001783f
C3599 VDD.n2970 GND 0.001783f
C3600 VDD.n2971 GND 0.001783f
C3601 VDD.n2972 GND 0.001435f
C3602 VDD.n2973 GND 0.001783f
C3603 VDD.n2974 GND 0.001783f
C3604 VDD.n2975 GND 0.001783f
C3605 VDD.n2976 GND 0.001783f
C3606 VDD.n2977 GND 0.158648f
C3607 VDD.n2978 GND 0.001783f
C3608 VDD.n2979 GND 0.001783f
C3609 VDD.n2980 GND 0.001783f
C3610 VDD.n2981 GND 0.001783f
C3611 VDD.n2982 GND 0.001783f
C3612 VDD.n2983 GND 0.001435f
C3613 VDD.n2984 GND 0.001783f
C3614 VDD.n2985 GND 0.001783f
C3615 VDD.n2986 GND 0.001783f
C3616 VDD.n2987 GND 0.001783f
C3617 VDD.n2988 GND 0.158648f
C3618 VDD.n2989 GND 0.001783f
C3619 VDD.n2990 GND 0.001783f
C3620 VDD.n2991 GND 0.001783f
C3621 VDD.n2992 GND 0.001783f
C3622 VDD.n2993 GND 0.001783f
C3623 VDD.n2994 GND 0.001191f
C3624 VDD.n2995 GND 0.003894f
C3625 VDD.n2996 GND 0.001783f
C3626 VDD.n2997 GND 0.003894f
C3627 VDD.n3031 GND 0.001783f
C3628 VDD.t93 GND 0.010031f
C3629 VDD.t92 GND 0.014304f
C3630 VDD.t91 GND 0.109243f
C3631 VDD.n3032 GND 0.024442f
C3632 VDD.n3033 GND 0.019628f
C3633 VDD.n3034 GND 0.002928f
C3634 VDD.n3035 GND 0.001783f
C3635 VDD.n3036 GND 0.001435f
C3636 VDD.n3037 GND 0.001783f
C3637 VDD.n3038 GND 0.001435f
C3638 VDD.n3039 GND 0.001783f
C3639 VDD.n3040 GND 0.001435f
C3640 VDD.n3041 GND 0.001783f
C3641 VDD.t87 GND 0.010031f
C3642 VDD.t86 GND 0.014304f
C3643 VDD.t85 GND 0.109243f
C3644 VDD.n3042 GND 0.024442f
C3645 VDD.n3043 GND 0.019628f
C3646 VDD.n3044 GND 0.001435f
C3647 VDD.n3045 GND 0.001783f
C3648 VDD.n3046 GND 0.001435f
C3649 VDD.n3047 GND 0.001783f
C3650 VDD.n3048 GND 0.001435f
C3651 VDD.n3049 GND 0.001783f
C3652 VDD.t33 GND 0.010031f
C3653 VDD.t32 GND 0.014304f
C3654 VDD.t31 GND 0.109243f
C3655 VDD.n3050 GND 0.024442f
C3656 VDD.n3051 GND 0.019628f
C3657 VDD.n3052 GND 0.001783f
C3658 VDD.n3053 GND 0.001435f
C3659 VDD.n3054 GND 0.001783f
C3660 VDD.n3055 GND 0.001435f
C3661 VDD.n3056 GND 0.001783f
C3662 VDD.n3057 GND 0.001435f
C3663 VDD.n3058 GND 0.001783f
C3664 VDD.t30 GND 0.010031f
C3665 VDD.t29 GND 0.014304f
C3666 VDD.t27 GND 0.109243f
C3667 VDD.n3059 GND 0.024442f
C3668 VDD.n3060 GND 0.019628f
C3669 VDD.n3061 GND 0.002928f
C3670 VDD.n3062 GND 0.001783f
C3671 VDD.n3063 GND 0.001435f
C3672 VDD.n3064 GND 0.001783f
C3673 VDD.n3065 GND 0.001435f
C3674 VDD.n3066 GND 0.001783f
C3675 VDD.n3067 GND 0.001435f
C3676 VDD.n3068 GND 0.001783f
C3677 VDD.t36 GND 0.010031f
C3678 VDD.t35 GND 0.014304f
C3679 VDD.t34 GND 0.109243f
C3680 VDD.n3069 GND 0.024442f
C3681 VDD.n3070 GND 0.019628f
C3682 VDD.n3071 GND 0.001435f
C3683 VDD.n3072 GND 0.001783f
C3684 VDD.n3073 GND 0.001435f
C3685 VDD.n3074 GND 0.001783f
C3686 VDD.n3075 GND 0.001435f
C3687 VDD.n3076 GND 0.003894f
C3688 VDD.n3077 GND 0.004059f
C3689 VDD.n3078 GND 0.001191f
C3690 VDD.n3079 GND 0.004059f
C3691 VDD.n3080 GND 0.001783f
C3692 VDD.n3081 GND 0.001783f
C3693 VDD.n3082 GND 0.001783f
C3694 VDD.n3083 GND 0.001783f
C3695 VDD.n3084 GND 0.001435f
C3696 VDD.n3085 GND 0.001435f
C3697 VDD.n3086 GND 0.001783f
C3698 VDD.n3087 GND 0.001783f
C3699 VDD.n3088 GND 0.001435f
C3700 VDD.n3089 GND 0.001783f
C3701 VDD.n3090 GND 0.001783f
C3702 VDD.n3091 GND 0.001783f
C3703 VDD.n3092 GND 0.001783f
C3704 VDD.n3093 GND 0.001783f
C3705 VDD.n3094 GND 0.001435f
C3706 VDD.n3095 GND 0.001435f
C3707 VDD.n3096 GND 0.001783f
C3708 VDD.n3097 GND 0.001783f
C3709 VDD.n3098 GND 0.001435f
C3710 VDD.n3099 GND 0.001783f
C3711 VDD.n3100 GND 0.001783f
C3712 VDD.n3101 GND 0.001783f
C3713 VDD.n3102 GND 0.001783f
C3714 VDD.n3103 GND 0.001783f
C3715 VDD.n3104 GND 0.001428f
C3716 VDD.n3105 GND 0.002928f
C3717 VDD.n3106 GND 0.001783f
C3718 VDD.n3107 GND 0.001783f
C3719 VDD.n3108 GND 9.69e-19
C3720 VDD.n3109 GND 0.001783f
C3721 VDD.n3110 GND 0.001783f
C3722 VDD.n3111 GND 0.001783f
C3723 VDD.n3112 GND 0.001783f
C3724 VDD.n3113 GND 0.001783f
C3725 VDD.n3114 GND 0.001435f
C3726 VDD.n3115 GND 0.001435f
C3727 VDD.n3116 GND 0.001783f
C3728 VDD.n3117 GND 0.001783f
C3729 VDD.n3118 GND 0.001435f
C3730 VDD.n3119 GND 0.001783f
C3731 VDD.n3120 GND 0.001783f
C3732 VDD.n3121 GND 0.001783f
C3733 VDD.n3122 GND 0.001783f
C3734 VDD.n3123 GND 0.001783f
C3735 VDD.n3124 GND 0.001435f
C3736 VDD.n3125 GND 0.001435f
C3737 VDD.n3126 GND 0.001783f
C3738 VDD.n3127 GND 0.001783f
C3739 VDD.n3128 GND 0.001435f
C3740 VDD.n3129 GND 0.001783f
C3741 VDD.n3130 GND 0.001783f
C3742 VDD.n3131 GND 0.001783f
C3743 VDD.n3132 GND 0.001783f
C3744 VDD.n3133 GND 0.001783f
C3745 VDD.n3134 GND 0.001435f
C3746 VDD.n3135 GND 0.001435f
C3747 VDD.n3136 GND 0.001783f
C3748 VDD.n3137 GND 0.001783f
C3749 VDD.n3138 GND 0.001198f
C3750 VDD.n3139 GND 0.001783f
C3751 VDD.n3140 GND 0.001783f
C3752 VDD.n3141 GND 0.001783f
C3753 VDD.n3142 GND 0.001783f
C3754 VDD.n3143 GND 0.001783f
C3755 VDD.n3144 GND 0.001198f
C3756 VDD.n3145 GND 0.001435f
C3757 VDD.n3146 GND 0.001783f
C3758 VDD.n3147 GND 0.001783f
C3759 VDD.n3148 GND 0.001435f
C3760 VDD.n3149 GND 0.001783f
C3761 VDD.n3150 GND 0.001783f
C3762 VDD.n3151 GND 0.001783f
C3763 VDD.n3152 GND 0.001783f
C3764 VDD.n3153 GND 0.001783f
C3765 VDD.n3154 GND 0.001435f
C3766 VDD.n3155 GND 0.001435f
C3767 VDD.n3156 GND 0.001783f
C3768 VDD.n3157 GND 0.001783f
C3769 VDD.n3158 GND 0.001435f
C3770 VDD.n3159 GND 0.001783f
C3771 VDD.n3160 GND 0.001783f
C3772 VDD.n3161 GND 0.001783f
C3773 VDD.n3162 GND 0.001783f
C3774 VDD.n3163 GND 0.001783f
C3775 VDD.n3164 GND 0.001435f
C3776 VDD.n3165 GND 0.001435f
C3777 VDD.n3166 GND 0.001783f
C3778 VDD.n3167 GND 0.001783f
C3779 VDD.n3168 GND 0.001435f
C3780 VDD.n3169 GND 0.001783f
C3781 VDD.n3170 GND 0.001783f
C3782 VDD.n3171 GND 0.001783f
C3783 VDD.n3172 GND 0.001783f
C3784 VDD.n3173 GND 0.001783f
C3785 VDD.n3174 GND 9.69e-19
C3786 VDD.n3175 GND 0.002928f
C3787 VDD.n3176 GND 0.001783f
C3788 VDD.n3177 GND 0.001783f
C3789 VDD.n3178 GND 0.001428f
C3790 VDD.n3179 GND 0.001783f
C3791 VDD.n3180 GND 0.001783f
C3792 VDD.n3181 GND 0.001435f
C3793 VDD.n3182 GND 0.001783f
C3794 VDD.n3183 GND 0.001783f
C3795 VDD.n3184 GND 0.001783f
C3796 VDD.n3185 GND 0.001435f
C3797 VDD.n3186 GND 0.001783f
C3798 VDD.n3187 GND 0.001783f
C3799 VDD.n3188 GND 0.001435f
C3800 VDD.n3189 GND 0.001783f
C3801 VDD.n3190 GND 0.001783f
C3802 VDD.n3191 GND 0.001435f
C3803 VDD.n3192 GND 0.001783f
C3804 VDD.n3193 GND 0.001783f
C3805 VDD.n3194 GND 0.001783f
C3806 VDD.n3195 GND 0.001435f
C3807 VDD.n3196 GND 0.001783f
C3808 VDD.n3197 GND 0.001783f
C3809 VDD.n3198 GND 0.001435f
C3810 VDD.n3199 GND 0.001783f
C3811 VDD.n3200 GND 0.001783f
C3812 VDD.n3201 GND 0.001435f
C3813 VDD.n3202 GND 0.001783f
C3814 VDD.n3203 GND 0.001783f
C3815 VDD.n3204 GND 0.001783f
C3816 VDD.n3205 GND 0.001435f
C3817 VDD.n3206 GND 0.001783f
C3818 VDD.n3207 GND 0.001783f
C3819 VDD.n3208 GND 7.39e-19
C3820 VDD.n3209 GND 0.00221f
C3821 VDD.n3210 GND 0.001783f
C3822 VDD.n3211 GND 0.001783f
C3823 VDD.n3212 GND 9.4e-19
C3824 VDD.n3213 GND 0.001783f
C3825 VDD.n3214 GND 0.001783f
C3826 VDD.n3215 GND 0.001783f
C3827 VDD.n3216 GND 0.001435f
C3828 VDD.n3217 GND 0.001783f
C3829 VDD.n3218 GND 0.001783f
C3830 VDD.n3219 GND 0.001435f
C3831 VDD.n3220 GND 0.001783f
C3832 VDD.n3221 GND 0.001783f
C3833 VDD.n3222 GND 0.001435f
C3834 VDD.n3223 GND 0.001783f
C3835 VDD.n3224 GND 0.001783f
C3836 VDD.n3225 GND 0.001783f
C3837 VDD.n3226 GND 0.001435f
C3838 VDD.n3227 GND 0.001783f
C3839 VDD.n3228 GND 0.001783f
C3840 VDD.n3229 GND 0.001435f
C3841 VDD.n3230 GND 0.001783f
C3842 VDD.n3231 GND 0.001783f
C3843 VDD.n3232 GND 0.001435f
C3844 VDD.n3233 GND 0.001783f
C3845 VDD.n3234 GND 0.001783f
C3846 VDD.n3235 GND 0.001783f
C3847 VDD.n3236 GND 0.001435f
C3848 VDD.n3237 GND 0.001783f
C3849 VDD.n3238 GND 0.001783f
C3850 VDD.n3239 GND 0.001435f
C3851 VDD.n3240 GND 0.001783f
C3852 VDD.n3241 GND 0.001227f
C3853 VDD.n3242 GND 0.001783f
C3854 VDD.n3243 GND 0.001783f
C3855 VDD.n3244 GND 0.001783f
C3856 VDD.n3245 GND 0.001435f
C3857 VDD.n3246 GND 0.001783f
C3858 VDD.n3247 GND 0.001435f
C3859 VDD.n3248 GND 0.001783f
C3860 VDD.n3249 GND 0.001783f
C3861 VDD.n3250 GND 0.001435f
C3862 VDD.n3251 GND 0.001435f
C3863 VDD.n3252 GND 0.001783f
C3864 VDD.n3253 GND 0.001783f
C3865 VDD.n3254 GND 0.001783f
C3866 VDD.n3255 GND 0.001783f
C3867 VDD.n3256 GND 0.001435f
C3868 VDD.n3257 GND 0.001435f
C3869 VDD.n3258 GND 0.001435f
C3870 VDD.n3259 GND 0.001783f
C3871 VDD.n3260 GND 0.001783f
C3872 VDD.n3261 GND 0.001783f
C3873 VDD.n3262 GND 0.001783f
C3874 VDD.n3263 GND 0.001435f
C3875 VDD.n3264 GND 0.001435f
C3876 VDD.n3265 GND 0.001191f
C3877 VDD.n3266 GND 0.003894f
C3878 VDD.n3267 GND 0.004059f
C3879 VDD.n3268 GND 9.26e-19
C3880 VDD.n3269 GND 0.004059f
C3881 VDD.n3271 GND 0.372029f
C3882 VDD.n3272 GND 0.22766f
C3883 VDD.n3273 GND 0.158648f
C3884 VDD.n3274 GND 0.001783f
C3885 VDD.n3275 GND 0.001435f
C3886 VDD.n3276 GND 0.001435f
C3887 VDD.n3277 GND 0.001435f
C3888 VDD.n3278 GND 0.001783f
C3889 VDD.n3279 GND 0.130091f
C3890 VDD.t28 GND 0.079324f
C3891 VDD.n3280 GND 0.107881f
C3892 VDD.n3281 GND 0.158648f
C3893 VDD.n3282 GND 0.001783f
C3894 VDD.n3283 GND 0.001435f
C3895 VDD.n3284 GND 0.001435f
C3896 VDD.n3285 GND 0.001435f
C3897 VDD.n3286 GND 0.001783f
C3898 VDD.n3287 GND 0.158648f
C3899 VDD.n3288 GND 0.158648f
C3900 VDD.n3289 GND 0.158648f
C3901 VDD.n3290 GND 0.001783f
C3902 VDD.n3291 GND 0.001435f
C3903 VDD.n3292 GND 0.001435f
C3904 VDD.n3293 GND 0.001435f
C3905 VDD.n3294 GND 0.001783f
C3906 VDD.n3295 GND 0.158648f
C3907 VDD.n3296 GND 0.001783f
C3908 VDD.n3297 GND 0.001435f
C3909 VDD.n3298 GND 0.001435f
C3910 VDD.n3299 GND 0.001435f
C3911 VDD.n3300 GND 0.001783f
C3912 VDD.t126 GND 0.158648f
C3913 VDD.n3301 GND 0.001783f
C3914 VDD.n3302 GND 0.001435f
C3915 VDD.n3303 GND 0.003335f
C3916 VDD.n3304 GND 0.001005f
C3917 VDD.n3305 GND 9.08e-19
C3918 VDD.n3306 GND 4.88e-19
C3919 VDD.n3307 GND 0.001153f
C3920 VDD.n3308 GND 5.17e-19
C3921 VDD.n3309 GND 0.003542f
C3922 VDD.t132 GND 0.002562f
C3923 VDD.n3310 GND 8.65e-19
C3924 VDD.n3311 GND 7.25e-19
C3925 VDD.n3312 GND 4.88e-19
C3926 VDD.n3313 GND 0.012395f
C3927 VDD.n3314 GND 9.08e-19
C3928 VDD.n3315 GND 4.88e-19
C3929 VDD.n3316 GND 5.17e-19
C3930 VDD.n3317 GND 0.001153f
C3931 VDD.n3318 GND 0.002818f
C3932 VDD.n3319 GND 5.17e-19
C3933 VDD.n3320 GND 4.88e-19
C3934 VDD.n3321 GND 0.002285f
C3935 VDD.n3322 GND 0.005604f
C3936 VDD.n3323 GND 0.001005f
C3937 VDD.n3324 GND 9.08e-19
C3938 VDD.n3325 GND 4.88e-19
C3939 VDD.n3326 GND 0.001153f
C3940 VDD.n3327 GND 5.17e-19
C3941 VDD.n3328 GND 0.003542f
C3942 VDD.t127 GND 0.002562f
C3943 VDD.n3329 GND 8.65e-19
C3944 VDD.n3330 GND 7.25e-19
C3945 VDD.n3331 GND 4.88e-19
C3946 VDD.n3332 GND 0.012395f
C3947 VDD.n3333 GND 9.08e-19
C3948 VDD.n3334 GND 4.88e-19
C3949 VDD.n3335 GND 5.17e-19
C3950 VDD.n3336 GND 0.001153f
C3951 VDD.n3337 GND 0.002818f
C3952 VDD.n3338 GND 5.17e-19
C3953 VDD.n3339 GND 4.88e-19
C3954 VDD.n3340 GND 0.002285f
C3955 VDD.n3341 GND 0.004299f
C3956 VDD.n3342 GND 0.097922f
C3957 VDD.n3343 GND 0.001005f
C3958 VDD.n3344 GND 9.08e-19
C3959 VDD.n3345 GND 4.88e-19
C3960 VDD.n3346 GND 0.001153f
C3961 VDD.n3347 GND 5.17e-19
C3962 VDD.n3348 GND 0.003542f
C3963 VDD.t138 GND 0.002562f
C3964 VDD.n3349 GND 8.65e-19
C3965 VDD.n3350 GND 7.25e-19
C3966 VDD.n3351 GND 4.88e-19
C3967 VDD.n3352 GND 0.012395f
C3968 VDD.n3353 GND 9.08e-19
C3969 VDD.n3354 GND 4.88e-19
C3970 VDD.n3355 GND 5.17e-19
C3971 VDD.n3356 GND 0.001153f
C3972 VDD.n3357 GND 0.002818f
C3973 VDD.n3358 GND 5.17e-19
C3974 VDD.n3359 GND 4.88e-19
C3975 VDD.n3360 GND 0.002285f
C3976 VDD.n3361 GND 0.004299f
C3977 VDD.n3362 GND 0.057698f
C3978 VDD.n3363 GND 0.001005f
C3979 VDD.n3364 GND 9.08e-19
C3980 VDD.n3365 GND 4.88e-19
C3981 VDD.n3366 GND 0.001153f
C3982 VDD.n3367 GND 5.17e-19
C3983 VDD.n3368 GND 0.003542f
C3984 VDD.t134 GND 0.002562f
C3985 VDD.n3369 GND 8.65e-19
C3986 VDD.n3370 GND 7.25e-19
C3987 VDD.n3371 GND 4.88e-19
C3988 VDD.n3372 GND 0.012395f
C3989 VDD.n3373 GND 9.08e-19
C3990 VDD.n3374 GND 4.88e-19
C3991 VDD.n3375 GND 5.17e-19
C3992 VDD.n3376 GND 0.001153f
C3993 VDD.n3377 GND 0.002818f
C3994 VDD.n3378 GND 5.17e-19
C3995 VDD.n3379 GND 4.88e-19
C3996 VDD.n3380 GND 0.002285f
C3997 VDD.n3381 GND 0.004299f
C3998 VDD.n3382 GND 0.057698f
C3999 VDD.n3383 GND 0.001005f
C4000 VDD.n3384 GND 9.08e-19
C4001 VDD.n3385 GND 4.88e-19
C4002 VDD.n3386 GND 0.001153f
C4003 VDD.n3387 GND 5.17e-19
C4004 VDD.n3388 GND 0.003542f
C4005 VDD.t137 GND 0.002562f
C4006 VDD.n3389 GND 8.65e-19
C4007 VDD.n3390 GND 7.25e-19
C4008 VDD.n3391 GND 4.88e-19
C4009 VDD.n3392 GND 0.012395f
C4010 VDD.n3393 GND 9.08e-19
C4011 VDD.n3394 GND 4.88e-19
C4012 VDD.n3395 GND 5.17e-19
C4013 VDD.n3396 GND 0.001153f
C4014 VDD.n3397 GND 0.002818f
C4015 VDD.n3398 GND 5.17e-19
C4016 VDD.n3399 GND 4.88e-19
C4017 VDD.n3400 GND 0.002285f
C4018 VDD.n3401 GND 0.004299f
C4019 VDD.n3402 GND 0.054622f
C4020 VDD.n3403 GND 0.40987f
C4021 VOUT.n0 GND 0.005628f
C4022 VOUT.n1 GND 0.005082f
C4023 VOUT.n2 GND 0.002731f
C4024 VOUT.n3 GND 0.006455f
C4025 VOUT.n4 GND 0.002892f
C4026 VOUT.n5 GND 0.019824f
C4027 VOUT.t37 GND 0.014336f
C4028 VOUT.n6 GND 0.004841f
C4029 VOUT.n7 GND 0.00406f
C4030 VOUT.n8 GND 0.002731f
C4031 VOUT.n9 GND 0.069373f
C4032 VOUT.n10 GND 0.005082f
C4033 VOUT.n11 GND 0.002731f
C4034 VOUT.n12 GND 0.002892f
C4035 VOUT.n13 GND 0.006455f
C4036 VOUT.n14 GND 0.015774f
C4037 VOUT.n15 GND 0.002892f
C4038 VOUT.n16 GND 0.002731f
C4039 VOUT.n17 GND 0.012788f
C4040 VOUT.n18 GND 0.032586f
C4041 VOUT.n19 GND 0.005628f
C4042 VOUT.n20 GND 0.005082f
C4043 VOUT.n21 GND 0.002731f
C4044 VOUT.n22 GND 0.006455f
C4045 VOUT.n23 GND 0.002892f
C4046 VOUT.n24 GND 0.019824f
C4047 VOUT.t35 GND 0.014336f
C4048 VOUT.n25 GND 0.004841f
C4049 VOUT.n26 GND 0.00406f
C4050 VOUT.n27 GND 0.002731f
C4051 VOUT.n28 GND 0.069373f
C4052 VOUT.n29 GND 0.005082f
C4053 VOUT.n30 GND 0.002731f
C4054 VOUT.n31 GND 0.002892f
C4055 VOUT.n32 GND 0.006455f
C4056 VOUT.n33 GND 0.015774f
C4057 VOUT.n34 GND 0.002892f
C4058 VOUT.n35 GND 0.002731f
C4059 VOUT.n36 GND 0.012788f
C4060 VOUT.n37 GND 0.027192f
C4061 VOUT.n38 GND 0.634581f
C4062 VOUT.n39 GND 0.005628f
C4063 VOUT.n40 GND 0.005082f
C4064 VOUT.n41 GND 0.002731f
C4065 VOUT.n42 GND 0.006455f
C4066 VOUT.n43 GND 0.002892f
C4067 VOUT.n44 GND 0.019824f
C4068 VOUT.t36 GND 0.014336f
C4069 VOUT.n45 GND 0.004841f
C4070 VOUT.n46 GND 0.00406f
C4071 VOUT.n47 GND 0.002731f
C4072 VOUT.n48 GND 0.069373f
C4073 VOUT.n49 GND 0.005082f
C4074 VOUT.n50 GND 0.002731f
C4075 VOUT.n51 GND 0.002892f
C4076 VOUT.n52 GND 0.006455f
C4077 VOUT.n53 GND 0.015774f
C4078 VOUT.n54 GND 0.002892f
C4079 VOUT.n55 GND 0.002731f
C4080 VOUT.n56 GND 0.012788f
C4081 VOUT.n57 GND 0.027192f
C4082 VOUT.n58 GND 0.365232f
C4083 VOUT.n59 GND 0.005628f
C4084 VOUT.n60 GND 0.005082f
C4085 VOUT.n61 GND 0.002731f
C4086 VOUT.n62 GND 0.006455f
C4087 VOUT.n63 GND 0.002892f
C4088 VOUT.n64 GND 0.019824f
C4089 VOUT.t39 GND 0.014336f
C4090 VOUT.n65 GND 0.004841f
C4091 VOUT.n66 GND 0.00406f
C4092 VOUT.n67 GND 0.002731f
C4093 VOUT.n68 GND 0.069373f
C4094 VOUT.n69 GND 0.005082f
C4095 VOUT.n70 GND 0.002731f
C4096 VOUT.n71 GND 0.002892f
C4097 VOUT.n72 GND 0.006455f
C4098 VOUT.n73 GND 0.015774f
C4099 VOUT.n74 GND 0.002892f
C4100 VOUT.n75 GND 0.002731f
C4101 VOUT.n76 GND 0.012788f
C4102 VOUT.n77 GND 0.027192f
C4103 VOUT.n78 GND 0.365232f
C4104 VOUT.n79 GND 0.005628f
C4105 VOUT.n80 GND 0.005082f
C4106 VOUT.n81 GND 0.002731f
C4107 VOUT.n82 GND 0.006455f
C4108 VOUT.n83 GND 0.002892f
C4109 VOUT.n84 GND 0.019824f
C4110 VOUT.t33 GND 0.014336f
C4111 VOUT.n85 GND 0.004841f
C4112 VOUT.n86 GND 0.00406f
C4113 VOUT.n87 GND 0.002731f
C4114 VOUT.n88 GND 0.069373f
C4115 VOUT.n89 GND 0.005082f
C4116 VOUT.n90 GND 0.002731f
C4117 VOUT.n91 GND 0.002892f
C4118 VOUT.n92 GND 0.006455f
C4119 VOUT.n93 GND 0.015774f
C4120 VOUT.n94 GND 0.002892f
C4121 VOUT.n95 GND 0.002731f
C4122 VOUT.n96 GND 0.012788f
C4123 VOUT.n97 GND 0.027192f
C4124 VOUT.n98 GND 0.495718f
C4125 VOUT.n99 GND 7.14075f
C4126 VOUT.n100 GND 1.27609f
C4127 VOUT.n101 GND 0.880022f
C4128 VOUT.n102 GND 0.880022f
C4129 VOUT.t42 GND 2.87235f
C4130 VOUT.t43 GND 2.7501f
C4131 VOUT.t46 GND 2.7501f
C4132 VOUT.t47 GND 2.88687f
C4133 VOUT.n103 GND 2.24058f
C4134 VOUT.n104 GND 1.14793f
C4135 VOUT.n105 GND 0.880022f
C4136 VOUT.n106 GND 1.01131f
C4137 VOUT.n107 GND 1.05329f
C4138 VOUT.n108 GND 0.880022f
C4139 VOUT.n109 GND 1.10735f
C4140 VOUT.n110 GND 2.67324f
C4141 VOUT.t44 GND 2.87235f
C4142 VOUT.n111 GND 2.67324f
C4143 VOUT.n112 GND 1.10735f
C4144 VOUT.t45 GND 2.7501f
C4145 VOUT.n113 GND 1.05329f
C4146 VOUT.n114 GND 1.01131f
C4147 VOUT.t40 GND 2.7501f
C4148 VOUT.n115 GND 1.05329f
C4149 VOUT.n116 GND 1.01131f
C4150 VOUT.t41 GND 2.7501f
C4151 VOUT.n117 GND 2.2274f
C4152 VOUT.n118 GND 1.49332f
C4153 VOUT.n119 GND 0.005628f
C4154 VOUT.n120 GND 0.005082f
C4155 VOUT.n121 GND 0.002731f
C4156 VOUT.n122 GND 0.006455f
C4157 VOUT.n123 GND 0.002892f
C4158 VOUT.n124 GND 0.019824f
C4159 VOUT.t34 GND 0.014336f
C4160 VOUT.n125 GND 0.004841f
C4161 VOUT.n126 GND 0.00406f
C4162 VOUT.n127 GND 0.002731f
C4163 VOUT.n128 GND 0.069373f
C4164 VOUT.n129 GND 0.005082f
C4165 VOUT.n130 GND 0.002731f
C4166 VOUT.n131 GND 0.002892f
C4167 VOUT.n132 GND 0.006455f
C4168 VOUT.n133 GND 0.015774f
C4169 VOUT.n134 GND 0.002892f
C4170 VOUT.n135 GND 0.002731f
C4171 VOUT.n136 GND 0.012788f
C4172 VOUT.n137 GND 0.033086f
C4173 VOUT.n138 GND 0.005628f
C4174 VOUT.n139 GND 0.005082f
C4175 VOUT.n140 GND 0.002731f
C4176 VOUT.n141 GND 0.006455f
C4177 VOUT.n142 GND 0.002892f
C4178 VOUT.n143 GND 0.019824f
C4179 VOUT.t38 GND 0.014336f
C4180 VOUT.n144 GND 0.004841f
C4181 VOUT.n145 GND 0.00406f
C4182 VOUT.n146 GND 0.002731f
C4183 VOUT.n147 GND 0.069373f
C4184 VOUT.n148 GND 0.005082f
C4185 VOUT.n149 GND 0.002731f
C4186 VOUT.n150 GND 0.002892f
C4187 VOUT.n151 GND 0.006455f
C4188 VOUT.n152 GND 0.015774f
C4189 VOUT.n153 GND 0.002892f
C4190 VOUT.n154 GND 0.002731f
C4191 VOUT.n155 GND 0.012788f
C4192 VOUT.n156 GND 0.027758f
C4193 VOUT.n157 GND 0.633516f
C4194 VOUT.n158 GND 0.005628f
C4195 VOUT.n159 GND 0.005082f
C4196 VOUT.n160 GND 0.002731f
C4197 VOUT.n161 GND 0.006455f
C4198 VOUT.n162 GND 0.002892f
C4199 VOUT.n163 GND 0.019824f
C4200 VOUT.t32 GND 0.014336f
C4201 VOUT.n164 GND 0.004841f
C4202 VOUT.n165 GND 0.00406f
C4203 VOUT.n166 GND 0.002731f
C4204 VOUT.n167 GND 0.069373f
C4205 VOUT.n168 GND 0.005082f
C4206 VOUT.n169 GND 0.002731f
C4207 VOUT.n170 GND 0.002892f
C4208 VOUT.n171 GND 0.006455f
C4209 VOUT.n172 GND 0.015774f
C4210 VOUT.n173 GND 0.002892f
C4211 VOUT.n174 GND 0.002731f
C4212 VOUT.n175 GND 0.012788f
C4213 VOUT.n176 GND 0.027758f
C4214 VOUT.n177 GND 0.364667f
C4215 VOUT.n178 GND 0.005628f
C4216 VOUT.n179 GND 0.005082f
C4217 VOUT.n180 GND 0.002731f
C4218 VOUT.n181 GND 0.006455f
C4219 VOUT.n182 GND 0.002892f
C4220 VOUT.n183 GND 0.019824f
C4221 VOUT.t30 GND 0.014336f
C4222 VOUT.n184 GND 0.004841f
C4223 VOUT.n185 GND 0.00406f
C4224 VOUT.n186 GND 0.002731f
C4225 VOUT.n187 GND 0.069373f
C4226 VOUT.n188 GND 0.005082f
C4227 VOUT.n189 GND 0.002731f
C4228 VOUT.n190 GND 0.002892f
C4229 VOUT.n191 GND 0.006455f
C4230 VOUT.n192 GND 0.015774f
C4231 VOUT.n193 GND 0.002892f
C4232 VOUT.n194 GND 0.002731f
C4233 VOUT.n195 GND 0.012788f
C4234 VOUT.n196 GND 0.027758f
C4235 VOUT.n197 GND 0.364667f
C4236 VOUT.n198 GND 0.005628f
C4237 VOUT.n199 GND 0.005082f
C4238 VOUT.n200 GND 0.002731f
C4239 VOUT.n201 GND 0.006455f
C4240 VOUT.n202 GND 0.002892f
C4241 VOUT.n203 GND 0.019824f
C4242 VOUT.t31 GND 0.014336f
C4243 VOUT.n204 GND 0.004841f
C4244 VOUT.n205 GND 0.00406f
C4245 VOUT.n206 GND 0.002731f
C4246 VOUT.n207 GND 0.069373f
C4247 VOUT.n208 GND 0.005082f
C4248 VOUT.n209 GND 0.002731f
C4249 VOUT.n210 GND 0.002892f
C4250 VOUT.n211 GND 0.006455f
C4251 VOUT.n212 GND 0.015774f
C4252 VOUT.n213 GND 0.002892f
C4253 VOUT.n214 GND 0.002731f
C4254 VOUT.n215 GND 0.012788f
C4255 VOUT.n216 GND 0.027758f
C4256 VOUT.n217 GND 0.495152f
C4257 VOUT.n218 GND 9.24917f
C4258 VOUT.n219 GND 0.007521f
C4259 VOUT.n220 GND 0.044654f
C4260 VOUT.n221 GND 0.002731f
C4261 VOUT.t19 GND 0.01182f
C4262 VOUT.n222 GND 0.01922f
C4263 VOUT.n223 GND 0.00442f
C4264 VOUT.n224 GND 0.004841f
C4265 VOUT.n225 GND 0.014641f
C4266 VOUT.n226 GND 0.002892f
C4267 VOUT.n227 GND 0.002731f
C4268 VOUT.n228 GND 0.0114f
C4269 VOUT.n229 GND 0.016896f
C4270 VOUT.t0 GND 0.010883f
C4271 VOUT.t3 GND 0.010883f
C4272 VOUT.n230 GND 0.0837f
C4273 VOUT.n231 GND 0.28196f
C4274 VOUT.t11 GND 0.010883f
C4275 VOUT.t21 GND 0.010883f
C4276 VOUT.n232 GND 0.0837f
C4277 VOUT.n233 GND 0.262721f
C4278 VOUT.n234 GND 0.007521f
C4279 VOUT.n235 GND 0.044654f
C4280 VOUT.n236 GND 0.002731f
C4281 VOUT.t18 GND 0.01182f
C4282 VOUT.n237 GND 0.01922f
C4283 VOUT.n238 GND 0.00442f
C4284 VOUT.n239 GND 0.004841f
C4285 VOUT.n240 GND 0.014641f
C4286 VOUT.n241 GND 0.002892f
C4287 VOUT.n242 GND 0.002731f
C4288 VOUT.n243 GND 0.0114f
C4289 VOUT.n244 GND 0.016896f
C4290 VOUT.t5 GND 0.010883f
C4291 VOUT.t23 GND 0.010883f
C4292 VOUT.n245 GND 0.0837f
C4293 VOUT.n246 GND 0.28196f
C4294 VOUT.t10 GND 0.010883f
C4295 VOUT.t27 GND 0.010883f
C4296 VOUT.n247 GND 0.0837f
C4297 VOUT.n248 GND 0.245196f
C4298 VOUT.n249 GND 0.252216f
C4299 VOUT.n250 GND 0.007521f
C4300 VOUT.n251 GND 0.044654f
C4301 VOUT.n252 GND 0.002731f
C4302 VOUT.t2 GND 0.01182f
C4303 VOUT.n253 GND 0.01922f
C4304 VOUT.n254 GND 0.00442f
C4305 VOUT.n255 GND 0.004841f
C4306 VOUT.n256 GND 0.014641f
C4307 VOUT.n257 GND 0.002892f
C4308 VOUT.n258 GND 0.002731f
C4309 VOUT.n259 GND 0.0114f
C4310 VOUT.n260 GND 0.016896f
C4311 VOUT.t14 GND 0.010883f
C4312 VOUT.t17 GND 0.010883f
C4313 VOUT.n261 GND 0.0837f
C4314 VOUT.n262 GND 0.28196f
C4315 VOUT.t26 GND 0.010883f
C4316 VOUT.t8 GND 0.010883f
C4317 VOUT.n263 GND 0.0837f
C4318 VOUT.n264 GND 0.245196f
C4319 VOUT.n265 GND 0.443045f
C4320 VOUT.n266 GND 9.06613f
C4321 VOUT.t4 GND 0.010883f
C4322 VOUT.t1 GND 0.010883f
C4323 VOUT.n267 GND 0.085908f
C4324 VOUT.t22 GND 0.010883f
C4325 VOUT.t13 GND 0.010883f
C4326 VOUT.n268 GND 0.0837f
C4327 VOUT.n269 GND 0.386366f
C4328 VOUT.n270 GND 0.007521f
C4329 VOUT.n271 GND 0.044654f
C4330 VOUT.n272 GND 0.002731f
C4331 VOUT.t25 GND 0.01182f
C4332 VOUT.n273 GND 0.01922f
C4333 VOUT.n274 GND 0.00442f
C4334 VOUT.n275 GND 0.004841f
C4335 VOUT.n276 GND 0.014641f
C4336 VOUT.n277 GND 0.002892f
C4337 VOUT.n278 GND 0.002731f
C4338 VOUT.n279 GND 0.0114f
C4339 VOUT.n280 GND 0.015284f
C4340 VOUT.n281 GND 0.167971f
C4341 VOUT.t28 GND 0.010883f
C4342 VOUT.t6 GND 0.010883f
C4343 VOUT.n282 GND 0.085908f
C4344 VOUT.t29 GND 0.010883f
C4345 VOUT.t12 GND 0.010883f
C4346 VOUT.n283 GND 0.0837f
C4347 VOUT.n284 GND 0.386366f
C4348 VOUT.n285 GND 0.007521f
C4349 VOUT.n286 GND 0.044654f
C4350 VOUT.n287 GND 0.002731f
C4351 VOUT.t20 GND 0.01182f
C4352 VOUT.n288 GND 0.01922f
C4353 VOUT.n289 GND 0.00442f
C4354 VOUT.n290 GND 0.004841f
C4355 VOUT.n291 GND 0.014641f
C4356 VOUT.n292 GND 0.002892f
C4357 VOUT.n293 GND 0.002731f
C4358 VOUT.n294 GND 0.0114f
C4359 VOUT.n295 GND 0.015284f
C4360 VOUT.n296 GND 0.150865f
C4361 VOUT.n297 GND 0.231292f
C4362 VOUT.t16 GND 0.010883f
C4363 VOUT.t15 GND 0.010883f
C4364 VOUT.n298 GND 0.085908f
C4365 VOUT.t7 GND 0.010883f
C4366 VOUT.t24 GND 0.010883f
C4367 VOUT.n299 GND 0.0837f
C4368 VOUT.n300 GND 0.386366f
C4369 VOUT.n301 GND 0.007521f
C4370 VOUT.n302 GND 0.044654f
C4371 VOUT.n303 GND 0.002731f
C4372 VOUT.t9 GND 0.01182f
C4373 VOUT.n304 GND 0.01922f
C4374 VOUT.n305 GND 0.00442f
C4375 VOUT.n306 GND 0.004841f
C4376 VOUT.n307 GND 0.014641f
C4377 VOUT.n308 GND 0.002892f
C4378 VOUT.n309 GND 0.002731f
C4379 VOUT.n310 GND 0.0114f
C4380 VOUT.n311 GND 0.015284f
C4381 VOUT.n312 GND 0.150865f
C4382 VOUT.n313 GND 0.432373f
C4383 VOUT.n314 GND 6.48825f
C4384 VOUT.n315 GND 4.74034f
C4385 CS_BIAS.n0 GND 0.008903f
C4386 CS_BIAS.t30 GND 0.106594f
C4387 CS_BIAS.n1 GND 0.008917f
C4388 CS_BIAS.n2 GND 0.006753f
C4389 CS_BIAS.t49 GND 0.106594f
C4390 CS_BIAS.n3 GND 0.046728f
C4391 CS_BIAS.n4 GND 0.006753f
C4392 CS_BIAS.n5 GND 0.013528f
C4393 CS_BIAS.n6 GND 0.008903f
C4394 CS_BIAS.t2 GND 0.106594f
C4395 CS_BIAS.n7 GND 0.008917f
C4396 CS_BIAS.n8 GND 0.006753f
C4397 CS_BIAS.t12 GND 0.106594f
C4398 CS_BIAS.n9 GND 0.046728f
C4399 CS_BIAS.n10 GND 0.006753f
C4400 CS_BIAS.n11 GND 0.013528f
C4401 CS_BIAS.n12 GND 0.006753f
C4402 CS_BIAS.t0 GND 0.106594f
C4403 CS_BIAS.n13 GND 0.006379f
C4404 CS_BIAS.n14 GND 0.06363f
C4405 CS_BIAS.t4 GND 0.106594f
C4406 CS_BIAS.t14 GND 0.153124f
C4407 CS_BIAS.n15 GND 0.062334f
C4408 CS_BIAS.n16 GND 0.067978f
C4409 CS_BIAS.n17 GND 0.011964f
C4410 CS_BIAS.n18 GND 0.012394f
C4411 CS_BIAS.n19 GND 0.006753f
C4412 CS_BIAS.n20 GND 0.006753f
C4413 CS_BIAS.n21 GND 0.006753f
C4414 CS_BIAS.n22 GND 0.013528f
C4415 CS_BIAS.n23 GND 0.009479f
C4416 CS_BIAS.n24 GND 0.046728f
C4417 CS_BIAS.n25 GND 0.009479f
C4418 CS_BIAS.n26 GND 0.006753f
C4419 CS_BIAS.n27 GND 0.006753f
C4420 CS_BIAS.n28 GND 0.006753f
C4421 CS_BIAS.n29 GND 0.006379f
C4422 CS_BIAS.n30 GND 0.012394f
C4423 CS_BIAS.n31 GND 0.011964f
C4424 CS_BIAS.n32 GND 0.006753f
C4425 CS_BIAS.n33 GND 0.006753f
C4426 CS_BIAS.n34 GND 0.006993f
C4427 CS_BIAS.n35 GND 0.012585f
C4428 CS_BIAS.n36 GND 0.010799f
C4429 CS_BIAS.n37 GND 0.006753f
C4430 CS_BIAS.n38 GND 0.006753f
C4431 CS_BIAS.n39 GND 0.006753f
C4432 CS_BIAS.n40 GND 0.012585f
C4433 CS_BIAS.n41 GND 0.008236f
C4434 CS_BIAS.n42 GND 0.066322f
C4435 CS_BIAS.n43 GND 0.053866f
C4436 CS_BIAS.n44 GND 0.003898f
C4437 CS_BIAS.n45 GND 0.023146f
C4438 CS_BIAS.n46 GND 0.001416f
C4439 CS_BIAS.t3 GND 0.006127f
C4440 CS_BIAS.n47 GND 0.009963f
C4441 CS_BIAS.n48 GND 0.002291f
C4442 CS_BIAS.n49 GND 0.002509f
C4443 CS_BIAS.n50 GND 0.007589f
C4444 CS_BIAS.n51 GND 0.001499f
C4445 CS_BIAS.n52 GND 0.001416f
C4446 CS_BIAS.n53 GND 0.005909f
C4447 CS_BIAS.n54 GND 0.007922f
C4448 CS_BIAS.n55 GND 0.080701f
C4449 CS_BIAS.t13 GND 0.005641f
C4450 CS_BIAS.t1 GND 0.005641f
C4451 CS_BIAS.n56 GND 0.043385f
C4452 CS_BIAS.n57 GND 0.07001f
C4453 CS_BIAS.t5 GND 0.005641f
C4454 CS_BIAS.t15 GND 0.005641f
C4455 CS_BIAS.n58 GND 0.044162f
C4456 CS_BIAS.n59 GND 0.170994f
C4457 CS_BIAS.n60 GND 0.043703f
C4458 CS_BIAS.t46 GND 0.106594f
C4459 CS_BIAS.n61 GND 0.013528f
C4460 CS_BIAS.n62 GND 0.006753f
C4461 CS_BIAS.t38 GND 0.106594f
C4462 CS_BIAS.n63 GND 0.067978f
C4463 CS_BIAS.t28 GND 0.153124f
C4464 CS_BIAS.n64 GND 0.062334f
C4465 CS_BIAS.n65 GND 0.06363f
C4466 CS_BIAS.n66 GND 0.011964f
C4467 CS_BIAS.n67 GND 0.012394f
C4468 CS_BIAS.n68 GND 0.006379f
C4469 CS_BIAS.n69 GND 0.006753f
C4470 CS_BIAS.n70 GND 0.006753f
C4471 CS_BIAS.n71 GND 0.005899f
C4472 CS_BIAS.n72 GND 0.009479f
C4473 CS_BIAS.n73 GND 0.046728f
C4474 CS_BIAS.n74 GND 0.009479f
C4475 CS_BIAS.n75 GND 0.005899f
C4476 CS_BIAS.n76 GND 0.006753f
C4477 CS_BIAS.n77 GND 0.006753f
C4478 CS_BIAS.n78 GND 0.006379f
C4479 CS_BIAS.n79 GND 0.012394f
C4480 CS_BIAS.n80 GND 0.011964f
C4481 CS_BIAS.n81 GND 0.006753f
C4482 CS_BIAS.n82 GND 0.006753f
C4483 CS_BIAS.n83 GND 0.006993f
C4484 CS_BIAS.n84 GND 0.012585f
C4485 CS_BIAS.n85 GND 0.010799f
C4486 CS_BIAS.n86 GND 0.006753f
C4487 CS_BIAS.n87 GND 0.006753f
C4488 CS_BIAS.n88 GND 0.006753f
C4489 CS_BIAS.n89 GND 0.012585f
C4490 CS_BIAS.n90 GND 0.008236f
C4491 CS_BIAS.n91 GND 0.066322f
C4492 CS_BIAS.n92 GND 0.034412f
C4493 CS_BIAS.n93 GND 0.008903f
C4494 CS_BIAS.t31 GND 0.106594f
C4495 CS_BIAS.n94 GND 0.008917f
C4496 CS_BIAS.n95 GND 0.006753f
C4497 CS_BIAS.t44 GND 0.106594f
C4498 CS_BIAS.n96 GND 0.046728f
C4499 CS_BIAS.n97 GND 0.006753f
C4500 CS_BIAS.n98 GND 0.013528f
C4501 CS_BIAS.n99 GND 0.006753f
C4502 CS_BIAS.t26 GND 0.106594f
C4503 CS_BIAS.n100 GND 0.006379f
C4504 CS_BIAS.n101 GND 0.06363f
C4505 CS_BIAS.t39 GND 0.106594f
C4506 CS_BIAS.t22 GND 0.153124f
C4507 CS_BIAS.n102 GND 0.062334f
C4508 CS_BIAS.n103 GND 0.067978f
C4509 CS_BIAS.n104 GND 0.011964f
C4510 CS_BIAS.n105 GND 0.012394f
C4511 CS_BIAS.n106 GND 0.006753f
C4512 CS_BIAS.n107 GND 0.006753f
C4513 CS_BIAS.n108 GND 0.006753f
C4514 CS_BIAS.n109 GND 0.013528f
C4515 CS_BIAS.n110 GND 0.009479f
C4516 CS_BIAS.n111 GND 0.046728f
C4517 CS_BIAS.n112 GND 0.009479f
C4518 CS_BIAS.n113 GND 0.006753f
C4519 CS_BIAS.n114 GND 0.006753f
C4520 CS_BIAS.n115 GND 0.006753f
C4521 CS_BIAS.n116 GND 0.006379f
C4522 CS_BIAS.n117 GND 0.012394f
C4523 CS_BIAS.n118 GND 0.011964f
C4524 CS_BIAS.n119 GND 0.006753f
C4525 CS_BIAS.n120 GND 0.006753f
C4526 CS_BIAS.n121 GND 0.006993f
C4527 CS_BIAS.n122 GND 0.012585f
C4528 CS_BIAS.n123 GND 0.010799f
C4529 CS_BIAS.n124 GND 0.006753f
C4530 CS_BIAS.n125 GND 0.006753f
C4531 CS_BIAS.n126 GND 0.006753f
C4532 CS_BIAS.n127 GND 0.012585f
C4533 CS_BIAS.n128 GND 0.008236f
C4534 CS_BIAS.n129 GND 0.066322f
C4535 CS_BIAS.n130 GND 0.026515f
C4536 CS_BIAS.n131 GND 0.067576f
C4537 CS_BIAS.n132 GND 0.008903f
C4538 CS_BIAS.t47 GND 0.106594f
C4539 CS_BIAS.n133 GND 0.008917f
C4540 CS_BIAS.n134 GND 0.006753f
C4541 CS_BIAS.t35 GND 0.106594f
C4542 CS_BIAS.n135 GND 0.046728f
C4543 CS_BIAS.n136 GND 0.006753f
C4544 CS_BIAS.n137 GND 0.013528f
C4545 CS_BIAS.n138 GND 0.006753f
C4546 CS_BIAS.t32 GND 0.106594f
C4547 CS_BIAS.n139 GND 0.006379f
C4548 CS_BIAS.n140 GND 0.06363f
C4549 CS_BIAS.t23 GND 0.106594f
C4550 CS_BIAS.t41 GND 0.153124f
C4551 CS_BIAS.n141 GND 0.062334f
C4552 CS_BIAS.n142 GND 0.067978f
C4553 CS_BIAS.n143 GND 0.011964f
C4554 CS_BIAS.n144 GND 0.012394f
C4555 CS_BIAS.n145 GND 0.006753f
C4556 CS_BIAS.n146 GND 0.006753f
C4557 CS_BIAS.n147 GND 0.006753f
C4558 CS_BIAS.n148 GND 0.013528f
C4559 CS_BIAS.n149 GND 0.009479f
C4560 CS_BIAS.n150 GND 0.046728f
C4561 CS_BIAS.n151 GND 0.009479f
C4562 CS_BIAS.n152 GND 0.006753f
C4563 CS_BIAS.n153 GND 0.006753f
C4564 CS_BIAS.n154 GND 0.006753f
C4565 CS_BIAS.n155 GND 0.006379f
C4566 CS_BIAS.n156 GND 0.012394f
C4567 CS_BIAS.n157 GND 0.011964f
C4568 CS_BIAS.n158 GND 0.006753f
C4569 CS_BIAS.n159 GND 0.006753f
C4570 CS_BIAS.n160 GND 0.006993f
C4571 CS_BIAS.n161 GND 0.012585f
C4572 CS_BIAS.n162 GND 0.010799f
C4573 CS_BIAS.n163 GND 0.006753f
C4574 CS_BIAS.n164 GND 0.006753f
C4575 CS_BIAS.n165 GND 0.006753f
C4576 CS_BIAS.n166 GND 0.012585f
C4577 CS_BIAS.n167 GND 0.008236f
C4578 CS_BIAS.n168 GND 0.066322f
C4579 CS_BIAS.n169 GND 0.026515f
C4580 CS_BIAS.n170 GND 0.714858f
C4581 CS_BIAS.n171 GND 0.008903f
C4582 CS_BIAS.t48 GND 0.106594f
C4583 CS_BIAS.n172 GND 0.008917f
C4584 CS_BIAS.n173 GND 0.006753f
C4585 CS_BIAS.t45 GND 0.106594f
C4586 CS_BIAS.n174 GND 0.046728f
C4587 CS_BIAS.n175 GND 0.006753f
C4588 CS_BIAS.n176 GND 0.013528f
C4589 CS_BIAS.n177 GND 0.003898f
C4590 CS_BIAS.n178 GND 0.023146f
C4591 CS_BIAS.n179 GND 0.001416f
C4592 CS_BIAS.t9 GND 0.006127f
C4593 CS_BIAS.n180 GND 0.009963f
C4594 CS_BIAS.n181 GND 0.002291f
C4595 CS_BIAS.n182 GND 0.002509f
C4596 CS_BIAS.n183 GND 0.007589f
C4597 CS_BIAS.n184 GND 0.001499f
C4598 CS_BIAS.n185 GND 0.001416f
C4599 CS_BIAS.n186 GND 0.005909f
C4600 CS_BIAS.n187 GND 0.008758f
C4601 CS_BIAS.t19 GND 0.005641f
C4602 CS_BIAS.t11 GND 0.005641f
C4603 CS_BIAS.n188 GND 0.043385f
C4604 CS_BIAS.n189 GND 0.116514f
C4605 CS_BIAS.n190 GND 0.008903f
C4606 CS_BIAS.t16 GND 0.106594f
C4607 CS_BIAS.n191 GND 0.008917f
C4608 CS_BIAS.n192 GND 0.006753f
C4609 CS_BIAS.t6 GND 0.106594f
C4610 CS_BIAS.n193 GND 0.046728f
C4611 CS_BIAS.n194 GND 0.006753f
C4612 CS_BIAS.n195 GND 0.013528f
C4613 CS_BIAS.n196 GND 0.006753f
C4614 CS_BIAS.t10 GND 0.106594f
C4615 CS_BIAS.n197 GND 0.006379f
C4616 CS_BIAS.n198 GND 0.06363f
C4617 CS_BIAS.t18 GND 0.106594f
C4618 CS_BIAS.t8 GND 0.153124f
C4619 CS_BIAS.n199 GND 0.062334f
C4620 CS_BIAS.n200 GND 0.067978f
C4621 CS_BIAS.n201 GND 0.011964f
C4622 CS_BIAS.n202 GND 0.012394f
C4623 CS_BIAS.n203 GND 0.006753f
C4624 CS_BIAS.n204 GND 0.006753f
C4625 CS_BIAS.n205 GND 0.006753f
C4626 CS_BIAS.n206 GND 0.013528f
C4627 CS_BIAS.n207 GND 0.009479f
C4628 CS_BIAS.n208 GND 0.046728f
C4629 CS_BIAS.n209 GND 0.009479f
C4630 CS_BIAS.n210 GND 0.006753f
C4631 CS_BIAS.n211 GND 0.006753f
C4632 CS_BIAS.n212 GND 0.006753f
C4633 CS_BIAS.n213 GND 0.006379f
C4634 CS_BIAS.n214 GND 0.012394f
C4635 CS_BIAS.n215 GND 0.011964f
C4636 CS_BIAS.n216 GND 0.006753f
C4637 CS_BIAS.n217 GND 0.006753f
C4638 CS_BIAS.n218 GND 0.006993f
C4639 CS_BIAS.n219 GND 0.012585f
C4640 CS_BIAS.n220 GND 0.010799f
C4641 CS_BIAS.n221 GND 0.006753f
C4642 CS_BIAS.n222 GND 0.006753f
C4643 CS_BIAS.n223 GND 0.006753f
C4644 CS_BIAS.n224 GND 0.012585f
C4645 CS_BIAS.n225 GND 0.008236f
C4646 CS_BIAS.n226 GND 0.066322f
C4647 CS_BIAS.n227 GND 0.056569f
C4648 CS_BIAS.t7 GND 0.005641f
C4649 CS_BIAS.t17 GND 0.005641f
C4650 CS_BIAS.n228 GND 0.043385f
C4651 CS_BIAS.n229 GND 0.122546f
C4652 CS_BIAS.n230 GND 0.079882f
C4653 CS_BIAS.n231 GND 0.043703f
C4654 CS_BIAS.t36 GND 0.106594f
C4655 CS_BIAS.n232 GND 0.013528f
C4656 CS_BIAS.n233 GND 0.006753f
C4657 CS_BIAS.t27 GND 0.106594f
C4658 CS_BIAS.n234 GND 0.067978f
C4659 CS_BIAS.t24 GND 0.153124f
C4660 CS_BIAS.n235 GND 0.062334f
C4661 CS_BIAS.n236 GND 0.06363f
C4662 CS_BIAS.n237 GND 0.011964f
C4663 CS_BIAS.n238 GND 0.012394f
C4664 CS_BIAS.n239 GND 0.006379f
C4665 CS_BIAS.n240 GND 0.006753f
C4666 CS_BIAS.n241 GND 0.006753f
C4667 CS_BIAS.n242 GND 0.005899f
C4668 CS_BIAS.n243 GND 0.009479f
C4669 CS_BIAS.n244 GND 0.046728f
C4670 CS_BIAS.n245 GND 0.009479f
C4671 CS_BIAS.n246 GND 0.005899f
C4672 CS_BIAS.n247 GND 0.006753f
C4673 CS_BIAS.n248 GND 0.006753f
C4674 CS_BIAS.n249 GND 0.006379f
C4675 CS_BIAS.n250 GND 0.012394f
C4676 CS_BIAS.n251 GND 0.011964f
C4677 CS_BIAS.n252 GND 0.006753f
C4678 CS_BIAS.n253 GND 0.006753f
C4679 CS_BIAS.n254 GND 0.006993f
C4680 CS_BIAS.n255 GND 0.012585f
C4681 CS_BIAS.n256 GND 0.010799f
C4682 CS_BIAS.n257 GND 0.006753f
C4683 CS_BIAS.n258 GND 0.006753f
C4684 CS_BIAS.n259 GND 0.006753f
C4685 CS_BIAS.n260 GND 0.012585f
C4686 CS_BIAS.n261 GND 0.008236f
C4687 CS_BIAS.n262 GND 0.066322f
C4688 CS_BIAS.n263 GND 0.034412f
C4689 CS_BIAS.n264 GND 0.008903f
C4690 CS_BIAS.t43 GND 0.106594f
C4691 CS_BIAS.n265 GND 0.008917f
C4692 CS_BIAS.n266 GND 0.006753f
C4693 CS_BIAS.t21 GND 0.106594f
C4694 CS_BIAS.n267 GND 0.046728f
C4695 CS_BIAS.n268 GND 0.006753f
C4696 CS_BIAS.n269 GND 0.013528f
C4697 CS_BIAS.n270 GND 0.006753f
C4698 CS_BIAS.t37 GND 0.106594f
C4699 CS_BIAS.n271 GND 0.006379f
C4700 CS_BIAS.n272 GND 0.06363f
C4701 CS_BIAS.t20 GND 0.106594f
C4702 CS_BIAS.t29 GND 0.153124f
C4703 CS_BIAS.n273 GND 0.062334f
C4704 CS_BIAS.n274 GND 0.067978f
C4705 CS_BIAS.n275 GND 0.011964f
C4706 CS_BIAS.n276 GND 0.012394f
C4707 CS_BIAS.n277 GND 0.006753f
C4708 CS_BIAS.n278 GND 0.006753f
C4709 CS_BIAS.n279 GND 0.006753f
C4710 CS_BIAS.n280 GND 0.013528f
C4711 CS_BIAS.n281 GND 0.009479f
C4712 CS_BIAS.n282 GND 0.046728f
C4713 CS_BIAS.n283 GND 0.009479f
C4714 CS_BIAS.n284 GND 0.006753f
C4715 CS_BIAS.n285 GND 0.006753f
C4716 CS_BIAS.n286 GND 0.006753f
C4717 CS_BIAS.n287 GND 0.006379f
C4718 CS_BIAS.n288 GND 0.012394f
C4719 CS_BIAS.n289 GND 0.011964f
C4720 CS_BIAS.n290 GND 0.006753f
C4721 CS_BIAS.n291 GND 0.006753f
C4722 CS_BIAS.n292 GND 0.006993f
C4723 CS_BIAS.n293 GND 0.012585f
C4724 CS_BIAS.n294 GND 0.010799f
C4725 CS_BIAS.n295 GND 0.006753f
C4726 CS_BIAS.n296 GND 0.006753f
C4727 CS_BIAS.n297 GND 0.006753f
C4728 CS_BIAS.n298 GND 0.012585f
C4729 CS_BIAS.n299 GND 0.008236f
C4730 CS_BIAS.n300 GND 0.066322f
C4731 CS_BIAS.n301 GND 0.026515f
C4732 CS_BIAS.n302 GND 0.067576f
C4733 CS_BIAS.n303 GND 0.008903f
C4734 CS_BIAS.t34 GND 0.106594f
C4735 CS_BIAS.n304 GND 0.008917f
C4736 CS_BIAS.n305 GND 0.006753f
C4737 CS_BIAS.t33 GND 0.106594f
C4738 CS_BIAS.n306 GND 0.046728f
C4739 CS_BIAS.n307 GND 0.006753f
C4740 CS_BIAS.n308 GND 0.013528f
C4741 CS_BIAS.n309 GND 0.006753f
C4742 CS_BIAS.t25 GND 0.106594f
C4743 CS_BIAS.n310 GND 0.006379f
C4744 CS_BIAS.n311 GND 0.06363f
C4745 CS_BIAS.t42 GND 0.106594f
C4746 CS_BIAS.t40 GND 0.153124f
C4747 CS_BIAS.n312 GND 0.062334f
C4748 CS_BIAS.n313 GND 0.067978f
C4749 CS_BIAS.n314 GND 0.011964f
C4750 CS_BIAS.n315 GND 0.012394f
C4751 CS_BIAS.n316 GND 0.006753f
C4752 CS_BIAS.n317 GND 0.006753f
C4753 CS_BIAS.n318 GND 0.006753f
C4754 CS_BIAS.n319 GND 0.013528f
C4755 CS_BIAS.n320 GND 0.009479f
C4756 CS_BIAS.n321 GND 0.046728f
C4757 CS_BIAS.n322 GND 0.009479f
C4758 CS_BIAS.n323 GND 0.006753f
C4759 CS_BIAS.n324 GND 0.006753f
C4760 CS_BIAS.n325 GND 0.006753f
C4761 CS_BIAS.n326 GND 0.006379f
C4762 CS_BIAS.n327 GND 0.012394f
C4763 CS_BIAS.n328 GND 0.011964f
C4764 CS_BIAS.n329 GND 0.006753f
C4765 CS_BIAS.n330 GND 0.006753f
C4766 CS_BIAS.n331 GND 0.006993f
C4767 CS_BIAS.n332 GND 0.012585f
C4768 CS_BIAS.n333 GND 0.010799f
C4769 CS_BIAS.n334 GND 0.006753f
C4770 CS_BIAS.n335 GND 0.006753f
C4771 CS_BIAS.n336 GND 0.006753f
C4772 CS_BIAS.n337 GND 0.012585f
C4773 CS_BIAS.n338 GND 0.008236f
C4774 CS_BIAS.n339 GND 0.066322f
C4775 CS_BIAS.n340 GND 0.026515f
C4776 CS_BIAS.n341 GND 0.134813f
C4777 CS_BIAS.n342 GND 5.41392f
.ends

