* NGSPICE file created from diff_pair_sample_0581.ext - technology: sky130A

.subckt diff_pair_sample_0581 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t5 VN.t0 VDD2.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5015 pd=8.48 as=0.63525 ps=4.18 w=3.85 l=3.82
X1 VTAIL.t7 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5015 pd=8.48 as=0.63525 ps=4.18 w=3.85 l=3.82
X2 VTAIL.t4 VN.t1 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5015 pd=8.48 as=0.63525 ps=4.18 w=3.85 l=3.82
X3 VDD2.t3 VN.t2 VTAIL.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=0.63525 pd=4.18 as=1.5015 ps=8.48 w=3.85 l=3.82
X4 VDD1.t2 VP.t1 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=0.63525 pd=4.18 as=1.5015 ps=8.48 w=3.85 l=3.82
X5 VDD2.t1 VN.t3 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.63525 pd=4.18 as=1.5015 ps=8.48 w=3.85 l=3.82
X6 VDD1.t1 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.63525 pd=4.18 as=1.5015 ps=8.48 w=3.85 l=3.82
X7 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=1.5015 pd=8.48 as=0 ps=0 w=3.85 l=3.82
X8 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5015 pd=8.48 as=0 ps=0 w=3.85 l=3.82
X9 VTAIL.t0 VP.t3 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5015 pd=8.48 as=0.63525 ps=4.18 w=3.85 l=3.82
X10 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.5015 pd=8.48 as=0 ps=0 w=3.85 l=3.82
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5015 pd=8.48 as=0 ps=0 w=3.85 l=3.82
R0 VN.n0 VN.t0 58.3545
R1 VN.n1 VN.t3 58.3545
R2 VN.n0 VN.t2 56.9995
R3 VN.n1 VN.t1 56.9995
R4 VN VN.n1 45.952
R5 VN VN.n0 1.84216
R6 VDD2.n2 VDD2.n0 111.424
R7 VDD2.n2 VDD2.n1 73.6579
R8 VDD2.n1 VDD2.t0 5.14336
R9 VDD2.n1 VDD2.t1 5.14336
R10 VDD2.n0 VDD2.t2 5.14336
R11 VDD2.n0 VDD2.t3 5.14336
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n154 VTAIL.n140 289.615
R14 VTAIL.n14 VTAIL.n0 289.615
R15 VTAIL.n34 VTAIL.n20 289.615
R16 VTAIL.n54 VTAIL.n40 289.615
R17 VTAIL.n134 VTAIL.n120 289.615
R18 VTAIL.n114 VTAIL.n100 289.615
R19 VTAIL.n94 VTAIL.n80 289.615
R20 VTAIL.n74 VTAIL.n60 289.615
R21 VTAIL.n147 VTAIL.n146 185
R22 VTAIL.n144 VTAIL.n143 185
R23 VTAIL.n153 VTAIL.n152 185
R24 VTAIL.n155 VTAIL.n154 185
R25 VTAIL.n7 VTAIL.n6 185
R26 VTAIL.n4 VTAIL.n3 185
R27 VTAIL.n13 VTAIL.n12 185
R28 VTAIL.n15 VTAIL.n14 185
R29 VTAIL.n27 VTAIL.n26 185
R30 VTAIL.n24 VTAIL.n23 185
R31 VTAIL.n33 VTAIL.n32 185
R32 VTAIL.n35 VTAIL.n34 185
R33 VTAIL.n47 VTAIL.n46 185
R34 VTAIL.n44 VTAIL.n43 185
R35 VTAIL.n53 VTAIL.n52 185
R36 VTAIL.n55 VTAIL.n54 185
R37 VTAIL.n135 VTAIL.n134 185
R38 VTAIL.n133 VTAIL.n132 185
R39 VTAIL.n124 VTAIL.n123 185
R40 VTAIL.n127 VTAIL.n126 185
R41 VTAIL.n115 VTAIL.n114 185
R42 VTAIL.n113 VTAIL.n112 185
R43 VTAIL.n104 VTAIL.n103 185
R44 VTAIL.n107 VTAIL.n106 185
R45 VTAIL.n95 VTAIL.n94 185
R46 VTAIL.n93 VTAIL.n92 185
R47 VTAIL.n84 VTAIL.n83 185
R48 VTAIL.n87 VTAIL.n86 185
R49 VTAIL.n75 VTAIL.n74 185
R50 VTAIL.n73 VTAIL.n72 185
R51 VTAIL.n64 VTAIL.n63 185
R52 VTAIL.n67 VTAIL.n66 185
R53 VTAIL.t3 VTAIL.n145 147.888
R54 VTAIL.t5 VTAIL.n5 147.888
R55 VTAIL.t1 VTAIL.n25 147.888
R56 VTAIL.t7 VTAIL.n45 147.888
R57 VTAIL.t6 VTAIL.n125 147.888
R58 VTAIL.t0 VTAIL.n105 147.888
R59 VTAIL.t2 VTAIL.n85 147.888
R60 VTAIL.t4 VTAIL.n65 147.888
R61 VTAIL.n146 VTAIL.n143 104.615
R62 VTAIL.n153 VTAIL.n143 104.615
R63 VTAIL.n154 VTAIL.n153 104.615
R64 VTAIL.n6 VTAIL.n3 104.615
R65 VTAIL.n13 VTAIL.n3 104.615
R66 VTAIL.n14 VTAIL.n13 104.615
R67 VTAIL.n26 VTAIL.n23 104.615
R68 VTAIL.n33 VTAIL.n23 104.615
R69 VTAIL.n34 VTAIL.n33 104.615
R70 VTAIL.n46 VTAIL.n43 104.615
R71 VTAIL.n53 VTAIL.n43 104.615
R72 VTAIL.n54 VTAIL.n53 104.615
R73 VTAIL.n134 VTAIL.n133 104.615
R74 VTAIL.n133 VTAIL.n123 104.615
R75 VTAIL.n126 VTAIL.n123 104.615
R76 VTAIL.n114 VTAIL.n113 104.615
R77 VTAIL.n113 VTAIL.n103 104.615
R78 VTAIL.n106 VTAIL.n103 104.615
R79 VTAIL.n94 VTAIL.n93 104.615
R80 VTAIL.n93 VTAIL.n83 104.615
R81 VTAIL.n86 VTAIL.n83 104.615
R82 VTAIL.n74 VTAIL.n73 104.615
R83 VTAIL.n73 VTAIL.n63 104.615
R84 VTAIL.n66 VTAIL.n63 104.615
R85 VTAIL.n146 VTAIL.t3 52.3082
R86 VTAIL.n6 VTAIL.t5 52.3082
R87 VTAIL.n26 VTAIL.t1 52.3082
R88 VTAIL.n46 VTAIL.t7 52.3082
R89 VTAIL.n126 VTAIL.t6 52.3082
R90 VTAIL.n106 VTAIL.t0 52.3082
R91 VTAIL.n86 VTAIL.t2 52.3082
R92 VTAIL.n66 VTAIL.t4 52.3082
R93 VTAIL.n159 VTAIL.n158 32.3793
R94 VTAIL.n19 VTAIL.n18 32.3793
R95 VTAIL.n39 VTAIL.n38 32.3793
R96 VTAIL.n59 VTAIL.n58 32.3793
R97 VTAIL.n139 VTAIL.n138 32.3793
R98 VTAIL.n119 VTAIL.n118 32.3793
R99 VTAIL.n99 VTAIL.n98 32.3793
R100 VTAIL.n79 VTAIL.n78 32.3793
R101 VTAIL.n159 VTAIL.n139 19.2634
R102 VTAIL.n79 VTAIL.n59 19.2634
R103 VTAIL.n147 VTAIL.n145 15.6496
R104 VTAIL.n7 VTAIL.n5 15.6496
R105 VTAIL.n27 VTAIL.n25 15.6496
R106 VTAIL.n47 VTAIL.n45 15.6496
R107 VTAIL.n127 VTAIL.n125 15.6496
R108 VTAIL.n107 VTAIL.n105 15.6496
R109 VTAIL.n87 VTAIL.n85 15.6496
R110 VTAIL.n67 VTAIL.n65 15.6496
R111 VTAIL.n148 VTAIL.n144 12.8005
R112 VTAIL.n8 VTAIL.n4 12.8005
R113 VTAIL.n28 VTAIL.n24 12.8005
R114 VTAIL.n48 VTAIL.n44 12.8005
R115 VTAIL.n128 VTAIL.n124 12.8005
R116 VTAIL.n108 VTAIL.n104 12.8005
R117 VTAIL.n88 VTAIL.n84 12.8005
R118 VTAIL.n68 VTAIL.n64 12.8005
R119 VTAIL.n152 VTAIL.n151 12.0247
R120 VTAIL.n12 VTAIL.n11 12.0247
R121 VTAIL.n32 VTAIL.n31 12.0247
R122 VTAIL.n52 VTAIL.n51 12.0247
R123 VTAIL.n132 VTAIL.n131 12.0247
R124 VTAIL.n112 VTAIL.n111 12.0247
R125 VTAIL.n92 VTAIL.n91 12.0247
R126 VTAIL.n72 VTAIL.n71 12.0247
R127 VTAIL.n155 VTAIL.n142 11.249
R128 VTAIL.n15 VTAIL.n2 11.249
R129 VTAIL.n35 VTAIL.n22 11.249
R130 VTAIL.n55 VTAIL.n42 11.249
R131 VTAIL.n135 VTAIL.n122 11.249
R132 VTAIL.n115 VTAIL.n102 11.249
R133 VTAIL.n95 VTAIL.n82 11.249
R134 VTAIL.n75 VTAIL.n62 11.249
R135 VTAIL.n156 VTAIL.n140 10.4732
R136 VTAIL.n16 VTAIL.n0 10.4732
R137 VTAIL.n36 VTAIL.n20 10.4732
R138 VTAIL.n56 VTAIL.n40 10.4732
R139 VTAIL.n136 VTAIL.n120 10.4732
R140 VTAIL.n116 VTAIL.n100 10.4732
R141 VTAIL.n96 VTAIL.n80 10.4732
R142 VTAIL.n76 VTAIL.n60 10.4732
R143 VTAIL.n158 VTAIL.n157 9.45567
R144 VTAIL.n18 VTAIL.n17 9.45567
R145 VTAIL.n38 VTAIL.n37 9.45567
R146 VTAIL.n58 VTAIL.n57 9.45567
R147 VTAIL.n138 VTAIL.n137 9.45567
R148 VTAIL.n118 VTAIL.n117 9.45567
R149 VTAIL.n98 VTAIL.n97 9.45567
R150 VTAIL.n78 VTAIL.n77 9.45567
R151 VTAIL.n157 VTAIL.n156 9.3005
R152 VTAIL.n142 VTAIL.n141 9.3005
R153 VTAIL.n151 VTAIL.n150 9.3005
R154 VTAIL.n149 VTAIL.n148 9.3005
R155 VTAIL.n17 VTAIL.n16 9.3005
R156 VTAIL.n2 VTAIL.n1 9.3005
R157 VTAIL.n11 VTAIL.n10 9.3005
R158 VTAIL.n9 VTAIL.n8 9.3005
R159 VTAIL.n37 VTAIL.n36 9.3005
R160 VTAIL.n22 VTAIL.n21 9.3005
R161 VTAIL.n31 VTAIL.n30 9.3005
R162 VTAIL.n29 VTAIL.n28 9.3005
R163 VTAIL.n57 VTAIL.n56 9.3005
R164 VTAIL.n42 VTAIL.n41 9.3005
R165 VTAIL.n51 VTAIL.n50 9.3005
R166 VTAIL.n49 VTAIL.n48 9.3005
R167 VTAIL.n137 VTAIL.n136 9.3005
R168 VTAIL.n122 VTAIL.n121 9.3005
R169 VTAIL.n131 VTAIL.n130 9.3005
R170 VTAIL.n129 VTAIL.n128 9.3005
R171 VTAIL.n117 VTAIL.n116 9.3005
R172 VTAIL.n102 VTAIL.n101 9.3005
R173 VTAIL.n111 VTAIL.n110 9.3005
R174 VTAIL.n109 VTAIL.n108 9.3005
R175 VTAIL.n97 VTAIL.n96 9.3005
R176 VTAIL.n82 VTAIL.n81 9.3005
R177 VTAIL.n91 VTAIL.n90 9.3005
R178 VTAIL.n89 VTAIL.n88 9.3005
R179 VTAIL.n77 VTAIL.n76 9.3005
R180 VTAIL.n62 VTAIL.n61 9.3005
R181 VTAIL.n71 VTAIL.n70 9.3005
R182 VTAIL.n69 VTAIL.n68 9.3005
R183 VTAIL.n149 VTAIL.n145 4.40546
R184 VTAIL.n9 VTAIL.n5 4.40546
R185 VTAIL.n29 VTAIL.n25 4.40546
R186 VTAIL.n49 VTAIL.n45 4.40546
R187 VTAIL.n129 VTAIL.n125 4.40546
R188 VTAIL.n109 VTAIL.n105 4.40546
R189 VTAIL.n89 VTAIL.n85 4.40546
R190 VTAIL.n69 VTAIL.n65 4.40546
R191 VTAIL.n99 VTAIL.n79 3.57809
R192 VTAIL.n139 VTAIL.n119 3.57809
R193 VTAIL.n59 VTAIL.n39 3.57809
R194 VTAIL.n158 VTAIL.n140 3.49141
R195 VTAIL.n18 VTAIL.n0 3.49141
R196 VTAIL.n38 VTAIL.n20 3.49141
R197 VTAIL.n58 VTAIL.n40 3.49141
R198 VTAIL.n138 VTAIL.n120 3.49141
R199 VTAIL.n118 VTAIL.n100 3.49141
R200 VTAIL.n98 VTAIL.n80 3.49141
R201 VTAIL.n78 VTAIL.n60 3.49141
R202 VTAIL.n156 VTAIL.n155 2.71565
R203 VTAIL.n16 VTAIL.n15 2.71565
R204 VTAIL.n36 VTAIL.n35 2.71565
R205 VTAIL.n56 VTAIL.n55 2.71565
R206 VTAIL.n136 VTAIL.n135 2.71565
R207 VTAIL.n116 VTAIL.n115 2.71565
R208 VTAIL.n96 VTAIL.n95 2.71565
R209 VTAIL.n76 VTAIL.n75 2.71565
R210 VTAIL.n152 VTAIL.n142 1.93989
R211 VTAIL.n12 VTAIL.n2 1.93989
R212 VTAIL.n32 VTAIL.n22 1.93989
R213 VTAIL.n52 VTAIL.n42 1.93989
R214 VTAIL.n132 VTAIL.n122 1.93989
R215 VTAIL.n112 VTAIL.n102 1.93989
R216 VTAIL.n92 VTAIL.n82 1.93989
R217 VTAIL.n72 VTAIL.n62 1.93989
R218 VTAIL VTAIL.n19 1.84748
R219 VTAIL VTAIL.n159 1.7311
R220 VTAIL.n151 VTAIL.n144 1.16414
R221 VTAIL.n11 VTAIL.n4 1.16414
R222 VTAIL.n31 VTAIL.n24 1.16414
R223 VTAIL.n51 VTAIL.n44 1.16414
R224 VTAIL.n131 VTAIL.n124 1.16414
R225 VTAIL.n111 VTAIL.n104 1.16414
R226 VTAIL.n91 VTAIL.n84 1.16414
R227 VTAIL.n71 VTAIL.n64 1.16414
R228 VTAIL.n119 VTAIL.n99 0.470328
R229 VTAIL.n39 VTAIL.n19 0.470328
R230 VTAIL.n148 VTAIL.n147 0.388379
R231 VTAIL.n8 VTAIL.n7 0.388379
R232 VTAIL.n28 VTAIL.n27 0.388379
R233 VTAIL.n48 VTAIL.n47 0.388379
R234 VTAIL.n128 VTAIL.n127 0.388379
R235 VTAIL.n108 VTAIL.n107 0.388379
R236 VTAIL.n88 VTAIL.n87 0.388379
R237 VTAIL.n68 VTAIL.n67 0.388379
R238 VTAIL.n150 VTAIL.n149 0.155672
R239 VTAIL.n150 VTAIL.n141 0.155672
R240 VTAIL.n157 VTAIL.n141 0.155672
R241 VTAIL.n10 VTAIL.n9 0.155672
R242 VTAIL.n10 VTAIL.n1 0.155672
R243 VTAIL.n17 VTAIL.n1 0.155672
R244 VTAIL.n30 VTAIL.n29 0.155672
R245 VTAIL.n30 VTAIL.n21 0.155672
R246 VTAIL.n37 VTAIL.n21 0.155672
R247 VTAIL.n50 VTAIL.n49 0.155672
R248 VTAIL.n50 VTAIL.n41 0.155672
R249 VTAIL.n57 VTAIL.n41 0.155672
R250 VTAIL.n137 VTAIL.n121 0.155672
R251 VTAIL.n130 VTAIL.n121 0.155672
R252 VTAIL.n130 VTAIL.n129 0.155672
R253 VTAIL.n117 VTAIL.n101 0.155672
R254 VTAIL.n110 VTAIL.n101 0.155672
R255 VTAIL.n110 VTAIL.n109 0.155672
R256 VTAIL.n97 VTAIL.n81 0.155672
R257 VTAIL.n90 VTAIL.n81 0.155672
R258 VTAIL.n90 VTAIL.n89 0.155672
R259 VTAIL.n77 VTAIL.n61 0.155672
R260 VTAIL.n70 VTAIL.n61 0.155672
R261 VTAIL.n70 VTAIL.n69 0.155672
R262 B.n593 B.n592 585
R263 B.n594 B.n593 585
R264 B.n197 B.n106 585
R265 B.n196 B.n195 585
R266 B.n194 B.n193 585
R267 B.n192 B.n191 585
R268 B.n190 B.n189 585
R269 B.n188 B.n187 585
R270 B.n186 B.n185 585
R271 B.n184 B.n183 585
R272 B.n182 B.n181 585
R273 B.n180 B.n179 585
R274 B.n178 B.n177 585
R275 B.n176 B.n175 585
R276 B.n174 B.n173 585
R277 B.n172 B.n171 585
R278 B.n170 B.n169 585
R279 B.n168 B.n167 585
R280 B.n166 B.n165 585
R281 B.n163 B.n162 585
R282 B.n161 B.n160 585
R283 B.n159 B.n158 585
R284 B.n157 B.n156 585
R285 B.n155 B.n154 585
R286 B.n153 B.n152 585
R287 B.n151 B.n150 585
R288 B.n149 B.n148 585
R289 B.n147 B.n146 585
R290 B.n145 B.n144 585
R291 B.n143 B.n142 585
R292 B.n141 B.n140 585
R293 B.n139 B.n138 585
R294 B.n137 B.n136 585
R295 B.n135 B.n134 585
R296 B.n133 B.n132 585
R297 B.n131 B.n130 585
R298 B.n129 B.n128 585
R299 B.n127 B.n126 585
R300 B.n125 B.n124 585
R301 B.n123 B.n122 585
R302 B.n121 B.n120 585
R303 B.n119 B.n118 585
R304 B.n117 B.n116 585
R305 B.n115 B.n114 585
R306 B.n113 B.n112 585
R307 B.n82 B.n81 585
R308 B.n591 B.n83 585
R309 B.n595 B.n83 585
R310 B.n590 B.n589 585
R311 B.n589 B.n79 585
R312 B.n588 B.n78 585
R313 B.n601 B.n78 585
R314 B.n587 B.n77 585
R315 B.n602 B.n77 585
R316 B.n586 B.n76 585
R317 B.n603 B.n76 585
R318 B.n585 B.n584 585
R319 B.n584 B.n72 585
R320 B.n583 B.n71 585
R321 B.n609 B.n71 585
R322 B.n582 B.n70 585
R323 B.n610 B.n70 585
R324 B.n581 B.n69 585
R325 B.n611 B.n69 585
R326 B.n580 B.n579 585
R327 B.n579 B.n68 585
R328 B.n578 B.n64 585
R329 B.n617 B.n64 585
R330 B.n577 B.n63 585
R331 B.n618 B.n63 585
R332 B.n576 B.n62 585
R333 B.n619 B.n62 585
R334 B.n575 B.n574 585
R335 B.n574 B.n58 585
R336 B.n573 B.n57 585
R337 B.n625 B.n57 585
R338 B.n572 B.n56 585
R339 B.n626 B.n56 585
R340 B.n571 B.n55 585
R341 B.n627 B.n55 585
R342 B.n570 B.n569 585
R343 B.n569 B.n51 585
R344 B.n568 B.n50 585
R345 B.n633 B.n50 585
R346 B.n567 B.n49 585
R347 B.n634 B.n49 585
R348 B.n566 B.n48 585
R349 B.n635 B.n48 585
R350 B.n565 B.n564 585
R351 B.n564 B.n44 585
R352 B.n563 B.n43 585
R353 B.n641 B.n43 585
R354 B.n562 B.n42 585
R355 B.n642 B.n42 585
R356 B.n561 B.n41 585
R357 B.n643 B.n41 585
R358 B.n560 B.n559 585
R359 B.n559 B.n37 585
R360 B.n558 B.n36 585
R361 B.n649 B.n36 585
R362 B.n557 B.n35 585
R363 B.n650 B.n35 585
R364 B.n556 B.n34 585
R365 B.n651 B.n34 585
R366 B.n555 B.n554 585
R367 B.n554 B.n30 585
R368 B.n553 B.n29 585
R369 B.n657 B.n29 585
R370 B.n552 B.n28 585
R371 B.n658 B.n28 585
R372 B.n551 B.n27 585
R373 B.n659 B.n27 585
R374 B.n550 B.n549 585
R375 B.n549 B.n23 585
R376 B.n548 B.n22 585
R377 B.n665 B.n22 585
R378 B.n547 B.n21 585
R379 B.n666 B.n21 585
R380 B.n546 B.n20 585
R381 B.n667 B.n20 585
R382 B.n545 B.n544 585
R383 B.n544 B.n16 585
R384 B.n543 B.n15 585
R385 B.n673 B.n15 585
R386 B.n542 B.n14 585
R387 B.n674 B.n14 585
R388 B.n541 B.n13 585
R389 B.n675 B.n13 585
R390 B.n540 B.n539 585
R391 B.n539 B.n12 585
R392 B.n538 B.n537 585
R393 B.n538 B.n8 585
R394 B.n536 B.n7 585
R395 B.n682 B.n7 585
R396 B.n535 B.n6 585
R397 B.n683 B.n6 585
R398 B.n534 B.n5 585
R399 B.n684 B.n5 585
R400 B.n533 B.n532 585
R401 B.n532 B.n4 585
R402 B.n531 B.n198 585
R403 B.n531 B.n530 585
R404 B.n521 B.n199 585
R405 B.n200 B.n199 585
R406 B.n523 B.n522 585
R407 B.n524 B.n523 585
R408 B.n520 B.n205 585
R409 B.n205 B.n204 585
R410 B.n519 B.n518 585
R411 B.n518 B.n517 585
R412 B.n207 B.n206 585
R413 B.n208 B.n207 585
R414 B.n510 B.n509 585
R415 B.n511 B.n510 585
R416 B.n508 B.n213 585
R417 B.n213 B.n212 585
R418 B.n507 B.n506 585
R419 B.n506 B.n505 585
R420 B.n215 B.n214 585
R421 B.n216 B.n215 585
R422 B.n498 B.n497 585
R423 B.n499 B.n498 585
R424 B.n496 B.n221 585
R425 B.n221 B.n220 585
R426 B.n495 B.n494 585
R427 B.n494 B.n493 585
R428 B.n223 B.n222 585
R429 B.n224 B.n223 585
R430 B.n486 B.n485 585
R431 B.n487 B.n486 585
R432 B.n484 B.n229 585
R433 B.n229 B.n228 585
R434 B.n483 B.n482 585
R435 B.n482 B.n481 585
R436 B.n231 B.n230 585
R437 B.n232 B.n231 585
R438 B.n474 B.n473 585
R439 B.n475 B.n474 585
R440 B.n472 B.n237 585
R441 B.n237 B.n236 585
R442 B.n471 B.n470 585
R443 B.n470 B.n469 585
R444 B.n239 B.n238 585
R445 B.n240 B.n239 585
R446 B.n462 B.n461 585
R447 B.n463 B.n462 585
R448 B.n460 B.n245 585
R449 B.n245 B.n244 585
R450 B.n459 B.n458 585
R451 B.n458 B.n457 585
R452 B.n247 B.n246 585
R453 B.n248 B.n247 585
R454 B.n450 B.n449 585
R455 B.n451 B.n450 585
R456 B.n448 B.n253 585
R457 B.n253 B.n252 585
R458 B.n447 B.n446 585
R459 B.n446 B.n445 585
R460 B.n255 B.n254 585
R461 B.n256 B.n255 585
R462 B.n438 B.n437 585
R463 B.n439 B.n438 585
R464 B.n436 B.n261 585
R465 B.n261 B.n260 585
R466 B.n435 B.n434 585
R467 B.n434 B.n433 585
R468 B.n263 B.n262 585
R469 B.n426 B.n263 585
R470 B.n425 B.n424 585
R471 B.n427 B.n425 585
R472 B.n423 B.n268 585
R473 B.n268 B.n267 585
R474 B.n422 B.n421 585
R475 B.n421 B.n420 585
R476 B.n270 B.n269 585
R477 B.n271 B.n270 585
R478 B.n413 B.n412 585
R479 B.n414 B.n413 585
R480 B.n411 B.n276 585
R481 B.n276 B.n275 585
R482 B.n410 B.n409 585
R483 B.n409 B.n408 585
R484 B.n278 B.n277 585
R485 B.n279 B.n278 585
R486 B.n401 B.n400 585
R487 B.n402 B.n401 585
R488 B.n282 B.n281 585
R489 B.n311 B.n309 585
R490 B.n312 B.n308 585
R491 B.n312 B.n283 585
R492 B.n315 B.n314 585
R493 B.n316 B.n307 585
R494 B.n318 B.n317 585
R495 B.n320 B.n306 585
R496 B.n323 B.n322 585
R497 B.n324 B.n305 585
R498 B.n326 B.n325 585
R499 B.n328 B.n304 585
R500 B.n331 B.n330 585
R501 B.n332 B.n303 585
R502 B.n334 B.n333 585
R503 B.n336 B.n302 585
R504 B.n339 B.n338 585
R505 B.n340 B.n301 585
R506 B.n345 B.n344 585
R507 B.n347 B.n300 585
R508 B.n350 B.n349 585
R509 B.n351 B.n299 585
R510 B.n353 B.n352 585
R511 B.n355 B.n298 585
R512 B.n358 B.n357 585
R513 B.n359 B.n297 585
R514 B.n361 B.n360 585
R515 B.n363 B.n296 585
R516 B.n366 B.n365 585
R517 B.n367 B.n292 585
R518 B.n369 B.n368 585
R519 B.n371 B.n291 585
R520 B.n374 B.n373 585
R521 B.n375 B.n290 585
R522 B.n377 B.n376 585
R523 B.n379 B.n289 585
R524 B.n382 B.n381 585
R525 B.n383 B.n288 585
R526 B.n385 B.n384 585
R527 B.n387 B.n287 585
R528 B.n390 B.n389 585
R529 B.n391 B.n286 585
R530 B.n393 B.n392 585
R531 B.n395 B.n285 585
R532 B.n398 B.n397 585
R533 B.n399 B.n284 585
R534 B.n404 B.n403 585
R535 B.n403 B.n402 585
R536 B.n405 B.n280 585
R537 B.n280 B.n279 585
R538 B.n407 B.n406 585
R539 B.n408 B.n407 585
R540 B.n274 B.n273 585
R541 B.n275 B.n274 585
R542 B.n416 B.n415 585
R543 B.n415 B.n414 585
R544 B.n417 B.n272 585
R545 B.n272 B.n271 585
R546 B.n419 B.n418 585
R547 B.n420 B.n419 585
R548 B.n266 B.n265 585
R549 B.n267 B.n266 585
R550 B.n429 B.n428 585
R551 B.n428 B.n427 585
R552 B.n430 B.n264 585
R553 B.n426 B.n264 585
R554 B.n432 B.n431 585
R555 B.n433 B.n432 585
R556 B.n259 B.n258 585
R557 B.n260 B.n259 585
R558 B.n441 B.n440 585
R559 B.n440 B.n439 585
R560 B.n442 B.n257 585
R561 B.n257 B.n256 585
R562 B.n444 B.n443 585
R563 B.n445 B.n444 585
R564 B.n251 B.n250 585
R565 B.n252 B.n251 585
R566 B.n453 B.n452 585
R567 B.n452 B.n451 585
R568 B.n454 B.n249 585
R569 B.n249 B.n248 585
R570 B.n456 B.n455 585
R571 B.n457 B.n456 585
R572 B.n243 B.n242 585
R573 B.n244 B.n243 585
R574 B.n465 B.n464 585
R575 B.n464 B.n463 585
R576 B.n466 B.n241 585
R577 B.n241 B.n240 585
R578 B.n468 B.n467 585
R579 B.n469 B.n468 585
R580 B.n235 B.n234 585
R581 B.n236 B.n235 585
R582 B.n477 B.n476 585
R583 B.n476 B.n475 585
R584 B.n478 B.n233 585
R585 B.n233 B.n232 585
R586 B.n480 B.n479 585
R587 B.n481 B.n480 585
R588 B.n227 B.n226 585
R589 B.n228 B.n227 585
R590 B.n489 B.n488 585
R591 B.n488 B.n487 585
R592 B.n490 B.n225 585
R593 B.n225 B.n224 585
R594 B.n492 B.n491 585
R595 B.n493 B.n492 585
R596 B.n219 B.n218 585
R597 B.n220 B.n219 585
R598 B.n501 B.n500 585
R599 B.n500 B.n499 585
R600 B.n502 B.n217 585
R601 B.n217 B.n216 585
R602 B.n504 B.n503 585
R603 B.n505 B.n504 585
R604 B.n211 B.n210 585
R605 B.n212 B.n211 585
R606 B.n513 B.n512 585
R607 B.n512 B.n511 585
R608 B.n514 B.n209 585
R609 B.n209 B.n208 585
R610 B.n516 B.n515 585
R611 B.n517 B.n516 585
R612 B.n203 B.n202 585
R613 B.n204 B.n203 585
R614 B.n526 B.n525 585
R615 B.n525 B.n524 585
R616 B.n527 B.n201 585
R617 B.n201 B.n200 585
R618 B.n529 B.n528 585
R619 B.n530 B.n529 585
R620 B.n3 B.n0 585
R621 B.n4 B.n3 585
R622 B.n681 B.n1 585
R623 B.n682 B.n681 585
R624 B.n680 B.n679 585
R625 B.n680 B.n8 585
R626 B.n678 B.n9 585
R627 B.n12 B.n9 585
R628 B.n677 B.n676 585
R629 B.n676 B.n675 585
R630 B.n11 B.n10 585
R631 B.n674 B.n11 585
R632 B.n672 B.n671 585
R633 B.n673 B.n672 585
R634 B.n670 B.n17 585
R635 B.n17 B.n16 585
R636 B.n669 B.n668 585
R637 B.n668 B.n667 585
R638 B.n19 B.n18 585
R639 B.n666 B.n19 585
R640 B.n664 B.n663 585
R641 B.n665 B.n664 585
R642 B.n662 B.n24 585
R643 B.n24 B.n23 585
R644 B.n661 B.n660 585
R645 B.n660 B.n659 585
R646 B.n26 B.n25 585
R647 B.n658 B.n26 585
R648 B.n656 B.n655 585
R649 B.n657 B.n656 585
R650 B.n654 B.n31 585
R651 B.n31 B.n30 585
R652 B.n653 B.n652 585
R653 B.n652 B.n651 585
R654 B.n33 B.n32 585
R655 B.n650 B.n33 585
R656 B.n648 B.n647 585
R657 B.n649 B.n648 585
R658 B.n646 B.n38 585
R659 B.n38 B.n37 585
R660 B.n645 B.n644 585
R661 B.n644 B.n643 585
R662 B.n40 B.n39 585
R663 B.n642 B.n40 585
R664 B.n640 B.n639 585
R665 B.n641 B.n640 585
R666 B.n638 B.n45 585
R667 B.n45 B.n44 585
R668 B.n637 B.n636 585
R669 B.n636 B.n635 585
R670 B.n47 B.n46 585
R671 B.n634 B.n47 585
R672 B.n632 B.n631 585
R673 B.n633 B.n632 585
R674 B.n630 B.n52 585
R675 B.n52 B.n51 585
R676 B.n629 B.n628 585
R677 B.n628 B.n627 585
R678 B.n54 B.n53 585
R679 B.n626 B.n54 585
R680 B.n624 B.n623 585
R681 B.n625 B.n624 585
R682 B.n622 B.n59 585
R683 B.n59 B.n58 585
R684 B.n621 B.n620 585
R685 B.n620 B.n619 585
R686 B.n61 B.n60 585
R687 B.n618 B.n61 585
R688 B.n616 B.n615 585
R689 B.n617 B.n616 585
R690 B.n614 B.n65 585
R691 B.n68 B.n65 585
R692 B.n613 B.n612 585
R693 B.n612 B.n611 585
R694 B.n67 B.n66 585
R695 B.n610 B.n67 585
R696 B.n608 B.n607 585
R697 B.n609 B.n608 585
R698 B.n606 B.n73 585
R699 B.n73 B.n72 585
R700 B.n605 B.n604 585
R701 B.n604 B.n603 585
R702 B.n75 B.n74 585
R703 B.n602 B.n75 585
R704 B.n600 B.n599 585
R705 B.n601 B.n600 585
R706 B.n598 B.n80 585
R707 B.n80 B.n79 585
R708 B.n597 B.n596 585
R709 B.n596 B.n595 585
R710 B.n685 B.n684 585
R711 B.n683 B.n2 585
R712 B.n596 B.n82 526.135
R713 B.n593 B.n83 526.135
R714 B.n401 B.n284 526.135
R715 B.n403 B.n282 526.135
R716 B.n594 B.n105 256.663
R717 B.n594 B.n104 256.663
R718 B.n594 B.n103 256.663
R719 B.n594 B.n102 256.663
R720 B.n594 B.n101 256.663
R721 B.n594 B.n100 256.663
R722 B.n594 B.n99 256.663
R723 B.n594 B.n98 256.663
R724 B.n594 B.n97 256.663
R725 B.n594 B.n96 256.663
R726 B.n594 B.n95 256.663
R727 B.n594 B.n94 256.663
R728 B.n594 B.n93 256.663
R729 B.n594 B.n92 256.663
R730 B.n594 B.n91 256.663
R731 B.n594 B.n90 256.663
R732 B.n594 B.n89 256.663
R733 B.n594 B.n88 256.663
R734 B.n594 B.n87 256.663
R735 B.n594 B.n86 256.663
R736 B.n594 B.n85 256.663
R737 B.n594 B.n84 256.663
R738 B.n310 B.n283 256.663
R739 B.n313 B.n283 256.663
R740 B.n319 B.n283 256.663
R741 B.n321 B.n283 256.663
R742 B.n327 B.n283 256.663
R743 B.n329 B.n283 256.663
R744 B.n335 B.n283 256.663
R745 B.n337 B.n283 256.663
R746 B.n346 B.n283 256.663
R747 B.n348 B.n283 256.663
R748 B.n354 B.n283 256.663
R749 B.n356 B.n283 256.663
R750 B.n362 B.n283 256.663
R751 B.n364 B.n283 256.663
R752 B.n370 B.n283 256.663
R753 B.n372 B.n283 256.663
R754 B.n378 B.n283 256.663
R755 B.n380 B.n283 256.663
R756 B.n386 B.n283 256.663
R757 B.n388 B.n283 256.663
R758 B.n394 B.n283 256.663
R759 B.n396 B.n283 256.663
R760 B.n687 B.n686 256.663
R761 B.n109 B.t15 233.649
R762 B.n107 B.t8 233.649
R763 B.n293 B.t12 233.649
R764 B.n341 B.t4 233.649
R765 B.n107 B.t10 222.835
R766 B.n293 B.t14 222.835
R767 B.n109 B.t16 222.835
R768 B.n341 B.t7 222.835
R769 B.n402 B.n283 167.562
R770 B.n595 B.n594 167.562
R771 B.n114 B.n113 163.367
R772 B.n118 B.n117 163.367
R773 B.n122 B.n121 163.367
R774 B.n126 B.n125 163.367
R775 B.n130 B.n129 163.367
R776 B.n134 B.n133 163.367
R777 B.n138 B.n137 163.367
R778 B.n142 B.n141 163.367
R779 B.n146 B.n145 163.367
R780 B.n150 B.n149 163.367
R781 B.n154 B.n153 163.367
R782 B.n158 B.n157 163.367
R783 B.n162 B.n161 163.367
R784 B.n167 B.n166 163.367
R785 B.n171 B.n170 163.367
R786 B.n175 B.n174 163.367
R787 B.n179 B.n178 163.367
R788 B.n183 B.n182 163.367
R789 B.n187 B.n186 163.367
R790 B.n191 B.n190 163.367
R791 B.n195 B.n194 163.367
R792 B.n593 B.n106 163.367
R793 B.n401 B.n278 163.367
R794 B.n409 B.n278 163.367
R795 B.n409 B.n276 163.367
R796 B.n413 B.n276 163.367
R797 B.n413 B.n270 163.367
R798 B.n421 B.n270 163.367
R799 B.n421 B.n268 163.367
R800 B.n425 B.n268 163.367
R801 B.n425 B.n263 163.367
R802 B.n434 B.n263 163.367
R803 B.n434 B.n261 163.367
R804 B.n438 B.n261 163.367
R805 B.n438 B.n255 163.367
R806 B.n446 B.n255 163.367
R807 B.n446 B.n253 163.367
R808 B.n450 B.n253 163.367
R809 B.n450 B.n247 163.367
R810 B.n458 B.n247 163.367
R811 B.n458 B.n245 163.367
R812 B.n462 B.n245 163.367
R813 B.n462 B.n239 163.367
R814 B.n470 B.n239 163.367
R815 B.n470 B.n237 163.367
R816 B.n474 B.n237 163.367
R817 B.n474 B.n231 163.367
R818 B.n482 B.n231 163.367
R819 B.n482 B.n229 163.367
R820 B.n486 B.n229 163.367
R821 B.n486 B.n223 163.367
R822 B.n494 B.n223 163.367
R823 B.n494 B.n221 163.367
R824 B.n498 B.n221 163.367
R825 B.n498 B.n215 163.367
R826 B.n506 B.n215 163.367
R827 B.n506 B.n213 163.367
R828 B.n510 B.n213 163.367
R829 B.n510 B.n207 163.367
R830 B.n518 B.n207 163.367
R831 B.n518 B.n205 163.367
R832 B.n523 B.n205 163.367
R833 B.n523 B.n199 163.367
R834 B.n531 B.n199 163.367
R835 B.n532 B.n531 163.367
R836 B.n532 B.n5 163.367
R837 B.n6 B.n5 163.367
R838 B.n7 B.n6 163.367
R839 B.n538 B.n7 163.367
R840 B.n539 B.n538 163.367
R841 B.n539 B.n13 163.367
R842 B.n14 B.n13 163.367
R843 B.n15 B.n14 163.367
R844 B.n544 B.n15 163.367
R845 B.n544 B.n20 163.367
R846 B.n21 B.n20 163.367
R847 B.n22 B.n21 163.367
R848 B.n549 B.n22 163.367
R849 B.n549 B.n27 163.367
R850 B.n28 B.n27 163.367
R851 B.n29 B.n28 163.367
R852 B.n554 B.n29 163.367
R853 B.n554 B.n34 163.367
R854 B.n35 B.n34 163.367
R855 B.n36 B.n35 163.367
R856 B.n559 B.n36 163.367
R857 B.n559 B.n41 163.367
R858 B.n42 B.n41 163.367
R859 B.n43 B.n42 163.367
R860 B.n564 B.n43 163.367
R861 B.n564 B.n48 163.367
R862 B.n49 B.n48 163.367
R863 B.n50 B.n49 163.367
R864 B.n569 B.n50 163.367
R865 B.n569 B.n55 163.367
R866 B.n56 B.n55 163.367
R867 B.n57 B.n56 163.367
R868 B.n574 B.n57 163.367
R869 B.n574 B.n62 163.367
R870 B.n63 B.n62 163.367
R871 B.n64 B.n63 163.367
R872 B.n579 B.n64 163.367
R873 B.n579 B.n69 163.367
R874 B.n70 B.n69 163.367
R875 B.n71 B.n70 163.367
R876 B.n584 B.n71 163.367
R877 B.n584 B.n76 163.367
R878 B.n77 B.n76 163.367
R879 B.n78 B.n77 163.367
R880 B.n589 B.n78 163.367
R881 B.n589 B.n83 163.367
R882 B.n312 B.n311 163.367
R883 B.n314 B.n312 163.367
R884 B.n318 B.n307 163.367
R885 B.n322 B.n320 163.367
R886 B.n326 B.n305 163.367
R887 B.n330 B.n328 163.367
R888 B.n334 B.n303 163.367
R889 B.n338 B.n336 163.367
R890 B.n345 B.n301 163.367
R891 B.n349 B.n347 163.367
R892 B.n353 B.n299 163.367
R893 B.n357 B.n355 163.367
R894 B.n361 B.n297 163.367
R895 B.n365 B.n363 163.367
R896 B.n369 B.n292 163.367
R897 B.n373 B.n371 163.367
R898 B.n377 B.n290 163.367
R899 B.n381 B.n379 163.367
R900 B.n385 B.n288 163.367
R901 B.n389 B.n387 163.367
R902 B.n393 B.n286 163.367
R903 B.n397 B.n395 163.367
R904 B.n403 B.n280 163.367
R905 B.n407 B.n280 163.367
R906 B.n407 B.n274 163.367
R907 B.n415 B.n274 163.367
R908 B.n415 B.n272 163.367
R909 B.n419 B.n272 163.367
R910 B.n419 B.n266 163.367
R911 B.n428 B.n266 163.367
R912 B.n428 B.n264 163.367
R913 B.n432 B.n264 163.367
R914 B.n432 B.n259 163.367
R915 B.n440 B.n259 163.367
R916 B.n440 B.n257 163.367
R917 B.n444 B.n257 163.367
R918 B.n444 B.n251 163.367
R919 B.n452 B.n251 163.367
R920 B.n452 B.n249 163.367
R921 B.n456 B.n249 163.367
R922 B.n456 B.n243 163.367
R923 B.n464 B.n243 163.367
R924 B.n464 B.n241 163.367
R925 B.n468 B.n241 163.367
R926 B.n468 B.n235 163.367
R927 B.n476 B.n235 163.367
R928 B.n476 B.n233 163.367
R929 B.n480 B.n233 163.367
R930 B.n480 B.n227 163.367
R931 B.n488 B.n227 163.367
R932 B.n488 B.n225 163.367
R933 B.n492 B.n225 163.367
R934 B.n492 B.n219 163.367
R935 B.n500 B.n219 163.367
R936 B.n500 B.n217 163.367
R937 B.n504 B.n217 163.367
R938 B.n504 B.n211 163.367
R939 B.n512 B.n211 163.367
R940 B.n512 B.n209 163.367
R941 B.n516 B.n209 163.367
R942 B.n516 B.n203 163.367
R943 B.n525 B.n203 163.367
R944 B.n525 B.n201 163.367
R945 B.n529 B.n201 163.367
R946 B.n529 B.n3 163.367
R947 B.n685 B.n3 163.367
R948 B.n681 B.n2 163.367
R949 B.n681 B.n680 163.367
R950 B.n680 B.n9 163.367
R951 B.n676 B.n9 163.367
R952 B.n676 B.n11 163.367
R953 B.n672 B.n11 163.367
R954 B.n672 B.n17 163.367
R955 B.n668 B.n17 163.367
R956 B.n668 B.n19 163.367
R957 B.n664 B.n19 163.367
R958 B.n664 B.n24 163.367
R959 B.n660 B.n24 163.367
R960 B.n660 B.n26 163.367
R961 B.n656 B.n26 163.367
R962 B.n656 B.n31 163.367
R963 B.n652 B.n31 163.367
R964 B.n652 B.n33 163.367
R965 B.n648 B.n33 163.367
R966 B.n648 B.n38 163.367
R967 B.n644 B.n38 163.367
R968 B.n644 B.n40 163.367
R969 B.n640 B.n40 163.367
R970 B.n640 B.n45 163.367
R971 B.n636 B.n45 163.367
R972 B.n636 B.n47 163.367
R973 B.n632 B.n47 163.367
R974 B.n632 B.n52 163.367
R975 B.n628 B.n52 163.367
R976 B.n628 B.n54 163.367
R977 B.n624 B.n54 163.367
R978 B.n624 B.n59 163.367
R979 B.n620 B.n59 163.367
R980 B.n620 B.n61 163.367
R981 B.n616 B.n61 163.367
R982 B.n616 B.n65 163.367
R983 B.n612 B.n65 163.367
R984 B.n612 B.n67 163.367
R985 B.n608 B.n67 163.367
R986 B.n608 B.n73 163.367
R987 B.n604 B.n73 163.367
R988 B.n604 B.n75 163.367
R989 B.n600 B.n75 163.367
R990 B.n600 B.n80 163.367
R991 B.n596 B.n80 163.367
R992 B.n108 B.t11 142.351
R993 B.n294 B.t13 142.351
R994 B.n110 B.t17 142.351
R995 B.n342 B.t6 142.351
R996 B.n402 B.n279 81.9731
R997 B.n408 B.n279 81.9731
R998 B.n408 B.n275 81.9731
R999 B.n414 B.n275 81.9731
R1000 B.n414 B.n271 81.9731
R1001 B.n420 B.n271 81.9731
R1002 B.n420 B.n267 81.9731
R1003 B.n427 B.n267 81.9731
R1004 B.n427 B.n426 81.9731
R1005 B.n433 B.n260 81.9731
R1006 B.n439 B.n260 81.9731
R1007 B.n439 B.n256 81.9731
R1008 B.n445 B.n256 81.9731
R1009 B.n445 B.n252 81.9731
R1010 B.n451 B.n252 81.9731
R1011 B.n451 B.n248 81.9731
R1012 B.n457 B.n248 81.9731
R1013 B.n457 B.n244 81.9731
R1014 B.n463 B.n244 81.9731
R1015 B.n463 B.n240 81.9731
R1016 B.n469 B.n240 81.9731
R1017 B.n469 B.n236 81.9731
R1018 B.n475 B.n236 81.9731
R1019 B.n481 B.n232 81.9731
R1020 B.n481 B.n228 81.9731
R1021 B.n487 B.n228 81.9731
R1022 B.n487 B.n224 81.9731
R1023 B.n493 B.n224 81.9731
R1024 B.n493 B.n220 81.9731
R1025 B.n499 B.n220 81.9731
R1026 B.n499 B.n216 81.9731
R1027 B.n505 B.n216 81.9731
R1028 B.n505 B.n212 81.9731
R1029 B.n511 B.n212 81.9731
R1030 B.n517 B.n208 81.9731
R1031 B.n517 B.n204 81.9731
R1032 B.n524 B.n204 81.9731
R1033 B.n524 B.n200 81.9731
R1034 B.n530 B.n200 81.9731
R1035 B.n530 B.n4 81.9731
R1036 B.n684 B.n4 81.9731
R1037 B.n684 B.n683 81.9731
R1038 B.n683 B.n682 81.9731
R1039 B.n682 B.n8 81.9731
R1040 B.n12 B.n8 81.9731
R1041 B.n675 B.n12 81.9731
R1042 B.n675 B.n674 81.9731
R1043 B.n674 B.n673 81.9731
R1044 B.n673 B.n16 81.9731
R1045 B.n667 B.n666 81.9731
R1046 B.n666 B.n665 81.9731
R1047 B.n665 B.n23 81.9731
R1048 B.n659 B.n23 81.9731
R1049 B.n659 B.n658 81.9731
R1050 B.n658 B.n657 81.9731
R1051 B.n657 B.n30 81.9731
R1052 B.n651 B.n30 81.9731
R1053 B.n651 B.n650 81.9731
R1054 B.n650 B.n649 81.9731
R1055 B.n649 B.n37 81.9731
R1056 B.n643 B.n642 81.9731
R1057 B.n642 B.n641 81.9731
R1058 B.n641 B.n44 81.9731
R1059 B.n635 B.n44 81.9731
R1060 B.n635 B.n634 81.9731
R1061 B.n634 B.n633 81.9731
R1062 B.n633 B.n51 81.9731
R1063 B.n627 B.n51 81.9731
R1064 B.n627 B.n626 81.9731
R1065 B.n626 B.n625 81.9731
R1066 B.n625 B.n58 81.9731
R1067 B.n619 B.n58 81.9731
R1068 B.n619 B.n618 81.9731
R1069 B.n618 B.n617 81.9731
R1070 B.n611 B.n68 81.9731
R1071 B.n611 B.n610 81.9731
R1072 B.n610 B.n609 81.9731
R1073 B.n609 B.n72 81.9731
R1074 B.n603 B.n72 81.9731
R1075 B.n603 B.n602 81.9731
R1076 B.n602 B.n601 81.9731
R1077 B.n601 B.n79 81.9731
R1078 B.n595 B.n79 81.9731
R1079 B.n110 B.n109 80.4853
R1080 B.n108 B.n107 80.4853
R1081 B.n294 B.n293 80.4853
R1082 B.n342 B.n341 80.4853
R1083 B.n84 B.n82 71.676
R1084 B.n114 B.n85 71.676
R1085 B.n118 B.n86 71.676
R1086 B.n122 B.n87 71.676
R1087 B.n126 B.n88 71.676
R1088 B.n130 B.n89 71.676
R1089 B.n134 B.n90 71.676
R1090 B.n138 B.n91 71.676
R1091 B.n142 B.n92 71.676
R1092 B.n146 B.n93 71.676
R1093 B.n150 B.n94 71.676
R1094 B.n154 B.n95 71.676
R1095 B.n158 B.n96 71.676
R1096 B.n162 B.n97 71.676
R1097 B.n167 B.n98 71.676
R1098 B.n171 B.n99 71.676
R1099 B.n175 B.n100 71.676
R1100 B.n179 B.n101 71.676
R1101 B.n183 B.n102 71.676
R1102 B.n187 B.n103 71.676
R1103 B.n191 B.n104 71.676
R1104 B.n195 B.n105 71.676
R1105 B.n106 B.n105 71.676
R1106 B.n194 B.n104 71.676
R1107 B.n190 B.n103 71.676
R1108 B.n186 B.n102 71.676
R1109 B.n182 B.n101 71.676
R1110 B.n178 B.n100 71.676
R1111 B.n174 B.n99 71.676
R1112 B.n170 B.n98 71.676
R1113 B.n166 B.n97 71.676
R1114 B.n161 B.n96 71.676
R1115 B.n157 B.n95 71.676
R1116 B.n153 B.n94 71.676
R1117 B.n149 B.n93 71.676
R1118 B.n145 B.n92 71.676
R1119 B.n141 B.n91 71.676
R1120 B.n137 B.n90 71.676
R1121 B.n133 B.n89 71.676
R1122 B.n129 B.n88 71.676
R1123 B.n125 B.n87 71.676
R1124 B.n121 B.n86 71.676
R1125 B.n117 B.n85 71.676
R1126 B.n113 B.n84 71.676
R1127 B.n310 B.n282 71.676
R1128 B.n314 B.n313 71.676
R1129 B.n319 B.n318 71.676
R1130 B.n322 B.n321 71.676
R1131 B.n327 B.n326 71.676
R1132 B.n330 B.n329 71.676
R1133 B.n335 B.n334 71.676
R1134 B.n338 B.n337 71.676
R1135 B.n346 B.n345 71.676
R1136 B.n349 B.n348 71.676
R1137 B.n354 B.n353 71.676
R1138 B.n357 B.n356 71.676
R1139 B.n362 B.n361 71.676
R1140 B.n365 B.n364 71.676
R1141 B.n370 B.n369 71.676
R1142 B.n373 B.n372 71.676
R1143 B.n378 B.n377 71.676
R1144 B.n381 B.n380 71.676
R1145 B.n386 B.n385 71.676
R1146 B.n389 B.n388 71.676
R1147 B.n394 B.n393 71.676
R1148 B.n397 B.n396 71.676
R1149 B.n311 B.n310 71.676
R1150 B.n313 B.n307 71.676
R1151 B.n320 B.n319 71.676
R1152 B.n321 B.n305 71.676
R1153 B.n328 B.n327 71.676
R1154 B.n329 B.n303 71.676
R1155 B.n336 B.n335 71.676
R1156 B.n337 B.n301 71.676
R1157 B.n347 B.n346 71.676
R1158 B.n348 B.n299 71.676
R1159 B.n355 B.n354 71.676
R1160 B.n356 B.n297 71.676
R1161 B.n363 B.n362 71.676
R1162 B.n364 B.n292 71.676
R1163 B.n371 B.n370 71.676
R1164 B.n372 B.n290 71.676
R1165 B.n379 B.n378 71.676
R1166 B.n380 B.n288 71.676
R1167 B.n387 B.n386 71.676
R1168 B.n388 B.n286 71.676
R1169 B.n395 B.n394 71.676
R1170 B.n396 B.n284 71.676
R1171 B.n686 B.n685 71.676
R1172 B.n686 B.n2 71.676
R1173 B.n433 B.t5 67.5074
R1174 B.n617 B.t9 67.5074
R1175 B.n511 B.t1 65.0964
R1176 B.n667 B.t0 65.0964
R1177 B.n111 B.n110 59.5399
R1178 B.n164 B.n108 59.5399
R1179 B.n295 B.n294 59.5399
R1180 B.n343 B.n342 59.5399
R1181 B.n475 B.t3 48.2197
R1182 B.n643 B.t2 48.2197
R1183 B.n404 B.n281 34.1859
R1184 B.n400 B.n399 34.1859
R1185 B.n592 B.n591 34.1859
R1186 B.n597 B.n81 34.1859
R1187 B.t3 B.n232 33.7539
R1188 B.t2 B.n37 33.7539
R1189 B B.n687 18.0485
R1190 B.t1 B.n208 16.8772
R1191 B.t0 B.n16 16.8772
R1192 B.n426 B.t5 14.4663
R1193 B.n68 B.t9 14.4663
R1194 B.n405 B.n404 10.6151
R1195 B.n406 B.n405 10.6151
R1196 B.n406 B.n273 10.6151
R1197 B.n416 B.n273 10.6151
R1198 B.n417 B.n416 10.6151
R1199 B.n418 B.n417 10.6151
R1200 B.n418 B.n265 10.6151
R1201 B.n429 B.n265 10.6151
R1202 B.n430 B.n429 10.6151
R1203 B.n431 B.n430 10.6151
R1204 B.n431 B.n258 10.6151
R1205 B.n441 B.n258 10.6151
R1206 B.n442 B.n441 10.6151
R1207 B.n443 B.n442 10.6151
R1208 B.n443 B.n250 10.6151
R1209 B.n453 B.n250 10.6151
R1210 B.n454 B.n453 10.6151
R1211 B.n455 B.n454 10.6151
R1212 B.n455 B.n242 10.6151
R1213 B.n465 B.n242 10.6151
R1214 B.n466 B.n465 10.6151
R1215 B.n467 B.n466 10.6151
R1216 B.n467 B.n234 10.6151
R1217 B.n477 B.n234 10.6151
R1218 B.n478 B.n477 10.6151
R1219 B.n479 B.n478 10.6151
R1220 B.n479 B.n226 10.6151
R1221 B.n489 B.n226 10.6151
R1222 B.n490 B.n489 10.6151
R1223 B.n491 B.n490 10.6151
R1224 B.n491 B.n218 10.6151
R1225 B.n501 B.n218 10.6151
R1226 B.n502 B.n501 10.6151
R1227 B.n503 B.n502 10.6151
R1228 B.n503 B.n210 10.6151
R1229 B.n513 B.n210 10.6151
R1230 B.n514 B.n513 10.6151
R1231 B.n515 B.n514 10.6151
R1232 B.n515 B.n202 10.6151
R1233 B.n526 B.n202 10.6151
R1234 B.n527 B.n526 10.6151
R1235 B.n528 B.n527 10.6151
R1236 B.n528 B.n0 10.6151
R1237 B.n309 B.n281 10.6151
R1238 B.n309 B.n308 10.6151
R1239 B.n315 B.n308 10.6151
R1240 B.n316 B.n315 10.6151
R1241 B.n317 B.n316 10.6151
R1242 B.n317 B.n306 10.6151
R1243 B.n323 B.n306 10.6151
R1244 B.n324 B.n323 10.6151
R1245 B.n325 B.n324 10.6151
R1246 B.n325 B.n304 10.6151
R1247 B.n331 B.n304 10.6151
R1248 B.n332 B.n331 10.6151
R1249 B.n333 B.n332 10.6151
R1250 B.n333 B.n302 10.6151
R1251 B.n339 B.n302 10.6151
R1252 B.n340 B.n339 10.6151
R1253 B.n344 B.n340 10.6151
R1254 B.n350 B.n300 10.6151
R1255 B.n351 B.n350 10.6151
R1256 B.n352 B.n351 10.6151
R1257 B.n352 B.n298 10.6151
R1258 B.n358 B.n298 10.6151
R1259 B.n359 B.n358 10.6151
R1260 B.n360 B.n359 10.6151
R1261 B.n360 B.n296 10.6151
R1262 B.n367 B.n366 10.6151
R1263 B.n368 B.n367 10.6151
R1264 B.n368 B.n291 10.6151
R1265 B.n374 B.n291 10.6151
R1266 B.n375 B.n374 10.6151
R1267 B.n376 B.n375 10.6151
R1268 B.n376 B.n289 10.6151
R1269 B.n382 B.n289 10.6151
R1270 B.n383 B.n382 10.6151
R1271 B.n384 B.n383 10.6151
R1272 B.n384 B.n287 10.6151
R1273 B.n390 B.n287 10.6151
R1274 B.n391 B.n390 10.6151
R1275 B.n392 B.n391 10.6151
R1276 B.n392 B.n285 10.6151
R1277 B.n398 B.n285 10.6151
R1278 B.n399 B.n398 10.6151
R1279 B.n400 B.n277 10.6151
R1280 B.n410 B.n277 10.6151
R1281 B.n411 B.n410 10.6151
R1282 B.n412 B.n411 10.6151
R1283 B.n412 B.n269 10.6151
R1284 B.n422 B.n269 10.6151
R1285 B.n423 B.n422 10.6151
R1286 B.n424 B.n423 10.6151
R1287 B.n424 B.n262 10.6151
R1288 B.n435 B.n262 10.6151
R1289 B.n436 B.n435 10.6151
R1290 B.n437 B.n436 10.6151
R1291 B.n437 B.n254 10.6151
R1292 B.n447 B.n254 10.6151
R1293 B.n448 B.n447 10.6151
R1294 B.n449 B.n448 10.6151
R1295 B.n449 B.n246 10.6151
R1296 B.n459 B.n246 10.6151
R1297 B.n460 B.n459 10.6151
R1298 B.n461 B.n460 10.6151
R1299 B.n461 B.n238 10.6151
R1300 B.n471 B.n238 10.6151
R1301 B.n472 B.n471 10.6151
R1302 B.n473 B.n472 10.6151
R1303 B.n473 B.n230 10.6151
R1304 B.n483 B.n230 10.6151
R1305 B.n484 B.n483 10.6151
R1306 B.n485 B.n484 10.6151
R1307 B.n485 B.n222 10.6151
R1308 B.n495 B.n222 10.6151
R1309 B.n496 B.n495 10.6151
R1310 B.n497 B.n496 10.6151
R1311 B.n497 B.n214 10.6151
R1312 B.n507 B.n214 10.6151
R1313 B.n508 B.n507 10.6151
R1314 B.n509 B.n508 10.6151
R1315 B.n509 B.n206 10.6151
R1316 B.n519 B.n206 10.6151
R1317 B.n520 B.n519 10.6151
R1318 B.n522 B.n520 10.6151
R1319 B.n522 B.n521 10.6151
R1320 B.n521 B.n198 10.6151
R1321 B.n533 B.n198 10.6151
R1322 B.n534 B.n533 10.6151
R1323 B.n535 B.n534 10.6151
R1324 B.n536 B.n535 10.6151
R1325 B.n537 B.n536 10.6151
R1326 B.n540 B.n537 10.6151
R1327 B.n541 B.n540 10.6151
R1328 B.n542 B.n541 10.6151
R1329 B.n543 B.n542 10.6151
R1330 B.n545 B.n543 10.6151
R1331 B.n546 B.n545 10.6151
R1332 B.n547 B.n546 10.6151
R1333 B.n548 B.n547 10.6151
R1334 B.n550 B.n548 10.6151
R1335 B.n551 B.n550 10.6151
R1336 B.n552 B.n551 10.6151
R1337 B.n553 B.n552 10.6151
R1338 B.n555 B.n553 10.6151
R1339 B.n556 B.n555 10.6151
R1340 B.n557 B.n556 10.6151
R1341 B.n558 B.n557 10.6151
R1342 B.n560 B.n558 10.6151
R1343 B.n561 B.n560 10.6151
R1344 B.n562 B.n561 10.6151
R1345 B.n563 B.n562 10.6151
R1346 B.n565 B.n563 10.6151
R1347 B.n566 B.n565 10.6151
R1348 B.n567 B.n566 10.6151
R1349 B.n568 B.n567 10.6151
R1350 B.n570 B.n568 10.6151
R1351 B.n571 B.n570 10.6151
R1352 B.n572 B.n571 10.6151
R1353 B.n573 B.n572 10.6151
R1354 B.n575 B.n573 10.6151
R1355 B.n576 B.n575 10.6151
R1356 B.n577 B.n576 10.6151
R1357 B.n578 B.n577 10.6151
R1358 B.n580 B.n578 10.6151
R1359 B.n581 B.n580 10.6151
R1360 B.n582 B.n581 10.6151
R1361 B.n583 B.n582 10.6151
R1362 B.n585 B.n583 10.6151
R1363 B.n586 B.n585 10.6151
R1364 B.n587 B.n586 10.6151
R1365 B.n588 B.n587 10.6151
R1366 B.n590 B.n588 10.6151
R1367 B.n591 B.n590 10.6151
R1368 B.n679 B.n1 10.6151
R1369 B.n679 B.n678 10.6151
R1370 B.n678 B.n677 10.6151
R1371 B.n677 B.n10 10.6151
R1372 B.n671 B.n10 10.6151
R1373 B.n671 B.n670 10.6151
R1374 B.n670 B.n669 10.6151
R1375 B.n669 B.n18 10.6151
R1376 B.n663 B.n18 10.6151
R1377 B.n663 B.n662 10.6151
R1378 B.n662 B.n661 10.6151
R1379 B.n661 B.n25 10.6151
R1380 B.n655 B.n25 10.6151
R1381 B.n655 B.n654 10.6151
R1382 B.n654 B.n653 10.6151
R1383 B.n653 B.n32 10.6151
R1384 B.n647 B.n32 10.6151
R1385 B.n647 B.n646 10.6151
R1386 B.n646 B.n645 10.6151
R1387 B.n645 B.n39 10.6151
R1388 B.n639 B.n39 10.6151
R1389 B.n639 B.n638 10.6151
R1390 B.n638 B.n637 10.6151
R1391 B.n637 B.n46 10.6151
R1392 B.n631 B.n46 10.6151
R1393 B.n631 B.n630 10.6151
R1394 B.n630 B.n629 10.6151
R1395 B.n629 B.n53 10.6151
R1396 B.n623 B.n53 10.6151
R1397 B.n623 B.n622 10.6151
R1398 B.n622 B.n621 10.6151
R1399 B.n621 B.n60 10.6151
R1400 B.n615 B.n60 10.6151
R1401 B.n615 B.n614 10.6151
R1402 B.n614 B.n613 10.6151
R1403 B.n613 B.n66 10.6151
R1404 B.n607 B.n66 10.6151
R1405 B.n607 B.n606 10.6151
R1406 B.n606 B.n605 10.6151
R1407 B.n605 B.n74 10.6151
R1408 B.n599 B.n74 10.6151
R1409 B.n599 B.n598 10.6151
R1410 B.n598 B.n597 10.6151
R1411 B.n112 B.n81 10.6151
R1412 B.n115 B.n112 10.6151
R1413 B.n116 B.n115 10.6151
R1414 B.n119 B.n116 10.6151
R1415 B.n120 B.n119 10.6151
R1416 B.n123 B.n120 10.6151
R1417 B.n124 B.n123 10.6151
R1418 B.n127 B.n124 10.6151
R1419 B.n128 B.n127 10.6151
R1420 B.n131 B.n128 10.6151
R1421 B.n132 B.n131 10.6151
R1422 B.n135 B.n132 10.6151
R1423 B.n136 B.n135 10.6151
R1424 B.n139 B.n136 10.6151
R1425 B.n140 B.n139 10.6151
R1426 B.n143 B.n140 10.6151
R1427 B.n144 B.n143 10.6151
R1428 B.n148 B.n147 10.6151
R1429 B.n151 B.n148 10.6151
R1430 B.n152 B.n151 10.6151
R1431 B.n155 B.n152 10.6151
R1432 B.n156 B.n155 10.6151
R1433 B.n159 B.n156 10.6151
R1434 B.n160 B.n159 10.6151
R1435 B.n163 B.n160 10.6151
R1436 B.n168 B.n165 10.6151
R1437 B.n169 B.n168 10.6151
R1438 B.n172 B.n169 10.6151
R1439 B.n173 B.n172 10.6151
R1440 B.n176 B.n173 10.6151
R1441 B.n177 B.n176 10.6151
R1442 B.n180 B.n177 10.6151
R1443 B.n181 B.n180 10.6151
R1444 B.n184 B.n181 10.6151
R1445 B.n185 B.n184 10.6151
R1446 B.n188 B.n185 10.6151
R1447 B.n189 B.n188 10.6151
R1448 B.n192 B.n189 10.6151
R1449 B.n193 B.n192 10.6151
R1450 B.n196 B.n193 10.6151
R1451 B.n197 B.n196 10.6151
R1452 B.n592 B.n197 10.6151
R1453 B.n687 B.n0 8.11757
R1454 B.n687 B.n1 8.11757
R1455 B.n343 B.n300 6.5566
R1456 B.n296 B.n295 6.5566
R1457 B.n147 B.n111 6.5566
R1458 B.n164 B.n163 6.5566
R1459 B.n344 B.n343 4.05904
R1460 B.n366 B.n295 4.05904
R1461 B.n144 B.n111 4.05904
R1462 B.n165 B.n164 4.05904
R1463 VP.n21 VP.n20 161.3
R1464 VP.n19 VP.n1 161.3
R1465 VP.n18 VP.n17 161.3
R1466 VP.n16 VP.n2 161.3
R1467 VP.n15 VP.n14 161.3
R1468 VP.n13 VP.n3 161.3
R1469 VP.n12 VP.n11 161.3
R1470 VP.n10 VP.n4 161.3
R1471 VP.n9 VP.n8 161.3
R1472 VP.n7 VP.n6 86.3974
R1473 VP.n22 VP.n0 86.3974
R1474 VP.n5 VP.t3 58.3543
R1475 VP.n5 VP.t1 56.9995
R1476 VP.n6 VP.n5 45.7866
R1477 VP.n14 VP.n13 40.4934
R1478 VP.n14 VP.n2 40.4934
R1479 VP.n8 VP.n4 24.4675
R1480 VP.n12 VP.n4 24.4675
R1481 VP.n13 VP.n12 24.4675
R1482 VP.n18 VP.n2 24.4675
R1483 VP.n19 VP.n18 24.4675
R1484 VP.n20 VP.n19 24.4675
R1485 VP.n7 VP.t0 24.2898
R1486 VP.n0 VP.t2 24.2898
R1487 VP.n8 VP.n7 3.67055
R1488 VP.n20 VP.n0 3.67055
R1489 VP.n9 VP.n6 0.354971
R1490 VP.n22 VP.n21 0.354971
R1491 VP VP.n22 0.26696
R1492 VP.n10 VP.n9 0.189894
R1493 VP.n11 VP.n10 0.189894
R1494 VP.n11 VP.n3 0.189894
R1495 VP.n15 VP.n3 0.189894
R1496 VP.n16 VP.n15 0.189894
R1497 VP.n17 VP.n16 0.189894
R1498 VP.n17 VP.n1 0.189894
R1499 VP.n21 VP.n1 0.189894
R1500 VDD1 VDD1.n1 111.95
R1501 VDD1 VDD1.n0 73.7161
R1502 VDD1.n0 VDD1.t0 5.14336
R1503 VDD1.n0 VDD1.t2 5.14336
R1504 VDD1.n1 VDD1.t3 5.14336
R1505 VDD1.n1 VDD1.t1 5.14336
C0 VP VTAIL 2.53758f
C1 VP VDD2 0.476682f
C2 VDD1 VTAIL 4.06202f
C3 VP VN 5.5665f
C4 VDD2 VDD1 1.32288f
C5 VDD1 VN 0.154313f
C6 VDD2 VTAIL 4.1244f
C7 VTAIL VN 2.52348f
C8 VDD2 VN 1.84888f
C9 VP VDD1 2.16958f
C10 VDD2 B 3.725367f
C11 VDD1 B 7.8311f
C12 VTAIL B 5.421374f
C13 VN B 12.18005f
C14 VP B 10.760204f
C15 VDD1.t0 B 0.092356f
C16 VDD1.t2 B 0.092356f
C17 VDD1.n0 B 0.721996f
C18 VDD1.t3 B 0.092356f
C19 VDD1.t1 B 0.092356f
C20 VDD1.n1 B 1.20642f
C21 VP.t2 B 1.01753f
C22 VP.n0 B 0.499289f
C23 VP.n1 B 0.027028f
C24 VP.n2 B 0.053718f
C25 VP.n3 B 0.027028f
C26 VP.n4 B 0.050373f
C27 VP.t3 B 1.37977f
C28 VP.t1 B 1.36531f
C29 VP.n5 B 2.33839f
C30 VP.n6 B 1.3772f
C31 VP.t0 B 1.01753f
C32 VP.n7 B 0.499289f
C33 VP.n8 B 0.029233f
C34 VP.n9 B 0.043623f
C35 VP.n10 B 0.027028f
C36 VP.n11 B 0.027028f
C37 VP.n12 B 0.050373f
C38 VP.n13 B 0.053718f
C39 VP.n14 B 0.02185f
C40 VP.n15 B 0.027028f
C41 VP.n16 B 0.027028f
C42 VP.n17 B 0.027028f
C43 VP.n18 B 0.050373f
C44 VP.n19 B 0.050373f
C45 VP.n20 B 0.029233f
C46 VP.n21 B 0.043623f
C47 VP.n22 B 0.082689f
C48 VTAIL.n0 B 0.032014f
C49 VTAIL.n1 B 0.024046f
C50 VTAIL.n2 B 0.012921f
C51 VTAIL.n3 B 0.030541f
C52 VTAIL.n4 B 0.013681f
C53 VTAIL.n5 B 0.091362f
C54 VTAIL.t5 B 0.050454f
C55 VTAIL.n6 B 0.022906f
C56 VTAIL.n7 B 0.017975f
C57 VTAIL.n8 B 0.012921f
C58 VTAIL.n9 B 0.332996f
C59 VTAIL.n10 B 0.024046f
C60 VTAIL.n11 B 0.012921f
C61 VTAIL.n12 B 0.013681f
C62 VTAIL.n13 B 0.030541f
C63 VTAIL.n14 B 0.06296f
C64 VTAIL.n15 B 0.013681f
C65 VTAIL.n16 B 0.012921f
C66 VTAIL.n17 B 0.055909f
C67 VTAIL.n18 B 0.034914f
C68 VTAIL.n19 B 0.20023f
C69 VTAIL.n20 B 0.032014f
C70 VTAIL.n21 B 0.024046f
C71 VTAIL.n22 B 0.012921f
C72 VTAIL.n23 B 0.030541f
C73 VTAIL.n24 B 0.013681f
C74 VTAIL.n25 B 0.091362f
C75 VTAIL.t1 B 0.050454f
C76 VTAIL.n26 B 0.022906f
C77 VTAIL.n27 B 0.017975f
C78 VTAIL.n28 B 0.012921f
C79 VTAIL.n29 B 0.332996f
C80 VTAIL.n30 B 0.024046f
C81 VTAIL.n31 B 0.012921f
C82 VTAIL.n32 B 0.013681f
C83 VTAIL.n33 B 0.030541f
C84 VTAIL.n34 B 0.06296f
C85 VTAIL.n35 B 0.013681f
C86 VTAIL.n36 B 0.012921f
C87 VTAIL.n37 B 0.055909f
C88 VTAIL.n38 B 0.034914f
C89 VTAIL.n39 B 0.334319f
C90 VTAIL.n40 B 0.032014f
C91 VTAIL.n41 B 0.024046f
C92 VTAIL.n42 B 0.012921f
C93 VTAIL.n43 B 0.030541f
C94 VTAIL.n44 B 0.013681f
C95 VTAIL.n45 B 0.091362f
C96 VTAIL.t7 B 0.050454f
C97 VTAIL.n46 B 0.022906f
C98 VTAIL.n47 B 0.017975f
C99 VTAIL.n48 B 0.012921f
C100 VTAIL.n49 B 0.332996f
C101 VTAIL.n50 B 0.024046f
C102 VTAIL.n51 B 0.012921f
C103 VTAIL.n52 B 0.013681f
C104 VTAIL.n53 B 0.030541f
C105 VTAIL.n54 B 0.06296f
C106 VTAIL.n55 B 0.013681f
C107 VTAIL.n56 B 0.012921f
C108 VTAIL.n57 B 0.055909f
C109 VTAIL.n58 B 0.034914f
C110 VTAIL.n59 B 1.1589f
C111 VTAIL.n60 B 0.032014f
C112 VTAIL.n61 B 0.024046f
C113 VTAIL.n62 B 0.012921f
C114 VTAIL.n63 B 0.030541f
C115 VTAIL.n64 B 0.013681f
C116 VTAIL.n65 B 0.091362f
C117 VTAIL.t4 B 0.050454f
C118 VTAIL.n66 B 0.022906f
C119 VTAIL.n67 B 0.017975f
C120 VTAIL.n68 B 0.012921f
C121 VTAIL.n69 B 0.332996f
C122 VTAIL.n70 B 0.024046f
C123 VTAIL.n71 B 0.012921f
C124 VTAIL.n72 B 0.013681f
C125 VTAIL.n73 B 0.030541f
C126 VTAIL.n74 B 0.06296f
C127 VTAIL.n75 B 0.013681f
C128 VTAIL.n76 B 0.012921f
C129 VTAIL.n77 B 0.055909f
C130 VTAIL.n78 B 0.034914f
C131 VTAIL.n79 B 1.1589f
C132 VTAIL.n80 B 0.032014f
C133 VTAIL.n81 B 0.024046f
C134 VTAIL.n82 B 0.012921f
C135 VTAIL.n83 B 0.030541f
C136 VTAIL.n84 B 0.013681f
C137 VTAIL.n85 B 0.091362f
C138 VTAIL.t2 B 0.050454f
C139 VTAIL.n86 B 0.022906f
C140 VTAIL.n87 B 0.017975f
C141 VTAIL.n88 B 0.012921f
C142 VTAIL.n89 B 0.332996f
C143 VTAIL.n90 B 0.024046f
C144 VTAIL.n91 B 0.012921f
C145 VTAIL.n92 B 0.013681f
C146 VTAIL.n93 B 0.030541f
C147 VTAIL.n94 B 0.06296f
C148 VTAIL.n95 B 0.013681f
C149 VTAIL.n96 B 0.012921f
C150 VTAIL.n97 B 0.055909f
C151 VTAIL.n98 B 0.034914f
C152 VTAIL.n99 B 0.334319f
C153 VTAIL.n100 B 0.032014f
C154 VTAIL.n101 B 0.024046f
C155 VTAIL.n102 B 0.012921f
C156 VTAIL.n103 B 0.030541f
C157 VTAIL.n104 B 0.013681f
C158 VTAIL.n105 B 0.091362f
C159 VTAIL.t0 B 0.050454f
C160 VTAIL.n106 B 0.022906f
C161 VTAIL.n107 B 0.017975f
C162 VTAIL.n108 B 0.012921f
C163 VTAIL.n109 B 0.332996f
C164 VTAIL.n110 B 0.024046f
C165 VTAIL.n111 B 0.012921f
C166 VTAIL.n112 B 0.013681f
C167 VTAIL.n113 B 0.030541f
C168 VTAIL.n114 B 0.06296f
C169 VTAIL.n115 B 0.013681f
C170 VTAIL.n116 B 0.012921f
C171 VTAIL.n117 B 0.055909f
C172 VTAIL.n118 B 0.034914f
C173 VTAIL.n119 B 0.334319f
C174 VTAIL.n120 B 0.032014f
C175 VTAIL.n121 B 0.024046f
C176 VTAIL.n122 B 0.012921f
C177 VTAIL.n123 B 0.030541f
C178 VTAIL.n124 B 0.013681f
C179 VTAIL.n125 B 0.091362f
C180 VTAIL.t6 B 0.050454f
C181 VTAIL.n126 B 0.022906f
C182 VTAIL.n127 B 0.017975f
C183 VTAIL.n128 B 0.012921f
C184 VTAIL.n129 B 0.332996f
C185 VTAIL.n130 B 0.024046f
C186 VTAIL.n131 B 0.012921f
C187 VTAIL.n132 B 0.013681f
C188 VTAIL.n133 B 0.030541f
C189 VTAIL.n134 B 0.06296f
C190 VTAIL.n135 B 0.013681f
C191 VTAIL.n136 B 0.012921f
C192 VTAIL.n137 B 0.055909f
C193 VTAIL.n138 B 0.034914f
C194 VTAIL.n139 B 1.1589f
C195 VTAIL.n140 B 0.032014f
C196 VTAIL.n141 B 0.024046f
C197 VTAIL.n142 B 0.012921f
C198 VTAIL.n143 B 0.030541f
C199 VTAIL.n144 B 0.013681f
C200 VTAIL.n145 B 0.091362f
C201 VTAIL.t3 B 0.050454f
C202 VTAIL.n146 B 0.022906f
C203 VTAIL.n147 B 0.017975f
C204 VTAIL.n148 B 0.012921f
C205 VTAIL.n149 B 0.332996f
C206 VTAIL.n150 B 0.024046f
C207 VTAIL.n151 B 0.012921f
C208 VTAIL.n152 B 0.013681f
C209 VTAIL.n153 B 0.030541f
C210 VTAIL.n154 B 0.06296f
C211 VTAIL.n155 B 0.013681f
C212 VTAIL.n156 B 0.012921f
C213 VTAIL.n157 B 0.055909f
C214 VTAIL.n158 B 0.034914f
C215 VTAIL.n159 B 1.01579f
C216 VDD2.t2 B 0.061194f
C217 VDD2.t3 B 0.061194f
C218 VDD2.n0 B 0.782834f
C219 VDD2.t0 B 0.061194f
C220 VDD2.t1 B 0.061194f
C221 VDD2.n1 B 0.478069f
C222 VDD2.n2 B 2.35813f
C223 VN.t2 B 1.06974f
C224 VN.t0 B 1.08107f
C225 VN.n0 B 0.655841f
C226 VN.t1 B 1.06974f
C227 VN.t3 B 1.08107f
C228 VN.n1 B 1.84107f
.ends

