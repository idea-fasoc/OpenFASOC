* NGSPICE file created from diff_pair_sample_1433.ext - technology: sky130A

.subckt diff_pair_sample_1433 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=1.8282 ps=11.41 w=11.08 l=1.18
X1 VDD1.t8 VP.t1 VTAIL.t16 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=4.3212 ps=22.94 w=11.08 l=1.18
X2 VDD1.t7 VP.t2 VTAIL.t14 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=1.8282 ps=11.41 w=11.08 l=1.18
X3 B.t11 B.t9 B.t10 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=0 ps=0 w=11.08 l=1.18
X4 VTAIL.t9 VP.t3 VDD1.t6 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X5 B.t8 B.t6 B.t7 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=0 ps=0 w=11.08 l=1.18
X6 VTAIL.t18 VP.t4 VDD1.t5 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X7 VTAIL.t10 VP.t5 VDD1.t4 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X8 B.t5 B.t3 B.t4 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=0 ps=0 w=11.08 l=1.18
X9 VDD2.t9 VN.t0 VTAIL.t3 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=1.8282 ps=11.41 w=11.08 l=1.18
X10 VDD1.t3 VP.t6 VTAIL.t11 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X11 VDD2.t8 VN.t1 VTAIL.t7 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X12 VDD2.t7 VN.t2 VTAIL.t8 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=4.3212 ps=22.94 w=11.08 l=1.18
X13 VTAIL.t12 VP.t7 VDD1.t2 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X14 VDD2.t6 VN.t3 VTAIL.t4 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X15 VDD2.t5 VN.t4 VTAIL.t0 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=1.8282 ps=11.41 w=11.08 l=1.18
X16 B.t2 B.t0 B.t1 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=4.3212 pd=22.94 as=0 ps=0 w=11.08 l=1.18
X17 VDD1.t1 VP.t8 VTAIL.t17 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=4.3212 ps=22.94 w=11.08 l=1.18
X18 VTAIL.t6 VN.t5 VDD2.t4 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X19 VTAIL.t2 VN.t6 VDD2.t3 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X20 VDD1.t0 VP.t9 VTAIL.t13 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X21 VTAIL.t19 VN.t7 VDD2.t2 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X22 VTAIL.t1 VN.t8 VDD2.t1 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=1.8282 ps=11.41 w=11.08 l=1.18
X23 VDD2.t0 VN.t9 VTAIL.t5 w_n2782_n3184# sky130_fd_pr__pfet_01v8 ad=1.8282 pd=11.41 as=4.3212 ps=22.94 w=11.08 l=1.18
R0 VP.n14 VP.t0 257.159
R1 VP.n7 VP.t2 226.296
R2 VP.n5 VP.t4 226.296
R3 VP.n3 VP.t6 226.296
R4 VP.n46 VP.t3 226.296
R5 VP.n53 VP.t1 226.296
R6 VP.n30 VP.t8 226.296
R7 VP.n23 VP.t5 226.296
R8 VP.n11 VP.t9 226.296
R9 VP.n13 VP.t7 226.296
R10 VP.n32 VP.n7 172.613
R11 VP.n54 VP.n53 172.613
R12 VP.n31 VP.n30 172.613
R13 VP.n16 VP.n15 161.3
R14 VP.n17 VP.n12 161.3
R15 VP.n19 VP.n18 161.3
R16 VP.n21 VP.n20 161.3
R17 VP.n22 VP.n10 161.3
R18 VP.n25 VP.n24 161.3
R19 VP.n26 VP.n9 161.3
R20 VP.n28 VP.n27 161.3
R21 VP.n29 VP.n8 161.3
R22 VP.n52 VP.n0 161.3
R23 VP.n51 VP.n50 161.3
R24 VP.n49 VP.n1 161.3
R25 VP.n48 VP.n47 161.3
R26 VP.n45 VP.n2 161.3
R27 VP.n44 VP.n43 161.3
R28 VP.n42 VP.n41 161.3
R29 VP.n40 VP.n4 161.3
R30 VP.n39 VP.n38 161.3
R31 VP.n37 VP.n36 161.3
R32 VP.n35 VP.n6 161.3
R33 VP.n34 VP.n33 161.3
R34 VP.n14 VP.n13 50.8823
R35 VP.n32 VP.n31 44.5952
R36 VP.n35 VP.n34 42.0302
R37 VP.n52 VP.n51 42.0302
R38 VP.n29 VP.n28 42.0302
R39 VP.n40 VP.n39 41.0614
R40 VP.n47 VP.n45 41.0614
R41 VP.n24 VP.n22 41.0614
R42 VP.n17 VP.n16 41.0614
R43 VP.n41 VP.n40 40.0926
R44 VP.n45 VP.n44 40.0926
R45 VP.n22 VP.n21 40.0926
R46 VP.n18 VP.n17 40.0926
R47 VP.n36 VP.n35 39.1239
R48 VP.n51 VP.n1 39.1239
R49 VP.n28 VP.n9 39.1239
R50 VP.n15 VP.n14 26.821
R51 VP.n34 VP.n7 13.2801
R52 VP.n53 VP.n52 13.2801
R53 VP.n30 VP.n29 13.2801
R54 VP.n39 VP.n5 12.7883
R55 VP.n47 VP.n46 12.7883
R56 VP.n24 VP.n23 12.7883
R57 VP.n16 VP.n13 12.7883
R58 VP.n41 VP.n3 12.2964
R59 VP.n44 VP.n3 12.2964
R60 VP.n18 VP.n11 12.2964
R61 VP.n21 VP.n11 12.2964
R62 VP.n36 VP.n5 11.8046
R63 VP.n46 VP.n1 11.8046
R64 VP.n23 VP.n9 11.8046
R65 VP.n15 VP.n12 0.189894
R66 VP.n19 VP.n12 0.189894
R67 VP.n20 VP.n19 0.189894
R68 VP.n20 VP.n10 0.189894
R69 VP.n25 VP.n10 0.189894
R70 VP.n26 VP.n25 0.189894
R71 VP.n27 VP.n26 0.189894
R72 VP.n27 VP.n8 0.189894
R73 VP.n31 VP.n8 0.189894
R74 VP.n33 VP.n32 0.189894
R75 VP.n33 VP.n6 0.189894
R76 VP.n37 VP.n6 0.189894
R77 VP.n38 VP.n37 0.189894
R78 VP.n38 VP.n4 0.189894
R79 VP.n42 VP.n4 0.189894
R80 VP.n43 VP.n42 0.189894
R81 VP.n43 VP.n2 0.189894
R82 VP.n48 VP.n2 0.189894
R83 VP.n49 VP.n48 0.189894
R84 VP.n50 VP.n49 0.189894
R85 VP.n50 VP.n0 0.189894
R86 VP.n54 VP.n0 0.189894
R87 VP VP.n54 0.0516364
R88 VTAIL.n11 VTAIL.t8 62.3356
R89 VTAIL.n17 VTAIL.t5 62.3355
R90 VTAIL.n2 VTAIL.t16 62.3355
R91 VTAIL.n16 VTAIL.t17 62.3355
R92 VTAIL.n15 VTAIL.n14 59.402
R93 VTAIL.n13 VTAIL.n12 59.402
R94 VTAIL.n10 VTAIL.n9 59.402
R95 VTAIL.n8 VTAIL.n7 59.402
R96 VTAIL.n19 VTAIL.n18 59.4018
R97 VTAIL.n1 VTAIL.n0 59.4018
R98 VTAIL.n4 VTAIL.n3 59.4018
R99 VTAIL.n6 VTAIL.n5 59.4018
R100 VTAIL.n8 VTAIL.n6 24.5221
R101 VTAIL.n17 VTAIL.n16 23.2203
R102 VTAIL.n18 VTAIL.t4 2.93416
R103 VTAIL.n18 VTAIL.t6 2.93416
R104 VTAIL.n0 VTAIL.t0 2.93416
R105 VTAIL.n0 VTAIL.t2 2.93416
R106 VTAIL.n3 VTAIL.t11 2.93416
R107 VTAIL.n3 VTAIL.t9 2.93416
R108 VTAIL.n5 VTAIL.t14 2.93416
R109 VTAIL.n5 VTAIL.t18 2.93416
R110 VTAIL.n14 VTAIL.t13 2.93416
R111 VTAIL.n14 VTAIL.t10 2.93416
R112 VTAIL.n12 VTAIL.t15 2.93416
R113 VTAIL.n12 VTAIL.t12 2.93416
R114 VTAIL.n9 VTAIL.t7 2.93416
R115 VTAIL.n9 VTAIL.t19 2.93416
R116 VTAIL.n7 VTAIL.t3 2.93416
R117 VTAIL.n7 VTAIL.t1 2.93416
R118 VTAIL.n10 VTAIL.n8 1.30222
R119 VTAIL.n11 VTAIL.n10 1.30222
R120 VTAIL.n15 VTAIL.n13 1.30222
R121 VTAIL.n16 VTAIL.n15 1.30222
R122 VTAIL.n6 VTAIL.n4 1.30222
R123 VTAIL.n4 VTAIL.n2 1.30222
R124 VTAIL.n19 VTAIL.n17 1.30222
R125 VTAIL.n13 VTAIL.n11 1.12119
R126 VTAIL.n2 VTAIL.n1 1.12119
R127 VTAIL VTAIL.n1 1.03498
R128 VTAIL VTAIL.n19 0.267741
R129 VDD1.n1 VDD1.t9 80.3161
R130 VDD1.n3 VDD1.t7 80.316
R131 VDD1.n5 VDD1.n4 77.0015
R132 VDD1.n1 VDD1.n0 76.0808
R133 VDD1.n7 VDD1.n6 76.0806
R134 VDD1.n3 VDD1.n2 76.0806
R135 VDD1.n7 VDD1.n5 40.6841
R136 VDD1.n6 VDD1.t4 2.93416
R137 VDD1.n6 VDD1.t1 2.93416
R138 VDD1.n0 VDD1.t2 2.93416
R139 VDD1.n0 VDD1.t0 2.93416
R140 VDD1.n4 VDD1.t6 2.93416
R141 VDD1.n4 VDD1.t8 2.93416
R142 VDD1.n2 VDD1.t5 2.93416
R143 VDD1.n2 VDD1.t3 2.93416
R144 VDD1 VDD1.n7 0.918603
R145 VDD1 VDD1.n1 0.384121
R146 VDD1.n5 VDD1.n3 0.270585
R147 B.n348 B.n347 585
R148 B.n346 B.n103 585
R149 B.n345 B.n344 585
R150 B.n343 B.n104 585
R151 B.n342 B.n341 585
R152 B.n340 B.n105 585
R153 B.n339 B.n338 585
R154 B.n337 B.n106 585
R155 B.n336 B.n335 585
R156 B.n334 B.n107 585
R157 B.n333 B.n332 585
R158 B.n331 B.n108 585
R159 B.n330 B.n329 585
R160 B.n328 B.n109 585
R161 B.n327 B.n326 585
R162 B.n325 B.n110 585
R163 B.n324 B.n323 585
R164 B.n322 B.n111 585
R165 B.n321 B.n320 585
R166 B.n319 B.n112 585
R167 B.n318 B.n317 585
R168 B.n316 B.n113 585
R169 B.n315 B.n314 585
R170 B.n313 B.n114 585
R171 B.n312 B.n311 585
R172 B.n310 B.n115 585
R173 B.n309 B.n308 585
R174 B.n307 B.n116 585
R175 B.n306 B.n305 585
R176 B.n304 B.n117 585
R177 B.n303 B.n302 585
R178 B.n301 B.n118 585
R179 B.n300 B.n299 585
R180 B.n298 B.n119 585
R181 B.n297 B.n296 585
R182 B.n295 B.n120 585
R183 B.n294 B.n293 585
R184 B.n292 B.n121 585
R185 B.n291 B.n290 585
R186 B.n288 B.n122 585
R187 B.n287 B.n286 585
R188 B.n285 B.n125 585
R189 B.n284 B.n283 585
R190 B.n282 B.n126 585
R191 B.n281 B.n280 585
R192 B.n279 B.n127 585
R193 B.n278 B.n277 585
R194 B.n276 B.n128 585
R195 B.n274 B.n273 585
R196 B.n272 B.n131 585
R197 B.n271 B.n270 585
R198 B.n269 B.n132 585
R199 B.n268 B.n267 585
R200 B.n266 B.n133 585
R201 B.n265 B.n264 585
R202 B.n263 B.n134 585
R203 B.n262 B.n261 585
R204 B.n260 B.n135 585
R205 B.n259 B.n258 585
R206 B.n257 B.n136 585
R207 B.n256 B.n255 585
R208 B.n254 B.n137 585
R209 B.n253 B.n252 585
R210 B.n251 B.n138 585
R211 B.n250 B.n249 585
R212 B.n248 B.n139 585
R213 B.n247 B.n246 585
R214 B.n245 B.n140 585
R215 B.n244 B.n243 585
R216 B.n242 B.n141 585
R217 B.n241 B.n240 585
R218 B.n239 B.n142 585
R219 B.n238 B.n237 585
R220 B.n236 B.n143 585
R221 B.n235 B.n234 585
R222 B.n233 B.n144 585
R223 B.n232 B.n231 585
R224 B.n230 B.n145 585
R225 B.n229 B.n228 585
R226 B.n227 B.n146 585
R227 B.n226 B.n225 585
R228 B.n224 B.n147 585
R229 B.n223 B.n222 585
R230 B.n221 B.n148 585
R231 B.n220 B.n219 585
R232 B.n218 B.n149 585
R233 B.n217 B.n216 585
R234 B.n349 B.n102 585
R235 B.n351 B.n350 585
R236 B.n352 B.n101 585
R237 B.n354 B.n353 585
R238 B.n355 B.n100 585
R239 B.n357 B.n356 585
R240 B.n358 B.n99 585
R241 B.n360 B.n359 585
R242 B.n361 B.n98 585
R243 B.n363 B.n362 585
R244 B.n364 B.n97 585
R245 B.n366 B.n365 585
R246 B.n367 B.n96 585
R247 B.n369 B.n368 585
R248 B.n370 B.n95 585
R249 B.n372 B.n371 585
R250 B.n373 B.n94 585
R251 B.n375 B.n374 585
R252 B.n376 B.n93 585
R253 B.n378 B.n377 585
R254 B.n379 B.n92 585
R255 B.n381 B.n380 585
R256 B.n382 B.n91 585
R257 B.n384 B.n383 585
R258 B.n385 B.n90 585
R259 B.n387 B.n386 585
R260 B.n388 B.n89 585
R261 B.n390 B.n389 585
R262 B.n391 B.n88 585
R263 B.n393 B.n392 585
R264 B.n394 B.n87 585
R265 B.n396 B.n395 585
R266 B.n397 B.n86 585
R267 B.n399 B.n398 585
R268 B.n400 B.n85 585
R269 B.n402 B.n401 585
R270 B.n403 B.n84 585
R271 B.n405 B.n404 585
R272 B.n406 B.n83 585
R273 B.n408 B.n407 585
R274 B.n409 B.n82 585
R275 B.n411 B.n410 585
R276 B.n412 B.n81 585
R277 B.n414 B.n413 585
R278 B.n415 B.n80 585
R279 B.n417 B.n416 585
R280 B.n418 B.n79 585
R281 B.n420 B.n419 585
R282 B.n421 B.n78 585
R283 B.n423 B.n422 585
R284 B.n424 B.n77 585
R285 B.n426 B.n425 585
R286 B.n427 B.n76 585
R287 B.n429 B.n428 585
R288 B.n430 B.n75 585
R289 B.n432 B.n431 585
R290 B.n433 B.n74 585
R291 B.n435 B.n434 585
R292 B.n436 B.n73 585
R293 B.n438 B.n437 585
R294 B.n439 B.n72 585
R295 B.n441 B.n440 585
R296 B.n442 B.n71 585
R297 B.n444 B.n443 585
R298 B.n445 B.n70 585
R299 B.n447 B.n446 585
R300 B.n448 B.n69 585
R301 B.n450 B.n449 585
R302 B.n451 B.n68 585
R303 B.n453 B.n452 585
R304 B.n584 B.n19 585
R305 B.n583 B.n582 585
R306 B.n581 B.n20 585
R307 B.n580 B.n579 585
R308 B.n578 B.n21 585
R309 B.n577 B.n576 585
R310 B.n575 B.n22 585
R311 B.n574 B.n573 585
R312 B.n572 B.n23 585
R313 B.n571 B.n570 585
R314 B.n569 B.n24 585
R315 B.n568 B.n567 585
R316 B.n566 B.n25 585
R317 B.n565 B.n564 585
R318 B.n563 B.n26 585
R319 B.n562 B.n561 585
R320 B.n560 B.n27 585
R321 B.n559 B.n558 585
R322 B.n557 B.n28 585
R323 B.n556 B.n555 585
R324 B.n554 B.n29 585
R325 B.n553 B.n552 585
R326 B.n551 B.n30 585
R327 B.n550 B.n549 585
R328 B.n548 B.n31 585
R329 B.n547 B.n546 585
R330 B.n545 B.n32 585
R331 B.n544 B.n543 585
R332 B.n542 B.n33 585
R333 B.n541 B.n540 585
R334 B.n539 B.n34 585
R335 B.n538 B.n537 585
R336 B.n536 B.n35 585
R337 B.n535 B.n534 585
R338 B.n533 B.n36 585
R339 B.n532 B.n531 585
R340 B.n530 B.n37 585
R341 B.n529 B.n528 585
R342 B.n527 B.n38 585
R343 B.n526 B.n525 585
R344 B.n524 B.n39 585
R345 B.n523 B.n522 585
R346 B.n521 B.n43 585
R347 B.n520 B.n519 585
R348 B.n518 B.n44 585
R349 B.n517 B.n516 585
R350 B.n515 B.n45 585
R351 B.n514 B.n513 585
R352 B.n511 B.n46 585
R353 B.n510 B.n509 585
R354 B.n508 B.n49 585
R355 B.n507 B.n506 585
R356 B.n505 B.n50 585
R357 B.n504 B.n503 585
R358 B.n502 B.n51 585
R359 B.n501 B.n500 585
R360 B.n499 B.n52 585
R361 B.n498 B.n497 585
R362 B.n496 B.n53 585
R363 B.n495 B.n494 585
R364 B.n493 B.n54 585
R365 B.n492 B.n491 585
R366 B.n490 B.n55 585
R367 B.n489 B.n488 585
R368 B.n487 B.n56 585
R369 B.n486 B.n485 585
R370 B.n484 B.n57 585
R371 B.n483 B.n482 585
R372 B.n481 B.n58 585
R373 B.n480 B.n479 585
R374 B.n478 B.n59 585
R375 B.n477 B.n476 585
R376 B.n475 B.n60 585
R377 B.n474 B.n473 585
R378 B.n472 B.n61 585
R379 B.n471 B.n470 585
R380 B.n469 B.n62 585
R381 B.n468 B.n467 585
R382 B.n466 B.n63 585
R383 B.n465 B.n464 585
R384 B.n463 B.n64 585
R385 B.n462 B.n461 585
R386 B.n460 B.n65 585
R387 B.n459 B.n458 585
R388 B.n457 B.n66 585
R389 B.n456 B.n455 585
R390 B.n454 B.n67 585
R391 B.n586 B.n585 585
R392 B.n587 B.n18 585
R393 B.n589 B.n588 585
R394 B.n590 B.n17 585
R395 B.n592 B.n591 585
R396 B.n593 B.n16 585
R397 B.n595 B.n594 585
R398 B.n596 B.n15 585
R399 B.n598 B.n597 585
R400 B.n599 B.n14 585
R401 B.n601 B.n600 585
R402 B.n602 B.n13 585
R403 B.n604 B.n603 585
R404 B.n605 B.n12 585
R405 B.n607 B.n606 585
R406 B.n608 B.n11 585
R407 B.n610 B.n609 585
R408 B.n611 B.n10 585
R409 B.n613 B.n612 585
R410 B.n614 B.n9 585
R411 B.n616 B.n615 585
R412 B.n617 B.n8 585
R413 B.n619 B.n618 585
R414 B.n620 B.n7 585
R415 B.n622 B.n621 585
R416 B.n623 B.n6 585
R417 B.n625 B.n624 585
R418 B.n626 B.n5 585
R419 B.n628 B.n627 585
R420 B.n629 B.n4 585
R421 B.n631 B.n630 585
R422 B.n632 B.n3 585
R423 B.n634 B.n633 585
R424 B.n635 B.n0 585
R425 B.n2 B.n1 585
R426 B.n167 B.n166 585
R427 B.n169 B.n168 585
R428 B.n170 B.n165 585
R429 B.n172 B.n171 585
R430 B.n173 B.n164 585
R431 B.n175 B.n174 585
R432 B.n176 B.n163 585
R433 B.n178 B.n177 585
R434 B.n179 B.n162 585
R435 B.n181 B.n180 585
R436 B.n182 B.n161 585
R437 B.n184 B.n183 585
R438 B.n185 B.n160 585
R439 B.n187 B.n186 585
R440 B.n188 B.n159 585
R441 B.n190 B.n189 585
R442 B.n191 B.n158 585
R443 B.n193 B.n192 585
R444 B.n194 B.n157 585
R445 B.n196 B.n195 585
R446 B.n197 B.n156 585
R447 B.n199 B.n198 585
R448 B.n200 B.n155 585
R449 B.n202 B.n201 585
R450 B.n203 B.n154 585
R451 B.n205 B.n204 585
R452 B.n206 B.n153 585
R453 B.n208 B.n207 585
R454 B.n209 B.n152 585
R455 B.n211 B.n210 585
R456 B.n212 B.n151 585
R457 B.n214 B.n213 585
R458 B.n215 B.n150 585
R459 B.n217 B.n150 574.183
R460 B.n347 B.n102 574.183
R461 B.n454 B.n453 574.183
R462 B.n586 B.n19 574.183
R463 B.n129 B.t0 430.307
R464 B.n123 B.t9 430.307
R465 B.n47 B.t6 430.307
R466 B.n40 B.t3 430.307
R467 B.n637 B.n636 256.663
R468 B.n636 B.n635 235.042
R469 B.n636 B.n2 235.042
R470 B.n218 B.n217 163.367
R471 B.n219 B.n218 163.367
R472 B.n219 B.n148 163.367
R473 B.n223 B.n148 163.367
R474 B.n224 B.n223 163.367
R475 B.n225 B.n224 163.367
R476 B.n225 B.n146 163.367
R477 B.n229 B.n146 163.367
R478 B.n230 B.n229 163.367
R479 B.n231 B.n230 163.367
R480 B.n231 B.n144 163.367
R481 B.n235 B.n144 163.367
R482 B.n236 B.n235 163.367
R483 B.n237 B.n236 163.367
R484 B.n237 B.n142 163.367
R485 B.n241 B.n142 163.367
R486 B.n242 B.n241 163.367
R487 B.n243 B.n242 163.367
R488 B.n243 B.n140 163.367
R489 B.n247 B.n140 163.367
R490 B.n248 B.n247 163.367
R491 B.n249 B.n248 163.367
R492 B.n249 B.n138 163.367
R493 B.n253 B.n138 163.367
R494 B.n254 B.n253 163.367
R495 B.n255 B.n254 163.367
R496 B.n255 B.n136 163.367
R497 B.n259 B.n136 163.367
R498 B.n260 B.n259 163.367
R499 B.n261 B.n260 163.367
R500 B.n261 B.n134 163.367
R501 B.n265 B.n134 163.367
R502 B.n266 B.n265 163.367
R503 B.n267 B.n266 163.367
R504 B.n267 B.n132 163.367
R505 B.n271 B.n132 163.367
R506 B.n272 B.n271 163.367
R507 B.n273 B.n272 163.367
R508 B.n273 B.n128 163.367
R509 B.n278 B.n128 163.367
R510 B.n279 B.n278 163.367
R511 B.n280 B.n279 163.367
R512 B.n280 B.n126 163.367
R513 B.n284 B.n126 163.367
R514 B.n285 B.n284 163.367
R515 B.n286 B.n285 163.367
R516 B.n286 B.n122 163.367
R517 B.n291 B.n122 163.367
R518 B.n292 B.n291 163.367
R519 B.n293 B.n292 163.367
R520 B.n293 B.n120 163.367
R521 B.n297 B.n120 163.367
R522 B.n298 B.n297 163.367
R523 B.n299 B.n298 163.367
R524 B.n299 B.n118 163.367
R525 B.n303 B.n118 163.367
R526 B.n304 B.n303 163.367
R527 B.n305 B.n304 163.367
R528 B.n305 B.n116 163.367
R529 B.n309 B.n116 163.367
R530 B.n310 B.n309 163.367
R531 B.n311 B.n310 163.367
R532 B.n311 B.n114 163.367
R533 B.n315 B.n114 163.367
R534 B.n316 B.n315 163.367
R535 B.n317 B.n316 163.367
R536 B.n317 B.n112 163.367
R537 B.n321 B.n112 163.367
R538 B.n322 B.n321 163.367
R539 B.n323 B.n322 163.367
R540 B.n323 B.n110 163.367
R541 B.n327 B.n110 163.367
R542 B.n328 B.n327 163.367
R543 B.n329 B.n328 163.367
R544 B.n329 B.n108 163.367
R545 B.n333 B.n108 163.367
R546 B.n334 B.n333 163.367
R547 B.n335 B.n334 163.367
R548 B.n335 B.n106 163.367
R549 B.n339 B.n106 163.367
R550 B.n340 B.n339 163.367
R551 B.n341 B.n340 163.367
R552 B.n341 B.n104 163.367
R553 B.n345 B.n104 163.367
R554 B.n346 B.n345 163.367
R555 B.n347 B.n346 163.367
R556 B.n453 B.n68 163.367
R557 B.n449 B.n68 163.367
R558 B.n449 B.n448 163.367
R559 B.n448 B.n447 163.367
R560 B.n447 B.n70 163.367
R561 B.n443 B.n70 163.367
R562 B.n443 B.n442 163.367
R563 B.n442 B.n441 163.367
R564 B.n441 B.n72 163.367
R565 B.n437 B.n72 163.367
R566 B.n437 B.n436 163.367
R567 B.n436 B.n435 163.367
R568 B.n435 B.n74 163.367
R569 B.n431 B.n74 163.367
R570 B.n431 B.n430 163.367
R571 B.n430 B.n429 163.367
R572 B.n429 B.n76 163.367
R573 B.n425 B.n76 163.367
R574 B.n425 B.n424 163.367
R575 B.n424 B.n423 163.367
R576 B.n423 B.n78 163.367
R577 B.n419 B.n78 163.367
R578 B.n419 B.n418 163.367
R579 B.n418 B.n417 163.367
R580 B.n417 B.n80 163.367
R581 B.n413 B.n80 163.367
R582 B.n413 B.n412 163.367
R583 B.n412 B.n411 163.367
R584 B.n411 B.n82 163.367
R585 B.n407 B.n82 163.367
R586 B.n407 B.n406 163.367
R587 B.n406 B.n405 163.367
R588 B.n405 B.n84 163.367
R589 B.n401 B.n84 163.367
R590 B.n401 B.n400 163.367
R591 B.n400 B.n399 163.367
R592 B.n399 B.n86 163.367
R593 B.n395 B.n86 163.367
R594 B.n395 B.n394 163.367
R595 B.n394 B.n393 163.367
R596 B.n393 B.n88 163.367
R597 B.n389 B.n88 163.367
R598 B.n389 B.n388 163.367
R599 B.n388 B.n387 163.367
R600 B.n387 B.n90 163.367
R601 B.n383 B.n90 163.367
R602 B.n383 B.n382 163.367
R603 B.n382 B.n381 163.367
R604 B.n381 B.n92 163.367
R605 B.n377 B.n92 163.367
R606 B.n377 B.n376 163.367
R607 B.n376 B.n375 163.367
R608 B.n375 B.n94 163.367
R609 B.n371 B.n94 163.367
R610 B.n371 B.n370 163.367
R611 B.n370 B.n369 163.367
R612 B.n369 B.n96 163.367
R613 B.n365 B.n96 163.367
R614 B.n365 B.n364 163.367
R615 B.n364 B.n363 163.367
R616 B.n363 B.n98 163.367
R617 B.n359 B.n98 163.367
R618 B.n359 B.n358 163.367
R619 B.n358 B.n357 163.367
R620 B.n357 B.n100 163.367
R621 B.n353 B.n100 163.367
R622 B.n353 B.n352 163.367
R623 B.n352 B.n351 163.367
R624 B.n351 B.n102 163.367
R625 B.n582 B.n19 163.367
R626 B.n582 B.n581 163.367
R627 B.n581 B.n580 163.367
R628 B.n580 B.n21 163.367
R629 B.n576 B.n21 163.367
R630 B.n576 B.n575 163.367
R631 B.n575 B.n574 163.367
R632 B.n574 B.n23 163.367
R633 B.n570 B.n23 163.367
R634 B.n570 B.n569 163.367
R635 B.n569 B.n568 163.367
R636 B.n568 B.n25 163.367
R637 B.n564 B.n25 163.367
R638 B.n564 B.n563 163.367
R639 B.n563 B.n562 163.367
R640 B.n562 B.n27 163.367
R641 B.n558 B.n27 163.367
R642 B.n558 B.n557 163.367
R643 B.n557 B.n556 163.367
R644 B.n556 B.n29 163.367
R645 B.n552 B.n29 163.367
R646 B.n552 B.n551 163.367
R647 B.n551 B.n550 163.367
R648 B.n550 B.n31 163.367
R649 B.n546 B.n31 163.367
R650 B.n546 B.n545 163.367
R651 B.n545 B.n544 163.367
R652 B.n544 B.n33 163.367
R653 B.n540 B.n33 163.367
R654 B.n540 B.n539 163.367
R655 B.n539 B.n538 163.367
R656 B.n538 B.n35 163.367
R657 B.n534 B.n35 163.367
R658 B.n534 B.n533 163.367
R659 B.n533 B.n532 163.367
R660 B.n532 B.n37 163.367
R661 B.n528 B.n37 163.367
R662 B.n528 B.n527 163.367
R663 B.n527 B.n526 163.367
R664 B.n526 B.n39 163.367
R665 B.n522 B.n39 163.367
R666 B.n522 B.n521 163.367
R667 B.n521 B.n520 163.367
R668 B.n520 B.n44 163.367
R669 B.n516 B.n44 163.367
R670 B.n516 B.n515 163.367
R671 B.n515 B.n514 163.367
R672 B.n514 B.n46 163.367
R673 B.n509 B.n46 163.367
R674 B.n509 B.n508 163.367
R675 B.n508 B.n507 163.367
R676 B.n507 B.n50 163.367
R677 B.n503 B.n50 163.367
R678 B.n503 B.n502 163.367
R679 B.n502 B.n501 163.367
R680 B.n501 B.n52 163.367
R681 B.n497 B.n52 163.367
R682 B.n497 B.n496 163.367
R683 B.n496 B.n495 163.367
R684 B.n495 B.n54 163.367
R685 B.n491 B.n54 163.367
R686 B.n491 B.n490 163.367
R687 B.n490 B.n489 163.367
R688 B.n489 B.n56 163.367
R689 B.n485 B.n56 163.367
R690 B.n485 B.n484 163.367
R691 B.n484 B.n483 163.367
R692 B.n483 B.n58 163.367
R693 B.n479 B.n58 163.367
R694 B.n479 B.n478 163.367
R695 B.n478 B.n477 163.367
R696 B.n477 B.n60 163.367
R697 B.n473 B.n60 163.367
R698 B.n473 B.n472 163.367
R699 B.n472 B.n471 163.367
R700 B.n471 B.n62 163.367
R701 B.n467 B.n62 163.367
R702 B.n467 B.n466 163.367
R703 B.n466 B.n465 163.367
R704 B.n465 B.n64 163.367
R705 B.n461 B.n64 163.367
R706 B.n461 B.n460 163.367
R707 B.n460 B.n459 163.367
R708 B.n459 B.n66 163.367
R709 B.n455 B.n66 163.367
R710 B.n455 B.n454 163.367
R711 B.n587 B.n586 163.367
R712 B.n588 B.n587 163.367
R713 B.n588 B.n17 163.367
R714 B.n592 B.n17 163.367
R715 B.n593 B.n592 163.367
R716 B.n594 B.n593 163.367
R717 B.n594 B.n15 163.367
R718 B.n598 B.n15 163.367
R719 B.n599 B.n598 163.367
R720 B.n600 B.n599 163.367
R721 B.n600 B.n13 163.367
R722 B.n604 B.n13 163.367
R723 B.n605 B.n604 163.367
R724 B.n606 B.n605 163.367
R725 B.n606 B.n11 163.367
R726 B.n610 B.n11 163.367
R727 B.n611 B.n610 163.367
R728 B.n612 B.n611 163.367
R729 B.n612 B.n9 163.367
R730 B.n616 B.n9 163.367
R731 B.n617 B.n616 163.367
R732 B.n618 B.n617 163.367
R733 B.n618 B.n7 163.367
R734 B.n622 B.n7 163.367
R735 B.n623 B.n622 163.367
R736 B.n624 B.n623 163.367
R737 B.n624 B.n5 163.367
R738 B.n628 B.n5 163.367
R739 B.n629 B.n628 163.367
R740 B.n630 B.n629 163.367
R741 B.n630 B.n3 163.367
R742 B.n634 B.n3 163.367
R743 B.n635 B.n634 163.367
R744 B.n166 B.n2 163.367
R745 B.n169 B.n166 163.367
R746 B.n170 B.n169 163.367
R747 B.n171 B.n170 163.367
R748 B.n171 B.n164 163.367
R749 B.n175 B.n164 163.367
R750 B.n176 B.n175 163.367
R751 B.n177 B.n176 163.367
R752 B.n177 B.n162 163.367
R753 B.n181 B.n162 163.367
R754 B.n182 B.n181 163.367
R755 B.n183 B.n182 163.367
R756 B.n183 B.n160 163.367
R757 B.n187 B.n160 163.367
R758 B.n188 B.n187 163.367
R759 B.n189 B.n188 163.367
R760 B.n189 B.n158 163.367
R761 B.n193 B.n158 163.367
R762 B.n194 B.n193 163.367
R763 B.n195 B.n194 163.367
R764 B.n195 B.n156 163.367
R765 B.n199 B.n156 163.367
R766 B.n200 B.n199 163.367
R767 B.n201 B.n200 163.367
R768 B.n201 B.n154 163.367
R769 B.n205 B.n154 163.367
R770 B.n206 B.n205 163.367
R771 B.n207 B.n206 163.367
R772 B.n207 B.n152 163.367
R773 B.n211 B.n152 163.367
R774 B.n212 B.n211 163.367
R775 B.n213 B.n212 163.367
R776 B.n213 B.n150 163.367
R777 B.n123 B.t10 140.501
R778 B.n47 B.t8 140.501
R779 B.n129 B.t1 140.488
R780 B.n40 B.t5 140.488
R781 B.n124 B.t11 111.216
R782 B.n48 B.t7 111.216
R783 B.n130 B.t2 111.204
R784 B.n41 B.t4 111.204
R785 B.n275 B.n130 59.5399
R786 B.n289 B.n124 59.5399
R787 B.n512 B.n48 59.5399
R788 B.n42 B.n41 59.5399
R789 B.n585 B.n584 37.3078
R790 B.n452 B.n67 37.3078
R791 B.n349 B.n348 37.3078
R792 B.n216 B.n215 37.3078
R793 B.n130 B.n129 29.2853
R794 B.n124 B.n123 29.2853
R795 B.n48 B.n47 29.2853
R796 B.n41 B.n40 29.2853
R797 B B.n637 18.0485
R798 B.n585 B.n18 10.6151
R799 B.n589 B.n18 10.6151
R800 B.n590 B.n589 10.6151
R801 B.n591 B.n590 10.6151
R802 B.n591 B.n16 10.6151
R803 B.n595 B.n16 10.6151
R804 B.n596 B.n595 10.6151
R805 B.n597 B.n596 10.6151
R806 B.n597 B.n14 10.6151
R807 B.n601 B.n14 10.6151
R808 B.n602 B.n601 10.6151
R809 B.n603 B.n602 10.6151
R810 B.n603 B.n12 10.6151
R811 B.n607 B.n12 10.6151
R812 B.n608 B.n607 10.6151
R813 B.n609 B.n608 10.6151
R814 B.n609 B.n10 10.6151
R815 B.n613 B.n10 10.6151
R816 B.n614 B.n613 10.6151
R817 B.n615 B.n614 10.6151
R818 B.n615 B.n8 10.6151
R819 B.n619 B.n8 10.6151
R820 B.n620 B.n619 10.6151
R821 B.n621 B.n620 10.6151
R822 B.n621 B.n6 10.6151
R823 B.n625 B.n6 10.6151
R824 B.n626 B.n625 10.6151
R825 B.n627 B.n626 10.6151
R826 B.n627 B.n4 10.6151
R827 B.n631 B.n4 10.6151
R828 B.n632 B.n631 10.6151
R829 B.n633 B.n632 10.6151
R830 B.n633 B.n0 10.6151
R831 B.n584 B.n583 10.6151
R832 B.n583 B.n20 10.6151
R833 B.n579 B.n20 10.6151
R834 B.n579 B.n578 10.6151
R835 B.n578 B.n577 10.6151
R836 B.n577 B.n22 10.6151
R837 B.n573 B.n22 10.6151
R838 B.n573 B.n572 10.6151
R839 B.n572 B.n571 10.6151
R840 B.n571 B.n24 10.6151
R841 B.n567 B.n24 10.6151
R842 B.n567 B.n566 10.6151
R843 B.n566 B.n565 10.6151
R844 B.n565 B.n26 10.6151
R845 B.n561 B.n26 10.6151
R846 B.n561 B.n560 10.6151
R847 B.n560 B.n559 10.6151
R848 B.n559 B.n28 10.6151
R849 B.n555 B.n28 10.6151
R850 B.n555 B.n554 10.6151
R851 B.n554 B.n553 10.6151
R852 B.n553 B.n30 10.6151
R853 B.n549 B.n30 10.6151
R854 B.n549 B.n548 10.6151
R855 B.n548 B.n547 10.6151
R856 B.n547 B.n32 10.6151
R857 B.n543 B.n32 10.6151
R858 B.n543 B.n542 10.6151
R859 B.n542 B.n541 10.6151
R860 B.n541 B.n34 10.6151
R861 B.n537 B.n34 10.6151
R862 B.n537 B.n536 10.6151
R863 B.n536 B.n535 10.6151
R864 B.n535 B.n36 10.6151
R865 B.n531 B.n36 10.6151
R866 B.n531 B.n530 10.6151
R867 B.n530 B.n529 10.6151
R868 B.n529 B.n38 10.6151
R869 B.n525 B.n524 10.6151
R870 B.n524 B.n523 10.6151
R871 B.n523 B.n43 10.6151
R872 B.n519 B.n43 10.6151
R873 B.n519 B.n518 10.6151
R874 B.n518 B.n517 10.6151
R875 B.n517 B.n45 10.6151
R876 B.n513 B.n45 10.6151
R877 B.n511 B.n510 10.6151
R878 B.n510 B.n49 10.6151
R879 B.n506 B.n49 10.6151
R880 B.n506 B.n505 10.6151
R881 B.n505 B.n504 10.6151
R882 B.n504 B.n51 10.6151
R883 B.n500 B.n51 10.6151
R884 B.n500 B.n499 10.6151
R885 B.n499 B.n498 10.6151
R886 B.n498 B.n53 10.6151
R887 B.n494 B.n53 10.6151
R888 B.n494 B.n493 10.6151
R889 B.n493 B.n492 10.6151
R890 B.n492 B.n55 10.6151
R891 B.n488 B.n55 10.6151
R892 B.n488 B.n487 10.6151
R893 B.n487 B.n486 10.6151
R894 B.n486 B.n57 10.6151
R895 B.n482 B.n57 10.6151
R896 B.n482 B.n481 10.6151
R897 B.n481 B.n480 10.6151
R898 B.n480 B.n59 10.6151
R899 B.n476 B.n59 10.6151
R900 B.n476 B.n475 10.6151
R901 B.n475 B.n474 10.6151
R902 B.n474 B.n61 10.6151
R903 B.n470 B.n61 10.6151
R904 B.n470 B.n469 10.6151
R905 B.n469 B.n468 10.6151
R906 B.n468 B.n63 10.6151
R907 B.n464 B.n63 10.6151
R908 B.n464 B.n463 10.6151
R909 B.n463 B.n462 10.6151
R910 B.n462 B.n65 10.6151
R911 B.n458 B.n65 10.6151
R912 B.n458 B.n457 10.6151
R913 B.n457 B.n456 10.6151
R914 B.n456 B.n67 10.6151
R915 B.n452 B.n451 10.6151
R916 B.n451 B.n450 10.6151
R917 B.n450 B.n69 10.6151
R918 B.n446 B.n69 10.6151
R919 B.n446 B.n445 10.6151
R920 B.n445 B.n444 10.6151
R921 B.n444 B.n71 10.6151
R922 B.n440 B.n71 10.6151
R923 B.n440 B.n439 10.6151
R924 B.n439 B.n438 10.6151
R925 B.n438 B.n73 10.6151
R926 B.n434 B.n73 10.6151
R927 B.n434 B.n433 10.6151
R928 B.n433 B.n432 10.6151
R929 B.n432 B.n75 10.6151
R930 B.n428 B.n75 10.6151
R931 B.n428 B.n427 10.6151
R932 B.n427 B.n426 10.6151
R933 B.n426 B.n77 10.6151
R934 B.n422 B.n77 10.6151
R935 B.n422 B.n421 10.6151
R936 B.n421 B.n420 10.6151
R937 B.n420 B.n79 10.6151
R938 B.n416 B.n79 10.6151
R939 B.n416 B.n415 10.6151
R940 B.n415 B.n414 10.6151
R941 B.n414 B.n81 10.6151
R942 B.n410 B.n81 10.6151
R943 B.n410 B.n409 10.6151
R944 B.n409 B.n408 10.6151
R945 B.n408 B.n83 10.6151
R946 B.n404 B.n83 10.6151
R947 B.n404 B.n403 10.6151
R948 B.n403 B.n402 10.6151
R949 B.n402 B.n85 10.6151
R950 B.n398 B.n85 10.6151
R951 B.n398 B.n397 10.6151
R952 B.n397 B.n396 10.6151
R953 B.n396 B.n87 10.6151
R954 B.n392 B.n87 10.6151
R955 B.n392 B.n391 10.6151
R956 B.n391 B.n390 10.6151
R957 B.n390 B.n89 10.6151
R958 B.n386 B.n89 10.6151
R959 B.n386 B.n385 10.6151
R960 B.n385 B.n384 10.6151
R961 B.n384 B.n91 10.6151
R962 B.n380 B.n91 10.6151
R963 B.n380 B.n379 10.6151
R964 B.n379 B.n378 10.6151
R965 B.n378 B.n93 10.6151
R966 B.n374 B.n93 10.6151
R967 B.n374 B.n373 10.6151
R968 B.n373 B.n372 10.6151
R969 B.n372 B.n95 10.6151
R970 B.n368 B.n95 10.6151
R971 B.n368 B.n367 10.6151
R972 B.n367 B.n366 10.6151
R973 B.n366 B.n97 10.6151
R974 B.n362 B.n97 10.6151
R975 B.n362 B.n361 10.6151
R976 B.n361 B.n360 10.6151
R977 B.n360 B.n99 10.6151
R978 B.n356 B.n99 10.6151
R979 B.n356 B.n355 10.6151
R980 B.n355 B.n354 10.6151
R981 B.n354 B.n101 10.6151
R982 B.n350 B.n101 10.6151
R983 B.n350 B.n349 10.6151
R984 B.n167 B.n1 10.6151
R985 B.n168 B.n167 10.6151
R986 B.n168 B.n165 10.6151
R987 B.n172 B.n165 10.6151
R988 B.n173 B.n172 10.6151
R989 B.n174 B.n173 10.6151
R990 B.n174 B.n163 10.6151
R991 B.n178 B.n163 10.6151
R992 B.n179 B.n178 10.6151
R993 B.n180 B.n179 10.6151
R994 B.n180 B.n161 10.6151
R995 B.n184 B.n161 10.6151
R996 B.n185 B.n184 10.6151
R997 B.n186 B.n185 10.6151
R998 B.n186 B.n159 10.6151
R999 B.n190 B.n159 10.6151
R1000 B.n191 B.n190 10.6151
R1001 B.n192 B.n191 10.6151
R1002 B.n192 B.n157 10.6151
R1003 B.n196 B.n157 10.6151
R1004 B.n197 B.n196 10.6151
R1005 B.n198 B.n197 10.6151
R1006 B.n198 B.n155 10.6151
R1007 B.n202 B.n155 10.6151
R1008 B.n203 B.n202 10.6151
R1009 B.n204 B.n203 10.6151
R1010 B.n204 B.n153 10.6151
R1011 B.n208 B.n153 10.6151
R1012 B.n209 B.n208 10.6151
R1013 B.n210 B.n209 10.6151
R1014 B.n210 B.n151 10.6151
R1015 B.n214 B.n151 10.6151
R1016 B.n215 B.n214 10.6151
R1017 B.n216 B.n149 10.6151
R1018 B.n220 B.n149 10.6151
R1019 B.n221 B.n220 10.6151
R1020 B.n222 B.n221 10.6151
R1021 B.n222 B.n147 10.6151
R1022 B.n226 B.n147 10.6151
R1023 B.n227 B.n226 10.6151
R1024 B.n228 B.n227 10.6151
R1025 B.n228 B.n145 10.6151
R1026 B.n232 B.n145 10.6151
R1027 B.n233 B.n232 10.6151
R1028 B.n234 B.n233 10.6151
R1029 B.n234 B.n143 10.6151
R1030 B.n238 B.n143 10.6151
R1031 B.n239 B.n238 10.6151
R1032 B.n240 B.n239 10.6151
R1033 B.n240 B.n141 10.6151
R1034 B.n244 B.n141 10.6151
R1035 B.n245 B.n244 10.6151
R1036 B.n246 B.n245 10.6151
R1037 B.n246 B.n139 10.6151
R1038 B.n250 B.n139 10.6151
R1039 B.n251 B.n250 10.6151
R1040 B.n252 B.n251 10.6151
R1041 B.n252 B.n137 10.6151
R1042 B.n256 B.n137 10.6151
R1043 B.n257 B.n256 10.6151
R1044 B.n258 B.n257 10.6151
R1045 B.n258 B.n135 10.6151
R1046 B.n262 B.n135 10.6151
R1047 B.n263 B.n262 10.6151
R1048 B.n264 B.n263 10.6151
R1049 B.n264 B.n133 10.6151
R1050 B.n268 B.n133 10.6151
R1051 B.n269 B.n268 10.6151
R1052 B.n270 B.n269 10.6151
R1053 B.n270 B.n131 10.6151
R1054 B.n274 B.n131 10.6151
R1055 B.n277 B.n276 10.6151
R1056 B.n277 B.n127 10.6151
R1057 B.n281 B.n127 10.6151
R1058 B.n282 B.n281 10.6151
R1059 B.n283 B.n282 10.6151
R1060 B.n283 B.n125 10.6151
R1061 B.n287 B.n125 10.6151
R1062 B.n288 B.n287 10.6151
R1063 B.n290 B.n121 10.6151
R1064 B.n294 B.n121 10.6151
R1065 B.n295 B.n294 10.6151
R1066 B.n296 B.n295 10.6151
R1067 B.n296 B.n119 10.6151
R1068 B.n300 B.n119 10.6151
R1069 B.n301 B.n300 10.6151
R1070 B.n302 B.n301 10.6151
R1071 B.n302 B.n117 10.6151
R1072 B.n306 B.n117 10.6151
R1073 B.n307 B.n306 10.6151
R1074 B.n308 B.n307 10.6151
R1075 B.n308 B.n115 10.6151
R1076 B.n312 B.n115 10.6151
R1077 B.n313 B.n312 10.6151
R1078 B.n314 B.n313 10.6151
R1079 B.n314 B.n113 10.6151
R1080 B.n318 B.n113 10.6151
R1081 B.n319 B.n318 10.6151
R1082 B.n320 B.n319 10.6151
R1083 B.n320 B.n111 10.6151
R1084 B.n324 B.n111 10.6151
R1085 B.n325 B.n324 10.6151
R1086 B.n326 B.n325 10.6151
R1087 B.n326 B.n109 10.6151
R1088 B.n330 B.n109 10.6151
R1089 B.n331 B.n330 10.6151
R1090 B.n332 B.n331 10.6151
R1091 B.n332 B.n107 10.6151
R1092 B.n336 B.n107 10.6151
R1093 B.n337 B.n336 10.6151
R1094 B.n338 B.n337 10.6151
R1095 B.n338 B.n105 10.6151
R1096 B.n342 B.n105 10.6151
R1097 B.n343 B.n342 10.6151
R1098 B.n344 B.n343 10.6151
R1099 B.n344 B.n103 10.6151
R1100 B.n348 B.n103 10.6151
R1101 B.n637 B.n0 8.11757
R1102 B.n637 B.n1 8.11757
R1103 B.n525 B.n42 6.5566
R1104 B.n513 B.n512 6.5566
R1105 B.n276 B.n275 6.5566
R1106 B.n289 B.n288 6.5566
R1107 B.n42 B.n38 4.05904
R1108 B.n512 B.n511 4.05904
R1109 B.n275 B.n274 4.05904
R1110 B.n290 B.n289 4.05904
R1111 VN.n6 VN.t4 257.159
R1112 VN.n31 VN.t2 257.159
R1113 VN.n5 VN.t6 226.296
R1114 VN.n3 VN.t3 226.296
R1115 VN.n15 VN.t5 226.296
R1116 VN.n22 VN.t9 226.296
R1117 VN.n30 VN.t7 226.296
R1118 VN.n28 VN.t1 226.296
R1119 VN.n27 VN.t8 226.296
R1120 VN.n46 VN.t0 226.296
R1121 VN.n23 VN.n22 172.613
R1122 VN.n47 VN.n46 172.613
R1123 VN.n45 VN.n24 161.3
R1124 VN.n44 VN.n43 161.3
R1125 VN.n42 VN.n25 161.3
R1126 VN.n41 VN.n40 161.3
R1127 VN.n39 VN.n26 161.3
R1128 VN.n38 VN.n37 161.3
R1129 VN.n36 VN.n35 161.3
R1130 VN.n34 VN.n29 161.3
R1131 VN.n33 VN.n32 161.3
R1132 VN.n21 VN.n0 161.3
R1133 VN.n20 VN.n19 161.3
R1134 VN.n18 VN.n1 161.3
R1135 VN.n17 VN.n16 161.3
R1136 VN.n14 VN.n2 161.3
R1137 VN.n13 VN.n12 161.3
R1138 VN.n11 VN.n10 161.3
R1139 VN.n9 VN.n4 161.3
R1140 VN.n8 VN.n7 161.3
R1141 VN.n6 VN.n5 50.8823
R1142 VN.n31 VN.n30 50.8823
R1143 VN VN.n47 44.9759
R1144 VN.n21 VN.n20 42.0302
R1145 VN.n45 VN.n44 42.0302
R1146 VN.n9 VN.n8 41.0614
R1147 VN.n16 VN.n14 41.0614
R1148 VN.n34 VN.n33 41.0614
R1149 VN.n40 VN.n39 41.0614
R1150 VN.n10 VN.n9 40.0926
R1151 VN.n14 VN.n13 40.0926
R1152 VN.n35 VN.n34 40.0926
R1153 VN.n39 VN.n38 40.0926
R1154 VN.n20 VN.n1 39.1239
R1155 VN.n44 VN.n25 39.1239
R1156 VN.n32 VN.n31 26.821
R1157 VN.n7 VN.n6 26.821
R1158 VN.n22 VN.n21 13.2801
R1159 VN.n46 VN.n45 13.2801
R1160 VN.n8 VN.n5 12.7883
R1161 VN.n16 VN.n15 12.7883
R1162 VN.n33 VN.n30 12.7883
R1163 VN.n40 VN.n27 12.7883
R1164 VN.n10 VN.n3 12.2964
R1165 VN.n13 VN.n3 12.2964
R1166 VN.n38 VN.n28 12.2964
R1167 VN.n35 VN.n28 12.2964
R1168 VN.n15 VN.n1 11.8046
R1169 VN.n27 VN.n25 11.8046
R1170 VN.n47 VN.n24 0.189894
R1171 VN.n43 VN.n24 0.189894
R1172 VN.n43 VN.n42 0.189894
R1173 VN.n42 VN.n41 0.189894
R1174 VN.n41 VN.n26 0.189894
R1175 VN.n37 VN.n26 0.189894
R1176 VN.n37 VN.n36 0.189894
R1177 VN.n36 VN.n29 0.189894
R1178 VN.n32 VN.n29 0.189894
R1179 VN.n7 VN.n4 0.189894
R1180 VN.n11 VN.n4 0.189894
R1181 VN.n12 VN.n11 0.189894
R1182 VN.n12 VN.n2 0.189894
R1183 VN.n17 VN.n2 0.189894
R1184 VN.n18 VN.n17 0.189894
R1185 VN.n19 VN.n18 0.189894
R1186 VN.n19 VN.n0 0.189894
R1187 VN.n23 VN.n0 0.189894
R1188 VN VN.n23 0.0516364
R1189 VDD2.n1 VDD2.t5 80.316
R1190 VDD2.n4 VDD2.t9 79.0144
R1191 VDD2.n3 VDD2.n2 77.0015
R1192 VDD2 VDD2.n7 76.9987
R1193 VDD2.n6 VDD2.n5 76.0808
R1194 VDD2.n1 VDD2.n0 76.0806
R1195 VDD2.n4 VDD2.n3 39.4502
R1196 VDD2.n7 VDD2.t2 2.93416
R1197 VDD2.n7 VDD2.t7 2.93416
R1198 VDD2.n5 VDD2.t1 2.93416
R1199 VDD2.n5 VDD2.t8 2.93416
R1200 VDD2.n2 VDD2.t4 2.93416
R1201 VDD2.n2 VDD2.t0 2.93416
R1202 VDD2.n0 VDD2.t3 2.93416
R1203 VDD2.n0 VDD2.t6 2.93416
R1204 VDD2.n6 VDD2.n4 1.30222
R1205 VDD2 VDD2.n6 0.384121
R1206 VDD2.n3 VDD2.n1 0.270585
C0 w_n2782_n3184# B 7.90073f
C1 VP VDD1 8.143229f
C2 VN B 0.913579f
C3 VTAIL VDD1 10.9917f
C4 VN w_n2782_n3184# 5.51078f
C5 VDD2 B 1.90231f
C6 VDD2 w_n2782_n3184# 2.23844f
C7 VN VDD2 7.89484f
C8 VP B 1.50744f
C9 VTAIL B 2.85647f
C10 VP w_n2782_n3184# 5.8686f
C11 VP VN 6.13296f
C12 VTAIL w_n2782_n3184# 2.8964f
C13 VN VTAIL 7.97867f
C14 VP VDD2 0.402414f
C15 VDD2 VTAIL 11.031f
C16 VP VTAIL 7.99312f
C17 B VDD1 1.83962f
C18 w_n2782_n3184# VDD1 2.16872f
C19 VN VDD1 0.150017f
C20 VDD2 VDD1 1.26404f
C21 VDD2 VSUBS 1.536314f
C22 VDD1 VSUBS 1.325738f
C23 VTAIL VSUBS 0.903668f
C24 VN VSUBS 5.43699f
C25 VP VSUBS 2.382498f
C26 B VSUBS 3.526258f
C27 w_n2782_n3184# VSUBS 0.109199p
C28 VDD2.t5 VSUBS 2.26817f
C29 VDD2.t3 VSUBS 0.223888f
C30 VDD2.t6 VSUBS 0.223888f
C31 VDD2.n0 VSUBS 1.72519f
C32 VDD2.n1 VSUBS 1.25729f
C33 VDD2.t4 VSUBS 0.223888f
C34 VDD2.t0 VSUBS 0.223888f
C35 VDD2.n2 VSUBS 1.73313f
C36 VDD2.n3 VSUBS 2.4083f
C37 VDD2.t9 VSUBS 2.25739f
C38 VDD2.n4 VSUBS 2.82932f
C39 VDD2.t1 VSUBS 0.223888f
C40 VDD2.t8 VSUBS 0.223888f
C41 VDD2.n5 VSUBS 1.72519f
C42 VDD2.n6 VSUBS 0.609064f
C43 VDD2.t2 VSUBS 0.223888f
C44 VDD2.t7 VSUBS 0.223888f
C45 VDD2.n7 VSUBS 1.73309f
C46 VN.n0 VSUBS 0.04269f
C47 VN.t9 VSUBS 1.51714f
C48 VN.n1 VSUBS 0.064649f
C49 VN.n2 VSUBS 0.04269f
C50 VN.t3 VSUBS 1.51714f
C51 VN.n3 VSUBS 0.56048f
C52 VN.n4 VSUBS 0.04269f
C53 VN.t6 VSUBS 1.51714f
C54 VN.n5 VSUBS 0.623565f
C55 VN.t4 VSUBS 1.59939f
C56 VN.n6 VSUBS 0.652595f
C57 VN.n7 VSUBS 0.22203f
C58 VN.n8 VSUBS 0.065422f
C59 VN.n9 VSUBS 0.034493f
C60 VN.n10 VSUBS 0.065064f
C61 VN.n11 VSUBS 0.04269f
C62 VN.n12 VSUBS 0.04269f
C63 VN.n13 VSUBS 0.065064f
C64 VN.n14 VSUBS 0.034493f
C65 VN.t5 VSUBS 1.51714f
C66 VN.n15 VSUBS 0.56048f
C67 VN.n16 VSUBS 0.065422f
C68 VN.n17 VSUBS 0.04269f
C69 VN.n18 VSUBS 0.04269f
C70 VN.n19 VSUBS 0.04269f
C71 VN.n20 VSUBS 0.034602f
C72 VN.n21 VSUBS 0.065728f
C73 VN.n22 VSUBS 0.630805f
C74 VN.n23 VSUBS 0.038015f
C75 VN.n24 VSUBS 0.04269f
C76 VN.t0 VSUBS 1.51714f
C77 VN.n25 VSUBS 0.064649f
C78 VN.n26 VSUBS 0.04269f
C79 VN.t8 VSUBS 1.51714f
C80 VN.n27 VSUBS 0.56048f
C81 VN.t1 VSUBS 1.51714f
C82 VN.n28 VSUBS 0.56048f
C83 VN.n29 VSUBS 0.04269f
C84 VN.t7 VSUBS 1.51714f
C85 VN.n30 VSUBS 0.623565f
C86 VN.t2 VSUBS 1.59939f
C87 VN.n31 VSUBS 0.652595f
C88 VN.n32 VSUBS 0.22203f
C89 VN.n33 VSUBS 0.065422f
C90 VN.n34 VSUBS 0.034493f
C91 VN.n35 VSUBS 0.065064f
C92 VN.n36 VSUBS 0.04269f
C93 VN.n37 VSUBS 0.04269f
C94 VN.n38 VSUBS 0.065064f
C95 VN.n39 VSUBS 0.034493f
C96 VN.n40 VSUBS 0.065422f
C97 VN.n41 VSUBS 0.04269f
C98 VN.n42 VSUBS 0.04269f
C99 VN.n43 VSUBS 0.04269f
C100 VN.n44 VSUBS 0.034602f
C101 VN.n45 VSUBS 0.065728f
C102 VN.n46 VSUBS 0.630805f
C103 VN.n47 VSUBS 1.97632f
C104 B.n0 VSUBS 0.006245f
C105 B.n1 VSUBS 0.006245f
C106 B.n2 VSUBS 0.009236f
C107 B.n3 VSUBS 0.007077f
C108 B.n4 VSUBS 0.007077f
C109 B.n5 VSUBS 0.007077f
C110 B.n6 VSUBS 0.007077f
C111 B.n7 VSUBS 0.007077f
C112 B.n8 VSUBS 0.007077f
C113 B.n9 VSUBS 0.007077f
C114 B.n10 VSUBS 0.007077f
C115 B.n11 VSUBS 0.007077f
C116 B.n12 VSUBS 0.007077f
C117 B.n13 VSUBS 0.007077f
C118 B.n14 VSUBS 0.007077f
C119 B.n15 VSUBS 0.007077f
C120 B.n16 VSUBS 0.007077f
C121 B.n17 VSUBS 0.007077f
C122 B.n18 VSUBS 0.007077f
C123 B.n19 VSUBS 0.018494f
C124 B.n20 VSUBS 0.007077f
C125 B.n21 VSUBS 0.007077f
C126 B.n22 VSUBS 0.007077f
C127 B.n23 VSUBS 0.007077f
C128 B.n24 VSUBS 0.007077f
C129 B.n25 VSUBS 0.007077f
C130 B.n26 VSUBS 0.007077f
C131 B.n27 VSUBS 0.007077f
C132 B.n28 VSUBS 0.007077f
C133 B.n29 VSUBS 0.007077f
C134 B.n30 VSUBS 0.007077f
C135 B.n31 VSUBS 0.007077f
C136 B.n32 VSUBS 0.007077f
C137 B.n33 VSUBS 0.007077f
C138 B.n34 VSUBS 0.007077f
C139 B.n35 VSUBS 0.007077f
C140 B.n36 VSUBS 0.007077f
C141 B.n37 VSUBS 0.007077f
C142 B.n38 VSUBS 0.004892f
C143 B.n39 VSUBS 0.007077f
C144 B.t4 VSUBS 0.361833f
C145 B.t5 VSUBS 0.373605f
C146 B.t3 VSUBS 0.570503f
C147 B.n40 VSUBS 0.156173f
C148 B.n41 VSUBS 0.066567f
C149 B.n42 VSUBS 0.016398f
C150 B.n43 VSUBS 0.007077f
C151 B.n44 VSUBS 0.007077f
C152 B.n45 VSUBS 0.007077f
C153 B.n46 VSUBS 0.007077f
C154 B.t7 VSUBS 0.361827f
C155 B.t8 VSUBS 0.373599f
C156 B.t6 VSUBS 0.570503f
C157 B.n47 VSUBS 0.156178f
C158 B.n48 VSUBS 0.066573f
C159 B.n49 VSUBS 0.007077f
C160 B.n50 VSUBS 0.007077f
C161 B.n51 VSUBS 0.007077f
C162 B.n52 VSUBS 0.007077f
C163 B.n53 VSUBS 0.007077f
C164 B.n54 VSUBS 0.007077f
C165 B.n55 VSUBS 0.007077f
C166 B.n56 VSUBS 0.007077f
C167 B.n57 VSUBS 0.007077f
C168 B.n58 VSUBS 0.007077f
C169 B.n59 VSUBS 0.007077f
C170 B.n60 VSUBS 0.007077f
C171 B.n61 VSUBS 0.007077f
C172 B.n62 VSUBS 0.007077f
C173 B.n63 VSUBS 0.007077f
C174 B.n64 VSUBS 0.007077f
C175 B.n65 VSUBS 0.007077f
C176 B.n66 VSUBS 0.007077f
C177 B.n67 VSUBS 0.018494f
C178 B.n68 VSUBS 0.007077f
C179 B.n69 VSUBS 0.007077f
C180 B.n70 VSUBS 0.007077f
C181 B.n71 VSUBS 0.007077f
C182 B.n72 VSUBS 0.007077f
C183 B.n73 VSUBS 0.007077f
C184 B.n74 VSUBS 0.007077f
C185 B.n75 VSUBS 0.007077f
C186 B.n76 VSUBS 0.007077f
C187 B.n77 VSUBS 0.007077f
C188 B.n78 VSUBS 0.007077f
C189 B.n79 VSUBS 0.007077f
C190 B.n80 VSUBS 0.007077f
C191 B.n81 VSUBS 0.007077f
C192 B.n82 VSUBS 0.007077f
C193 B.n83 VSUBS 0.007077f
C194 B.n84 VSUBS 0.007077f
C195 B.n85 VSUBS 0.007077f
C196 B.n86 VSUBS 0.007077f
C197 B.n87 VSUBS 0.007077f
C198 B.n88 VSUBS 0.007077f
C199 B.n89 VSUBS 0.007077f
C200 B.n90 VSUBS 0.007077f
C201 B.n91 VSUBS 0.007077f
C202 B.n92 VSUBS 0.007077f
C203 B.n93 VSUBS 0.007077f
C204 B.n94 VSUBS 0.007077f
C205 B.n95 VSUBS 0.007077f
C206 B.n96 VSUBS 0.007077f
C207 B.n97 VSUBS 0.007077f
C208 B.n98 VSUBS 0.007077f
C209 B.n99 VSUBS 0.007077f
C210 B.n100 VSUBS 0.007077f
C211 B.n101 VSUBS 0.007077f
C212 B.n102 VSUBS 0.017726f
C213 B.n103 VSUBS 0.007077f
C214 B.n104 VSUBS 0.007077f
C215 B.n105 VSUBS 0.007077f
C216 B.n106 VSUBS 0.007077f
C217 B.n107 VSUBS 0.007077f
C218 B.n108 VSUBS 0.007077f
C219 B.n109 VSUBS 0.007077f
C220 B.n110 VSUBS 0.007077f
C221 B.n111 VSUBS 0.007077f
C222 B.n112 VSUBS 0.007077f
C223 B.n113 VSUBS 0.007077f
C224 B.n114 VSUBS 0.007077f
C225 B.n115 VSUBS 0.007077f
C226 B.n116 VSUBS 0.007077f
C227 B.n117 VSUBS 0.007077f
C228 B.n118 VSUBS 0.007077f
C229 B.n119 VSUBS 0.007077f
C230 B.n120 VSUBS 0.007077f
C231 B.n121 VSUBS 0.007077f
C232 B.n122 VSUBS 0.007077f
C233 B.t11 VSUBS 0.361827f
C234 B.t10 VSUBS 0.373599f
C235 B.t9 VSUBS 0.570503f
C236 B.n123 VSUBS 0.156178f
C237 B.n124 VSUBS 0.066573f
C238 B.n125 VSUBS 0.007077f
C239 B.n126 VSUBS 0.007077f
C240 B.n127 VSUBS 0.007077f
C241 B.n128 VSUBS 0.007077f
C242 B.t2 VSUBS 0.361833f
C243 B.t1 VSUBS 0.373605f
C244 B.t0 VSUBS 0.570503f
C245 B.n129 VSUBS 0.156173f
C246 B.n130 VSUBS 0.066567f
C247 B.n131 VSUBS 0.007077f
C248 B.n132 VSUBS 0.007077f
C249 B.n133 VSUBS 0.007077f
C250 B.n134 VSUBS 0.007077f
C251 B.n135 VSUBS 0.007077f
C252 B.n136 VSUBS 0.007077f
C253 B.n137 VSUBS 0.007077f
C254 B.n138 VSUBS 0.007077f
C255 B.n139 VSUBS 0.007077f
C256 B.n140 VSUBS 0.007077f
C257 B.n141 VSUBS 0.007077f
C258 B.n142 VSUBS 0.007077f
C259 B.n143 VSUBS 0.007077f
C260 B.n144 VSUBS 0.007077f
C261 B.n145 VSUBS 0.007077f
C262 B.n146 VSUBS 0.007077f
C263 B.n147 VSUBS 0.007077f
C264 B.n148 VSUBS 0.007077f
C265 B.n149 VSUBS 0.007077f
C266 B.n150 VSUBS 0.017726f
C267 B.n151 VSUBS 0.007077f
C268 B.n152 VSUBS 0.007077f
C269 B.n153 VSUBS 0.007077f
C270 B.n154 VSUBS 0.007077f
C271 B.n155 VSUBS 0.007077f
C272 B.n156 VSUBS 0.007077f
C273 B.n157 VSUBS 0.007077f
C274 B.n158 VSUBS 0.007077f
C275 B.n159 VSUBS 0.007077f
C276 B.n160 VSUBS 0.007077f
C277 B.n161 VSUBS 0.007077f
C278 B.n162 VSUBS 0.007077f
C279 B.n163 VSUBS 0.007077f
C280 B.n164 VSUBS 0.007077f
C281 B.n165 VSUBS 0.007077f
C282 B.n166 VSUBS 0.007077f
C283 B.n167 VSUBS 0.007077f
C284 B.n168 VSUBS 0.007077f
C285 B.n169 VSUBS 0.007077f
C286 B.n170 VSUBS 0.007077f
C287 B.n171 VSUBS 0.007077f
C288 B.n172 VSUBS 0.007077f
C289 B.n173 VSUBS 0.007077f
C290 B.n174 VSUBS 0.007077f
C291 B.n175 VSUBS 0.007077f
C292 B.n176 VSUBS 0.007077f
C293 B.n177 VSUBS 0.007077f
C294 B.n178 VSUBS 0.007077f
C295 B.n179 VSUBS 0.007077f
C296 B.n180 VSUBS 0.007077f
C297 B.n181 VSUBS 0.007077f
C298 B.n182 VSUBS 0.007077f
C299 B.n183 VSUBS 0.007077f
C300 B.n184 VSUBS 0.007077f
C301 B.n185 VSUBS 0.007077f
C302 B.n186 VSUBS 0.007077f
C303 B.n187 VSUBS 0.007077f
C304 B.n188 VSUBS 0.007077f
C305 B.n189 VSUBS 0.007077f
C306 B.n190 VSUBS 0.007077f
C307 B.n191 VSUBS 0.007077f
C308 B.n192 VSUBS 0.007077f
C309 B.n193 VSUBS 0.007077f
C310 B.n194 VSUBS 0.007077f
C311 B.n195 VSUBS 0.007077f
C312 B.n196 VSUBS 0.007077f
C313 B.n197 VSUBS 0.007077f
C314 B.n198 VSUBS 0.007077f
C315 B.n199 VSUBS 0.007077f
C316 B.n200 VSUBS 0.007077f
C317 B.n201 VSUBS 0.007077f
C318 B.n202 VSUBS 0.007077f
C319 B.n203 VSUBS 0.007077f
C320 B.n204 VSUBS 0.007077f
C321 B.n205 VSUBS 0.007077f
C322 B.n206 VSUBS 0.007077f
C323 B.n207 VSUBS 0.007077f
C324 B.n208 VSUBS 0.007077f
C325 B.n209 VSUBS 0.007077f
C326 B.n210 VSUBS 0.007077f
C327 B.n211 VSUBS 0.007077f
C328 B.n212 VSUBS 0.007077f
C329 B.n213 VSUBS 0.007077f
C330 B.n214 VSUBS 0.007077f
C331 B.n215 VSUBS 0.017726f
C332 B.n216 VSUBS 0.018494f
C333 B.n217 VSUBS 0.018494f
C334 B.n218 VSUBS 0.007077f
C335 B.n219 VSUBS 0.007077f
C336 B.n220 VSUBS 0.007077f
C337 B.n221 VSUBS 0.007077f
C338 B.n222 VSUBS 0.007077f
C339 B.n223 VSUBS 0.007077f
C340 B.n224 VSUBS 0.007077f
C341 B.n225 VSUBS 0.007077f
C342 B.n226 VSUBS 0.007077f
C343 B.n227 VSUBS 0.007077f
C344 B.n228 VSUBS 0.007077f
C345 B.n229 VSUBS 0.007077f
C346 B.n230 VSUBS 0.007077f
C347 B.n231 VSUBS 0.007077f
C348 B.n232 VSUBS 0.007077f
C349 B.n233 VSUBS 0.007077f
C350 B.n234 VSUBS 0.007077f
C351 B.n235 VSUBS 0.007077f
C352 B.n236 VSUBS 0.007077f
C353 B.n237 VSUBS 0.007077f
C354 B.n238 VSUBS 0.007077f
C355 B.n239 VSUBS 0.007077f
C356 B.n240 VSUBS 0.007077f
C357 B.n241 VSUBS 0.007077f
C358 B.n242 VSUBS 0.007077f
C359 B.n243 VSUBS 0.007077f
C360 B.n244 VSUBS 0.007077f
C361 B.n245 VSUBS 0.007077f
C362 B.n246 VSUBS 0.007077f
C363 B.n247 VSUBS 0.007077f
C364 B.n248 VSUBS 0.007077f
C365 B.n249 VSUBS 0.007077f
C366 B.n250 VSUBS 0.007077f
C367 B.n251 VSUBS 0.007077f
C368 B.n252 VSUBS 0.007077f
C369 B.n253 VSUBS 0.007077f
C370 B.n254 VSUBS 0.007077f
C371 B.n255 VSUBS 0.007077f
C372 B.n256 VSUBS 0.007077f
C373 B.n257 VSUBS 0.007077f
C374 B.n258 VSUBS 0.007077f
C375 B.n259 VSUBS 0.007077f
C376 B.n260 VSUBS 0.007077f
C377 B.n261 VSUBS 0.007077f
C378 B.n262 VSUBS 0.007077f
C379 B.n263 VSUBS 0.007077f
C380 B.n264 VSUBS 0.007077f
C381 B.n265 VSUBS 0.007077f
C382 B.n266 VSUBS 0.007077f
C383 B.n267 VSUBS 0.007077f
C384 B.n268 VSUBS 0.007077f
C385 B.n269 VSUBS 0.007077f
C386 B.n270 VSUBS 0.007077f
C387 B.n271 VSUBS 0.007077f
C388 B.n272 VSUBS 0.007077f
C389 B.n273 VSUBS 0.007077f
C390 B.n274 VSUBS 0.004892f
C391 B.n275 VSUBS 0.016398f
C392 B.n276 VSUBS 0.005724f
C393 B.n277 VSUBS 0.007077f
C394 B.n278 VSUBS 0.007077f
C395 B.n279 VSUBS 0.007077f
C396 B.n280 VSUBS 0.007077f
C397 B.n281 VSUBS 0.007077f
C398 B.n282 VSUBS 0.007077f
C399 B.n283 VSUBS 0.007077f
C400 B.n284 VSUBS 0.007077f
C401 B.n285 VSUBS 0.007077f
C402 B.n286 VSUBS 0.007077f
C403 B.n287 VSUBS 0.007077f
C404 B.n288 VSUBS 0.005724f
C405 B.n289 VSUBS 0.016398f
C406 B.n290 VSUBS 0.004892f
C407 B.n291 VSUBS 0.007077f
C408 B.n292 VSUBS 0.007077f
C409 B.n293 VSUBS 0.007077f
C410 B.n294 VSUBS 0.007077f
C411 B.n295 VSUBS 0.007077f
C412 B.n296 VSUBS 0.007077f
C413 B.n297 VSUBS 0.007077f
C414 B.n298 VSUBS 0.007077f
C415 B.n299 VSUBS 0.007077f
C416 B.n300 VSUBS 0.007077f
C417 B.n301 VSUBS 0.007077f
C418 B.n302 VSUBS 0.007077f
C419 B.n303 VSUBS 0.007077f
C420 B.n304 VSUBS 0.007077f
C421 B.n305 VSUBS 0.007077f
C422 B.n306 VSUBS 0.007077f
C423 B.n307 VSUBS 0.007077f
C424 B.n308 VSUBS 0.007077f
C425 B.n309 VSUBS 0.007077f
C426 B.n310 VSUBS 0.007077f
C427 B.n311 VSUBS 0.007077f
C428 B.n312 VSUBS 0.007077f
C429 B.n313 VSUBS 0.007077f
C430 B.n314 VSUBS 0.007077f
C431 B.n315 VSUBS 0.007077f
C432 B.n316 VSUBS 0.007077f
C433 B.n317 VSUBS 0.007077f
C434 B.n318 VSUBS 0.007077f
C435 B.n319 VSUBS 0.007077f
C436 B.n320 VSUBS 0.007077f
C437 B.n321 VSUBS 0.007077f
C438 B.n322 VSUBS 0.007077f
C439 B.n323 VSUBS 0.007077f
C440 B.n324 VSUBS 0.007077f
C441 B.n325 VSUBS 0.007077f
C442 B.n326 VSUBS 0.007077f
C443 B.n327 VSUBS 0.007077f
C444 B.n328 VSUBS 0.007077f
C445 B.n329 VSUBS 0.007077f
C446 B.n330 VSUBS 0.007077f
C447 B.n331 VSUBS 0.007077f
C448 B.n332 VSUBS 0.007077f
C449 B.n333 VSUBS 0.007077f
C450 B.n334 VSUBS 0.007077f
C451 B.n335 VSUBS 0.007077f
C452 B.n336 VSUBS 0.007077f
C453 B.n337 VSUBS 0.007077f
C454 B.n338 VSUBS 0.007077f
C455 B.n339 VSUBS 0.007077f
C456 B.n340 VSUBS 0.007077f
C457 B.n341 VSUBS 0.007077f
C458 B.n342 VSUBS 0.007077f
C459 B.n343 VSUBS 0.007077f
C460 B.n344 VSUBS 0.007077f
C461 B.n345 VSUBS 0.007077f
C462 B.n346 VSUBS 0.007077f
C463 B.n347 VSUBS 0.018494f
C464 B.n348 VSUBS 0.017762f
C465 B.n349 VSUBS 0.018458f
C466 B.n350 VSUBS 0.007077f
C467 B.n351 VSUBS 0.007077f
C468 B.n352 VSUBS 0.007077f
C469 B.n353 VSUBS 0.007077f
C470 B.n354 VSUBS 0.007077f
C471 B.n355 VSUBS 0.007077f
C472 B.n356 VSUBS 0.007077f
C473 B.n357 VSUBS 0.007077f
C474 B.n358 VSUBS 0.007077f
C475 B.n359 VSUBS 0.007077f
C476 B.n360 VSUBS 0.007077f
C477 B.n361 VSUBS 0.007077f
C478 B.n362 VSUBS 0.007077f
C479 B.n363 VSUBS 0.007077f
C480 B.n364 VSUBS 0.007077f
C481 B.n365 VSUBS 0.007077f
C482 B.n366 VSUBS 0.007077f
C483 B.n367 VSUBS 0.007077f
C484 B.n368 VSUBS 0.007077f
C485 B.n369 VSUBS 0.007077f
C486 B.n370 VSUBS 0.007077f
C487 B.n371 VSUBS 0.007077f
C488 B.n372 VSUBS 0.007077f
C489 B.n373 VSUBS 0.007077f
C490 B.n374 VSUBS 0.007077f
C491 B.n375 VSUBS 0.007077f
C492 B.n376 VSUBS 0.007077f
C493 B.n377 VSUBS 0.007077f
C494 B.n378 VSUBS 0.007077f
C495 B.n379 VSUBS 0.007077f
C496 B.n380 VSUBS 0.007077f
C497 B.n381 VSUBS 0.007077f
C498 B.n382 VSUBS 0.007077f
C499 B.n383 VSUBS 0.007077f
C500 B.n384 VSUBS 0.007077f
C501 B.n385 VSUBS 0.007077f
C502 B.n386 VSUBS 0.007077f
C503 B.n387 VSUBS 0.007077f
C504 B.n388 VSUBS 0.007077f
C505 B.n389 VSUBS 0.007077f
C506 B.n390 VSUBS 0.007077f
C507 B.n391 VSUBS 0.007077f
C508 B.n392 VSUBS 0.007077f
C509 B.n393 VSUBS 0.007077f
C510 B.n394 VSUBS 0.007077f
C511 B.n395 VSUBS 0.007077f
C512 B.n396 VSUBS 0.007077f
C513 B.n397 VSUBS 0.007077f
C514 B.n398 VSUBS 0.007077f
C515 B.n399 VSUBS 0.007077f
C516 B.n400 VSUBS 0.007077f
C517 B.n401 VSUBS 0.007077f
C518 B.n402 VSUBS 0.007077f
C519 B.n403 VSUBS 0.007077f
C520 B.n404 VSUBS 0.007077f
C521 B.n405 VSUBS 0.007077f
C522 B.n406 VSUBS 0.007077f
C523 B.n407 VSUBS 0.007077f
C524 B.n408 VSUBS 0.007077f
C525 B.n409 VSUBS 0.007077f
C526 B.n410 VSUBS 0.007077f
C527 B.n411 VSUBS 0.007077f
C528 B.n412 VSUBS 0.007077f
C529 B.n413 VSUBS 0.007077f
C530 B.n414 VSUBS 0.007077f
C531 B.n415 VSUBS 0.007077f
C532 B.n416 VSUBS 0.007077f
C533 B.n417 VSUBS 0.007077f
C534 B.n418 VSUBS 0.007077f
C535 B.n419 VSUBS 0.007077f
C536 B.n420 VSUBS 0.007077f
C537 B.n421 VSUBS 0.007077f
C538 B.n422 VSUBS 0.007077f
C539 B.n423 VSUBS 0.007077f
C540 B.n424 VSUBS 0.007077f
C541 B.n425 VSUBS 0.007077f
C542 B.n426 VSUBS 0.007077f
C543 B.n427 VSUBS 0.007077f
C544 B.n428 VSUBS 0.007077f
C545 B.n429 VSUBS 0.007077f
C546 B.n430 VSUBS 0.007077f
C547 B.n431 VSUBS 0.007077f
C548 B.n432 VSUBS 0.007077f
C549 B.n433 VSUBS 0.007077f
C550 B.n434 VSUBS 0.007077f
C551 B.n435 VSUBS 0.007077f
C552 B.n436 VSUBS 0.007077f
C553 B.n437 VSUBS 0.007077f
C554 B.n438 VSUBS 0.007077f
C555 B.n439 VSUBS 0.007077f
C556 B.n440 VSUBS 0.007077f
C557 B.n441 VSUBS 0.007077f
C558 B.n442 VSUBS 0.007077f
C559 B.n443 VSUBS 0.007077f
C560 B.n444 VSUBS 0.007077f
C561 B.n445 VSUBS 0.007077f
C562 B.n446 VSUBS 0.007077f
C563 B.n447 VSUBS 0.007077f
C564 B.n448 VSUBS 0.007077f
C565 B.n449 VSUBS 0.007077f
C566 B.n450 VSUBS 0.007077f
C567 B.n451 VSUBS 0.007077f
C568 B.n452 VSUBS 0.017726f
C569 B.n453 VSUBS 0.017726f
C570 B.n454 VSUBS 0.018494f
C571 B.n455 VSUBS 0.007077f
C572 B.n456 VSUBS 0.007077f
C573 B.n457 VSUBS 0.007077f
C574 B.n458 VSUBS 0.007077f
C575 B.n459 VSUBS 0.007077f
C576 B.n460 VSUBS 0.007077f
C577 B.n461 VSUBS 0.007077f
C578 B.n462 VSUBS 0.007077f
C579 B.n463 VSUBS 0.007077f
C580 B.n464 VSUBS 0.007077f
C581 B.n465 VSUBS 0.007077f
C582 B.n466 VSUBS 0.007077f
C583 B.n467 VSUBS 0.007077f
C584 B.n468 VSUBS 0.007077f
C585 B.n469 VSUBS 0.007077f
C586 B.n470 VSUBS 0.007077f
C587 B.n471 VSUBS 0.007077f
C588 B.n472 VSUBS 0.007077f
C589 B.n473 VSUBS 0.007077f
C590 B.n474 VSUBS 0.007077f
C591 B.n475 VSUBS 0.007077f
C592 B.n476 VSUBS 0.007077f
C593 B.n477 VSUBS 0.007077f
C594 B.n478 VSUBS 0.007077f
C595 B.n479 VSUBS 0.007077f
C596 B.n480 VSUBS 0.007077f
C597 B.n481 VSUBS 0.007077f
C598 B.n482 VSUBS 0.007077f
C599 B.n483 VSUBS 0.007077f
C600 B.n484 VSUBS 0.007077f
C601 B.n485 VSUBS 0.007077f
C602 B.n486 VSUBS 0.007077f
C603 B.n487 VSUBS 0.007077f
C604 B.n488 VSUBS 0.007077f
C605 B.n489 VSUBS 0.007077f
C606 B.n490 VSUBS 0.007077f
C607 B.n491 VSUBS 0.007077f
C608 B.n492 VSUBS 0.007077f
C609 B.n493 VSUBS 0.007077f
C610 B.n494 VSUBS 0.007077f
C611 B.n495 VSUBS 0.007077f
C612 B.n496 VSUBS 0.007077f
C613 B.n497 VSUBS 0.007077f
C614 B.n498 VSUBS 0.007077f
C615 B.n499 VSUBS 0.007077f
C616 B.n500 VSUBS 0.007077f
C617 B.n501 VSUBS 0.007077f
C618 B.n502 VSUBS 0.007077f
C619 B.n503 VSUBS 0.007077f
C620 B.n504 VSUBS 0.007077f
C621 B.n505 VSUBS 0.007077f
C622 B.n506 VSUBS 0.007077f
C623 B.n507 VSUBS 0.007077f
C624 B.n508 VSUBS 0.007077f
C625 B.n509 VSUBS 0.007077f
C626 B.n510 VSUBS 0.007077f
C627 B.n511 VSUBS 0.004892f
C628 B.n512 VSUBS 0.016398f
C629 B.n513 VSUBS 0.005724f
C630 B.n514 VSUBS 0.007077f
C631 B.n515 VSUBS 0.007077f
C632 B.n516 VSUBS 0.007077f
C633 B.n517 VSUBS 0.007077f
C634 B.n518 VSUBS 0.007077f
C635 B.n519 VSUBS 0.007077f
C636 B.n520 VSUBS 0.007077f
C637 B.n521 VSUBS 0.007077f
C638 B.n522 VSUBS 0.007077f
C639 B.n523 VSUBS 0.007077f
C640 B.n524 VSUBS 0.007077f
C641 B.n525 VSUBS 0.005724f
C642 B.n526 VSUBS 0.007077f
C643 B.n527 VSUBS 0.007077f
C644 B.n528 VSUBS 0.007077f
C645 B.n529 VSUBS 0.007077f
C646 B.n530 VSUBS 0.007077f
C647 B.n531 VSUBS 0.007077f
C648 B.n532 VSUBS 0.007077f
C649 B.n533 VSUBS 0.007077f
C650 B.n534 VSUBS 0.007077f
C651 B.n535 VSUBS 0.007077f
C652 B.n536 VSUBS 0.007077f
C653 B.n537 VSUBS 0.007077f
C654 B.n538 VSUBS 0.007077f
C655 B.n539 VSUBS 0.007077f
C656 B.n540 VSUBS 0.007077f
C657 B.n541 VSUBS 0.007077f
C658 B.n542 VSUBS 0.007077f
C659 B.n543 VSUBS 0.007077f
C660 B.n544 VSUBS 0.007077f
C661 B.n545 VSUBS 0.007077f
C662 B.n546 VSUBS 0.007077f
C663 B.n547 VSUBS 0.007077f
C664 B.n548 VSUBS 0.007077f
C665 B.n549 VSUBS 0.007077f
C666 B.n550 VSUBS 0.007077f
C667 B.n551 VSUBS 0.007077f
C668 B.n552 VSUBS 0.007077f
C669 B.n553 VSUBS 0.007077f
C670 B.n554 VSUBS 0.007077f
C671 B.n555 VSUBS 0.007077f
C672 B.n556 VSUBS 0.007077f
C673 B.n557 VSUBS 0.007077f
C674 B.n558 VSUBS 0.007077f
C675 B.n559 VSUBS 0.007077f
C676 B.n560 VSUBS 0.007077f
C677 B.n561 VSUBS 0.007077f
C678 B.n562 VSUBS 0.007077f
C679 B.n563 VSUBS 0.007077f
C680 B.n564 VSUBS 0.007077f
C681 B.n565 VSUBS 0.007077f
C682 B.n566 VSUBS 0.007077f
C683 B.n567 VSUBS 0.007077f
C684 B.n568 VSUBS 0.007077f
C685 B.n569 VSUBS 0.007077f
C686 B.n570 VSUBS 0.007077f
C687 B.n571 VSUBS 0.007077f
C688 B.n572 VSUBS 0.007077f
C689 B.n573 VSUBS 0.007077f
C690 B.n574 VSUBS 0.007077f
C691 B.n575 VSUBS 0.007077f
C692 B.n576 VSUBS 0.007077f
C693 B.n577 VSUBS 0.007077f
C694 B.n578 VSUBS 0.007077f
C695 B.n579 VSUBS 0.007077f
C696 B.n580 VSUBS 0.007077f
C697 B.n581 VSUBS 0.007077f
C698 B.n582 VSUBS 0.007077f
C699 B.n583 VSUBS 0.007077f
C700 B.n584 VSUBS 0.018494f
C701 B.n585 VSUBS 0.017726f
C702 B.n586 VSUBS 0.017726f
C703 B.n587 VSUBS 0.007077f
C704 B.n588 VSUBS 0.007077f
C705 B.n589 VSUBS 0.007077f
C706 B.n590 VSUBS 0.007077f
C707 B.n591 VSUBS 0.007077f
C708 B.n592 VSUBS 0.007077f
C709 B.n593 VSUBS 0.007077f
C710 B.n594 VSUBS 0.007077f
C711 B.n595 VSUBS 0.007077f
C712 B.n596 VSUBS 0.007077f
C713 B.n597 VSUBS 0.007077f
C714 B.n598 VSUBS 0.007077f
C715 B.n599 VSUBS 0.007077f
C716 B.n600 VSUBS 0.007077f
C717 B.n601 VSUBS 0.007077f
C718 B.n602 VSUBS 0.007077f
C719 B.n603 VSUBS 0.007077f
C720 B.n604 VSUBS 0.007077f
C721 B.n605 VSUBS 0.007077f
C722 B.n606 VSUBS 0.007077f
C723 B.n607 VSUBS 0.007077f
C724 B.n608 VSUBS 0.007077f
C725 B.n609 VSUBS 0.007077f
C726 B.n610 VSUBS 0.007077f
C727 B.n611 VSUBS 0.007077f
C728 B.n612 VSUBS 0.007077f
C729 B.n613 VSUBS 0.007077f
C730 B.n614 VSUBS 0.007077f
C731 B.n615 VSUBS 0.007077f
C732 B.n616 VSUBS 0.007077f
C733 B.n617 VSUBS 0.007077f
C734 B.n618 VSUBS 0.007077f
C735 B.n619 VSUBS 0.007077f
C736 B.n620 VSUBS 0.007077f
C737 B.n621 VSUBS 0.007077f
C738 B.n622 VSUBS 0.007077f
C739 B.n623 VSUBS 0.007077f
C740 B.n624 VSUBS 0.007077f
C741 B.n625 VSUBS 0.007077f
C742 B.n626 VSUBS 0.007077f
C743 B.n627 VSUBS 0.007077f
C744 B.n628 VSUBS 0.007077f
C745 B.n629 VSUBS 0.007077f
C746 B.n630 VSUBS 0.007077f
C747 B.n631 VSUBS 0.007077f
C748 B.n632 VSUBS 0.007077f
C749 B.n633 VSUBS 0.007077f
C750 B.n634 VSUBS 0.007077f
C751 B.n635 VSUBS 0.009236f
C752 B.n636 VSUBS 0.009838f
C753 B.n637 VSUBS 0.019565f
C754 VDD1.t9 VSUBS 2.27948f
C755 VDD1.t2 VSUBS 0.225003f
C756 VDD1.t0 VSUBS 0.225003f
C757 VDD1.n0 VSUBS 1.73378f
C758 VDD1.n1 VSUBS 1.27073f
C759 VDD1.t7 VSUBS 2.27947f
C760 VDD1.t5 VSUBS 0.225003f
C761 VDD1.t3 VSUBS 0.225003f
C762 VDD1.n2 VSUBS 1.73378f
C763 VDD1.n3 VSUBS 1.26355f
C764 VDD1.t6 VSUBS 0.225003f
C765 VDD1.t8 VSUBS 0.225003f
C766 VDD1.n4 VSUBS 1.74176f
C767 VDD1.n5 VSUBS 2.51083f
C768 VDD1.t4 VSUBS 0.225003f
C769 VDD1.t1 VSUBS 0.225003f
C770 VDD1.n6 VSUBS 1.73378f
C771 VDD1.n7 VSUBS 2.84502f
C772 VTAIL.t0 VSUBS 0.250042f
C773 VTAIL.t2 VSUBS 0.250042f
C774 VTAIL.n0 VSUBS 1.7808f
C775 VTAIL.n1 VSUBS 0.830558f
C776 VTAIL.t16 VSUBS 2.35859f
C777 VTAIL.n2 VSUBS 0.959289f
C778 VTAIL.t11 VSUBS 0.250042f
C779 VTAIL.t9 VSUBS 0.250042f
C780 VTAIL.n3 VSUBS 1.7808f
C781 VTAIL.n4 VSUBS 0.871807f
C782 VTAIL.t14 VSUBS 0.250042f
C783 VTAIL.t18 VSUBS 0.250042f
C784 VTAIL.n5 VSUBS 1.7808f
C785 VTAIL.n6 VSUBS 2.25845f
C786 VTAIL.t3 VSUBS 0.250042f
C787 VTAIL.t1 VSUBS 0.250042f
C788 VTAIL.n7 VSUBS 1.7808f
C789 VTAIL.n8 VSUBS 2.25844f
C790 VTAIL.t7 VSUBS 0.250042f
C791 VTAIL.t19 VSUBS 0.250042f
C792 VTAIL.n9 VSUBS 1.7808f
C793 VTAIL.n10 VSUBS 0.8718f
C794 VTAIL.t8 VSUBS 2.35861f
C795 VTAIL.n11 VSUBS 0.959272f
C796 VTAIL.t15 VSUBS 0.250042f
C797 VTAIL.t12 VSUBS 0.250042f
C798 VTAIL.n12 VSUBS 1.7808f
C799 VTAIL.n13 VSUBS 0.855141f
C800 VTAIL.t13 VSUBS 0.250042f
C801 VTAIL.t10 VSUBS 0.250042f
C802 VTAIL.n14 VSUBS 1.7808f
C803 VTAIL.n15 VSUBS 0.8718f
C804 VTAIL.t17 VSUBS 2.35859f
C805 VTAIL.n16 VSUBS 2.2428f
C806 VTAIL.t5 VSUBS 2.35859f
C807 VTAIL.n17 VSUBS 2.2428f
C808 VTAIL.t4 VSUBS 0.250042f
C809 VTAIL.t6 VSUBS 0.250042f
C810 VTAIL.n18 VSUBS 1.7808f
C811 VTAIL.n19 VSUBS 0.776616f
C812 VP.n0 VSUBS 0.043717f
C813 VP.t1 VSUBS 1.55363f
C814 VP.n1 VSUBS 0.066204f
C815 VP.n2 VSUBS 0.043717f
C816 VP.t6 VSUBS 1.55363f
C817 VP.n3 VSUBS 0.573961f
C818 VP.n4 VSUBS 0.043717f
C819 VP.t4 VSUBS 1.55363f
C820 VP.n5 VSUBS 0.573961f
C821 VP.n6 VSUBS 0.043717f
C822 VP.t2 VSUBS 1.55363f
C823 VP.n7 VSUBS 0.645978f
C824 VP.n8 VSUBS 0.043717f
C825 VP.t8 VSUBS 1.55363f
C826 VP.n9 VSUBS 0.066204f
C827 VP.n10 VSUBS 0.043717f
C828 VP.t9 VSUBS 1.55363f
C829 VP.n11 VSUBS 0.573961f
C830 VP.n12 VSUBS 0.043717f
C831 VP.t7 VSUBS 1.55363f
C832 VP.n13 VSUBS 0.638563f
C833 VP.t0 VSUBS 1.63786f
C834 VP.n14 VSUBS 0.668291f
C835 VP.n15 VSUBS 0.22737f
C836 VP.n16 VSUBS 0.066996f
C837 VP.n17 VSUBS 0.035323f
C838 VP.n18 VSUBS 0.066629f
C839 VP.n19 VSUBS 0.043717f
C840 VP.n20 VSUBS 0.043717f
C841 VP.n21 VSUBS 0.066629f
C842 VP.n22 VSUBS 0.035323f
C843 VP.t5 VSUBS 1.55363f
C844 VP.n23 VSUBS 0.573961f
C845 VP.n24 VSUBS 0.066996f
C846 VP.n25 VSUBS 0.043717f
C847 VP.n26 VSUBS 0.043717f
C848 VP.n27 VSUBS 0.043717f
C849 VP.n28 VSUBS 0.035434f
C850 VP.n29 VSUBS 0.067309f
C851 VP.n30 VSUBS 0.645978f
C852 VP.n31 VSUBS 1.99526f
C853 VP.n32 VSUBS 2.0306f
C854 VP.n33 VSUBS 0.043717f
C855 VP.n34 VSUBS 0.067309f
C856 VP.n35 VSUBS 0.035434f
C857 VP.n36 VSUBS 0.066204f
C858 VP.n37 VSUBS 0.043717f
C859 VP.n38 VSUBS 0.043717f
C860 VP.n39 VSUBS 0.066996f
C861 VP.n40 VSUBS 0.035323f
C862 VP.n41 VSUBS 0.066629f
C863 VP.n42 VSUBS 0.043717f
C864 VP.n43 VSUBS 0.043717f
C865 VP.n44 VSUBS 0.066629f
C866 VP.n45 VSUBS 0.035323f
C867 VP.t3 VSUBS 1.55363f
C868 VP.n46 VSUBS 0.573961f
C869 VP.n47 VSUBS 0.066996f
C870 VP.n48 VSUBS 0.043717f
C871 VP.n49 VSUBS 0.043717f
C872 VP.n50 VSUBS 0.043717f
C873 VP.n51 VSUBS 0.035434f
C874 VP.n52 VSUBS 0.067309f
C875 VP.n53 VSUBS 0.645978f
C876 VP.n54 VSUBS 0.03893f
.ends

