* NGSPICE file created from diff_pair_sample_0603.ext - technology: sky130A

.subckt diff_pair_sample_0603 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=1.15
X1 VTAIL.t7 VN.t0 VDD2.t0 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0.49335 ps=3.32 w=2.99 l=1.15
X2 B.t8 B.t6 B.t7 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=1.15
X3 B.t5 B.t3 B.t4 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=1.15
X4 VDD2.t1 VN.t1 VTAIL.t6 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=1.1661 ps=6.76 w=2.99 l=1.15
X5 VDD1.t3 VP.t0 VTAIL.t2 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=1.1661 ps=6.76 w=2.99 l=1.15
X6 VDD2.t2 VN.t2 VTAIL.t5 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=1.1661 ps=6.76 w=2.99 l=1.15
X7 VDD1.t2 VP.t1 VTAIL.t3 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=0.49335 pd=3.32 as=1.1661 ps=6.76 w=2.99 l=1.15
X8 VTAIL.t1 VP.t2 VDD1.t1 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0.49335 ps=3.32 w=2.99 l=1.15
X9 B.t2 B.t0 B.t1 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0 ps=0 w=2.99 l=1.15
X10 VTAIL.t4 VN.t3 VDD2.t3 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0.49335 ps=3.32 w=2.99 l=1.15
X11 VTAIL.t0 VP.t3 VDD1.t0 w_n1858_n1566# sky130_fd_pr__pfet_01v8 ad=1.1661 pd=6.76 as=0.49335 ps=3.32 w=2.99 l=1.15
R0 B.n250 B.n249 585
R1 B.n251 B.n36 585
R2 B.n253 B.n252 585
R3 B.n254 B.n35 585
R4 B.n256 B.n255 585
R5 B.n257 B.n34 585
R6 B.n259 B.n258 585
R7 B.n260 B.n33 585
R8 B.n262 B.n261 585
R9 B.n263 B.n32 585
R10 B.n265 B.n264 585
R11 B.n266 B.n31 585
R12 B.n268 B.n267 585
R13 B.n269 B.n30 585
R14 B.n271 B.n270 585
R15 B.n273 B.n27 585
R16 B.n275 B.n274 585
R17 B.n276 B.n26 585
R18 B.n278 B.n277 585
R19 B.n279 B.n25 585
R20 B.n281 B.n280 585
R21 B.n282 B.n24 585
R22 B.n284 B.n283 585
R23 B.n285 B.n23 585
R24 B.n287 B.n286 585
R25 B.n289 B.n288 585
R26 B.n290 B.n19 585
R27 B.n292 B.n291 585
R28 B.n293 B.n18 585
R29 B.n295 B.n294 585
R30 B.n296 B.n17 585
R31 B.n298 B.n297 585
R32 B.n299 B.n16 585
R33 B.n301 B.n300 585
R34 B.n302 B.n15 585
R35 B.n304 B.n303 585
R36 B.n305 B.n14 585
R37 B.n307 B.n306 585
R38 B.n308 B.n13 585
R39 B.n310 B.n309 585
R40 B.n248 B.n37 585
R41 B.n247 B.n246 585
R42 B.n245 B.n38 585
R43 B.n244 B.n243 585
R44 B.n242 B.n39 585
R45 B.n241 B.n240 585
R46 B.n239 B.n40 585
R47 B.n238 B.n237 585
R48 B.n236 B.n41 585
R49 B.n235 B.n234 585
R50 B.n233 B.n42 585
R51 B.n232 B.n231 585
R52 B.n230 B.n43 585
R53 B.n229 B.n228 585
R54 B.n227 B.n44 585
R55 B.n226 B.n225 585
R56 B.n224 B.n45 585
R57 B.n223 B.n222 585
R58 B.n221 B.n46 585
R59 B.n220 B.n219 585
R60 B.n218 B.n47 585
R61 B.n217 B.n216 585
R62 B.n215 B.n48 585
R63 B.n214 B.n213 585
R64 B.n212 B.n49 585
R65 B.n211 B.n210 585
R66 B.n209 B.n50 585
R67 B.n208 B.n207 585
R68 B.n206 B.n51 585
R69 B.n205 B.n204 585
R70 B.n203 B.n52 585
R71 B.n202 B.n201 585
R72 B.n200 B.n53 585
R73 B.n199 B.n198 585
R74 B.n197 B.n54 585
R75 B.n196 B.n195 585
R76 B.n194 B.n55 585
R77 B.n193 B.n192 585
R78 B.n191 B.n56 585
R79 B.n190 B.n189 585
R80 B.n188 B.n57 585
R81 B.n187 B.n186 585
R82 B.n185 B.n58 585
R83 B.n124 B.n123 585
R84 B.n125 B.n82 585
R85 B.n127 B.n126 585
R86 B.n128 B.n81 585
R87 B.n130 B.n129 585
R88 B.n131 B.n80 585
R89 B.n133 B.n132 585
R90 B.n134 B.n79 585
R91 B.n136 B.n135 585
R92 B.n137 B.n78 585
R93 B.n139 B.n138 585
R94 B.n140 B.n77 585
R95 B.n142 B.n141 585
R96 B.n143 B.n76 585
R97 B.n145 B.n144 585
R98 B.n147 B.n73 585
R99 B.n149 B.n148 585
R100 B.n150 B.n72 585
R101 B.n152 B.n151 585
R102 B.n153 B.n71 585
R103 B.n155 B.n154 585
R104 B.n156 B.n70 585
R105 B.n158 B.n157 585
R106 B.n159 B.n69 585
R107 B.n161 B.n160 585
R108 B.n163 B.n162 585
R109 B.n164 B.n65 585
R110 B.n166 B.n165 585
R111 B.n167 B.n64 585
R112 B.n169 B.n168 585
R113 B.n170 B.n63 585
R114 B.n172 B.n171 585
R115 B.n173 B.n62 585
R116 B.n175 B.n174 585
R117 B.n176 B.n61 585
R118 B.n178 B.n177 585
R119 B.n179 B.n60 585
R120 B.n181 B.n180 585
R121 B.n182 B.n59 585
R122 B.n184 B.n183 585
R123 B.n122 B.n83 585
R124 B.n121 B.n120 585
R125 B.n119 B.n84 585
R126 B.n118 B.n117 585
R127 B.n116 B.n85 585
R128 B.n115 B.n114 585
R129 B.n113 B.n86 585
R130 B.n112 B.n111 585
R131 B.n110 B.n87 585
R132 B.n109 B.n108 585
R133 B.n107 B.n88 585
R134 B.n106 B.n105 585
R135 B.n104 B.n89 585
R136 B.n103 B.n102 585
R137 B.n101 B.n90 585
R138 B.n100 B.n99 585
R139 B.n98 B.n91 585
R140 B.n97 B.n96 585
R141 B.n95 B.n92 585
R142 B.n94 B.n93 585
R143 B.n2 B.n0 585
R144 B.n341 B.n1 585
R145 B.n340 B.n339 585
R146 B.n338 B.n3 585
R147 B.n337 B.n336 585
R148 B.n335 B.n4 585
R149 B.n334 B.n333 585
R150 B.n332 B.n5 585
R151 B.n331 B.n330 585
R152 B.n329 B.n6 585
R153 B.n328 B.n327 585
R154 B.n326 B.n7 585
R155 B.n325 B.n324 585
R156 B.n323 B.n8 585
R157 B.n322 B.n321 585
R158 B.n320 B.n9 585
R159 B.n319 B.n318 585
R160 B.n317 B.n10 585
R161 B.n316 B.n315 585
R162 B.n314 B.n11 585
R163 B.n313 B.n312 585
R164 B.n311 B.n12 585
R165 B.n343 B.n342 585
R166 B.n124 B.n83 511.721
R167 B.n311 B.n310 511.721
R168 B.n185 B.n184 511.721
R169 B.n250 B.n37 511.721
R170 B.n66 B.t6 266.509
R171 B.n74 B.t0 266.509
R172 B.n20 B.t3 266.509
R173 B.n28 B.t9 266.509
R174 B.n66 B.t8 173.768
R175 B.n28 B.t10 173.768
R176 B.n74 B.t2 173.767
R177 B.n20 B.t4 173.767
R178 B.n120 B.n83 163.367
R179 B.n120 B.n119 163.367
R180 B.n119 B.n118 163.367
R181 B.n118 B.n85 163.367
R182 B.n114 B.n85 163.367
R183 B.n114 B.n113 163.367
R184 B.n113 B.n112 163.367
R185 B.n112 B.n87 163.367
R186 B.n108 B.n87 163.367
R187 B.n108 B.n107 163.367
R188 B.n107 B.n106 163.367
R189 B.n106 B.n89 163.367
R190 B.n102 B.n89 163.367
R191 B.n102 B.n101 163.367
R192 B.n101 B.n100 163.367
R193 B.n100 B.n91 163.367
R194 B.n96 B.n91 163.367
R195 B.n96 B.n95 163.367
R196 B.n95 B.n94 163.367
R197 B.n94 B.n2 163.367
R198 B.n342 B.n2 163.367
R199 B.n342 B.n341 163.367
R200 B.n341 B.n340 163.367
R201 B.n340 B.n3 163.367
R202 B.n336 B.n3 163.367
R203 B.n336 B.n335 163.367
R204 B.n335 B.n334 163.367
R205 B.n334 B.n5 163.367
R206 B.n330 B.n5 163.367
R207 B.n330 B.n329 163.367
R208 B.n329 B.n328 163.367
R209 B.n328 B.n7 163.367
R210 B.n324 B.n7 163.367
R211 B.n324 B.n323 163.367
R212 B.n323 B.n322 163.367
R213 B.n322 B.n9 163.367
R214 B.n318 B.n9 163.367
R215 B.n318 B.n317 163.367
R216 B.n317 B.n316 163.367
R217 B.n316 B.n11 163.367
R218 B.n312 B.n11 163.367
R219 B.n312 B.n311 163.367
R220 B.n125 B.n124 163.367
R221 B.n126 B.n125 163.367
R222 B.n126 B.n81 163.367
R223 B.n130 B.n81 163.367
R224 B.n131 B.n130 163.367
R225 B.n132 B.n131 163.367
R226 B.n132 B.n79 163.367
R227 B.n136 B.n79 163.367
R228 B.n137 B.n136 163.367
R229 B.n138 B.n137 163.367
R230 B.n138 B.n77 163.367
R231 B.n142 B.n77 163.367
R232 B.n143 B.n142 163.367
R233 B.n144 B.n143 163.367
R234 B.n144 B.n73 163.367
R235 B.n149 B.n73 163.367
R236 B.n150 B.n149 163.367
R237 B.n151 B.n150 163.367
R238 B.n151 B.n71 163.367
R239 B.n155 B.n71 163.367
R240 B.n156 B.n155 163.367
R241 B.n157 B.n156 163.367
R242 B.n157 B.n69 163.367
R243 B.n161 B.n69 163.367
R244 B.n162 B.n161 163.367
R245 B.n162 B.n65 163.367
R246 B.n166 B.n65 163.367
R247 B.n167 B.n166 163.367
R248 B.n168 B.n167 163.367
R249 B.n168 B.n63 163.367
R250 B.n172 B.n63 163.367
R251 B.n173 B.n172 163.367
R252 B.n174 B.n173 163.367
R253 B.n174 B.n61 163.367
R254 B.n178 B.n61 163.367
R255 B.n179 B.n178 163.367
R256 B.n180 B.n179 163.367
R257 B.n180 B.n59 163.367
R258 B.n184 B.n59 163.367
R259 B.n186 B.n185 163.367
R260 B.n186 B.n57 163.367
R261 B.n190 B.n57 163.367
R262 B.n191 B.n190 163.367
R263 B.n192 B.n191 163.367
R264 B.n192 B.n55 163.367
R265 B.n196 B.n55 163.367
R266 B.n197 B.n196 163.367
R267 B.n198 B.n197 163.367
R268 B.n198 B.n53 163.367
R269 B.n202 B.n53 163.367
R270 B.n203 B.n202 163.367
R271 B.n204 B.n203 163.367
R272 B.n204 B.n51 163.367
R273 B.n208 B.n51 163.367
R274 B.n209 B.n208 163.367
R275 B.n210 B.n209 163.367
R276 B.n210 B.n49 163.367
R277 B.n214 B.n49 163.367
R278 B.n215 B.n214 163.367
R279 B.n216 B.n215 163.367
R280 B.n216 B.n47 163.367
R281 B.n220 B.n47 163.367
R282 B.n221 B.n220 163.367
R283 B.n222 B.n221 163.367
R284 B.n222 B.n45 163.367
R285 B.n226 B.n45 163.367
R286 B.n227 B.n226 163.367
R287 B.n228 B.n227 163.367
R288 B.n228 B.n43 163.367
R289 B.n232 B.n43 163.367
R290 B.n233 B.n232 163.367
R291 B.n234 B.n233 163.367
R292 B.n234 B.n41 163.367
R293 B.n238 B.n41 163.367
R294 B.n239 B.n238 163.367
R295 B.n240 B.n239 163.367
R296 B.n240 B.n39 163.367
R297 B.n244 B.n39 163.367
R298 B.n245 B.n244 163.367
R299 B.n246 B.n245 163.367
R300 B.n246 B.n37 163.367
R301 B.n310 B.n13 163.367
R302 B.n306 B.n13 163.367
R303 B.n306 B.n305 163.367
R304 B.n305 B.n304 163.367
R305 B.n304 B.n15 163.367
R306 B.n300 B.n15 163.367
R307 B.n300 B.n299 163.367
R308 B.n299 B.n298 163.367
R309 B.n298 B.n17 163.367
R310 B.n294 B.n17 163.367
R311 B.n294 B.n293 163.367
R312 B.n293 B.n292 163.367
R313 B.n292 B.n19 163.367
R314 B.n288 B.n19 163.367
R315 B.n288 B.n287 163.367
R316 B.n287 B.n23 163.367
R317 B.n283 B.n23 163.367
R318 B.n283 B.n282 163.367
R319 B.n282 B.n281 163.367
R320 B.n281 B.n25 163.367
R321 B.n277 B.n25 163.367
R322 B.n277 B.n276 163.367
R323 B.n276 B.n275 163.367
R324 B.n275 B.n27 163.367
R325 B.n270 B.n27 163.367
R326 B.n270 B.n269 163.367
R327 B.n269 B.n268 163.367
R328 B.n268 B.n31 163.367
R329 B.n264 B.n31 163.367
R330 B.n264 B.n263 163.367
R331 B.n263 B.n262 163.367
R332 B.n262 B.n33 163.367
R333 B.n258 B.n33 163.367
R334 B.n258 B.n257 163.367
R335 B.n257 B.n256 163.367
R336 B.n256 B.n35 163.367
R337 B.n252 B.n35 163.367
R338 B.n252 B.n251 163.367
R339 B.n251 B.n250 163.367
R340 B.n67 B.t7 145.065
R341 B.n29 B.t11 145.065
R342 B.n75 B.t1 145.064
R343 B.n21 B.t5 145.064
R344 B.n68 B.n67 59.5399
R345 B.n146 B.n75 59.5399
R346 B.n22 B.n21 59.5399
R347 B.n272 B.n29 59.5399
R348 B.n309 B.n12 33.2493
R349 B.n249 B.n248 33.2493
R350 B.n183 B.n58 33.2493
R351 B.n123 B.n122 33.2493
R352 B.n67 B.n66 28.7035
R353 B.n75 B.n74 28.7035
R354 B.n21 B.n20 28.7035
R355 B.n29 B.n28 28.7035
R356 B B.n343 18.0485
R357 B.n309 B.n308 10.6151
R358 B.n308 B.n307 10.6151
R359 B.n307 B.n14 10.6151
R360 B.n303 B.n14 10.6151
R361 B.n303 B.n302 10.6151
R362 B.n302 B.n301 10.6151
R363 B.n301 B.n16 10.6151
R364 B.n297 B.n16 10.6151
R365 B.n297 B.n296 10.6151
R366 B.n296 B.n295 10.6151
R367 B.n295 B.n18 10.6151
R368 B.n291 B.n18 10.6151
R369 B.n291 B.n290 10.6151
R370 B.n290 B.n289 10.6151
R371 B.n286 B.n285 10.6151
R372 B.n285 B.n284 10.6151
R373 B.n284 B.n24 10.6151
R374 B.n280 B.n24 10.6151
R375 B.n280 B.n279 10.6151
R376 B.n279 B.n278 10.6151
R377 B.n278 B.n26 10.6151
R378 B.n274 B.n26 10.6151
R379 B.n274 B.n273 10.6151
R380 B.n271 B.n30 10.6151
R381 B.n267 B.n30 10.6151
R382 B.n267 B.n266 10.6151
R383 B.n266 B.n265 10.6151
R384 B.n265 B.n32 10.6151
R385 B.n261 B.n32 10.6151
R386 B.n261 B.n260 10.6151
R387 B.n260 B.n259 10.6151
R388 B.n259 B.n34 10.6151
R389 B.n255 B.n34 10.6151
R390 B.n255 B.n254 10.6151
R391 B.n254 B.n253 10.6151
R392 B.n253 B.n36 10.6151
R393 B.n249 B.n36 10.6151
R394 B.n187 B.n58 10.6151
R395 B.n188 B.n187 10.6151
R396 B.n189 B.n188 10.6151
R397 B.n189 B.n56 10.6151
R398 B.n193 B.n56 10.6151
R399 B.n194 B.n193 10.6151
R400 B.n195 B.n194 10.6151
R401 B.n195 B.n54 10.6151
R402 B.n199 B.n54 10.6151
R403 B.n200 B.n199 10.6151
R404 B.n201 B.n200 10.6151
R405 B.n201 B.n52 10.6151
R406 B.n205 B.n52 10.6151
R407 B.n206 B.n205 10.6151
R408 B.n207 B.n206 10.6151
R409 B.n207 B.n50 10.6151
R410 B.n211 B.n50 10.6151
R411 B.n212 B.n211 10.6151
R412 B.n213 B.n212 10.6151
R413 B.n213 B.n48 10.6151
R414 B.n217 B.n48 10.6151
R415 B.n218 B.n217 10.6151
R416 B.n219 B.n218 10.6151
R417 B.n219 B.n46 10.6151
R418 B.n223 B.n46 10.6151
R419 B.n224 B.n223 10.6151
R420 B.n225 B.n224 10.6151
R421 B.n225 B.n44 10.6151
R422 B.n229 B.n44 10.6151
R423 B.n230 B.n229 10.6151
R424 B.n231 B.n230 10.6151
R425 B.n231 B.n42 10.6151
R426 B.n235 B.n42 10.6151
R427 B.n236 B.n235 10.6151
R428 B.n237 B.n236 10.6151
R429 B.n237 B.n40 10.6151
R430 B.n241 B.n40 10.6151
R431 B.n242 B.n241 10.6151
R432 B.n243 B.n242 10.6151
R433 B.n243 B.n38 10.6151
R434 B.n247 B.n38 10.6151
R435 B.n248 B.n247 10.6151
R436 B.n123 B.n82 10.6151
R437 B.n127 B.n82 10.6151
R438 B.n128 B.n127 10.6151
R439 B.n129 B.n128 10.6151
R440 B.n129 B.n80 10.6151
R441 B.n133 B.n80 10.6151
R442 B.n134 B.n133 10.6151
R443 B.n135 B.n134 10.6151
R444 B.n135 B.n78 10.6151
R445 B.n139 B.n78 10.6151
R446 B.n140 B.n139 10.6151
R447 B.n141 B.n140 10.6151
R448 B.n141 B.n76 10.6151
R449 B.n145 B.n76 10.6151
R450 B.n148 B.n147 10.6151
R451 B.n148 B.n72 10.6151
R452 B.n152 B.n72 10.6151
R453 B.n153 B.n152 10.6151
R454 B.n154 B.n153 10.6151
R455 B.n154 B.n70 10.6151
R456 B.n158 B.n70 10.6151
R457 B.n159 B.n158 10.6151
R458 B.n160 B.n159 10.6151
R459 B.n164 B.n163 10.6151
R460 B.n165 B.n164 10.6151
R461 B.n165 B.n64 10.6151
R462 B.n169 B.n64 10.6151
R463 B.n170 B.n169 10.6151
R464 B.n171 B.n170 10.6151
R465 B.n171 B.n62 10.6151
R466 B.n175 B.n62 10.6151
R467 B.n176 B.n175 10.6151
R468 B.n177 B.n176 10.6151
R469 B.n177 B.n60 10.6151
R470 B.n181 B.n60 10.6151
R471 B.n182 B.n181 10.6151
R472 B.n183 B.n182 10.6151
R473 B.n122 B.n121 10.6151
R474 B.n121 B.n84 10.6151
R475 B.n117 B.n84 10.6151
R476 B.n117 B.n116 10.6151
R477 B.n116 B.n115 10.6151
R478 B.n115 B.n86 10.6151
R479 B.n111 B.n86 10.6151
R480 B.n111 B.n110 10.6151
R481 B.n110 B.n109 10.6151
R482 B.n109 B.n88 10.6151
R483 B.n105 B.n88 10.6151
R484 B.n105 B.n104 10.6151
R485 B.n104 B.n103 10.6151
R486 B.n103 B.n90 10.6151
R487 B.n99 B.n90 10.6151
R488 B.n99 B.n98 10.6151
R489 B.n98 B.n97 10.6151
R490 B.n97 B.n92 10.6151
R491 B.n93 B.n92 10.6151
R492 B.n93 B.n0 10.6151
R493 B.n339 B.n1 10.6151
R494 B.n339 B.n338 10.6151
R495 B.n338 B.n337 10.6151
R496 B.n337 B.n4 10.6151
R497 B.n333 B.n4 10.6151
R498 B.n333 B.n332 10.6151
R499 B.n332 B.n331 10.6151
R500 B.n331 B.n6 10.6151
R501 B.n327 B.n6 10.6151
R502 B.n327 B.n326 10.6151
R503 B.n326 B.n325 10.6151
R504 B.n325 B.n8 10.6151
R505 B.n321 B.n8 10.6151
R506 B.n321 B.n320 10.6151
R507 B.n320 B.n319 10.6151
R508 B.n319 B.n10 10.6151
R509 B.n315 B.n10 10.6151
R510 B.n315 B.n314 10.6151
R511 B.n314 B.n313 10.6151
R512 B.n313 B.n12 10.6151
R513 B.n289 B.n22 9.36635
R514 B.n272 B.n271 9.36635
R515 B.n146 B.n145 9.36635
R516 B.n163 B.n68 9.36635
R517 B.n343 B.n0 2.81026
R518 B.n343 B.n1 2.81026
R519 B.n286 B.n22 1.24928
R520 B.n273 B.n272 1.24928
R521 B.n147 B.n146 1.24928
R522 B.n160 B.n68 1.24928
R523 VN.n0 VN.t0 97.9935
R524 VN.n1 VN.t2 97.9935
R525 VN.n0 VN.t1 97.7783
R526 VN.n1 VN.t3 97.7783
R527 VN VN.n1 54.0096
R528 VN VN.n0 18.771
R529 VDD2.n2 VDD2.n0 172.65
R530 VDD2.n2 VDD2.n1 142.53
R531 VDD2.n1 VDD2.t3 10.8717
R532 VDD2.n1 VDD2.t2 10.8717
R533 VDD2.n0 VDD2.t0 10.8717
R534 VDD2.n0 VDD2.t1 10.8717
R535 VDD2 VDD2.n2 0.0586897
R536 VTAIL.n5 VTAIL.t0 136.724
R537 VTAIL.n4 VTAIL.t5 136.724
R538 VTAIL.n3 VTAIL.t4 136.724
R539 VTAIL.n6 VTAIL.t2 136.722
R540 VTAIL.n7 VTAIL.t6 136.722
R541 VTAIL.n0 VTAIL.t7 136.722
R542 VTAIL.n1 VTAIL.t3 136.722
R543 VTAIL.n2 VTAIL.t1 136.722
R544 VTAIL.n7 VTAIL.n6 16.2203
R545 VTAIL.n3 VTAIL.n2 16.2203
R546 VTAIL.n4 VTAIL.n3 1.27636
R547 VTAIL.n6 VTAIL.n5 1.27636
R548 VTAIL.n2 VTAIL.n1 1.27636
R549 VTAIL VTAIL.n0 0.696621
R550 VTAIL VTAIL.n7 0.580241
R551 VTAIL.n5 VTAIL.n4 0.470328
R552 VTAIL.n1 VTAIL.n0 0.470328
R553 VP.n4 VP.n3 174.024
R554 VP.n10 VP.n9 174.024
R555 VP.n8 VP.n0 161.3
R556 VP.n7 VP.n6 161.3
R557 VP.n5 VP.n1 161.3
R558 VP.n2 VP.t3 97.9935
R559 VP.n2 VP.t0 97.7783
R560 VP.n3 VP.t2 62.6605
R561 VP.n9 VP.t1 62.6605
R562 VP.n4 VP.n2 53.6289
R563 VP.n7 VP.n1 40.4934
R564 VP.n8 VP.n7 40.4934
R565 VP.n3 VP.n1 11.7447
R566 VP.n9 VP.n8 11.7447
R567 VP.n5 VP.n4 0.189894
R568 VP.n6 VP.n5 0.189894
R569 VP.n6 VP.n0 0.189894
R570 VP.n10 VP.n0 0.189894
R571 VP VP.n10 0.0516364
R572 VDD1 VDD1.n1 173.175
R573 VDD1 VDD1.n0 142.589
R574 VDD1.n0 VDD1.t0 10.8717
R575 VDD1.n0 VDD1.t3 10.8717
R576 VDD1.n1 VDD1.t1 10.8717
R577 VDD1.n1 VDD1.t2 10.8717
C0 VDD1 VDD2 0.672372f
C1 VDD2 VP 0.30727f
C2 VDD2 w_n1858_n1566# 0.938548f
C3 B VTAIL 1.51315f
C4 VN B 0.720229f
C5 VDD1 B 0.762355f
C6 VP B 1.10333f
C7 B w_n1858_n1566# 4.93479f
C8 VN VTAIL 1.33595f
C9 VDD1 VTAIL 2.74343f
C10 VP VTAIL 1.35005f
C11 VTAIL w_n1858_n1566# 1.8239f
C12 VDD1 VN 0.152408f
C13 VN VP 3.488f
C14 VDD2 B 0.791007f
C15 VDD1 VP 1.34285f
C16 VN w_n1858_n1566# 2.70599f
C17 VDD1 w_n1858_n1566# 0.91507f
C18 VP w_n1858_n1566# 2.93883f
C19 VDD2 VTAIL 2.78792f
C20 VDD2 VN 1.1889f
C21 VDD2 VSUBS 0.475608f
C22 VDD1 VSUBS 2.589143f
C23 VTAIL VSUBS 0.374695f
C24 VN VSUBS 3.98627f
C25 VP VSUBS 1.068554f
C26 B VSUBS 2.14356f
C27 w_n1858_n1566# VSUBS 36.8553f
C28 VDD1.t0 VSUBS 0.042524f
C29 VDD1.t3 VSUBS 0.042524f
C30 VDD1.n0 VSUBS 0.22205f
C31 VDD1.t1 VSUBS 0.042524f
C32 VDD1.t2 VSUBS 0.042524f
C33 VDD1.n1 VSUBS 0.361708f
C34 VP.n0 VSUBS 0.047917f
C35 VP.t1 VSUBS 0.410268f
C36 VP.n1 VSUBS 0.072308f
C37 VP.t3 VSUBS 0.533742f
C38 VP.t0 VSUBS 0.532932f
C39 VP.n2 VSUBS 1.54126f
C40 VP.t2 VSUBS 0.410268f
C41 VP.n3 VSUBS 0.271792f
C42 VP.n4 VSUBS 2.04326f
C43 VP.n5 VSUBS 0.047917f
C44 VP.n6 VSUBS 0.047917f
C45 VP.n7 VSUBS 0.038737f
C46 VP.n8 VSUBS 0.072308f
C47 VP.n9 VSUBS 0.271792f
C48 VP.n10 VSUBS 0.042954f
C49 VTAIL.t7 VSUBS 0.228464f
C50 VTAIL.n0 VSUBS 0.256835f
C51 VTAIL.t3 VSUBS 0.228464f
C52 VTAIL.n1 VSUBS 0.283602f
C53 VTAIL.t1 VSUBS 0.228464f
C54 VTAIL.n2 VSUBS 0.634469f
C55 VTAIL.t4 VSUBS 0.228465f
C56 VTAIL.n3 VSUBS 0.634468f
C57 VTAIL.t5 VSUBS 0.228465f
C58 VTAIL.n4 VSUBS 0.283602f
C59 VTAIL.t0 VSUBS 0.228465f
C60 VTAIL.n5 VSUBS 0.283602f
C61 VTAIL.t2 VSUBS 0.228464f
C62 VTAIL.n6 VSUBS 0.634469f
C63 VTAIL.t6 VSUBS 0.228464f
C64 VTAIL.n7 VSUBS 0.602328f
C65 VDD2.t0 VSUBS 0.045212f
C66 VDD2.t1 VSUBS 0.045212f
C67 VDD2.n0 VSUBS 0.37561f
C68 VDD2.t3 VSUBS 0.045212f
C69 VDD2.t2 VSUBS 0.045212f
C70 VDD2.n1 VSUBS 0.235951f
C71 VDD2.n2 VSUBS 1.92481f
C72 VN.t0 VSUBS 0.511677f
C73 VN.t1 VSUBS 0.510901f
C74 VN.n0 VSUBS 0.463803f
C75 VN.t2 VSUBS 0.511677f
C76 VN.t3 VSUBS 0.510901f
C77 VN.n1 VSUBS 1.50133f
C78 B.n0 VSUBS 0.005031f
C79 B.n1 VSUBS 0.005031f
C80 B.n2 VSUBS 0.007956f
C81 B.n3 VSUBS 0.007956f
C82 B.n4 VSUBS 0.007956f
C83 B.n5 VSUBS 0.007956f
C84 B.n6 VSUBS 0.007956f
C85 B.n7 VSUBS 0.007956f
C86 B.n8 VSUBS 0.007956f
C87 B.n9 VSUBS 0.007956f
C88 B.n10 VSUBS 0.007956f
C89 B.n11 VSUBS 0.007956f
C90 B.n12 VSUBS 0.018196f
C91 B.n13 VSUBS 0.007956f
C92 B.n14 VSUBS 0.007956f
C93 B.n15 VSUBS 0.007956f
C94 B.n16 VSUBS 0.007956f
C95 B.n17 VSUBS 0.007956f
C96 B.n18 VSUBS 0.007956f
C97 B.n19 VSUBS 0.007956f
C98 B.t5 VSUBS 0.081501f
C99 B.t4 VSUBS 0.090777f
C100 B.t3 VSUBS 0.184236f
C101 B.n20 VSUBS 0.079053f
C102 B.n21 VSUBS 0.067505f
C103 B.n22 VSUBS 0.018434f
C104 B.n23 VSUBS 0.007956f
C105 B.n24 VSUBS 0.007956f
C106 B.n25 VSUBS 0.007956f
C107 B.n26 VSUBS 0.007956f
C108 B.n27 VSUBS 0.007956f
C109 B.t11 VSUBS 0.081501f
C110 B.t10 VSUBS 0.090777f
C111 B.t9 VSUBS 0.184236f
C112 B.n28 VSUBS 0.079053f
C113 B.n29 VSUBS 0.067505f
C114 B.n30 VSUBS 0.007956f
C115 B.n31 VSUBS 0.007956f
C116 B.n32 VSUBS 0.007956f
C117 B.n33 VSUBS 0.007956f
C118 B.n34 VSUBS 0.007956f
C119 B.n35 VSUBS 0.007956f
C120 B.n36 VSUBS 0.007956f
C121 B.n37 VSUBS 0.018196f
C122 B.n38 VSUBS 0.007956f
C123 B.n39 VSUBS 0.007956f
C124 B.n40 VSUBS 0.007956f
C125 B.n41 VSUBS 0.007956f
C126 B.n42 VSUBS 0.007956f
C127 B.n43 VSUBS 0.007956f
C128 B.n44 VSUBS 0.007956f
C129 B.n45 VSUBS 0.007956f
C130 B.n46 VSUBS 0.007956f
C131 B.n47 VSUBS 0.007956f
C132 B.n48 VSUBS 0.007956f
C133 B.n49 VSUBS 0.007956f
C134 B.n50 VSUBS 0.007956f
C135 B.n51 VSUBS 0.007956f
C136 B.n52 VSUBS 0.007956f
C137 B.n53 VSUBS 0.007956f
C138 B.n54 VSUBS 0.007956f
C139 B.n55 VSUBS 0.007956f
C140 B.n56 VSUBS 0.007956f
C141 B.n57 VSUBS 0.007956f
C142 B.n58 VSUBS 0.018196f
C143 B.n59 VSUBS 0.007956f
C144 B.n60 VSUBS 0.007956f
C145 B.n61 VSUBS 0.007956f
C146 B.n62 VSUBS 0.007956f
C147 B.n63 VSUBS 0.007956f
C148 B.n64 VSUBS 0.007956f
C149 B.n65 VSUBS 0.007956f
C150 B.t7 VSUBS 0.081501f
C151 B.t8 VSUBS 0.090777f
C152 B.t6 VSUBS 0.184236f
C153 B.n66 VSUBS 0.079053f
C154 B.n67 VSUBS 0.067505f
C155 B.n68 VSUBS 0.018434f
C156 B.n69 VSUBS 0.007956f
C157 B.n70 VSUBS 0.007956f
C158 B.n71 VSUBS 0.007956f
C159 B.n72 VSUBS 0.007956f
C160 B.n73 VSUBS 0.007956f
C161 B.t1 VSUBS 0.081501f
C162 B.t2 VSUBS 0.090777f
C163 B.t0 VSUBS 0.184236f
C164 B.n74 VSUBS 0.079053f
C165 B.n75 VSUBS 0.067505f
C166 B.n76 VSUBS 0.007956f
C167 B.n77 VSUBS 0.007956f
C168 B.n78 VSUBS 0.007956f
C169 B.n79 VSUBS 0.007956f
C170 B.n80 VSUBS 0.007956f
C171 B.n81 VSUBS 0.007956f
C172 B.n82 VSUBS 0.007956f
C173 B.n83 VSUBS 0.018196f
C174 B.n84 VSUBS 0.007956f
C175 B.n85 VSUBS 0.007956f
C176 B.n86 VSUBS 0.007956f
C177 B.n87 VSUBS 0.007956f
C178 B.n88 VSUBS 0.007956f
C179 B.n89 VSUBS 0.007956f
C180 B.n90 VSUBS 0.007956f
C181 B.n91 VSUBS 0.007956f
C182 B.n92 VSUBS 0.007956f
C183 B.n93 VSUBS 0.007956f
C184 B.n94 VSUBS 0.007956f
C185 B.n95 VSUBS 0.007956f
C186 B.n96 VSUBS 0.007956f
C187 B.n97 VSUBS 0.007956f
C188 B.n98 VSUBS 0.007956f
C189 B.n99 VSUBS 0.007956f
C190 B.n100 VSUBS 0.007956f
C191 B.n101 VSUBS 0.007956f
C192 B.n102 VSUBS 0.007956f
C193 B.n103 VSUBS 0.007956f
C194 B.n104 VSUBS 0.007956f
C195 B.n105 VSUBS 0.007956f
C196 B.n106 VSUBS 0.007956f
C197 B.n107 VSUBS 0.007956f
C198 B.n108 VSUBS 0.007956f
C199 B.n109 VSUBS 0.007956f
C200 B.n110 VSUBS 0.007956f
C201 B.n111 VSUBS 0.007956f
C202 B.n112 VSUBS 0.007956f
C203 B.n113 VSUBS 0.007956f
C204 B.n114 VSUBS 0.007956f
C205 B.n115 VSUBS 0.007956f
C206 B.n116 VSUBS 0.007956f
C207 B.n117 VSUBS 0.007956f
C208 B.n118 VSUBS 0.007956f
C209 B.n119 VSUBS 0.007956f
C210 B.n120 VSUBS 0.007956f
C211 B.n121 VSUBS 0.007956f
C212 B.n122 VSUBS 0.018196f
C213 B.n123 VSUBS 0.01948f
C214 B.n124 VSUBS 0.01948f
C215 B.n125 VSUBS 0.007956f
C216 B.n126 VSUBS 0.007956f
C217 B.n127 VSUBS 0.007956f
C218 B.n128 VSUBS 0.007956f
C219 B.n129 VSUBS 0.007956f
C220 B.n130 VSUBS 0.007956f
C221 B.n131 VSUBS 0.007956f
C222 B.n132 VSUBS 0.007956f
C223 B.n133 VSUBS 0.007956f
C224 B.n134 VSUBS 0.007956f
C225 B.n135 VSUBS 0.007956f
C226 B.n136 VSUBS 0.007956f
C227 B.n137 VSUBS 0.007956f
C228 B.n138 VSUBS 0.007956f
C229 B.n139 VSUBS 0.007956f
C230 B.n140 VSUBS 0.007956f
C231 B.n141 VSUBS 0.007956f
C232 B.n142 VSUBS 0.007956f
C233 B.n143 VSUBS 0.007956f
C234 B.n144 VSUBS 0.007956f
C235 B.n145 VSUBS 0.007488f
C236 B.n146 VSUBS 0.018434f
C237 B.n147 VSUBS 0.004446f
C238 B.n148 VSUBS 0.007956f
C239 B.n149 VSUBS 0.007956f
C240 B.n150 VSUBS 0.007956f
C241 B.n151 VSUBS 0.007956f
C242 B.n152 VSUBS 0.007956f
C243 B.n153 VSUBS 0.007956f
C244 B.n154 VSUBS 0.007956f
C245 B.n155 VSUBS 0.007956f
C246 B.n156 VSUBS 0.007956f
C247 B.n157 VSUBS 0.007956f
C248 B.n158 VSUBS 0.007956f
C249 B.n159 VSUBS 0.007956f
C250 B.n160 VSUBS 0.004446f
C251 B.n161 VSUBS 0.007956f
C252 B.n162 VSUBS 0.007956f
C253 B.n163 VSUBS 0.007488f
C254 B.n164 VSUBS 0.007956f
C255 B.n165 VSUBS 0.007956f
C256 B.n166 VSUBS 0.007956f
C257 B.n167 VSUBS 0.007956f
C258 B.n168 VSUBS 0.007956f
C259 B.n169 VSUBS 0.007956f
C260 B.n170 VSUBS 0.007956f
C261 B.n171 VSUBS 0.007956f
C262 B.n172 VSUBS 0.007956f
C263 B.n173 VSUBS 0.007956f
C264 B.n174 VSUBS 0.007956f
C265 B.n175 VSUBS 0.007956f
C266 B.n176 VSUBS 0.007956f
C267 B.n177 VSUBS 0.007956f
C268 B.n178 VSUBS 0.007956f
C269 B.n179 VSUBS 0.007956f
C270 B.n180 VSUBS 0.007956f
C271 B.n181 VSUBS 0.007956f
C272 B.n182 VSUBS 0.007956f
C273 B.n183 VSUBS 0.01948f
C274 B.n184 VSUBS 0.01948f
C275 B.n185 VSUBS 0.018196f
C276 B.n186 VSUBS 0.007956f
C277 B.n187 VSUBS 0.007956f
C278 B.n188 VSUBS 0.007956f
C279 B.n189 VSUBS 0.007956f
C280 B.n190 VSUBS 0.007956f
C281 B.n191 VSUBS 0.007956f
C282 B.n192 VSUBS 0.007956f
C283 B.n193 VSUBS 0.007956f
C284 B.n194 VSUBS 0.007956f
C285 B.n195 VSUBS 0.007956f
C286 B.n196 VSUBS 0.007956f
C287 B.n197 VSUBS 0.007956f
C288 B.n198 VSUBS 0.007956f
C289 B.n199 VSUBS 0.007956f
C290 B.n200 VSUBS 0.007956f
C291 B.n201 VSUBS 0.007956f
C292 B.n202 VSUBS 0.007956f
C293 B.n203 VSUBS 0.007956f
C294 B.n204 VSUBS 0.007956f
C295 B.n205 VSUBS 0.007956f
C296 B.n206 VSUBS 0.007956f
C297 B.n207 VSUBS 0.007956f
C298 B.n208 VSUBS 0.007956f
C299 B.n209 VSUBS 0.007956f
C300 B.n210 VSUBS 0.007956f
C301 B.n211 VSUBS 0.007956f
C302 B.n212 VSUBS 0.007956f
C303 B.n213 VSUBS 0.007956f
C304 B.n214 VSUBS 0.007956f
C305 B.n215 VSUBS 0.007956f
C306 B.n216 VSUBS 0.007956f
C307 B.n217 VSUBS 0.007956f
C308 B.n218 VSUBS 0.007956f
C309 B.n219 VSUBS 0.007956f
C310 B.n220 VSUBS 0.007956f
C311 B.n221 VSUBS 0.007956f
C312 B.n222 VSUBS 0.007956f
C313 B.n223 VSUBS 0.007956f
C314 B.n224 VSUBS 0.007956f
C315 B.n225 VSUBS 0.007956f
C316 B.n226 VSUBS 0.007956f
C317 B.n227 VSUBS 0.007956f
C318 B.n228 VSUBS 0.007956f
C319 B.n229 VSUBS 0.007956f
C320 B.n230 VSUBS 0.007956f
C321 B.n231 VSUBS 0.007956f
C322 B.n232 VSUBS 0.007956f
C323 B.n233 VSUBS 0.007956f
C324 B.n234 VSUBS 0.007956f
C325 B.n235 VSUBS 0.007956f
C326 B.n236 VSUBS 0.007956f
C327 B.n237 VSUBS 0.007956f
C328 B.n238 VSUBS 0.007956f
C329 B.n239 VSUBS 0.007956f
C330 B.n240 VSUBS 0.007956f
C331 B.n241 VSUBS 0.007956f
C332 B.n242 VSUBS 0.007956f
C333 B.n243 VSUBS 0.007956f
C334 B.n244 VSUBS 0.007956f
C335 B.n245 VSUBS 0.007956f
C336 B.n246 VSUBS 0.007956f
C337 B.n247 VSUBS 0.007956f
C338 B.n248 VSUBS 0.019119f
C339 B.n249 VSUBS 0.018556f
C340 B.n250 VSUBS 0.01948f
C341 B.n251 VSUBS 0.007956f
C342 B.n252 VSUBS 0.007956f
C343 B.n253 VSUBS 0.007956f
C344 B.n254 VSUBS 0.007956f
C345 B.n255 VSUBS 0.007956f
C346 B.n256 VSUBS 0.007956f
C347 B.n257 VSUBS 0.007956f
C348 B.n258 VSUBS 0.007956f
C349 B.n259 VSUBS 0.007956f
C350 B.n260 VSUBS 0.007956f
C351 B.n261 VSUBS 0.007956f
C352 B.n262 VSUBS 0.007956f
C353 B.n263 VSUBS 0.007956f
C354 B.n264 VSUBS 0.007956f
C355 B.n265 VSUBS 0.007956f
C356 B.n266 VSUBS 0.007956f
C357 B.n267 VSUBS 0.007956f
C358 B.n268 VSUBS 0.007956f
C359 B.n269 VSUBS 0.007956f
C360 B.n270 VSUBS 0.007956f
C361 B.n271 VSUBS 0.007488f
C362 B.n272 VSUBS 0.018434f
C363 B.n273 VSUBS 0.004446f
C364 B.n274 VSUBS 0.007956f
C365 B.n275 VSUBS 0.007956f
C366 B.n276 VSUBS 0.007956f
C367 B.n277 VSUBS 0.007956f
C368 B.n278 VSUBS 0.007956f
C369 B.n279 VSUBS 0.007956f
C370 B.n280 VSUBS 0.007956f
C371 B.n281 VSUBS 0.007956f
C372 B.n282 VSUBS 0.007956f
C373 B.n283 VSUBS 0.007956f
C374 B.n284 VSUBS 0.007956f
C375 B.n285 VSUBS 0.007956f
C376 B.n286 VSUBS 0.004446f
C377 B.n287 VSUBS 0.007956f
C378 B.n288 VSUBS 0.007956f
C379 B.n289 VSUBS 0.007488f
C380 B.n290 VSUBS 0.007956f
C381 B.n291 VSUBS 0.007956f
C382 B.n292 VSUBS 0.007956f
C383 B.n293 VSUBS 0.007956f
C384 B.n294 VSUBS 0.007956f
C385 B.n295 VSUBS 0.007956f
C386 B.n296 VSUBS 0.007956f
C387 B.n297 VSUBS 0.007956f
C388 B.n298 VSUBS 0.007956f
C389 B.n299 VSUBS 0.007956f
C390 B.n300 VSUBS 0.007956f
C391 B.n301 VSUBS 0.007956f
C392 B.n302 VSUBS 0.007956f
C393 B.n303 VSUBS 0.007956f
C394 B.n304 VSUBS 0.007956f
C395 B.n305 VSUBS 0.007956f
C396 B.n306 VSUBS 0.007956f
C397 B.n307 VSUBS 0.007956f
C398 B.n308 VSUBS 0.007956f
C399 B.n309 VSUBS 0.01948f
C400 B.n310 VSUBS 0.01948f
C401 B.n311 VSUBS 0.018196f
C402 B.n312 VSUBS 0.007956f
C403 B.n313 VSUBS 0.007956f
C404 B.n314 VSUBS 0.007956f
C405 B.n315 VSUBS 0.007956f
C406 B.n316 VSUBS 0.007956f
C407 B.n317 VSUBS 0.007956f
C408 B.n318 VSUBS 0.007956f
C409 B.n319 VSUBS 0.007956f
C410 B.n320 VSUBS 0.007956f
C411 B.n321 VSUBS 0.007956f
C412 B.n322 VSUBS 0.007956f
C413 B.n323 VSUBS 0.007956f
C414 B.n324 VSUBS 0.007956f
C415 B.n325 VSUBS 0.007956f
C416 B.n326 VSUBS 0.007956f
C417 B.n327 VSUBS 0.007956f
C418 B.n328 VSUBS 0.007956f
C419 B.n329 VSUBS 0.007956f
C420 B.n330 VSUBS 0.007956f
C421 B.n331 VSUBS 0.007956f
C422 B.n332 VSUBS 0.007956f
C423 B.n333 VSUBS 0.007956f
C424 B.n334 VSUBS 0.007956f
C425 B.n335 VSUBS 0.007956f
C426 B.n336 VSUBS 0.007956f
C427 B.n337 VSUBS 0.007956f
C428 B.n338 VSUBS 0.007956f
C429 B.n339 VSUBS 0.007956f
C430 B.n340 VSUBS 0.007956f
C431 B.n341 VSUBS 0.007956f
C432 B.n342 VSUBS 0.007956f
C433 B.n343 VSUBS 0.018016f
.ends

