* NGSPICE file created from diff_pair_sample_0847.ext - technology: sky130A

.subckt diff_pair_sample_0847 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X1 VDD2.t8 VN.t1 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=5.6706 pd=29.86 as=2.3991 ps=14.87 w=14.54 l=0.91
X2 VDD1.t9 VP.t0 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=5.6706 ps=29.86 w=14.54 l=0.91
X3 VDD1.t8 VP.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X4 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=5.6706 pd=29.86 as=0 ps=0 w=14.54 l=0.91
X5 VTAIL.t16 VN.t2 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X6 VTAIL.t5 VP.t2 VDD1.t7 B.t5 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X7 VDD1.t6 VP.t3 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=5.6706 ps=29.86 w=14.54 l=0.91
X8 VDD2.t6 VN.t3 VTAIL.t12 B.t7 sky130_fd_pr__nfet_01v8 ad=5.6706 pd=29.86 as=2.3991 ps=14.87 w=14.54 l=0.91
X9 VTAIL.t10 VN.t4 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X10 VTAIL.t4 VP.t4 VDD1.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X11 VTAIL.t14 VN.t5 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X12 VTAIL.t2 VP.t5 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X13 VTAIL.t13 VN.t6 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X14 VDD2.t2 VN.t7 VTAIL.t19 B.t3 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X15 VTAIL.t0 VP.t6 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X16 VDD1.t2 VP.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=2.3991 ps=14.87 w=14.54 l=0.91
X17 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=5.6706 pd=29.86 as=0 ps=0 w=14.54 l=0.91
X18 VDD2.t1 VN.t8 VTAIL.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=5.6706 ps=29.86 w=14.54 l=0.91
X19 VDD1.t1 VP.t8 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=5.6706 pd=29.86 as=2.3991 ps=14.87 w=14.54 l=0.91
X20 VDD1.t0 VP.t9 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.6706 pd=29.86 as=2.3991 ps=14.87 w=14.54 l=0.91
X21 VDD2.t0 VN.t9 VTAIL.t18 B.t8 sky130_fd_pr__nfet_01v8 ad=2.3991 pd=14.87 as=5.6706 ps=29.86 w=14.54 l=0.91
X22 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=5.6706 pd=29.86 as=0 ps=0 w=14.54 l=0.91
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.6706 pd=29.86 as=0 ps=0 w=14.54 l=0.91
R0 VN.n4 VN.t1 445.101
R1 VN.n23 VN.t8 445.101
R2 VN.n17 VN.t9 428.238
R3 VN.n36 VN.t3 428.238
R4 VN.n10 VN.t0 385.07
R5 VN.n5 VN.t5 385.07
R6 VN.n1 VN.t4 385.07
R7 VN.n29 VN.t7 385.07
R8 VN.n24 VN.t6 385.07
R9 VN.n20 VN.t2 385.07
R10 VN.n18 VN.n17 161.3
R11 VN.n37 VN.n36 161.3
R12 VN.n35 VN.n19 161.3
R13 VN.n34 VN.n33 161.3
R14 VN.n32 VN.n31 161.3
R15 VN.n30 VN.n21 161.3
R16 VN.n29 VN.n28 161.3
R17 VN.n27 VN.n22 161.3
R18 VN.n26 VN.n25 161.3
R19 VN.n16 VN.n0 161.3
R20 VN.n15 VN.n14 161.3
R21 VN.n13 VN.n12 161.3
R22 VN.n11 VN.n2 161.3
R23 VN.n10 VN.n9 161.3
R24 VN.n8 VN.n3 161.3
R25 VN.n7 VN.n6 161.3
R26 VN.n16 VN.n15 54.1398
R27 VN.n35 VN.n34 54.1398
R28 VN.n6 VN.n3 52.2023
R29 VN.n12 VN.n11 52.2023
R30 VN.n25 VN.n22 52.2023
R31 VN.n31 VN.n30 52.2023
R32 VN VN.n37 46.2221
R33 VN.n26 VN.n23 43.5964
R34 VN.n7 VN.n4 43.5964
R35 VN.n5 VN.n4 43.1485
R36 VN.n24 VN.n23 43.1485
R37 VN.n10 VN.n3 28.9518
R38 VN.n11 VN.n10 28.9518
R39 VN.n29 VN.n22 28.9518
R40 VN.n30 VN.n29 28.9518
R41 VN.n15 VN.n1 12.7883
R42 VN.n34 VN.n20 12.7883
R43 VN.n6 VN.n5 11.8046
R44 VN.n12 VN.n1 11.8046
R45 VN.n25 VN.n24 11.8046
R46 VN.n31 VN.n20 11.8046
R47 VN.n17 VN.n16 3.65202
R48 VN.n36 VN.n35 3.65202
R49 VN.n37 VN.n19 0.189894
R50 VN.n33 VN.n19 0.189894
R51 VN.n33 VN.n32 0.189894
R52 VN.n32 VN.n21 0.189894
R53 VN.n28 VN.n21 0.189894
R54 VN.n28 VN.n27 0.189894
R55 VN.n27 VN.n26 0.189894
R56 VN.n8 VN.n7 0.189894
R57 VN.n9 VN.n8 0.189894
R58 VN.n9 VN.n2 0.189894
R59 VN.n13 VN.n2 0.189894
R60 VN.n14 VN.n13 0.189894
R61 VN.n14 VN.n0 0.189894
R62 VN.n18 VN.n0 0.189894
R63 VN VN.n18 0.0516364
R64 VTAIL.n11 VTAIL.t17 44.1161
R65 VTAIL.n16 VTAIL.t8 44.116
R66 VTAIL.n17 VTAIL.t18 44.1158
R67 VTAIL.n2 VTAIL.t9 44.1158
R68 VTAIL.n15 VTAIL.n14 42.7543
R69 VTAIL.n13 VTAIL.n12 42.7543
R70 VTAIL.n10 VTAIL.n9 42.7543
R71 VTAIL.n8 VTAIL.n7 42.7543
R72 VTAIL.n19 VTAIL.n18 42.7543
R73 VTAIL.n1 VTAIL.n0 42.7543
R74 VTAIL.n4 VTAIL.n3 42.7543
R75 VTAIL.n6 VTAIL.n5 42.7543
R76 VTAIL.n8 VTAIL.n6 27.0393
R77 VTAIL.n17 VTAIL.n16 25.9703
R78 VTAIL.n18 VTAIL.t15 1.36226
R79 VTAIL.n18 VTAIL.t10 1.36226
R80 VTAIL.n0 VTAIL.t11 1.36226
R81 VTAIL.n0 VTAIL.t14 1.36226
R82 VTAIL.n3 VTAIL.t3 1.36226
R83 VTAIL.n3 VTAIL.t2 1.36226
R84 VTAIL.n5 VTAIL.t7 1.36226
R85 VTAIL.n5 VTAIL.t4 1.36226
R86 VTAIL.n14 VTAIL.t6 1.36226
R87 VTAIL.n14 VTAIL.t5 1.36226
R88 VTAIL.n12 VTAIL.t1 1.36226
R89 VTAIL.n12 VTAIL.t0 1.36226
R90 VTAIL.n9 VTAIL.t19 1.36226
R91 VTAIL.n9 VTAIL.t13 1.36226
R92 VTAIL.n7 VTAIL.t12 1.36226
R93 VTAIL.n7 VTAIL.t16 1.36226
R94 VTAIL.n10 VTAIL.n8 1.06947
R95 VTAIL.n11 VTAIL.n10 1.06947
R96 VTAIL.n15 VTAIL.n13 1.06947
R97 VTAIL.n16 VTAIL.n15 1.06947
R98 VTAIL.n6 VTAIL.n4 1.06947
R99 VTAIL.n4 VTAIL.n2 1.06947
R100 VTAIL.n19 VTAIL.n17 1.06947
R101 VTAIL.n13 VTAIL.n11 1.00481
R102 VTAIL.n2 VTAIL.n1 1.00481
R103 VTAIL VTAIL.n1 0.860414
R104 VTAIL VTAIL.n19 0.209552
R105 VDD2.n1 VDD2.t8 61.8636
R106 VDD2.n4 VDD2.t6 60.7948
R107 VDD2.n3 VDD2.n2 60.1794
R108 VDD2 VDD2.n7 60.1766
R109 VDD2.n6 VDD2.n5 59.4331
R110 VDD2.n1 VDD2.n0 59.433
R111 VDD2.n4 VDD2.n3 41.3274
R112 VDD2.n7 VDD2.t3 1.36226
R113 VDD2.n7 VDD2.t1 1.36226
R114 VDD2.n5 VDD2.t7 1.36226
R115 VDD2.n5 VDD2.t2 1.36226
R116 VDD2.n2 VDD2.t5 1.36226
R117 VDD2.n2 VDD2.t0 1.36226
R118 VDD2.n0 VDD2.t4 1.36226
R119 VDD2.n0 VDD2.t9 1.36226
R120 VDD2.n6 VDD2.n4 1.06947
R121 VDD2 VDD2.n6 0.325931
R122 VDD2.n3 VDD2.n1 0.212395
R123 B.n206 B.t21 587.346
R124 B.n198 B.t14 587.346
R125 B.n83 B.t18 587.346
R126 B.n91 B.t10 587.346
R127 B.n579 B.n578 585
R128 B.n581 B.n116 585
R129 B.n584 B.n583 585
R130 B.n585 B.n115 585
R131 B.n587 B.n586 585
R132 B.n589 B.n114 585
R133 B.n592 B.n591 585
R134 B.n593 B.n113 585
R135 B.n595 B.n594 585
R136 B.n597 B.n112 585
R137 B.n600 B.n599 585
R138 B.n601 B.n111 585
R139 B.n603 B.n602 585
R140 B.n605 B.n110 585
R141 B.n608 B.n607 585
R142 B.n609 B.n109 585
R143 B.n611 B.n610 585
R144 B.n613 B.n108 585
R145 B.n616 B.n615 585
R146 B.n617 B.n107 585
R147 B.n619 B.n618 585
R148 B.n621 B.n106 585
R149 B.n624 B.n623 585
R150 B.n625 B.n105 585
R151 B.n627 B.n626 585
R152 B.n629 B.n104 585
R153 B.n632 B.n631 585
R154 B.n633 B.n103 585
R155 B.n635 B.n634 585
R156 B.n637 B.n102 585
R157 B.n640 B.n639 585
R158 B.n641 B.n101 585
R159 B.n643 B.n642 585
R160 B.n645 B.n100 585
R161 B.n648 B.n647 585
R162 B.n649 B.n99 585
R163 B.n651 B.n650 585
R164 B.n653 B.n98 585
R165 B.n656 B.n655 585
R166 B.n657 B.n97 585
R167 B.n659 B.n658 585
R168 B.n661 B.n96 585
R169 B.n664 B.n663 585
R170 B.n665 B.n95 585
R171 B.n667 B.n666 585
R172 B.n669 B.n94 585
R173 B.n672 B.n671 585
R174 B.n673 B.n90 585
R175 B.n675 B.n674 585
R176 B.n677 B.n89 585
R177 B.n680 B.n679 585
R178 B.n681 B.n88 585
R179 B.n683 B.n682 585
R180 B.n685 B.n87 585
R181 B.n688 B.n687 585
R182 B.n689 B.n86 585
R183 B.n691 B.n690 585
R184 B.n693 B.n85 585
R185 B.n696 B.n695 585
R186 B.n698 B.n82 585
R187 B.n700 B.n699 585
R188 B.n702 B.n81 585
R189 B.n705 B.n704 585
R190 B.n706 B.n80 585
R191 B.n708 B.n707 585
R192 B.n710 B.n79 585
R193 B.n713 B.n712 585
R194 B.n714 B.n78 585
R195 B.n716 B.n715 585
R196 B.n718 B.n77 585
R197 B.n721 B.n720 585
R198 B.n722 B.n76 585
R199 B.n724 B.n723 585
R200 B.n726 B.n75 585
R201 B.n729 B.n728 585
R202 B.n730 B.n74 585
R203 B.n732 B.n731 585
R204 B.n734 B.n73 585
R205 B.n737 B.n736 585
R206 B.n738 B.n72 585
R207 B.n740 B.n739 585
R208 B.n742 B.n71 585
R209 B.n745 B.n744 585
R210 B.n746 B.n70 585
R211 B.n748 B.n747 585
R212 B.n750 B.n69 585
R213 B.n753 B.n752 585
R214 B.n754 B.n68 585
R215 B.n756 B.n755 585
R216 B.n758 B.n67 585
R217 B.n761 B.n760 585
R218 B.n762 B.n66 585
R219 B.n764 B.n763 585
R220 B.n766 B.n65 585
R221 B.n769 B.n768 585
R222 B.n770 B.n64 585
R223 B.n772 B.n771 585
R224 B.n774 B.n63 585
R225 B.n777 B.n776 585
R226 B.n778 B.n62 585
R227 B.n780 B.n779 585
R228 B.n782 B.n61 585
R229 B.n785 B.n784 585
R230 B.n786 B.n60 585
R231 B.n788 B.n787 585
R232 B.n790 B.n59 585
R233 B.n793 B.n792 585
R234 B.n794 B.n58 585
R235 B.n577 B.n56 585
R236 B.n797 B.n56 585
R237 B.n576 B.n55 585
R238 B.n798 B.n55 585
R239 B.n575 B.n54 585
R240 B.n799 B.n54 585
R241 B.n574 B.n573 585
R242 B.n573 B.n50 585
R243 B.n572 B.n49 585
R244 B.n805 B.n49 585
R245 B.n571 B.n48 585
R246 B.n806 B.n48 585
R247 B.n570 B.n47 585
R248 B.n807 B.n47 585
R249 B.n569 B.n568 585
R250 B.n568 B.n43 585
R251 B.n567 B.n42 585
R252 B.n813 B.n42 585
R253 B.n566 B.n41 585
R254 B.n814 B.n41 585
R255 B.n565 B.n40 585
R256 B.n815 B.n40 585
R257 B.n564 B.n563 585
R258 B.n563 B.n39 585
R259 B.n562 B.n35 585
R260 B.n821 B.n35 585
R261 B.n561 B.n34 585
R262 B.n822 B.n34 585
R263 B.n560 B.n33 585
R264 B.n823 B.n33 585
R265 B.n559 B.n558 585
R266 B.n558 B.n32 585
R267 B.n557 B.n28 585
R268 B.n829 B.n28 585
R269 B.n556 B.n27 585
R270 B.n830 B.n27 585
R271 B.n555 B.n26 585
R272 B.n831 B.n26 585
R273 B.n554 B.n553 585
R274 B.n553 B.n25 585
R275 B.n552 B.n21 585
R276 B.n837 B.n21 585
R277 B.n551 B.n20 585
R278 B.n838 B.n20 585
R279 B.n550 B.n19 585
R280 B.n839 B.n19 585
R281 B.n549 B.n548 585
R282 B.n548 B.n15 585
R283 B.n547 B.n14 585
R284 B.n845 B.n14 585
R285 B.n546 B.n13 585
R286 B.n846 B.n13 585
R287 B.n545 B.n12 585
R288 B.n847 B.n12 585
R289 B.n544 B.n543 585
R290 B.n543 B.n8 585
R291 B.n542 B.n7 585
R292 B.n853 B.n7 585
R293 B.n541 B.n6 585
R294 B.n854 B.n6 585
R295 B.n540 B.n5 585
R296 B.n855 B.n5 585
R297 B.n539 B.n538 585
R298 B.n538 B.n4 585
R299 B.n537 B.n117 585
R300 B.n537 B.n536 585
R301 B.n527 B.n118 585
R302 B.n119 B.n118 585
R303 B.n529 B.n528 585
R304 B.n530 B.n529 585
R305 B.n526 B.n124 585
R306 B.n124 B.n123 585
R307 B.n525 B.n524 585
R308 B.n524 B.n523 585
R309 B.n126 B.n125 585
R310 B.n127 B.n126 585
R311 B.n516 B.n515 585
R312 B.n517 B.n516 585
R313 B.n514 B.n132 585
R314 B.n132 B.n131 585
R315 B.n513 B.n512 585
R316 B.n512 B.n511 585
R317 B.n134 B.n133 585
R318 B.n504 B.n134 585
R319 B.n503 B.n502 585
R320 B.n505 B.n503 585
R321 B.n501 B.n139 585
R322 B.n139 B.n138 585
R323 B.n500 B.n499 585
R324 B.n499 B.n498 585
R325 B.n141 B.n140 585
R326 B.n491 B.n141 585
R327 B.n490 B.n489 585
R328 B.n492 B.n490 585
R329 B.n488 B.n146 585
R330 B.n146 B.n145 585
R331 B.n487 B.n486 585
R332 B.n486 B.n485 585
R333 B.n148 B.n147 585
R334 B.n478 B.n148 585
R335 B.n477 B.n476 585
R336 B.n479 B.n477 585
R337 B.n475 B.n153 585
R338 B.n153 B.n152 585
R339 B.n474 B.n473 585
R340 B.n473 B.n472 585
R341 B.n155 B.n154 585
R342 B.n156 B.n155 585
R343 B.n465 B.n464 585
R344 B.n466 B.n465 585
R345 B.n463 B.n160 585
R346 B.n164 B.n160 585
R347 B.n462 B.n461 585
R348 B.n461 B.n460 585
R349 B.n162 B.n161 585
R350 B.n163 B.n162 585
R351 B.n453 B.n452 585
R352 B.n454 B.n453 585
R353 B.n451 B.n169 585
R354 B.n169 B.n168 585
R355 B.n450 B.n449 585
R356 B.n449 B.n448 585
R357 B.n445 B.n173 585
R358 B.n444 B.n443 585
R359 B.n441 B.n174 585
R360 B.n441 B.n172 585
R361 B.n440 B.n439 585
R362 B.n438 B.n437 585
R363 B.n436 B.n176 585
R364 B.n434 B.n433 585
R365 B.n432 B.n177 585
R366 B.n431 B.n430 585
R367 B.n428 B.n178 585
R368 B.n426 B.n425 585
R369 B.n424 B.n179 585
R370 B.n423 B.n422 585
R371 B.n420 B.n180 585
R372 B.n418 B.n417 585
R373 B.n416 B.n181 585
R374 B.n415 B.n414 585
R375 B.n412 B.n182 585
R376 B.n410 B.n409 585
R377 B.n408 B.n183 585
R378 B.n407 B.n406 585
R379 B.n404 B.n184 585
R380 B.n402 B.n401 585
R381 B.n400 B.n185 585
R382 B.n399 B.n398 585
R383 B.n396 B.n186 585
R384 B.n394 B.n393 585
R385 B.n392 B.n187 585
R386 B.n391 B.n390 585
R387 B.n388 B.n188 585
R388 B.n386 B.n385 585
R389 B.n384 B.n189 585
R390 B.n383 B.n382 585
R391 B.n380 B.n190 585
R392 B.n378 B.n377 585
R393 B.n376 B.n191 585
R394 B.n375 B.n374 585
R395 B.n372 B.n192 585
R396 B.n370 B.n369 585
R397 B.n368 B.n193 585
R398 B.n367 B.n366 585
R399 B.n364 B.n194 585
R400 B.n362 B.n361 585
R401 B.n360 B.n195 585
R402 B.n359 B.n358 585
R403 B.n356 B.n196 585
R404 B.n354 B.n353 585
R405 B.n352 B.n197 585
R406 B.n351 B.n350 585
R407 B.n348 B.n347 585
R408 B.n346 B.n345 585
R409 B.n344 B.n202 585
R410 B.n342 B.n341 585
R411 B.n340 B.n203 585
R412 B.n339 B.n338 585
R413 B.n336 B.n204 585
R414 B.n334 B.n333 585
R415 B.n332 B.n205 585
R416 B.n331 B.n330 585
R417 B.n328 B.n327 585
R418 B.n326 B.n325 585
R419 B.n324 B.n210 585
R420 B.n322 B.n321 585
R421 B.n320 B.n211 585
R422 B.n319 B.n318 585
R423 B.n316 B.n212 585
R424 B.n314 B.n313 585
R425 B.n312 B.n213 585
R426 B.n311 B.n310 585
R427 B.n308 B.n214 585
R428 B.n306 B.n305 585
R429 B.n304 B.n215 585
R430 B.n303 B.n302 585
R431 B.n300 B.n216 585
R432 B.n298 B.n297 585
R433 B.n296 B.n217 585
R434 B.n295 B.n294 585
R435 B.n292 B.n218 585
R436 B.n290 B.n289 585
R437 B.n288 B.n219 585
R438 B.n287 B.n286 585
R439 B.n284 B.n220 585
R440 B.n282 B.n281 585
R441 B.n280 B.n221 585
R442 B.n279 B.n278 585
R443 B.n276 B.n222 585
R444 B.n274 B.n273 585
R445 B.n272 B.n223 585
R446 B.n271 B.n270 585
R447 B.n268 B.n224 585
R448 B.n266 B.n265 585
R449 B.n264 B.n225 585
R450 B.n263 B.n262 585
R451 B.n260 B.n226 585
R452 B.n258 B.n257 585
R453 B.n256 B.n227 585
R454 B.n255 B.n254 585
R455 B.n252 B.n228 585
R456 B.n250 B.n249 585
R457 B.n248 B.n229 585
R458 B.n247 B.n246 585
R459 B.n244 B.n230 585
R460 B.n242 B.n241 585
R461 B.n240 B.n231 585
R462 B.n239 B.n238 585
R463 B.n236 B.n232 585
R464 B.n234 B.n233 585
R465 B.n171 B.n170 585
R466 B.n172 B.n171 585
R467 B.n447 B.n446 585
R468 B.n448 B.n447 585
R469 B.n167 B.n166 585
R470 B.n168 B.n167 585
R471 B.n456 B.n455 585
R472 B.n455 B.n454 585
R473 B.n457 B.n165 585
R474 B.n165 B.n163 585
R475 B.n459 B.n458 585
R476 B.n460 B.n459 585
R477 B.n159 B.n158 585
R478 B.n164 B.n159 585
R479 B.n468 B.n467 585
R480 B.n467 B.n466 585
R481 B.n469 B.n157 585
R482 B.n157 B.n156 585
R483 B.n471 B.n470 585
R484 B.n472 B.n471 585
R485 B.n151 B.n150 585
R486 B.n152 B.n151 585
R487 B.n481 B.n480 585
R488 B.n480 B.n479 585
R489 B.n482 B.n149 585
R490 B.n478 B.n149 585
R491 B.n484 B.n483 585
R492 B.n485 B.n484 585
R493 B.n144 B.n143 585
R494 B.n145 B.n144 585
R495 B.n494 B.n493 585
R496 B.n493 B.n492 585
R497 B.n495 B.n142 585
R498 B.n491 B.n142 585
R499 B.n497 B.n496 585
R500 B.n498 B.n497 585
R501 B.n137 B.n136 585
R502 B.n138 B.n137 585
R503 B.n507 B.n506 585
R504 B.n506 B.n505 585
R505 B.n508 B.n135 585
R506 B.n504 B.n135 585
R507 B.n510 B.n509 585
R508 B.n511 B.n510 585
R509 B.n130 B.n129 585
R510 B.n131 B.n130 585
R511 B.n519 B.n518 585
R512 B.n518 B.n517 585
R513 B.n520 B.n128 585
R514 B.n128 B.n127 585
R515 B.n522 B.n521 585
R516 B.n523 B.n522 585
R517 B.n122 B.n121 585
R518 B.n123 B.n122 585
R519 B.n532 B.n531 585
R520 B.n531 B.n530 585
R521 B.n533 B.n120 585
R522 B.n120 B.n119 585
R523 B.n535 B.n534 585
R524 B.n536 B.n535 585
R525 B.n2 B.n0 585
R526 B.n4 B.n2 585
R527 B.n3 B.n1 585
R528 B.n854 B.n3 585
R529 B.n852 B.n851 585
R530 B.n853 B.n852 585
R531 B.n850 B.n9 585
R532 B.n9 B.n8 585
R533 B.n849 B.n848 585
R534 B.n848 B.n847 585
R535 B.n11 B.n10 585
R536 B.n846 B.n11 585
R537 B.n844 B.n843 585
R538 B.n845 B.n844 585
R539 B.n842 B.n16 585
R540 B.n16 B.n15 585
R541 B.n841 B.n840 585
R542 B.n840 B.n839 585
R543 B.n18 B.n17 585
R544 B.n838 B.n18 585
R545 B.n836 B.n835 585
R546 B.n837 B.n836 585
R547 B.n834 B.n22 585
R548 B.n25 B.n22 585
R549 B.n833 B.n832 585
R550 B.n832 B.n831 585
R551 B.n24 B.n23 585
R552 B.n830 B.n24 585
R553 B.n828 B.n827 585
R554 B.n829 B.n828 585
R555 B.n826 B.n29 585
R556 B.n32 B.n29 585
R557 B.n825 B.n824 585
R558 B.n824 B.n823 585
R559 B.n31 B.n30 585
R560 B.n822 B.n31 585
R561 B.n820 B.n819 585
R562 B.n821 B.n820 585
R563 B.n818 B.n36 585
R564 B.n39 B.n36 585
R565 B.n817 B.n816 585
R566 B.n816 B.n815 585
R567 B.n38 B.n37 585
R568 B.n814 B.n38 585
R569 B.n812 B.n811 585
R570 B.n813 B.n812 585
R571 B.n810 B.n44 585
R572 B.n44 B.n43 585
R573 B.n809 B.n808 585
R574 B.n808 B.n807 585
R575 B.n46 B.n45 585
R576 B.n806 B.n46 585
R577 B.n804 B.n803 585
R578 B.n805 B.n804 585
R579 B.n802 B.n51 585
R580 B.n51 B.n50 585
R581 B.n801 B.n800 585
R582 B.n800 B.n799 585
R583 B.n53 B.n52 585
R584 B.n798 B.n53 585
R585 B.n796 B.n795 585
R586 B.n797 B.n796 585
R587 B.n857 B.n856 585
R588 B.n856 B.n855 585
R589 B.n447 B.n173 478.086
R590 B.n796 B.n58 478.086
R591 B.n449 B.n171 478.086
R592 B.n579 B.n56 478.086
R593 B.n580 B.n57 256.663
R594 B.n582 B.n57 256.663
R595 B.n588 B.n57 256.663
R596 B.n590 B.n57 256.663
R597 B.n596 B.n57 256.663
R598 B.n598 B.n57 256.663
R599 B.n604 B.n57 256.663
R600 B.n606 B.n57 256.663
R601 B.n612 B.n57 256.663
R602 B.n614 B.n57 256.663
R603 B.n620 B.n57 256.663
R604 B.n622 B.n57 256.663
R605 B.n628 B.n57 256.663
R606 B.n630 B.n57 256.663
R607 B.n636 B.n57 256.663
R608 B.n638 B.n57 256.663
R609 B.n644 B.n57 256.663
R610 B.n646 B.n57 256.663
R611 B.n652 B.n57 256.663
R612 B.n654 B.n57 256.663
R613 B.n660 B.n57 256.663
R614 B.n662 B.n57 256.663
R615 B.n668 B.n57 256.663
R616 B.n670 B.n57 256.663
R617 B.n676 B.n57 256.663
R618 B.n678 B.n57 256.663
R619 B.n684 B.n57 256.663
R620 B.n686 B.n57 256.663
R621 B.n692 B.n57 256.663
R622 B.n694 B.n57 256.663
R623 B.n701 B.n57 256.663
R624 B.n703 B.n57 256.663
R625 B.n709 B.n57 256.663
R626 B.n711 B.n57 256.663
R627 B.n717 B.n57 256.663
R628 B.n719 B.n57 256.663
R629 B.n725 B.n57 256.663
R630 B.n727 B.n57 256.663
R631 B.n733 B.n57 256.663
R632 B.n735 B.n57 256.663
R633 B.n741 B.n57 256.663
R634 B.n743 B.n57 256.663
R635 B.n749 B.n57 256.663
R636 B.n751 B.n57 256.663
R637 B.n757 B.n57 256.663
R638 B.n759 B.n57 256.663
R639 B.n765 B.n57 256.663
R640 B.n767 B.n57 256.663
R641 B.n773 B.n57 256.663
R642 B.n775 B.n57 256.663
R643 B.n781 B.n57 256.663
R644 B.n783 B.n57 256.663
R645 B.n789 B.n57 256.663
R646 B.n791 B.n57 256.663
R647 B.n442 B.n172 256.663
R648 B.n175 B.n172 256.663
R649 B.n435 B.n172 256.663
R650 B.n429 B.n172 256.663
R651 B.n427 B.n172 256.663
R652 B.n421 B.n172 256.663
R653 B.n419 B.n172 256.663
R654 B.n413 B.n172 256.663
R655 B.n411 B.n172 256.663
R656 B.n405 B.n172 256.663
R657 B.n403 B.n172 256.663
R658 B.n397 B.n172 256.663
R659 B.n395 B.n172 256.663
R660 B.n389 B.n172 256.663
R661 B.n387 B.n172 256.663
R662 B.n381 B.n172 256.663
R663 B.n379 B.n172 256.663
R664 B.n373 B.n172 256.663
R665 B.n371 B.n172 256.663
R666 B.n365 B.n172 256.663
R667 B.n363 B.n172 256.663
R668 B.n357 B.n172 256.663
R669 B.n355 B.n172 256.663
R670 B.n349 B.n172 256.663
R671 B.n201 B.n172 256.663
R672 B.n343 B.n172 256.663
R673 B.n337 B.n172 256.663
R674 B.n335 B.n172 256.663
R675 B.n329 B.n172 256.663
R676 B.n209 B.n172 256.663
R677 B.n323 B.n172 256.663
R678 B.n317 B.n172 256.663
R679 B.n315 B.n172 256.663
R680 B.n309 B.n172 256.663
R681 B.n307 B.n172 256.663
R682 B.n301 B.n172 256.663
R683 B.n299 B.n172 256.663
R684 B.n293 B.n172 256.663
R685 B.n291 B.n172 256.663
R686 B.n285 B.n172 256.663
R687 B.n283 B.n172 256.663
R688 B.n277 B.n172 256.663
R689 B.n275 B.n172 256.663
R690 B.n269 B.n172 256.663
R691 B.n267 B.n172 256.663
R692 B.n261 B.n172 256.663
R693 B.n259 B.n172 256.663
R694 B.n253 B.n172 256.663
R695 B.n251 B.n172 256.663
R696 B.n245 B.n172 256.663
R697 B.n243 B.n172 256.663
R698 B.n237 B.n172 256.663
R699 B.n235 B.n172 256.663
R700 B.n447 B.n167 163.367
R701 B.n455 B.n167 163.367
R702 B.n455 B.n165 163.367
R703 B.n459 B.n165 163.367
R704 B.n459 B.n159 163.367
R705 B.n467 B.n159 163.367
R706 B.n467 B.n157 163.367
R707 B.n471 B.n157 163.367
R708 B.n471 B.n151 163.367
R709 B.n480 B.n151 163.367
R710 B.n480 B.n149 163.367
R711 B.n484 B.n149 163.367
R712 B.n484 B.n144 163.367
R713 B.n493 B.n144 163.367
R714 B.n493 B.n142 163.367
R715 B.n497 B.n142 163.367
R716 B.n497 B.n137 163.367
R717 B.n506 B.n137 163.367
R718 B.n506 B.n135 163.367
R719 B.n510 B.n135 163.367
R720 B.n510 B.n130 163.367
R721 B.n518 B.n130 163.367
R722 B.n518 B.n128 163.367
R723 B.n522 B.n128 163.367
R724 B.n522 B.n122 163.367
R725 B.n531 B.n122 163.367
R726 B.n531 B.n120 163.367
R727 B.n535 B.n120 163.367
R728 B.n535 B.n2 163.367
R729 B.n856 B.n2 163.367
R730 B.n856 B.n3 163.367
R731 B.n852 B.n3 163.367
R732 B.n852 B.n9 163.367
R733 B.n848 B.n9 163.367
R734 B.n848 B.n11 163.367
R735 B.n844 B.n11 163.367
R736 B.n844 B.n16 163.367
R737 B.n840 B.n16 163.367
R738 B.n840 B.n18 163.367
R739 B.n836 B.n18 163.367
R740 B.n836 B.n22 163.367
R741 B.n832 B.n22 163.367
R742 B.n832 B.n24 163.367
R743 B.n828 B.n24 163.367
R744 B.n828 B.n29 163.367
R745 B.n824 B.n29 163.367
R746 B.n824 B.n31 163.367
R747 B.n820 B.n31 163.367
R748 B.n820 B.n36 163.367
R749 B.n816 B.n36 163.367
R750 B.n816 B.n38 163.367
R751 B.n812 B.n38 163.367
R752 B.n812 B.n44 163.367
R753 B.n808 B.n44 163.367
R754 B.n808 B.n46 163.367
R755 B.n804 B.n46 163.367
R756 B.n804 B.n51 163.367
R757 B.n800 B.n51 163.367
R758 B.n800 B.n53 163.367
R759 B.n796 B.n53 163.367
R760 B.n443 B.n441 163.367
R761 B.n441 B.n440 163.367
R762 B.n437 B.n436 163.367
R763 B.n434 B.n177 163.367
R764 B.n430 B.n428 163.367
R765 B.n426 B.n179 163.367
R766 B.n422 B.n420 163.367
R767 B.n418 B.n181 163.367
R768 B.n414 B.n412 163.367
R769 B.n410 B.n183 163.367
R770 B.n406 B.n404 163.367
R771 B.n402 B.n185 163.367
R772 B.n398 B.n396 163.367
R773 B.n394 B.n187 163.367
R774 B.n390 B.n388 163.367
R775 B.n386 B.n189 163.367
R776 B.n382 B.n380 163.367
R777 B.n378 B.n191 163.367
R778 B.n374 B.n372 163.367
R779 B.n370 B.n193 163.367
R780 B.n366 B.n364 163.367
R781 B.n362 B.n195 163.367
R782 B.n358 B.n356 163.367
R783 B.n354 B.n197 163.367
R784 B.n350 B.n348 163.367
R785 B.n345 B.n344 163.367
R786 B.n342 B.n203 163.367
R787 B.n338 B.n336 163.367
R788 B.n334 B.n205 163.367
R789 B.n330 B.n328 163.367
R790 B.n325 B.n324 163.367
R791 B.n322 B.n211 163.367
R792 B.n318 B.n316 163.367
R793 B.n314 B.n213 163.367
R794 B.n310 B.n308 163.367
R795 B.n306 B.n215 163.367
R796 B.n302 B.n300 163.367
R797 B.n298 B.n217 163.367
R798 B.n294 B.n292 163.367
R799 B.n290 B.n219 163.367
R800 B.n286 B.n284 163.367
R801 B.n282 B.n221 163.367
R802 B.n278 B.n276 163.367
R803 B.n274 B.n223 163.367
R804 B.n270 B.n268 163.367
R805 B.n266 B.n225 163.367
R806 B.n262 B.n260 163.367
R807 B.n258 B.n227 163.367
R808 B.n254 B.n252 163.367
R809 B.n250 B.n229 163.367
R810 B.n246 B.n244 163.367
R811 B.n242 B.n231 163.367
R812 B.n238 B.n236 163.367
R813 B.n234 B.n171 163.367
R814 B.n449 B.n169 163.367
R815 B.n453 B.n169 163.367
R816 B.n453 B.n162 163.367
R817 B.n461 B.n162 163.367
R818 B.n461 B.n160 163.367
R819 B.n465 B.n160 163.367
R820 B.n465 B.n155 163.367
R821 B.n473 B.n155 163.367
R822 B.n473 B.n153 163.367
R823 B.n477 B.n153 163.367
R824 B.n477 B.n148 163.367
R825 B.n486 B.n148 163.367
R826 B.n486 B.n146 163.367
R827 B.n490 B.n146 163.367
R828 B.n490 B.n141 163.367
R829 B.n499 B.n141 163.367
R830 B.n499 B.n139 163.367
R831 B.n503 B.n139 163.367
R832 B.n503 B.n134 163.367
R833 B.n512 B.n134 163.367
R834 B.n512 B.n132 163.367
R835 B.n516 B.n132 163.367
R836 B.n516 B.n126 163.367
R837 B.n524 B.n126 163.367
R838 B.n524 B.n124 163.367
R839 B.n529 B.n124 163.367
R840 B.n529 B.n118 163.367
R841 B.n537 B.n118 163.367
R842 B.n538 B.n537 163.367
R843 B.n538 B.n5 163.367
R844 B.n6 B.n5 163.367
R845 B.n7 B.n6 163.367
R846 B.n543 B.n7 163.367
R847 B.n543 B.n12 163.367
R848 B.n13 B.n12 163.367
R849 B.n14 B.n13 163.367
R850 B.n548 B.n14 163.367
R851 B.n548 B.n19 163.367
R852 B.n20 B.n19 163.367
R853 B.n21 B.n20 163.367
R854 B.n553 B.n21 163.367
R855 B.n553 B.n26 163.367
R856 B.n27 B.n26 163.367
R857 B.n28 B.n27 163.367
R858 B.n558 B.n28 163.367
R859 B.n558 B.n33 163.367
R860 B.n34 B.n33 163.367
R861 B.n35 B.n34 163.367
R862 B.n563 B.n35 163.367
R863 B.n563 B.n40 163.367
R864 B.n41 B.n40 163.367
R865 B.n42 B.n41 163.367
R866 B.n568 B.n42 163.367
R867 B.n568 B.n47 163.367
R868 B.n48 B.n47 163.367
R869 B.n49 B.n48 163.367
R870 B.n573 B.n49 163.367
R871 B.n573 B.n54 163.367
R872 B.n55 B.n54 163.367
R873 B.n56 B.n55 163.367
R874 B.n792 B.n790 163.367
R875 B.n788 B.n60 163.367
R876 B.n784 B.n782 163.367
R877 B.n780 B.n62 163.367
R878 B.n776 B.n774 163.367
R879 B.n772 B.n64 163.367
R880 B.n768 B.n766 163.367
R881 B.n764 B.n66 163.367
R882 B.n760 B.n758 163.367
R883 B.n756 B.n68 163.367
R884 B.n752 B.n750 163.367
R885 B.n748 B.n70 163.367
R886 B.n744 B.n742 163.367
R887 B.n740 B.n72 163.367
R888 B.n736 B.n734 163.367
R889 B.n732 B.n74 163.367
R890 B.n728 B.n726 163.367
R891 B.n724 B.n76 163.367
R892 B.n720 B.n718 163.367
R893 B.n716 B.n78 163.367
R894 B.n712 B.n710 163.367
R895 B.n708 B.n80 163.367
R896 B.n704 B.n702 163.367
R897 B.n700 B.n82 163.367
R898 B.n695 B.n693 163.367
R899 B.n691 B.n86 163.367
R900 B.n687 B.n685 163.367
R901 B.n683 B.n88 163.367
R902 B.n679 B.n677 163.367
R903 B.n675 B.n90 163.367
R904 B.n671 B.n669 163.367
R905 B.n667 B.n95 163.367
R906 B.n663 B.n661 163.367
R907 B.n659 B.n97 163.367
R908 B.n655 B.n653 163.367
R909 B.n651 B.n99 163.367
R910 B.n647 B.n645 163.367
R911 B.n643 B.n101 163.367
R912 B.n639 B.n637 163.367
R913 B.n635 B.n103 163.367
R914 B.n631 B.n629 163.367
R915 B.n627 B.n105 163.367
R916 B.n623 B.n621 163.367
R917 B.n619 B.n107 163.367
R918 B.n615 B.n613 163.367
R919 B.n611 B.n109 163.367
R920 B.n607 B.n605 163.367
R921 B.n603 B.n111 163.367
R922 B.n599 B.n597 163.367
R923 B.n595 B.n113 163.367
R924 B.n591 B.n589 163.367
R925 B.n587 B.n115 163.367
R926 B.n583 B.n581 163.367
R927 B.n206 B.t23 96.5961
R928 B.n91 B.t12 96.5961
R929 B.n198 B.t17 96.5773
R930 B.n83 B.t19 96.5773
R931 B.n207 B.t22 72.5476
R932 B.n92 B.t13 72.5476
R933 B.n199 B.t16 72.5288
R934 B.n84 B.t20 72.5288
R935 B.n442 B.n173 71.676
R936 B.n440 B.n175 71.676
R937 B.n436 B.n435 71.676
R938 B.n429 B.n177 71.676
R939 B.n428 B.n427 71.676
R940 B.n421 B.n179 71.676
R941 B.n420 B.n419 71.676
R942 B.n413 B.n181 71.676
R943 B.n412 B.n411 71.676
R944 B.n405 B.n183 71.676
R945 B.n404 B.n403 71.676
R946 B.n397 B.n185 71.676
R947 B.n396 B.n395 71.676
R948 B.n389 B.n187 71.676
R949 B.n388 B.n387 71.676
R950 B.n381 B.n189 71.676
R951 B.n380 B.n379 71.676
R952 B.n373 B.n191 71.676
R953 B.n372 B.n371 71.676
R954 B.n365 B.n193 71.676
R955 B.n364 B.n363 71.676
R956 B.n357 B.n195 71.676
R957 B.n356 B.n355 71.676
R958 B.n349 B.n197 71.676
R959 B.n348 B.n201 71.676
R960 B.n344 B.n343 71.676
R961 B.n337 B.n203 71.676
R962 B.n336 B.n335 71.676
R963 B.n329 B.n205 71.676
R964 B.n328 B.n209 71.676
R965 B.n324 B.n323 71.676
R966 B.n317 B.n211 71.676
R967 B.n316 B.n315 71.676
R968 B.n309 B.n213 71.676
R969 B.n308 B.n307 71.676
R970 B.n301 B.n215 71.676
R971 B.n300 B.n299 71.676
R972 B.n293 B.n217 71.676
R973 B.n292 B.n291 71.676
R974 B.n285 B.n219 71.676
R975 B.n284 B.n283 71.676
R976 B.n277 B.n221 71.676
R977 B.n276 B.n275 71.676
R978 B.n269 B.n223 71.676
R979 B.n268 B.n267 71.676
R980 B.n261 B.n225 71.676
R981 B.n260 B.n259 71.676
R982 B.n253 B.n227 71.676
R983 B.n252 B.n251 71.676
R984 B.n245 B.n229 71.676
R985 B.n244 B.n243 71.676
R986 B.n237 B.n231 71.676
R987 B.n236 B.n235 71.676
R988 B.n791 B.n58 71.676
R989 B.n790 B.n789 71.676
R990 B.n783 B.n60 71.676
R991 B.n782 B.n781 71.676
R992 B.n775 B.n62 71.676
R993 B.n774 B.n773 71.676
R994 B.n767 B.n64 71.676
R995 B.n766 B.n765 71.676
R996 B.n759 B.n66 71.676
R997 B.n758 B.n757 71.676
R998 B.n751 B.n68 71.676
R999 B.n750 B.n749 71.676
R1000 B.n743 B.n70 71.676
R1001 B.n742 B.n741 71.676
R1002 B.n735 B.n72 71.676
R1003 B.n734 B.n733 71.676
R1004 B.n727 B.n74 71.676
R1005 B.n726 B.n725 71.676
R1006 B.n719 B.n76 71.676
R1007 B.n718 B.n717 71.676
R1008 B.n711 B.n78 71.676
R1009 B.n710 B.n709 71.676
R1010 B.n703 B.n80 71.676
R1011 B.n702 B.n701 71.676
R1012 B.n694 B.n82 71.676
R1013 B.n693 B.n692 71.676
R1014 B.n686 B.n86 71.676
R1015 B.n685 B.n684 71.676
R1016 B.n678 B.n88 71.676
R1017 B.n677 B.n676 71.676
R1018 B.n670 B.n90 71.676
R1019 B.n669 B.n668 71.676
R1020 B.n662 B.n95 71.676
R1021 B.n661 B.n660 71.676
R1022 B.n654 B.n97 71.676
R1023 B.n653 B.n652 71.676
R1024 B.n646 B.n99 71.676
R1025 B.n645 B.n644 71.676
R1026 B.n638 B.n101 71.676
R1027 B.n637 B.n636 71.676
R1028 B.n630 B.n103 71.676
R1029 B.n629 B.n628 71.676
R1030 B.n622 B.n105 71.676
R1031 B.n621 B.n620 71.676
R1032 B.n614 B.n107 71.676
R1033 B.n613 B.n612 71.676
R1034 B.n606 B.n109 71.676
R1035 B.n605 B.n604 71.676
R1036 B.n598 B.n111 71.676
R1037 B.n597 B.n596 71.676
R1038 B.n590 B.n113 71.676
R1039 B.n589 B.n588 71.676
R1040 B.n582 B.n115 71.676
R1041 B.n581 B.n580 71.676
R1042 B.n580 B.n579 71.676
R1043 B.n583 B.n582 71.676
R1044 B.n588 B.n587 71.676
R1045 B.n591 B.n590 71.676
R1046 B.n596 B.n595 71.676
R1047 B.n599 B.n598 71.676
R1048 B.n604 B.n603 71.676
R1049 B.n607 B.n606 71.676
R1050 B.n612 B.n611 71.676
R1051 B.n615 B.n614 71.676
R1052 B.n620 B.n619 71.676
R1053 B.n623 B.n622 71.676
R1054 B.n628 B.n627 71.676
R1055 B.n631 B.n630 71.676
R1056 B.n636 B.n635 71.676
R1057 B.n639 B.n638 71.676
R1058 B.n644 B.n643 71.676
R1059 B.n647 B.n646 71.676
R1060 B.n652 B.n651 71.676
R1061 B.n655 B.n654 71.676
R1062 B.n660 B.n659 71.676
R1063 B.n663 B.n662 71.676
R1064 B.n668 B.n667 71.676
R1065 B.n671 B.n670 71.676
R1066 B.n676 B.n675 71.676
R1067 B.n679 B.n678 71.676
R1068 B.n684 B.n683 71.676
R1069 B.n687 B.n686 71.676
R1070 B.n692 B.n691 71.676
R1071 B.n695 B.n694 71.676
R1072 B.n701 B.n700 71.676
R1073 B.n704 B.n703 71.676
R1074 B.n709 B.n708 71.676
R1075 B.n712 B.n711 71.676
R1076 B.n717 B.n716 71.676
R1077 B.n720 B.n719 71.676
R1078 B.n725 B.n724 71.676
R1079 B.n728 B.n727 71.676
R1080 B.n733 B.n732 71.676
R1081 B.n736 B.n735 71.676
R1082 B.n741 B.n740 71.676
R1083 B.n744 B.n743 71.676
R1084 B.n749 B.n748 71.676
R1085 B.n752 B.n751 71.676
R1086 B.n757 B.n756 71.676
R1087 B.n760 B.n759 71.676
R1088 B.n765 B.n764 71.676
R1089 B.n768 B.n767 71.676
R1090 B.n773 B.n772 71.676
R1091 B.n776 B.n775 71.676
R1092 B.n781 B.n780 71.676
R1093 B.n784 B.n783 71.676
R1094 B.n789 B.n788 71.676
R1095 B.n792 B.n791 71.676
R1096 B.n443 B.n442 71.676
R1097 B.n437 B.n175 71.676
R1098 B.n435 B.n434 71.676
R1099 B.n430 B.n429 71.676
R1100 B.n427 B.n426 71.676
R1101 B.n422 B.n421 71.676
R1102 B.n419 B.n418 71.676
R1103 B.n414 B.n413 71.676
R1104 B.n411 B.n410 71.676
R1105 B.n406 B.n405 71.676
R1106 B.n403 B.n402 71.676
R1107 B.n398 B.n397 71.676
R1108 B.n395 B.n394 71.676
R1109 B.n390 B.n389 71.676
R1110 B.n387 B.n386 71.676
R1111 B.n382 B.n381 71.676
R1112 B.n379 B.n378 71.676
R1113 B.n374 B.n373 71.676
R1114 B.n371 B.n370 71.676
R1115 B.n366 B.n365 71.676
R1116 B.n363 B.n362 71.676
R1117 B.n358 B.n357 71.676
R1118 B.n355 B.n354 71.676
R1119 B.n350 B.n349 71.676
R1120 B.n345 B.n201 71.676
R1121 B.n343 B.n342 71.676
R1122 B.n338 B.n337 71.676
R1123 B.n335 B.n334 71.676
R1124 B.n330 B.n329 71.676
R1125 B.n325 B.n209 71.676
R1126 B.n323 B.n322 71.676
R1127 B.n318 B.n317 71.676
R1128 B.n315 B.n314 71.676
R1129 B.n310 B.n309 71.676
R1130 B.n307 B.n306 71.676
R1131 B.n302 B.n301 71.676
R1132 B.n299 B.n298 71.676
R1133 B.n294 B.n293 71.676
R1134 B.n291 B.n290 71.676
R1135 B.n286 B.n285 71.676
R1136 B.n283 B.n282 71.676
R1137 B.n278 B.n277 71.676
R1138 B.n275 B.n274 71.676
R1139 B.n270 B.n269 71.676
R1140 B.n267 B.n266 71.676
R1141 B.n262 B.n261 71.676
R1142 B.n259 B.n258 71.676
R1143 B.n254 B.n253 71.676
R1144 B.n251 B.n250 71.676
R1145 B.n246 B.n245 71.676
R1146 B.n243 B.n242 71.676
R1147 B.n238 B.n237 71.676
R1148 B.n235 B.n234 71.676
R1149 B.n448 B.n172 68.2821
R1150 B.n797 B.n57 68.2821
R1151 B.n208 B.n207 59.5399
R1152 B.n200 B.n199 59.5399
R1153 B.n697 B.n84 59.5399
R1154 B.n93 B.n92 59.5399
R1155 B.n448 B.n168 37.7497
R1156 B.n454 B.n168 37.7497
R1157 B.n454 B.n163 37.7497
R1158 B.n460 B.n163 37.7497
R1159 B.n460 B.n164 37.7497
R1160 B.n466 B.n156 37.7497
R1161 B.n472 B.n156 37.7497
R1162 B.n472 B.n152 37.7497
R1163 B.n479 B.n152 37.7497
R1164 B.n479 B.n478 37.7497
R1165 B.n485 B.n145 37.7497
R1166 B.n492 B.n145 37.7497
R1167 B.n492 B.n491 37.7497
R1168 B.n498 B.n138 37.7497
R1169 B.n505 B.n138 37.7497
R1170 B.n505 B.n504 37.7497
R1171 B.n511 B.n131 37.7497
R1172 B.n517 B.n131 37.7497
R1173 B.n523 B.n127 37.7497
R1174 B.n523 B.n123 37.7497
R1175 B.n530 B.n123 37.7497
R1176 B.n536 B.n119 37.7497
R1177 B.n536 B.n4 37.7497
R1178 B.n855 B.n4 37.7497
R1179 B.n855 B.n854 37.7497
R1180 B.n854 B.n853 37.7497
R1181 B.n853 B.n8 37.7497
R1182 B.n847 B.n846 37.7497
R1183 B.n846 B.n845 37.7497
R1184 B.n845 B.n15 37.7497
R1185 B.n839 B.n838 37.7497
R1186 B.n838 B.n837 37.7497
R1187 B.n831 B.n25 37.7497
R1188 B.n831 B.n830 37.7497
R1189 B.n830 B.n829 37.7497
R1190 B.n823 B.n32 37.7497
R1191 B.n823 B.n822 37.7497
R1192 B.n822 B.n821 37.7497
R1193 B.n815 B.n39 37.7497
R1194 B.n815 B.n814 37.7497
R1195 B.n814 B.n813 37.7497
R1196 B.n813 B.n43 37.7497
R1197 B.n807 B.n43 37.7497
R1198 B.n806 B.n805 37.7497
R1199 B.n805 B.n50 37.7497
R1200 B.n799 B.n50 37.7497
R1201 B.n799 B.n798 37.7497
R1202 B.n798 B.n797 37.7497
R1203 B.n478 B.t7 37.1945
R1204 B.n39 B.t8 37.1945
R1205 B.n517 B.t2 34.974
R1206 B.n839 B.t0 34.974
R1207 B.n466 B.t15 32.7535
R1208 B.n807 B.t11 32.7535
R1209 B.n795 B.n794 31.0639
R1210 B.n578 B.n577 31.0639
R1211 B.n450 B.n170 31.0639
R1212 B.n446 B.n445 31.0639
R1213 B.n511 B.t3 27.2021
R1214 B.n837 B.t6 27.2021
R1215 B.n207 B.n206 24.049
R1216 B.n199 B.n198 24.049
R1217 B.n84 B.n83 24.049
R1218 B.n92 B.n91 24.049
R1219 B.n491 B.t4 23.8713
R1220 B.n32 B.t5 23.8713
R1221 B.n530 B.t9 21.6508
R1222 B.n847 B.t1 21.6508
R1223 B B.n857 18.0485
R1224 B.t9 B.n119 16.0994
R1225 B.t1 B.n8 16.0994
R1226 B.n498 B.t4 13.8789
R1227 B.n829 B.t5 13.8789
R1228 B.n794 B.n793 10.6151
R1229 B.n793 B.n59 10.6151
R1230 B.n787 B.n59 10.6151
R1231 B.n787 B.n786 10.6151
R1232 B.n786 B.n785 10.6151
R1233 B.n785 B.n61 10.6151
R1234 B.n779 B.n61 10.6151
R1235 B.n779 B.n778 10.6151
R1236 B.n778 B.n777 10.6151
R1237 B.n777 B.n63 10.6151
R1238 B.n771 B.n63 10.6151
R1239 B.n771 B.n770 10.6151
R1240 B.n770 B.n769 10.6151
R1241 B.n769 B.n65 10.6151
R1242 B.n763 B.n65 10.6151
R1243 B.n763 B.n762 10.6151
R1244 B.n762 B.n761 10.6151
R1245 B.n761 B.n67 10.6151
R1246 B.n755 B.n67 10.6151
R1247 B.n755 B.n754 10.6151
R1248 B.n754 B.n753 10.6151
R1249 B.n753 B.n69 10.6151
R1250 B.n747 B.n69 10.6151
R1251 B.n747 B.n746 10.6151
R1252 B.n746 B.n745 10.6151
R1253 B.n745 B.n71 10.6151
R1254 B.n739 B.n71 10.6151
R1255 B.n739 B.n738 10.6151
R1256 B.n738 B.n737 10.6151
R1257 B.n737 B.n73 10.6151
R1258 B.n731 B.n73 10.6151
R1259 B.n731 B.n730 10.6151
R1260 B.n730 B.n729 10.6151
R1261 B.n729 B.n75 10.6151
R1262 B.n723 B.n75 10.6151
R1263 B.n723 B.n722 10.6151
R1264 B.n722 B.n721 10.6151
R1265 B.n721 B.n77 10.6151
R1266 B.n715 B.n77 10.6151
R1267 B.n715 B.n714 10.6151
R1268 B.n714 B.n713 10.6151
R1269 B.n713 B.n79 10.6151
R1270 B.n707 B.n79 10.6151
R1271 B.n707 B.n706 10.6151
R1272 B.n706 B.n705 10.6151
R1273 B.n705 B.n81 10.6151
R1274 B.n699 B.n81 10.6151
R1275 B.n699 B.n698 10.6151
R1276 B.n696 B.n85 10.6151
R1277 B.n690 B.n85 10.6151
R1278 B.n690 B.n689 10.6151
R1279 B.n689 B.n688 10.6151
R1280 B.n688 B.n87 10.6151
R1281 B.n682 B.n87 10.6151
R1282 B.n682 B.n681 10.6151
R1283 B.n681 B.n680 10.6151
R1284 B.n680 B.n89 10.6151
R1285 B.n674 B.n673 10.6151
R1286 B.n673 B.n672 10.6151
R1287 B.n672 B.n94 10.6151
R1288 B.n666 B.n94 10.6151
R1289 B.n666 B.n665 10.6151
R1290 B.n665 B.n664 10.6151
R1291 B.n664 B.n96 10.6151
R1292 B.n658 B.n96 10.6151
R1293 B.n658 B.n657 10.6151
R1294 B.n657 B.n656 10.6151
R1295 B.n656 B.n98 10.6151
R1296 B.n650 B.n98 10.6151
R1297 B.n650 B.n649 10.6151
R1298 B.n649 B.n648 10.6151
R1299 B.n648 B.n100 10.6151
R1300 B.n642 B.n100 10.6151
R1301 B.n642 B.n641 10.6151
R1302 B.n641 B.n640 10.6151
R1303 B.n640 B.n102 10.6151
R1304 B.n634 B.n102 10.6151
R1305 B.n634 B.n633 10.6151
R1306 B.n633 B.n632 10.6151
R1307 B.n632 B.n104 10.6151
R1308 B.n626 B.n104 10.6151
R1309 B.n626 B.n625 10.6151
R1310 B.n625 B.n624 10.6151
R1311 B.n624 B.n106 10.6151
R1312 B.n618 B.n106 10.6151
R1313 B.n618 B.n617 10.6151
R1314 B.n617 B.n616 10.6151
R1315 B.n616 B.n108 10.6151
R1316 B.n610 B.n108 10.6151
R1317 B.n610 B.n609 10.6151
R1318 B.n609 B.n608 10.6151
R1319 B.n608 B.n110 10.6151
R1320 B.n602 B.n110 10.6151
R1321 B.n602 B.n601 10.6151
R1322 B.n601 B.n600 10.6151
R1323 B.n600 B.n112 10.6151
R1324 B.n594 B.n112 10.6151
R1325 B.n594 B.n593 10.6151
R1326 B.n593 B.n592 10.6151
R1327 B.n592 B.n114 10.6151
R1328 B.n586 B.n114 10.6151
R1329 B.n586 B.n585 10.6151
R1330 B.n585 B.n584 10.6151
R1331 B.n584 B.n116 10.6151
R1332 B.n578 B.n116 10.6151
R1333 B.n451 B.n450 10.6151
R1334 B.n452 B.n451 10.6151
R1335 B.n452 B.n161 10.6151
R1336 B.n462 B.n161 10.6151
R1337 B.n463 B.n462 10.6151
R1338 B.n464 B.n463 10.6151
R1339 B.n464 B.n154 10.6151
R1340 B.n474 B.n154 10.6151
R1341 B.n475 B.n474 10.6151
R1342 B.n476 B.n475 10.6151
R1343 B.n476 B.n147 10.6151
R1344 B.n487 B.n147 10.6151
R1345 B.n488 B.n487 10.6151
R1346 B.n489 B.n488 10.6151
R1347 B.n489 B.n140 10.6151
R1348 B.n500 B.n140 10.6151
R1349 B.n501 B.n500 10.6151
R1350 B.n502 B.n501 10.6151
R1351 B.n502 B.n133 10.6151
R1352 B.n513 B.n133 10.6151
R1353 B.n514 B.n513 10.6151
R1354 B.n515 B.n514 10.6151
R1355 B.n515 B.n125 10.6151
R1356 B.n525 B.n125 10.6151
R1357 B.n526 B.n525 10.6151
R1358 B.n528 B.n526 10.6151
R1359 B.n528 B.n527 10.6151
R1360 B.n527 B.n117 10.6151
R1361 B.n539 B.n117 10.6151
R1362 B.n540 B.n539 10.6151
R1363 B.n541 B.n540 10.6151
R1364 B.n542 B.n541 10.6151
R1365 B.n544 B.n542 10.6151
R1366 B.n545 B.n544 10.6151
R1367 B.n546 B.n545 10.6151
R1368 B.n547 B.n546 10.6151
R1369 B.n549 B.n547 10.6151
R1370 B.n550 B.n549 10.6151
R1371 B.n551 B.n550 10.6151
R1372 B.n552 B.n551 10.6151
R1373 B.n554 B.n552 10.6151
R1374 B.n555 B.n554 10.6151
R1375 B.n556 B.n555 10.6151
R1376 B.n557 B.n556 10.6151
R1377 B.n559 B.n557 10.6151
R1378 B.n560 B.n559 10.6151
R1379 B.n561 B.n560 10.6151
R1380 B.n562 B.n561 10.6151
R1381 B.n564 B.n562 10.6151
R1382 B.n565 B.n564 10.6151
R1383 B.n566 B.n565 10.6151
R1384 B.n567 B.n566 10.6151
R1385 B.n569 B.n567 10.6151
R1386 B.n570 B.n569 10.6151
R1387 B.n571 B.n570 10.6151
R1388 B.n572 B.n571 10.6151
R1389 B.n574 B.n572 10.6151
R1390 B.n575 B.n574 10.6151
R1391 B.n576 B.n575 10.6151
R1392 B.n577 B.n576 10.6151
R1393 B.n445 B.n444 10.6151
R1394 B.n444 B.n174 10.6151
R1395 B.n439 B.n174 10.6151
R1396 B.n439 B.n438 10.6151
R1397 B.n438 B.n176 10.6151
R1398 B.n433 B.n176 10.6151
R1399 B.n433 B.n432 10.6151
R1400 B.n432 B.n431 10.6151
R1401 B.n431 B.n178 10.6151
R1402 B.n425 B.n178 10.6151
R1403 B.n425 B.n424 10.6151
R1404 B.n424 B.n423 10.6151
R1405 B.n423 B.n180 10.6151
R1406 B.n417 B.n180 10.6151
R1407 B.n417 B.n416 10.6151
R1408 B.n416 B.n415 10.6151
R1409 B.n415 B.n182 10.6151
R1410 B.n409 B.n182 10.6151
R1411 B.n409 B.n408 10.6151
R1412 B.n408 B.n407 10.6151
R1413 B.n407 B.n184 10.6151
R1414 B.n401 B.n184 10.6151
R1415 B.n401 B.n400 10.6151
R1416 B.n400 B.n399 10.6151
R1417 B.n399 B.n186 10.6151
R1418 B.n393 B.n186 10.6151
R1419 B.n393 B.n392 10.6151
R1420 B.n392 B.n391 10.6151
R1421 B.n391 B.n188 10.6151
R1422 B.n385 B.n188 10.6151
R1423 B.n385 B.n384 10.6151
R1424 B.n384 B.n383 10.6151
R1425 B.n383 B.n190 10.6151
R1426 B.n377 B.n190 10.6151
R1427 B.n377 B.n376 10.6151
R1428 B.n376 B.n375 10.6151
R1429 B.n375 B.n192 10.6151
R1430 B.n369 B.n192 10.6151
R1431 B.n369 B.n368 10.6151
R1432 B.n368 B.n367 10.6151
R1433 B.n367 B.n194 10.6151
R1434 B.n361 B.n194 10.6151
R1435 B.n361 B.n360 10.6151
R1436 B.n360 B.n359 10.6151
R1437 B.n359 B.n196 10.6151
R1438 B.n353 B.n196 10.6151
R1439 B.n353 B.n352 10.6151
R1440 B.n352 B.n351 10.6151
R1441 B.n347 B.n346 10.6151
R1442 B.n346 B.n202 10.6151
R1443 B.n341 B.n202 10.6151
R1444 B.n341 B.n340 10.6151
R1445 B.n340 B.n339 10.6151
R1446 B.n339 B.n204 10.6151
R1447 B.n333 B.n204 10.6151
R1448 B.n333 B.n332 10.6151
R1449 B.n332 B.n331 10.6151
R1450 B.n327 B.n326 10.6151
R1451 B.n326 B.n210 10.6151
R1452 B.n321 B.n210 10.6151
R1453 B.n321 B.n320 10.6151
R1454 B.n320 B.n319 10.6151
R1455 B.n319 B.n212 10.6151
R1456 B.n313 B.n212 10.6151
R1457 B.n313 B.n312 10.6151
R1458 B.n312 B.n311 10.6151
R1459 B.n311 B.n214 10.6151
R1460 B.n305 B.n214 10.6151
R1461 B.n305 B.n304 10.6151
R1462 B.n304 B.n303 10.6151
R1463 B.n303 B.n216 10.6151
R1464 B.n297 B.n216 10.6151
R1465 B.n297 B.n296 10.6151
R1466 B.n296 B.n295 10.6151
R1467 B.n295 B.n218 10.6151
R1468 B.n289 B.n218 10.6151
R1469 B.n289 B.n288 10.6151
R1470 B.n288 B.n287 10.6151
R1471 B.n287 B.n220 10.6151
R1472 B.n281 B.n220 10.6151
R1473 B.n281 B.n280 10.6151
R1474 B.n280 B.n279 10.6151
R1475 B.n279 B.n222 10.6151
R1476 B.n273 B.n222 10.6151
R1477 B.n273 B.n272 10.6151
R1478 B.n272 B.n271 10.6151
R1479 B.n271 B.n224 10.6151
R1480 B.n265 B.n224 10.6151
R1481 B.n265 B.n264 10.6151
R1482 B.n264 B.n263 10.6151
R1483 B.n263 B.n226 10.6151
R1484 B.n257 B.n226 10.6151
R1485 B.n257 B.n256 10.6151
R1486 B.n256 B.n255 10.6151
R1487 B.n255 B.n228 10.6151
R1488 B.n249 B.n228 10.6151
R1489 B.n249 B.n248 10.6151
R1490 B.n248 B.n247 10.6151
R1491 B.n247 B.n230 10.6151
R1492 B.n241 B.n230 10.6151
R1493 B.n241 B.n240 10.6151
R1494 B.n240 B.n239 10.6151
R1495 B.n239 B.n232 10.6151
R1496 B.n233 B.n232 10.6151
R1497 B.n233 B.n170 10.6151
R1498 B.n446 B.n166 10.6151
R1499 B.n456 B.n166 10.6151
R1500 B.n457 B.n456 10.6151
R1501 B.n458 B.n457 10.6151
R1502 B.n458 B.n158 10.6151
R1503 B.n468 B.n158 10.6151
R1504 B.n469 B.n468 10.6151
R1505 B.n470 B.n469 10.6151
R1506 B.n470 B.n150 10.6151
R1507 B.n481 B.n150 10.6151
R1508 B.n482 B.n481 10.6151
R1509 B.n483 B.n482 10.6151
R1510 B.n483 B.n143 10.6151
R1511 B.n494 B.n143 10.6151
R1512 B.n495 B.n494 10.6151
R1513 B.n496 B.n495 10.6151
R1514 B.n496 B.n136 10.6151
R1515 B.n507 B.n136 10.6151
R1516 B.n508 B.n507 10.6151
R1517 B.n509 B.n508 10.6151
R1518 B.n509 B.n129 10.6151
R1519 B.n519 B.n129 10.6151
R1520 B.n520 B.n519 10.6151
R1521 B.n521 B.n520 10.6151
R1522 B.n521 B.n121 10.6151
R1523 B.n532 B.n121 10.6151
R1524 B.n533 B.n532 10.6151
R1525 B.n534 B.n533 10.6151
R1526 B.n534 B.n0 10.6151
R1527 B.n851 B.n1 10.6151
R1528 B.n851 B.n850 10.6151
R1529 B.n850 B.n849 10.6151
R1530 B.n849 B.n10 10.6151
R1531 B.n843 B.n10 10.6151
R1532 B.n843 B.n842 10.6151
R1533 B.n842 B.n841 10.6151
R1534 B.n841 B.n17 10.6151
R1535 B.n835 B.n17 10.6151
R1536 B.n835 B.n834 10.6151
R1537 B.n834 B.n833 10.6151
R1538 B.n833 B.n23 10.6151
R1539 B.n827 B.n23 10.6151
R1540 B.n827 B.n826 10.6151
R1541 B.n826 B.n825 10.6151
R1542 B.n825 B.n30 10.6151
R1543 B.n819 B.n30 10.6151
R1544 B.n819 B.n818 10.6151
R1545 B.n818 B.n817 10.6151
R1546 B.n817 B.n37 10.6151
R1547 B.n811 B.n37 10.6151
R1548 B.n811 B.n810 10.6151
R1549 B.n810 B.n809 10.6151
R1550 B.n809 B.n45 10.6151
R1551 B.n803 B.n45 10.6151
R1552 B.n803 B.n802 10.6151
R1553 B.n802 B.n801 10.6151
R1554 B.n801 B.n52 10.6151
R1555 B.n795 B.n52 10.6151
R1556 B.n504 B.t3 10.5481
R1557 B.n25 B.t6 10.5481
R1558 B.n698 B.n697 9.36635
R1559 B.n674 B.n93 9.36635
R1560 B.n351 B.n200 9.36635
R1561 B.n327 B.n208 9.36635
R1562 B.n164 B.t15 4.99671
R1563 B.t11 B.n806 4.99671
R1564 B.n857 B.n0 2.81026
R1565 B.n857 B.n1 2.81026
R1566 B.t2 B.n127 2.77618
R1567 B.t0 B.n15 2.77618
R1568 B.n697 B.n696 1.24928
R1569 B.n93 B.n89 1.24928
R1570 B.n347 B.n200 1.24928
R1571 B.n331 B.n208 1.24928
R1572 B.n485 B.t7 0.555635
R1573 B.n821 B.t8 0.555635
R1574 VP.n10 VP.t9 445.101
R1575 VP.n5 VP.t8 428.238
R1576 VP.n41 VP.t0 428.238
R1577 VP.n23 VP.t3 428.238
R1578 VP.n34 VP.t1 385.07
R1579 VP.n29 VP.t4 385.07
R1580 VP.n1 VP.t5 385.07
R1581 VP.n16 VP.t7 385.07
R1582 VP.n7 VP.t2 385.07
R1583 VP.n11 VP.t6 385.07
R1584 VP.n42 VP.n41 161.3
R1585 VP.n13 VP.n12 161.3
R1586 VP.n14 VP.n9 161.3
R1587 VP.n16 VP.n15 161.3
R1588 VP.n17 VP.n8 161.3
R1589 VP.n19 VP.n18 161.3
R1590 VP.n21 VP.n20 161.3
R1591 VP.n22 VP.n6 161.3
R1592 VP.n24 VP.n23 161.3
R1593 VP.n40 VP.n0 161.3
R1594 VP.n39 VP.n38 161.3
R1595 VP.n37 VP.n36 161.3
R1596 VP.n35 VP.n2 161.3
R1597 VP.n34 VP.n33 161.3
R1598 VP.n32 VP.n3 161.3
R1599 VP.n31 VP.n30 161.3
R1600 VP.n28 VP.n4 161.3
R1601 VP.n27 VP.n26 161.3
R1602 VP.n25 VP.n5 161.3
R1603 VP.n28 VP.n27 54.1398
R1604 VP.n40 VP.n39 54.1398
R1605 VP.n22 VP.n21 54.1398
R1606 VP.n30 VP.n3 52.2023
R1607 VP.n36 VP.n35 52.2023
R1608 VP.n18 VP.n17 52.2023
R1609 VP.n12 VP.n9 52.2023
R1610 VP.n25 VP.n24 45.8414
R1611 VP.n13 VP.n10 43.5964
R1612 VP.n11 VP.n10 43.1485
R1613 VP.n34 VP.n3 28.9518
R1614 VP.n35 VP.n34 28.9518
R1615 VP.n17 VP.n16 28.9518
R1616 VP.n16 VP.n9 28.9518
R1617 VP.n29 VP.n28 12.7883
R1618 VP.n39 VP.n1 12.7883
R1619 VP.n21 VP.n7 12.7883
R1620 VP.n30 VP.n29 11.8046
R1621 VP.n36 VP.n1 11.8046
R1622 VP.n18 VP.n7 11.8046
R1623 VP.n12 VP.n11 11.8046
R1624 VP.n27 VP.n5 3.65202
R1625 VP.n41 VP.n40 3.65202
R1626 VP.n23 VP.n22 3.65202
R1627 VP.n14 VP.n13 0.189894
R1628 VP.n15 VP.n14 0.189894
R1629 VP.n15 VP.n8 0.189894
R1630 VP.n19 VP.n8 0.189894
R1631 VP.n20 VP.n19 0.189894
R1632 VP.n20 VP.n6 0.189894
R1633 VP.n24 VP.n6 0.189894
R1634 VP.n26 VP.n25 0.189894
R1635 VP.n26 VP.n4 0.189894
R1636 VP.n31 VP.n4 0.189894
R1637 VP.n32 VP.n31 0.189894
R1638 VP.n33 VP.n32 0.189894
R1639 VP.n33 VP.n2 0.189894
R1640 VP.n37 VP.n2 0.189894
R1641 VP.n38 VP.n37 0.189894
R1642 VP.n38 VP.n0 0.189894
R1643 VP.n42 VP.n0 0.189894
R1644 VP VP.n42 0.0516364
R1645 VDD1.n1 VDD1.t0 61.8638
R1646 VDD1.n3 VDD1.t1 61.8636
R1647 VDD1.n5 VDD1.n4 60.1794
R1648 VDD1.n7 VDD1.n6 59.4331
R1649 VDD1.n1 VDD1.n0 59.4331
R1650 VDD1.n3 VDD1.n2 59.433
R1651 VDD1.n7 VDD1.n5 42.4449
R1652 VDD1.n6 VDD1.t7 1.36226
R1653 VDD1.n6 VDD1.t6 1.36226
R1654 VDD1.n0 VDD1.t3 1.36226
R1655 VDD1.n0 VDD1.t2 1.36226
R1656 VDD1.n4 VDD1.t4 1.36226
R1657 VDD1.n4 VDD1.t9 1.36226
R1658 VDD1.n2 VDD1.t5 1.36226
R1659 VDD1.n2 VDD1.t8 1.36226
R1660 VDD1 VDD1.n7 0.744035
R1661 VDD1 VDD1.n1 0.325931
R1662 VDD1.n5 VDD1.n3 0.212395
C0 VP VDD1 9.34736f
C1 VDD1 VDD2 1.10499f
C2 VTAIL VDD1 14.870501f
C3 VN VDD1 0.149819f
C4 VP VDD2 0.368954f
C5 VTAIL VP 8.983251f
C6 VTAIL VDD2 14.9056f
C7 VP VN 6.373509f
C8 VTAIL VN 8.96861f
C9 VN VDD2 9.13351f
C10 VDD2 B 5.673996f
C11 VDD1 B 5.609646f
C12 VTAIL B 7.66624f
C13 VN B 10.6402f
C14 VP B 8.678586f
C15 VDD1.t0 B 3.1171f
C16 VDD1.t3 B 0.270919f
C17 VDD1.t2 B 0.270919f
C18 VDD1.n0 B 2.43714f
C19 VDD1.n1 B 0.656935f
C20 VDD1.t1 B 3.11709f
C21 VDD1.t5 B 0.270919f
C22 VDD1.t8 B 0.270919f
C23 VDD1.n2 B 2.43715f
C24 VDD1.n3 B 0.650892f
C25 VDD1.t4 B 0.270919f
C26 VDD1.t9 B 0.270919f
C27 VDD1.n4 B 2.44147f
C28 VDD1.n5 B 2.13232f
C29 VDD1.t7 B 0.270919f
C30 VDD1.t6 B 0.270919f
C31 VDD1.n6 B 2.43714f
C32 VDD1.n7 B 2.52419f
C33 VP.n0 B 0.038632f
C34 VP.t5 B 1.39964f
C35 VP.n1 B 0.51286f
C36 VP.n2 B 0.038632f
C37 VP.t1 B 1.39964f
C38 VP.n3 B 0.038927f
C39 VP.n4 B 0.038632f
C40 VP.t4 B 1.39964f
C41 VP.t8 B 1.45317f
C42 VP.n5 B 0.5542f
C43 VP.n6 B 0.038632f
C44 VP.t3 B 1.45317f
C45 VP.t2 B 1.39964f
C46 VP.n7 B 0.51286f
C47 VP.n8 B 0.038632f
C48 VP.t7 B 1.39964f
C49 VP.n9 B 0.038927f
C50 VP.t9 B 1.47458f
C51 VP.n10 B 0.560741f
C52 VP.t6 B 1.39964f
C53 VP.n11 B 0.548619f
C54 VP.n12 B 0.05063f
C55 VP.n13 B 0.162539f
C56 VP.n14 B 0.038632f
C57 VP.n15 B 0.038632f
C58 VP.n16 B 0.557867f
C59 VP.n17 B 0.038927f
C60 VP.n18 B 0.05063f
C61 VP.n19 B 0.038632f
C62 VP.n20 B 0.038632f
C63 VP.n21 B 0.050417f
C64 VP.n22 B 0.012497f
C65 VP.n23 B 0.5542f
C66 VP.n24 B 1.83748f
C67 VP.n25 B 1.86786f
C68 VP.n26 B 0.038632f
C69 VP.n27 B 0.012497f
C70 VP.n28 B 0.050417f
C71 VP.n29 B 0.51286f
C72 VP.n30 B 0.05063f
C73 VP.n31 B 0.038632f
C74 VP.n32 B 0.038632f
C75 VP.n33 B 0.038632f
C76 VP.n34 B 0.557867f
C77 VP.n35 B 0.038927f
C78 VP.n36 B 0.05063f
C79 VP.n37 B 0.038632f
C80 VP.n38 B 0.038632f
C81 VP.n39 B 0.050417f
C82 VP.n40 B 0.012497f
C83 VP.t0 B 1.45317f
C84 VP.n41 B 0.5542f
C85 VP.n42 B 0.029938f
C86 VDD2.t8 B 3.1025f
C87 VDD2.t4 B 0.26965f
C88 VDD2.t9 B 0.26965f
C89 VDD2.n0 B 2.42573f
C90 VDD2.n1 B 0.647844f
C91 VDD2.t5 B 0.26965f
C92 VDD2.t0 B 0.26965f
C93 VDD2.n2 B 2.43004f
C94 VDD2.n3 B 2.04457f
C95 VDD2.t6 B 3.09637f
C96 VDD2.n4 B 2.512f
C97 VDD2.t7 B 0.26965f
C98 VDD2.t2 B 0.26965f
C99 VDD2.n5 B 2.42573f
C100 VDD2.n6 B 0.305189f
C101 VDD2.t3 B 0.26965f
C102 VDD2.t1 B 0.26965f
C103 VDD2.n7 B 2.43001f
C104 VTAIL.t11 B 0.283108f
C105 VTAIL.t14 B 0.283108f
C106 VTAIL.n0 B 2.46682f
C107 VTAIL.n1 B 0.404213f
C108 VTAIL.t9 B 3.14768f
C109 VTAIL.n2 B 0.51206f
C110 VTAIL.t3 B 0.283108f
C111 VTAIL.t2 B 0.283108f
C112 VTAIL.n3 B 2.46682f
C113 VTAIL.n4 B 0.425944f
C114 VTAIL.t7 B 0.283108f
C115 VTAIL.t4 B 0.283108f
C116 VTAIL.n5 B 2.46682f
C117 VTAIL.n6 B 1.84068f
C118 VTAIL.t12 B 0.283108f
C119 VTAIL.t16 B 0.283108f
C120 VTAIL.n7 B 2.46682f
C121 VTAIL.n8 B 1.84068f
C122 VTAIL.t19 B 0.283108f
C123 VTAIL.t13 B 0.283108f
C124 VTAIL.n9 B 2.46682f
C125 VTAIL.n10 B 0.425945f
C126 VTAIL.t17 B 3.14769f
C127 VTAIL.n11 B 0.512052f
C128 VTAIL.t1 B 0.283108f
C129 VTAIL.t0 B 0.283108f
C130 VTAIL.n12 B 2.46682f
C131 VTAIL.n13 B 0.420812f
C132 VTAIL.t6 B 0.283108f
C133 VTAIL.t5 B 0.283108f
C134 VTAIL.n14 B 2.46682f
C135 VTAIL.n15 B 0.425945f
C136 VTAIL.t8 B 3.14769f
C137 VTAIL.n16 B 1.84705f
C138 VTAIL.t18 B 3.14768f
C139 VTAIL.n17 B 1.84706f
C140 VTAIL.t15 B 0.283108f
C141 VTAIL.t10 B 0.283108f
C142 VTAIL.n18 B 2.46682f
C143 VTAIL.n19 B 0.357671f
C144 VN.n0 B 0.038235f
C145 VN.t4 B 1.38526f
C146 VN.n1 B 0.507592f
C147 VN.n2 B 0.038235f
C148 VN.t0 B 1.38526f
C149 VN.n3 B 0.038527f
C150 VN.t1 B 1.45944f
C151 VN.n4 B 0.554981f
C152 VN.t5 B 1.38526f
C153 VN.n5 B 0.542983f
C154 VN.n6 B 0.050109f
C155 VN.n7 B 0.160869f
C156 VN.n8 B 0.038235f
C157 VN.n9 B 0.038235f
C158 VN.n10 B 0.552136f
C159 VN.n11 B 0.038527f
C160 VN.n12 B 0.050109f
C161 VN.n13 B 0.038235f
C162 VN.n14 B 0.038235f
C163 VN.n15 B 0.049899f
C164 VN.n16 B 0.012368f
C165 VN.t9 B 1.43824f
C166 VN.n17 B 0.548506f
C167 VN.n18 B 0.02963f
C168 VN.n19 B 0.038235f
C169 VN.t2 B 1.38526f
C170 VN.n20 B 0.507592f
C171 VN.n21 B 0.038235f
C172 VN.t7 B 1.38526f
C173 VN.n22 B 0.038527f
C174 VN.t8 B 1.45944f
C175 VN.n23 B 0.554981f
C176 VN.t6 B 1.38526f
C177 VN.n24 B 0.542983f
C178 VN.n25 B 0.050109f
C179 VN.n26 B 0.160869f
C180 VN.n27 B 0.038235f
C181 VN.n28 B 0.038235f
C182 VN.n29 B 0.552136f
C183 VN.n30 B 0.038527f
C184 VN.n31 B 0.050109f
C185 VN.n32 B 0.038235f
C186 VN.n33 B 0.038235f
C187 VN.n34 B 0.049899f
C188 VN.n35 B 0.012368f
C189 VN.t3 B 1.43824f
C190 VN.n36 B 0.548506f
C191 VN.n37 B 1.84358f
.ends

