* NGSPICE file created from diff_pair_sample_0168.ext - technology: sky130A

.subckt diff_pair_sample_0168 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t9 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=0.5775 pd=3.83 as=1.365 ps=7.78 w=3.5 l=1.06
X1 VTAIL.t4 VP.t0 VDD1.t5 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=0.5775 pd=3.83 as=0.5775 ps=3.83 w=3.5 l=1.06
X2 B.t11 B.t9 B.t10 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=1.365 pd=7.78 as=0 ps=0 w=3.5 l=1.06
X3 VDD2.t4 VN.t1 VTAIL.t7 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=1.365 pd=7.78 as=0.5775 ps=3.83 w=3.5 l=1.06
X4 VDD1.t4 VP.t1 VTAIL.t1 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=0.5775 pd=3.83 as=1.365 ps=7.78 w=3.5 l=1.06
X5 VDD1.t3 VP.t2 VTAIL.t3 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=1.365 pd=7.78 as=0.5775 ps=3.83 w=3.5 l=1.06
X6 VDD2.t3 VN.t2 VTAIL.t6 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=0.5775 pd=3.83 as=1.365 ps=7.78 w=3.5 l=1.06
X7 B.t8 B.t6 B.t7 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=1.365 pd=7.78 as=0 ps=0 w=3.5 l=1.06
X8 VTAIL.t2 VP.t3 VDD1.t2 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=0.5775 pd=3.83 as=0.5775 ps=3.83 w=3.5 l=1.06
X9 VTAIL.t8 VN.t3 VDD2.t2 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=0.5775 pd=3.83 as=0.5775 ps=3.83 w=3.5 l=1.06
X10 VDD2.t1 VN.t4 VTAIL.t11 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=1.365 pd=7.78 as=0.5775 ps=3.83 w=3.5 l=1.06
X11 B.t5 B.t3 B.t4 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=1.365 pd=7.78 as=0 ps=0 w=3.5 l=1.06
X12 VDD1.t1 VP.t4 VTAIL.t5 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=1.365 pd=7.78 as=0.5775 ps=3.83 w=3.5 l=1.06
X13 VDD1.t0 VP.t5 VTAIL.t0 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=0.5775 pd=3.83 as=1.365 ps=7.78 w=3.5 l=1.06
X14 VTAIL.t10 VN.t5 VDD2.t0 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=0.5775 pd=3.83 as=0.5775 ps=3.83 w=3.5 l=1.06
X15 B.t2 B.t0 B.t1 w_n2082_n1668# sky130_fd_pr__pfet_01v8 ad=1.365 pd=7.78 as=0 ps=0 w=3.5 l=1.06
R0 VN.n9 VN.n6 161.3
R1 VN.n3 VN.n0 161.3
R2 VN.n1 VN.t1 139.452
R3 VN.n7 VN.t2 139.452
R4 VN.n4 VN.t0 116.635
R5 VN.n10 VN.t4 116.635
R6 VN.n11 VN.n10 80.6037
R7 VN.n5 VN.n4 80.6037
R8 VN.n2 VN.t5 79.576
R9 VN.n8 VN.t3 79.576
R10 VN.n4 VN.n3 49.676
R11 VN.n10 VN.n9 49.676
R12 VN VN.n11 36.6316
R13 VN.n2 VN.n1 32.5096
R14 VN.n8 VN.n7 32.5096
R15 VN.n7 VN.n6 28.2313
R16 VN.n1 VN.n0 28.2313
R17 VN.n3 VN.n2 24.5923
R18 VN.n9 VN.n8 24.5923
R19 VN.n11 VN.n6 0.285035
R20 VN.n5 VN.n0 0.285035
R21 VN VN.n5 0.146778
R22 VTAIL.n7 VTAIL.t6 112.904
R23 VTAIL.n11 VTAIL.t9 112.904
R24 VTAIL.n2 VTAIL.t0 112.904
R25 VTAIL.n10 VTAIL.t1 112.904
R26 VTAIL.n9 VTAIL.n8 103.618
R27 VTAIL.n6 VTAIL.n5 103.618
R28 VTAIL.n1 VTAIL.n0 103.618
R29 VTAIL.n4 VTAIL.n3 103.618
R30 VTAIL.n6 VTAIL.n4 17.7807
R31 VTAIL.n11 VTAIL.n10 16.5824
R32 VTAIL.n0 VTAIL.t7 9.28764
R33 VTAIL.n0 VTAIL.t10 9.28764
R34 VTAIL.n3 VTAIL.t3 9.28764
R35 VTAIL.n3 VTAIL.t2 9.28764
R36 VTAIL.n8 VTAIL.t5 9.28764
R37 VTAIL.n8 VTAIL.t4 9.28764
R38 VTAIL.n5 VTAIL.t11 9.28764
R39 VTAIL.n5 VTAIL.t8 9.28764
R40 VTAIL.n7 VTAIL.n6 1.19878
R41 VTAIL.n10 VTAIL.n9 1.19878
R42 VTAIL.n4 VTAIL.n2 1.19878
R43 VTAIL.n9 VTAIL.n7 1.06947
R44 VTAIL.n2 VTAIL.n1 1.06947
R45 VTAIL VTAIL.n11 0.841017
R46 VTAIL VTAIL.n1 0.358259
R47 VDD2.n1 VDD2.t4 130.427
R48 VDD2.n2 VDD2.t1 129.583
R49 VDD2.n1 VDD2.n0 120.54
R50 VDD2 VDD2.n3 120.537
R51 VDD2.n2 VDD2.n1 30.6269
R52 VDD2.n3 VDD2.t2 9.28764
R53 VDD2.n3 VDD2.t3 9.28764
R54 VDD2.n0 VDD2.t0 9.28764
R55 VDD2.n0 VDD2.t5 9.28764
R56 VDD2 VDD2.n2 0.957397
R57 VP.n5 VP.n2 161.3
R58 VP.n13 VP.n0 161.3
R59 VP.n12 VP.n11 161.3
R60 VP.n10 VP.n1 161.3
R61 VP.n3 VP.t4 139.452
R62 VP.n8 VP.t2 116.635
R63 VP.n14 VP.t5 116.635
R64 VP.n6 VP.t1 116.635
R65 VP.n7 VP.n6 80.6037
R66 VP.n15 VP.n14 80.6037
R67 VP.n9 VP.n8 80.6037
R68 VP.n12 VP.t3 79.576
R69 VP.n4 VP.t0 79.576
R70 VP.n8 VP.n1 49.676
R71 VP.n14 VP.n13 49.676
R72 VP.n6 VP.n5 49.676
R73 VP.n9 VP.n7 36.3461
R74 VP.n4 VP.n3 32.5096
R75 VP.n3 VP.n2 28.2313
R76 VP.n12 VP.n1 24.5923
R77 VP.n13 VP.n12 24.5923
R78 VP.n5 VP.n4 24.5923
R79 VP.n7 VP.n2 0.285035
R80 VP.n10 VP.n9 0.285035
R81 VP.n15 VP.n0 0.285035
R82 VP.n11 VP.n10 0.189894
R83 VP.n11 VP.n0 0.189894
R84 VP VP.n15 0.146778
R85 VDD1 VDD1.t1 130.541
R86 VDD1.n1 VDD1.t3 130.427
R87 VDD1.n1 VDD1.n0 120.54
R88 VDD1.n3 VDD1.n2 120.296
R89 VDD1.n3 VDD1.n1 31.8091
R90 VDD1.n2 VDD1.t5 9.28764
R91 VDD1.n2 VDD1.t4 9.28764
R92 VDD1.n0 VDD1.t2 9.28764
R93 VDD1.n0 VDD1.t0 9.28764
R94 VDD1 VDD1.n3 0.241879
R95 B.n203 B.n202 585
R96 B.n201 B.n66 585
R97 B.n200 B.n199 585
R98 B.n198 B.n67 585
R99 B.n197 B.n196 585
R100 B.n195 B.n68 585
R101 B.n194 B.n193 585
R102 B.n192 B.n69 585
R103 B.n191 B.n190 585
R104 B.n189 B.n70 585
R105 B.n188 B.n187 585
R106 B.n186 B.n71 585
R107 B.n185 B.n184 585
R108 B.n183 B.n72 585
R109 B.n182 B.n181 585
R110 B.n180 B.n73 585
R111 B.n179 B.n178 585
R112 B.n176 B.n74 585
R113 B.n175 B.n174 585
R114 B.n173 B.n77 585
R115 B.n172 B.n171 585
R116 B.n170 B.n78 585
R117 B.n169 B.n168 585
R118 B.n167 B.n79 585
R119 B.n166 B.n165 585
R120 B.n164 B.n80 585
R121 B.n162 B.n161 585
R122 B.n160 B.n83 585
R123 B.n159 B.n158 585
R124 B.n157 B.n84 585
R125 B.n156 B.n155 585
R126 B.n154 B.n85 585
R127 B.n153 B.n152 585
R128 B.n151 B.n86 585
R129 B.n150 B.n149 585
R130 B.n148 B.n87 585
R131 B.n147 B.n146 585
R132 B.n145 B.n88 585
R133 B.n144 B.n143 585
R134 B.n142 B.n89 585
R135 B.n141 B.n140 585
R136 B.n139 B.n90 585
R137 B.n138 B.n137 585
R138 B.n204 B.n65 585
R139 B.n206 B.n205 585
R140 B.n207 B.n64 585
R141 B.n209 B.n208 585
R142 B.n210 B.n63 585
R143 B.n212 B.n211 585
R144 B.n213 B.n62 585
R145 B.n215 B.n214 585
R146 B.n216 B.n61 585
R147 B.n218 B.n217 585
R148 B.n219 B.n60 585
R149 B.n221 B.n220 585
R150 B.n222 B.n59 585
R151 B.n224 B.n223 585
R152 B.n225 B.n58 585
R153 B.n227 B.n226 585
R154 B.n228 B.n57 585
R155 B.n230 B.n229 585
R156 B.n231 B.n56 585
R157 B.n233 B.n232 585
R158 B.n234 B.n55 585
R159 B.n236 B.n235 585
R160 B.n237 B.n54 585
R161 B.n239 B.n238 585
R162 B.n240 B.n53 585
R163 B.n242 B.n241 585
R164 B.n243 B.n52 585
R165 B.n245 B.n244 585
R166 B.n246 B.n51 585
R167 B.n248 B.n247 585
R168 B.n249 B.n50 585
R169 B.n251 B.n250 585
R170 B.n252 B.n49 585
R171 B.n254 B.n253 585
R172 B.n255 B.n48 585
R173 B.n257 B.n256 585
R174 B.n258 B.n47 585
R175 B.n260 B.n259 585
R176 B.n261 B.n46 585
R177 B.n263 B.n262 585
R178 B.n264 B.n45 585
R179 B.n266 B.n265 585
R180 B.n267 B.n44 585
R181 B.n269 B.n268 585
R182 B.n270 B.n43 585
R183 B.n272 B.n271 585
R184 B.n273 B.n42 585
R185 B.n275 B.n274 585
R186 B.n276 B.n41 585
R187 B.n278 B.n277 585
R188 B.n343 B.n14 585
R189 B.n342 B.n341 585
R190 B.n340 B.n15 585
R191 B.n339 B.n338 585
R192 B.n337 B.n16 585
R193 B.n336 B.n335 585
R194 B.n334 B.n17 585
R195 B.n333 B.n332 585
R196 B.n331 B.n18 585
R197 B.n330 B.n329 585
R198 B.n328 B.n19 585
R199 B.n327 B.n326 585
R200 B.n325 B.n20 585
R201 B.n324 B.n323 585
R202 B.n322 B.n21 585
R203 B.n321 B.n320 585
R204 B.n319 B.n22 585
R205 B.n318 B.n317 585
R206 B.n316 B.n23 585
R207 B.n315 B.n314 585
R208 B.n313 B.n27 585
R209 B.n312 B.n311 585
R210 B.n310 B.n28 585
R211 B.n309 B.n308 585
R212 B.n307 B.n29 585
R213 B.n306 B.n305 585
R214 B.n303 B.n30 585
R215 B.n302 B.n301 585
R216 B.n300 B.n33 585
R217 B.n299 B.n298 585
R218 B.n297 B.n34 585
R219 B.n296 B.n295 585
R220 B.n294 B.n35 585
R221 B.n293 B.n292 585
R222 B.n291 B.n36 585
R223 B.n290 B.n289 585
R224 B.n288 B.n37 585
R225 B.n287 B.n286 585
R226 B.n285 B.n38 585
R227 B.n284 B.n283 585
R228 B.n282 B.n39 585
R229 B.n281 B.n280 585
R230 B.n279 B.n40 585
R231 B.n345 B.n344 585
R232 B.n346 B.n13 585
R233 B.n348 B.n347 585
R234 B.n349 B.n12 585
R235 B.n351 B.n350 585
R236 B.n352 B.n11 585
R237 B.n354 B.n353 585
R238 B.n355 B.n10 585
R239 B.n357 B.n356 585
R240 B.n358 B.n9 585
R241 B.n360 B.n359 585
R242 B.n361 B.n8 585
R243 B.n363 B.n362 585
R244 B.n364 B.n7 585
R245 B.n366 B.n365 585
R246 B.n367 B.n6 585
R247 B.n369 B.n368 585
R248 B.n370 B.n5 585
R249 B.n372 B.n371 585
R250 B.n373 B.n4 585
R251 B.n375 B.n374 585
R252 B.n376 B.n3 585
R253 B.n378 B.n377 585
R254 B.n379 B.n0 585
R255 B.n2 B.n1 585
R256 B.n103 B.n102 585
R257 B.n105 B.n104 585
R258 B.n106 B.n101 585
R259 B.n108 B.n107 585
R260 B.n109 B.n100 585
R261 B.n111 B.n110 585
R262 B.n112 B.n99 585
R263 B.n114 B.n113 585
R264 B.n115 B.n98 585
R265 B.n117 B.n116 585
R266 B.n118 B.n97 585
R267 B.n120 B.n119 585
R268 B.n121 B.n96 585
R269 B.n123 B.n122 585
R270 B.n124 B.n95 585
R271 B.n126 B.n125 585
R272 B.n127 B.n94 585
R273 B.n129 B.n128 585
R274 B.n130 B.n93 585
R275 B.n132 B.n131 585
R276 B.n133 B.n92 585
R277 B.n135 B.n134 585
R278 B.n136 B.n91 585
R279 B.n137 B.n136 478.086
R280 B.n204 B.n203 478.086
R281 B.n277 B.n40 478.086
R282 B.n344 B.n343 478.086
R283 B.n81 B.t9 282.892
R284 B.n75 B.t3 282.892
R285 B.n31 B.t0 282.892
R286 B.n24 B.t6 282.892
R287 B.n381 B.n380 256.663
R288 B.n380 B.n379 235.042
R289 B.n380 B.n2 235.042
R290 B.n137 B.n90 163.367
R291 B.n141 B.n90 163.367
R292 B.n142 B.n141 163.367
R293 B.n143 B.n142 163.367
R294 B.n143 B.n88 163.367
R295 B.n147 B.n88 163.367
R296 B.n148 B.n147 163.367
R297 B.n149 B.n148 163.367
R298 B.n149 B.n86 163.367
R299 B.n153 B.n86 163.367
R300 B.n154 B.n153 163.367
R301 B.n155 B.n154 163.367
R302 B.n155 B.n84 163.367
R303 B.n159 B.n84 163.367
R304 B.n160 B.n159 163.367
R305 B.n161 B.n160 163.367
R306 B.n161 B.n80 163.367
R307 B.n166 B.n80 163.367
R308 B.n167 B.n166 163.367
R309 B.n168 B.n167 163.367
R310 B.n168 B.n78 163.367
R311 B.n172 B.n78 163.367
R312 B.n173 B.n172 163.367
R313 B.n174 B.n173 163.367
R314 B.n174 B.n74 163.367
R315 B.n179 B.n74 163.367
R316 B.n180 B.n179 163.367
R317 B.n181 B.n180 163.367
R318 B.n181 B.n72 163.367
R319 B.n185 B.n72 163.367
R320 B.n186 B.n185 163.367
R321 B.n187 B.n186 163.367
R322 B.n187 B.n70 163.367
R323 B.n191 B.n70 163.367
R324 B.n192 B.n191 163.367
R325 B.n193 B.n192 163.367
R326 B.n193 B.n68 163.367
R327 B.n197 B.n68 163.367
R328 B.n198 B.n197 163.367
R329 B.n199 B.n198 163.367
R330 B.n199 B.n66 163.367
R331 B.n203 B.n66 163.367
R332 B.n277 B.n276 163.367
R333 B.n276 B.n275 163.367
R334 B.n275 B.n42 163.367
R335 B.n271 B.n42 163.367
R336 B.n271 B.n270 163.367
R337 B.n270 B.n269 163.367
R338 B.n269 B.n44 163.367
R339 B.n265 B.n44 163.367
R340 B.n265 B.n264 163.367
R341 B.n264 B.n263 163.367
R342 B.n263 B.n46 163.367
R343 B.n259 B.n46 163.367
R344 B.n259 B.n258 163.367
R345 B.n258 B.n257 163.367
R346 B.n257 B.n48 163.367
R347 B.n253 B.n48 163.367
R348 B.n253 B.n252 163.367
R349 B.n252 B.n251 163.367
R350 B.n251 B.n50 163.367
R351 B.n247 B.n50 163.367
R352 B.n247 B.n246 163.367
R353 B.n246 B.n245 163.367
R354 B.n245 B.n52 163.367
R355 B.n241 B.n52 163.367
R356 B.n241 B.n240 163.367
R357 B.n240 B.n239 163.367
R358 B.n239 B.n54 163.367
R359 B.n235 B.n54 163.367
R360 B.n235 B.n234 163.367
R361 B.n234 B.n233 163.367
R362 B.n233 B.n56 163.367
R363 B.n229 B.n56 163.367
R364 B.n229 B.n228 163.367
R365 B.n228 B.n227 163.367
R366 B.n227 B.n58 163.367
R367 B.n223 B.n58 163.367
R368 B.n223 B.n222 163.367
R369 B.n222 B.n221 163.367
R370 B.n221 B.n60 163.367
R371 B.n217 B.n60 163.367
R372 B.n217 B.n216 163.367
R373 B.n216 B.n215 163.367
R374 B.n215 B.n62 163.367
R375 B.n211 B.n62 163.367
R376 B.n211 B.n210 163.367
R377 B.n210 B.n209 163.367
R378 B.n209 B.n64 163.367
R379 B.n205 B.n64 163.367
R380 B.n205 B.n204 163.367
R381 B.n343 B.n342 163.367
R382 B.n342 B.n15 163.367
R383 B.n338 B.n15 163.367
R384 B.n338 B.n337 163.367
R385 B.n337 B.n336 163.367
R386 B.n336 B.n17 163.367
R387 B.n332 B.n17 163.367
R388 B.n332 B.n331 163.367
R389 B.n331 B.n330 163.367
R390 B.n330 B.n19 163.367
R391 B.n326 B.n19 163.367
R392 B.n326 B.n325 163.367
R393 B.n325 B.n324 163.367
R394 B.n324 B.n21 163.367
R395 B.n320 B.n21 163.367
R396 B.n320 B.n319 163.367
R397 B.n319 B.n318 163.367
R398 B.n318 B.n23 163.367
R399 B.n314 B.n23 163.367
R400 B.n314 B.n313 163.367
R401 B.n313 B.n312 163.367
R402 B.n312 B.n28 163.367
R403 B.n308 B.n28 163.367
R404 B.n308 B.n307 163.367
R405 B.n307 B.n306 163.367
R406 B.n306 B.n30 163.367
R407 B.n301 B.n30 163.367
R408 B.n301 B.n300 163.367
R409 B.n300 B.n299 163.367
R410 B.n299 B.n34 163.367
R411 B.n295 B.n34 163.367
R412 B.n295 B.n294 163.367
R413 B.n294 B.n293 163.367
R414 B.n293 B.n36 163.367
R415 B.n289 B.n36 163.367
R416 B.n289 B.n288 163.367
R417 B.n288 B.n287 163.367
R418 B.n287 B.n38 163.367
R419 B.n283 B.n38 163.367
R420 B.n283 B.n282 163.367
R421 B.n282 B.n281 163.367
R422 B.n281 B.n40 163.367
R423 B.n344 B.n13 163.367
R424 B.n348 B.n13 163.367
R425 B.n349 B.n348 163.367
R426 B.n350 B.n349 163.367
R427 B.n350 B.n11 163.367
R428 B.n354 B.n11 163.367
R429 B.n355 B.n354 163.367
R430 B.n356 B.n355 163.367
R431 B.n356 B.n9 163.367
R432 B.n360 B.n9 163.367
R433 B.n361 B.n360 163.367
R434 B.n362 B.n361 163.367
R435 B.n362 B.n7 163.367
R436 B.n366 B.n7 163.367
R437 B.n367 B.n366 163.367
R438 B.n368 B.n367 163.367
R439 B.n368 B.n5 163.367
R440 B.n372 B.n5 163.367
R441 B.n373 B.n372 163.367
R442 B.n374 B.n373 163.367
R443 B.n374 B.n3 163.367
R444 B.n378 B.n3 163.367
R445 B.n379 B.n378 163.367
R446 B.n102 B.n2 163.367
R447 B.n105 B.n102 163.367
R448 B.n106 B.n105 163.367
R449 B.n107 B.n106 163.367
R450 B.n107 B.n100 163.367
R451 B.n111 B.n100 163.367
R452 B.n112 B.n111 163.367
R453 B.n113 B.n112 163.367
R454 B.n113 B.n98 163.367
R455 B.n117 B.n98 163.367
R456 B.n118 B.n117 163.367
R457 B.n119 B.n118 163.367
R458 B.n119 B.n96 163.367
R459 B.n123 B.n96 163.367
R460 B.n124 B.n123 163.367
R461 B.n125 B.n124 163.367
R462 B.n125 B.n94 163.367
R463 B.n129 B.n94 163.367
R464 B.n130 B.n129 163.367
R465 B.n131 B.n130 163.367
R466 B.n131 B.n92 163.367
R467 B.n135 B.n92 163.367
R468 B.n136 B.n135 163.367
R469 B.n75 B.t4 155.252
R470 B.n31 B.t2 155.252
R471 B.n81 B.t10 155.25
R472 B.n24 B.t8 155.25
R473 B.n76 B.t5 128.296
R474 B.n32 B.t1 128.296
R475 B.n82 B.t11 128.292
R476 B.n25 B.t7 128.292
R477 B.n163 B.n82 59.5399
R478 B.n177 B.n76 59.5399
R479 B.n304 B.n32 59.5399
R480 B.n26 B.n25 59.5399
R481 B.n345 B.n14 31.0639
R482 B.n279 B.n278 31.0639
R483 B.n202 B.n65 31.0639
R484 B.n138 B.n91 31.0639
R485 B.n82 B.n81 26.9581
R486 B.n76 B.n75 26.9581
R487 B.n32 B.n31 26.9581
R488 B.n25 B.n24 26.9581
R489 B B.n381 18.0485
R490 B.n346 B.n345 10.6151
R491 B.n347 B.n346 10.6151
R492 B.n347 B.n12 10.6151
R493 B.n351 B.n12 10.6151
R494 B.n352 B.n351 10.6151
R495 B.n353 B.n352 10.6151
R496 B.n353 B.n10 10.6151
R497 B.n357 B.n10 10.6151
R498 B.n358 B.n357 10.6151
R499 B.n359 B.n358 10.6151
R500 B.n359 B.n8 10.6151
R501 B.n363 B.n8 10.6151
R502 B.n364 B.n363 10.6151
R503 B.n365 B.n364 10.6151
R504 B.n365 B.n6 10.6151
R505 B.n369 B.n6 10.6151
R506 B.n370 B.n369 10.6151
R507 B.n371 B.n370 10.6151
R508 B.n371 B.n4 10.6151
R509 B.n375 B.n4 10.6151
R510 B.n376 B.n375 10.6151
R511 B.n377 B.n376 10.6151
R512 B.n377 B.n0 10.6151
R513 B.n341 B.n14 10.6151
R514 B.n341 B.n340 10.6151
R515 B.n340 B.n339 10.6151
R516 B.n339 B.n16 10.6151
R517 B.n335 B.n16 10.6151
R518 B.n335 B.n334 10.6151
R519 B.n334 B.n333 10.6151
R520 B.n333 B.n18 10.6151
R521 B.n329 B.n18 10.6151
R522 B.n329 B.n328 10.6151
R523 B.n328 B.n327 10.6151
R524 B.n327 B.n20 10.6151
R525 B.n323 B.n20 10.6151
R526 B.n323 B.n322 10.6151
R527 B.n322 B.n321 10.6151
R528 B.n321 B.n22 10.6151
R529 B.n317 B.n316 10.6151
R530 B.n316 B.n315 10.6151
R531 B.n315 B.n27 10.6151
R532 B.n311 B.n27 10.6151
R533 B.n311 B.n310 10.6151
R534 B.n310 B.n309 10.6151
R535 B.n309 B.n29 10.6151
R536 B.n305 B.n29 10.6151
R537 B.n303 B.n302 10.6151
R538 B.n302 B.n33 10.6151
R539 B.n298 B.n33 10.6151
R540 B.n298 B.n297 10.6151
R541 B.n297 B.n296 10.6151
R542 B.n296 B.n35 10.6151
R543 B.n292 B.n35 10.6151
R544 B.n292 B.n291 10.6151
R545 B.n291 B.n290 10.6151
R546 B.n290 B.n37 10.6151
R547 B.n286 B.n37 10.6151
R548 B.n286 B.n285 10.6151
R549 B.n285 B.n284 10.6151
R550 B.n284 B.n39 10.6151
R551 B.n280 B.n39 10.6151
R552 B.n280 B.n279 10.6151
R553 B.n278 B.n41 10.6151
R554 B.n274 B.n41 10.6151
R555 B.n274 B.n273 10.6151
R556 B.n273 B.n272 10.6151
R557 B.n272 B.n43 10.6151
R558 B.n268 B.n43 10.6151
R559 B.n268 B.n267 10.6151
R560 B.n267 B.n266 10.6151
R561 B.n266 B.n45 10.6151
R562 B.n262 B.n45 10.6151
R563 B.n262 B.n261 10.6151
R564 B.n261 B.n260 10.6151
R565 B.n260 B.n47 10.6151
R566 B.n256 B.n47 10.6151
R567 B.n256 B.n255 10.6151
R568 B.n255 B.n254 10.6151
R569 B.n254 B.n49 10.6151
R570 B.n250 B.n49 10.6151
R571 B.n250 B.n249 10.6151
R572 B.n249 B.n248 10.6151
R573 B.n248 B.n51 10.6151
R574 B.n244 B.n51 10.6151
R575 B.n244 B.n243 10.6151
R576 B.n243 B.n242 10.6151
R577 B.n242 B.n53 10.6151
R578 B.n238 B.n53 10.6151
R579 B.n238 B.n237 10.6151
R580 B.n237 B.n236 10.6151
R581 B.n236 B.n55 10.6151
R582 B.n232 B.n55 10.6151
R583 B.n232 B.n231 10.6151
R584 B.n231 B.n230 10.6151
R585 B.n230 B.n57 10.6151
R586 B.n226 B.n57 10.6151
R587 B.n226 B.n225 10.6151
R588 B.n225 B.n224 10.6151
R589 B.n224 B.n59 10.6151
R590 B.n220 B.n59 10.6151
R591 B.n220 B.n219 10.6151
R592 B.n219 B.n218 10.6151
R593 B.n218 B.n61 10.6151
R594 B.n214 B.n61 10.6151
R595 B.n214 B.n213 10.6151
R596 B.n213 B.n212 10.6151
R597 B.n212 B.n63 10.6151
R598 B.n208 B.n63 10.6151
R599 B.n208 B.n207 10.6151
R600 B.n207 B.n206 10.6151
R601 B.n206 B.n65 10.6151
R602 B.n103 B.n1 10.6151
R603 B.n104 B.n103 10.6151
R604 B.n104 B.n101 10.6151
R605 B.n108 B.n101 10.6151
R606 B.n109 B.n108 10.6151
R607 B.n110 B.n109 10.6151
R608 B.n110 B.n99 10.6151
R609 B.n114 B.n99 10.6151
R610 B.n115 B.n114 10.6151
R611 B.n116 B.n115 10.6151
R612 B.n116 B.n97 10.6151
R613 B.n120 B.n97 10.6151
R614 B.n121 B.n120 10.6151
R615 B.n122 B.n121 10.6151
R616 B.n122 B.n95 10.6151
R617 B.n126 B.n95 10.6151
R618 B.n127 B.n126 10.6151
R619 B.n128 B.n127 10.6151
R620 B.n128 B.n93 10.6151
R621 B.n132 B.n93 10.6151
R622 B.n133 B.n132 10.6151
R623 B.n134 B.n133 10.6151
R624 B.n134 B.n91 10.6151
R625 B.n139 B.n138 10.6151
R626 B.n140 B.n139 10.6151
R627 B.n140 B.n89 10.6151
R628 B.n144 B.n89 10.6151
R629 B.n145 B.n144 10.6151
R630 B.n146 B.n145 10.6151
R631 B.n146 B.n87 10.6151
R632 B.n150 B.n87 10.6151
R633 B.n151 B.n150 10.6151
R634 B.n152 B.n151 10.6151
R635 B.n152 B.n85 10.6151
R636 B.n156 B.n85 10.6151
R637 B.n157 B.n156 10.6151
R638 B.n158 B.n157 10.6151
R639 B.n158 B.n83 10.6151
R640 B.n162 B.n83 10.6151
R641 B.n165 B.n164 10.6151
R642 B.n165 B.n79 10.6151
R643 B.n169 B.n79 10.6151
R644 B.n170 B.n169 10.6151
R645 B.n171 B.n170 10.6151
R646 B.n171 B.n77 10.6151
R647 B.n175 B.n77 10.6151
R648 B.n176 B.n175 10.6151
R649 B.n178 B.n73 10.6151
R650 B.n182 B.n73 10.6151
R651 B.n183 B.n182 10.6151
R652 B.n184 B.n183 10.6151
R653 B.n184 B.n71 10.6151
R654 B.n188 B.n71 10.6151
R655 B.n189 B.n188 10.6151
R656 B.n190 B.n189 10.6151
R657 B.n190 B.n69 10.6151
R658 B.n194 B.n69 10.6151
R659 B.n195 B.n194 10.6151
R660 B.n196 B.n195 10.6151
R661 B.n196 B.n67 10.6151
R662 B.n200 B.n67 10.6151
R663 B.n201 B.n200 10.6151
R664 B.n202 B.n201 10.6151
R665 B.n381 B.n0 8.11757
R666 B.n381 B.n1 8.11757
R667 B.n317 B.n26 6.5566
R668 B.n305 B.n304 6.5566
R669 B.n164 B.n163 6.5566
R670 B.n177 B.n176 6.5566
R671 B.n26 B.n22 4.05904
R672 B.n304 B.n303 4.05904
R673 B.n163 B.n162 4.05904
R674 B.n178 B.n177 4.05904
C0 VDD1 VP 1.94242f
C1 w_n2082_n1668# VDD1 1.28876f
C2 VDD2 VN 1.76576f
C3 VDD1 VTAIL 4.04779f
C4 VDD1 B 1.03368f
C5 VN VP 3.85952f
C6 w_n2082_n1668# VN 3.39768f
C7 VDD2 VP 0.332398f
C8 w_n2082_n1668# VDD2 1.32384f
C9 VTAIL VN 1.9928f
C10 VN B 0.745221f
C11 w_n2082_n1668# VP 3.66099f
C12 VDD2 VTAIL 4.08939f
C13 VDD2 B 1.07122f
C14 VTAIL VP 2.00702f
C15 B VP 1.17941f
C16 w_n2082_n1668# VTAIL 1.60115f
C17 w_n2082_n1668# B 5.16735f
C18 VDD1 VN 0.15369f
C19 VTAIL B 1.29587f
C20 VDD2 VDD1 0.841103f
C21 VDD2 VSUBS 0.817243f
C22 VDD1 VSUBS 1.101222f
C23 VTAIL VSUBS 0.389892f
C24 VN VSUBS 3.45142f
C25 VP VSUBS 1.327984f
C26 B VSUBS 2.278767f
C27 w_n2082_n1668# VSUBS 43.846897f
C28 B.n0 VSUBS 0.006725f
C29 B.n1 VSUBS 0.006725f
C30 B.n2 VSUBS 0.009946f
C31 B.n3 VSUBS 0.007622f
C32 B.n4 VSUBS 0.007622f
C33 B.n5 VSUBS 0.007622f
C34 B.n6 VSUBS 0.007622f
C35 B.n7 VSUBS 0.007622f
C36 B.n8 VSUBS 0.007622f
C37 B.n9 VSUBS 0.007622f
C38 B.n10 VSUBS 0.007622f
C39 B.n11 VSUBS 0.007622f
C40 B.n12 VSUBS 0.007622f
C41 B.n13 VSUBS 0.007622f
C42 B.n14 VSUBS 0.017758f
C43 B.n15 VSUBS 0.007622f
C44 B.n16 VSUBS 0.007622f
C45 B.n17 VSUBS 0.007622f
C46 B.n18 VSUBS 0.007622f
C47 B.n19 VSUBS 0.007622f
C48 B.n20 VSUBS 0.007622f
C49 B.n21 VSUBS 0.007622f
C50 B.n22 VSUBS 0.005268f
C51 B.n23 VSUBS 0.007622f
C52 B.t7 VSUBS 0.096309f
C53 B.t8 VSUBS 0.105901f
C54 B.t6 VSUBS 0.187582f
C55 B.n24 VSUBS 0.079416f
C56 B.n25 VSUBS 0.06611f
C57 B.n26 VSUBS 0.01766f
C58 B.n27 VSUBS 0.007622f
C59 B.n28 VSUBS 0.007622f
C60 B.n29 VSUBS 0.007622f
C61 B.n30 VSUBS 0.007622f
C62 B.t1 VSUBS 0.096309f
C63 B.t2 VSUBS 0.105901f
C64 B.t0 VSUBS 0.187582f
C65 B.n31 VSUBS 0.079416f
C66 B.n32 VSUBS 0.066109f
C67 B.n33 VSUBS 0.007622f
C68 B.n34 VSUBS 0.007622f
C69 B.n35 VSUBS 0.007622f
C70 B.n36 VSUBS 0.007622f
C71 B.n37 VSUBS 0.007622f
C72 B.n38 VSUBS 0.007622f
C73 B.n39 VSUBS 0.007622f
C74 B.n40 VSUBS 0.017758f
C75 B.n41 VSUBS 0.007622f
C76 B.n42 VSUBS 0.007622f
C77 B.n43 VSUBS 0.007622f
C78 B.n44 VSUBS 0.007622f
C79 B.n45 VSUBS 0.007622f
C80 B.n46 VSUBS 0.007622f
C81 B.n47 VSUBS 0.007622f
C82 B.n48 VSUBS 0.007622f
C83 B.n49 VSUBS 0.007622f
C84 B.n50 VSUBS 0.007622f
C85 B.n51 VSUBS 0.007622f
C86 B.n52 VSUBS 0.007622f
C87 B.n53 VSUBS 0.007622f
C88 B.n54 VSUBS 0.007622f
C89 B.n55 VSUBS 0.007622f
C90 B.n56 VSUBS 0.007622f
C91 B.n57 VSUBS 0.007622f
C92 B.n58 VSUBS 0.007622f
C93 B.n59 VSUBS 0.007622f
C94 B.n60 VSUBS 0.007622f
C95 B.n61 VSUBS 0.007622f
C96 B.n62 VSUBS 0.007622f
C97 B.n63 VSUBS 0.007622f
C98 B.n64 VSUBS 0.007622f
C99 B.n65 VSUBS 0.017712f
C100 B.n66 VSUBS 0.007622f
C101 B.n67 VSUBS 0.007622f
C102 B.n68 VSUBS 0.007622f
C103 B.n69 VSUBS 0.007622f
C104 B.n70 VSUBS 0.007622f
C105 B.n71 VSUBS 0.007622f
C106 B.n72 VSUBS 0.007622f
C107 B.n73 VSUBS 0.007622f
C108 B.n74 VSUBS 0.007622f
C109 B.t5 VSUBS 0.096309f
C110 B.t4 VSUBS 0.105901f
C111 B.t3 VSUBS 0.187582f
C112 B.n75 VSUBS 0.079416f
C113 B.n76 VSUBS 0.066109f
C114 B.n77 VSUBS 0.007622f
C115 B.n78 VSUBS 0.007622f
C116 B.n79 VSUBS 0.007622f
C117 B.n80 VSUBS 0.007622f
C118 B.t11 VSUBS 0.096309f
C119 B.t10 VSUBS 0.105901f
C120 B.t9 VSUBS 0.187582f
C121 B.n81 VSUBS 0.079416f
C122 B.n82 VSUBS 0.06611f
C123 B.n83 VSUBS 0.007622f
C124 B.n84 VSUBS 0.007622f
C125 B.n85 VSUBS 0.007622f
C126 B.n86 VSUBS 0.007622f
C127 B.n87 VSUBS 0.007622f
C128 B.n88 VSUBS 0.007622f
C129 B.n89 VSUBS 0.007622f
C130 B.n90 VSUBS 0.007622f
C131 B.n91 VSUBS 0.016765f
C132 B.n92 VSUBS 0.007622f
C133 B.n93 VSUBS 0.007622f
C134 B.n94 VSUBS 0.007622f
C135 B.n95 VSUBS 0.007622f
C136 B.n96 VSUBS 0.007622f
C137 B.n97 VSUBS 0.007622f
C138 B.n98 VSUBS 0.007622f
C139 B.n99 VSUBS 0.007622f
C140 B.n100 VSUBS 0.007622f
C141 B.n101 VSUBS 0.007622f
C142 B.n102 VSUBS 0.007622f
C143 B.n103 VSUBS 0.007622f
C144 B.n104 VSUBS 0.007622f
C145 B.n105 VSUBS 0.007622f
C146 B.n106 VSUBS 0.007622f
C147 B.n107 VSUBS 0.007622f
C148 B.n108 VSUBS 0.007622f
C149 B.n109 VSUBS 0.007622f
C150 B.n110 VSUBS 0.007622f
C151 B.n111 VSUBS 0.007622f
C152 B.n112 VSUBS 0.007622f
C153 B.n113 VSUBS 0.007622f
C154 B.n114 VSUBS 0.007622f
C155 B.n115 VSUBS 0.007622f
C156 B.n116 VSUBS 0.007622f
C157 B.n117 VSUBS 0.007622f
C158 B.n118 VSUBS 0.007622f
C159 B.n119 VSUBS 0.007622f
C160 B.n120 VSUBS 0.007622f
C161 B.n121 VSUBS 0.007622f
C162 B.n122 VSUBS 0.007622f
C163 B.n123 VSUBS 0.007622f
C164 B.n124 VSUBS 0.007622f
C165 B.n125 VSUBS 0.007622f
C166 B.n126 VSUBS 0.007622f
C167 B.n127 VSUBS 0.007622f
C168 B.n128 VSUBS 0.007622f
C169 B.n129 VSUBS 0.007622f
C170 B.n130 VSUBS 0.007622f
C171 B.n131 VSUBS 0.007622f
C172 B.n132 VSUBS 0.007622f
C173 B.n133 VSUBS 0.007622f
C174 B.n134 VSUBS 0.007622f
C175 B.n135 VSUBS 0.007622f
C176 B.n136 VSUBS 0.016765f
C177 B.n137 VSUBS 0.017758f
C178 B.n138 VSUBS 0.017758f
C179 B.n139 VSUBS 0.007622f
C180 B.n140 VSUBS 0.007622f
C181 B.n141 VSUBS 0.007622f
C182 B.n142 VSUBS 0.007622f
C183 B.n143 VSUBS 0.007622f
C184 B.n144 VSUBS 0.007622f
C185 B.n145 VSUBS 0.007622f
C186 B.n146 VSUBS 0.007622f
C187 B.n147 VSUBS 0.007622f
C188 B.n148 VSUBS 0.007622f
C189 B.n149 VSUBS 0.007622f
C190 B.n150 VSUBS 0.007622f
C191 B.n151 VSUBS 0.007622f
C192 B.n152 VSUBS 0.007622f
C193 B.n153 VSUBS 0.007622f
C194 B.n154 VSUBS 0.007622f
C195 B.n155 VSUBS 0.007622f
C196 B.n156 VSUBS 0.007622f
C197 B.n157 VSUBS 0.007622f
C198 B.n158 VSUBS 0.007622f
C199 B.n159 VSUBS 0.007622f
C200 B.n160 VSUBS 0.007622f
C201 B.n161 VSUBS 0.007622f
C202 B.n162 VSUBS 0.005268f
C203 B.n163 VSUBS 0.01766f
C204 B.n164 VSUBS 0.006165f
C205 B.n165 VSUBS 0.007622f
C206 B.n166 VSUBS 0.007622f
C207 B.n167 VSUBS 0.007622f
C208 B.n168 VSUBS 0.007622f
C209 B.n169 VSUBS 0.007622f
C210 B.n170 VSUBS 0.007622f
C211 B.n171 VSUBS 0.007622f
C212 B.n172 VSUBS 0.007622f
C213 B.n173 VSUBS 0.007622f
C214 B.n174 VSUBS 0.007622f
C215 B.n175 VSUBS 0.007622f
C216 B.n176 VSUBS 0.006165f
C217 B.n177 VSUBS 0.01766f
C218 B.n178 VSUBS 0.005268f
C219 B.n179 VSUBS 0.007622f
C220 B.n180 VSUBS 0.007622f
C221 B.n181 VSUBS 0.007622f
C222 B.n182 VSUBS 0.007622f
C223 B.n183 VSUBS 0.007622f
C224 B.n184 VSUBS 0.007622f
C225 B.n185 VSUBS 0.007622f
C226 B.n186 VSUBS 0.007622f
C227 B.n187 VSUBS 0.007622f
C228 B.n188 VSUBS 0.007622f
C229 B.n189 VSUBS 0.007622f
C230 B.n190 VSUBS 0.007622f
C231 B.n191 VSUBS 0.007622f
C232 B.n192 VSUBS 0.007622f
C233 B.n193 VSUBS 0.007622f
C234 B.n194 VSUBS 0.007622f
C235 B.n195 VSUBS 0.007622f
C236 B.n196 VSUBS 0.007622f
C237 B.n197 VSUBS 0.007622f
C238 B.n198 VSUBS 0.007622f
C239 B.n199 VSUBS 0.007622f
C240 B.n200 VSUBS 0.007622f
C241 B.n201 VSUBS 0.007622f
C242 B.n202 VSUBS 0.016812f
C243 B.n203 VSUBS 0.017758f
C244 B.n204 VSUBS 0.016765f
C245 B.n205 VSUBS 0.007622f
C246 B.n206 VSUBS 0.007622f
C247 B.n207 VSUBS 0.007622f
C248 B.n208 VSUBS 0.007622f
C249 B.n209 VSUBS 0.007622f
C250 B.n210 VSUBS 0.007622f
C251 B.n211 VSUBS 0.007622f
C252 B.n212 VSUBS 0.007622f
C253 B.n213 VSUBS 0.007622f
C254 B.n214 VSUBS 0.007622f
C255 B.n215 VSUBS 0.007622f
C256 B.n216 VSUBS 0.007622f
C257 B.n217 VSUBS 0.007622f
C258 B.n218 VSUBS 0.007622f
C259 B.n219 VSUBS 0.007622f
C260 B.n220 VSUBS 0.007622f
C261 B.n221 VSUBS 0.007622f
C262 B.n222 VSUBS 0.007622f
C263 B.n223 VSUBS 0.007622f
C264 B.n224 VSUBS 0.007622f
C265 B.n225 VSUBS 0.007622f
C266 B.n226 VSUBS 0.007622f
C267 B.n227 VSUBS 0.007622f
C268 B.n228 VSUBS 0.007622f
C269 B.n229 VSUBS 0.007622f
C270 B.n230 VSUBS 0.007622f
C271 B.n231 VSUBS 0.007622f
C272 B.n232 VSUBS 0.007622f
C273 B.n233 VSUBS 0.007622f
C274 B.n234 VSUBS 0.007622f
C275 B.n235 VSUBS 0.007622f
C276 B.n236 VSUBS 0.007622f
C277 B.n237 VSUBS 0.007622f
C278 B.n238 VSUBS 0.007622f
C279 B.n239 VSUBS 0.007622f
C280 B.n240 VSUBS 0.007622f
C281 B.n241 VSUBS 0.007622f
C282 B.n242 VSUBS 0.007622f
C283 B.n243 VSUBS 0.007622f
C284 B.n244 VSUBS 0.007622f
C285 B.n245 VSUBS 0.007622f
C286 B.n246 VSUBS 0.007622f
C287 B.n247 VSUBS 0.007622f
C288 B.n248 VSUBS 0.007622f
C289 B.n249 VSUBS 0.007622f
C290 B.n250 VSUBS 0.007622f
C291 B.n251 VSUBS 0.007622f
C292 B.n252 VSUBS 0.007622f
C293 B.n253 VSUBS 0.007622f
C294 B.n254 VSUBS 0.007622f
C295 B.n255 VSUBS 0.007622f
C296 B.n256 VSUBS 0.007622f
C297 B.n257 VSUBS 0.007622f
C298 B.n258 VSUBS 0.007622f
C299 B.n259 VSUBS 0.007622f
C300 B.n260 VSUBS 0.007622f
C301 B.n261 VSUBS 0.007622f
C302 B.n262 VSUBS 0.007622f
C303 B.n263 VSUBS 0.007622f
C304 B.n264 VSUBS 0.007622f
C305 B.n265 VSUBS 0.007622f
C306 B.n266 VSUBS 0.007622f
C307 B.n267 VSUBS 0.007622f
C308 B.n268 VSUBS 0.007622f
C309 B.n269 VSUBS 0.007622f
C310 B.n270 VSUBS 0.007622f
C311 B.n271 VSUBS 0.007622f
C312 B.n272 VSUBS 0.007622f
C313 B.n273 VSUBS 0.007622f
C314 B.n274 VSUBS 0.007622f
C315 B.n275 VSUBS 0.007622f
C316 B.n276 VSUBS 0.007622f
C317 B.n277 VSUBS 0.016765f
C318 B.n278 VSUBS 0.016765f
C319 B.n279 VSUBS 0.017758f
C320 B.n280 VSUBS 0.007622f
C321 B.n281 VSUBS 0.007622f
C322 B.n282 VSUBS 0.007622f
C323 B.n283 VSUBS 0.007622f
C324 B.n284 VSUBS 0.007622f
C325 B.n285 VSUBS 0.007622f
C326 B.n286 VSUBS 0.007622f
C327 B.n287 VSUBS 0.007622f
C328 B.n288 VSUBS 0.007622f
C329 B.n289 VSUBS 0.007622f
C330 B.n290 VSUBS 0.007622f
C331 B.n291 VSUBS 0.007622f
C332 B.n292 VSUBS 0.007622f
C333 B.n293 VSUBS 0.007622f
C334 B.n294 VSUBS 0.007622f
C335 B.n295 VSUBS 0.007622f
C336 B.n296 VSUBS 0.007622f
C337 B.n297 VSUBS 0.007622f
C338 B.n298 VSUBS 0.007622f
C339 B.n299 VSUBS 0.007622f
C340 B.n300 VSUBS 0.007622f
C341 B.n301 VSUBS 0.007622f
C342 B.n302 VSUBS 0.007622f
C343 B.n303 VSUBS 0.005268f
C344 B.n304 VSUBS 0.01766f
C345 B.n305 VSUBS 0.006165f
C346 B.n306 VSUBS 0.007622f
C347 B.n307 VSUBS 0.007622f
C348 B.n308 VSUBS 0.007622f
C349 B.n309 VSUBS 0.007622f
C350 B.n310 VSUBS 0.007622f
C351 B.n311 VSUBS 0.007622f
C352 B.n312 VSUBS 0.007622f
C353 B.n313 VSUBS 0.007622f
C354 B.n314 VSUBS 0.007622f
C355 B.n315 VSUBS 0.007622f
C356 B.n316 VSUBS 0.007622f
C357 B.n317 VSUBS 0.006165f
C358 B.n318 VSUBS 0.007622f
C359 B.n319 VSUBS 0.007622f
C360 B.n320 VSUBS 0.007622f
C361 B.n321 VSUBS 0.007622f
C362 B.n322 VSUBS 0.007622f
C363 B.n323 VSUBS 0.007622f
C364 B.n324 VSUBS 0.007622f
C365 B.n325 VSUBS 0.007622f
C366 B.n326 VSUBS 0.007622f
C367 B.n327 VSUBS 0.007622f
C368 B.n328 VSUBS 0.007622f
C369 B.n329 VSUBS 0.007622f
C370 B.n330 VSUBS 0.007622f
C371 B.n331 VSUBS 0.007622f
C372 B.n332 VSUBS 0.007622f
C373 B.n333 VSUBS 0.007622f
C374 B.n334 VSUBS 0.007622f
C375 B.n335 VSUBS 0.007622f
C376 B.n336 VSUBS 0.007622f
C377 B.n337 VSUBS 0.007622f
C378 B.n338 VSUBS 0.007622f
C379 B.n339 VSUBS 0.007622f
C380 B.n340 VSUBS 0.007622f
C381 B.n341 VSUBS 0.007622f
C382 B.n342 VSUBS 0.007622f
C383 B.n343 VSUBS 0.017758f
C384 B.n344 VSUBS 0.016765f
C385 B.n345 VSUBS 0.016765f
C386 B.n346 VSUBS 0.007622f
C387 B.n347 VSUBS 0.007622f
C388 B.n348 VSUBS 0.007622f
C389 B.n349 VSUBS 0.007622f
C390 B.n350 VSUBS 0.007622f
C391 B.n351 VSUBS 0.007622f
C392 B.n352 VSUBS 0.007622f
C393 B.n353 VSUBS 0.007622f
C394 B.n354 VSUBS 0.007622f
C395 B.n355 VSUBS 0.007622f
C396 B.n356 VSUBS 0.007622f
C397 B.n357 VSUBS 0.007622f
C398 B.n358 VSUBS 0.007622f
C399 B.n359 VSUBS 0.007622f
C400 B.n360 VSUBS 0.007622f
C401 B.n361 VSUBS 0.007622f
C402 B.n362 VSUBS 0.007622f
C403 B.n363 VSUBS 0.007622f
C404 B.n364 VSUBS 0.007622f
C405 B.n365 VSUBS 0.007622f
C406 B.n366 VSUBS 0.007622f
C407 B.n367 VSUBS 0.007622f
C408 B.n368 VSUBS 0.007622f
C409 B.n369 VSUBS 0.007622f
C410 B.n370 VSUBS 0.007622f
C411 B.n371 VSUBS 0.007622f
C412 B.n372 VSUBS 0.007622f
C413 B.n373 VSUBS 0.007622f
C414 B.n374 VSUBS 0.007622f
C415 B.n375 VSUBS 0.007622f
C416 B.n376 VSUBS 0.007622f
C417 B.n377 VSUBS 0.007622f
C418 B.n378 VSUBS 0.007622f
C419 B.n379 VSUBS 0.009946f
C420 B.n380 VSUBS 0.010596f
C421 B.n381 VSUBS 0.02107f
C422 VDD1.t1 VSUBS 0.330891f
C423 VDD1.t3 VSUBS 0.330614f
C424 VDD1.t2 VSUBS 0.042246f
C425 VDD1.t0 VSUBS 0.042246f
C426 VDD1.n0 VSUBS 0.236318f
C427 VDD1.n1 VSUBS 1.25391f
C428 VDD1.t5 VSUBS 0.042246f
C429 VDD1.t4 VSUBS 0.042246f
C430 VDD1.n2 VSUBS 0.235743f
C431 VDD1.n3 VSUBS 1.10615f
C432 VP.n0 VSUBS 0.07145f
C433 VP.t3 VSUBS 0.503703f
C434 VP.n1 VSUBS 0.066642f
C435 VP.n2 VSUBS 0.294276f
C436 VP.t1 VSUBS 0.590127f
C437 VP.t0 VSUBS 0.503703f
C438 VP.t4 VSUBS 0.644764f
C439 VP.n3 VSUBS 0.300245f
C440 VP.n4 VSUBS 0.320024f
C441 VP.n5 VSUBS 0.066642f
C442 VP.n6 VSUBS 0.320811f
C443 VP.n7 VSUBS 1.73285f
C444 VP.t2 VSUBS 0.590127f
C445 VP.n8 VSUBS 0.320811f
C446 VP.n9 VSUBS 1.78596f
C447 VP.n10 VSUBS 0.07145f
C448 VP.n11 VSUBS 0.053546f
C449 VP.n12 VSUBS 0.28487f
C450 VP.n13 VSUBS 0.066642f
C451 VP.t5 VSUBS 0.590127f
C452 VP.n14 VSUBS 0.320811f
C453 VP.n15 VSUBS 0.050148f
C454 VDD2.t4 VSUBS 0.343727f
C455 VDD2.t0 VSUBS 0.043922f
C456 VDD2.t5 VSUBS 0.043922f
C457 VDD2.n0 VSUBS 0.245691f
C458 VDD2.n1 VSUBS 1.25257f
C459 VDD2.t1 VSUBS 0.341877f
C460 VDD2.n2 VSUBS 1.14075f
C461 VDD2.t2 VSUBS 0.043922f
C462 VDD2.t3 VSUBS 0.043922f
C463 VDD2.n3 VSUBS 0.24568f
C464 VTAIL.t7 VSUBS 0.064458f
C465 VTAIL.t10 VSUBS 0.064458f
C466 VTAIL.n0 VSUBS 0.310036f
C467 VTAIL.n1 VSUBS 0.43806f
C468 VTAIL.t0 VSUBS 0.45117f
C469 VTAIL.n2 VSUBS 0.53584f
C470 VTAIL.t3 VSUBS 0.064458f
C471 VTAIL.t2 VSUBS 0.064458f
C472 VTAIL.n3 VSUBS 0.310036f
C473 VTAIL.n4 VSUBS 1.14403f
C474 VTAIL.t11 VSUBS 0.064458f
C475 VTAIL.t8 VSUBS 0.064458f
C476 VTAIL.n5 VSUBS 0.310037f
C477 VTAIL.n6 VSUBS 1.14403f
C478 VTAIL.t6 VSUBS 0.451172f
C479 VTAIL.n7 VSUBS 0.535837f
C480 VTAIL.t5 VSUBS 0.064458f
C481 VTAIL.t4 VSUBS 0.064458f
C482 VTAIL.n8 VSUBS 0.310037f
C483 VTAIL.n9 VSUBS 0.501177f
C484 VTAIL.t1 VSUBS 0.45117f
C485 VTAIL.n10 VSUBS 1.08871f
C486 VTAIL.t9 VSUBS 0.45117f
C487 VTAIL.n11 VSUBS 1.06184f
C488 VN.n0 VSUBS 0.222031f
C489 VN.t5 VSUBS 0.380044f
C490 VN.t1 VSUBS 0.486475f
C491 VN.n1 VSUBS 0.226535f
C492 VN.n2 VSUBS 0.241458f
C493 VN.n3 VSUBS 0.050281f
C494 VN.t0 VSUBS 0.445252f
C495 VN.n4 VSUBS 0.242052f
C496 VN.n5 VSUBS 0.037836f
C497 VN.n6 VSUBS 0.222031f
C498 VN.t3 VSUBS 0.380044f
C499 VN.t2 VSUBS 0.486475f
C500 VN.n7 VSUBS 0.226535f
C501 VN.n8 VSUBS 0.241458f
C502 VN.n9 VSUBS 0.050281f
C503 VN.t4 VSUBS 0.445252f
C504 VN.n10 VSUBS 0.242052f
C505 VN.n11 VSUBS 1.33073f
.ends

