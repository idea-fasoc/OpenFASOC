* NGSPICE file created from diff_pair_sample_0718.ext - technology: sky130A

.subckt diff_pair_sample_0718 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t4 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=2.69775 pd=16.68 as=2.69775 ps=16.68 w=16.35 l=3.18
X1 VDD2.t5 VN.t0 VTAIL.t3 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=6.3765 pd=33.48 as=2.69775 ps=16.68 w=16.35 l=3.18
X2 VDD2.t4 VN.t1 VTAIL.t4 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=6.3765 pd=33.48 as=2.69775 ps=16.68 w=16.35 l=3.18
X3 B.t11 B.t9 B.t10 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=6.3765 pd=33.48 as=0 ps=0 w=16.35 l=3.18
X4 VDD1.t3 VP.t1 VTAIL.t10 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=6.3765 pd=33.48 as=2.69775 ps=16.68 w=16.35 l=3.18
X5 VDD2.t3 VN.t2 VTAIL.t0 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=2.69775 pd=16.68 as=6.3765 ps=33.48 w=16.35 l=3.18
X6 VDD2.t2 VN.t3 VTAIL.t5 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=2.69775 pd=16.68 as=6.3765 ps=33.48 w=16.35 l=3.18
X7 B.t8 B.t6 B.t7 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=6.3765 pd=33.48 as=0 ps=0 w=16.35 l=3.18
X8 VTAIL.t9 VP.t2 VDD1.t2 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=2.69775 pd=16.68 as=2.69775 ps=16.68 w=16.35 l=3.18
X9 VTAIL.t2 VN.t4 VDD2.t1 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=2.69775 pd=16.68 as=2.69775 ps=16.68 w=16.35 l=3.18
X10 B.t5 B.t3 B.t4 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=6.3765 pd=33.48 as=0 ps=0 w=16.35 l=3.18
X11 B.t2 B.t0 B.t1 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=6.3765 pd=33.48 as=0 ps=0 w=16.35 l=3.18
X12 VDD1.t0 VP.t3 VTAIL.t8 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=6.3765 pd=33.48 as=2.69775 ps=16.68 w=16.35 l=3.18
X13 VTAIL.t1 VN.t5 VDD2.t0 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=2.69775 pd=16.68 as=2.69775 ps=16.68 w=16.35 l=3.18
X14 VDD1.t5 VP.t4 VTAIL.t7 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=2.69775 pd=16.68 as=6.3765 ps=33.48 w=16.35 l=3.18
X15 VDD1.t1 VP.t5 VTAIL.t6 w_n3778_n4238# sky130_fd_pr__pfet_01v8 ad=2.69775 pd=16.68 as=6.3765 ps=33.48 w=16.35 l=3.18
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n23 VP.n10 161.3
R6 VP.n25 VP.n24 161.3
R7 VP.n49 VP.n48 161.3
R8 VP.n47 VP.n1 161.3
R9 VP.n46 VP.n45 161.3
R10 VP.n44 VP.n2 161.3
R11 VP.n43 VP.n42 161.3
R12 VP.n41 VP.n3 161.3
R13 VP.n40 VP.n39 161.3
R14 VP.n38 VP.n37 161.3
R15 VP.n36 VP.n5 161.3
R16 VP.n35 VP.n34 161.3
R17 VP.n33 VP.n6 161.3
R18 VP.n32 VP.n31 161.3
R19 VP.n30 VP.n7 161.3
R20 VP.n29 VP.n28 161.3
R21 VP.n14 VP.t3 156.618
R22 VP.n8 VP.t1 123.91
R23 VP.n4 VP.t2 123.91
R24 VP.n0 VP.t4 123.91
R25 VP.n9 VP.t5 123.91
R26 VP.n13 VP.t0 123.91
R27 VP.n27 VP.n8 77.3446
R28 VP.n50 VP.n0 77.3446
R29 VP.n26 VP.n9 77.3446
R30 VP.n14 VP.n13 62.0352
R31 VP.n27 VP.n26 54.2986
R32 VP.n31 VP.n6 40.979
R33 VP.n46 VP.n2 40.979
R34 VP.n22 VP.n11 40.979
R35 VP.n35 VP.n6 40.0078
R36 VP.n42 VP.n2 40.0078
R37 VP.n18 VP.n11 40.0078
R38 VP.n30 VP.n29 24.4675
R39 VP.n31 VP.n30 24.4675
R40 VP.n36 VP.n35 24.4675
R41 VP.n37 VP.n36 24.4675
R42 VP.n41 VP.n40 24.4675
R43 VP.n42 VP.n41 24.4675
R44 VP.n47 VP.n46 24.4675
R45 VP.n48 VP.n47 24.4675
R46 VP.n23 VP.n22 24.4675
R47 VP.n24 VP.n23 24.4675
R48 VP.n17 VP.n16 24.4675
R49 VP.n18 VP.n17 24.4675
R50 VP.n29 VP.n8 12.7233
R51 VP.n48 VP.n0 12.7233
R52 VP.n24 VP.n9 12.7233
R53 VP.n37 VP.n4 12.234
R54 VP.n40 VP.n4 12.234
R55 VP.n16 VP.n13 12.234
R56 VP.n15 VP.n14 4.25366
R57 VP.n26 VP.n25 0.354971
R58 VP.n28 VP.n27 0.354971
R59 VP.n50 VP.n49 0.354971
R60 VP VP.n50 0.26696
R61 VP.n15 VP.n12 0.189894
R62 VP.n19 VP.n12 0.189894
R63 VP.n20 VP.n19 0.189894
R64 VP.n21 VP.n20 0.189894
R65 VP.n21 VP.n10 0.189894
R66 VP.n25 VP.n10 0.189894
R67 VP.n28 VP.n7 0.189894
R68 VP.n32 VP.n7 0.189894
R69 VP.n33 VP.n32 0.189894
R70 VP.n34 VP.n33 0.189894
R71 VP.n34 VP.n5 0.189894
R72 VP.n38 VP.n5 0.189894
R73 VP.n39 VP.n38 0.189894
R74 VP.n39 VP.n3 0.189894
R75 VP.n43 VP.n3 0.189894
R76 VP.n44 VP.n43 0.189894
R77 VP.n45 VP.n44 0.189894
R78 VP.n45 VP.n1 0.189894
R79 VP.n49 VP.n1 0.189894
R80 VDD1 VDD1.t0 72.1617
R81 VDD1.n1 VDD1.t3 72.0479
R82 VDD1.n1 VDD1.n0 68.5469
R83 VDD1.n3 VDD1.n2 67.8458
R84 VDD1.n3 VDD1.n1 49.7401
R85 VDD1.n2 VDD1.t4 1.98857
R86 VDD1.n2 VDD1.t1 1.98857
R87 VDD1.n0 VDD1.t2 1.98857
R88 VDD1.n0 VDD1.t5 1.98857
R89 VDD1 VDD1.n3 0.698776
R90 VTAIL.n7 VTAIL.t5 53.1553
R91 VTAIL.n11 VTAIL.t0 53.1551
R92 VTAIL.n2 VTAIL.t7 53.1551
R93 VTAIL.n10 VTAIL.t6 53.1551
R94 VTAIL.n9 VTAIL.n8 51.1672
R95 VTAIL.n6 VTAIL.n5 51.1672
R96 VTAIL.n1 VTAIL.n0 51.167
R97 VTAIL.n4 VTAIL.n3 51.167
R98 VTAIL.n6 VTAIL.n4 32.5134
R99 VTAIL.n11 VTAIL.n10 29.4876
R100 VTAIL.n7 VTAIL.n6 3.02636
R101 VTAIL.n10 VTAIL.n9 3.02636
R102 VTAIL.n4 VTAIL.n2 3.02636
R103 VTAIL VTAIL.n11 2.21171
R104 VTAIL.n0 VTAIL.t4 1.98857
R105 VTAIL.n0 VTAIL.t1 1.98857
R106 VTAIL.n3 VTAIL.t10 1.98857
R107 VTAIL.n3 VTAIL.t9 1.98857
R108 VTAIL.n8 VTAIL.t8 1.98857
R109 VTAIL.n8 VTAIL.t11 1.98857
R110 VTAIL.n5 VTAIL.t3 1.98857
R111 VTAIL.n5 VTAIL.t2 1.98857
R112 VTAIL.n9 VTAIL.n7 1.98326
R113 VTAIL.n2 VTAIL.n1 1.98326
R114 VTAIL VTAIL.n1 0.815155
R115 VN.n34 VN.n33 161.3
R116 VN.n32 VN.n19 161.3
R117 VN.n31 VN.n30 161.3
R118 VN.n29 VN.n20 161.3
R119 VN.n28 VN.n27 161.3
R120 VN.n26 VN.n21 161.3
R121 VN.n25 VN.n24 161.3
R122 VN.n16 VN.n15 161.3
R123 VN.n14 VN.n1 161.3
R124 VN.n13 VN.n12 161.3
R125 VN.n11 VN.n2 161.3
R126 VN.n10 VN.n9 161.3
R127 VN.n8 VN.n3 161.3
R128 VN.n7 VN.n6 161.3
R129 VN.n23 VN.t3 156.618
R130 VN.n5 VN.t1 156.618
R131 VN.n4 VN.t5 123.91
R132 VN.n0 VN.t2 123.91
R133 VN.n22 VN.t4 123.91
R134 VN.n18 VN.t0 123.91
R135 VN.n17 VN.n0 77.3446
R136 VN.n35 VN.n18 77.3446
R137 VN.n5 VN.n4 62.0351
R138 VN.n23 VN.n22 62.0351
R139 VN VN.n35 54.4639
R140 VN.n13 VN.n2 40.979
R141 VN.n31 VN.n20 40.979
R142 VN.n9 VN.n2 40.0078
R143 VN.n27 VN.n20 40.0078
R144 VN.n8 VN.n7 24.4675
R145 VN.n9 VN.n8 24.4675
R146 VN.n14 VN.n13 24.4675
R147 VN.n15 VN.n14 24.4675
R148 VN.n27 VN.n26 24.4675
R149 VN.n26 VN.n25 24.4675
R150 VN.n33 VN.n32 24.4675
R151 VN.n32 VN.n31 24.4675
R152 VN.n15 VN.n0 12.7233
R153 VN.n33 VN.n18 12.7233
R154 VN.n7 VN.n4 12.234
R155 VN.n25 VN.n22 12.234
R156 VN.n24 VN.n23 4.25368
R157 VN.n6 VN.n5 4.25368
R158 VN.n35 VN.n34 0.354971
R159 VN.n17 VN.n16 0.354971
R160 VN VN.n17 0.26696
R161 VN.n34 VN.n19 0.189894
R162 VN.n30 VN.n19 0.189894
R163 VN.n30 VN.n29 0.189894
R164 VN.n29 VN.n28 0.189894
R165 VN.n28 VN.n21 0.189894
R166 VN.n24 VN.n21 0.189894
R167 VN.n6 VN.n3 0.189894
R168 VN.n10 VN.n3 0.189894
R169 VN.n11 VN.n10 0.189894
R170 VN.n12 VN.n11 0.189894
R171 VN.n12 VN.n1 0.189894
R172 VN.n16 VN.n1 0.189894
R173 VDD2.n1 VDD2.t4 72.0479
R174 VDD2.n2 VDD2.t5 69.8341
R175 VDD2.n1 VDD2.n0 68.5469
R176 VDD2 VDD2.n3 68.5441
R177 VDD2.n2 VDD2.n1 47.6442
R178 VDD2 VDD2.n2 2.32809
R179 VDD2.n3 VDD2.t1 1.98857
R180 VDD2.n3 VDD2.t2 1.98857
R181 VDD2.n0 VDD2.t0 1.98857
R182 VDD2.n0 VDD2.t3 1.98857
R183 B.n478 B.n477 585
R184 B.n476 B.n141 585
R185 B.n475 B.n474 585
R186 B.n473 B.n142 585
R187 B.n472 B.n471 585
R188 B.n470 B.n143 585
R189 B.n469 B.n468 585
R190 B.n467 B.n144 585
R191 B.n466 B.n465 585
R192 B.n464 B.n145 585
R193 B.n463 B.n462 585
R194 B.n461 B.n146 585
R195 B.n460 B.n459 585
R196 B.n458 B.n147 585
R197 B.n457 B.n456 585
R198 B.n455 B.n148 585
R199 B.n454 B.n453 585
R200 B.n452 B.n149 585
R201 B.n451 B.n450 585
R202 B.n449 B.n150 585
R203 B.n448 B.n447 585
R204 B.n446 B.n151 585
R205 B.n445 B.n444 585
R206 B.n443 B.n152 585
R207 B.n442 B.n441 585
R208 B.n440 B.n153 585
R209 B.n439 B.n438 585
R210 B.n437 B.n154 585
R211 B.n436 B.n435 585
R212 B.n434 B.n155 585
R213 B.n433 B.n432 585
R214 B.n431 B.n156 585
R215 B.n430 B.n429 585
R216 B.n428 B.n157 585
R217 B.n427 B.n426 585
R218 B.n425 B.n158 585
R219 B.n424 B.n423 585
R220 B.n422 B.n159 585
R221 B.n421 B.n420 585
R222 B.n419 B.n160 585
R223 B.n418 B.n417 585
R224 B.n416 B.n161 585
R225 B.n415 B.n414 585
R226 B.n413 B.n162 585
R227 B.n412 B.n411 585
R228 B.n410 B.n163 585
R229 B.n409 B.n408 585
R230 B.n407 B.n164 585
R231 B.n406 B.n405 585
R232 B.n404 B.n165 585
R233 B.n403 B.n402 585
R234 B.n401 B.n166 585
R235 B.n400 B.n399 585
R236 B.n398 B.n167 585
R237 B.n397 B.n396 585
R238 B.n392 B.n168 585
R239 B.n391 B.n390 585
R240 B.n389 B.n169 585
R241 B.n388 B.n387 585
R242 B.n386 B.n170 585
R243 B.n385 B.n384 585
R244 B.n383 B.n171 585
R245 B.n382 B.n381 585
R246 B.n380 B.n172 585
R247 B.n378 B.n377 585
R248 B.n376 B.n175 585
R249 B.n375 B.n374 585
R250 B.n373 B.n176 585
R251 B.n372 B.n371 585
R252 B.n370 B.n177 585
R253 B.n369 B.n368 585
R254 B.n367 B.n178 585
R255 B.n366 B.n365 585
R256 B.n364 B.n179 585
R257 B.n363 B.n362 585
R258 B.n361 B.n180 585
R259 B.n360 B.n359 585
R260 B.n358 B.n181 585
R261 B.n357 B.n356 585
R262 B.n355 B.n182 585
R263 B.n354 B.n353 585
R264 B.n352 B.n183 585
R265 B.n351 B.n350 585
R266 B.n349 B.n184 585
R267 B.n348 B.n347 585
R268 B.n346 B.n185 585
R269 B.n345 B.n344 585
R270 B.n343 B.n186 585
R271 B.n342 B.n341 585
R272 B.n340 B.n187 585
R273 B.n339 B.n338 585
R274 B.n337 B.n188 585
R275 B.n336 B.n335 585
R276 B.n334 B.n189 585
R277 B.n333 B.n332 585
R278 B.n331 B.n190 585
R279 B.n330 B.n329 585
R280 B.n328 B.n191 585
R281 B.n327 B.n326 585
R282 B.n325 B.n192 585
R283 B.n324 B.n323 585
R284 B.n322 B.n193 585
R285 B.n321 B.n320 585
R286 B.n319 B.n194 585
R287 B.n318 B.n317 585
R288 B.n316 B.n195 585
R289 B.n315 B.n314 585
R290 B.n313 B.n196 585
R291 B.n312 B.n311 585
R292 B.n310 B.n197 585
R293 B.n309 B.n308 585
R294 B.n307 B.n198 585
R295 B.n306 B.n305 585
R296 B.n304 B.n199 585
R297 B.n303 B.n302 585
R298 B.n301 B.n200 585
R299 B.n300 B.n299 585
R300 B.n298 B.n201 585
R301 B.n479 B.n140 585
R302 B.n481 B.n480 585
R303 B.n482 B.n139 585
R304 B.n484 B.n483 585
R305 B.n485 B.n138 585
R306 B.n487 B.n486 585
R307 B.n488 B.n137 585
R308 B.n490 B.n489 585
R309 B.n491 B.n136 585
R310 B.n493 B.n492 585
R311 B.n494 B.n135 585
R312 B.n496 B.n495 585
R313 B.n497 B.n134 585
R314 B.n499 B.n498 585
R315 B.n500 B.n133 585
R316 B.n502 B.n501 585
R317 B.n503 B.n132 585
R318 B.n505 B.n504 585
R319 B.n506 B.n131 585
R320 B.n508 B.n507 585
R321 B.n509 B.n130 585
R322 B.n511 B.n510 585
R323 B.n512 B.n129 585
R324 B.n514 B.n513 585
R325 B.n515 B.n128 585
R326 B.n517 B.n516 585
R327 B.n518 B.n127 585
R328 B.n520 B.n519 585
R329 B.n521 B.n126 585
R330 B.n523 B.n522 585
R331 B.n524 B.n125 585
R332 B.n526 B.n525 585
R333 B.n527 B.n124 585
R334 B.n529 B.n528 585
R335 B.n530 B.n123 585
R336 B.n532 B.n531 585
R337 B.n533 B.n122 585
R338 B.n535 B.n534 585
R339 B.n536 B.n121 585
R340 B.n538 B.n537 585
R341 B.n539 B.n120 585
R342 B.n541 B.n540 585
R343 B.n542 B.n119 585
R344 B.n544 B.n543 585
R345 B.n545 B.n118 585
R346 B.n547 B.n546 585
R347 B.n548 B.n117 585
R348 B.n550 B.n549 585
R349 B.n551 B.n116 585
R350 B.n553 B.n552 585
R351 B.n554 B.n115 585
R352 B.n556 B.n555 585
R353 B.n557 B.n114 585
R354 B.n559 B.n558 585
R355 B.n560 B.n113 585
R356 B.n562 B.n561 585
R357 B.n563 B.n112 585
R358 B.n565 B.n564 585
R359 B.n566 B.n111 585
R360 B.n568 B.n567 585
R361 B.n569 B.n110 585
R362 B.n571 B.n570 585
R363 B.n572 B.n109 585
R364 B.n574 B.n573 585
R365 B.n575 B.n108 585
R366 B.n577 B.n576 585
R367 B.n578 B.n107 585
R368 B.n580 B.n579 585
R369 B.n581 B.n106 585
R370 B.n583 B.n582 585
R371 B.n584 B.n105 585
R372 B.n586 B.n585 585
R373 B.n587 B.n104 585
R374 B.n589 B.n588 585
R375 B.n590 B.n103 585
R376 B.n592 B.n591 585
R377 B.n593 B.n102 585
R378 B.n595 B.n594 585
R379 B.n596 B.n101 585
R380 B.n598 B.n597 585
R381 B.n599 B.n100 585
R382 B.n601 B.n600 585
R383 B.n602 B.n99 585
R384 B.n604 B.n603 585
R385 B.n605 B.n98 585
R386 B.n607 B.n606 585
R387 B.n608 B.n97 585
R388 B.n610 B.n609 585
R389 B.n611 B.n96 585
R390 B.n613 B.n612 585
R391 B.n614 B.n95 585
R392 B.n616 B.n615 585
R393 B.n617 B.n94 585
R394 B.n619 B.n618 585
R395 B.n620 B.n93 585
R396 B.n622 B.n621 585
R397 B.n623 B.n92 585
R398 B.n625 B.n624 585
R399 B.n626 B.n91 585
R400 B.n628 B.n627 585
R401 B.n806 B.n805 585
R402 B.n804 B.n27 585
R403 B.n803 B.n802 585
R404 B.n801 B.n28 585
R405 B.n800 B.n799 585
R406 B.n798 B.n29 585
R407 B.n797 B.n796 585
R408 B.n795 B.n30 585
R409 B.n794 B.n793 585
R410 B.n792 B.n31 585
R411 B.n791 B.n790 585
R412 B.n789 B.n32 585
R413 B.n788 B.n787 585
R414 B.n786 B.n33 585
R415 B.n785 B.n784 585
R416 B.n783 B.n34 585
R417 B.n782 B.n781 585
R418 B.n780 B.n35 585
R419 B.n779 B.n778 585
R420 B.n777 B.n36 585
R421 B.n776 B.n775 585
R422 B.n774 B.n37 585
R423 B.n773 B.n772 585
R424 B.n771 B.n38 585
R425 B.n770 B.n769 585
R426 B.n768 B.n39 585
R427 B.n767 B.n766 585
R428 B.n765 B.n40 585
R429 B.n764 B.n763 585
R430 B.n762 B.n41 585
R431 B.n761 B.n760 585
R432 B.n759 B.n42 585
R433 B.n758 B.n757 585
R434 B.n756 B.n43 585
R435 B.n755 B.n754 585
R436 B.n753 B.n44 585
R437 B.n752 B.n751 585
R438 B.n750 B.n45 585
R439 B.n749 B.n748 585
R440 B.n747 B.n46 585
R441 B.n746 B.n745 585
R442 B.n744 B.n47 585
R443 B.n743 B.n742 585
R444 B.n741 B.n48 585
R445 B.n740 B.n739 585
R446 B.n738 B.n49 585
R447 B.n737 B.n736 585
R448 B.n735 B.n50 585
R449 B.n734 B.n733 585
R450 B.n732 B.n51 585
R451 B.n731 B.n730 585
R452 B.n729 B.n52 585
R453 B.n728 B.n727 585
R454 B.n726 B.n53 585
R455 B.n724 B.n723 585
R456 B.n722 B.n56 585
R457 B.n721 B.n720 585
R458 B.n719 B.n57 585
R459 B.n718 B.n717 585
R460 B.n716 B.n58 585
R461 B.n715 B.n714 585
R462 B.n713 B.n59 585
R463 B.n712 B.n711 585
R464 B.n710 B.n60 585
R465 B.n709 B.n708 585
R466 B.n707 B.n61 585
R467 B.n706 B.n705 585
R468 B.n704 B.n65 585
R469 B.n703 B.n702 585
R470 B.n701 B.n66 585
R471 B.n700 B.n699 585
R472 B.n698 B.n67 585
R473 B.n697 B.n696 585
R474 B.n695 B.n68 585
R475 B.n694 B.n693 585
R476 B.n692 B.n69 585
R477 B.n691 B.n690 585
R478 B.n689 B.n70 585
R479 B.n688 B.n687 585
R480 B.n686 B.n71 585
R481 B.n685 B.n684 585
R482 B.n683 B.n72 585
R483 B.n682 B.n681 585
R484 B.n680 B.n73 585
R485 B.n679 B.n678 585
R486 B.n677 B.n74 585
R487 B.n676 B.n675 585
R488 B.n674 B.n75 585
R489 B.n673 B.n672 585
R490 B.n671 B.n76 585
R491 B.n670 B.n669 585
R492 B.n668 B.n77 585
R493 B.n667 B.n666 585
R494 B.n665 B.n78 585
R495 B.n664 B.n663 585
R496 B.n662 B.n79 585
R497 B.n661 B.n660 585
R498 B.n659 B.n80 585
R499 B.n658 B.n657 585
R500 B.n656 B.n81 585
R501 B.n655 B.n654 585
R502 B.n653 B.n82 585
R503 B.n652 B.n651 585
R504 B.n650 B.n83 585
R505 B.n649 B.n648 585
R506 B.n647 B.n84 585
R507 B.n646 B.n645 585
R508 B.n644 B.n85 585
R509 B.n643 B.n642 585
R510 B.n641 B.n86 585
R511 B.n640 B.n639 585
R512 B.n638 B.n87 585
R513 B.n637 B.n636 585
R514 B.n635 B.n88 585
R515 B.n634 B.n633 585
R516 B.n632 B.n89 585
R517 B.n631 B.n630 585
R518 B.n629 B.n90 585
R519 B.n807 B.n26 585
R520 B.n809 B.n808 585
R521 B.n810 B.n25 585
R522 B.n812 B.n811 585
R523 B.n813 B.n24 585
R524 B.n815 B.n814 585
R525 B.n816 B.n23 585
R526 B.n818 B.n817 585
R527 B.n819 B.n22 585
R528 B.n821 B.n820 585
R529 B.n822 B.n21 585
R530 B.n824 B.n823 585
R531 B.n825 B.n20 585
R532 B.n827 B.n826 585
R533 B.n828 B.n19 585
R534 B.n830 B.n829 585
R535 B.n831 B.n18 585
R536 B.n833 B.n832 585
R537 B.n834 B.n17 585
R538 B.n836 B.n835 585
R539 B.n837 B.n16 585
R540 B.n839 B.n838 585
R541 B.n840 B.n15 585
R542 B.n842 B.n841 585
R543 B.n843 B.n14 585
R544 B.n845 B.n844 585
R545 B.n846 B.n13 585
R546 B.n848 B.n847 585
R547 B.n849 B.n12 585
R548 B.n851 B.n850 585
R549 B.n852 B.n11 585
R550 B.n854 B.n853 585
R551 B.n855 B.n10 585
R552 B.n857 B.n856 585
R553 B.n858 B.n9 585
R554 B.n860 B.n859 585
R555 B.n861 B.n8 585
R556 B.n863 B.n862 585
R557 B.n864 B.n7 585
R558 B.n866 B.n865 585
R559 B.n867 B.n6 585
R560 B.n869 B.n868 585
R561 B.n870 B.n5 585
R562 B.n872 B.n871 585
R563 B.n873 B.n4 585
R564 B.n875 B.n874 585
R565 B.n876 B.n3 585
R566 B.n878 B.n877 585
R567 B.n879 B.n0 585
R568 B.n2 B.n1 585
R569 B.n226 B.n225 585
R570 B.n228 B.n227 585
R571 B.n229 B.n224 585
R572 B.n231 B.n230 585
R573 B.n232 B.n223 585
R574 B.n234 B.n233 585
R575 B.n235 B.n222 585
R576 B.n237 B.n236 585
R577 B.n238 B.n221 585
R578 B.n240 B.n239 585
R579 B.n241 B.n220 585
R580 B.n243 B.n242 585
R581 B.n244 B.n219 585
R582 B.n246 B.n245 585
R583 B.n247 B.n218 585
R584 B.n249 B.n248 585
R585 B.n250 B.n217 585
R586 B.n252 B.n251 585
R587 B.n253 B.n216 585
R588 B.n255 B.n254 585
R589 B.n256 B.n215 585
R590 B.n258 B.n257 585
R591 B.n259 B.n214 585
R592 B.n261 B.n260 585
R593 B.n262 B.n213 585
R594 B.n264 B.n263 585
R595 B.n265 B.n212 585
R596 B.n267 B.n266 585
R597 B.n268 B.n211 585
R598 B.n270 B.n269 585
R599 B.n271 B.n210 585
R600 B.n273 B.n272 585
R601 B.n274 B.n209 585
R602 B.n276 B.n275 585
R603 B.n277 B.n208 585
R604 B.n279 B.n278 585
R605 B.n280 B.n207 585
R606 B.n282 B.n281 585
R607 B.n283 B.n206 585
R608 B.n285 B.n284 585
R609 B.n286 B.n205 585
R610 B.n288 B.n287 585
R611 B.n289 B.n204 585
R612 B.n291 B.n290 585
R613 B.n292 B.n203 585
R614 B.n294 B.n293 585
R615 B.n295 B.n202 585
R616 B.n297 B.n296 585
R617 B.n298 B.n297 516.524
R618 B.n477 B.n140 516.524
R619 B.n627 B.n90 516.524
R620 B.n807 B.n806 516.524
R621 B.n173 B.t3 332.692
R622 B.n393 B.t9 332.692
R623 B.n62 B.t0 332.692
R624 B.n54 B.t6 332.692
R625 B.n881 B.n880 256.663
R626 B.n880 B.n879 235.042
R627 B.n880 B.n2 235.042
R628 B.n393 B.t10 175.038
R629 B.n62 B.t2 175.038
R630 B.n173 B.t4 175.018
R631 B.n54 B.t8 175.018
R632 B.n299 B.n298 163.367
R633 B.n299 B.n200 163.367
R634 B.n303 B.n200 163.367
R635 B.n304 B.n303 163.367
R636 B.n305 B.n304 163.367
R637 B.n305 B.n198 163.367
R638 B.n309 B.n198 163.367
R639 B.n310 B.n309 163.367
R640 B.n311 B.n310 163.367
R641 B.n311 B.n196 163.367
R642 B.n315 B.n196 163.367
R643 B.n316 B.n315 163.367
R644 B.n317 B.n316 163.367
R645 B.n317 B.n194 163.367
R646 B.n321 B.n194 163.367
R647 B.n322 B.n321 163.367
R648 B.n323 B.n322 163.367
R649 B.n323 B.n192 163.367
R650 B.n327 B.n192 163.367
R651 B.n328 B.n327 163.367
R652 B.n329 B.n328 163.367
R653 B.n329 B.n190 163.367
R654 B.n333 B.n190 163.367
R655 B.n334 B.n333 163.367
R656 B.n335 B.n334 163.367
R657 B.n335 B.n188 163.367
R658 B.n339 B.n188 163.367
R659 B.n340 B.n339 163.367
R660 B.n341 B.n340 163.367
R661 B.n341 B.n186 163.367
R662 B.n345 B.n186 163.367
R663 B.n346 B.n345 163.367
R664 B.n347 B.n346 163.367
R665 B.n347 B.n184 163.367
R666 B.n351 B.n184 163.367
R667 B.n352 B.n351 163.367
R668 B.n353 B.n352 163.367
R669 B.n353 B.n182 163.367
R670 B.n357 B.n182 163.367
R671 B.n358 B.n357 163.367
R672 B.n359 B.n358 163.367
R673 B.n359 B.n180 163.367
R674 B.n363 B.n180 163.367
R675 B.n364 B.n363 163.367
R676 B.n365 B.n364 163.367
R677 B.n365 B.n178 163.367
R678 B.n369 B.n178 163.367
R679 B.n370 B.n369 163.367
R680 B.n371 B.n370 163.367
R681 B.n371 B.n176 163.367
R682 B.n375 B.n176 163.367
R683 B.n376 B.n375 163.367
R684 B.n377 B.n376 163.367
R685 B.n377 B.n172 163.367
R686 B.n382 B.n172 163.367
R687 B.n383 B.n382 163.367
R688 B.n384 B.n383 163.367
R689 B.n384 B.n170 163.367
R690 B.n388 B.n170 163.367
R691 B.n389 B.n388 163.367
R692 B.n390 B.n389 163.367
R693 B.n390 B.n168 163.367
R694 B.n397 B.n168 163.367
R695 B.n398 B.n397 163.367
R696 B.n399 B.n398 163.367
R697 B.n399 B.n166 163.367
R698 B.n403 B.n166 163.367
R699 B.n404 B.n403 163.367
R700 B.n405 B.n404 163.367
R701 B.n405 B.n164 163.367
R702 B.n409 B.n164 163.367
R703 B.n410 B.n409 163.367
R704 B.n411 B.n410 163.367
R705 B.n411 B.n162 163.367
R706 B.n415 B.n162 163.367
R707 B.n416 B.n415 163.367
R708 B.n417 B.n416 163.367
R709 B.n417 B.n160 163.367
R710 B.n421 B.n160 163.367
R711 B.n422 B.n421 163.367
R712 B.n423 B.n422 163.367
R713 B.n423 B.n158 163.367
R714 B.n427 B.n158 163.367
R715 B.n428 B.n427 163.367
R716 B.n429 B.n428 163.367
R717 B.n429 B.n156 163.367
R718 B.n433 B.n156 163.367
R719 B.n434 B.n433 163.367
R720 B.n435 B.n434 163.367
R721 B.n435 B.n154 163.367
R722 B.n439 B.n154 163.367
R723 B.n440 B.n439 163.367
R724 B.n441 B.n440 163.367
R725 B.n441 B.n152 163.367
R726 B.n445 B.n152 163.367
R727 B.n446 B.n445 163.367
R728 B.n447 B.n446 163.367
R729 B.n447 B.n150 163.367
R730 B.n451 B.n150 163.367
R731 B.n452 B.n451 163.367
R732 B.n453 B.n452 163.367
R733 B.n453 B.n148 163.367
R734 B.n457 B.n148 163.367
R735 B.n458 B.n457 163.367
R736 B.n459 B.n458 163.367
R737 B.n459 B.n146 163.367
R738 B.n463 B.n146 163.367
R739 B.n464 B.n463 163.367
R740 B.n465 B.n464 163.367
R741 B.n465 B.n144 163.367
R742 B.n469 B.n144 163.367
R743 B.n470 B.n469 163.367
R744 B.n471 B.n470 163.367
R745 B.n471 B.n142 163.367
R746 B.n475 B.n142 163.367
R747 B.n476 B.n475 163.367
R748 B.n477 B.n476 163.367
R749 B.n627 B.n626 163.367
R750 B.n626 B.n625 163.367
R751 B.n625 B.n92 163.367
R752 B.n621 B.n92 163.367
R753 B.n621 B.n620 163.367
R754 B.n620 B.n619 163.367
R755 B.n619 B.n94 163.367
R756 B.n615 B.n94 163.367
R757 B.n615 B.n614 163.367
R758 B.n614 B.n613 163.367
R759 B.n613 B.n96 163.367
R760 B.n609 B.n96 163.367
R761 B.n609 B.n608 163.367
R762 B.n608 B.n607 163.367
R763 B.n607 B.n98 163.367
R764 B.n603 B.n98 163.367
R765 B.n603 B.n602 163.367
R766 B.n602 B.n601 163.367
R767 B.n601 B.n100 163.367
R768 B.n597 B.n100 163.367
R769 B.n597 B.n596 163.367
R770 B.n596 B.n595 163.367
R771 B.n595 B.n102 163.367
R772 B.n591 B.n102 163.367
R773 B.n591 B.n590 163.367
R774 B.n590 B.n589 163.367
R775 B.n589 B.n104 163.367
R776 B.n585 B.n104 163.367
R777 B.n585 B.n584 163.367
R778 B.n584 B.n583 163.367
R779 B.n583 B.n106 163.367
R780 B.n579 B.n106 163.367
R781 B.n579 B.n578 163.367
R782 B.n578 B.n577 163.367
R783 B.n577 B.n108 163.367
R784 B.n573 B.n108 163.367
R785 B.n573 B.n572 163.367
R786 B.n572 B.n571 163.367
R787 B.n571 B.n110 163.367
R788 B.n567 B.n110 163.367
R789 B.n567 B.n566 163.367
R790 B.n566 B.n565 163.367
R791 B.n565 B.n112 163.367
R792 B.n561 B.n112 163.367
R793 B.n561 B.n560 163.367
R794 B.n560 B.n559 163.367
R795 B.n559 B.n114 163.367
R796 B.n555 B.n114 163.367
R797 B.n555 B.n554 163.367
R798 B.n554 B.n553 163.367
R799 B.n553 B.n116 163.367
R800 B.n549 B.n116 163.367
R801 B.n549 B.n548 163.367
R802 B.n548 B.n547 163.367
R803 B.n547 B.n118 163.367
R804 B.n543 B.n118 163.367
R805 B.n543 B.n542 163.367
R806 B.n542 B.n541 163.367
R807 B.n541 B.n120 163.367
R808 B.n537 B.n120 163.367
R809 B.n537 B.n536 163.367
R810 B.n536 B.n535 163.367
R811 B.n535 B.n122 163.367
R812 B.n531 B.n122 163.367
R813 B.n531 B.n530 163.367
R814 B.n530 B.n529 163.367
R815 B.n529 B.n124 163.367
R816 B.n525 B.n124 163.367
R817 B.n525 B.n524 163.367
R818 B.n524 B.n523 163.367
R819 B.n523 B.n126 163.367
R820 B.n519 B.n126 163.367
R821 B.n519 B.n518 163.367
R822 B.n518 B.n517 163.367
R823 B.n517 B.n128 163.367
R824 B.n513 B.n128 163.367
R825 B.n513 B.n512 163.367
R826 B.n512 B.n511 163.367
R827 B.n511 B.n130 163.367
R828 B.n507 B.n130 163.367
R829 B.n507 B.n506 163.367
R830 B.n506 B.n505 163.367
R831 B.n505 B.n132 163.367
R832 B.n501 B.n132 163.367
R833 B.n501 B.n500 163.367
R834 B.n500 B.n499 163.367
R835 B.n499 B.n134 163.367
R836 B.n495 B.n134 163.367
R837 B.n495 B.n494 163.367
R838 B.n494 B.n493 163.367
R839 B.n493 B.n136 163.367
R840 B.n489 B.n136 163.367
R841 B.n489 B.n488 163.367
R842 B.n488 B.n487 163.367
R843 B.n487 B.n138 163.367
R844 B.n483 B.n138 163.367
R845 B.n483 B.n482 163.367
R846 B.n482 B.n481 163.367
R847 B.n481 B.n140 163.367
R848 B.n806 B.n27 163.367
R849 B.n802 B.n27 163.367
R850 B.n802 B.n801 163.367
R851 B.n801 B.n800 163.367
R852 B.n800 B.n29 163.367
R853 B.n796 B.n29 163.367
R854 B.n796 B.n795 163.367
R855 B.n795 B.n794 163.367
R856 B.n794 B.n31 163.367
R857 B.n790 B.n31 163.367
R858 B.n790 B.n789 163.367
R859 B.n789 B.n788 163.367
R860 B.n788 B.n33 163.367
R861 B.n784 B.n33 163.367
R862 B.n784 B.n783 163.367
R863 B.n783 B.n782 163.367
R864 B.n782 B.n35 163.367
R865 B.n778 B.n35 163.367
R866 B.n778 B.n777 163.367
R867 B.n777 B.n776 163.367
R868 B.n776 B.n37 163.367
R869 B.n772 B.n37 163.367
R870 B.n772 B.n771 163.367
R871 B.n771 B.n770 163.367
R872 B.n770 B.n39 163.367
R873 B.n766 B.n39 163.367
R874 B.n766 B.n765 163.367
R875 B.n765 B.n764 163.367
R876 B.n764 B.n41 163.367
R877 B.n760 B.n41 163.367
R878 B.n760 B.n759 163.367
R879 B.n759 B.n758 163.367
R880 B.n758 B.n43 163.367
R881 B.n754 B.n43 163.367
R882 B.n754 B.n753 163.367
R883 B.n753 B.n752 163.367
R884 B.n752 B.n45 163.367
R885 B.n748 B.n45 163.367
R886 B.n748 B.n747 163.367
R887 B.n747 B.n746 163.367
R888 B.n746 B.n47 163.367
R889 B.n742 B.n47 163.367
R890 B.n742 B.n741 163.367
R891 B.n741 B.n740 163.367
R892 B.n740 B.n49 163.367
R893 B.n736 B.n49 163.367
R894 B.n736 B.n735 163.367
R895 B.n735 B.n734 163.367
R896 B.n734 B.n51 163.367
R897 B.n730 B.n51 163.367
R898 B.n730 B.n729 163.367
R899 B.n729 B.n728 163.367
R900 B.n728 B.n53 163.367
R901 B.n723 B.n53 163.367
R902 B.n723 B.n722 163.367
R903 B.n722 B.n721 163.367
R904 B.n721 B.n57 163.367
R905 B.n717 B.n57 163.367
R906 B.n717 B.n716 163.367
R907 B.n716 B.n715 163.367
R908 B.n715 B.n59 163.367
R909 B.n711 B.n59 163.367
R910 B.n711 B.n710 163.367
R911 B.n710 B.n709 163.367
R912 B.n709 B.n61 163.367
R913 B.n705 B.n61 163.367
R914 B.n705 B.n704 163.367
R915 B.n704 B.n703 163.367
R916 B.n703 B.n66 163.367
R917 B.n699 B.n66 163.367
R918 B.n699 B.n698 163.367
R919 B.n698 B.n697 163.367
R920 B.n697 B.n68 163.367
R921 B.n693 B.n68 163.367
R922 B.n693 B.n692 163.367
R923 B.n692 B.n691 163.367
R924 B.n691 B.n70 163.367
R925 B.n687 B.n70 163.367
R926 B.n687 B.n686 163.367
R927 B.n686 B.n685 163.367
R928 B.n685 B.n72 163.367
R929 B.n681 B.n72 163.367
R930 B.n681 B.n680 163.367
R931 B.n680 B.n679 163.367
R932 B.n679 B.n74 163.367
R933 B.n675 B.n74 163.367
R934 B.n675 B.n674 163.367
R935 B.n674 B.n673 163.367
R936 B.n673 B.n76 163.367
R937 B.n669 B.n76 163.367
R938 B.n669 B.n668 163.367
R939 B.n668 B.n667 163.367
R940 B.n667 B.n78 163.367
R941 B.n663 B.n78 163.367
R942 B.n663 B.n662 163.367
R943 B.n662 B.n661 163.367
R944 B.n661 B.n80 163.367
R945 B.n657 B.n80 163.367
R946 B.n657 B.n656 163.367
R947 B.n656 B.n655 163.367
R948 B.n655 B.n82 163.367
R949 B.n651 B.n82 163.367
R950 B.n651 B.n650 163.367
R951 B.n650 B.n649 163.367
R952 B.n649 B.n84 163.367
R953 B.n645 B.n84 163.367
R954 B.n645 B.n644 163.367
R955 B.n644 B.n643 163.367
R956 B.n643 B.n86 163.367
R957 B.n639 B.n86 163.367
R958 B.n639 B.n638 163.367
R959 B.n638 B.n637 163.367
R960 B.n637 B.n88 163.367
R961 B.n633 B.n88 163.367
R962 B.n633 B.n632 163.367
R963 B.n632 B.n631 163.367
R964 B.n631 B.n90 163.367
R965 B.n808 B.n807 163.367
R966 B.n808 B.n25 163.367
R967 B.n812 B.n25 163.367
R968 B.n813 B.n812 163.367
R969 B.n814 B.n813 163.367
R970 B.n814 B.n23 163.367
R971 B.n818 B.n23 163.367
R972 B.n819 B.n818 163.367
R973 B.n820 B.n819 163.367
R974 B.n820 B.n21 163.367
R975 B.n824 B.n21 163.367
R976 B.n825 B.n824 163.367
R977 B.n826 B.n825 163.367
R978 B.n826 B.n19 163.367
R979 B.n830 B.n19 163.367
R980 B.n831 B.n830 163.367
R981 B.n832 B.n831 163.367
R982 B.n832 B.n17 163.367
R983 B.n836 B.n17 163.367
R984 B.n837 B.n836 163.367
R985 B.n838 B.n837 163.367
R986 B.n838 B.n15 163.367
R987 B.n842 B.n15 163.367
R988 B.n843 B.n842 163.367
R989 B.n844 B.n843 163.367
R990 B.n844 B.n13 163.367
R991 B.n848 B.n13 163.367
R992 B.n849 B.n848 163.367
R993 B.n850 B.n849 163.367
R994 B.n850 B.n11 163.367
R995 B.n854 B.n11 163.367
R996 B.n855 B.n854 163.367
R997 B.n856 B.n855 163.367
R998 B.n856 B.n9 163.367
R999 B.n860 B.n9 163.367
R1000 B.n861 B.n860 163.367
R1001 B.n862 B.n861 163.367
R1002 B.n862 B.n7 163.367
R1003 B.n866 B.n7 163.367
R1004 B.n867 B.n866 163.367
R1005 B.n868 B.n867 163.367
R1006 B.n868 B.n5 163.367
R1007 B.n872 B.n5 163.367
R1008 B.n873 B.n872 163.367
R1009 B.n874 B.n873 163.367
R1010 B.n874 B.n3 163.367
R1011 B.n878 B.n3 163.367
R1012 B.n879 B.n878 163.367
R1013 B.n226 B.n2 163.367
R1014 B.n227 B.n226 163.367
R1015 B.n227 B.n224 163.367
R1016 B.n231 B.n224 163.367
R1017 B.n232 B.n231 163.367
R1018 B.n233 B.n232 163.367
R1019 B.n233 B.n222 163.367
R1020 B.n237 B.n222 163.367
R1021 B.n238 B.n237 163.367
R1022 B.n239 B.n238 163.367
R1023 B.n239 B.n220 163.367
R1024 B.n243 B.n220 163.367
R1025 B.n244 B.n243 163.367
R1026 B.n245 B.n244 163.367
R1027 B.n245 B.n218 163.367
R1028 B.n249 B.n218 163.367
R1029 B.n250 B.n249 163.367
R1030 B.n251 B.n250 163.367
R1031 B.n251 B.n216 163.367
R1032 B.n255 B.n216 163.367
R1033 B.n256 B.n255 163.367
R1034 B.n257 B.n256 163.367
R1035 B.n257 B.n214 163.367
R1036 B.n261 B.n214 163.367
R1037 B.n262 B.n261 163.367
R1038 B.n263 B.n262 163.367
R1039 B.n263 B.n212 163.367
R1040 B.n267 B.n212 163.367
R1041 B.n268 B.n267 163.367
R1042 B.n269 B.n268 163.367
R1043 B.n269 B.n210 163.367
R1044 B.n273 B.n210 163.367
R1045 B.n274 B.n273 163.367
R1046 B.n275 B.n274 163.367
R1047 B.n275 B.n208 163.367
R1048 B.n279 B.n208 163.367
R1049 B.n280 B.n279 163.367
R1050 B.n281 B.n280 163.367
R1051 B.n281 B.n206 163.367
R1052 B.n285 B.n206 163.367
R1053 B.n286 B.n285 163.367
R1054 B.n287 B.n286 163.367
R1055 B.n287 B.n204 163.367
R1056 B.n291 B.n204 163.367
R1057 B.n292 B.n291 163.367
R1058 B.n293 B.n292 163.367
R1059 B.n293 B.n202 163.367
R1060 B.n297 B.n202 163.367
R1061 B.n394 B.t11 106.966
R1062 B.n63 B.t1 106.966
R1063 B.n174 B.t5 106.945
R1064 B.n55 B.t7 106.945
R1065 B.n174 B.n173 68.0732
R1066 B.n394 B.n393 68.0732
R1067 B.n63 B.n62 68.0732
R1068 B.n55 B.n54 68.0732
R1069 B.n379 B.n174 59.5399
R1070 B.n395 B.n394 59.5399
R1071 B.n64 B.n63 59.5399
R1072 B.n725 B.n55 59.5399
R1073 B.n805 B.n26 33.5615
R1074 B.n629 B.n628 33.5615
R1075 B.n479 B.n478 33.5615
R1076 B.n296 B.n201 33.5615
R1077 B B.n881 18.0485
R1078 B.n809 B.n26 10.6151
R1079 B.n810 B.n809 10.6151
R1080 B.n811 B.n810 10.6151
R1081 B.n811 B.n24 10.6151
R1082 B.n815 B.n24 10.6151
R1083 B.n816 B.n815 10.6151
R1084 B.n817 B.n816 10.6151
R1085 B.n817 B.n22 10.6151
R1086 B.n821 B.n22 10.6151
R1087 B.n822 B.n821 10.6151
R1088 B.n823 B.n822 10.6151
R1089 B.n823 B.n20 10.6151
R1090 B.n827 B.n20 10.6151
R1091 B.n828 B.n827 10.6151
R1092 B.n829 B.n828 10.6151
R1093 B.n829 B.n18 10.6151
R1094 B.n833 B.n18 10.6151
R1095 B.n834 B.n833 10.6151
R1096 B.n835 B.n834 10.6151
R1097 B.n835 B.n16 10.6151
R1098 B.n839 B.n16 10.6151
R1099 B.n840 B.n839 10.6151
R1100 B.n841 B.n840 10.6151
R1101 B.n841 B.n14 10.6151
R1102 B.n845 B.n14 10.6151
R1103 B.n846 B.n845 10.6151
R1104 B.n847 B.n846 10.6151
R1105 B.n847 B.n12 10.6151
R1106 B.n851 B.n12 10.6151
R1107 B.n852 B.n851 10.6151
R1108 B.n853 B.n852 10.6151
R1109 B.n853 B.n10 10.6151
R1110 B.n857 B.n10 10.6151
R1111 B.n858 B.n857 10.6151
R1112 B.n859 B.n858 10.6151
R1113 B.n859 B.n8 10.6151
R1114 B.n863 B.n8 10.6151
R1115 B.n864 B.n863 10.6151
R1116 B.n865 B.n864 10.6151
R1117 B.n865 B.n6 10.6151
R1118 B.n869 B.n6 10.6151
R1119 B.n870 B.n869 10.6151
R1120 B.n871 B.n870 10.6151
R1121 B.n871 B.n4 10.6151
R1122 B.n875 B.n4 10.6151
R1123 B.n876 B.n875 10.6151
R1124 B.n877 B.n876 10.6151
R1125 B.n877 B.n0 10.6151
R1126 B.n805 B.n804 10.6151
R1127 B.n804 B.n803 10.6151
R1128 B.n803 B.n28 10.6151
R1129 B.n799 B.n28 10.6151
R1130 B.n799 B.n798 10.6151
R1131 B.n798 B.n797 10.6151
R1132 B.n797 B.n30 10.6151
R1133 B.n793 B.n30 10.6151
R1134 B.n793 B.n792 10.6151
R1135 B.n792 B.n791 10.6151
R1136 B.n791 B.n32 10.6151
R1137 B.n787 B.n32 10.6151
R1138 B.n787 B.n786 10.6151
R1139 B.n786 B.n785 10.6151
R1140 B.n785 B.n34 10.6151
R1141 B.n781 B.n34 10.6151
R1142 B.n781 B.n780 10.6151
R1143 B.n780 B.n779 10.6151
R1144 B.n779 B.n36 10.6151
R1145 B.n775 B.n36 10.6151
R1146 B.n775 B.n774 10.6151
R1147 B.n774 B.n773 10.6151
R1148 B.n773 B.n38 10.6151
R1149 B.n769 B.n38 10.6151
R1150 B.n769 B.n768 10.6151
R1151 B.n768 B.n767 10.6151
R1152 B.n767 B.n40 10.6151
R1153 B.n763 B.n40 10.6151
R1154 B.n763 B.n762 10.6151
R1155 B.n762 B.n761 10.6151
R1156 B.n761 B.n42 10.6151
R1157 B.n757 B.n42 10.6151
R1158 B.n757 B.n756 10.6151
R1159 B.n756 B.n755 10.6151
R1160 B.n755 B.n44 10.6151
R1161 B.n751 B.n44 10.6151
R1162 B.n751 B.n750 10.6151
R1163 B.n750 B.n749 10.6151
R1164 B.n749 B.n46 10.6151
R1165 B.n745 B.n46 10.6151
R1166 B.n745 B.n744 10.6151
R1167 B.n744 B.n743 10.6151
R1168 B.n743 B.n48 10.6151
R1169 B.n739 B.n48 10.6151
R1170 B.n739 B.n738 10.6151
R1171 B.n738 B.n737 10.6151
R1172 B.n737 B.n50 10.6151
R1173 B.n733 B.n50 10.6151
R1174 B.n733 B.n732 10.6151
R1175 B.n732 B.n731 10.6151
R1176 B.n731 B.n52 10.6151
R1177 B.n727 B.n52 10.6151
R1178 B.n727 B.n726 10.6151
R1179 B.n724 B.n56 10.6151
R1180 B.n720 B.n56 10.6151
R1181 B.n720 B.n719 10.6151
R1182 B.n719 B.n718 10.6151
R1183 B.n718 B.n58 10.6151
R1184 B.n714 B.n58 10.6151
R1185 B.n714 B.n713 10.6151
R1186 B.n713 B.n712 10.6151
R1187 B.n712 B.n60 10.6151
R1188 B.n708 B.n707 10.6151
R1189 B.n707 B.n706 10.6151
R1190 B.n706 B.n65 10.6151
R1191 B.n702 B.n65 10.6151
R1192 B.n702 B.n701 10.6151
R1193 B.n701 B.n700 10.6151
R1194 B.n700 B.n67 10.6151
R1195 B.n696 B.n67 10.6151
R1196 B.n696 B.n695 10.6151
R1197 B.n695 B.n694 10.6151
R1198 B.n694 B.n69 10.6151
R1199 B.n690 B.n69 10.6151
R1200 B.n690 B.n689 10.6151
R1201 B.n689 B.n688 10.6151
R1202 B.n688 B.n71 10.6151
R1203 B.n684 B.n71 10.6151
R1204 B.n684 B.n683 10.6151
R1205 B.n683 B.n682 10.6151
R1206 B.n682 B.n73 10.6151
R1207 B.n678 B.n73 10.6151
R1208 B.n678 B.n677 10.6151
R1209 B.n677 B.n676 10.6151
R1210 B.n676 B.n75 10.6151
R1211 B.n672 B.n75 10.6151
R1212 B.n672 B.n671 10.6151
R1213 B.n671 B.n670 10.6151
R1214 B.n670 B.n77 10.6151
R1215 B.n666 B.n77 10.6151
R1216 B.n666 B.n665 10.6151
R1217 B.n665 B.n664 10.6151
R1218 B.n664 B.n79 10.6151
R1219 B.n660 B.n79 10.6151
R1220 B.n660 B.n659 10.6151
R1221 B.n659 B.n658 10.6151
R1222 B.n658 B.n81 10.6151
R1223 B.n654 B.n81 10.6151
R1224 B.n654 B.n653 10.6151
R1225 B.n653 B.n652 10.6151
R1226 B.n652 B.n83 10.6151
R1227 B.n648 B.n83 10.6151
R1228 B.n648 B.n647 10.6151
R1229 B.n647 B.n646 10.6151
R1230 B.n646 B.n85 10.6151
R1231 B.n642 B.n85 10.6151
R1232 B.n642 B.n641 10.6151
R1233 B.n641 B.n640 10.6151
R1234 B.n640 B.n87 10.6151
R1235 B.n636 B.n87 10.6151
R1236 B.n636 B.n635 10.6151
R1237 B.n635 B.n634 10.6151
R1238 B.n634 B.n89 10.6151
R1239 B.n630 B.n89 10.6151
R1240 B.n630 B.n629 10.6151
R1241 B.n628 B.n91 10.6151
R1242 B.n624 B.n91 10.6151
R1243 B.n624 B.n623 10.6151
R1244 B.n623 B.n622 10.6151
R1245 B.n622 B.n93 10.6151
R1246 B.n618 B.n93 10.6151
R1247 B.n618 B.n617 10.6151
R1248 B.n617 B.n616 10.6151
R1249 B.n616 B.n95 10.6151
R1250 B.n612 B.n95 10.6151
R1251 B.n612 B.n611 10.6151
R1252 B.n611 B.n610 10.6151
R1253 B.n610 B.n97 10.6151
R1254 B.n606 B.n97 10.6151
R1255 B.n606 B.n605 10.6151
R1256 B.n605 B.n604 10.6151
R1257 B.n604 B.n99 10.6151
R1258 B.n600 B.n99 10.6151
R1259 B.n600 B.n599 10.6151
R1260 B.n599 B.n598 10.6151
R1261 B.n598 B.n101 10.6151
R1262 B.n594 B.n101 10.6151
R1263 B.n594 B.n593 10.6151
R1264 B.n593 B.n592 10.6151
R1265 B.n592 B.n103 10.6151
R1266 B.n588 B.n103 10.6151
R1267 B.n588 B.n587 10.6151
R1268 B.n587 B.n586 10.6151
R1269 B.n586 B.n105 10.6151
R1270 B.n582 B.n105 10.6151
R1271 B.n582 B.n581 10.6151
R1272 B.n581 B.n580 10.6151
R1273 B.n580 B.n107 10.6151
R1274 B.n576 B.n107 10.6151
R1275 B.n576 B.n575 10.6151
R1276 B.n575 B.n574 10.6151
R1277 B.n574 B.n109 10.6151
R1278 B.n570 B.n109 10.6151
R1279 B.n570 B.n569 10.6151
R1280 B.n569 B.n568 10.6151
R1281 B.n568 B.n111 10.6151
R1282 B.n564 B.n111 10.6151
R1283 B.n564 B.n563 10.6151
R1284 B.n563 B.n562 10.6151
R1285 B.n562 B.n113 10.6151
R1286 B.n558 B.n113 10.6151
R1287 B.n558 B.n557 10.6151
R1288 B.n557 B.n556 10.6151
R1289 B.n556 B.n115 10.6151
R1290 B.n552 B.n115 10.6151
R1291 B.n552 B.n551 10.6151
R1292 B.n551 B.n550 10.6151
R1293 B.n550 B.n117 10.6151
R1294 B.n546 B.n117 10.6151
R1295 B.n546 B.n545 10.6151
R1296 B.n545 B.n544 10.6151
R1297 B.n544 B.n119 10.6151
R1298 B.n540 B.n119 10.6151
R1299 B.n540 B.n539 10.6151
R1300 B.n539 B.n538 10.6151
R1301 B.n538 B.n121 10.6151
R1302 B.n534 B.n121 10.6151
R1303 B.n534 B.n533 10.6151
R1304 B.n533 B.n532 10.6151
R1305 B.n532 B.n123 10.6151
R1306 B.n528 B.n123 10.6151
R1307 B.n528 B.n527 10.6151
R1308 B.n527 B.n526 10.6151
R1309 B.n526 B.n125 10.6151
R1310 B.n522 B.n125 10.6151
R1311 B.n522 B.n521 10.6151
R1312 B.n521 B.n520 10.6151
R1313 B.n520 B.n127 10.6151
R1314 B.n516 B.n127 10.6151
R1315 B.n516 B.n515 10.6151
R1316 B.n515 B.n514 10.6151
R1317 B.n514 B.n129 10.6151
R1318 B.n510 B.n129 10.6151
R1319 B.n510 B.n509 10.6151
R1320 B.n509 B.n508 10.6151
R1321 B.n508 B.n131 10.6151
R1322 B.n504 B.n131 10.6151
R1323 B.n504 B.n503 10.6151
R1324 B.n503 B.n502 10.6151
R1325 B.n502 B.n133 10.6151
R1326 B.n498 B.n133 10.6151
R1327 B.n498 B.n497 10.6151
R1328 B.n497 B.n496 10.6151
R1329 B.n496 B.n135 10.6151
R1330 B.n492 B.n135 10.6151
R1331 B.n492 B.n491 10.6151
R1332 B.n491 B.n490 10.6151
R1333 B.n490 B.n137 10.6151
R1334 B.n486 B.n137 10.6151
R1335 B.n486 B.n485 10.6151
R1336 B.n485 B.n484 10.6151
R1337 B.n484 B.n139 10.6151
R1338 B.n480 B.n139 10.6151
R1339 B.n480 B.n479 10.6151
R1340 B.n225 B.n1 10.6151
R1341 B.n228 B.n225 10.6151
R1342 B.n229 B.n228 10.6151
R1343 B.n230 B.n229 10.6151
R1344 B.n230 B.n223 10.6151
R1345 B.n234 B.n223 10.6151
R1346 B.n235 B.n234 10.6151
R1347 B.n236 B.n235 10.6151
R1348 B.n236 B.n221 10.6151
R1349 B.n240 B.n221 10.6151
R1350 B.n241 B.n240 10.6151
R1351 B.n242 B.n241 10.6151
R1352 B.n242 B.n219 10.6151
R1353 B.n246 B.n219 10.6151
R1354 B.n247 B.n246 10.6151
R1355 B.n248 B.n247 10.6151
R1356 B.n248 B.n217 10.6151
R1357 B.n252 B.n217 10.6151
R1358 B.n253 B.n252 10.6151
R1359 B.n254 B.n253 10.6151
R1360 B.n254 B.n215 10.6151
R1361 B.n258 B.n215 10.6151
R1362 B.n259 B.n258 10.6151
R1363 B.n260 B.n259 10.6151
R1364 B.n260 B.n213 10.6151
R1365 B.n264 B.n213 10.6151
R1366 B.n265 B.n264 10.6151
R1367 B.n266 B.n265 10.6151
R1368 B.n266 B.n211 10.6151
R1369 B.n270 B.n211 10.6151
R1370 B.n271 B.n270 10.6151
R1371 B.n272 B.n271 10.6151
R1372 B.n272 B.n209 10.6151
R1373 B.n276 B.n209 10.6151
R1374 B.n277 B.n276 10.6151
R1375 B.n278 B.n277 10.6151
R1376 B.n278 B.n207 10.6151
R1377 B.n282 B.n207 10.6151
R1378 B.n283 B.n282 10.6151
R1379 B.n284 B.n283 10.6151
R1380 B.n284 B.n205 10.6151
R1381 B.n288 B.n205 10.6151
R1382 B.n289 B.n288 10.6151
R1383 B.n290 B.n289 10.6151
R1384 B.n290 B.n203 10.6151
R1385 B.n294 B.n203 10.6151
R1386 B.n295 B.n294 10.6151
R1387 B.n296 B.n295 10.6151
R1388 B.n300 B.n201 10.6151
R1389 B.n301 B.n300 10.6151
R1390 B.n302 B.n301 10.6151
R1391 B.n302 B.n199 10.6151
R1392 B.n306 B.n199 10.6151
R1393 B.n307 B.n306 10.6151
R1394 B.n308 B.n307 10.6151
R1395 B.n308 B.n197 10.6151
R1396 B.n312 B.n197 10.6151
R1397 B.n313 B.n312 10.6151
R1398 B.n314 B.n313 10.6151
R1399 B.n314 B.n195 10.6151
R1400 B.n318 B.n195 10.6151
R1401 B.n319 B.n318 10.6151
R1402 B.n320 B.n319 10.6151
R1403 B.n320 B.n193 10.6151
R1404 B.n324 B.n193 10.6151
R1405 B.n325 B.n324 10.6151
R1406 B.n326 B.n325 10.6151
R1407 B.n326 B.n191 10.6151
R1408 B.n330 B.n191 10.6151
R1409 B.n331 B.n330 10.6151
R1410 B.n332 B.n331 10.6151
R1411 B.n332 B.n189 10.6151
R1412 B.n336 B.n189 10.6151
R1413 B.n337 B.n336 10.6151
R1414 B.n338 B.n337 10.6151
R1415 B.n338 B.n187 10.6151
R1416 B.n342 B.n187 10.6151
R1417 B.n343 B.n342 10.6151
R1418 B.n344 B.n343 10.6151
R1419 B.n344 B.n185 10.6151
R1420 B.n348 B.n185 10.6151
R1421 B.n349 B.n348 10.6151
R1422 B.n350 B.n349 10.6151
R1423 B.n350 B.n183 10.6151
R1424 B.n354 B.n183 10.6151
R1425 B.n355 B.n354 10.6151
R1426 B.n356 B.n355 10.6151
R1427 B.n356 B.n181 10.6151
R1428 B.n360 B.n181 10.6151
R1429 B.n361 B.n360 10.6151
R1430 B.n362 B.n361 10.6151
R1431 B.n362 B.n179 10.6151
R1432 B.n366 B.n179 10.6151
R1433 B.n367 B.n366 10.6151
R1434 B.n368 B.n367 10.6151
R1435 B.n368 B.n177 10.6151
R1436 B.n372 B.n177 10.6151
R1437 B.n373 B.n372 10.6151
R1438 B.n374 B.n373 10.6151
R1439 B.n374 B.n175 10.6151
R1440 B.n378 B.n175 10.6151
R1441 B.n381 B.n380 10.6151
R1442 B.n381 B.n171 10.6151
R1443 B.n385 B.n171 10.6151
R1444 B.n386 B.n385 10.6151
R1445 B.n387 B.n386 10.6151
R1446 B.n387 B.n169 10.6151
R1447 B.n391 B.n169 10.6151
R1448 B.n392 B.n391 10.6151
R1449 B.n396 B.n392 10.6151
R1450 B.n400 B.n167 10.6151
R1451 B.n401 B.n400 10.6151
R1452 B.n402 B.n401 10.6151
R1453 B.n402 B.n165 10.6151
R1454 B.n406 B.n165 10.6151
R1455 B.n407 B.n406 10.6151
R1456 B.n408 B.n407 10.6151
R1457 B.n408 B.n163 10.6151
R1458 B.n412 B.n163 10.6151
R1459 B.n413 B.n412 10.6151
R1460 B.n414 B.n413 10.6151
R1461 B.n414 B.n161 10.6151
R1462 B.n418 B.n161 10.6151
R1463 B.n419 B.n418 10.6151
R1464 B.n420 B.n419 10.6151
R1465 B.n420 B.n159 10.6151
R1466 B.n424 B.n159 10.6151
R1467 B.n425 B.n424 10.6151
R1468 B.n426 B.n425 10.6151
R1469 B.n426 B.n157 10.6151
R1470 B.n430 B.n157 10.6151
R1471 B.n431 B.n430 10.6151
R1472 B.n432 B.n431 10.6151
R1473 B.n432 B.n155 10.6151
R1474 B.n436 B.n155 10.6151
R1475 B.n437 B.n436 10.6151
R1476 B.n438 B.n437 10.6151
R1477 B.n438 B.n153 10.6151
R1478 B.n442 B.n153 10.6151
R1479 B.n443 B.n442 10.6151
R1480 B.n444 B.n443 10.6151
R1481 B.n444 B.n151 10.6151
R1482 B.n448 B.n151 10.6151
R1483 B.n449 B.n448 10.6151
R1484 B.n450 B.n449 10.6151
R1485 B.n450 B.n149 10.6151
R1486 B.n454 B.n149 10.6151
R1487 B.n455 B.n454 10.6151
R1488 B.n456 B.n455 10.6151
R1489 B.n456 B.n147 10.6151
R1490 B.n460 B.n147 10.6151
R1491 B.n461 B.n460 10.6151
R1492 B.n462 B.n461 10.6151
R1493 B.n462 B.n145 10.6151
R1494 B.n466 B.n145 10.6151
R1495 B.n467 B.n466 10.6151
R1496 B.n468 B.n467 10.6151
R1497 B.n468 B.n143 10.6151
R1498 B.n472 B.n143 10.6151
R1499 B.n473 B.n472 10.6151
R1500 B.n474 B.n473 10.6151
R1501 B.n474 B.n141 10.6151
R1502 B.n478 B.n141 10.6151
R1503 B.n726 B.n725 9.36635
R1504 B.n708 B.n64 9.36635
R1505 B.n379 B.n378 9.36635
R1506 B.n395 B.n167 9.36635
R1507 B.n881 B.n0 8.11757
R1508 B.n881 B.n1 8.11757
R1509 B.n725 B.n724 1.24928
R1510 B.n64 B.n60 1.24928
R1511 B.n380 B.n379 1.24928
R1512 B.n396 B.n395 1.24928
C0 B VN 1.34061f
C1 VDD2 VP 0.50759f
C2 VTAIL VN 9.44892f
C3 w_n3778_n4238# VDD1 2.72786f
C4 B VDD1 2.59266f
C5 VTAIL VDD1 9.35747f
C6 VN VP 8.30016f
C7 VDD2 VN 9.35079f
C8 w_n3778_n4238# B 11.6969f
C9 w_n3778_n4238# VTAIL 3.61253f
C10 B VTAIL 4.92833f
C11 VDD1 VP 9.703321f
C12 VDD2 VDD1 1.63219f
C13 w_n3778_n4238# VP 7.88375f
C14 B VP 2.16173f
C15 w_n3778_n4238# VDD2 2.83146f
C16 B VDD2 2.68067f
C17 VDD1 VN 0.15133f
C18 VTAIL VP 9.46321f
C19 VDD2 VTAIL 9.411901f
C20 w_n3778_n4238# VN 7.39369f
C21 VDD2 VSUBS 2.18619f
C22 VDD1 VSUBS 2.72874f
C23 VTAIL VSUBS 1.461925f
C24 VN VSUBS 6.55481f
C25 VP VSUBS 3.54659f
C26 B VSUBS 5.578545f
C27 w_n3778_n4238# VSUBS 0.196078p
C28 B.n0 VSUBS 0.006814f
C29 B.n1 VSUBS 0.006814f
C30 B.n2 VSUBS 0.010078f
C31 B.n3 VSUBS 0.007723f
C32 B.n4 VSUBS 0.007723f
C33 B.n5 VSUBS 0.007723f
C34 B.n6 VSUBS 0.007723f
C35 B.n7 VSUBS 0.007723f
C36 B.n8 VSUBS 0.007723f
C37 B.n9 VSUBS 0.007723f
C38 B.n10 VSUBS 0.007723f
C39 B.n11 VSUBS 0.007723f
C40 B.n12 VSUBS 0.007723f
C41 B.n13 VSUBS 0.007723f
C42 B.n14 VSUBS 0.007723f
C43 B.n15 VSUBS 0.007723f
C44 B.n16 VSUBS 0.007723f
C45 B.n17 VSUBS 0.007723f
C46 B.n18 VSUBS 0.007723f
C47 B.n19 VSUBS 0.007723f
C48 B.n20 VSUBS 0.007723f
C49 B.n21 VSUBS 0.007723f
C50 B.n22 VSUBS 0.007723f
C51 B.n23 VSUBS 0.007723f
C52 B.n24 VSUBS 0.007723f
C53 B.n25 VSUBS 0.007723f
C54 B.n26 VSUBS 0.018193f
C55 B.n27 VSUBS 0.007723f
C56 B.n28 VSUBS 0.007723f
C57 B.n29 VSUBS 0.007723f
C58 B.n30 VSUBS 0.007723f
C59 B.n31 VSUBS 0.007723f
C60 B.n32 VSUBS 0.007723f
C61 B.n33 VSUBS 0.007723f
C62 B.n34 VSUBS 0.007723f
C63 B.n35 VSUBS 0.007723f
C64 B.n36 VSUBS 0.007723f
C65 B.n37 VSUBS 0.007723f
C66 B.n38 VSUBS 0.007723f
C67 B.n39 VSUBS 0.007723f
C68 B.n40 VSUBS 0.007723f
C69 B.n41 VSUBS 0.007723f
C70 B.n42 VSUBS 0.007723f
C71 B.n43 VSUBS 0.007723f
C72 B.n44 VSUBS 0.007723f
C73 B.n45 VSUBS 0.007723f
C74 B.n46 VSUBS 0.007723f
C75 B.n47 VSUBS 0.007723f
C76 B.n48 VSUBS 0.007723f
C77 B.n49 VSUBS 0.007723f
C78 B.n50 VSUBS 0.007723f
C79 B.n51 VSUBS 0.007723f
C80 B.n52 VSUBS 0.007723f
C81 B.n53 VSUBS 0.007723f
C82 B.t7 VSUBS 0.60465f
C83 B.t8 VSUBS 0.632327f
C84 B.t6 VSUBS 2.59808f
C85 B.n54 VSUBS 0.363984f
C86 B.n55 VSUBS 0.082175f
C87 B.n56 VSUBS 0.007723f
C88 B.n57 VSUBS 0.007723f
C89 B.n58 VSUBS 0.007723f
C90 B.n59 VSUBS 0.007723f
C91 B.n60 VSUBS 0.004316f
C92 B.n61 VSUBS 0.007723f
C93 B.t1 VSUBS 0.60463f
C94 B.t2 VSUBS 0.632312f
C95 B.t0 VSUBS 2.59808f
C96 B.n62 VSUBS 0.363999f
C97 B.n63 VSUBS 0.082195f
C98 B.n64 VSUBS 0.017893f
C99 B.n65 VSUBS 0.007723f
C100 B.n66 VSUBS 0.007723f
C101 B.n67 VSUBS 0.007723f
C102 B.n68 VSUBS 0.007723f
C103 B.n69 VSUBS 0.007723f
C104 B.n70 VSUBS 0.007723f
C105 B.n71 VSUBS 0.007723f
C106 B.n72 VSUBS 0.007723f
C107 B.n73 VSUBS 0.007723f
C108 B.n74 VSUBS 0.007723f
C109 B.n75 VSUBS 0.007723f
C110 B.n76 VSUBS 0.007723f
C111 B.n77 VSUBS 0.007723f
C112 B.n78 VSUBS 0.007723f
C113 B.n79 VSUBS 0.007723f
C114 B.n80 VSUBS 0.007723f
C115 B.n81 VSUBS 0.007723f
C116 B.n82 VSUBS 0.007723f
C117 B.n83 VSUBS 0.007723f
C118 B.n84 VSUBS 0.007723f
C119 B.n85 VSUBS 0.007723f
C120 B.n86 VSUBS 0.007723f
C121 B.n87 VSUBS 0.007723f
C122 B.n88 VSUBS 0.007723f
C123 B.n89 VSUBS 0.007723f
C124 B.n90 VSUBS 0.018604f
C125 B.n91 VSUBS 0.007723f
C126 B.n92 VSUBS 0.007723f
C127 B.n93 VSUBS 0.007723f
C128 B.n94 VSUBS 0.007723f
C129 B.n95 VSUBS 0.007723f
C130 B.n96 VSUBS 0.007723f
C131 B.n97 VSUBS 0.007723f
C132 B.n98 VSUBS 0.007723f
C133 B.n99 VSUBS 0.007723f
C134 B.n100 VSUBS 0.007723f
C135 B.n101 VSUBS 0.007723f
C136 B.n102 VSUBS 0.007723f
C137 B.n103 VSUBS 0.007723f
C138 B.n104 VSUBS 0.007723f
C139 B.n105 VSUBS 0.007723f
C140 B.n106 VSUBS 0.007723f
C141 B.n107 VSUBS 0.007723f
C142 B.n108 VSUBS 0.007723f
C143 B.n109 VSUBS 0.007723f
C144 B.n110 VSUBS 0.007723f
C145 B.n111 VSUBS 0.007723f
C146 B.n112 VSUBS 0.007723f
C147 B.n113 VSUBS 0.007723f
C148 B.n114 VSUBS 0.007723f
C149 B.n115 VSUBS 0.007723f
C150 B.n116 VSUBS 0.007723f
C151 B.n117 VSUBS 0.007723f
C152 B.n118 VSUBS 0.007723f
C153 B.n119 VSUBS 0.007723f
C154 B.n120 VSUBS 0.007723f
C155 B.n121 VSUBS 0.007723f
C156 B.n122 VSUBS 0.007723f
C157 B.n123 VSUBS 0.007723f
C158 B.n124 VSUBS 0.007723f
C159 B.n125 VSUBS 0.007723f
C160 B.n126 VSUBS 0.007723f
C161 B.n127 VSUBS 0.007723f
C162 B.n128 VSUBS 0.007723f
C163 B.n129 VSUBS 0.007723f
C164 B.n130 VSUBS 0.007723f
C165 B.n131 VSUBS 0.007723f
C166 B.n132 VSUBS 0.007723f
C167 B.n133 VSUBS 0.007723f
C168 B.n134 VSUBS 0.007723f
C169 B.n135 VSUBS 0.007723f
C170 B.n136 VSUBS 0.007723f
C171 B.n137 VSUBS 0.007723f
C172 B.n138 VSUBS 0.007723f
C173 B.n139 VSUBS 0.007723f
C174 B.n140 VSUBS 0.018193f
C175 B.n141 VSUBS 0.007723f
C176 B.n142 VSUBS 0.007723f
C177 B.n143 VSUBS 0.007723f
C178 B.n144 VSUBS 0.007723f
C179 B.n145 VSUBS 0.007723f
C180 B.n146 VSUBS 0.007723f
C181 B.n147 VSUBS 0.007723f
C182 B.n148 VSUBS 0.007723f
C183 B.n149 VSUBS 0.007723f
C184 B.n150 VSUBS 0.007723f
C185 B.n151 VSUBS 0.007723f
C186 B.n152 VSUBS 0.007723f
C187 B.n153 VSUBS 0.007723f
C188 B.n154 VSUBS 0.007723f
C189 B.n155 VSUBS 0.007723f
C190 B.n156 VSUBS 0.007723f
C191 B.n157 VSUBS 0.007723f
C192 B.n158 VSUBS 0.007723f
C193 B.n159 VSUBS 0.007723f
C194 B.n160 VSUBS 0.007723f
C195 B.n161 VSUBS 0.007723f
C196 B.n162 VSUBS 0.007723f
C197 B.n163 VSUBS 0.007723f
C198 B.n164 VSUBS 0.007723f
C199 B.n165 VSUBS 0.007723f
C200 B.n166 VSUBS 0.007723f
C201 B.n167 VSUBS 0.007269f
C202 B.n168 VSUBS 0.007723f
C203 B.n169 VSUBS 0.007723f
C204 B.n170 VSUBS 0.007723f
C205 B.n171 VSUBS 0.007723f
C206 B.n172 VSUBS 0.007723f
C207 B.t5 VSUBS 0.60465f
C208 B.t4 VSUBS 0.632327f
C209 B.t3 VSUBS 2.59808f
C210 B.n173 VSUBS 0.363984f
C211 B.n174 VSUBS 0.082175f
C212 B.n175 VSUBS 0.007723f
C213 B.n176 VSUBS 0.007723f
C214 B.n177 VSUBS 0.007723f
C215 B.n178 VSUBS 0.007723f
C216 B.n179 VSUBS 0.007723f
C217 B.n180 VSUBS 0.007723f
C218 B.n181 VSUBS 0.007723f
C219 B.n182 VSUBS 0.007723f
C220 B.n183 VSUBS 0.007723f
C221 B.n184 VSUBS 0.007723f
C222 B.n185 VSUBS 0.007723f
C223 B.n186 VSUBS 0.007723f
C224 B.n187 VSUBS 0.007723f
C225 B.n188 VSUBS 0.007723f
C226 B.n189 VSUBS 0.007723f
C227 B.n190 VSUBS 0.007723f
C228 B.n191 VSUBS 0.007723f
C229 B.n192 VSUBS 0.007723f
C230 B.n193 VSUBS 0.007723f
C231 B.n194 VSUBS 0.007723f
C232 B.n195 VSUBS 0.007723f
C233 B.n196 VSUBS 0.007723f
C234 B.n197 VSUBS 0.007723f
C235 B.n198 VSUBS 0.007723f
C236 B.n199 VSUBS 0.007723f
C237 B.n200 VSUBS 0.007723f
C238 B.n201 VSUBS 0.018604f
C239 B.n202 VSUBS 0.007723f
C240 B.n203 VSUBS 0.007723f
C241 B.n204 VSUBS 0.007723f
C242 B.n205 VSUBS 0.007723f
C243 B.n206 VSUBS 0.007723f
C244 B.n207 VSUBS 0.007723f
C245 B.n208 VSUBS 0.007723f
C246 B.n209 VSUBS 0.007723f
C247 B.n210 VSUBS 0.007723f
C248 B.n211 VSUBS 0.007723f
C249 B.n212 VSUBS 0.007723f
C250 B.n213 VSUBS 0.007723f
C251 B.n214 VSUBS 0.007723f
C252 B.n215 VSUBS 0.007723f
C253 B.n216 VSUBS 0.007723f
C254 B.n217 VSUBS 0.007723f
C255 B.n218 VSUBS 0.007723f
C256 B.n219 VSUBS 0.007723f
C257 B.n220 VSUBS 0.007723f
C258 B.n221 VSUBS 0.007723f
C259 B.n222 VSUBS 0.007723f
C260 B.n223 VSUBS 0.007723f
C261 B.n224 VSUBS 0.007723f
C262 B.n225 VSUBS 0.007723f
C263 B.n226 VSUBS 0.007723f
C264 B.n227 VSUBS 0.007723f
C265 B.n228 VSUBS 0.007723f
C266 B.n229 VSUBS 0.007723f
C267 B.n230 VSUBS 0.007723f
C268 B.n231 VSUBS 0.007723f
C269 B.n232 VSUBS 0.007723f
C270 B.n233 VSUBS 0.007723f
C271 B.n234 VSUBS 0.007723f
C272 B.n235 VSUBS 0.007723f
C273 B.n236 VSUBS 0.007723f
C274 B.n237 VSUBS 0.007723f
C275 B.n238 VSUBS 0.007723f
C276 B.n239 VSUBS 0.007723f
C277 B.n240 VSUBS 0.007723f
C278 B.n241 VSUBS 0.007723f
C279 B.n242 VSUBS 0.007723f
C280 B.n243 VSUBS 0.007723f
C281 B.n244 VSUBS 0.007723f
C282 B.n245 VSUBS 0.007723f
C283 B.n246 VSUBS 0.007723f
C284 B.n247 VSUBS 0.007723f
C285 B.n248 VSUBS 0.007723f
C286 B.n249 VSUBS 0.007723f
C287 B.n250 VSUBS 0.007723f
C288 B.n251 VSUBS 0.007723f
C289 B.n252 VSUBS 0.007723f
C290 B.n253 VSUBS 0.007723f
C291 B.n254 VSUBS 0.007723f
C292 B.n255 VSUBS 0.007723f
C293 B.n256 VSUBS 0.007723f
C294 B.n257 VSUBS 0.007723f
C295 B.n258 VSUBS 0.007723f
C296 B.n259 VSUBS 0.007723f
C297 B.n260 VSUBS 0.007723f
C298 B.n261 VSUBS 0.007723f
C299 B.n262 VSUBS 0.007723f
C300 B.n263 VSUBS 0.007723f
C301 B.n264 VSUBS 0.007723f
C302 B.n265 VSUBS 0.007723f
C303 B.n266 VSUBS 0.007723f
C304 B.n267 VSUBS 0.007723f
C305 B.n268 VSUBS 0.007723f
C306 B.n269 VSUBS 0.007723f
C307 B.n270 VSUBS 0.007723f
C308 B.n271 VSUBS 0.007723f
C309 B.n272 VSUBS 0.007723f
C310 B.n273 VSUBS 0.007723f
C311 B.n274 VSUBS 0.007723f
C312 B.n275 VSUBS 0.007723f
C313 B.n276 VSUBS 0.007723f
C314 B.n277 VSUBS 0.007723f
C315 B.n278 VSUBS 0.007723f
C316 B.n279 VSUBS 0.007723f
C317 B.n280 VSUBS 0.007723f
C318 B.n281 VSUBS 0.007723f
C319 B.n282 VSUBS 0.007723f
C320 B.n283 VSUBS 0.007723f
C321 B.n284 VSUBS 0.007723f
C322 B.n285 VSUBS 0.007723f
C323 B.n286 VSUBS 0.007723f
C324 B.n287 VSUBS 0.007723f
C325 B.n288 VSUBS 0.007723f
C326 B.n289 VSUBS 0.007723f
C327 B.n290 VSUBS 0.007723f
C328 B.n291 VSUBS 0.007723f
C329 B.n292 VSUBS 0.007723f
C330 B.n293 VSUBS 0.007723f
C331 B.n294 VSUBS 0.007723f
C332 B.n295 VSUBS 0.007723f
C333 B.n296 VSUBS 0.018193f
C334 B.n297 VSUBS 0.018193f
C335 B.n298 VSUBS 0.018604f
C336 B.n299 VSUBS 0.007723f
C337 B.n300 VSUBS 0.007723f
C338 B.n301 VSUBS 0.007723f
C339 B.n302 VSUBS 0.007723f
C340 B.n303 VSUBS 0.007723f
C341 B.n304 VSUBS 0.007723f
C342 B.n305 VSUBS 0.007723f
C343 B.n306 VSUBS 0.007723f
C344 B.n307 VSUBS 0.007723f
C345 B.n308 VSUBS 0.007723f
C346 B.n309 VSUBS 0.007723f
C347 B.n310 VSUBS 0.007723f
C348 B.n311 VSUBS 0.007723f
C349 B.n312 VSUBS 0.007723f
C350 B.n313 VSUBS 0.007723f
C351 B.n314 VSUBS 0.007723f
C352 B.n315 VSUBS 0.007723f
C353 B.n316 VSUBS 0.007723f
C354 B.n317 VSUBS 0.007723f
C355 B.n318 VSUBS 0.007723f
C356 B.n319 VSUBS 0.007723f
C357 B.n320 VSUBS 0.007723f
C358 B.n321 VSUBS 0.007723f
C359 B.n322 VSUBS 0.007723f
C360 B.n323 VSUBS 0.007723f
C361 B.n324 VSUBS 0.007723f
C362 B.n325 VSUBS 0.007723f
C363 B.n326 VSUBS 0.007723f
C364 B.n327 VSUBS 0.007723f
C365 B.n328 VSUBS 0.007723f
C366 B.n329 VSUBS 0.007723f
C367 B.n330 VSUBS 0.007723f
C368 B.n331 VSUBS 0.007723f
C369 B.n332 VSUBS 0.007723f
C370 B.n333 VSUBS 0.007723f
C371 B.n334 VSUBS 0.007723f
C372 B.n335 VSUBS 0.007723f
C373 B.n336 VSUBS 0.007723f
C374 B.n337 VSUBS 0.007723f
C375 B.n338 VSUBS 0.007723f
C376 B.n339 VSUBS 0.007723f
C377 B.n340 VSUBS 0.007723f
C378 B.n341 VSUBS 0.007723f
C379 B.n342 VSUBS 0.007723f
C380 B.n343 VSUBS 0.007723f
C381 B.n344 VSUBS 0.007723f
C382 B.n345 VSUBS 0.007723f
C383 B.n346 VSUBS 0.007723f
C384 B.n347 VSUBS 0.007723f
C385 B.n348 VSUBS 0.007723f
C386 B.n349 VSUBS 0.007723f
C387 B.n350 VSUBS 0.007723f
C388 B.n351 VSUBS 0.007723f
C389 B.n352 VSUBS 0.007723f
C390 B.n353 VSUBS 0.007723f
C391 B.n354 VSUBS 0.007723f
C392 B.n355 VSUBS 0.007723f
C393 B.n356 VSUBS 0.007723f
C394 B.n357 VSUBS 0.007723f
C395 B.n358 VSUBS 0.007723f
C396 B.n359 VSUBS 0.007723f
C397 B.n360 VSUBS 0.007723f
C398 B.n361 VSUBS 0.007723f
C399 B.n362 VSUBS 0.007723f
C400 B.n363 VSUBS 0.007723f
C401 B.n364 VSUBS 0.007723f
C402 B.n365 VSUBS 0.007723f
C403 B.n366 VSUBS 0.007723f
C404 B.n367 VSUBS 0.007723f
C405 B.n368 VSUBS 0.007723f
C406 B.n369 VSUBS 0.007723f
C407 B.n370 VSUBS 0.007723f
C408 B.n371 VSUBS 0.007723f
C409 B.n372 VSUBS 0.007723f
C410 B.n373 VSUBS 0.007723f
C411 B.n374 VSUBS 0.007723f
C412 B.n375 VSUBS 0.007723f
C413 B.n376 VSUBS 0.007723f
C414 B.n377 VSUBS 0.007723f
C415 B.n378 VSUBS 0.007269f
C416 B.n379 VSUBS 0.017893f
C417 B.n380 VSUBS 0.004316f
C418 B.n381 VSUBS 0.007723f
C419 B.n382 VSUBS 0.007723f
C420 B.n383 VSUBS 0.007723f
C421 B.n384 VSUBS 0.007723f
C422 B.n385 VSUBS 0.007723f
C423 B.n386 VSUBS 0.007723f
C424 B.n387 VSUBS 0.007723f
C425 B.n388 VSUBS 0.007723f
C426 B.n389 VSUBS 0.007723f
C427 B.n390 VSUBS 0.007723f
C428 B.n391 VSUBS 0.007723f
C429 B.n392 VSUBS 0.007723f
C430 B.t11 VSUBS 0.60463f
C431 B.t10 VSUBS 0.632312f
C432 B.t9 VSUBS 2.59808f
C433 B.n393 VSUBS 0.363999f
C434 B.n394 VSUBS 0.082195f
C435 B.n395 VSUBS 0.017893f
C436 B.n396 VSUBS 0.004316f
C437 B.n397 VSUBS 0.007723f
C438 B.n398 VSUBS 0.007723f
C439 B.n399 VSUBS 0.007723f
C440 B.n400 VSUBS 0.007723f
C441 B.n401 VSUBS 0.007723f
C442 B.n402 VSUBS 0.007723f
C443 B.n403 VSUBS 0.007723f
C444 B.n404 VSUBS 0.007723f
C445 B.n405 VSUBS 0.007723f
C446 B.n406 VSUBS 0.007723f
C447 B.n407 VSUBS 0.007723f
C448 B.n408 VSUBS 0.007723f
C449 B.n409 VSUBS 0.007723f
C450 B.n410 VSUBS 0.007723f
C451 B.n411 VSUBS 0.007723f
C452 B.n412 VSUBS 0.007723f
C453 B.n413 VSUBS 0.007723f
C454 B.n414 VSUBS 0.007723f
C455 B.n415 VSUBS 0.007723f
C456 B.n416 VSUBS 0.007723f
C457 B.n417 VSUBS 0.007723f
C458 B.n418 VSUBS 0.007723f
C459 B.n419 VSUBS 0.007723f
C460 B.n420 VSUBS 0.007723f
C461 B.n421 VSUBS 0.007723f
C462 B.n422 VSUBS 0.007723f
C463 B.n423 VSUBS 0.007723f
C464 B.n424 VSUBS 0.007723f
C465 B.n425 VSUBS 0.007723f
C466 B.n426 VSUBS 0.007723f
C467 B.n427 VSUBS 0.007723f
C468 B.n428 VSUBS 0.007723f
C469 B.n429 VSUBS 0.007723f
C470 B.n430 VSUBS 0.007723f
C471 B.n431 VSUBS 0.007723f
C472 B.n432 VSUBS 0.007723f
C473 B.n433 VSUBS 0.007723f
C474 B.n434 VSUBS 0.007723f
C475 B.n435 VSUBS 0.007723f
C476 B.n436 VSUBS 0.007723f
C477 B.n437 VSUBS 0.007723f
C478 B.n438 VSUBS 0.007723f
C479 B.n439 VSUBS 0.007723f
C480 B.n440 VSUBS 0.007723f
C481 B.n441 VSUBS 0.007723f
C482 B.n442 VSUBS 0.007723f
C483 B.n443 VSUBS 0.007723f
C484 B.n444 VSUBS 0.007723f
C485 B.n445 VSUBS 0.007723f
C486 B.n446 VSUBS 0.007723f
C487 B.n447 VSUBS 0.007723f
C488 B.n448 VSUBS 0.007723f
C489 B.n449 VSUBS 0.007723f
C490 B.n450 VSUBS 0.007723f
C491 B.n451 VSUBS 0.007723f
C492 B.n452 VSUBS 0.007723f
C493 B.n453 VSUBS 0.007723f
C494 B.n454 VSUBS 0.007723f
C495 B.n455 VSUBS 0.007723f
C496 B.n456 VSUBS 0.007723f
C497 B.n457 VSUBS 0.007723f
C498 B.n458 VSUBS 0.007723f
C499 B.n459 VSUBS 0.007723f
C500 B.n460 VSUBS 0.007723f
C501 B.n461 VSUBS 0.007723f
C502 B.n462 VSUBS 0.007723f
C503 B.n463 VSUBS 0.007723f
C504 B.n464 VSUBS 0.007723f
C505 B.n465 VSUBS 0.007723f
C506 B.n466 VSUBS 0.007723f
C507 B.n467 VSUBS 0.007723f
C508 B.n468 VSUBS 0.007723f
C509 B.n469 VSUBS 0.007723f
C510 B.n470 VSUBS 0.007723f
C511 B.n471 VSUBS 0.007723f
C512 B.n472 VSUBS 0.007723f
C513 B.n473 VSUBS 0.007723f
C514 B.n474 VSUBS 0.007723f
C515 B.n475 VSUBS 0.007723f
C516 B.n476 VSUBS 0.007723f
C517 B.n477 VSUBS 0.018604f
C518 B.n478 VSUBS 0.017716f
C519 B.n479 VSUBS 0.019081f
C520 B.n480 VSUBS 0.007723f
C521 B.n481 VSUBS 0.007723f
C522 B.n482 VSUBS 0.007723f
C523 B.n483 VSUBS 0.007723f
C524 B.n484 VSUBS 0.007723f
C525 B.n485 VSUBS 0.007723f
C526 B.n486 VSUBS 0.007723f
C527 B.n487 VSUBS 0.007723f
C528 B.n488 VSUBS 0.007723f
C529 B.n489 VSUBS 0.007723f
C530 B.n490 VSUBS 0.007723f
C531 B.n491 VSUBS 0.007723f
C532 B.n492 VSUBS 0.007723f
C533 B.n493 VSUBS 0.007723f
C534 B.n494 VSUBS 0.007723f
C535 B.n495 VSUBS 0.007723f
C536 B.n496 VSUBS 0.007723f
C537 B.n497 VSUBS 0.007723f
C538 B.n498 VSUBS 0.007723f
C539 B.n499 VSUBS 0.007723f
C540 B.n500 VSUBS 0.007723f
C541 B.n501 VSUBS 0.007723f
C542 B.n502 VSUBS 0.007723f
C543 B.n503 VSUBS 0.007723f
C544 B.n504 VSUBS 0.007723f
C545 B.n505 VSUBS 0.007723f
C546 B.n506 VSUBS 0.007723f
C547 B.n507 VSUBS 0.007723f
C548 B.n508 VSUBS 0.007723f
C549 B.n509 VSUBS 0.007723f
C550 B.n510 VSUBS 0.007723f
C551 B.n511 VSUBS 0.007723f
C552 B.n512 VSUBS 0.007723f
C553 B.n513 VSUBS 0.007723f
C554 B.n514 VSUBS 0.007723f
C555 B.n515 VSUBS 0.007723f
C556 B.n516 VSUBS 0.007723f
C557 B.n517 VSUBS 0.007723f
C558 B.n518 VSUBS 0.007723f
C559 B.n519 VSUBS 0.007723f
C560 B.n520 VSUBS 0.007723f
C561 B.n521 VSUBS 0.007723f
C562 B.n522 VSUBS 0.007723f
C563 B.n523 VSUBS 0.007723f
C564 B.n524 VSUBS 0.007723f
C565 B.n525 VSUBS 0.007723f
C566 B.n526 VSUBS 0.007723f
C567 B.n527 VSUBS 0.007723f
C568 B.n528 VSUBS 0.007723f
C569 B.n529 VSUBS 0.007723f
C570 B.n530 VSUBS 0.007723f
C571 B.n531 VSUBS 0.007723f
C572 B.n532 VSUBS 0.007723f
C573 B.n533 VSUBS 0.007723f
C574 B.n534 VSUBS 0.007723f
C575 B.n535 VSUBS 0.007723f
C576 B.n536 VSUBS 0.007723f
C577 B.n537 VSUBS 0.007723f
C578 B.n538 VSUBS 0.007723f
C579 B.n539 VSUBS 0.007723f
C580 B.n540 VSUBS 0.007723f
C581 B.n541 VSUBS 0.007723f
C582 B.n542 VSUBS 0.007723f
C583 B.n543 VSUBS 0.007723f
C584 B.n544 VSUBS 0.007723f
C585 B.n545 VSUBS 0.007723f
C586 B.n546 VSUBS 0.007723f
C587 B.n547 VSUBS 0.007723f
C588 B.n548 VSUBS 0.007723f
C589 B.n549 VSUBS 0.007723f
C590 B.n550 VSUBS 0.007723f
C591 B.n551 VSUBS 0.007723f
C592 B.n552 VSUBS 0.007723f
C593 B.n553 VSUBS 0.007723f
C594 B.n554 VSUBS 0.007723f
C595 B.n555 VSUBS 0.007723f
C596 B.n556 VSUBS 0.007723f
C597 B.n557 VSUBS 0.007723f
C598 B.n558 VSUBS 0.007723f
C599 B.n559 VSUBS 0.007723f
C600 B.n560 VSUBS 0.007723f
C601 B.n561 VSUBS 0.007723f
C602 B.n562 VSUBS 0.007723f
C603 B.n563 VSUBS 0.007723f
C604 B.n564 VSUBS 0.007723f
C605 B.n565 VSUBS 0.007723f
C606 B.n566 VSUBS 0.007723f
C607 B.n567 VSUBS 0.007723f
C608 B.n568 VSUBS 0.007723f
C609 B.n569 VSUBS 0.007723f
C610 B.n570 VSUBS 0.007723f
C611 B.n571 VSUBS 0.007723f
C612 B.n572 VSUBS 0.007723f
C613 B.n573 VSUBS 0.007723f
C614 B.n574 VSUBS 0.007723f
C615 B.n575 VSUBS 0.007723f
C616 B.n576 VSUBS 0.007723f
C617 B.n577 VSUBS 0.007723f
C618 B.n578 VSUBS 0.007723f
C619 B.n579 VSUBS 0.007723f
C620 B.n580 VSUBS 0.007723f
C621 B.n581 VSUBS 0.007723f
C622 B.n582 VSUBS 0.007723f
C623 B.n583 VSUBS 0.007723f
C624 B.n584 VSUBS 0.007723f
C625 B.n585 VSUBS 0.007723f
C626 B.n586 VSUBS 0.007723f
C627 B.n587 VSUBS 0.007723f
C628 B.n588 VSUBS 0.007723f
C629 B.n589 VSUBS 0.007723f
C630 B.n590 VSUBS 0.007723f
C631 B.n591 VSUBS 0.007723f
C632 B.n592 VSUBS 0.007723f
C633 B.n593 VSUBS 0.007723f
C634 B.n594 VSUBS 0.007723f
C635 B.n595 VSUBS 0.007723f
C636 B.n596 VSUBS 0.007723f
C637 B.n597 VSUBS 0.007723f
C638 B.n598 VSUBS 0.007723f
C639 B.n599 VSUBS 0.007723f
C640 B.n600 VSUBS 0.007723f
C641 B.n601 VSUBS 0.007723f
C642 B.n602 VSUBS 0.007723f
C643 B.n603 VSUBS 0.007723f
C644 B.n604 VSUBS 0.007723f
C645 B.n605 VSUBS 0.007723f
C646 B.n606 VSUBS 0.007723f
C647 B.n607 VSUBS 0.007723f
C648 B.n608 VSUBS 0.007723f
C649 B.n609 VSUBS 0.007723f
C650 B.n610 VSUBS 0.007723f
C651 B.n611 VSUBS 0.007723f
C652 B.n612 VSUBS 0.007723f
C653 B.n613 VSUBS 0.007723f
C654 B.n614 VSUBS 0.007723f
C655 B.n615 VSUBS 0.007723f
C656 B.n616 VSUBS 0.007723f
C657 B.n617 VSUBS 0.007723f
C658 B.n618 VSUBS 0.007723f
C659 B.n619 VSUBS 0.007723f
C660 B.n620 VSUBS 0.007723f
C661 B.n621 VSUBS 0.007723f
C662 B.n622 VSUBS 0.007723f
C663 B.n623 VSUBS 0.007723f
C664 B.n624 VSUBS 0.007723f
C665 B.n625 VSUBS 0.007723f
C666 B.n626 VSUBS 0.007723f
C667 B.n627 VSUBS 0.018193f
C668 B.n628 VSUBS 0.018193f
C669 B.n629 VSUBS 0.018604f
C670 B.n630 VSUBS 0.007723f
C671 B.n631 VSUBS 0.007723f
C672 B.n632 VSUBS 0.007723f
C673 B.n633 VSUBS 0.007723f
C674 B.n634 VSUBS 0.007723f
C675 B.n635 VSUBS 0.007723f
C676 B.n636 VSUBS 0.007723f
C677 B.n637 VSUBS 0.007723f
C678 B.n638 VSUBS 0.007723f
C679 B.n639 VSUBS 0.007723f
C680 B.n640 VSUBS 0.007723f
C681 B.n641 VSUBS 0.007723f
C682 B.n642 VSUBS 0.007723f
C683 B.n643 VSUBS 0.007723f
C684 B.n644 VSUBS 0.007723f
C685 B.n645 VSUBS 0.007723f
C686 B.n646 VSUBS 0.007723f
C687 B.n647 VSUBS 0.007723f
C688 B.n648 VSUBS 0.007723f
C689 B.n649 VSUBS 0.007723f
C690 B.n650 VSUBS 0.007723f
C691 B.n651 VSUBS 0.007723f
C692 B.n652 VSUBS 0.007723f
C693 B.n653 VSUBS 0.007723f
C694 B.n654 VSUBS 0.007723f
C695 B.n655 VSUBS 0.007723f
C696 B.n656 VSUBS 0.007723f
C697 B.n657 VSUBS 0.007723f
C698 B.n658 VSUBS 0.007723f
C699 B.n659 VSUBS 0.007723f
C700 B.n660 VSUBS 0.007723f
C701 B.n661 VSUBS 0.007723f
C702 B.n662 VSUBS 0.007723f
C703 B.n663 VSUBS 0.007723f
C704 B.n664 VSUBS 0.007723f
C705 B.n665 VSUBS 0.007723f
C706 B.n666 VSUBS 0.007723f
C707 B.n667 VSUBS 0.007723f
C708 B.n668 VSUBS 0.007723f
C709 B.n669 VSUBS 0.007723f
C710 B.n670 VSUBS 0.007723f
C711 B.n671 VSUBS 0.007723f
C712 B.n672 VSUBS 0.007723f
C713 B.n673 VSUBS 0.007723f
C714 B.n674 VSUBS 0.007723f
C715 B.n675 VSUBS 0.007723f
C716 B.n676 VSUBS 0.007723f
C717 B.n677 VSUBS 0.007723f
C718 B.n678 VSUBS 0.007723f
C719 B.n679 VSUBS 0.007723f
C720 B.n680 VSUBS 0.007723f
C721 B.n681 VSUBS 0.007723f
C722 B.n682 VSUBS 0.007723f
C723 B.n683 VSUBS 0.007723f
C724 B.n684 VSUBS 0.007723f
C725 B.n685 VSUBS 0.007723f
C726 B.n686 VSUBS 0.007723f
C727 B.n687 VSUBS 0.007723f
C728 B.n688 VSUBS 0.007723f
C729 B.n689 VSUBS 0.007723f
C730 B.n690 VSUBS 0.007723f
C731 B.n691 VSUBS 0.007723f
C732 B.n692 VSUBS 0.007723f
C733 B.n693 VSUBS 0.007723f
C734 B.n694 VSUBS 0.007723f
C735 B.n695 VSUBS 0.007723f
C736 B.n696 VSUBS 0.007723f
C737 B.n697 VSUBS 0.007723f
C738 B.n698 VSUBS 0.007723f
C739 B.n699 VSUBS 0.007723f
C740 B.n700 VSUBS 0.007723f
C741 B.n701 VSUBS 0.007723f
C742 B.n702 VSUBS 0.007723f
C743 B.n703 VSUBS 0.007723f
C744 B.n704 VSUBS 0.007723f
C745 B.n705 VSUBS 0.007723f
C746 B.n706 VSUBS 0.007723f
C747 B.n707 VSUBS 0.007723f
C748 B.n708 VSUBS 0.007269f
C749 B.n709 VSUBS 0.007723f
C750 B.n710 VSUBS 0.007723f
C751 B.n711 VSUBS 0.007723f
C752 B.n712 VSUBS 0.007723f
C753 B.n713 VSUBS 0.007723f
C754 B.n714 VSUBS 0.007723f
C755 B.n715 VSUBS 0.007723f
C756 B.n716 VSUBS 0.007723f
C757 B.n717 VSUBS 0.007723f
C758 B.n718 VSUBS 0.007723f
C759 B.n719 VSUBS 0.007723f
C760 B.n720 VSUBS 0.007723f
C761 B.n721 VSUBS 0.007723f
C762 B.n722 VSUBS 0.007723f
C763 B.n723 VSUBS 0.007723f
C764 B.n724 VSUBS 0.004316f
C765 B.n725 VSUBS 0.017893f
C766 B.n726 VSUBS 0.007269f
C767 B.n727 VSUBS 0.007723f
C768 B.n728 VSUBS 0.007723f
C769 B.n729 VSUBS 0.007723f
C770 B.n730 VSUBS 0.007723f
C771 B.n731 VSUBS 0.007723f
C772 B.n732 VSUBS 0.007723f
C773 B.n733 VSUBS 0.007723f
C774 B.n734 VSUBS 0.007723f
C775 B.n735 VSUBS 0.007723f
C776 B.n736 VSUBS 0.007723f
C777 B.n737 VSUBS 0.007723f
C778 B.n738 VSUBS 0.007723f
C779 B.n739 VSUBS 0.007723f
C780 B.n740 VSUBS 0.007723f
C781 B.n741 VSUBS 0.007723f
C782 B.n742 VSUBS 0.007723f
C783 B.n743 VSUBS 0.007723f
C784 B.n744 VSUBS 0.007723f
C785 B.n745 VSUBS 0.007723f
C786 B.n746 VSUBS 0.007723f
C787 B.n747 VSUBS 0.007723f
C788 B.n748 VSUBS 0.007723f
C789 B.n749 VSUBS 0.007723f
C790 B.n750 VSUBS 0.007723f
C791 B.n751 VSUBS 0.007723f
C792 B.n752 VSUBS 0.007723f
C793 B.n753 VSUBS 0.007723f
C794 B.n754 VSUBS 0.007723f
C795 B.n755 VSUBS 0.007723f
C796 B.n756 VSUBS 0.007723f
C797 B.n757 VSUBS 0.007723f
C798 B.n758 VSUBS 0.007723f
C799 B.n759 VSUBS 0.007723f
C800 B.n760 VSUBS 0.007723f
C801 B.n761 VSUBS 0.007723f
C802 B.n762 VSUBS 0.007723f
C803 B.n763 VSUBS 0.007723f
C804 B.n764 VSUBS 0.007723f
C805 B.n765 VSUBS 0.007723f
C806 B.n766 VSUBS 0.007723f
C807 B.n767 VSUBS 0.007723f
C808 B.n768 VSUBS 0.007723f
C809 B.n769 VSUBS 0.007723f
C810 B.n770 VSUBS 0.007723f
C811 B.n771 VSUBS 0.007723f
C812 B.n772 VSUBS 0.007723f
C813 B.n773 VSUBS 0.007723f
C814 B.n774 VSUBS 0.007723f
C815 B.n775 VSUBS 0.007723f
C816 B.n776 VSUBS 0.007723f
C817 B.n777 VSUBS 0.007723f
C818 B.n778 VSUBS 0.007723f
C819 B.n779 VSUBS 0.007723f
C820 B.n780 VSUBS 0.007723f
C821 B.n781 VSUBS 0.007723f
C822 B.n782 VSUBS 0.007723f
C823 B.n783 VSUBS 0.007723f
C824 B.n784 VSUBS 0.007723f
C825 B.n785 VSUBS 0.007723f
C826 B.n786 VSUBS 0.007723f
C827 B.n787 VSUBS 0.007723f
C828 B.n788 VSUBS 0.007723f
C829 B.n789 VSUBS 0.007723f
C830 B.n790 VSUBS 0.007723f
C831 B.n791 VSUBS 0.007723f
C832 B.n792 VSUBS 0.007723f
C833 B.n793 VSUBS 0.007723f
C834 B.n794 VSUBS 0.007723f
C835 B.n795 VSUBS 0.007723f
C836 B.n796 VSUBS 0.007723f
C837 B.n797 VSUBS 0.007723f
C838 B.n798 VSUBS 0.007723f
C839 B.n799 VSUBS 0.007723f
C840 B.n800 VSUBS 0.007723f
C841 B.n801 VSUBS 0.007723f
C842 B.n802 VSUBS 0.007723f
C843 B.n803 VSUBS 0.007723f
C844 B.n804 VSUBS 0.007723f
C845 B.n805 VSUBS 0.018604f
C846 B.n806 VSUBS 0.018604f
C847 B.n807 VSUBS 0.018193f
C848 B.n808 VSUBS 0.007723f
C849 B.n809 VSUBS 0.007723f
C850 B.n810 VSUBS 0.007723f
C851 B.n811 VSUBS 0.007723f
C852 B.n812 VSUBS 0.007723f
C853 B.n813 VSUBS 0.007723f
C854 B.n814 VSUBS 0.007723f
C855 B.n815 VSUBS 0.007723f
C856 B.n816 VSUBS 0.007723f
C857 B.n817 VSUBS 0.007723f
C858 B.n818 VSUBS 0.007723f
C859 B.n819 VSUBS 0.007723f
C860 B.n820 VSUBS 0.007723f
C861 B.n821 VSUBS 0.007723f
C862 B.n822 VSUBS 0.007723f
C863 B.n823 VSUBS 0.007723f
C864 B.n824 VSUBS 0.007723f
C865 B.n825 VSUBS 0.007723f
C866 B.n826 VSUBS 0.007723f
C867 B.n827 VSUBS 0.007723f
C868 B.n828 VSUBS 0.007723f
C869 B.n829 VSUBS 0.007723f
C870 B.n830 VSUBS 0.007723f
C871 B.n831 VSUBS 0.007723f
C872 B.n832 VSUBS 0.007723f
C873 B.n833 VSUBS 0.007723f
C874 B.n834 VSUBS 0.007723f
C875 B.n835 VSUBS 0.007723f
C876 B.n836 VSUBS 0.007723f
C877 B.n837 VSUBS 0.007723f
C878 B.n838 VSUBS 0.007723f
C879 B.n839 VSUBS 0.007723f
C880 B.n840 VSUBS 0.007723f
C881 B.n841 VSUBS 0.007723f
C882 B.n842 VSUBS 0.007723f
C883 B.n843 VSUBS 0.007723f
C884 B.n844 VSUBS 0.007723f
C885 B.n845 VSUBS 0.007723f
C886 B.n846 VSUBS 0.007723f
C887 B.n847 VSUBS 0.007723f
C888 B.n848 VSUBS 0.007723f
C889 B.n849 VSUBS 0.007723f
C890 B.n850 VSUBS 0.007723f
C891 B.n851 VSUBS 0.007723f
C892 B.n852 VSUBS 0.007723f
C893 B.n853 VSUBS 0.007723f
C894 B.n854 VSUBS 0.007723f
C895 B.n855 VSUBS 0.007723f
C896 B.n856 VSUBS 0.007723f
C897 B.n857 VSUBS 0.007723f
C898 B.n858 VSUBS 0.007723f
C899 B.n859 VSUBS 0.007723f
C900 B.n860 VSUBS 0.007723f
C901 B.n861 VSUBS 0.007723f
C902 B.n862 VSUBS 0.007723f
C903 B.n863 VSUBS 0.007723f
C904 B.n864 VSUBS 0.007723f
C905 B.n865 VSUBS 0.007723f
C906 B.n866 VSUBS 0.007723f
C907 B.n867 VSUBS 0.007723f
C908 B.n868 VSUBS 0.007723f
C909 B.n869 VSUBS 0.007723f
C910 B.n870 VSUBS 0.007723f
C911 B.n871 VSUBS 0.007723f
C912 B.n872 VSUBS 0.007723f
C913 B.n873 VSUBS 0.007723f
C914 B.n874 VSUBS 0.007723f
C915 B.n875 VSUBS 0.007723f
C916 B.n876 VSUBS 0.007723f
C917 B.n877 VSUBS 0.007723f
C918 B.n878 VSUBS 0.007723f
C919 B.n879 VSUBS 0.010078f
C920 B.n880 VSUBS 0.010736f
C921 B.n881 VSUBS 0.021349f
C922 VDD2.t4 VSUBS 3.79314f
C923 VDD2.t0 VSUBS 0.35449f
C924 VDD2.t3 VSUBS 0.35449f
C925 VDD2.n0 VSUBS 2.90927f
C926 VDD2.n1 VSUBS 4.41143f
C927 VDD2.t5 VSUBS 3.76703f
C928 VDD2.n2 VSUBS 3.95054f
C929 VDD2.t1 VSUBS 0.35449f
C930 VDD2.t2 VSUBS 0.35449f
C931 VDD2.n3 VSUBS 2.90922f
C932 VN.t2 VSUBS 3.56243f
C933 VN.n0 VSUBS 1.32717f
C934 VN.n1 VSUBS 0.024958f
C935 VN.n2 VSUBS 0.020185f
C936 VN.n3 VSUBS 0.024958f
C937 VN.t5 VSUBS 3.56243f
C938 VN.n4 VSUBS 1.31705f
C939 VN.t1 VSUBS 3.85649f
C940 VN.n5 VSUBS 1.26621f
C941 VN.n6 VSUBS 0.290329f
C942 VN.n7 VSUBS 0.035033f
C943 VN.n8 VSUBS 0.046515f
C944 VN.n9 VSUBS 0.049726f
C945 VN.n10 VSUBS 0.024958f
C946 VN.n11 VSUBS 0.024958f
C947 VN.n12 VSUBS 0.024958f
C948 VN.n13 VSUBS 0.049476f
C949 VN.n14 VSUBS 0.046515f
C950 VN.n15 VSUBS 0.035492f
C951 VN.n16 VSUBS 0.040281f
C952 VN.n17 VSUBS 0.060971f
C953 VN.t0 VSUBS 3.56243f
C954 VN.n18 VSUBS 1.32717f
C955 VN.n19 VSUBS 0.024958f
C956 VN.n20 VSUBS 0.020185f
C957 VN.n21 VSUBS 0.024958f
C958 VN.t4 VSUBS 3.56243f
C959 VN.n22 VSUBS 1.31705f
C960 VN.t3 VSUBS 3.85649f
C961 VN.n23 VSUBS 1.26621f
C962 VN.n24 VSUBS 0.290329f
C963 VN.n25 VSUBS 0.035033f
C964 VN.n26 VSUBS 0.046515f
C965 VN.n27 VSUBS 0.049726f
C966 VN.n28 VSUBS 0.024958f
C967 VN.n29 VSUBS 0.024958f
C968 VN.n30 VSUBS 0.024958f
C969 VN.n31 VSUBS 0.049476f
C970 VN.n32 VSUBS 0.046515f
C971 VN.n33 VSUBS 0.035492f
C972 VN.n34 VSUBS 0.040281f
C973 VN.n35 VSUBS 1.60401f
C974 VTAIL.t4 VSUBS 0.365007f
C975 VTAIL.t1 VSUBS 0.365007f
C976 VTAIL.n0 VSUBS 2.80591f
C977 VTAIL.n1 VSUBS 0.955322f
C978 VTAIL.t7 VSUBS 3.67285f
C979 VTAIL.n2 VSUBS 1.28513f
C980 VTAIL.t10 VSUBS 0.365007f
C981 VTAIL.t9 VSUBS 0.365007f
C982 VTAIL.n3 VSUBS 2.80591f
C983 VTAIL.n4 VSUBS 3.19381f
C984 VTAIL.t3 VSUBS 0.365007f
C985 VTAIL.t2 VSUBS 0.365007f
C986 VTAIL.n5 VSUBS 2.80591f
C987 VTAIL.n6 VSUBS 3.19381f
C988 VTAIL.t5 VSUBS 3.67286f
C989 VTAIL.n7 VSUBS 1.28513f
C990 VTAIL.t8 VSUBS 0.365007f
C991 VTAIL.t11 VSUBS 0.365007f
C992 VTAIL.n8 VSUBS 2.80591f
C993 VTAIL.n9 VSUBS 1.1566f
C994 VTAIL.t6 VSUBS 3.67285f
C995 VTAIL.n10 VSUBS 3.04689f
C996 VTAIL.t0 VSUBS 3.67285f
C997 VTAIL.n11 VSUBS 2.97274f
C998 VDD1.t0 VSUBS 3.79454f
C999 VDD1.t3 VSUBS 3.79293f
C1000 VDD1.t2 VSUBS 0.35447f
C1001 VDD1.t5 VSUBS 0.35447f
C1002 VDD1.n0 VSUBS 2.90911f
C1003 VDD1.n1 VSUBS 4.5679f
C1004 VDD1.t4 VSUBS 0.35447f
C1005 VDD1.t1 VSUBS 0.35447f
C1006 VDD1.n2 VSUBS 2.90006f
C1007 VDD1.n3 VSUBS 3.91842f
C1008 VP.t4 VSUBS 3.88648f
C1009 VP.n0 VSUBS 1.4479f
C1010 VP.n1 VSUBS 0.027228f
C1011 VP.n2 VSUBS 0.022021f
C1012 VP.n3 VSUBS 0.027228f
C1013 VP.t2 VSUBS 3.88648f
C1014 VP.n4 VSUBS 1.34751f
C1015 VP.n5 VSUBS 0.027228f
C1016 VP.n6 VSUBS 0.022021f
C1017 VP.n7 VSUBS 0.027228f
C1018 VP.t1 VSUBS 3.88648f
C1019 VP.n8 VSUBS 1.4479f
C1020 VP.t5 VSUBS 3.88648f
C1021 VP.n9 VSUBS 1.4479f
C1022 VP.n10 VSUBS 0.027228f
C1023 VP.n11 VSUBS 0.022021f
C1024 VP.n12 VSUBS 0.027228f
C1025 VP.t0 VSUBS 3.88648f
C1026 VP.n13 VSUBS 1.43686f
C1027 VP.t3 VSUBS 4.2073f
C1028 VP.n14 VSUBS 1.38139f
C1029 VP.n15 VSUBS 0.316739f
C1030 VP.n16 VSUBS 0.038219f
C1031 VP.n17 VSUBS 0.050746f
C1032 VP.n18 VSUBS 0.05425f
C1033 VP.n19 VSUBS 0.027228f
C1034 VP.n20 VSUBS 0.027228f
C1035 VP.n21 VSUBS 0.027228f
C1036 VP.n22 VSUBS 0.053977f
C1037 VP.n23 VSUBS 0.050746f
C1038 VP.n24 VSUBS 0.03872f
C1039 VP.n25 VSUBS 0.043945f
C1040 VP.n26 VSUBS 1.73908f
C1041 VP.n27 VSUBS 1.7571f
C1042 VP.n28 VSUBS 0.043945f
C1043 VP.n29 VSUBS 0.03872f
C1044 VP.n30 VSUBS 0.050746f
C1045 VP.n31 VSUBS 0.053977f
C1046 VP.n32 VSUBS 0.027228f
C1047 VP.n33 VSUBS 0.027228f
C1048 VP.n34 VSUBS 0.027228f
C1049 VP.n35 VSUBS 0.05425f
C1050 VP.n36 VSUBS 0.050746f
C1051 VP.n37 VSUBS 0.038219f
C1052 VP.n38 VSUBS 0.027228f
C1053 VP.n39 VSUBS 0.027228f
C1054 VP.n40 VSUBS 0.038219f
C1055 VP.n41 VSUBS 0.050746f
C1056 VP.n42 VSUBS 0.05425f
C1057 VP.n43 VSUBS 0.027228f
C1058 VP.n44 VSUBS 0.027228f
C1059 VP.n45 VSUBS 0.027228f
C1060 VP.n46 VSUBS 0.053977f
C1061 VP.n47 VSUBS 0.050746f
C1062 VP.n48 VSUBS 0.03872f
C1063 VP.n49 VSUBS 0.043945f
C1064 VP.n50 VSUBS 0.066517f
.ends

