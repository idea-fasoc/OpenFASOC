* NGSPICE file created from diff_pair_sample_1420.ext - technology: sky130A

.subckt diff_pair_sample_1420 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9718 pd=16.02 as=1.2573 ps=7.95 w=7.62 l=0.86
X1 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=2.9718 pd=16.02 as=0 ps=0 w=7.62 l=0.86
X2 VTAIL.t10 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2573 pd=7.95 as=1.2573 ps=7.95 w=7.62 l=0.86
X3 VTAIL.t5 VN.t0 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2573 pd=7.95 as=1.2573 ps=7.95 w=7.62 l=0.86
X4 VDD1.t3 VP.t2 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2573 pd=7.95 as=2.9718 ps=16.02 w=7.62 l=0.86
X5 VDD1.t2 VP.t3 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2573 pd=7.95 as=2.9718 ps=16.02 w=7.62 l=0.86
X6 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9718 pd=16.02 as=0 ps=0 w=7.62 l=0.86
X7 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.9718 pd=16.02 as=0 ps=0 w=7.62 l=0.86
X8 VDD2.t4 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2573 pd=7.95 as=2.9718 ps=16.02 w=7.62 l=0.86
X9 VTAIL.t1 VN.t2 VDD2.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2573 pd=7.95 as=1.2573 ps=7.95 w=7.62 l=0.86
X10 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9718 pd=16.02 as=1.2573 ps=7.95 w=7.62 l=0.86
X11 VDD2.t1 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2573 pd=7.95 as=2.9718 ps=16.02 w=7.62 l=0.86
X12 VTAIL.t9 VP.t4 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2573 pd=7.95 as=1.2573 ps=7.95 w=7.62 l=0.86
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9718 pd=16.02 as=0 ps=0 w=7.62 l=0.86
X14 VDD1.t0 VP.t5 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9718 pd=16.02 as=1.2573 ps=7.95 w=7.62 l=0.86
X15 VDD2.t0 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9718 pd=16.02 as=1.2573 ps=7.95 w=7.62 l=0.86
R0 VP.n5 VP.t0 275.695
R1 VP.n12 VP.t5 259.776
R2 VP.n19 VP.t3 259.776
R3 VP.n9 VP.t2 259.776
R4 VP.n1 VP.t4 213.537
R5 VP.n4 VP.t1 213.537
R6 VP.n20 VP.n19 161.3
R7 VP.n7 VP.n6 161.3
R8 VP.n8 VP.n3 161.3
R9 VP.n10 VP.n9 161.3
R10 VP.n18 VP.n0 161.3
R11 VP.n17 VP.n16 161.3
R12 VP.n15 VP.n14 161.3
R13 VP.n13 VP.n2 161.3
R14 VP.n12 VP.n11 161.3
R15 VP.n14 VP.n13 55.5035
R16 VP.n18 VP.n17 55.5035
R17 VP.n8 VP.n7 55.5035
R18 VP.n6 VP.n5 43.768
R19 VP.n5 VP.n4 42.6032
R20 VP.n11 VP.n10 38.4816
R21 VP.n14 VP.n1 12.1722
R22 VP.n17 VP.n1 12.1722
R23 VP.n7 VP.n4 12.1722
R24 VP.n13 VP.n12 1.46111
R25 VP.n19 VP.n18 1.46111
R26 VP.n9 VP.n8 1.46111
R27 VP.n6 VP.n3 0.189894
R28 VP.n10 VP.n3 0.189894
R29 VP.n11 VP.n2 0.189894
R30 VP.n15 VP.n2 0.189894
R31 VP.n16 VP.n15 0.189894
R32 VP.n16 VP.n0 0.189894
R33 VP.n20 VP.n0 0.189894
R34 VP VP.n20 0.0516364
R35 VTAIL.n7 VTAIL.t4 53.7018
R36 VTAIL.n11 VTAIL.t3 53.7016
R37 VTAIL.n2 VTAIL.t7 53.7016
R38 VTAIL.n10 VTAIL.t11 53.7016
R39 VTAIL.n9 VTAIL.n8 51.1034
R40 VTAIL.n6 VTAIL.n5 51.1034
R41 VTAIL.n1 VTAIL.n0 51.1032
R42 VTAIL.n4 VTAIL.n3 51.1032
R43 VTAIL.n6 VTAIL.n4 20.9876
R44 VTAIL.n11 VTAIL.n10 19.9617
R45 VTAIL.n0 VTAIL.t2 2.59893
R46 VTAIL.n0 VTAIL.t5 2.59893
R47 VTAIL.n3 VTAIL.t6 2.59893
R48 VTAIL.n3 VTAIL.t9 2.59893
R49 VTAIL.n8 VTAIL.t8 2.59893
R50 VTAIL.n8 VTAIL.t10 2.59893
R51 VTAIL.n5 VTAIL.t0 2.59893
R52 VTAIL.n5 VTAIL.t1 2.59893
R53 VTAIL.n7 VTAIL.n6 1.02636
R54 VTAIL.n10 VTAIL.n9 1.02636
R55 VTAIL.n4 VTAIL.n2 1.02636
R56 VTAIL.n9 VTAIL.n7 0.983259
R57 VTAIL.n2 VTAIL.n1 0.983259
R58 VTAIL VTAIL.n11 0.711707
R59 VTAIL VTAIL.n1 0.315155
R60 VDD1 VDD1.t5 71.2082
R61 VDD1.n1 VDD1.t0 71.0945
R62 VDD1.n1 VDD1.n0 67.9831
R63 VDD1.n3 VDD1.n2 67.782
R64 VDD1.n3 VDD1.n1 34.7143
R65 VDD1.n2 VDD1.t4 2.59893
R66 VDD1.n2 VDD1.t3 2.59893
R67 VDD1.n0 VDD1.t1 2.59893
R68 VDD1.n0 VDD1.t2 2.59893
R69 VDD1 VDD1.n3 0.198776
R70 B.n392 B.n82 585
R71 B.n82 B.n43 585
R72 B.n394 B.n393 585
R73 B.n396 B.n81 585
R74 B.n399 B.n398 585
R75 B.n400 B.n80 585
R76 B.n402 B.n401 585
R77 B.n404 B.n79 585
R78 B.n407 B.n406 585
R79 B.n408 B.n78 585
R80 B.n410 B.n409 585
R81 B.n412 B.n77 585
R82 B.n415 B.n414 585
R83 B.n416 B.n76 585
R84 B.n418 B.n417 585
R85 B.n420 B.n75 585
R86 B.n423 B.n422 585
R87 B.n424 B.n74 585
R88 B.n426 B.n425 585
R89 B.n428 B.n73 585
R90 B.n431 B.n430 585
R91 B.n432 B.n72 585
R92 B.n434 B.n433 585
R93 B.n436 B.n71 585
R94 B.n439 B.n438 585
R95 B.n440 B.n70 585
R96 B.n442 B.n441 585
R97 B.n444 B.n69 585
R98 B.n446 B.n445 585
R99 B.n448 B.n447 585
R100 B.n451 B.n450 585
R101 B.n452 B.n64 585
R102 B.n454 B.n453 585
R103 B.n456 B.n63 585
R104 B.n459 B.n458 585
R105 B.n460 B.n62 585
R106 B.n462 B.n461 585
R107 B.n464 B.n61 585
R108 B.n467 B.n466 585
R109 B.n469 B.n58 585
R110 B.n471 B.n470 585
R111 B.n473 B.n57 585
R112 B.n476 B.n475 585
R113 B.n477 B.n56 585
R114 B.n479 B.n478 585
R115 B.n481 B.n55 585
R116 B.n484 B.n483 585
R117 B.n485 B.n54 585
R118 B.n487 B.n486 585
R119 B.n489 B.n53 585
R120 B.n492 B.n491 585
R121 B.n493 B.n52 585
R122 B.n495 B.n494 585
R123 B.n497 B.n51 585
R124 B.n500 B.n499 585
R125 B.n501 B.n50 585
R126 B.n503 B.n502 585
R127 B.n505 B.n49 585
R128 B.n508 B.n507 585
R129 B.n509 B.n48 585
R130 B.n511 B.n510 585
R131 B.n513 B.n47 585
R132 B.n516 B.n515 585
R133 B.n517 B.n46 585
R134 B.n519 B.n518 585
R135 B.n521 B.n45 585
R136 B.n524 B.n523 585
R137 B.n525 B.n44 585
R138 B.n391 B.n42 585
R139 B.n528 B.n42 585
R140 B.n390 B.n41 585
R141 B.n529 B.n41 585
R142 B.n389 B.n40 585
R143 B.n530 B.n40 585
R144 B.n388 B.n387 585
R145 B.n387 B.n36 585
R146 B.n386 B.n35 585
R147 B.n536 B.n35 585
R148 B.n385 B.n34 585
R149 B.n537 B.n34 585
R150 B.n384 B.n33 585
R151 B.n538 B.n33 585
R152 B.n383 B.n382 585
R153 B.n382 B.n29 585
R154 B.n381 B.n28 585
R155 B.n544 B.n28 585
R156 B.n380 B.n27 585
R157 B.n545 B.n27 585
R158 B.n379 B.n26 585
R159 B.n546 B.n26 585
R160 B.n378 B.n377 585
R161 B.n377 B.n25 585
R162 B.n376 B.n21 585
R163 B.n552 B.n21 585
R164 B.n375 B.n20 585
R165 B.n553 B.n20 585
R166 B.n374 B.n19 585
R167 B.n554 B.n19 585
R168 B.n373 B.n372 585
R169 B.n372 B.n18 585
R170 B.n371 B.n14 585
R171 B.n560 B.n14 585
R172 B.n370 B.n13 585
R173 B.n561 B.n13 585
R174 B.n369 B.n12 585
R175 B.n562 B.n12 585
R176 B.n368 B.n367 585
R177 B.n367 B.n8 585
R178 B.n366 B.n7 585
R179 B.n568 B.n7 585
R180 B.n365 B.n6 585
R181 B.n569 B.n6 585
R182 B.n364 B.n5 585
R183 B.n570 B.n5 585
R184 B.n363 B.n362 585
R185 B.n362 B.n4 585
R186 B.n361 B.n83 585
R187 B.n361 B.n360 585
R188 B.n351 B.n84 585
R189 B.n85 B.n84 585
R190 B.n353 B.n352 585
R191 B.n354 B.n353 585
R192 B.n350 B.n90 585
R193 B.n90 B.n89 585
R194 B.n349 B.n348 585
R195 B.n348 B.n347 585
R196 B.n92 B.n91 585
R197 B.n340 B.n92 585
R198 B.n339 B.n338 585
R199 B.n341 B.n339 585
R200 B.n337 B.n97 585
R201 B.n97 B.n96 585
R202 B.n336 B.n335 585
R203 B.n335 B.n334 585
R204 B.n99 B.n98 585
R205 B.n327 B.n99 585
R206 B.n326 B.n325 585
R207 B.n328 B.n326 585
R208 B.n324 B.n104 585
R209 B.n104 B.n103 585
R210 B.n323 B.n322 585
R211 B.n322 B.n321 585
R212 B.n106 B.n105 585
R213 B.n107 B.n106 585
R214 B.n314 B.n313 585
R215 B.n315 B.n314 585
R216 B.n312 B.n112 585
R217 B.n112 B.n111 585
R218 B.n311 B.n310 585
R219 B.n310 B.n309 585
R220 B.n114 B.n113 585
R221 B.n115 B.n114 585
R222 B.n302 B.n301 585
R223 B.n303 B.n302 585
R224 B.n300 B.n120 585
R225 B.n120 B.n119 585
R226 B.n299 B.n298 585
R227 B.n298 B.n297 585
R228 B.n294 B.n124 585
R229 B.n293 B.n292 585
R230 B.n290 B.n125 585
R231 B.n290 B.n123 585
R232 B.n289 B.n288 585
R233 B.n287 B.n286 585
R234 B.n285 B.n127 585
R235 B.n283 B.n282 585
R236 B.n281 B.n128 585
R237 B.n280 B.n279 585
R238 B.n277 B.n129 585
R239 B.n275 B.n274 585
R240 B.n273 B.n130 585
R241 B.n272 B.n271 585
R242 B.n269 B.n131 585
R243 B.n267 B.n266 585
R244 B.n265 B.n132 585
R245 B.n264 B.n263 585
R246 B.n261 B.n133 585
R247 B.n259 B.n258 585
R248 B.n257 B.n134 585
R249 B.n256 B.n255 585
R250 B.n253 B.n135 585
R251 B.n251 B.n250 585
R252 B.n249 B.n136 585
R253 B.n248 B.n247 585
R254 B.n245 B.n137 585
R255 B.n243 B.n242 585
R256 B.n241 B.n138 585
R257 B.n240 B.n239 585
R258 B.n237 B.n236 585
R259 B.n235 B.n234 585
R260 B.n233 B.n143 585
R261 B.n231 B.n230 585
R262 B.n229 B.n144 585
R263 B.n228 B.n227 585
R264 B.n225 B.n145 585
R265 B.n223 B.n222 585
R266 B.n221 B.n146 585
R267 B.n219 B.n218 585
R268 B.n216 B.n149 585
R269 B.n214 B.n213 585
R270 B.n212 B.n150 585
R271 B.n211 B.n210 585
R272 B.n208 B.n151 585
R273 B.n206 B.n205 585
R274 B.n204 B.n152 585
R275 B.n203 B.n202 585
R276 B.n200 B.n153 585
R277 B.n198 B.n197 585
R278 B.n196 B.n154 585
R279 B.n195 B.n194 585
R280 B.n192 B.n155 585
R281 B.n190 B.n189 585
R282 B.n188 B.n156 585
R283 B.n187 B.n186 585
R284 B.n184 B.n157 585
R285 B.n182 B.n181 585
R286 B.n180 B.n158 585
R287 B.n179 B.n178 585
R288 B.n176 B.n159 585
R289 B.n174 B.n173 585
R290 B.n172 B.n160 585
R291 B.n171 B.n170 585
R292 B.n168 B.n161 585
R293 B.n166 B.n165 585
R294 B.n164 B.n163 585
R295 B.n122 B.n121 585
R296 B.n296 B.n295 585
R297 B.n297 B.n296 585
R298 B.n118 B.n117 585
R299 B.n119 B.n118 585
R300 B.n305 B.n304 585
R301 B.n304 B.n303 585
R302 B.n306 B.n116 585
R303 B.n116 B.n115 585
R304 B.n308 B.n307 585
R305 B.n309 B.n308 585
R306 B.n110 B.n109 585
R307 B.n111 B.n110 585
R308 B.n317 B.n316 585
R309 B.n316 B.n315 585
R310 B.n318 B.n108 585
R311 B.n108 B.n107 585
R312 B.n320 B.n319 585
R313 B.n321 B.n320 585
R314 B.n102 B.n101 585
R315 B.n103 B.n102 585
R316 B.n330 B.n329 585
R317 B.n329 B.n328 585
R318 B.n331 B.n100 585
R319 B.n327 B.n100 585
R320 B.n333 B.n332 585
R321 B.n334 B.n333 585
R322 B.n95 B.n94 585
R323 B.n96 B.n95 585
R324 B.n343 B.n342 585
R325 B.n342 B.n341 585
R326 B.n344 B.n93 585
R327 B.n340 B.n93 585
R328 B.n346 B.n345 585
R329 B.n347 B.n346 585
R330 B.n88 B.n87 585
R331 B.n89 B.n88 585
R332 B.n356 B.n355 585
R333 B.n355 B.n354 585
R334 B.n357 B.n86 585
R335 B.n86 B.n85 585
R336 B.n359 B.n358 585
R337 B.n360 B.n359 585
R338 B.n2 B.n0 585
R339 B.n4 B.n2 585
R340 B.n3 B.n1 585
R341 B.n569 B.n3 585
R342 B.n567 B.n566 585
R343 B.n568 B.n567 585
R344 B.n565 B.n9 585
R345 B.n9 B.n8 585
R346 B.n564 B.n563 585
R347 B.n563 B.n562 585
R348 B.n11 B.n10 585
R349 B.n561 B.n11 585
R350 B.n559 B.n558 585
R351 B.n560 B.n559 585
R352 B.n557 B.n15 585
R353 B.n18 B.n15 585
R354 B.n556 B.n555 585
R355 B.n555 B.n554 585
R356 B.n17 B.n16 585
R357 B.n553 B.n17 585
R358 B.n551 B.n550 585
R359 B.n552 B.n551 585
R360 B.n549 B.n22 585
R361 B.n25 B.n22 585
R362 B.n548 B.n547 585
R363 B.n547 B.n546 585
R364 B.n24 B.n23 585
R365 B.n545 B.n24 585
R366 B.n543 B.n542 585
R367 B.n544 B.n543 585
R368 B.n541 B.n30 585
R369 B.n30 B.n29 585
R370 B.n540 B.n539 585
R371 B.n539 B.n538 585
R372 B.n32 B.n31 585
R373 B.n537 B.n32 585
R374 B.n535 B.n534 585
R375 B.n536 B.n535 585
R376 B.n533 B.n37 585
R377 B.n37 B.n36 585
R378 B.n532 B.n531 585
R379 B.n531 B.n530 585
R380 B.n39 B.n38 585
R381 B.n529 B.n39 585
R382 B.n527 B.n526 585
R383 B.n528 B.n527 585
R384 B.n572 B.n571 585
R385 B.n571 B.n570 585
R386 B.n296 B.n124 521.33
R387 B.n527 B.n44 521.33
R388 B.n298 B.n122 521.33
R389 B.n82 B.n42 521.33
R390 B.n147 B.t17 416.051
R391 B.n65 B.t14 416.051
R392 B.n139 B.t10 415.44
R393 B.n59 B.t6 415.44
R394 B.n395 B.n43 256.663
R395 B.n397 B.n43 256.663
R396 B.n403 B.n43 256.663
R397 B.n405 B.n43 256.663
R398 B.n411 B.n43 256.663
R399 B.n413 B.n43 256.663
R400 B.n419 B.n43 256.663
R401 B.n421 B.n43 256.663
R402 B.n427 B.n43 256.663
R403 B.n429 B.n43 256.663
R404 B.n435 B.n43 256.663
R405 B.n437 B.n43 256.663
R406 B.n443 B.n43 256.663
R407 B.n68 B.n43 256.663
R408 B.n449 B.n43 256.663
R409 B.n455 B.n43 256.663
R410 B.n457 B.n43 256.663
R411 B.n463 B.n43 256.663
R412 B.n465 B.n43 256.663
R413 B.n472 B.n43 256.663
R414 B.n474 B.n43 256.663
R415 B.n480 B.n43 256.663
R416 B.n482 B.n43 256.663
R417 B.n488 B.n43 256.663
R418 B.n490 B.n43 256.663
R419 B.n496 B.n43 256.663
R420 B.n498 B.n43 256.663
R421 B.n504 B.n43 256.663
R422 B.n506 B.n43 256.663
R423 B.n512 B.n43 256.663
R424 B.n514 B.n43 256.663
R425 B.n520 B.n43 256.663
R426 B.n522 B.n43 256.663
R427 B.n291 B.n123 256.663
R428 B.n126 B.n123 256.663
R429 B.n284 B.n123 256.663
R430 B.n278 B.n123 256.663
R431 B.n276 B.n123 256.663
R432 B.n270 B.n123 256.663
R433 B.n268 B.n123 256.663
R434 B.n262 B.n123 256.663
R435 B.n260 B.n123 256.663
R436 B.n254 B.n123 256.663
R437 B.n252 B.n123 256.663
R438 B.n246 B.n123 256.663
R439 B.n244 B.n123 256.663
R440 B.n238 B.n123 256.663
R441 B.n142 B.n123 256.663
R442 B.n232 B.n123 256.663
R443 B.n226 B.n123 256.663
R444 B.n224 B.n123 256.663
R445 B.n217 B.n123 256.663
R446 B.n215 B.n123 256.663
R447 B.n209 B.n123 256.663
R448 B.n207 B.n123 256.663
R449 B.n201 B.n123 256.663
R450 B.n199 B.n123 256.663
R451 B.n193 B.n123 256.663
R452 B.n191 B.n123 256.663
R453 B.n185 B.n123 256.663
R454 B.n183 B.n123 256.663
R455 B.n177 B.n123 256.663
R456 B.n175 B.n123 256.663
R457 B.n169 B.n123 256.663
R458 B.n167 B.n123 256.663
R459 B.n162 B.n123 256.663
R460 B.n296 B.n118 163.367
R461 B.n304 B.n118 163.367
R462 B.n304 B.n116 163.367
R463 B.n308 B.n116 163.367
R464 B.n308 B.n110 163.367
R465 B.n316 B.n110 163.367
R466 B.n316 B.n108 163.367
R467 B.n320 B.n108 163.367
R468 B.n320 B.n102 163.367
R469 B.n329 B.n102 163.367
R470 B.n329 B.n100 163.367
R471 B.n333 B.n100 163.367
R472 B.n333 B.n95 163.367
R473 B.n342 B.n95 163.367
R474 B.n342 B.n93 163.367
R475 B.n346 B.n93 163.367
R476 B.n346 B.n88 163.367
R477 B.n355 B.n88 163.367
R478 B.n355 B.n86 163.367
R479 B.n359 B.n86 163.367
R480 B.n359 B.n2 163.367
R481 B.n571 B.n2 163.367
R482 B.n571 B.n3 163.367
R483 B.n567 B.n3 163.367
R484 B.n567 B.n9 163.367
R485 B.n563 B.n9 163.367
R486 B.n563 B.n11 163.367
R487 B.n559 B.n11 163.367
R488 B.n559 B.n15 163.367
R489 B.n555 B.n15 163.367
R490 B.n555 B.n17 163.367
R491 B.n551 B.n17 163.367
R492 B.n551 B.n22 163.367
R493 B.n547 B.n22 163.367
R494 B.n547 B.n24 163.367
R495 B.n543 B.n24 163.367
R496 B.n543 B.n30 163.367
R497 B.n539 B.n30 163.367
R498 B.n539 B.n32 163.367
R499 B.n535 B.n32 163.367
R500 B.n535 B.n37 163.367
R501 B.n531 B.n37 163.367
R502 B.n531 B.n39 163.367
R503 B.n527 B.n39 163.367
R504 B.n292 B.n290 163.367
R505 B.n290 B.n289 163.367
R506 B.n286 B.n285 163.367
R507 B.n283 B.n128 163.367
R508 B.n279 B.n277 163.367
R509 B.n275 B.n130 163.367
R510 B.n271 B.n269 163.367
R511 B.n267 B.n132 163.367
R512 B.n263 B.n261 163.367
R513 B.n259 B.n134 163.367
R514 B.n255 B.n253 163.367
R515 B.n251 B.n136 163.367
R516 B.n247 B.n245 163.367
R517 B.n243 B.n138 163.367
R518 B.n239 B.n237 163.367
R519 B.n234 B.n233 163.367
R520 B.n231 B.n144 163.367
R521 B.n227 B.n225 163.367
R522 B.n223 B.n146 163.367
R523 B.n218 B.n216 163.367
R524 B.n214 B.n150 163.367
R525 B.n210 B.n208 163.367
R526 B.n206 B.n152 163.367
R527 B.n202 B.n200 163.367
R528 B.n198 B.n154 163.367
R529 B.n194 B.n192 163.367
R530 B.n190 B.n156 163.367
R531 B.n186 B.n184 163.367
R532 B.n182 B.n158 163.367
R533 B.n178 B.n176 163.367
R534 B.n174 B.n160 163.367
R535 B.n170 B.n168 163.367
R536 B.n166 B.n163 163.367
R537 B.n298 B.n120 163.367
R538 B.n302 B.n120 163.367
R539 B.n302 B.n114 163.367
R540 B.n310 B.n114 163.367
R541 B.n310 B.n112 163.367
R542 B.n314 B.n112 163.367
R543 B.n314 B.n106 163.367
R544 B.n322 B.n106 163.367
R545 B.n322 B.n104 163.367
R546 B.n326 B.n104 163.367
R547 B.n326 B.n99 163.367
R548 B.n335 B.n99 163.367
R549 B.n335 B.n97 163.367
R550 B.n339 B.n97 163.367
R551 B.n339 B.n92 163.367
R552 B.n348 B.n92 163.367
R553 B.n348 B.n90 163.367
R554 B.n353 B.n90 163.367
R555 B.n353 B.n84 163.367
R556 B.n361 B.n84 163.367
R557 B.n362 B.n361 163.367
R558 B.n362 B.n5 163.367
R559 B.n6 B.n5 163.367
R560 B.n7 B.n6 163.367
R561 B.n367 B.n7 163.367
R562 B.n367 B.n12 163.367
R563 B.n13 B.n12 163.367
R564 B.n14 B.n13 163.367
R565 B.n372 B.n14 163.367
R566 B.n372 B.n19 163.367
R567 B.n20 B.n19 163.367
R568 B.n21 B.n20 163.367
R569 B.n377 B.n21 163.367
R570 B.n377 B.n26 163.367
R571 B.n27 B.n26 163.367
R572 B.n28 B.n27 163.367
R573 B.n382 B.n28 163.367
R574 B.n382 B.n33 163.367
R575 B.n34 B.n33 163.367
R576 B.n35 B.n34 163.367
R577 B.n387 B.n35 163.367
R578 B.n387 B.n40 163.367
R579 B.n41 B.n40 163.367
R580 B.n42 B.n41 163.367
R581 B.n523 B.n521 163.367
R582 B.n519 B.n46 163.367
R583 B.n515 B.n513 163.367
R584 B.n511 B.n48 163.367
R585 B.n507 B.n505 163.367
R586 B.n503 B.n50 163.367
R587 B.n499 B.n497 163.367
R588 B.n495 B.n52 163.367
R589 B.n491 B.n489 163.367
R590 B.n487 B.n54 163.367
R591 B.n483 B.n481 163.367
R592 B.n479 B.n56 163.367
R593 B.n475 B.n473 163.367
R594 B.n471 B.n58 163.367
R595 B.n466 B.n464 163.367
R596 B.n462 B.n62 163.367
R597 B.n458 B.n456 163.367
R598 B.n454 B.n64 163.367
R599 B.n450 B.n448 163.367
R600 B.n445 B.n444 163.367
R601 B.n442 B.n70 163.367
R602 B.n438 B.n436 163.367
R603 B.n434 B.n72 163.367
R604 B.n430 B.n428 163.367
R605 B.n426 B.n74 163.367
R606 B.n422 B.n420 163.367
R607 B.n418 B.n76 163.367
R608 B.n414 B.n412 163.367
R609 B.n410 B.n78 163.367
R610 B.n406 B.n404 163.367
R611 B.n402 B.n80 163.367
R612 B.n398 B.n396 163.367
R613 B.n394 B.n82 163.367
R614 B.n297 B.n123 111.749
R615 B.n528 B.n43 111.749
R616 B.n147 B.t19 94.7211
R617 B.n65 B.t15 94.7211
R618 B.n139 B.t13 94.7124
R619 B.n59 B.t8 94.7124
R620 B.n291 B.n124 71.676
R621 B.n289 B.n126 71.676
R622 B.n285 B.n284 71.676
R623 B.n278 B.n128 71.676
R624 B.n277 B.n276 71.676
R625 B.n270 B.n130 71.676
R626 B.n269 B.n268 71.676
R627 B.n262 B.n132 71.676
R628 B.n261 B.n260 71.676
R629 B.n254 B.n134 71.676
R630 B.n253 B.n252 71.676
R631 B.n246 B.n136 71.676
R632 B.n245 B.n244 71.676
R633 B.n238 B.n138 71.676
R634 B.n237 B.n142 71.676
R635 B.n233 B.n232 71.676
R636 B.n226 B.n144 71.676
R637 B.n225 B.n224 71.676
R638 B.n217 B.n146 71.676
R639 B.n216 B.n215 71.676
R640 B.n209 B.n150 71.676
R641 B.n208 B.n207 71.676
R642 B.n201 B.n152 71.676
R643 B.n200 B.n199 71.676
R644 B.n193 B.n154 71.676
R645 B.n192 B.n191 71.676
R646 B.n185 B.n156 71.676
R647 B.n184 B.n183 71.676
R648 B.n177 B.n158 71.676
R649 B.n176 B.n175 71.676
R650 B.n169 B.n160 71.676
R651 B.n168 B.n167 71.676
R652 B.n163 B.n162 71.676
R653 B.n522 B.n44 71.676
R654 B.n521 B.n520 71.676
R655 B.n514 B.n46 71.676
R656 B.n513 B.n512 71.676
R657 B.n506 B.n48 71.676
R658 B.n505 B.n504 71.676
R659 B.n498 B.n50 71.676
R660 B.n497 B.n496 71.676
R661 B.n490 B.n52 71.676
R662 B.n489 B.n488 71.676
R663 B.n482 B.n54 71.676
R664 B.n481 B.n480 71.676
R665 B.n474 B.n56 71.676
R666 B.n473 B.n472 71.676
R667 B.n465 B.n58 71.676
R668 B.n464 B.n463 71.676
R669 B.n457 B.n62 71.676
R670 B.n456 B.n455 71.676
R671 B.n449 B.n64 71.676
R672 B.n448 B.n68 71.676
R673 B.n444 B.n443 71.676
R674 B.n437 B.n70 71.676
R675 B.n436 B.n435 71.676
R676 B.n429 B.n72 71.676
R677 B.n428 B.n427 71.676
R678 B.n421 B.n74 71.676
R679 B.n420 B.n419 71.676
R680 B.n413 B.n76 71.676
R681 B.n412 B.n411 71.676
R682 B.n405 B.n78 71.676
R683 B.n404 B.n403 71.676
R684 B.n397 B.n80 71.676
R685 B.n396 B.n395 71.676
R686 B.n395 B.n394 71.676
R687 B.n398 B.n397 71.676
R688 B.n403 B.n402 71.676
R689 B.n406 B.n405 71.676
R690 B.n411 B.n410 71.676
R691 B.n414 B.n413 71.676
R692 B.n419 B.n418 71.676
R693 B.n422 B.n421 71.676
R694 B.n427 B.n426 71.676
R695 B.n430 B.n429 71.676
R696 B.n435 B.n434 71.676
R697 B.n438 B.n437 71.676
R698 B.n443 B.n442 71.676
R699 B.n445 B.n68 71.676
R700 B.n450 B.n449 71.676
R701 B.n455 B.n454 71.676
R702 B.n458 B.n457 71.676
R703 B.n463 B.n462 71.676
R704 B.n466 B.n465 71.676
R705 B.n472 B.n471 71.676
R706 B.n475 B.n474 71.676
R707 B.n480 B.n479 71.676
R708 B.n483 B.n482 71.676
R709 B.n488 B.n487 71.676
R710 B.n491 B.n490 71.676
R711 B.n496 B.n495 71.676
R712 B.n499 B.n498 71.676
R713 B.n504 B.n503 71.676
R714 B.n507 B.n506 71.676
R715 B.n512 B.n511 71.676
R716 B.n515 B.n514 71.676
R717 B.n520 B.n519 71.676
R718 B.n523 B.n522 71.676
R719 B.n292 B.n291 71.676
R720 B.n286 B.n126 71.676
R721 B.n284 B.n283 71.676
R722 B.n279 B.n278 71.676
R723 B.n276 B.n275 71.676
R724 B.n271 B.n270 71.676
R725 B.n268 B.n267 71.676
R726 B.n263 B.n262 71.676
R727 B.n260 B.n259 71.676
R728 B.n255 B.n254 71.676
R729 B.n252 B.n251 71.676
R730 B.n247 B.n246 71.676
R731 B.n244 B.n243 71.676
R732 B.n239 B.n238 71.676
R733 B.n234 B.n142 71.676
R734 B.n232 B.n231 71.676
R735 B.n227 B.n226 71.676
R736 B.n224 B.n223 71.676
R737 B.n218 B.n217 71.676
R738 B.n215 B.n214 71.676
R739 B.n210 B.n209 71.676
R740 B.n207 B.n206 71.676
R741 B.n202 B.n201 71.676
R742 B.n199 B.n198 71.676
R743 B.n194 B.n193 71.676
R744 B.n191 B.n190 71.676
R745 B.n186 B.n185 71.676
R746 B.n183 B.n182 71.676
R747 B.n178 B.n177 71.676
R748 B.n175 B.n174 71.676
R749 B.n170 B.n169 71.676
R750 B.n167 B.n166 71.676
R751 B.n162 B.n122 71.676
R752 B.n148 B.t18 71.6423
R753 B.n66 B.t16 71.6423
R754 B.n140 B.t12 71.6336
R755 B.n60 B.t9 71.6336
R756 B.n220 B.n148 59.5399
R757 B.n141 B.n140 59.5399
R758 B.n468 B.n60 59.5399
R759 B.n67 B.n66 59.5399
R760 B.n297 B.n119 58.0075
R761 B.n303 B.n119 58.0075
R762 B.n303 B.n115 58.0075
R763 B.n309 B.n115 58.0075
R764 B.n315 B.n111 58.0075
R765 B.n315 B.n107 58.0075
R766 B.n321 B.n107 58.0075
R767 B.n321 B.n103 58.0075
R768 B.n328 B.n103 58.0075
R769 B.n328 B.n327 58.0075
R770 B.n334 B.n96 58.0075
R771 B.n341 B.n96 58.0075
R772 B.n341 B.n340 58.0075
R773 B.n347 B.n89 58.0075
R774 B.n354 B.n89 58.0075
R775 B.n360 B.n85 58.0075
R776 B.n360 B.n4 58.0075
R777 B.n570 B.n4 58.0075
R778 B.n570 B.n569 58.0075
R779 B.n569 B.n568 58.0075
R780 B.n568 B.n8 58.0075
R781 B.n562 B.n561 58.0075
R782 B.n561 B.n560 58.0075
R783 B.n554 B.n18 58.0075
R784 B.n554 B.n553 58.0075
R785 B.n553 B.n552 58.0075
R786 B.n546 B.n25 58.0075
R787 B.n546 B.n545 58.0075
R788 B.n545 B.n544 58.0075
R789 B.n544 B.n29 58.0075
R790 B.n538 B.n29 58.0075
R791 B.n538 B.n537 58.0075
R792 B.n536 B.n36 58.0075
R793 B.n530 B.n36 58.0075
R794 B.n530 B.n529 58.0075
R795 B.n529 B.n528 58.0075
R796 B.n309 B.t11 54.5953
R797 B.t7 B.n536 54.5953
R798 B.n347 B.t1 49.477
R799 B.n560 B.t5 49.477
R800 B.n327 B.t0 37.5344
R801 B.n354 B.t4 37.5344
R802 B.n562 B.t2 37.5344
R803 B.n25 B.t3 37.5344
R804 B.n526 B.n525 33.8737
R805 B.n392 B.n391 33.8737
R806 B.n299 B.n121 33.8737
R807 B.n295 B.n294 33.8737
R808 B.n148 B.n147 23.0793
R809 B.n140 B.n139 23.0793
R810 B.n60 B.n59 23.0793
R811 B.n66 B.n65 23.0793
R812 B.n334 B.t0 20.4736
R813 B.t4 B.n85 20.4736
R814 B.t2 B.n8 20.4736
R815 B.n552 B.t3 20.4736
R816 B B.n572 18.0485
R817 B.n525 B.n524 10.6151
R818 B.n524 B.n45 10.6151
R819 B.n518 B.n45 10.6151
R820 B.n518 B.n517 10.6151
R821 B.n517 B.n516 10.6151
R822 B.n516 B.n47 10.6151
R823 B.n510 B.n47 10.6151
R824 B.n510 B.n509 10.6151
R825 B.n509 B.n508 10.6151
R826 B.n508 B.n49 10.6151
R827 B.n502 B.n49 10.6151
R828 B.n502 B.n501 10.6151
R829 B.n501 B.n500 10.6151
R830 B.n500 B.n51 10.6151
R831 B.n494 B.n51 10.6151
R832 B.n494 B.n493 10.6151
R833 B.n493 B.n492 10.6151
R834 B.n492 B.n53 10.6151
R835 B.n486 B.n53 10.6151
R836 B.n486 B.n485 10.6151
R837 B.n485 B.n484 10.6151
R838 B.n484 B.n55 10.6151
R839 B.n478 B.n55 10.6151
R840 B.n478 B.n477 10.6151
R841 B.n477 B.n476 10.6151
R842 B.n476 B.n57 10.6151
R843 B.n470 B.n57 10.6151
R844 B.n470 B.n469 10.6151
R845 B.n467 B.n61 10.6151
R846 B.n461 B.n61 10.6151
R847 B.n461 B.n460 10.6151
R848 B.n460 B.n459 10.6151
R849 B.n459 B.n63 10.6151
R850 B.n453 B.n63 10.6151
R851 B.n453 B.n452 10.6151
R852 B.n452 B.n451 10.6151
R853 B.n447 B.n446 10.6151
R854 B.n446 B.n69 10.6151
R855 B.n441 B.n69 10.6151
R856 B.n441 B.n440 10.6151
R857 B.n440 B.n439 10.6151
R858 B.n439 B.n71 10.6151
R859 B.n433 B.n71 10.6151
R860 B.n433 B.n432 10.6151
R861 B.n432 B.n431 10.6151
R862 B.n431 B.n73 10.6151
R863 B.n425 B.n73 10.6151
R864 B.n425 B.n424 10.6151
R865 B.n424 B.n423 10.6151
R866 B.n423 B.n75 10.6151
R867 B.n417 B.n75 10.6151
R868 B.n417 B.n416 10.6151
R869 B.n416 B.n415 10.6151
R870 B.n415 B.n77 10.6151
R871 B.n409 B.n77 10.6151
R872 B.n409 B.n408 10.6151
R873 B.n408 B.n407 10.6151
R874 B.n407 B.n79 10.6151
R875 B.n401 B.n79 10.6151
R876 B.n401 B.n400 10.6151
R877 B.n400 B.n399 10.6151
R878 B.n399 B.n81 10.6151
R879 B.n393 B.n81 10.6151
R880 B.n393 B.n392 10.6151
R881 B.n300 B.n299 10.6151
R882 B.n301 B.n300 10.6151
R883 B.n301 B.n113 10.6151
R884 B.n311 B.n113 10.6151
R885 B.n312 B.n311 10.6151
R886 B.n313 B.n312 10.6151
R887 B.n313 B.n105 10.6151
R888 B.n323 B.n105 10.6151
R889 B.n324 B.n323 10.6151
R890 B.n325 B.n324 10.6151
R891 B.n325 B.n98 10.6151
R892 B.n336 B.n98 10.6151
R893 B.n337 B.n336 10.6151
R894 B.n338 B.n337 10.6151
R895 B.n338 B.n91 10.6151
R896 B.n349 B.n91 10.6151
R897 B.n350 B.n349 10.6151
R898 B.n352 B.n350 10.6151
R899 B.n352 B.n351 10.6151
R900 B.n351 B.n83 10.6151
R901 B.n363 B.n83 10.6151
R902 B.n364 B.n363 10.6151
R903 B.n365 B.n364 10.6151
R904 B.n366 B.n365 10.6151
R905 B.n368 B.n366 10.6151
R906 B.n369 B.n368 10.6151
R907 B.n370 B.n369 10.6151
R908 B.n371 B.n370 10.6151
R909 B.n373 B.n371 10.6151
R910 B.n374 B.n373 10.6151
R911 B.n375 B.n374 10.6151
R912 B.n376 B.n375 10.6151
R913 B.n378 B.n376 10.6151
R914 B.n379 B.n378 10.6151
R915 B.n380 B.n379 10.6151
R916 B.n381 B.n380 10.6151
R917 B.n383 B.n381 10.6151
R918 B.n384 B.n383 10.6151
R919 B.n385 B.n384 10.6151
R920 B.n386 B.n385 10.6151
R921 B.n388 B.n386 10.6151
R922 B.n389 B.n388 10.6151
R923 B.n390 B.n389 10.6151
R924 B.n391 B.n390 10.6151
R925 B.n294 B.n293 10.6151
R926 B.n293 B.n125 10.6151
R927 B.n288 B.n125 10.6151
R928 B.n288 B.n287 10.6151
R929 B.n287 B.n127 10.6151
R930 B.n282 B.n127 10.6151
R931 B.n282 B.n281 10.6151
R932 B.n281 B.n280 10.6151
R933 B.n280 B.n129 10.6151
R934 B.n274 B.n129 10.6151
R935 B.n274 B.n273 10.6151
R936 B.n273 B.n272 10.6151
R937 B.n272 B.n131 10.6151
R938 B.n266 B.n131 10.6151
R939 B.n266 B.n265 10.6151
R940 B.n265 B.n264 10.6151
R941 B.n264 B.n133 10.6151
R942 B.n258 B.n133 10.6151
R943 B.n258 B.n257 10.6151
R944 B.n257 B.n256 10.6151
R945 B.n256 B.n135 10.6151
R946 B.n250 B.n135 10.6151
R947 B.n250 B.n249 10.6151
R948 B.n249 B.n248 10.6151
R949 B.n248 B.n137 10.6151
R950 B.n242 B.n137 10.6151
R951 B.n242 B.n241 10.6151
R952 B.n241 B.n240 10.6151
R953 B.n236 B.n235 10.6151
R954 B.n235 B.n143 10.6151
R955 B.n230 B.n143 10.6151
R956 B.n230 B.n229 10.6151
R957 B.n229 B.n228 10.6151
R958 B.n228 B.n145 10.6151
R959 B.n222 B.n145 10.6151
R960 B.n222 B.n221 10.6151
R961 B.n219 B.n149 10.6151
R962 B.n213 B.n149 10.6151
R963 B.n213 B.n212 10.6151
R964 B.n212 B.n211 10.6151
R965 B.n211 B.n151 10.6151
R966 B.n205 B.n151 10.6151
R967 B.n205 B.n204 10.6151
R968 B.n204 B.n203 10.6151
R969 B.n203 B.n153 10.6151
R970 B.n197 B.n153 10.6151
R971 B.n197 B.n196 10.6151
R972 B.n196 B.n195 10.6151
R973 B.n195 B.n155 10.6151
R974 B.n189 B.n155 10.6151
R975 B.n189 B.n188 10.6151
R976 B.n188 B.n187 10.6151
R977 B.n187 B.n157 10.6151
R978 B.n181 B.n157 10.6151
R979 B.n181 B.n180 10.6151
R980 B.n180 B.n179 10.6151
R981 B.n179 B.n159 10.6151
R982 B.n173 B.n159 10.6151
R983 B.n173 B.n172 10.6151
R984 B.n172 B.n171 10.6151
R985 B.n171 B.n161 10.6151
R986 B.n165 B.n161 10.6151
R987 B.n165 B.n164 10.6151
R988 B.n164 B.n121 10.6151
R989 B.n295 B.n117 10.6151
R990 B.n305 B.n117 10.6151
R991 B.n306 B.n305 10.6151
R992 B.n307 B.n306 10.6151
R993 B.n307 B.n109 10.6151
R994 B.n317 B.n109 10.6151
R995 B.n318 B.n317 10.6151
R996 B.n319 B.n318 10.6151
R997 B.n319 B.n101 10.6151
R998 B.n330 B.n101 10.6151
R999 B.n331 B.n330 10.6151
R1000 B.n332 B.n331 10.6151
R1001 B.n332 B.n94 10.6151
R1002 B.n343 B.n94 10.6151
R1003 B.n344 B.n343 10.6151
R1004 B.n345 B.n344 10.6151
R1005 B.n345 B.n87 10.6151
R1006 B.n356 B.n87 10.6151
R1007 B.n357 B.n356 10.6151
R1008 B.n358 B.n357 10.6151
R1009 B.n358 B.n0 10.6151
R1010 B.n566 B.n1 10.6151
R1011 B.n566 B.n565 10.6151
R1012 B.n565 B.n564 10.6151
R1013 B.n564 B.n10 10.6151
R1014 B.n558 B.n10 10.6151
R1015 B.n558 B.n557 10.6151
R1016 B.n557 B.n556 10.6151
R1017 B.n556 B.n16 10.6151
R1018 B.n550 B.n16 10.6151
R1019 B.n550 B.n549 10.6151
R1020 B.n549 B.n548 10.6151
R1021 B.n548 B.n23 10.6151
R1022 B.n542 B.n23 10.6151
R1023 B.n542 B.n541 10.6151
R1024 B.n541 B.n540 10.6151
R1025 B.n540 B.n31 10.6151
R1026 B.n534 B.n31 10.6151
R1027 B.n534 B.n533 10.6151
R1028 B.n533 B.n532 10.6151
R1029 B.n532 B.n38 10.6151
R1030 B.n526 B.n38 10.6151
R1031 B.n340 B.t1 8.53094
R1032 B.n18 B.t5 8.53094
R1033 B.n468 B.n467 6.4005
R1034 B.n451 B.n67 6.4005
R1035 B.n236 B.n141 6.4005
R1036 B.n221 B.n220 6.4005
R1037 B.n469 B.n468 4.21513
R1038 B.n447 B.n67 4.21513
R1039 B.n240 B.n141 4.21513
R1040 B.n220 B.n219 4.21513
R1041 B.t11 B.n111 3.41268
R1042 B.n537 B.t7 3.41268
R1043 B.n572 B.n0 2.81026
R1044 B.n572 B.n1 2.81026
R1045 VN.n2 VN.t3 275.695
R1046 VN.n10 VN.t1 275.695
R1047 VN.n6 VN.t4 259.776
R1048 VN.n14 VN.t5 259.776
R1049 VN.n1 VN.t0 213.537
R1050 VN.n9 VN.t2 213.537
R1051 VN.n7 VN.n6 161.3
R1052 VN.n15 VN.n14 161.3
R1053 VN.n13 VN.n8 161.3
R1054 VN.n12 VN.n11 161.3
R1055 VN.n5 VN.n0 161.3
R1056 VN.n4 VN.n3 161.3
R1057 VN.n5 VN.n4 55.5035
R1058 VN.n13 VN.n12 55.5035
R1059 VN.n11 VN.n10 43.768
R1060 VN.n3 VN.n2 43.768
R1061 VN.n2 VN.n1 42.6032
R1062 VN.n10 VN.n9 42.6032
R1063 VN VN.n15 38.8622
R1064 VN.n4 VN.n1 12.1722
R1065 VN.n12 VN.n9 12.1722
R1066 VN.n6 VN.n5 1.46111
R1067 VN.n14 VN.n13 1.46111
R1068 VN.n15 VN.n8 0.189894
R1069 VN.n11 VN.n8 0.189894
R1070 VN.n3 VN.n0 0.189894
R1071 VN.n7 VN.n0 0.189894
R1072 VN VN.n7 0.0516364
R1073 VDD2.n1 VDD2.t2 71.0945
R1074 VDD2.n2 VDD2.t0 70.3806
R1075 VDD2.n1 VDD2.n0 67.9831
R1076 VDD2 VDD2.n3 67.9803
R1077 VDD2.n2 VDD2.n1 33.6183
R1078 VDD2.n3 VDD2.t3 2.59893
R1079 VDD2.n3 VDD2.t4 2.59893
R1080 VDD2.n0 VDD2.t5 2.59893
R1081 VDD2.n0 VDD2.t1 2.59893
R1082 VDD2 VDD2.n2 0.828086
C0 VP VTAIL 3.07452f
C1 VDD1 VTAIL 6.59427f
C2 VN VDD2 3.15401f
C3 VP VDD2 0.310207f
C4 VP VN 4.42993f
C5 VDD1 VDD2 0.76804f
C6 VDD1 VN 0.148071f
C7 VDD1 VP 3.31325f
C8 VDD2 VTAIL 6.63224f
C9 VN VTAIL 3.06012f
C10 VDD2 B 3.827258f
C11 VDD1 B 4.060594f
C12 VTAIL B 4.908561f
C13 VN B 7.635591f
C14 VP B 5.958216f
C15 VDD2.t2 B 1.51325f
C16 VDD2.t5 B 0.137611f
C17 VDD2.t1 B 0.137611f
C18 VDD2.n0 B 1.18844f
C19 VDD2.n1 B 1.70552f
C20 VDD2.t0 B 1.51028f
C21 VDD2.n2 B 1.78964f
C22 VDD2.t3 B 0.137611f
C23 VDD2.t4 B 0.137611f
C24 VDD2.n3 B 1.18842f
C25 VN.n0 B 0.04338f
C26 VN.t0 B 0.761126f
C27 VN.n1 B 0.345007f
C28 VN.t3 B 0.839434f
C29 VN.n2 B 0.356441f
C30 VN.n3 B 0.17907f
C31 VN.n4 B 0.054889f
C32 VN.n5 B 0.013476f
C33 VN.t4 B 0.818629f
C34 VN.n6 B 0.347347f
C35 VN.n7 B 0.033618f
C36 VN.n8 B 0.04338f
C37 VN.t2 B 0.761126f
C38 VN.n9 B 0.345007f
C39 VN.t1 B 0.839434f
C40 VN.n10 B 0.356441f
C41 VN.n11 B 0.17907f
C42 VN.n12 B 0.054889f
C43 VN.n13 B 0.013476f
C44 VN.t5 B 0.818629f
C45 VN.n14 B 0.347347f
C46 VN.n15 B 1.56915f
C47 VDD1.t5 B 1.51619f
C48 VDD1.t0 B 1.51563f
C49 VDD1.t1 B 0.137828f
C50 VDD1.t2 B 0.137828f
C51 VDD1.n0 B 1.19031f
C52 VDD1.n1 B 1.78045f
C53 VDD1.t4 B 0.137828f
C54 VDD1.t3 B 0.137828f
C55 VDD1.n2 B 1.18947f
C56 VDD1.n3 B 1.78131f
C57 VTAIL.t2 B 0.149832f
C58 VTAIL.t5 B 0.149832f
C59 VTAIL.n0 B 1.23067f
C60 VTAIL.n1 B 0.328524f
C61 VTAIL.t7 B 1.56723f
C62 VTAIL.n2 B 0.457618f
C63 VTAIL.t6 B 0.149832f
C64 VTAIL.t9 B 0.149832f
C65 VTAIL.n3 B 1.23067f
C66 VTAIL.n4 B 1.33594f
C67 VTAIL.t0 B 0.149832f
C68 VTAIL.t1 B 0.149832f
C69 VTAIL.n5 B 1.23067f
C70 VTAIL.n6 B 1.33594f
C71 VTAIL.t4 B 1.56724f
C72 VTAIL.n7 B 0.457615f
C73 VTAIL.t8 B 0.149832f
C74 VTAIL.t10 B 0.149832f
C75 VTAIL.n8 B 1.23067f
C76 VTAIL.n9 B 0.385544f
C77 VTAIL.t11 B 1.56723f
C78 VTAIL.n10 B 1.32576f
C79 VTAIL.t3 B 1.56723f
C80 VTAIL.n11 B 1.30053f
C81 VP.n0 B 0.044036f
C82 VP.t4 B 0.772643f
C83 VP.n1 B 0.310301f
C84 VP.n2 B 0.044036f
C85 VP.n3 B 0.044036f
C86 VP.t2 B 0.831015f
C87 VP.t1 B 0.772643f
C88 VP.n4 B 0.350227f
C89 VP.t0 B 0.852136f
C90 VP.n5 B 0.361834f
C91 VP.n6 B 0.18178f
C92 VP.n7 B 0.055719f
C93 VP.n8 B 0.013679f
C94 VP.n9 B 0.352602f
C95 VP.n10 B 1.56382f
C96 VP.n11 B 1.60484f
C97 VP.t5 B 0.831015f
C98 VP.n12 B 0.352602f
C99 VP.n13 B 0.013679f
C100 VP.n14 B 0.055719f
C101 VP.n15 B 0.044036f
C102 VP.n16 B 0.044036f
C103 VP.n17 B 0.055719f
C104 VP.n18 B 0.013679f
C105 VP.t3 B 0.831015f
C106 VP.n19 B 0.352602f
C107 VP.n20 B 0.034126f
.ends

