* NGSPICE file created from diff_pair_sample_0650.ext - technology: sky130A

.subckt diff_pair_sample_0650 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1314_n4656# sky130_fd_pr__pfet_01v8 ad=7.1838 pd=37.62 as=0 ps=0 w=18.42 l=0.53
X1 VDD1.t1 VP.t0 VTAIL.t2 w_n1314_n4656# sky130_fd_pr__pfet_01v8 ad=7.1838 pd=37.62 as=7.1838 ps=37.62 w=18.42 l=0.53
X2 VDD1.t0 VP.t1 VTAIL.t3 w_n1314_n4656# sky130_fd_pr__pfet_01v8 ad=7.1838 pd=37.62 as=7.1838 ps=37.62 w=18.42 l=0.53
X3 B.t8 B.t6 B.t7 w_n1314_n4656# sky130_fd_pr__pfet_01v8 ad=7.1838 pd=37.62 as=0 ps=0 w=18.42 l=0.53
X4 B.t5 B.t3 B.t4 w_n1314_n4656# sky130_fd_pr__pfet_01v8 ad=7.1838 pd=37.62 as=0 ps=0 w=18.42 l=0.53
X5 VDD2.t1 VN.t0 VTAIL.t1 w_n1314_n4656# sky130_fd_pr__pfet_01v8 ad=7.1838 pd=37.62 as=7.1838 ps=37.62 w=18.42 l=0.53
X6 VDD2.t0 VN.t1 VTAIL.t0 w_n1314_n4656# sky130_fd_pr__pfet_01v8 ad=7.1838 pd=37.62 as=7.1838 ps=37.62 w=18.42 l=0.53
X7 B.t2 B.t0 B.t1 w_n1314_n4656# sky130_fd_pr__pfet_01v8 ad=7.1838 pd=37.62 as=0 ps=0 w=18.42 l=0.53
R0 B.n122 B.t9 1043.31
R1 B.n130 B.t0 1043.31
R2 B.n40 B.t6 1043.31
R3 B.n46 B.t3 1043.31
R4 B.n425 B.n424 585
R5 B.n426 B.n77 585
R6 B.n428 B.n427 585
R7 B.n429 B.n76 585
R8 B.n431 B.n430 585
R9 B.n432 B.n75 585
R10 B.n434 B.n433 585
R11 B.n435 B.n74 585
R12 B.n437 B.n436 585
R13 B.n438 B.n73 585
R14 B.n440 B.n439 585
R15 B.n441 B.n72 585
R16 B.n443 B.n442 585
R17 B.n444 B.n71 585
R18 B.n446 B.n445 585
R19 B.n447 B.n70 585
R20 B.n449 B.n448 585
R21 B.n450 B.n69 585
R22 B.n452 B.n451 585
R23 B.n453 B.n68 585
R24 B.n455 B.n454 585
R25 B.n456 B.n67 585
R26 B.n458 B.n457 585
R27 B.n459 B.n66 585
R28 B.n461 B.n460 585
R29 B.n462 B.n65 585
R30 B.n464 B.n463 585
R31 B.n465 B.n64 585
R32 B.n467 B.n466 585
R33 B.n468 B.n63 585
R34 B.n470 B.n469 585
R35 B.n471 B.n62 585
R36 B.n473 B.n472 585
R37 B.n474 B.n61 585
R38 B.n476 B.n475 585
R39 B.n477 B.n60 585
R40 B.n479 B.n478 585
R41 B.n480 B.n59 585
R42 B.n482 B.n481 585
R43 B.n483 B.n58 585
R44 B.n485 B.n484 585
R45 B.n486 B.n57 585
R46 B.n488 B.n487 585
R47 B.n489 B.n56 585
R48 B.n491 B.n490 585
R49 B.n492 B.n55 585
R50 B.n494 B.n493 585
R51 B.n495 B.n54 585
R52 B.n497 B.n496 585
R53 B.n498 B.n53 585
R54 B.n500 B.n499 585
R55 B.n501 B.n52 585
R56 B.n503 B.n502 585
R57 B.n504 B.n51 585
R58 B.n506 B.n505 585
R59 B.n507 B.n50 585
R60 B.n509 B.n508 585
R61 B.n510 B.n49 585
R62 B.n512 B.n511 585
R63 B.n513 B.n48 585
R64 B.n515 B.n514 585
R65 B.n517 B.n45 585
R66 B.n519 B.n518 585
R67 B.n520 B.n44 585
R68 B.n522 B.n521 585
R69 B.n523 B.n43 585
R70 B.n525 B.n524 585
R71 B.n526 B.n42 585
R72 B.n528 B.n527 585
R73 B.n529 B.n39 585
R74 B.n532 B.n531 585
R75 B.n533 B.n38 585
R76 B.n535 B.n534 585
R77 B.n536 B.n37 585
R78 B.n538 B.n537 585
R79 B.n539 B.n36 585
R80 B.n541 B.n540 585
R81 B.n542 B.n35 585
R82 B.n544 B.n543 585
R83 B.n545 B.n34 585
R84 B.n547 B.n546 585
R85 B.n548 B.n33 585
R86 B.n550 B.n549 585
R87 B.n551 B.n32 585
R88 B.n553 B.n552 585
R89 B.n554 B.n31 585
R90 B.n556 B.n555 585
R91 B.n557 B.n30 585
R92 B.n559 B.n558 585
R93 B.n560 B.n29 585
R94 B.n562 B.n561 585
R95 B.n563 B.n28 585
R96 B.n565 B.n564 585
R97 B.n566 B.n27 585
R98 B.n568 B.n567 585
R99 B.n569 B.n26 585
R100 B.n571 B.n570 585
R101 B.n572 B.n25 585
R102 B.n574 B.n573 585
R103 B.n575 B.n24 585
R104 B.n577 B.n576 585
R105 B.n578 B.n23 585
R106 B.n580 B.n579 585
R107 B.n581 B.n22 585
R108 B.n583 B.n582 585
R109 B.n584 B.n21 585
R110 B.n586 B.n585 585
R111 B.n587 B.n20 585
R112 B.n589 B.n588 585
R113 B.n590 B.n19 585
R114 B.n592 B.n591 585
R115 B.n593 B.n18 585
R116 B.n595 B.n594 585
R117 B.n596 B.n17 585
R118 B.n598 B.n597 585
R119 B.n599 B.n16 585
R120 B.n601 B.n600 585
R121 B.n602 B.n15 585
R122 B.n604 B.n603 585
R123 B.n605 B.n14 585
R124 B.n607 B.n606 585
R125 B.n608 B.n13 585
R126 B.n610 B.n609 585
R127 B.n611 B.n12 585
R128 B.n613 B.n612 585
R129 B.n614 B.n11 585
R130 B.n616 B.n615 585
R131 B.n617 B.n10 585
R132 B.n619 B.n618 585
R133 B.n620 B.n9 585
R134 B.n622 B.n621 585
R135 B.n423 B.n78 585
R136 B.n422 B.n421 585
R137 B.n420 B.n79 585
R138 B.n419 B.n418 585
R139 B.n417 B.n80 585
R140 B.n416 B.n415 585
R141 B.n414 B.n81 585
R142 B.n413 B.n412 585
R143 B.n411 B.n82 585
R144 B.n410 B.n409 585
R145 B.n408 B.n83 585
R146 B.n407 B.n406 585
R147 B.n405 B.n84 585
R148 B.n404 B.n403 585
R149 B.n402 B.n85 585
R150 B.n401 B.n400 585
R151 B.n399 B.n86 585
R152 B.n398 B.n397 585
R153 B.n396 B.n87 585
R154 B.n395 B.n394 585
R155 B.n393 B.n88 585
R156 B.n392 B.n391 585
R157 B.n390 B.n89 585
R158 B.n389 B.n388 585
R159 B.n387 B.n90 585
R160 B.n386 B.n385 585
R161 B.n384 B.n91 585
R162 B.n186 B.n161 585
R163 B.n188 B.n187 585
R164 B.n189 B.n160 585
R165 B.n191 B.n190 585
R166 B.n192 B.n159 585
R167 B.n194 B.n193 585
R168 B.n195 B.n158 585
R169 B.n197 B.n196 585
R170 B.n198 B.n157 585
R171 B.n200 B.n199 585
R172 B.n201 B.n156 585
R173 B.n203 B.n202 585
R174 B.n204 B.n155 585
R175 B.n206 B.n205 585
R176 B.n207 B.n154 585
R177 B.n209 B.n208 585
R178 B.n210 B.n153 585
R179 B.n212 B.n211 585
R180 B.n213 B.n152 585
R181 B.n215 B.n214 585
R182 B.n216 B.n151 585
R183 B.n218 B.n217 585
R184 B.n219 B.n150 585
R185 B.n221 B.n220 585
R186 B.n222 B.n149 585
R187 B.n224 B.n223 585
R188 B.n225 B.n148 585
R189 B.n227 B.n226 585
R190 B.n228 B.n147 585
R191 B.n230 B.n229 585
R192 B.n231 B.n146 585
R193 B.n233 B.n232 585
R194 B.n234 B.n145 585
R195 B.n236 B.n235 585
R196 B.n237 B.n144 585
R197 B.n239 B.n238 585
R198 B.n240 B.n143 585
R199 B.n242 B.n241 585
R200 B.n243 B.n142 585
R201 B.n245 B.n244 585
R202 B.n246 B.n141 585
R203 B.n248 B.n247 585
R204 B.n249 B.n140 585
R205 B.n251 B.n250 585
R206 B.n252 B.n139 585
R207 B.n254 B.n253 585
R208 B.n255 B.n138 585
R209 B.n257 B.n256 585
R210 B.n258 B.n137 585
R211 B.n260 B.n259 585
R212 B.n261 B.n136 585
R213 B.n263 B.n262 585
R214 B.n264 B.n135 585
R215 B.n266 B.n265 585
R216 B.n267 B.n134 585
R217 B.n269 B.n268 585
R218 B.n270 B.n133 585
R219 B.n272 B.n271 585
R220 B.n273 B.n132 585
R221 B.n275 B.n274 585
R222 B.n276 B.n129 585
R223 B.n279 B.n278 585
R224 B.n280 B.n128 585
R225 B.n282 B.n281 585
R226 B.n283 B.n127 585
R227 B.n285 B.n284 585
R228 B.n286 B.n126 585
R229 B.n288 B.n287 585
R230 B.n289 B.n125 585
R231 B.n291 B.n290 585
R232 B.n293 B.n292 585
R233 B.n294 B.n121 585
R234 B.n296 B.n295 585
R235 B.n297 B.n120 585
R236 B.n299 B.n298 585
R237 B.n300 B.n119 585
R238 B.n302 B.n301 585
R239 B.n303 B.n118 585
R240 B.n305 B.n304 585
R241 B.n306 B.n117 585
R242 B.n308 B.n307 585
R243 B.n309 B.n116 585
R244 B.n311 B.n310 585
R245 B.n312 B.n115 585
R246 B.n314 B.n313 585
R247 B.n315 B.n114 585
R248 B.n317 B.n316 585
R249 B.n318 B.n113 585
R250 B.n320 B.n319 585
R251 B.n321 B.n112 585
R252 B.n323 B.n322 585
R253 B.n324 B.n111 585
R254 B.n326 B.n325 585
R255 B.n327 B.n110 585
R256 B.n329 B.n328 585
R257 B.n330 B.n109 585
R258 B.n332 B.n331 585
R259 B.n333 B.n108 585
R260 B.n335 B.n334 585
R261 B.n336 B.n107 585
R262 B.n338 B.n337 585
R263 B.n339 B.n106 585
R264 B.n341 B.n340 585
R265 B.n342 B.n105 585
R266 B.n344 B.n343 585
R267 B.n345 B.n104 585
R268 B.n347 B.n346 585
R269 B.n348 B.n103 585
R270 B.n350 B.n349 585
R271 B.n351 B.n102 585
R272 B.n353 B.n352 585
R273 B.n354 B.n101 585
R274 B.n356 B.n355 585
R275 B.n357 B.n100 585
R276 B.n359 B.n358 585
R277 B.n360 B.n99 585
R278 B.n362 B.n361 585
R279 B.n363 B.n98 585
R280 B.n365 B.n364 585
R281 B.n366 B.n97 585
R282 B.n368 B.n367 585
R283 B.n369 B.n96 585
R284 B.n371 B.n370 585
R285 B.n372 B.n95 585
R286 B.n374 B.n373 585
R287 B.n375 B.n94 585
R288 B.n377 B.n376 585
R289 B.n378 B.n93 585
R290 B.n380 B.n379 585
R291 B.n381 B.n92 585
R292 B.n383 B.n382 585
R293 B.n185 B.n184 585
R294 B.n183 B.n162 585
R295 B.n182 B.n181 585
R296 B.n180 B.n163 585
R297 B.n179 B.n178 585
R298 B.n177 B.n164 585
R299 B.n176 B.n175 585
R300 B.n174 B.n165 585
R301 B.n173 B.n172 585
R302 B.n171 B.n166 585
R303 B.n170 B.n169 585
R304 B.n168 B.n167 585
R305 B.n2 B.n0 585
R306 B.n641 B.n1 585
R307 B.n640 B.n639 585
R308 B.n638 B.n3 585
R309 B.n637 B.n636 585
R310 B.n635 B.n4 585
R311 B.n634 B.n633 585
R312 B.n632 B.n5 585
R313 B.n631 B.n630 585
R314 B.n629 B.n6 585
R315 B.n628 B.n627 585
R316 B.n626 B.n7 585
R317 B.n625 B.n624 585
R318 B.n623 B.n8 585
R319 B.n643 B.n642 585
R320 B.n184 B.n161 502.111
R321 B.n623 B.n622 502.111
R322 B.n382 B.n91 502.111
R323 B.n424 B.n423 502.111
R324 B.n184 B.n183 163.367
R325 B.n183 B.n182 163.367
R326 B.n182 B.n163 163.367
R327 B.n178 B.n163 163.367
R328 B.n178 B.n177 163.367
R329 B.n177 B.n176 163.367
R330 B.n176 B.n165 163.367
R331 B.n172 B.n165 163.367
R332 B.n172 B.n171 163.367
R333 B.n171 B.n170 163.367
R334 B.n170 B.n167 163.367
R335 B.n167 B.n2 163.367
R336 B.n642 B.n2 163.367
R337 B.n642 B.n641 163.367
R338 B.n641 B.n640 163.367
R339 B.n640 B.n3 163.367
R340 B.n636 B.n3 163.367
R341 B.n636 B.n635 163.367
R342 B.n635 B.n634 163.367
R343 B.n634 B.n5 163.367
R344 B.n630 B.n5 163.367
R345 B.n630 B.n629 163.367
R346 B.n629 B.n628 163.367
R347 B.n628 B.n7 163.367
R348 B.n624 B.n7 163.367
R349 B.n624 B.n623 163.367
R350 B.n188 B.n161 163.367
R351 B.n189 B.n188 163.367
R352 B.n190 B.n189 163.367
R353 B.n190 B.n159 163.367
R354 B.n194 B.n159 163.367
R355 B.n195 B.n194 163.367
R356 B.n196 B.n195 163.367
R357 B.n196 B.n157 163.367
R358 B.n200 B.n157 163.367
R359 B.n201 B.n200 163.367
R360 B.n202 B.n201 163.367
R361 B.n202 B.n155 163.367
R362 B.n206 B.n155 163.367
R363 B.n207 B.n206 163.367
R364 B.n208 B.n207 163.367
R365 B.n208 B.n153 163.367
R366 B.n212 B.n153 163.367
R367 B.n213 B.n212 163.367
R368 B.n214 B.n213 163.367
R369 B.n214 B.n151 163.367
R370 B.n218 B.n151 163.367
R371 B.n219 B.n218 163.367
R372 B.n220 B.n219 163.367
R373 B.n220 B.n149 163.367
R374 B.n224 B.n149 163.367
R375 B.n225 B.n224 163.367
R376 B.n226 B.n225 163.367
R377 B.n226 B.n147 163.367
R378 B.n230 B.n147 163.367
R379 B.n231 B.n230 163.367
R380 B.n232 B.n231 163.367
R381 B.n232 B.n145 163.367
R382 B.n236 B.n145 163.367
R383 B.n237 B.n236 163.367
R384 B.n238 B.n237 163.367
R385 B.n238 B.n143 163.367
R386 B.n242 B.n143 163.367
R387 B.n243 B.n242 163.367
R388 B.n244 B.n243 163.367
R389 B.n244 B.n141 163.367
R390 B.n248 B.n141 163.367
R391 B.n249 B.n248 163.367
R392 B.n250 B.n249 163.367
R393 B.n250 B.n139 163.367
R394 B.n254 B.n139 163.367
R395 B.n255 B.n254 163.367
R396 B.n256 B.n255 163.367
R397 B.n256 B.n137 163.367
R398 B.n260 B.n137 163.367
R399 B.n261 B.n260 163.367
R400 B.n262 B.n261 163.367
R401 B.n262 B.n135 163.367
R402 B.n266 B.n135 163.367
R403 B.n267 B.n266 163.367
R404 B.n268 B.n267 163.367
R405 B.n268 B.n133 163.367
R406 B.n272 B.n133 163.367
R407 B.n273 B.n272 163.367
R408 B.n274 B.n273 163.367
R409 B.n274 B.n129 163.367
R410 B.n279 B.n129 163.367
R411 B.n280 B.n279 163.367
R412 B.n281 B.n280 163.367
R413 B.n281 B.n127 163.367
R414 B.n285 B.n127 163.367
R415 B.n286 B.n285 163.367
R416 B.n287 B.n286 163.367
R417 B.n287 B.n125 163.367
R418 B.n291 B.n125 163.367
R419 B.n292 B.n291 163.367
R420 B.n292 B.n121 163.367
R421 B.n296 B.n121 163.367
R422 B.n297 B.n296 163.367
R423 B.n298 B.n297 163.367
R424 B.n298 B.n119 163.367
R425 B.n302 B.n119 163.367
R426 B.n303 B.n302 163.367
R427 B.n304 B.n303 163.367
R428 B.n304 B.n117 163.367
R429 B.n308 B.n117 163.367
R430 B.n309 B.n308 163.367
R431 B.n310 B.n309 163.367
R432 B.n310 B.n115 163.367
R433 B.n314 B.n115 163.367
R434 B.n315 B.n314 163.367
R435 B.n316 B.n315 163.367
R436 B.n316 B.n113 163.367
R437 B.n320 B.n113 163.367
R438 B.n321 B.n320 163.367
R439 B.n322 B.n321 163.367
R440 B.n322 B.n111 163.367
R441 B.n326 B.n111 163.367
R442 B.n327 B.n326 163.367
R443 B.n328 B.n327 163.367
R444 B.n328 B.n109 163.367
R445 B.n332 B.n109 163.367
R446 B.n333 B.n332 163.367
R447 B.n334 B.n333 163.367
R448 B.n334 B.n107 163.367
R449 B.n338 B.n107 163.367
R450 B.n339 B.n338 163.367
R451 B.n340 B.n339 163.367
R452 B.n340 B.n105 163.367
R453 B.n344 B.n105 163.367
R454 B.n345 B.n344 163.367
R455 B.n346 B.n345 163.367
R456 B.n346 B.n103 163.367
R457 B.n350 B.n103 163.367
R458 B.n351 B.n350 163.367
R459 B.n352 B.n351 163.367
R460 B.n352 B.n101 163.367
R461 B.n356 B.n101 163.367
R462 B.n357 B.n356 163.367
R463 B.n358 B.n357 163.367
R464 B.n358 B.n99 163.367
R465 B.n362 B.n99 163.367
R466 B.n363 B.n362 163.367
R467 B.n364 B.n363 163.367
R468 B.n364 B.n97 163.367
R469 B.n368 B.n97 163.367
R470 B.n369 B.n368 163.367
R471 B.n370 B.n369 163.367
R472 B.n370 B.n95 163.367
R473 B.n374 B.n95 163.367
R474 B.n375 B.n374 163.367
R475 B.n376 B.n375 163.367
R476 B.n376 B.n93 163.367
R477 B.n380 B.n93 163.367
R478 B.n381 B.n380 163.367
R479 B.n382 B.n381 163.367
R480 B.n386 B.n91 163.367
R481 B.n387 B.n386 163.367
R482 B.n388 B.n387 163.367
R483 B.n388 B.n89 163.367
R484 B.n392 B.n89 163.367
R485 B.n393 B.n392 163.367
R486 B.n394 B.n393 163.367
R487 B.n394 B.n87 163.367
R488 B.n398 B.n87 163.367
R489 B.n399 B.n398 163.367
R490 B.n400 B.n399 163.367
R491 B.n400 B.n85 163.367
R492 B.n404 B.n85 163.367
R493 B.n405 B.n404 163.367
R494 B.n406 B.n405 163.367
R495 B.n406 B.n83 163.367
R496 B.n410 B.n83 163.367
R497 B.n411 B.n410 163.367
R498 B.n412 B.n411 163.367
R499 B.n412 B.n81 163.367
R500 B.n416 B.n81 163.367
R501 B.n417 B.n416 163.367
R502 B.n418 B.n417 163.367
R503 B.n418 B.n79 163.367
R504 B.n422 B.n79 163.367
R505 B.n423 B.n422 163.367
R506 B.n622 B.n9 163.367
R507 B.n618 B.n9 163.367
R508 B.n618 B.n617 163.367
R509 B.n617 B.n616 163.367
R510 B.n616 B.n11 163.367
R511 B.n612 B.n11 163.367
R512 B.n612 B.n611 163.367
R513 B.n611 B.n610 163.367
R514 B.n610 B.n13 163.367
R515 B.n606 B.n13 163.367
R516 B.n606 B.n605 163.367
R517 B.n605 B.n604 163.367
R518 B.n604 B.n15 163.367
R519 B.n600 B.n15 163.367
R520 B.n600 B.n599 163.367
R521 B.n599 B.n598 163.367
R522 B.n598 B.n17 163.367
R523 B.n594 B.n17 163.367
R524 B.n594 B.n593 163.367
R525 B.n593 B.n592 163.367
R526 B.n592 B.n19 163.367
R527 B.n588 B.n19 163.367
R528 B.n588 B.n587 163.367
R529 B.n587 B.n586 163.367
R530 B.n586 B.n21 163.367
R531 B.n582 B.n21 163.367
R532 B.n582 B.n581 163.367
R533 B.n581 B.n580 163.367
R534 B.n580 B.n23 163.367
R535 B.n576 B.n23 163.367
R536 B.n576 B.n575 163.367
R537 B.n575 B.n574 163.367
R538 B.n574 B.n25 163.367
R539 B.n570 B.n25 163.367
R540 B.n570 B.n569 163.367
R541 B.n569 B.n568 163.367
R542 B.n568 B.n27 163.367
R543 B.n564 B.n27 163.367
R544 B.n564 B.n563 163.367
R545 B.n563 B.n562 163.367
R546 B.n562 B.n29 163.367
R547 B.n558 B.n29 163.367
R548 B.n558 B.n557 163.367
R549 B.n557 B.n556 163.367
R550 B.n556 B.n31 163.367
R551 B.n552 B.n31 163.367
R552 B.n552 B.n551 163.367
R553 B.n551 B.n550 163.367
R554 B.n550 B.n33 163.367
R555 B.n546 B.n33 163.367
R556 B.n546 B.n545 163.367
R557 B.n545 B.n544 163.367
R558 B.n544 B.n35 163.367
R559 B.n540 B.n35 163.367
R560 B.n540 B.n539 163.367
R561 B.n539 B.n538 163.367
R562 B.n538 B.n37 163.367
R563 B.n534 B.n37 163.367
R564 B.n534 B.n533 163.367
R565 B.n533 B.n532 163.367
R566 B.n532 B.n39 163.367
R567 B.n527 B.n39 163.367
R568 B.n527 B.n526 163.367
R569 B.n526 B.n525 163.367
R570 B.n525 B.n43 163.367
R571 B.n521 B.n43 163.367
R572 B.n521 B.n520 163.367
R573 B.n520 B.n519 163.367
R574 B.n519 B.n45 163.367
R575 B.n514 B.n45 163.367
R576 B.n514 B.n513 163.367
R577 B.n513 B.n512 163.367
R578 B.n512 B.n49 163.367
R579 B.n508 B.n49 163.367
R580 B.n508 B.n507 163.367
R581 B.n507 B.n506 163.367
R582 B.n506 B.n51 163.367
R583 B.n502 B.n51 163.367
R584 B.n502 B.n501 163.367
R585 B.n501 B.n500 163.367
R586 B.n500 B.n53 163.367
R587 B.n496 B.n53 163.367
R588 B.n496 B.n495 163.367
R589 B.n495 B.n494 163.367
R590 B.n494 B.n55 163.367
R591 B.n490 B.n55 163.367
R592 B.n490 B.n489 163.367
R593 B.n489 B.n488 163.367
R594 B.n488 B.n57 163.367
R595 B.n484 B.n57 163.367
R596 B.n484 B.n483 163.367
R597 B.n483 B.n482 163.367
R598 B.n482 B.n59 163.367
R599 B.n478 B.n59 163.367
R600 B.n478 B.n477 163.367
R601 B.n477 B.n476 163.367
R602 B.n476 B.n61 163.367
R603 B.n472 B.n61 163.367
R604 B.n472 B.n471 163.367
R605 B.n471 B.n470 163.367
R606 B.n470 B.n63 163.367
R607 B.n466 B.n63 163.367
R608 B.n466 B.n465 163.367
R609 B.n465 B.n464 163.367
R610 B.n464 B.n65 163.367
R611 B.n460 B.n65 163.367
R612 B.n460 B.n459 163.367
R613 B.n459 B.n458 163.367
R614 B.n458 B.n67 163.367
R615 B.n454 B.n67 163.367
R616 B.n454 B.n453 163.367
R617 B.n453 B.n452 163.367
R618 B.n452 B.n69 163.367
R619 B.n448 B.n69 163.367
R620 B.n448 B.n447 163.367
R621 B.n447 B.n446 163.367
R622 B.n446 B.n71 163.367
R623 B.n442 B.n71 163.367
R624 B.n442 B.n441 163.367
R625 B.n441 B.n440 163.367
R626 B.n440 B.n73 163.367
R627 B.n436 B.n73 163.367
R628 B.n436 B.n435 163.367
R629 B.n435 B.n434 163.367
R630 B.n434 B.n75 163.367
R631 B.n430 B.n75 163.367
R632 B.n430 B.n429 163.367
R633 B.n429 B.n428 163.367
R634 B.n428 B.n77 163.367
R635 B.n424 B.n77 163.367
R636 B.n122 B.t11 124.005
R637 B.n46 B.t4 124.005
R638 B.n130 B.t2 123.983
R639 B.n40 B.t7 123.983
R640 B.n123 B.t10 107.328
R641 B.n47 B.t5 107.328
R642 B.n131 B.t1 107.303
R643 B.n41 B.t8 107.303
R644 B.n124 B.n123 59.5399
R645 B.n277 B.n131 59.5399
R646 B.n530 B.n41 59.5399
R647 B.n516 B.n47 59.5399
R648 B.n621 B.n8 32.6249
R649 B.n425 B.n78 32.6249
R650 B.n384 B.n383 32.6249
R651 B.n186 B.n185 32.6249
R652 B B.n643 18.0485
R653 B.n123 B.n122 16.6793
R654 B.n131 B.n130 16.6793
R655 B.n41 B.n40 16.6793
R656 B.n47 B.n46 16.6793
R657 B.n621 B.n620 10.6151
R658 B.n620 B.n619 10.6151
R659 B.n619 B.n10 10.6151
R660 B.n615 B.n10 10.6151
R661 B.n615 B.n614 10.6151
R662 B.n614 B.n613 10.6151
R663 B.n613 B.n12 10.6151
R664 B.n609 B.n12 10.6151
R665 B.n609 B.n608 10.6151
R666 B.n608 B.n607 10.6151
R667 B.n607 B.n14 10.6151
R668 B.n603 B.n14 10.6151
R669 B.n603 B.n602 10.6151
R670 B.n602 B.n601 10.6151
R671 B.n601 B.n16 10.6151
R672 B.n597 B.n16 10.6151
R673 B.n597 B.n596 10.6151
R674 B.n596 B.n595 10.6151
R675 B.n595 B.n18 10.6151
R676 B.n591 B.n18 10.6151
R677 B.n591 B.n590 10.6151
R678 B.n590 B.n589 10.6151
R679 B.n589 B.n20 10.6151
R680 B.n585 B.n20 10.6151
R681 B.n585 B.n584 10.6151
R682 B.n584 B.n583 10.6151
R683 B.n583 B.n22 10.6151
R684 B.n579 B.n22 10.6151
R685 B.n579 B.n578 10.6151
R686 B.n578 B.n577 10.6151
R687 B.n577 B.n24 10.6151
R688 B.n573 B.n24 10.6151
R689 B.n573 B.n572 10.6151
R690 B.n572 B.n571 10.6151
R691 B.n571 B.n26 10.6151
R692 B.n567 B.n26 10.6151
R693 B.n567 B.n566 10.6151
R694 B.n566 B.n565 10.6151
R695 B.n565 B.n28 10.6151
R696 B.n561 B.n28 10.6151
R697 B.n561 B.n560 10.6151
R698 B.n560 B.n559 10.6151
R699 B.n559 B.n30 10.6151
R700 B.n555 B.n30 10.6151
R701 B.n555 B.n554 10.6151
R702 B.n554 B.n553 10.6151
R703 B.n553 B.n32 10.6151
R704 B.n549 B.n32 10.6151
R705 B.n549 B.n548 10.6151
R706 B.n548 B.n547 10.6151
R707 B.n547 B.n34 10.6151
R708 B.n543 B.n34 10.6151
R709 B.n543 B.n542 10.6151
R710 B.n542 B.n541 10.6151
R711 B.n541 B.n36 10.6151
R712 B.n537 B.n36 10.6151
R713 B.n537 B.n536 10.6151
R714 B.n536 B.n535 10.6151
R715 B.n535 B.n38 10.6151
R716 B.n531 B.n38 10.6151
R717 B.n529 B.n528 10.6151
R718 B.n528 B.n42 10.6151
R719 B.n524 B.n42 10.6151
R720 B.n524 B.n523 10.6151
R721 B.n523 B.n522 10.6151
R722 B.n522 B.n44 10.6151
R723 B.n518 B.n44 10.6151
R724 B.n518 B.n517 10.6151
R725 B.n515 B.n48 10.6151
R726 B.n511 B.n48 10.6151
R727 B.n511 B.n510 10.6151
R728 B.n510 B.n509 10.6151
R729 B.n509 B.n50 10.6151
R730 B.n505 B.n50 10.6151
R731 B.n505 B.n504 10.6151
R732 B.n504 B.n503 10.6151
R733 B.n503 B.n52 10.6151
R734 B.n499 B.n52 10.6151
R735 B.n499 B.n498 10.6151
R736 B.n498 B.n497 10.6151
R737 B.n497 B.n54 10.6151
R738 B.n493 B.n54 10.6151
R739 B.n493 B.n492 10.6151
R740 B.n492 B.n491 10.6151
R741 B.n491 B.n56 10.6151
R742 B.n487 B.n56 10.6151
R743 B.n487 B.n486 10.6151
R744 B.n486 B.n485 10.6151
R745 B.n485 B.n58 10.6151
R746 B.n481 B.n58 10.6151
R747 B.n481 B.n480 10.6151
R748 B.n480 B.n479 10.6151
R749 B.n479 B.n60 10.6151
R750 B.n475 B.n60 10.6151
R751 B.n475 B.n474 10.6151
R752 B.n474 B.n473 10.6151
R753 B.n473 B.n62 10.6151
R754 B.n469 B.n62 10.6151
R755 B.n469 B.n468 10.6151
R756 B.n468 B.n467 10.6151
R757 B.n467 B.n64 10.6151
R758 B.n463 B.n64 10.6151
R759 B.n463 B.n462 10.6151
R760 B.n462 B.n461 10.6151
R761 B.n461 B.n66 10.6151
R762 B.n457 B.n66 10.6151
R763 B.n457 B.n456 10.6151
R764 B.n456 B.n455 10.6151
R765 B.n455 B.n68 10.6151
R766 B.n451 B.n68 10.6151
R767 B.n451 B.n450 10.6151
R768 B.n450 B.n449 10.6151
R769 B.n449 B.n70 10.6151
R770 B.n445 B.n70 10.6151
R771 B.n445 B.n444 10.6151
R772 B.n444 B.n443 10.6151
R773 B.n443 B.n72 10.6151
R774 B.n439 B.n72 10.6151
R775 B.n439 B.n438 10.6151
R776 B.n438 B.n437 10.6151
R777 B.n437 B.n74 10.6151
R778 B.n433 B.n74 10.6151
R779 B.n433 B.n432 10.6151
R780 B.n432 B.n431 10.6151
R781 B.n431 B.n76 10.6151
R782 B.n427 B.n76 10.6151
R783 B.n427 B.n426 10.6151
R784 B.n426 B.n425 10.6151
R785 B.n385 B.n384 10.6151
R786 B.n385 B.n90 10.6151
R787 B.n389 B.n90 10.6151
R788 B.n390 B.n389 10.6151
R789 B.n391 B.n390 10.6151
R790 B.n391 B.n88 10.6151
R791 B.n395 B.n88 10.6151
R792 B.n396 B.n395 10.6151
R793 B.n397 B.n396 10.6151
R794 B.n397 B.n86 10.6151
R795 B.n401 B.n86 10.6151
R796 B.n402 B.n401 10.6151
R797 B.n403 B.n402 10.6151
R798 B.n403 B.n84 10.6151
R799 B.n407 B.n84 10.6151
R800 B.n408 B.n407 10.6151
R801 B.n409 B.n408 10.6151
R802 B.n409 B.n82 10.6151
R803 B.n413 B.n82 10.6151
R804 B.n414 B.n413 10.6151
R805 B.n415 B.n414 10.6151
R806 B.n415 B.n80 10.6151
R807 B.n419 B.n80 10.6151
R808 B.n420 B.n419 10.6151
R809 B.n421 B.n420 10.6151
R810 B.n421 B.n78 10.6151
R811 B.n187 B.n186 10.6151
R812 B.n187 B.n160 10.6151
R813 B.n191 B.n160 10.6151
R814 B.n192 B.n191 10.6151
R815 B.n193 B.n192 10.6151
R816 B.n193 B.n158 10.6151
R817 B.n197 B.n158 10.6151
R818 B.n198 B.n197 10.6151
R819 B.n199 B.n198 10.6151
R820 B.n199 B.n156 10.6151
R821 B.n203 B.n156 10.6151
R822 B.n204 B.n203 10.6151
R823 B.n205 B.n204 10.6151
R824 B.n205 B.n154 10.6151
R825 B.n209 B.n154 10.6151
R826 B.n210 B.n209 10.6151
R827 B.n211 B.n210 10.6151
R828 B.n211 B.n152 10.6151
R829 B.n215 B.n152 10.6151
R830 B.n216 B.n215 10.6151
R831 B.n217 B.n216 10.6151
R832 B.n217 B.n150 10.6151
R833 B.n221 B.n150 10.6151
R834 B.n222 B.n221 10.6151
R835 B.n223 B.n222 10.6151
R836 B.n223 B.n148 10.6151
R837 B.n227 B.n148 10.6151
R838 B.n228 B.n227 10.6151
R839 B.n229 B.n228 10.6151
R840 B.n229 B.n146 10.6151
R841 B.n233 B.n146 10.6151
R842 B.n234 B.n233 10.6151
R843 B.n235 B.n234 10.6151
R844 B.n235 B.n144 10.6151
R845 B.n239 B.n144 10.6151
R846 B.n240 B.n239 10.6151
R847 B.n241 B.n240 10.6151
R848 B.n241 B.n142 10.6151
R849 B.n245 B.n142 10.6151
R850 B.n246 B.n245 10.6151
R851 B.n247 B.n246 10.6151
R852 B.n247 B.n140 10.6151
R853 B.n251 B.n140 10.6151
R854 B.n252 B.n251 10.6151
R855 B.n253 B.n252 10.6151
R856 B.n253 B.n138 10.6151
R857 B.n257 B.n138 10.6151
R858 B.n258 B.n257 10.6151
R859 B.n259 B.n258 10.6151
R860 B.n259 B.n136 10.6151
R861 B.n263 B.n136 10.6151
R862 B.n264 B.n263 10.6151
R863 B.n265 B.n264 10.6151
R864 B.n265 B.n134 10.6151
R865 B.n269 B.n134 10.6151
R866 B.n270 B.n269 10.6151
R867 B.n271 B.n270 10.6151
R868 B.n271 B.n132 10.6151
R869 B.n275 B.n132 10.6151
R870 B.n276 B.n275 10.6151
R871 B.n278 B.n128 10.6151
R872 B.n282 B.n128 10.6151
R873 B.n283 B.n282 10.6151
R874 B.n284 B.n283 10.6151
R875 B.n284 B.n126 10.6151
R876 B.n288 B.n126 10.6151
R877 B.n289 B.n288 10.6151
R878 B.n290 B.n289 10.6151
R879 B.n294 B.n293 10.6151
R880 B.n295 B.n294 10.6151
R881 B.n295 B.n120 10.6151
R882 B.n299 B.n120 10.6151
R883 B.n300 B.n299 10.6151
R884 B.n301 B.n300 10.6151
R885 B.n301 B.n118 10.6151
R886 B.n305 B.n118 10.6151
R887 B.n306 B.n305 10.6151
R888 B.n307 B.n306 10.6151
R889 B.n307 B.n116 10.6151
R890 B.n311 B.n116 10.6151
R891 B.n312 B.n311 10.6151
R892 B.n313 B.n312 10.6151
R893 B.n313 B.n114 10.6151
R894 B.n317 B.n114 10.6151
R895 B.n318 B.n317 10.6151
R896 B.n319 B.n318 10.6151
R897 B.n319 B.n112 10.6151
R898 B.n323 B.n112 10.6151
R899 B.n324 B.n323 10.6151
R900 B.n325 B.n324 10.6151
R901 B.n325 B.n110 10.6151
R902 B.n329 B.n110 10.6151
R903 B.n330 B.n329 10.6151
R904 B.n331 B.n330 10.6151
R905 B.n331 B.n108 10.6151
R906 B.n335 B.n108 10.6151
R907 B.n336 B.n335 10.6151
R908 B.n337 B.n336 10.6151
R909 B.n337 B.n106 10.6151
R910 B.n341 B.n106 10.6151
R911 B.n342 B.n341 10.6151
R912 B.n343 B.n342 10.6151
R913 B.n343 B.n104 10.6151
R914 B.n347 B.n104 10.6151
R915 B.n348 B.n347 10.6151
R916 B.n349 B.n348 10.6151
R917 B.n349 B.n102 10.6151
R918 B.n353 B.n102 10.6151
R919 B.n354 B.n353 10.6151
R920 B.n355 B.n354 10.6151
R921 B.n355 B.n100 10.6151
R922 B.n359 B.n100 10.6151
R923 B.n360 B.n359 10.6151
R924 B.n361 B.n360 10.6151
R925 B.n361 B.n98 10.6151
R926 B.n365 B.n98 10.6151
R927 B.n366 B.n365 10.6151
R928 B.n367 B.n366 10.6151
R929 B.n367 B.n96 10.6151
R930 B.n371 B.n96 10.6151
R931 B.n372 B.n371 10.6151
R932 B.n373 B.n372 10.6151
R933 B.n373 B.n94 10.6151
R934 B.n377 B.n94 10.6151
R935 B.n378 B.n377 10.6151
R936 B.n379 B.n378 10.6151
R937 B.n379 B.n92 10.6151
R938 B.n383 B.n92 10.6151
R939 B.n185 B.n162 10.6151
R940 B.n181 B.n162 10.6151
R941 B.n181 B.n180 10.6151
R942 B.n180 B.n179 10.6151
R943 B.n179 B.n164 10.6151
R944 B.n175 B.n164 10.6151
R945 B.n175 B.n174 10.6151
R946 B.n174 B.n173 10.6151
R947 B.n173 B.n166 10.6151
R948 B.n169 B.n166 10.6151
R949 B.n169 B.n168 10.6151
R950 B.n168 B.n0 10.6151
R951 B.n639 B.n1 10.6151
R952 B.n639 B.n638 10.6151
R953 B.n638 B.n637 10.6151
R954 B.n637 B.n4 10.6151
R955 B.n633 B.n4 10.6151
R956 B.n633 B.n632 10.6151
R957 B.n632 B.n631 10.6151
R958 B.n631 B.n6 10.6151
R959 B.n627 B.n6 10.6151
R960 B.n627 B.n626 10.6151
R961 B.n626 B.n625 10.6151
R962 B.n625 B.n8 10.6151
R963 B.n530 B.n529 7.18099
R964 B.n517 B.n516 7.18099
R965 B.n278 B.n277 7.18099
R966 B.n290 B.n124 7.18099
R967 B.n531 B.n530 3.43465
R968 B.n516 B.n515 3.43465
R969 B.n277 B.n276 3.43465
R970 B.n293 B.n124 3.43465
R971 B.n643 B.n0 2.81026
R972 B.n643 B.n1 2.81026
R973 VP.n0 VP.t1 1117.96
R974 VP.n0 VP.t0 1073.92
R975 VP VP.n0 0.0516364
R976 VTAIL.n1 VTAIL.t0 56.7865
R977 VTAIL.n3 VTAIL.t1 56.7855
R978 VTAIL.n0 VTAIL.t2 56.7855
R979 VTAIL.n2 VTAIL.t3 56.7854
R980 VTAIL.n1 VTAIL.n0 29.7462
R981 VTAIL.n3 VTAIL.n2 29.0048
R982 VTAIL.n2 VTAIL.n1 0.841017
R983 VTAIL VTAIL.n0 0.713862
R984 VTAIL VTAIL.n3 0.127655
R985 VDD1 VDD1.t1 115.213
R986 VDD1 VDD1.t0 73.7077
R987 VN VN.t1 1118.34
R988 VN VN.t0 1073.97
R989 VDD2.n0 VDD2.t1 114.504
R990 VDD2.n0 VDD2.t0 73.4642
R991 VDD2 VDD2.n0 0.244034
C0 VTAIL w_n1314_n4656# 4.04994f
C1 B w_n1314_n4656# 8.3757f
C2 VP VDD1 2.72095f
C3 VDD2 VDD1 0.448327f
C4 VN w_n1314_n4656# 1.76542f
C5 VTAIL VDD1 8.61253f
C6 VP VDD2 0.24866f
C7 VDD1 B 1.84471f
C8 VP VTAIL 1.81183f
C9 VTAIL VDD2 8.64055f
C10 VP B 1.03084f
C11 VDD2 B 1.85807f
C12 VN VDD1 0.148178f
C13 VTAIL B 3.76611f
C14 VN VP 5.67578f
C15 VN VDD2 2.62751f
C16 VDD1 w_n1314_n4656# 2.03195f
C17 VN VTAIL 1.79687f
C18 VP w_n1314_n4656# 1.92834f
C19 VN B 0.771309f
C20 VDD2 w_n1314_n4656# 2.03489f
C21 VDD2 VSUBS 0.963842f
C22 VDD1 VSUBS 5.53753f
C23 VTAIL VSUBS 0.261859f
C24 VN VSUBS 7.10172f
C25 VP VSUBS 1.30056f
C26 B VSUBS 2.915124f
C27 w_n1314_n4656# VSUBS 74.787605f
C28 VDD2.t1 VSUBS 4.79114f
C29 VDD2.t0 VSUBS 3.9891f
C30 VDD2.n0 VSUBS 4.3692f
C31 VN.t0 VSUBS 1.44869f
C32 VN.t1 VSUBS 1.55507f
C33 VDD1.t0 VSUBS 3.99315f
C34 VDD1.t1 VSUBS 4.82468f
C35 VTAIL.t2 VSUBS 3.78809f
C36 VTAIL.n0 VSUBS 2.48149f
C37 VTAIL.t0 VSUBS 3.78809f
C38 VTAIL.n1 VSUBS 2.49171f
C39 VTAIL.t3 VSUBS 3.78808f
C40 VTAIL.n2 VSUBS 2.43212f
C41 VTAIL.t1 VSUBS 3.78809f
C42 VTAIL.n3 VSUBS 2.37475f
C43 VP.t1 VSUBS 1.58493f
C44 VP.t0 VSUBS 1.47853f
C45 VP.n0 VSUBS 5.32421f
C46 B.n0 VSUBS 0.004463f
C47 B.n1 VSUBS 0.004463f
C48 B.n2 VSUBS 0.007058f
C49 B.n3 VSUBS 0.007058f
C50 B.n4 VSUBS 0.007058f
C51 B.n5 VSUBS 0.007058f
C52 B.n6 VSUBS 0.007058f
C53 B.n7 VSUBS 0.007058f
C54 B.n8 VSUBS 0.015882f
C55 B.n9 VSUBS 0.007058f
C56 B.n10 VSUBS 0.007058f
C57 B.n11 VSUBS 0.007058f
C58 B.n12 VSUBS 0.007058f
C59 B.n13 VSUBS 0.007058f
C60 B.n14 VSUBS 0.007058f
C61 B.n15 VSUBS 0.007058f
C62 B.n16 VSUBS 0.007058f
C63 B.n17 VSUBS 0.007058f
C64 B.n18 VSUBS 0.007058f
C65 B.n19 VSUBS 0.007058f
C66 B.n20 VSUBS 0.007058f
C67 B.n21 VSUBS 0.007058f
C68 B.n22 VSUBS 0.007058f
C69 B.n23 VSUBS 0.007058f
C70 B.n24 VSUBS 0.007058f
C71 B.n25 VSUBS 0.007058f
C72 B.n26 VSUBS 0.007058f
C73 B.n27 VSUBS 0.007058f
C74 B.n28 VSUBS 0.007058f
C75 B.n29 VSUBS 0.007058f
C76 B.n30 VSUBS 0.007058f
C77 B.n31 VSUBS 0.007058f
C78 B.n32 VSUBS 0.007058f
C79 B.n33 VSUBS 0.007058f
C80 B.n34 VSUBS 0.007058f
C81 B.n35 VSUBS 0.007058f
C82 B.n36 VSUBS 0.007058f
C83 B.n37 VSUBS 0.007058f
C84 B.n38 VSUBS 0.007058f
C85 B.n39 VSUBS 0.007058f
C86 B.t8 VSUBS 0.627973f
C87 B.t7 VSUBS 0.635243f
C88 B.t6 VSUBS 0.390459f
C89 B.n40 VSUBS 0.163297f
C90 B.n41 VSUBS 0.064106f
C91 B.n42 VSUBS 0.007058f
C92 B.n43 VSUBS 0.007058f
C93 B.n44 VSUBS 0.007058f
C94 B.n45 VSUBS 0.007058f
C95 B.t5 VSUBS 0.627948f
C96 B.t4 VSUBS 0.63522f
C97 B.t3 VSUBS 0.390459f
C98 B.n46 VSUBS 0.16332f
C99 B.n47 VSUBS 0.06413f
C100 B.n48 VSUBS 0.007058f
C101 B.n49 VSUBS 0.007058f
C102 B.n50 VSUBS 0.007058f
C103 B.n51 VSUBS 0.007058f
C104 B.n52 VSUBS 0.007058f
C105 B.n53 VSUBS 0.007058f
C106 B.n54 VSUBS 0.007058f
C107 B.n55 VSUBS 0.007058f
C108 B.n56 VSUBS 0.007058f
C109 B.n57 VSUBS 0.007058f
C110 B.n58 VSUBS 0.007058f
C111 B.n59 VSUBS 0.007058f
C112 B.n60 VSUBS 0.007058f
C113 B.n61 VSUBS 0.007058f
C114 B.n62 VSUBS 0.007058f
C115 B.n63 VSUBS 0.007058f
C116 B.n64 VSUBS 0.007058f
C117 B.n65 VSUBS 0.007058f
C118 B.n66 VSUBS 0.007058f
C119 B.n67 VSUBS 0.007058f
C120 B.n68 VSUBS 0.007058f
C121 B.n69 VSUBS 0.007058f
C122 B.n70 VSUBS 0.007058f
C123 B.n71 VSUBS 0.007058f
C124 B.n72 VSUBS 0.007058f
C125 B.n73 VSUBS 0.007058f
C126 B.n74 VSUBS 0.007058f
C127 B.n75 VSUBS 0.007058f
C128 B.n76 VSUBS 0.007058f
C129 B.n77 VSUBS 0.007058f
C130 B.n78 VSUBS 0.016717f
C131 B.n79 VSUBS 0.007058f
C132 B.n80 VSUBS 0.007058f
C133 B.n81 VSUBS 0.007058f
C134 B.n82 VSUBS 0.007058f
C135 B.n83 VSUBS 0.007058f
C136 B.n84 VSUBS 0.007058f
C137 B.n85 VSUBS 0.007058f
C138 B.n86 VSUBS 0.007058f
C139 B.n87 VSUBS 0.007058f
C140 B.n88 VSUBS 0.007058f
C141 B.n89 VSUBS 0.007058f
C142 B.n90 VSUBS 0.007058f
C143 B.n91 VSUBS 0.015882f
C144 B.n92 VSUBS 0.007058f
C145 B.n93 VSUBS 0.007058f
C146 B.n94 VSUBS 0.007058f
C147 B.n95 VSUBS 0.007058f
C148 B.n96 VSUBS 0.007058f
C149 B.n97 VSUBS 0.007058f
C150 B.n98 VSUBS 0.007058f
C151 B.n99 VSUBS 0.007058f
C152 B.n100 VSUBS 0.007058f
C153 B.n101 VSUBS 0.007058f
C154 B.n102 VSUBS 0.007058f
C155 B.n103 VSUBS 0.007058f
C156 B.n104 VSUBS 0.007058f
C157 B.n105 VSUBS 0.007058f
C158 B.n106 VSUBS 0.007058f
C159 B.n107 VSUBS 0.007058f
C160 B.n108 VSUBS 0.007058f
C161 B.n109 VSUBS 0.007058f
C162 B.n110 VSUBS 0.007058f
C163 B.n111 VSUBS 0.007058f
C164 B.n112 VSUBS 0.007058f
C165 B.n113 VSUBS 0.007058f
C166 B.n114 VSUBS 0.007058f
C167 B.n115 VSUBS 0.007058f
C168 B.n116 VSUBS 0.007058f
C169 B.n117 VSUBS 0.007058f
C170 B.n118 VSUBS 0.007058f
C171 B.n119 VSUBS 0.007058f
C172 B.n120 VSUBS 0.007058f
C173 B.n121 VSUBS 0.007058f
C174 B.t10 VSUBS 0.627948f
C175 B.t11 VSUBS 0.63522f
C176 B.t9 VSUBS 0.390459f
C177 B.n122 VSUBS 0.16332f
C178 B.n123 VSUBS 0.06413f
C179 B.n124 VSUBS 0.016353f
C180 B.n125 VSUBS 0.007058f
C181 B.n126 VSUBS 0.007058f
C182 B.n127 VSUBS 0.007058f
C183 B.n128 VSUBS 0.007058f
C184 B.n129 VSUBS 0.007058f
C185 B.t1 VSUBS 0.627973f
C186 B.t2 VSUBS 0.635243f
C187 B.t0 VSUBS 0.390459f
C188 B.n130 VSUBS 0.163297f
C189 B.n131 VSUBS 0.064106f
C190 B.n132 VSUBS 0.007058f
C191 B.n133 VSUBS 0.007058f
C192 B.n134 VSUBS 0.007058f
C193 B.n135 VSUBS 0.007058f
C194 B.n136 VSUBS 0.007058f
C195 B.n137 VSUBS 0.007058f
C196 B.n138 VSUBS 0.007058f
C197 B.n139 VSUBS 0.007058f
C198 B.n140 VSUBS 0.007058f
C199 B.n141 VSUBS 0.007058f
C200 B.n142 VSUBS 0.007058f
C201 B.n143 VSUBS 0.007058f
C202 B.n144 VSUBS 0.007058f
C203 B.n145 VSUBS 0.007058f
C204 B.n146 VSUBS 0.007058f
C205 B.n147 VSUBS 0.007058f
C206 B.n148 VSUBS 0.007058f
C207 B.n149 VSUBS 0.007058f
C208 B.n150 VSUBS 0.007058f
C209 B.n151 VSUBS 0.007058f
C210 B.n152 VSUBS 0.007058f
C211 B.n153 VSUBS 0.007058f
C212 B.n154 VSUBS 0.007058f
C213 B.n155 VSUBS 0.007058f
C214 B.n156 VSUBS 0.007058f
C215 B.n157 VSUBS 0.007058f
C216 B.n158 VSUBS 0.007058f
C217 B.n159 VSUBS 0.007058f
C218 B.n160 VSUBS 0.007058f
C219 B.n161 VSUBS 0.017124f
C220 B.n162 VSUBS 0.007058f
C221 B.n163 VSUBS 0.007058f
C222 B.n164 VSUBS 0.007058f
C223 B.n165 VSUBS 0.007058f
C224 B.n166 VSUBS 0.007058f
C225 B.n167 VSUBS 0.007058f
C226 B.n168 VSUBS 0.007058f
C227 B.n169 VSUBS 0.007058f
C228 B.n170 VSUBS 0.007058f
C229 B.n171 VSUBS 0.007058f
C230 B.n172 VSUBS 0.007058f
C231 B.n173 VSUBS 0.007058f
C232 B.n174 VSUBS 0.007058f
C233 B.n175 VSUBS 0.007058f
C234 B.n176 VSUBS 0.007058f
C235 B.n177 VSUBS 0.007058f
C236 B.n178 VSUBS 0.007058f
C237 B.n179 VSUBS 0.007058f
C238 B.n180 VSUBS 0.007058f
C239 B.n181 VSUBS 0.007058f
C240 B.n182 VSUBS 0.007058f
C241 B.n183 VSUBS 0.007058f
C242 B.n184 VSUBS 0.015882f
C243 B.n185 VSUBS 0.015882f
C244 B.n186 VSUBS 0.017124f
C245 B.n187 VSUBS 0.007058f
C246 B.n188 VSUBS 0.007058f
C247 B.n189 VSUBS 0.007058f
C248 B.n190 VSUBS 0.007058f
C249 B.n191 VSUBS 0.007058f
C250 B.n192 VSUBS 0.007058f
C251 B.n193 VSUBS 0.007058f
C252 B.n194 VSUBS 0.007058f
C253 B.n195 VSUBS 0.007058f
C254 B.n196 VSUBS 0.007058f
C255 B.n197 VSUBS 0.007058f
C256 B.n198 VSUBS 0.007058f
C257 B.n199 VSUBS 0.007058f
C258 B.n200 VSUBS 0.007058f
C259 B.n201 VSUBS 0.007058f
C260 B.n202 VSUBS 0.007058f
C261 B.n203 VSUBS 0.007058f
C262 B.n204 VSUBS 0.007058f
C263 B.n205 VSUBS 0.007058f
C264 B.n206 VSUBS 0.007058f
C265 B.n207 VSUBS 0.007058f
C266 B.n208 VSUBS 0.007058f
C267 B.n209 VSUBS 0.007058f
C268 B.n210 VSUBS 0.007058f
C269 B.n211 VSUBS 0.007058f
C270 B.n212 VSUBS 0.007058f
C271 B.n213 VSUBS 0.007058f
C272 B.n214 VSUBS 0.007058f
C273 B.n215 VSUBS 0.007058f
C274 B.n216 VSUBS 0.007058f
C275 B.n217 VSUBS 0.007058f
C276 B.n218 VSUBS 0.007058f
C277 B.n219 VSUBS 0.007058f
C278 B.n220 VSUBS 0.007058f
C279 B.n221 VSUBS 0.007058f
C280 B.n222 VSUBS 0.007058f
C281 B.n223 VSUBS 0.007058f
C282 B.n224 VSUBS 0.007058f
C283 B.n225 VSUBS 0.007058f
C284 B.n226 VSUBS 0.007058f
C285 B.n227 VSUBS 0.007058f
C286 B.n228 VSUBS 0.007058f
C287 B.n229 VSUBS 0.007058f
C288 B.n230 VSUBS 0.007058f
C289 B.n231 VSUBS 0.007058f
C290 B.n232 VSUBS 0.007058f
C291 B.n233 VSUBS 0.007058f
C292 B.n234 VSUBS 0.007058f
C293 B.n235 VSUBS 0.007058f
C294 B.n236 VSUBS 0.007058f
C295 B.n237 VSUBS 0.007058f
C296 B.n238 VSUBS 0.007058f
C297 B.n239 VSUBS 0.007058f
C298 B.n240 VSUBS 0.007058f
C299 B.n241 VSUBS 0.007058f
C300 B.n242 VSUBS 0.007058f
C301 B.n243 VSUBS 0.007058f
C302 B.n244 VSUBS 0.007058f
C303 B.n245 VSUBS 0.007058f
C304 B.n246 VSUBS 0.007058f
C305 B.n247 VSUBS 0.007058f
C306 B.n248 VSUBS 0.007058f
C307 B.n249 VSUBS 0.007058f
C308 B.n250 VSUBS 0.007058f
C309 B.n251 VSUBS 0.007058f
C310 B.n252 VSUBS 0.007058f
C311 B.n253 VSUBS 0.007058f
C312 B.n254 VSUBS 0.007058f
C313 B.n255 VSUBS 0.007058f
C314 B.n256 VSUBS 0.007058f
C315 B.n257 VSUBS 0.007058f
C316 B.n258 VSUBS 0.007058f
C317 B.n259 VSUBS 0.007058f
C318 B.n260 VSUBS 0.007058f
C319 B.n261 VSUBS 0.007058f
C320 B.n262 VSUBS 0.007058f
C321 B.n263 VSUBS 0.007058f
C322 B.n264 VSUBS 0.007058f
C323 B.n265 VSUBS 0.007058f
C324 B.n266 VSUBS 0.007058f
C325 B.n267 VSUBS 0.007058f
C326 B.n268 VSUBS 0.007058f
C327 B.n269 VSUBS 0.007058f
C328 B.n270 VSUBS 0.007058f
C329 B.n271 VSUBS 0.007058f
C330 B.n272 VSUBS 0.007058f
C331 B.n273 VSUBS 0.007058f
C332 B.n274 VSUBS 0.007058f
C333 B.n275 VSUBS 0.007058f
C334 B.n276 VSUBS 0.004671f
C335 B.n277 VSUBS 0.016353f
C336 B.n278 VSUBS 0.005916f
C337 B.n279 VSUBS 0.007058f
C338 B.n280 VSUBS 0.007058f
C339 B.n281 VSUBS 0.007058f
C340 B.n282 VSUBS 0.007058f
C341 B.n283 VSUBS 0.007058f
C342 B.n284 VSUBS 0.007058f
C343 B.n285 VSUBS 0.007058f
C344 B.n286 VSUBS 0.007058f
C345 B.n287 VSUBS 0.007058f
C346 B.n288 VSUBS 0.007058f
C347 B.n289 VSUBS 0.007058f
C348 B.n290 VSUBS 0.005916f
C349 B.n291 VSUBS 0.007058f
C350 B.n292 VSUBS 0.007058f
C351 B.n293 VSUBS 0.004671f
C352 B.n294 VSUBS 0.007058f
C353 B.n295 VSUBS 0.007058f
C354 B.n296 VSUBS 0.007058f
C355 B.n297 VSUBS 0.007058f
C356 B.n298 VSUBS 0.007058f
C357 B.n299 VSUBS 0.007058f
C358 B.n300 VSUBS 0.007058f
C359 B.n301 VSUBS 0.007058f
C360 B.n302 VSUBS 0.007058f
C361 B.n303 VSUBS 0.007058f
C362 B.n304 VSUBS 0.007058f
C363 B.n305 VSUBS 0.007058f
C364 B.n306 VSUBS 0.007058f
C365 B.n307 VSUBS 0.007058f
C366 B.n308 VSUBS 0.007058f
C367 B.n309 VSUBS 0.007058f
C368 B.n310 VSUBS 0.007058f
C369 B.n311 VSUBS 0.007058f
C370 B.n312 VSUBS 0.007058f
C371 B.n313 VSUBS 0.007058f
C372 B.n314 VSUBS 0.007058f
C373 B.n315 VSUBS 0.007058f
C374 B.n316 VSUBS 0.007058f
C375 B.n317 VSUBS 0.007058f
C376 B.n318 VSUBS 0.007058f
C377 B.n319 VSUBS 0.007058f
C378 B.n320 VSUBS 0.007058f
C379 B.n321 VSUBS 0.007058f
C380 B.n322 VSUBS 0.007058f
C381 B.n323 VSUBS 0.007058f
C382 B.n324 VSUBS 0.007058f
C383 B.n325 VSUBS 0.007058f
C384 B.n326 VSUBS 0.007058f
C385 B.n327 VSUBS 0.007058f
C386 B.n328 VSUBS 0.007058f
C387 B.n329 VSUBS 0.007058f
C388 B.n330 VSUBS 0.007058f
C389 B.n331 VSUBS 0.007058f
C390 B.n332 VSUBS 0.007058f
C391 B.n333 VSUBS 0.007058f
C392 B.n334 VSUBS 0.007058f
C393 B.n335 VSUBS 0.007058f
C394 B.n336 VSUBS 0.007058f
C395 B.n337 VSUBS 0.007058f
C396 B.n338 VSUBS 0.007058f
C397 B.n339 VSUBS 0.007058f
C398 B.n340 VSUBS 0.007058f
C399 B.n341 VSUBS 0.007058f
C400 B.n342 VSUBS 0.007058f
C401 B.n343 VSUBS 0.007058f
C402 B.n344 VSUBS 0.007058f
C403 B.n345 VSUBS 0.007058f
C404 B.n346 VSUBS 0.007058f
C405 B.n347 VSUBS 0.007058f
C406 B.n348 VSUBS 0.007058f
C407 B.n349 VSUBS 0.007058f
C408 B.n350 VSUBS 0.007058f
C409 B.n351 VSUBS 0.007058f
C410 B.n352 VSUBS 0.007058f
C411 B.n353 VSUBS 0.007058f
C412 B.n354 VSUBS 0.007058f
C413 B.n355 VSUBS 0.007058f
C414 B.n356 VSUBS 0.007058f
C415 B.n357 VSUBS 0.007058f
C416 B.n358 VSUBS 0.007058f
C417 B.n359 VSUBS 0.007058f
C418 B.n360 VSUBS 0.007058f
C419 B.n361 VSUBS 0.007058f
C420 B.n362 VSUBS 0.007058f
C421 B.n363 VSUBS 0.007058f
C422 B.n364 VSUBS 0.007058f
C423 B.n365 VSUBS 0.007058f
C424 B.n366 VSUBS 0.007058f
C425 B.n367 VSUBS 0.007058f
C426 B.n368 VSUBS 0.007058f
C427 B.n369 VSUBS 0.007058f
C428 B.n370 VSUBS 0.007058f
C429 B.n371 VSUBS 0.007058f
C430 B.n372 VSUBS 0.007058f
C431 B.n373 VSUBS 0.007058f
C432 B.n374 VSUBS 0.007058f
C433 B.n375 VSUBS 0.007058f
C434 B.n376 VSUBS 0.007058f
C435 B.n377 VSUBS 0.007058f
C436 B.n378 VSUBS 0.007058f
C437 B.n379 VSUBS 0.007058f
C438 B.n380 VSUBS 0.007058f
C439 B.n381 VSUBS 0.007058f
C440 B.n382 VSUBS 0.017124f
C441 B.n383 VSUBS 0.017124f
C442 B.n384 VSUBS 0.015882f
C443 B.n385 VSUBS 0.007058f
C444 B.n386 VSUBS 0.007058f
C445 B.n387 VSUBS 0.007058f
C446 B.n388 VSUBS 0.007058f
C447 B.n389 VSUBS 0.007058f
C448 B.n390 VSUBS 0.007058f
C449 B.n391 VSUBS 0.007058f
C450 B.n392 VSUBS 0.007058f
C451 B.n393 VSUBS 0.007058f
C452 B.n394 VSUBS 0.007058f
C453 B.n395 VSUBS 0.007058f
C454 B.n396 VSUBS 0.007058f
C455 B.n397 VSUBS 0.007058f
C456 B.n398 VSUBS 0.007058f
C457 B.n399 VSUBS 0.007058f
C458 B.n400 VSUBS 0.007058f
C459 B.n401 VSUBS 0.007058f
C460 B.n402 VSUBS 0.007058f
C461 B.n403 VSUBS 0.007058f
C462 B.n404 VSUBS 0.007058f
C463 B.n405 VSUBS 0.007058f
C464 B.n406 VSUBS 0.007058f
C465 B.n407 VSUBS 0.007058f
C466 B.n408 VSUBS 0.007058f
C467 B.n409 VSUBS 0.007058f
C468 B.n410 VSUBS 0.007058f
C469 B.n411 VSUBS 0.007058f
C470 B.n412 VSUBS 0.007058f
C471 B.n413 VSUBS 0.007058f
C472 B.n414 VSUBS 0.007058f
C473 B.n415 VSUBS 0.007058f
C474 B.n416 VSUBS 0.007058f
C475 B.n417 VSUBS 0.007058f
C476 B.n418 VSUBS 0.007058f
C477 B.n419 VSUBS 0.007058f
C478 B.n420 VSUBS 0.007058f
C479 B.n421 VSUBS 0.007058f
C480 B.n422 VSUBS 0.007058f
C481 B.n423 VSUBS 0.015882f
C482 B.n424 VSUBS 0.017124f
C483 B.n425 VSUBS 0.016289f
C484 B.n426 VSUBS 0.007058f
C485 B.n427 VSUBS 0.007058f
C486 B.n428 VSUBS 0.007058f
C487 B.n429 VSUBS 0.007058f
C488 B.n430 VSUBS 0.007058f
C489 B.n431 VSUBS 0.007058f
C490 B.n432 VSUBS 0.007058f
C491 B.n433 VSUBS 0.007058f
C492 B.n434 VSUBS 0.007058f
C493 B.n435 VSUBS 0.007058f
C494 B.n436 VSUBS 0.007058f
C495 B.n437 VSUBS 0.007058f
C496 B.n438 VSUBS 0.007058f
C497 B.n439 VSUBS 0.007058f
C498 B.n440 VSUBS 0.007058f
C499 B.n441 VSUBS 0.007058f
C500 B.n442 VSUBS 0.007058f
C501 B.n443 VSUBS 0.007058f
C502 B.n444 VSUBS 0.007058f
C503 B.n445 VSUBS 0.007058f
C504 B.n446 VSUBS 0.007058f
C505 B.n447 VSUBS 0.007058f
C506 B.n448 VSUBS 0.007058f
C507 B.n449 VSUBS 0.007058f
C508 B.n450 VSUBS 0.007058f
C509 B.n451 VSUBS 0.007058f
C510 B.n452 VSUBS 0.007058f
C511 B.n453 VSUBS 0.007058f
C512 B.n454 VSUBS 0.007058f
C513 B.n455 VSUBS 0.007058f
C514 B.n456 VSUBS 0.007058f
C515 B.n457 VSUBS 0.007058f
C516 B.n458 VSUBS 0.007058f
C517 B.n459 VSUBS 0.007058f
C518 B.n460 VSUBS 0.007058f
C519 B.n461 VSUBS 0.007058f
C520 B.n462 VSUBS 0.007058f
C521 B.n463 VSUBS 0.007058f
C522 B.n464 VSUBS 0.007058f
C523 B.n465 VSUBS 0.007058f
C524 B.n466 VSUBS 0.007058f
C525 B.n467 VSUBS 0.007058f
C526 B.n468 VSUBS 0.007058f
C527 B.n469 VSUBS 0.007058f
C528 B.n470 VSUBS 0.007058f
C529 B.n471 VSUBS 0.007058f
C530 B.n472 VSUBS 0.007058f
C531 B.n473 VSUBS 0.007058f
C532 B.n474 VSUBS 0.007058f
C533 B.n475 VSUBS 0.007058f
C534 B.n476 VSUBS 0.007058f
C535 B.n477 VSUBS 0.007058f
C536 B.n478 VSUBS 0.007058f
C537 B.n479 VSUBS 0.007058f
C538 B.n480 VSUBS 0.007058f
C539 B.n481 VSUBS 0.007058f
C540 B.n482 VSUBS 0.007058f
C541 B.n483 VSUBS 0.007058f
C542 B.n484 VSUBS 0.007058f
C543 B.n485 VSUBS 0.007058f
C544 B.n486 VSUBS 0.007058f
C545 B.n487 VSUBS 0.007058f
C546 B.n488 VSUBS 0.007058f
C547 B.n489 VSUBS 0.007058f
C548 B.n490 VSUBS 0.007058f
C549 B.n491 VSUBS 0.007058f
C550 B.n492 VSUBS 0.007058f
C551 B.n493 VSUBS 0.007058f
C552 B.n494 VSUBS 0.007058f
C553 B.n495 VSUBS 0.007058f
C554 B.n496 VSUBS 0.007058f
C555 B.n497 VSUBS 0.007058f
C556 B.n498 VSUBS 0.007058f
C557 B.n499 VSUBS 0.007058f
C558 B.n500 VSUBS 0.007058f
C559 B.n501 VSUBS 0.007058f
C560 B.n502 VSUBS 0.007058f
C561 B.n503 VSUBS 0.007058f
C562 B.n504 VSUBS 0.007058f
C563 B.n505 VSUBS 0.007058f
C564 B.n506 VSUBS 0.007058f
C565 B.n507 VSUBS 0.007058f
C566 B.n508 VSUBS 0.007058f
C567 B.n509 VSUBS 0.007058f
C568 B.n510 VSUBS 0.007058f
C569 B.n511 VSUBS 0.007058f
C570 B.n512 VSUBS 0.007058f
C571 B.n513 VSUBS 0.007058f
C572 B.n514 VSUBS 0.007058f
C573 B.n515 VSUBS 0.004671f
C574 B.n516 VSUBS 0.016353f
C575 B.n517 VSUBS 0.005916f
C576 B.n518 VSUBS 0.007058f
C577 B.n519 VSUBS 0.007058f
C578 B.n520 VSUBS 0.007058f
C579 B.n521 VSUBS 0.007058f
C580 B.n522 VSUBS 0.007058f
C581 B.n523 VSUBS 0.007058f
C582 B.n524 VSUBS 0.007058f
C583 B.n525 VSUBS 0.007058f
C584 B.n526 VSUBS 0.007058f
C585 B.n527 VSUBS 0.007058f
C586 B.n528 VSUBS 0.007058f
C587 B.n529 VSUBS 0.005916f
C588 B.n530 VSUBS 0.016353f
C589 B.n531 VSUBS 0.004671f
C590 B.n532 VSUBS 0.007058f
C591 B.n533 VSUBS 0.007058f
C592 B.n534 VSUBS 0.007058f
C593 B.n535 VSUBS 0.007058f
C594 B.n536 VSUBS 0.007058f
C595 B.n537 VSUBS 0.007058f
C596 B.n538 VSUBS 0.007058f
C597 B.n539 VSUBS 0.007058f
C598 B.n540 VSUBS 0.007058f
C599 B.n541 VSUBS 0.007058f
C600 B.n542 VSUBS 0.007058f
C601 B.n543 VSUBS 0.007058f
C602 B.n544 VSUBS 0.007058f
C603 B.n545 VSUBS 0.007058f
C604 B.n546 VSUBS 0.007058f
C605 B.n547 VSUBS 0.007058f
C606 B.n548 VSUBS 0.007058f
C607 B.n549 VSUBS 0.007058f
C608 B.n550 VSUBS 0.007058f
C609 B.n551 VSUBS 0.007058f
C610 B.n552 VSUBS 0.007058f
C611 B.n553 VSUBS 0.007058f
C612 B.n554 VSUBS 0.007058f
C613 B.n555 VSUBS 0.007058f
C614 B.n556 VSUBS 0.007058f
C615 B.n557 VSUBS 0.007058f
C616 B.n558 VSUBS 0.007058f
C617 B.n559 VSUBS 0.007058f
C618 B.n560 VSUBS 0.007058f
C619 B.n561 VSUBS 0.007058f
C620 B.n562 VSUBS 0.007058f
C621 B.n563 VSUBS 0.007058f
C622 B.n564 VSUBS 0.007058f
C623 B.n565 VSUBS 0.007058f
C624 B.n566 VSUBS 0.007058f
C625 B.n567 VSUBS 0.007058f
C626 B.n568 VSUBS 0.007058f
C627 B.n569 VSUBS 0.007058f
C628 B.n570 VSUBS 0.007058f
C629 B.n571 VSUBS 0.007058f
C630 B.n572 VSUBS 0.007058f
C631 B.n573 VSUBS 0.007058f
C632 B.n574 VSUBS 0.007058f
C633 B.n575 VSUBS 0.007058f
C634 B.n576 VSUBS 0.007058f
C635 B.n577 VSUBS 0.007058f
C636 B.n578 VSUBS 0.007058f
C637 B.n579 VSUBS 0.007058f
C638 B.n580 VSUBS 0.007058f
C639 B.n581 VSUBS 0.007058f
C640 B.n582 VSUBS 0.007058f
C641 B.n583 VSUBS 0.007058f
C642 B.n584 VSUBS 0.007058f
C643 B.n585 VSUBS 0.007058f
C644 B.n586 VSUBS 0.007058f
C645 B.n587 VSUBS 0.007058f
C646 B.n588 VSUBS 0.007058f
C647 B.n589 VSUBS 0.007058f
C648 B.n590 VSUBS 0.007058f
C649 B.n591 VSUBS 0.007058f
C650 B.n592 VSUBS 0.007058f
C651 B.n593 VSUBS 0.007058f
C652 B.n594 VSUBS 0.007058f
C653 B.n595 VSUBS 0.007058f
C654 B.n596 VSUBS 0.007058f
C655 B.n597 VSUBS 0.007058f
C656 B.n598 VSUBS 0.007058f
C657 B.n599 VSUBS 0.007058f
C658 B.n600 VSUBS 0.007058f
C659 B.n601 VSUBS 0.007058f
C660 B.n602 VSUBS 0.007058f
C661 B.n603 VSUBS 0.007058f
C662 B.n604 VSUBS 0.007058f
C663 B.n605 VSUBS 0.007058f
C664 B.n606 VSUBS 0.007058f
C665 B.n607 VSUBS 0.007058f
C666 B.n608 VSUBS 0.007058f
C667 B.n609 VSUBS 0.007058f
C668 B.n610 VSUBS 0.007058f
C669 B.n611 VSUBS 0.007058f
C670 B.n612 VSUBS 0.007058f
C671 B.n613 VSUBS 0.007058f
C672 B.n614 VSUBS 0.007058f
C673 B.n615 VSUBS 0.007058f
C674 B.n616 VSUBS 0.007058f
C675 B.n617 VSUBS 0.007058f
C676 B.n618 VSUBS 0.007058f
C677 B.n619 VSUBS 0.007058f
C678 B.n620 VSUBS 0.007058f
C679 B.n621 VSUBS 0.017124f
C680 B.n622 VSUBS 0.017124f
C681 B.n623 VSUBS 0.015882f
C682 B.n624 VSUBS 0.007058f
C683 B.n625 VSUBS 0.007058f
C684 B.n626 VSUBS 0.007058f
C685 B.n627 VSUBS 0.007058f
C686 B.n628 VSUBS 0.007058f
C687 B.n629 VSUBS 0.007058f
C688 B.n630 VSUBS 0.007058f
C689 B.n631 VSUBS 0.007058f
C690 B.n632 VSUBS 0.007058f
C691 B.n633 VSUBS 0.007058f
C692 B.n634 VSUBS 0.007058f
C693 B.n635 VSUBS 0.007058f
C694 B.n636 VSUBS 0.007058f
C695 B.n637 VSUBS 0.007058f
C696 B.n638 VSUBS 0.007058f
C697 B.n639 VSUBS 0.007058f
C698 B.n640 VSUBS 0.007058f
C699 B.n641 VSUBS 0.007058f
C700 B.n642 VSUBS 0.007058f
C701 B.n643 VSUBS 0.015982f
.ends

