* NGSPICE file created from diff_pair_sample_1743.ext - technology: sky130A

.subckt diff_pair_sample_1743 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.4446 pd=3.06 as=0 ps=0 w=1.14 l=3.04
X1 VTAIL.t15 VP.t0 VDD1.t2 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.1881 ps=1.47 w=1.14 l=3.04
X2 VTAIL.t6 VN.t0 VDD2.t7 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.4446 pd=3.06 as=0.1881 ps=1.47 w=1.14 l=3.04
X3 VTAIL.t5 VN.t1 VDD2.t6 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.4446 pd=3.06 as=0.1881 ps=1.47 w=1.14 l=3.04
X4 VDD1.t7 VP.t1 VTAIL.t14 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.1881 ps=1.47 w=1.14 l=3.04
X5 VDD1.t4 VP.t2 VTAIL.t13 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.1881 ps=1.47 w=1.14 l=3.04
X6 VDD2.t5 VN.t2 VTAIL.t2 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.4446 ps=3.06 w=1.14 l=3.04
X7 VTAIL.t4 VN.t3 VDD2.t4 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.1881 ps=1.47 w=1.14 l=3.04
X8 VDD1.t0 VP.t3 VTAIL.t12 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.4446 ps=3.06 w=1.14 l=3.04
X9 VDD1.t6 VP.t4 VTAIL.t11 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.4446 ps=3.06 w=1.14 l=3.04
X10 VDD2.t3 VN.t4 VTAIL.t3 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.1881 ps=1.47 w=1.14 l=3.04
X11 VTAIL.t10 VP.t5 VDD1.t5 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.1881 ps=1.47 w=1.14 l=3.04
X12 B.t8 B.t6 B.t7 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.4446 pd=3.06 as=0 ps=0 w=1.14 l=3.04
X13 B.t5 B.t3 B.t4 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.4446 pd=3.06 as=0 ps=0 w=1.14 l=3.04
X14 B.t2 B.t0 B.t1 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.4446 pd=3.06 as=0 ps=0 w=1.14 l=3.04
X15 VTAIL.t7 VN.t5 VDD2.t2 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.1881 ps=1.47 w=1.14 l=3.04
X16 VDD2.t1 VN.t6 VTAIL.t1 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.4446 ps=3.06 w=1.14 l=3.04
X17 VTAIL.t9 VP.t6 VDD1.t1 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.4446 pd=3.06 as=0.1881 ps=1.47 w=1.14 l=3.04
X18 VTAIL.t8 VP.t7 VDD1.t3 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.4446 pd=3.06 as=0.1881 ps=1.47 w=1.14 l=3.04
X19 VDD2.t0 VN.t7 VTAIL.t0 w_n4340_n1196# sky130_fd_pr__pfet_01v8 ad=0.1881 pd=1.47 as=0.1881 ps=1.47 w=1.14 l=3.04
R0 B.n283 B.n282 585
R1 B.n281 B.n108 585
R2 B.n280 B.n279 585
R3 B.n278 B.n109 585
R4 B.n277 B.n276 585
R5 B.n275 B.n110 585
R6 B.n274 B.n273 585
R7 B.n272 B.n111 585
R8 B.n271 B.n270 585
R9 B.n269 B.n112 585
R10 B.n268 B.n267 585
R11 B.n263 B.n113 585
R12 B.n262 B.n261 585
R13 B.n260 B.n114 585
R14 B.n259 B.n258 585
R15 B.n257 B.n115 585
R16 B.n256 B.n255 585
R17 B.n254 B.n116 585
R18 B.n253 B.n252 585
R19 B.n250 B.n117 585
R20 B.n249 B.n248 585
R21 B.n247 B.n120 585
R22 B.n246 B.n245 585
R23 B.n244 B.n121 585
R24 B.n243 B.n242 585
R25 B.n241 B.n122 585
R26 B.n240 B.n239 585
R27 B.n238 B.n123 585
R28 B.n237 B.n236 585
R29 B.n284 B.n107 585
R30 B.n286 B.n285 585
R31 B.n287 B.n106 585
R32 B.n289 B.n288 585
R33 B.n290 B.n105 585
R34 B.n292 B.n291 585
R35 B.n293 B.n104 585
R36 B.n295 B.n294 585
R37 B.n296 B.n103 585
R38 B.n298 B.n297 585
R39 B.n299 B.n102 585
R40 B.n301 B.n300 585
R41 B.n302 B.n101 585
R42 B.n304 B.n303 585
R43 B.n305 B.n100 585
R44 B.n307 B.n306 585
R45 B.n308 B.n99 585
R46 B.n310 B.n309 585
R47 B.n311 B.n98 585
R48 B.n313 B.n312 585
R49 B.n314 B.n97 585
R50 B.n316 B.n315 585
R51 B.n317 B.n96 585
R52 B.n319 B.n318 585
R53 B.n320 B.n95 585
R54 B.n322 B.n321 585
R55 B.n323 B.n94 585
R56 B.n325 B.n324 585
R57 B.n326 B.n93 585
R58 B.n328 B.n327 585
R59 B.n329 B.n92 585
R60 B.n331 B.n330 585
R61 B.n332 B.n91 585
R62 B.n334 B.n333 585
R63 B.n335 B.n90 585
R64 B.n337 B.n336 585
R65 B.n338 B.n89 585
R66 B.n340 B.n339 585
R67 B.n341 B.n88 585
R68 B.n343 B.n342 585
R69 B.n344 B.n87 585
R70 B.n346 B.n345 585
R71 B.n347 B.n86 585
R72 B.n349 B.n348 585
R73 B.n350 B.n85 585
R74 B.n352 B.n351 585
R75 B.n353 B.n84 585
R76 B.n355 B.n354 585
R77 B.n356 B.n83 585
R78 B.n358 B.n357 585
R79 B.n359 B.n82 585
R80 B.n361 B.n360 585
R81 B.n362 B.n81 585
R82 B.n364 B.n363 585
R83 B.n365 B.n80 585
R84 B.n367 B.n366 585
R85 B.n368 B.n79 585
R86 B.n370 B.n369 585
R87 B.n371 B.n78 585
R88 B.n373 B.n372 585
R89 B.n374 B.n77 585
R90 B.n376 B.n375 585
R91 B.n377 B.n76 585
R92 B.n379 B.n378 585
R93 B.n380 B.n75 585
R94 B.n382 B.n381 585
R95 B.n383 B.n74 585
R96 B.n385 B.n384 585
R97 B.n386 B.n73 585
R98 B.n388 B.n387 585
R99 B.n389 B.n72 585
R100 B.n391 B.n390 585
R101 B.n392 B.n71 585
R102 B.n394 B.n393 585
R103 B.n395 B.n70 585
R104 B.n397 B.n396 585
R105 B.n398 B.n69 585
R106 B.n400 B.n399 585
R107 B.n401 B.n68 585
R108 B.n403 B.n402 585
R109 B.n404 B.n67 585
R110 B.n406 B.n405 585
R111 B.n407 B.n66 585
R112 B.n409 B.n408 585
R113 B.n410 B.n65 585
R114 B.n412 B.n411 585
R115 B.n413 B.n64 585
R116 B.n415 B.n414 585
R117 B.n416 B.n63 585
R118 B.n418 B.n417 585
R119 B.n419 B.n62 585
R120 B.n421 B.n420 585
R121 B.n422 B.n61 585
R122 B.n424 B.n423 585
R123 B.n425 B.n60 585
R124 B.n427 B.n426 585
R125 B.n428 B.n59 585
R126 B.n430 B.n429 585
R127 B.n431 B.n58 585
R128 B.n433 B.n432 585
R129 B.n434 B.n57 585
R130 B.n436 B.n435 585
R131 B.n437 B.n56 585
R132 B.n439 B.n438 585
R133 B.n440 B.n55 585
R134 B.n442 B.n441 585
R135 B.n443 B.n54 585
R136 B.n445 B.n444 585
R137 B.n446 B.n53 585
R138 B.n448 B.n447 585
R139 B.n449 B.n52 585
R140 B.n451 B.n450 585
R141 B.n452 B.n51 585
R142 B.n454 B.n453 585
R143 B.n455 B.n50 585
R144 B.n457 B.n456 585
R145 B.n502 B.n501 585
R146 B.n500 B.n31 585
R147 B.n499 B.n498 585
R148 B.n497 B.n32 585
R149 B.n496 B.n495 585
R150 B.n494 B.n33 585
R151 B.n493 B.n492 585
R152 B.n491 B.n34 585
R153 B.n490 B.n489 585
R154 B.n488 B.n35 585
R155 B.n486 B.n485 585
R156 B.n484 B.n38 585
R157 B.n483 B.n482 585
R158 B.n481 B.n39 585
R159 B.n480 B.n479 585
R160 B.n478 B.n40 585
R161 B.n477 B.n476 585
R162 B.n475 B.n41 585
R163 B.n474 B.n473 585
R164 B.n472 B.n471 585
R165 B.n470 B.n45 585
R166 B.n469 B.n468 585
R167 B.n467 B.n46 585
R168 B.n466 B.n465 585
R169 B.n464 B.n47 585
R170 B.n463 B.n462 585
R171 B.n461 B.n48 585
R172 B.n460 B.n459 585
R173 B.n458 B.n49 585
R174 B.n503 B.n30 585
R175 B.n505 B.n504 585
R176 B.n506 B.n29 585
R177 B.n508 B.n507 585
R178 B.n509 B.n28 585
R179 B.n511 B.n510 585
R180 B.n512 B.n27 585
R181 B.n514 B.n513 585
R182 B.n515 B.n26 585
R183 B.n517 B.n516 585
R184 B.n518 B.n25 585
R185 B.n520 B.n519 585
R186 B.n521 B.n24 585
R187 B.n523 B.n522 585
R188 B.n524 B.n23 585
R189 B.n526 B.n525 585
R190 B.n527 B.n22 585
R191 B.n529 B.n528 585
R192 B.n530 B.n21 585
R193 B.n532 B.n531 585
R194 B.n533 B.n20 585
R195 B.n535 B.n534 585
R196 B.n536 B.n19 585
R197 B.n538 B.n537 585
R198 B.n539 B.n18 585
R199 B.n541 B.n540 585
R200 B.n542 B.n17 585
R201 B.n544 B.n543 585
R202 B.n545 B.n16 585
R203 B.n547 B.n546 585
R204 B.n548 B.n15 585
R205 B.n550 B.n549 585
R206 B.n551 B.n14 585
R207 B.n553 B.n552 585
R208 B.n554 B.n13 585
R209 B.n556 B.n555 585
R210 B.n557 B.n12 585
R211 B.n559 B.n558 585
R212 B.n560 B.n11 585
R213 B.n562 B.n561 585
R214 B.n563 B.n10 585
R215 B.n565 B.n564 585
R216 B.n566 B.n9 585
R217 B.n568 B.n567 585
R218 B.n569 B.n8 585
R219 B.n571 B.n570 585
R220 B.n572 B.n7 585
R221 B.n574 B.n573 585
R222 B.n575 B.n6 585
R223 B.n577 B.n576 585
R224 B.n578 B.n5 585
R225 B.n580 B.n579 585
R226 B.n581 B.n4 585
R227 B.n583 B.n582 585
R228 B.n584 B.n3 585
R229 B.n586 B.n585 585
R230 B.n587 B.n0 585
R231 B.n2 B.n1 585
R232 B.n153 B.n152 585
R233 B.n154 B.n151 585
R234 B.n156 B.n155 585
R235 B.n157 B.n150 585
R236 B.n159 B.n158 585
R237 B.n160 B.n149 585
R238 B.n162 B.n161 585
R239 B.n163 B.n148 585
R240 B.n165 B.n164 585
R241 B.n166 B.n147 585
R242 B.n168 B.n167 585
R243 B.n169 B.n146 585
R244 B.n171 B.n170 585
R245 B.n172 B.n145 585
R246 B.n174 B.n173 585
R247 B.n175 B.n144 585
R248 B.n177 B.n176 585
R249 B.n178 B.n143 585
R250 B.n180 B.n179 585
R251 B.n181 B.n142 585
R252 B.n183 B.n182 585
R253 B.n184 B.n141 585
R254 B.n186 B.n185 585
R255 B.n187 B.n140 585
R256 B.n189 B.n188 585
R257 B.n190 B.n139 585
R258 B.n192 B.n191 585
R259 B.n193 B.n138 585
R260 B.n195 B.n194 585
R261 B.n196 B.n137 585
R262 B.n198 B.n197 585
R263 B.n199 B.n136 585
R264 B.n201 B.n200 585
R265 B.n202 B.n135 585
R266 B.n204 B.n203 585
R267 B.n205 B.n134 585
R268 B.n207 B.n206 585
R269 B.n208 B.n133 585
R270 B.n210 B.n209 585
R271 B.n211 B.n132 585
R272 B.n213 B.n212 585
R273 B.n214 B.n131 585
R274 B.n216 B.n215 585
R275 B.n217 B.n130 585
R276 B.n219 B.n218 585
R277 B.n220 B.n129 585
R278 B.n222 B.n221 585
R279 B.n223 B.n128 585
R280 B.n225 B.n224 585
R281 B.n226 B.n127 585
R282 B.n228 B.n227 585
R283 B.n229 B.n126 585
R284 B.n231 B.n230 585
R285 B.n232 B.n125 585
R286 B.n234 B.n233 585
R287 B.n235 B.n124 585
R288 B.n236 B.n235 521.33
R289 B.n282 B.n107 521.33
R290 B.n456 B.n49 521.33
R291 B.n503 B.n502 521.33
R292 B.n118 B.t10 429.272
R293 B.n264 B.t4 429.272
R294 B.n42 B.t2 429.272
R295 B.n36 B.t8 429.272
R296 B.n119 B.t11 363.914
R297 B.n265 B.t5 363.914
R298 B.n43 B.t1 363.914
R299 B.n37 B.t7 363.914
R300 B.n589 B.n588 256.663
R301 B.n588 B.n587 235.042
R302 B.n588 B.n2 235.042
R303 B.n118 B.t9 209.327
R304 B.n264 B.t3 209.327
R305 B.n42 B.t0 209.327
R306 B.n36 B.t6 209.327
R307 B.n236 B.n123 163.367
R308 B.n240 B.n123 163.367
R309 B.n241 B.n240 163.367
R310 B.n242 B.n241 163.367
R311 B.n242 B.n121 163.367
R312 B.n246 B.n121 163.367
R313 B.n247 B.n246 163.367
R314 B.n248 B.n247 163.367
R315 B.n248 B.n117 163.367
R316 B.n253 B.n117 163.367
R317 B.n254 B.n253 163.367
R318 B.n255 B.n254 163.367
R319 B.n255 B.n115 163.367
R320 B.n259 B.n115 163.367
R321 B.n260 B.n259 163.367
R322 B.n261 B.n260 163.367
R323 B.n261 B.n113 163.367
R324 B.n268 B.n113 163.367
R325 B.n269 B.n268 163.367
R326 B.n270 B.n269 163.367
R327 B.n270 B.n111 163.367
R328 B.n274 B.n111 163.367
R329 B.n275 B.n274 163.367
R330 B.n276 B.n275 163.367
R331 B.n276 B.n109 163.367
R332 B.n280 B.n109 163.367
R333 B.n281 B.n280 163.367
R334 B.n282 B.n281 163.367
R335 B.n456 B.n455 163.367
R336 B.n455 B.n454 163.367
R337 B.n454 B.n51 163.367
R338 B.n450 B.n51 163.367
R339 B.n450 B.n449 163.367
R340 B.n449 B.n448 163.367
R341 B.n448 B.n53 163.367
R342 B.n444 B.n53 163.367
R343 B.n444 B.n443 163.367
R344 B.n443 B.n442 163.367
R345 B.n442 B.n55 163.367
R346 B.n438 B.n55 163.367
R347 B.n438 B.n437 163.367
R348 B.n437 B.n436 163.367
R349 B.n436 B.n57 163.367
R350 B.n432 B.n57 163.367
R351 B.n432 B.n431 163.367
R352 B.n431 B.n430 163.367
R353 B.n430 B.n59 163.367
R354 B.n426 B.n59 163.367
R355 B.n426 B.n425 163.367
R356 B.n425 B.n424 163.367
R357 B.n424 B.n61 163.367
R358 B.n420 B.n61 163.367
R359 B.n420 B.n419 163.367
R360 B.n419 B.n418 163.367
R361 B.n418 B.n63 163.367
R362 B.n414 B.n63 163.367
R363 B.n414 B.n413 163.367
R364 B.n413 B.n412 163.367
R365 B.n412 B.n65 163.367
R366 B.n408 B.n65 163.367
R367 B.n408 B.n407 163.367
R368 B.n407 B.n406 163.367
R369 B.n406 B.n67 163.367
R370 B.n402 B.n67 163.367
R371 B.n402 B.n401 163.367
R372 B.n401 B.n400 163.367
R373 B.n400 B.n69 163.367
R374 B.n396 B.n69 163.367
R375 B.n396 B.n395 163.367
R376 B.n395 B.n394 163.367
R377 B.n394 B.n71 163.367
R378 B.n390 B.n71 163.367
R379 B.n390 B.n389 163.367
R380 B.n389 B.n388 163.367
R381 B.n388 B.n73 163.367
R382 B.n384 B.n73 163.367
R383 B.n384 B.n383 163.367
R384 B.n383 B.n382 163.367
R385 B.n382 B.n75 163.367
R386 B.n378 B.n75 163.367
R387 B.n378 B.n377 163.367
R388 B.n377 B.n376 163.367
R389 B.n376 B.n77 163.367
R390 B.n372 B.n77 163.367
R391 B.n372 B.n371 163.367
R392 B.n371 B.n370 163.367
R393 B.n370 B.n79 163.367
R394 B.n366 B.n79 163.367
R395 B.n366 B.n365 163.367
R396 B.n365 B.n364 163.367
R397 B.n364 B.n81 163.367
R398 B.n360 B.n81 163.367
R399 B.n360 B.n359 163.367
R400 B.n359 B.n358 163.367
R401 B.n358 B.n83 163.367
R402 B.n354 B.n83 163.367
R403 B.n354 B.n353 163.367
R404 B.n353 B.n352 163.367
R405 B.n352 B.n85 163.367
R406 B.n348 B.n85 163.367
R407 B.n348 B.n347 163.367
R408 B.n347 B.n346 163.367
R409 B.n346 B.n87 163.367
R410 B.n342 B.n87 163.367
R411 B.n342 B.n341 163.367
R412 B.n341 B.n340 163.367
R413 B.n340 B.n89 163.367
R414 B.n336 B.n89 163.367
R415 B.n336 B.n335 163.367
R416 B.n335 B.n334 163.367
R417 B.n334 B.n91 163.367
R418 B.n330 B.n91 163.367
R419 B.n330 B.n329 163.367
R420 B.n329 B.n328 163.367
R421 B.n328 B.n93 163.367
R422 B.n324 B.n93 163.367
R423 B.n324 B.n323 163.367
R424 B.n323 B.n322 163.367
R425 B.n322 B.n95 163.367
R426 B.n318 B.n95 163.367
R427 B.n318 B.n317 163.367
R428 B.n317 B.n316 163.367
R429 B.n316 B.n97 163.367
R430 B.n312 B.n97 163.367
R431 B.n312 B.n311 163.367
R432 B.n311 B.n310 163.367
R433 B.n310 B.n99 163.367
R434 B.n306 B.n99 163.367
R435 B.n306 B.n305 163.367
R436 B.n305 B.n304 163.367
R437 B.n304 B.n101 163.367
R438 B.n300 B.n101 163.367
R439 B.n300 B.n299 163.367
R440 B.n299 B.n298 163.367
R441 B.n298 B.n103 163.367
R442 B.n294 B.n103 163.367
R443 B.n294 B.n293 163.367
R444 B.n293 B.n292 163.367
R445 B.n292 B.n105 163.367
R446 B.n288 B.n105 163.367
R447 B.n288 B.n287 163.367
R448 B.n287 B.n286 163.367
R449 B.n286 B.n107 163.367
R450 B.n502 B.n31 163.367
R451 B.n498 B.n31 163.367
R452 B.n498 B.n497 163.367
R453 B.n497 B.n496 163.367
R454 B.n496 B.n33 163.367
R455 B.n492 B.n33 163.367
R456 B.n492 B.n491 163.367
R457 B.n491 B.n490 163.367
R458 B.n490 B.n35 163.367
R459 B.n485 B.n35 163.367
R460 B.n485 B.n484 163.367
R461 B.n484 B.n483 163.367
R462 B.n483 B.n39 163.367
R463 B.n479 B.n39 163.367
R464 B.n479 B.n478 163.367
R465 B.n478 B.n477 163.367
R466 B.n477 B.n41 163.367
R467 B.n473 B.n41 163.367
R468 B.n473 B.n472 163.367
R469 B.n472 B.n45 163.367
R470 B.n468 B.n45 163.367
R471 B.n468 B.n467 163.367
R472 B.n467 B.n466 163.367
R473 B.n466 B.n47 163.367
R474 B.n462 B.n47 163.367
R475 B.n462 B.n461 163.367
R476 B.n461 B.n460 163.367
R477 B.n460 B.n49 163.367
R478 B.n504 B.n503 163.367
R479 B.n504 B.n29 163.367
R480 B.n508 B.n29 163.367
R481 B.n509 B.n508 163.367
R482 B.n510 B.n509 163.367
R483 B.n510 B.n27 163.367
R484 B.n514 B.n27 163.367
R485 B.n515 B.n514 163.367
R486 B.n516 B.n515 163.367
R487 B.n516 B.n25 163.367
R488 B.n520 B.n25 163.367
R489 B.n521 B.n520 163.367
R490 B.n522 B.n521 163.367
R491 B.n522 B.n23 163.367
R492 B.n526 B.n23 163.367
R493 B.n527 B.n526 163.367
R494 B.n528 B.n527 163.367
R495 B.n528 B.n21 163.367
R496 B.n532 B.n21 163.367
R497 B.n533 B.n532 163.367
R498 B.n534 B.n533 163.367
R499 B.n534 B.n19 163.367
R500 B.n538 B.n19 163.367
R501 B.n539 B.n538 163.367
R502 B.n540 B.n539 163.367
R503 B.n540 B.n17 163.367
R504 B.n544 B.n17 163.367
R505 B.n545 B.n544 163.367
R506 B.n546 B.n545 163.367
R507 B.n546 B.n15 163.367
R508 B.n550 B.n15 163.367
R509 B.n551 B.n550 163.367
R510 B.n552 B.n551 163.367
R511 B.n552 B.n13 163.367
R512 B.n556 B.n13 163.367
R513 B.n557 B.n556 163.367
R514 B.n558 B.n557 163.367
R515 B.n558 B.n11 163.367
R516 B.n562 B.n11 163.367
R517 B.n563 B.n562 163.367
R518 B.n564 B.n563 163.367
R519 B.n564 B.n9 163.367
R520 B.n568 B.n9 163.367
R521 B.n569 B.n568 163.367
R522 B.n570 B.n569 163.367
R523 B.n570 B.n7 163.367
R524 B.n574 B.n7 163.367
R525 B.n575 B.n574 163.367
R526 B.n576 B.n575 163.367
R527 B.n576 B.n5 163.367
R528 B.n580 B.n5 163.367
R529 B.n581 B.n580 163.367
R530 B.n582 B.n581 163.367
R531 B.n582 B.n3 163.367
R532 B.n586 B.n3 163.367
R533 B.n587 B.n586 163.367
R534 B.n152 B.n2 163.367
R535 B.n152 B.n151 163.367
R536 B.n156 B.n151 163.367
R537 B.n157 B.n156 163.367
R538 B.n158 B.n157 163.367
R539 B.n158 B.n149 163.367
R540 B.n162 B.n149 163.367
R541 B.n163 B.n162 163.367
R542 B.n164 B.n163 163.367
R543 B.n164 B.n147 163.367
R544 B.n168 B.n147 163.367
R545 B.n169 B.n168 163.367
R546 B.n170 B.n169 163.367
R547 B.n170 B.n145 163.367
R548 B.n174 B.n145 163.367
R549 B.n175 B.n174 163.367
R550 B.n176 B.n175 163.367
R551 B.n176 B.n143 163.367
R552 B.n180 B.n143 163.367
R553 B.n181 B.n180 163.367
R554 B.n182 B.n181 163.367
R555 B.n182 B.n141 163.367
R556 B.n186 B.n141 163.367
R557 B.n187 B.n186 163.367
R558 B.n188 B.n187 163.367
R559 B.n188 B.n139 163.367
R560 B.n192 B.n139 163.367
R561 B.n193 B.n192 163.367
R562 B.n194 B.n193 163.367
R563 B.n194 B.n137 163.367
R564 B.n198 B.n137 163.367
R565 B.n199 B.n198 163.367
R566 B.n200 B.n199 163.367
R567 B.n200 B.n135 163.367
R568 B.n204 B.n135 163.367
R569 B.n205 B.n204 163.367
R570 B.n206 B.n205 163.367
R571 B.n206 B.n133 163.367
R572 B.n210 B.n133 163.367
R573 B.n211 B.n210 163.367
R574 B.n212 B.n211 163.367
R575 B.n212 B.n131 163.367
R576 B.n216 B.n131 163.367
R577 B.n217 B.n216 163.367
R578 B.n218 B.n217 163.367
R579 B.n218 B.n129 163.367
R580 B.n222 B.n129 163.367
R581 B.n223 B.n222 163.367
R582 B.n224 B.n223 163.367
R583 B.n224 B.n127 163.367
R584 B.n228 B.n127 163.367
R585 B.n229 B.n228 163.367
R586 B.n230 B.n229 163.367
R587 B.n230 B.n125 163.367
R588 B.n234 B.n125 163.367
R589 B.n235 B.n234 163.367
R590 B.n119 B.n118 65.3581
R591 B.n265 B.n264 65.3581
R592 B.n43 B.n42 65.3581
R593 B.n37 B.n36 65.3581
R594 B.n251 B.n119 59.5399
R595 B.n266 B.n265 59.5399
R596 B.n44 B.n43 59.5399
R597 B.n487 B.n37 59.5399
R598 B.n501 B.n30 33.8737
R599 B.n458 B.n457 33.8737
R600 B.n284 B.n283 33.8737
R601 B.n237 B.n124 33.8737
R602 B B.n589 18.0485
R603 B.n505 B.n30 10.6151
R604 B.n506 B.n505 10.6151
R605 B.n507 B.n506 10.6151
R606 B.n507 B.n28 10.6151
R607 B.n511 B.n28 10.6151
R608 B.n512 B.n511 10.6151
R609 B.n513 B.n512 10.6151
R610 B.n513 B.n26 10.6151
R611 B.n517 B.n26 10.6151
R612 B.n518 B.n517 10.6151
R613 B.n519 B.n518 10.6151
R614 B.n519 B.n24 10.6151
R615 B.n523 B.n24 10.6151
R616 B.n524 B.n523 10.6151
R617 B.n525 B.n524 10.6151
R618 B.n525 B.n22 10.6151
R619 B.n529 B.n22 10.6151
R620 B.n530 B.n529 10.6151
R621 B.n531 B.n530 10.6151
R622 B.n531 B.n20 10.6151
R623 B.n535 B.n20 10.6151
R624 B.n536 B.n535 10.6151
R625 B.n537 B.n536 10.6151
R626 B.n537 B.n18 10.6151
R627 B.n541 B.n18 10.6151
R628 B.n542 B.n541 10.6151
R629 B.n543 B.n542 10.6151
R630 B.n543 B.n16 10.6151
R631 B.n547 B.n16 10.6151
R632 B.n548 B.n547 10.6151
R633 B.n549 B.n548 10.6151
R634 B.n549 B.n14 10.6151
R635 B.n553 B.n14 10.6151
R636 B.n554 B.n553 10.6151
R637 B.n555 B.n554 10.6151
R638 B.n555 B.n12 10.6151
R639 B.n559 B.n12 10.6151
R640 B.n560 B.n559 10.6151
R641 B.n561 B.n560 10.6151
R642 B.n561 B.n10 10.6151
R643 B.n565 B.n10 10.6151
R644 B.n566 B.n565 10.6151
R645 B.n567 B.n566 10.6151
R646 B.n567 B.n8 10.6151
R647 B.n571 B.n8 10.6151
R648 B.n572 B.n571 10.6151
R649 B.n573 B.n572 10.6151
R650 B.n573 B.n6 10.6151
R651 B.n577 B.n6 10.6151
R652 B.n578 B.n577 10.6151
R653 B.n579 B.n578 10.6151
R654 B.n579 B.n4 10.6151
R655 B.n583 B.n4 10.6151
R656 B.n584 B.n583 10.6151
R657 B.n585 B.n584 10.6151
R658 B.n585 B.n0 10.6151
R659 B.n501 B.n500 10.6151
R660 B.n500 B.n499 10.6151
R661 B.n499 B.n32 10.6151
R662 B.n495 B.n32 10.6151
R663 B.n495 B.n494 10.6151
R664 B.n494 B.n493 10.6151
R665 B.n493 B.n34 10.6151
R666 B.n489 B.n34 10.6151
R667 B.n489 B.n488 10.6151
R668 B.n486 B.n38 10.6151
R669 B.n482 B.n38 10.6151
R670 B.n482 B.n481 10.6151
R671 B.n481 B.n480 10.6151
R672 B.n480 B.n40 10.6151
R673 B.n476 B.n40 10.6151
R674 B.n476 B.n475 10.6151
R675 B.n475 B.n474 10.6151
R676 B.n471 B.n470 10.6151
R677 B.n470 B.n469 10.6151
R678 B.n469 B.n46 10.6151
R679 B.n465 B.n46 10.6151
R680 B.n465 B.n464 10.6151
R681 B.n464 B.n463 10.6151
R682 B.n463 B.n48 10.6151
R683 B.n459 B.n48 10.6151
R684 B.n459 B.n458 10.6151
R685 B.n457 B.n50 10.6151
R686 B.n453 B.n50 10.6151
R687 B.n453 B.n452 10.6151
R688 B.n452 B.n451 10.6151
R689 B.n451 B.n52 10.6151
R690 B.n447 B.n52 10.6151
R691 B.n447 B.n446 10.6151
R692 B.n446 B.n445 10.6151
R693 B.n445 B.n54 10.6151
R694 B.n441 B.n54 10.6151
R695 B.n441 B.n440 10.6151
R696 B.n440 B.n439 10.6151
R697 B.n439 B.n56 10.6151
R698 B.n435 B.n56 10.6151
R699 B.n435 B.n434 10.6151
R700 B.n434 B.n433 10.6151
R701 B.n433 B.n58 10.6151
R702 B.n429 B.n58 10.6151
R703 B.n429 B.n428 10.6151
R704 B.n428 B.n427 10.6151
R705 B.n427 B.n60 10.6151
R706 B.n423 B.n60 10.6151
R707 B.n423 B.n422 10.6151
R708 B.n422 B.n421 10.6151
R709 B.n421 B.n62 10.6151
R710 B.n417 B.n62 10.6151
R711 B.n417 B.n416 10.6151
R712 B.n416 B.n415 10.6151
R713 B.n415 B.n64 10.6151
R714 B.n411 B.n64 10.6151
R715 B.n411 B.n410 10.6151
R716 B.n410 B.n409 10.6151
R717 B.n409 B.n66 10.6151
R718 B.n405 B.n66 10.6151
R719 B.n405 B.n404 10.6151
R720 B.n404 B.n403 10.6151
R721 B.n403 B.n68 10.6151
R722 B.n399 B.n68 10.6151
R723 B.n399 B.n398 10.6151
R724 B.n398 B.n397 10.6151
R725 B.n397 B.n70 10.6151
R726 B.n393 B.n70 10.6151
R727 B.n393 B.n392 10.6151
R728 B.n392 B.n391 10.6151
R729 B.n391 B.n72 10.6151
R730 B.n387 B.n72 10.6151
R731 B.n387 B.n386 10.6151
R732 B.n386 B.n385 10.6151
R733 B.n385 B.n74 10.6151
R734 B.n381 B.n74 10.6151
R735 B.n381 B.n380 10.6151
R736 B.n380 B.n379 10.6151
R737 B.n379 B.n76 10.6151
R738 B.n375 B.n76 10.6151
R739 B.n375 B.n374 10.6151
R740 B.n374 B.n373 10.6151
R741 B.n373 B.n78 10.6151
R742 B.n369 B.n78 10.6151
R743 B.n369 B.n368 10.6151
R744 B.n368 B.n367 10.6151
R745 B.n367 B.n80 10.6151
R746 B.n363 B.n80 10.6151
R747 B.n363 B.n362 10.6151
R748 B.n362 B.n361 10.6151
R749 B.n361 B.n82 10.6151
R750 B.n357 B.n82 10.6151
R751 B.n357 B.n356 10.6151
R752 B.n356 B.n355 10.6151
R753 B.n355 B.n84 10.6151
R754 B.n351 B.n84 10.6151
R755 B.n351 B.n350 10.6151
R756 B.n350 B.n349 10.6151
R757 B.n349 B.n86 10.6151
R758 B.n345 B.n86 10.6151
R759 B.n345 B.n344 10.6151
R760 B.n344 B.n343 10.6151
R761 B.n343 B.n88 10.6151
R762 B.n339 B.n88 10.6151
R763 B.n339 B.n338 10.6151
R764 B.n338 B.n337 10.6151
R765 B.n337 B.n90 10.6151
R766 B.n333 B.n90 10.6151
R767 B.n333 B.n332 10.6151
R768 B.n332 B.n331 10.6151
R769 B.n331 B.n92 10.6151
R770 B.n327 B.n92 10.6151
R771 B.n327 B.n326 10.6151
R772 B.n326 B.n325 10.6151
R773 B.n325 B.n94 10.6151
R774 B.n321 B.n94 10.6151
R775 B.n321 B.n320 10.6151
R776 B.n320 B.n319 10.6151
R777 B.n319 B.n96 10.6151
R778 B.n315 B.n96 10.6151
R779 B.n315 B.n314 10.6151
R780 B.n314 B.n313 10.6151
R781 B.n313 B.n98 10.6151
R782 B.n309 B.n98 10.6151
R783 B.n309 B.n308 10.6151
R784 B.n308 B.n307 10.6151
R785 B.n307 B.n100 10.6151
R786 B.n303 B.n100 10.6151
R787 B.n303 B.n302 10.6151
R788 B.n302 B.n301 10.6151
R789 B.n301 B.n102 10.6151
R790 B.n297 B.n102 10.6151
R791 B.n297 B.n296 10.6151
R792 B.n296 B.n295 10.6151
R793 B.n295 B.n104 10.6151
R794 B.n291 B.n104 10.6151
R795 B.n291 B.n290 10.6151
R796 B.n290 B.n289 10.6151
R797 B.n289 B.n106 10.6151
R798 B.n285 B.n106 10.6151
R799 B.n285 B.n284 10.6151
R800 B.n153 B.n1 10.6151
R801 B.n154 B.n153 10.6151
R802 B.n155 B.n154 10.6151
R803 B.n155 B.n150 10.6151
R804 B.n159 B.n150 10.6151
R805 B.n160 B.n159 10.6151
R806 B.n161 B.n160 10.6151
R807 B.n161 B.n148 10.6151
R808 B.n165 B.n148 10.6151
R809 B.n166 B.n165 10.6151
R810 B.n167 B.n166 10.6151
R811 B.n167 B.n146 10.6151
R812 B.n171 B.n146 10.6151
R813 B.n172 B.n171 10.6151
R814 B.n173 B.n172 10.6151
R815 B.n173 B.n144 10.6151
R816 B.n177 B.n144 10.6151
R817 B.n178 B.n177 10.6151
R818 B.n179 B.n178 10.6151
R819 B.n179 B.n142 10.6151
R820 B.n183 B.n142 10.6151
R821 B.n184 B.n183 10.6151
R822 B.n185 B.n184 10.6151
R823 B.n185 B.n140 10.6151
R824 B.n189 B.n140 10.6151
R825 B.n190 B.n189 10.6151
R826 B.n191 B.n190 10.6151
R827 B.n191 B.n138 10.6151
R828 B.n195 B.n138 10.6151
R829 B.n196 B.n195 10.6151
R830 B.n197 B.n196 10.6151
R831 B.n197 B.n136 10.6151
R832 B.n201 B.n136 10.6151
R833 B.n202 B.n201 10.6151
R834 B.n203 B.n202 10.6151
R835 B.n203 B.n134 10.6151
R836 B.n207 B.n134 10.6151
R837 B.n208 B.n207 10.6151
R838 B.n209 B.n208 10.6151
R839 B.n209 B.n132 10.6151
R840 B.n213 B.n132 10.6151
R841 B.n214 B.n213 10.6151
R842 B.n215 B.n214 10.6151
R843 B.n215 B.n130 10.6151
R844 B.n219 B.n130 10.6151
R845 B.n220 B.n219 10.6151
R846 B.n221 B.n220 10.6151
R847 B.n221 B.n128 10.6151
R848 B.n225 B.n128 10.6151
R849 B.n226 B.n225 10.6151
R850 B.n227 B.n226 10.6151
R851 B.n227 B.n126 10.6151
R852 B.n231 B.n126 10.6151
R853 B.n232 B.n231 10.6151
R854 B.n233 B.n232 10.6151
R855 B.n233 B.n124 10.6151
R856 B.n238 B.n237 10.6151
R857 B.n239 B.n238 10.6151
R858 B.n239 B.n122 10.6151
R859 B.n243 B.n122 10.6151
R860 B.n244 B.n243 10.6151
R861 B.n245 B.n244 10.6151
R862 B.n245 B.n120 10.6151
R863 B.n249 B.n120 10.6151
R864 B.n250 B.n249 10.6151
R865 B.n252 B.n116 10.6151
R866 B.n256 B.n116 10.6151
R867 B.n257 B.n256 10.6151
R868 B.n258 B.n257 10.6151
R869 B.n258 B.n114 10.6151
R870 B.n262 B.n114 10.6151
R871 B.n263 B.n262 10.6151
R872 B.n267 B.n263 10.6151
R873 B.n271 B.n112 10.6151
R874 B.n272 B.n271 10.6151
R875 B.n273 B.n272 10.6151
R876 B.n273 B.n110 10.6151
R877 B.n277 B.n110 10.6151
R878 B.n278 B.n277 10.6151
R879 B.n279 B.n278 10.6151
R880 B.n279 B.n108 10.6151
R881 B.n283 B.n108 10.6151
R882 B.n589 B.n0 8.11757
R883 B.n589 B.n1 8.11757
R884 B.n487 B.n486 6.5566
R885 B.n474 B.n44 6.5566
R886 B.n252 B.n251 6.5566
R887 B.n267 B.n266 6.5566
R888 B.n488 B.n487 4.05904
R889 B.n471 B.n44 4.05904
R890 B.n251 B.n250 4.05904
R891 B.n266 B.n112 4.05904
R892 VP.n21 VP.n18 161.3
R893 VP.n23 VP.n22 161.3
R894 VP.n24 VP.n17 161.3
R895 VP.n26 VP.n25 161.3
R896 VP.n27 VP.n16 161.3
R897 VP.n29 VP.n28 161.3
R898 VP.n31 VP.n30 161.3
R899 VP.n32 VP.n14 161.3
R900 VP.n34 VP.n33 161.3
R901 VP.n35 VP.n13 161.3
R902 VP.n37 VP.n36 161.3
R903 VP.n38 VP.n12 161.3
R904 VP.n40 VP.n39 161.3
R905 VP.n75 VP.n74 161.3
R906 VP.n73 VP.n1 161.3
R907 VP.n72 VP.n71 161.3
R908 VP.n70 VP.n2 161.3
R909 VP.n69 VP.n68 161.3
R910 VP.n67 VP.n3 161.3
R911 VP.n66 VP.n65 161.3
R912 VP.n64 VP.n63 161.3
R913 VP.n62 VP.n5 161.3
R914 VP.n61 VP.n60 161.3
R915 VP.n59 VP.n6 161.3
R916 VP.n58 VP.n57 161.3
R917 VP.n56 VP.n7 161.3
R918 VP.n54 VP.n53 161.3
R919 VP.n52 VP.n8 161.3
R920 VP.n51 VP.n50 161.3
R921 VP.n49 VP.n9 161.3
R922 VP.n48 VP.n47 161.3
R923 VP.n46 VP.n10 161.3
R924 VP.n45 VP.n44 161.3
R925 VP.n43 VP.n42 75.2445
R926 VP.n76 VP.n0 75.2445
R927 VP.n41 VP.n11 75.2445
R928 VP.n61 VP.n6 56.5617
R929 VP.n26 VP.n17 56.5617
R930 VP.n20 VP.n19 52.6903
R931 VP.n49 VP.n48 52.2023
R932 VP.n72 VP.n2 52.2023
R933 VP.n37 VP.n13 52.2023
R934 VP.n42 VP.n41 44.7799
R935 VP.n19 VP.t7 42.1945
R936 VP.n50 VP.n49 28.9518
R937 VP.n68 VP.n2 28.9518
R938 VP.n33 VP.n13 28.9518
R939 VP.n44 VP.n10 24.5923
R940 VP.n48 VP.n10 24.5923
R941 VP.n50 VP.n8 24.5923
R942 VP.n54 VP.n8 24.5923
R943 VP.n57 VP.n56 24.5923
R944 VP.n57 VP.n6 24.5923
R945 VP.n62 VP.n61 24.5923
R946 VP.n63 VP.n62 24.5923
R947 VP.n67 VP.n66 24.5923
R948 VP.n68 VP.n67 24.5923
R949 VP.n73 VP.n72 24.5923
R950 VP.n74 VP.n73 24.5923
R951 VP.n38 VP.n37 24.5923
R952 VP.n39 VP.n38 24.5923
R953 VP.n27 VP.n26 24.5923
R954 VP.n28 VP.n27 24.5923
R955 VP.n32 VP.n31 24.5923
R956 VP.n33 VP.n32 24.5923
R957 VP.n22 VP.n21 24.5923
R958 VP.n22 VP.n17 24.5923
R959 VP.n56 VP.n55 21.3954
R960 VP.n63 VP.n4 21.3954
R961 VP.n28 VP.n15 21.3954
R962 VP.n21 VP.n20 21.3954
R963 VP.n44 VP.n43 15.0015
R964 VP.n74 VP.n0 15.0015
R965 VP.n39 VP.n11 15.0015
R966 VP.n43 VP.t6 9.038
R967 VP.n55 VP.t2 9.038
R968 VP.n4 VP.t5 9.038
R969 VP.n0 VP.t4 9.038
R970 VP.n11 VP.t3 9.038
R971 VP.n15 VP.t0 9.038
R972 VP.n20 VP.t1 9.038
R973 VP.n19 VP.n18 4.13669
R974 VP.n55 VP.n54 3.19744
R975 VP.n66 VP.n4 3.19744
R976 VP.n31 VP.n15 3.19744
R977 VP.n41 VP.n40 0.354861
R978 VP.n45 VP.n42 0.354861
R979 VP.n76 VP.n75 0.354861
R980 VP VP.n76 0.267071
R981 VP.n23 VP.n18 0.189894
R982 VP.n24 VP.n23 0.189894
R983 VP.n25 VP.n24 0.189894
R984 VP.n25 VP.n16 0.189894
R985 VP.n29 VP.n16 0.189894
R986 VP.n30 VP.n29 0.189894
R987 VP.n30 VP.n14 0.189894
R988 VP.n34 VP.n14 0.189894
R989 VP.n35 VP.n34 0.189894
R990 VP.n36 VP.n35 0.189894
R991 VP.n36 VP.n12 0.189894
R992 VP.n40 VP.n12 0.189894
R993 VP.n46 VP.n45 0.189894
R994 VP.n47 VP.n46 0.189894
R995 VP.n47 VP.n9 0.189894
R996 VP.n51 VP.n9 0.189894
R997 VP.n52 VP.n51 0.189894
R998 VP.n53 VP.n52 0.189894
R999 VP.n53 VP.n7 0.189894
R1000 VP.n58 VP.n7 0.189894
R1001 VP.n59 VP.n58 0.189894
R1002 VP.n60 VP.n59 0.189894
R1003 VP.n60 VP.n5 0.189894
R1004 VP.n64 VP.n5 0.189894
R1005 VP.n65 VP.n64 0.189894
R1006 VP.n65 VP.n3 0.189894
R1007 VP.n69 VP.n3 0.189894
R1008 VP.n70 VP.n69 0.189894
R1009 VP.n71 VP.n70 0.189894
R1010 VP.n71 VP.n1 0.189894
R1011 VP.n75 VP.n1 0.189894
R1012 VDD1 VDD1.n0 348.55
R1013 VDD1.n3 VDD1.n2 348.437
R1014 VDD1.n3 VDD1.n1 348.437
R1015 VDD1.n5 VDD1.n4 347.039
R1016 VDD1.n5 VDD1.n3 38.3543
R1017 VDD1.n4 VDD1.t2 28.5137
R1018 VDD1.n4 VDD1.t0 28.5137
R1019 VDD1.n0 VDD1.t3 28.5137
R1020 VDD1.n0 VDD1.t7 28.5137
R1021 VDD1.n2 VDD1.t5 28.5137
R1022 VDD1.n2 VDD1.t6 28.5137
R1023 VDD1.n1 VDD1.t1 28.5137
R1024 VDD1.n1 VDD1.t4 28.5137
R1025 VDD1 VDD1.n5 1.3949
R1026 VTAIL.n15 VTAIL.t1 373.298
R1027 VTAIL.n2 VTAIL.t5 373.298
R1028 VTAIL.n3 VTAIL.t11 373.298
R1029 VTAIL.n6 VTAIL.t9 373.298
R1030 VTAIL.n14 VTAIL.t12 373.298
R1031 VTAIL.n11 VTAIL.t8 373.298
R1032 VTAIL.n10 VTAIL.t2 373.298
R1033 VTAIL.n7 VTAIL.t6 373.298
R1034 VTAIL.n1 VTAIL.n0 330.361
R1035 VTAIL.n5 VTAIL.n4 330.361
R1036 VTAIL.n13 VTAIL.n12 330.36
R1037 VTAIL.n9 VTAIL.n8 330.36
R1038 VTAIL.n0 VTAIL.t3 28.5137
R1039 VTAIL.n0 VTAIL.t4 28.5137
R1040 VTAIL.n4 VTAIL.t13 28.5137
R1041 VTAIL.n4 VTAIL.t10 28.5137
R1042 VTAIL.n12 VTAIL.t14 28.5137
R1043 VTAIL.n12 VTAIL.t15 28.5137
R1044 VTAIL.n8 VTAIL.t0 28.5137
R1045 VTAIL.n8 VTAIL.t7 28.5137
R1046 VTAIL.n15 VTAIL.n14 16.2548
R1047 VTAIL.n7 VTAIL.n6 16.2548
R1048 VTAIL.n9 VTAIL.n7 2.90567
R1049 VTAIL.n10 VTAIL.n9 2.90567
R1050 VTAIL.n13 VTAIL.n11 2.90567
R1051 VTAIL.n14 VTAIL.n13 2.90567
R1052 VTAIL.n6 VTAIL.n5 2.90567
R1053 VTAIL.n5 VTAIL.n3 2.90567
R1054 VTAIL.n2 VTAIL.n1 2.90567
R1055 VTAIL VTAIL.n15 2.84748
R1056 VTAIL.n11 VTAIL.n10 0.470328
R1057 VTAIL.n3 VTAIL.n2 0.470328
R1058 VTAIL VTAIL.n1 0.0586897
R1059 VN.n60 VN.n59 161.3
R1060 VN.n58 VN.n32 161.3
R1061 VN.n57 VN.n56 161.3
R1062 VN.n55 VN.n33 161.3
R1063 VN.n54 VN.n53 161.3
R1064 VN.n52 VN.n34 161.3
R1065 VN.n51 VN.n50 161.3
R1066 VN.n49 VN.n48 161.3
R1067 VN.n47 VN.n36 161.3
R1068 VN.n46 VN.n45 161.3
R1069 VN.n44 VN.n37 161.3
R1070 VN.n43 VN.n42 161.3
R1071 VN.n41 VN.n38 161.3
R1072 VN.n29 VN.n28 161.3
R1073 VN.n27 VN.n1 161.3
R1074 VN.n26 VN.n25 161.3
R1075 VN.n24 VN.n2 161.3
R1076 VN.n23 VN.n22 161.3
R1077 VN.n21 VN.n3 161.3
R1078 VN.n20 VN.n19 161.3
R1079 VN.n18 VN.n17 161.3
R1080 VN.n16 VN.n5 161.3
R1081 VN.n15 VN.n14 161.3
R1082 VN.n13 VN.n6 161.3
R1083 VN.n12 VN.n11 161.3
R1084 VN.n10 VN.n7 161.3
R1085 VN.n30 VN.n0 75.2445
R1086 VN.n61 VN.n31 75.2445
R1087 VN.n15 VN.n6 56.5617
R1088 VN.n46 VN.n37 56.5617
R1089 VN.n9 VN.n8 52.6903
R1090 VN.n40 VN.n39 52.6903
R1091 VN.n26 VN.n2 52.2023
R1092 VN.n57 VN.n33 52.2023
R1093 VN VN.n61 44.9451
R1094 VN.n39 VN.t2 42.1947
R1095 VN.n8 VN.t1 42.1947
R1096 VN.n22 VN.n2 28.9518
R1097 VN.n53 VN.n33 28.9518
R1098 VN.n11 VN.n10 24.5923
R1099 VN.n11 VN.n6 24.5923
R1100 VN.n16 VN.n15 24.5923
R1101 VN.n17 VN.n16 24.5923
R1102 VN.n21 VN.n20 24.5923
R1103 VN.n22 VN.n21 24.5923
R1104 VN.n27 VN.n26 24.5923
R1105 VN.n28 VN.n27 24.5923
R1106 VN.n42 VN.n37 24.5923
R1107 VN.n42 VN.n41 24.5923
R1108 VN.n53 VN.n52 24.5923
R1109 VN.n52 VN.n51 24.5923
R1110 VN.n48 VN.n47 24.5923
R1111 VN.n47 VN.n46 24.5923
R1112 VN.n59 VN.n58 24.5923
R1113 VN.n58 VN.n57 24.5923
R1114 VN.n10 VN.n9 21.3954
R1115 VN.n17 VN.n4 21.3954
R1116 VN.n41 VN.n40 21.3954
R1117 VN.n48 VN.n35 21.3954
R1118 VN.n28 VN.n0 15.0015
R1119 VN.n59 VN.n31 15.0015
R1120 VN.n9 VN.t4 9.038
R1121 VN.n4 VN.t3 9.038
R1122 VN.n0 VN.t6 9.038
R1123 VN.n40 VN.t5 9.038
R1124 VN.n35 VN.t7 9.038
R1125 VN.n31 VN.t0 9.038
R1126 VN.n8 VN.n7 4.13672
R1127 VN.n39 VN.n38 4.13672
R1128 VN.n20 VN.n4 3.19744
R1129 VN.n51 VN.n35 3.19744
R1130 VN.n61 VN.n60 0.354861
R1131 VN.n30 VN.n29 0.354861
R1132 VN VN.n30 0.267071
R1133 VN.n60 VN.n32 0.189894
R1134 VN.n56 VN.n32 0.189894
R1135 VN.n56 VN.n55 0.189894
R1136 VN.n55 VN.n54 0.189894
R1137 VN.n54 VN.n34 0.189894
R1138 VN.n50 VN.n34 0.189894
R1139 VN.n50 VN.n49 0.189894
R1140 VN.n49 VN.n36 0.189894
R1141 VN.n45 VN.n36 0.189894
R1142 VN.n45 VN.n44 0.189894
R1143 VN.n44 VN.n43 0.189894
R1144 VN.n43 VN.n38 0.189894
R1145 VN.n12 VN.n7 0.189894
R1146 VN.n13 VN.n12 0.189894
R1147 VN.n14 VN.n13 0.189894
R1148 VN.n14 VN.n5 0.189894
R1149 VN.n18 VN.n5 0.189894
R1150 VN.n19 VN.n18 0.189894
R1151 VN.n19 VN.n3 0.189894
R1152 VN.n23 VN.n3 0.189894
R1153 VN.n24 VN.n23 0.189894
R1154 VN.n25 VN.n24 0.189894
R1155 VN.n25 VN.n1 0.189894
R1156 VN.n29 VN.n1 0.189894
R1157 VDD2.n2 VDD2.n1 348.437
R1158 VDD2.n2 VDD2.n0 348.437
R1159 VDD2 VDD2.n5 348.435
R1160 VDD2.n4 VDD2.n3 347.038
R1161 VDD2.n4 VDD2.n2 37.7713
R1162 VDD2.n5 VDD2.t2 28.5137
R1163 VDD2.n5 VDD2.t5 28.5137
R1164 VDD2.n3 VDD2.t7 28.5137
R1165 VDD2.n3 VDD2.t0 28.5137
R1166 VDD2.n1 VDD2.t4 28.5137
R1167 VDD2.n1 VDD2.t1 28.5137
R1168 VDD2.n0 VDD2.t6 28.5137
R1169 VDD2.n0 VDD2.t3 28.5137
R1170 VDD2 VDD2.n4 1.51128
C0 VP VDD1 1.68966f
C1 B VDD2 1.60052f
C2 VTAIL B 1.35375f
C3 w_n4340_n1196# B 7.83639f
C4 VN B 1.17722f
C5 VTAIL VDD2 4.90127f
C6 B VP 2.12507f
C7 w_n4340_n1196# VDD2 1.92909f
C8 VN VDD2 1.27783f
C9 VTAIL w_n4340_n1196# 1.77031f
C10 VTAIL VN 2.73325f
C11 B VDD1 1.49001f
C12 VN w_n4340_n1196# 8.790179f
C13 VDD2 VP 0.575625f
C14 VTAIL VP 2.74736f
C15 VDD2 VDD1 2.00625f
C16 w_n4340_n1196# VP 9.34762f
C17 VN VP 6.19694f
C18 VTAIL VDD1 4.8439f
C19 w_n4340_n1196# VDD1 1.79694f
C20 VN VDD1 0.159709f
C21 VDD2 VSUBS 1.471942f
C22 VDD1 VSUBS 2.165771f
C23 VTAIL VSUBS 0.581033f
C24 VN VSUBS 7.65802f
C25 VP VSUBS 3.392471f
C26 B VSUBS 4.290339f
C27 w_n4340_n1196# VSUBS 66.8186f
C28 VDD2.t6 VSUBS 0.024218f
C29 VDD2.t3 VSUBS 0.024218f
C30 VDD2.n0 VSUBS 0.082942f
C31 VDD2.t4 VSUBS 0.024218f
C32 VDD2.t1 VSUBS 0.024218f
C33 VDD2.n1 VSUBS 0.082942f
C34 VDD2.n2 VSUBS 3.10069f
C35 VDD2.t7 VSUBS 0.024218f
C36 VDD2.t0 VSUBS 0.024218f
C37 VDD2.n3 VSUBS 0.080526f
C38 VDD2.n4 VSUBS 2.42537f
C39 VDD2.t2 VSUBS 0.024218f
C40 VDD2.t5 VSUBS 0.024218f
C41 VDD2.n5 VSUBS 0.082934f
C42 VN.t6 VSUBS 0.384644f
C43 VN.n0 VSUBS 0.436418f
C44 VN.n1 VSUBS 0.055969f
C45 VN.n2 VSUBS 0.056398f
C46 VN.n3 VSUBS 0.055969f
C47 VN.t3 VSUBS 0.384644f
C48 VN.n4 VSUBS 0.232434f
C49 VN.n5 VSUBS 0.055969f
C50 VN.n6 VSUBS 0.08136f
C51 VN.n7 VSUBS 0.639348f
C52 VN.t4 VSUBS 0.384644f
C53 VN.t1 VSUBS 0.865733f
C54 VN.n8 VSUBS 0.446836f
C55 VN.n9 VSUBS 0.431029f
C56 VN.n10 VSUBS 0.097129f
C57 VN.n11 VSUBS 0.10379f
C58 VN.n12 VSUBS 0.055969f
C59 VN.n13 VSUBS 0.055969f
C60 VN.n14 VSUBS 0.055969f
C61 VN.n15 VSUBS 0.08136f
C62 VN.n16 VSUBS 0.10379f
C63 VN.n17 VSUBS 0.097129f
C64 VN.n18 VSUBS 0.055969f
C65 VN.n19 VSUBS 0.055969f
C66 VN.n20 VSUBS 0.059213f
C67 VN.n21 VSUBS 0.10379f
C68 VN.n22 VSUBS 0.110117f
C69 VN.n23 VSUBS 0.055969f
C70 VN.n24 VSUBS 0.055969f
C71 VN.n25 VSUBS 0.055969f
C72 VN.n26 VSUBS 0.099996f
C73 VN.n27 VSUBS 0.10379f
C74 VN.n28 VSUBS 0.083807f
C75 VN.n29 VSUBS 0.090319f
C76 VN.n30 VSUBS 0.12884f
C77 VN.t0 VSUBS 0.384644f
C78 VN.n31 VSUBS 0.436418f
C79 VN.n32 VSUBS 0.055969f
C80 VN.n33 VSUBS 0.056398f
C81 VN.n34 VSUBS 0.055969f
C82 VN.t7 VSUBS 0.384644f
C83 VN.n35 VSUBS 0.232434f
C84 VN.n36 VSUBS 0.055969f
C85 VN.n37 VSUBS 0.08136f
C86 VN.n38 VSUBS 0.639349f
C87 VN.t5 VSUBS 0.384644f
C88 VN.t2 VSUBS 0.865733f
C89 VN.n39 VSUBS 0.446836f
C90 VN.n40 VSUBS 0.431029f
C91 VN.n41 VSUBS 0.097129f
C92 VN.n42 VSUBS 0.10379f
C93 VN.n43 VSUBS 0.055969f
C94 VN.n44 VSUBS 0.055969f
C95 VN.n45 VSUBS 0.055969f
C96 VN.n46 VSUBS 0.08136f
C97 VN.n47 VSUBS 0.10379f
C98 VN.n48 VSUBS 0.097129f
C99 VN.n49 VSUBS 0.055969f
C100 VN.n50 VSUBS 0.055969f
C101 VN.n51 VSUBS 0.059213f
C102 VN.n52 VSUBS 0.10379f
C103 VN.n53 VSUBS 0.110117f
C104 VN.n54 VSUBS 0.055969f
C105 VN.n55 VSUBS 0.055969f
C106 VN.n56 VSUBS 0.055969f
C107 VN.n57 VSUBS 0.099996f
C108 VN.n58 VSUBS 0.10379f
C109 VN.n59 VSUBS 0.083807f
C110 VN.n60 VSUBS 0.090319f
C111 VN.n61 VSUBS 2.71858f
C112 VTAIL.t3 VSUBS 0.033652f
C113 VTAIL.t4 VSUBS 0.033652f
C114 VTAIL.n0 VSUBS 0.096937f
C115 VTAIL.n1 VSUBS 0.624234f
C116 VTAIL.t5 VSUBS 0.169738f
C117 VTAIL.n2 VSUBS 0.692758f
C118 VTAIL.t11 VSUBS 0.169738f
C119 VTAIL.n3 VSUBS 0.692758f
C120 VTAIL.t13 VSUBS 0.033652f
C121 VTAIL.t10 VSUBS 0.033652f
C122 VTAIL.n4 VSUBS 0.096937f
C123 VTAIL.n5 VSUBS 0.966916f
C124 VTAIL.t9 VSUBS 0.169738f
C125 VTAIL.n6 VSUBS 1.61161f
C126 VTAIL.t6 VSUBS 0.169738f
C127 VTAIL.n7 VSUBS 1.61161f
C128 VTAIL.t0 VSUBS 0.033652f
C129 VTAIL.t7 VSUBS 0.033652f
C130 VTAIL.n8 VSUBS 0.096936f
C131 VTAIL.n9 VSUBS 0.966916f
C132 VTAIL.t2 VSUBS 0.169738f
C133 VTAIL.n10 VSUBS 0.692758f
C134 VTAIL.t8 VSUBS 0.169738f
C135 VTAIL.n11 VSUBS 0.692758f
C136 VTAIL.t14 VSUBS 0.033652f
C137 VTAIL.t15 VSUBS 0.033652f
C138 VTAIL.n12 VSUBS 0.096936f
C139 VTAIL.n13 VSUBS 0.966916f
C140 VTAIL.t12 VSUBS 0.169738f
C141 VTAIL.n14 VSUBS 1.61161f
C142 VTAIL.t1 VSUBS 0.169738f
C143 VTAIL.n15 VSUBS 1.6046f
C144 VDD1.t3 VSUBS 0.023529f
C145 VDD1.t7 VSUBS 0.023529f
C146 VDD1.n0 VSUBS 0.080809f
C147 VDD1.t1 VSUBS 0.023529f
C148 VDD1.t4 VSUBS 0.023529f
C149 VDD1.n1 VSUBS 0.08058f
C150 VDD1.t5 VSUBS 0.023529f
C151 VDD1.t6 VSUBS 0.023529f
C152 VDD1.n2 VSUBS 0.08058f
C153 VDD1.n3 VSUBS 3.06677f
C154 VDD1.t2 VSUBS 0.023529f
C155 VDD1.t0 VSUBS 0.023529f
C156 VDD1.n4 VSUBS 0.078234f
C157 VDD1.n5 VSUBS 2.38862f
C158 VP.t4 VSUBS 0.443115f
C159 VP.n0 VSUBS 0.502759f
C160 VP.n1 VSUBS 0.064477f
C161 VP.n2 VSUBS 0.064971f
C162 VP.n3 VSUBS 0.064477f
C163 VP.t5 VSUBS 0.443115f
C164 VP.n4 VSUBS 0.267767f
C165 VP.n5 VSUBS 0.064477f
C166 VP.n6 VSUBS 0.093728f
C167 VP.n7 VSUBS 0.064477f
C168 VP.t2 VSUBS 0.443115f
C169 VP.n8 VSUBS 0.119568f
C170 VP.n9 VSUBS 0.064477f
C171 VP.n10 VSUBS 0.119568f
C172 VP.t3 VSUBS 0.443115f
C173 VP.n11 VSUBS 0.502759f
C174 VP.n12 VSUBS 0.064477f
C175 VP.n13 VSUBS 0.064971f
C176 VP.n14 VSUBS 0.064477f
C177 VP.t0 VSUBS 0.443115f
C178 VP.n15 VSUBS 0.267767f
C179 VP.n16 VSUBS 0.064477f
C180 VP.n17 VSUBS 0.093728f
C181 VP.n18 VSUBS 0.736539f
C182 VP.t1 VSUBS 0.443115f
C183 VP.t7 VSUBS 0.997335f
C184 VP.n19 VSUBS 0.514762f
C185 VP.n20 VSUBS 0.496552f
C186 VP.n21 VSUBS 0.111894f
C187 VP.n22 VSUBS 0.119568f
C188 VP.n23 VSUBS 0.064477f
C189 VP.n24 VSUBS 0.064477f
C190 VP.n25 VSUBS 0.064477f
C191 VP.n26 VSUBS 0.093728f
C192 VP.n27 VSUBS 0.119568f
C193 VP.n28 VSUBS 0.111894f
C194 VP.n29 VSUBS 0.064477f
C195 VP.n30 VSUBS 0.064477f
C196 VP.n31 VSUBS 0.068214f
C197 VP.n32 VSUBS 0.119568f
C198 VP.n33 VSUBS 0.126856f
C199 VP.n34 VSUBS 0.064477f
C200 VP.n35 VSUBS 0.064477f
C201 VP.n36 VSUBS 0.064477f
C202 VP.n37 VSUBS 0.115197f
C203 VP.n38 VSUBS 0.119568f
C204 VP.n39 VSUBS 0.096547f
C205 VP.n40 VSUBS 0.104049f
C206 VP.n41 VSUBS 3.10439f
C207 VP.n42 VSUBS 3.1563f
C208 VP.t6 VSUBS 0.443115f
C209 VP.n43 VSUBS 0.502759f
C210 VP.n44 VSUBS 0.096547f
C211 VP.n45 VSUBS 0.104049f
C212 VP.n46 VSUBS 0.064477f
C213 VP.n47 VSUBS 0.064477f
C214 VP.n48 VSUBS 0.115197f
C215 VP.n49 VSUBS 0.064971f
C216 VP.n50 VSUBS 0.126856f
C217 VP.n51 VSUBS 0.064477f
C218 VP.n52 VSUBS 0.064477f
C219 VP.n53 VSUBS 0.064477f
C220 VP.n54 VSUBS 0.068214f
C221 VP.n55 VSUBS 0.267767f
C222 VP.n56 VSUBS 0.111894f
C223 VP.n57 VSUBS 0.119568f
C224 VP.n58 VSUBS 0.064477f
C225 VP.n59 VSUBS 0.064477f
C226 VP.n60 VSUBS 0.064477f
C227 VP.n61 VSUBS 0.093728f
C228 VP.n62 VSUBS 0.119568f
C229 VP.n63 VSUBS 0.111894f
C230 VP.n64 VSUBS 0.064477f
C231 VP.n65 VSUBS 0.064477f
C232 VP.n66 VSUBS 0.068214f
C233 VP.n67 VSUBS 0.119568f
C234 VP.n68 VSUBS 0.126856f
C235 VP.n69 VSUBS 0.064477f
C236 VP.n70 VSUBS 0.064477f
C237 VP.n71 VSUBS 0.064477f
C238 VP.n72 VSUBS 0.115197f
C239 VP.n73 VSUBS 0.119568f
C240 VP.n74 VSUBS 0.096547f
C241 VP.n75 VSUBS 0.104049f
C242 VP.n76 VSUBS 0.148426f
C243 B.n0 VSUBS 0.01083f
C244 B.n1 VSUBS 0.01083f
C245 B.n2 VSUBS 0.016017f
C246 B.n3 VSUBS 0.012274f
C247 B.n4 VSUBS 0.012274f
C248 B.n5 VSUBS 0.012274f
C249 B.n6 VSUBS 0.012274f
C250 B.n7 VSUBS 0.012274f
C251 B.n8 VSUBS 0.012274f
C252 B.n9 VSUBS 0.012274f
C253 B.n10 VSUBS 0.012274f
C254 B.n11 VSUBS 0.012274f
C255 B.n12 VSUBS 0.012274f
C256 B.n13 VSUBS 0.012274f
C257 B.n14 VSUBS 0.012274f
C258 B.n15 VSUBS 0.012274f
C259 B.n16 VSUBS 0.012274f
C260 B.n17 VSUBS 0.012274f
C261 B.n18 VSUBS 0.012274f
C262 B.n19 VSUBS 0.012274f
C263 B.n20 VSUBS 0.012274f
C264 B.n21 VSUBS 0.012274f
C265 B.n22 VSUBS 0.012274f
C266 B.n23 VSUBS 0.012274f
C267 B.n24 VSUBS 0.012274f
C268 B.n25 VSUBS 0.012274f
C269 B.n26 VSUBS 0.012274f
C270 B.n27 VSUBS 0.012274f
C271 B.n28 VSUBS 0.012274f
C272 B.n29 VSUBS 0.012274f
C273 B.n30 VSUBS 0.028519f
C274 B.n31 VSUBS 0.012274f
C275 B.n32 VSUBS 0.012274f
C276 B.n33 VSUBS 0.012274f
C277 B.n34 VSUBS 0.012274f
C278 B.n35 VSUBS 0.012274f
C279 B.t7 VSUBS 0.037659f
C280 B.t8 VSUBS 0.048492f
C281 B.t6 VSUBS 0.306708f
C282 B.n36 VSUBS 0.11731f
C283 B.n37 VSUBS 0.088659f
C284 B.n38 VSUBS 0.012274f
C285 B.n39 VSUBS 0.012274f
C286 B.n40 VSUBS 0.012274f
C287 B.n41 VSUBS 0.012274f
C288 B.t1 VSUBS 0.037659f
C289 B.t2 VSUBS 0.048492f
C290 B.t0 VSUBS 0.306708f
C291 B.n42 VSUBS 0.11731f
C292 B.n43 VSUBS 0.088659f
C293 B.n44 VSUBS 0.028438f
C294 B.n45 VSUBS 0.012274f
C295 B.n46 VSUBS 0.012274f
C296 B.n47 VSUBS 0.012274f
C297 B.n48 VSUBS 0.012274f
C298 B.n49 VSUBS 0.030326f
C299 B.n50 VSUBS 0.012274f
C300 B.n51 VSUBS 0.012274f
C301 B.n52 VSUBS 0.012274f
C302 B.n53 VSUBS 0.012274f
C303 B.n54 VSUBS 0.012274f
C304 B.n55 VSUBS 0.012274f
C305 B.n56 VSUBS 0.012274f
C306 B.n57 VSUBS 0.012274f
C307 B.n58 VSUBS 0.012274f
C308 B.n59 VSUBS 0.012274f
C309 B.n60 VSUBS 0.012274f
C310 B.n61 VSUBS 0.012274f
C311 B.n62 VSUBS 0.012274f
C312 B.n63 VSUBS 0.012274f
C313 B.n64 VSUBS 0.012274f
C314 B.n65 VSUBS 0.012274f
C315 B.n66 VSUBS 0.012274f
C316 B.n67 VSUBS 0.012274f
C317 B.n68 VSUBS 0.012274f
C318 B.n69 VSUBS 0.012274f
C319 B.n70 VSUBS 0.012274f
C320 B.n71 VSUBS 0.012274f
C321 B.n72 VSUBS 0.012274f
C322 B.n73 VSUBS 0.012274f
C323 B.n74 VSUBS 0.012274f
C324 B.n75 VSUBS 0.012274f
C325 B.n76 VSUBS 0.012274f
C326 B.n77 VSUBS 0.012274f
C327 B.n78 VSUBS 0.012274f
C328 B.n79 VSUBS 0.012274f
C329 B.n80 VSUBS 0.012274f
C330 B.n81 VSUBS 0.012274f
C331 B.n82 VSUBS 0.012274f
C332 B.n83 VSUBS 0.012274f
C333 B.n84 VSUBS 0.012274f
C334 B.n85 VSUBS 0.012274f
C335 B.n86 VSUBS 0.012274f
C336 B.n87 VSUBS 0.012274f
C337 B.n88 VSUBS 0.012274f
C338 B.n89 VSUBS 0.012274f
C339 B.n90 VSUBS 0.012274f
C340 B.n91 VSUBS 0.012274f
C341 B.n92 VSUBS 0.012274f
C342 B.n93 VSUBS 0.012274f
C343 B.n94 VSUBS 0.012274f
C344 B.n95 VSUBS 0.012274f
C345 B.n96 VSUBS 0.012274f
C346 B.n97 VSUBS 0.012274f
C347 B.n98 VSUBS 0.012274f
C348 B.n99 VSUBS 0.012274f
C349 B.n100 VSUBS 0.012274f
C350 B.n101 VSUBS 0.012274f
C351 B.n102 VSUBS 0.012274f
C352 B.n103 VSUBS 0.012274f
C353 B.n104 VSUBS 0.012274f
C354 B.n105 VSUBS 0.012274f
C355 B.n106 VSUBS 0.012274f
C356 B.n107 VSUBS 0.028519f
C357 B.n108 VSUBS 0.012274f
C358 B.n109 VSUBS 0.012274f
C359 B.n110 VSUBS 0.012274f
C360 B.n111 VSUBS 0.012274f
C361 B.n112 VSUBS 0.008484f
C362 B.n113 VSUBS 0.012274f
C363 B.n114 VSUBS 0.012274f
C364 B.n115 VSUBS 0.012274f
C365 B.n116 VSUBS 0.012274f
C366 B.n117 VSUBS 0.012274f
C367 B.t11 VSUBS 0.037659f
C368 B.t10 VSUBS 0.048492f
C369 B.t9 VSUBS 0.306708f
C370 B.n118 VSUBS 0.11731f
C371 B.n119 VSUBS 0.088659f
C372 B.n120 VSUBS 0.012274f
C373 B.n121 VSUBS 0.012274f
C374 B.n122 VSUBS 0.012274f
C375 B.n123 VSUBS 0.012274f
C376 B.n124 VSUBS 0.028519f
C377 B.n125 VSUBS 0.012274f
C378 B.n126 VSUBS 0.012274f
C379 B.n127 VSUBS 0.012274f
C380 B.n128 VSUBS 0.012274f
C381 B.n129 VSUBS 0.012274f
C382 B.n130 VSUBS 0.012274f
C383 B.n131 VSUBS 0.012274f
C384 B.n132 VSUBS 0.012274f
C385 B.n133 VSUBS 0.012274f
C386 B.n134 VSUBS 0.012274f
C387 B.n135 VSUBS 0.012274f
C388 B.n136 VSUBS 0.012274f
C389 B.n137 VSUBS 0.012274f
C390 B.n138 VSUBS 0.012274f
C391 B.n139 VSUBS 0.012274f
C392 B.n140 VSUBS 0.012274f
C393 B.n141 VSUBS 0.012274f
C394 B.n142 VSUBS 0.012274f
C395 B.n143 VSUBS 0.012274f
C396 B.n144 VSUBS 0.012274f
C397 B.n145 VSUBS 0.012274f
C398 B.n146 VSUBS 0.012274f
C399 B.n147 VSUBS 0.012274f
C400 B.n148 VSUBS 0.012274f
C401 B.n149 VSUBS 0.012274f
C402 B.n150 VSUBS 0.012274f
C403 B.n151 VSUBS 0.012274f
C404 B.n152 VSUBS 0.012274f
C405 B.n153 VSUBS 0.012274f
C406 B.n154 VSUBS 0.012274f
C407 B.n155 VSUBS 0.012274f
C408 B.n156 VSUBS 0.012274f
C409 B.n157 VSUBS 0.012274f
C410 B.n158 VSUBS 0.012274f
C411 B.n159 VSUBS 0.012274f
C412 B.n160 VSUBS 0.012274f
C413 B.n161 VSUBS 0.012274f
C414 B.n162 VSUBS 0.012274f
C415 B.n163 VSUBS 0.012274f
C416 B.n164 VSUBS 0.012274f
C417 B.n165 VSUBS 0.012274f
C418 B.n166 VSUBS 0.012274f
C419 B.n167 VSUBS 0.012274f
C420 B.n168 VSUBS 0.012274f
C421 B.n169 VSUBS 0.012274f
C422 B.n170 VSUBS 0.012274f
C423 B.n171 VSUBS 0.012274f
C424 B.n172 VSUBS 0.012274f
C425 B.n173 VSUBS 0.012274f
C426 B.n174 VSUBS 0.012274f
C427 B.n175 VSUBS 0.012274f
C428 B.n176 VSUBS 0.012274f
C429 B.n177 VSUBS 0.012274f
C430 B.n178 VSUBS 0.012274f
C431 B.n179 VSUBS 0.012274f
C432 B.n180 VSUBS 0.012274f
C433 B.n181 VSUBS 0.012274f
C434 B.n182 VSUBS 0.012274f
C435 B.n183 VSUBS 0.012274f
C436 B.n184 VSUBS 0.012274f
C437 B.n185 VSUBS 0.012274f
C438 B.n186 VSUBS 0.012274f
C439 B.n187 VSUBS 0.012274f
C440 B.n188 VSUBS 0.012274f
C441 B.n189 VSUBS 0.012274f
C442 B.n190 VSUBS 0.012274f
C443 B.n191 VSUBS 0.012274f
C444 B.n192 VSUBS 0.012274f
C445 B.n193 VSUBS 0.012274f
C446 B.n194 VSUBS 0.012274f
C447 B.n195 VSUBS 0.012274f
C448 B.n196 VSUBS 0.012274f
C449 B.n197 VSUBS 0.012274f
C450 B.n198 VSUBS 0.012274f
C451 B.n199 VSUBS 0.012274f
C452 B.n200 VSUBS 0.012274f
C453 B.n201 VSUBS 0.012274f
C454 B.n202 VSUBS 0.012274f
C455 B.n203 VSUBS 0.012274f
C456 B.n204 VSUBS 0.012274f
C457 B.n205 VSUBS 0.012274f
C458 B.n206 VSUBS 0.012274f
C459 B.n207 VSUBS 0.012274f
C460 B.n208 VSUBS 0.012274f
C461 B.n209 VSUBS 0.012274f
C462 B.n210 VSUBS 0.012274f
C463 B.n211 VSUBS 0.012274f
C464 B.n212 VSUBS 0.012274f
C465 B.n213 VSUBS 0.012274f
C466 B.n214 VSUBS 0.012274f
C467 B.n215 VSUBS 0.012274f
C468 B.n216 VSUBS 0.012274f
C469 B.n217 VSUBS 0.012274f
C470 B.n218 VSUBS 0.012274f
C471 B.n219 VSUBS 0.012274f
C472 B.n220 VSUBS 0.012274f
C473 B.n221 VSUBS 0.012274f
C474 B.n222 VSUBS 0.012274f
C475 B.n223 VSUBS 0.012274f
C476 B.n224 VSUBS 0.012274f
C477 B.n225 VSUBS 0.012274f
C478 B.n226 VSUBS 0.012274f
C479 B.n227 VSUBS 0.012274f
C480 B.n228 VSUBS 0.012274f
C481 B.n229 VSUBS 0.012274f
C482 B.n230 VSUBS 0.012274f
C483 B.n231 VSUBS 0.012274f
C484 B.n232 VSUBS 0.012274f
C485 B.n233 VSUBS 0.012274f
C486 B.n234 VSUBS 0.012274f
C487 B.n235 VSUBS 0.028519f
C488 B.n236 VSUBS 0.030326f
C489 B.n237 VSUBS 0.030326f
C490 B.n238 VSUBS 0.012274f
C491 B.n239 VSUBS 0.012274f
C492 B.n240 VSUBS 0.012274f
C493 B.n241 VSUBS 0.012274f
C494 B.n242 VSUBS 0.012274f
C495 B.n243 VSUBS 0.012274f
C496 B.n244 VSUBS 0.012274f
C497 B.n245 VSUBS 0.012274f
C498 B.n246 VSUBS 0.012274f
C499 B.n247 VSUBS 0.012274f
C500 B.n248 VSUBS 0.012274f
C501 B.n249 VSUBS 0.012274f
C502 B.n250 VSUBS 0.008484f
C503 B.n251 VSUBS 0.028438f
C504 B.n252 VSUBS 0.009928f
C505 B.n253 VSUBS 0.012274f
C506 B.n254 VSUBS 0.012274f
C507 B.n255 VSUBS 0.012274f
C508 B.n256 VSUBS 0.012274f
C509 B.n257 VSUBS 0.012274f
C510 B.n258 VSUBS 0.012274f
C511 B.n259 VSUBS 0.012274f
C512 B.n260 VSUBS 0.012274f
C513 B.n261 VSUBS 0.012274f
C514 B.n262 VSUBS 0.012274f
C515 B.n263 VSUBS 0.012274f
C516 B.t5 VSUBS 0.037659f
C517 B.t4 VSUBS 0.048492f
C518 B.t3 VSUBS 0.306708f
C519 B.n264 VSUBS 0.11731f
C520 B.n265 VSUBS 0.088659f
C521 B.n266 VSUBS 0.028438f
C522 B.n267 VSUBS 0.009928f
C523 B.n268 VSUBS 0.012274f
C524 B.n269 VSUBS 0.012274f
C525 B.n270 VSUBS 0.012274f
C526 B.n271 VSUBS 0.012274f
C527 B.n272 VSUBS 0.012274f
C528 B.n273 VSUBS 0.012274f
C529 B.n274 VSUBS 0.012274f
C530 B.n275 VSUBS 0.012274f
C531 B.n276 VSUBS 0.012274f
C532 B.n277 VSUBS 0.012274f
C533 B.n278 VSUBS 0.012274f
C534 B.n279 VSUBS 0.012274f
C535 B.n280 VSUBS 0.012274f
C536 B.n281 VSUBS 0.012274f
C537 B.n282 VSUBS 0.030326f
C538 B.n283 VSUBS 0.028928f
C539 B.n284 VSUBS 0.029917f
C540 B.n285 VSUBS 0.012274f
C541 B.n286 VSUBS 0.012274f
C542 B.n287 VSUBS 0.012274f
C543 B.n288 VSUBS 0.012274f
C544 B.n289 VSUBS 0.012274f
C545 B.n290 VSUBS 0.012274f
C546 B.n291 VSUBS 0.012274f
C547 B.n292 VSUBS 0.012274f
C548 B.n293 VSUBS 0.012274f
C549 B.n294 VSUBS 0.012274f
C550 B.n295 VSUBS 0.012274f
C551 B.n296 VSUBS 0.012274f
C552 B.n297 VSUBS 0.012274f
C553 B.n298 VSUBS 0.012274f
C554 B.n299 VSUBS 0.012274f
C555 B.n300 VSUBS 0.012274f
C556 B.n301 VSUBS 0.012274f
C557 B.n302 VSUBS 0.012274f
C558 B.n303 VSUBS 0.012274f
C559 B.n304 VSUBS 0.012274f
C560 B.n305 VSUBS 0.012274f
C561 B.n306 VSUBS 0.012274f
C562 B.n307 VSUBS 0.012274f
C563 B.n308 VSUBS 0.012274f
C564 B.n309 VSUBS 0.012274f
C565 B.n310 VSUBS 0.012274f
C566 B.n311 VSUBS 0.012274f
C567 B.n312 VSUBS 0.012274f
C568 B.n313 VSUBS 0.012274f
C569 B.n314 VSUBS 0.012274f
C570 B.n315 VSUBS 0.012274f
C571 B.n316 VSUBS 0.012274f
C572 B.n317 VSUBS 0.012274f
C573 B.n318 VSUBS 0.012274f
C574 B.n319 VSUBS 0.012274f
C575 B.n320 VSUBS 0.012274f
C576 B.n321 VSUBS 0.012274f
C577 B.n322 VSUBS 0.012274f
C578 B.n323 VSUBS 0.012274f
C579 B.n324 VSUBS 0.012274f
C580 B.n325 VSUBS 0.012274f
C581 B.n326 VSUBS 0.012274f
C582 B.n327 VSUBS 0.012274f
C583 B.n328 VSUBS 0.012274f
C584 B.n329 VSUBS 0.012274f
C585 B.n330 VSUBS 0.012274f
C586 B.n331 VSUBS 0.012274f
C587 B.n332 VSUBS 0.012274f
C588 B.n333 VSUBS 0.012274f
C589 B.n334 VSUBS 0.012274f
C590 B.n335 VSUBS 0.012274f
C591 B.n336 VSUBS 0.012274f
C592 B.n337 VSUBS 0.012274f
C593 B.n338 VSUBS 0.012274f
C594 B.n339 VSUBS 0.012274f
C595 B.n340 VSUBS 0.012274f
C596 B.n341 VSUBS 0.012274f
C597 B.n342 VSUBS 0.012274f
C598 B.n343 VSUBS 0.012274f
C599 B.n344 VSUBS 0.012274f
C600 B.n345 VSUBS 0.012274f
C601 B.n346 VSUBS 0.012274f
C602 B.n347 VSUBS 0.012274f
C603 B.n348 VSUBS 0.012274f
C604 B.n349 VSUBS 0.012274f
C605 B.n350 VSUBS 0.012274f
C606 B.n351 VSUBS 0.012274f
C607 B.n352 VSUBS 0.012274f
C608 B.n353 VSUBS 0.012274f
C609 B.n354 VSUBS 0.012274f
C610 B.n355 VSUBS 0.012274f
C611 B.n356 VSUBS 0.012274f
C612 B.n357 VSUBS 0.012274f
C613 B.n358 VSUBS 0.012274f
C614 B.n359 VSUBS 0.012274f
C615 B.n360 VSUBS 0.012274f
C616 B.n361 VSUBS 0.012274f
C617 B.n362 VSUBS 0.012274f
C618 B.n363 VSUBS 0.012274f
C619 B.n364 VSUBS 0.012274f
C620 B.n365 VSUBS 0.012274f
C621 B.n366 VSUBS 0.012274f
C622 B.n367 VSUBS 0.012274f
C623 B.n368 VSUBS 0.012274f
C624 B.n369 VSUBS 0.012274f
C625 B.n370 VSUBS 0.012274f
C626 B.n371 VSUBS 0.012274f
C627 B.n372 VSUBS 0.012274f
C628 B.n373 VSUBS 0.012274f
C629 B.n374 VSUBS 0.012274f
C630 B.n375 VSUBS 0.012274f
C631 B.n376 VSUBS 0.012274f
C632 B.n377 VSUBS 0.012274f
C633 B.n378 VSUBS 0.012274f
C634 B.n379 VSUBS 0.012274f
C635 B.n380 VSUBS 0.012274f
C636 B.n381 VSUBS 0.012274f
C637 B.n382 VSUBS 0.012274f
C638 B.n383 VSUBS 0.012274f
C639 B.n384 VSUBS 0.012274f
C640 B.n385 VSUBS 0.012274f
C641 B.n386 VSUBS 0.012274f
C642 B.n387 VSUBS 0.012274f
C643 B.n388 VSUBS 0.012274f
C644 B.n389 VSUBS 0.012274f
C645 B.n390 VSUBS 0.012274f
C646 B.n391 VSUBS 0.012274f
C647 B.n392 VSUBS 0.012274f
C648 B.n393 VSUBS 0.012274f
C649 B.n394 VSUBS 0.012274f
C650 B.n395 VSUBS 0.012274f
C651 B.n396 VSUBS 0.012274f
C652 B.n397 VSUBS 0.012274f
C653 B.n398 VSUBS 0.012274f
C654 B.n399 VSUBS 0.012274f
C655 B.n400 VSUBS 0.012274f
C656 B.n401 VSUBS 0.012274f
C657 B.n402 VSUBS 0.012274f
C658 B.n403 VSUBS 0.012274f
C659 B.n404 VSUBS 0.012274f
C660 B.n405 VSUBS 0.012274f
C661 B.n406 VSUBS 0.012274f
C662 B.n407 VSUBS 0.012274f
C663 B.n408 VSUBS 0.012274f
C664 B.n409 VSUBS 0.012274f
C665 B.n410 VSUBS 0.012274f
C666 B.n411 VSUBS 0.012274f
C667 B.n412 VSUBS 0.012274f
C668 B.n413 VSUBS 0.012274f
C669 B.n414 VSUBS 0.012274f
C670 B.n415 VSUBS 0.012274f
C671 B.n416 VSUBS 0.012274f
C672 B.n417 VSUBS 0.012274f
C673 B.n418 VSUBS 0.012274f
C674 B.n419 VSUBS 0.012274f
C675 B.n420 VSUBS 0.012274f
C676 B.n421 VSUBS 0.012274f
C677 B.n422 VSUBS 0.012274f
C678 B.n423 VSUBS 0.012274f
C679 B.n424 VSUBS 0.012274f
C680 B.n425 VSUBS 0.012274f
C681 B.n426 VSUBS 0.012274f
C682 B.n427 VSUBS 0.012274f
C683 B.n428 VSUBS 0.012274f
C684 B.n429 VSUBS 0.012274f
C685 B.n430 VSUBS 0.012274f
C686 B.n431 VSUBS 0.012274f
C687 B.n432 VSUBS 0.012274f
C688 B.n433 VSUBS 0.012274f
C689 B.n434 VSUBS 0.012274f
C690 B.n435 VSUBS 0.012274f
C691 B.n436 VSUBS 0.012274f
C692 B.n437 VSUBS 0.012274f
C693 B.n438 VSUBS 0.012274f
C694 B.n439 VSUBS 0.012274f
C695 B.n440 VSUBS 0.012274f
C696 B.n441 VSUBS 0.012274f
C697 B.n442 VSUBS 0.012274f
C698 B.n443 VSUBS 0.012274f
C699 B.n444 VSUBS 0.012274f
C700 B.n445 VSUBS 0.012274f
C701 B.n446 VSUBS 0.012274f
C702 B.n447 VSUBS 0.012274f
C703 B.n448 VSUBS 0.012274f
C704 B.n449 VSUBS 0.012274f
C705 B.n450 VSUBS 0.012274f
C706 B.n451 VSUBS 0.012274f
C707 B.n452 VSUBS 0.012274f
C708 B.n453 VSUBS 0.012274f
C709 B.n454 VSUBS 0.012274f
C710 B.n455 VSUBS 0.012274f
C711 B.n456 VSUBS 0.028519f
C712 B.n457 VSUBS 0.028519f
C713 B.n458 VSUBS 0.030326f
C714 B.n459 VSUBS 0.012274f
C715 B.n460 VSUBS 0.012274f
C716 B.n461 VSUBS 0.012274f
C717 B.n462 VSUBS 0.012274f
C718 B.n463 VSUBS 0.012274f
C719 B.n464 VSUBS 0.012274f
C720 B.n465 VSUBS 0.012274f
C721 B.n466 VSUBS 0.012274f
C722 B.n467 VSUBS 0.012274f
C723 B.n468 VSUBS 0.012274f
C724 B.n469 VSUBS 0.012274f
C725 B.n470 VSUBS 0.012274f
C726 B.n471 VSUBS 0.008484f
C727 B.n472 VSUBS 0.012274f
C728 B.n473 VSUBS 0.012274f
C729 B.n474 VSUBS 0.009928f
C730 B.n475 VSUBS 0.012274f
C731 B.n476 VSUBS 0.012274f
C732 B.n477 VSUBS 0.012274f
C733 B.n478 VSUBS 0.012274f
C734 B.n479 VSUBS 0.012274f
C735 B.n480 VSUBS 0.012274f
C736 B.n481 VSUBS 0.012274f
C737 B.n482 VSUBS 0.012274f
C738 B.n483 VSUBS 0.012274f
C739 B.n484 VSUBS 0.012274f
C740 B.n485 VSUBS 0.012274f
C741 B.n486 VSUBS 0.009928f
C742 B.n487 VSUBS 0.028438f
C743 B.n488 VSUBS 0.008484f
C744 B.n489 VSUBS 0.012274f
C745 B.n490 VSUBS 0.012274f
C746 B.n491 VSUBS 0.012274f
C747 B.n492 VSUBS 0.012274f
C748 B.n493 VSUBS 0.012274f
C749 B.n494 VSUBS 0.012274f
C750 B.n495 VSUBS 0.012274f
C751 B.n496 VSUBS 0.012274f
C752 B.n497 VSUBS 0.012274f
C753 B.n498 VSUBS 0.012274f
C754 B.n499 VSUBS 0.012274f
C755 B.n500 VSUBS 0.012274f
C756 B.n501 VSUBS 0.030326f
C757 B.n502 VSUBS 0.030326f
C758 B.n503 VSUBS 0.028519f
C759 B.n504 VSUBS 0.012274f
C760 B.n505 VSUBS 0.012274f
C761 B.n506 VSUBS 0.012274f
C762 B.n507 VSUBS 0.012274f
C763 B.n508 VSUBS 0.012274f
C764 B.n509 VSUBS 0.012274f
C765 B.n510 VSUBS 0.012274f
C766 B.n511 VSUBS 0.012274f
C767 B.n512 VSUBS 0.012274f
C768 B.n513 VSUBS 0.012274f
C769 B.n514 VSUBS 0.012274f
C770 B.n515 VSUBS 0.012274f
C771 B.n516 VSUBS 0.012274f
C772 B.n517 VSUBS 0.012274f
C773 B.n518 VSUBS 0.012274f
C774 B.n519 VSUBS 0.012274f
C775 B.n520 VSUBS 0.012274f
C776 B.n521 VSUBS 0.012274f
C777 B.n522 VSUBS 0.012274f
C778 B.n523 VSUBS 0.012274f
C779 B.n524 VSUBS 0.012274f
C780 B.n525 VSUBS 0.012274f
C781 B.n526 VSUBS 0.012274f
C782 B.n527 VSUBS 0.012274f
C783 B.n528 VSUBS 0.012274f
C784 B.n529 VSUBS 0.012274f
C785 B.n530 VSUBS 0.012274f
C786 B.n531 VSUBS 0.012274f
C787 B.n532 VSUBS 0.012274f
C788 B.n533 VSUBS 0.012274f
C789 B.n534 VSUBS 0.012274f
C790 B.n535 VSUBS 0.012274f
C791 B.n536 VSUBS 0.012274f
C792 B.n537 VSUBS 0.012274f
C793 B.n538 VSUBS 0.012274f
C794 B.n539 VSUBS 0.012274f
C795 B.n540 VSUBS 0.012274f
C796 B.n541 VSUBS 0.012274f
C797 B.n542 VSUBS 0.012274f
C798 B.n543 VSUBS 0.012274f
C799 B.n544 VSUBS 0.012274f
C800 B.n545 VSUBS 0.012274f
C801 B.n546 VSUBS 0.012274f
C802 B.n547 VSUBS 0.012274f
C803 B.n548 VSUBS 0.012274f
C804 B.n549 VSUBS 0.012274f
C805 B.n550 VSUBS 0.012274f
C806 B.n551 VSUBS 0.012274f
C807 B.n552 VSUBS 0.012274f
C808 B.n553 VSUBS 0.012274f
C809 B.n554 VSUBS 0.012274f
C810 B.n555 VSUBS 0.012274f
C811 B.n556 VSUBS 0.012274f
C812 B.n557 VSUBS 0.012274f
C813 B.n558 VSUBS 0.012274f
C814 B.n559 VSUBS 0.012274f
C815 B.n560 VSUBS 0.012274f
C816 B.n561 VSUBS 0.012274f
C817 B.n562 VSUBS 0.012274f
C818 B.n563 VSUBS 0.012274f
C819 B.n564 VSUBS 0.012274f
C820 B.n565 VSUBS 0.012274f
C821 B.n566 VSUBS 0.012274f
C822 B.n567 VSUBS 0.012274f
C823 B.n568 VSUBS 0.012274f
C824 B.n569 VSUBS 0.012274f
C825 B.n570 VSUBS 0.012274f
C826 B.n571 VSUBS 0.012274f
C827 B.n572 VSUBS 0.012274f
C828 B.n573 VSUBS 0.012274f
C829 B.n574 VSUBS 0.012274f
C830 B.n575 VSUBS 0.012274f
C831 B.n576 VSUBS 0.012274f
C832 B.n577 VSUBS 0.012274f
C833 B.n578 VSUBS 0.012274f
C834 B.n579 VSUBS 0.012274f
C835 B.n580 VSUBS 0.012274f
C836 B.n581 VSUBS 0.012274f
C837 B.n582 VSUBS 0.012274f
C838 B.n583 VSUBS 0.012274f
C839 B.n584 VSUBS 0.012274f
C840 B.n585 VSUBS 0.012274f
C841 B.n586 VSUBS 0.012274f
C842 B.n587 VSUBS 0.016017f
C843 B.n588 VSUBS 0.017063f
C844 B.n589 VSUBS 0.03393f
.ends

