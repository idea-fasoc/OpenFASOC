* NGSPICE file created from diff_pair_sample_1414.ext - technology: sky130A

.subckt diff_pair_sample_1414 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t6 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=1.32165 ps=8.34 w=8.01 l=1.2
X1 B.t11 B.t9 B.t10 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=3.1239 pd=16.8 as=0 ps=0 w=8.01 l=1.2
X2 VDD1.t2 VP.t1 VTAIL.t14 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=3.1239 ps=16.8 w=8.01 l=1.2
X3 B.t8 B.t6 B.t7 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=3.1239 pd=16.8 as=0 ps=0 w=8.01 l=1.2
X4 VDD1.t3 VP.t2 VTAIL.t13 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=1.32165 ps=8.34 w=8.01 l=1.2
X5 VDD2.t7 VN.t0 VTAIL.t2 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=3.1239 ps=16.8 w=8.01 l=1.2
X6 VDD2.t6 VN.t1 VTAIL.t1 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=3.1239 ps=16.8 w=8.01 l=1.2
X7 VTAIL.t6 VN.t2 VDD2.t5 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=1.32165 ps=8.34 w=8.01 l=1.2
X8 VTAIL.t7 VN.t3 VDD2.t4 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=1.32165 ps=8.34 w=8.01 l=1.2
X9 B.t5 B.t3 B.t4 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=3.1239 pd=16.8 as=0 ps=0 w=8.01 l=1.2
X10 VTAIL.t12 VP.t3 VDD1.t1 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=3.1239 pd=16.8 as=1.32165 ps=8.34 w=8.01 l=1.2
X11 VTAIL.t11 VP.t4 VDD1.t0 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=1.32165 ps=8.34 w=8.01 l=1.2
X12 VDD2.t3 VN.t4 VTAIL.t4 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=1.32165 ps=8.34 w=8.01 l=1.2
X13 B.t2 B.t0 B.t1 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=3.1239 pd=16.8 as=0 ps=0 w=8.01 l=1.2
X14 VDD1.t7 VP.t5 VTAIL.t10 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=3.1239 ps=16.8 w=8.01 l=1.2
X15 VDD2.t2 VN.t5 VTAIL.t0 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=1.32165 ps=8.34 w=8.01 l=1.2
X16 VDD1.t5 VP.t6 VTAIL.t9 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=1.32165 pd=8.34 as=1.32165 ps=8.34 w=8.01 l=1.2
X17 VTAIL.t8 VP.t7 VDD1.t4 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=3.1239 pd=16.8 as=1.32165 ps=8.34 w=8.01 l=1.2
X18 VTAIL.t3 VN.t6 VDD2.t1 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=3.1239 pd=16.8 as=1.32165 ps=8.34 w=8.01 l=1.2
X19 VTAIL.t5 VN.t7 VDD2.t0 w_n2500_n2570# sky130_fd_pr__pfet_01v8 ad=3.1239 pd=16.8 as=1.32165 ps=8.34 w=8.01 l=1.2
R0 VP.n9 VP.t3 212.308
R1 VP.n21 VP.t7 193.804
R2 VP.n33 VP.t5 193.804
R3 VP.n18 VP.t1 193.804
R4 VP.n11 VP.n10 161.3
R5 VP.n12 VP.n7 161.3
R6 VP.n14 VP.n13 161.3
R7 VP.n16 VP.n15 161.3
R8 VP.n17 VP.n5 161.3
R9 VP.n32 VP.n0 161.3
R10 VP.n31 VP.n30 161.3
R11 VP.n29 VP.n28 161.3
R12 VP.n27 VP.n2 161.3
R13 VP.n26 VP.n25 161.3
R14 VP.n24 VP.n23 161.3
R15 VP.n22 VP.n4 161.3
R16 VP.n3 VP.t2 160.868
R17 VP.n1 VP.t4 160.868
R18 VP.n6 VP.t0 160.868
R19 VP.n8 VP.t6 160.868
R20 VP.n19 VP.n18 80.6037
R21 VP.n34 VP.n33 80.6037
R22 VP.n21 VP.n20 80.6037
R23 VP.n9 VP.n8 44.8004
R24 VP.n20 VP.n19 41.4332
R25 VP.n27 VP.n26 40.4934
R26 VP.n28 VP.n27 40.4934
R27 VP.n13 VP.n12 40.4934
R28 VP.n12 VP.n11 40.4934
R29 VP.n23 VP.n22 37.5796
R30 VP.n32 VP.n31 37.5796
R31 VP.n17 VP.n16 37.5796
R32 VP.n10 VP.n9 29.7304
R33 VP.n22 VP.n21 28.4823
R34 VP.n33 VP.n32 28.4823
R35 VP.n18 VP.n17 28.4823
R36 VP.n26 VP.n3 12.968
R37 VP.n28 VP.n1 12.968
R38 VP.n13 VP.n6 12.968
R39 VP.n11 VP.n8 12.968
R40 VP.n23 VP.n3 11.5
R41 VP.n31 VP.n1 11.5
R42 VP.n16 VP.n6 11.5
R43 VP.n19 VP.n5 0.285035
R44 VP.n20 VP.n4 0.285035
R45 VP.n34 VP.n0 0.285035
R46 VP.n10 VP.n7 0.189894
R47 VP.n14 VP.n7 0.189894
R48 VP.n15 VP.n14 0.189894
R49 VP.n15 VP.n5 0.189894
R50 VP.n24 VP.n4 0.189894
R51 VP.n25 VP.n24 0.189894
R52 VP.n25 VP.n2 0.189894
R53 VP.n29 VP.n2 0.189894
R54 VP.n30 VP.n29 0.189894
R55 VP.n30 VP.n0 0.189894
R56 VP VP.n34 0.146778
R57 VDD1 VDD1.n0 87.1496
R58 VDD1.n3 VDD1.n2 87.0359
R59 VDD1.n3 VDD1.n1 87.0359
R60 VDD1.n5 VDD1.n4 86.4318
R61 VDD1.n5 VDD1.n3 37.1388
R62 VDD1.n4 VDD1.t6 4.05855
R63 VDD1.n4 VDD1.t2 4.05855
R64 VDD1.n0 VDD1.t1 4.05855
R65 VDD1.n0 VDD1.t5 4.05855
R66 VDD1.n2 VDD1.t0 4.05855
R67 VDD1.n2 VDD1.t7 4.05855
R68 VDD1.n1 VDD1.t4 4.05855
R69 VDD1.n1 VDD1.t3 4.05855
R70 VDD1 VDD1.n5 0.601793
R71 VTAIL.n338 VTAIL.n302 756.745
R72 VTAIL.n38 VTAIL.n2 756.745
R73 VTAIL.n80 VTAIL.n44 756.745
R74 VTAIL.n124 VTAIL.n88 756.745
R75 VTAIL.n296 VTAIL.n260 756.745
R76 VTAIL.n252 VTAIL.n216 756.745
R77 VTAIL.n210 VTAIL.n174 756.745
R78 VTAIL.n166 VTAIL.n130 756.745
R79 VTAIL.n314 VTAIL.n313 585
R80 VTAIL.n319 VTAIL.n318 585
R81 VTAIL.n321 VTAIL.n320 585
R82 VTAIL.n310 VTAIL.n309 585
R83 VTAIL.n327 VTAIL.n326 585
R84 VTAIL.n329 VTAIL.n328 585
R85 VTAIL.n306 VTAIL.n305 585
R86 VTAIL.n336 VTAIL.n335 585
R87 VTAIL.n337 VTAIL.n304 585
R88 VTAIL.n339 VTAIL.n338 585
R89 VTAIL.n14 VTAIL.n13 585
R90 VTAIL.n19 VTAIL.n18 585
R91 VTAIL.n21 VTAIL.n20 585
R92 VTAIL.n10 VTAIL.n9 585
R93 VTAIL.n27 VTAIL.n26 585
R94 VTAIL.n29 VTAIL.n28 585
R95 VTAIL.n6 VTAIL.n5 585
R96 VTAIL.n36 VTAIL.n35 585
R97 VTAIL.n37 VTAIL.n4 585
R98 VTAIL.n39 VTAIL.n38 585
R99 VTAIL.n56 VTAIL.n55 585
R100 VTAIL.n61 VTAIL.n60 585
R101 VTAIL.n63 VTAIL.n62 585
R102 VTAIL.n52 VTAIL.n51 585
R103 VTAIL.n69 VTAIL.n68 585
R104 VTAIL.n71 VTAIL.n70 585
R105 VTAIL.n48 VTAIL.n47 585
R106 VTAIL.n78 VTAIL.n77 585
R107 VTAIL.n79 VTAIL.n46 585
R108 VTAIL.n81 VTAIL.n80 585
R109 VTAIL.n100 VTAIL.n99 585
R110 VTAIL.n105 VTAIL.n104 585
R111 VTAIL.n107 VTAIL.n106 585
R112 VTAIL.n96 VTAIL.n95 585
R113 VTAIL.n113 VTAIL.n112 585
R114 VTAIL.n115 VTAIL.n114 585
R115 VTAIL.n92 VTAIL.n91 585
R116 VTAIL.n122 VTAIL.n121 585
R117 VTAIL.n123 VTAIL.n90 585
R118 VTAIL.n125 VTAIL.n124 585
R119 VTAIL.n297 VTAIL.n296 585
R120 VTAIL.n295 VTAIL.n262 585
R121 VTAIL.n294 VTAIL.n293 585
R122 VTAIL.n265 VTAIL.n263 585
R123 VTAIL.n288 VTAIL.n287 585
R124 VTAIL.n286 VTAIL.n285 585
R125 VTAIL.n269 VTAIL.n268 585
R126 VTAIL.n280 VTAIL.n279 585
R127 VTAIL.n278 VTAIL.n277 585
R128 VTAIL.n273 VTAIL.n272 585
R129 VTAIL.n253 VTAIL.n252 585
R130 VTAIL.n251 VTAIL.n218 585
R131 VTAIL.n250 VTAIL.n249 585
R132 VTAIL.n221 VTAIL.n219 585
R133 VTAIL.n244 VTAIL.n243 585
R134 VTAIL.n242 VTAIL.n241 585
R135 VTAIL.n225 VTAIL.n224 585
R136 VTAIL.n236 VTAIL.n235 585
R137 VTAIL.n234 VTAIL.n233 585
R138 VTAIL.n229 VTAIL.n228 585
R139 VTAIL.n211 VTAIL.n210 585
R140 VTAIL.n209 VTAIL.n176 585
R141 VTAIL.n208 VTAIL.n207 585
R142 VTAIL.n179 VTAIL.n177 585
R143 VTAIL.n202 VTAIL.n201 585
R144 VTAIL.n200 VTAIL.n199 585
R145 VTAIL.n183 VTAIL.n182 585
R146 VTAIL.n194 VTAIL.n193 585
R147 VTAIL.n192 VTAIL.n191 585
R148 VTAIL.n187 VTAIL.n186 585
R149 VTAIL.n167 VTAIL.n166 585
R150 VTAIL.n165 VTAIL.n132 585
R151 VTAIL.n164 VTAIL.n163 585
R152 VTAIL.n135 VTAIL.n133 585
R153 VTAIL.n158 VTAIL.n157 585
R154 VTAIL.n156 VTAIL.n155 585
R155 VTAIL.n139 VTAIL.n138 585
R156 VTAIL.n150 VTAIL.n149 585
R157 VTAIL.n148 VTAIL.n147 585
R158 VTAIL.n143 VTAIL.n142 585
R159 VTAIL.n315 VTAIL.t1 329.043
R160 VTAIL.n15 VTAIL.t3 329.043
R161 VTAIL.n57 VTAIL.t10 329.043
R162 VTAIL.n101 VTAIL.t8 329.043
R163 VTAIL.n274 VTAIL.t14 329.043
R164 VTAIL.n230 VTAIL.t12 329.043
R165 VTAIL.n188 VTAIL.t2 329.043
R166 VTAIL.n144 VTAIL.t5 329.043
R167 VTAIL.n319 VTAIL.n313 171.744
R168 VTAIL.n320 VTAIL.n319 171.744
R169 VTAIL.n320 VTAIL.n309 171.744
R170 VTAIL.n327 VTAIL.n309 171.744
R171 VTAIL.n328 VTAIL.n327 171.744
R172 VTAIL.n328 VTAIL.n305 171.744
R173 VTAIL.n336 VTAIL.n305 171.744
R174 VTAIL.n337 VTAIL.n336 171.744
R175 VTAIL.n338 VTAIL.n337 171.744
R176 VTAIL.n19 VTAIL.n13 171.744
R177 VTAIL.n20 VTAIL.n19 171.744
R178 VTAIL.n20 VTAIL.n9 171.744
R179 VTAIL.n27 VTAIL.n9 171.744
R180 VTAIL.n28 VTAIL.n27 171.744
R181 VTAIL.n28 VTAIL.n5 171.744
R182 VTAIL.n36 VTAIL.n5 171.744
R183 VTAIL.n37 VTAIL.n36 171.744
R184 VTAIL.n38 VTAIL.n37 171.744
R185 VTAIL.n61 VTAIL.n55 171.744
R186 VTAIL.n62 VTAIL.n61 171.744
R187 VTAIL.n62 VTAIL.n51 171.744
R188 VTAIL.n69 VTAIL.n51 171.744
R189 VTAIL.n70 VTAIL.n69 171.744
R190 VTAIL.n70 VTAIL.n47 171.744
R191 VTAIL.n78 VTAIL.n47 171.744
R192 VTAIL.n79 VTAIL.n78 171.744
R193 VTAIL.n80 VTAIL.n79 171.744
R194 VTAIL.n105 VTAIL.n99 171.744
R195 VTAIL.n106 VTAIL.n105 171.744
R196 VTAIL.n106 VTAIL.n95 171.744
R197 VTAIL.n113 VTAIL.n95 171.744
R198 VTAIL.n114 VTAIL.n113 171.744
R199 VTAIL.n114 VTAIL.n91 171.744
R200 VTAIL.n122 VTAIL.n91 171.744
R201 VTAIL.n123 VTAIL.n122 171.744
R202 VTAIL.n124 VTAIL.n123 171.744
R203 VTAIL.n296 VTAIL.n295 171.744
R204 VTAIL.n295 VTAIL.n294 171.744
R205 VTAIL.n294 VTAIL.n263 171.744
R206 VTAIL.n287 VTAIL.n263 171.744
R207 VTAIL.n287 VTAIL.n286 171.744
R208 VTAIL.n286 VTAIL.n268 171.744
R209 VTAIL.n279 VTAIL.n268 171.744
R210 VTAIL.n279 VTAIL.n278 171.744
R211 VTAIL.n278 VTAIL.n272 171.744
R212 VTAIL.n252 VTAIL.n251 171.744
R213 VTAIL.n251 VTAIL.n250 171.744
R214 VTAIL.n250 VTAIL.n219 171.744
R215 VTAIL.n243 VTAIL.n219 171.744
R216 VTAIL.n243 VTAIL.n242 171.744
R217 VTAIL.n242 VTAIL.n224 171.744
R218 VTAIL.n235 VTAIL.n224 171.744
R219 VTAIL.n235 VTAIL.n234 171.744
R220 VTAIL.n234 VTAIL.n228 171.744
R221 VTAIL.n210 VTAIL.n209 171.744
R222 VTAIL.n209 VTAIL.n208 171.744
R223 VTAIL.n208 VTAIL.n177 171.744
R224 VTAIL.n201 VTAIL.n177 171.744
R225 VTAIL.n201 VTAIL.n200 171.744
R226 VTAIL.n200 VTAIL.n182 171.744
R227 VTAIL.n193 VTAIL.n182 171.744
R228 VTAIL.n193 VTAIL.n192 171.744
R229 VTAIL.n192 VTAIL.n186 171.744
R230 VTAIL.n166 VTAIL.n165 171.744
R231 VTAIL.n165 VTAIL.n164 171.744
R232 VTAIL.n164 VTAIL.n133 171.744
R233 VTAIL.n157 VTAIL.n133 171.744
R234 VTAIL.n157 VTAIL.n156 171.744
R235 VTAIL.n156 VTAIL.n138 171.744
R236 VTAIL.n149 VTAIL.n138 171.744
R237 VTAIL.n149 VTAIL.n148 171.744
R238 VTAIL.n148 VTAIL.n142 171.744
R239 VTAIL.t1 VTAIL.n313 85.8723
R240 VTAIL.t3 VTAIL.n13 85.8723
R241 VTAIL.t10 VTAIL.n55 85.8723
R242 VTAIL.t8 VTAIL.n99 85.8723
R243 VTAIL.t14 VTAIL.n272 85.8723
R244 VTAIL.t12 VTAIL.n228 85.8723
R245 VTAIL.t2 VTAIL.n186 85.8723
R246 VTAIL.t5 VTAIL.n142 85.8723
R247 VTAIL.n259 VTAIL.n258 69.7532
R248 VTAIL.n173 VTAIL.n172 69.7532
R249 VTAIL.n1 VTAIL.n0 69.753
R250 VTAIL.n87 VTAIL.n86 69.753
R251 VTAIL.n343 VTAIL.n342 36.2581
R252 VTAIL.n43 VTAIL.n42 36.2581
R253 VTAIL.n85 VTAIL.n84 36.2581
R254 VTAIL.n129 VTAIL.n128 36.2581
R255 VTAIL.n301 VTAIL.n300 36.2581
R256 VTAIL.n257 VTAIL.n256 36.2581
R257 VTAIL.n215 VTAIL.n214 36.2581
R258 VTAIL.n171 VTAIL.n170 36.2581
R259 VTAIL.n343 VTAIL.n301 20.591
R260 VTAIL.n171 VTAIL.n129 20.591
R261 VTAIL.n339 VTAIL.n304 13.1884
R262 VTAIL.n39 VTAIL.n4 13.1884
R263 VTAIL.n81 VTAIL.n46 13.1884
R264 VTAIL.n125 VTAIL.n90 13.1884
R265 VTAIL.n297 VTAIL.n262 13.1884
R266 VTAIL.n253 VTAIL.n218 13.1884
R267 VTAIL.n211 VTAIL.n176 13.1884
R268 VTAIL.n167 VTAIL.n132 13.1884
R269 VTAIL.n335 VTAIL.n334 12.8005
R270 VTAIL.n340 VTAIL.n302 12.8005
R271 VTAIL.n35 VTAIL.n34 12.8005
R272 VTAIL.n40 VTAIL.n2 12.8005
R273 VTAIL.n77 VTAIL.n76 12.8005
R274 VTAIL.n82 VTAIL.n44 12.8005
R275 VTAIL.n121 VTAIL.n120 12.8005
R276 VTAIL.n126 VTAIL.n88 12.8005
R277 VTAIL.n298 VTAIL.n260 12.8005
R278 VTAIL.n293 VTAIL.n264 12.8005
R279 VTAIL.n254 VTAIL.n216 12.8005
R280 VTAIL.n249 VTAIL.n220 12.8005
R281 VTAIL.n212 VTAIL.n174 12.8005
R282 VTAIL.n207 VTAIL.n178 12.8005
R283 VTAIL.n168 VTAIL.n130 12.8005
R284 VTAIL.n163 VTAIL.n134 12.8005
R285 VTAIL.n333 VTAIL.n306 12.0247
R286 VTAIL.n33 VTAIL.n6 12.0247
R287 VTAIL.n75 VTAIL.n48 12.0247
R288 VTAIL.n119 VTAIL.n92 12.0247
R289 VTAIL.n292 VTAIL.n265 12.0247
R290 VTAIL.n248 VTAIL.n221 12.0247
R291 VTAIL.n206 VTAIL.n179 12.0247
R292 VTAIL.n162 VTAIL.n135 12.0247
R293 VTAIL.n330 VTAIL.n329 11.249
R294 VTAIL.n30 VTAIL.n29 11.249
R295 VTAIL.n72 VTAIL.n71 11.249
R296 VTAIL.n116 VTAIL.n115 11.249
R297 VTAIL.n289 VTAIL.n288 11.249
R298 VTAIL.n245 VTAIL.n244 11.249
R299 VTAIL.n203 VTAIL.n202 11.249
R300 VTAIL.n159 VTAIL.n158 11.249
R301 VTAIL.n315 VTAIL.n314 10.7238
R302 VTAIL.n15 VTAIL.n14 10.7238
R303 VTAIL.n57 VTAIL.n56 10.7238
R304 VTAIL.n101 VTAIL.n100 10.7238
R305 VTAIL.n274 VTAIL.n273 10.7238
R306 VTAIL.n230 VTAIL.n229 10.7238
R307 VTAIL.n188 VTAIL.n187 10.7238
R308 VTAIL.n144 VTAIL.n143 10.7238
R309 VTAIL.n326 VTAIL.n308 10.4732
R310 VTAIL.n26 VTAIL.n8 10.4732
R311 VTAIL.n68 VTAIL.n50 10.4732
R312 VTAIL.n112 VTAIL.n94 10.4732
R313 VTAIL.n285 VTAIL.n267 10.4732
R314 VTAIL.n241 VTAIL.n223 10.4732
R315 VTAIL.n199 VTAIL.n181 10.4732
R316 VTAIL.n155 VTAIL.n137 10.4732
R317 VTAIL.n325 VTAIL.n310 9.69747
R318 VTAIL.n25 VTAIL.n10 9.69747
R319 VTAIL.n67 VTAIL.n52 9.69747
R320 VTAIL.n111 VTAIL.n96 9.69747
R321 VTAIL.n284 VTAIL.n269 9.69747
R322 VTAIL.n240 VTAIL.n225 9.69747
R323 VTAIL.n198 VTAIL.n183 9.69747
R324 VTAIL.n154 VTAIL.n139 9.69747
R325 VTAIL.n342 VTAIL.n341 9.45567
R326 VTAIL.n42 VTAIL.n41 9.45567
R327 VTAIL.n84 VTAIL.n83 9.45567
R328 VTAIL.n128 VTAIL.n127 9.45567
R329 VTAIL.n300 VTAIL.n299 9.45567
R330 VTAIL.n256 VTAIL.n255 9.45567
R331 VTAIL.n214 VTAIL.n213 9.45567
R332 VTAIL.n170 VTAIL.n169 9.45567
R333 VTAIL.n341 VTAIL.n340 9.3005
R334 VTAIL.n317 VTAIL.n316 9.3005
R335 VTAIL.n312 VTAIL.n311 9.3005
R336 VTAIL.n323 VTAIL.n322 9.3005
R337 VTAIL.n325 VTAIL.n324 9.3005
R338 VTAIL.n308 VTAIL.n307 9.3005
R339 VTAIL.n331 VTAIL.n330 9.3005
R340 VTAIL.n333 VTAIL.n332 9.3005
R341 VTAIL.n334 VTAIL.n303 9.3005
R342 VTAIL.n41 VTAIL.n40 9.3005
R343 VTAIL.n17 VTAIL.n16 9.3005
R344 VTAIL.n12 VTAIL.n11 9.3005
R345 VTAIL.n23 VTAIL.n22 9.3005
R346 VTAIL.n25 VTAIL.n24 9.3005
R347 VTAIL.n8 VTAIL.n7 9.3005
R348 VTAIL.n31 VTAIL.n30 9.3005
R349 VTAIL.n33 VTAIL.n32 9.3005
R350 VTAIL.n34 VTAIL.n3 9.3005
R351 VTAIL.n83 VTAIL.n82 9.3005
R352 VTAIL.n59 VTAIL.n58 9.3005
R353 VTAIL.n54 VTAIL.n53 9.3005
R354 VTAIL.n65 VTAIL.n64 9.3005
R355 VTAIL.n67 VTAIL.n66 9.3005
R356 VTAIL.n50 VTAIL.n49 9.3005
R357 VTAIL.n73 VTAIL.n72 9.3005
R358 VTAIL.n75 VTAIL.n74 9.3005
R359 VTAIL.n76 VTAIL.n45 9.3005
R360 VTAIL.n127 VTAIL.n126 9.3005
R361 VTAIL.n103 VTAIL.n102 9.3005
R362 VTAIL.n98 VTAIL.n97 9.3005
R363 VTAIL.n109 VTAIL.n108 9.3005
R364 VTAIL.n111 VTAIL.n110 9.3005
R365 VTAIL.n94 VTAIL.n93 9.3005
R366 VTAIL.n117 VTAIL.n116 9.3005
R367 VTAIL.n119 VTAIL.n118 9.3005
R368 VTAIL.n120 VTAIL.n89 9.3005
R369 VTAIL.n276 VTAIL.n275 9.3005
R370 VTAIL.n271 VTAIL.n270 9.3005
R371 VTAIL.n282 VTAIL.n281 9.3005
R372 VTAIL.n284 VTAIL.n283 9.3005
R373 VTAIL.n267 VTAIL.n266 9.3005
R374 VTAIL.n290 VTAIL.n289 9.3005
R375 VTAIL.n292 VTAIL.n291 9.3005
R376 VTAIL.n264 VTAIL.n261 9.3005
R377 VTAIL.n299 VTAIL.n298 9.3005
R378 VTAIL.n232 VTAIL.n231 9.3005
R379 VTAIL.n227 VTAIL.n226 9.3005
R380 VTAIL.n238 VTAIL.n237 9.3005
R381 VTAIL.n240 VTAIL.n239 9.3005
R382 VTAIL.n223 VTAIL.n222 9.3005
R383 VTAIL.n246 VTAIL.n245 9.3005
R384 VTAIL.n248 VTAIL.n247 9.3005
R385 VTAIL.n220 VTAIL.n217 9.3005
R386 VTAIL.n255 VTAIL.n254 9.3005
R387 VTAIL.n190 VTAIL.n189 9.3005
R388 VTAIL.n185 VTAIL.n184 9.3005
R389 VTAIL.n196 VTAIL.n195 9.3005
R390 VTAIL.n198 VTAIL.n197 9.3005
R391 VTAIL.n181 VTAIL.n180 9.3005
R392 VTAIL.n204 VTAIL.n203 9.3005
R393 VTAIL.n206 VTAIL.n205 9.3005
R394 VTAIL.n178 VTAIL.n175 9.3005
R395 VTAIL.n213 VTAIL.n212 9.3005
R396 VTAIL.n146 VTAIL.n145 9.3005
R397 VTAIL.n141 VTAIL.n140 9.3005
R398 VTAIL.n152 VTAIL.n151 9.3005
R399 VTAIL.n154 VTAIL.n153 9.3005
R400 VTAIL.n137 VTAIL.n136 9.3005
R401 VTAIL.n160 VTAIL.n159 9.3005
R402 VTAIL.n162 VTAIL.n161 9.3005
R403 VTAIL.n134 VTAIL.n131 9.3005
R404 VTAIL.n169 VTAIL.n168 9.3005
R405 VTAIL.n322 VTAIL.n321 8.92171
R406 VTAIL.n22 VTAIL.n21 8.92171
R407 VTAIL.n64 VTAIL.n63 8.92171
R408 VTAIL.n108 VTAIL.n107 8.92171
R409 VTAIL.n281 VTAIL.n280 8.92171
R410 VTAIL.n237 VTAIL.n236 8.92171
R411 VTAIL.n195 VTAIL.n194 8.92171
R412 VTAIL.n151 VTAIL.n150 8.92171
R413 VTAIL.n318 VTAIL.n312 8.14595
R414 VTAIL.n18 VTAIL.n12 8.14595
R415 VTAIL.n60 VTAIL.n54 8.14595
R416 VTAIL.n104 VTAIL.n98 8.14595
R417 VTAIL.n277 VTAIL.n271 8.14595
R418 VTAIL.n233 VTAIL.n227 8.14595
R419 VTAIL.n191 VTAIL.n185 8.14595
R420 VTAIL.n147 VTAIL.n141 8.14595
R421 VTAIL.n317 VTAIL.n314 7.3702
R422 VTAIL.n17 VTAIL.n14 7.3702
R423 VTAIL.n59 VTAIL.n56 7.3702
R424 VTAIL.n103 VTAIL.n100 7.3702
R425 VTAIL.n276 VTAIL.n273 7.3702
R426 VTAIL.n232 VTAIL.n229 7.3702
R427 VTAIL.n190 VTAIL.n187 7.3702
R428 VTAIL.n146 VTAIL.n143 7.3702
R429 VTAIL.n318 VTAIL.n317 5.81868
R430 VTAIL.n18 VTAIL.n17 5.81868
R431 VTAIL.n60 VTAIL.n59 5.81868
R432 VTAIL.n104 VTAIL.n103 5.81868
R433 VTAIL.n277 VTAIL.n276 5.81868
R434 VTAIL.n233 VTAIL.n232 5.81868
R435 VTAIL.n191 VTAIL.n190 5.81868
R436 VTAIL.n147 VTAIL.n146 5.81868
R437 VTAIL.n321 VTAIL.n312 5.04292
R438 VTAIL.n21 VTAIL.n12 5.04292
R439 VTAIL.n63 VTAIL.n54 5.04292
R440 VTAIL.n107 VTAIL.n98 5.04292
R441 VTAIL.n280 VTAIL.n271 5.04292
R442 VTAIL.n236 VTAIL.n227 5.04292
R443 VTAIL.n194 VTAIL.n185 5.04292
R444 VTAIL.n150 VTAIL.n141 5.04292
R445 VTAIL.n322 VTAIL.n310 4.26717
R446 VTAIL.n22 VTAIL.n10 4.26717
R447 VTAIL.n64 VTAIL.n52 4.26717
R448 VTAIL.n108 VTAIL.n96 4.26717
R449 VTAIL.n281 VTAIL.n269 4.26717
R450 VTAIL.n237 VTAIL.n225 4.26717
R451 VTAIL.n195 VTAIL.n183 4.26717
R452 VTAIL.n151 VTAIL.n139 4.26717
R453 VTAIL.n0 VTAIL.t0 4.05855
R454 VTAIL.n0 VTAIL.t6 4.05855
R455 VTAIL.n86 VTAIL.t13 4.05855
R456 VTAIL.n86 VTAIL.t11 4.05855
R457 VTAIL.n258 VTAIL.t9 4.05855
R458 VTAIL.n258 VTAIL.t15 4.05855
R459 VTAIL.n172 VTAIL.t4 4.05855
R460 VTAIL.n172 VTAIL.t7 4.05855
R461 VTAIL.n326 VTAIL.n325 3.49141
R462 VTAIL.n26 VTAIL.n25 3.49141
R463 VTAIL.n68 VTAIL.n67 3.49141
R464 VTAIL.n112 VTAIL.n111 3.49141
R465 VTAIL.n285 VTAIL.n284 3.49141
R466 VTAIL.n241 VTAIL.n240 3.49141
R467 VTAIL.n199 VTAIL.n198 3.49141
R468 VTAIL.n155 VTAIL.n154 3.49141
R469 VTAIL.n329 VTAIL.n308 2.71565
R470 VTAIL.n29 VTAIL.n8 2.71565
R471 VTAIL.n71 VTAIL.n50 2.71565
R472 VTAIL.n115 VTAIL.n94 2.71565
R473 VTAIL.n288 VTAIL.n267 2.71565
R474 VTAIL.n244 VTAIL.n223 2.71565
R475 VTAIL.n202 VTAIL.n181 2.71565
R476 VTAIL.n158 VTAIL.n137 2.71565
R477 VTAIL.n316 VTAIL.n315 2.4129
R478 VTAIL.n16 VTAIL.n15 2.4129
R479 VTAIL.n58 VTAIL.n57 2.4129
R480 VTAIL.n102 VTAIL.n101 2.4129
R481 VTAIL.n275 VTAIL.n274 2.4129
R482 VTAIL.n231 VTAIL.n230 2.4129
R483 VTAIL.n189 VTAIL.n188 2.4129
R484 VTAIL.n145 VTAIL.n144 2.4129
R485 VTAIL.n330 VTAIL.n306 1.93989
R486 VTAIL.n30 VTAIL.n6 1.93989
R487 VTAIL.n72 VTAIL.n48 1.93989
R488 VTAIL.n116 VTAIL.n92 1.93989
R489 VTAIL.n289 VTAIL.n265 1.93989
R490 VTAIL.n245 VTAIL.n221 1.93989
R491 VTAIL.n203 VTAIL.n179 1.93989
R492 VTAIL.n159 VTAIL.n135 1.93989
R493 VTAIL.n173 VTAIL.n171 1.31947
R494 VTAIL.n215 VTAIL.n173 1.31947
R495 VTAIL.n259 VTAIL.n257 1.31947
R496 VTAIL.n301 VTAIL.n259 1.31947
R497 VTAIL.n129 VTAIL.n87 1.31947
R498 VTAIL.n87 VTAIL.n85 1.31947
R499 VTAIL.n43 VTAIL.n1 1.31947
R500 VTAIL VTAIL.n343 1.26128
R501 VTAIL.n335 VTAIL.n333 1.16414
R502 VTAIL.n342 VTAIL.n302 1.16414
R503 VTAIL.n35 VTAIL.n33 1.16414
R504 VTAIL.n42 VTAIL.n2 1.16414
R505 VTAIL.n77 VTAIL.n75 1.16414
R506 VTAIL.n84 VTAIL.n44 1.16414
R507 VTAIL.n121 VTAIL.n119 1.16414
R508 VTAIL.n128 VTAIL.n88 1.16414
R509 VTAIL.n300 VTAIL.n260 1.16414
R510 VTAIL.n293 VTAIL.n292 1.16414
R511 VTAIL.n256 VTAIL.n216 1.16414
R512 VTAIL.n249 VTAIL.n248 1.16414
R513 VTAIL.n214 VTAIL.n174 1.16414
R514 VTAIL.n207 VTAIL.n206 1.16414
R515 VTAIL.n170 VTAIL.n130 1.16414
R516 VTAIL.n163 VTAIL.n162 1.16414
R517 VTAIL.n257 VTAIL.n215 0.470328
R518 VTAIL.n85 VTAIL.n43 0.470328
R519 VTAIL.n334 VTAIL.n304 0.388379
R520 VTAIL.n340 VTAIL.n339 0.388379
R521 VTAIL.n34 VTAIL.n4 0.388379
R522 VTAIL.n40 VTAIL.n39 0.388379
R523 VTAIL.n76 VTAIL.n46 0.388379
R524 VTAIL.n82 VTAIL.n81 0.388379
R525 VTAIL.n120 VTAIL.n90 0.388379
R526 VTAIL.n126 VTAIL.n125 0.388379
R527 VTAIL.n298 VTAIL.n297 0.388379
R528 VTAIL.n264 VTAIL.n262 0.388379
R529 VTAIL.n254 VTAIL.n253 0.388379
R530 VTAIL.n220 VTAIL.n218 0.388379
R531 VTAIL.n212 VTAIL.n211 0.388379
R532 VTAIL.n178 VTAIL.n176 0.388379
R533 VTAIL.n168 VTAIL.n167 0.388379
R534 VTAIL.n134 VTAIL.n132 0.388379
R535 VTAIL.n316 VTAIL.n311 0.155672
R536 VTAIL.n323 VTAIL.n311 0.155672
R537 VTAIL.n324 VTAIL.n323 0.155672
R538 VTAIL.n324 VTAIL.n307 0.155672
R539 VTAIL.n331 VTAIL.n307 0.155672
R540 VTAIL.n332 VTAIL.n331 0.155672
R541 VTAIL.n332 VTAIL.n303 0.155672
R542 VTAIL.n341 VTAIL.n303 0.155672
R543 VTAIL.n16 VTAIL.n11 0.155672
R544 VTAIL.n23 VTAIL.n11 0.155672
R545 VTAIL.n24 VTAIL.n23 0.155672
R546 VTAIL.n24 VTAIL.n7 0.155672
R547 VTAIL.n31 VTAIL.n7 0.155672
R548 VTAIL.n32 VTAIL.n31 0.155672
R549 VTAIL.n32 VTAIL.n3 0.155672
R550 VTAIL.n41 VTAIL.n3 0.155672
R551 VTAIL.n58 VTAIL.n53 0.155672
R552 VTAIL.n65 VTAIL.n53 0.155672
R553 VTAIL.n66 VTAIL.n65 0.155672
R554 VTAIL.n66 VTAIL.n49 0.155672
R555 VTAIL.n73 VTAIL.n49 0.155672
R556 VTAIL.n74 VTAIL.n73 0.155672
R557 VTAIL.n74 VTAIL.n45 0.155672
R558 VTAIL.n83 VTAIL.n45 0.155672
R559 VTAIL.n102 VTAIL.n97 0.155672
R560 VTAIL.n109 VTAIL.n97 0.155672
R561 VTAIL.n110 VTAIL.n109 0.155672
R562 VTAIL.n110 VTAIL.n93 0.155672
R563 VTAIL.n117 VTAIL.n93 0.155672
R564 VTAIL.n118 VTAIL.n117 0.155672
R565 VTAIL.n118 VTAIL.n89 0.155672
R566 VTAIL.n127 VTAIL.n89 0.155672
R567 VTAIL.n299 VTAIL.n261 0.155672
R568 VTAIL.n291 VTAIL.n261 0.155672
R569 VTAIL.n291 VTAIL.n290 0.155672
R570 VTAIL.n290 VTAIL.n266 0.155672
R571 VTAIL.n283 VTAIL.n266 0.155672
R572 VTAIL.n283 VTAIL.n282 0.155672
R573 VTAIL.n282 VTAIL.n270 0.155672
R574 VTAIL.n275 VTAIL.n270 0.155672
R575 VTAIL.n255 VTAIL.n217 0.155672
R576 VTAIL.n247 VTAIL.n217 0.155672
R577 VTAIL.n247 VTAIL.n246 0.155672
R578 VTAIL.n246 VTAIL.n222 0.155672
R579 VTAIL.n239 VTAIL.n222 0.155672
R580 VTAIL.n239 VTAIL.n238 0.155672
R581 VTAIL.n238 VTAIL.n226 0.155672
R582 VTAIL.n231 VTAIL.n226 0.155672
R583 VTAIL.n213 VTAIL.n175 0.155672
R584 VTAIL.n205 VTAIL.n175 0.155672
R585 VTAIL.n205 VTAIL.n204 0.155672
R586 VTAIL.n204 VTAIL.n180 0.155672
R587 VTAIL.n197 VTAIL.n180 0.155672
R588 VTAIL.n197 VTAIL.n196 0.155672
R589 VTAIL.n196 VTAIL.n184 0.155672
R590 VTAIL.n189 VTAIL.n184 0.155672
R591 VTAIL.n169 VTAIL.n131 0.155672
R592 VTAIL.n161 VTAIL.n131 0.155672
R593 VTAIL.n161 VTAIL.n160 0.155672
R594 VTAIL.n160 VTAIL.n136 0.155672
R595 VTAIL.n153 VTAIL.n136 0.155672
R596 VTAIL.n153 VTAIL.n152 0.155672
R597 VTAIL.n152 VTAIL.n140 0.155672
R598 VTAIL.n145 VTAIL.n140 0.155672
R599 VTAIL VTAIL.n1 0.0586897
R600 B.n288 B.n87 585
R601 B.n287 B.n286 585
R602 B.n285 B.n88 585
R603 B.n284 B.n283 585
R604 B.n282 B.n89 585
R605 B.n281 B.n280 585
R606 B.n279 B.n90 585
R607 B.n278 B.n277 585
R608 B.n276 B.n91 585
R609 B.n275 B.n274 585
R610 B.n273 B.n92 585
R611 B.n272 B.n271 585
R612 B.n270 B.n93 585
R613 B.n269 B.n268 585
R614 B.n267 B.n94 585
R615 B.n266 B.n265 585
R616 B.n264 B.n95 585
R617 B.n263 B.n262 585
R618 B.n261 B.n96 585
R619 B.n260 B.n259 585
R620 B.n258 B.n97 585
R621 B.n257 B.n256 585
R622 B.n255 B.n98 585
R623 B.n254 B.n253 585
R624 B.n252 B.n99 585
R625 B.n251 B.n250 585
R626 B.n249 B.n100 585
R627 B.n248 B.n247 585
R628 B.n246 B.n101 585
R629 B.n245 B.n244 585
R630 B.n243 B.n242 585
R631 B.n241 B.n105 585
R632 B.n240 B.n239 585
R633 B.n238 B.n106 585
R634 B.n237 B.n236 585
R635 B.n235 B.n107 585
R636 B.n234 B.n233 585
R637 B.n232 B.n108 585
R638 B.n231 B.n230 585
R639 B.n228 B.n109 585
R640 B.n227 B.n226 585
R641 B.n225 B.n112 585
R642 B.n224 B.n223 585
R643 B.n222 B.n113 585
R644 B.n221 B.n220 585
R645 B.n219 B.n114 585
R646 B.n218 B.n217 585
R647 B.n216 B.n115 585
R648 B.n215 B.n214 585
R649 B.n213 B.n116 585
R650 B.n212 B.n211 585
R651 B.n210 B.n117 585
R652 B.n209 B.n208 585
R653 B.n207 B.n118 585
R654 B.n206 B.n205 585
R655 B.n204 B.n119 585
R656 B.n203 B.n202 585
R657 B.n201 B.n120 585
R658 B.n200 B.n199 585
R659 B.n198 B.n121 585
R660 B.n197 B.n196 585
R661 B.n195 B.n122 585
R662 B.n194 B.n193 585
R663 B.n192 B.n123 585
R664 B.n191 B.n190 585
R665 B.n189 B.n124 585
R666 B.n188 B.n187 585
R667 B.n186 B.n125 585
R668 B.n185 B.n184 585
R669 B.n290 B.n289 585
R670 B.n291 B.n86 585
R671 B.n293 B.n292 585
R672 B.n294 B.n85 585
R673 B.n296 B.n295 585
R674 B.n297 B.n84 585
R675 B.n299 B.n298 585
R676 B.n300 B.n83 585
R677 B.n302 B.n301 585
R678 B.n303 B.n82 585
R679 B.n305 B.n304 585
R680 B.n306 B.n81 585
R681 B.n308 B.n307 585
R682 B.n309 B.n80 585
R683 B.n311 B.n310 585
R684 B.n312 B.n79 585
R685 B.n314 B.n313 585
R686 B.n315 B.n78 585
R687 B.n317 B.n316 585
R688 B.n318 B.n77 585
R689 B.n320 B.n319 585
R690 B.n321 B.n76 585
R691 B.n323 B.n322 585
R692 B.n324 B.n75 585
R693 B.n326 B.n325 585
R694 B.n327 B.n74 585
R695 B.n329 B.n328 585
R696 B.n330 B.n73 585
R697 B.n332 B.n331 585
R698 B.n333 B.n72 585
R699 B.n335 B.n334 585
R700 B.n336 B.n71 585
R701 B.n338 B.n337 585
R702 B.n339 B.n70 585
R703 B.n341 B.n340 585
R704 B.n342 B.n69 585
R705 B.n344 B.n343 585
R706 B.n345 B.n68 585
R707 B.n347 B.n346 585
R708 B.n348 B.n67 585
R709 B.n350 B.n349 585
R710 B.n351 B.n66 585
R711 B.n353 B.n352 585
R712 B.n354 B.n65 585
R713 B.n356 B.n355 585
R714 B.n357 B.n64 585
R715 B.n359 B.n358 585
R716 B.n360 B.n63 585
R717 B.n362 B.n361 585
R718 B.n363 B.n62 585
R719 B.n365 B.n364 585
R720 B.n366 B.n61 585
R721 B.n368 B.n367 585
R722 B.n369 B.n60 585
R723 B.n371 B.n370 585
R724 B.n372 B.n59 585
R725 B.n374 B.n373 585
R726 B.n375 B.n58 585
R727 B.n377 B.n376 585
R728 B.n378 B.n57 585
R729 B.n380 B.n379 585
R730 B.n381 B.n56 585
R731 B.n486 B.n17 585
R732 B.n485 B.n484 585
R733 B.n483 B.n18 585
R734 B.n482 B.n481 585
R735 B.n480 B.n19 585
R736 B.n479 B.n478 585
R737 B.n477 B.n20 585
R738 B.n476 B.n475 585
R739 B.n474 B.n21 585
R740 B.n473 B.n472 585
R741 B.n471 B.n22 585
R742 B.n470 B.n469 585
R743 B.n468 B.n23 585
R744 B.n467 B.n466 585
R745 B.n465 B.n24 585
R746 B.n464 B.n463 585
R747 B.n462 B.n25 585
R748 B.n461 B.n460 585
R749 B.n459 B.n26 585
R750 B.n458 B.n457 585
R751 B.n456 B.n27 585
R752 B.n455 B.n454 585
R753 B.n453 B.n28 585
R754 B.n452 B.n451 585
R755 B.n450 B.n29 585
R756 B.n449 B.n448 585
R757 B.n447 B.n30 585
R758 B.n446 B.n445 585
R759 B.n444 B.n31 585
R760 B.n443 B.n442 585
R761 B.n441 B.n440 585
R762 B.n439 B.n35 585
R763 B.n438 B.n437 585
R764 B.n436 B.n36 585
R765 B.n435 B.n434 585
R766 B.n433 B.n37 585
R767 B.n432 B.n431 585
R768 B.n430 B.n38 585
R769 B.n429 B.n428 585
R770 B.n426 B.n39 585
R771 B.n425 B.n424 585
R772 B.n423 B.n42 585
R773 B.n422 B.n421 585
R774 B.n420 B.n43 585
R775 B.n419 B.n418 585
R776 B.n417 B.n44 585
R777 B.n416 B.n415 585
R778 B.n414 B.n45 585
R779 B.n413 B.n412 585
R780 B.n411 B.n46 585
R781 B.n410 B.n409 585
R782 B.n408 B.n47 585
R783 B.n407 B.n406 585
R784 B.n405 B.n48 585
R785 B.n404 B.n403 585
R786 B.n402 B.n49 585
R787 B.n401 B.n400 585
R788 B.n399 B.n50 585
R789 B.n398 B.n397 585
R790 B.n396 B.n51 585
R791 B.n395 B.n394 585
R792 B.n393 B.n52 585
R793 B.n392 B.n391 585
R794 B.n390 B.n53 585
R795 B.n389 B.n388 585
R796 B.n387 B.n54 585
R797 B.n386 B.n385 585
R798 B.n384 B.n55 585
R799 B.n383 B.n382 585
R800 B.n488 B.n487 585
R801 B.n489 B.n16 585
R802 B.n491 B.n490 585
R803 B.n492 B.n15 585
R804 B.n494 B.n493 585
R805 B.n495 B.n14 585
R806 B.n497 B.n496 585
R807 B.n498 B.n13 585
R808 B.n500 B.n499 585
R809 B.n501 B.n12 585
R810 B.n503 B.n502 585
R811 B.n504 B.n11 585
R812 B.n506 B.n505 585
R813 B.n507 B.n10 585
R814 B.n509 B.n508 585
R815 B.n510 B.n9 585
R816 B.n512 B.n511 585
R817 B.n513 B.n8 585
R818 B.n515 B.n514 585
R819 B.n516 B.n7 585
R820 B.n518 B.n517 585
R821 B.n519 B.n6 585
R822 B.n521 B.n520 585
R823 B.n522 B.n5 585
R824 B.n524 B.n523 585
R825 B.n525 B.n4 585
R826 B.n527 B.n526 585
R827 B.n528 B.n3 585
R828 B.n530 B.n529 585
R829 B.n531 B.n0 585
R830 B.n2 B.n1 585
R831 B.n141 B.n140 585
R832 B.n143 B.n142 585
R833 B.n144 B.n139 585
R834 B.n146 B.n145 585
R835 B.n147 B.n138 585
R836 B.n149 B.n148 585
R837 B.n150 B.n137 585
R838 B.n152 B.n151 585
R839 B.n153 B.n136 585
R840 B.n155 B.n154 585
R841 B.n156 B.n135 585
R842 B.n158 B.n157 585
R843 B.n159 B.n134 585
R844 B.n161 B.n160 585
R845 B.n162 B.n133 585
R846 B.n164 B.n163 585
R847 B.n165 B.n132 585
R848 B.n167 B.n166 585
R849 B.n168 B.n131 585
R850 B.n170 B.n169 585
R851 B.n171 B.n130 585
R852 B.n173 B.n172 585
R853 B.n174 B.n129 585
R854 B.n176 B.n175 585
R855 B.n177 B.n128 585
R856 B.n179 B.n178 585
R857 B.n180 B.n127 585
R858 B.n182 B.n181 585
R859 B.n183 B.n126 585
R860 B.n184 B.n183 545.355
R861 B.n290 B.n87 545.355
R862 B.n382 B.n381 545.355
R863 B.n488 B.n17 545.355
R864 B.n110 B.t9 364.985
R865 B.n102 B.t6 364.985
R866 B.n40 B.t0 364.985
R867 B.n32 B.t3 364.985
R868 B.n102 B.t7 333.557
R869 B.n40 B.t2 333.557
R870 B.n110 B.t10 333.557
R871 B.n32 B.t5 333.557
R872 B.n103 B.t8 303.885
R873 B.n41 B.t1 303.885
R874 B.n111 B.t11 303.885
R875 B.n33 B.t4 303.885
R876 B.n533 B.n532 256.663
R877 B.n532 B.n531 235.042
R878 B.n532 B.n2 235.042
R879 B.n184 B.n125 163.367
R880 B.n188 B.n125 163.367
R881 B.n189 B.n188 163.367
R882 B.n190 B.n189 163.367
R883 B.n190 B.n123 163.367
R884 B.n194 B.n123 163.367
R885 B.n195 B.n194 163.367
R886 B.n196 B.n195 163.367
R887 B.n196 B.n121 163.367
R888 B.n200 B.n121 163.367
R889 B.n201 B.n200 163.367
R890 B.n202 B.n201 163.367
R891 B.n202 B.n119 163.367
R892 B.n206 B.n119 163.367
R893 B.n207 B.n206 163.367
R894 B.n208 B.n207 163.367
R895 B.n208 B.n117 163.367
R896 B.n212 B.n117 163.367
R897 B.n213 B.n212 163.367
R898 B.n214 B.n213 163.367
R899 B.n214 B.n115 163.367
R900 B.n218 B.n115 163.367
R901 B.n219 B.n218 163.367
R902 B.n220 B.n219 163.367
R903 B.n220 B.n113 163.367
R904 B.n224 B.n113 163.367
R905 B.n225 B.n224 163.367
R906 B.n226 B.n225 163.367
R907 B.n226 B.n109 163.367
R908 B.n231 B.n109 163.367
R909 B.n232 B.n231 163.367
R910 B.n233 B.n232 163.367
R911 B.n233 B.n107 163.367
R912 B.n237 B.n107 163.367
R913 B.n238 B.n237 163.367
R914 B.n239 B.n238 163.367
R915 B.n239 B.n105 163.367
R916 B.n243 B.n105 163.367
R917 B.n244 B.n243 163.367
R918 B.n244 B.n101 163.367
R919 B.n248 B.n101 163.367
R920 B.n249 B.n248 163.367
R921 B.n250 B.n249 163.367
R922 B.n250 B.n99 163.367
R923 B.n254 B.n99 163.367
R924 B.n255 B.n254 163.367
R925 B.n256 B.n255 163.367
R926 B.n256 B.n97 163.367
R927 B.n260 B.n97 163.367
R928 B.n261 B.n260 163.367
R929 B.n262 B.n261 163.367
R930 B.n262 B.n95 163.367
R931 B.n266 B.n95 163.367
R932 B.n267 B.n266 163.367
R933 B.n268 B.n267 163.367
R934 B.n268 B.n93 163.367
R935 B.n272 B.n93 163.367
R936 B.n273 B.n272 163.367
R937 B.n274 B.n273 163.367
R938 B.n274 B.n91 163.367
R939 B.n278 B.n91 163.367
R940 B.n279 B.n278 163.367
R941 B.n280 B.n279 163.367
R942 B.n280 B.n89 163.367
R943 B.n284 B.n89 163.367
R944 B.n285 B.n284 163.367
R945 B.n286 B.n285 163.367
R946 B.n286 B.n87 163.367
R947 B.n381 B.n380 163.367
R948 B.n380 B.n57 163.367
R949 B.n376 B.n57 163.367
R950 B.n376 B.n375 163.367
R951 B.n375 B.n374 163.367
R952 B.n374 B.n59 163.367
R953 B.n370 B.n59 163.367
R954 B.n370 B.n369 163.367
R955 B.n369 B.n368 163.367
R956 B.n368 B.n61 163.367
R957 B.n364 B.n61 163.367
R958 B.n364 B.n363 163.367
R959 B.n363 B.n362 163.367
R960 B.n362 B.n63 163.367
R961 B.n358 B.n63 163.367
R962 B.n358 B.n357 163.367
R963 B.n357 B.n356 163.367
R964 B.n356 B.n65 163.367
R965 B.n352 B.n65 163.367
R966 B.n352 B.n351 163.367
R967 B.n351 B.n350 163.367
R968 B.n350 B.n67 163.367
R969 B.n346 B.n67 163.367
R970 B.n346 B.n345 163.367
R971 B.n345 B.n344 163.367
R972 B.n344 B.n69 163.367
R973 B.n340 B.n69 163.367
R974 B.n340 B.n339 163.367
R975 B.n339 B.n338 163.367
R976 B.n338 B.n71 163.367
R977 B.n334 B.n71 163.367
R978 B.n334 B.n333 163.367
R979 B.n333 B.n332 163.367
R980 B.n332 B.n73 163.367
R981 B.n328 B.n73 163.367
R982 B.n328 B.n327 163.367
R983 B.n327 B.n326 163.367
R984 B.n326 B.n75 163.367
R985 B.n322 B.n75 163.367
R986 B.n322 B.n321 163.367
R987 B.n321 B.n320 163.367
R988 B.n320 B.n77 163.367
R989 B.n316 B.n77 163.367
R990 B.n316 B.n315 163.367
R991 B.n315 B.n314 163.367
R992 B.n314 B.n79 163.367
R993 B.n310 B.n79 163.367
R994 B.n310 B.n309 163.367
R995 B.n309 B.n308 163.367
R996 B.n308 B.n81 163.367
R997 B.n304 B.n81 163.367
R998 B.n304 B.n303 163.367
R999 B.n303 B.n302 163.367
R1000 B.n302 B.n83 163.367
R1001 B.n298 B.n83 163.367
R1002 B.n298 B.n297 163.367
R1003 B.n297 B.n296 163.367
R1004 B.n296 B.n85 163.367
R1005 B.n292 B.n85 163.367
R1006 B.n292 B.n291 163.367
R1007 B.n291 B.n290 163.367
R1008 B.n484 B.n17 163.367
R1009 B.n484 B.n483 163.367
R1010 B.n483 B.n482 163.367
R1011 B.n482 B.n19 163.367
R1012 B.n478 B.n19 163.367
R1013 B.n478 B.n477 163.367
R1014 B.n477 B.n476 163.367
R1015 B.n476 B.n21 163.367
R1016 B.n472 B.n21 163.367
R1017 B.n472 B.n471 163.367
R1018 B.n471 B.n470 163.367
R1019 B.n470 B.n23 163.367
R1020 B.n466 B.n23 163.367
R1021 B.n466 B.n465 163.367
R1022 B.n465 B.n464 163.367
R1023 B.n464 B.n25 163.367
R1024 B.n460 B.n25 163.367
R1025 B.n460 B.n459 163.367
R1026 B.n459 B.n458 163.367
R1027 B.n458 B.n27 163.367
R1028 B.n454 B.n27 163.367
R1029 B.n454 B.n453 163.367
R1030 B.n453 B.n452 163.367
R1031 B.n452 B.n29 163.367
R1032 B.n448 B.n29 163.367
R1033 B.n448 B.n447 163.367
R1034 B.n447 B.n446 163.367
R1035 B.n446 B.n31 163.367
R1036 B.n442 B.n31 163.367
R1037 B.n442 B.n441 163.367
R1038 B.n441 B.n35 163.367
R1039 B.n437 B.n35 163.367
R1040 B.n437 B.n436 163.367
R1041 B.n436 B.n435 163.367
R1042 B.n435 B.n37 163.367
R1043 B.n431 B.n37 163.367
R1044 B.n431 B.n430 163.367
R1045 B.n430 B.n429 163.367
R1046 B.n429 B.n39 163.367
R1047 B.n424 B.n39 163.367
R1048 B.n424 B.n423 163.367
R1049 B.n423 B.n422 163.367
R1050 B.n422 B.n43 163.367
R1051 B.n418 B.n43 163.367
R1052 B.n418 B.n417 163.367
R1053 B.n417 B.n416 163.367
R1054 B.n416 B.n45 163.367
R1055 B.n412 B.n45 163.367
R1056 B.n412 B.n411 163.367
R1057 B.n411 B.n410 163.367
R1058 B.n410 B.n47 163.367
R1059 B.n406 B.n47 163.367
R1060 B.n406 B.n405 163.367
R1061 B.n405 B.n404 163.367
R1062 B.n404 B.n49 163.367
R1063 B.n400 B.n49 163.367
R1064 B.n400 B.n399 163.367
R1065 B.n399 B.n398 163.367
R1066 B.n398 B.n51 163.367
R1067 B.n394 B.n51 163.367
R1068 B.n394 B.n393 163.367
R1069 B.n393 B.n392 163.367
R1070 B.n392 B.n53 163.367
R1071 B.n388 B.n53 163.367
R1072 B.n388 B.n387 163.367
R1073 B.n387 B.n386 163.367
R1074 B.n386 B.n55 163.367
R1075 B.n382 B.n55 163.367
R1076 B.n489 B.n488 163.367
R1077 B.n490 B.n489 163.367
R1078 B.n490 B.n15 163.367
R1079 B.n494 B.n15 163.367
R1080 B.n495 B.n494 163.367
R1081 B.n496 B.n495 163.367
R1082 B.n496 B.n13 163.367
R1083 B.n500 B.n13 163.367
R1084 B.n501 B.n500 163.367
R1085 B.n502 B.n501 163.367
R1086 B.n502 B.n11 163.367
R1087 B.n506 B.n11 163.367
R1088 B.n507 B.n506 163.367
R1089 B.n508 B.n507 163.367
R1090 B.n508 B.n9 163.367
R1091 B.n512 B.n9 163.367
R1092 B.n513 B.n512 163.367
R1093 B.n514 B.n513 163.367
R1094 B.n514 B.n7 163.367
R1095 B.n518 B.n7 163.367
R1096 B.n519 B.n518 163.367
R1097 B.n520 B.n519 163.367
R1098 B.n520 B.n5 163.367
R1099 B.n524 B.n5 163.367
R1100 B.n525 B.n524 163.367
R1101 B.n526 B.n525 163.367
R1102 B.n526 B.n3 163.367
R1103 B.n530 B.n3 163.367
R1104 B.n531 B.n530 163.367
R1105 B.n141 B.n2 163.367
R1106 B.n142 B.n141 163.367
R1107 B.n142 B.n139 163.367
R1108 B.n146 B.n139 163.367
R1109 B.n147 B.n146 163.367
R1110 B.n148 B.n147 163.367
R1111 B.n148 B.n137 163.367
R1112 B.n152 B.n137 163.367
R1113 B.n153 B.n152 163.367
R1114 B.n154 B.n153 163.367
R1115 B.n154 B.n135 163.367
R1116 B.n158 B.n135 163.367
R1117 B.n159 B.n158 163.367
R1118 B.n160 B.n159 163.367
R1119 B.n160 B.n133 163.367
R1120 B.n164 B.n133 163.367
R1121 B.n165 B.n164 163.367
R1122 B.n166 B.n165 163.367
R1123 B.n166 B.n131 163.367
R1124 B.n170 B.n131 163.367
R1125 B.n171 B.n170 163.367
R1126 B.n172 B.n171 163.367
R1127 B.n172 B.n129 163.367
R1128 B.n176 B.n129 163.367
R1129 B.n177 B.n176 163.367
R1130 B.n178 B.n177 163.367
R1131 B.n178 B.n127 163.367
R1132 B.n182 B.n127 163.367
R1133 B.n183 B.n182 163.367
R1134 B.n229 B.n111 59.5399
R1135 B.n104 B.n103 59.5399
R1136 B.n427 B.n41 59.5399
R1137 B.n34 B.n33 59.5399
R1138 B.n487 B.n486 35.4346
R1139 B.n383 B.n56 35.4346
R1140 B.n185 B.n126 35.4346
R1141 B.n289 B.n288 35.4346
R1142 B.n111 B.n110 29.6732
R1143 B.n103 B.n102 29.6732
R1144 B.n41 B.n40 29.6732
R1145 B.n33 B.n32 29.6732
R1146 B B.n533 18.0485
R1147 B.n487 B.n16 10.6151
R1148 B.n491 B.n16 10.6151
R1149 B.n492 B.n491 10.6151
R1150 B.n493 B.n492 10.6151
R1151 B.n493 B.n14 10.6151
R1152 B.n497 B.n14 10.6151
R1153 B.n498 B.n497 10.6151
R1154 B.n499 B.n498 10.6151
R1155 B.n499 B.n12 10.6151
R1156 B.n503 B.n12 10.6151
R1157 B.n504 B.n503 10.6151
R1158 B.n505 B.n504 10.6151
R1159 B.n505 B.n10 10.6151
R1160 B.n509 B.n10 10.6151
R1161 B.n510 B.n509 10.6151
R1162 B.n511 B.n510 10.6151
R1163 B.n511 B.n8 10.6151
R1164 B.n515 B.n8 10.6151
R1165 B.n516 B.n515 10.6151
R1166 B.n517 B.n516 10.6151
R1167 B.n517 B.n6 10.6151
R1168 B.n521 B.n6 10.6151
R1169 B.n522 B.n521 10.6151
R1170 B.n523 B.n522 10.6151
R1171 B.n523 B.n4 10.6151
R1172 B.n527 B.n4 10.6151
R1173 B.n528 B.n527 10.6151
R1174 B.n529 B.n528 10.6151
R1175 B.n529 B.n0 10.6151
R1176 B.n486 B.n485 10.6151
R1177 B.n485 B.n18 10.6151
R1178 B.n481 B.n18 10.6151
R1179 B.n481 B.n480 10.6151
R1180 B.n480 B.n479 10.6151
R1181 B.n479 B.n20 10.6151
R1182 B.n475 B.n20 10.6151
R1183 B.n475 B.n474 10.6151
R1184 B.n474 B.n473 10.6151
R1185 B.n473 B.n22 10.6151
R1186 B.n469 B.n22 10.6151
R1187 B.n469 B.n468 10.6151
R1188 B.n468 B.n467 10.6151
R1189 B.n467 B.n24 10.6151
R1190 B.n463 B.n24 10.6151
R1191 B.n463 B.n462 10.6151
R1192 B.n462 B.n461 10.6151
R1193 B.n461 B.n26 10.6151
R1194 B.n457 B.n26 10.6151
R1195 B.n457 B.n456 10.6151
R1196 B.n456 B.n455 10.6151
R1197 B.n455 B.n28 10.6151
R1198 B.n451 B.n28 10.6151
R1199 B.n451 B.n450 10.6151
R1200 B.n450 B.n449 10.6151
R1201 B.n449 B.n30 10.6151
R1202 B.n445 B.n30 10.6151
R1203 B.n445 B.n444 10.6151
R1204 B.n444 B.n443 10.6151
R1205 B.n440 B.n439 10.6151
R1206 B.n439 B.n438 10.6151
R1207 B.n438 B.n36 10.6151
R1208 B.n434 B.n36 10.6151
R1209 B.n434 B.n433 10.6151
R1210 B.n433 B.n432 10.6151
R1211 B.n432 B.n38 10.6151
R1212 B.n428 B.n38 10.6151
R1213 B.n426 B.n425 10.6151
R1214 B.n425 B.n42 10.6151
R1215 B.n421 B.n42 10.6151
R1216 B.n421 B.n420 10.6151
R1217 B.n420 B.n419 10.6151
R1218 B.n419 B.n44 10.6151
R1219 B.n415 B.n44 10.6151
R1220 B.n415 B.n414 10.6151
R1221 B.n414 B.n413 10.6151
R1222 B.n413 B.n46 10.6151
R1223 B.n409 B.n46 10.6151
R1224 B.n409 B.n408 10.6151
R1225 B.n408 B.n407 10.6151
R1226 B.n407 B.n48 10.6151
R1227 B.n403 B.n48 10.6151
R1228 B.n403 B.n402 10.6151
R1229 B.n402 B.n401 10.6151
R1230 B.n401 B.n50 10.6151
R1231 B.n397 B.n50 10.6151
R1232 B.n397 B.n396 10.6151
R1233 B.n396 B.n395 10.6151
R1234 B.n395 B.n52 10.6151
R1235 B.n391 B.n52 10.6151
R1236 B.n391 B.n390 10.6151
R1237 B.n390 B.n389 10.6151
R1238 B.n389 B.n54 10.6151
R1239 B.n385 B.n54 10.6151
R1240 B.n385 B.n384 10.6151
R1241 B.n384 B.n383 10.6151
R1242 B.n379 B.n56 10.6151
R1243 B.n379 B.n378 10.6151
R1244 B.n378 B.n377 10.6151
R1245 B.n377 B.n58 10.6151
R1246 B.n373 B.n58 10.6151
R1247 B.n373 B.n372 10.6151
R1248 B.n372 B.n371 10.6151
R1249 B.n371 B.n60 10.6151
R1250 B.n367 B.n60 10.6151
R1251 B.n367 B.n366 10.6151
R1252 B.n366 B.n365 10.6151
R1253 B.n365 B.n62 10.6151
R1254 B.n361 B.n62 10.6151
R1255 B.n361 B.n360 10.6151
R1256 B.n360 B.n359 10.6151
R1257 B.n359 B.n64 10.6151
R1258 B.n355 B.n64 10.6151
R1259 B.n355 B.n354 10.6151
R1260 B.n354 B.n353 10.6151
R1261 B.n353 B.n66 10.6151
R1262 B.n349 B.n66 10.6151
R1263 B.n349 B.n348 10.6151
R1264 B.n348 B.n347 10.6151
R1265 B.n347 B.n68 10.6151
R1266 B.n343 B.n68 10.6151
R1267 B.n343 B.n342 10.6151
R1268 B.n342 B.n341 10.6151
R1269 B.n341 B.n70 10.6151
R1270 B.n337 B.n70 10.6151
R1271 B.n337 B.n336 10.6151
R1272 B.n336 B.n335 10.6151
R1273 B.n335 B.n72 10.6151
R1274 B.n331 B.n72 10.6151
R1275 B.n331 B.n330 10.6151
R1276 B.n330 B.n329 10.6151
R1277 B.n329 B.n74 10.6151
R1278 B.n325 B.n74 10.6151
R1279 B.n325 B.n324 10.6151
R1280 B.n324 B.n323 10.6151
R1281 B.n323 B.n76 10.6151
R1282 B.n319 B.n76 10.6151
R1283 B.n319 B.n318 10.6151
R1284 B.n318 B.n317 10.6151
R1285 B.n317 B.n78 10.6151
R1286 B.n313 B.n78 10.6151
R1287 B.n313 B.n312 10.6151
R1288 B.n312 B.n311 10.6151
R1289 B.n311 B.n80 10.6151
R1290 B.n307 B.n80 10.6151
R1291 B.n307 B.n306 10.6151
R1292 B.n306 B.n305 10.6151
R1293 B.n305 B.n82 10.6151
R1294 B.n301 B.n82 10.6151
R1295 B.n301 B.n300 10.6151
R1296 B.n300 B.n299 10.6151
R1297 B.n299 B.n84 10.6151
R1298 B.n295 B.n84 10.6151
R1299 B.n295 B.n294 10.6151
R1300 B.n294 B.n293 10.6151
R1301 B.n293 B.n86 10.6151
R1302 B.n289 B.n86 10.6151
R1303 B.n140 B.n1 10.6151
R1304 B.n143 B.n140 10.6151
R1305 B.n144 B.n143 10.6151
R1306 B.n145 B.n144 10.6151
R1307 B.n145 B.n138 10.6151
R1308 B.n149 B.n138 10.6151
R1309 B.n150 B.n149 10.6151
R1310 B.n151 B.n150 10.6151
R1311 B.n151 B.n136 10.6151
R1312 B.n155 B.n136 10.6151
R1313 B.n156 B.n155 10.6151
R1314 B.n157 B.n156 10.6151
R1315 B.n157 B.n134 10.6151
R1316 B.n161 B.n134 10.6151
R1317 B.n162 B.n161 10.6151
R1318 B.n163 B.n162 10.6151
R1319 B.n163 B.n132 10.6151
R1320 B.n167 B.n132 10.6151
R1321 B.n168 B.n167 10.6151
R1322 B.n169 B.n168 10.6151
R1323 B.n169 B.n130 10.6151
R1324 B.n173 B.n130 10.6151
R1325 B.n174 B.n173 10.6151
R1326 B.n175 B.n174 10.6151
R1327 B.n175 B.n128 10.6151
R1328 B.n179 B.n128 10.6151
R1329 B.n180 B.n179 10.6151
R1330 B.n181 B.n180 10.6151
R1331 B.n181 B.n126 10.6151
R1332 B.n186 B.n185 10.6151
R1333 B.n187 B.n186 10.6151
R1334 B.n187 B.n124 10.6151
R1335 B.n191 B.n124 10.6151
R1336 B.n192 B.n191 10.6151
R1337 B.n193 B.n192 10.6151
R1338 B.n193 B.n122 10.6151
R1339 B.n197 B.n122 10.6151
R1340 B.n198 B.n197 10.6151
R1341 B.n199 B.n198 10.6151
R1342 B.n199 B.n120 10.6151
R1343 B.n203 B.n120 10.6151
R1344 B.n204 B.n203 10.6151
R1345 B.n205 B.n204 10.6151
R1346 B.n205 B.n118 10.6151
R1347 B.n209 B.n118 10.6151
R1348 B.n210 B.n209 10.6151
R1349 B.n211 B.n210 10.6151
R1350 B.n211 B.n116 10.6151
R1351 B.n215 B.n116 10.6151
R1352 B.n216 B.n215 10.6151
R1353 B.n217 B.n216 10.6151
R1354 B.n217 B.n114 10.6151
R1355 B.n221 B.n114 10.6151
R1356 B.n222 B.n221 10.6151
R1357 B.n223 B.n222 10.6151
R1358 B.n223 B.n112 10.6151
R1359 B.n227 B.n112 10.6151
R1360 B.n228 B.n227 10.6151
R1361 B.n230 B.n108 10.6151
R1362 B.n234 B.n108 10.6151
R1363 B.n235 B.n234 10.6151
R1364 B.n236 B.n235 10.6151
R1365 B.n236 B.n106 10.6151
R1366 B.n240 B.n106 10.6151
R1367 B.n241 B.n240 10.6151
R1368 B.n242 B.n241 10.6151
R1369 B.n246 B.n245 10.6151
R1370 B.n247 B.n246 10.6151
R1371 B.n247 B.n100 10.6151
R1372 B.n251 B.n100 10.6151
R1373 B.n252 B.n251 10.6151
R1374 B.n253 B.n252 10.6151
R1375 B.n253 B.n98 10.6151
R1376 B.n257 B.n98 10.6151
R1377 B.n258 B.n257 10.6151
R1378 B.n259 B.n258 10.6151
R1379 B.n259 B.n96 10.6151
R1380 B.n263 B.n96 10.6151
R1381 B.n264 B.n263 10.6151
R1382 B.n265 B.n264 10.6151
R1383 B.n265 B.n94 10.6151
R1384 B.n269 B.n94 10.6151
R1385 B.n270 B.n269 10.6151
R1386 B.n271 B.n270 10.6151
R1387 B.n271 B.n92 10.6151
R1388 B.n275 B.n92 10.6151
R1389 B.n276 B.n275 10.6151
R1390 B.n277 B.n276 10.6151
R1391 B.n277 B.n90 10.6151
R1392 B.n281 B.n90 10.6151
R1393 B.n282 B.n281 10.6151
R1394 B.n283 B.n282 10.6151
R1395 B.n283 B.n88 10.6151
R1396 B.n287 B.n88 10.6151
R1397 B.n288 B.n287 10.6151
R1398 B.n533 B.n0 8.11757
R1399 B.n533 B.n1 8.11757
R1400 B.n440 B.n34 6.5566
R1401 B.n428 B.n427 6.5566
R1402 B.n230 B.n229 6.5566
R1403 B.n242 B.n104 6.5566
R1404 B.n443 B.n34 4.05904
R1405 B.n427 B.n426 4.05904
R1406 B.n229 B.n228 4.05904
R1407 B.n245 B.n104 4.05904
R1408 VN.n4 VN.t6 212.308
R1409 VN.n19 VN.t0 212.308
R1410 VN.n13 VN.t1 193.804
R1411 VN.n28 VN.t7 193.804
R1412 VN.n27 VN.n15 161.3
R1413 VN.n26 VN.n25 161.3
R1414 VN.n24 VN.n23 161.3
R1415 VN.n22 VN.n17 161.3
R1416 VN.n21 VN.n20 161.3
R1417 VN.n12 VN.n0 161.3
R1418 VN.n11 VN.n10 161.3
R1419 VN.n9 VN.n8 161.3
R1420 VN.n7 VN.n2 161.3
R1421 VN.n6 VN.n5 161.3
R1422 VN.n3 VN.t5 160.868
R1423 VN.n1 VN.t2 160.868
R1424 VN.n18 VN.t3 160.868
R1425 VN.n16 VN.t4 160.868
R1426 VN.n29 VN.n28 80.6037
R1427 VN.n14 VN.n13 80.6037
R1428 VN.n4 VN.n3 44.8004
R1429 VN.n19 VN.n18 44.8004
R1430 VN VN.n29 41.7187
R1431 VN.n7 VN.n6 40.4934
R1432 VN.n8 VN.n7 40.4934
R1433 VN.n22 VN.n21 40.4934
R1434 VN.n23 VN.n22 40.4934
R1435 VN.n12 VN.n11 37.5796
R1436 VN.n27 VN.n26 37.5796
R1437 VN.n20 VN.n19 29.7304
R1438 VN.n5 VN.n4 29.7304
R1439 VN.n13 VN.n12 28.4823
R1440 VN.n28 VN.n27 28.4823
R1441 VN.n6 VN.n3 12.968
R1442 VN.n8 VN.n1 12.968
R1443 VN.n21 VN.n18 12.968
R1444 VN.n23 VN.n16 12.968
R1445 VN.n11 VN.n1 11.5
R1446 VN.n26 VN.n16 11.5
R1447 VN.n29 VN.n15 0.285035
R1448 VN.n14 VN.n0 0.285035
R1449 VN.n25 VN.n15 0.189894
R1450 VN.n25 VN.n24 0.189894
R1451 VN.n24 VN.n17 0.189894
R1452 VN.n20 VN.n17 0.189894
R1453 VN.n5 VN.n2 0.189894
R1454 VN.n9 VN.n2 0.189894
R1455 VN.n10 VN.n9 0.189894
R1456 VN.n10 VN.n0 0.189894
R1457 VN VN.n14 0.146778
R1458 VDD2.n2 VDD2.n1 87.0359
R1459 VDD2.n2 VDD2.n0 87.0359
R1460 VDD2 VDD2.n5 87.0331
R1461 VDD2.n4 VDD2.n3 86.432
R1462 VDD2.n4 VDD2.n2 36.5558
R1463 VDD2.n5 VDD2.t4 4.05855
R1464 VDD2.n5 VDD2.t7 4.05855
R1465 VDD2.n3 VDD2.t0 4.05855
R1466 VDD2.n3 VDD2.t3 4.05855
R1467 VDD2.n1 VDD2.t5 4.05855
R1468 VDD2.n1 VDD2.t6 4.05855
R1469 VDD2.n0 VDD2.t1 4.05855
R1470 VDD2.n0 VDD2.t2 4.05855
R1471 VDD2 VDD2.n4 0.718172
C0 B VDD2 1.16749f
C1 VDD1 VDD2 1.07356f
C2 w_n2500_n2570# VTAIL 3.1931f
C3 VN VP 5.21299f
C4 B VDD1 1.11534f
C5 VN VTAIL 4.91129f
C6 w_n2500_n2570# VN 4.63268f
C7 VP VDD2 0.370259f
C8 VP B 1.38168f
C9 VP VDD1 5.03743f
C10 VTAIL VDD2 6.91802f
C11 B VTAIL 3.05038f
C12 VTAIL VDD1 6.87299f
C13 w_n2500_n2570# VDD2 1.4283f
C14 w_n2500_n2570# B 6.85354f
C15 w_n2500_n2570# VDD1 1.37246f
C16 VN VDD2 4.81662f
C17 VN B 0.851998f
C18 VN VDD1 0.14876f
C19 VP VTAIL 4.92539f
C20 w_n2500_n2570# VP 4.9531f
C21 VDD2 VSUBS 1.275083f
C22 VDD1 VSUBS 1.67389f
C23 VTAIL VSUBS 0.873978f
C24 VN VSUBS 4.88727f
C25 VP VSUBS 2.019571f
C26 B VSUBS 3.105534f
C27 w_n2500_n2570# VSUBS 79.71f
C28 VDD2.t1 VSUBS 0.159915f
C29 VDD2.t2 VSUBS 0.159915f
C30 VDD2.n0 VSUBS 1.16638f
C31 VDD2.t5 VSUBS 0.159915f
C32 VDD2.t6 VSUBS 0.159915f
C33 VDD2.n1 VSUBS 1.16638f
C34 VDD2.n2 VSUBS 2.67501f
C35 VDD2.t0 VSUBS 0.159915f
C36 VDD2.t3 VSUBS 0.159915f
C37 VDD2.n3 VSUBS 1.16228f
C38 VDD2.n4 VSUBS 2.39087f
C39 VDD2.t4 VSUBS 0.159915f
C40 VDD2.t7 VSUBS 0.159915f
C41 VDD2.n5 VSUBS 1.16635f
C42 VN.n0 VSUBS 0.062047f
C43 VN.t2 VSUBS 1.20044f
C44 VN.n1 VSUBS 0.460303f
C45 VN.n2 VSUBS 0.046499f
C46 VN.t5 VSUBS 1.20044f
C47 VN.n3 VSUBS 0.519265f
C48 VN.t6 VSUBS 1.33438f
C49 VN.n4 VSUBS 0.537964f
C50 VN.n5 VSUBS 0.238699f
C51 VN.n6 VSUBS 0.072305f
C52 VN.n7 VSUBS 0.03759f
C53 VN.n8 VSUBS 0.072305f
C54 VN.n9 VSUBS 0.046499f
C55 VN.n10 VSUBS 0.046499f
C56 VN.n11 VSUBS 0.070848f
C57 VN.n12 VSUBS 0.027235f
C58 VN.t1 VSUBS 1.28593f
C59 VN.n13 VSUBS 0.545182f
C60 VN.n14 VSUBS 0.043548f
C61 VN.n15 VSUBS 0.062047f
C62 VN.t4 VSUBS 1.20044f
C63 VN.n16 VSUBS 0.460303f
C64 VN.n17 VSUBS 0.046499f
C65 VN.t3 VSUBS 1.20044f
C66 VN.n18 VSUBS 0.519265f
C67 VN.t0 VSUBS 1.33438f
C68 VN.n19 VSUBS 0.537964f
C69 VN.n20 VSUBS 0.238699f
C70 VN.n21 VSUBS 0.072305f
C71 VN.n22 VSUBS 0.03759f
C72 VN.n23 VSUBS 0.072305f
C73 VN.n24 VSUBS 0.046499f
C74 VN.n25 VSUBS 0.046499f
C75 VN.n26 VSUBS 0.070848f
C76 VN.n27 VSUBS 0.027235f
C77 VN.t7 VSUBS 1.28593f
C78 VN.n28 VSUBS 0.545182f
C79 VN.n29 VSUBS 1.91888f
C80 B.n0 VSUBS 0.007386f
C81 B.n1 VSUBS 0.007386f
C82 B.n2 VSUBS 0.010924f
C83 B.n3 VSUBS 0.008371f
C84 B.n4 VSUBS 0.008371f
C85 B.n5 VSUBS 0.008371f
C86 B.n6 VSUBS 0.008371f
C87 B.n7 VSUBS 0.008371f
C88 B.n8 VSUBS 0.008371f
C89 B.n9 VSUBS 0.008371f
C90 B.n10 VSUBS 0.008371f
C91 B.n11 VSUBS 0.008371f
C92 B.n12 VSUBS 0.008371f
C93 B.n13 VSUBS 0.008371f
C94 B.n14 VSUBS 0.008371f
C95 B.n15 VSUBS 0.008371f
C96 B.n16 VSUBS 0.008371f
C97 B.n17 VSUBS 0.021071f
C98 B.n18 VSUBS 0.008371f
C99 B.n19 VSUBS 0.008371f
C100 B.n20 VSUBS 0.008371f
C101 B.n21 VSUBS 0.008371f
C102 B.n22 VSUBS 0.008371f
C103 B.n23 VSUBS 0.008371f
C104 B.n24 VSUBS 0.008371f
C105 B.n25 VSUBS 0.008371f
C106 B.n26 VSUBS 0.008371f
C107 B.n27 VSUBS 0.008371f
C108 B.n28 VSUBS 0.008371f
C109 B.n29 VSUBS 0.008371f
C110 B.n30 VSUBS 0.008371f
C111 B.n31 VSUBS 0.008371f
C112 B.t4 VSUBS 0.151711f
C113 B.t5 VSUBS 0.170431f
C114 B.t3 VSUBS 0.508265f
C115 B.n32 VSUBS 0.282371f
C116 B.n33 VSUBS 0.222369f
C117 B.n34 VSUBS 0.019395f
C118 B.n35 VSUBS 0.008371f
C119 B.n36 VSUBS 0.008371f
C120 B.n37 VSUBS 0.008371f
C121 B.n38 VSUBS 0.008371f
C122 B.n39 VSUBS 0.008371f
C123 B.t1 VSUBS 0.151714f
C124 B.t2 VSUBS 0.170433f
C125 B.t0 VSUBS 0.508265f
C126 B.n40 VSUBS 0.282368f
C127 B.n41 VSUBS 0.222366f
C128 B.n42 VSUBS 0.008371f
C129 B.n43 VSUBS 0.008371f
C130 B.n44 VSUBS 0.008371f
C131 B.n45 VSUBS 0.008371f
C132 B.n46 VSUBS 0.008371f
C133 B.n47 VSUBS 0.008371f
C134 B.n48 VSUBS 0.008371f
C135 B.n49 VSUBS 0.008371f
C136 B.n50 VSUBS 0.008371f
C137 B.n51 VSUBS 0.008371f
C138 B.n52 VSUBS 0.008371f
C139 B.n53 VSUBS 0.008371f
C140 B.n54 VSUBS 0.008371f
C141 B.n55 VSUBS 0.008371f
C142 B.n56 VSUBS 0.020293f
C143 B.n57 VSUBS 0.008371f
C144 B.n58 VSUBS 0.008371f
C145 B.n59 VSUBS 0.008371f
C146 B.n60 VSUBS 0.008371f
C147 B.n61 VSUBS 0.008371f
C148 B.n62 VSUBS 0.008371f
C149 B.n63 VSUBS 0.008371f
C150 B.n64 VSUBS 0.008371f
C151 B.n65 VSUBS 0.008371f
C152 B.n66 VSUBS 0.008371f
C153 B.n67 VSUBS 0.008371f
C154 B.n68 VSUBS 0.008371f
C155 B.n69 VSUBS 0.008371f
C156 B.n70 VSUBS 0.008371f
C157 B.n71 VSUBS 0.008371f
C158 B.n72 VSUBS 0.008371f
C159 B.n73 VSUBS 0.008371f
C160 B.n74 VSUBS 0.008371f
C161 B.n75 VSUBS 0.008371f
C162 B.n76 VSUBS 0.008371f
C163 B.n77 VSUBS 0.008371f
C164 B.n78 VSUBS 0.008371f
C165 B.n79 VSUBS 0.008371f
C166 B.n80 VSUBS 0.008371f
C167 B.n81 VSUBS 0.008371f
C168 B.n82 VSUBS 0.008371f
C169 B.n83 VSUBS 0.008371f
C170 B.n84 VSUBS 0.008371f
C171 B.n85 VSUBS 0.008371f
C172 B.n86 VSUBS 0.008371f
C173 B.n87 VSUBS 0.021071f
C174 B.n88 VSUBS 0.008371f
C175 B.n89 VSUBS 0.008371f
C176 B.n90 VSUBS 0.008371f
C177 B.n91 VSUBS 0.008371f
C178 B.n92 VSUBS 0.008371f
C179 B.n93 VSUBS 0.008371f
C180 B.n94 VSUBS 0.008371f
C181 B.n95 VSUBS 0.008371f
C182 B.n96 VSUBS 0.008371f
C183 B.n97 VSUBS 0.008371f
C184 B.n98 VSUBS 0.008371f
C185 B.n99 VSUBS 0.008371f
C186 B.n100 VSUBS 0.008371f
C187 B.n101 VSUBS 0.008371f
C188 B.t8 VSUBS 0.151714f
C189 B.t7 VSUBS 0.170433f
C190 B.t6 VSUBS 0.508265f
C191 B.n102 VSUBS 0.282368f
C192 B.n103 VSUBS 0.222366f
C193 B.n104 VSUBS 0.019395f
C194 B.n105 VSUBS 0.008371f
C195 B.n106 VSUBS 0.008371f
C196 B.n107 VSUBS 0.008371f
C197 B.n108 VSUBS 0.008371f
C198 B.n109 VSUBS 0.008371f
C199 B.t11 VSUBS 0.151711f
C200 B.t10 VSUBS 0.170431f
C201 B.t9 VSUBS 0.508265f
C202 B.n110 VSUBS 0.282371f
C203 B.n111 VSUBS 0.222369f
C204 B.n112 VSUBS 0.008371f
C205 B.n113 VSUBS 0.008371f
C206 B.n114 VSUBS 0.008371f
C207 B.n115 VSUBS 0.008371f
C208 B.n116 VSUBS 0.008371f
C209 B.n117 VSUBS 0.008371f
C210 B.n118 VSUBS 0.008371f
C211 B.n119 VSUBS 0.008371f
C212 B.n120 VSUBS 0.008371f
C213 B.n121 VSUBS 0.008371f
C214 B.n122 VSUBS 0.008371f
C215 B.n123 VSUBS 0.008371f
C216 B.n124 VSUBS 0.008371f
C217 B.n125 VSUBS 0.008371f
C218 B.n126 VSUBS 0.020293f
C219 B.n127 VSUBS 0.008371f
C220 B.n128 VSUBS 0.008371f
C221 B.n129 VSUBS 0.008371f
C222 B.n130 VSUBS 0.008371f
C223 B.n131 VSUBS 0.008371f
C224 B.n132 VSUBS 0.008371f
C225 B.n133 VSUBS 0.008371f
C226 B.n134 VSUBS 0.008371f
C227 B.n135 VSUBS 0.008371f
C228 B.n136 VSUBS 0.008371f
C229 B.n137 VSUBS 0.008371f
C230 B.n138 VSUBS 0.008371f
C231 B.n139 VSUBS 0.008371f
C232 B.n140 VSUBS 0.008371f
C233 B.n141 VSUBS 0.008371f
C234 B.n142 VSUBS 0.008371f
C235 B.n143 VSUBS 0.008371f
C236 B.n144 VSUBS 0.008371f
C237 B.n145 VSUBS 0.008371f
C238 B.n146 VSUBS 0.008371f
C239 B.n147 VSUBS 0.008371f
C240 B.n148 VSUBS 0.008371f
C241 B.n149 VSUBS 0.008371f
C242 B.n150 VSUBS 0.008371f
C243 B.n151 VSUBS 0.008371f
C244 B.n152 VSUBS 0.008371f
C245 B.n153 VSUBS 0.008371f
C246 B.n154 VSUBS 0.008371f
C247 B.n155 VSUBS 0.008371f
C248 B.n156 VSUBS 0.008371f
C249 B.n157 VSUBS 0.008371f
C250 B.n158 VSUBS 0.008371f
C251 B.n159 VSUBS 0.008371f
C252 B.n160 VSUBS 0.008371f
C253 B.n161 VSUBS 0.008371f
C254 B.n162 VSUBS 0.008371f
C255 B.n163 VSUBS 0.008371f
C256 B.n164 VSUBS 0.008371f
C257 B.n165 VSUBS 0.008371f
C258 B.n166 VSUBS 0.008371f
C259 B.n167 VSUBS 0.008371f
C260 B.n168 VSUBS 0.008371f
C261 B.n169 VSUBS 0.008371f
C262 B.n170 VSUBS 0.008371f
C263 B.n171 VSUBS 0.008371f
C264 B.n172 VSUBS 0.008371f
C265 B.n173 VSUBS 0.008371f
C266 B.n174 VSUBS 0.008371f
C267 B.n175 VSUBS 0.008371f
C268 B.n176 VSUBS 0.008371f
C269 B.n177 VSUBS 0.008371f
C270 B.n178 VSUBS 0.008371f
C271 B.n179 VSUBS 0.008371f
C272 B.n180 VSUBS 0.008371f
C273 B.n181 VSUBS 0.008371f
C274 B.n182 VSUBS 0.008371f
C275 B.n183 VSUBS 0.020293f
C276 B.n184 VSUBS 0.021071f
C277 B.n185 VSUBS 0.021071f
C278 B.n186 VSUBS 0.008371f
C279 B.n187 VSUBS 0.008371f
C280 B.n188 VSUBS 0.008371f
C281 B.n189 VSUBS 0.008371f
C282 B.n190 VSUBS 0.008371f
C283 B.n191 VSUBS 0.008371f
C284 B.n192 VSUBS 0.008371f
C285 B.n193 VSUBS 0.008371f
C286 B.n194 VSUBS 0.008371f
C287 B.n195 VSUBS 0.008371f
C288 B.n196 VSUBS 0.008371f
C289 B.n197 VSUBS 0.008371f
C290 B.n198 VSUBS 0.008371f
C291 B.n199 VSUBS 0.008371f
C292 B.n200 VSUBS 0.008371f
C293 B.n201 VSUBS 0.008371f
C294 B.n202 VSUBS 0.008371f
C295 B.n203 VSUBS 0.008371f
C296 B.n204 VSUBS 0.008371f
C297 B.n205 VSUBS 0.008371f
C298 B.n206 VSUBS 0.008371f
C299 B.n207 VSUBS 0.008371f
C300 B.n208 VSUBS 0.008371f
C301 B.n209 VSUBS 0.008371f
C302 B.n210 VSUBS 0.008371f
C303 B.n211 VSUBS 0.008371f
C304 B.n212 VSUBS 0.008371f
C305 B.n213 VSUBS 0.008371f
C306 B.n214 VSUBS 0.008371f
C307 B.n215 VSUBS 0.008371f
C308 B.n216 VSUBS 0.008371f
C309 B.n217 VSUBS 0.008371f
C310 B.n218 VSUBS 0.008371f
C311 B.n219 VSUBS 0.008371f
C312 B.n220 VSUBS 0.008371f
C313 B.n221 VSUBS 0.008371f
C314 B.n222 VSUBS 0.008371f
C315 B.n223 VSUBS 0.008371f
C316 B.n224 VSUBS 0.008371f
C317 B.n225 VSUBS 0.008371f
C318 B.n226 VSUBS 0.008371f
C319 B.n227 VSUBS 0.008371f
C320 B.n228 VSUBS 0.005786f
C321 B.n229 VSUBS 0.019395f
C322 B.n230 VSUBS 0.006771f
C323 B.n231 VSUBS 0.008371f
C324 B.n232 VSUBS 0.008371f
C325 B.n233 VSUBS 0.008371f
C326 B.n234 VSUBS 0.008371f
C327 B.n235 VSUBS 0.008371f
C328 B.n236 VSUBS 0.008371f
C329 B.n237 VSUBS 0.008371f
C330 B.n238 VSUBS 0.008371f
C331 B.n239 VSUBS 0.008371f
C332 B.n240 VSUBS 0.008371f
C333 B.n241 VSUBS 0.008371f
C334 B.n242 VSUBS 0.006771f
C335 B.n243 VSUBS 0.008371f
C336 B.n244 VSUBS 0.008371f
C337 B.n245 VSUBS 0.005786f
C338 B.n246 VSUBS 0.008371f
C339 B.n247 VSUBS 0.008371f
C340 B.n248 VSUBS 0.008371f
C341 B.n249 VSUBS 0.008371f
C342 B.n250 VSUBS 0.008371f
C343 B.n251 VSUBS 0.008371f
C344 B.n252 VSUBS 0.008371f
C345 B.n253 VSUBS 0.008371f
C346 B.n254 VSUBS 0.008371f
C347 B.n255 VSUBS 0.008371f
C348 B.n256 VSUBS 0.008371f
C349 B.n257 VSUBS 0.008371f
C350 B.n258 VSUBS 0.008371f
C351 B.n259 VSUBS 0.008371f
C352 B.n260 VSUBS 0.008371f
C353 B.n261 VSUBS 0.008371f
C354 B.n262 VSUBS 0.008371f
C355 B.n263 VSUBS 0.008371f
C356 B.n264 VSUBS 0.008371f
C357 B.n265 VSUBS 0.008371f
C358 B.n266 VSUBS 0.008371f
C359 B.n267 VSUBS 0.008371f
C360 B.n268 VSUBS 0.008371f
C361 B.n269 VSUBS 0.008371f
C362 B.n270 VSUBS 0.008371f
C363 B.n271 VSUBS 0.008371f
C364 B.n272 VSUBS 0.008371f
C365 B.n273 VSUBS 0.008371f
C366 B.n274 VSUBS 0.008371f
C367 B.n275 VSUBS 0.008371f
C368 B.n276 VSUBS 0.008371f
C369 B.n277 VSUBS 0.008371f
C370 B.n278 VSUBS 0.008371f
C371 B.n279 VSUBS 0.008371f
C372 B.n280 VSUBS 0.008371f
C373 B.n281 VSUBS 0.008371f
C374 B.n282 VSUBS 0.008371f
C375 B.n283 VSUBS 0.008371f
C376 B.n284 VSUBS 0.008371f
C377 B.n285 VSUBS 0.008371f
C378 B.n286 VSUBS 0.008371f
C379 B.n287 VSUBS 0.008371f
C380 B.n288 VSUBS 0.02016f
C381 B.n289 VSUBS 0.021205f
C382 B.n290 VSUBS 0.020293f
C383 B.n291 VSUBS 0.008371f
C384 B.n292 VSUBS 0.008371f
C385 B.n293 VSUBS 0.008371f
C386 B.n294 VSUBS 0.008371f
C387 B.n295 VSUBS 0.008371f
C388 B.n296 VSUBS 0.008371f
C389 B.n297 VSUBS 0.008371f
C390 B.n298 VSUBS 0.008371f
C391 B.n299 VSUBS 0.008371f
C392 B.n300 VSUBS 0.008371f
C393 B.n301 VSUBS 0.008371f
C394 B.n302 VSUBS 0.008371f
C395 B.n303 VSUBS 0.008371f
C396 B.n304 VSUBS 0.008371f
C397 B.n305 VSUBS 0.008371f
C398 B.n306 VSUBS 0.008371f
C399 B.n307 VSUBS 0.008371f
C400 B.n308 VSUBS 0.008371f
C401 B.n309 VSUBS 0.008371f
C402 B.n310 VSUBS 0.008371f
C403 B.n311 VSUBS 0.008371f
C404 B.n312 VSUBS 0.008371f
C405 B.n313 VSUBS 0.008371f
C406 B.n314 VSUBS 0.008371f
C407 B.n315 VSUBS 0.008371f
C408 B.n316 VSUBS 0.008371f
C409 B.n317 VSUBS 0.008371f
C410 B.n318 VSUBS 0.008371f
C411 B.n319 VSUBS 0.008371f
C412 B.n320 VSUBS 0.008371f
C413 B.n321 VSUBS 0.008371f
C414 B.n322 VSUBS 0.008371f
C415 B.n323 VSUBS 0.008371f
C416 B.n324 VSUBS 0.008371f
C417 B.n325 VSUBS 0.008371f
C418 B.n326 VSUBS 0.008371f
C419 B.n327 VSUBS 0.008371f
C420 B.n328 VSUBS 0.008371f
C421 B.n329 VSUBS 0.008371f
C422 B.n330 VSUBS 0.008371f
C423 B.n331 VSUBS 0.008371f
C424 B.n332 VSUBS 0.008371f
C425 B.n333 VSUBS 0.008371f
C426 B.n334 VSUBS 0.008371f
C427 B.n335 VSUBS 0.008371f
C428 B.n336 VSUBS 0.008371f
C429 B.n337 VSUBS 0.008371f
C430 B.n338 VSUBS 0.008371f
C431 B.n339 VSUBS 0.008371f
C432 B.n340 VSUBS 0.008371f
C433 B.n341 VSUBS 0.008371f
C434 B.n342 VSUBS 0.008371f
C435 B.n343 VSUBS 0.008371f
C436 B.n344 VSUBS 0.008371f
C437 B.n345 VSUBS 0.008371f
C438 B.n346 VSUBS 0.008371f
C439 B.n347 VSUBS 0.008371f
C440 B.n348 VSUBS 0.008371f
C441 B.n349 VSUBS 0.008371f
C442 B.n350 VSUBS 0.008371f
C443 B.n351 VSUBS 0.008371f
C444 B.n352 VSUBS 0.008371f
C445 B.n353 VSUBS 0.008371f
C446 B.n354 VSUBS 0.008371f
C447 B.n355 VSUBS 0.008371f
C448 B.n356 VSUBS 0.008371f
C449 B.n357 VSUBS 0.008371f
C450 B.n358 VSUBS 0.008371f
C451 B.n359 VSUBS 0.008371f
C452 B.n360 VSUBS 0.008371f
C453 B.n361 VSUBS 0.008371f
C454 B.n362 VSUBS 0.008371f
C455 B.n363 VSUBS 0.008371f
C456 B.n364 VSUBS 0.008371f
C457 B.n365 VSUBS 0.008371f
C458 B.n366 VSUBS 0.008371f
C459 B.n367 VSUBS 0.008371f
C460 B.n368 VSUBS 0.008371f
C461 B.n369 VSUBS 0.008371f
C462 B.n370 VSUBS 0.008371f
C463 B.n371 VSUBS 0.008371f
C464 B.n372 VSUBS 0.008371f
C465 B.n373 VSUBS 0.008371f
C466 B.n374 VSUBS 0.008371f
C467 B.n375 VSUBS 0.008371f
C468 B.n376 VSUBS 0.008371f
C469 B.n377 VSUBS 0.008371f
C470 B.n378 VSUBS 0.008371f
C471 B.n379 VSUBS 0.008371f
C472 B.n380 VSUBS 0.008371f
C473 B.n381 VSUBS 0.020293f
C474 B.n382 VSUBS 0.021071f
C475 B.n383 VSUBS 0.021071f
C476 B.n384 VSUBS 0.008371f
C477 B.n385 VSUBS 0.008371f
C478 B.n386 VSUBS 0.008371f
C479 B.n387 VSUBS 0.008371f
C480 B.n388 VSUBS 0.008371f
C481 B.n389 VSUBS 0.008371f
C482 B.n390 VSUBS 0.008371f
C483 B.n391 VSUBS 0.008371f
C484 B.n392 VSUBS 0.008371f
C485 B.n393 VSUBS 0.008371f
C486 B.n394 VSUBS 0.008371f
C487 B.n395 VSUBS 0.008371f
C488 B.n396 VSUBS 0.008371f
C489 B.n397 VSUBS 0.008371f
C490 B.n398 VSUBS 0.008371f
C491 B.n399 VSUBS 0.008371f
C492 B.n400 VSUBS 0.008371f
C493 B.n401 VSUBS 0.008371f
C494 B.n402 VSUBS 0.008371f
C495 B.n403 VSUBS 0.008371f
C496 B.n404 VSUBS 0.008371f
C497 B.n405 VSUBS 0.008371f
C498 B.n406 VSUBS 0.008371f
C499 B.n407 VSUBS 0.008371f
C500 B.n408 VSUBS 0.008371f
C501 B.n409 VSUBS 0.008371f
C502 B.n410 VSUBS 0.008371f
C503 B.n411 VSUBS 0.008371f
C504 B.n412 VSUBS 0.008371f
C505 B.n413 VSUBS 0.008371f
C506 B.n414 VSUBS 0.008371f
C507 B.n415 VSUBS 0.008371f
C508 B.n416 VSUBS 0.008371f
C509 B.n417 VSUBS 0.008371f
C510 B.n418 VSUBS 0.008371f
C511 B.n419 VSUBS 0.008371f
C512 B.n420 VSUBS 0.008371f
C513 B.n421 VSUBS 0.008371f
C514 B.n422 VSUBS 0.008371f
C515 B.n423 VSUBS 0.008371f
C516 B.n424 VSUBS 0.008371f
C517 B.n425 VSUBS 0.008371f
C518 B.n426 VSUBS 0.005786f
C519 B.n427 VSUBS 0.019395f
C520 B.n428 VSUBS 0.006771f
C521 B.n429 VSUBS 0.008371f
C522 B.n430 VSUBS 0.008371f
C523 B.n431 VSUBS 0.008371f
C524 B.n432 VSUBS 0.008371f
C525 B.n433 VSUBS 0.008371f
C526 B.n434 VSUBS 0.008371f
C527 B.n435 VSUBS 0.008371f
C528 B.n436 VSUBS 0.008371f
C529 B.n437 VSUBS 0.008371f
C530 B.n438 VSUBS 0.008371f
C531 B.n439 VSUBS 0.008371f
C532 B.n440 VSUBS 0.006771f
C533 B.n441 VSUBS 0.008371f
C534 B.n442 VSUBS 0.008371f
C535 B.n443 VSUBS 0.005786f
C536 B.n444 VSUBS 0.008371f
C537 B.n445 VSUBS 0.008371f
C538 B.n446 VSUBS 0.008371f
C539 B.n447 VSUBS 0.008371f
C540 B.n448 VSUBS 0.008371f
C541 B.n449 VSUBS 0.008371f
C542 B.n450 VSUBS 0.008371f
C543 B.n451 VSUBS 0.008371f
C544 B.n452 VSUBS 0.008371f
C545 B.n453 VSUBS 0.008371f
C546 B.n454 VSUBS 0.008371f
C547 B.n455 VSUBS 0.008371f
C548 B.n456 VSUBS 0.008371f
C549 B.n457 VSUBS 0.008371f
C550 B.n458 VSUBS 0.008371f
C551 B.n459 VSUBS 0.008371f
C552 B.n460 VSUBS 0.008371f
C553 B.n461 VSUBS 0.008371f
C554 B.n462 VSUBS 0.008371f
C555 B.n463 VSUBS 0.008371f
C556 B.n464 VSUBS 0.008371f
C557 B.n465 VSUBS 0.008371f
C558 B.n466 VSUBS 0.008371f
C559 B.n467 VSUBS 0.008371f
C560 B.n468 VSUBS 0.008371f
C561 B.n469 VSUBS 0.008371f
C562 B.n470 VSUBS 0.008371f
C563 B.n471 VSUBS 0.008371f
C564 B.n472 VSUBS 0.008371f
C565 B.n473 VSUBS 0.008371f
C566 B.n474 VSUBS 0.008371f
C567 B.n475 VSUBS 0.008371f
C568 B.n476 VSUBS 0.008371f
C569 B.n477 VSUBS 0.008371f
C570 B.n478 VSUBS 0.008371f
C571 B.n479 VSUBS 0.008371f
C572 B.n480 VSUBS 0.008371f
C573 B.n481 VSUBS 0.008371f
C574 B.n482 VSUBS 0.008371f
C575 B.n483 VSUBS 0.008371f
C576 B.n484 VSUBS 0.008371f
C577 B.n485 VSUBS 0.008371f
C578 B.n486 VSUBS 0.021071f
C579 B.n487 VSUBS 0.020293f
C580 B.n488 VSUBS 0.020293f
C581 B.n489 VSUBS 0.008371f
C582 B.n490 VSUBS 0.008371f
C583 B.n491 VSUBS 0.008371f
C584 B.n492 VSUBS 0.008371f
C585 B.n493 VSUBS 0.008371f
C586 B.n494 VSUBS 0.008371f
C587 B.n495 VSUBS 0.008371f
C588 B.n496 VSUBS 0.008371f
C589 B.n497 VSUBS 0.008371f
C590 B.n498 VSUBS 0.008371f
C591 B.n499 VSUBS 0.008371f
C592 B.n500 VSUBS 0.008371f
C593 B.n501 VSUBS 0.008371f
C594 B.n502 VSUBS 0.008371f
C595 B.n503 VSUBS 0.008371f
C596 B.n504 VSUBS 0.008371f
C597 B.n505 VSUBS 0.008371f
C598 B.n506 VSUBS 0.008371f
C599 B.n507 VSUBS 0.008371f
C600 B.n508 VSUBS 0.008371f
C601 B.n509 VSUBS 0.008371f
C602 B.n510 VSUBS 0.008371f
C603 B.n511 VSUBS 0.008371f
C604 B.n512 VSUBS 0.008371f
C605 B.n513 VSUBS 0.008371f
C606 B.n514 VSUBS 0.008371f
C607 B.n515 VSUBS 0.008371f
C608 B.n516 VSUBS 0.008371f
C609 B.n517 VSUBS 0.008371f
C610 B.n518 VSUBS 0.008371f
C611 B.n519 VSUBS 0.008371f
C612 B.n520 VSUBS 0.008371f
C613 B.n521 VSUBS 0.008371f
C614 B.n522 VSUBS 0.008371f
C615 B.n523 VSUBS 0.008371f
C616 B.n524 VSUBS 0.008371f
C617 B.n525 VSUBS 0.008371f
C618 B.n526 VSUBS 0.008371f
C619 B.n527 VSUBS 0.008371f
C620 B.n528 VSUBS 0.008371f
C621 B.n529 VSUBS 0.008371f
C622 B.n530 VSUBS 0.008371f
C623 B.n531 VSUBS 0.010924f
C624 B.n532 VSUBS 0.011637f
C625 B.n533 VSUBS 0.023141f
C626 VTAIL.t0 VSUBS 0.163141f
C627 VTAIL.t6 VSUBS 0.163141f
C628 VTAIL.n0 VSUBS 1.08356f
C629 VTAIL.n1 VSUBS 0.613674f
C630 VTAIL.n2 VSUBS 0.027884f
C631 VTAIL.n3 VSUBS 0.025774f
C632 VTAIL.n4 VSUBS 0.014257f
C633 VTAIL.n5 VSUBS 0.032736f
C634 VTAIL.n6 VSUBS 0.014664f
C635 VTAIL.n7 VSUBS 0.025774f
C636 VTAIL.n8 VSUBS 0.01385f
C637 VTAIL.n9 VSUBS 0.032736f
C638 VTAIL.n10 VSUBS 0.014664f
C639 VTAIL.n11 VSUBS 0.025774f
C640 VTAIL.n12 VSUBS 0.01385f
C641 VTAIL.n13 VSUBS 0.024552f
C642 VTAIL.n14 VSUBS 0.024625f
C643 VTAIL.t3 VSUBS 0.070333f
C644 VTAIL.n15 VSUBS 0.156601f
C645 VTAIL.n16 VSUBS 0.815494f
C646 VTAIL.n17 VSUBS 0.01385f
C647 VTAIL.n18 VSUBS 0.014664f
C648 VTAIL.n19 VSUBS 0.032736f
C649 VTAIL.n20 VSUBS 0.032736f
C650 VTAIL.n21 VSUBS 0.014664f
C651 VTAIL.n22 VSUBS 0.01385f
C652 VTAIL.n23 VSUBS 0.025774f
C653 VTAIL.n24 VSUBS 0.025774f
C654 VTAIL.n25 VSUBS 0.01385f
C655 VTAIL.n26 VSUBS 0.014664f
C656 VTAIL.n27 VSUBS 0.032736f
C657 VTAIL.n28 VSUBS 0.032736f
C658 VTAIL.n29 VSUBS 0.014664f
C659 VTAIL.n30 VSUBS 0.01385f
C660 VTAIL.n31 VSUBS 0.025774f
C661 VTAIL.n32 VSUBS 0.025774f
C662 VTAIL.n33 VSUBS 0.01385f
C663 VTAIL.n34 VSUBS 0.01385f
C664 VTAIL.n35 VSUBS 0.014664f
C665 VTAIL.n36 VSUBS 0.032736f
C666 VTAIL.n37 VSUBS 0.032736f
C667 VTAIL.n38 VSUBS 0.077766f
C668 VTAIL.n39 VSUBS 0.014257f
C669 VTAIL.n40 VSUBS 0.01385f
C670 VTAIL.n41 VSUBS 0.066969f
C671 VTAIL.n42 VSUBS 0.039257f
C672 VTAIL.n43 VSUBS 0.174754f
C673 VTAIL.n44 VSUBS 0.027884f
C674 VTAIL.n45 VSUBS 0.025774f
C675 VTAIL.n46 VSUBS 0.014257f
C676 VTAIL.n47 VSUBS 0.032736f
C677 VTAIL.n48 VSUBS 0.014664f
C678 VTAIL.n49 VSUBS 0.025774f
C679 VTAIL.n50 VSUBS 0.01385f
C680 VTAIL.n51 VSUBS 0.032736f
C681 VTAIL.n52 VSUBS 0.014664f
C682 VTAIL.n53 VSUBS 0.025774f
C683 VTAIL.n54 VSUBS 0.01385f
C684 VTAIL.n55 VSUBS 0.024552f
C685 VTAIL.n56 VSUBS 0.024625f
C686 VTAIL.t10 VSUBS 0.070333f
C687 VTAIL.n57 VSUBS 0.156601f
C688 VTAIL.n58 VSUBS 0.815494f
C689 VTAIL.n59 VSUBS 0.01385f
C690 VTAIL.n60 VSUBS 0.014664f
C691 VTAIL.n61 VSUBS 0.032736f
C692 VTAIL.n62 VSUBS 0.032736f
C693 VTAIL.n63 VSUBS 0.014664f
C694 VTAIL.n64 VSUBS 0.01385f
C695 VTAIL.n65 VSUBS 0.025774f
C696 VTAIL.n66 VSUBS 0.025774f
C697 VTAIL.n67 VSUBS 0.01385f
C698 VTAIL.n68 VSUBS 0.014664f
C699 VTAIL.n69 VSUBS 0.032736f
C700 VTAIL.n70 VSUBS 0.032736f
C701 VTAIL.n71 VSUBS 0.014664f
C702 VTAIL.n72 VSUBS 0.01385f
C703 VTAIL.n73 VSUBS 0.025774f
C704 VTAIL.n74 VSUBS 0.025774f
C705 VTAIL.n75 VSUBS 0.01385f
C706 VTAIL.n76 VSUBS 0.01385f
C707 VTAIL.n77 VSUBS 0.014664f
C708 VTAIL.n78 VSUBS 0.032736f
C709 VTAIL.n79 VSUBS 0.032736f
C710 VTAIL.n80 VSUBS 0.077766f
C711 VTAIL.n81 VSUBS 0.014257f
C712 VTAIL.n82 VSUBS 0.01385f
C713 VTAIL.n83 VSUBS 0.066969f
C714 VTAIL.n84 VSUBS 0.039257f
C715 VTAIL.n85 VSUBS 0.174754f
C716 VTAIL.t13 VSUBS 0.163141f
C717 VTAIL.t11 VSUBS 0.163141f
C718 VTAIL.n86 VSUBS 1.08356f
C719 VTAIL.n87 VSUBS 0.718379f
C720 VTAIL.n88 VSUBS 0.027884f
C721 VTAIL.n89 VSUBS 0.025774f
C722 VTAIL.n90 VSUBS 0.014257f
C723 VTAIL.n91 VSUBS 0.032736f
C724 VTAIL.n92 VSUBS 0.014664f
C725 VTAIL.n93 VSUBS 0.025774f
C726 VTAIL.n94 VSUBS 0.01385f
C727 VTAIL.n95 VSUBS 0.032736f
C728 VTAIL.n96 VSUBS 0.014664f
C729 VTAIL.n97 VSUBS 0.025774f
C730 VTAIL.n98 VSUBS 0.01385f
C731 VTAIL.n99 VSUBS 0.024552f
C732 VTAIL.n100 VSUBS 0.024625f
C733 VTAIL.t8 VSUBS 0.070333f
C734 VTAIL.n101 VSUBS 0.156601f
C735 VTAIL.n102 VSUBS 0.815494f
C736 VTAIL.n103 VSUBS 0.01385f
C737 VTAIL.n104 VSUBS 0.014664f
C738 VTAIL.n105 VSUBS 0.032736f
C739 VTAIL.n106 VSUBS 0.032736f
C740 VTAIL.n107 VSUBS 0.014664f
C741 VTAIL.n108 VSUBS 0.01385f
C742 VTAIL.n109 VSUBS 0.025774f
C743 VTAIL.n110 VSUBS 0.025774f
C744 VTAIL.n111 VSUBS 0.01385f
C745 VTAIL.n112 VSUBS 0.014664f
C746 VTAIL.n113 VSUBS 0.032736f
C747 VTAIL.n114 VSUBS 0.032736f
C748 VTAIL.n115 VSUBS 0.014664f
C749 VTAIL.n116 VSUBS 0.01385f
C750 VTAIL.n117 VSUBS 0.025774f
C751 VTAIL.n118 VSUBS 0.025774f
C752 VTAIL.n119 VSUBS 0.01385f
C753 VTAIL.n120 VSUBS 0.01385f
C754 VTAIL.n121 VSUBS 0.014664f
C755 VTAIL.n122 VSUBS 0.032736f
C756 VTAIL.n123 VSUBS 0.032736f
C757 VTAIL.n124 VSUBS 0.077766f
C758 VTAIL.n125 VSUBS 0.014257f
C759 VTAIL.n126 VSUBS 0.01385f
C760 VTAIL.n127 VSUBS 0.066969f
C761 VTAIL.n128 VSUBS 0.039257f
C762 VTAIL.n129 VSUBS 1.16884f
C763 VTAIL.n130 VSUBS 0.027884f
C764 VTAIL.n131 VSUBS 0.025774f
C765 VTAIL.n132 VSUBS 0.014257f
C766 VTAIL.n133 VSUBS 0.032736f
C767 VTAIL.n134 VSUBS 0.01385f
C768 VTAIL.n135 VSUBS 0.014664f
C769 VTAIL.n136 VSUBS 0.025774f
C770 VTAIL.n137 VSUBS 0.01385f
C771 VTAIL.n138 VSUBS 0.032736f
C772 VTAIL.n139 VSUBS 0.014664f
C773 VTAIL.n140 VSUBS 0.025774f
C774 VTAIL.n141 VSUBS 0.01385f
C775 VTAIL.n142 VSUBS 0.024552f
C776 VTAIL.n143 VSUBS 0.024625f
C777 VTAIL.t5 VSUBS 0.070333f
C778 VTAIL.n144 VSUBS 0.156601f
C779 VTAIL.n145 VSUBS 0.815494f
C780 VTAIL.n146 VSUBS 0.01385f
C781 VTAIL.n147 VSUBS 0.014664f
C782 VTAIL.n148 VSUBS 0.032736f
C783 VTAIL.n149 VSUBS 0.032736f
C784 VTAIL.n150 VSUBS 0.014664f
C785 VTAIL.n151 VSUBS 0.01385f
C786 VTAIL.n152 VSUBS 0.025774f
C787 VTAIL.n153 VSUBS 0.025774f
C788 VTAIL.n154 VSUBS 0.01385f
C789 VTAIL.n155 VSUBS 0.014664f
C790 VTAIL.n156 VSUBS 0.032736f
C791 VTAIL.n157 VSUBS 0.032736f
C792 VTAIL.n158 VSUBS 0.014664f
C793 VTAIL.n159 VSUBS 0.01385f
C794 VTAIL.n160 VSUBS 0.025774f
C795 VTAIL.n161 VSUBS 0.025774f
C796 VTAIL.n162 VSUBS 0.01385f
C797 VTAIL.n163 VSUBS 0.014664f
C798 VTAIL.n164 VSUBS 0.032736f
C799 VTAIL.n165 VSUBS 0.032736f
C800 VTAIL.n166 VSUBS 0.077766f
C801 VTAIL.n167 VSUBS 0.014257f
C802 VTAIL.n168 VSUBS 0.01385f
C803 VTAIL.n169 VSUBS 0.066969f
C804 VTAIL.n170 VSUBS 0.039257f
C805 VTAIL.n171 VSUBS 1.16884f
C806 VTAIL.t4 VSUBS 0.163141f
C807 VTAIL.t7 VSUBS 0.163141f
C808 VTAIL.n172 VSUBS 1.08356f
C809 VTAIL.n173 VSUBS 0.718372f
C810 VTAIL.n174 VSUBS 0.027884f
C811 VTAIL.n175 VSUBS 0.025774f
C812 VTAIL.n176 VSUBS 0.014257f
C813 VTAIL.n177 VSUBS 0.032736f
C814 VTAIL.n178 VSUBS 0.01385f
C815 VTAIL.n179 VSUBS 0.014664f
C816 VTAIL.n180 VSUBS 0.025774f
C817 VTAIL.n181 VSUBS 0.01385f
C818 VTAIL.n182 VSUBS 0.032736f
C819 VTAIL.n183 VSUBS 0.014664f
C820 VTAIL.n184 VSUBS 0.025774f
C821 VTAIL.n185 VSUBS 0.01385f
C822 VTAIL.n186 VSUBS 0.024552f
C823 VTAIL.n187 VSUBS 0.024625f
C824 VTAIL.t2 VSUBS 0.070333f
C825 VTAIL.n188 VSUBS 0.156601f
C826 VTAIL.n189 VSUBS 0.815494f
C827 VTAIL.n190 VSUBS 0.01385f
C828 VTAIL.n191 VSUBS 0.014664f
C829 VTAIL.n192 VSUBS 0.032736f
C830 VTAIL.n193 VSUBS 0.032736f
C831 VTAIL.n194 VSUBS 0.014664f
C832 VTAIL.n195 VSUBS 0.01385f
C833 VTAIL.n196 VSUBS 0.025774f
C834 VTAIL.n197 VSUBS 0.025774f
C835 VTAIL.n198 VSUBS 0.01385f
C836 VTAIL.n199 VSUBS 0.014664f
C837 VTAIL.n200 VSUBS 0.032736f
C838 VTAIL.n201 VSUBS 0.032736f
C839 VTAIL.n202 VSUBS 0.014664f
C840 VTAIL.n203 VSUBS 0.01385f
C841 VTAIL.n204 VSUBS 0.025774f
C842 VTAIL.n205 VSUBS 0.025774f
C843 VTAIL.n206 VSUBS 0.01385f
C844 VTAIL.n207 VSUBS 0.014664f
C845 VTAIL.n208 VSUBS 0.032736f
C846 VTAIL.n209 VSUBS 0.032736f
C847 VTAIL.n210 VSUBS 0.077766f
C848 VTAIL.n211 VSUBS 0.014257f
C849 VTAIL.n212 VSUBS 0.01385f
C850 VTAIL.n213 VSUBS 0.066969f
C851 VTAIL.n214 VSUBS 0.039257f
C852 VTAIL.n215 VSUBS 0.174754f
C853 VTAIL.n216 VSUBS 0.027884f
C854 VTAIL.n217 VSUBS 0.025774f
C855 VTAIL.n218 VSUBS 0.014257f
C856 VTAIL.n219 VSUBS 0.032736f
C857 VTAIL.n220 VSUBS 0.01385f
C858 VTAIL.n221 VSUBS 0.014664f
C859 VTAIL.n222 VSUBS 0.025774f
C860 VTAIL.n223 VSUBS 0.01385f
C861 VTAIL.n224 VSUBS 0.032736f
C862 VTAIL.n225 VSUBS 0.014664f
C863 VTAIL.n226 VSUBS 0.025774f
C864 VTAIL.n227 VSUBS 0.01385f
C865 VTAIL.n228 VSUBS 0.024552f
C866 VTAIL.n229 VSUBS 0.024625f
C867 VTAIL.t12 VSUBS 0.070333f
C868 VTAIL.n230 VSUBS 0.156601f
C869 VTAIL.n231 VSUBS 0.815494f
C870 VTAIL.n232 VSUBS 0.01385f
C871 VTAIL.n233 VSUBS 0.014664f
C872 VTAIL.n234 VSUBS 0.032736f
C873 VTAIL.n235 VSUBS 0.032736f
C874 VTAIL.n236 VSUBS 0.014664f
C875 VTAIL.n237 VSUBS 0.01385f
C876 VTAIL.n238 VSUBS 0.025774f
C877 VTAIL.n239 VSUBS 0.025774f
C878 VTAIL.n240 VSUBS 0.01385f
C879 VTAIL.n241 VSUBS 0.014664f
C880 VTAIL.n242 VSUBS 0.032736f
C881 VTAIL.n243 VSUBS 0.032736f
C882 VTAIL.n244 VSUBS 0.014664f
C883 VTAIL.n245 VSUBS 0.01385f
C884 VTAIL.n246 VSUBS 0.025774f
C885 VTAIL.n247 VSUBS 0.025774f
C886 VTAIL.n248 VSUBS 0.01385f
C887 VTAIL.n249 VSUBS 0.014664f
C888 VTAIL.n250 VSUBS 0.032736f
C889 VTAIL.n251 VSUBS 0.032736f
C890 VTAIL.n252 VSUBS 0.077766f
C891 VTAIL.n253 VSUBS 0.014257f
C892 VTAIL.n254 VSUBS 0.01385f
C893 VTAIL.n255 VSUBS 0.066969f
C894 VTAIL.n256 VSUBS 0.039257f
C895 VTAIL.n257 VSUBS 0.174754f
C896 VTAIL.t9 VSUBS 0.163141f
C897 VTAIL.t15 VSUBS 0.163141f
C898 VTAIL.n258 VSUBS 1.08356f
C899 VTAIL.n259 VSUBS 0.718372f
C900 VTAIL.n260 VSUBS 0.027884f
C901 VTAIL.n261 VSUBS 0.025774f
C902 VTAIL.n262 VSUBS 0.014257f
C903 VTAIL.n263 VSUBS 0.032736f
C904 VTAIL.n264 VSUBS 0.01385f
C905 VTAIL.n265 VSUBS 0.014664f
C906 VTAIL.n266 VSUBS 0.025774f
C907 VTAIL.n267 VSUBS 0.01385f
C908 VTAIL.n268 VSUBS 0.032736f
C909 VTAIL.n269 VSUBS 0.014664f
C910 VTAIL.n270 VSUBS 0.025774f
C911 VTAIL.n271 VSUBS 0.01385f
C912 VTAIL.n272 VSUBS 0.024552f
C913 VTAIL.n273 VSUBS 0.024625f
C914 VTAIL.t14 VSUBS 0.070333f
C915 VTAIL.n274 VSUBS 0.156601f
C916 VTAIL.n275 VSUBS 0.815494f
C917 VTAIL.n276 VSUBS 0.01385f
C918 VTAIL.n277 VSUBS 0.014664f
C919 VTAIL.n278 VSUBS 0.032736f
C920 VTAIL.n279 VSUBS 0.032736f
C921 VTAIL.n280 VSUBS 0.014664f
C922 VTAIL.n281 VSUBS 0.01385f
C923 VTAIL.n282 VSUBS 0.025774f
C924 VTAIL.n283 VSUBS 0.025774f
C925 VTAIL.n284 VSUBS 0.01385f
C926 VTAIL.n285 VSUBS 0.014664f
C927 VTAIL.n286 VSUBS 0.032736f
C928 VTAIL.n287 VSUBS 0.032736f
C929 VTAIL.n288 VSUBS 0.014664f
C930 VTAIL.n289 VSUBS 0.01385f
C931 VTAIL.n290 VSUBS 0.025774f
C932 VTAIL.n291 VSUBS 0.025774f
C933 VTAIL.n292 VSUBS 0.01385f
C934 VTAIL.n293 VSUBS 0.014664f
C935 VTAIL.n294 VSUBS 0.032736f
C936 VTAIL.n295 VSUBS 0.032736f
C937 VTAIL.n296 VSUBS 0.077766f
C938 VTAIL.n297 VSUBS 0.014257f
C939 VTAIL.n298 VSUBS 0.01385f
C940 VTAIL.n299 VSUBS 0.066969f
C941 VTAIL.n300 VSUBS 0.039257f
C942 VTAIL.n301 VSUBS 1.16884f
C943 VTAIL.n302 VSUBS 0.027884f
C944 VTAIL.n303 VSUBS 0.025774f
C945 VTAIL.n304 VSUBS 0.014257f
C946 VTAIL.n305 VSUBS 0.032736f
C947 VTAIL.n306 VSUBS 0.014664f
C948 VTAIL.n307 VSUBS 0.025774f
C949 VTAIL.n308 VSUBS 0.01385f
C950 VTAIL.n309 VSUBS 0.032736f
C951 VTAIL.n310 VSUBS 0.014664f
C952 VTAIL.n311 VSUBS 0.025774f
C953 VTAIL.n312 VSUBS 0.01385f
C954 VTAIL.n313 VSUBS 0.024552f
C955 VTAIL.n314 VSUBS 0.024625f
C956 VTAIL.t1 VSUBS 0.070333f
C957 VTAIL.n315 VSUBS 0.156601f
C958 VTAIL.n316 VSUBS 0.815494f
C959 VTAIL.n317 VSUBS 0.01385f
C960 VTAIL.n318 VSUBS 0.014664f
C961 VTAIL.n319 VSUBS 0.032736f
C962 VTAIL.n320 VSUBS 0.032736f
C963 VTAIL.n321 VSUBS 0.014664f
C964 VTAIL.n322 VSUBS 0.01385f
C965 VTAIL.n323 VSUBS 0.025774f
C966 VTAIL.n324 VSUBS 0.025774f
C967 VTAIL.n325 VSUBS 0.01385f
C968 VTAIL.n326 VSUBS 0.014664f
C969 VTAIL.n327 VSUBS 0.032736f
C970 VTAIL.n328 VSUBS 0.032736f
C971 VTAIL.n329 VSUBS 0.014664f
C972 VTAIL.n330 VSUBS 0.01385f
C973 VTAIL.n331 VSUBS 0.025774f
C974 VTAIL.n332 VSUBS 0.025774f
C975 VTAIL.n333 VSUBS 0.01385f
C976 VTAIL.n334 VSUBS 0.01385f
C977 VTAIL.n335 VSUBS 0.014664f
C978 VTAIL.n336 VSUBS 0.032736f
C979 VTAIL.n337 VSUBS 0.032736f
C980 VTAIL.n338 VSUBS 0.077766f
C981 VTAIL.n339 VSUBS 0.014257f
C982 VTAIL.n340 VSUBS 0.01385f
C983 VTAIL.n341 VSUBS 0.066969f
C984 VTAIL.n342 VSUBS 0.039257f
C985 VTAIL.n343 VSUBS 1.16401f
C986 VDD1.t1 VSUBS 0.161361f
C987 VDD1.t5 VSUBS 0.161361f
C988 VDD1.n0 VSUBS 1.17778f
C989 VDD1.t4 VSUBS 0.161361f
C990 VDD1.t3 VSUBS 0.161361f
C991 VDD1.n1 VSUBS 1.17693f
C992 VDD1.t0 VSUBS 0.161361f
C993 VDD1.t7 VSUBS 0.161361f
C994 VDD1.n2 VSUBS 1.17693f
C995 VDD1.n3 VSUBS 2.75338f
C996 VDD1.t6 VSUBS 0.161361f
C997 VDD1.t2 VSUBS 0.161361f
C998 VDD1.n4 VSUBS 1.17279f
C999 VDD1.n5 VSUBS 2.44292f
C1000 VP.n0 VSUBS 0.064172f
C1001 VP.t4 VSUBS 1.24154f
C1002 VP.n1 VSUBS 0.476062f
C1003 VP.n2 VSUBS 0.048091f
C1004 VP.t2 VSUBS 1.24154f
C1005 VP.n3 VSUBS 0.476062f
C1006 VP.n4 VSUBS 0.064172f
C1007 VP.n5 VSUBS 0.064172f
C1008 VP.t1 VSUBS 1.32995f
C1009 VP.t0 VSUBS 1.24154f
C1010 VP.n6 VSUBS 0.476062f
C1011 VP.n7 VSUBS 0.048091f
C1012 VP.t6 VSUBS 1.24154f
C1013 VP.n8 VSUBS 0.537042f
C1014 VP.t3 VSUBS 1.38006f
C1015 VP.n9 VSUBS 0.556382f
C1016 VP.n10 VSUBS 0.246871f
C1017 VP.n11 VSUBS 0.074781f
C1018 VP.n12 VSUBS 0.038877f
C1019 VP.n13 VSUBS 0.074781f
C1020 VP.n14 VSUBS 0.048091f
C1021 VP.n15 VSUBS 0.048091f
C1022 VP.n16 VSUBS 0.073274f
C1023 VP.n17 VSUBS 0.028168f
C1024 VP.n18 VSUBS 0.563846f
C1025 VP.n19 VSUBS 1.95752f
C1026 VP.n20 VSUBS 1.99925f
C1027 VP.t7 VSUBS 1.32995f
C1028 VP.n21 VSUBS 0.563846f
C1029 VP.n22 VSUBS 0.028168f
C1030 VP.n23 VSUBS 0.073274f
C1031 VP.n24 VSUBS 0.048091f
C1032 VP.n25 VSUBS 0.048091f
C1033 VP.n26 VSUBS 0.074781f
C1034 VP.n27 VSUBS 0.038877f
C1035 VP.n28 VSUBS 0.074781f
C1036 VP.n29 VSUBS 0.048091f
C1037 VP.n30 VSUBS 0.048091f
C1038 VP.n31 VSUBS 0.073274f
C1039 VP.n32 VSUBS 0.028168f
C1040 VP.t5 VSUBS 1.32995f
C1041 VP.n33 VSUBS 0.563846f
C1042 VP.n34 VSUBS 0.045039f
.ends

