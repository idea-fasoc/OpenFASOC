* NGSPICE file created from diff_pair_sample_1156.ext - technology: sky130A

.subckt diff_pair_sample_1156 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t18 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=5.0427 ps=26.64 w=12.93 l=2.11
X1 VTAIL.t0 VN.t0 VDD2.t9 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X2 VDD1.t8 VP.t1 VTAIL.t19 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=5.0427 pd=26.64 as=2.13345 ps=13.26 w=12.93 l=2.11
X3 VTAIL.t1 VN.t1 VDD2.t8 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X4 VTAIL.t13 VP.t2 VDD1.t7 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X5 VDD1.t6 VP.t3 VTAIL.t16 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=5.0427 ps=26.64 w=12.93 l=2.11
X6 VTAIL.t11 VP.t4 VDD1.t5 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X7 VDD2.t7 VN.t2 VTAIL.t3 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X8 VTAIL.t14 VP.t5 VDD1.t4 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X9 VDD2.t6 VN.t3 VTAIL.t2 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=5.0427 ps=26.64 w=12.93 l=2.11
X10 VDD2.t5 VN.t4 VTAIL.t7 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=5.0427 ps=26.64 w=12.93 l=2.11
X11 VDD2.t4 VN.t5 VTAIL.t5 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=5.0427 pd=26.64 as=2.13345 ps=13.26 w=12.93 l=2.11
X12 B.t11 B.t9 B.t10 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=5.0427 pd=26.64 as=0 ps=0 w=12.93 l=2.11
X13 VDD1.t3 VP.t6 VTAIL.t12 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X14 VTAIL.t4 VN.t6 VDD2.t3 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X15 VTAIL.t6 VN.t7 VDD2.t2 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X16 VDD1.t2 VP.t7 VTAIL.t10 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X17 B.t8 B.t6 B.t7 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=5.0427 pd=26.64 as=0 ps=0 w=12.93 l=2.11
X18 B.t5 B.t3 B.t4 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=5.0427 pd=26.64 as=0 ps=0 w=12.93 l=2.11
X19 VDD2.t1 VN.t8 VTAIL.t9 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X20 VDD2.t0 VN.t9 VTAIL.t8 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=5.0427 pd=26.64 as=2.13345 ps=13.26 w=12.93 l=2.11
X21 VTAIL.t17 VP.t8 VDD1.t1 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=2.13345 pd=13.26 as=2.13345 ps=13.26 w=12.93 l=2.11
X22 B.t2 B.t0 B.t1 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=5.0427 pd=26.64 as=0 ps=0 w=12.93 l=2.11
X23 VDD1.t0 VP.t9 VTAIL.t15 w_n3898_n3554# sky130_fd_pr__pfet_01v8 ad=5.0427 pd=26.64 as=2.13345 ps=13.26 w=12.93 l=2.11
R0 VP.n18 VP.t9 181.585
R1 VP.n20 VP.n19 161.3
R2 VP.n21 VP.n16 161.3
R3 VP.n23 VP.n22 161.3
R4 VP.n24 VP.n15 161.3
R5 VP.n26 VP.n25 161.3
R6 VP.n27 VP.n14 161.3
R7 VP.n29 VP.n28 161.3
R8 VP.n30 VP.n13 161.3
R9 VP.n32 VP.n31 161.3
R10 VP.n34 VP.n12 161.3
R11 VP.n36 VP.n35 161.3
R12 VP.n37 VP.n11 161.3
R13 VP.n39 VP.n38 161.3
R14 VP.n40 VP.n10 161.3
R15 VP.n74 VP.n0 161.3
R16 VP.n73 VP.n72 161.3
R17 VP.n71 VP.n1 161.3
R18 VP.n70 VP.n69 161.3
R19 VP.n68 VP.n2 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n64 VP.n3 161.3
R22 VP.n63 VP.n62 161.3
R23 VP.n61 VP.n4 161.3
R24 VP.n60 VP.n59 161.3
R25 VP.n58 VP.n5 161.3
R26 VP.n57 VP.n56 161.3
R27 VP.n55 VP.n6 161.3
R28 VP.n54 VP.n53 161.3
R29 VP.n52 VP.n51 161.3
R30 VP.n50 VP.n8 161.3
R31 VP.n49 VP.n48 161.3
R32 VP.n47 VP.n9 161.3
R33 VP.n46 VP.n45 161.3
R34 VP.n60 VP.t7 147.685
R35 VP.n44 VP.t1 147.685
R36 VP.n7 VP.t2 147.685
R37 VP.n67 VP.t5 147.685
R38 VP.n75 VP.t0 147.685
R39 VP.n26 VP.t6 147.685
R40 VP.n41 VP.t3 147.685
R41 VP.n33 VP.t8 147.685
R42 VP.n17 VP.t4 147.685
R43 VP.n44 VP.n43 92.1615
R44 VP.n76 VP.n75 92.1615
R45 VP.n42 VP.n41 92.1615
R46 VP.n56 VP.n55 56.5193
R47 VP.n62 VP.n3 56.5193
R48 VP.n28 VP.n13 56.5193
R49 VP.n22 VP.n21 56.5193
R50 VP.n49 VP.n9 56.0336
R51 VP.n73 VP.n1 56.0336
R52 VP.n39 VP.n11 56.0336
R53 VP.n43 VP.n42 51.189
R54 VP.n18 VP.n17 48.9316
R55 VP.n50 VP.n49 24.9531
R56 VP.n69 VP.n1 24.9531
R57 VP.n35 VP.n11 24.9531
R58 VP.n45 VP.n9 24.4675
R59 VP.n51 VP.n50 24.4675
R60 VP.n55 VP.n54 24.4675
R61 VP.n56 VP.n5 24.4675
R62 VP.n60 VP.n5 24.4675
R63 VP.n61 VP.n60 24.4675
R64 VP.n62 VP.n61 24.4675
R65 VP.n66 VP.n3 24.4675
R66 VP.n69 VP.n68 24.4675
R67 VP.n74 VP.n73 24.4675
R68 VP.n40 VP.n39 24.4675
R69 VP.n32 VP.n13 24.4675
R70 VP.n35 VP.n34 24.4675
R71 VP.n22 VP.n15 24.4675
R72 VP.n26 VP.n15 24.4675
R73 VP.n27 VP.n26 24.4675
R74 VP.n28 VP.n27 24.4675
R75 VP.n21 VP.n20 24.4675
R76 VP.n54 VP.n7 21.5315
R77 VP.n67 VP.n66 21.5315
R78 VP.n33 VP.n32 21.5315
R79 VP.n20 VP.n17 21.5315
R80 VP.n45 VP.n44 18.5954
R81 VP.n75 VP.n74 18.5954
R82 VP.n41 VP.n40 18.5954
R83 VP.n19 VP.n18 9.10118
R84 VP.n51 VP.n7 2.93654
R85 VP.n68 VP.n67 2.93654
R86 VP.n34 VP.n33 2.93654
R87 VP.n42 VP.n10 0.278367
R88 VP.n46 VP.n43 0.278367
R89 VP.n76 VP.n0 0.278367
R90 VP.n19 VP.n16 0.189894
R91 VP.n23 VP.n16 0.189894
R92 VP.n24 VP.n23 0.189894
R93 VP.n25 VP.n24 0.189894
R94 VP.n25 VP.n14 0.189894
R95 VP.n29 VP.n14 0.189894
R96 VP.n30 VP.n29 0.189894
R97 VP.n31 VP.n30 0.189894
R98 VP.n31 VP.n12 0.189894
R99 VP.n36 VP.n12 0.189894
R100 VP.n37 VP.n36 0.189894
R101 VP.n38 VP.n37 0.189894
R102 VP.n38 VP.n10 0.189894
R103 VP.n47 VP.n46 0.189894
R104 VP.n48 VP.n47 0.189894
R105 VP.n48 VP.n8 0.189894
R106 VP.n52 VP.n8 0.189894
R107 VP.n53 VP.n52 0.189894
R108 VP.n53 VP.n6 0.189894
R109 VP.n57 VP.n6 0.189894
R110 VP.n58 VP.n57 0.189894
R111 VP.n59 VP.n58 0.189894
R112 VP.n59 VP.n4 0.189894
R113 VP.n63 VP.n4 0.189894
R114 VP.n64 VP.n63 0.189894
R115 VP.n65 VP.n64 0.189894
R116 VP.n65 VP.n2 0.189894
R117 VP.n70 VP.n2 0.189894
R118 VP.n71 VP.n70 0.189894
R119 VP.n72 VP.n71 0.189894
R120 VP.n72 VP.n0 0.189894
R121 VP VP.n76 0.153454
R122 VTAIL.n11 VTAIL.t2 59.8903
R123 VTAIL.n17 VTAIL.t7 59.8892
R124 VTAIL.n2 VTAIL.t18 59.8892
R125 VTAIL.n16 VTAIL.t16 59.8892
R126 VTAIL.n15 VTAIL.n14 57.3765
R127 VTAIL.n13 VTAIL.n12 57.3765
R128 VTAIL.n10 VTAIL.n9 57.3765
R129 VTAIL.n8 VTAIL.n7 57.3765
R130 VTAIL.n19 VTAIL.n18 57.3753
R131 VTAIL.n1 VTAIL.n0 57.3753
R132 VTAIL.n4 VTAIL.n3 57.3753
R133 VTAIL.n6 VTAIL.n5 57.3753
R134 VTAIL.n8 VTAIL.n6 27.7203
R135 VTAIL.n17 VTAIL.n16 25.6169
R136 VTAIL.n18 VTAIL.t9 2.51442
R137 VTAIL.n18 VTAIL.t0 2.51442
R138 VTAIL.n0 VTAIL.t8 2.51442
R139 VTAIL.n0 VTAIL.t1 2.51442
R140 VTAIL.n3 VTAIL.t10 2.51442
R141 VTAIL.n3 VTAIL.t14 2.51442
R142 VTAIL.n5 VTAIL.t19 2.51442
R143 VTAIL.n5 VTAIL.t13 2.51442
R144 VTAIL.n14 VTAIL.t12 2.51442
R145 VTAIL.n14 VTAIL.t17 2.51442
R146 VTAIL.n12 VTAIL.t15 2.51442
R147 VTAIL.n12 VTAIL.t11 2.51442
R148 VTAIL.n9 VTAIL.t3 2.51442
R149 VTAIL.n9 VTAIL.t6 2.51442
R150 VTAIL.n7 VTAIL.t5 2.51442
R151 VTAIL.n7 VTAIL.t4 2.51442
R152 VTAIL.n10 VTAIL.n8 2.10395
R153 VTAIL.n11 VTAIL.n10 2.10395
R154 VTAIL.n15 VTAIL.n13 2.10395
R155 VTAIL.n16 VTAIL.n15 2.10395
R156 VTAIL.n6 VTAIL.n4 2.10395
R157 VTAIL.n4 VTAIL.n2 2.10395
R158 VTAIL.n19 VTAIL.n17 2.10395
R159 VTAIL VTAIL.n1 1.63628
R160 VTAIL.n13 VTAIL.n11 1.52205
R161 VTAIL.n2 VTAIL.n1 1.52205
R162 VTAIL VTAIL.n19 0.468172
R163 VDD1.n1 VDD1.t0 78.6726
R164 VDD1.n3 VDD1.t8 78.6714
R165 VDD1.n5 VDD1.n4 75.5763
R166 VDD1.n1 VDD1.n0 74.0552
R167 VDD1.n7 VDD1.n6 74.0541
R168 VDD1.n3 VDD1.n2 74.054
R169 VDD1.n7 VDD1.n5 46.488
R170 VDD1.n6 VDD1.t1 2.51442
R171 VDD1.n6 VDD1.t6 2.51442
R172 VDD1.n0 VDD1.t5 2.51442
R173 VDD1.n0 VDD1.t3 2.51442
R174 VDD1.n4 VDD1.t4 2.51442
R175 VDD1.n4 VDD1.t9 2.51442
R176 VDD1.n2 VDD1.t7 2.51442
R177 VDD1.n2 VDD1.t2 2.51442
R178 VDD1 VDD1.n7 1.5199
R179 VDD1 VDD1.n1 0.584552
R180 VDD1.n5 VDD1.n3 0.471016
R181 VN.n8 VN.t9 181.585
R182 VN.n41 VN.t3 181.585
R183 VN.n63 VN.n33 161.3
R184 VN.n62 VN.n61 161.3
R185 VN.n60 VN.n34 161.3
R186 VN.n59 VN.n58 161.3
R187 VN.n57 VN.n35 161.3
R188 VN.n55 VN.n54 161.3
R189 VN.n53 VN.n36 161.3
R190 VN.n52 VN.n51 161.3
R191 VN.n50 VN.n37 161.3
R192 VN.n49 VN.n48 161.3
R193 VN.n47 VN.n38 161.3
R194 VN.n46 VN.n45 161.3
R195 VN.n44 VN.n39 161.3
R196 VN.n43 VN.n42 161.3
R197 VN.n30 VN.n0 161.3
R198 VN.n29 VN.n28 161.3
R199 VN.n27 VN.n1 161.3
R200 VN.n26 VN.n25 161.3
R201 VN.n24 VN.n2 161.3
R202 VN.n22 VN.n21 161.3
R203 VN.n20 VN.n3 161.3
R204 VN.n19 VN.n18 161.3
R205 VN.n17 VN.n4 161.3
R206 VN.n16 VN.n15 161.3
R207 VN.n14 VN.n5 161.3
R208 VN.n13 VN.n12 161.3
R209 VN.n11 VN.n6 161.3
R210 VN.n10 VN.n9 161.3
R211 VN.n16 VN.t8 147.685
R212 VN.n7 VN.t1 147.685
R213 VN.n23 VN.t0 147.685
R214 VN.n31 VN.t4 147.685
R215 VN.n49 VN.t2 147.685
R216 VN.n40 VN.t7 147.685
R217 VN.n56 VN.t6 147.685
R218 VN.n64 VN.t5 147.685
R219 VN.n32 VN.n31 92.1615
R220 VN.n65 VN.n64 92.1615
R221 VN.n12 VN.n11 56.5193
R222 VN.n18 VN.n3 56.5193
R223 VN.n45 VN.n44 56.5193
R224 VN.n51 VN.n36 56.5193
R225 VN.n29 VN.n1 56.0336
R226 VN.n62 VN.n34 56.0336
R227 VN VN.n65 51.4678
R228 VN.n8 VN.n7 48.9316
R229 VN.n41 VN.n40 48.9316
R230 VN.n25 VN.n1 24.9531
R231 VN.n58 VN.n34 24.9531
R232 VN.n11 VN.n10 24.4675
R233 VN.n12 VN.n5 24.4675
R234 VN.n16 VN.n5 24.4675
R235 VN.n17 VN.n16 24.4675
R236 VN.n18 VN.n17 24.4675
R237 VN.n22 VN.n3 24.4675
R238 VN.n25 VN.n24 24.4675
R239 VN.n30 VN.n29 24.4675
R240 VN.n44 VN.n43 24.4675
R241 VN.n51 VN.n50 24.4675
R242 VN.n50 VN.n49 24.4675
R243 VN.n49 VN.n38 24.4675
R244 VN.n45 VN.n38 24.4675
R245 VN.n58 VN.n57 24.4675
R246 VN.n55 VN.n36 24.4675
R247 VN.n63 VN.n62 24.4675
R248 VN.n10 VN.n7 21.5315
R249 VN.n23 VN.n22 21.5315
R250 VN.n43 VN.n40 21.5315
R251 VN.n56 VN.n55 21.5315
R252 VN.n31 VN.n30 18.5954
R253 VN.n64 VN.n63 18.5954
R254 VN.n42 VN.n41 9.10118
R255 VN.n9 VN.n8 9.10118
R256 VN.n24 VN.n23 2.93654
R257 VN.n57 VN.n56 2.93654
R258 VN.n65 VN.n33 0.278367
R259 VN.n32 VN.n0 0.278367
R260 VN.n61 VN.n33 0.189894
R261 VN.n61 VN.n60 0.189894
R262 VN.n60 VN.n59 0.189894
R263 VN.n59 VN.n35 0.189894
R264 VN.n54 VN.n35 0.189894
R265 VN.n54 VN.n53 0.189894
R266 VN.n53 VN.n52 0.189894
R267 VN.n52 VN.n37 0.189894
R268 VN.n48 VN.n37 0.189894
R269 VN.n48 VN.n47 0.189894
R270 VN.n47 VN.n46 0.189894
R271 VN.n46 VN.n39 0.189894
R272 VN.n42 VN.n39 0.189894
R273 VN.n9 VN.n6 0.189894
R274 VN.n13 VN.n6 0.189894
R275 VN.n14 VN.n13 0.189894
R276 VN.n15 VN.n14 0.189894
R277 VN.n15 VN.n4 0.189894
R278 VN.n19 VN.n4 0.189894
R279 VN.n20 VN.n19 0.189894
R280 VN.n21 VN.n20 0.189894
R281 VN.n21 VN.n2 0.189894
R282 VN.n26 VN.n2 0.189894
R283 VN.n27 VN.n26 0.189894
R284 VN.n28 VN.n27 0.189894
R285 VN.n28 VN.n0 0.189894
R286 VN VN.n32 0.153454
R287 VDD2.n1 VDD2.t0 78.6714
R288 VDD2.n4 VDD2.t4 76.5691
R289 VDD2.n3 VDD2.n2 75.5763
R290 VDD2 VDD2.n7 75.5735
R291 VDD2.n6 VDD2.n5 74.0552
R292 VDD2.n1 VDD2.n0 74.054
R293 VDD2.n4 VDD2.n3 44.8532
R294 VDD2.n7 VDD2.t2 2.51442
R295 VDD2.n7 VDD2.t6 2.51442
R296 VDD2.n5 VDD2.t3 2.51442
R297 VDD2.n5 VDD2.t7 2.51442
R298 VDD2.n2 VDD2.t9 2.51442
R299 VDD2.n2 VDD2.t5 2.51442
R300 VDD2.n0 VDD2.t8 2.51442
R301 VDD2.n0 VDD2.t1 2.51442
R302 VDD2.n6 VDD2.n4 2.10395
R303 VDD2 VDD2.n6 0.584552
R304 VDD2.n3 VDD2.n1 0.471016
R305 B.n590 B.n81 585
R306 B.n592 B.n591 585
R307 B.n593 B.n80 585
R308 B.n595 B.n594 585
R309 B.n596 B.n79 585
R310 B.n598 B.n597 585
R311 B.n599 B.n78 585
R312 B.n601 B.n600 585
R313 B.n602 B.n77 585
R314 B.n604 B.n603 585
R315 B.n605 B.n76 585
R316 B.n607 B.n606 585
R317 B.n608 B.n75 585
R318 B.n610 B.n609 585
R319 B.n611 B.n74 585
R320 B.n613 B.n612 585
R321 B.n614 B.n73 585
R322 B.n616 B.n615 585
R323 B.n617 B.n72 585
R324 B.n619 B.n618 585
R325 B.n620 B.n71 585
R326 B.n622 B.n621 585
R327 B.n623 B.n70 585
R328 B.n625 B.n624 585
R329 B.n626 B.n69 585
R330 B.n628 B.n627 585
R331 B.n629 B.n68 585
R332 B.n631 B.n630 585
R333 B.n632 B.n67 585
R334 B.n634 B.n633 585
R335 B.n635 B.n66 585
R336 B.n637 B.n636 585
R337 B.n638 B.n65 585
R338 B.n640 B.n639 585
R339 B.n641 B.n64 585
R340 B.n643 B.n642 585
R341 B.n644 B.n63 585
R342 B.n646 B.n645 585
R343 B.n647 B.n62 585
R344 B.n649 B.n648 585
R345 B.n650 B.n61 585
R346 B.n652 B.n651 585
R347 B.n653 B.n57 585
R348 B.n655 B.n654 585
R349 B.n656 B.n56 585
R350 B.n658 B.n657 585
R351 B.n659 B.n55 585
R352 B.n661 B.n660 585
R353 B.n662 B.n54 585
R354 B.n664 B.n663 585
R355 B.n665 B.n53 585
R356 B.n667 B.n666 585
R357 B.n668 B.n52 585
R358 B.n670 B.n669 585
R359 B.n672 B.n49 585
R360 B.n674 B.n673 585
R361 B.n675 B.n48 585
R362 B.n677 B.n676 585
R363 B.n678 B.n47 585
R364 B.n680 B.n679 585
R365 B.n681 B.n46 585
R366 B.n683 B.n682 585
R367 B.n684 B.n45 585
R368 B.n686 B.n685 585
R369 B.n687 B.n44 585
R370 B.n689 B.n688 585
R371 B.n690 B.n43 585
R372 B.n692 B.n691 585
R373 B.n693 B.n42 585
R374 B.n695 B.n694 585
R375 B.n696 B.n41 585
R376 B.n698 B.n697 585
R377 B.n699 B.n40 585
R378 B.n701 B.n700 585
R379 B.n702 B.n39 585
R380 B.n704 B.n703 585
R381 B.n705 B.n38 585
R382 B.n707 B.n706 585
R383 B.n708 B.n37 585
R384 B.n710 B.n709 585
R385 B.n711 B.n36 585
R386 B.n713 B.n712 585
R387 B.n714 B.n35 585
R388 B.n716 B.n715 585
R389 B.n717 B.n34 585
R390 B.n719 B.n718 585
R391 B.n720 B.n33 585
R392 B.n722 B.n721 585
R393 B.n723 B.n32 585
R394 B.n725 B.n724 585
R395 B.n726 B.n31 585
R396 B.n728 B.n727 585
R397 B.n729 B.n30 585
R398 B.n731 B.n730 585
R399 B.n732 B.n29 585
R400 B.n734 B.n733 585
R401 B.n735 B.n28 585
R402 B.n737 B.n736 585
R403 B.n589 B.n588 585
R404 B.n587 B.n82 585
R405 B.n586 B.n585 585
R406 B.n584 B.n83 585
R407 B.n583 B.n582 585
R408 B.n581 B.n84 585
R409 B.n580 B.n579 585
R410 B.n578 B.n85 585
R411 B.n577 B.n576 585
R412 B.n575 B.n86 585
R413 B.n574 B.n573 585
R414 B.n572 B.n87 585
R415 B.n571 B.n570 585
R416 B.n569 B.n88 585
R417 B.n568 B.n567 585
R418 B.n566 B.n89 585
R419 B.n565 B.n564 585
R420 B.n563 B.n90 585
R421 B.n562 B.n561 585
R422 B.n560 B.n91 585
R423 B.n559 B.n558 585
R424 B.n557 B.n92 585
R425 B.n556 B.n555 585
R426 B.n554 B.n93 585
R427 B.n553 B.n552 585
R428 B.n551 B.n94 585
R429 B.n550 B.n549 585
R430 B.n548 B.n95 585
R431 B.n547 B.n546 585
R432 B.n545 B.n96 585
R433 B.n544 B.n543 585
R434 B.n542 B.n97 585
R435 B.n541 B.n540 585
R436 B.n539 B.n98 585
R437 B.n538 B.n537 585
R438 B.n536 B.n99 585
R439 B.n535 B.n534 585
R440 B.n533 B.n100 585
R441 B.n532 B.n531 585
R442 B.n530 B.n101 585
R443 B.n529 B.n528 585
R444 B.n527 B.n102 585
R445 B.n526 B.n525 585
R446 B.n524 B.n103 585
R447 B.n523 B.n522 585
R448 B.n521 B.n104 585
R449 B.n520 B.n519 585
R450 B.n518 B.n105 585
R451 B.n517 B.n516 585
R452 B.n515 B.n106 585
R453 B.n514 B.n513 585
R454 B.n512 B.n107 585
R455 B.n511 B.n510 585
R456 B.n509 B.n108 585
R457 B.n508 B.n507 585
R458 B.n506 B.n109 585
R459 B.n505 B.n504 585
R460 B.n503 B.n110 585
R461 B.n502 B.n501 585
R462 B.n500 B.n111 585
R463 B.n499 B.n498 585
R464 B.n497 B.n112 585
R465 B.n496 B.n495 585
R466 B.n494 B.n113 585
R467 B.n493 B.n492 585
R468 B.n491 B.n114 585
R469 B.n490 B.n489 585
R470 B.n488 B.n115 585
R471 B.n487 B.n486 585
R472 B.n485 B.n116 585
R473 B.n484 B.n483 585
R474 B.n482 B.n117 585
R475 B.n481 B.n480 585
R476 B.n479 B.n118 585
R477 B.n478 B.n477 585
R478 B.n476 B.n119 585
R479 B.n475 B.n474 585
R480 B.n473 B.n120 585
R481 B.n472 B.n471 585
R482 B.n470 B.n121 585
R483 B.n469 B.n468 585
R484 B.n467 B.n122 585
R485 B.n466 B.n465 585
R486 B.n464 B.n123 585
R487 B.n463 B.n462 585
R488 B.n461 B.n124 585
R489 B.n460 B.n459 585
R490 B.n458 B.n125 585
R491 B.n457 B.n456 585
R492 B.n455 B.n126 585
R493 B.n454 B.n453 585
R494 B.n452 B.n127 585
R495 B.n451 B.n450 585
R496 B.n449 B.n128 585
R497 B.n448 B.n447 585
R498 B.n446 B.n129 585
R499 B.n445 B.n444 585
R500 B.n443 B.n130 585
R501 B.n442 B.n441 585
R502 B.n440 B.n131 585
R503 B.n439 B.n438 585
R504 B.n437 B.n132 585
R505 B.n436 B.n435 585
R506 B.n287 B.n186 585
R507 B.n289 B.n288 585
R508 B.n290 B.n185 585
R509 B.n292 B.n291 585
R510 B.n293 B.n184 585
R511 B.n295 B.n294 585
R512 B.n296 B.n183 585
R513 B.n298 B.n297 585
R514 B.n299 B.n182 585
R515 B.n301 B.n300 585
R516 B.n302 B.n181 585
R517 B.n304 B.n303 585
R518 B.n305 B.n180 585
R519 B.n307 B.n306 585
R520 B.n308 B.n179 585
R521 B.n310 B.n309 585
R522 B.n311 B.n178 585
R523 B.n313 B.n312 585
R524 B.n314 B.n177 585
R525 B.n316 B.n315 585
R526 B.n317 B.n176 585
R527 B.n319 B.n318 585
R528 B.n320 B.n175 585
R529 B.n322 B.n321 585
R530 B.n323 B.n174 585
R531 B.n325 B.n324 585
R532 B.n326 B.n173 585
R533 B.n328 B.n327 585
R534 B.n329 B.n172 585
R535 B.n331 B.n330 585
R536 B.n332 B.n171 585
R537 B.n334 B.n333 585
R538 B.n335 B.n170 585
R539 B.n337 B.n336 585
R540 B.n338 B.n169 585
R541 B.n340 B.n339 585
R542 B.n341 B.n168 585
R543 B.n343 B.n342 585
R544 B.n344 B.n167 585
R545 B.n346 B.n345 585
R546 B.n347 B.n166 585
R547 B.n349 B.n348 585
R548 B.n350 B.n165 585
R549 B.n352 B.n351 585
R550 B.n354 B.n162 585
R551 B.n356 B.n355 585
R552 B.n357 B.n161 585
R553 B.n359 B.n358 585
R554 B.n360 B.n160 585
R555 B.n362 B.n361 585
R556 B.n363 B.n159 585
R557 B.n365 B.n364 585
R558 B.n366 B.n158 585
R559 B.n368 B.n367 585
R560 B.n370 B.n369 585
R561 B.n371 B.n154 585
R562 B.n373 B.n372 585
R563 B.n374 B.n153 585
R564 B.n376 B.n375 585
R565 B.n377 B.n152 585
R566 B.n379 B.n378 585
R567 B.n380 B.n151 585
R568 B.n382 B.n381 585
R569 B.n383 B.n150 585
R570 B.n385 B.n384 585
R571 B.n386 B.n149 585
R572 B.n388 B.n387 585
R573 B.n389 B.n148 585
R574 B.n391 B.n390 585
R575 B.n392 B.n147 585
R576 B.n394 B.n393 585
R577 B.n395 B.n146 585
R578 B.n397 B.n396 585
R579 B.n398 B.n145 585
R580 B.n400 B.n399 585
R581 B.n401 B.n144 585
R582 B.n403 B.n402 585
R583 B.n404 B.n143 585
R584 B.n406 B.n405 585
R585 B.n407 B.n142 585
R586 B.n409 B.n408 585
R587 B.n410 B.n141 585
R588 B.n412 B.n411 585
R589 B.n413 B.n140 585
R590 B.n415 B.n414 585
R591 B.n416 B.n139 585
R592 B.n418 B.n417 585
R593 B.n419 B.n138 585
R594 B.n421 B.n420 585
R595 B.n422 B.n137 585
R596 B.n424 B.n423 585
R597 B.n425 B.n136 585
R598 B.n427 B.n426 585
R599 B.n428 B.n135 585
R600 B.n430 B.n429 585
R601 B.n431 B.n134 585
R602 B.n433 B.n432 585
R603 B.n434 B.n133 585
R604 B.n286 B.n285 585
R605 B.n284 B.n187 585
R606 B.n283 B.n282 585
R607 B.n281 B.n188 585
R608 B.n280 B.n279 585
R609 B.n278 B.n189 585
R610 B.n277 B.n276 585
R611 B.n275 B.n190 585
R612 B.n274 B.n273 585
R613 B.n272 B.n191 585
R614 B.n271 B.n270 585
R615 B.n269 B.n192 585
R616 B.n268 B.n267 585
R617 B.n266 B.n193 585
R618 B.n265 B.n264 585
R619 B.n263 B.n194 585
R620 B.n262 B.n261 585
R621 B.n260 B.n195 585
R622 B.n259 B.n258 585
R623 B.n257 B.n196 585
R624 B.n256 B.n255 585
R625 B.n254 B.n197 585
R626 B.n253 B.n252 585
R627 B.n251 B.n198 585
R628 B.n250 B.n249 585
R629 B.n248 B.n199 585
R630 B.n247 B.n246 585
R631 B.n245 B.n200 585
R632 B.n244 B.n243 585
R633 B.n242 B.n201 585
R634 B.n241 B.n240 585
R635 B.n239 B.n202 585
R636 B.n238 B.n237 585
R637 B.n236 B.n203 585
R638 B.n235 B.n234 585
R639 B.n233 B.n204 585
R640 B.n232 B.n231 585
R641 B.n230 B.n205 585
R642 B.n229 B.n228 585
R643 B.n227 B.n206 585
R644 B.n226 B.n225 585
R645 B.n224 B.n207 585
R646 B.n223 B.n222 585
R647 B.n221 B.n208 585
R648 B.n220 B.n219 585
R649 B.n218 B.n209 585
R650 B.n217 B.n216 585
R651 B.n215 B.n210 585
R652 B.n214 B.n213 585
R653 B.n212 B.n211 585
R654 B.n2 B.n0 585
R655 B.n813 B.n1 585
R656 B.n812 B.n811 585
R657 B.n810 B.n3 585
R658 B.n809 B.n808 585
R659 B.n807 B.n4 585
R660 B.n806 B.n805 585
R661 B.n804 B.n5 585
R662 B.n803 B.n802 585
R663 B.n801 B.n6 585
R664 B.n800 B.n799 585
R665 B.n798 B.n7 585
R666 B.n797 B.n796 585
R667 B.n795 B.n8 585
R668 B.n794 B.n793 585
R669 B.n792 B.n9 585
R670 B.n791 B.n790 585
R671 B.n789 B.n10 585
R672 B.n788 B.n787 585
R673 B.n786 B.n11 585
R674 B.n785 B.n784 585
R675 B.n783 B.n12 585
R676 B.n782 B.n781 585
R677 B.n780 B.n13 585
R678 B.n779 B.n778 585
R679 B.n777 B.n14 585
R680 B.n776 B.n775 585
R681 B.n774 B.n15 585
R682 B.n773 B.n772 585
R683 B.n771 B.n16 585
R684 B.n770 B.n769 585
R685 B.n768 B.n17 585
R686 B.n767 B.n766 585
R687 B.n765 B.n18 585
R688 B.n764 B.n763 585
R689 B.n762 B.n19 585
R690 B.n761 B.n760 585
R691 B.n759 B.n20 585
R692 B.n758 B.n757 585
R693 B.n756 B.n21 585
R694 B.n755 B.n754 585
R695 B.n753 B.n22 585
R696 B.n752 B.n751 585
R697 B.n750 B.n23 585
R698 B.n749 B.n748 585
R699 B.n747 B.n24 585
R700 B.n746 B.n745 585
R701 B.n744 B.n25 585
R702 B.n743 B.n742 585
R703 B.n741 B.n26 585
R704 B.n740 B.n739 585
R705 B.n738 B.n27 585
R706 B.n815 B.n814 585
R707 B.n285 B.n186 550.159
R708 B.n736 B.n27 550.159
R709 B.n435 B.n434 550.159
R710 B.n590 B.n589 550.159
R711 B.n155 B.t6 354.849
R712 B.n163 B.t3 354.849
R713 B.n50 B.t0 354.849
R714 B.n58 B.t9 354.849
R715 B.n285 B.n284 163.367
R716 B.n284 B.n283 163.367
R717 B.n283 B.n188 163.367
R718 B.n279 B.n188 163.367
R719 B.n279 B.n278 163.367
R720 B.n278 B.n277 163.367
R721 B.n277 B.n190 163.367
R722 B.n273 B.n190 163.367
R723 B.n273 B.n272 163.367
R724 B.n272 B.n271 163.367
R725 B.n271 B.n192 163.367
R726 B.n267 B.n192 163.367
R727 B.n267 B.n266 163.367
R728 B.n266 B.n265 163.367
R729 B.n265 B.n194 163.367
R730 B.n261 B.n194 163.367
R731 B.n261 B.n260 163.367
R732 B.n260 B.n259 163.367
R733 B.n259 B.n196 163.367
R734 B.n255 B.n196 163.367
R735 B.n255 B.n254 163.367
R736 B.n254 B.n253 163.367
R737 B.n253 B.n198 163.367
R738 B.n249 B.n198 163.367
R739 B.n249 B.n248 163.367
R740 B.n248 B.n247 163.367
R741 B.n247 B.n200 163.367
R742 B.n243 B.n200 163.367
R743 B.n243 B.n242 163.367
R744 B.n242 B.n241 163.367
R745 B.n241 B.n202 163.367
R746 B.n237 B.n202 163.367
R747 B.n237 B.n236 163.367
R748 B.n236 B.n235 163.367
R749 B.n235 B.n204 163.367
R750 B.n231 B.n204 163.367
R751 B.n231 B.n230 163.367
R752 B.n230 B.n229 163.367
R753 B.n229 B.n206 163.367
R754 B.n225 B.n206 163.367
R755 B.n225 B.n224 163.367
R756 B.n224 B.n223 163.367
R757 B.n223 B.n208 163.367
R758 B.n219 B.n208 163.367
R759 B.n219 B.n218 163.367
R760 B.n218 B.n217 163.367
R761 B.n217 B.n210 163.367
R762 B.n213 B.n210 163.367
R763 B.n213 B.n212 163.367
R764 B.n212 B.n2 163.367
R765 B.n814 B.n2 163.367
R766 B.n814 B.n813 163.367
R767 B.n813 B.n812 163.367
R768 B.n812 B.n3 163.367
R769 B.n808 B.n3 163.367
R770 B.n808 B.n807 163.367
R771 B.n807 B.n806 163.367
R772 B.n806 B.n5 163.367
R773 B.n802 B.n5 163.367
R774 B.n802 B.n801 163.367
R775 B.n801 B.n800 163.367
R776 B.n800 B.n7 163.367
R777 B.n796 B.n7 163.367
R778 B.n796 B.n795 163.367
R779 B.n795 B.n794 163.367
R780 B.n794 B.n9 163.367
R781 B.n790 B.n9 163.367
R782 B.n790 B.n789 163.367
R783 B.n789 B.n788 163.367
R784 B.n788 B.n11 163.367
R785 B.n784 B.n11 163.367
R786 B.n784 B.n783 163.367
R787 B.n783 B.n782 163.367
R788 B.n782 B.n13 163.367
R789 B.n778 B.n13 163.367
R790 B.n778 B.n777 163.367
R791 B.n777 B.n776 163.367
R792 B.n776 B.n15 163.367
R793 B.n772 B.n15 163.367
R794 B.n772 B.n771 163.367
R795 B.n771 B.n770 163.367
R796 B.n770 B.n17 163.367
R797 B.n766 B.n17 163.367
R798 B.n766 B.n765 163.367
R799 B.n765 B.n764 163.367
R800 B.n764 B.n19 163.367
R801 B.n760 B.n19 163.367
R802 B.n760 B.n759 163.367
R803 B.n759 B.n758 163.367
R804 B.n758 B.n21 163.367
R805 B.n754 B.n21 163.367
R806 B.n754 B.n753 163.367
R807 B.n753 B.n752 163.367
R808 B.n752 B.n23 163.367
R809 B.n748 B.n23 163.367
R810 B.n748 B.n747 163.367
R811 B.n747 B.n746 163.367
R812 B.n746 B.n25 163.367
R813 B.n742 B.n25 163.367
R814 B.n742 B.n741 163.367
R815 B.n741 B.n740 163.367
R816 B.n740 B.n27 163.367
R817 B.n289 B.n186 163.367
R818 B.n290 B.n289 163.367
R819 B.n291 B.n290 163.367
R820 B.n291 B.n184 163.367
R821 B.n295 B.n184 163.367
R822 B.n296 B.n295 163.367
R823 B.n297 B.n296 163.367
R824 B.n297 B.n182 163.367
R825 B.n301 B.n182 163.367
R826 B.n302 B.n301 163.367
R827 B.n303 B.n302 163.367
R828 B.n303 B.n180 163.367
R829 B.n307 B.n180 163.367
R830 B.n308 B.n307 163.367
R831 B.n309 B.n308 163.367
R832 B.n309 B.n178 163.367
R833 B.n313 B.n178 163.367
R834 B.n314 B.n313 163.367
R835 B.n315 B.n314 163.367
R836 B.n315 B.n176 163.367
R837 B.n319 B.n176 163.367
R838 B.n320 B.n319 163.367
R839 B.n321 B.n320 163.367
R840 B.n321 B.n174 163.367
R841 B.n325 B.n174 163.367
R842 B.n326 B.n325 163.367
R843 B.n327 B.n326 163.367
R844 B.n327 B.n172 163.367
R845 B.n331 B.n172 163.367
R846 B.n332 B.n331 163.367
R847 B.n333 B.n332 163.367
R848 B.n333 B.n170 163.367
R849 B.n337 B.n170 163.367
R850 B.n338 B.n337 163.367
R851 B.n339 B.n338 163.367
R852 B.n339 B.n168 163.367
R853 B.n343 B.n168 163.367
R854 B.n344 B.n343 163.367
R855 B.n345 B.n344 163.367
R856 B.n345 B.n166 163.367
R857 B.n349 B.n166 163.367
R858 B.n350 B.n349 163.367
R859 B.n351 B.n350 163.367
R860 B.n351 B.n162 163.367
R861 B.n356 B.n162 163.367
R862 B.n357 B.n356 163.367
R863 B.n358 B.n357 163.367
R864 B.n358 B.n160 163.367
R865 B.n362 B.n160 163.367
R866 B.n363 B.n362 163.367
R867 B.n364 B.n363 163.367
R868 B.n364 B.n158 163.367
R869 B.n368 B.n158 163.367
R870 B.n369 B.n368 163.367
R871 B.n369 B.n154 163.367
R872 B.n373 B.n154 163.367
R873 B.n374 B.n373 163.367
R874 B.n375 B.n374 163.367
R875 B.n375 B.n152 163.367
R876 B.n379 B.n152 163.367
R877 B.n380 B.n379 163.367
R878 B.n381 B.n380 163.367
R879 B.n381 B.n150 163.367
R880 B.n385 B.n150 163.367
R881 B.n386 B.n385 163.367
R882 B.n387 B.n386 163.367
R883 B.n387 B.n148 163.367
R884 B.n391 B.n148 163.367
R885 B.n392 B.n391 163.367
R886 B.n393 B.n392 163.367
R887 B.n393 B.n146 163.367
R888 B.n397 B.n146 163.367
R889 B.n398 B.n397 163.367
R890 B.n399 B.n398 163.367
R891 B.n399 B.n144 163.367
R892 B.n403 B.n144 163.367
R893 B.n404 B.n403 163.367
R894 B.n405 B.n404 163.367
R895 B.n405 B.n142 163.367
R896 B.n409 B.n142 163.367
R897 B.n410 B.n409 163.367
R898 B.n411 B.n410 163.367
R899 B.n411 B.n140 163.367
R900 B.n415 B.n140 163.367
R901 B.n416 B.n415 163.367
R902 B.n417 B.n416 163.367
R903 B.n417 B.n138 163.367
R904 B.n421 B.n138 163.367
R905 B.n422 B.n421 163.367
R906 B.n423 B.n422 163.367
R907 B.n423 B.n136 163.367
R908 B.n427 B.n136 163.367
R909 B.n428 B.n427 163.367
R910 B.n429 B.n428 163.367
R911 B.n429 B.n134 163.367
R912 B.n433 B.n134 163.367
R913 B.n434 B.n433 163.367
R914 B.n435 B.n132 163.367
R915 B.n439 B.n132 163.367
R916 B.n440 B.n439 163.367
R917 B.n441 B.n440 163.367
R918 B.n441 B.n130 163.367
R919 B.n445 B.n130 163.367
R920 B.n446 B.n445 163.367
R921 B.n447 B.n446 163.367
R922 B.n447 B.n128 163.367
R923 B.n451 B.n128 163.367
R924 B.n452 B.n451 163.367
R925 B.n453 B.n452 163.367
R926 B.n453 B.n126 163.367
R927 B.n457 B.n126 163.367
R928 B.n458 B.n457 163.367
R929 B.n459 B.n458 163.367
R930 B.n459 B.n124 163.367
R931 B.n463 B.n124 163.367
R932 B.n464 B.n463 163.367
R933 B.n465 B.n464 163.367
R934 B.n465 B.n122 163.367
R935 B.n469 B.n122 163.367
R936 B.n470 B.n469 163.367
R937 B.n471 B.n470 163.367
R938 B.n471 B.n120 163.367
R939 B.n475 B.n120 163.367
R940 B.n476 B.n475 163.367
R941 B.n477 B.n476 163.367
R942 B.n477 B.n118 163.367
R943 B.n481 B.n118 163.367
R944 B.n482 B.n481 163.367
R945 B.n483 B.n482 163.367
R946 B.n483 B.n116 163.367
R947 B.n487 B.n116 163.367
R948 B.n488 B.n487 163.367
R949 B.n489 B.n488 163.367
R950 B.n489 B.n114 163.367
R951 B.n493 B.n114 163.367
R952 B.n494 B.n493 163.367
R953 B.n495 B.n494 163.367
R954 B.n495 B.n112 163.367
R955 B.n499 B.n112 163.367
R956 B.n500 B.n499 163.367
R957 B.n501 B.n500 163.367
R958 B.n501 B.n110 163.367
R959 B.n505 B.n110 163.367
R960 B.n506 B.n505 163.367
R961 B.n507 B.n506 163.367
R962 B.n507 B.n108 163.367
R963 B.n511 B.n108 163.367
R964 B.n512 B.n511 163.367
R965 B.n513 B.n512 163.367
R966 B.n513 B.n106 163.367
R967 B.n517 B.n106 163.367
R968 B.n518 B.n517 163.367
R969 B.n519 B.n518 163.367
R970 B.n519 B.n104 163.367
R971 B.n523 B.n104 163.367
R972 B.n524 B.n523 163.367
R973 B.n525 B.n524 163.367
R974 B.n525 B.n102 163.367
R975 B.n529 B.n102 163.367
R976 B.n530 B.n529 163.367
R977 B.n531 B.n530 163.367
R978 B.n531 B.n100 163.367
R979 B.n535 B.n100 163.367
R980 B.n536 B.n535 163.367
R981 B.n537 B.n536 163.367
R982 B.n537 B.n98 163.367
R983 B.n541 B.n98 163.367
R984 B.n542 B.n541 163.367
R985 B.n543 B.n542 163.367
R986 B.n543 B.n96 163.367
R987 B.n547 B.n96 163.367
R988 B.n548 B.n547 163.367
R989 B.n549 B.n548 163.367
R990 B.n549 B.n94 163.367
R991 B.n553 B.n94 163.367
R992 B.n554 B.n553 163.367
R993 B.n555 B.n554 163.367
R994 B.n555 B.n92 163.367
R995 B.n559 B.n92 163.367
R996 B.n560 B.n559 163.367
R997 B.n561 B.n560 163.367
R998 B.n561 B.n90 163.367
R999 B.n565 B.n90 163.367
R1000 B.n566 B.n565 163.367
R1001 B.n567 B.n566 163.367
R1002 B.n567 B.n88 163.367
R1003 B.n571 B.n88 163.367
R1004 B.n572 B.n571 163.367
R1005 B.n573 B.n572 163.367
R1006 B.n573 B.n86 163.367
R1007 B.n577 B.n86 163.367
R1008 B.n578 B.n577 163.367
R1009 B.n579 B.n578 163.367
R1010 B.n579 B.n84 163.367
R1011 B.n583 B.n84 163.367
R1012 B.n584 B.n583 163.367
R1013 B.n585 B.n584 163.367
R1014 B.n585 B.n82 163.367
R1015 B.n589 B.n82 163.367
R1016 B.n736 B.n735 163.367
R1017 B.n735 B.n734 163.367
R1018 B.n734 B.n29 163.367
R1019 B.n730 B.n29 163.367
R1020 B.n730 B.n729 163.367
R1021 B.n729 B.n728 163.367
R1022 B.n728 B.n31 163.367
R1023 B.n724 B.n31 163.367
R1024 B.n724 B.n723 163.367
R1025 B.n723 B.n722 163.367
R1026 B.n722 B.n33 163.367
R1027 B.n718 B.n33 163.367
R1028 B.n718 B.n717 163.367
R1029 B.n717 B.n716 163.367
R1030 B.n716 B.n35 163.367
R1031 B.n712 B.n35 163.367
R1032 B.n712 B.n711 163.367
R1033 B.n711 B.n710 163.367
R1034 B.n710 B.n37 163.367
R1035 B.n706 B.n37 163.367
R1036 B.n706 B.n705 163.367
R1037 B.n705 B.n704 163.367
R1038 B.n704 B.n39 163.367
R1039 B.n700 B.n39 163.367
R1040 B.n700 B.n699 163.367
R1041 B.n699 B.n698 163.367
R1042 B.n698 B.n41 163.367
R1043 B.n694 B.n41 163.367
R1044 B.n694 B.n693 163.367
R1045 B.n693 B.n692 163.367
R1046 B.n692 B.n43 163.367
R1047 B.n688 B.n43 163.367
R1048 B.n688 B.n687 163.367
R1049 B.n687 B.n686 163.367
R1050 B.n686 B.n45 163.367
R1051 B.n682 B.n45 163.367
R1052 B.n682 B.n681 163.367
R1053 B.n681 B.n680 163.367
R1054 B.n680 B.n47 163.367
R1055 B.n676 B.n47 163.367
R1056 B.n676 B.n675 163.367
R1057 B.n675 B.n674 163.367
R1058 B.n674 B.n49 163.367
R1059 B.n669 B.n49 163.367
R1060 B.n669 B.n668 163.367
R1061 B.n668 B.n667 163.367
R1062 B.n667 B.n53 163.367
R1063 B.n663 B.n53 163.367
R1064 B.n663 B.n662 163.367
R1065 B.n662 B.n661 163.367
R1066 B.n661 B.n55 163.367
R1067 B.n657 B.n55 163.367
R1068 B.n657 B.n656 163.367
R1069 B.n656 B.n655 163.367
R1070 B.n655 B.n57 163.367
R1071 B.n651 B.n57 163.367
R1072 B.n651 B.n650 163.367
R1073 B.n650 B.n649 163.367
R1074 B.n649 B.n62 163.367
R1075 B.n645 B.n62 163.367
R1076 B.n645 B.n644 163.367
R1077 B.n644 B.n643 163.367
R1078 B.n643 B.n64 163.367
R1079 B.n639 B.n64 163.367
R1080 B.n639 B.n638 163.367
R1081 B.n638 B.n637 163.367
R1082 B.n637 B.n66 163.367
R1083 B.n633 B.n66 163.367
R1084 B.n633 B.n632 163.367
R1085 B.n632 B.n631 163.367
R1086 B.n631 B.n68 163.367
R1087 B.n627 B.n68 163.367
R1088 B.n627 B.n626 163.367
R1089 B.n626 B.n625 163.367
R1090 B.n625 B.n70 163.367
R1091 B.n621 B.n70 163.367
R1092 B.n621 B.n620 163.367
R1093 B.n620 B.n619 163.367
R1094 B.n619 B.n72 163.367
R1095 B.n615 B.n72 163.367
R1096 B.n615 B.n614 163.367
R1097 B.n614 B.n613 163.367
R1098 B.n613 B.n74 163.367
R1099 B.n609 B.n74 163.367
R1100 B.n609 B.n608 163.367
R1101 B.n608 B.n607 163.367
R1102 B.n607 B.n76 163.367
R1103 B.n603 B.n76 163.367
R1104 B.n603 B.n602 163.367
R1105 B.n602 B.n601 163.367
R1106 B.n601 B.n78 163.367
R1107 B.n597 B.n78 163.367
R1108 B.n597 B.n596 163.367
R1109 B.n596 B.n595 163.367
R1110 B.n595 B.n80 163.367
R1111 B.n591 B.n80 163.367
R1112 B.n591 B.n590 163.367
R1113 B.n155 B.t8 154.423
R1114 B.n58 B.t10 154.423
R1115 B.n163 B.t5 154.406
R1116 B.n50 B.t1 154.406
R1117 B.n156 B.t7 107.102
R1118 B.n59 B.t11 107.102
R1119 B.n164 B.t4 107.085
R1120 B.n51 B.t2 107.085
R1121 B.n157 B.n156 59.5399
R1122 B.n353 B.n164 59.5399
R1123 B.n671 B.n51 59.5399
R1124 B.n60 B.n59 59.5399
R1125 B.n156 B.n155 47.3217
R1126 B.n164 B.n163 47.3217
R1127 B.n51 B.n50 47.3217
R1128 B.n59 B.n58 47.3217
R1129 B.n738 B.n737 35.7468
R1130 B.n588 B.n81 35.7468
R1131 B.n436 B.n133 35.7468
R1132 B.n287 B.n286 35.7468
R1133 B B.n815 18.0485
R1134 B.n737 B.n28 10.6151
R1135 B.n733 B.n28 10.6151
R1136 B.n733 B.n732 10.6151
R1137 B.n732 B.n731 10.6151
R1138 B.n731 B.n30 10.6151
R1139 B.n727 B.n30 10.6151
R1140 B.n727 B.n726 10.6151
R1141 B.n726 B.n725 10.6151
R1142 B.n725 B.n32 10.6151
R1143 B.n721 B.n32 10.6151
R1144 B.n721 B.n720 10.6151
R1145 B.n720 B.n719 10.6151
R1146 B.n719 B.n34 10.6151
R1147 B.n715 B.n34 10.6151
R1148 B.n715 B.n714 10.6151
R1149 B.n714 B.n713 10.6151
R1150 B.n713 B.n36 10.6151
R1151 B.n709 B.n36 10.6151
R1152 B.n709 B.n708 10.6151
R1153 B.n708 B.n707 10.6151
R1154 B.n707 B.n38 10.6151
R1155 B.n703 B.n38 10.6151
R1156 B.n703 B.n702 10.6151
R1157 B.n702 B.n701 10.6151
R1158 B.n701 B.n40 10.6151
R1159 B.n697 B.n40 10.6151
R1160 B.n697 B.n696 10.6151
R1161 B.n696 B.n695 10.6151
R1162 B.n695 B.n42 10.6151
R1163 B.n691 B.n42 10.6151
R1164 B.n691 B.n690 10.6151
R1165 B.n690 B.n689 10.6151
R1166 B.n689 B.n44 10.6151
R1167 B.n685 B.n44 10.6151
R1168 B.n685 B.n684 10.6151
R1169 B.n684 B.n683 10.6151
R1170 B.n683 B.n46 10.6151
R1171 B.n679 B.n46 10.6151
R1172 B.n679 B.n678 10.6151
R1173 B.n678 B.n677 10.6151
R1174 B.n677 B.n48 10.6151
R1175 B.n673 B.n48 10.6151
R1176 B.n673 B.n672 10.6151
R1177 B.n670 B.n52 10.6151
R1178 B.n666 B.n52 10.6151
R1179 B.n666 B.n665 10.6151
R1180 B.n665 B.n664 10.6151
R1181 B.n664 B.n54 10.6151
R1182 B.n660 B.n54 10.6151
R1183 B.n660 B.n659 10.6151
R1184 B.n659 B.n658 10.6151
R1185 B.n658 B.n56 10.6151
R1186 B.n654 B.n653 10.6151
R1187 B.n653 B.n652 10.6151
R1188 B.n652 B.n61 10.6151
R1189 B.n648 B.n61 10.6151
R1190 B.n648 B.n647 10.6151
R1191 B.n647 B.n646 10.6151
R1192 B.n646 B.n63 10.6151
R1193 B.n642 B.n63 10.6151
R1194 B.n642 B.n641 10.6151
R1195 B.n641 B.n640 10.6151
R1196 B.n640 B.n65 10.6151
R1197 B.n636 B.n65 10.6151
R1198 B.n636 B.n635 10.6151
R1199 B.n635 B.n634 10.6151
R1200 B.n634 B.n67 10.6151
R1201 B.n630 B.n67 10.6151
R1202 B.n630 B.n629 10.6151
R1203 B.n629 B.n628 10.6151
R1204 B.n628 B.n69 10.6151
R1205 B.n624 B.n69 10.6151
R1206 B.n624 B.n623 10.6151
R1207 B.n623 B.n622 10.6151
R1208 B.n622 B.n71 10.6151
R1209 B.n618 B.n71 10.6151
R1210 B.n618 B.n617 10.6151
R1211 B.n617 B.n616 10.6151
R1212 B.n616 B.n73 10.6151
R1213 B.n612 B.n73 10.6151
R1214 B.n612 B.n611 10.6151
R1215 B.n611 B.n610 10.6151
R1216 B.n610 B.n75 10.6151
R1217 B.n606 B.n75 10.6151
R1218 B.n606 B.n605 10.6151
R1219 B.n605 B.n604 10.6151
R1220 B.n604 B.n77 10.6151
R1221 B.n600 B.n77 10.6151
R1222 B.n600 B.n599 10.6151
R1223 B.n599 B.n598 10.6151
R1224 B.n598 B.n79 10.6151
R1225 B.n594 B.n79 10.6151
R1226 B.n594 B.n593 10.6151
R1227 B.n593 B.n592 10.6151
R1228 B.n592 B.n81 10.6151
R1229 B.n437 B.n436 10.6151
R1230 B.n438 B.n437 10.6151
R1231 B.n438 B.n131 10.6151
R1232 B.n442 B.n131 10.6151
R1233 B.n443 B.n442 10.6151
R1234 B.n444 B.n443 10.6151
R1235 B.n444 B.n129 10.6151
R1236 B.n448 B.n129 10.6151
R1237 B.n449 B.n448 10.6151
R1238 B.n450 B.n449 10.6151
R1239 B.n450 B.n127 10.6151
R1240 B.n454 B.n127 10.6151
R1241 B.n455 B.n454 10.6151
R1242 B.n456 B.n455 10.6151
R1243 B.n456 B.n125 10.6151
R1244 B.n460 B.n125 10.6151
R1245 B.n461 B.n460 10.6151
R1246 B.n462 B.n461 10.6151
R1247 B.n462 B.n123 10.6151
R1248 B.n466 B.n123 10.6151
R1249 B.n467 B.n466 10.6151
R1250 B.n468 B.n467 10.6151
R1251 B.n468 B.n121 10.6151
R1252 B.n472 B.n121 10.6151
R1253 B.n473 B.n472 10.6151
R1254 B.n474 B.n473 10.6151
R1255 B.n474 B.n119 10.6151
R1256 B.n478 B.n119 10.6151
R1257 B.n479 B.n478 10.6151
R1258 B.n480 B.n479 10.6151
R1259 B.n480 B.n117 10.6151
R1260 B.n484 B.n117 10.6151
R1261 B.n485 B.n484 10.6151
R1262 B.n486 B.n485 10.6151
R1263 B.n486 B.n115 10.6151
R1264 B.n490 B.n115 10.6151
R1265 B.n491 B.n490 10.6151
R1266 B.n492 B.n491 10.6151
R1267 B.n492 B.n113 10.6151
R1268 B.n496 B.n113 10.6151
R1269 B.n497 B.n496 10.6151
R1270 B.n498 B.n497 10.6151
R1271 B.n498 B.n111 10.6151
R1272 B.n502 B.n111 10.6151
R1273 B.n503 B.n502 10.6151
R1274 B.n504 B.n503 10.6151
R1275 B.n504 B.n109 10.6151
R1276 B.n508 B.n109 10.6151
R1277 B.n509 B.n508 10.6151
R1278 B.n510 B.n509 10.6151
R1279 B.n510 B.n107 10.6151
R1280 B.n514 B.n107 10.6151
R1281 B.n515 B.n514 10.6151
R1282 B.n516 B.n515 10.6151
R1283 B.n516 B.n105 10.6151
R1284 B.n520 B.n105 10.6151
R1285 B.n521 B.n520 10.6151
R1286 B.n522 B.n521 10.6151
R1287 B.n522 B.n103 10.6151
R1288 B.n526 B.n103 10.6151
R1289 B.n527 B.n526 10.6151
R1290 B.n528 B.n527 10.6151
R1291 B.n528 B.n101 10.6151
R1292 B.n532 B.n101 10.6151
R1293 B.n533 B.n532 10.6151
R1294 B.n534 B.n533 10.6151
R1295 B.n534 B.n99 10.6151
R1296 B.n538 B.n99 10.6151
R1297 B.n539 B.n538 10.6151
R1298 B.n540 B.n539 10.6151
R1299 B.n540 B.n97 10.6151
R1300 B.n544 B.n97 10.6151
R1301 B.n545 B.n544 10.6151
R1302 B.n546 B.n545 10.6151
R1303 B.n546 B.n95 10.6151
R1304 B.n550 B.n95 10.6151
R1305 B.n551 B.n550 10.6151
R1306 B.n552 B.n551 10.6151
R1307 B.n552 B.n93 10.6151
R1308 B.n556 B.n93 10.6151
R1309 B.n557 B.n556 10.6151
R1310 B.n558 B.n557 10.6151
R1311 B.n558 B.n91 10.6151
R1312 B.n562 B.n91 10.6151
R1313 B.n563 B.n562 10.6151
R1314 B.n564 B.n563 10.6151
R1315 B.n564 B.n89 10.6151
R1316 B.n568 B.n89 10.6151
R1317 B.n569 B.n568 10.6151
R1318 B.n570 B.n569 10.6151
R1319 B.n570 B.n87 10.6151
R1320 B.n574 B.n87 10.6151
R1321 B.n575 B.n574 10.6151
R1322 B.n576 B.n575 10.6151
R1323 B.n576 B.n85 10.6151
R1324 B.n580 B.n85 10.6151
R1325 B.n581 B.n580 10.6151
R1326 B.n582 B.n581 10.6151
R1327 B.n582 B.n83 10.6151
R1328 B.n586 B.n83 10.6151
R1329 B.n587 B.n586 10.6151
R1330 B.n588 B.n587 10.6151
R1331 B.n288 B.n287 10.6151
R1332 B.n288 B.n185 10.6151
R1333 B.n292 B.n185 10.6151
R1334 B.n293 B.n292 10.6151
R1335 B.n294 B.n293 10.6151
R1336 B.n294 B.n183 10.6151
R1337 B.n298 B.n183 10.6151
R1338 B.n299 B.n298 10.6151
R1339 B.n300 B.n299 10.6151
R1340 B.n300 B.n181 10.6151
R1341 B.n304 B.n181 10.6151
R1342 B.n305 B.n304 10.6151
R1343 B.n306 B.n305 10.6151
R1344 B.n306 B.n179 10.6151
R1345 B.n310 B.n179 10.6151
R1346 B.n311 B.n310 10.6151
R1347 B.n312 B.n311 10.6151
R1348 B.n312 B.n177 10.6151
R1349 B.n316 B.n177 10.6151
R1350 B.n317 B.n316 10.6151
R1351 B.n318 B.n317 10.6151
R1352 B.n318 B.n175 10.6151
R1353 B.n322 B.n175 10.6151
R1354 B.n323 B.n322 10.6151
R1355 B.n324 B.n323 10.6151
R1356 B.n324 B.n173 10.6151
R1357 B.n328 B.n173 10.6151
R1358 B.n329 B.n328 10.6151
R1359 B.n330 B.n329 10.6151
R1360 B.n330 B.n171 10.6151
R1361 B.n334 B.n171 10.6151
R1362 B.n335 B.n334 10.6151
R1363 B.n336 B.n335 10.6151
R1364 B.n336 B.n169 10.6151
R1365 B.n340 B.n169 10.6151
R1366 B.n341 B.n340 10.6151
R1367 B.n342 B.n341 10.6151
R1368 B.n342 B.n167 10.6151
R1369 B.n346 B.n167 10.6151
R1370 B.n347 B.n346 10.6151
R1371 B.n348 B.n347 10.6151
R1372 B.n348 B.n165 10.6151
R1373 B.n352 B.n165 10.6151
R1374 B.n355 B.n354 10.6151
R1375 B.n355 B.n161 10.6151
R1376 B.n359 B.n161 10.6151
R1377 B.n360 B.n359 10.6151
R1378 B.n361 B.n360 10.6151
R1379 B.n361 B.n159 10.6151
R1380 B.n365 B.n159 10.6151
R1381 B.n366 B.n365 10.6151
R1382 B.n367 B.n366 10.6151
R1383 B.n371 B.n370 10.6151
R1384 B.n372 B.n371 10.6151
R1385 B.n372 B.n153 10.6151
R1386 B.n376 B.n153 10.6151
R1387 B.n377 B.n376 10.6151
R1388 B.n378 B.n377 10.6151
R1389 B.n378 B.n151 10.6151
R1390 B.n382 B.n151 10.6151
R1391 B.n383 B.n382 10.6151
R1392 B.n384 B.n383 10.6151
R1393 B.n384 B.n149 10.6151
R1394 B.n388 B.n149 10.6151
R1395 B.n389 B.n388 10.6151
R1396 B.n390 B.n389 10.6151
R1397 B.n390 B.n147 10.6151
R1398 B.n394 B.n147 10.6151
R1399 B.n395 B.n394 10.6151
R1400 B.n396 B.n395 10.6151
R1401 B.n396 B.n145 10.6151
R1402 B.n400 B.n145 10.6151
R1403 B.n401 B.n400 10.6151
R1404 B.n402 B.n401 10.6151
R1405 B.n402 B.n143 10.6151
R1406 B.n406 B.n143 10.6151
R1407 B.n407 B.n406 10.6151
R1408 B.n408 B.n407 10.6151
R1409 B.n408 B.n141 10.6151
R1410 B.n412 B.n141 10.6151
R1411 B.n413 B.n412 10.6151
R1412 B.n414 B.n413 10.6151
R1413 B.n414 B.n139 10.6151
R1414 B.n418 B.n139 10.6151
R1415 B.n419 B.n418 10.6151
R1416 B.n420 B.n419 10.6151
R1417 B.n420 B.n137 10.6151
R1418 B.n424 B.n137 10.6151
R1419 B.n425 B.n424 10.6151
R1420 B.n426 B.n425 10.6151
R1421 B.n426 B.n135 10.6151
R1422 B.n430 B.n135 10.6151
R1423 B.n431 B.n430 10.6151
R1424 B.n432 B.n431 10.6151
R1425 B.n432 B.n133 10.6151
R1426 B.n286 B.n187 10.6151
R1427 B.n282 B.n187 10.6151
R1428 B.n282 B.n281 10.6151
R1429 B.n281 B.n280 10.6151
R1430 B.n280 B.n189 10.6151
R1431 B.n276 B.n189 10.6151
R1432 B.n276 B.n275 10.6151
R1433 B.n275 B.n274 10.6151
R1434 B.n274 B.n191 10.6151
R1435 B.n270 B.n191 10.6151
R1436 B.n270 B.n269 10.6151
R1437 B.n269 B.n268 10.6151
R1438 B.n268 B.n193 10.6151
R1439 B.n264 B.n193 10.6151
R1440 B.n264 B.n263 10.6151
R1441 B.n263 B.n262 10.6151
R1442 B.n262 B.n195 10.6151
R1443 B.n258 B.n195 10.6151
R1444 B.n258 B.n257 10.6151
R1445 B.n257 B.n256 10.6151
R1446 B.n256 B.n197 10.6151
R1447 B.n252 B.n197 10.6151
R1448 B.n252 B.n251 10.6151
R1449 B.n251 B.n250 10.6151
R1450 B.n250 B.n199 10.6151
R1451 B.n246 B.n199 10.6151
R1452 B.n246 B.n245 10.6151
R1453 B.n245 B.n244 10.6151
R1454 B.n244 B.n201 10.6151
R1455 B.n240 B.n201 10.6151
R1456 B.n240 B.n239 10.6151
R1457 B.n239 B.n238 10.6151
R1458 B.n238 B.n203 10.6151
R1459 B.n234 B.n203 10.6151
R1460 B.n234 B.n233 10.6151
R1461 B.n233 B.n232 10.6151
R1462 B.n232 B.n205 10.6151
R1463 B.n228 B.n205 10.6151
R1464 B.n228 B.n227 10.6151
R1465 B.n227 B.n226 10.6151
R1466 B.n226 B.n207 10.6151
R1467 B.n222 B.n207 10.6151
R1468 B.n222 B.n221 10.6151
R1469 B.n221 B.n220 10.6151
R1470 B.n220 B.n209 10.6151
R1471 B.n216 B.n209 10.6151
R1472 B.n216 B.n215 10.6151
R1473 B.n215 B.n214 10.6151
R1474 B.n214 B.n211 10.6151
R1475 B.n211 B.n0 10.6151
R1476 B.n811 B.n1 10.6151
R1477 B.n811 B.n810 10.6151
R1478 B.n810 B.n809 10.6151
R1479 B.n809 B.n4 10.6151
R1480 B.n805 B.n4 10.6151
R1481 B.n805 B.n804 10.6151
R1482 B.n804 B.n803 10.6151
R1483 B.n803 B.n6 10.6151
R1484 B.n799 B.n6 10.6151
R1485 B.n799 B.n798 10.6151
R1486 B.n798 B.n797 10.6151
R1487 B.n797 B.n8 10.6151
R1488 B.n793 B.n8 10.6151
R1489 B.n793 B.n792 10.6151
R1490 B.n792 B.n791 10.6151
R1491 B.n791 B.n10 10.6151
R1492 B.n787 B.n10 10.6151
R1493 B.n787 B.n786 10.6151
R1494 B.n786 B.n785 10.6151
R1495 B.n785 B.n12 10.6151
R1496 B.n781 B.n12 10.6151
R1497 B.n781 B.n780 10.6151
R1498 B.n780 B.n779 10.6151
R1499 B.n779 B.n14 10.6151
R1500 B.n775 B.n14 10.6151
R1501 B.n775 B.n774 10.6151
R1502 B.n774 B.n773 10.6151
R1503 B.n773 B.n16 10.6151
R1504 B.n769 B.n16 10.6151
R1505 B.n769 B.n768 10.6151
R1506 B.n768 B.n767 10.6151
R1507 B.n767 B.n18 10.6151
R1508 B.n763 B.n18 10.6151
R1509 B.n763 B.n762 10.6151
R1510 B.n762 B.n761 10.6151
R1511 B.n761 B.n20 10.6151
R1512 B.n757 B.n20 10.6151
R1513 B.n757 B.n756 10.6151
R1514 B.n756 B.n755 10.6151
R1515 B.n755 B.n22 10.6151
R1516 B.n751 B.n22 10.6151
R1517 B.n751 B.n750 10.6151
R1518 B.n750 B.n749 10.6151
R1519 B.n749 B.n24 10.6151
R1520 B.n745 B.n24 10.6151
R1521 B.n745 B.n744 10.6151
R1522 B.n744 B.n743 10.6151
R1523 B.n743 B.n26 10.6151
R1524 B.n739 B.n26 10.6151
R1525 B.n739 B.n738 10.6151
R1526 B.n672 B.n671 9.36635
R1527 B.n654 B.n60 9.36635
R1528 B.n353 B.n352 9.36635
R1529 B.n370 B.n157 9.36635
R1530 B.n815 B.n0 2.81026
R1531 B.n815 B.n1 2.81026
R1532 B.n671 B.n670 1.24928
R1533 B.n60 B.n56 1.24928
R1534 B.n354 B.n353 1.24928
R1535 B.n367 B.n157 1.24928
C0 VP B 2.0178f
C1 VN w_n3898_n3554# 8.20265f
C2 VTAIL w_n3898_n3554# 3.28457f
C3 VN B 1.16966f
C4 VDD1 w_n3898_n3554# 2.67019f
C5 VTAIL B 3.7176f
C6 VN VP 7.8491f
C7 VTAIL VP 11.3475f
C8 VDD1 B 2.36019f
C9 VDD2 w_n3898_n3554# 2.78837f
C10 VDD1 VP 11.2998f
C11 VDD2 B 2.45903f
C12 VTAIL VN 11.333099f
C13 VDD2 VP 0.521316f
C14 VDD1 VN 0.152373f
C15 VDD2 VN 10.9349f
C16 VDD1 VTAIL 10.882299f
C17 VDD2 VTAIL 10.929099f
C18 VDD2 VDD1 1.85666f
C19 B w_n3898_n3554# 9.98351f
C20 VP w_n3898_n3554# 8.70864f
C21 VDD2 VSUBS 1.94234f
C22 VDD1 VSUBS 1.772333f
C23 VTAIL VSUBS 1.215547f
C24 VN VSUBS 6.91711f
C25 VP VSUBS 3.65397f
C26 B VSUBS 4.836993f
C27 w_n3898_n3554# VSUBS 0.170311p
C28 B.n0 VSUBS 0.005938f
C29 B.n1 VSUBS 0.005938f
C30 B.n2 VSUBS 0.00939f
C31 B.n3 VSUBS 0.00939f
C32 B.n4 VSUBS 0.00939f
C33 B.n5 VSUBS 0.00939f
C34 B.n6 VSUBS 0.00939f
C35 B.n7 VSUBS 0.00939f
C36 B.n8 VSUBS 0.00939f
C37 B.n9 VSUBS 0.00939f
C38 B.n10 VSUBS 0.00939f
C39 B.n11 VSUBS 0.00939f
C40 B.n12 VSUBS 0.00939f
C41 B.n13 VSUBS 0.00939f
C42 B.n14 VSUBS 0.00939f
C43 B.n15 VSUBS 0.00939f
C44 B.n16 VSUBS 0.00939f
C45 B.n17 VSUBS 0.00939f
C46 B.n18 VSUBS 0.00939f
C47 B.n19 VSUBS 0.00939f
C48 B.n20 VSUBS 0.00939f
C49 B.n21 VSUBS 0.00939f
C50 B.n22 VSUBS 0.00939f
C51 B.n23 VSUBS 0.00939f
C52 B.n24 VSUBS 0.00939f
C53 B.n25 VSUBS 0.00939f
C54 B.n26 VSUBS 0.00939f
C55 B.n27 VSUBS 0.022831f
C56 B.n28 VSUBS 0.00939f
C57 B.n29 VSUBS 0.00939f
C58 B.n30 VSUBS 0.00939f
C59 B.n31 VSUBS 0.00939f
C60 B.n32 VSUBS 0.00939f
C61 B.n33 VSUBS 0.00939f
C62 B.n34 VSUBS 0.00939f
C63 B.n35 VSUBS 0.00939f
C64 B.n36 VSUBS 0.00939f
C65 B.n37 VSUBS 0.00939f
C66 B.n38 VSUBS 0.00939f
C67 B.n39 VSUBS 0.00939f
C68 B.n40 VSUBS 0.00939f
C69 B.n41 VSUBS 0.00939f
C70 B.n42 VSUBS 0.00939f
C71 B.n43 VSUBS 0.00939f
C72 B.n44 VSUBS 0.00939f
C73 B.n45 VSUBS 0.00939f
C74 B.n46 VSUBS 0.00939f
C75 B.n47 VSUBS 0.00939f
C76 B.n48 VSUBS 0.00939f
C77 B.n49 VSUBS 0.00939f
C78 B.t2 VSUBS 0.569583f
C79 B.t1 VSUBS 0.5942f
C80 B.t0 VSUBS 1.63458f
C81 B.n50 VSUBS 0.293396f
C82 B.n51 VSUBS 0.093717f
C83 B.n52 VSUBS 0.00939f
C84 B.n53 VSUBS 0.00939f
C85 B.n54 VSUBS 0.00939f
C86 B.n55 VSUBS 0.00939f
C87 B.n56 VSUBS 0.005248f
C88 B.n57 VSUBS 0.00939f
C89 B.t11 VSUBS 0.56957f
C90 B.t10 VSUBS 0.594188f
C91 B.t9 VSUBS 1.63458f
C92 B.n58 VSUBS 0.293408f
C93 B.n59 VSUBS 0.09373f
C94 B.n60 VSUBS 0.021757f
C95 B.n61 VSUBS 0.00939f
C96 B.n62 VSUBS 0.00939f
C97 B.n63 VSUBS 0.00939f
C98 B.n64 VSUBS 0.00939f
C99 B.n65 VSUBS 0.00939f
C100 B.n66 VSUBS 0.00939f
C101 B.n67 VSUBS 0.00939f
C102 B.n68 VSUBS 0.00939f
C103 B.n69 VSUBS 0.00939f
C104 B.n70 VSUBS 0.00939f
C105 B.n71 VSUBS 0.00939f
C106 B.n72 VSUBS 0.00939f
C107 B.n73 VSUBS 0.00939f
C108 B.n74 VSUBS 0.00939f
C109 B.n75 VSUBS 0.00939f
C110 B.n76 VSUBS 0.00939f
C111 B.n77 VSUBS 0.00939f
C112 B.n78 VSUBS 0.00939f
C113 B.n79 VSUBS 0.00939f
C114 B.n80 VSUBS 0.00939f
C115 B.n81 VSUBS 0.022831f
C116 B.n82 VSUBS 0.00939f
C117 B.n83 VSUBS 0.00939f
C118 B.n84 VSUBS 0.00939f
C119 B.n85 VSUBS 0.00939f
C120 B.n86 VSUBS 0.00939f
C121 B.n87 VSUBS 0.00939f
C122 B.n88 VSUBS 0.00939f
C123 B.n89 VSUBS 0.00939f
C124 B.n90 VSUBS 0.00939f
C125 B.n91 VSUBS 0.00939f
C126 B.n92 VSUBS 0.00939f
C127 B.n93 VSUBS 0.00939f
C128 B.n94 VSUBS 0.00939f
C129 B.n95 VSUBS 0.00939f
C130 B.n96 VSUBS 0.00939f
C131 B.n97 VSUBS 0.00939f
C132 B.n98 VSUBS 0.00939f
C133 B.n99 VSUBS 0.00939f
C134 B.n100 VSUBS 0.00939f
C135 B.n101 VSUBS 0.00939f
C136 B.n102 VSUBS 0.00939f
C137 B.n103 VSUBS 0.00939f
C138 B.n104 VSUBS 0.00939f
C139 B.n105 VSUBS 0.00939f
C140 B.n106 VSUBS 0.00939f
C141 B.n107 VSUBS 0.00939f
C142 B.n108 VSUBS 0.00939f
C143 B.n109 VSUBS 0.00939f
C144 B.n110 VSUBS 0.00939f
C145 B.n111 VSUBS 0.00939f
C146 B.n112 VSUBS 0.00939f
C147 B.n113 VSUBS 0.00939f
C148 B.n114 VSUBS 0.00939f
C149 B.n115 VSUBS 0.00939f
C150 B.n116 VSUBS 0.00939f
C151 B.n117 VSUBS 0.00939f
C152 B.n118 VSUBS 0.00939f
C153 B.n119 VSUBS 0.00939f
C154 B.n120 VSUBS 0.00939f
C155 B.n121 VSUBS 0.00939f
C156 B.n122 VSUBS 0.00939f
C157 B.n123 VSUBS 0.00939f
C158 B.n124 VSUBS 0.00939f
C159 B.n125 VSUBS 0.00939f
C160 B.n126 VSUBS 0.00939f
C161 B.n127 VSUBS 0.00939f
C162 B.n128 VSUBS 0.00939f
C163 B.n129 VSUBS 0.00939f
C164 B.n130 VSUBS 0.00939f
C165 B.n131 VSUBS 0.00939f
C166 B.n132 VSUBS 0.00939f
C167 B.n133 VSUBS 0.023845f
C168 B.n134 VSUBS 0.00939f
C169 B.n135 VSUBS 0.00939f
C170 B.n136 VSUBS 0.00939f
C171 B.n137 VSUBS 0.00939f
C172 B.n138 VSUBS 0.00939f
C173 B.n139 VSUBS 0.00939f
C174 B.n140 VSUBS 0.00939f
C175 B.n141 VSUBS 0.00939f
C176 B.n142 VSUBS 0.00939f
C177 B.n143 VSUBS 0.00939f
C178 B.n144 VSUBS 0.00939f
C179 B.n145 VSUBS 0.00939f
C180 B.n146 VSUBS 0.00939f
C181 B.n147 VSUBS 0.00939f
C182 B.n148 VSUBS 0.00939f
C183 B.n149 VSUBS 0.00939f
C184 B.n150 VSUBS 0.00939f
C185 B.n151 VSUBS 0.00939f
C186 B.n152 VSUBS 0.00939f
C187 B.n153 VSUBS 0.00939f
C188 B.n154 VSUBS 0.00939f
C189 B.t7 VSUBS 0.56957f
C190 B.t8 VSUBS 0.594188f
C191 B.t6 VSUBS 1.63458f
C192 B.n155 VSUBS 0.293408f
C193 B.n156 VSUBS 0.09373f
C194 B.n157 VSUBS 0.021757f
C195 B.n158 VSUBS 0.00939f
C196 B.n159 VSUBS 0.00939f
C197 B.n160 VSUBS 0.00939f
C198 B.n161 VSUBS 0.00939f
C199 B.n162 VSUBS 0.00939f
C200 B.t4 VSUBS 0.569583f
C201 B.t5 VSUBS 0.5942f
C202 B.t3 VSUBS 1.63458f
C203 B.n163 VSUBS 0.293396f
C204 B.n164 VSUBS 0.093717f
C205 B.n165 VSUBS 0.00939f
C206 B.n166 VSUBS 0.00939f
C207 B.n167 VSUBS 0.00939f
C208 B.n168 VSUBS 0.00939f
C209 B.n169 VSUBS 0.00939f
C210 B.n170 VSUBS 0.00939f
C211 B.n171 VSUBS 0.00939f
C212 B.n172 VSUBS 0.00939f
C213 B.n173 VSUBS 0.00939f
C214 B.n174 VSUBS 0.00939f
C215 B.n175 VSUBS 0.00939f
C216 B.n176 VSUBS 0.00939f
C217 B.n177 VSUBS 0.00939f
C218 B.n178 VSUBS 0.00939f
C219 B.n179 VSUBS 0.00939f
C220 B.n180 VSUBS 0.00939f
C221 B.n181 VSUBS 0.00939f
C222 B.n182 VSUBS 0.00939f
C223 B.n183 VSUBS 0.00939f
C224 B.n184 VSUBS 0.00939f
C225 B.n185 VSUBS 0.00939f
C226 B.n186 VSUBS 0.023845f
C227 B.n187 VSUBS 0.00939f
C228 B.n188 VSUBS 0.00939f
C229 B.n189 VSUBS 0.00939f
C230 B.n190 VSUBS 0.00939f
C231 B.n191 VSUBS 0.00939f
C232 B.n192 VSUBS 0.00939f
C233 B.n193 VSUBS 0.00939f
C234 B.n194 VSUBS 0.00939f
C235 B.n195 VSUBS 0.00939f
C236 B.n196 VSUBS 0.00939f
C237 B.n197 VSUBS 0.00939f
C238 B.n198 VSUBS 0.00939f
C239 B.n199 VSUBS 0.00939f
C240 B.n200 VSUBS 0.00939f
C241 B.n201 VSUBS 0.00939f
C242 B.n202 VSUBS 0.00939f
C243 B.n203 VSUBS 0.00939f
C244 B.n204 VSUBS 0.00939f
C245 B.n205 VSUBS 0.00939f
C246 B.n206 VSUBS 0.00939f
C247 B.n207 VSUBS 0.00939f
C248 B.n208 VSUBS 0.00939f
C249 B.n209 VSUBS 0.00939f
C250 B.n210 VSUBS 0.00939f
C251 B.n211 VSUBS 0.00939f
C252 B.n212 VSUBS 0.00939f
C253 B.n213 VSUBS 0.00939f
C254 B.n214 VSUBS 0.00939f
C255 B.n215 VSUBS 0.00939f
C256 B.n216 VSUBS 0.00939f
C257 B.n217 VSUBS 0.00939f
C258 B.n218 VSUBS 0.00939f
C259 B.n219 VSUBS 0.00939f
C260 B.n220 VSUBS 0.00939f
C261 B.n221 VSUBS 0.00939f
C262 B.n222 VSUBS 0.00939f
C263 B.n223 VSUBS 0.00939f
C264 B.n224 VSUBS 0.00939f
C265 B.n225 VSUBS 0.00939f
C266 B.n226 VSUBS 0.00939f
C267 B.n227 VSUBS 0.00939f
C268 B.n228 VSUBS 0.00939f
C269 B.n229 VSUBS 0.00939f
C270 B.n230 VSUBS 0.00939f
C271 B.n231 VSUBS 0.00939f
C272 B.n232 VSUBS 0.00939f
C273 B.n233 VSUBS 0.00939f
C274 B.n234 VSUBS 0.00939f
C275 B.n235 VSUBS 0.00939f
C276 B.n236 VSUBS 0.00939f
C277 B.n237 VSUBS 0.00939f
C278 B.n238 VSUBS 0.00939f
C279 B.n239 VSUBS 0.00939f
C280 B.n240 VSUBS 0.00939f
C281 B.n241 VSUBS 0.00939f
C282 B.n242 VSUBS 0.00939f
C283 B.n243 VSUBS 0.00939f
C284 B.n244 VSUBS 0.00939f
C285 B.n245 VSUBS 0.00939f
C286 B.n246 VSUBS 0.00939f
C287 B.n247 VSUBS 0.00939f
C288 B.n248 VSUBS 0.00939f
C289 B.n249 VSUBS 0.00939f
C290 B.n250 VSUBS 0.00939f
C291 B.n251 VSUBS 0.00939f
C292 B.n252 VSUBS 0.00939f
C293 B.n253 VSUBS 0.00939f
C294 B.n254 VSUBS 0.00939f
C295 B.n255 VSUBS 0.00939f
C296 B.n256 VSUBS 0.00939f
C297 B.n257 VSUBS 0.00939f
C298 B.n258 VSUBS 0.00939f
C299 B.n259 VSUBS 0.00939f
C300 B.n260 VSUBS 0.00939f
C301 B.n261 VSUBS 0.00939f
C302 B.n262 VSUBS 0.00939f
C303 B.n263 VSUBS 0.00939f
C304 B.n264 VSUBS 0.00939f
C305 B.n265 VSUBS 0.00939f
C306 B.n266 VSUBS 0.00939f
C307 B.n267 VSUBS 0.00939f
C308 B.n268 VSUBS 0.00939f
C309 B.n269 VSUBS 0.00939f
C310 B.n270 VSUBS 0.00939f
C311 B.n271 VSUBS 0.00939f
C312 B.n272 VSUBS 0.00939f
C313 B.n273 VSUBS 0.00939f
C314 B.n274 VSUBS 0.00939f
C315 B.n275 VSUBS 0.00939f
C316 B.n276 VSUBS 0.00939f
C317 B.n277 VSUBS 0.00939f
C318 B.n278 VSUBS 0.00939f
C319 B.n279 VSUBS 0.00939f
C320 B.n280 VSUBS 0.00939f
C321 B.n281 VSUBS 0.00939f
C322 B.n282 VSUBS 0.00939f
C323 B.n283 VSUBS 0.00939f
C324 B.n284 VSUBS 0.00939f
C325 B.n285 VSUBS 0.022831f
C326 B.n286 VSUBS 0.022831f
C327 B.n287 VSUBS 0.023845f
C328 B.n288 VSUBS 0.00939f
C329 B.n289 VSUBS 0.00939f
C330 B.n290 VSUBS 0.00939f
C331 B.n291 VSUBS 0.00939f
C332 B.n292 VSUBS 0.00939f
C333 B.n293 VSUBS 0.00939f
C334 B.n294 VSUBS 0.00939f
C335 B.n295 VSUBS 0.00939f
C336 B.n296 VSUBS 0.00939f
C337 B.n297 VSUBS 0.00939f
C338 B.n298 VSUBS 0.00939f
C339 B.n299 VSUBS 0.00939f
C340 B.n300 VSUBS 0.00939f
C341 B.n301 VSUBS 0.00939f
C342 B.n302 VSUBS 0.00939f
C343 B.n303 VSUBS 0.00939f
C344 B.n304 VSUBS 0.00939f
C345 B.n305 VSUBS 0.00939f
C346 B.n306 VSUBS 0.00939f
C347 B.n307 VSUBS 0.00939f
C348 B.n308 VSUBS 0.00939f
C349 B.n309 VSUBS 0.00939f
C350 B.n310 VSUBS 0.00939f
C351 B.n311 VSUBS 0.00939f
C352 B.n312 VSUBS 0.00939f
C353 B.n313 VSUBS 0.00939f
C354 B.n314 VSUBS 0.00939f
C355 B.n315 VSUBS 0.00939f
C356 B.n316 VSUBS 0.00939f
C357 B.n317 VSUBS 0.00939f
C358 B.n318 VSUBS 0.00939f
C359 B.n319 VSUBS 0.00939f
C360 B.n320 VSUBS 0.00939f
C361 B.n321 VSUBS 0.00939f
C362 B.n322 VSUBS 0.00939f
C363 B.n323 VSUBS 0.00939f
C364 B.n324 VSUBS 0.00939f
C365 B.n325 VSUBS 0.00939f
C366 B.n326 VSUBS 0.00939f
C367 B.n327 VSUBS 0.00939f
C368 B.n328 VSUBS 0.00939f
C369 B.n329 VSUBS 0.00939f
C370 B.n330 VSUBS 0.00939f
C371 B.n331 VSUBS 0.00939f
C372 B.n332 VSUBS 0.00939f
C373 B.n333 VSUBS 0.00939f
C374 B.n334 VSUBS 0.00939f
C375 B.n335 VSUBS 0.00939f
C376 B.n336 VSUBS 0.00939f
C377 B.n337 VSUBS 0.00939f
C378 B.n338 VSUBS 0.00939f
C379 B.n339 VSUBS 0.00939f
C380 B.n340 VSUBS 0.00939f
C381 B.n341 VSUBS 0.00939f
C382 B.n342 VSUBS 0.00939f
C383 B.n343 VSUBS 0.00939f
C384 B.n344 VSUBS 0.00939f
C385 B.n345 VSUBS 0.00939f
C386 B.n346 VSUBS 0.00939f
C387 B.n347 VSUBS 0.00939f
C388 B.n348 VSUBS 0.00939f
C389 B.n349 VSUBS 0.00939f
C390 B.n350 VSUBS 0.00939f
C391 B.n351 VSUBS 0.00939f
C392 B.n352 VSUBS 0.008838f
C393 B.n353 VSUBS 0.021757f
C394 B.n354 VSUBS 0.005248f
C395 B.n355 VSUBS 0.00939f
C396 B.n356 VSUBS 0.00939f
C397 B.n357 VSUBS 0.00939f
C398 B.n358 VSUBS 0.00939f
C399 B.n359 VSUBS 0.00939f
C400 B.n360 VSUBS 0.00939f
C401 B.n361 VSUBS 0.00939f
C402 B.n362 VSUBS 0.00939f
C403 B.n363 VSUBS 0.00939f
C404 B.n364 VSUBS 0.00939f
C405 B.n365 VSUBS 0.00939f
C406 B.n366 VSUBS 0.00939f
C407 B.n367 VSUBS 0.005248f
C408 B.n368 VSUBS 0.00939f
C409 B.n369 VSUBS 0.00939f
C410 B.n370 VSUBS 0.008838f
C411 B.n371 VSUBS 0.00939f
C412 B.n372 VSUBS 0.00939f
C413 B.n373 VSUBS 0.00939f
C414 B.n374 VSUBS 0.00939f
C415 B.n375 VSUBS 0.00939f
C416 B.n376 VSUBS 0.00939f
C417 B.n377 VSUBS 0.00939f
C418 B.n378 VSUBS 0.00939f
C419 B.n379 VSUBS 0.00939f
C420 B.n380 VSUBS 0.00939f
C421 B.n381 VSUBS 0.00939f
C422 B.n382 VSUBS 0.00939f
C423 B.n383 VSUBS 0.00939f
C424 B.n384 VSUBS 0.00939f
C425 B.n385 VSUBS 0.00939f
C426 B.n386 VSUBS 0.00939f
C427 B.n387 VSUBS 0.00939f
C428 B.n388 VSUBS 0.00939f
C429 B.n389 VSUBS 0.00939f
C430 B.n390 VSUBS 0.00939f
C431 B.n391 VSUBS 0.00939f
C432 B.n392 VSUBS 0.00939f
C433 B.n393 VSUBS 0.00939f
C434 B.n394 VSUBS 0.00939f
C435 B.n395 VSUBS 0.00939f
C436 B.n396 VSUBS 0.00939f
C437 B.n397 VSUBS 0.00939f
C438 B.n398 VSUBS 0.00939f
C439 B.n399 VSUBS 0.00939f
C440 B.n400 VSUBS 0.00939f
C441 B.n401 VSUBS 0.00939f
C442 B.n402 VSUBS 0.00939f
C443 B.n403 VSUBS 0.00939f
C444 B.n404 VSUBS 0.00939f
C445 B.n405 VSUBS 0.00939f
C446 B.n406 VSUBS 0.00939f
C447 B.n407 VSUBS 0.00939f
C448 B.n408 VSUBS 0.00939f
C449 B.n409 VSUBS 0.00939f
C450 B.n410 VSUBS 0.00939f
C451 B.n411 VSUBS 0.00939f
C452 B.n412 VSUBS 0.00939f
C453 B.n413 VSUBS 0.00939f
C454 B.n414 VSUBS 0.00939f
C455 B.n415 VSUBS 0.00939f
C456 B.n416 VSUBS 0.00939f
C457 B.n417 VSUBS 0.00939f
C458 B.n418 VSUBS 0.00939f
C459 B.n419 VSUBS 0.00939f
C460 B.n420 VSUBS 0.00939f
C461 B.n421 VSUBS 0.00939f
C462 B.n422 VSUBS 0.00939f
C463 B.n423 VSUBS 0.00939f
C464 B.n424 VSUBS 0.00939f
C465 B.n425 VSUBS 0.00939f
C466 B.n426 VSUBS 0.00939f
C467 B.n427 VSUBS 0.00939f
C468 B.n428 VSUBS 0.00939f
C469 B.n429 VSUBS 0.00939f
C470 B.n430 VSUBS 0.00939f
C471 B.n431 VSUBS 0.00939f
C472 B.n432 VSUBS 0.00939f
C473 B.n433 VSUBS 0.00939f
C474 B.n434 VSUBS 0.023845f
C475 B.n435 VSUBS 0.022831f
C476 B.n436 VSUBS 0.022831f
C477 B.n437 VSUBS 0.00939f
C478 B.n438 VSUBS 0.00939f
C479 B.n439 VSUBS 0.00939f
C480 B.n440 VSUBS 0.00939f
C481 B.n441 VSUBS 0.00939f
C482 B.n442 VSUBS 0.00939f
C483 B.n443 VSUBS 0.00939f
C484 B.n444 VSUBS 0.00939f
C485 B.n445 VSUBS 0.00939f
C486 B.n446 VSUBS 0.00939f
C487 B.n447 VSUBS 0.00939f
C488 B.n448 VSUBS 0.00939f
C489 B.n449 VSUBS 0.00939f
C490 B.n450 VSUBS 0.00939f
C491 B.n451 VSUBS 0.00939f
C492 B.n452 VSUBS 0.00939f
C493 B.n453 VSUBS 0.00939f
C494 B.n454 VSUBS 0.00939f
C495 B.n455 VSUBS 0.00939f
C496 B.n456 VSUBS 0.00939f
C497 B.n457 VSUBS 0.00939f
C498 B.n458 VSUBS 0.00939f
C499 B.n459 VSUBS 0.00939f
C500 B.n460 VSUBS 0.00939f
C501 B.n461 VSUBS 0.00939f
C502 B.n462 VSUBS 0.00939f
C503 B.n463 VSUBS 0.00939f
C504 B.n464 VSUBS 0.00939f
C505 B.n465 VSUBS 0.00939f
C506 B.n466 VSUBS 0.00939f
C507 B.n467 VSUBS 0.00939f
C508 B.n468 VSUBS 0.00939f
C509 B.n469 VSUBS 0.00939f
C510 B.n470 VSUBS 0.00939f
C511 B.n471 VSUBS 0.00939f
C512 B.n472 VSUBS 0.00939f
C513 B.n473 VSUBS 0.00939f
C514 B.n474 VSUBS 0.00939f
C515 B.n475 VSUBS 0.00939f
C516 B.n476 VSUBS 0.00939f
C517 B.n477 VSUBS 0.00939f
C518 B.n478 VSUBS 0.00939f
C519 B.n479 VSUBS 0.00939f
C520 B.n480 VSUBS 0.00939f
C521 B.n481 VSUBS 0.00939f
C522 B.n482 VSUBS 0.00939f
C523 B.n483 VSUBS 0.00939f
C524 B.n484 VSUBS 0.00939f
C525 B.n485 VSUBS 0.00939f
C526 B.n486 VSUBS 0.00939f
C527 B.n487 VSUBS 0.00939f
C528 B.n488 VSUBS 0.00939f
C529 B.n489 VSUBS 0.00939f
C530 B.n490 VSUBS 0.00939f
C531 B.n491 VSUBS 0.00939f
C532 B.n492 VSUBS 0.00939f
C533 B.n493 VSUBS 0.00939f
C534 B.n494 VSUBS 0.00939f
C535 B.n495 VSUBS 0.00939f
C536 B.n496 VSUBS 0.00939f
C537 B.n497 VSUBS 0.00939f
C538 B.n498 VSUBS 0.00939f
C539 B.n499 VSUBS 0.00939f
C540 B.n500 VSUBS 0.00939f
C541 B.n501 VSUBS 0.00939f
C542 B.n502 VSUBS 0.00939f
C543 B.n503 VSUBS 0.00939f
C544 B.n504 VSUBS 0.00939f
C545 B.n505 VSUBS 0.00939f
C546 B.n506 VSUBS 0.00939f
C547 B.n507 VSUBS 0.00939f
C548 B.n508 VSUBS 0.00939f
C549 B.n509 VSUBS 0.00939f
C550 B.n510 VSUBS 0.00939f
C551 B.n511 VSUBS 0.00939f
C552 B.n512 VSUBS 0.00939f
C553 B.n513 VSUBS 0.00939f
C554 B.n514 VSUBS 0.00939f
C555 B.n515 VSUBS 0.00939f
C556 B.n516 VSUBS 0.00939f
C557 B.n517 VSUBS 0.00939f
C558 B.n518 VSUBS 0.00939f
C559 B.n519 VSUBS 0.00939f
C560 B.n520 VSUBS 0.00939f
C561 B.n521 VSUBS 0.00939f
C562 B.n522 VSUBS 0.00939f
C563 B.n523 VSUBS 0.00939f
C564 B.n524 VSUBS 0.00939f
C565 B.n525 VSUBS 0.00939f
C566 B.n526 VSUBS 0.00939f
C567 B.n527 VSUBS 0.00939f
C568 B.n528 VSUBS 0.00939f
C569 B.n529 VSUBS 0.00939f
C570 B.n530 VSUBS 0.00939f
C571 B.n531 VSUBS 0.00939f
C572 B.n532 VSUBS 0.00939f
C573 B.n533 VSUBS 0.00939f
C574 B.n534 VSUBS 0.00939f
C575 B.n535 VSUBS 0.00939f
C576 B.n536 VSUBS 0.00939f
C577 B.n537 VSUBS 0.00939f
C578 B.n538 VSUBS 0.00939f
C579 B.n539 VSUBS 0.00939f
C580 B.n540 VSUBS 0.00939f
C581 B.n541 VSUBS 0.00939f
C582 B.n542 VSUBS 0.00939f
C583 B.n543 VSUBS 0.00939f
C584 B.n544 VSUBS 0.00939f
C585 B.n545 VSUBS 0.00939f
C586 B.n546 VSUBS 0.00939f
C587 B.n547 VSUBS 0.00939f
C588 B.n548 VSUBS 0.00939f
C589 B.n549 VSUBS 0.00939f
C590 B.n550 VSUBS 0.00939f
C591 B.n551 VSUBS 0.00939f
C592 B.n552 VSUBS 0.00939f
C593 B.n553 VSUBS 0.00939f
C594 B.n554 VSUBS 0.00939f
C595 B.n555 VSUBS 0.00939f
C596 B.n556 VSUBS 0.00939f
C597 B.n557 VSUBS 0.00939f
C598 B.n558 VSUBS 0.00939f
C599 B.n559 VSUBS 0.00939f
C600 B.n560 VSUBS 0.00939f
C601 B.n561 VSUBS 0.00939f
C602 B.n562 VSUBS 0.00939f
C603 B.n563 VSUBS 0.00939f
C604 B.n564 VSUBS 0.00939f
C605 B.n565 VSUBS 0.00939f
C606 B.n566 VSUBS 0.00939f
C607 B.n567 VSUBS 0.00939f
C608 B.n568 VSUBS 0.00939f
C609 B.n569 VSUBS 0.00939f
C610 B.n570 VSUBS 0.00939f
C611 B.n571 VSUBS 0.00939f
C612 B.n572 VSUBS 0.00939f
C613 B.n573 VSUBS 0.00939f
C614 B.n574 VSUBS 0.00939f
C615 B.n575 VSUBS 0.00939f
C616 B.n576 VSUBS 0.00939f
C617 B.n577 VSUBS 0.00939f
C618 B.n578 VSUBS 0.00939f
C619 B.n579 VSUBS 0.00939f
C620 B.n580 VSUBS 0.00939f
C621 B.n581 VSUBS 0.00939f
C622 B.n582 VSUBS 0.00939f
C623 B.n583 VSUBS 0.00939f
C624 B.n584 VSUBS 0.00939f
C625 B.n585 VSUBS 0.00939f
C626 B.n586 VSUBS 0.00939f
C627 B.n587 VSUBS 0.00939f
C628 B.n588 VSUBS 0.023845f
C629 B.n589 VSUBS 0.022831f
C630 B.n590 VSUBS 0.023845f
C631 B.n591 VSUBS 0.00939f
C632 B.n592 VSUBS 0.00939f
C633 B.n593 VSUBS 0.00939f
C634 B.n594 VSUBS 0.00939f
C635 B.n595 VSUBS 0.00939f
C636 B.n596 VSUBS 0.00939f
C637 B.n597 VSUBS 0.00939f
C638 B.n598 VSUBS 0.00939f
C639 B.n599 VSUBS 0.00939f
C640 B.n600 VSUBS 0.00939f
C641 B.n601 VSUBS 0.00939f
C642 B.n602 VSUBS 0.00939f
C643 B.n603 VSUBS 0.00939f
C644 B.n604 VSUBS 0.00939f
C645 B.n605 VSUBS 0.00939f
C646 B.n606 VSUBS 0.00939f
C647 B.n607 VSUBS 0.00939f
C648 B.n608 VSUBS 0.00939f
C649 B.n609 VSUBS 0.00939f
C650 B.n610 VSUBS 0.00939f
C651 B.n611 VSUBS 0.00939f
C652 B.n612 VSUBS 0.00939f
C653 B.n613 VSUBS 0.00939f
C654 B.n614 VSUBS 0.00939f
C655 B.n615 VSUBS 0.00939f
C656 B.n616 VSUBS 0.00939f
C657 B.n617 VSUBS 0.00939f
C658 B.n618 VSUBS 0.00939f
C659 B.n619 VSUBS 0.00939f
C660 B.n620 VSUBS 0.00939f
C661 B.n621 VSUBS 0.00939f
C662 B.n622 VSUBS 0.00939f
C663 B.n623 VSUBS 0.00939f
C664 B.n624 VSUBS 0.00939f
C665 B.n625 VSUBS 0.00939f
C666 B.n626 VSUBS 0.00939f
C667 B.n627 VSUBS 0.00939f
C668 B.n628 VSUBS 0.00939f
C669 B.n629 VSUBS 0.00939f
C670 B.n630 VSUBS 0.00939f
C671 B.n631 VSUBS 0.00939f
C672 B.n632 VSUBS 0.00939f
C673 B.n633 VSUBS 0.00939f
C674 B.n634 VSUBS 0.00939f
C675 B.n635 VSUBS 0.00939f
C676 B.n636 VSUBS 0.00939f
C677 B.n637 VSUBS 0.00939f
C678 B.n638 VSUBS 0.00939f
C679 B.n639 VSUBS 0.00939f
C680 B.n640 VSUBS 0.00939f
C681 B.n641 VSUBS 0.00939f
C682 B.n642 VSUBS 0.00939f
C683 B.n643 VSUBS 0.00939f
C684 B.n644 VSUBS 0.00939f
C685 B.n645 VSUBS 0.00939f
C686 B.n646 VSUBS 0.00939f
C687 B.n647 VSUBS 0.00939f
C688 B.n648 VSUBS 0.00939f
C689 B.n649 VSUBS 0.00939f
C690 B.n650 VSUBS 0.00939f
C691 B.n651 VSUBS 0.00939f
C692 B.n652 VSUBS 0.00939f
C693 B.n653 VSUBS 0.00939f
C694 B.n654 VSUBS 0.008838f
C695 B.n655 VSUBS 0.00939f
C696 B.n656 VSUBS 0.00939f
C697 B.n657 VSUBS 0.00939f
C698 B.n658 VSUBS 0.00939f
C699 B.n659 VSUBS 0.00939f
C700 B.n660 VSUBS 0.00939f
C701 B.n661 VSUBS 0.00939f
C702 B.n662 VSUBS 0.00939f
C703 B.n663 VSUBS 0.00939f
C704 B.n664 VSUBS 0.00939f
C705 B.n665 VSUBS 0.00939f
C706 B.n666 VSUBS 0.00939f
C707 B.n667 VSUBS 0.00939f
C708 B.n668 VSUBS 0.00939f
C709 B.n669 VSUBS 0.00939f
C710 B.n670 VSUBS 0.005248f
C711 B.n671 VSUBS 0.021757f
C712 B.n672 VSUBS 0.008838f
C713 B.n673 VSUBS 0.00939f
C714 B.n674 VSUBS 0.00939f
C715 B.n675 VSUBS 0.00939f
C716 B.n676 VSUBS 0.00939f
C717 B.n677 VSUBS 0.00939f
C718 B.n678 VSUBS 0.00939f
C719 B.n679 VSUBS 0.00939f
C720 B.n680 VSUBS 0.00939f
C721 B.n681 VSUBS 0.00939f
C722 B.n682 VSUBS 0.00939f
C723 B.n683 VSUBS 0.00939f
C724 B.n684 VSUBS 0.00939f
C725 B.n685 VSUBS 0.00939f
C726 B.n686 VSUBS 0.00939f
C727 B.n687 VSUBS 0.00939f
C728 B.n688 VSUBS 0.00939f
C729 B.n689 VSUBS 0.00939f
C730 B.n690 VSUBS 0.00939f
C731 B.n691 VSUBS 0.00939f
C732 B.n692 VSUBS 0.00939f
C733 B.n693 VSUBS 0.00939f
C734 B.n694 VSUBS 0.00939f
C735 B.n695 VSUBS 0.00939f
C736 B.n696 VSUBS 0.00939f
C737 B.n697 VSUBS 0.00939f
C738 B.n698 VSUBS 0.00939f
C739 B.n699 VSUBS 0.00939f
C740 B.n700 VSUBS 0.00939f
C741 B.n701 VSUBS 0.00939f
C742 B.n702 VSUBS 0.00939f
C743 B.n703 VSUBS 0.00939f
C744 B.n704 VSUBS 0.00939f
C745 B.n705 VSUBS 0.00939f
C746 B.n706 VSUBS 0.00939f
C747 B.n707 VSUBS 0.00939f
C748 B.n708 VSUBS 0.00939f
C749 B.n709 VSUBS 0.00939f
C750 B.n710 VSUBS 0.00939f
C751 B.n711 VSUBS 0.00939f
C752 B.n712 VSUBS 0.00939f
C753 B.n713 VSUBS 0.00939f
C754 B.n714 VSUBS 0.00939f
C755 B.n715 VSUBS 0.00939f
C756 B.n716 VSUBS 0.00939f
C757 B.n717 VSUBS 0.00939f
C758 B.n718 VSUBS 0.00939f
C759 B.n719 VSUBS 0.00939f
C760 B.n720 VSUBS 0.00939f
C761 B.n721 VSUBS 0.00939f
C762 B.n722 VSUBS 0.00939f
C763 B.n723 VSUBS 0.00939f
C764 B.n724 VSUBS 0.00939f
C765 B.n725 VSUBS 0.00939f
C766 B.n726 VSUBS 0.00939f
C767 B.n727 VSUBS 0.00939f
C768 B.n728 VSUBS 0.00939f
C769 B.n729 VSUBS 0.00939f
C770 B.n730 VSUBS 0.00939f
C771 B.n731 VSUBS 0.00939f
C772 B.n732 VSUBS 0.00939f
C773 B.n733 VSUBS 0.00939f
C774 B.n734 VSUBS 0.00939f
C775 B.n735 VSUBS 0.00939f
C776 B.n736 VSUBS 0.023845f
C777 B.n737 VSUBS 0.023845f
C778 B.n738 VSUBS 0.022831f
C779 B.n739 VSUBS 0.00939f
C780 B.n740 VSUBS 0.00939f
C781 B.n741 VSUBS 0.00939f
C782 B.n742 VSUBS 0.00939f
C783 B.n743 VSUBS 0.00939f
C784 B.n744 VSUBS 0.00939f
C785 B.n745 VSUBS 0.00939f
C786 B.n746 VSUBS 0.00939f
C787 B.n747 VSUBS 0.00939f
C788 B.n748 VSUBS 0.00939f
C789 B.n749 VSUBS 0.00939f
C790 B.n750 VSUBS 0.00939f
C791 B.n751 VSUBS 0.00939f
C792 B.n752 VSUBS 0.00939f
C793 B.n753 VSUBS 0.00939f
C794 B.n754 VSUBS 0.00939f
C795 B.n755 VSUBS 0.00939f
C796 B.n756 VSUBS 0.00939f
C797 B.n757 VSUBS 0.00939f
C798 B.n758 VSUBS 0.00939f
C799 B.n759 VSUBS 0.00939f
C800 B.n760 VSUBS 0.00939f
C801 B.n761 VSUBS 0.00939f
C802 B.n762 VSUBS 0.00939f
C803 B.n763 VSUBS 0.00939f
C804 B.n764 VSUBS 0.00939f
C805 B.n765 VSUBS 0.00939f
C806 B.n766 VSUBS 0.00939f
C807 B.n767 VSUBS 0.00939f
C808 B.n768 VSUBS 0.00939f
C809 B.n769 VSUBS 0.00939f
C810 B.n770 VSUBS 0.00939f
C811 B.n771 VSUBS 0.00939f
C812 B.n772 VSUBS 0.00939f
C813 B.n773 VSUBS 0.00939f
C814 B.n774 VSUBS 0.00939f
C815 B.n775 VSUBS 0.00939f
C816 B.n776 VSUBS 0.00939f
C817 B.n777 VSUBS 0.00939f
C818 B.n778 VSUBS 0.00939f
C819 B.n779 VSUBS 0.00939f
C820 B.n780 VSUBS 0.00939f
C821 B.n781 VSUBS 0.00939f
C822 B.n782 VSUBS 0.00939f
C823 B.n783 VSUBS 0.00939f
C824 B.n784 VSUBS 0.00939f
C825 B.n785 VSUBS 0.00939f
C826 B.n786 VSUBS 0.00939f
C827 B.n787 VSUBS 0.00939f
C828 B.n788 VSUBS 0.00939f
C829 B.n789 VSUBS 0.00939f
C830 B.n790 VSUBS 0.00939f
C831 B.n791 VSUBS 0.00939f
C832 B.n792 VSUBS 0.00939f
C833 B.n793 VSUBS 0.00939f
C834 B.n794 VSUBS 0.00939f
C835 B.n795 VSUBS 0.00939f
C836 B.n796 VSUBS 0.00939f
C837 B.n797 VSUBS 0.00939f
C838 B.n798 VSUBS 0.00939f
C839 B.n799 VSUBS 0.00939f
C840 B.n800 VSUBS 0.00939f
C841 B.n801 VSUBS 0.00939f
C842 B.n802 VSUBS 0.00939f
C843 B.n803 VSUBS 0.00939f
C844 B.n804 VSUBS 0.00939f
C845 B.n805 VSUBS 0.00939f
C846 B.n806 VSUBS 0.00939f
C847 B.n807 VSUBS 0.00939f
C848 B.n808 VSUBS 0.00939f
C849 B.n809 VSUBS 0.00939f
C850 B.n810 VSUBS 0.00939f
C851 B.n811 VSUBS 0.00939f
C852 B.n812 VSUBS 0.00939f
C853 B.n813 VSUBS 0.00939f
C854 B.n814 VSUBS 0.00939f
C855 B.n815 VSUBS 0.021263f
C856 VDD2.t0 VSUBS 2.92526f
C857 VDD2.t8 VSUBS 0.279991f
C858 VDD2.t1 VSUBS 0.279991f
C859 VDD2.n0 VSUBS 2.2296f
C860 VDD2.n1 VSUBS 1.5019f
C861 VDD2.t9 VSUBS 0.279991f
C862 VDD2.t5 VSUBS 0.279991f
C863 VDD2.n2 VSUBS 2.24644f
C864 VDD2.n3 VSUBS 3.24157f
C865 VDD2.t4 VSUBS 2.90415f
C866 VDD2.n4 VSUBS 3.58943f
C867 VDD2.t3 VSUBS 0.279991f
C868 VDD2.t7 VSUBS 0.279991f
C869 VDD2.n5 VSUBS 2.22962f
C870 VDD2.n6 VSUBS 0.741565f
C871 VDD2.t2 VSUBS 0.279991f
C872 VDD2.t6 VSUBS 0.279991f
C873 VDD2.n7 VSUBS 2.24639f
C874 VN.n0 VSUBS 0.040607f
C875 VN.t4 VSUBS 2.29422f
C876 VN.n1 VSUBS 0.036775f
C877 VN.n2 VSUBS 0.0308f
C878 VN.t0 VSUBS 2.29422f
C879 VN.n3 VSUBS 0.047538f
C880 VN.n4 VSUBS 0.0308f
C881 VN.t8 VSUBS 2.29422f
C882 VN.n5 VSUBS 0.057404f
C883 VN.n6 VSUBS 0.0308f
C884 VN.t1 VSUBS 2.29422f
C885 VN.n7 VSUBS 0.90156f
C886 VN.t9 VSUBS 2.47695f
C887 VN.n8 VSUBS 0.880809f
C888 VN.n9 VSUBS 0.259615f
C889 VN.n10 VSUBS 0.054003f
C890 VN.n11 VSUBS 0.047538f
C891 VN.n12 VSUBS 0.042388f
C892 VN.n13 VSUBS 0.0308f
C893 VN.n14 VSUBS 0.0308f
C894 VN.n15 VSUBS 0.0308f
C895 VN.n16 VSUBS 0.842382f
C896 VN.n17 VSUBS 0.057404f
C897 VN.n18 VSUBS 0.042388f
C898 VN.n19 VSUBS 0.0308f
C899 VN.n20 VSUBS 0.0308f
C900 VN.n21 VSUBS 0.0308f
C901 VN.n22 VSUBS 0.054003f
C902 VN.n23 VSUBS 0.813319f
C903 VN.n24 VSUBS 0.032464f
C904 VN.n25 VSUBS 0.057943f
C905 VN.n26 VSUBS 0.0308f
C906 VN.n27 VSUBS 0.0308f
C907 VN.n28 VSUBS 0.0308f
C908 VN.n29 VSUBS 0.052612f
C909 VN.n30 VSUBS 0.050602f
C910 VN.n31 VSUBS 0.910616f
C911 VN.n32 VSUBS 0.039046f
C912 VN.n33 VSUBS 0.040607f
C913 VN.t5 VSUBS 2.29422f
C914 VN.n34 VSUBS 0.036775f
C915 VN.n35 VSUBS 0.0308f
C916 VN.t6 VSUBS 2.29422f
C917 VN.n36 VSUBS 0.047538f
C918 VN.n37 VSUBS 0.0308f
C919 VN.t2 VSUBS 2.29422f
C920 VN.n38 VSUBS 0.057404f
C921 VN.n39 VSUBS 0.0308f
C922 VN.t7 VSUBS 2.29422f
C923 VN.n40 VSUBS 0.90156f
C924 VN.t3 VSUBS 2.47695f
C925 VN.n41 VSUBS 0.880809f
C926 VN.n42 VSUBS 0.259615f
C927 VN.n43 VSUBS 0.054003f
C928 VN.n44 VSUBS 0.047538f
C929 VN.n45 VSUBS 0.042388f
C930 VN.n46 VSUBS 0.0308f
C931 VN.n47 VSUBS 0.0308f
C932 VN.n48 VSUBS 0.0308f
C933 VN.n49 VSUBS 0.842382f
C934 VN.n50 VSUBS 0.057404f
C935 VN.n51 VSUBS 0.042388f
C936 VN.n52 VSUBS 0.0308f
C937 VN.n53 VSUBS 0.0308f
C938 VN.n54 VSUBS 0.0308f
C939 VN.n55 VSUBS 0.054003f
C940 VN.n56 VSUBS 0.813319f
C941 VN.n57 VSUBS 0.032464f
C942 VN.n58 VSUBS 0.057943f
C943 VN.n59 VSUBS 0.0308f
C944 VN.n60 VSUBS 0.0308f
C945 VN.n61 VSUBS 0.0308f
C946 VN.n62 VSUBS 0.052612f
C947 VN.n63 VSUBS 0.050602f
C948 VN.n64 VSUBS 0.910616f
C949 VN.n65 VSUBS 1.7786f
C950 VDD1.t0 VSUBS 2.9359f
C951 VDD1.t5 VSUBS 0.281008f
C952 VDD1.t3 VSUBS 0.281008f
C953 VDD1.n0 VSUBS 2.23771f
C954 VDD1.n1 VSUBS 1.51604f
C955 VDD1.t8 VSUBS 2.93588f
C956 VDD1.t7 VSUBS 0.281008f
C957 VDD1.t2 VSUBS 0.281008f
C958 VDD1.n2 VSUBS 2.2377f
C959 VDD1.n3 VSUBS 1.50736f
C960 VDD1.t4 VSUBS 0.281008f
C961 VDD1.t9 VSUBS 0.281008f
C962 VDD1.n4 VSUBS 2.2546f
C963 VDD1.n5 VSUBS 3.37726f
C964 VDD1.t1 VSUBS 0.281008f
C965 VDD1.t6 VSUBS 0.281008f
C966 VDD1.n6 VSUBS 2.2377f
C967 VDD1.n7 VSUBS 3.62539f
C968 VTAIL.t8 VSUBS 0.288158f
C969 VTAIL.t1 VSUBS 0.288158f
C970 VTAIL.n0 VSUBS 2.14533f
C971 VTAIL.n1 VSUBS 0.91688f
C972 VTAIL.t18 VSUBS 2.82027f
C973 VTAIL.n2 VSUBS 1.07033f
C974 VTAIL.t10 VSUBS 0.288158f
C975 VTAIL.t14 VSUBS 0.288158f
C976 VTAIL.n3 VSUBS 2.14533f
C977 VTAIL.n4 VSUBS 1.01226f
C978 VTAIL.t19 VSUBS 0.288158f
C979 VTAIL.t13 VSUBS 0.288158f
C980 VTAIL.n5 VSUBS 2.14533f
C981 VTAIL.n6 VSUBS 2.59941f
C982 VTAIL.t5 VSUBS 0.288158f
C983 VTAIL.t4 VSUBS 0.288158f
C984 VTAIL.n7 VSUBS 2.14535f
C985 VTAIL.n8 VSUBS 2.59939f
C986 VTAIL.t3 VSUBS 0.288158f
C987 VTAIL.t6 VSUBS 0.288158f
C988 VTAIL.n9 VSUBS 2.14535f
C989 VTAIL.n10 VSUBS 1.01224f
C990 VTAIL.t2 VSUBS 2.8203f
C991 VTAIL.n11 VSUBS 1.0703f
C992 VTAIL.t15 VSUBS 0.288158f
C993 VTAIL.t11 VSUBS 0.288158f
C994 VTAIL.n12 VSUBS 2.14535f
C995 VTAIL.n13 VSUBS 0.959359f
C996 VTAIL.t12 VSUBS 0.288158f
C997 VTAIL.t17 VSUBS 0.288158f
C998 VTAIL.n14 VSUBS 2.14535f
C999 VTAIL.n15 VSUBS 1.01224f
C1000 VTAIL.t16 VSUBS 2.82027f
C1001 VTAIL.n16 VSUBS 2.51922f
C1002 VTAIL.t7 VSUBS 2.82027f
C1003 VTAIL.n17 VSUBS 2.51922f
C1004 VTAIL.t9 VSUBS 0.288158f
C1005 VTAIL.t0 VSUBS 0.288158f
C1006 VTAIL.n18 VSUBS 2.14533f
C1007 VTAIL.n19 VSUBS 0.863609f
C1008 VP.n0 VSUBS 0.04374f
C1009 VP.t0 VSUBS 2.47119f
C1010 VP.n1 VSUBS 0.039612f
C1011 VP.n2 VSUBS 0.033176f
C1012 VP.t5 VSUBS 2.47119f
C1013 VP.n3 VSUBS 0.051205f
C1014 VP.n4 VSUBS 0.033176f
C1015 VP.t7 VSUBS 2.47119f
C1016 VP.n5 VSUBS 0.061832f
C1017 VP.n6 VSUBS 0.033176f
C1018 VP.t2 VSUBS 2.47119f
C1019 VP.n7 VSUBS 0.876056f
C1020 VP.n8 VSUBS 0.033176f
C1021 VP.n9 VSUBS 0.05667f
C1022 VP.n10 VSUBS 0.04374f
C1023 VP.t3 VSUBS 2.47119f
C1024 VP.n11 VSUBS 0.039612f
C1025 VP.n12 VSUBS 0.033176f
C1026 VP.t8 VSUBS 2.47119f
C1027 VP.n13 VSUBS 0.051205f
C1028 VP.n14 VSUBS 0.033176f
C1029 VP.t6 VSUBS 2.47119f
C1030 VP.n15 VSUBS 0.061832f
C1031 VP.n16 VSUBS 0.033176f
C1032 VP.t4 VSUBS 2.47119f
C1033 VP.n17 VSUBS 0.971104f
C1034 VP.t9 VSUBS 2.66801f
C1035 VP.n18 VSUBS 0.948752f
C1036 VP.n19 VSUBS 0.279641f
C1037 VP.n20 VSUBS 0.058169f
C1038 VP.n21 VSUBS 0.051205f
C1039 VP.n22 VSUBS 0.045658f
C1040 VP.n23 VSUBS 0.033176f
C1041 VP.n24 VSUBS 0.033176f
C1042 VP.n25 VSUBS 0.033176f
C1043 VP.n26 VSUBS 0.907361f
C1044 VP.n27 VSUBS 0.061832f
C1045 VP.n28 VSUBS 0.045658f
C1046 VP.n29 VSUBS 0.033176f
C1047 VP.n30 VSUBS 0.033176f
C1048 VP.n31 VSUBS 0.033176f
C1049 VP.n32 VSUBS 0.058169f
C1050 VP.n33 VSUBS 0.876056f
C1051 VP.n34 VSUBS 0.034969f
C1052 VP.n35 VSUBS 0.062413f
C1053 VP.n36 VSUBS 0.033176f
C1054 VP.n37 VSUBS 0.033176f
C1055 VP.n38 VSUBS 0.033176f
C1056 VP.n39 VSUBS 0.05667f
C1057 VP.n40 VSUBS 0.054506f
C1058 VP.n41 VSUBS 0.980859f
C1059 VP.n42 VSUBS 1.89804f
C1060 VP.n43 VSUBS 1.92134f
C1061 VP.t1 VSUBS 2.47119f
C1062 VP.n44 VSUBS 0.980859f
C1063 VP.n45 VSUBS 0.054506f
C1064 VP.n46 VSUBS 0.04374f
C1065 VP.n47 VSUBS 0.033176f
C1066 VP.n48 VSUBS 0.033176f
C1067 VP.n49 VSUBS 0.039612f
C1068 VP.n50 VSUBS 0.062413f
C1069 VP.n51 VSUBS 0.034969f
C1070 VP.n52 VSUBS 0.033176f
C1071 VP.n53 VSUBS 0.033176f
C1072 VP.n54 VSUBS 0.058169f
C1073 VP.n55 VSUBS 0.051205f
C1074 VP.n56 VSUBS 0.045658f
C1075 VP.n57 VSUBS 0.033176f
C1076 VP.n58 VSUBS 0.033176f
C1077 VP.n59 VSUBS 0.033176f
C1078 VP.n60 VSUBS 0.907361f
C1079 VP.n61 VSUBS 0.061832f
C1080 VP.n62 VSUBS 0.045658f
C1081 VP.n63 VSUBS 0.033176f
C1082 VP.n64 VSUBS 0.033176f
C1083 VP.n65 VSUBS 0.033176f
C1084 VP.n66 VSUBS 0.058169f
C1085 VP.n67 VSUBS 0.876056f
C1086 VP.n68 VSUBS 0.034969f
C1087 VP.n69 VSUBS 0.062413f
C1088 VP.n70 VSUBS 0.033176f
C1089 VP.n71 VSUBS 0.033176f
C1090 VP.n72 VSUBS 0.033176f
C1091 VP.n73 VSUBS 0.05667f
C1092 VP.n74 VSUBS 0.054506f
C1093 VP.n75 VSUBS 0.980859f
C1094 VP.n76 VSUBS 0.042058f
.ends

