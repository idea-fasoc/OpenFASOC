* NGSPICE file created from diff_pair_sample_0877.ext - technology: sky130A

.subckt diff_pair_sample_0877 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t18 B.t0 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
X1 VTAIL.t2 VN.t0 VDD2.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
X2 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=4.0209 pd=21.4 as=0 ps=0 w=10.31 l=0.7
X3 VDD1.t8 VP.t1 VTAIL.t15 B.t6 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=4.0209 ps=21.4 w=10.31 l=0.7
X4 VDD1.t7 VP.t2 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=4.0209 pd=21.4 as=1.70115 ps=10.64 w=10.31 l=0.7
X5 VTAIL.t17 VP.t3 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
X6 VDD1.t5 VP.t4 VTAIL.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=4.0209 pd=21.4 as=1.70115 ps=10.64 w=10.31 l=0.7
X7 VDD2.t8 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=4.0209 pd=21.4 as=1.70115 ps=10.64 w=10.31 l=0.7
X8 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=4.0209 pd=21.4 as=0 ps=0 w=10.31 l=0.7
X9 VDD1.t4 VP.t5 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
X10 VDD2.t7 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
X11 VTAIL.t12 VP.t6 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
X12 VDD2.t6 VN.t3 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=4.0209 ps=21.4 w=10.31 l=0.7
X13 VTAIL.t10 VP.t7 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
X14 VDD1.t1 VP.t8 VTAIL.t11 B.t9 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=4.0209 ps=21.4 w=10.31 l=0.7
X15 VTAIL.t4 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
X16 VDD2.t4 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
X17 VTAIL.t9 VP.t9 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
X18 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=4.0209 pd=21.4 as=0 ps=0 w=10.31 l=0.7
X19 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.0209 pd=21.4 as=0 ps=0 w=10.31 l=0.7
X20 VDD2.t3 VN.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=4.0209 ps=21.4 w=10.31 l=0.7
X21 VDD2.t2 VN.t7 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=4.0209 pd=21.4 as=1.70115 ps=10.64 w=10.31 l=0.7
X22 VTAIL.t7 VN.t8 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
X23 VTAIL.t3 VN.t9 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.70115 pd=10.64 as=1.70115 ps=10.64 w=10.31 l=0.7
R0 VP.n7 VP.t2 434.17
R1 VP.n18 VP.t4 411.421
R2 VP.n22 VP.t3 411.421
R3 VP.n24 VP.t5 411.421
R4 VP.n28 VP.t9 411.421
R5 VP.n30 VP.t8 411.421
R6 VP.n16 VP.t1 411.421
R7 VP.n14 VP.t6 411.421
R8 VP.n6 VP.t0 411.421
R9 VP.n8 VP.t7 411.421
R10 VP.n31 VP.n30 161.3
R11 VP.n10 VP.n9 161.3
R12 VP.n11 VP.n6 161.3
R13 VP.n13 VP.n12 161.3
R14 VP.n14 VP.n5 161.3
R15 VP.n15 VP.n4 161.3
R16 VP.n17 VP.n16 161.3
R17 VP.n29 VP.n0 161.3
R18 VP.n28 VP.n27 161.3
R19 VP.n26 VP.n1 161.3
R20 VP.n25 VP.n24 161.3
R21 VP.n23 VP.n2 161.3
R22 VP.n22 VP.n21 161.3
R23 VP.n20 VP.n3 161.3
R24 VP.n19 VP.n18 161.3
R25 VP.n10 VP.n7 44.8741
R26 VP.n19 VP.n17 41.5043
R27 VP.n18 VP.n3 30.6732
R28 VP.n30 VP.n29 30.6732
R29 VP.n16 VP.n15 30.6732
R30 VP.n23 VP.n22 26.2914
R31 VP.n28 VP.n1 26.2914
R32 VP.n14 VP.n13 26.2914
R33 VP.n9 VP.n8 26.2914
R34 VP.n24 VP.n23 21.9096
R35 VP.n24 VP.n1 21.9096
R36 VP.n13 VP.n6 21.9096
R37 VP.n9 VP.n6 21.9096
R38 VP.n8 VP.n7 19.0667
R39 VP.n22 VP.n3 17.5278
R40 VP.n29 VP.n28 17.5278
R41 VP.n15 VP.n14 17.5278
R42 VP.n11 VP.n10 0.189894
R43 VP.n12 VP.n11 0.189894
R44 VP.n12 VP.n5 0.189894
R45 VP.n5 VP.n4 0.189894
R46 VP.n17 VP.n4 0.189894
R47 VP.n20 VP.n19 0.189894
R48 VP.n21 VP.n20 0.189894
R49 VP.n21 VP.n2 0.189894
R50 VP.n25 VP.n2 0.189894
R51 VP.n26 VP.n25 0.189894
R52 VP.n27 VP.n26 0.189894
R53 VP.n27 VP.n0 0.189894
R54 VP.n31 VP.n0 0.189894
R55 VP VP.n31 0.0516364
R56 VTAIL.n11 VTAIL.t19 47.5307
R57 VTAIL.n17 VTAIL.t6 47.5305
R58 VTAIL.n2 VTAIL.t11 47.5305
R59 VTAIL.n16 VTAIL.t15 47.5305
R60 VTAIL.n15 VTAIL.n14 45.6103
R61 VTAIL.n13 VTAIL.n12 45.6103
R62 VTAIL.n10 VTAIL.n9 45.6103
R63 VTAIL.n8 VTAIL.n7 45.6103
R64 VTAIL.n19 VTAIL.n18 45.61
R65 VTAIL.n1 VTAIL.n0 45.61
R66 VTAIL.n4 VTAIL.n3 45.61
R67 VTAIL.n6 VTAIL.n5 45.61
R68 VTAIL.n8 VTAIL.n6 23.0307
R69 VTAIL.n17 VTAIL.n16 22.1427
R70 VTAIL.n18 VTAIL.t0 1.92097
R71 VTAIL.n18 VTAIL.t4 1.92097
R72 VTAIL.n0 VTAIL.t8 1.92097
R73 VTAIL.n0 VTAIL.t3 1.92097
R74 VTAIL.n3 VTAIL.t14 1.92097
R75 VTAIL.n3 VTAIL.t9 1.92097
R76 VTAIL.n5 VTAIL.t13 1.92097
R77 VTAIL.n5 VTAIL.t17 1.92097
R78 VTAIL.n14 VTAIL.t18 1.92097
R79 VTAIL.n14 VTAIL.t12 1.92097
R80 VTAIL.n12 VTAIL.t16 1.92097
R81 VTAIL.n12 VTAIL.t10 1.92097
R82 VTAIL.n9 VTAIL.t1 1.92097
R83 VTAIL.n9 VTAIL.t2 1.92097
R84 VTAIL.n7 VTAIL.t5 1.92097
R85 VTAIL.n7 VTAIL.t7 1.92097
R86 VTAIL.n13 VTAIL.n11 0.914293
R87 VTAIL.n2 VTAIL.n1 0.914293
R88 VTAIL.n10 VTAIL.n8 0.888431
R89 VTAIL.n11 VTAIL.n10 0.888431
R90 VTAIL.n15 VTAIL.n13 0.888431
R91 VTAIL.n16 VTAIL.n15 0.888431
R92 VTAIL.n6 VTAIL.n4 0.888431
R93 VTAIL.n4 VTAIL.n2 0.888431
R94 VTAIL.n19 VTAIL.n17 0.888431
R95 VTAIL VTAIL.n1 0.724638
R96 VTAIL VTAIL.n19 0.164293
R97 VDD1.n1 VDD1.t7 65.0974
R98 VDD1.n3 VDD1.t5 65.0972
R99 VDD1.n5 VDD1.n4 62.8994
R100 VDD1.n1 VDD1.n0 62.2891
R101 VDD1.n7 VDD1.n6 62.2889
R102 VDD1.n3 VDD1.n2 62.2888
R103 VDD1.n7 VDD1.n5 37.8479
R104 VDD1.n6 VDD1.t3 1.92097
R105 VDD1.n6 VDD1.t8 1.92097
R106 VDD1.n0 VDD1.t2 1.92097
R107 VDD1.n0 VDD1.t9 1.92097
R108 VDD1.n4 VDD1.t0 1.92097
R109 VDD1.n4 VDD1.t1 1.92097
R110 VDD1.n2 VDD1.t6 1.92097
R111 VDD1.n2 VDD1.t4 1.92097
R112 VDD1 VDD1.n7 0.608259
R113 VDD1 VDD1.n1 0.280672
R114 VDD1.n5 VDD1.n3 0.167137
R115 B.n472 B.n97 585
R116 B.n97 B.n50 585
R117 B.n474 B.n473 585
R118 B.n476 B.n96 585
R119 B.n479 B.n478 585
R120 B.n480 B.n95 585
R121 B.n482 B.n481 585
R122 B.n484 B.n94 585
R123 B.n487 B.n486 585
R124 B.n488 B.n93 585
R125 B.n490 B.n489 585
R126 B.n492 B.n92 585
R127 B.n495 B.n494 585
R128 B.n496 B.n91 585
R129 B.n498 B.n497 585
R130 B.n500 B.n90 585
R131 B.n503 B.n502 585
R132 B.n504 B.n89 585
R133 B.n506 B.n505 585
R134 B.n508 B.n88 585
R135 B.n511 B.n510 585
R136 B.n512 B.n87 585
R137 B.n514 B.n513 585
R138 B.n516 B.n86 585
R139 B.n519 B.n518 585
R140 B.n520 B.n85 585
R141 B.n522 B.n521 585
R142 B.n524 B.n84 585
R143 B.n527 B.n526 585
R144 B.n528 B.n83 585
R145 B.n530 B.n529 585
R146 B.n532 B.n82 585
R147 B.n535 B.n534 585
R148 B.n536 B.n81 585
R149 B.n538 B.n537 585
R150 B.n540 B.n80 585
R151 B.n542 B.n541 585
R152 B.n544 B.n543 585
R153 B.n547 B.n546 585
R154 B.n548 B.n75 585
R155 B.n550 B.n549 585
R156 B.n552 B.n74 585
R157 B.n555 B.n554 585
R158 B.n556 B.n73 585
R159 B.n558 B.n557 585
R160 B.n560 B.n72 585
R161 B.n563 B.n562 585
R162 B.n565 B.n69 585
R163 B.n567 B.n566 585
R164 B.n569 B.n68 585
R165 B.n572 B.n571 585
R166 B.n573 B.n67 585
R167 B.n575 B.n574 585
R168 B.n577 B.n66 585
R169 B.n580 B.n579 585
R170 B.n581 B.n65 585
R171 B.n583 B.n582 585
R172 B.n585 B.n64 585
R173 B.n588 B.n587 585
R174 B.n589 B.n63 585
R175 B.n591 B.n590 585
R176 B.n593 B.n62 585
R177 B.n596 B.n595 585
R178 B.n597 B.n61 585
R179 B.n599 B.n598 585
R180 B.n601 B.n60 585
R181 B.n604 B.n603 585
R182 B.n605 B.n59 585
R183 B.n607 B.n606 585
R184 B.n609 B.n58 585
R185 B.n612 B.n611 585
R186 B.n613 B.n57 585
R187 B.n615 B.n614 585
R188 B.n617 B.n56 585
R189 B.n620 B.n619 585
R190 B.n621 B.n55 585
R191 B.n623 B.n622 585
R192 B.n625 B.n54 585
R193 B.n628 B.n627 585
R194 B.n629 B.n53 585
R195 B.n631 B.n630 585
R196 B.n633 B.n52 585
R197 B.n636 B.n635 585
R198 B.n637 B.n51 585
R199 B.n471 B.n49 585
R200 B.n640 B.n49 585
R201 B.n470 B.n48 585
R202 B.n641 B.n48 585
R203 B.n469 B.n47 585
R204 B.n642 B.n47 585
R205 B.n468 B.n467 585
R206 B.n467 B.n43 585
R207 B.n466 B.n42 585
R208 B.n648 B.n42 585
R209 B.n465 B.n41 585
R210 B.n649 B.n41 585
R211 B.n464 B.n40 585
R212 B.n650 B.n40 585
R213 B.n463 B.n462 585
R214 B.n462 B.n36 585
R215 B.n461 B.n35 585
R216 B.n656 B.n35 585
R217 B.n460 B.n34 585
R218 B.n657 B.n34 585
R219 B.n459 B.n33 585
R220 B.n658 B.n33 585
R221 B.n458 B.n457 585
R222 B.n457 B.n29 585
R223 B.n456 B.n28 585
R224 B.n664 B.n28 585
R225 B.n455 B.n27 585
R226 B.n665 B.n27 585
R227 B.n454 B.n26 585
R228 B.n666 B.n26 585
R229 B.n453 B.n452 585
R230 B.n452 B.n22 585
R231 B.n451 B.n21 585
R232 B.n672 B.n21 585
R233 B.n450 B.n20 585
R234 B.n673 B.n20 585
R235 B.n449 B.n19 585
R236 B.n674 B.n19 585
R237 B.n448 B.n447 585
R238 B.n447 B.n18 585
R239 B.n446 B.n14 585
R240 B.n680 B.n14 585
R241 B.n445 B.n13 585
R242 B.n681 B.n13 585
R243 B.n444 B.n12 585
R244 B.n682 B.n12 585
R245 B.n443 B.n442 585
R246 B.n442 B.n8 585
R247 B.n441 B.n7 585
R248 B.n688 B.n7 585
R249 B.n440 B.n6 585
R250 B.n689 B.n6 585
R251 B.n439 B.n5 585
R252 B.n690 B.n5 585
R253 B.n438 B.n437 585
R254 B.n437 B.n4 585
R255 B.n436 B.n98 585
R256 B.n436 B.n435 585
R257 B.n426 B.n99 585
R258 B.n100 B.n99 585
R259 B.n428 B.n427 585
R260 B.n429 B.n428 585
R261 B.n425 B.n105 585
R262 B.n105 B.n104 585
R263 B.n424 B.n423 585
R264 B.n423 B.n422 585
R265 B.n107 B.n106 585
R266 B.n415 B.n107 585
R267 B.n414 B.n413 585
R268 B.n416 B.n414 585
R269 B.n412 B.n112 585
R270 B.n112 B.n111 585
R271 B.n411 B.n410 585
R272 B.n410 B.n409 585
R273 B.n114 B.n113 585
R274 B.n115 B.n114 585
R275 B.n402 B.n401 585
R276 B.n403 B.n402 585
R277 B.n400 B.n119 585
R278 B.n123 B.n119 585
R279 B.n399 B.n398 585
R280 B.n398 B.n397 585
R281 B.n121 B.n120 585
R282 B.n122 B.n121 585
R283 B.n390 B.n389 585
R284 B.n391 B.n390 585
R285 B.n388 B.n128 585
R286 B.n128 B.n127 585
R287 B.n387 B.n386 585
R288 B.n386 B.n385 585
R289 B.n130 B.n129 585
R290 B.n131 B.n130 585
R291 B.n378 B.n377 585
R292 B.n379 B.n378 585
R293 B.n376 B.n136 585
R294 B.n136 B.n135 585
R295 B.n375 B.n374 585
R296 B.n374 B.n373 585
R297 B.n138 B.n137 585
R298 B.n139 B.n138 585
R299 B.n366 B.n365 585
R300 B.n367 B.n366 585
R301 B.n364 B.n144 585
R302 B.n144 B.n143 585
R303 B.n363 B.n362 585
R304 B.n362 B.n361 585
R305 B.n358 B.n148 585
R306 B.n357 B.n356 585
R307 B.n354 B.n149 585
R308 B.n354 B.n147 585
R309 B.n353 B.n352 585
R310 B.n351 B.n350 585
R311 B.n349 B.n151 585
R312 B.n347 B.n346 585
R313 B.n345 B.n152 585
R314 B.n344 B.n343 585
R315 B.n341 B.n153 585
R316 B.n339 B.n338 585
R317 B.n337 B.n154 585
R318 B.n336 B.n335 585
R319 B.n333 B.n155 585
R320 B.n331 B.n330 585
R321 B.n329 B.n156 585
R322 B.n328 B.n327 585
R323 B.n325 B.n157 585
R324 B.n323 B.n322 585
R325 B.n321 B.n158 585
R326 B.n320 B.n319 585
R327 B.n317 B.n159 585
R328 B.n315 B.n314 585
R329 B.n313 B.n160 585
R330 B.n312 B.n311 585
R331 B.n309 B.n161 585
R332 B.n307 B.n306 585
R333 B.n305 B.n162 585
R334 B.n304 B.n303 585
R335 B.n301 B.n163 585
R336 B.n299 B.n298 585
R337 B.n297 B.n164 585
R338 B.n296 B.n295 585
R339 B.n293 B.n165 585
R340 B.n291 B.n290 585
R341 B.n289 B.n166 585
R342 B.n288 B.n287 585
R343 B.n285 B.n284 585
R344 B.n283 B.n282 585
R345 B.n281 B.n171 585
R346 B.n279 B.n278 585
R347 B.n277 B.n172 585
R348 B.n276 B.n275 585
R349 B.n273 B.n173 585
R350 B.n271 B.n270 585
R351 B.n269 B.n174 585
R352 B.n267 B.n266 585
R353 B.n264 B.n177 585
R354 B.n262 B.n261 585
R355 B.n260 B.n178 585
R356 B.n259 B.n258 585
R357 B.n256 B.n179 585
R358 B.n254 B.n253 585
R359 B.n252 B.n180 585
R360 B.n251 B.n250 585
R361 B.n248 B.n181 585
R362 B.n246 B.n245 585
R363 B.n244 B.n182 585
R364 B.n243 B.n242 585
R365 B.n240 B.n183 585
R366 B.n238 B.n237 585
R367 B.n236 B.n184 585
R368 B.n235 B.n234 585
R369 B.n232 B.n185 585
R370 B.n230 B.n229 585
R371 B.n228 B.n186 585
R372 B.n227 B.n226 585
R373 B.n224 B.n187 585
R374 B.n222 B.n221 585
R375 B.n220 B.n188 585
R376 B.n219 B.n218 585
R377 B.n216 B.n189 585
R378 B.n214 B.n213 585
R379 B.n212 B.n190 585
R380 B.n211 B.n210 585
R381 B.n208 B.n191 585
R382 B.n206 B.n205 585
R383 B.n204 B.n192 585
R384 B.n203 B.n202 585
R385 B.n200 B.n193 585
R386 B.n198 B.n197 585
R387 B.n196 B.n195 585
R388 B.n146 B.n145 585
R389 B.n360 B.n359 585
R390 B.n361 B.n360 585
R391 B.n142 B.n141 585
R392 B.n143 B.n142 585
R393 B.n369 B.n368 585
R394 B.n368 B.n367 585
R395 B.n370 B.n140 585
R396 B.n140 B.n139 585
R397 B.n372 B.n371 585
R398 B.n373 B.n372 585
R399 B.n134 B.n133 585
R400 B.n135 B.n134 585
R401 B.n381 B.n380 585
R402 B.n380 B.n379 585
R403 B.n382 B.n132 585
R404 B.n132 B.n131 585
R405 B.n384 B.n383 585
R406 B.n385 B.n384 585
R407 B.n126 B.n125 585
R408 B.n127 B.n126 585
R409 B.n393 B.n392 585
R410 B.n392 B.n391 585
R411 B.n394 B.n124 585
R412 B.n124 B.n122 585
R413 B.n396 B.n395 585
R414 B.n397 B.n396 585
R415 B.n118 B.n117 585
R416 B.n123 B.n118 585
R417 B.n405 B.n404 585
R418 B.n404 B.n403 585
R419 B.n406 B.n116 585
R420 B.n116 B.n115 585
R421 B.n408 B.n407 585
R422 B.n409 B.n408 585
R423 B.n110 B.n109 585
R424 B.n111 B.n110 585
R425 B.n418 B.n417 585
R426 B.n417 B.n416 585
R427 B.n419 B.n108 585
R428 B.n415 B.n108 585
R429 B.n421 B.n420 585
R430 B.n422 B.n421 585
R431 B.n103 B.n102 585
R432 B.n104 B.n103 585
R433 B.n431 B.n430 585
R434 B.n430 B.n429 585
R435 B.n432 B.n101 585
R436 B.n101 B.n100 585
R437 B.n434 B.n433 585
R438 B.n435 B.n434 585
R439 B.n2 B.n0 585
R440 B.n4 B.n2 585
R441 B.n3 B.n1 585
R442 B.n689 B.n3 585
R443 B.n687 B.n686 585
R444 B.n688 B.n687 585
R445 B.n685 B.n9 585
R446 B.n9 B.n8 585
R447 B.n684 B.n683 585
R448 B.n683 B.n682 585
R449 B.n11 B.n10 585
R450 B.n681 B.n11 585
R451 B.n679 B.n678 585
R452 B.n680 B.n679 585
R453 B.n677 B.n15 585
R454 B.n18 B.n15 585
R455 B.n676 B.n675 585
R456 B.n675 B.n674 585
R457 B.n17 B.n16 585
R458 B.n673 B.n17 585
R459 B.n671 B.n670 585
R460 B.n672 B.n671 585
R461 B.n669 B.n23 585
R462 B.n23 B.n22 585
R463 B.n668 B.n667 585
R464 B.n667 B.n666 585
R465 B.n25 B.n24 585
R466 B.n665 B.n25 585
R467 B.n663 B.n662 585
R468 B.n664 B.n663 585
R469 B.n661 B.n30 585
R470 B.n30 B.n29 585
R471 B.n660 B.n659 585
R472 B.n659 B.n658 585
R473 B.n32 B.n31 585
R474 B.n657 B.n32 585
R475 B.n655 B.n654 585
R476 B.n656 B.n655 585
R477 B.n653 B.n37 585
R478 B.n37 B.n36 585
R479 B.n652 B.n651 585
R480 B.n651 B.n650 585
R481 B.n39 B.n38 585
R482 B.n649 B.n39 585
R483 B.n647 B.n646 585
R484 B.n648 B.n647 585
R485 B.n645 B.n44 585
R486 B.n44 B.n43 585
R487 B.n644 B.n643 585
R488 B.n643 B.n642 585
R489 B.n46 B.n45 585
R490 B.n641 B.n46 585
R491 B.n639 B.n638 585
R492 B.n640 B.n639 585
R493 B.n692 B.n691 585
R494 B.n691 B.n690 585
R495 B.n175 B.t10 557.923
R496 B.n167 B.t18 557.923
R497 B.n70 B.t21 557.923
R498 B.n76 B.t14 557.923
R499 B.n360 B.n148 535.745
R500 B.n639 B.n51 535.745
R501 B.n362 B.n146 535.745
R502 B.n97 B.n49 535.745
R503 B.n475 B.n50 256.663
R504 B.n477 B.n50 256.663
R505 B.n483 B.n50 256.663
R506 B.n485 B.n50 256.663
R507 B.n491 B.n50 256.663
R508 B.n493 B.n50 256.663
R509 B.n499 B.n50 256.663
R510 B.n501 B.n50 256.663
R511 B.n507 B.n50 256.663
R512 B.n509 B.n50 256.663
R513 B.n515 B.n50 256.663
R514 B.n517 B.n50 256.663
R515 B.n523 B.n50 256.663
R516 B.n525 B.n50 256.663
R517 B.n531 B.n50 256.663
R518 B.n533 B.n50 256.663
R519 B.n539 B.n50 256.663
R520 B.n79 B.n50 256.663
R521 B.n545 B.n50 256.663
R522 B.n551 B.n50 256.663
R523 B.n553 B.n50 256.663
R524 B.n559 B.n50 256.663
R525 B.n561 B.n50 256.663
R526 B.n568 B.n50 256.663
R527 B.n570 B.n50 256.663
R528 B.n576 B.n50 256.663
R529 B.n578 B.n50 256.663
R530 B.n584 B.n50 256.663
R531 B.n586 B.n50 256.663
R532 B.n592 B.n50 256.663
R533 B.n594 B.n50 256.663
R534 B.n600 B.n50 256.663
R535 B.n602 B.n50 256.663
R536 B.n608 B.n50 256.663
R537 B.n610 B.n50 256.663
R538 B.n616 B.n50 256.663
R539 B.n618 B.n50 256.663
R540 B.n624 B.n50 256.663
R541 B.n626 B.n50 256.663
R542 B.n632 B.n50 256.663
R543 B.n634 B.n50 256.663
R544 B.n355 B.n147 256.663
R545 B.n150 B.n147 256.663
R546 B.n348 B.n147 256.663
R547 B.n342 B.n147 256.663
R548 B.n340 B.n147 256.663
R549 B.n334 B.n147 256.663
R550 B.n332 B.n147 256.663
R551 B.n326 B.n147 256.663
R552 B.n324 B.n147 256.663
R553 B.n318 B.n147 256.663
R554 B.n316 B.n147 256.663
R555 B.n310 B.n147 256.663
R556 B.n308 B.n147 256.663
R557 B.n302 B.n147 256.663
R558 B.n300 B.n147 256.663
R559 B.n294 B.n147 256.663
R560 B.n292 B.n147 256.663
R561 B.n286 B.n147 256.663
R562 B.n170 B.n147 256.663
R563 B.n280 B.n147 256.663
R564 B.n274 B.n147 256.663
R565 B.n272 B.n147 256.663
R566 B.n265 B.n147 256.663
R567 B.n263 B.n147 256.663
R568 B.n257 B.n147 256.663
R569 B.n255 B.n147 256.663
R570 B.n249 B.n147 256.663
R571 B.n247 B.n147 256.663
R572 B.n241 B.n147 256.663
R573 B.n239 B.n147 256.663
R574 B.n233 B.n147 256.663
R575 B.n231 B.n147 256.663
R576 B.n225 B.n147 256.663
R577 B.n223 B.n147 256.663
R578 B.n217 B.n147 256.663
R579 B.n215 B.n147 256.663
R580 B.n209 B.n147 256.663
R581 B.n207 B.n147 256.663
R582 B.n201 B.n147 256.663
R583 B.n199 B.n147 256.663
R584 B.n194 B.n147 256.663
R585 B.n360 B.n142 163.367
R586 B.n368 B.n142 163.367
R587 B.n368 B.n140 163.367
R588 B.n372 B.n140 163.367
R589 B.n372 B.n134 163.367
R590 B.n380 B.n134 163.367
R591 B.n380 B.n132 163.367
R592 B.n384 B.n132 163.367
R593 B.n384 B.n126 163.367
R594 B.n392 B.n126 163.367
R595 B.n392 B.n124 163.367
R596 B.n396 B.n124 163.367
R597 B.n396 B.n118 163.367
R598 B.n404 B.n118 163.367
R599 B.n404 B.n116 163.367
R600 B.n408 B.n116 163.367
R601 B.n408 B.n110 163.367
R602 B.n417 B.n110 163.367
R603 B.n417 B.n108 163.367
R604 B.n421 B.n108 163.367
R605 B.n421 B.n103 163.367
R606 B.n430 B.n103 163.367
R607 B.n430 B.n101 163.367
R608 B.n434 B.n101 163.367
R609 B.n434 B.n2 163.367
R610 B.n691 B.n2 163.367
R611 B.n691 B.n3 163.367
R612 B.n687 B.n3 163.367
R613 B.n687 B.n9 163.367
R614 B.n683 B.n9 163.367
R615 B.n683 B.n11 163.367
R616 B.n679 B.n11 163.367
R617 B.n679 B.n15 163.367
R618 B.n675 B.n15 163.367
R619 B.n675 B.n17 163.367
R620 B.n671 B.n17 163.367
R621 B.n671 B.n23 163.367
R622 B.n667 B.n23 163.367
R623 B.n667 B.n25 163.367
R624 B.n663 B.n25 163.367
R625 B.n663 B.n30 163.367
R626 B.n659 B.n30 163.367
R627 B.n659 B.n32 163.367
R628 B.n655 B.n32 163.367
R629 B.n655 B.n37 163.367
R630 B.n651 B.n37 163.367
R631 B.n651 B.n39 163.367
R632 B.n647 B.n39 163.367
R633 B.n647 B.n44 163.367
R634 B.n643 B.n44 163.367
R635 B.n643 B.n46 163.367
R636 B.n639 B.n46 163.367
R637 B.n356 B.n354 163.367
R638 B.n354 B.n353 163.367
R639 B.n350 B.n349 163.367
R640 B.n347 B.n152 163.367
R641 B.n343 B.n341 163.367
R642 B.n339 B.n154 163.367
R643 B.n335 B.n333 163.367
R644 B.n331 B.n156 163.367
R645 B.n327 B.n325 163.367
R646 B.n323 B.n158 163.367
R647 B.n319 B.n317 163.367
R648 B.n315 B.n160 163.367
R649 B.n311 B.n309 163.367
R650 B.n307 B.n162 163.367
R651 B.n303 B.n301 163.367
R652 B.n299 B.n164 163.367
R653 B.n295 B.n293 163.367
R654 B.n291 B.n166 163.367
R655 B.n287 B.n285 163.367
R656 B.n282 B.n281 163.367
R657 B.n279 B.n172 163.367
R658 B.n275 B.n273 163.367
R659 B.n271 B.n174 163.367
R660 B.n266 B.n264 163.367
R661 B.n262 B.n178 163.367
R662 B.n258 B.n256 163.367
R663 B.n254 B.n180 163.367
R664 B.n250 B.n248 163.367
R665 B.n246 B.n182 163.367
R666 B.n242 B.n240 163.367
R667 B.n238 B.n184 163.367
R668 B.n234 B.n232 163.367
R669 B.n230 B.n186 163.367
R670 B.n226 B.n224 163.367
R671 B.n222 B.n188 163.367
R672 B.n218 B.n216 163.367
R673 B.n214 B.n190 163.367
R674 B.n210 B.n208 163.367
R675 B.n206 B.n192 163.367
R676 B.n202 B.n200 163.367
R677 B.n198 B.n195 163.367
R678 B.n362 B.n144 163.367
R679 B.n366 B.n144 163.367
R680 B.n366 B.n138 163.367
R681 B.n374 B.n138 163.367
R682 B.n374 B.n136 163.367
R683 B.n378 B.n136 163.367
R684 B.n378 B.n130 163.367
R685 B.n386 B.n130 163.367
R686 B.n386 B.n128 163.367
R687 B.n390 B.n128 163.367
R688 B.n390 B.n121 163.367
R689 B.n398 B.n121 163.367
R690 B.n398 B.n119 163.367
R691 B.n402 B.n119 163.367
R692 B.n402 B.n114 163.367
R693 B.n410 B.n114 163.367
R694 B.n410 B.n112 163.367
R695 B.n414 B.n112 163.367
R696 B.n414 B.n107 163.367
R697 B.n423 B.n107 163.367
R698 B.n423 B.n105 163.367
R699 B.n428 B.n105 163.367
R700 B.n428 B.n99 163.367
R701 B.n436 B.n99 163.367
R702 B.n437 B.n436 163.367
R703 B.n437 B.n5 163.367
R704 B.n6 B.n5 163.367
R705 B.n7 B.n6 163.367
R706 B.n442 B.n7 163.367
R707 B.n442 B.n12 163.367
R708 B.n13 B.n12 163.367
R709 B.n14 B.n13 163.367
R710 B.n447 B.n14 163.367
R711 B.n447 B.n19 163.367
R712 B.n20 B.n19 163.367
R713 B.n21 B.n20 163.367
R714 B.n452 B.n21 163.367
R715 B.n452 B.n26 163.367
R716 B.n27 B.n26 163.367
R717 B.n28 B.n27 163.367
R718 B.n457 B.n28 163.367
R719 B.n457 B.n33 163.367
R720 B.n34 B.n33 163.367
R721 B.n35 B.n34 163.367
R722 B.n462 B.n35 163.367
R723 B.n462 B.n40 163.367
R724 B.n41 B.n40 163.367
R725 B.n42 B.n41 163.367
R726 B.n467 B.n42 163.367
R727 B.n467 B.n47 163.367
R728 B.n48 B.n47 163.367
R729 B.n49 B.n48 163.367
R730 B.n635 B.n633 163.367
R731 B.n631 B.n53 163.367
R732 B.n627 B.n625 163.367
R733 B.n623 B.n55 163.367
R734 B.n619 B.n617 163.367
R735 B.n615 B.n57 163.367
R736 B.n611 B.n609 163.367
R737 B.n607 B.n59 163.367
R738 B.n603 B.n601 163.367
R739 B.n599 B.n61 163.367
R740 B.n595 B.n593 163.367
R741 B.n591 B.n63 163.367
R742 B.n587 B.n585 163.367
R743 B.n583 B.n65 163.367
R744 B.n579 B.n577 163.367
R745 B.n575 B.n67 163.367
R746 B.n571 B.n569 163.367
R747 B.n567 B.n69 163.367
R748 B.n562 B.n560 163.367
R749 B.n558 B.n73 163.367
R750 B.n554 B.n552 163.367
R751 B.n550 B.n75 163.367
R752 B.n546 B.n544 163.367
R753 B.n541 B.n540 163.367
R754 B.n538 B.n81 163.367
R755 B.n534 B.n532 163.367
R756 B.n530 B.n83 163.367
R757 B.n526 B.n524 163.367
R758 B.n522 B.n85 163.367
R759 B.n518 B.n516 163.367
R760 B.n514 B.n87 163.367
R761 B.n510 B.n508 163.367
R762 B.n506 B.n89 163.367
R763 B.n502 B.n500 163.367
R764 B.n498 B.n91 163.367
R765 B.n494 B.n492 163.367
R766 B.n490 B.n93 163.367
R767 B.n486 B.n484 163.367
R768 B.n482 B.n95 163.367
R769 B.n478 B.n476 163.367
R770 B.n474 B.n97 163.367
R771 B.n361 B.n147 100.93
R772 B.n640 B.n50 100.93
R773 B.n175 B.t13 90.167
R774 B.n76 B.t16 90.167
R775 B.n167 B.t20 90.1542
R776 B.n70 B.t22 90.1542
R777 B.n355 B.n148 71.676
R778 B.n353 B.n150 71.676
R779 B.n349 B.n348 71.676
R780 B.n342 B.n152 71.676
R781 B.n341 B.n340 71.676
R782 B.n334 B.n154 71.676
R783 B.n333 B.n332 71.676
R784 B.n326 B.n156 71.676
R785 B.n325 B.n324 71.676
R786 B.n318 B.n158 71.676
R787 B.n317 B.n316 71.676
R788 B.n310 B.n160 71.676
R789 B.n309 B.n308 71.676
R790 B.n302 B.n162 71.676
R791 B.n301 B.n300 71.676
R792 B.n294 B.n164 71.676
R793 B.n293 B.n292 71.676
R794 B.n286 B.n166 71.676
R795 B.n285 B.n170 71.676
R796 B.n281 B.n280 71.676
R797 B.n274 B.n172 71.676
R798 B.n273 B.n272 71.676
R799 B.n265 B.n174 71.676
R800 B.n264 B.n263 71.676
R801 B.n257 B.n178 71.676
R802 B.n256 B.n255 71.676
R803 B.n249 B.n180 71.676
R804 B.n248 B.n247 71.676
R805 B.n241 B.n182 71.676
R806 B.n240 B.n239 71.676
R807 B.n233 B.n184 71.676
R808 B.n232 B.n231 71.676
R809 B.n225 B.n186 71.676
R810 B.n224 B.n223 71.676
R811 B.n217 B.n188 71.676
R812 B.n216 B.n215 71.676
R813 B.n209 B.n190 71.676
R814 B.n208 B.n207 71.676
R815 B.n201 B.n192 71.676
R816 B.n200 B.n199 71.676
R817 B.n195 B.n194 71.676
R818 B.n634 B.n51 71.676
R819 B.n633 B.n632 71.676
R820 B.n626 B.n53 71.676
R821 B.n625 B.n624 71.676
R822 B.n618 B.n55 71.676
R823 B.n617 B.n616 71.676
R824 B.n610 B.n57 71.676
R825 B.n609 B.n608 71.676
R826 B.n602 B.n59 71.676
R827 B.n601 B.n600 71.676
R828 B.n594 B.n61 71.676
R829 B.n593 B.n592 71.676
R830 B.n586 B.n63 71.676
R831 B.n585 B.n584 71.676
R832 B.n578 B.n65 71.676
R833 B.n577 B.n576 71.676
R834 B.n570 B.n67 71.676
R835 B.n569 B.n568 71.676
R836 B.n561 B.n69 71.676
R837 B.n560 B.n559 71.676
R838 B.n553 B.n73 71.676
R839 B.n552 B.n551 71.676
R840 B.n545 B.n75 71.676
R841 B.n544 B.n79 71.676
R842 B.n540 B.n539 71.676
R843 B.n533 B.n81 71.676
R844 B.n532 B.n531 71.676
R845 B.n525 B.n83 71.676
R846 B.n524 B.n523 71.676
R847 B.n517 B.n85 71.676
R848 B.n516 B.n515 71.676
R849 B.n509 B.n87 71.676
R850 B.n508 B.n507 71.676
R851 B.n501 B.n89 71.676
R852 B.n500 B.n499 71.676
R853 B.n493 B.n91 71.676
R854 B.n492 B.n491 71.676
R855 B.n485 B.n93 71.676
R856 B.n484 B.n483 71.676
R857 B.n477 B.n95 71.676
R858 B.n476 B.n475 71.676
R859 B.n475 B.n474 71.676
R860 B.n478 B.n477 71.676
R861 B.n483 B.n482 71.676
R862 B.n486 B.n485 71.676
R863 B.n491 B.n490 71.676
R864 B.n494 B.n493 71.676
R865 B.n499 B.n498 71.676
R866 B.n502 B.n501 71.676
R867 B.n507 B.n506 71.676
R868 B.n510 B.n509 71.676
R869 B.n515 B.n514 71.676
R870 B.n518 B.n517 71.676
R871 B.n523 B.n522 71.676
R872 B.n526 B.n525 71.676
R873 B.n531 B.n530 71.676
R874 B.n534 B.n533 71.676
R875 B.n539 B.n538 71.676
R876 B.n541 B.n79 71.676
R877 B.n546 B.n545 71.676
R878 B.n551 B.n550 71.676
R879 B.n554 B.n553 71.676
R880 B.n559 B.n558 71.676
R881 B.n562 B.n561 71.676
R882 B.n568 B.n567 71.676
R883 B.n571 B.n570 71.676
R884 B.n576 B.n575 71.676
R885 B.n579 B.n578 71.676
R886 B.n584 B.n583 71.676
R887 B.n587 B.n586 71.676
R888 B.n592 B.n591 71.676
R889 B.n595 B.n594 71.676
R890 B.n600 B.n599 71.676
R891 B.n603 B.n602 71.676
R892 B.n608 B.n607 71.676
R893 B.n611 B.n610 71.676
R894 B.n616 B.n615 71.676
R895 B.n619 B.n618 71.676
R896 B.n624 B.n623 71.676
R897 B.n627 B.n626 71.676
R898 B.n632 B.n631 71.676
R899 B.n635 B.n634 71.676
R900 B.n356 B.n355 71.676
R901 B.n350 B.n150 71.676
R902 B.n348 B.n347 71.676
R903 B.n343 B.n342 71.676
R904 B.n340 B.n339 71.676
R905 B.n335 B.n334 71.676
R906 B.n332 B.n331 71.676
R907 B.n327 B.n326 71.676
R908 B.n324 B.n323 71.676
R909 B.n319 B.n318 71.676
R910 B.n316 B.n315 71.676
R911 B.n311 B.n310 71.676
R912 B.n308 B.n307 71.676
R913 B.n303 B.n302 71.676
R914 B.n300 B.n299 71.676
R915 B.n295 B.n294 71.676
R916 B.n292 B.n291 71.676
R917 B.n287 B.n286 71.676
R918 B.n282 B.n170 71.676
R919 B.n280 B.n279 71.676
R920 B.n275 B.n274 71.676
R921 B.n272 B.n271 71.676
R922 B.n266 B.n265 71.676
R923 B.n263 B.n262 71.676
R924 B.n258 B.n257 71.676
R925 B.n255 B.n254 71.676
R926 B.n250 B.n249 71.676
R927 B.n247 B.n246 71.676
R928 B.n242 B.n241 71.676
R929 B.n239 B.n238 71.676
R930 B.n234 B.n233 71.676
R931 B.n231 B.n230 71.676
R932 B.n226 B.n225 71.676
R933 B.n223 B.n222 71.676
R934 B.n218 B.n217 71.676
R935 B.n215 B.n214 71.676
R936 B.n210 B.n209 71.676
R937 B.n207 B.n206 71.676
R938 B.n202 B.n201 71.676
R939 B.n199 B.n198 71.676
R940 B.n194 B.n146 71.676
R941 B.n176 B.t12 70.1912
R942 B.n77 B.t17 70.1912
R943 B.n168 B.t19 70.1785
R944 B.n71 B.t23 70.1785
R945 B.n268 B.n176 59.5399
R946 B.n169 B.n168 59.5399
R947 B.n564 B.n71 59.5399
R948 B.n78 B.n77 59.5399
R949 B.n361 B.n143 47.9954
R950 B.n367 B.n143 47.9954
R951 B.n367 B.n139 47.9954
R952 B.n373 B.n139 47.9954
R953 B.n379 B.n135 47.9954
R954 B.n379 B.n131 47.9954
R955 B.n385 B.n131 47.9954
R956 B.n385 B.n127 47.9954
R957 B.n391 B.n127 47.9954
R958 B.n397 B.n122 47.9954
R959 B.n397 B.n123 47.9954
R960 B.n403 B.n115 47.9954
R961 B.n409 B.n115 47.9954
R962 B.n416 B.n111 47.9954
R963 B.n416 B.n415 47.9954
R964 B.n422 B.n104 47.9954
R965 B.n429 B.n104 47.9954
R966 B.n435 B.n100 47.9954
R967 B.n435 B.n4 47.9954
R968 B.n690 B.n4 47.9954
R969 B.n690 B.n689 47.9954
R970 B.n689 B.n688 47.9954
R971 B.n688 B.n8 47.9954
R972 B.n682 B.n681 47.9954
R973 B.n681 B.n680 47.9954
R974 B.n674 B.n18 47.9954
R975 B.n674 B.n673 47.9954
R976 B.n672 B.n22 47.9954
R977 B.n666 B.n22 47.9954
R978 B.n665 B.n664 47.9954
R979 B.n664 B.n29 47.9954
R980 B.n658 B.n657 47.9954
R981 B.n657 B.n656 47.9954
R982 B.n656 B.n36 47.9954
R983 B.n650 B.n36 47.9954
R984 B.n650 B.n649 47.9954
R985 B.n648 B.n43 47.9954
R986 B.n642 B.n43 47.9954
R987 B.n642 B.n641 47.9954
R988 B.n641 B.n640 47.9954
R989 B.n429 B.t9 42.3489
R990 B.n682 B.t8 42.3489
R991 B.n415 B.t2 40.9373
R992 B.n18 B.t3 40.9373
R993 B.n409 B.t1 39.5257
R994 B.t0 B.n672 39.5257
R995 B.n123 B.t7 38.1141
R996 B.t4 B.n665 38.1141
R997 B.n391 B.t5 36.7025
R998 B.n658 B.t6 36.7025
R999 B.n638 B.n637 34.8103
R1000 B.n472 B.n471 34.8103
R1001 B.n363 B.n145 34.8103
R1002 B.n359 B.n358 34.8103
R1003 B.n373 B.t11 25.4095
R1004 B.t15 B.n648 25.4095
R1005 B.t11 B.n135 22.5863
R1006 B.n649 B.t15 22.5863
R1007 B.n176 B.n175 19.9763
R1008 B.n168 B.n167 19.9763
R1009 B.n71 B.n70 19.9763
R1010 B.n77 B.n76 19.9763
R1011 B B.n692 18.0485
R1012 B.t5 B.n122 11.2934
R1013 B.t6 B.n29 11.2934
R1014 B.n637 B.n636 10.6151
R1015 B.n636 B.n52 10.6151
R1016 B.n630 B.n52 10.6151
R1017 B.n630 B.n629 10.6151
R1018 B.n629 B.n628 10.6151
R1019 B.n628 B.n54 10.6151
R1020 B.n622 B.n54 10.6151
R1021 B.n622 B.n621 10.6151
R1022 B.n621 B.n620 10.6151
R1023 B.n620 B.n56 10.6151
R1024 B.n614 B.n56 10.6151
R1025 B.n614 B.n613 10.6151
R1026 B.n613 B.n612 10.6151
R1027 B.n612 B.n58 10.6151
R1028 B.n606 B.n58 10.6151
R1029 B.n606 B.n605 10.6151
R1030 B.n605 B.n604 10.6151
R1031 B.n604 B.n60 10.6151
R1032 B.n598 B.n60 10.6151
R1033 B.n598 B.n597 10.6151
R1034 B.n597 B.n596 10.6151
R1035 B.n596 B.n62 10.6151
R1036 B.n590 B.n62 10.6151
R1037 B.n590 B.n589 10.6151
R1038 B.n589 B.n588 10.6151
R1039 B.n588 B.n64 10.6151
R1040 B.n582 B.n64 10.6151
R1041 B.n582 B.n581 10.6151
R1042 B.n581 B.n580 10.6151
R1043 B.n580 B.n66 10.6151
R1044 B.n574 B.n66 10.6151
R1045 B.n574 B.n573 10.6151
R1046 B.n573 B.n572 10.6151
R1047 B.n572 B.n68 10.6151
R1048 B.n566 B.n68 10.6151
R1049 B.n566 B.n565 10.6151
R1050 B.n563 B.n72 10.6151
R1051 B.n557 B.n72 10.6151
R1052 B.n557 B.n556 10.6151
R1053 B.n556 B.n555 10.6151
R1054 B.n555 B.n74 10.6151
R1055 B.n549 B.n74 10.6151
R1056 B.n549 B.n548 10.6151
R1057 B.n548 B.n547 10.6151
R1058 B.n543 B.n542 10.6151
R1059 B.n542 B.n80 10.6151
R1060 B.n537 B.n80 10.6151
R1061 B.n537 B.n536 10.6151
R1062 B.n536 B.n535 10.6151
R1063 B.n535 B.n82 10.6151
R1064 B.n529 B.n82 10.6151
R1065 B.n529 B.n528 10.6151
R1066 B.n528 B.n527 10.6151
R1067 B.n527 B.n84 10.6151
R1068 B.n521 B.n84 10.6151
R1069 B.n521 B.n520 10.6151
R1070 B.n520 B.n519 10.6151
R1071 B.n519 B.n86 10.6151
R1072 B.n513 B.n86 10.6151
R1073 B.n513 B.n512 10.6151
R1074 B.n512 B.n511 10.6151
R1075 B.n511 B.n88 10.6151
R1076 B.n505 B.n88 10.6151
R1077 B.n505 B.n504 10.6151
R1078 B.n504 B.n503 10.6151
R1079 B.n503 B.n90 10.6151
R1080 B.n497 B.n90 10.6151
R1081 B.n497 B.n496 10.6151
R1082 B.n496 B.n495 10.6151
R1083 B.n495 B.n92 10.6151
R1084 B.n489 B.n92 10.6151
R1085 B.n489 B.n488 10.6151
R1086 B.n488 B.n487 10.6151
R1087 B.n487 B.n94 10.6151
R1088 B.n481 B.n94 10.6151
R1089 B.n481 B.n480 10.6151
R1090 B.n480 B.n479 10.6151
R1091 B.n479 B.n96 10.6151
R1092 B.n473 B.n96 10.6151
R1093 B.n473 B.n472 10.6151
R1094 B.n364 B.n363 10.6151
R1095 B.n365 B.n364 10.6151
R1096 B.n365 B.n137 10.6151
R1097 B.n375 B.n137 10.6151
R1098 B.n376 B.n375 10.6151
R1099 B.n377 B.n376 10.6151
R1100 B.n377 B.n129 10.6151
R1101 B.n387 B.n129 10.6151
R1102 B.n388 B.n387 10.6151
R1103 B.n389 B.n388 10.6151
R1104 B.n389 B.n120 10.6151
R1105 B.n399 B.n120 10.6151
R1106 B.n400 B.n399 10.6151
R1107 B.n401 B.n400 10.6151
R1108 B.n401 B.n113 10.6151
R1109 B.n411 B.n113 10.6151
R1110 B.n412 B.n411 10.6151
R1111 B.n413 B.n412 10.6151
R1112 B.n413 B.n106 10.6151
R1113 B.n424 B.n106 10.6151
R1114 B.n425 B.n424 10.6151
R1115 B.n427 B.n425 10.6151
R1116 B.n427 B.n426 10.6151
R1117 B.n426 B.n98 10.6151
R1118 B.n438 B.n98 10.6151
R1119 B.n439 B.n438 10.6151
R1120 B.n440 B.n439 10.6151
R1121 B.n441 B.n440 10.6151
R1122 B.n443 B.n441 10.6151
R1123 B.n444 B.n443 10.6151
R1124 B.n445 B.n444 10.6151
R1125 B.n446 B.n445 10.6151
R1126 B.n448 B.n446 10.6151
R1127 B.n449 B.n448 10.6151
R1128 B.n450 B.n449 10.6151
R1129 B.n451 B.n450 10.6151
R1130 B.n453 B.n451 10.6151
R1131 B.n454 B.n453 10.6151
R1132 B.n455 B.n454 10.6151
R1133 B.n456 B.n455 10.6151
R1134 B.n458 B.n456 10.6151
R1135 B.n459 B.n458 10.6151
R1136 B.n460 B.n459 10.6151
R1137 B.n461 B.n460 10.6151
R1138 B.n463 B.n461 10.6151
R1139 B.n464 B.n463 10.6151
R1140 B.n465 B.n464 10.6151
R1141 B.n466 B.n465 10.6151
R1142 B.n468 B.n466 10.6151
R1143 B.n469 B.n468 10.6151
R1144 B.n470 B.n469 10.6151
R1145 B.n471 B.n470 10.6151
R1146 B.n358 B.n357 10.6151
R1147 B.n357 B.n149 10.6151
R1148 B.n352 B.n149 10.6151
R1149 B.n352 B.n351 10.6151
R1150 B.n351 B.n151 10.6151
R1151 B.n346 B.n151 10.6151
R1152 B.n346 B.n345 10.6151
R1153 B.n345 B.n344 10.6151
R1154 B.n344 B.n153 10.6151
R1155 B.n338 B.n153 10.6151
R1156 B.n338 B.n337 10.6151
R1157 B.n337 B.n336 10.6151
R1158 B.n336 B.n155 10.6151
R1159 B.n330 B.n155 10.6151
R1160 B.n330 B.n329 10.6151
R1161 B.n329 B.n328 10.6151
R1162 B.n328 B.n157 10.6151
R1163 B.n322 B.n157 10.6151
R1164 B.n322 B.n321 10.6151
R1165 B.n321 B.n320 10.6151
R1166 B.n320 B.n159 10.6151
R1167 B.n314 B.n159 10.6151
R1168 B.n314 B.n313 10.6151
R1169 B.n313 B.n312 10.6151
R1170 B.n312 B.n161 10.6151
R1171 B.n306 B.n161 10.6151
R1172 B.n306 B.n305 10.6151
R1173 B.n305 B.n304 10.6151
R1174 B.n304 B.n163 10.6151
R1175 B.n298 B.n163 10.6151
R1176 B.n298 B.n297 10.6151
R1177 B.n297 B.n296 10.6151
R1178 B.n296 B.n165 10.6151
R1179 B.n290 B.n165 10.6151
R1180 B.n290 B.n289 10.6151
R1181 B.n289 B.n288 10.6151
R1182 B.n284 B.n283 10.6151
R1183 B.n283 B.n171 10.6151
R1184 B.n278 B.n171 10.6151
R1185 B.n278 B.n277 10.6151
R1186 B.n277 B.n276 10.6151
R1187 B.n276 B.n173 10.6151
R1188 B.n270 B.n173 10.6151
R1189 B.n270 B.n269 10.6151
R1190 B.n267 B.n177 10.6151
R1191 B.n261 B.n177 10.6151
R1192 B.n261 B.n260 10.6151
R1193 B.n260 B.n259 10.6151
R1194 B.n259 B.n179 10.6151
R1195 B.n253 B.n179 10.6151
R1196 B.n253 B.n252 10.6151
R1197 B.n252 B.n251 10.6151
R1198 B.n251 B.n181 10.6151
R1199 B.n245 B.n181 10.6151
R1200 B.n245 B.n244 10.6151
R1201 B.n244 B.n243 10.6151
R1202 B.n243 B.n183 10.6151
R1203 B.n237 B.n183 10.6151
R1204 B.n237 B.n236 10.6151
R1205 B.n236 B.n235 10.6151
R1206 B.n235 B.n185 10.6151
R1207 B.n229 B.n185 10.6151
R1208 B.n229 B.n228 10.6151
R1209 B.n228 B.n227 10.6151
R1210 B.n227 B.n187 10.6151
R1211 B.n221 B.n187 10.6151
R1212 B.n221 B.n220 10.6151
R1213 B.n220 B.n219 10.6151
R1214 B.n219 B.n189 10.6151
R1215 B.n213 B.n189 10.6151
R1216 B.n213 B.n212 10.6151
R1217 B.n212 B.n211 10.6151
R1218 B.n211 B.n191 10.6151
R1219 B.n205 B.n191 10.6151
R1220 B.n205 B.n204 10.6151
R1221 B.n204 B.n203 10.6151
R1222 B.n203 B.n193 10.6151
R1223 B.n197 B.n193 10.6151
R1224 B.n197 B.n196 10.6151
R1225 B.n196 B.n145 10.6151
R1226 B.n359 B.n141 10.6151
R1227 B.n369 B.n141 10.6151
R1228 B.n370 B.n369 10.6151
R1229 B.n371 B.n370 10.6151
R1230 B.n371 B.n133 10.6151
R1231 B.n381 B.n133 10.6151
R1232 B.n382 B.n381 10.6151
R1233 B.n383 B.n382 10.6151
R1234 B.n383 B.n125 10.6151
R1235 B.n393 B.n125 10.6151
R1236 B.n394 B.n393 10.6151
R1237 B.n395 B.n394 10.6151
R1238 B.n395 B.n117 10.6151
R1239 B.n405 B.n117 10.6151
R1240 B.n406 B.n405 10.6151
R1241 B.n407 B.n406 10.6151
R1242 B.n407 B.n109 10.6151
R1243 B.n418 B.n109 10.6151
R1244 B.n419 B.n418 10.6151
R1245 B.n420 B.n419 10.6151
R1246 B.n420 B.n102 10.6151
R1247 B.n431 B.n102 10.6151
R1248 B.n432 B.n431 10.6151
R1249 B.n433 B.n432 10.6151
R1250 B.n433 B.n0 10.6151
R1251 B.n686 B.n1 10.6151
R1252 B.n686 B.n685 10.6151
R1253 B.n685 B.n684 10.6151
R1254 B.n684 B.n10 10.6151
R1255 B.n678 B.n10 10.6151
R1256 B.n678 B.n677 10.6151
R1257 B.n677 B.n676 10.6151
R1258 B.n676 B.n16 10.6151
R1259 B.n670 B.n16 10.6151
R1260 B.n670 B.n669 10.6151
R1261 B.n669 B.n668 10.6151
R1262 B.n668 B.n24 10.6151
R1263 B.n662 B.n24 10.6151
R1264 B.n662 B.n661 10.6151
R1265 B.n661 B.n660 10.6151
R1266 B.n660 B.n31 10.6151
R1267 B.n654 B.n31 10.6151
R1268 B.n654 B.n653 10.6151
R1269 B.n653 B.n652 10.6151
R1270 B.n652 B.n38 10.6151
R1271 B.n646 B.n38 10.6151
R1272 B.n646 B.n645 10.6151
R1273 B.n645 B.n644 10.6151
R1274 B.n644 B.n45 10.6151
R1275 B.n638 B.n45 10.6151
R1276 B.n403 B.t7 9.8818
R1277 B.n666 B.t4 9.8818
R1278 B.t1 B.n111 8.47018
R1279 B.n673 B.t0 8.47018
R1280 B.n422 B.t2 7.05857
R1281 B.n680 B.t3 7.05857
R1282 B.n564 B.n563 6.5566
R1283 B.n547 B.n78 6.5566
R1284 B.n284 B.n169 6.5566
R1285 B.n269 B.n268 6.5566
R1286 B.t9 B.n100 5.64696
R1287 B.t8 B.n8 5.64696
R1288 B.n565 B.n564 4.05904
R1289 B.n543 B.n78 4.05904
R1290 B.n288 B.n169 4.05904
R1291 B.n268 B.n267 4.05904
R1292 B.n692 B.n0 2.81026
R1293 B.n692 B.n1 2.81026
R1294 VN.n3 VN.t7 434.17
R1295 VN.n17 VN.t3 434.17
R1296 VN.n4 VN.t9 411.421
R1297 VN.n6 VN.t5 411.421
R1298 VN.n10 VN.t4 411.421
R1299 VN.n12 VN.t6 411.421
R1300 VN.n18 VN.t0 411.421
R1301 VN.n20 VN.t2 411.421
R1302 VN.n24 VN.t8 411.421
R1303 VN.n26 VN.t1 411.421
R1304 VN.n13 VN.n12 161.3
R1305 VN.n27 VN.n26 161.3
R1306 VN.n25 VN.n14 161.3
R1307 VN.n24 VN.n23 161.3
R1308 VN.n22 VN.n15 161.3
R1309 VN.n21 VN.n20 161.3
R1310 VN.n19 VN.n16 161.3
R1311 VN.n11 VN.n0 161.3
R1312 VN.n10 VN.n9 161.3
R1313 VN.n8 VN.n1 161.3
R1314 VN.n7 VN.n6 161.3
R1315 VN.n5 VN.n2 161.3
R1316 VN.n17 VN.n16 44.8741
R1317 VN.n3 VN.n2 44.8741
R1318 VN VN.n27 41.885
R1319 VN.n12 VN.n11 30.6732
R1320 VN.n26 VN.n25 30.6732
R1321 VN.n5 VN.n4 26.2914
R1322 VN.n10 VN.n1 26.2914
R1323 VN.n19 VN.n18 26.2914
R1324 VN.n24 VN.n15 26.2914
R1325 VN.n6 VN.n5 21.9096
R1326 VN.n6 VN.n1 21.9096
R1327 VN.n20 VN.n19 21.9096
R1328 VN.n20 VN.n15 21.9096
R1329 VN.n4 VN.n3 19.0667
R1330 VN.n18 VN.n17 19.0667
R1331 VN.n11 VN.n10 17.5278
R1332 VN.n25 VN.n24 17.5278
R1333 VN.n27 VN.n14 0.189894
R1334 VN.n23 VN.n14 0.189894
R1335 VN.n23 VN.n22 0.189894
R1336 VN.n22 VN.n21 0.189894
R1337 VN.n21 VN.n16 0.189894
R1338 VN.n7 VN.n2 0.189894
R1339 VN.n8 VN.n7 0.189894
R1340 VN.n9 VN.n8 0.189894
R1341 VN.n9 VN.n0 0.189894
R1342 VN.n13 VN.n0 0.189894
R1343 VN VN.n13 0.0516364
R1344 VDD2.n1 VDD2.t2 65.0972
R1345 VDD2.n4 VDD2.t8 64.2095
R1346 VDD2.n3 VDD2.n2 62.8994
R1347 VDD2 VDD2.n7 62.8966
R1348 VDD2.n6 VDD2.n5 62.2891
R1349 VDD2.n1 VDD2.n0 62.2888
R1350 VDD2.n4 VDD2.n3 36.8209
R1351 VDD2.n7 VDD2.t9 1.92097
R1352 VDD2.n7 VDD2.t6 1.92097
R1353 VDD2.n5 VDD2.t1 1.92097
R1354 VDD2.n5 VDD2.t7 1.92097
R1355 VDD2.n2 VDD2.t5 1.92097
R1356 VDD2.n2 VDD2.t3 1.92097
R1357 VDD2.n0 VDD2.t0 1.92097
R1358 VDD2.n0 VDD2.t4 1.92097
R1359 VDD2.n6 VDD2.n4 0.888431
R1360 VDD2 VDD2.n6 0.280672
R1361 VDD2.n3 VDD2.n1 0.167137
C0 VDD2 VDD1 0.969442f
C1 VP VTAIL 5.73108f
C2 VN VTAIL 5.71654f
C3 VN VP 5.2851f
C4 VDD2 VTAIL 12.6016f
C5 VDD1 VTAIL 12.566501f
C6 VDD2 VP 0.340953f
C7 VDD1 VP 6.00241f
C8 VDD2 VN 5.81423f
C9 VDD1 VN 0.14865f
C10 VDD2 B 4.668561f
C11 VDD1 B 4.594674f
C12 VTAIL B 5.881037f
C13 VN B 9.265349f
C14 VP B 7.390994f
C15 VDD2.t2 B 2.24434f
C16 VDD2.t0 B 0.199356f
C17 VDD2.t4 B 0.199356f
C18 VDD2.n0 B 1.75887f
C19 VDD2.n1 B 0.625235f
C20 VDD2.t5 B 0.199356f
C21 VDD2.t3 B 0.199356f
C22 VDD2.n2 B 1.76207f
C23 VDD2.n3 B 1.7616f
C24 VDD2.t8 B 2.23967f
C25 VDD2.n4 B 2.20513f
C26 VDD2.t1 B 0.199356f
C27 VDD2.t7 B 0.199356f
C28 VDD2.n5 B 1.75888f
C29 VDD2.n6 B 0.292391f
C30 VDD2.t9 B 0.199356f
C31 VDD2.t6 B 0.199356f
C32 VDD2.n7 B 1.76204f
C33 VN.n0 B 0.042838f
C34 VN.n1 B 0.009721f
C35 VN.n2 B 0.178927f
C36 VN.t7 B 0.903321f
C37 VN.n3 B 0.347104f
C38 VN.t9 B 0.884353f
C39 VN.n4 B 0.366482f
C40 VN.n5 B 0.009721f
C41 VN.t5 B 0.884353f
C42 VN.n6 B 0.362166f
C43 VN.n7 B 0.042838f
C44 VN.n8 B 0.042838f
C45 VN.n9 B 0.042838f
C46 VN.t4 B 0.884353f
C47 VN.n10 B 0.362166f
C48 VN.n11 B 0.009721f
C49 VN.t6 B 0.884353f
C50 VN.n12 B 0.359789f
C51 VN.n13 B 0.033198f
C52 VN.n14 B 0.042838f
C53 VN.n15 B 0.009721f
C54 VN.t8 B 0.884353f
C55 VN.n16 B 0.178927f
C56 VN.t3 B 0.903321f
C57 VN.n17 B 0.347104f
C58 VN.t0 B 0.884353f
C59 VN.n18 B 0.366482f
C60 VN.n19 B 0.009721f
C61 VN.t2 B 0.884353f
C62 VN.n20 B 0.362166f
C63 VN.n21 B 0.042838f
C64 VN.n22 B 0.042838f
C65 VN.n23 B 0.042838f
C66 VN.n24 B 0.362166f
C67 VN.n25 B 0.009721f
C68 VN.t1 B 0.884353f
C69 VN.n26 B 0.359789f
C70 VN.n27 B 1.7616f
C71 VDD1.t7 B 2.25765f
C72 VDD1.t2 B 0.200538f
C73 VDD1.t9 B 0.200538f
C74 VDD1.n0 B 1.7693f
C75 VDD1.n1 B 0.634515f
C76 VDD1.t5 B 2.25765f
C77 VDD1.t6 B 0.200538f
C78 VDD1.t4 B 0.200538f
C79 VDD1.n2 B 1.7693f
C80 VDD1.n3 B 0.628942f
C81 VDD1.t0 B 0.200538f
C82 VDD1.t1 B 0.200538f
C83 VDD1.n4 B 1.77252f
C84 VDD1.n5 B 1.8473f
C85 VDD1.t3 B 0.200538f
C86 VDD1.t8 B 0.200538f
C87 VDD1.n6 B 1.7693f
C88 VDD1.n7 B 2.2188f
C89 VTAIL.t8 B 0.211882f
C90 VTAIL.t3 B 0.211882f
C91 VTAIL.n0 B 1.79334f
C92 VTAIL.n1 B 0.390825f
C93 VTAIL.t11 B 2.28395f
C94 VTAIL.n2 B 0.491799f
C95 VTAIL.t14 B 0.211882f
C96 VTAIL.t9 B 0.211882f
C97 VTAIL.n3 B 1.79334f
C98 VTAIL.n4 B 0.402384f
C99 VTAIL.t13 B 0.211882f
C100 VTAIL.t17 B 0.211882f
C101 VTAIL.n5 B 1.79334f
C102 VTAIL.n6 B 1.57485f
C103 VTAIL.t5 B 0.211882f
C104 VTAIL.t7 B 0.211882f
C105 VTAIL.n7 B 1.79335f
C106 VTAIL.n8 B 1.57485f
C107 VTAIL.t1 B 0.211882f
C108 VTAIL.t2 B 0.211882f
C109 VTAIL.n9 B 1.79335f
C110 VTAIL.n10 B 0.402378f
C111 VTAIL.t19 B 2.28396f
C112 VTAIL.n11 B 0.491793f
C113 VTAIL.t16 B 0.211882f
C114 VTAIL.t10 B 0.211882f
C115 VTAIL.n12 B 1.79335f
C116 VTAIL.n13 B 0.404545f
C117 VTAIL.t18 B 0.211882f
C118 VTAIL.t12 B 0.211882f
C119 VTAIL.n14 B 1.79335f
C120 VTAIL.n15 B 0.402378f
C121 VTAIL.t15 B 2.28395f
C122 VTAIL.n16 B 1.58769f
C123 VTAIL.t6 B 2.28395f
C124 VTAIL.n17 B 1.58769f
C125 VTAIL.t0 B 0.211882f
C126 VTAIL.t4 B 0.211882f
C127 VTAIL.n18 B 1.79334f
C128 VTAIL.n19 B 0.341702f
C129 VP.n0 B 0.043504f
C130 VP.n1 B 0.009872f
C131 VP.n2 B 0.043504f
C132 VP.n3 B 0.009872f
C133 VP.n4 B 0.043504f
C134 VP.t1 B 0.898101f
C135 VP.t6 B 0.898101f
C136 VP.n5 B 0.043504f
C137 VP.t0 B 0.898101f
C138 VP.n6 B 0.367796f
C139 VP.t2 B 0.917363f
C140 VP.n7 B 0.3525f
C141 VP.t7 B 0.898101f
C142 VP.n8 B 0.372179f
C143 VP.n9 B 0.009872f
C144 VP.n10 B 0.181709f
C145 VP.n11 B 0.043504f
C146 VP.n12 B 0.043504f
C147 VP.n13 B 0.009872f
C148 VP.n14 B 0.367796f
C149 VP.n15 B 0.009872f
C150 VP.n16 B 0.365382f
C151 VP.n17 B 1.7604f
C152 VP.t4 B 0.898101f
C153 VP.n18 B 0.365382f
C154 VP.n19 B 1.79808f
C155 VP.n20 B 0.043504f
C156 VP.n21 B 0.043504f
C157 VP.t3 B 0.898101f
C158 VP.n22 B 0.367796f
C159 VP.n23 B 0.009872f
C160 VP.t5 B 0.898101f
C161 VP.n24 B 0.367796f
C162 VP.n25 B 0.043504f
C163 VP.n26 B 0.043504f
C164 VP.n27 B 0.043504f
C165 VP.t9 B 0.898101f
C166 VP.n28 B 0.367796f
C167 VP.n29 B 0.009872f
C168 VP.t8 B 0.898101f
C169 VP.n30 B 0.365382f
C170 VP.n31 B 0.033714f
.ends

