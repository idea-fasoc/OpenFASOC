* NGSPICE file created from diff_pair_sample_1795.ext - technology: sky130A

.subckt diff_pair_sample_1795 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=6.5715 pd=34.48 as=0 ps=0 w=16.85 l=0.58
X1 VTAIL.t11 VP.t0 VDD1.t3 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=2.78025 pd=17.18 as=2.78025 ps=17.18 w=16.85 l=0.58
X2 VTAIL.t10 VP.t1 VDD1.t2 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=2.78025 pd=17.18 as=2.78025 ps=17.18 w=16.85 l=0.58
X3 VDD1.t5 VP.t2 VTAIL.t9 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=2.78025 pd=17.18 as=6.5715 ps=34.48 w=16.85 l=0.58
X4 VDD2.t5 VN.t0 VTAIL.t3 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=2.78025 pd=17.18 as=6.5715 ps=34.48 w=16.85 l=0.58
X5 VTAIL.t4 VN.t1 VDD2.t4 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=2.78025 pd=17.18 as=2.78025 ps=17.18 w=16.85 l=0.58
X6 B.t8 B.t6 B.t7 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=6.5715 pd=34.48 as=0 ps=0 w=16.85 l=0.58
X7 VDD1.t4 VP.t3 VTAIL.t8 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=2.78025 pd=17.18 as=6.5715 ps=34.48 w=16.85 l=0.58
X8 B.t5 B.t3 B.t4 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=6.5715 pd=34.48 as=0 ps=0 w=16.85 l=0.58
X9 VTAIL.t5 VN.t2 VDD2.t3 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=2.78025 pd=17.18 as=2.78025 ps=17.18 w=16.85 l=0.58
X10 VDD2.t2 VN.t3 VTAIL.t2 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=6.5715 pd=34.48 as=2.78025 ps=17.18 w=16.85 l=0.58
X11 B.t2 B.t0 B.t1 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=6.5715 pd=34.48 as=0 ps=0 w=16.85 l=0.58
X12 VDD1.t0 VP.t4 VTAIL.t7 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=6.5715 pd=34.48 as=2.78025 ps=17.18 w=16.85 l=0.58
X13 VDD2.t1 VN.t4 VTAIL.t0 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=2.78025 pd=17.18 as=6.5715 ps=34.48 w=16.85 l=0.58
X14 VDD1.t1 VP.t5 VTAIL.t6 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=6.5715 pd=34.48 as=2.78025 ps=17.18 w=16.85 l=0.58
X15 VDD2.t0 VN.t5 VTAIL.t1 w_n1698_n4338# sky130_fd_pr__pfet_01v8 ad=6.5715 pd=34.48 as=2.78025 ps=17.18 w=16.85 l=0.58
R0 B.n124 B.t3 904.893
R1 B.n132 B.t0 904.893
R2 B.n40 B.t9 904.893
R3 B.n46 B.t6 904.893
R4 B.n439 B.n76 585
R5 B.n441 B.n440 585
R6 B.n442 B.n75 585
R7 B.n444 B.n443 585
R8 B.n445 B.n74 585
R9 B.n447 B.n446 585
R10 B.n448 B.n73 585
R11 B.n450 B.n449 585
R12 B.n451 B.n72 585
R13 B.n453 B.n452 585
R14 B.n454 B.n71 585
R15 B.n456 B.n455 585
R16 B.n457 B.n70 585
R17 B.n459 B.n458 585
R18 B.n460 B.n69 585
R19 B.n462 B.n461 585
R20 B.n463 B.n68 585
R21 B.n465 B.n464 585
R22 B.n466 B.n67 585
R23 B.n468 B.n467 585
R24 B.n469 B.n66 585
R25 B.n471 B.n470 585
R26 B.n472 B.n65 585
R27 B.n474 B.n473 585
R28 B.n475 B.n64 585
R29 B.n477 B.n476 585
R30 B.n478 B.n63 585
R31 B.n480 B.n479 585
R32 B.n481 B.n62 585
R33 B.n483 B.n482 585
R34 B.n484 B.n61 585
R35 B.n486 B.n485 585
R36 B.n487 B.n60 585
R37 B.n489 B.n488 585
R38 B.n490 B.n59 585
R39 B.n492 B.n491 585
R40 B.n493 B.n58 585
R41 B.n495 B.n494 585
R42 B.n496 B.n57 585
R43 B.n498 B.n497 585
R44 B.n499 B.n56 585
R45 B.n501 B.n500 585
R46 B.n502 B.n55 585
R47 B.n504 B.n503 585
R48 B.n505 B.n54 585
R49 B.n507 B.n506 585
R50 B.n508 B.n53 585
R51 B.n510 B.n509 585
R52 B.n511 B.n52 585
R53 B.n513 B.n512 585
R54 B.n514 B.n51 585
R55 B.n516 B.n515 585
R56 B.n517 B.n50 585
R57 B.n519 B.n518 585
R58 B.n520 B.n49 585
R59 B.n522 B.n521 585
R60 B.n524 B.n523 585
R61 B.n525 B.n45 585
R62 B.n527 B.n526 585
R63 B.n528 B.n44 585
R64 B.n530 B.n529 585
R65 B.n531 B.n43 585
R66 B.n533 B.n532 585
R67 B.n534 B.n42 585
R68 B.n536 B.n535 585
R69 B.n538 B.n39 585
R70 B.n540 B.n539 585
R71 B.n541 B.n38 585
R72 B.n543 B.n542 585
R73 B.n544 B.n37 585
R74 B.n546 B.n545 585
R75 B.n547 B.n36 585
R76 B.n549 B.n548 585
R77 B.n550 B.n35 585
R78 B.n552 B.n551 585
R79 B.n553 B.n34 585
R80 B.n555 B.n554 585
R81 B.n556 B.n33 585
R82 B.n558 B.n557 585
R83 B.n559 B.n32 585
R84 B.n561 B.n560 585
R85 B.n562 B.n31 585
R86 B.n564 B.n563 585
R87 B.n565 B.n30 585
R88 B.n567 B.n566 585
R89 B.n568 B.n29 585
R90 B.n570 B.n569 585
R91 B.n571 B.n28 585
R92 B.n573 B.n572 585
R93 B.n574 B.n27 585
R94 B.n576 B.n575 585
R95 B.n577 B.n26 585
R96 B.n579 B.n578 585
R97 B.n580 B.n25 585
R98 B.n582 B.n581 585
R99 B.n583 B.n24 585
R100 B.n585 B.n584 585
R101 B.n586 B.n23 585
R102 B.n588 B.n587 585
R103 B.n589 B.n22 585
R104 B.n591 B.n590 585
R105 B.n592 B.n21 585
R106 B.n594 B.n593 585
R107 B.n595 B.n20 585
R108 B.n597 B.n596 585
R109 B.n598 B.n19 585
R110 B.n600 B.n599 585
R111 B.n601 B.n18 585
R112 B.n603 B.n602 585
R113 B.n604 B.n17 585
R114 B.n606 B.n605 585
R115 B.n607 B.n16 585
R116 B.n609 B.n608 585
R117 B.n610 B.n15 585
R118 B.n612 B.n611 585
R119 B.n613 B.n14 585
R120 B.n615 B.n614 585
R121 B.n616 B.n13 585
R122 B.n618 B.n617 585
R123 B.n619 B.n12 585
R124 B.n621 B.n620 585
R125 B.n438 B.n437 585
R126 B.n436 B.n77 585
R127 B.n435 B.n434 585
R128 B.n433 B.n78 585
R129 B.n432 B.n431 585
R130 B.n430 B.n79 585
R131 B.n429 B.n428 585
R132 B.n427 B.n80 585
R133 B.n426 B.n425 585
R134 B.n424 B.n81 585
R135 B.n423 B.n422 585
R136 B.n421 B.n82 585
R137 B.n420 B.n419 585
R138 B.n418 B.n83 585
R139 B.n417 B.n416 585
R140 B.n415 B.n84 585
R141 B.n414 B.n413 585
R142 B.n412 B.n85 585
R143 B.n411 B.n410 585
R144 B.n409 B.n86 585
R145 B.n408 B.n407 585
R146 B.n406 B.n87 585
R147 B.n405 B.n404 585
R148 B.n403 B.n88 585
R149 B.n402 B.n401 585
R150 B.n400 B.n89 585
R151 B.n399 B.n398 585
R152 B.n397 B.n90 585
R153 B.n396 B.n395 585
R154 B.n394 B.n91 585
R155 B.n393 B.n392 585
R156 B.n391 B.n92 585
R157 B.n390 B.n389 585
R158 B.n388 B.n93 585
R159 B.n387 B.n386 585
R160 B.n385 B.n94 585
R161 B.n384 B.n383 585
R162 B.n382 B.n95 585
R163 B.n381 B.n380 585
R164 B.n198 B.n197 585
R165 B.n199 B.n160 585
R166 B.n201 B.n200 585
R167 B.n202 B.n159 585
R168 B.n204 B.n203 585
R169 B.n205 B.n158 585
R170 B.n207 B.n206 585
R171 B.n208 B.n157 585
R172 B.n210 B.n209 585
R173 B.n211 B.n156 585
R174 B.n213 B.n212 585
R175 B.n214 B.n155 585
R176 B.n216 B.n215 585
R177 B.n217 B.n154 585
R178 B.n219 B.n218 585
R179 B.n220 B.n153 585
R180 B.n222 B.n221 585
R181 B.n223 B.n152 585
R182 B.n225 B.n224 585
R183 B.n226 B.n151 585
R184 B.n228 B.n227 585
R185 B.n229 B.n150 585
R186 B.n231 B.n230 585
R187 B.n232 B.n149 585
R188 B.n234 B.n233 585
R189 B.n235 B.n148 585
R190 B.n237 B.n236 585
R191 B.n238 B.n147 585
R192 B.n240 B.n239 585
R193 B.n241 B.n146 585
R194 B.n243 B.n242 585
R195 B.n244 B.n145 585
R196 B.n246 B.n245 585
R197 B.n247 B.n144 585
R198 B.n249 B.n248 585
R199 B.n250 B.n143 585
R200 B.n252 B.n251 585
R201 B.n253 B.n142 585
R202 B.n255 B.n254 585
R203 B.n256 B.n141 585
R204 B.n258 B.n257 585
R205 B.n259 B.n140 585
R206 B.n261 B.n260 585
R207 B.n262 B.n139 585
R208 B.n264 B.n263 585
R209 B.n265 B.n138 585
R210 B.n267 B.n266 585
R211 B.n268 B.n137 585
R212 B.n270 B.n269 585
R213 B.n271 B.n136 585
R214 B.n273 B.n272 585
R215 B.n274 B.n135 585
R216 B.n276 B.n275 585
R217 B.n277 B.n134 585
R218 B.n279 B.n278 585
R219 B.n280 B.n131 585
R220 B.n283 B.n282 585
R221 B.n284 B.n130 585
R222 B.n286 B.n285 585
R223 B.n287 B.n129 585
R224 B.n289 B.n288 585
R225 B.n290 B.n128 585
R226 B.n292 B.n291 585
R227 B.n293 B.n127 585
R228 B.n295 B.n294 585
R229 B.n297 B.n296 585
R230 B.n298 B.n123 585
R231 B.n300 B.n299 585
R232 B.n301 B.n122 585
R233 B.n303 B.n302 585
R234 B.n304 B.n121 585
R235 B.n306 B.n305 585
R236 B.n307 B.n120 585
R237 B.n309 B.n308 585
R238 B.n310 B.n119 585
R239 B.n312 B.n311 585
R240 B.n313 B.n118 585
R241 B.n315 B.n314 585
R242 B.n316 B.n117 585
R243 B.n318 B.n317 585
R244 B.n319 B.n116 585
R245 B.n321 B.n320 585
R246 B.n322 B.n115 585
R247 B.n324 B.n323 585
R248 B.n325 B.n114 585
R249 B.n327 B.n326 585
R250 B.n328 B.n113 585
R251 B.n330 B.n329 585
R252 B.n331 B.n112 585
R253 B.n333 B.n332 585
R254 B.n334 B.n111 585
R255 B.n336 B.n335 585
R256 B.n337 B.n110 585
R257 B.n339 B.n338 585
R258 B.n340 B.n109 585
R259 B.n342 B.n341 585
R260 B.n343 B.n108 585
R261 B.n345 B.n344 585
R262 B.n346 B.n107 585
R263 B.n348 B.n347 585
R264 B.n349 B.n106 585
R265 B.n351 B.n350 585
R266 B.n352 B.n105 585
R267 B.n354 B.n353 585
R268 B.n355 B.n104 585
R269 B.n357 B.n356 585
R270 B.n358 B.n103 585
R271 B.n360 B.n359 585
R272 B.n361 B.n102 585
R273 B.n363 B.n362 585
R274 B.n364 B.n101 585
R275 B.n366 B.n365 585
R276 B.n367 B.n100 585
R277 B.n369 B.n368 585
R278 B.n370 B.n99 585
R279 B.n372 B.n371 585
R280 B.n373 B.n98 585
R281 B.n375 B.n374 585
R282 B.n376 B.n97 585
R283 B.n378 B.n377 585
R284 B.n379 B.n96 585
R285 B.n196 B.n161 585
R286 B.n195 B.n194 585
R287 B.n193 B.n162 585
R288 B.n192 B.n191 585
R289 B.n190 B.n163 585
R290 B.n189 B.n188 585
R291 B.n187 B.n164 585
R292 B.n186 B.n185 585
R293 B.n184 B.n165 585
R294 B.n183 B.n182 585
R295 B.n181 B.n166 585
R296 B.n180 B.n179 585
R297 B.n178 B.n167 585
R298 B.n177 B.n176 585
R299 B.n175 B.n168 585
R300 B.n174 B.n173 585
R301 B.n172 B.n169 585
R302 B.n171 B.n170 585
R303 B.n2 B.n0 585
R304 B.n649 B.n1 585
R305 B.n648 B.n647 585
R306 B.n646 B.n3 585
R307 B.n645 B.n644 585
R308 B.n643 B.n4 585
R309 B.n642 B.n641 585
R310 B.n640 B.n5 585
R311 B.n639 B.n638 585
R312 B.n637 B.n6 585
R313 B.n636 B.n635 585
R314 B.n634 B.n7 585
R315 B.n633 B.n632 585
R316 B.n631 B.n8 585
R317 B.n630 B.n629 585
R318 B.n628 B.n9 585
R319 B.n627 B.n626 585
R320 B.n625 B.n10 585
R321 B.n624 B.n623 585
R322 B.n622 B.n11 585
R323 B.n651 B.n650 585
R324 B.n198 B.n161 497.305
R325 B.n620 B.n11 497.305
R326 B.n380 B.n379 497.305
R327 B.n439 B.n438 497.305
R328 B.n124 B.t5 480.659
R329 B.n46 B.t7 480.659
R330 B.n132 B.t2 480.659
R331 B.n40 B.t10 480.659
R332 B.n125 B.t4 463.01
R333 B.n47 B.t8 463.01
R334 B.n133 B.t1 463.01
R335 B.n41 B.t11 463.01
R336 B.n194 B.n161 163.367
R337 B.n194 B.n193 163.367
R338 B.n193 B.n192 163.367
R339 B.n192 B.n163 163.367
R340 B.n188 B.n163 163.367
R341 B.n188 B.n187 163.367
R342 B.n187 B.n186 163.367
R343 B.n186 B.n165 163.367
R344 B.n182 B.n165 163.367
R345 B.n182 B.n181 163.367
R346 B.n181 B.n180 163.367
R347 B.n180 B.n167 163.367
R348 B.n176 B.n167 163.367
R349 B.n176 B.n175 163.367
R350 B.n175 B.n174 163.367
R351 B.n174 B.n169 163.367
R352 B.n170 B.n169 163.367
R353 B.n170 B.n2 163.367
R354 B.n650 B.n2 163.367
R355 B.n650 B.n649 163.367
R356 B.n649 B.n648 163.367
R357 B.n648 B.n3 163.367
R358 B.n644 B.n3 163.367
R359 B.n644 B.n643 163.367
R360 B.n643 B.n642 163.367
R361 B.n642 B.n5 163.367
R362 B.n638 B.n5 163.367
R363 B.n638 B.n637 163.367
R364 B.n637 B.n636 163.367
R365 B.n636 B.n7 163.367
R366 B.n632 B.n7 163.367
R367 B.n632 B.n631 163.367
R368 B.n631 B.n630 163.367
R369 B.n630 B.n9 163.367
R370 B.n626 B.n9 163.367
R371 B.n626 B.n625 163.367
R372 B.n625 B.n624 163.367
R373 B.n624 B.n11 163.367
R374 B.n199 B.n198 163.367
R375 B.n200 B.n199 163.367
R376 B.n200 B.n159 163.367
R377 B.n204 B.n159 163.367
R378 B.n205 B.n204 163.367
R379 B.n206 B.n205 163.367
R380 B.n206 B.n157 163.367
R381 B.n210 B.n157 163.367
R382 B.n211 B.n210 163.367
R383 B.n212 B.n211 163.367
R384 B.n212 B.n155 163.367
R385 B.n216 B.n155 163.367
R386 B.n217 B.n216 163.367
R387 B.n218 B.n217 163.367
R388 B.n218 B.n153 163.367
R389 B.n222 B.n153 163.367
R390 B.n223 B.n222 163.367
R391 B.n224 B.n223 163.367
R392 B.n224 B.n151 163.367
R393 B.n228 B.n151 163.367
R394 B.n229 B.n228 163.367
R395 B.n230 B.n229 163.367
R396 B.n230 B.n149 163.367
R397 B.n234 B.n149 163.367
R398 B.n235 B.n234 163.367
R399 B.n236 B.n235 163.367
R400 B.n236 B.n147 163.367
R401 B.n240 B.n147 163.367
R402 B.n241 B.n240 163.367
R403 B.n242 B.n241 163.367
R404 B.n242 B.n145 163.367
R405 B.n246 B.n145 163.367
R406 B.n247 B.n246 163.367
R407 B.n248 B.n247 163.367
R408 B.n248 B.n143 163.367
R409 B.n252 B.n143 163.367
R410 B.n253 B.n252 163.367
R411 B.n254 B.n253 163.367
R412 B.n254 B.n141 163.367
R413 B.n258 B.n141 163.367
R414 B.n259 B.n258 163.367
R415 B.n260 B.n259 163.367
R416 B.n260 B.n139 163.367
R417 B.n264 B.n139 163.367
R418 B.n265 B.n264 163.367
R419 B.n266 B.n265 163.367
R420 B.n266 B.n137 163.367
R421 B.n270 B.n137 163.367
R422 B.n271 B.n270 163.367
R423 B.n272 B.n271 163.367
R424 B.n272 B.n135 163.367
R425 B.n276 B.n135 163.367
R426 B.n277 B.n276 163.367
R427 B.n278 B.n277 163.367
R428 B.n278 B.n131 163.367
R429 B.n283 B.n131 163.367
R430 B.n284 B.n283 163.367
R431 B.n285 B.n284 163.367
R432 B.n285 B.n129 163.367
R433 B.n289 B.n129 163.367
R434 B.n290 B.n289 163.367
R435 B.n291 B.n290 163.367
R436 B.n291 B.n127 163.367
R437 B.n295 B.n127 163.367
R438 B.n296 B.n295 163.367
R439 B.n296 B.n123 163.367
R440 B.n300 B.n123 163.367
R441 B.n301 B.n300 163.367
R442 B.n302 B.n301 163.367
R443 B.n302 B.n121 163.367
R444 B.n306 B.n121 163.367
R445 B.n307 B.n306 163.367
R446 B.n308 B.n307 163.367
R447 B.n308 B.n119 163.367
R448 B.n312 B.n119 163.367
R449 B.n313 B.n312 163.367
R450 B.n314 B.n313 163.367
R451 B.n314 B.n117 163.367
R452 B.n318 B.n117 163.367
R453 B.n319 B.n318 163.367
R454 B.n320 B.n319 163.367
R455 B.n320 B.n115 163.367
R456 B.n324 B.n115 163.367
R457 B.n325 B.n324 163.367
R458 B.n326 B.n325 163.367
R459 B.n326 B.n113 163.367
R460 B.n330 B.n113 163.367
R461 B.n331 B.n330 163.367
R462 B.n332 B.n331 163.367
R463 B.n332 B.n111 163.367
R464 B.n336 B.n111 163.367
R465 B.n337 B.n336 163.367
R466 B.n338 B.n337 163.367
R467 B.n338 B.n109 163.367
R468 B.n342 B.n109 163.367
R469 B.n343 B.n342 163.367
R470 B.n344 B.n343 163.367
R471 B.n344 B.n107 163.367
R472 B.n348 B.n107 163.367
R473 B.n349 B.n348 163.367
R474 B.n350 B.n349 163.367
R475 B.n350 B.n105 163.367
R476 B.n354 B.n105 163.367
R477 B.n355 B.n354 163.367
R478 B.n356 B.n355 163.367
R479 B.n356 B.n103 163.367
R480 B.n360 B.n103 163.367
R481 B.n361 B.n360 163.367
R482 B.n362 B.n361 163.367
R483 B.n362 B.n101 163.367
R484 B.n366 B.n101 163.367
R485 B.n367 B.n366 163.367
R486 B.n368 B.n367 163.367
R487 B.n368 B.n99 163.367
R488 B.n372 B.n99 163.367
R489 B.n373 B.n372 163.367
R490 B.n374 B.n373 163.367
R491 B.n374 B.n97 163.367
R492 B.n378 B.n97 163.367
R493 B.n379 B.n378 163.367
R494 B.n380 B.n95 163.367
R495 B.n384 B.n95 163.367
R496 B.n385 B.n384 163.367
R497 B.n386 B.n385 163.367
R498 B.n386 B.n93 163.367
R499 B.n390 B.n93 163.367
R500 B.n391 B.n390 163.367
R501 B.n392 B.n391 163.367
R502 B.n392 B.n91 163.367
R503 B.n396 B.n91 163.367
R504 B.n397 B.n396 163.367
R505 B.n398 B.n397 163.367
R506 B.n398 B.n89 163.367
R507 B.n402 B.n89 163.367
R508 B.n403 B.n402 163.367
R509 B.n404 B.n403 163.367
R510 B.n404 B.n87 163.367
R511 B.n408 B.n87 163.367
R512 B.n409 B.n408 163.367
R513 B.n410 B.n409 163.367
R514 B.n410 B.n85 163.367
R515 B.n414 B.n85 163.367
R516 B.n415 B.n414 163.367
R517 B.n416 B.n415 163.367
R518 B.n416 B.n83 163.367
R519 B.n420 B.n83 163.367
R520 B.n421 B.n420 163.367
R521 B.n422 B.n421 163.367
R522 B.n422 B.n81 163.367
R523 B.n426 B.n81 163.367
R524 B.n427 B.n426 163.367
R525 B.n428 B.n427 163.367
R526 B.n428 B.n79 163.367
R527 B.n432 B.n79 163.367
R528 B.n433 B.n432 163.367
R529 B.n434 B.n433 163.367
R530 B.n434 B.n77 163.367
R531 B.n438 B.n77 163.367
R532 B.n620 B.n619 163.367
R533 B.n619 B.n618 163.367
R534 B.n618 B.n13 163.367
R535 B.n614 B.n13 163.367
R536 B.n614 B.n613 163.367
R537 B.n613 B.n612 163.367
R538 B.n612 B.n15 163.367
R539 B.n608 B.n15 163.367
R540 B.n608 B.n607 163.367
R541 B.n607 B.n606 163.367
R542 B.n606 B.n17 163.367
R543 B.n602 B.n17 163.367
R544 B.n602 B.n601 163.367
R545 B.n601 B.n600 163.367
R546 B.n600 B.n19 163.367
R547 B.n596 B.n19 163.367
R548 B.n596 B.n595 163.367
R549 B.n595 B.n594 163.367
R550 B.n594 B.n21 163.367
R551 B.n590 B.n21 163.367
R552 B.n590 B.n589 163.367
R553 B.n589 B.n588 163.367
R554 B.n588 B.n23 163.367
R555 B.n584 B.n23 163.367
R556 B.n584 B.n583 163.367
R557 B.n583 B.n582 163.367
R558 B.n582 B.n25 163.367
R559 B.n578 B.n25 163.367
R560 B.n578 B.n577 163.367
R561 B.n577 B.n576 163.367
R562 B.n576 B.n27 163.367
R563 B.n572 B.n27 163.367
R564 B.n572 B.n571 163.367
R565 B.n571 B.n570 163.367
R566 B.n570 B.n29 163.367
R567 B.n566 B.n29 163.367
R568 B.n566 B.n565 163.367
R569 B.n565 B.n564 163.367
R570 B.n564 B.n31 163.367
R571 B.n560 B.n31 163.367
R572 B.n560 B.n559 163.367
R573 B.n559 B.n558 163.367
R574 B.n558 B.n33 163.367
R575 B.n554 B.n33 163.367
R576 B.n554 B.n553 163.367
R577 B.n553 B.n552 163.367
R578 B.n552 B.n35 163.367
R579 B.n548 B.n35 163.367
R580 B.n548 B.n547 163.367
R581 B.n547 B.n546 163.367
R582 B.n546 B.n37 163.367
R583 B.n542 B.n37 163.367
R584 B.n542 B.n541 163.367
R585 B.n541 B.n540 163.367
R586 B.n540 B.n39 163.367
R587 B.n535 B.n39 163.367
R588 B.n535 B.n534 163.367
R589 B.n534 B.n533 163.367
R590 B.n533 B.n43 163.367
R591 B.n529 B.n43 163.367
R592 B.n529 B.n528 163.367
R593 B.n528 B.n527 163.367
R594 B.n527 B.n45 163.367
R595 B.n523 B.n45 163.367
R596 B.n523 B.n522 163.367
R597 B.n522 B.n49 163.367
R598 B.n518 B.n49 163.367
R599 B.n518 B.n517 163.367
R600 B.n517 B.n516 163.367
R601 B.n516 B.n51 163.367
R602 B.n512 B.n51 163.367
R603 B.n512 B.n511 163.367
R604 B.n511 B.n510 163.367
R605 B.n510 B.n53 163.367
R606 B.n506 B.n53 163.367
R607 B.n506 B.n505 163.367
R608 B.n505 B.n504 163.367
R609 B.n504 B.n55 163.367
R610 B.n500 B.n55 163.367
R611 B.n500 B.n499 163.367
R612 B.n499 B.n498 163.367
R613 B.n498 B.n57 163.367
R614 B.n494 B.n57 163.367
R615 B.n494 B.n493 163.367
R616 B.n493 B.n492 163.367
R617 B.n492 B.n59 163.367
R618 B.n488 B.n59 163.367
R619 B.n488 B.n487 163.367
R620 B.n487 B.n486 163.367
R621 B.n486 B.n61 163.367
R622 B.n482 B.n61 163.367
R623 B.n482 B.n481 163.367
R624 B.n481 B.n480 163.367
R625 B.n480 B.n63 163.367
R626 B.n476 B.n63 163.367
R627 B.n476 B.n475 163.367
R628 B.n475 B.n474 163.367
R629 B.n474 B.n65 163.367
R630 B.n470 B.n65 163.367
R631 B.n470 B.n469 163.367
R632 B.n469 B.n468 163.367
R633 B.n468 B.n67 163.367
R634 B.n464 B.n67 163.367
R635 B.n464 B.n463 163.367
R636 B.n463 B.n462 163.367
R637 B.n462 B.n69 163.367
R638 B.n458 B.n69 163.367
R639 B.n458 B.n457 163.367
R640 B.n457 B.n456 163.367
R641 B.n456 B.n71 163.367
R642 B.n452 B.n71 163.367
R643 B.n452 B.n451 163.367
R644 B.n451 B.n450 163.367
R645 B.n450 B.n73 163.367
R646 B.n446 B.n73 163.367
R647 B.n446 B.n445 163.367
R648 B.n445 B.n444 163.367
R649 B.n444 B.n75 163.367
R650 B.n440 B.n75 163.367
R651 B.n440 B.n439 163.367
R652 B.n126 B.n125 59.5399
R653 B.n281 B.n133 59.5399
R654 B.n537 B.n41 59.5399
R655 B.n48 B.n47 59.5399
R656 B.n622 B.n621 32.3127
R657 B.n437 B.n76 32.3127
R658 B.n381 B.n96 32.3127
R659 B.n197 B.n196 32.3127
R660 B B.n651 18.0485
R661 B.n125 B.n124 17.649
R662 B.n133 B.n132 17.649
R663 B.n41 B.n40 17.649
R664 B.n47 B.n46 17.649
R665 B.n621 B.n12 10.6151
R666 B.n617 B.n12 10.6151
R667 B.n617 B.n616 10.6151
R668 B.n616 B.n615 10.6151
R669 B.n615 B.n14 10.6151
R670 B.n611 B.n14 10.6151
R671 B.n611 B.n610 10.6151
R672 B.n610 B.n609 10.6151
R673 B.n609 B.n16 10.6151
R674 B.n605 B.n16 10.6151
R675 B.n605 B.n604 10.6151
R676 B.n604 B.n603 10.6151
R677 B.n603 B.n18 10.6151
R678 B.n599 B.n18 10.6151
R679 B.n599 B.n598 10.6151
R680 B.n598 B.n597 10.6151
R681 B.n597 B.n20 10.6151
R682 B.n593 B.n20 10.6151
R683 B.n593 B.n592 10.6151
R684 B.n592 B.n591 10.6151
R685 B.n591 B.n22 10.6151
R686 B.n587 B.n22 10.6151
R687 B.n587 B.n586 10.6151
R688 B.n586 B.n585 10.6151
R689 B.n585 B.n24 10.6151
R690 B.n581 B.n24 10.6151
R691 B.n581 B.n580 10.6151
R692 B.n580 B.n579 10.6151
R693 B.n579 B.n26 10.6151
R694 B.n575 B.n26 10.6151
R695 B.n575 B.n574 10.6151
R696 B.n574 B.n573 10.6151
R697 B.n573 B.n28 10.6151
R698 B.n569 B.n28 10.6151
R699 B.n569 B.n568 10.6151
R700 B.n568 B.n567 10.6151
R701 B.n567 B.n30 10.6151
R702 B.n563 B.n30 10.6151
R703 B.n563 B.n562 10.6151
R704 B.n562 B.n561 10.6151
R705 B.n561 B.n32 10.6151
R706 B.n557 B.n32 10.6151
R707 B.n557 B.n556 10.6151
R708 B.n556 B.n555 10.6151
R709 B.n555 B.n34 10.6151
R710 B.n551 B.n34 10.6151
R711 B.n551 B.n550 10.6151
R712 B.n550 B.n549 10.6151
R713 B.n549 B.n36 10.6151
R714 B.n545 B.n36 10.6151
R715 B.n545 B.n544 10.6151
R716 B.n544 B.n543 10.6151
R717 B.n543 B.n38 10.6151
R718 B.n539 B.n38 10.6151
R719 B.n539 B.n538 10.6151
R720 B.n536 B.n42 10.6151
R721 B.n532 B.n42 10.6151
R722 B.n532 B.n531 10.6151
R723 B.n531 B.n530 10.6151
R724 B.n530 B.n44 10.6151
R725 B.n526 B.n44 10.6151
R726 B.n526 B.n525 10.6151
R727 B.n525 B.n524 10.6151
R728 B.n521 B.n520 10.6151
R729 B.n520 B.n519 10.6151
R730 B.n519 B.n50 10.6151
R731 B.n515 B.n50 10.6151
R732 B.n515 B.n514 10.6151
R733 B.n514 B.n513 10.6151
R734 B.n513 B.n52 10.6151
R735 B.n509 B.n52 10.6151
R736 B.n509 B.n508 10.6151
R737 B.n508 B.n507 10.6151
R738 B.n507 B.n54 10.6151
R739 B.n503 B.n54 10.6151
R740 B.n503 B.n502 10.6151
R741 B.n502 B.n501 10.6151
R742 B.n501 B.n56 10.6151
R743 B.n497 B.n56 10.6151
R744 B.n497 B.n496 10.6151
R745 B.n496 B.n495 10.6151
R746 B.n495 B.n58 10.6151
R747 B.n491 B.n58 10.6151
R748 B.n491 B.n490 10.6151
R749 B.n490 B.n489 10.6151
R750 B.n489 B.n60 10.6151
R751 B.n485 B.n60 10.6151
R752 B.n485 B.n484 10.6151
R753 B.n484 B.n483 10.6151
R754 B.n483 B.n62 10.6151
R755 B.n479 B.n62 10.6151
R756 B.n479 B.n478 10.6151
R757 B.n478 B.n477 10.6151
R758 B.n477 B.n64 10.6151
R759 B.n473 B.n64 10.6151
R760 B.n473 B.n472 10.6151
R761 B.n472 B.n471 10.6151
R762 B.n471 B.n66 10.6151
R763 B.n467 B.n66 10.6151
R764 B.n467 B.n466 10.6151
R765 B.n466 B.n465 10.6151
R766 B.n465 B.n68 10.6151
R767 B.n461 B.n68 10.6151
R768 B.n461 B.n460 10.6151
R769 B.n460 B.n459 10.6151
R770 B.n459 B.n70 10.6151
R771 B.n455 B.n70 10.6151
R772 B.n455 B.n454 10.6151
R773 B.n454 B.n453 10.6151
R774 B.n453 B.n72 10.6151
R775 B.n449 B.n72 10.6151
R776 B.n449 B.n448 10.6151
R777 B.n448 B.n447 10.6151
R778 B.n447 B.n74 10.6151
R779 B.n443 B.n74 10.6151
R780 B.n443 B.n442 10.6151
R781 B.n442 B.n441 10.6151
R782 B.n441 B.n76 10.6151
R783 B.n382 B.n381 10.6151
R784 B.n383 B.n382 10.6151
R785 B.n383 B.n94 10.6151
R786 B.n387 B.n94 10.6151
R787 B.n388 B.n387 10.6151
R788 B.n389 B.n388 10.6151
R789 B.n389 B.n92 10.6151
R790 B.n393 B.n92 10.6151
R791 B.n394 B.n393 10.6151
R792 B.n395 B.n394 10.6151
R793 B.n395 B.n90 10.6151
R794 B.n399 B.n90 10.6151
R795 B.n400 B.n399 10.6151
R796 B.n401 B.n400 10.6151
R797 B.n401 B.n88 10.6151
R798 B.n405 B.n88 10.6151
R799 B.n406 B.n405 10.6151
R800 B.n407 B.n406 10.6151
R801 B.n407 B.n86 10.6151
R802 B.n411 B.n86 10.6151
R803 B.n412 B.n411 10.6151
R804 B.n413 B.n412 10.6151
R805 B.n413 B.n84 10.6151
R806 B.n417 B.n84 10.6151
R807 B.n418 B.n417 10.6151
R808 B.n419 B.n418 10.6151
R809 B.n419 B.n82 10.6151
R810 B.n423 B.n82 10.6151
R811 B.n424 B.n423 10.6151
R812 B.n425 B.n424 10.6151
R813 B.n425 B.n80 10.6151
R814 B.n429 B.n80 10.6151
R815 B.n430 B.n429 10.6151
R816 B.n431 B.n430 10.6151
R817 B.n431 B.n78 10.6151
R818 B.n435 B.n78 10.6151
R819 B.n436 B.n435 10.6151
R820 B.n437 B.n436 10.6151
R821 B.n197 B.n160 10.6151
R822 B.n201 B.n160 10.6151
R823 B.n202 B.n201 10.6151
R824 B.n203 B.n202 10.6151
R825 B.n203 B.n158 10.6151
R826 B.n207 B.n158 10.6151
R827 B.n208 B.n207 10.6151
R828 B.n209 B.n208 10.6151
R829 B.n209 B.n156 10.6151
R830 B.n213 B.n156 10.6151
R831 B.n214 B.n213 10.6151
R832 B.n215 B.n214 10.6151
R833 B.n215 B.n154 10.6151
R834 B.n219 B.n154 10.6151
R835 B.n220 B.n219 10.6151
R836 B.n221 B.n220 10.6151
R837 B.n221 B.n152 10.6151
R838 B.n225 B.n152 10.6151
R839 B.n226 B.n225 10.6151
R840 B.n227 B.n226 10.6151
R841 B.n227 B.n150 10.6151
R842 B.n231 B.n150 10.6151
R843 B.n232 B.n231 10.6151
R844 B.n233 B.n232 10.6151
R845 B.n233 B.n148 10.6151
R846 B.n237 B.n148 10.6151
R847 B.n238 B.n237 10.6151
R848 B.n239 B.n238 10.6151
R849 B.n239 B.n146 10.6151
R850 B.n243 B.n146 10.6151
R851 B.n244 B.n243 10.6151
R852 B.n245 B.n244 10.6151
R853 B.n245 B.n144 10.6151
R854 B.n249 B.n144 10.6151
R855 B.n250 B.n249 10.6151
R856 B.n251 B.n250 10.6151
R857 B.n251 B.n142 10.6151
R858 B.n255 B.n142 10.6151
R859 B.n256 B.n255 10.6151
R860 B.n257 B.n256 10.6151
R861 B.n257 B.n140 10.6151
R862 B.n261 B.n140 10.6151
R863 B.n262 B.n261 10.6151
R864 B.n263 B.n262 10.6151
R865 B.n263 B.n138 10.6151
R866 B.n267 B.n138 10.6151
R867 B.n268 B.n267 10.6151
R868 B.n269 B.n268 10.6151
R869 B.n269 B.n136 10.6151
R870 B.n273 B.n136 10.6151
R871 B.n274 B.n273 10.6151
R872 B.n275 B.n274 10.6151
R873 B.n275 B.n134 10.6151
R874 B.n279 B.n134 10.6151
R875 B.n280 B.n279 10.6151
R876 B.n282 B.n130 10.6151
R877 B.n286 B.n130 10.6151
R878 B.n287 B.n286 10.6151
R879 B.n288 B.n287 10.6151
R880 B.n288 B.n128 10.6151
R881 B.n292 B.n128 10.6151
R882 B.n293 B.n292 10.6151
R883 B.n294 B.n293 10.6151
R884 B.n298 B.n297 10.6151
R885 B.n299 B.n298 10.6151
R886 B.n299 B.n122 10.6151
R887 B.n303 B.n122 10.6151
R888 B.n304 B.n303 10.6151
R889 B.n305 B.n304 10.6151
R890 B.n305 B.n120 10.6151
R891 B.n309 B.n120 10.6151
R892 B.n310 B.n309 10.6151
R893 B.n311 B.n310 10.6151
R894 B.n311 B.n118 10.6151
R895 B.n315 B.n118 10.6151
R896 B.n316 B.n315 10.6151
R897 B.n317 B.n316 10.6151
R898 B.n317 B.n116 10.6151
R899 B.n321 B.n116 10.6151
R900 B.n322 B.n321 10.6151
R901 B.n323 B.n322 10.6151
R902 B.n323 B.n114 10.6151
R903 B.n327 B.n114 10.6151
R904 B.n328 B.n327 10.6151
R905 B.n329 B.n328 10.6151
R906 B.n329 B.n112 10.6151
R907 B.n333 B.n112 10.6151
R908 B.n334 B.n333 10.6151
R909 B.n335 B.n334 10.6151
R910 B.n335 B.n110 10.6151
R911 B.n339 B.n110 10.6151
R912 B.n340 B.n339 10.6151
R913 B.n341 B.n340 10.6151
R914 B.n341 B.n108 10.6151
R915 B.n345 B.n108 10.6151
R916 B.n346 B.n345 10.6151
R917 B.n347 B.n346 10.6151
R918 B.n347 B.n106 10.6151
R919 B.n351 B.n106 10.6151
R920 B.n352 B.n351 10.6151
R921 B.n353 B.n352 10.6151
R922 B.n353 B.n104 10.6151
R923 B.n357 B.n104 10.6151
R924 B.n358 B.n357 10.6151
R925 B.n359 B.n358 10.6151
R926 B.n359 B.n102 10.6151
R927 B.n363 B.n102 10.6151
R928 B.n364 B.n363 10.6151
R929 B.n365 B.n364 10.6151
R930 B.n365 B.n100 10.6151
R931 B.n369 B.n100 10.6151
R932 B.n370 B.n369 10.6151
R933 B.n371 B.n370 10.6151
R934 B.n371 B.n98 10.6151
R935 B.n375 B.n98 10.6151
R936 B.n376 B.n375 10.6151
R937 B.n377 B.n376 10.6151
R938 B.n377 B.n96 10.6151
R939 B.n196 B.n195 10.6151
R940 B.n195 B.n162 10.6151
R941 B.n191 B.n162 10.6151
R942 B.n191 B.n190 10.6151
R943 B.n190 B.n189 10.6151
R944 B.n189 B.n164 10.6151
R945 B.n185 B.n164 10.6151
R946 B.n185 B.n184 10.6151
R947 B.n184 B.n183 10.6151
R948 B.n183 B.n166 10.6151
R949 B.n179 B.n166 10.6151
R950 B.n179 B.n178 10.6151
R951 B.n178 B.n177 10.6151
R952 B.n177 B.n168 10.6151
R953 B.n173 B.n168 10.6151
R954 B.n173 B.n172 10.6151
R955 B.n172 B.n171 10.6151
R956 B.n171 B.n0 10.6151
R957 B.n647 B.n1 10.6151
R958 B.n647 B.n646 10.6151
R959 B.n646 B.n645 10.6151
R960 B.n645 B.n4 10.6151
R961 B.n641 B.n4 10.6151
R962 B.n641 B.n640 10.6151
R963 B.n640 B.n639 10.6151
R964 B.n639 B.n6 10.6151
R965 B.n635 B.n6 10.6151
R966 B.n635 B.n634 10.6151
R967 B.n634 B.n633 10.6151
R968 B.n633 B.n8 10.6151
R969 B.n629 B.n8 10.6151
R970 B.n629 B.n628 10.6151
R971 B.n628 B.n627 10.6151
R972 B.n627 B.n10 10.6151
R973 B.n623 B.n10 10.6151
R974 B.n623 B.n622 10.6151
R975 B.n537 B.n536 6.5566
R976 B.n524 B.n48 6.5566
R977 B.n282 B.n281 6.5566
R978 B.n294 B.n126 6.5566
R979 B.n538 B.n537 4.05904
R980 B.n521 B.n48 4.05904
R981 B.n281 B.n280 4.05904
R982 B.n297 B.n126 4.05904
R983 B.n651 B.n0 2.81026
R984 B.n651 B.n1 2.81026
R985 VP.n1 VP.t4 795.112
R986 VP.n6 VP.t5 768.292
R987 VP.n7 VP.t1 768.292
R988 VP.n8 VP.t3 768.292
R989 VP.n3 VP.t2 768.292
R990 VP.n2 VP.t0 768.292
R991 VP.n9 VP.n8 161.3
R992 VP.n4 VP.n3 161.3
R993 VP.n6 VP.n5 161.3
R994 VP.n7 VP.n0 80.6037
R995 VP.n7 VP.n6 48.2005
R996 VP.n8 VP.n7 48.2005
R997 VP.n3 VP.n2 48.2005
R998 VP.n4 VP.n1 45.1367
R999 VP.n5 VP.n4 44.474
R1000 VP.n2 VP.n1 13.3799
R1001 VP.n5 VP.n0 0.285035
R1002 VP.n9 VP.n0 0.285035
R1003 VP VP.n9 0.0516364
R1004 VDD1.n88 VDD1.n0 756.745
R1005 VDD1.n181 VDD1.n93 756.745
R1006 VDD1.n89 VDD1.n88 585
R1007 VDD1.n87 VDD1.n86 585
R1008 VDD1.n4 VDD1.n3 585
R1009 VDD1.n81 VDD1.n80 585
R1010 VDD1.n79 VDD1.n78 585
R1011 VDD1.n77 VDD1.n7 585
R1012 VDD1.n11 VDD1.n8 585
R1013 VDD1.n72 VDD1.n71 585
R1014 VDD1.n70 VDD1.n69 585
R1015 VDD1.n13 VDD1.n12 585
R1016 VDD1.n64 VDD1.n63 585
R1017 VDD1.n62 VDD1.n61 585
R1018 VDD1.n17 VDD1.n16 585
R1019 VDD1.n56 VDD1.n55 585
R1020 VDD1.n54 VDD1.n53 585
R1021 VDD1.n21 VDD1.n20 585
R1022 VDD1.n48 VDD1.n47 585
R1023 VDD1.n46 VDD1.n45 585
R1024 VDD1.n25 VDD1.n24 585
R1025 VDD1.n40 VDD1.n39 585
R1026 VDD1.n38 VDD1.n37 585
R1027 VDD1.n29 VDD1.n28 585
R1028 VDD1.n32 VDD1.n31 585
R1029 VDD1.n124 VDD1.n123 585
R1030 VDD1.n121 VDD1.n120 585
R1031 VDD1.n130 VDD1.n129 585
R1032 VDD1.n132 VDD1.n131 585
R1033 VDD1.n117 VDD1.n116 585
R1034 VDD1.n138 VDD1.n137 585
R1035 VDD1.n140 VDD1.n139 585
R1036 VDD1.n113 VDD1.n112 585
R1037 VDD1.n146 VDD1.n145 585
R1038 VDD1.n148 VDD1.n147 585
R1039 VDD1.n109 VDD1.n108 585
R1040 VDD1.n154 VDD1.n153 585
R1041 VDD1.n156 VDD1.n155 585
R1042 VDD1.n105 VDD1.n104 585
R1043 VDD1.n162 VDD1.n161 585
R1044 VDD1.n165 VDD1.n164 585
R1045 VDD1.n163 VDD1.n101 585
R1046 VDD1.n170 VDD1.n100 585
R1047 VDD1.n172 VDD1.n171 585
R1048 VDD1.n174 VDD1.n173 585
R1049 VDD1.n97 VDD1.n96 585
R1050 VDD1.n180 VDD1.n179 585
R1051 VDD1.n182 VDD1.n181 585
R1052 VDD1.t0 VDD1.n30 327.466
R1053 VDD1.t1 VDD1.n122 327.466
R1054 VDD1.n88 VDD1.n87 171.744
R1055 VDD1.n87 VDD1.n3 171.744
R1056 VDD1.n80 VDD1.n3 171.744
R1057 VDD1.n80 VDD1.n79 171.744
R1058 VDD1.n79 VDD1.n7 171.744
R1059 VDD1.n11 VDD1.n7 171.744
R1060 VDD1.n71 VDD1.n11 171.744
R1061 VDD1.n71 VDD1.n70 171.744
R1062 VDD1.n70 VDD1.n12 171.744
R1063 VDD1.n63 VDD1.n12 171.744
R1064 VDD1.n63 VDD1.n62 171.744
R1065 VDD1.n62 VDD1.n16 171.744
R1066 VDD1.n55 VDD1.n16 171.744
R1067 VDD1.n55 VDD1.n54 171.744
R1068 VDD1.n54 VDD1.n20 171.744
R1069 VDD1.n47 VDD1.n20 171.744
R1070 VDD1.n47 VDD1.n46 171.744
R1071 VDD1.n46 VDD1.n24 171.744
R1072 VDD1.n39 VDD1.n24 171.744
R1073 VDD1.n39 VDD1.n38 171.744
R1074 VDD1.n38 VDD1.n28 171.744
R1075 VDD1.n31 VDD1.n28 171.744
R1076 VDD1.n123 VDD1.n120 171.744
R1077 VDD1.n130 VDD1.n120 171.744
R1078 VDD1.n131 VDD1.n130 171.744
R1079 VDD1.n131 VDD1.n116 171.744
R1080 VDD1.n138 VDD1.n116 171.744
R1081 VDD1.n139 VDD1.n138 171.744
R1082 VDD1.n139 VDD1.n112 171.744
R1083 VDD1.n146 VDD1.n112 171.744
R1084 VDD1.n147 VDD1.n146 171.744
R1085 VDD1.n147 VDD1.n108 171.744
R1086 VDD1.n154 VDD1.n108 171.744
R1087 VDD1.n155 VDD1.n154 171.744
R1088 VDD1.n155 VDD1.n104 171.744
R1089 VDD1.n162 VDD1.n104 171.744
R1090 VDD1.n164 VDD1.n162 171.744
R1091 VDD1.n164 VDD1.n163 171.744
R1092 VDD1.n163 VDD1.n100 171.744
R1093 VDD1.n172 VDD1.n100 171.744
R1094 VDD1.n173 VDD1.n172 171.744
R1095 VDD1.n173 VDD1.n96 171.744
R1096 VDD1.n180 VDD1.n96 171.744
R1097 VDD1.n181 VDD1.n180 171.744
R1098 VDD1.n31 VDD1.t0 85.8723
R1099 VDD1.n123 VDD1.t1 85.8723
R1100 VDD1.n187 VDD1.n186 70.5023
R1101 VDD1.n189 VDD1.n188 70.3615
R1102 VDD1 VDD1.n92 50.4804
R1103 VDD1.n187 VDD1.n185 50.3668
R1104 VDD1.n189 VDD1.n187 41.766
R1105 VDD1.n32 VDD1.n30 16.3895
R1106 VDD1.n124 VDD1.n122 16.3895
R1107 VDD1.n78 VDD1.n77 13.1884
R1108 VDD1.n171 VDD1.n170 13.1884
R1109 VDD1.n81 VDD1.n6 12.8005
R1110 VDD1.n76 VDD1.n8 12.8005
R1111 VDD1.n33 VDD1.n29 12.8005
R1112 VDD1.n125 VDD1.n121 12.8005
R1113 VDD1.n169 VDD1.n101 12.8005
R1114 VDD1.n174 VDD1.n99 12.8005
R1115 VDD1.n82 VDD1.n4 12.0247
R1116 VDD1.n73 VDD1.n72 12.0247
R1117 VDD1.n37 VDD1.n36 12.0247
R1118 VDD1.n129 VDD1.n128 12.0247
R1119 VDD1.n166 VDD1.n165 12.0247
R1120 VDD1.n175 VDD1.n97 12.0247
R1121 VDD1.n86 VDD1.n85 11.249
R1122 VDD1.n69 VDD1.n10 11.249
R1123 VDD1.n40 VDD1.n27 11.249
R1124 VDD1.n132 VDD1.n119 11.249
R1125 VDD1.n161 VDD1.n103 11.249
R1126 VDD1.n179 VDD1.n178 11.249
R1127 VDD1.n89 VDD1.n2 10.4732
R1128 VDD1.n68 VDD1.n13 10.4732
R1129 VDD1.n41 VDD1.n25 10.4732
R1130 VDD1.n133 VDD1.n117 10.4732
R1131 VDD1.n160 VDD1.n105 10.4732
R1132 VDD1.n182 VDD1.n95 10.4732
R1133 VDD1.n90 VDD1.n0 9.69747
R1134 VDD1.n65 VDD1.n64 9.69747
R1135 VDD1.n45 VDD1.n44 9.69747
R1136 VDD1.n137 VDD1.n136 9.69747
R1137 VDD1.n157 VDD1.n156 9.69747
R1138 VDD1.n183 VDD1.n93 9.69747
R1139 VDD1.n92 VDD1.n91 9.45567
R1140 VDD1.n185 VDD1.n184 9.45567
R1141 VDD1.n58 VDD1.n57 9.3005
R1142 VDD1.n60 VDD1.n59 9.3005
R1143 VDD1.n15 VDD1.n14 9.3005
R1144 VDD1.n66 VDD1.n65 9.3005
R1145 VDD1.n68 VDD1.n67 9.3005
R1146 VDD1.n10 VDD1.n9 9.3005
R1147 VDD1.n74 VDD1.n73 9.3005
R1148 VDD1.n76 VDD1.n75 9.3005
R1149 VDD1.n91 VDD1.n90 9.3005
R1150 VDD1.n2 VDD1.n1 9.3005
R1151 VDD1.n85 VDD1.n84 9.3005
R1152 VDD1.n83 VDD1.n82 9.3005
R1153 VDD1.n6 VDD1.n5 9.3005
R1154 VDD1.n19 VDD1.n18 9.3005
R1155 VDD1.n52 VDD1.n51 9.3005
R1156 VDD1.n50 VDD1.n49 9.3005
R1157 VDD1.n23 VDD1.n22 9.3005
R1158 VDD1.n44 VDD1.n43 9.3005
R1159 VDD1.n42 VDD1.n41 9.3005
R1160 VDD1.n27 VDD1.n26 9.3005
R1161 VDD1.n36 VDD1.n35 9.3005
R1162 VDD1.n34 VDD1.n33 9.3005
R1163 VDD1.n184 VDD1.n183 9.3005
R1164 VDD1.n95 VDD1.n94 9.3005
R1165 VDD1.n178 VDD1.n177 9.3005
R1166 VDD1.n176 VDD1.n175 9.3005
R1167 VDD1.n99 VDD1.n98 9.3005
R1168 VDD1.n144 VDD1.n143 9.3005
R1169 VDD1.n142 VDD1.n141 9.3005
R1170 VDD1.n115 VDD1.n114 9.3005
R1171 VDD1.n136 VDD1.n135 9.3005
R1172 VDD1.n134 VDD1.n133 9.3005
R1173 VDD1.n119 VDD1.n118 9.3005
R1174 VDD1.n128 VDD1.n127 9.3005
R1175 VDD1.n126 VDD1.n125 9.3005
R1176 VDD1.n111 VDD1.n110 9.3005
R1177 VDD1.n150 VDD1.n149 9.3005
R1178 VDD1.n152 VDD1.n151 9.3005
R1179 VDD1.n107 VDD1.n106 9.3005
R1180 VDD1.n158 VDD1.n157 9.3005
R1181 VDD1.n160 VDD1.n159 9.3005
R1182 VDD1.n103 VDD1.n102 9.3005
R1183 VDD1.n167 VDD1.n166 9.3005
R1184 VDD1.n169 VDD1.n168 9.3005
R1185 VDD1.n61 VDD1.n15 8.92171
R1186 VDD1.n48 VDD1.n23 8.92171
R1187 VDD1.n140 VDD1.n115 8.92171
R1188 VDD1.n153 VDD1.n107 8.92171
R1189 VDD1.n60 VDD1.n17 8.14595
R1190 VDD1.n49 VDD1.n21 8.14595
R1191 VDD1.n141 VDD1.n113 8.14595
R1192 VDD1.n152 VDD1.n109 8.14595
R1193 VDD1.n57 VDD1.n56 7.3702
R1194 VDD1.n53 VDD1.n52 7.3702
R1195 VDD1.n145 VDD1.n144 7.3702
R1196 VDD1.n149 VDD1.n148 7.3702
R1197 VDD1.n56 VDD1.n19 6.59444
R1198 VDD1.n53 VDD1.n19 6.59444
R1199 VDD1.n145 VDD1.n111 6.59444
R1200 VDD1.n148 VDD1.n111 6.59444
R1201 VDD1.n57 VDD1.n17 5.81868
R1202 VDD1.n52 VDD1.n21 5.81868
R1203 VDD1.n144 VDD1.n113 5.81868
R1204 VDD1.n149 VDD1.n109 5.81868
R1205 VDD1.n61 VDD1.n60 5.04292
R1206 VDD1.n49 VDD1.n48 5.04292
R1207 VDD1.n141 VDD1.n140 5.04292
R1208 VDD1.n153 VDD1.n152 5.04292
R1209 VDD1.n92 VDD1.n0 4.26717
R1210 VDD1.n64 VDD1.n15 4.26717
R1211 VDD1.n45 VDD1.n23 4.26717
R1212 VDD1.n137 VDD1.n115 4.26717
R1213 VDD1.n156 VDD1.n107 4.26717
R1214 VDD1.n185 VDD1.n93 4.26717
R1215 VDD1.n34 VDD1.n30 3.70982
R1216 VDD1.n126 VDD1.n122 3.70982
R1217 VDD1.n90 VDD1.n89 3.49141
R1218 VDD1.n65 VDD1.n13 3.49141
R1219 VDD1.n44 VDD1.n25 3.49141
R1220 VDD1.n136 VDD1.n117 3.49141
R1221 VDD1.n157 VDD1.n105 3.49141
R1222 VDD1.n183 VDD1.n182 3.49141
R1223 VDD1.n86 VDD1.n2 2.71565
R1224 VDD1.n69 VDD1.n68 2.71565
R1225 VDD1.n41 VDD1.n40 2.71565
R1226 VDD1.n133 VDD1.n132 2.71565
R1227 VDD1.n161 VDD1.n160 2.71565
R1228 VDD1.n179 VDD1.n95 2.71565
R1229 VDD1.n85 VDD1.n4 1.93989
R1230 VDD1.n72 VDD1.n10 1.93989
R1231 VDD1.n37 VDD1.n27 1.93989
R1232 VDD1.n129 VDD1.n119 1.93989
R1233 VDD1.n165 VDD1.n103 1.93989
R1234 VDD1.n178 VDD1.n97 1.93989
R1235 VDD1.n188 VDD1.t3 1.92958
R1236 VDD1.n188 VDD1.t5 1.92958
R1237 VDD1.n186 VDD1.t2 1.92958
R1238 VDD1.n186 VDD1.t4 1.92958
R1239 VDD1.n82 VDD1.n81 1.16414
R1240 VDD1.n73 VDD1.n8 1.16414
R1241 VDD1.n36 VDD1.n29 1.16414
R1242 VDD1.n128 VDD1.n121 1.16414
R1243 VDD1.n166 VDD1.n101 1.16414
R1244 VDD1.n175 VDD1.n174 1.16414
R1245 VDD1.n78 VDD1.n6 0.388379
R1246 VDD1.n77 VDD1.n76 0.388379
R1247 VDD1.n33 VDD1.n32 0.388379
R1248 VDD1.n125 VDD1.n124 0.388379
R1249 VDD1.n170 VDD1.n169 0.388379
R1250 VDD1.n171 VDD1.n99 0.388379
R1251 VDD1.n91 VDD1.n1 0.155672
R1252 VDD1.n84 VDD1.n1 0.155672
R1253 VDD1.n84 VDD1.n83 0.155672
R1254 VDD1.n83 VDD1.n5 0.155672
R1255 VDD1.n75 VDD1.n5 0.155672
R1256 VDD1.n75 VDD1.n74 0.155672
R1257 VDD1.n74 VDD1.n9 0.155672
R1258 VDD1.n67 VDD1.n9 0.155672
R1259 VDD1.n67 VDD1.n66 0.155672
R1260 VDD1.n66 VDD1.n14 0.155672
R1261 VDD1.n59 VDD1.n14 0.155672
R1262 VDD1.n59 VDD1.n58 0.155672
R1263 VDD1.n58 VDD1.n18 0.155672
R1264 VDD1.n51 VDD1.n18 0.155672
R1265 VDD1.n51 VDD1.n50 0.155672
R1266 VDD1.n50 VDD1.n22 0.155672
R1267 VDD1.n43 VDD1.n22 0.155672
R1268 VDD1.n43 VDD1.n42 0.155672
R1269 VDD1.n42 VDD1.n26 0.155672
R1270 VDD1.n35 VDD1.n26 0.155672
R1271 VDD1.n35 VDD1.n34 0.155672
R1272 VDD1.n127 VDD1.n126 0.155672
R1273 VDD1.n127 VDD1.n118 0.155672
R1274 VDD1.n134 VDD1.n118 0.155672
R1275 VDD1.n135 VDD1.n134 0.155672
R1276 VDD1.n135 VDD1.n114 0.155672
R1277 VDD1.n142 VDD1.n114 0.155672
R1278 VDD1.n143 VDD1.n142 0.155672
R1279 VDD1.n143 VDD1.n110 0.155672
R1280 VDD1.n150 VDD1.n110 0.155672
R1281 VDD1.n151 VDD1.n150 0.155672
R1282 VDD1.n151 VDD1.n106 0.155672
R1283 VDD1.n158 VDD1.n106 0.155672
R1284 VDD1.n159 VDD1.n158 0.155672
R1285 VDD1.n159 VDD1.n102 0.155672
R1286 VDD1.n167 VDD1.n102 0.155672
R1287 VDD1.n168 VDD1.n167 0.155672
R1288 VDD1.n168 VDD1.n98 0.155672
R1289 VDD1.n176 VDD1.n98 0.155672
R1290 VDD1.n177 VDD1.n176 0.155672
R1291 VDD1.n177 VDD1.n94 0.155672
R1292 VDD1.n184 VDD1.n94 0.155672
R1293 VDD1 VDD1.n189 0.138431
R1294 VTAIL.n378 VTAIL.n290 756.745
R1295 VTAIL.n90 VTAIL.n2 756.745
R1296 VTAIL.n284 VTAIL.n196 756.745
R1297 VTAIL.n188 VTAIL.n100 756.745
R1298 VTAIL.n321 VTAIL.n320 585
R1299 VTAIL.n318 VTAIL.n317 585
R1300 VTAIL.n327 VTAIL.n326 585
R1301 VTAIL.n329 VTAIL.n328 585
R1302 VTAIL.n314 VTAIL.n313 585
R1303 VTAIL.n335 VTAIL.n334 585
R1304 VTAIL.n337 VTAIL.n336 585
R1305 VTAIL.n310 VTAIL.n309 585
R1306 VTAIL.n343 VTAIL.n342 585
R1307 VTAIL.n345 VTAIL.n344 585
R1308 VTAIL.n306 VTAIL.n305 585
R1309 VTAIL.n351 VTAIL.n350 585
R1310 VTAIL.n353 VTAIL.n352 585
R1311 VTAIL.n302 VTAIL.n301 585
R1312 VTAIL.n359 VTAIL.n358 585
R1313 VTAIL.n362 VTAIL.n361 585
R1314 VTAIL.n360 VTAIL.n298 585
R1315 VTAIL.n367 VTAIL.n297 585
R1316 VTAIL.n369 VTAIL.n368 585
R1317 VTAIL.n371 VTAIL.n370 585
R1318 VTAIL.n294 VTAIL.n293 585
R1319 VTAIL.n377 VTAIL.n376 585
R1320 VTAIL.n379 VTAIL.n378 585
R1321 VTAIL.n33 VTAIL.n32 585
R1322 VTAIL.n30 VTAIL.n29 585
R1323 VTAIL.n39 VTAIL.n38 585
R1324 VTAIL.n41 VTAIL.n40 585
R1325 VTAIL.n26 VTAIL.n25 585
R1326 VTAIL.n47 VTAIL.n46 585
R1327 VTAIL.n49 VTAIL.n48 585
R1328 VTAIL.n22 VTAIL.n21 585
R1329 VTAIL.n55 VTAIL.n54 585
R1330 VTAIL.n57 VTAIL.n56 585
R1331 VTAIL.n18 VTAIL.n17 585
R1332 VTAIL.n63 VTAIL.n62 585
R1333 VTAIL.n65 VTAIL.n64 585
R1334 VTAIL.n14 VTAIL.n13 585
R1335 VTAIL.n71 VTAIL.n70 585
R1336 VTAIL.n74 VTAIL.n73 585
R1337 VTAIL.n72 VTAIL.n10 585
R1338 VTAIL.n79 VTAIL.n9 585
R1339 VTAIL.n81 VTAIL.n80 585
R1340 VTAIL.n83 VTAIL.n82 585
R1341 VTAIL.n6 VTAIL.n5 585
R1342 VTAIL.n89 VTAIL.n88 585
R1343 VTAIL.n91 VTAIL.n90 585
R1344 VTAIL.n285 VTAIL.n284 585
R1345 VTAIL.n283 VTAIL.n282 585
R1346 VTAIL.n200 VTAIL.n199 585
R1347 VTAIL.n277 VTAIL.n276 585
R1348 VTAIL.n275 VTAIL.n274 585
R1349 VTAIL.n273 VTAIL.n203 585
R1350 VTAIL.n207 VTAIL.n204 585
R1351 VTAIL.n268 VTAIL.n267 585
R1352 VTAIL.n266 VTAIL.n265 585
R1353 VTAIL.n209 VTAIL.n208 585
R1354 VTAIL.n260 VTAIL.n259 585
R1355 VTAIL.n258 VTAIL.n257 585
R1356 VTAIL.n213 VTAIL.n212 585
R1357 VTAIL.n252 VTAIL.n251 585
R1358 VTAIL.n250 VTAIL.n249 585
R1359 VTAIL.n217 VTAIL.n216 585
R1360 VTAIL.n244 VTAIL.n243 585
R1361 VTAIL.n242 VTAIL.n241 585
R1362 VTAIL.n221 VTAIL.n220 585
R1363 VTAIL.n236 VTAIL.n235 585
R1364 VTAIL.n234 VTAIL.n233 585
R1365 VTAIL.n225 VTAIL.n224 585
R1366 VTAIL.n228 VTAIL.n227 585
R1367 VTAIL.n189 VTAIL.n188 585
R1368 VTAIL.n187 VTAIL.n186 585
R1369 VTAIL.n104 VTAIL.n103 585
R1370 VTAIL.n181 VTAIL.n180 585
R1371 VTAIL.n179 VTAIL.n178 585
R1372 VTAIL.n177 VTAIL.n107 585
R1373 VTAIL.n111 VTAIL.n108 585
R1374 VTAIL.n172 VTAIL.n171 585
R1375 VTAIL.n170 VTAIL.n169 585
R1376 VTAIL.n113 VTAIL.n112 585
R1377 VTAIL.n164 VTAIL.n163 585
R1378 VTAIL.n162 VTAIL.n161 585
R1379 VTAIL.n117 VTAIL.n116 585
R1380 VTAIL.n156 VTAIL.n155 585
R1381 VTAIL.n154 VTAIL.n153 585
R1382 VTAIL.n121 VTAIL.n120 585
R1383 VTAIL.n148 VTAIL.n147 585
R1384 VTAIL.n146 VTAIL.n145 585
R1385 VTAIL.n125 VTAIL.n124 585
R1386 VTAIL.n140 VTAIL.n139 585
R1387 VTAIL.n138 VTAIL.n137 585
R1388 VTAIL.n129 VTAIL.n128 585
R1389 VTAIL.n132 VTAIL.n131 585
R1390 VTAIL.t9 VTAIL.n226 327.466
R1391 VTAIL.t3 VTAIL.n130 327.466
R1392 VTAIL.t0 VTAIL.n319 327.466
R1393 VTAIL.t8 VTAIL.n31 327.466
R1394 VTAIL.n320 VTAIL.n317 171.744
R1395 VTAIL.n327 VTAIL.n317 171.744
R1396 VTAIL.n328 VTAIL.n327 171.744
R1397 VTAIL.n328 VTAIL.n313 171.744
R1398 VTAIL.n335 VTAIL.n313 171.744
R1399 VTAIL.n336 VTAIL.n335 171.744
R1400 VTAIL.n336 VTAIL.n309 171.744
R1401 VTAIL.n343 VTAIL.n309 171.744
R1402 VTAIL.n344 VTAIL.n343 171.744
R1403 VTAIL.n344 VTAIL.n305 171.744
R1404 VTAIL.n351 VTAIL.n305 171.744
R1405 VTAIL.n352 VTAIL.n351 171.744
R1406 VTAIL.n352 VTAIL.n301 171.744
R1407 VTAIL.n359 VTAIL.n301 171.744
R1408 VTAIL.n361 VTAIL.n359 171.744
R1409 VTAIL.n361 VTAIL.n360 171.744
R1410 VTAIL.n360 VTAIL.n297 171.744
R1411 VTAIL.n369 VTAIL.n297 171.744
R1412 VTAIL.n370 VTAIL.n369 171.744
R1413 VTAIL.n370 VTAIL.n293 171.744
R1414 VTAIL.n377 VTAIL.n293 171.744
R1415 VTAIL.n378 VTAIL.n377 171.744
R1416 VTAIL.n32 VTAIL.n29 171.744
R1417 VTAIL.n39 VTAIL.n29 171.744
R1418 VTAIL.n40 VTAIL.n39 171.744
R1419 VTAIL.n40 VTAIL.n25 171.744
R1420 VTAIL.n47 VTAIL.n25 171.744
R1421 VTAIL.n48 VTAIL.n47 171.744
R1422 VTAIL.n48 VTAIL.n21 171.744
R1423 VTAIL.n55 VTAIL.n21 171.744
R1424 VTAIL.n56 VTAIL.n55 171.744
R1425 VTAIL.n56 VTAIL.n17 171.744
R1426 VTAIL.n63 VTAIL.n17 171.744
R1427 VTAIL.n64 VTAIL.n63 171.744
R1428 VTAIL.n64 VTAIL.n13 171.744
R1429 VTAIL.n71 VTAIL.n13 171.744
R1430 VTAIL.n73 VTAIL.n71 171.744
R1431 VTAIL.n73 VTAIL.n72 171.744
R1432 VTAIL.n72 VTAIL.n9 171.744
R1433 VTAIL.n81 VTAIL.n9 171.744
R1434 VTAIL.n82 VTAIL.n81 171.744
R1435 VTAIL.n82 VTAIL.n5 171.744
R1436 VTAIL.n89 VTAIL.n5 171.744
R1437 VTAIL.n90 VTAIL.n89 171.744
R1438 VTAIL.n284 VTAIL.n283 171.744
R1439 VTAIL.n283 VTAIL.n199 171.744
R1440 VTAIL.n276 VTAIL.n199 171.744
R1441 VTAIL.n276 VTAIL.n275 171.744
R1442 VTAIL.n275 VTAIL.n203 171.744
R1443 VTAIL.n207 VTAIL.n203 171.744
R1444 VTAIL.n267 VTAIL.n207 171.744
R1445 VTAIL.n267 VTAIL.n266 171.744
R1446 VTAIL.n266 VTAIL.n208 171.744
R1447 VTAIL.n259 VTAIL.n208 171.744
R1448 VTAIL.n259 VTAIL.n258 171.744
R1449 VTAIL.n258 VTAIL.n212 171.744
R1450 VTAIL.n251 VTAIL.n212 171.744
R1451 VTAIL.n251 VTAIL.n250 171.744
R1452 VTAIL.n250 VTAIL.n216 171.744
R1453 VTAIL.n243 VTAIL.n216 171.744
R1454 VTAIL.n243 VTAIL.n242 171.744
R1455 VTAIL.n242 VTAIL.n220 171.744
R1456 VTAIL.n235 VTAIL.n220 171.744
R1457 VTAIL.n235 VTAIL.n234 171.744
R1458 VTAIL.n234 VTAIL.n224 171.744
R1459 VTAIL.n227 VTAIL.n224 171.744
R1460 VTAIL.n188 VTAIL.n187 171.744
R1461 VTAIL.n187 VTAIL.n103 171.744
R1462 VTAIL.n180 VTAIL.n103 171.744
R1463 VTAIL.n180 VTAIL.n179 171.744
R1464 VTAIL.n179 VTAIL.n107 171.744
R1465 VTAIL.n111 VTAIL.n107 171.744
R1466 VTAIL.n171 VTAIL.n111 171.744
R1467 VTAIL.n171 VTAIL.n170 171.744
R1468 VTAIL.n170 VTAIL.n112 171.744
R1469 VTAIL.n163 VTAIL.n112 171.744
R1470 VTAIL.n163 VTAIL.n162 171.744
R1471 VTAIL.n162 VTAIL.n116 171.744
R1472 VTAIL.n155 VTAIL.n116 171.744
R1473 VTAIL.n155 VTAIL.n154 171.744
R1474 VTAIL.n154 VTAIL.n120 171.744
R1475 VTAIL.n147 VTAIL.n120 171.744
R1476 VTAIL.n147 VTAIL.n146 171.744
R1477 VTAIL.n146 VTAIL.n124 171.744
R1478 VTAIL.n139 VTAIL.n124 171.744
R1479 VTAIL.n139 VTAIL.n138 171.744
R1480 VTAIL.n138 VTAIL.n128 171.744
R1481 VTAIL.n131 VTAIL.n128 171.744
R1482 VTAIL.n320 VTAIL.t0 85.8723
R1483 VTAIL.n32 VTAIL.t8 85.8723
R1484 VTAIL.n227 VTAIL.t9 85.8723
R1485 VTAIL.n131 VTAIL.t3 85.8723
R1486 VTAIL.n195 VTAIL.n194 53.683
R1487 VTAIL.n99 VTAIL.n98 53.683
R1488 VTAIL.n1 VTAIL.n0 53.6828
R1489 VTAIL.n97 VTAIL.n96 53.6828
R1490 VTAIL.n383 VTAIL.n382 33.155
R1491 VTAIL.n95 VTAIL.n94 33.155
R1492 VTAIL.n289 VTAIL.n288 33.155
R1493 VTAIL.n193 VTAIL.n192 33.155
R1494 VTAIL.n99 VTAIL.n97 28.4617
R1495 VTAIL.n383 VTAIL.n289 27.6772
R1496 VTAIL.n321 VTAIL.n319 16.3895
R1497 VTAIL.n33 VTAIL.n31 16.3895
R1498 VTAIL.n228 VTAIL.n226 16.3895
R1499 VTAIL.n132 VTAIL.n130 16.3895
R1500 VTAIL.n368 VTAIL.n367 13.1884
R1501 VTAIL.n80 VTAIL.n79 13.1884
R1502 VTAIL.n274 VTAIL.n273 13.1884
R1503 VTAIL.n178 VTAIL.n177 13.1884
R1504 VTAIL.n322 VTAIL.n318 12.8005
R1505 VTAIL.n366 VTAIL.n298 12.8005
R1506 VTAIL.n371 VTAIL.n296 12.8005
R1507 VTAIL.n34 VTAIL.n30 12.8005
R1508 VTAIL.n78 VTAIL.n10 12.8005
R1509 VTAIL.n83 VTAIL.n8 12.8005
R1510 VTAIL.n277 VTAIL.n202 12.8005
R1511 VTAIL.n272 VTAIL.n204 12.8005
R1512 VTAIL.n229 VTAIL.n225 12.8005
R1513 VTAIL.n181 VTAIL.n106 12.8005
R1514 VTAIL.n176 VTAIL.n108 12.8005
R1515 VTAIL.n133 VTAIL.n129 12.8005
R1516 VTAIL.n326 VTAIL.n325 12.0247
R1517 VTAIL.n363 VTAIL.n362 12.0247
R1518 VTAIL.n372 VTAIL.n294 12.0247
R1519 VTAIL.n38 VTAIL.n37 12.0247
R1520 VTAIL.n75 VTAIL.n74 12.0247
R1521 VTAIL.n84 VTAIL.n6 12.0247
R1522 VTAIL.n278 VTAIL.n200 12.0247
R1523 VTAIL.n269 VTAIL.n268 12.0247
R1524 VTAIL.n233 VTAIL.n232 12.0247
R1525 VTAIL.n182 VTAIL.n104 12.0247
R1526 VTAIL.n173 VTAIL.n172 12.0247
R1527 VTAIL.n137 VTAIL.n136 12.0247
R1528 VTAIL.n329 VTAIL.n316 11.249
R1529 VTAIL.n358 VTAIL.n300 11.249
R1530 VTAIL.n376 VTAIL.n375 11.249
R1531 VTAIL.n41 VTAIL.n28 11.249
R1532 VTAIL.n70 VTAIL.n12 11.249
R1533 VTAIL.n88 VTAIL.n87 11.249
R1534 VTAIL.n282 VTAIL.n281 11.249
R1535 VTAIL.n265 VTAIL.n206 11.249
R1536 VTAIL.n236 VTAIL.n223 11.249
R1537 VTAIL.n186 VTAIL.n185 11.249
R1538 VTAIL.n169 VTAIL.n110 11.249
R1539 VTAIL.n140 VTAIL.n127 11.249
R1540 VTAIL.n330 VTAIL.n314 10.4732
R1541 VTAIL.n357 VTAIL.n302 10.4732
R1542 VTAIL.n379 VTAIL.n292 10.4732
R1543 VTAIL.n42 VTAIL.n26 10.4732
R1544 VTAIL.n69 VTAIL.n14 10.4732
R1545 VTAIL.n91 VTAIL.n4 10.4732
R1546 VTAIL.n285 VTAIL.n198 10.4732
R1547 VTAIL.n264 VTAIL.n209 10.4732
R1548 VTAIL.n237 VTAIL.n221 10.4732
R1549 VTAIL.n189 VTAIL.n102 10.4732
R1550 VTAIL.n168 VTAIL.n113 10.4732
R1551 VTAIL.n141 VTAIL.n125 10.4732
R1552 VTAIL.n334 VTAIL.n333 9.69747
R1553 VTAIL.n354 VTAIL.n353 9.69747
R1554 VTAIL.n380 VTAIL.n290 9.69747
R1555 VTAIL.n46 VTAIL.n45 9.69747
R1556 VTAIL.n66 VTAIL.n65 9.69747
R1557 VTAIL.n92 VTAIL.n2 9.69747
R1558 VTAIL.n286 VTAIL.n196 9.69747
R1559 VTAIL.n261 VTAIL.n260 9.69747
R1560 VTAIL.n241 VTAIL.n240 9.69747
R1561 VTAIL.n190 VTAIL.n100 9.69747
R1562 VTAIL.n165 VTAIL.n164 9.69747
R1563 VTAIL.n145 VTAIL.n144 9.69747
R1564 VTAIL.n382 VTAIL.n381 9.45567
R1565 VTAIL.n94 VTAIL.n93 9.45567
R1566 VTAIL.n288 VTAIL.n287 9.45567
R1567 VTAIL.n192 VTAIL.n191 9.45567
R1568 VTAIL.n381 VTAIL.n380 9.3005
R1569 VTAIL.n292 VTAIL.n291 9.3005
R1570 VTAIL.n375 VTAIL.n374 9.3005
R1571 VTAIL.n373 VTAIL.n372 9.3005
R1572 VTAIL.n296 VTAIL.n295 9.3005
R1573 VTAIL.n341 VTAIL.n340 9.3005
R1574 VTAIL.n339 VTAIL.n338 9.3005
R1575 VTAIL.n312 VTAIL.n311 9.3005
R1576 VTAIL.n333 VTAIL.n332 9.3005
R1577 VTAIL.n331 VTAIL.n330 9.3005
R1578 VTAIL.n316 VTAIL.n315 9.3005
R1579 VTAIL.n325 VTAIL.n324 9.3005
R1580 VTAIL.n323 VTAIL.n322 9.3005
R1581 VTAIL.n308 VTAIL.n307 9.3005
R1582 VTAIL.n347 VTAIL.n346 9.3005
R1583 VTAIL.n349 VTAIL.n348 9.3005
R1584 VTAIL.n304 VTAIL.n303 9.3005
R1585 VTAIL.n355 VTAIL.n354 9.3005
R1586 VTAIL.n357 VTAIL.n356 9.3005
R1587 VTAIL.n300 VTAIL.n299 9.3005
R1588 VTAIL.n364 VTAIL.n363 9.3005
R1589 VTAIL.n366 VTAIL.n365 9.3005
R1590 VTAIL.n93 VTAIL.n92 9.3005
R1591 VTAIL.n4 VTAIL.n3 9.3005
R1592 VTAIL.n87 VTAIL.n86 9.3005
R1593 VTAIL.n85 VTAIL.n84 9.3005
R1594 VTAIL.n8 VTAIL.n7 9.3005
R1595 VTAIL.n53 VTAIL.n52 9.3005
R1596 VTAIL.n51 VTAIL.n50 9.3005
R1597 VTAIL.n24 VTAIL.n23 9.3005
R1598 VTAIL.n45 VTAIL.n44 9.3005
R1599 VTAIL.n43 VTAIL.n42 9.3005
R1600 VTAIL.n28 VTAIL.n27 9.3005
R1601 VTAIL.n37 VTAIL.n36 9.3005
R1602 VTAIL.n35 VTAIL.n34 9.3005
R1603 VTAIL.n20 VTAIL.n19 9.3005
R1604 VTAIL.n59 VTAIL.n58 9.3005
R1605 VTAIL.n61 VTAIL.n60 9.3005
R1606 VTAIL.n16 VTAIL.n15 9.3005
R1607 VTAIL.n67 VTAIL.n66 9.3005
R1608 VTAIL.n69 VTAIL.n68 9.3005
R1609 VTAIL.n12 VTAIL.n11 9.3005
R1610 VTAIL.n76 VTAIL.n75 9.3005
R1611 VTAIL.n78 VTAIL.n77 9.3005
R1612 VTAIL.n254 VTAIL.n253 9.3005
R1613 VTAIL.n256 VTAIL.n255 9.3005
R1614 VTAIL.n211 VTAIL.n210 9.3005
R1615 VTAIL.n262 VTAIL.n261 9.3005
R1616 VTAIL.n264 VTAIL.n263 9.3005
R1617 VTAIL.n206 VTAIL.n205 9.3005
R1618 VTAIL.n270 VTAIL.n269 9.3005
R1619 VTAIL.n272 VTAIL.n271 9.3005
R1620 VTAIL.n287 VTAIL.n286 9.3005
R1621 VTAIL.n198 VTAIL.n197 9.3005
R1622 VTAIL.n281 VTAIL.n280 9.3005
R1623 VTAIL.n279 VTAIL.n278 9.3005
R1624 VTAIL.n202 VTAIL.n201 9.3005
R1625 VTAIL.n215 VTAIL.n214 9.3005
R1626 VTAIL.n248 VTAIL.n247 9.3005
R1627 VTAIL.n246 VTAIL.n245 9.3005
R1628 VTAIL.n219 VTAIL.n218 9.3005
R1629 VTAIL.n240 VTAIL.n239 9.3005
R1630 VTAIL.n238 VTAIL.n237 9.3005
R1631 VTAIL.n223 VTAIL.n222 9.3005
R1632 VTAIL.n232 VTAIL.n231 9.3005
R1633 VTAIL.n230 VTAIL.n229 9.3005
R1634 VTAIL.n158 VTAIL.n157 9.3005
R1635 VTAIL.n160 VTAIL.n159 9.3005
R1636 VTAIL.n115 VTAIL.n114 9.3005
R1637 VTAIL.n166 VTAIL.n165 9.3005
R1638 VTAIL.n168 VTAIL.n167 9.3005
R1639 VTAIL.n110 VTAIL.n109 9.3005
R1640 VTAIL.n174 VTAIL.n173 9.3005
R1641 VTAIL.n176 VTAIL.n175 9.3005
R1642 VTAIL.n191 VTAIL.n190 9.3005
R1643 VTAIL.n102 VTAIL.n101 9.3005
R1644 VTAIL.n185 VTAIL.n184 9.3005
R1645 VTAIL.n183 VTAIL.n182 9.3005
R1646 VTAIL.n106 VTAIL.n105 9.3005
R1647 VTAIL.n119 VTAIL.n118 9.3005
R1648 VTAIL.n152 VTAIL.n151 9.3005
R1649 VTAIL.n150 VTAIL.n149 9.3005
R1650 VTAIL.n123 VTAIL.n122 9.3005
R1651 VTAIL.n144 VTAIL.n143 9.3005
R1652 VTAIL.n142 VTAIL.n141 9.3005
R1653 VTAIL.n127 VTAIL.n126 9.3005
R1654 VTAIL.n136 VTAIL.n135 9.3005
R1655 VTAIL.n134 VTAIL.n133 9.3005
R1656 VTAIL.n337 VTAIL.n312 8.92171
R1657 VTAIL.n350 VTAIL.n304 8.92171
R1658 VTAIL.n49 VTAIL.n24 8.92171
R1659 VTAIL.n62 VTAIL.n16 8.92171
R1660 VTAIL.n257 VTAIL.n211 8.92171
R1661 VTAIL.n244 VTAIL.n219 8.92171
R1662 VTAIL.n161 VTAIL.n115 8.92171
R1663 VTAIL.n148 VTAIL.n123 8.92171
R1664 VTAIL.n338 VTAIL.n310 8.14595
R1665 VTAIL.n349 VTAIL.n306 8.14595
R1666 VTAIL.n50 VTAIL.n22 8.14595
R1667 VTAIL.n61 VTAIL.n18 8.14595
R1668 VTAIL.n256 VTAIL.n213 8.14595
R1669 VTAIL.n245 VTAIL.n217 8.14595
R1670 VTAIL.n160 VTAIL.n117 8.14595
R1671 VTAIL.n149 VTAIL.n121 8.14595
R1672 VTAIL.n342 VTAIL.n341 7.3702
R1673 VTAIL.n346 VTAIL.n345 7.3702
R1674 VTAIL.n54 VTAIL.n53 7.3702
R1675 VTAIL.n58 VTAIL.n57 7.3702
R1676 VTAIL.n253 VTAIL.n252 7.3702
R1677 VTAIL.n249 VTAIL.n248 7.3702
R1678 VTAIL.n157 VTAIL.n156 7.3702
R1679 VTAIL.n153 VTAIL.n152 7.3702
R1680 VTAIL.n342 VTAIL.n308 6.59444
R1681 VTAIL.n345 VTAIL.n308 6.59444
R1682 VTAIL.n54 VTAIL.n20 6.59444
R1683 VTAIL.n57 VTAIL.n20 6.59444
R1684 VTAIL.n252 VTAIL.n215 6.59444
R1685 VTAIL.n249 VTAIL.n215 6.59444
R1686 VTAIL.n156 VTAIL.n119 6.59444
R1687 VTAIL.n153 VTAIL.n119 6.59444
R1688 VTAIL.n341 VTAIL.n310 5.81868
R1689 VTAIL.n346 VTAIL.n306 5.81868
R1690 VTAIL.n53 VTAIL.n22 5.81868
R1691 VTAIL.n58 VTAIL.n18 5.81868
R1692 VTAIL.n253 VTAIL.n213 5.81868
R1693 VTAIL.n248 VTAIL.n217 5.81868
R1694 VTAIL.n157 VTAIL.n117 5.81868
R1695 VTAIL.n152 VTAIL.n121 5.81868
R1696 VTAIL.n338 VTAIL.n337 5.04292
R1697 VTAIL.n350 VTAIL.n349 5.04292
R1698 VTAIL.n50 VTAIL.n49 5.04292
R1699 VTAIL.n62 VTAIL.n61 5.04292
R1700 VTAIL.n257 VTAIL.n256 5.04292
R1701 VTAIL.n245 VTAIL.n244 5.04292
R1702 VTAIL.n161 VTAIL.n160 5.04292
R1703 VTAIL.n149 VTAIL.n148 5.04292
R1704 VTAIL.n334 VTAIL.n312 4.26717
R1705 VTAIL.n353 VTAIL.n304 4.26717
R1706 VTAIL.n382 VTAIL.n290 4.26717
R1707 VTAIL.n46 VTAIL.n24 4.26717
R1708 VTAIL.n65 VTAIL.n16 4.26717
R1709 VTAIL.n94 VTAIL.n2 4.26717
R1710 VTAIL.n288 VTAIL.n196 4.26717
R1711 VTAIL.n260 VTAIL.n211 4.26717
R1712 VTAIL.n241 VTAIL.n219 4.26717
R1713 VTAIL.n192 VTAIL.n100 4.26717
R1714 VTAIL.n164 VTAIL.n115 4.26717
R1715 VTAIL.n145 VTAIL.n123 4.26717
R1716 VTAIL.n323 VTAIL.n319 3.70982
R1717 VTAIL.n35 VTAIL.n31 3.70982
R1718 VTAIL.n230 VTAIL.n226 3.70982
R1719 VTAIL.n134 VTAIL.n130 3.70982
R1720 VTAIL.n333 VTAIL.n314 3.49141
R1721 VTAIL.n354 VTAIL.n302 3.49141
R1722 VTAIL.n380 VTAIL.n379 3.49141
R1723 VTAIL.n45 VTAIL.n26 3.49141
R1724 VTAIL.n66 VTAIL.n14 3.49141
R1725 VTAIL.n92 VTAIL.n91 3.49141
R1726 VTAIL.n286 VTAIL.n285 3.49141
R1727 VTAIL.n261 VTAIL.n209 3.49141
R1728 VTAIL.n240 VTAIL.n221 3.49141
R1729 VTAIL.n190 VTAIL.n189 3.49141
R1730 VTAIL.n165 VTAIL.n113 3.49141
R1731 VTAIL.n144 VTAIL.n125 3.49141
R1732 VTAIL.n330 VTAIL.n329 2.71565
R1733 VTAIL.n358 VTAIL.n357 2.71565
R1734 VTAIL.n376 VTAIL.n292 2.71565
R1735 VTAIL.n42 VTAIL.n41 2.71565
R1736 VTAIL.n70 VTAIL.n69 2.71565
R1737 VTAIL.n88 VTAIL.n4 2.71565
R1738 VTAIL.n282 VTAIL.n198 2.71565
R1739 VTAIL.n265 VTAIL.n264 2.71565
R1740 VTAIL.n237 VTAIL.n236 2.71565
R1741 VTAIL.n186 VTAIL.n102 2.71565
R1742 VTAIL.n169 VTAIL.n168 2.71565
R1743 VTAIL.n141 VTAIL.n140 2.71565
R1744 VTAIL.n326 VTAIL.n316 1.93989
R1745 VTAIL.n362 VTAIL.n300 1.93989
R1746 VTAIL.n375 VTAIL.n294 1.93989
R1747 VTAIL.n38 VTAIL.n28 1.93989
R1748 VTAIL.n74 VTAIL.n12 1.93989
R1749 VTAIL.n87 VTAIL.n6 1.93989
R1750 VTAIL.n281 VTAIL.n200 1.93989
R1751 VTAIL.n268 VTAIL.n206 1.93989
R1752 VTAIL.n233 VTAIL.n223 1.93989
R1753 VTAIL.n185 VTAIL.n104 1.93989
R1754 VTAIL.n172 VTAIL.n110 1.93989
R1755 VTAIL.n137 VTAIL.n127 1.93989
R1756 VTAIL.n0 VTAIL.t2 1.92958
R1757 VTAIL.n0 VTAIL.t4 1.92958
R1758 VTAIL.n96 VTAIL.t6 1.92958
R1759 VTAIL.n96 VTAIL.t10 1.92958
R1760 VTAIL.n194 VTAIL.t7 1.92958
R1761 VTAIL.n194 VTAIL.t11 1.92958
R1762 VTAIL.n98 VTAIL.t1 1.92958
R1763 VTAIL.n98 VTAIL.t5 1.92958
R1764 VTAIL.n325 VTAIL.n318 1.16414
R1765 VTAIL.n363 VTAIL.n298 1.16414
R1766 VTAIL.n372 VTAIL.n371 1.16414
R1767 VTAIL.n37 VTAIL.n30 1.16414
R1768 VTAIL.n75 VTAIL.n10 1.16414
R1769 VTAIL.n84 VTAIL.n83 1.16414
R1770 VTAIL.n278 VTAIL.n277 1.16414
R1771 VTAIL.n269 VTAIL.n204 1.16414
R1772 VTAIL.n232 VTAIL.n225 1.16414
R1773 VTAIL.n182 VTAIL.n181 1.16414
R1774 VTAIL.n173 VTAIL.n108 1.16414
R1775 VTAIL.n136 VTAIL.n129 1.16414
R1776 VTAIL.n195 VTAIL.n193 0.862569
R1777 VTAIL.n95 VTAIL.n1 0.862569
R1778 VTAIL.n193 VTAIL.n99 0.784983
R1779 VTAIL.n289 VTAIL.n195 0.784983
R1780 VTAIL.n97 VTAIL.n95 0.784983
R1781 VTAIL VTAIL.n383 0.530672
R1782 VTAIL.n322 VTAIL.n321 0.388379
R1783 VTAIL.n367 VTAIL.n366 0.388379
R1784 VTAIL.n368 VTAIL.n296 0.388379
R1785 VTAIL.n34 VTAIL.n33 0.388379
R1786 VTAIL.n79 VTAIL.n78 0.388379
R1787 VTAIL.n80 VTAIL.n8 0.388379
R1788 VTAIL.n274 VTAIL.n202 0.388379
R1789 VTAIL.n273 VTAIL.n272 0.388379
R1790 VTAIL.n229 VTAIL.n228 0.388379
R1791 VTAIL.n178 VTAIL.n106 0.388379
R1792 VTAIL.n177 VTAIL.n176 0.388379
R1793 VTAIL.n133 VTAIL.n132 0.388379
R1794 VTAIL VTAIL.n1 0.25481
R1795 VTAIL.n324 VTAIL.n323 0.155672
R1796 VTAIL.n324 VTAIL.n315 0.155672
R1797 VTAIL.n331 VTAIL.n315 0.155672
R1798 VTAIL.n332 VTAIL.n331 0.155672
R1799 VTAIL.n332 VTAIL.n311 0.155672
R1800 VTAIL.n339 VTAIL.n311 0.155672
R1801 VTAIL.n340 VTAIL.n339 0.155672
R1802 VTAIL.n340 VTAIL.n307 0.155672
R1803 VTAIL.n347 VTAIL.n307 0.155672
R1804 VTAIL.n348 VTAIL.n347 0.155672
R1805 VTAIL.n348 VTAIL.n303 0.155672
R1806 VTAIL.n355 VTAIL.n303 0.155672
R1807 VTAIL.n356 VTAIL.n355 0.155672
R1808 VTAIL.n356 VTAIL.n299 0.155672
R1809 VTAIL.n364 VTAIL.n299 0.155672
R1810 VTAIL.n365 VTAIL.n364 0.155672
R1811 VTAIL.n365 VTAIL.n295 0.155672
R1812 VTAIL.n373 VTAIL.n295 0.155672
R1813 VTAIL.n374 VTAIL.n373 0.155672
R1814 VTAIL.n374 VTAIL.n291 0.155672
R1815 VTAIL.n381 VTAIL.n291 0.155672
R1816 VTAIL.n36 VTAIL.n35 0.155672
R1817 VTAIL.n36 VTAIL.n27 0.155672
R1818 VTAIL.n43 VTAIL.n27 0.155672
R1819 VTAIL.n44 VTAIL.n43 0.155672
R1820 VTAIL.n44 VTAIL.n23 0.155672
R1821 VTAIL.n51 VTAIL.n23 0.155672
R1822 VTAIL.n52 VTAIL.n51 0.155672
R1823 VTAIL.n52 VTAIL.n19 0.155672
R1824 VTAIL.n59 VTAIL.n19 0.155672
R1825 VTAIL.n60 VTAIL.n59 0.155672
R1826 VTAIL.n60 VTAIL.n15 0.155672
R1827 VTAIL.n67 VTAIL.n15 0.155672
R1828 VTAIL.n68 VTAIL.n67 0.155672
R1829 VTAIL.n68 VTAIL.n11 0.155672
R1830 VTAIL.n76 VTAIL.n11 0.155672
R1831 VTAIL.n77 VTAIL.n76 0.155672
R1832 VTAIL.n77 VTAIL.n7 0.155672
R1833 VTAIL.n85 VTAIL.n7 0.155672
R1834 VTAIL.n86 VTAIL.n85 0.155672
R1835 VTAIL.n86 VTAIL.n3 0.155672
R1836 VTAIL.n93 VTAIL.n3 0.155672
R1837 VTAIL.n287 VTAIL.n197 0.155672
R1838 VTAIL.n280 VTAIL.n197 0.155672
R1839 VTAIL.n280 VTAIL.n279 0.155672
R1840 VTAIL.n279 VTAIL.n201 0.155672
R1841 VTAIL.n271 VTAIL.n201 0.155672
R1842 VTAIL.n271 VTAIL.n270 0.155672
R1843 VTAIL.n270 VTAIL.n205 0.155672
R1844 VTAIL.n263 VTAIL.n205 0.155672
R1845 VTAIL.n263 VTAIL.n262 0.155672
R1846 VTAIL.n262 VTAIL.n210 0.155672
R1847 VTAIL.n255 VTAIL.n210 0.155672
R1848 VTAIL.n255 VTAIL.n254 0.155672
R1849 VTAIL.n254 VTAIL.n214 0.155672
R1850 VTAIL.n247 VTAIL.n214 0.155672
R1851 VTAIL.n247 VTAIL.n246 0.155672
R1852 VTAIL.n246 VTAIL.n218 0.155672
R1853 VTAIL.n239 VTAIL.n218 0.155672
R1854 VTAIL.n239 VTAIL.n238 0.155672
R1855 VTAIL.n238 VTAIL.n222 0.155672
R1856 VTAIL.n231 VTAIL.n222 0.155672
R1857 VTAIL.n231 VTAIL.n230 0.155672
R1858 VTAIL.n191 VTAIL.n101 0.155672
R1859 VTAIL.n184 VTAIL.n101 0.155672
R1860 VTAIL.n184 VTAIL.n183 0.155672
R1861 VTAIL.n183 VTAIL.n105 0.155672
R1862 VTAIL.n175 VTAIL.n105 0.155672
R1863 VTAIL.n175 VTAIL.n174 0.155672
R1864 VTAIL.n174 VTAIL.n109 0.155672
R1865 VTAIL.n167 VTAIL.n109 0.155672
R1866 VTAIL.n167 VTAIL.n166 0.155672
R1867 VTAIL.n166 VTAIL.n114 0.155672
R1868 VTAIL.n159 VTAIL.n114 0.155672
R1869 VTAIL.n159 VTAIL.n158 0.155672
R1870 VTAIL.n158 VTAIL.n118 0.155672
R1871 VTAIL.n151 VTAIL.n118 0.155672
R1872 VTAIL.n151 VTAIL.n150 0.155672
R1873 VTAIL.n150 VTAIL.n122 0.155672
R1874 VTAIL.n143 VTAIL.n122 0.155672
R1875 VTAIL.n143 VTAIL.n142 0.155672
R1876 VTAIL.n142 VTAIL.n126 0.155672
R1877 VTAIL.n135 VTAIL.n126 0.155672
R1878 VTAIL.n135 VTAIL.n134 0.155672
R1879 VN.n0 VN.t3 795.112
R1880 VN.n4 VN.t0 795.112
R1881 VN.n1 VN.t1 768.292
R1882 VN.n2 VN.t4 768.292
R1883 VN.n5 VN.t2 768.292
R1884 VN.n6 VN.t5 768.292
R1885 VN.n3 VN.n2 161.3
R1886 VN.n7 VN.n6 161.3
R1887 VN.n2 VN.n1 48.2005
R1888 VN.n6 VN.n5 48.2005
R1889 VN.n7 VN.n4 45.1367
R1890 VN.n3 VN.n0 45.1367
R1891 VN VN.n7 44.8547
R1892 VN.n5 VN.n4 13.3799
R1893 VN.n1 VN.n0 13.3799
R1894 VN VN.n3 0.0516364
R1895 VDD2.n183 VDD2.n95 756.745
R1896 VDD2.n88 VDD2.n0 756.745
R1897 VDD2.n184 VDD2.n183 585
R1898 VDD2.n182 VDD2.n181 585
R1899 VDD2.n99 VDD2.n98 585
R1900 VDD2.n176 VDD2.n175 585
R1901 VDD2.n174 VDD2.n173 585
R1902 VDD2.n172 VDD2.n102 585
R1903 VDD2.n106 VDD2.n103 585
R1904 VDD2.n167 VDD2.n166 585
R1905 VDD2.n165 VDD2.n164 585
R1906 VDD2.n108 VDD2.n107 585
R1907 VDD2.n159 VDD2.n158 585
R1908 VDD2.n157 VDD2.n156 585
R1909 VDD2.n112 VDD2.n111 585
R1910 VDD2.n151 VDD2.n150 585
R1911 VDD2.n149 VDD2.n148 585
R1912 VDD2.n116 VDD2.n115 585
R1913 VDD2.n143 VDD2.n142 585
R1914 VDD2.n141 VDD2.n140 585
R1915 VDD2.n120 VDD2.n119 585
R1916 VDD2.n135 VDD2.n134 585
R1917 VDD2.n133 VDD2.n132 585
R1918 VDD2.n124 VDD2.n123 585
R1919 VDD2.n127 VDD2.n126 585
R1920 VDD2.n31 VDD2.n30 585
R1921 VDD2.n28 VDD2.n27 585
R1922 VDD2.n37 VDD2.n36 585
R1923 VDD2.n39 VDD2.n38 585
R1924 VDD2.n24 VDD2.n23 585
R1925 VDD2.n45 VDD2.n44 585
R1926 VDD2.n47 VDD2.n46 585
R1927 VDD2.n20 VDD2.n19 585
R1928 VDD2.n53 VDD2.n52 585
R1929 VDD2.n55 VDD2.n54 585
R1930 VDD2.n16 VDD2.n15 585
R1931 VDD2.n61 VDD2.n60 585
R1932 VDD2.n63 VDD2.n62 585
R1933 VDD2.n12 VDD2.n11 585
R1934 VDD2.n69 VDD2.n68 585
R1935 VDD2.n72 VDD2.n71 585
R1936 VDD2.n70 VDD2.n8 585
R1937 VDD2.n77 VDD2.n7 585
R1938 VDD2.n79 VDD2.n78 585
R1939 VDD2.n81 VDD2.n80 585
R1940 VDD2.n4 VDD2.n3 585
R1941 VDD2.n87 VDD2.n86 585
R1942 VDD2.n89 VDD2.n88 585
R1943 VDD2.t0 VDD2.n125 327.466
R1944 VDD2.t2 VDD2.n29 327.466
R1945 VDD2.n183 VDD2.n182 171.744
R1946 VDD2.n182 VDD2.n98 171.744
R1947 VDD2.n175 VDD2.n98 171.744
R1948 VDD2.n175 VDD2.n174 171.744
R1949 VDD2.n174 VDD2.n102 171.744
R1950 VDD2.n106 VDD2.n102 171.744
R1951 VDD2.n166 VDD2.n106 171.744
R1952 VDD2.n166 VDD2.n165 171.744
R1953 VDD2.n165 VDD2.n107 171.744
R1954 VDD2.n158 VDD2.n107 171.744
R1955 VDD2.n158 VDD2.n157 171.744
R1956 VDD2.n157 VDD2.n111 171.744
R1957 VDD2.n150 VDD2.n111 171.744
R1958 VDD2.n150 VDD2.n149 171.744
R1959 VDD2.n149 VDD2.n115 171.744
R1960 VDD2.n142 VDD2.n115 171.744
R1961 VDD2.n142 VDD2.n141 171.744
R1962 VDD2.n141 VDD2.n119 171.744
R1963 VDD2.n134 VDD2.n119 171.744
R1964 VDD2.n134 VDD2.n133 171.744
R1965 VDD2.n133 VDD2.n123 171.744
R1966 VDD2.n126 VDD2.n123 171.744
R1967 VDD2.n30 VDD2.n27 171.744
R1968 VDD2.n37 VDD2.n27 171.744
R1969 VDD2.n38 VDD2.n37 171.744
R1970 VDD2.n38 VDD2.n23 171.744
R1971 VDD2.n45 VDD2.n23 171.744
R1972 VDD2.n46 VDD2.n45 171.744
R1973 VDD2.n46 VDD2.n19 171.744
R1974 VDD2.n53 VDD2.n19 171.744
R1975 VDD2.n54 VDD2.n53 171.744
R1976 VDD2.n54 VDD2.n15 171.744
R1977 VDD2.n61 VDD2.n15 171.744
R1978 VDD2.n62 VDD2.n61 171.744
R1979 VDD2.n62 VDD2.n11 171.744
R1980 VDD2.n69 VDD2.n11 171.744
R1981 VDD2.n71 VDD2.n69 171.744
R1982 VDD2.n71 VDD2.n70 171.744
R1983 VDD2.n70 VDD2.n7 171.744
R1984 VDD2.n79 VDD2.n7 171.744
R1985 VDD2.n80 VDD2.n79 171.744
R1986 VDD2.n80 VDD2.n3 171.744
R1987 VDD2.n87 VDD2.n3 171.744
R1988 VDD2.n88 VDD2.n87 171.744
R1989 VDD2.n126 VDD2.t0 85.8723
R1990 VDD2.n30 VDD2.t2 85.8723
R1991 VDD2.n94 VDD2.n93 70.5023
R1992 VDD2 VDD2.n189 70.4995
R1993 VDD2.n94 VDD2.n92 50.3668
R1994 VDD2.n188 VDD2.n187 49.8338
R1995 VDD2.n188 VDD2.n94 40.7907
R1996 VDD2.n127 VDD2.n125 16.3895
R1997 VDD2.n31 VDD2.n29 16.3895
R1998 VDD2.n173 VDD2.n172 13.1884
R1999 VDD2.n78 VDD2.n77 13.1884
R2000 VDD2.n176 VDD2.n101 12.8005
R2001 VDD2.n171 VDD2.n103 12.8005
R2002 VDD2.n128 VDD2.n124 12.8005
R2003 VDD2.n32 VDD2.n28 12.8005
R2004 VDD2.n76 VDD2.n8 12.8005
R2005 VDD2.n81 VDD2.n6 12.8005
R2006 VDD2.n177 VDD2.n99 12.0247
R2007 VDD2.n168 VDD2.n167 12.0247
R2008 VDD2.n132 VDD2.n131 12.0247
R2009 VDD2.n36 VDD2.n35 12.0247
R2010 VDD2.n73 VDD2.n72 12.0247
R2011 VDD2.n82 VDD2.n4 12.0247
R2012 VDD2.n181 VDD2.n180 11.249
R2013 VDD2.n164 VDD2.n105 11.249
R2014 VDD2.n135 VDD2.n122 11.249
R2015 VDD2.n39 VDD2.n26 11.249
R2016 VDD2.n68 VDD2.n10 11.249
R2017 VDD2.n86 VDD2.n85 11.249
R2018 VDD2.n184 VDD2.n97 10.4732
R2019 VDD2.n163 VDD2.n108 10.4732
R2020 VDD2.n136 VDD2.n120 10.4732
R2021 VDD2.n40 VDD2.n24 10.4732
R2022 VDD2.n67 VDD2.n12 10.4732
R2023 VDD2.n89 VDD2.n2 10.4732
R2024 VDD2.n185 VDD2.n95 9.69747
R2025 VDD2.n160 VDD2.n159 9.69747
R2026 VDD2.n140 VDD2.n139 9.69747
R2027 VDD2.n44 VDD2.n43 9.69747
R2028 VDD2.n64 VDD2.n63 9.69747
R2029 VDD2.n90 VDD2.n0 9.69747
R2030 VDD2.n187 VDD2.n186 9.45567
R2031 VDD2.n92 VDD2.n91 9.45567
R2032 VDD2.n153 VDD2.n152 9.3005
R2033 VDD2.n155 VDD2.n154 9.3005
R2034 VDD2.n110 VDD2.n109 9.3005
R2035 VDD2.n161 VDD2.n160 9.3005
R2036 VDD2.n163 VDD2.n162 9.3005
R2037 VDD2.n105 VDD2.n104 9.3005
R2038 VDD2.n169 VDD2.n168 9.3005
R2039 VDD2.n171 VDD2.n170 9.3005
R2040 VDD2.n186 VDD2.n185 9.3005
R2041 VDD2.n97 VDD2.n96 9.3005
R2042 VDD2.n180 VDD2.n179 9.3005
R2043 VDD2.n178 VDD2.n177 9.3005
R2044 VDD2.n101 VDD2.n100 9.3005
R2045 VDD2.n114 VDD2.n113 9.3005
R2046 VDD2.n147 VDD2.n146 9.3005
R2047 VDD2.n145 VDD2.n144 9.3005
R2048 VDD2.n118 VDD2.n117 9.3005
R2049 VDD2.n139 VDD2.n138 9.3005
R2050 VDD2.n137 VDD2.n136 9.3005
R2051 VDD2.n122 VDD2.n121 9.3005
R2052 VDD2.n131 VDD2.n130 9.3005
R2053 VDD2.n129 VDD2.n128 9.3005
R2054 VDD2.n91 VDD2.n90 9.3005
R2055 VDD2.n2 VDD2.n1 9.3005
R2056 VDD2.n85 VDD2.n84 9.3005
R2057 VDD2.n83 VDD2.n82 9.3005
R2058 VDD2.n6 VDD2.n5 9.3005
R2059 VDD2.n51 VDD2.n50 9.3005
R2060 VDD2.n49 VDD2.n48 9.3005
R2061 VDD2.n22 VDD2.n21 9.3005
R2062 VDD2.n43 VDD2.n42 9.3005
R2063 VDD2.n41 VDD2.n40 9.3005
R2064 VDD2.n26 VDD2.n25 9.3005
R2065 VDD2.n35 VDD2.n34 9.3005
R2066 VDD2.n33 VDD2.n32 9.3005
R2067 VDD2.n18 VDD2.n17 9.3005
R2068 VDD2.n57 VDD2.n56 9.3005
R2069 VDD2.n59 VDD2.n58 9.3005
R2070 VDD2.n14 VDD2.n13 9.3005
R2071 VDD2.n65 VDD2.n64 9.3005
R2072 VDD2.n67 VDD2.n66 9.3005
R2073 VDD2.n10 VDD2.n9 9.3005
R2074 VDD2.n74 VDD2.n73 9.3005
R2075 VDD2.n76 VDD2.n75 9.3005
R2076 VDD2.n156 VDD2.n110 8.92171
R2077 VDD2.n143 VDD2.n118 8.92171
R2078 VDD2.n47 VDD2.n22 8.92171
R2079 VDD2.n60 VDD2.n14 8.92171
R2080 VDD2.n155 VDD2.n112 8.14595
R2081 VDD2.n144 VDD2.n116 8.14595
R2082 VDD2.n48 VDD2.n20 8.14595
R2083 VDD2.n59 VDD2.n16 8.14595
R2084 VDD2.n152 VDD2.n151 7.3702
R2085 VDD2.n148 VDD2.n147 7.3702
R2086 VDD2.n52 VDD2.n51 7.3702
R2087 VDD2.n56 VDD2.n55 7.3702
R2088 VDD2.n151 VDD2.n114 6.59444
R2089 VDD2.n148 VDD2.n114 6.59444
R2090 VDD2.n52 VDD2.n18 6.59444
R2091 VDD2.n55 VDD2.n18 6.59444
R2092 VDD2.n152 VDD2.n112 5.81868
R2093 VDD2.n147 VDD2.n116 5.81868
R2094 VDD2.n51 VDD2.n20 5.81868
R2095 VDD2.n56 VDD2.n16 5.81868
R2096 VDD2.n156 VDD2.n155 5.04292
R2097 VDD2.n144 VDD2.n143 5.04292
R2098 VDD2.n48 VDD2.n47 5.04292
R2099 VDD2.n60 VDD2.n59 5.04292
R2100 VDD2.n187 VDD2.n95 4.26717
R2101 VDD2.n159 VDD2.n110 4.26717
R2102 VDD2.n140 VDD2.n118 4.26717
R2103 VDD2.n44 VDD2.n22 4.26717
R2104 VDD2.n63 VDD2.n14 4.26717
R2105 VDD2.n92 VDD2.n0 4.26717
R2106 VDD2.n129 VDD2.n125 3.70982
R2107 VDD2.n33 VDD2.n29 3.70982
R2108 VDD2.n185 VDD2.n184 3.49141
R2109 VDD2.n160 VDD2.n108 3.49141
R2110 VDD2.n139 VDD2.n120 3.49141
R2111 VDD2.n43 VDD2.n24 3.49141
R2112 VDD2.n64 VDD2.n12 3.49141
R2113 VDD2.n90 VDD2.n89 3.49141
R2114 VDD2.n181 VDD2.n97 2.71565
R2115 VDD2.n164 VDD2.n163 2.71565
R2116 VDD2.n136 VDD2.n135 2.71565
R2117 VDD2.n40 VDD2.n39 2.71565
R2118 VDD2.n68 VDD2.n67 2.71565
R2119 VDD2.n86 VDD2.n2 2.71565
R2120 VDD2.n180 VDD2.n99 1.93989
R2121 VDD2.n167 VDD2.n105 1.93989
R2122 VDD2.n132 VDD2.n122 1.93989
R2123 VDD2.n36 VDD2.n26 1.93989
R2124 VDD2.n72 VDD2.n10 1.93989
R2125 VDD2.n85 VDD2.n4 1.93989
R2126 VDD2.n189 VDD2.t3 1.92958
R2127 VDD2.n189 VDD2.t5 1.92958
R2128 VDD2.n93 VDD2.t4 1.92958
R2129 VDD2.n93 VDD2.t1 1.92958
R2130 VDD2.n177 VDD2.n176 1.16414
R2131 VDD2.n168 VDD2.n103 1.16414
R2132 VDD2.n131 VDD2.n124 1.16414
R2133 VDD2.n35 VDD2.n28 1.16414
R2134 VDD2.n73 VDD2.n8 1.16414
R2135 VDD2.n82 VDD2.n81 1.16414
R2136 VDD2 VDD2.n188 0.647052
R2137 VDD2.n173 VDD2.n101 0.388379
R2138 VDD2.n172 VDD2.n171 0.388379
R2139 VDD2.n128 VDD2.n127 0.388379
R2140 VDD2.n32 VDD2.n31 0.388379
R2141 VDD2.n77 VDD2.n76 0.388379
R2142 VDD2.n78 VDD2.n6 0.388379
R2143 VDD2.n186 VDD2.n96 0.155672
R2144 VDD2.n179 VDD2.n96 0.155672
R2145 VDD2.n179 VDD2.n178 0.155672
R2146 VDD2.n178 VDD2.n100 0.155672
R2147 VDD2.n170 VDD2.n100 0.155672
R2148 VDD2.n170 VDD2.n169 0.155672
R2149 VDD2.n169 VDD2.n104 0.155672
R2150 VDD2.n162 VDD2.n104 0.155672
R2151 VDD2.n162 VDD2.n161 0.155672
R2152 VDD2.n161 VDD2.n109 0.155672
R2153 VDD2.n154 VDD2.n109 0.155672
R2154 VDD2.n154 VDD2.n153 0.155672
R2155 VDD2.n153 VDD2.n113 0.155672
R2156 VDD2.n146 VDD2.n113 0.155672
R2157 VDD2.n146 VDD2.n145 0.155672
R2158 VDD2.n145 VDD2.n117 0.155672
R2159 VDD2.n138 VDD2.n117 0.155672
R2160 VDD2.n138 VDD2.n137 0.155672
R2161 VDD2.n137 VDD2.n121 0.155672
R2162 VDD2.n130 VDD2.n121 0.155672
R2163 VDD2.n130 VDD2.n129 0.155672
R2164 VDD2.n34 VDD2.n33 0.155672
R2165 VDD2.n34 VDD2.n25 0.155672
R2166 VDD2.n41 VDD2.n25 0.155672
R2167 VDD2.n42 VDD2.n41 0.155672
R2168 VDD2.n42 VDD2.n21 0.155672
R2169 VDD2.n49 VDD2.n21 0.155672
R2170 VDD2.n50 VDD2.n49 0.155672
R2171 VDD2.n50 VDD2.n17 0.155672
R2172 VDD2.n57 VDD2.n17 0.155672
R2173 VDD2.n58 VDD2.n57 0.155672
R2174 VDD2.n58 VDD2.n13 0.155672
R2175 VDD2.n65 VDD2.n13 0.155672
R2176 VDD2.n66 VDD2.n65 0.155672
R2177 VDD2.n66 VDD2.n9 0.155672
R2178 VDD2.n74 VDD2.n9 0.155672
R2179 VDD2.n75 VDD2.n74 0.155672
R2180 VDD2.n75 VDD2.n5 0.155672
R2181 VDD2.n83 VDD2.n5 0.155672
R2182 VDD2.n84 VDD2.n83 0.155672
R2183 VDD2.n84 VDD2.n1 0.155672
R2184 VDD2.n91 VDD2.n1 0.155672
C0 VN B 0.795248f
C1 VDD1 VP 5.53353f
C2 VTAIL VDD1 14.2665f
C3 VN VP 5.86117f
C4 VN VTAIL 4.85512f
C5 B VP 1.1422f
C6 VTAIL B 3.46935f
C7 VDD2 w_n1698_n4338# 2.15912f
C8 VTAIL VP 4.86998f
C9 VDD1 VDD2 0.66973f
C10 VN VDD2 5.39968f
C11 VDD1 w_n1698_n4338# 2.13879f
C12 VN w_n1698_n4338# 2.81356f
C13 VDD2 B 1.89794f
C14 VN VDD1 0.148034f
C15 VDD2 VP 0.288344f
C16 VTAIL VDD2 14.2963f
C17 w_n1698_n4338# B 8.24817f
C18 VDD1 B 1.87178f
C19 w_n1698_n4338# VP 3.02745f
C20 VTAIL w_n1698_n4338# 3.72763f
C21 VDD2 VSUBS 1.551827f
C22 VDD1 VSUBS 1.286031f
C23 VTAIL VSUBS 0.856193f
C24 VN VSUBS 4.85827f
C25 VP VSUBS 1.561846f
C26 B VSUBS 3.045006f
C27 w_n1698_n4338# VSUBS 90.163795f
C28 VDD2.n0 VSUBS 0.029002f
C29 VDD2.n1 VSUBS 0.026807f
C30 VDD2.n2 VSUBS 0.014405f
C31 VDD2.n3 VSUBS 0.034048f
C32 VDD2.n4 VSUBS 0.015252f
C33 VDD2.n5 VSUBS 0.026807f
C34 VDD2.n6 VSUBS 0.014405f
C35 VDD2.n7 VSUBS 0.034048f
C36 VDD2.n8 VSUBS 0.015252f
C37 VDD2.n9 VSUBS 0.026807f
C38 VDD2.n10 VSUBS 0.014405f
C39 VDD2.n11 VSUBS 0.034048f
C40 VDD2.n12 VSUBS 0.015252f
C41 VDD2.n13 VSUBS 0.026807f
C42 VDD2.n14 VSUBS 0.014405f
C43 VDD2.n15 VSUBS 0.034048f
C44 VDD2.n16 VSUBS 0.015252f
C45 VDD2.n17 VSUBS 0.026807f
C46 VDD2.n18 VSUBS 0.014405f
C47 VDD2.n19 VSUBS 0.034048f
C48 VDD2.n20 VSUBS 0.015252f
C49 VDD2.n21 VSUBS 0.026807f
C50 VDD2.n22 VSUBS 0.014405f
C51 VDD2.n23 VSUBS 0.034048f
C52 VDD2.n24 VSUBS 0.015252f
C53 VDD2.n25 VSUBS 0.026807f
C54 VDD2.n26 VSUBS 0.014405f
C55 VDD2.n27 VSUBS 0.034048f
C56 VDD2.n28 VSUBS 0.015252f
C57 VDD2.n29 VSUBS 0.203594f
C58 VDD2.t2 VSUBS 0.073013f
C59 VDD2.n30 VSUBS 0.025536f
C60 VDD2.n31 VSUBS 0.02166f
C61 VDD2.n32 VSUBS 0.014405f
C62 VDD2.n33 VSUBS 1.93683f
C63 VDD2.n34 VSUBS 0.026807f
C64 VDD2.n35 VSUBS 0.014405f
C65 VDD2.n36 VSUBS 0.015252f
C66 VDD2.n37 VSUBS 0.034048f
C67 VDD2.n38 VSUBS 0.034048f
C68 VDD2.n39 VSUBS 0.015252f
C69 VDD2.n40 VSUBS 0.014405f
C70 VDD2.n41 VSUBS 0.026807f
C71 VDD2.n42 VSUBS 0.026807f
C72 VDD2.n43 VSUBS 0.014405f
C73 VDD2.n44 VSUBS 0.015252f
C74 VDD2.n45 VSUBS 0.034048f
C75 VDD2.n46 VSUBS 0.034048f
C76 VDD2.n47 VSUBS 0.015252f
C77 VDD2.n48 VSUBS 0.014405f
C78 VDD2.n49 VSUBS 0.026807f
C79 VDD2.n50 VSUBS 0.026807f
C80 VDD2.n51 VSUBS 0.014405f
C81 VDD2.n52 VSUBS 0.015252f
C82 VDD2.n53 VSUBS 0.034048f
C83 VDD2.n54 VSUBS 0.034048f
C84 VDD2.n55 VSUBS 0.015252f
C85 VDD2.n56 VSUBS 0.014405f
C86 VDD2.n57 VSUBS 0.026807f
C87 VDD2.n58 VSUBS 0.026807f
C88 VDD2.n59 VSUBS 0.014405f
C89 VDD2.n60 VSUBS 0.015252f
C90 VDD2.n61 VSUBS 0.034048f
C91 VDD2.n62 VSUBS 0.034048f
C92 VDD2.n63 VSUBS 0.015252f
C93 VDD2.n64 VSUBS 0.014405f
C94 VDD2.n65 VSUBS 0.026807f
C95 VDD2.n66 VSUBS 0.026807f
C96 VDD2.n67 VSUBS 0.014405f
C97 VDD2.n68 VSUBS 0.015252f
C98 VDD2.n69 VSUBS 0.034048f
C99 VDD2.n70 VSUBS 0.034048f
C100 VDD2.n71 VSUBS 0.034048f
C101 VDD2.n72 VSUBS 0.015252f
C102 VDD2.n73 VSUBS 0.014405f
C103 VDD2.n74 VSUBS 0.026807f
C104 VDD2.n75 VSUBS 0.026807f
C105 VDD2.n76 VSUBS 0.014405f
C106 VDD2.n77 VSUBS 0.014829f
C107 VDD2.n78 VSUBS 0.014829f
C108 VDD2.n79 VSUBS 0.034048f
C109 VDD2.n80 VSUBS 0.034048f
C110 VDD2.n81 VSUBS 0.015252f
C111 VDD2.n82 VSUBS 0.014405f
C112 VDD2.n83 VSUBS 0.026807f
C113 VDD2.n84 VSUBS 0.026807f
C114 VDD2.n85 VSUBS 0.014405f
C115 VDD2.n86 VSUBS 0.015252f
C116 VDD2.n87 VSUBS 0.034048f
C117 VDD2.n88 VSUBS 0.080884f
C118 VDD2.n89 VSUBS 0.015252f
C119 VDD2.n90 VSUBS 0.014405f
C120 VDD2.n91 VSUBS 0.063794f
C121 VDD2.n92 VSUBS 0.060215f
C122 VDD2.t4 VSUBS 0.356946f
C123 VDD2.t1 VSUBS 0.356946f
C124 VDD2.n93 VSUBS 2.94613f
C125 VDD2.n94 VSUBS 2.54988f
C126 VDD2.n95 VSUBS 0.029002f
C127 VDD2.n96 VSUBS 0.026807f
C128 VDD2.n97 VSUBS 0.014405f
C129 VDD2.n98 VSUBS 0.034048f
C130 VDD2.n99 VSUBS 0.015252f
C131 VDD2.n100 VSUBS 0.026807f
C132 VDD2.n101 VSUBS 0.014405f
C133 VDD2.n102 VSUBS 0.034048f
C134 VDD2.n103 VSUBS 0.015252f
C135 VDD2.n104 VSUBS 0.026807f
C136 VDD2.n105 VSUBS 0.014405f
C137 VDD2.n106 VSUBS 0.034048f
C138 VDD2.n107 VSUBS 0.034048f
C139 VDD2.n108 VSUBS 0.015252f
C140 VDD2.n109 VSUBS 0.026807f
C141 VDD2.n110 VSUBS 0.014405f
C142 VDD2.n111 VSUBS 0.034048f
C143 VDD2.n112 VSUBS 0.015252f
C144 VDD2.n113 VSUBS 0.026807f
C145 VDD2.n114 VSUBS 0.014405f
C146 VDD2.n115 VSUBS 0.034048f
C147 VDD2.n116 VSUBS 0.015252f
C148 VDD2.n117 VSUBS 0.026807f
C149 VDD2.n118 VSUBS 0.014405f
C150 VDD2.n119 VSUBS 0.034048f
C151 VDD2.n120 VSUBS 0.015252f
C152 VDD2.n121 VSUBS 0.026807f
C153 VDD2.n122 VSUBS 0.014405f
C154 VDD2.n123 VSUBS 0.034048f
C155 VDD2.n124 VSUBS 0.015252f
C156 VDD2.n125 VSUBS 0.203594f
C157 VDD2.t0 VSUBS 0.073013f
C158 VDD2.n126 VSUBS 0.025536f
C159 VDD2.n127 VSUBS 0.02166f
C160 VDD2.n128 VSUBS 0.014405f
C161 VDD2.n129 VSUBS 1.93683f
C162 VDD2.n130 VSUBS 0.026807f
C163 VDD2.n131 VSUBS 0.014405f
C164 VDD2.n132 VSUBS 0.015252f
C165 VDD2.n133 VSUBS 0.034048f
C166 VDD2.n134 VSUBS 0.034048f
C167 VDD2.n135 VSUBS 0.015252f
C168 VDD2.n136 VSUBS 0.014405f
C169 VDD2.n137 VSUBS 0.026807f
C170 VDD2.n138 VSUBS 0.026807f
C171 VDD2.n139 VSUBS 0.014405f
C172 VDD2.n140 VSUBS 0.015252f
C173 VDD2.n141 VSUBS 0.034048f
C174 VDD2.n142 VSUBS 0.034048f
C175 VDD2.n143 VSUBS 0.015252f
C176 VDD2.n144 VSUBS 0.014405f
C177 VDD2.n145 VSUBS 0.026807f
C178 VDD2.n146 VSUBS 0.026807f
C179 VDD2.n147 VSUBS 0.014405f
C180 VDD2.n148 VSUBS 0.015252f
C181 VDD2.n149 VSUBS 0.034048f
C182 VDD2.n150 VSUBS 0.034048f
C183 VDD2.n151 VSUBS 0.015252f
C184 VDD2.n152 VSUBS 0.014405f
C185 VDD2.n153 VSUBS 0.026807f
C186 VDD2.n154 VSUBS 0.026807f
C187 VDD2.n155 VSUBS 0.014405f
C188 VDD2.n156 VSUBS 0.015252f
C189 VDD2.n157 VSUBS 0.034048f
C190 VDD2.n158 VSUBS 0.034048f
C191 VDD2.n159 VSUBS 0.015252f
C192 VDD2.n160 VSUBS 0.014405f
C193 VDD2.n161 VSUBS 0.026807f
C194 VDD2.n162 VSUBS 0.026807f
C195 VDD2.n163 VSUBS 0.014405f
C196 VDD2.n164 VSUBS 0.015252f
C197 VDD2.n165 VSUBS 0.034048f
C198 VDD2.n166 VSUBS 0.034048f
C199 VDD2.n167 VSUBS 0.015252f
C200 VDD2.n168 VSUBS 0.014405f
C201 VDD2.n169 VSUBS 0.026807f
C202 VDD2.n170 VSUBS 0.026807f
C203 VDD2.n171 VSUBS 0.014405f
C204 VDD2.n172 VSUBS 0.014829f
C205 VDD2.n173 VSUBS 0.014829f
C206 VDD2.n174 VSUBS 0.034048f
C207 VDD2.n175 VSUBS 0.034048f
C208 VDD2.n176 VSUBS 0.015252f
C209 VDD2.n177 VSUBS 0.014405f
C210 VDD2.n178 VSUBS 0.026807f
C211 VDD2.n179 VSUBS 0.026807f
C212 VDD2.n180 VSUBS 0.014405f
C213 VDD2.n181 VSUBS 0.015252f
C214 VDD2.n182 VSUBS 0.034048f
C215 VDD2.n183 VSUBS 0.080884f
C216 VDD2.n184 VSUBS 0.015252f
C217 VDD2.n185 VSUBS 0.014405f
C218 VDD2.n186 VSUBS 0.063794f
C219 VDD2.n187 VSUBS 0.059158f
C220 VDD2.n188 VSUBS 2.55984f
C221 VDD2.t3 VSUBS 0.356946f
C222 VDD2.t5 VSUBS 0.356946f
C223 VDD2.n189 VSUBS 2.94609f
C224 VN.t3 VSUBS 1.61825f
C225 VN.n0 VSUBS 0.591352f
C226 VN.t1 VSUBS 1.59764f
C227 VN.n1 VSUBS 0.623813f
C228 VN.t4 VSUBS 1.59764f
C229 VN.n2 VSUBS 0.610742f
C230 VN.n3 VSUBS 0.230438f
C231 VN.t0 VSUBS 1.61825f
C232 VN.n4 VSUBS 0.591352f
C233 VN.t2 VSUBS 1.59764f
C234 VN.n5 VSUBS 0.623813f
C235 VN.t5 VSUBS 1.59764f
C236 VN.n6 VSUBS 0.610742f
C237 VN.n7 VSUBS 2.83449f
C238 VTAIL.t2 VSUBS 0.388495f
C239 VTAIL.t4 VSUBS 0.388495f
C240 VTAIL.n0 VSUBS 3.03117f
C241 VTAIL.n1 VSUBS 0.804966f
C242 VTAIL.n2 VSUBS 0.031566f
C243 VTAIL.n3 VSUBS 0.029176f
C244 VTAIL.n4 VSUBS 0.015678f
C245 VTAIL.n5 VSUBS 0.037057f
C246 VTAIL.n6 VSUBS 0.0166f
C247 VTAIL.n7 VSUBS 0.029176f
C248 VTAIL.n8 VSUBS 0.015678f
C249 VTAIL.n9 VSUBS 0.037057f
C250 VTAIL.n10 VSUBS 0.0166f
C251 VTAIL.n11 VSUBS 0.029176f
C252 VTAIL.n12 VSUBS 0.015678f
C253 VTAIL.n13 VSUBS 0.037057f
C254 VTAIL.n14 VSUBS 0.0166f
C255 VTAIL.n15 VSUBS 0.029176f
C256 VTAIL.n16 VSUBS 0.015678f
C257 VTAIL.n17 VSUBS 0.037057f
C258 VTAIL.n18 VSUBS 0.0166f
C259 VTAIL.n19 VSUBS 0.029176f
C260 VTAIL.n20 VSUBS 0.015678f
C261 VTAIL.n21 VSUBS 0.037057f
C262 VTAIL.n22 VSUBS 0.0166f
C263 VTAIL.n23 VSUBS 0.029176f
C264 VTAIL.n24 VSUBS 0.015678f
C265 VTAIL.n25 VSUBS 0.037057f
C266 VTAIL.n26 VSUBS 0.0166f
C267 VTAIL.n27 VSUBS 0.029176f
C268 VTAIL.n28 VSUBS 0.015678f
C269 VTAIL.n29 VSUBS 0.037057f
C270 VTAIL.n30 VSUBS 0.0166f
C271 VTAIL.n31 VSUBS 0.221589f
C272 VTAIL.t8 VSUBS 0.079467f
C273 VTAIL.n32 VSUBS 0.027793f
C274 VTAIL.n33 VSUBS 0.023574f
C275 VTAIL.n34 VSUBS 0.015678f
C276 VTAIL.n35 VSUBS 2.10801f
C277 VTAIL.n36 VSUBS 0.029176f
C278 VTAIL.n37 VSUBS 0.015678f
C279 VTAIL.n38 VSUBS 0.0166f
C280 VTAIL.n39 VSUBS 0.037057f
C281 VTAIL.n40 VSUBS 0.037057f
C282 VTAIL.n41 VSUBS 0.0166f
C283 VTAIL.n42 VSUBS 0.015678f
C284 VTAIL.n43 VSUBS 0.029176f
C285 VTAIL.n44 VSUBS 0.029176f
C286 VTAIL.n45 VSUBS 0.015678f
C287 VTAIL.n46 VSUBS 0.0166f
C288 VTAIL.n47 VSUBS 0.037057f
C289 VTAIL.n48 VSUBS 0.037057f
C290 VTAIL.n49 VSUBS 0.0166f
C291 VTAIL.n50 VSUBS 0.015678f
C292 VTAIL.n51 VSUBS 0.029176f
C293 VTAIL.n52 VSUBS 0.029176f
C294 VTAIL.n53 VSUBS 0.015678f
C295 VTAIL.n54 VSUBS 0.0166f
C296 VTAIL.n55 VSUBS 0.037057f
C297 VTAIL.n56 VSUBS 0.037057f
C298 VTAIL.n57 VSUBS 0.0166f
C299 VTAIL.n58 VSUBS 0.015678f
C300 VTAIL.n59 VSUBS 0.029176f
C301 VTAIL.n60 VSUBS 0.029176f
C302 VTAIL.n61 VSUBS 0.015678f
C303 VTAIL.n62 VSUBS 0.0166f
C304 VTAIL.n63 VSUBS 0.037057f
C305 VTAIL.n64 VSUBS 0.037057f
C306 VTAIL.n65 VSUBS 0.0166f
C307 VTAIL.n66 VSUBS 0.015678f
C308 VTAIL.n67 VSUBS 0.029176f
C309 VTAIL.n68 VSUBS 0.029176f
C310 VTAIL.n69 VSUBS 0.015678f
C311 VTAIL.n70 VSUBS 0.0166f
C312 VTAIL.n71 VSUBS 0.037057f
C313 VTAIL.n72 VSUBS 0.037057f
C314 VTAIL.n73 VSUBS 0.037057f
C315 VTAIL.n74 VSUBS 0.0166f
C316 VTAIL.n75 VSUBS 0.015678f
C317 VTAIL.n76 VSUBS 0.029176f
C318 VTAIL.n77 VSUBS 0.029176f
C319 VTAIL.n78 VSUBS 0.015678f
C320 VTAIL.n79 VSUBS 0.016139f
C321 VTAIL.n80 VSUBS 0.016139f
C322 VTAIL.n81 VSUBS 0.037057f
C323 VTAIL.n82 VSUBS 0.037057f
C324 VTAIL.n83 VSUBS 0.0166f
C325 VTAIL.n84 VSUBS 0.015678f
C326 VTAIL.n85 VSUBS 0.029176f
C327 VTAIL.n86 VSUBS 0.029176f
C328 VTAIL.n87 VSUBS 0.015678f
C329 VTAIL.n88 VSUBS 0.0166f
C330 VTAIL.n89 VSUBS 0.037057f
C331 VTAIL.n90 VSUBS 0.088033f
C332 VTAIL.n91 VSUBS 0.0166f
C333 VTAIL.n92 VSUBS 0.015678f
C334 VTAIL.n93 VSUBS 0.069433f
C335 VTAIL.n94 VSUBS 0.044257f
C336 VTAIL.n95 VSUBS 0.180842f
C337 VTAIL.t6 VSUBS 0.388495f
C338 VTAIL.t10 VSUBS 0.388495f
C339 VTAIL.n96 VSUBS 3.03117f
C340 VTAIL.n97 VSUBS 2.68321f
C341 VTAIL.t1 VSUBS 0.388495f
C342 VTAIL.t5 VSUBS 0.388495f
C343 VTAIL.n98 VSUBS 3.03118f
C344 VTAIL.n99 VSUBS 2.6832f
C345 VTAIL.n100 VSUBS 0.031566f
C346 VTAIL.n101 VSUBS 0.029176f
C347 VTAIL.n102 VSUBS 0.015678f
C348 VTAIL.n103 VSUBS 0.037057f
C349 VTAIL.n104 VSUBS 0.0166f
C350 VTAIL.n105 VSUBS 0.029176f
C351 VTAIL.n106 VSUBS 0.015678f
C352 VTAIL.n107 VSUBS 0.037057f
C353 VTAIL.n108 VSUBS 0.0166f
C354 VTAIL.n109 VSUBS 0.029176f
C355 VTAIL.n110 VSUBS 0.015678f
C356 VTAIL.n111 VSUBS 0.037057f
C357 VTAIL.n112 VSUBS 0.037057f
C358 VTAIL.n113 VSUBS 0.0166f
C359 VTAIL.n114 VSUBS 0.029176f
C360 VTAIL.n115 VSUBS 0.015678f
C361 VTAIL.n116 VSUBS 0.037057f
C362 VTAIL.n117 VSUBS 0.0166f
C363 VTAIL.n118 VSUBS 0.029176f
C364 VTAIL.n119 VSUBS 0.015678f
C365 VTAIL.n120 VSUBS 0.037057f
C366 VTAIL.n121 VSUBS 0.0166f
C367 VTAIL.n122 VSUBS 0.029176f
C368 VTAIL.n123 VSUBS 0.015678f
C369 VTAIL.n124 VSUBS 0.037057f
C370 VTAIL.n125 VSUBS 0.0166f
C371 VTAIL.n126 VSUBS 0.029176f
C372 VTAIL.n127 VSUBS 0.015678f
C373 VTAIL.n128 VSUBS 0.037057f
C374 VTAIL.n129 VSUBS 0.0166f
C375 VTAIL.n130 VSUBS 0.221589f
C376 VTAIL.t3 VSUBS 0.079467f
C377 VTAIL.n131 VSUBS 0.027793f
C378 VTAIL.n132 VSUBS 0.023574f
C379 VTAIL.n133 VSUBS 0.015678f
C380 VTAIL.n134 VSUBS 2.10801f
C381 VTAIL.n135 VSUBS 0.029176f
C382 VTAIL.n136 VSUBS 0.015678f
C383 VTAIL.n137 VSUBS 0.0166f
C384 VTAIL.n138 VSUBS 0.037057f
C385 VTAIL.n139 VSUBS 0.037057f
C386 VTAIL.n140 VSUBS 0.0166f
C387 VTAIL.n141 VSUBS 0.015678f
C388 VTAIL.n142 VSUBS 0.029176f
C389 VTAIL.n143 VSUBS 0.029176f
C390 VTAIL.n144 VSUBS 0.015678f
C391 VTAIL.n145 VSUBS 0.0166f
C392 VTAIL.n146 VSUBS 0.037057f
C393 VTAIL.n147 VSUBS 0.037057f
C394 VTAIL.n148 VSUBS 0.0166f
C395 VTAIL.n149 VSUBS 0.015678f
C396 VTAIL.n150 VSUBS 0.029176f
C397 VTAIL.n151 VSUBS 0.029176f
C398 VTAIL.n152 VSUBS 0.015678f
C399 VTAIL.n153 VSUBS 0.0166f
C400 VTAIL.n154 VSUBS 0.037057f
C401 VTAIL.n155 VSUBS 0.037057f
C402 VTAIL.n156 VSUBS 0.0166f
C403 VTAIL.n157 VSUBS 0.015678f
C404 VTAIL.n158 VSUBS 0.029176f
C405 VTAIL.n159 VSUBS 0.029176f
C406 VTAIL.n160 VSUBS 0.015678f
C407 VTAIL.n161 VSUBS 0.0166f
C408 VTAIL.n162 VSUBS 0.037057f
C409 VTAIL.n163 VSUBS 0.037057f
C410 VTAIL.n164 VSUBS 0.0166f
C411 VTAIL.n165 VSUBS 0.015678f
C412 VTAIL.n166 VSUBS 0.029176f
C413 VTAIL.n167 VSUBS 0.029176f
C414 VTAIL.n168 VSUBS 0.015678f
C415 VTAIL.n169 VSUBS 0.0166f
C416 VTAIL.n170 VSUBS 0.037057f
C417 VTAIL.n171 VSUBS 0.037057f
C418 VTAIL.n172 VSUBS 0.0166f
C419 VTAIL.n173 VSUBS 0.015678f
C420 VTAIL.n174 VSUBS 0.029176f
C421 VTAIL.n175 VSUBS 0.029176f
C422 VTAIL.n176 VSUBS 0.015678f
C423 VTAIL.n177 VSUBS 0.016139f
C424 VTAIL.n178 VSUBS 0.016139f
C425 VTAIL.n179 VSUBS 0.037057f
C426 VTAIL.n180 VSUBS 0.037057f
C427 VTAIL.n181 VSUBS 0.0166f
C428 VTAIL.n182 VSUBS 0.015678f
C429 VTAIL.n183 VSUBS 0.029176f
C430 VTAIL.n184 VSUBS 0.029176f
C431 VTAIL.n185 VSUBS 0.015678f
C432 VTAIL.n186 VSUBS 0.0166f
C433 VTAIL.n187 VSUBS 0.037057f
C434 VTAIL.n188 VSUBS 0.088033f
C435 VTAIL.n189 VSUBS 0.0166f
C436 VTAIL.n190 VSUBS 0.015678f
C437 VTAIL.n191 VSUBS 0.069433f
C438 VTAIL.n192 VSUBS 0.044257f
C439 VTAIL.n193 VSUBS 0.180842f
C440 VTAIL.t7 VSUBS 0.388495f
C441 VTAIL.t11 VSUBS 0.388495f
C442 VTAIL.n194 VSUBS 3.03118f
C443 VTAIL.n195 VSUBS 0.854791f
C444 VTAIL.n196 VSUBS 0.031566f
C445 VTAIL.n197 VSUBS 0.029176f
C446 VTAIL.n198 VSUBS 0.015678f
C447 VTAIL.n199 VSUBS 0.037057f
C448 VTAIL.n200 VSUBS 0.0166f
C449 VTAIL.n201 VSUBS 0.029176f
C450 VTAIL.n202 VSUBS 0.015678f
C451 VTAIL.n203 VSUBS 0.037057f
C452 VTAIL.n204 VSUBS 0.0166f
C453 VTAIL.n205 VSUBS 0.029176f
C454 VTAIL.n206 VSUBS 0.015678f
C455 VTAIL.n207 VSUBS 0.037057f
C456 VTAIL.n208 VSUBS 0.037057f
C457 VTAIL.n209 VSUBS 0.0166f
C458 VTAIL.n210 VSUBS 0.029176f
C459 VTAIL.n211 VSUBS 0.015678f
C460 VTAIL.n212 VSUBS 0.037057f
C461 VTAIL.n213 VSUBS 0.0166f
C462 VTAIL.n214 VSUBS 0.029176f
C463 VTAIL.n215 VSUBS 0.015678f
C464 VTAIL.n216 VSUBS 0.037057f
C465 VTAIL.n217 VSUBS 0.0166f
C466 VTAIL.n218 VSUBS 0.029176f
C467 VTAIL.n219 VSUBS 0.015678f
C468 VTAIL.n220 VSUBS 0.037057f
C469 VTAIL.n221 VSUBS 0.0166f
C470 VTAIL.n222 VSUBS 0.029176f
C471 VTAIL.n223 VSUBS 0.015678f
C472 VTAIL.n224 VSUBS 0.037057f
C473 VTAIL.n225 VSUBS 0.0166f
C474 VTAIL.n226 VSUBS 0.221589f
C475 VTAIL.t9 VSUBS 0.079467f
C476 VTAIL.n227 VSUBS 0.027793f
C477 VTAIL.n228 VSUBS 0.023574f
C478 VTAIL.n229 VSUBS 0.015678f
C479 VTAIL.n230 VSUBS 2.10801f
C480 VTAIL.n231 VSUBS 0.029176f
C481 VTAIL.n232 VSUBS 0.015678f
C482 VTAIL.n233 VSUBS 0.0166f
C483 VTAIL.n234 VSUBS 0.037057f
C484 VTAIL.n235 VSUBS 0.037057f
C485 VTAIL.n236 VSUBS 0.0166f
C486 VTAIL.n237 VSUBS 0.015678f
C487 VTAIL.n238 VSUBS 0.029176f
C488 VTAIL.n239 VSUBS 0.029176f
C489 VTAIL.n240 VSUBS 0.015678f
C490 VTAIL.n241 VSUBS 0.0166f
C491 VTAIL.n242 VSUBS 0.037057f
C492 VTAIL.n243 VSUBS 0.037057f
C493 VTAIL.n244 VSUBS 0.0166f
C494 VTAIL.n245 VSUBS 0.015678f
C495 VTAIL.n246 VSUBS 0.029176f
C496 VTAIL.n247 VSUBS 0.029176f
C497 VTAIL.n248 VSUBS 0.015678f
C498 VTAIL.n249 VSUBS 0.0166f
C499 VTAIL.n250 VSUBS 0.037057f
C500 VTAIL.n251 VSUBS 0.037057f
C501 VTAIL.n252 VSUBS 0.0166f
C502 VTAIL.n253 VSUBS 0.015678f
C503 VTAIL.n254 VSUBS 0.029176f
C504 VTAIL.n255 VSUBS 0.029176f
C505 VTAIL.n256 VSUBS 0.015678f
C506 VTAIL.n257 VSUBS 0.0166f
C507 VTAIL.n258 VSUBS 0.037057f
C508 VTAIL.n259 VSUBS 0.037057f
C509 VTAIL.n260 VSUBS 0.0166f
C510 VTAIL.n261 VSUBS 0.015678f
C511 VTAIL.n262 VSUBS 0.029176f
C512 VTAIL.n263 VSUBS 0.029176f
C513 VTAIL.n264 VSUBS 0.015678f
C514 VTAIL.n265 VSUBS 0.0166f
C515 VTAIL.n266 VSUBS 0.037057f
C516 VTAIL.n267 VSUBS 0.037057f
C517 VTAIL.n268 VSUBS 0.0166f
C518 VTAIL.n269 VSUBS 0.015678f
C519 VTAIL.n270 VSUBS 0.029176f
C520 VTAIL.n271 VSUBS 0.029176f
C521 VTAIL.n272 VSUBS 0.015678f
C522 VTAIL.n273 VSUBS 0.016139f
C523 VTAIL.n274 VSUBS 0.016139f
C524 VTAIL.n275 VSUBS 0.037057f
C525 VTAIL.n276 VSUBS 0.037057f
C526 VTAIL.n277 VSUBS 0.0166f
C527 VTAIL.n278 VSUBS 0.015678f
C528 VTAIL.n279 VSUBS 0.029176f
C529 VTAIL.n280 VSUBS 0.029176f
C530 VTAIL.n281 VSUBS 0.015678f
C531 VTAIL.n282 VSUBS 0.0166f
C532 VTAIL.n283 VSUBS 0.037057f
C533 VTAIL.n284 VSUBS 0.088033f
C534 VTAIL.n285 VSUBS 0.0166f
C535 VTAIL.n286 VSUBS 0.015678f
C536 VTAIL.n287 VSUBS 0.069433f
C537 VTAIL.n288 VSUBS 0.044257f
C538 VTAIL.n289 VSUBS 1.9355f
C539 VTAIL.n290 VSUBS 0.031566f
C540 VTAIL.n291 VSUBS 0.029176f
C541 VTAIL.n292 VSUBS 0.015678f
C542 VTAIL.n293 VSUBS 0.037057f
C543 VTAIL.n294 VSUBS 0.0166f
C544 VTAIL.n295 VSUBS 0.029176f
C545 VTAIL.n296 VSUBS 0.015678f
C546 VTAIL.n297 VSUBS 0.037057f
C547 VTAIL.n298 VSUBS 0.0166f
C548 VTAIL.n299 VSUBS 0.029176f
C549 VTAIL.n300 VSUBS 0.015678f
C550 VTAIL.n301 VSUBS 0.037057f
C551 VTAIL.n302 VSUBS 0.0166f
C552 VTAIL.n303 VSUBS 0.029176f
C553 VTAIL.n304 VSUBS 0.015678f
C554 VTAIL.n305 VSUBS 0.037057f
C555 VTAIL.n306 VSUBS 0.0166f
C556 VTAIL.n307 VSUBS 0.029176f
C557 VTAIL.n308 VSUBS 0.015678f
C558 VTAIL.n309 VSUBS 0.037057f
C559 VTAIL.n310 VSUBS 0.0166f
C560 VTAIL.n311 VSUBS 0.029176f
C561 VTAIL.n312 VSUBS 0.015678f
C562 VTAIL.n313 VSUBS 0.037057f
C563 VTAIL.n314 VSUBS 0.0166f
C564 VTAIL.n315 VSUBS 0.029176f
C565 VTAIL.n316 VSUBS 0.015678f
C566 VTAIL.n317 VSUBS 0.037057f
C567 VTAIL.n318 VSUBS 0.0166f
C568 VTAIL.n319 VSUBS 0.221589f
C569 VTAIL.t0 VSUBS 0.079467f
C570 VTAIL.n320 VSUBS 0.027793f
C571 VTAIL.n321 VSUBS 0.023574f
C572 VTAIL.n322 VSUBS 0.015678f
C573 VTAIL.n323 VSUBS 2.10801f
C574 VTAIL.n324 VSUBS 0.029176f
C575 VTAIL.n325 VSUBS 0.015678f
C576 VTAIL.n326 VSUBS 0.0166f
C577 VTAIL.n327 VSUBS 0.037057f
C578 VTAIL.n328 VSUBS 0.037057f
C579 VTAIL.n329 VSUBS 0.0166f
C580 VTAIL.n330 VSUBS 0.015678f
C581 VTAIL.n331 VSUBS 0.029176f
C582 VTAIL.n332 VSUBS 0.029176f
C583 VTAIL.n333 VSUBS 0.015678f
C584 VTAIL.n334 VSUBS 0.0166f
C585 VTAIL.n335 VSUBS 0.037057f
C586 VTAIL.n336 VSUBS 0.037057f
C587 VTAIL.n337 VSUBS 0.0166f
C588 VTAIL.n338 VSUBS 0.015678f
C589 VTAIL.n339 VSUBS 0.029176f
C590 VTAIL.n340 VSUBS 0.029176f
C591 VTAIL.n341 VSUBS 0.015678f
C592 VTAIL.n342 VSUBS 0.0166f
C593 VTAIL.n343 VSUBS 0.037057f
C594 VTAIL.n344 VSUBS 0.037057f
C595 VTAIL.n345 VSUBS 0.0166f
C596 VTAIL.n346 VSUBS 0.015678f
C597 VTAIL.n347 VSUBS 0.029176f
C598 VTAIL.n348 VSUBS 0.029176f
C599 VTAIL.n349 VSUBS 0.015678f
C600 VTAIL.n350 VSUBS 0.0166f
C601 VTAIL.n351 VSUBS 0.037057f
C602 VTAIL.n352 VSUBS 0.037057f
C603 VTAIL.n353 VSUBS 0.0166f
C604 VTAIL.n354 VSUBS 0.015678f
C605 VTAIL.n355 VSUBS 0.029176f
C606 VTAIL.n356 VSUBS 0.029176f
C607 VTAIL.n357 VSUBS 0.015678f
C608 VTAIL.n358 VSUBS 0.0166f
C609 VTAIL.n359 VSUBS 0.037057f
C610 VTAIL.n360 VSUBS 0.037057f
C611 VTAIL.n361 VSUBS 0.037057f
C612 VTAIL.n362 VSUBS 0.0166f
C613 VTAIL.n363 VSUBS 0.015678f
C614 VTAIL.n364 VSUBS 0.029176f
C615 VTAIL.n365 VSUBS 0.029176f
C616 VTAIL.n366 VSUBS 0.015678f
C617 VTAIL.n367 VSUBS 0.016139f
C618 VTAIL.n368 VSUBS 0.016139f
C619 VTAIL.n369 VSUBS 0.037057f
C620 VTAIL.n370 VSUBS 0.037057f
C621 VTAIL.n371 VSUBS 0.0166f
C622 VTAIL.n372 VSUBS 0.015678f
C623 VTAIL.n373 VSUBS 0.029176f
C624 VTAIL.n374 VSUBS 0.029176f
C625 VTAIL.n375 VSUBS 0.015678f
C626 VTAIL.n376 VSUBS 0.0166f
C627 VTAIL.n377 VSUBS 0.037057f
C628 VTAIL.n378 VSUBS 0.088033f
C629 VTAIL.n379 VSUBS 0.0166f
C630 VTAIL.n380 VSUBS 0.015678f
C631 VTAIL.n381 VSUBS 0.069433f
C632 VTAIL.n382 VSUBS 0.044257f
C633 VTAIL.n383 VSUBS 1.91159f
C634 VDD1.n0 VSUBS 0.028872f
C635 VDD1.n1 VSUBS 0.026686f
C636 VDD1.n2 VSUBS 0.01434f
C637 VDD1.n3 VSUBS 0.033895f
C638 VDD1.n4 VSUBS 0.015184f
C639 VDD1.n5 VSUBS 0.026686f
C640 VDD1.n6 VSUBS 0.01434f
C641 VDD1.n7 VSUBS 0.033895f
C642 VDD1.n8 VSUBS 0.015184f
C643 VDD1.n9 VSUBS 0.026686f
C644 VDD1.n10 VSUBS 0.01434f
C645 VDD1.n11 VSUBS 0.033895f
C646 VDD1.n12 VSUBS 0.033895f
C647 VDD1.n13 VSUBS 0.015184f
C648 VDD1.n14 VSUBS 0.026686f
C649 VDD1.n15 VSUBS 0.01434f
C650 VDD1.n16 VSUBS 0.033895f
C651 VDD1.n17 VSUBS 0.015184f
C652 VDD1.n18 VSUBS 0.026686f
C653 VDD1.n19 VSUBS 0.01434f
C654 VDD1.n20 VSUBS 0.033895f
C655 VDD1.n21 VSUBS 0.015184f
C656 VDD1.n22 VSUBS 0.026686f
C657 VDD1.n23 VSUBS 0.01434f
C658 VDD1.n24 VSUBS 0.033895f
C659 VDD1.n25 VSUBS 0.015184f
C660 VDD1.n26 VSUBS 0.026686f
C661 VDD1.n27 VSUBS 0.01434f
C662 VDD1.n28 VSUBS 0.033895f
C663 VDD1.n29 VSUBS 0.015184f
C664 VDD1.n30 VSUBS 0.202678f
C665 VDD1.t0 VSUBS 0.072685f
C666 VDD1.n31 VSUBS 0.025421f
C667 VDD1.n32 VSUBS 0.021562f
C668 VDD1.n33 VSUBS 0.01434f
C669 VDD1.n34 VSUBS 1.92811f
C670 VDD1.n35 VSUBS 0.026686f
C671 VDD1.n36 VSUBS 0.01434f
C672 VDD1.n37 VSUBS 0.015184f
C673 VDD1.n38 VSUBS 0.033895f
C674 VDD1.n39 VSUBS 0.033895f
C675 VDD1.n40 VSUBS 0.015184f
C676 VDD1.n41 VSUBS 0.01434f
C677 VDD1.n42 VSUBS 0.026686f
C678 VDD1.n43 VSUBS 0.026686f
C679 VDD1.n44 VSUBS 0.01434f
C680 VDD1.n45 VSUBS 0.015184f
C681 VDD1.n46 VSUBS 0.033895f
C682 VDD1.n47 VSUBS 0.033895f
C683 VDD1.n48 VSUBS 0.015184f
C684 VDD1.n49 VSUBS 0.01434f
C685 VDD1.n50 VSUBS 0.026686f
C686 VDD1.n51 VSUBS 0.026686f
C687 VDD1.n52 VSUBS 0.01434f
C688 VDD1.n53 VSUBS 0.015184f
C689 VDD1.n54 VSUBS 0.033895f
C690 VDD1.n55 VSUBS 0.033895f
C691 VDD1.n56 VSUBS 0.015184f
C692 VDD1.n57 VSUBS 0.01434f
C693 VDD1.n58 VSUBS 0.026686f
C694 VDD1.n59 VSUBS 0.026686f
C695 VDD1.n60 VSUBS 0.01434f
C696 VDD1.n61 VSUBS 0.015184f
C697 VDD1.n62 VSUBS 0.033895f
C698 VDD1.n63 VSUBS 0.033895f
C699 VDD1.n64 VSUBS 0.015184f
C700 VDD1.n65 VSUBS 0.01434f
C701 VDD1.n66 VSUBS 0.026686f
C702 VDD1.n67 VSUBS 0.026686f
C703 VDD1.n68 VSUBS 0.01434f
C704 VDD1.n69 VSUBS 0.015184f
C705 VDD1.n70 VSUBS 0.033895f
C706 VDD1.n71 VSUBS 0.033895f
C707 VDD1.n72 VSUBS 0.015184f
C708 VDD1.n73 VSUBS 0.01434f
C709 VDD1.n74 VSUBS 0.026686f
C710 VDD1.n75 VSUBS 0.026686f
C711 VDD1.n76 VSUBS 0.01434f
C712 VDD1.n77 VSUBS 0.014762f
C713 VDD1.n78 VSUBS 0.014762f
C714 VDD1.n79 VSUBS 0.033895f
C715 VDD1.n80 VSUBS 0.033895f
C716 VDD1.n81 VSUBS 0.015184f
C717 VDD1.n82 VSUBS 0.01434f
C718 VDD1.n83 VSUBS 0.026686f
C719 VDD1.n84 VSUBS 0.026686f
C720 VDD1.n85 VSUBS 0.01434f
C721 VDD1.n86 VSUBS 0.015184f
C722 VDD1.n87 VSUBS 0.033895f
C723 VDD1.n88 VSUBS 0.08052f
C724 VDD1.n89 VSUBS 0.015184f
C725 VDD1.n90 VSUBS 0.01434f
C726 VDD1.n91 VSUBS 0.063507f
C727 VDD1.n92 VSUBS 0.060276f
C728 VDD1.n93 VSUBS 0.028872f
C729 VDD1.n94 VSUBS 0.026686f
C730 VDD1.n95 VSUBS 0.01434f
C731 VDD1.n96 VSUBS 0.033895f
C732 VDD1.n97 VSUBS 0.015184f
C733 VDD1.n98 VSUBS 0.026686f
C734 VDD1.n99 VSUBS 0.01434f
C735 VDD1.n100 VSUBS 0.033895f
C736 VDD1.n101 VSUBS 0.015184f
C737 VDD1.n102 VSUBS 0.026686f
C738 VDD1.n103 VSUBS 0.01434f
C739 VDD1.n104 VSUBS 0.033895f
C740 VDD1.n105 VSUBS 0.015184f
C741 VDD1.n106 VSUBS 0.026686f
C742 VDD1.n107 VSUBS 0.01434f
C743 VDD1.n108 VSUBS 0.033895f
C744 VDD1.n109 VSUBS 0.015184f
C745 VDD1.n110 VSUBS 0.026686f
C746 VDD1.n111 VSUBS 0.01434f
C747 VDD1.n112 VSUBS 0.033895f
C748 VDD1.n113 VSUBS 0.015184f
C749 VDD1.n114 VSUBS 0.026686f
C750 VDD1.n115 VSUBS 0.01434f
C751 VDD1.n116 VSUBS 0.033895f
C752 VDD1.n117 VSUBS 0.015184f
C753 VDD1.n118 VSUBS 0.026686f
C754 VDD1.n119 VSUBS 0.01434f
C755 VDD1.n120 VSUBS 0.033895f
C756 VDD1.n121 VSUBS 0.015184f
C757 VDD1.n122 VSUBS 0.202678f
C758 VDD1.t1 VSUBS 0.072685f
C759 VDD1.n123 VSUBS 0.025421f
C760 VDD1.n124 VSUBS 0.021562f
C761 VDD1.n125 VSUBS 0.01434f
C762 VDD1.n126 VSUBS 1.92811f
C763 VDD1.n127 VSUBS 0.026686f
C764 VDD1.n128 VSUBS 0.01434f
C765 VDD1.n129 VSUBS 0.015184f
C766 VDD1.n130 VSUBS 0.033895f
C767 VDD1.n131 VSUBS 0.033895f
C768 VDD1.n132 VSUBS 0.015184f
C769 VDD1.n133 VSUBS 0.01434f
C770 VDD1.n134 VSUBS 0.026686f
C771 VDD1.n135 VSUBS 0.026686f
C772 VDD1.n136 VSUBS 0.01434f
C773 VDD1.n137 VSUBS 0.015184f
C774 VDD1.n138 VSUBS 0.033895f
C775 VDD1.n139 VSUBS 0.033895f
C776 VDD1.n140 VSUBS 0.015184f
C777 VDD1.n141 VSUBS 0.01434f
C778 VDD1.n142 VSUBS 0.026686f
C779 VDD1.n143 VSUBS 0.026686f
C780 VDD1.n144 VSUBS 0.01434f
C781 VDD1.n145 VSUBS 0.015184f
C782 VDD1.n146 VSUBS 0.033895f
C783 VDD1.n147 VSUBS 0.033895f
C784 VDD1.n148 VSUBS 0.015184f
C785 VDD1.n149 VSUBS 0.01434f
C786 VDD1.n150 VSUBS 0.026686f
C787 VDD1.n151 VSUBS 0.026686f
C788 VDD1.n152 VSUBS 0.01434f
C789 VDD1.n153 VSUBS 0.015184f
C790 VDD1.n154 VSUBS 0.033895f
C791 VDD1.n155 VSUBS 0.033895f
C792 VDD1.n156 VSUBS 0.015184f
C793 VDD1.n157 VSUBS 0.01434f
C794 VDD1.n158 VSUBS 0.026686f
C795 VDD1.n159 VSUBS 0.026686f
C796 VDD1.n160 VSUBS 0.01434f
C797 VDD1.n161 VSUBS 0.015184f
C798 VDD1.n162 VSUBS 0.033895f
C799 VDD1.n163 VSUBS 0.033895f
C800 VDD1.n164 VSUBS 0.033895f
C801 VDD1.n165 VSUBS 0.015184f
C802 VDD1.n166 VSUBS 0.01434f
C803 VDD1.n167 VSUBS 0.026686f
C804 VDD1.n168 VSUBS 0.026686f
C805 VDD1.n169 VSUBS 0.01434f
C806 VDD1.n170 VSUBS 0.014762f
C807 VDD1.n171 VSUBS 0.014762f
C808 VDD1.n172 VSUBS 0.033895f
C809 VDD1.n173 VSUBS 0.033895f
C810 VDD1.n174 VSUBS 0.015184f
C811 VDD1.n175 VSUBS 0.01434f
C812 VDD1.n176 VSUBS 0.026686f
C813 VDD1.n177 VSUBS 0.026686f
C814 VDD1.n178 VSUBS 0.01434f
C815 VDD1.n179 VSUBS 0.015184f
C816 VDD1.n180 VSUBS 0.033895f
C817 VDD1.n181 VSUBS 0.08052f
C818 VDD1.n182 VSUBS 0.015184f
C819 VDD1.n183 VSUBS 0.01434f
C820 VDD1.n184 VSUBS 0.063507f
C821 VDD1.n185 VSUBS 0.059944f
C822 VDD1.t2 VSUBS 0.35534f
C823 VDD1.t4 VSUBS 0.35534f
C824 VDD1.n186 VSUBS 2.93287f
C825 VDD1.n187 VSUBS 2.61899f
C826 VDD1.t3 VSUBS 0.35534f
C827 VDD1.t5 VSUBS 0.35534f
C828 VDD1.n188 VSUBS 2.93164f
C829 VDD1.n189 VSUBS 3.06571f
C830 VP.n0 VSUBS 0.078228f
C831 VP.t4 VSUBS 1.65083f
C832 VP.n1 VSUBS 0.60326f
C833 VP.t2 VSUBS 1.62981f
C834 VP.t0 VSUBS 1.62981f
C835 VP.n2 VSUBS 0.636375f
C836 VP.n3 VSUBS 0.623041f
C837 VP.n4 VSUBS 2.85313f
C838 VP.n5 VSUBS 2.73073f
C839 VP.t5 VSUBS 1.62981f
C840 VP.n6 VSUBS 0.623041f
C841 VP.t1 VSUBS 1.62981f
C842 VP.n7 VSUBS 0.636375f
C843 VP.t3 VSUBS 1.62981f
C844 VP.n8 VSUBS 0.623041f
C845 VP.n9 VSUBS 0.065188f
C846 B.n0 VSUBS 0.004424f
C847 B.n1 VSUBS 0.004424f
C848 B.n2 VSUBS 0.006997f
C849 B.n3 VSUBS 0.006997f
C850 B.n4 VSUBS 0.006997f
C851 B.n5 VSUBS 0.006997f
C852 B.n6 VSUBS 0.006997f
C853 B.n7 VSUBS 0.006997f
C854 B.n8 VSUBS 0.006997f
C855 B.n9 VSUBS 0.006997f
C856 B.n10 VSUBS 0.006997f
C857 B.n11 VSUBS 0.016104f
C858 B.n12 VSUBS 0.006997f
C859 B.n13 VSUBS 0.006997f
C860 B.n14 VSUBS 0.006997f
C861 B.n15 VSUBS 0.006997f
C862 B.n16 VSUBS 0.006997f
C863 B.n17 VSUBS 0.006997f
C864 B.n18 VSUBS 0.006997f
C865 B.n19 VSUBS 0.006997f
C866 B.n20 VSUBS 0.006997f
C867 B.n21 VSUBS 0.006997f
C868 B.n22 VSUBS 0.006997f
C869 B.n23 VSUBS 0.006997f
C870 B.n24 VSUBS 0.006997f
C871 B.n25 VSUBS 0.006997f
C872 B.n26 VSUBS 0.006997f
C873 B.n27 VSUBS 0.006997f
C874 B.n28 VSUBS 0.006997f
C875 B.n29 VSUBS 0.006997f
C876 B.n30 VSUBS 0.006997f
C877 B.n31 VSUBS 0.006997f
C878 B.n32 VSUBS 0.006997f
C879 B.n33 VSUBS 0.006997f
C880 B.n34 VSUBS 0.006997f
C881 B.n35 VSUBS 0.006997f
C882 B.n36 VSUBS 0.006997f
C883 B.n37 VSUBS 0.006997f
C884 B.n38 VSUBS 0.006997f
C885 B.n39 VSUBS 0.006997f
C886 B.t11 VSUBS 0.323285f
C887 B.t10 VSUBS 0.334164f
C888 B.t9 VSUBS 0.390878f
C889 B.n40 VSUBS 0.398047f
C890 B.n41 VSUBS 0.306261f
C891 B.n42 VSUBS 0.006997f
C892 B.n43 VSUBS 0.006997f
C893 B.n44 VSUBS 0.006997f
C894 B.n45 VSUBS 0.006997f
C895 B.t8 VSUBS 0.323288f
C896 B.t7 VSUBS 0.334167f
C897 B.t6 VSUBS 0.390878f
C898 B.n46 VSUBS 0.398044f
C899 B.n47 VSUBS 0.306258f
C900 B.n48 VSUBS 0.016211f
C901 B.n49 VSUBS 0.006997f
C902 B.n50 VSUBS 0.006997f
C903 B.n51 VSUBS 0.006997f
C904 B.n52 VSUBS 0.006997f
C905 B.n53 VSUBS 0.006997f
C906 B.n54 VSUBS 0.006997f
C907 B.n55 VSUBS 0.006997f
C908 B.n56 VSUBS 0.006997f
C909 B.n57 VSUBS 0.006997f
C910 B.n58 VSUBS 0.006997f
C911 B.n59 VSUBS 0.006997f
C912 B.n60 VSUBS 0.006997f
C913 B.n61 VSUBS 0.006997f
C914 B.n62 VSUBS 0.006997f
C915 B.n63 VSUBS 0.006997f
C916 B.n64 VSUBS 0.006997f
C917 B.n65 VSUBS 0.006997f
C918 B.n66 VSUBS 0.006997f
C919 B.n67 VSUBS 0.006997f
C920 B.n68 VSUBS 0.006997f
C921 B.n69 VSUBS 0.006997f
C922 B.n70 VSUBS 0.006997f
C923 B.n71 VSUBS 0.006997f
C924 B.n72 VSUBS 0.006997f
C925 B.n73 VSUBS 0.006997f
C926 B.n74 VSUBS 0.006997f
C927 B.n75 VSUBS 0.006997f
C928 B.n76 VSUBS 0.015574f
C929 B.n77 VSUBS 0.006997f
C930 B.n78 VSUBS 0.006997f
C931 B.n79 VSUBS 0.006997f
C932 B.n80 VSUBS 0.006997f
C933 B.n81 VSUBS 0.006997f
C934 B.n82 VSUBS 0.006997f
C935 B.n83 VSUBS 0.006997f
C936 B.n84 VSUBS 0.006997f
C937 B.n85 VSUBS 0.006997f
C938 B.n86 VSUBS 0.006997f
C939 B.n87 VSUBS 0.006997f
C940 B.n88 VSUBS 0.006997f
C941 B.n89 VSUBS 0.006997f
C942 B.n90 VSUBS 0.006997f
C943 B.n91 VSUBS 0.006997f
C944 B.n92 VSUBS 0.006997f
C945 B.n93 VSUBS 0.006997f
C946 B.n94 VSUBS 0.006997f
C947 B.n95 VSUBS 0.006997f
C948 B.n96 VSUBS 0.01641f
C949 B.n97 VSUBS 0.006997f
C950 B.n98 VSUBS 0.006997f
C951 B.n99 VSUBS 0.006997f
C952 B.n100 VSUBS 0.006997f
C953 B.n101 VSUBS 0.006997f
C954 B.n102 VSUBS 0.006997f
C955 B.n103 VSUBS 0.006997f
C956 B.n104 VSUBS 0.006997f
C957 B.n105 VSUBS 0.006997f
C958 B.n106 VSUBS 0.006997f
C959 B.n107 VSUBS 0.006997f
C960 B.n108 VSUBS 0.006997f
C961 B.n109 VSUBS 0.006997f
C962 B.n110 VSUBS 0.006997f
C963 B.n111 VSUBS 0.006997f
C964 B.n112 VSUBS 0.006997f
C965 B.n113 VSUBS 0.006997f
C966 B.n114 VSUBS 0.006997f
C967 B.n115 VSUBS 0.006997f
C968 B.n116 VSUBS 0.006997f
C969 B.n117 VSUBS 0.006997f
C970 B.n118 VSUBS 0.006997f
C971 B.n119 VSUBS 0.006997f
C972 B.n120 VSUBS 0.006997f
C973 B.n121 VSUBS 0.006997f
C974 B.n122 VSUBS 0.006997f
C975 B.n123 VSUBS 0.006997f
C976 B.t4 VSUBS 0.323288f
C977 B.t5 VSUBS 0.334167f
C978 B.t3 VSUBS 0.390878f
C979 B.n124 VSUBS 0.398044f
C980 B.n125 VSUBS 0.306258f
C981 B.n126 VSUBS 0.016211f
C982 B.n127 VSUBS 0.006997f
C983 B.n128 VSUBS 0.006997f
C984 B.n129 VSUBS 0.006997f
C985 B.n130 VSUBS 0.006997f
C986 B.n131 VSUBS 0.006997f
C987 B.t1 VSUBS 0.323285f
C988 B.t2 VSUBS 0.334164f
C989 B.t0 VSUBS 0.390878f
C990 B.n132 VSUBS 0.398047f
C991 B.n133 VSUBS 0.306261f
C992 B.n134 VSUBS 0.006997f
C993 B.n135 VSUBS 0.006997f
C994 B.n136 VSUBS 0.006997f
C995 B.n137 VSUBS 0.006997f
C996 B.n138 VSUBS 0.006997f
C997 B.n139 VSUBS 0.006997f
C998 B.n140 VSUBS 0.006997f
C999 B.n141 VSUBS 0.006997f
C1000 B.n142 VSUBS 0.006997f
C1001 B.n143 VSUBS 0.006997f
C1002 B.n144 VSUBS 0.006997f
C1003 B.n145 VSUBS 0.006997f
C1004 B.n146 VSUBS 0.006997f
C1005 B.n147 VSUBS 0.006997f
C1006 B.n148 VSUBS 0.006997f
C1007 B.n149 VSUBS 0.006997f
C1008 B.n150 VSUBS 0.006997f
C1009 B.n151 VSUBS 0.006997f
C1010 B.n152 VSUBS 0.006997f
C1011 B.n153 VSUBS 0.006997f
C1012 B.n154 VSUBS 0.006997f
C1013 B.n155 VSUBS 0.006997f
C1014 B.n156 VSUBS 0.006997f
C1015 B.n157 VSUBS 0.006997f
C1016 B.n158 VSUBS 0.006997f
C1017 B.n159 VSUBS 0.006997f
C1018 B.n160 VSUBS 0.006997f
C1019 B.n161 VSUBS 0.016104f
C1020 B.n162 VSUBS 0.006997f
C1021 B.n163 VSUBS 0.006997f
C1022 B.n164 VSUBS 0.006997f
C1023 B.n165 VSUBS 0.006997f
C1024 B.n166 VSUBS 0.006997f
C1025 B.n167 VSUBS 0.006997f
C1026 B.n168 VSUBS 0.006997f
C1027 B.n169 VSUBS 0.006997f
C1028 B.n170 VSUBS 0.006997f
C1029 B.n171 VSUBS 0.006997f
C1030 B.n172 VSUBS 0.006997f
C1031 B.n173 VSUBS 0.006997f
C1032 B.n174 VSUBS 0.006997f
C1033 B.n175 VSUBS 0.006997f
C1034 B.n176 VSUBS 0.006997f
C1035 B.n177 VSUBS 0.006997f
C1036 B.n178 VSUBS 0.006997f
C1037 B.n179 VSUBS 0.006997f
C1038 B.n180 VSUBS 0.006997f
C1039 B.n181 VSUBS 0.006997f
C1040 B.n182 VSUBS 0.006997f
C1041 B.n183 VSUBS 0.006997f
C1042 B.n184 VSUBS 0.006997f
C1043 B.n185 VSUBS 0.006997f
C1044 B.n186 VSUBS 0.006997f
C1045 B.n187 VSUBS 0.006997f
C1046 B.n188 VSUBS 0.006997f
C1047 B.n189 VSUBS 0.006997f
C1048 B.n190 VSUBS 0.006997f
C1049 B.n191 VSUBS 0.006997f
C1050 B.n192 VSUBS 0.006997f
C1051 B.n193 VSUBS 0.006997f
C1052 B.n194 VSUBS 0.006997f
C1053 B.n195 VSUBS 0.006997f
C1054 B.n196 VSUBS 0.016104f
C1055 B.n197 VSUBS 0.01641f
C1056 B.n198 VSUBS 0.01641f
C1057 B.n199 VSUBS 0.006997f
C1058 B.n200 VSUBS 0.006997f
C1059 B.n201 VSUBS 0.006997f
C1060 B.n202 VSUBS 0.006997f
C1061 B.n203 VSUBS 0.006997f
C1062 B.n204 VSUBS 0.006997f
C1063 B.n205 VSUBS 0.006997f
C1064 B.n206 VSUBS 0.006997f
C1065 B.n207 VSUBS 0.006997f
C1066 B.n208 VSUBS 0.006997f
C1067 B.n209 VSUBS 0.006997f
C1068 B.n210 VSUBS 0.006997f
C1069 B.n211 VSUBS 0.006997f
C1070 B.n212 VSUBS 0.006997f
C1071 B.n213 VSUBS 0.006997f
C1072 B.n214 VSUBS 0.006997f
C1073 B.n215 VSUBS 0.006997f
C1074 B.n216 VSUBS 0.006997f
C1075 B.n217 VSUBS 0.006997f
C1076 B.n218 VSUBS 0.006997f
C1077 B.n219 VSUBS 0.006997f
C1078 B.n220 VSUBS 0.006997f
C1079 B.n221 VSUBS 0.006997f
C1080 B.n222 VSUBS 0.006997f
C1081 B.n223 VSUBS 0.006997f
C1082 B.n224 VSUBS 0.006997f
C1083 B.n225 VSUBS 0.006997f
C1084 B.n226 VSUBS 0.006997f
C1085 B.n227 VSUBS 0.006997f
C1086 B.n228 VSUBS 0.006997f
C1087 B.n229 VSUBS 0.006997f
C1088 B.n230 VSUBS 0.006997f
C1089 B.n231 VSUBS 0.006997f
C1090 B.n232 VSUBS 0.006997f
C1091 B.n233 VSUBS 0.006997f
C1092 B.n234 VSUBS 0.006997f
C1093 B.n235 VSUBS 0.006997f
C1094 B.n236 VSUBS 0.006997f
C1095 B.n237 VSUBS 0.006997f
C1096 B.n238 VSUBS 0.006997f
C1097 B.n239 VSUBS 0.006997f
C1098 B.n240 VSUBS 0.006997f
C1099 B.n241 VSUBS 0.006997f
C1100 B.n242 VSUBS 0.006997f
C1101 B.n243 VSUBS 0.006997f
C1102 B.n244 VSUBS 0.006997f
C1103 B.n245 VSUBS 0.006997f
C1104 B.n246 VSUBS 0.006997f
C1105 B.n247 VSUBS 0.006997f
C1106 B.n248 VSUBS 0.006997f
C1107 B.n249 VSUBS 0.006997f
C1108 B.n250 VSUBS 0.006997f
C1109 B.n251 VSUBS 0.006997f
C1110 B.n252 VSUBS 0.006997f
C1111 B.n253 VSUBS 0.006997f
C1112 B.n254 VSUBS 0.006997f
C1113 B.n255 VSUBS 0.006997f
C1114 B.n256 VSUBS 0.006997f
C1115 B.n257 VSUBS 0.006997f
C1116 B.n258 VSUBS 0.006997f
C1117 B.n259 VSUBS 0.006997f
C1118 B.n260 VSUBS 0.006997f
C1119 B.n261 VSUBS 0.006997f
C1120 B.n262 VSUBS 0.006997f
C1121 B.n263 VSUBS 0.006997f
C1122 B.n264 VSUBS 0.006997f
C1123 B.n265 VSUBS 0.006997f
C1124 B.n266 VSUBS 0.006997f
C1125 B.n267 VSUBS 0.006997f
C1126 B.n268 VSUBS 0.006997f
C1127 B.n269 VSUBS 0.006997f
C1128 B.n270 VSUBS 0.006997f
C1129 B.n271 VSUBS 0.006997f
C1130 B.n272 VSUBS 0.006997f
C1131 B.n273 VSUBS 0.006997f
C1132 B.n274 VSUBS 0.006997f
C1133 B.n275 VSUBS 0.006997f
C1134 B.n276 VSUBS 0.006997f
C1135 B.n277 VSUBS 0.006997f
C1136 B.n278 VSUBS 0.006997f
C1137 B.n279 VSUBS 0.006997f
C1138 B.n280 VSUBS 0.004836f
C1139 B.n281 VSUBS 0.016211f
C1140 B.n282 VSUBS 0.005659f
C1141 B.n283 VSUBS 0.006997f
C1142 B.n284 VSUBS 0.006997f
C1143 B.n285 VSUBS 0.006997f
C1144 B.n286 VSUBS 0.006997f
C1145 B.n287 VSUBS 0.006997f
C1146 B.n288 VSUBS 0.006997f
C1147 B.n289 VSUBS 0.006997f
C1148 B.n290 VSUBS 0.006997f
C1149 B.n291 VSUBS 0.006997f
C1150 B.n292 VSUBS 0.006997f
C1151 B.n293 VSUBS 0.006997f
C1152 B.n294 VSUBS 0.005659f
C1153 B.n295 VSUBS 0.006997f
C1154 B.n296 VSUBS 0.006997f
C1155 B.n297 VSUBS 0.004836f
C1156 B.n298 VSUBS 0.006997f
C1157 B.n299 VSUBS 0.006997f
C1158 B.n300 VSUBS 0.006997f
C1159 B.n301 VSUBS 0.006997f
C1160 B.n302 VSUBS 0.006997f
C1161 B.n303 VSUBS 0.006997f
C1162 B.n304 VSUBS 0.006997f
C1163 B.n305 VSUBS 0.006997f
C1164 B.n306 VSUBS 0.006997f
C1165 B.n307 VSUBS 0.006997f
C1166 B.n308 VSUBS 0.006997f
C1167 B.n309 VSUBS 0.006997f
C1168 B.n310 VSUBS 0.006997f
C1169 B.n311 VSUBS 0.006997f
C1170 B.n312 VSUBS 0.006997f
C1171 B.n313 VSUBS 0.006997f
C1172 B.n314 VSUBS 0.006997f
C1173 B.n315 VSUBS 0.006997f
C1174 B.n316 VSUBS 0.006997f
C1175 B.n317 VSUBS 0.006997f
C1176 B.n318 VSUBS 0.006997f
C1177 B.n319 VSUBS 0.006997f
C1178 B.n320 VSUBS 0.006997f
C1179 B.n321 VSUBS 0.006997f
C1180 B.n322 VSUBS 0.006997f
C1181 B.n323 VSUBS 0.006997f
C1182 B.n324 VSUBS 0.006997f
C1183 B.n325 VSUBS 0.006997f
C1184 B.n326 VSUBS 0.006997f
C1185 B.n327 VSUBS 0.006997f
C1186 B.n328 VSUBS 0.006997f
C1187 B.n329 VSUBS 0.006997f
C1188 B.n330 VSUBS 0.006997f
C1189 B.n331 VSUBS 0.006997f
C1190 B.n332 VSUBS 0.006997f
C1191 B.n333 VSUBS 0.006997f
C1192 B.n334 VSUBS 0.006997f
C1193 B.n335 VSUBS 0.006997f
C1194 B.n336 VSUBS 0.006997f
C1195 B.n337 VSUBS 0.006997f
C1196 B.n338 VSUBS 0.006997f
C1197 B.n339 VSUBS 0.006997f
C1198 B.n340 VSUBS 0.006997f
C1199 B.n341 VSUBS 0.006997f
C1200 B.n342 VSUBS 0.006997f
C1201 B.n343 VSUBS 0.006997f
C1202 B.n344 VSUBS 0.006997f
C1203 B.n345 VSUBS 0.006997f
C1204 B.n346 VSUBS 0.006997f
C1205 B.n347 VSUBS 0.006997f
C1206 B.n348 VSUBS 0.006997f
C1207 B.n349 VSUBS 0.006997f
C1208 B.n350 VSUBS 0.006997f
C1209 B.n351 VSUBS 0.006997f
C1210 B.n352 VSUBS 0.006997f
C1211 B.n353 VSUBS 0.006997f
C1212 B.n354 VSUBS 0.006997f
C1213 B.n355 VSUBS 0.006997f
C1214 B.n356 VSUBS 0.006997f
C1215 B.n357 VSUBS 0.006997f
C1216 B.n358 VSUBS 0.006997f
C1217 B.n359 VSUBS 0.006997f
C1218 B.n360 VSUBS 0.006997f
C1219 B.n361 VSUBS 0.006997f
C1220 B.n362 VSUBS 0.006997f
C1221 B.n363 VSUBS 0.006997f
C1222 B.n364 VSUBS 0.006997f
C1223 B.n365 VSUBS 0.006997f
C1224 B.n366 VSUBS 0.006997f
C1225 B.n367 VSUBS 0.006997f
C1226 B.n368 VSUBS 0.006997f
C1227 B.n369 VSUBS 0.006997f
C1228 B.n370 VSUBS 0.006997f
C1229 B.n371 VSUBS 0.006997f
C1230 B.n372 VSUBS 0.006997f
C1231 B.n373 VSUBS 0.006997f
C1232 B.n374 VSUBS 0.006997f
C1233 B.n375 VSUBS 0.006997f
C1234 B.n376 VSUBS 0.006997f
C1235 B.n377 VSUBS 0.006997f
C1236 B.n378 VSUBS 0.006997f
C1237 B.n379 VSUBS 0.01641f
C1238 B.n380 VSUBS 0.016104f
C1239 B.n381 VSUBS 0.016104f
C1240 B.n382 VSUBS 0.006997f
C1241 B.n383 VSUBS 0.006997f
C1242 B.n384 VSUBS 0.006997f
C1243 B.n385 VSUBS 0.006997f
C1244 B.n386 VSUBS 0.006997f
C1245 B.n387 VSUBS 0.006997f
C1246 B.n388 VSUBS 0.006997f
C1247 B.n389 VSUBS 0.006997f
C1248 B.n390 VSUBS 0.006997f
C1249 B.n391 VSUBS 0.006997f
C1250 B.n392 VSUBS 0.006997f
C1251 B.n393 VSUBS 0.006997f
C1252 B.n394 VSUBS 0.006997f
C1253 B.n395 VSUBS 0.006997f
C1254 B.n396 VSUBS 0.006997f
C1255 B.n397 VSUBS 0.006997f
C1256 B.n398 VSUBS 0.006997f
C1257 B.n399 VSUBS 0.006997f
C1258 B.n400 VSUBS 0.006997f
C1259 B.n401 VSUBS 0.006997f
C1260 B.n402 VSUBS 0.006997f
C1261 B.n403 VSUBS 0.006997f
C1262 B.n404 VSUBS 0.006997f
C1263 B.n405 VSUBS 0.006997f
C1264 B.n406 VSUBS 0.006997f
C1265 B.n407 VSUBS 0.006997f
C1266 B.n408 VSUBS 0.006997f
C1267 B.n409 VSUBS 0.006997f
C1268 B.n410 VSUBS 0.006997f
C1269 B.n411 VSUBS 0.006997f
C1270 B.n412 VSUBS 0.006997f
C1271 B.n413 VSUBS 0.006997f
C1272 B.n414 VSUBS 0.006997f
C1273 B.n415 VSUBS 0.006997f
C1274 B.n416 VSUBS 0.006997f
C1275 B.n417 VSUBS 0.006997f
C1276 B.n418 VSUBS 0.006997f
C1277 B.n419 VSUBS 0.006997f
C1278 B.n420 VSUBS 0.006997f
C1279 B.n421 VSUBS 0.006997f
C1280 B.n422 VSUBS 0.006997f
C1281 B.n423 VSUBS 0.006997f
C1282 B.n424 VSUBS 0.006997f
C1283 B.n425 VSUBS 0.006997f
C1284 B.n426 VSUBS 0.006997f
C1285 B.n427 VSUBS 0.006997f
C1286 B.n428 VSUBS 0.006997f
C1287 B.n429 VSUBS 0.006997f
C1288 B.n430 VSUBS 0.006997f
C1289 B.n431 VSUBS 0.006997f
C1290 B.n432 VSUBS 0.006997f
C1291 B.n433 VSUBS 0.006997f
C1292 B.n434 VSUBS 0.006997f
C1293 B.n435 VSUBS 0.006997f
C1294 B.n436 VSUBS 0.006997f
C1295 B.n437 VSUBS 0.01694f
C1296 B.n438 VSUBS 0.016104f
C1297 B.n439 VSUBS 0.01641f
C1298 B.n440 VSUBS 0.006997f
C1299 B.n441 VSUBS 0.006997f
C1300 B.n442 VSUBS 0.006997f
C1301 B.n443 VSUBS 0.006997f
C1302 B.n444 VSUBS 0.006997f
C1303 B.n445 VSUBS 0.006997f
C1304 B.n446 VSUBS 0.006997f
C1305 B.n447 VSUBS 0.006997f
C1306 B.n448 VSUBS 0.006997f
C1307 B.n449 VSUBS 0.006997f
C1308 B.n450 VSUBS 0.006997f
C1309 B.n451 VSUBS 0.006997f
C1310 B.n452 VSUBS 0.006997f
C1311 B.n453 VSUBS 0.006997f
C1312 B.n454 VSUBS 0.006997f
C1313 B.n455 VSUBS 0.006997f
C1314 B.n456 VSUBS 0.006997f
C1315 B.n457 VSUBS 0.006997f
C1316 B.n458 VSUBS 0.006997f
C1317 B.n459 VSUBS 0.006997f
C1318 B.n460 VSUBS 0.006997f
C1319 B.n461 VSUBS 0.006997f
C1320 B.n462 VSUBS 0.006997f
C1321 B.n463 VSUBS 0.006997f
C1322 B.n464 VSUBS 0.006997f
C1323 B.n465 VSUBS 0.006997f
C1324 B.n466 VSUBS 0.006997f
C1325 B.n467 VSUBS 0.006997f
C1326 B.n468 VSUBS 0.006997f
C1327 B.n469 VSUBS 0.006997f
C1328 B.n470 VSUBS 0.006997f
C1329 B.n471 VSUBS 0.006997f
C1330 B.n472 VSUBS 0.006997f
C1331 B.n473 VSUBS 0.006997f
C1332 B.n474 VSUBS 0.006997f
C1333 B.n475 VSUBS 0.006997f
C1334 B.n476 VSUBS 0.006997f
C1335 B.n477 VSUBS 0.006997f
C1336 B.n478 VSUBS 0.006997f
C1337 B.n479 VSUBS 0.006997f
C1338 B.n480 VSUBS 0.006997f
C1339 B.n481 VSUBS 0.006997f
C1340 B.n482 VSUBS 0.006997f
C1341 B.n483 VSUBS 0.006997f
C1342 B.n484 VSUBS 0.006997f
C1343 B.n485 VSUBS 0.006997f
C1344 B.n486 VSUBS 0.006997f
C1345 B.n487 VSUBS 0.006997f
C1346 B.n488 VSUBS 0.006997f
C1347 B.n489 VSUBS 0.006997f
C1348 B.n490 VSUBS 0.006997f
C1349 B.n491 VSUBS 0.006997f
C1350 B.n492 VSUBS 0.006997f
C1351 B.n493 VSUBS 0.006997f
C1352 B.n494 VSUBS 0.006997f
C1353 B.n495 VSUBS 0.006997f
C1354 B.n496 VSUBS 0.006997f
C1355 B.n497 VSUBS 0.006997f
C1356 B.n498 VSUBS 0.006997f
C1357 B.n499 VSUBS 0.006997f
C1358 B.n500 VSUBS 0.006997f
C1359 B.n501 VSUBS 0.006997f
C1360 B.n502 VSUBS 0.006997f
C1361 B.n503 VSUBS 0.006997f
C1362 B.n504 VSUBS 0.006997f
C1363 B.n505 VSUBS 0.006997f
C1364 B.n506 VSUBS 0.006997f
C1365 B.n507 VSUBS 0.006997f
C1366 B.n508 VSUBS 0.006997f
C1367 B.n509 VSUBS 0.006997f
C1368 B.n510 VSUBS 0.006997f
C1369 B.n511 VSUBS 0.006997f
C1370 B.n512 VSUBS 0.006997f
C1371 B.n513 VSUBS 0.006997f
C1372 B.n514 VSUBS 0.006997f
C1373 B.n515 VSUBS 0.006997f
C1374 B.n516 VSUBS 0.006997f
C1375 B.n517 VSUBS 0.006997f
C1376 B.n518 VSUBS 0.006997f
C1377 B.n519 VSUBS 0.006997f
C1378 B.n520 VSUBS 0.006997f
C1379 B.n521 VSUBS 0.004836f
C1380 B.n522 VSUBS 0.006997f
C1381 B.n523 VSUBS 0.006997f
C1382 B.n524 VSUBS 0.005659f
C1383 B.n525 VSUBS 0.006997f
C1384 B.n526 VSUBS 0.006997f
C1385 B.n527 VSUBS 0.006997f
C1386 B.n528 VSUBS 0.006997f
C1387 B.n529 VSUBS 0.006997f
C1388 B.n530 VSUBS 0.006997f
C1389 B.n531 VSUBS 0.006997f
C1390 B.n532 VSUBS 0.006997f
C1391 B.n533 VSUBS 0.006997f
C1392 B.n534 VSUBS 0.006997f
C1393 B.n535 VSUBS 0.006997f
C1394 B.n536 VSUBS 0.005659f
C1395 B.n537 VSUBS 0.016211f
C1396 B.n538 VSUBS 0.004836f
C1397 B.n539 VSUBS 0.006997f
C1398 B.n540 VSUBS 0.006997f
C1399 B.n541 VSUBS 0.006997f
C1400 B.n542 VSUBS 0.006997f
C1401 B.n543 VSUBS 0.006997f
C1402 B.n544 VSUBS 0.006997f
C1403 B.n545 VSUBS 0.006997f
C1404 B.n546 VSUBS 0.006997f
C1405 B.n547 VSUBS 0.006997f
C1406 B.n548 VSUBS 0.006997f
C1407 B.n549 VSUBS 0.006997f
C1408 B.n550 VSUBS 0.006997f
C1409 B.n551 VSUBS 0.006997f
C1410 B.n552 VSUBS 0.006997f
C1411 B.n553 VSUBS 0.006997f
C1412 B.n554 VSUBS 0.006997f
C1413 B.n555 VSUBS 0.006997f
C1414 B.n556 VSUBS 0.006997f
C1415 B.n557 VSUBS 0.006997f
C1416 B.n558 VSUBS 0.006997f
C1417 B.n559 VSUBS 0.006997f
C1418 B.n560 VSUBS 0.006997f
C1419 B.n561 VSUBS 0.006997f
C1420 B.n562 VSUBS 0.006997f
C1421 B.n563 VSUBS 0.006997f
C1422 B.n564 VSUBS 0.006997f
C1423 B.n565 VSUBS 0.006997f
C1424 B.n566 VSUBS 0.006997f
C1425 B.n567 VSUBS 0.006997f
C1426 B.n568 VSUBS 0.006997f
C1427 B.n569 VSUBS 0.006997f
C1428 B.n570 VSUBS 0.006997f
C1429 B.n571 VSUBS 0.006997f
C1430 B.n572 VSUBS 0.006997f
C1431 B.n573 VSUBS 0.006997f
C1432 B.n574 VSUBS 0.006997f
C1433 B.n575 VSUBS 0.006997f
C1434 B.n576 VSUBS 0.006997f
C1435 B.n577 VSUBS 0.006997f
C1436 B.n578 VSUBS 0.006997f
C1437 B.n579 VSUBS 0.006997f
C1438 B.n580 VSUBS 0.006997f
C1439 B.n581 VSUBS 0.006997f
C1440 B.n582 VSUBS 0.006997f
C1441 B.n583 VSUBS 0.006997f
C1442 B.n584 VSUBS 0.006997f
C1443 B.n585 VSUBS 0.006997f
C1444 B.n586 VSUBS 0.006997f
C1445 B.n587 VSUBS 0.006997f
C1446 B.n588 VSUBS 0.006997f
C1447 B.n589 VSUBS 0.006997f
C1448 B.n590 VSUBS 0.006997f
C1449 B.n591 VSUBS 0.006997f
C1450 B.n592 VSUBS 0.006997f
C1451 B.n593 VSUBS 0.006997f
C1452 B.n594 VSUBS 0.006997f
C1453 B.n595 VSUBS 0.006997f
C1454 B.n596 VSUBS 0.006997f
C1455 B.n597 VSUBS 0.006997f
C1456 B.n598 VSUBS 0.006997f
C1457 B.n599 VSUBS 0.006997f
C1458 B.n600 VSUBS 0.006997f
C1459 B.n601 VSUBS 0.006997f
C1460 B.n602 VSUBS 0.006997f
C1461 B.n603 VSUBS 0.006997f
C1462 B.n604 VSUBS 0.006997f
C1463 B.n605 VSUBS 0.006997f
C1464 B.n606 VSUBS 0.006997f
C1465 B.n607 VSUBS 0.006997f
C1466 B.n608 VSUBS 0.006997f
C1467 B.n609 VSUBS 0.006997f
C1468 B.n610 VSUBS 0.006997f
C1469 B.n611 VSUBS 0.006997f
C1470 B.n612 VSUBS 0.006997f
C1471 B.n613 VSUBS 0.006997f
C1472 B.n614 VSUBS 0.006997f
C1473 B.n615 VSUBS 0.006997f
C1474 B.n616 VSUBS 0.006997f
C1475 B.n617 VSUBS 0.006997f
C1476 B.n618 VSUBS 0.006997f
C1477 B.n619 VSUBS 0.006997f
C1478 B.n620 VSUBS 0.01641f
C1479 B.n621 VSUBS 0.01641f
C1480 B.n622 VSUBS 0.016104f
C1481 B.n623 VSUBS 0.006997f
C1482 B.n624 VSUBS 0.006997f
C1483 B.n625 VSUBS 0.006997f
C1484 B.n626 VSUBS 0.006997f
C1485 B.n627 VSUBS 0.006997f
C1486 B.n628 VSUBS 0.006997f
C1487 B.n629 VSUBS 0.006997f
C1488 B.n630 VSUBS 0.006997f
C1489 B.n631 VSUBS 0.006997f
C1490 B.n632 VSUBS 0.006997f
C1491 B.n633 VSUBS 0.006997f
C1492 B.n634 VSUBS 0.006997f
C1493 B.n635 VSUBS 0.006997f
C1494 B.n636 VSUBS 0.006997f
C1495 B.n637 VSUBS 0.006997f
C1496 B.n638 VSUBS 0.006997f
C1497 B.n639 VSUBS 0.006997f
C1498 B.n640 VSUBS 0.006997f
C1499 B.n641 VSUBS 0.006997f
C1500 B.n642 VSUBS 0.006997f
C1501 B.n643 VSUBS 0.006997f
C1502 B.n644 VSUBS 0.006997f
C1503 B.n645 VSUBS 0.006997f
C1504 B.n646 VSUBS 0.006997f
C1505 B.n647 VSUBS 0.006997f
C1506 B.n648 VSUBS 0.006997f
C1507 B.n649 VSUBS 0.006997f
C1508 B.n650 VSUBS 0.006997f
C1509 B.n651 VSUBS 0.015843f
.ends

