* NGSPICE file created from diff_pair_sample_1799.ext - technology: sky130A

.subckt diff_pair_sample_1799 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t7 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=2.8545 pd=17.63 as=6.747 ps=35.38 w=17.3 l=2.88
X1 B.t11 B.t9 B.t10 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=6.747 pd=35.38 as=0 ps=0 w=17.3 l=2.88
X2 VTAIL.t4 VN.t1 VDD2.t2 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=6.747 pd=35.38 as=2.8545 ps=17.63 w=17.3 l=2.88
X3 VTAIL.t1 VP.t0 VDD1.t3 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=6.747 pd=35.38 as=2.8545 ps=17.63 w=17.3 l=2.88
X4 B.t8 B.t6 B.t7 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=6.747 pd=35.38 as=0 ps=0 w=17.3 l=2.88
X5 B.t5 B.t3 B.t4 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=6.747 pd=35.38 as=0 ps=0 w=17.3 l=2.88
X6 VDD2.t1 VN.t2 VTAIL.t6 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=2.8545 pd=17.63 as=6.747 ps=35.38 w=17.3 l=2.88
X7 VTAIL.t3 VP.t1 VDD1.t2 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=6.747 pd=35.38 as=2.8545 ps=17.63 w=17.3 l=2.88
X8 VDD1.t1 VP.t2 VTAIL.t2 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=2.8545 pd=17.63 as=6.747 ps=35.38 w=17.3 l=2.88
X9 VDD1.t0 VP.t3 VTAIL.t0 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=2.8545 pd=17.63 as=6.747 ps=35.38 w=17.3 l=2.88
X10 B.t2 B.t0 B.t1 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=6.747 pd=35.38 as=0 ps=0 w=17.3 l=2.88
X11 VTAIL.t5 VN.t3 VDD2.t0 w_n2896_n4428# sky130_fd_pr__pfet_01v8 ad=6.747 pd=35.38 as=2.8545 ps=17.63 w=17.3 l=2.88
R0 VN.n0 VN.t1 180.502
R1 VN.n1 VN.t2 180.502
R2 VN.n0 VN.t0 179.599
R3 VN.n1 VN.t3 179.599
R4 VN VN.n1 54.8787
R5 VN VN.n0 3.38246
R6 VTAIL.n5 VTAIL.t1 57.1174
R7 VTAIL.n4 VTAIL.t6 57.1174
R8 VTAIL.n3 VTAIL.t5 57.1174
R9 VTAIL.n7 VTAIL.t7 57.1173
R10 VTAIL.n0 VTAIL.t4 57.1173
R11 VTAIL.n1 VTAIL.t2 57.1173
R12 VTAIL.n2 VTAIL.t3 57.1173
R13 VTAIL.n6 VTAIL.t0 57.1173
R14 VTAIL.n7 VTAIL.n6 30.0479
R15 VTAIL.n3 VTAIL.n2 30.0479
R16 VTAIL.n4 VTAIL.n3 2.76774
R17 VTAIL.n6 VTAIL.n5 2.76774
R18 VTAIL.n2 VTAIL.n1 2.76774
R19 VTAIL VTAIL.n0 1.44231
R20 VTAIL VTAIL.n7 1.32593
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 118.847
R24 VDD2.n2 VDD2.n1 71.9171
R25 VDD2.n1 VDD2.t0 1.8794
R26 VDD2.n1 VDD2.t1 1.8794
R27 VDD2.n0 VDD2.t2 1.8794
R28 VDD2.n0 VDD2.t3 1.8794
R29 VDD2 VDD2.n2 0.0586897
R30 B.n447 B.n124 585
R31 B.n446 B.n445 585
R32 B.n444 B.n125 585
R33 B.n443 B.n442 585
R34 B.n441 B.n126 585
R35 B.n440 B.n439 585
R36 B.n438 B.n127 585
R37 B.n437 B.n436 585
R38 B.n435 B.n128 585
R39 B.n434 B.n433 585
R40 B.n432 B.n129 585
R41 B.n431 B.n430 585
R42 B.n429 B.n130 585
R43 B.n428 B.n427 585
R44 B.n426 B.n131 585
R45 B.n425 B.n424 585
R46 B.n423 B.n132 585
R47 B.n422 B.n421 585
R48 B.n420 B.n133 585
R49 B.n419 B.n418 585
R50 B.n417 B.n134 585
R51 B.n416 B.n415 585
R52 B.n414 B.n135 585
R53 B.n413 B.n412 585
R54 B.n411 B.n136 585
R55 B.n410 B.n409 585
R56 B.n408 B.n137 585
R57 B.n407 B.n406 585
R58 B.n405 B.n138 585
R59 B.n404 B.n403 585
R60 B.n402 B.n139 585
R61 B.n401 B.n400 585
R62 B.n399 B.n140 585
R63 B.n398 B.n397 585
R64 B.n396 B.n141 585
R65 B.n395 B.n394 585
R66 B.n393 B.n142 585
R67 B.n392 B.n391 585
R68 B.n390 B.n143 585
R69 B.n389 B.n388 585
R70 B.n387 B.n144 585
R71 B.n386 B.n385 585
R72 B.n384 B.n145 585
R73 B.n383 B.n382 585
R74 B.n381 B.n146 585
R75 B.n380 B.n379 585
R76 B.n378 B.n147 585
R77 B.n377 B.n376 585
R78 B.n375 B.n148 585
R79 B.n374 B.n373 585
R80 B.n372 B.n149 585
R81 B.n371 B.n370 585
R82 B.n369 B.n150 585
R83 B.n368 B.n367 585
R84 B.n366 B.n151 585
R85 B.n365 B.n364 585
R86 B.n363 B.n152 585
R87 B.n361 B.n360 585
R88 B.n359 B.n155 585
R89 B.n358 B.n357 585
R90 B.n356 B.n156 585
R91 B.n355 B.n354 585
R92 B.n353 B.n157 585
R93 B.n352 B.n351 585
R94 B.n350 B.n158 585
R95 B.n349 B.n348 585
R96 B.n347 B.n159 585
R97 B.n346 B.n345 585
R98 B.n341 B.n160 585
R99 B.n340 B.n339 585
R100 B.n338 B.n161 585
R101 B.n337 B.n336 585
R102 B.n335 B.n162 585
R103 B.n334 B.n333 585
R104 B.n332 B.n163 585
R105 B.n331 B.n330 585
R106 B.n329 B.n164 585
R107 B.n328 B.n327 585
R108 B.n326 B.n165 585
R109 B.n325 B.n324 585
R110 B.n323 B.n166 585
R111 B.n322 B.n321 585
R112 B.n320 B.n167 585
R113 B.n319 B.n318 585
R114 B.n317 B.n168 585
R115 B.n316 B.n315 585
R116 B.n314 B.n169 585
R117 B.n313 B.n312 585
R118 B.n311 B.n170 585
R119 B.n310 B.n309 585
R120 B.n308 B.n171 585
R121 B.n307 B.n306 585
R122 B.n305 B.n172 585
R123 B.n304 B.n303 585
R124 B.n302 B.n173 585
R125 B.n301 B.n300 585
R126 B.n299 B.n174 585
R127 B.n298 B.n297 585
R128 B.n296 B.n175 585
R129 B.n295 B.n294 585
R130 B.n293 B.n176 585
R131 B.n292 B.n291 585
R132 B.n290 B.n177 585
R133 B.n289 B.n288 585
R134 B.n287 B.n178 585
R135 B.n286 B.n285 585
R136 B.n284 B.n179 585
R137 B.n283 B.n282 585
R138 B.n281 B.n180 585
R139 B.n280 B.n279 585
R140 B.n278 B.n181 585
R141 B.n277 B.n276 585
R142 B.n275 B.n182 585
R143 B.n274 B.n273 585
R144 B.n272 B.n183 585
R145 B.n271 B.n270 585
R146 B.n269 B.n184 585
R147 B.n268 B.n267 585
R148 B.n266 B.n185 585
R149 B.n265 B.n264 585
R150 B.n263 B.n186 585
R151 B.n262 B.n261 585
R152 B.n260 B.n187 585
R153 B.n259 B.n258 585
R154 B.n449 B.n448 585
R155 B.n450 B.n123 585
R156 B.n452 B.n451 585
R157 B.n453 B.n122 585
R158 B.n455 B.n454 585
R159 B.n456 B.n121 585
R160 B.n458 B.n457 585
R161 B.n459 B.n120 585
R162 B.n461 B.n460 585
R163 B.n462 B.n119 585
R164 B.n464 B.n463 585
R165 B.n465 B.n118 585
R166 B.n467 B.n466 585
R167 B.n468 B.n117 585
R168 B.n470 B.n469 585
R169 B.n471 B.n116 585
R170 B.n473 B.n472 585
R171 B.n474 B.n115 585
R172 B.n476 B.n475 585
R173 B.n477 B.n114 585
R174 B.n479 B.n478 585
R175 B.n480 B.n113 585
R176 B.n482 B.n481 585
R177 B.n483 B.n112 585
R178 B.n485 B.n484 585
R179 B.n486 B.n111 585
R180 B.n488 B.n487 585
R181 B.n489 B.n110 585
R182 B.n491 B.n490 585
R183 B.n492 B.n109 585
R184 B.n494 B.n493 585
R185 B.n495 B.n108 585
R186 B.n497 B.n496 585
R187 B.n498 B.n107 585
R188 B.n500 B.n499 585
R189 B.n501 B.n106 585
R190 B.n503 B.n502 585
R191 B.n504 B.n105 585
R192 B.n506 B.n505 585
R193 B.n507 B.n104 585
R194 B.n509 B.n508 585
R195 B.n510 B.n103 585
R196 B.n512 B.n511 585
R197 B.n513 B.n102 585
R198 B.n515 B.n514 585
R199 B.n516 B.n101 585
R200 B.n518 B.n517 585
R201 B.n519 B.n100 585
R202 B.n521 B.n520 585
R203 B.n522 B.n99 585
R204 B.n524 B.n523 585
R205 B.n525 B.n98 585
R206 B.n527 B.n526 585
R207 B.n528 B.n97 585
R208 B.n530 B.n529 585
R209 B.n531 B.n96 585
R210 B.n533 B.n532 585
R211 B.n534 B.n95 585
R212 B.n536 B.n535 585
R213 B.n537 B.n94 585
R214 B.n539 B.n538 585
R215 B.n540 B.n93 585
R216 B.n542 B.n541 585
R217 B.n543 B.n92 585
R218 B.n545 B.n544 585
R219 B.n546 B.n91 585
R220 B.n548 B.n547 585
R221 B.n549 B.n90 585
R222 B.n551 B.n550 585
R223 B.n552 B.n89 585
R224 B.n554 B.n553 585
R225 B.n555 B.n88 585
R226 B.n557 B.n556 585
R227 B.n558 B.n87 585
R228 B.n745 B.n20 585
R229 B.n744 B.n743 585
R230 B.n742 B.n21 585
R231 B.n741 B.n740 585
R232 B.n739 B.n22 585
R233 B.n738 B.n737 585
R234 B.n736 B.n23 585
R235 B.n735 B.n734 585
R236 B.n733 B.n24 585
R237 B.n732 B.n731 585
R238 B.n730 B.n25 585
R239 B.n729 B.n728 585
R240 B.n727 B.n26 585
R241 B.n726 B.n725 585
R242 B.n724 B.n27 585
R243 B.n723 B.n722 585
R244 B.n721 B.n28 585
R245 B.n720 B.n719 585
R246 B.n718 B.n29 585
R247 B.n717 B.n716 585
R248 B.n715 B.n30 585
R249 B.n714 B.n713 585
R250 B.n712 B.n31 585
R251 B.n711 B.n710 585
R252 B.n709 B.n32 585
R253 B.n708 B.n707 585
R254 B.n706 B.n33 585
R255 B.n705 B.n704 585
R256 B.n703 B.n34 585
R257 B.n702 B.n701 585
R258 B.n700 B.n35 585
R259 B.n699 B.n698 585
R260 B.n697 B.n36 585
R261 B.n696 B.n695 585
R262 B.n694 B.n37 585
R263 B.n693 B.n692 585
R264 B.n691 B.n38 585
R265 B.n690 B.n689 585
R266 B.n688 B.n39 585
R267 B.n687 B.n686 585
R268 B.n685 B.n40 585
R269 B.n684 B.n683 585
R270 B.n682 B.n41 585
R271 B.n681 B.n680 585
R272 B.n679 B.n42 585
R273 B.n678 B.n677 585
R274 B.n676 B.n43 585
R275 B.n675 B.n674 585
R276 B.n673 B.n44 585
R277 B.n672 B.n671 585
R278 B.n670 B.n45 585
R279 B.n669 B.n668 585
R280 B.n667 B.n46 585
R281 B.n666 B.n665 585
R282 B.n664 B.n47 585
R283 B.n663 B.n662 585
R284 B.n661 B.n48 585
R285 B.n660 B.n659 585
R286 B.n658 B.n49 585
R287 B.n657 B.n656 585
R288 B.n655 B.n53 585
R289 B.n654 B.n653 585
R290 B.n652 B.n54 585
R291 B.n651 B.n650 585
R292 B.n649 B.n55 585
R293 B.n648 B.n647 585
R294 B.n646 B.n56 585
R295 B.n644 B.n643 585
R296 B.n642 B.n59 585
R297 B.n641 B.n640 585
R298 B.n639 B.n60 585
R299 B.n638 B.n637 585
R300 B.n636 B.n61 585
R301 B.n635 B.n634 585
R302 B.n633 B.n62 585
R303 B.n632 B.n631 585
R304 B.n630 B.n63 585
R305 B.n629 B.n628 585
R306 B.n627 B.n64 585
R307 B.n626 B.n625 585
R308 B.n624 B.n65 585
R309 B.n623 B.n622 585
R310 B.n621 B.n66 585
R311 B.n620 B.n619 585
R312 B.n618 B.n67 585
R313 B.n617 B.n616 585
R314 B.n615 B.n68 585
R315 B.n614 B.n613 585
R316 B.n612 B.n69 585
R317 B.n611 B.n610 585
R318 B.n609 B.n70 585
R319 B.n608 B.n607 585
R320 B.n606 B.n71 585
R321 B.n605 B.n604 585
R322 B.n603 B.n72 585
R323 B.n602 B.n601 585
R324 B.n600 B.n73 585
R325 B.n599 B.n598 585
R326 B.n597 B.n74 585
R327 B.n596 B.n595 585
R328 B.n594 B.n75 585
R329 B.n593 B.n592 585
R330 B.n591 B.n76 585
R331 B.n590 B.n589 585
R332 B.n588 B.n77 585
R333 B.n587 B.n586 585
R334 B.n585 B.n78 585
R335 B.n584 B.n583 585
R336 B.n582 B.n79 585
R337 B.n581 B.n580 585
R338 B.n579 B.n80 585
R339 B.n578 B.n577 585
R340 B.n576 B.n81 585
R341 B.n575 B.n574 585
R342 B.n573 B.n82 585
R343 B.n572 B.n571 585
R344 B.n570 B.n83 585
R345 B.n569 B.n568 585
R346 B.n567 B.n84 585
R347 B.n566 B.n565 585
R348 B.n564 B.n85 585
R349 B.n563 B.n562 585
R350 B.n561 B.n86 585
R351 B.n560 B.n559 585
R352 B.n747 B.n746 585
R353 B.n748 B.n19 585
R354 B.n750 B.n749 585
R355 B.n751 B.n18 585
R356 B.n753 B.n752 585
R357 B.n754 B.n17 585
R358 B.n756 B.n755 585
R359 B.n757 B.n16 585
R360 B.n759 B.n758 585
R361 B.n760 B.n15 585
R362 B.n762 B.n761 585
R363 B.n763 B.n14 585
R364 B.n765 B.n764 585
R365 B.n766 B.n13 585
R366 B.n768 B.n767 585
R367 B.n769 B.n12 585
R368 B.n771 B.n770 585
R369 B.n772 B.n11 585
R370 B.n774 B.n773 585
R371 B.n775 B.n10 585
R372 B.n777 B.n776 585
R373 B.n778 B.n9 585
R374 B.n780 B.n779 585
R375 B.n781 B.n8 585
R376 B.n783 B.n782 585
R377 B.n784 B.n7 585
R378 B.n786 B.n785 585
R379 B.n787 B.n6 585
R380 B.n789 B.n788 585
R381 B.n790 B.n5 585
R382 B.n792 B.n791 585
R383 B.n793 B.n4 585
R384 B.n795 B.n794 585
R385 B.n796 B.n3 585
R386 B.n798 B.n797 585
R387 B.n799 B.n0 585
R388 B.n2 B.n1 585
R389 B.n206 B.n205 585
R390 B.n208 B.n207 585
R391 B.n209 B.n204 585
R392 B.n211 B.n210 585
R393 B.n212 B.n203 585
R394 B.n214 B.n213 585
R395 B.n215 B.n202 585
R396 B.n217 B.n216 585
R397 B.n218 B.n201 585
R398 B.n220 B.n219 585
R399 B.n221 B.n200 585
R400 B.n223 B.n222 585
R401 B.n224 B.n199 585
R402 B.n226 B.n225 585
R403 B.n227 B.n198 585
R404 B.n229 B.n228 585
R405 B.n230 B.n197 585
R406 B.n232 B.n231 585
R407 B.n233 B.n196 585
R408 B.n235 B.n234 585
R409 B.n236 B.n195 585
R410 B.n238 B.n237 585
R411 B.n239 B.n194 585
R412 B.n241 B.n240 585
R413 B.n242 B.n193 585
R414 B.n244 B.n243 585
R415 B.n245 B.n192 585
R416 B.n247 B.n246 585
R417 B.n248 B.n191 585
R418 B.n250 B.n249 585
R419 B.n251 B.n190 585
R420 B.n253 B.n252 585
R421 B.n254 B.n189 585
R422 B.n256 B.n255 585
R423 B.n257 B.n188 585
R424 B.n259 B.n188 487.695
R425 B.n449 B.n124 487.695
R426 B.n559 B.n558 487.695
R427 B.n746 B.n745 487.695
R428 B.n342 B.t0 353.202
R429 B.n153 B.t9 353.202
R430 B.n57 B.t3 353.202
R431 B.n50 B.t6 353.202
R432 B.n801 B.n800 256.663
R433 B.n800 B.n799 235.042
R434 B.n800 B.n2 235.042
R435 B.n153 B.t10 174.349
R436 B.n57 B.t5 174.349
R437 B.n342 B.t1 174.327
R438 B.n50 B.t8 174.327
R439 B.n260 B.n259 163.367
R440 B.n261 B.n260 163.367
R441 B.n261 B.n186 163.367
R442 B.n265 B.n186 163.367
R443 B.n266 B.n265 163.367
R444 B.n267 B.n266 163.367
R445 B.n267 B.n184 163.367
R446 B.n271 B.n184 163.367
R447 B.n272 B.n271 163.367
R448 B.n273 B.n272 163.367
R449 B.n273 B.n182 163.367
R450 B.n277 B.n182 163.367
R451 B.n278 B.n277 163.367
R452 B.n279 B.n278 163.367
R453 B.n279 B.n180 163.367
R454 B.n283 B.n180 163.367
R455 B.n284 B.n283 163.367
R456 B.n285 B.n284 163.367
R457 B.n285 B.n178 163.367
R458 B.n289 B.n178 163.367
R459 B.n290 B.n289 163.367
R460 B.n291 B.n290 163.367
R461 B.n291 B.n176 163.367
R462 B.n295 B.n176 163.367
R463 B.n296 B.n295 163.367
R464 B.n297 B.n296 163.367
R465 B.n297 B.n174 163.367
R466 B.n301 B.n174 163.367
R467 B.n302 B.n301 163.367
R468 B.n303 B.n302 163.367
R469 B.n303 B.n172 163.367
R470 B.n307 B.n172 163.367
R471 B.n308 B.n307 163.367
R472 B.n309 B.n308 163.367
R473 B.n309 B.n170 163.367
R474 B.n313 B.n170 163.367
R475 B.n314 B.n313 163.367
R476 B.n315 B.n314 163.367
R477 B.n315 B.n168 163.367
R478 B.n319 B.n168 163.367
R479 B.n320 B.n319 163.367
R480 B.n321 B.n320 163.367
R481 B.n321 B.n166 163.367
R482 B.n325 B.n166 163.367
R483 B.n326 B.n325 163.367
R484 B.n327 B.n326 163.367
R485 B.n327 B.n164 163.367
R486 B.n331 B.n164 163.367
R487 B.n332 B.n331 163.367
R488 B.n333 B.n332 163.367
R489 B.n333 B.n162 163.367
R490 B.n337 B.n162 163.367
R491 B.n338 B.n337 163.367
R492 B.n339 B.n338 163.367
R493 B.n339 B.n160 163.367
R494 B.n346 B.n160 163.367
R495 B.n347 B.n346 163.367
R496 B.n348 B.n347 163.367
R497 B.n348 B.n158 163.367
R498 B.n352 B.n158 163.367
R499 B.n353 B.n352 163.367
R500 B.n354 B.n353 163.367
R501 B.n354 B.n156 163.367
R502 B.n358 B.n156 163.367
R503 B.n359 B.n358 163.367
R504 B.n360 B.n359 163.367
R505 B.n360 B.n152 163.367
R506 B.n365 B.n152 163.367
R507 B.n366 B.n365 163.367
R508 B.n367 B.n366 163.367
R509 B.n367 B.n150 163.367
R510 B.n371 B.n150 163.367
R511 B.n372 B.n371 163.367
R512 B.n373 B.n372 163.367
R513 B.n373 B.n148 163.367
R514 B.n377 B.n148 163.367
R515 B.n378 B.n377 163.367
R516 B.n379 B.n378 163.367
R517 B.n379 B.n146 163.367
R518 B.n383 B.n146 163.367
R519 B.n384 B.n383 163.367
R520 B.n385 B.n384 163.367
R521 B.n385 B.n144 163.367
R522 B.n389 B.n144 163.367
R523 B.n390 B.n389 163.367
R524 B.n391 B.n390 163.367
R525 B.n391 B.n142 163.367
R526 B.n395 B.n142 163.367
R527 B.n396 B.n395 163.367
R528 B.n397 B.n396 163.367
R529 B.n397 B.n140 163.367
R530 B.n401 B.n140 163.367
R531 B.n402 B.n401 163.367
R532 B.n403 B.n402 163.367
R533 B.n403 B.n138 163.367
R534 B.n407 B.n138 163.367
R535 B.n408 B.n407 163.367
R536 B.n409 B.n408 163.367
R537 B.n409 B.n136 163.367
R538 B.n413 B.n136 163.367
R539 B.n414 B.n413 163.367
R540 B.n415 B.n414 163.367
R541 B.n415 B.n134 163.367
R542 B.n419 B.n134 163.367
R543 B.n420 B.n419 163.367
R544 B.n421 B.n420 163.367
R545 B.n421 B.n132 163.367
R546 B.n425 B.n132 163.367
R547 B.n426 B.n425 163.367
R548 B.n427 B.n426 163.367
R549 B.n427 B.n130 163.367
R550 B.n431 B.n130 163.367
R551 B.n432 B.n431 163.367
R552 B.n433 B.n432 163.367
R553 B.n433 B.n128 163.367
R554 B.n437 B.n128 163.367
R555 B.n438 B.n437 163.367
R556 B.n439 B.n438 163.367
R557 B.n439 B.n126 163.367
R558 B.n443 B.n126 163.367
R559 B.n444 B.n443 163.367
R560 B.n445 B.n444 163.367
R561 B.n445 B.n124 163.367
R562 B.n558 B.n557 163.367
R563 B.n557 B.n88 163.367
R564 B.n553 B.n88 163.367
R565 B.n553 B.n552 163.367
R566 B.n552 B.n551 163.367
R567 B.n551 B.n90 163.367
R568 B.n547 B.n90 163.367
R569 B.n547 B.n546 163.367
R570 B.n546 B.n545 163.367
R571 B.n545 B.n92 163.367
R572 B.n541 B.n92 163.367
R573 B.n541 B.n540 163.367
R574 B.n540 B.n539 163.367
R575 B.n539 B.n94 163.367
R576 B.n535 B.n94 163.367
R577 B.n535 B.n534 163.367
R578 B.n534 B.n533 163.367
R579 B.n533 B.n96 163.367
R580 B.n529 B.n96 163.367
R581 B.n529 B.n528 163.367
R582 B.n528 B.n527 163.367
R583 B.n527 B.n98 163.367
R584 B.n523 B.n98 163.367
R585 B.n523 B.n522 163.367
R586 B.n522 B.n521 163.367
R587 B.n521 B.n100 163.367
R588 B.n517 B.n100 163.367
R589 B.n517 B.n516 163.367
R590 B.n516 B.n515 163.367
R591 B.n515 B.n102 163.367
R592 B.n511 B.n102 163.367
R593 B.n511 B.n510 163.367
R594 B.n510 B.n509 163.367
R595 B.n509 B.n104 163.367
R596 B.n505 B.n104 163.367
R597 B.n505 B.n504 163.367
R598 B.n504 B.n503 163.367
R599 B.n503 B.n106 163.367
R600 B.n499 B.n106 163.367
R601 B.n499 B.n498 163.367
R602 B.n498 B.n497 163.367
R603 B.n497 B.n108 163.367
R604 B.n493 B.n108 163.367
R605 B.n493 B.n492 163.367
R606 B.n492 B.n491 163.367
R607 B.n491 B.n110 163.367
R608 B.n487 B.n110 163.367
R609 B.n487 B.n486 163.367
R610 B.n486 B.n485 163.367
R611 B.n485 B.n112 163.367
R612 B.n481 B.n112 163.367
R613 B.n481 B.n480 163.367
R614 B.n480 B.n479 163.367
R615 B.n479 B.n114 163.367
R616 B.n475 B.n114 163.367
R617 B.n475 B.n474 163.367
R618 B.n474 B.n473 163.367
R619 B.n473 B.n116 163.367
R620 B.n469 B.n116 163.367
R621 B.n469 B.n468 163.367
R622 B.n468 B.n467 163.367
R623 B.n467 B.n118 163.367
R624 B.n463 B.n118 163.367
R625 B.n463 B.n462 163.367
R626 B.n462 B.n461 163.367
R627 B.n461 B.n120 163.367
R628 B.n457 B.n120 163.367
R629 B.n457 B.n456 163.367
R630 B.n456 B.n455 163.367
R631 B.n455 B.n122 163.367
R632 B.n451 B.n122 163.367
R633 B.n451 B.n450 163.367
R634 B.n450 B.n449 163.367
R635 B.n745 B.n744 163.367
R636 B.n744 B.n21 163.367
R637 B.n740 B.n21 163.367
R638 B.n740 B.n739 163.367
R639 B.n739 B.n738 163.367
R640 B.n738 B.n23 163.367
R641 B.n734 B.n23 163.367
R642 B.n734 B.n733 163.367
R643 B.n733 B.n732 163.367
R644 B.n732 B.n25 163.367
R645 B.n728 B.n25 163.367
R646 B.n728 B.n727 163.367
R647 B.n727 B.n726 163.367
R648 B.n726 B.n27 163.367
R649 B.n722 B.n27 163.367
R650 B.n722 B.n721 163.367
R651 B.n721 B.n720 163.367
R652 B.n720 B.n29 163.367
R653 B.n716 B.n29 163.367
R654 B.n716 B.n715 163.367
R655 B.n715 B.n714 163.367
R656 B.n714 B.n31 163.367
R657 B.n710 B.n31 163.367
R658 B.n710 B.n709 163.367
R659 B.n709 B.n708 163.367
R660 B.n708 B.n33 163.367
R661 B.n704 B.n33 163.367
R662 B.n704 B.n703 163.367
R663 B.n703 B.n702 163.367
R664 B.n702 B.n35 163.367
R665 B.n698 B.n35 163.367
R666 B.n698 B.n697 163.367
R667 B.n697 B.n696 163.367
R668 B.n696 B.n37 163.367
R669 B.n692 B.n37 163.367
R670 B.n692 B.n691 163.367
R671 B.n691 B.n690 163.367
R672 B.n690 B.n39 163.367
R673 B.n686 B.n39 163.367
R674 B.n686 B.n685 163.367
R675 B.n685 B.n684 163.367
R676 B.n684 B.n41 163.367
R677 B.n680 B.n41 163.367
R678 B.n680 B.n679 163.367
R679 B.n679 B.n678 163.367
R680 B.n678 B.n43 163.367
R681 B.n674 B.n43 163.367
R682 B.n674 B.n673 163.367
R683 B.n673 B.n672 163.367
R684 B.n672 B.n45 163.367
R685 B.n668 B.n45 163.367
R686 B.n668 B.n667 163.367
R687 B.n667 B.n666 163.367
R688 B.n666 B.n47 163.367
R689 B.n662 B.n47 163.367
R690 B.n662 B.n661 163.367
R691 B.n661 B.n660 163.367
R692 B.n660 B.n49 163.367
R693 B.n656 B.n49 163.367
R694 B.n656 B.n655 163.367
R695 B.n655 B.n654 163.367
R696 B.n654 B.n54 163.367
R697 B.n650 B.n54 163.367
R698 B.n650 B.n649 163.367
R699 B.n649 B.n648 163.367
R700 B.n648 B.n56 163.367
R701 B.n643 B.n56 163.367
R702 B.n643 B.n642 163.367
R703 B.n642 B.n641 163.367
R704 B.n641 B.n60 163.367
R705 B.n637 B.n60 163.367
R706 B.n637 B.n636 163.367
R707 B.n636 B.n635 163.367
R708 B.n635 B.n62 163.367
R709 B.n631 B.n62 163.367
R710 B.n631 B.n630 163.367
R711 B.n630 B.n629 163.367
R712 B.n629 B.n64 163.367
R713 B.n625 B.n64 163.367
R714 B.n625 B.n624 163.367
R715 B.n624 B.n623 163.367
R716 B.n623 B.n66 163.367
R717 B.n619 B.n66 163.367
R718 B.n619 B.n618 163.367
R719 B.n618 B.n617 163.367
R720 B.n617 B.n68 163.367
R721 B.n613 B.n68 163.367
R722 B.n613 B.n612 163.367
R723 B.n612 B.n611 163.367
R724 B.n611 B.n70 163.367
R725 B.n607 B.n70 163.367
R726 B.n607 B.n606 163.367
R727 B.n606 B.n605 163.367
R728 B.n605 B.n72 163.367
R729 B.n601 B.n72 163.367
R730 B.n601 B.n600 163.367
R731 B.n600 B.n599 163.367
R732 B.n599 B.n74 163.367
R733 B.n595 B.n74 163.367
R734 B.n595 B.n594 163.367
R735 B.n594 B.n593 163.367
R736 B.n593 B.n76 163.367
R737 B.n589 B.n76 163.367
R738 B.n589 B.n588 163.367
R739 B.n588 B.n587 163.367
R740 B.n587 B.n78 163.367
R741 B.n583 B.n78 163.367
R742 B.n583 B.n582 163.367
R743 B.n582 B.n581 163.367
R744 B.n581 B.n80 163.367
R745 B.n577 B.n80 163.367
R746 B.n577 B.n576 163.367
R747 B.n576 B.n575 163.367
R748 B.n575 B.n82 163.367
R749 B.n571 B.n82 163.367
R750 B.n571 B.n570 163.367
R751 B.n570 B.n569 163.367
R752 B.n569 B.n84 163.367
R753 B.n565 B.n84 163.367
R754 B.n565 B.n564 163.367
R755 B.n564 B.n563 163.367
R756 B.n563 B.n86 163.367
R757 B.n559 B.n86 163.367
R758 B.n746 B.n19 163.367
R759 B.n750 B.n19 163.367
R760 B.n751 B.n750 163.367
R761 B.n752 B.n751 163.367
R762 B.n752 B.n17 163.367
R763 B.n756 B.n17 163.367
R764 B.n757 B.n756 163.367
R765 B.n758 B.n757 163.367
R766 B.n758 B.n15 163.367
R767 B.n762 B.n15 163.367
R768 B.n763 B.n762 163.367
R769 B.n764 B.n763 163.367
R770 B.n764 B.n13 163.367
R771 B.n768 B.n13 163.367
R772 B.n769 B.n768 163.367
R773 B.n770 B.n769 163.367
R774 B.n770 B.n11 163.367
R775 B.n774 B.n11 163.367
R776 B.n775 B.n774 163.367
R777 B.n776 B.n775 163.367
R778 B.n776 B.n9 163.367
R779 B.n780 B.n9 163.367
R780 B.n781 B.n780 163.367
R781 B.n782 B.n781 163.367
R782 B.n782 B.n7 163.367
R783 B.n786 B.n7 163.367
R784 B.n787 B.n786 163.367
R785 B.n788 B.n787 163.367
R786 B.n788 B.n5 163.367
R787 B.n792 B.n5 163.367
R788 B.n793 B.n792 163.367
R789 B.n794 B.n793 163.367
R790 B.n794 B.n3 163.367
R791 B.n798 B.n3 163.367
R792 B.n799 B.n798 163.367
R793 B.n206 B.n2 163.367
R794 B.n207 B.n206 163.367
R795 B.n207 B.n204 163.367
R796 B.n211 B.n204 163.367
R797 B.n212 B.n211 163.367
R798 B.n213 B.n212 163.367
R799 B.n213 B.n202 163.367
R800 B.n217 B.n202 163.367
R801 B.n218 B.n217 163.367
R802 B.n219 B.n218 163.367
R803 B.n219 B.n200 163.367
R804 B.n223 B.n200 163.367
R805 B.n224 B.n223 163.367
R806 B.n225 B.n224 163.367
R807 B.n225 B.n198 163.367
R808 B.n229 B.n198 163.367
R809 B.n230 B.n229 163.367
R810 B.n231 B.n230 163.367
R811 B.n231 B.n196 163.367
R812 B.n235 B.n196 163.367
R813 B.n236 B.n235 163.367
R814 B.n237 B.n236 163.367
R815 B.n237 B.n194 163.367
R816 B.n241 B.n194 163.367
R817 B.n242 B.n241 163.367
R818 B.n243 B.n242 163.367
R819 B.n243 B.n192 163.367
R820 B.n247 B.n192 163.367
R821 B.n248 B.n247 163.367
R822 B.n249 B.n248 163.367
R823 B.n249 B.n190 163.367
R824 B.n253 B.n190 163.367
R825 B.n254 B.n253 163.367
R826 B.n255 B.n254 163.367
R827 B.n255 B.n188 163.367
R828 B.n154 B.t11 112.094
R829 B.n58 B.t4 112.094
R830 B.n343 B.t2 112.073
R831 B.n51 B.t7 112.073
R832 B.n343 B.n342 62.255
R833 B.n154 B.n153 62.255
R834 B.n58 B.n57 62.255
R835 B.n51 B.n50 62.255
R836 B.n344 B.n343 59.5399
R837 B.n362 B.n154 59.5399
R838 B.n645 B.n58 59.5399
R839 B.n52 B.n51 59.5399
R840 B.n747 B.n20 31.6883
R841 B.n560 B.n87 31.6883
R842 B.n448 B.n447 31.6883
R843 B.n258 B.n257 31.6883
R844 B B.n801 18.0485
R845 B.n748 B.n747 10.6151
R846 B.n749 B.n748 10.6151
R847 B.n749 B.n18 10.6151
R848 B.n753 B.n18 10.6151
R849 B.n754 B.n753 10.6151
R850 B.n755 B.n754 10.6151
R851 B.n755 B.n16 10.6151
R852 B.n759 B.n16 10.6151
R853 B.n760 B.n759 10.6151
R854 B.n761 B.n760 10.6151
R855 B.n761 B.n14 10.6151
R856 B.n765 B.n14 10.6151
R857 B.n766 B.n765 10.6151
R858 B.n767 B.n766 10.6151
R859 B.n767 B.n12 10.6151
R860 B.n771 B.n12 10.6151
R861 B.n772 B.n771 10.6151
R862 B.n773 B.n772 10.6151
R863 B.n773 B.n10 10.6151
R864 B.n777 B.n10 10.6151
R865 B.n778 B.n777 10.6151
R866 B.n779 B.n778 10.6151
R867 B.n779 B.n8 10.6151
R868 B.n783 B.n8 10.6151
R869 B.n784 B.n783 10.6151
R870 B.n785 B.n784 10.6151
R871 B.n785 B.n6 10.6151
R872 B.n789 B.n6 10.6151
R873 B.n790 B.n789 10.6151
R874 B.n791 B.n790 10.6151
R875 B.n791 B.n4 10.6151
R876 B.n795 B.n4 10.6151
R877 B.n796 B.n795 10.6151
R878 B.n797 B.n796 10.6151
R879 B.n797 B.n0 10.6151
R880 B.n743 B.n20 10.6151
R881 B.n743 B.n742 10.6151
R882 B.n742 B.n741 10.6151
R883 B.n741 B.n22 10.6151
R884 B.n737 B.n22 10.6151
R885 B.n737 B.n736 10.6151
R886 B.n736 B.n735 10.6151
R887 B.n735 B.n24 10.6151
R888 B.n731 B.n24 10.6151
R889 B.n731 B.n730 10.6151
R890 B.n730 B.n729 10.6151
R891 B.n729 B.n26 10.6151
R892 B.n725 B.n26 10.6151
R893 B.n725 B.n724 10.6151
R894 B.n724 B.n723 10.6151
R895 B.n723 B.n28 10.6151
R896 B.n719 B.n28 10.6151
R897 B.n719 B.n718 10.6151
R898 B.n718 B.n717 10.6151
R899 B.n717 B.n30 10.6151
R900 B.n713 B.n30 10.6151
R901 B.n713 B.n712 10.6151
R902 B.n712 B.n711 10.6151
R903 B.n711 B.n32 10.6151
R904 B.n707 B.n32 10.6151
R905 B.n707 B.n706 10.6151
R906 B.n706 B.n705 10.6151
R907 B.n705 B.n34 10.6151
R908 B.n701 B.n34 10.6151
R909 B.n701 B.n700 10.6151
R910 B.n700 B.n699 10.6151
R911 B.n699 B.n36 10.6151
R912 B.n695 B.n36 10.6151
R913 B.n695 B.n694 10.6151
R914 B.n694 B.n693 10.6151
R915 B.n693 B.n38 10.6151
R916 B.n689 B.n38 10.6151
R917 B.n689 B.n688 10.6151
R918 B.n688 B.n687 10.6151
R919 B.n687 B.n40 10.6151
R920 B.n683 B.n40 10.6151
R921 B.n683 B.n682 10.6151
R922 B.n682 B.n681 10.6151
R923 B.n681 B.n42 10.6151
R924 B.n677 B.n42 10.6151
R925 B.n677 B.n676 10.6151
R926 B.n676 B.n675 10.6151
R927 B.n675 B.n44 10.6151
R928 B.n671 B.n44 10.6151
R929 B.n671 B.n670 10.6151
R930 B.n670 B.n669 10.6151
R931 B.n669 B.n46 10.6151
R932 B.n665 B.n46 10.6151
R933 B.n665 B.n664 10.6151
R934 B.n664 B.n663 10.6151
R935 B.n663 B.n48 10.6151
R936 B.n659 B.n658 10.6151
R937 B.n658 B.n657 10.6151
R938 B.n657 B.n53 10.6151
R939 B.n653 B.n53 10.6151
R940 B.n653 B.n652 10.6151
R941 B.n652 B.n651 10.6151
R942 B.n651 B.n55 10.6151
R943 B.n647 B.n55 10.6151
R944 B.n647 B.n646 10.6151
R945 B.n644 B.n59 10.6151
R946 B.n640 B.n59 10.6151
R947 B.n640 B.n639 10.6151
R948 B.n639 B.n638 10.6151
R949 B.n638 B.n61 10.6151
R950 B.n634 B.n61 10.6151
R951 B.n634 B.n633 10.6151
R952 B.n633 B.n632 10.6151
R953 B.n632 B.n63 10.6151
R954 B.n628 B.n63 10.6151
R955 B.n628 B.n627 10.6151
R956 B.n627 B.n626 10.6151
R957 B.n626 B.n65 10.6151
R958 B.n622 B.n65 10.6151
R959 B.n622 B.n621 10.6151
R960 B.n621 B.n620 10.6151
R961 B.n620 B.n67 10.6151
R962 B.n616 B.n67 10.6151
R963 B.n616 B.n615 10.6151
R964 B.n615 B.n614 10.6151
R965 B.n614 B.n69 10.6151
R966 B.n610 B.n69 10.6151
R967 B.n610 B.n609 10.6151
R968 B.n609 B.n608 10.6151
R969 B.n608 B.n71 10.6151
R970 B.n604 B.n71 10.6151
R971 B.n604 B.n603 10.6151
R972 B.n603 B.n602 10.6151
R973 B.n602 B.n73 10.6151
R974 B.n598 B.n73 10.6151
R975 B.n598 B.n597 10.6151
R976 B.n597 B.n596 10.6151
R977 B.n596 B.n75 10.6151
R978 B.n592 B.n75 10.6151
R979 B.n592 B.n591 10.6151
R980 B.n591 B.n590 10.6151
R981 B.n590 B.n77 10.6151
R982 B.n586 B.n77 10.6151
R983 B.n586 B.n585 10.6151
R984 B.n585 B.n584 10.6151
R985 B.n584 B.n79 10.6151
R986 B.n580 B.n79 10.6151
R987 B.n580 B.n579 10.6151
R988 B.n579 B.n578 10.6151
R989 B.n578 B.n81 10.6151
R990 B.n574 B.n81 10.6151
R991 B.n574 B.n573 10.6151
R992 B.n573 B.n572 10.6151
R993 B.n572 B.n83 10.6151
R994 B.n568 B.n83 10.6151
R995 B.n568 B.n567 10.6151
R996 B.n567 B.n566 10.6151
R997 B.n566 B.n85 10.6151
R998 B.n562 B.n85 10.6151
R999 B.n562 B.n561 10.6151
R1000 B.n561 B.n560 10.6151
R1001 B.n556 B.n87 10.6151
R1002 B.n556 B.n555 10.6151
R1003 B.n555 B.n554 10.6151
R1004 B.n554 B.n89 10.6151
R1005 B.n550 B.n89 10.6151
R1006 B.n550 B.n549 10.6151
R1007 B.n549 B.n548 10.6151
R1008 B.n548 B.n91 10.6151
R1009 B.n544 B.n91 10.6151
R1010 B.n544 B.n543 10.6151
R1011 B.n543 B.n542 10.6151
R1012 B.n542 B.n93 10.6151
R1013 B.n538 B.n93 10.6151
R1014 B.n538 B.n537 10.6151
R1015 B.n537 B.n536 10.6151
R1016 B.n536 B.n95 10.6151
R1017 B.n532 B.n95 10.6151
R1018 B.n532 B.n531 10.6151
R1019 B.n531 B.n530 10.6151
R1020 B.n530 B.n97 10.6151
R1021 B.n526 B.n97 10.6151
R1022 B.n526 B.n525 10.6151
R1023 B.n525 B.n524 10.6151
R1024 B.n524 B.n99 10.6151
R1025 B.n520 B.n99 10.6151
R1026 B.n520 B.n519 10.6151
R1027 B.n519 B.n518 10.6151
R1028 B.n518 B.n101 10.6151
R1029 B.n514 B.n101 10.6151
R1030 B.n514 B.n513 10.6151
R1031 B.n513 B.n512 10.6151
R1032 B.n512 B.n103 10.6151
R1033 B.n508 B.n103 10.6151
R1034 B.n508 B.n507 10.6151
R1035 B.n507 B.n506 10.6151
R1036 B.n506 B.n105 10.6151
R1037 B.n502 B.n105 10.6151
R1038 B.n502 B.n501 10.6151
R1039 B.n501 B.n500 10.6151
R1040 B.n500 B.n107 10.6151
R1041 B.n496 B.n107 10.6151
R1042 B.n496 B.n495 10.6151
R1043 B.n495 B.n494 10.6151
R1044 B.n494 B.n109 10.6151
R1045 B.n490 B.n109 10.6151
R1046 B.n490 B.n489 10.6151
R1047 B.n489 B.n488 10.6151
R1048 B.n488 B.n111 10.6151
R1049 B.n484 B.n111 10.6151
R1050 B.n484 B.n483 10.6151
R1051 B.n483 B.n482 10.6151
R1052 B.n482 B.n113 10.6151
R1053 B.n478 B.n113 10.6151
R1054 B.n478 B.n477 10.6151
R1055 B.n477 B.n476 10.6151
R1056 B.n476 B.n115 10.6151
R1057 B.n472 B.n115 10.6151
R1058 B.n472 B.n471 10.6151
R1059 B.n471 B.n470 10.6151
R1060 B.n470 B.n117 10.6151
R1061 B.n466 B.n117 10.6151
R1062 B.n466 B.n465 10.6151
R1063 B.n465 B.n464 10.6151
R1064 B.n464 B.n119 10.6151
R1065 B.n460 B.n119 10.6151
R1066 B.n460 B.n459 10.6151
R1067 B.n459 B.n458 10.6151
R1068 B.n458 B.n121 10.6151
R1069 B.n454 B.n121 10.6151
R1070 B.n454 B.n453 10.6151
R1071 B.n453 B.n452 10.6151
R1072 B.n452 B.n123 10.6151
R1073 B.n448 B.n123 10.6151
R1074 B.n205 B.n1 10.6151
R1075 B.n208 B.n205 10.6151
R1076 B.n209 B.n208 10.6151
R1077 B.n210 B.n209 10.6151
R1078 B.n210 B.n203 10.6151
R1079 B.n214 B.n203 10.6151
R1080 B.n215 B.n214 10.6151
R1081 B.n216 B.n215 10.6151
R1082 B.n216 B.n201 10.6151
R1083 B.n220 B.n201 10.6151
R1084 B.n221 B.n220 10.6151
R1085 B.n222 B.n221 10.6151
R1086 B.n222 B.n199 10.6151
R1087 B.n226 B.n199 10.6151
R1088 B.n227 B.n226 10.6151
R1089 B.n228 B.n227 10.6151
R1090 B.n228 B.n197 10.6151
R1091 B.n232 B.n197 10.6151
R1092 B.n233 B.n232 10.6151
R1093 B.n234 B.n233 10.6151
R1094 B.n234 B.n195 10.6151
R1095 B.n238 B.n195 10.6151
R1096 B.n239 B.n238 10.6151
R1097 B.n240 B.n239 10.6151
R1098 B.n240 B.n193 10.6151
R1099 B.n244 B.n193 10.6151
R1100 B.n245 B.n244 10.6151
R1101 B.n246 B.n245 10.6151
R1102 B.n246 B.n191 10.6151
R1103 B.n250 B.n191 10.6151
R1104 B.n251 B.n250 10.6151
R1105 B.n252 B.n251 10.6151
R1106 B.n252 B.n189 10.6151
R1107 B.n256 B.n189 10.6151
R1108 B.n257 B.n256 10.6151
R1109 B.n258 B.n187 10.6151
R1110 B.n262 B.n187 10.6151
R1111 B.n263 B.n262 10.6151
R1112 B.n264 B.n263 10.6151
R1113 B.n264 B.n185 10.6151
R1114 B.n268 B.n185 10.6151
R1115 B.n269 B.n268 10.6151
R1116 B.n270 B.n269 10.6151
R1117 B.n270 B.n183 10.6151
R1118 B.n274 B.n183 10.6151
R1119 B.n275 B.n274 10.6151
R1120 B.n276 B.n275 10.6151
R1121 B.n276 B.n181 10.6151
R1122 B.n280 B.n181 10.6151
R1123 B.n281 B.n280 10.6151
R1124 B.n282 B.n281 10.6151
R1125 B.n282 B.n179 10.6151
R1126 B.n286 B.n179 10.6151
R1127 B.n287 B.n286 10.6151
R1128 B.n288 B.n287 10.6151
R1129 B.n288 B.n177 10.6151
R1130 B.n292 B.n177 10.6151
R1131 B.n293 B.n292 10.6151
R1132 B.n294 B.n293 10.6151
R1133 B.n294 B.n175 10.6151
R1134 B.n298 B.n175 10.6151
R1135 B.n299 B.n298 10.6151
R1136 B.n300 B.n299 10.6151
R1137 B.n300 B.n173 10.6151
R1138 B.n304 B.n173 10.6151
R1139 B.n305 B.n304 10.6151
R1140 B.n306 B.n305 10.6151
R1141 B.n306 B.n171 10.6151
R1142 B.n310 B.n171 10.6151
R1143 B.n311 B.n310 10.6151
R1144 B.n312 B.n311 10.6151
R1145 B.n312 B.n169 10.6151
R1146 B.n316 B.n169 10.6151
R1147 B.n317 B.n316 10.6151
R1148 B.n318 B.n317 10.6151
R1149 B.n318 B.n167 10.6151
R1150 B.n322 B.n167 10.6151
R1151 B.n323 B.n322 10.6151
R1152 B.n324 B.n323 10.6151
R1153 B.n324 B.n165 10.6151
R1154 B.n328 B.n165 10.6151
R1155 B.n329 B.n328 10.6151
R1156 B.n330 B.n329 10.6151
R1157 B.n330 B.n163 10.6151
R1158 B.n334 B.n163 10.6151
R1159 B.n335 B.n334 10.6151
R1160 B.n336 B.n335 10.6151
R1161 B.n336 B.n161 10.6151
R1162 B.n340 B.n161 10.6151
R1163 B.n341 B.n340 10.6151
R1164 B.n345 B.n341 10.6151
R1165 B.n349 B.n159 10.6151
R1166 B.n350 B.n349 10.6151
R1167 B.n351 B.n350 10.6151
R1168 B.n351 B.n157 10.6151
R1169 B.n355 B.n157 10.6151
R1170 B.n356 B.n355 10.6151
R1171 B.n357 B.n356 10.6151
R1172 B.n357 B.n155 10.6151
R1173 B.n361 B.n155 10.6151
R1174 B.n364 B.n363 10.6151
R1175 B.n364 B.n151 10.6151
R1176 B.n368 B.n151 10.6151
R1177 B.n369 B.n368 10.6151
R1178 B.n370 B.n369 10.6151
R1179 B.n370 B.n149 10.6151
R1180 B.n374 B.n149 10.6151
R1181 B.n375 B.n374 10.6151
R1182 B.n376 B.n375 10.6151
R1183 B.n376 B.n147 10.6151
R1184 B.n380 B.n147 10.6151
R1185 B.n381 B.n380 10.6151
R1186 B.n382 B.n381 10.6151
R1187 B.n382 B.n145 10.6151
R1188 B.n386 B.n145 10.6151
R1189 B.n387 B.n386 10.6151
R1190 B.n388 B.n387 10.6151
R1191 B.n388 B.n143 10.6151
R1192 B.n392 B.n143 10.6151
R1193 B.n393 B.n392 10.6151
R1194 B.n394 B.n393 10.6151
R1195 B.n394 B.n141 10.6151
R1196 B.n398 B.n141 10.6151
R1197 B.n399 B.n398 10.6151
R1198 B.n400 B.n399 10.6151
R1199 B.n400 B.n139 10.6151
R1200 B.n404 B.n139 10.6151
R1201 B.n405 B.n404 10.6151
R1202 B.n406 B.n405 10.6151
R1203 B.n406 B.n137 10.6151
R1204 B.n410 B.n137 10.6151
R1205 B.n411 B.n410 10.6151
R1206 B.n412 B.n411 10.6151
R1207 B.n412 B.n135 10.6151
R1208 B.n416 B.n135 10.6151
R1209 B.n417 B.n416 10.6151
R1210 B.n418 B.n417 10.6151
R1211 B.n418 B.n133 10.6151
R1212 B.n422 B.n133 10.6151
R1213 B.n423 B.n422 10.6151
R1214 B.n424 B.n423 10.6151
R1215 B.n424 B.n131 10.6151
R1216 B.n428 B.n131 10.6151
R1217 B.n429 B.n428 10.6151
R1218 B.n430 B.n429 10.6151
R1219 B.n430 B.n129 10.6151
R1220 B.n434 B.n129 10.6151
R1221 B.n435 B.n434 10.6151
R1222 B.n436 B.n435 10.6151
R1223 B.n436 B.n127 10.6151
R1224 B.n440 B.n127 10.6151
R1225 B.n441 B.n440 10.6151
R1226 B.n442 B.n441 10.6151
R1227 B.n442 B.n125 10.6151
R1228 B.n446 B.n125 10.6151
R1229 B.n447 B.n446 10.6151
R1230 B.n52 B.n48 9.36635
R1231 B.n645 B.n644 9.36635
R1232 B.n345 B.n344 9.36635
R1233 B.n363 B.n362 9.36635
R1234 B.n801 B.n0 8.11757
R1235 B.n801 B.n1 8.11757
R1236 B.n659 B.n52 1.24928
R1237 B.n646 B.n645 1.24928
R1238 B.n344 B.n159 1.24928
R1239 B.n362 B.n361 1.24928
R1240 VP.n4 VP.t0 180.502
R1241 VP.n4 VP.t3 179.599
R1242 VP.n16 VP.n0 161.3
R1243 VP.n15 VP.n14 161.3
R1244 VP.n13 VP.n1 161.3
R1245 VP.n12 VP.n11 161.3
R1246 VP.n10 VP.n2 161.3
R1247 VP.n9 VP.n8 161.3
R1248 VP.n7 VP.n3 161.3
R1249 VP.n5 VP.t1 144.768
R1250 VP.n17 VP.t2 144.768
R1251 VP.n6 VP.n5 105.743
R1252 VP.n18 VP.n17 105.743
R1253 VP.n6 VP.n4 54.5998
R1254 VP.n11 VP.n10 40.577
R1255 VP.n11 VP.n1 40.577
R1256 VP.n9 VP.n3 24.5923
R1257 VP.n10 VP.n9 24.5923
R1258 VP.n15 VP.n1 24.5923
R1259 VP.n16 VP.n15 24.5923
R1260 VP.n5 VP.n3 5.16479
R1261 VP.n17 VP.n16 5.16479
R1262 VP.n7 VP.n6 0.278335
R1263 VP.n18 VP.n0 0.278335
R1264 VP.n8 VP.n7 0.189894
R1265 VP.n8 VP.n2 0.189894
R1266 VP.n12 VP.n2 0.189894
R1267 VP.n13 VP.n12 0.189894
R1268 VP.n14 VP.n13 0.189894
R1269 VP.n14 VP.n0 0.189894
R1270 VP VP.n18 0.153485
R1271 VDD1 VDD1.n1 119.373
R1272 VDD1 VDD1.n0 71.9753
R1273 VDD1.n0 VDD1.t3 1.8794
R1274 VDD1.n0 VDD1.t0 1.8794
R1275 VDD1.n1 VDD1.t2 1.8794
R1276 VDD1.n1 VDD1.t1 1.8794
C0 VTAIL VP 6.55873f
C1 VDD1 VN 0.149427f
C2 VN B 1.22812f
C3 VDD2 VP 0.412296f
C4 VDD1 w_n2896_n4428# 1.64587f
C5 w_n2896_n4428# B 11.0762f
C6 VDD1 VTAIL 6.67292f
C7 VTAIL B 6.8354f
C8 VDD2 VDD1 1.09032f
C9 VDD2 B 1.51021f
C10 VDD1 VP 7.09587f
C11 VP B 1.8484f
C12 VDD1 B 1.45341f
C13 w_n2896_n4428# VN 5.04501f
C14 VTAIL VN 6.54462f
C15 w_n2896_n4428# VTAIL 5.16168f
C16 VDD2 VN 6.83381f
C17 VN VP 7.36743f
C18 VDD2 w_n2896_n4428# 1.7082f
C19 w_n2896_n4428# VP 5.41801f
C20 VDD2 VTAIL 6.72901f
C21 VDD2 VSUBS 1.118715f
C22 VDD1 VSUBS 6.570849f
C23 VTAIL VSUBS 1.496128f
C24 VN VSUBS 5.76974f
C25 VP VSUBS 2.618875f
C26 B VSUBS 4.965461f
C27 w_n2896_n4428# VSUBS 0.156905p
C28 VDD1.t3 VSUBS 0.367055f
C29 VDD1.t0 VSUBS 0.367055f
C30 VDD1.n0 VSUBS 3.04678f
C31 VDD1.t2 VSUBS 0.367055f
C32 VDD1.t1 VSUBS 0.367055f
C33 VDD1.n1 VSUBS 3.99991f
C34 VP.n0 VSUBS 0.038331f
C35 VP.t2 VSUBS 3.98156f
C36 VP.n1 VSUBS 0.057483f
C37 VP.n2 VSUBS 0.029075f
C38 VP.n3 VSUBS 0.03289f
C39 VP.t3 VSUBS 4.28752f
C40 VP.t0 VSUBS 4.29519f
C41 VP.n4 VSUBS 4.54045f
C42 VP.t1 VSUBS 3.98156f
C43 VP.n5 VSUBS 1.47976f
C44 VP.n6 VSUBS 1.82684f
C45 VP.n7 VSUBS 0.038331f
C46 VP.n8 VSUBS 0.029075f
C47 VP.n9 VSUBS 0.053917f
C48 VP.n10 VSUBS 0.057483f
C49 VP.n11 VSUBS 0.023483f
C50 VP.n12 VSUBS 0.029075f
C51 VP.n13 VSUBS 0.029075f
C52 VP.n14 VSUBS 0.029075f
C53 VP.n15 VSUBS 0.053917f
C54 VP.n16 VSUBS 0.03289f
C55 VP.n17 VSUBS 1.47976f
C56 VP.n18 VSUBS 0.053606f
C57 B.n0 VSUBS 0.005241f
C58 B.n1 VSUBS 0.005241f
C59 B.n2 VSUBS 0.007752f
C60 B.n3 VSUBS 0.00594f
C61 B.n4 VSUBS 0.00594f
C62 B.n5 VSUBS 0.00594f
C63 B.n6 VSUBS 0.00594f
C64 B.n7 VSUBS 0.00594f
C65 B.n8 VSUBS 0.00594f
C66 B.n9 VSUBS 0.00594f
C67 B.n10 VSUBS 0.00594f
C68 B.n11 VSUBS 0.00594f
C69 B.n12 VSUBS 0.00594f
C70 B.n13 VSUBS 0.00594f
C71 B.n14 VSUBS 0.00594f
C72 B.n15 VSUBS 0.00594f
C73 B.n16 VSUBS 0.00594f
C74 B.n17 VSUBS 0.00594f
C75 B.n18 VSUBS 0.00594f
C76 B.n19 VSUBS 0.00594f
C77 B.n20 VSUBS 0.013936f
C78 B.n21 VSUBS 0.00594f
C79 B.n22 VSUBS 0.00594f
C80 B.n23 VSUBS 0.00594f
C81 B.n24 VSUBS 0.00594f
C82 B.n25 VSUBS 0.00594f
C83 B.n26 VSUBS 0.00594f
C84 B.n27 VSUBS 0.00594f
C85 B.n28 VSUBS 0.00594f
C86 B.n29 VSUBS 0.00594f
C87 B.n30 VSUBS 0.00594f
C88 B.n31 VSUBS 0.00594f
C89 B.n32 VSUBS 0.00594f
C90 B.n33 VSUBS 0.00594f
C91 B.n34 VSUBS 0.00594f
C92 B.n35 VSUBS 0.00594f
C93 B.n36 VSUBS 0.00594f
C94 B.n37 VSUBS 0.00594f
C95 B.n38 VSUBS 0.00594f
C96 B.n39 VSUBS 0.00594f
C97 B.n40 VSUBS 0.00594f
C98 B.n41 VSUBS 0.00594f
C99 B.n42 VSUBS 0.00594f
C100 B.n43 VSUBS 0.00594f
C101 B.n44 VSUBS 0.00594f
C102 B.n45 VSUBS 0.00594f
C103 B.n46 VSUBS 0.00594f
C104 B.n47 VSUBS 0.00594f
C105 B.n48 VSUBS 0.005591f
C106 B.n49 VSUBS 0.00594f
C107 B.t7 VSUBS 0.49424f
C108 B.t8 VSUBS 0.513405f
C109 B.t6 VSUBS 1.89466f
C110 B.n50 VSUBS 0.290186f
C111 B.n51 VSUBS 0.062138f
C112 B.n52 VSUBS 0.013763f
C113 B.n53 VSUBS 0.00594f
C114 B.n54 VSUBS 0.00594f
C115 B.n55 VSUBS 0.00594f
C116 B.n56 VSUBS 0.00594f
C117 B.t4 VSUBS 0.494223f
C118 B.t5 VSUBS 0.513391f
C119 B.t3 VSUBS 1.89466f
C120 B.n57 VSUBS 0.290199f
C121 B.n58 VSUBS 0.062155f
C122 B.n59 VSUBS 0.00594f
C123 B.n60 VSUBS 0.00594f
C124 B.n61 VSUBS 0.00594f
C125 B.n62 VSUBS 0.00594f
C126 B.n63 VSUBS 0.00594f
C127 B.n64 VSUBS 0.00594f
C128 B.n65 VSUBS 0.00594f
C129 B.n66 VSUBS 0.00594f
C130 B.n67 VSUBS 0.00594f
C131 B.n68 VSUBS 0.00594f
C132 B.n69 VSUBS 0.00594f
C133 B.n70 VSUBS 0.00594f
C134 B.n71 VSUBS 0.00594f
C135 B.n72 VSUBS 0.00594f
C136 B.n73 VSUBS 0.00594f
C137 B.n74 VSUBS 0.00594f
C138 B.n75 VSUBS 0.00594f
C139 B.n76 VSUBS 0.00594f
C140 B.n77 VSUBS 0.00594f
C141 B.n78 VSUBS 0.00594f
C142 B.n79 VSUBS 0.00594f
C143 B.n80 VSUBS 0.00594f
C144 B.n81 VSUBS 0.00594f
C145 B.n82 VSUBS 0.00594f
C146 B.n83 VSUBS 0.00594f
C147 B.n84 VSUBS 0.00594f
C148 B.n85 VSUBS 0.00594f
C149 B.n86 VSUBS 0.00594f
C150 B.n87 VSUBS 0.013319f
C151 B.n88 VSUBS 0.00594f
C152 B.n89 VSUBS 0.00594f
C153 B.n90 VSUBS 0.00594f
C154 B.n91 VSUBS 0.00594f
C155 B.n92 VSUBS 0.00594f
C156 B.n93 VSUBS 0.00594f
C157 B.n94 VSUBS 0.00594f
C158 B.n95 VSUBS 0.00594f
C159 B.n96 VSUBS 0.00594f
C160 B.n97 VSUBS 0.00594f
C161 B.n98 VSUBS 0.00594f
C162 B.n99 VSUBS 0.00594f
C163 B.n100 VSUBS 0.00594f
C164 B.n101 VSUBS 0.00594f
C165 B.n102 VSUBS 0.00594f
C166 B.n103 VSUBS 0.00594f
C167 B.n104 VSUBS 0.00594f
C168 B.n105 VSUBS 0.00594f
C169 B.n106 VSUBS 0.00594f
C170 B.n107 VSUBS 0.00594f
C171 B.n108 VSUBS 0.00594f
C172 B.n109 VSUBS 0.00594f
C173 B.n110 VSUBS 0.00594f
C174 B.n111 VSUBS 0.00594f
C175 B.n112 VSUBS 0.00594f
C176 B.n113 VSUBS 0.00594f
C177 B.n114 VSUBS 0.00594f
C178 B.n115 VSUBS 0.00594f
C179 B.n116 VSUBS 0.00594f
C180 B.n117 VSUBS 0.00594f
C181 B.n118 VSUBS 0.00594f
C182 B.n119 VSUBS 0.00594f
C183 B.n120 VSUBS 0.00594f
C184 B.n121 VSUBS 0.00594f
C185 B.n122 VSUBS 0.00594f
C186 B.n123 VSUBS 0.00594f
C187 B.n124 VSUBS 0.013936f
C188 B.n125 VSUBS 0.00594f
C189 B.n126 VSUBS 0.00594f
C190 B.n127 VSUBS 0.00594f
C191 B.n128 VSUBS 0.00594f
C192 B.n129 VSUBS 0.00594f
C193 B.n130 VSUBS 0.00594f
C194 B.n131 VSUBS 0.00594f
C195 B.n132 VSUBS 0.00594f
C196 B.n133 VSUBS 0.00594f
C197 B.n134 VSUBS 0.00594f
C198 B.n135 VSUBS 0.00594f
C199 B.n136 VSUBS 0.00594f
C200 B.n137 VSUBS 0.00594f
C201 B.n138 VSUBS 0.00594f
C202 B.n139 VSUBS 0.00594f
C203 B.n140 VSUBS 0.00594f
C204 B.n141 VSUBS 0.00594f
C205 B.n142 VSUBS 0.00594f
C206 B.n143 VSUBS 0.00594f
C207 B.n144 VSUBS 0.00594f
C208 B.n145 VSUBS 0.00594f
C209 B.n146 VSUBS 0.00594f
C210 B.n147 VSUBS 0.00594f
C211 B.n148 VSUBS 0.00594f
C212 B.n149 VSUBS 0.00594f
C213 B.n150 VSUBS 0.00594f
C214 B.n151 VSUBS 0.00594f
C215 B.n152 VSUBS 0.00594f
C216 B.t11 VSUBS 0.494223f
C217 B.t10 VSUBS 0.513391f
C218 B.t9 VSUBS 1.89466f
C219 B.n153 VSUBS 0.290199f
C220 B.n154 VSUBS 0.062155f
C221 B.n155 VSUBS 0.00594f
C222 B.n156 VSUBS 0.00594f
C223 B.n157 VSUBS 0.00594f
C224 B.n158 VSUBS 0.00594f
C225 B.n159 VSUBS 0.00332f
C226 B.n160 VSUBS 0.00594f
C227 B.n161 VSUBS 0.00594f
C228 B.n162 VSUBS 0.00594f
C229 B.n163 VSUBS 0.00594f
C230 B.n164 VSUBS 0.00594f
C231 B.n165 VSUBS 0.00594f
C232 B.n166 VSUBS 0.00594f
C233 B.n167 VSUBS 0.00594f
C234 B.n168 VSUBS 0.00594f
C235 B.n169 VSUBS 0.00594f
C236 B.n170 VSUBS 0.00594f
C237 B.n171 VSUBS 0.00594f
C238 B.n172 VSUBS 0.00594f
C239 B.n173 VSUBS 0.00594f
C240 B.n174 VSUBS 0.00594f
C241 B.n175 VSUBS 0.00594f
C242 B.n176 VSUBS 0.00594f
C243 B.n177 VSUBS 0.00594f
C244 B.n178 VSUBS 0.00594f
C245 B.n179 VSUBS 0.00594f
C246 B.n180 VSUBS 0.00594f
C247 B.n181 VSUBS 0.00594f
C248 B.n182 VSUBS 0.00594f
C249 B.n183 VSUBS 0.00594f
C250 B.n184 VSUBS 0.00594f
C251 B.n185 VSUBS 0.00594f
C252 B.n186 VSUBS 0.00594f
C253 B.n187 VSUBS 0.00594f
C254 B.n188 VSUBS 0.013319f
C255 B.n189 VSUBS 0.00594f
C256 B.n190 VSUBS 0.00594f
C257 B.n191 VSUBS 0.00594f
C258 B.n192 VSUBS 0.00594f
C259 B.n193 VSUBS 0.00594f
C260 B.n194 VSUBS 0.00594f
C261 B.n195 VSUBS 0.00594f
C262 B.n196 VSUBS 0.00594f
C263 B.n197 VSUBS 0.00594f
C264 B.n198 VSUBS 0.00594f
C265 B.n199 VSUBS 0.00594f
C266 B.n200 VSUBS 0.00594f
C267 B.n201 VSUBS 0.00594f
C268 B.n202 VSUBS 0.00594f
C269 B.n203 VSUBS 0.00594f
C270 B.n204 VSUBS 0.00594f
C271 B.n205 VSUBS 0.00594f
C272 B.n206 VSUBS 0.00594f
C273 B.n207 VSUBS 0.00594f
C274 B.n208 VSUBS 0.00594f
C275 B.n209 VSUBS 0.00594f
C276 B.n210 VSUBS 0.00594f
C277 B.n211 VSUBS 0.00594f
C278 B.n212 VSUBS 0.00594f
C279 B.n213 VSUBS 0.00594f
C280 B.n214 VSUBS 0.00594f
C281 B.n215 VSUBS 0.00594f
C282 B.n216 VSUBS 0.00594f
C283 B.n217 VSUBS 0.00594f
C284 B.n218 VSUBS 0.00594f
C285 B.n219 VSUBS 0.00594f
C286 B.n220 VSUBS 0.00594f
C287 B.n221 VSUBS 0.00594f
C288 B.n222 VSUBS 0.00594f
C289 B.n223 VSUBS 0.00594f
C290 B.n224 VSUBS 0.00594f
C291 B.n225 VSUBS 0.00594f
C292 B.n226 VSUBS 0.00594f
C293 B.n227 VSUBS 0.00594f
C294 B.n228 VSUBS 0.00594f
C295 B.n229 VSUBS 0.00594f
C296 B.n230 VSUBS 0.00594f
C297 B.n231 VSUBS 0.00594f
C298 B.n232 VSUBS 0.00594f
C299 B.n233 VSUBS 0.00594f
C300 B.n234 VSUBS 0.00594f
C301 B.n235 VSUBS 0.00594f
C302 B.n236 VSUBS 0.00594f
C303 B.n237 VSUBS 0.00594f
C304 B.n238 VSUBS 0.00594f
C305 B.n239 VSUBS 0.00594f
C306 B.n240 VSUBS 0.00594f
C307 B.n241 VSUBS 0.00594f
C308 B.n242 VSUBS 0.00594f
C309 B.n243 VSUBS 0.00594f
C310 B.n244 VSUBS 0.00594f
C311 B.n245 VSUBS 0.00594f
C312 B.n246 VSUBS 0.00594f
C313 B.n247 VSUBS 0.00594f
C314 B.n248 VSUBS 0.00594f
C315 B.n249 VSUBS 0.00594f
C316 B.n250 VSUBS 0.00594f
C317 B.n251 VSUBS 0.00594f
C318 B.n252 VSUBS 0.00594f
C319 B.n253 VSUBS 0.00594f
C320 B.n254 VSUBS 0.00594f
C321 B.n255 VSUBS 0.00594f
C322 B.n256 VSUBS 0.00594f
C323 B.n257 VSUBS 0.013319f
C324 B.n258 VSUBS 0.013936f
C325 B.n259 VSUBS 0.013936f
C326 B.n260 VSUBS 0.00594f
C327 B.n261 VSUBS 0.00594f
C328 B.n262 VSUBS 0.00594f
C329 B.n263 VSUBS 0.00594f
C330 B.n264 VSUBS 0.00594f
C331 B.n265 VSUBS 0.00594f
C332 B.n266 VSUBS 0.00594f
C333 B.n267 VSUBS 0.00594f
C334 B.n268 VSUBS 0.00594f
C335 B.n269 VSUBS 0.00594f
C336 B.n270 VSUBS 0.00594f
C337 B.n271 VSUBS 0.00594f
C338 B.n272 VSUBS 0.00594f
C339 B.n273 VSUBS 0.00594f
C340 B.n274 VSUBS 0.00594f
C341 B.n275 VSUBS 0.00594f
C342 B.n276 VSUBS 0.00594f
C343 B.n277 VSUBS 0.00594f
C344 B.n278 VSUBS 0.00594f
C345 B.n279 VSUBS 0.00594f
C346 B.n280 VSUBS 0.00594f
C347 B.n281 VSUBS 0.00594f
C348 B.n282 VSUBS 0.00594f
C349 B.n283 VSUBS 0.00594f
C350 B.n284 VSUBS 0.00594f
C351 B.n285 VSUBS 0.00594f
C352 B.n286 VSUBS 0.00594f
C353 B.n287 VSUBS 0.00594f
C354 B.n288 VSUBS 0.00594f
C355 B.n289 VSUBS 0.00594f
C356 B.n290 VSUBS 0.00594f
C357 B.n291 VSUBS 0.00594f
C358 B.n292 VSUBS 0.00594f
C359 B.n293 VSUBS 0.00594f
C360 B.n294 VSUBS 0.00594f
C361 B.n295 VSUBS 0.00594f
C362 B.n296 VSUBS 0.00594f
C363 B.n297 VSUBS 0.00594f
C364 B.n298 VSUBS 0.00594f
C365 B.n299 VSUBS 0.00594f
C366 B.n300 VSUBS 0.00594f
C367 B.n301 VSUBS 0.00594f
C368 B.n302 VSUBS 0.00594f
C369 B.n303 VSUBS 0.00594f
C370 B.n304 VSUBS 0.00594f
C371 B.n305 VSUBS 0.00594f
C372 B.n306 VSUBS 0.00594f
C373 B.n307 VSUBS 0.00594f
C374 B.n308 VSUBS 0.00594f
C375 B.n309 VSUBS 0.00594f
C376 B.n310 VSUBS 0.00594f
C377 B.n311 VSUBS 0.00594f
C378 B.n312 VSUBS 0.00594f
C379 B.n313 VSUBS 0.00594f
C380 B.n314 VSUBS 0.00594f
C381 B.n315 VSUBS 0.00594f
C382 B.n316 VSUBS 0.00594f
C383 B.n317 VSUBS 0.00594f
C384 B.n318 VSUBS 0.00594f
C385 B.n319 VSUBS 0.00594f
C386 B.n320 VSUBS 0.00594f
C387 B.n321 VSUBS 0.00594f
C388 B.n322 VSUBS 0.00594f
C389 B.n323 VSUBS 0.00594f
C390 B.n324 VSUBS 0.00594f
C391 B.n325 VSUBS 0.00594f
C392 B.n326 VSUBS 0.00594f
C393 B.n327 VSUBS 0.00594f
C394 B.n328 VSUBS 0.00594f
C395 B.n329 VSUBS 0.00594f
C396 B.n330 VSUBS 0.00594f
C397 B.n331 VSUBS 0.00594f
C398 B.n332 VSUBS 0.00594f
C399 B.n333 VSUBS 0.00594f
C400 B.n334 VSUBS 0.00594f
C401 B.n335 VSUBS 0.00594f
C402 B.n336 VSUBS 0.00594f
C403 B.n337 VSUBS 0.00594f
C404 B.n338 VSUBS 0.00594f
C405 B.n339 VSUBS 0.00594f
C406 B.n340 VSUBS 0.00594f
C407 B.n341 VSUBS 0.00594f
C408 B.t2 VSUBS 0.49424f
C409 B.t1 VSUBS 0.513405f
C410 B.t0 VSUBS 1.89466f
C411 B.n342 VSUBS 0.290186f
C412 B.n343 VSUBS 0.062138f
C413 B.n344 VSUBS 0.013763f
C414 B.n345 VSUBS 0.005591f
C415 B.n346 VSUBS 0.00594f
C416 B.n347 VSUBS 0.00594f
C417 B.n348 VSUBS 0.00594f
C418 B.n349 VSUBS 0.00594f
C419 B.n350 VSUBS 0.00594f
C420 B.n351 VSUBS 0.00594f
C421 B.n352 VSUBS 0.00594f
C422 B.n353 VSUBS 0.00594f
C423 B.n354 VSUBS 0.00594f
C424 B.n355 VSUBS 0.00594f
C425 B.n356 VSUBS 0.00594f
C426 B.n357 VSUBS 0.00594f
C427 B.n358 VSUBS 0.00594f
C428 B.n359 VSUBS 0.00594f
C429 B.n360 VSUBS 0.00594f
C430 B.n361 VSUBS 0.00332f
C431 B.n362 VSUBS 0.013763f
C432 B.n363 VSUBS 0.005591f
C433 B.n364 VSUBS 0.00594f
C434 B.n365 VSUBS 0.00594f
C435 B.n366 VSUBS 0.00594f
C436 B.n367 VSUBS 0.00594f
C437 B.n368 VSUBS 0.00594f
C438 B.n369 VSUBS 0.00594f
C439 B.n370 VSUBS 0.00594f
C440 B.n371 VSUBS 0.00594f
C441 B.n372 VSUBS 0.00594f
C442 B.n373 VSUBS 0.00594f
C443 B.n374 VSUBS 0.00594f
C444 B.n375 VSUBS 0.00594f
C445 B.n376 VSUBS 0.00594f
C446 B.n377 VSUBS 0.00594f
C447 B.n378 VSUBS 0.00594f
C448 B.n379 VSUBS 0.00594f
C449 B.n380 VSUBS 0.00594f
C450 B.n381 VSUBS 0.00594f
C451 B.n382 VSUBS 0.00594f
C452 B.n383 VSUBS 0.00594f
C453 B.n384 VSUBS 0.00594f
C454 B.n385 VSUBS 0.00594f
C455 B.n386 VSUBS 0.00594f
C456 B.n387 VSUBS 0.00594f
C457 B.n388 VSUBS 0.00594f
C458 B.n389 VSUBS 0.00594f
C459 B.n390 VSUBS 0.00594f
C460 B.n391 VSUBS 0.00594f
C461 B.n392 VSUBS 0.00594f
C462 B.n393 VSUBS 0.00594f
C463 B.n394 VSUBS 0.00594f
C464 B.n395 VSUBS 0.00594f
C465 B.n396 VSUBS 0.00594f
C466 B.n397 VSUBS 0.00594f
C467 B.n398 VSUBS 0.00594f
C468 B.n399 VSUBS 0.00594f
C469 B.n400 VSUBS 0.00594f
C470 B.n401 VSUBS 0.00594f
C471 B.n402 VSUBS 0.00594f
C472 B.n403 VSUBS 0.00594f
C473 B.n404 VSUBS 0.00594f
C474 B.n405 VSUBS 0.00594f
C475 B.n406 VSUBS 0.00594f
C476 B.n407 VSUBS 0.00594f
C477 B.n408 VSUBS 0.00594f
C478 B.n409 VSUBS 0.00594f
C479 B.n410 VSUBS 0.00594f
C480 B.n411 VSUBS 0.00594f
C481 B.n412 VSUBS 0.00594f
C482 B.n413 VSUBS 0.00594f
C483 B.n414 VSUBS 0.00594f
C484 B.n415 VSUBS 0.00594f
C485 B.n416 VSUBS 0.00594f
C486 B.n417 VSUBS 0.00594f
C487 B.n418 VSUBS 0.00594f
C488 B.n419 VSUBS 0.00594f
C489 B.n420 VSUBS 0.00594f
C490 B.n421 VSUBS 0.00594f
C491 B.n422 VSUBS 0.00594f
C492 B.n423 VSUBS 0.00594f
C493 B.n424 VSUBS 0.00594f
C494 B.n425 VSUBS 0.00594f
C495 B.n426 VSUBS 0.00594f
C496 B.n427 VSUBS 0.00594f
C497 B.n428 VSUBS 0.00594f
C498 B.n429 VSUBS 0.00594f
C499 B.n430 VSUBS 0.00594f
C500 B.n431 VSUBS 0.00594f
C501 B.n432 VSUBS 0.00594f
C502 B.n433 VSUBS 0.00594f
C503 B.n434 VSUBS 0.00594f
C504 B.n435 VSUBS 0.00594f
C505 B.n436 VSUBS 0.00594f
C506 B.n437 VSUBS 0.00594f
C507 B.n438 VSUBS 0.00594f
C508 B.n439 VSUBS 0.00594f
C509 B.n440 VSUBS 0.00594f
C510 B.n441 VSUBS 0.00594f
C511 B.n442 VSUBS 0.00594f
C512 B.n443 VSUBS 0.00594f
C513 B.n444 VSUBS 0.00594f
C514 B.n445 VSUBS 0.00594f
C515 B.n446 VSUBS 0.00594f
C516 B.n447 VSUBS 0.013213f
C517 B.n448 VSUBS 0.014042f
C518 B.n449 VSUBS 0.013319f
C519 B.n450 VSUBS 0.00594f
C520 B.n451 VSUBS 0.00594f
C521 B.n452 VSUBS 0.00594f
C522 B.n453 VSUBS 0.00594f
C523 B.n454 VSUBS 0.00594f
C524 B.n455 VSUBS 0.00594f
C525 B.n456 VSUBS 0.00594f
C526 B.n457 VSUBS 0.00594f
C527 B.n458 VSUBS 0.00594f
C528 B.n459 VSUBS 0.00594f
C529 B.n460 VSUBS 0.00594f
C530 B.n461 VSUBS 0.00594f
C531 B.n462 VSUBS 0.00594f
C532 B.n463 VSUBS 0.00594f
C533 B.n464 VSUBS 0.00594f
C534 B.n465 VSUBS 0.00594f
C535 B.n466 VSUBS 0.00594f
C536 B.n467 VSUBS 0.00594f
C537 B.n468 VSUBS 0.00594f
C538 B.n469 VSUBS 0.00594f
C539 B.n470 VSUBS 0.00594f
C540 B.n471 VSUBS 0.00594f
C541 B.n472 VSUBS 0.00594f
C542 B.n473 VSUBS 0.00594f
C543 B.n474 VSUBS 0.00594f
C544 B.n475 VSUBS 0.00594f
C545 B.n476 VSUBS 0.00594f
C546 B.n477 VSUBS 0.00594f
C547 B.n478 VSUBS 0.00594f
C548 B.n479 VSUBS 0.00594f
C549 B.n480 VSUBS 0.00594f
C550 B.n481 VSUBS 0.00594f
C551 B.n482 VSUBS 0.00594f
C552 B.n483 VSUBS 0.00594f
C553 B.n484 VSUBS 0.00594f
C554 B.n485 VSUBS 0.00594f
C555 B.n486 VSUBS 0.00594f
C556 B.n487 VSUBS 0.00594f
C557 B.n488 VSUBS 0.00594f
C558 B.n489 VSUBS 0.00594f
C559 B.n490 VSUBS 0.00594f
C560 B.n491 VSUBS 0.00594f
C561 B.n492 VSUBS 0.00594f
C562 B.n493 VSUBS 0.00594f
C563 B.n494 VSUBS 0.00594f
C564 B.n495 VSUBS 0.00594f
C565 B.n496 VSUBS 0.00594f
C566 B.n497 VSUBS 0.00594f
C567 B.n498 VSUBS 0.00594f
C568 B.n499 VSUBS 0.00594f
C569 B.n500 VSUBS 0.00594f
C570 B.n501 VSUBS 0.00594f
C571 B.n502 VSUBS 0.00594f
C572 B.n503 VSUBS 0.00594f
C573 B.n504 VSUBS 0.00594f
C574 B.n505 VSUBS 0.00594f
C575 B.n506 VSUBS 0.00594f
C576 B.n507 VSUBS 0.00594f
C577 B.n508 VSUBS 0.00594f
C578 B.n509 VSUBS 0.00594f
C579 B.n510 VSUBS 0.00594f
C580 B.n511 VSUBS 0.00594f
C581 B.n512 VSUBS 0.00594f
C582 B.n513 VSUBS 0.00594f
C583 B.n514 VSUBS 0.00594f
C584 B.n515 VSUBS 0.00594f
C585 B.n516 VSUBS 0.00594f
C586 B.n517 VSUBS 0.00594f
C587 B.n518 VSUBS 0.00594f
C588 B.n519 VSUBS 0.00594f
C589 B.n520 VSUBS 0.00594f
C590 B.n521 VSUBS 0.00594f
C591 B.n522 VSUBS 0.00594f
C592 B.n523 VSUBS 0.00594f
C593 B.n524 VSUBS 0.00594f
C594 B.n525 VSUBS 0.00594f
C595 B.n526 VSUBS 0.00594f
C596 B.n527 VSUBS 0.00594f
C597 B.n528 VSUBS 0.00594f
C598 B.n529 VSUBS 0.00594f
C599 B.n530 VSUBS 0.00594f
C600 B.n531 VSUBS 0.00594f
C601 B.n532 VSUBS 0.00594f
C602 B.n533 VSUBS 0.00594f
C603 B.n534 VSUBS 0.00594f
C604 B.n535 VSUBS 0.00594f
C605 B.n536 VSUBS 0.00594f
C606 B.n537 VSUBS 0.00594f
C607 B.n538 VSUBS 0.00594f
C608 B.n539 VSUBS 0.00594f
C609 B.n540 VSUBS 0.00594f
C610 B.n541 VSUBS 0.00594f
C611 B.n542 VSUBS 0.00594f
C612 B.n543 VSUBS 0.00594f
C613 B.n544 VSUBS 0.00594f
C614 B.n545 VSUBS 0.00594f
C615 B.n546 VSUBS 0.00594f
C616 B.n547 VSUBS 0.00594f
C617 B.n548 VSUBS 0.00594f
C618 B.n549 VSUBS 0.00594f
C619 B.n550 VSUBS 0.00594f
C620 B.n551 VSUBS 0.00594f
C621 B.n552 VSUBS 0.00594f
C622 B.n553 VSUBS 0.00594f
C623 B.n554 VSUBS 0.00594f
C624 B.n555 VSUBS 0.00594f
C625 B.n556 VSUBS 0.00594f
C626 B.n557 VSUBS 0.00594f
C627 B.n558 VSUBS 0.013319f
C628 B.n559 VSUBS 0.013936f
C629 B.n560 VSUBS 0.013936f
C630 B.n561 VSUBS 0.00594f
C631 B.n562 VSUBS 0.00594f
C632 B.n563 VSUBS 0.00594f
C633 B.n564 VSUBS 0.00594f
C634 B.n565 VSUBS 0.00594f
C635 B.n566 VSUBS 0.00594f
C636 B.n567 VSUBS 0.00594f
C637 B.n568 VSUBS 0.00594f
C638 B.n569 VSUBS 0.00594f
C639 B.n570 VSUBS 0.00594f
C640 B.n571 VSUBS 0.00594f
C641 B.n572 VSUBS 0.00594f
C642 B.n573 VSUBS 0.00594f
C643 B.n574 VSUBS 0.00594f
C644 B.n575 VSUBS 0.00594f
C645 B.n576 VSUBS 0.00594f
C646 B.n577 VSUBS 0.00594f
C647 B.n578 VSUBS 0.00594f
C648 B.n579 VSUBS 0.00594f
C649 B.n580 VSUBS 0.00594f
C650 B.n581 VSUBS 0.00594f
C651 B.n582 VSUBS 0.00594f
C652 B.n583 VSUBS 0.00594f
C653 B.n584 VSUBS 0.00594f
C654 B.n585 VSUBS 0.00594f
C655 B.n586 VSUBS 0.00594f
C656 B.n587 VSUBS 0.00594f
C657 B.n588 VSUBS 0.00594f
C658 B.n589 VSUBS 0.00594f
C659 B.n590 VSUBS 0.00594f
C660 B.n591 VSUBS 0.00594f
C661 B.n592 VSUBS 0.00594f
C662 B.n593 VSUBS 0.00594f
C663 B.n594 VSUBS 0.00594f
C664 B.n595 VSUBS 0.00594f
C665 B.n596 VSUBS 0.00594f
C666 B.n597 VSUBS 0.00594f
C667 B.n598 VSUBS 0.00594f
C668 B.n599 VSUBS 0.00594f
C669 B.n600 VSUBS 0.00594f
C670 B.n601 VSUBS 0.00594f
C671 B.n602 VSUBS 0.00594f
C672 B.n603 VSUBS 0.00594f
C673 B.n604 VSUBS 0.00594f
C674 B.n605 VSUBS 0.00594f
C675 B.n606 VSUBS 0.00594f
C676 B.n607 VSUBS 0.00594f
C677 B.n608 VSUBS 0.00594f
C678 B.n609 VSUBS 0.00594f
C679 B.n610 VSUBS 0.00594f
C680 B.n611 VSUBS 0.00594f
C681 B.n612 VSUBS 0.00594f
C682 B.n613 VSUBS 0.00594f
C683 B.n614 VSUBS 0.00594f
C684 B.n615 VSUBS 0.00594f
C685 B.n616 VSUBS 0.00594f
C686 B.n617 VSUBS 0.00594f
C687 B.n618 VSUBS 0.00594f
C688 B.n619 VSUBS 0.00594f
C689 B.n620 VSUBS 0.00594f
C690 B.n621 VSUBS 0.00594f
C691 B.n622 VSUBS 0.00594f
C692 B.n623 VSUBS 0.00594f
C693 B.n624 VSUBS 0.00594f
C694 B.n625 VSUBS 0.00594f
C695 B.n626 VSUBS 0.00594f
C696 B.n627 VSUBS 0.00594f
C697 B.n628 VSUBS 0.00594f
C698 B.n629 VSUBS 0.00594f
C699 B.n630 VSUBS 0.00594f
C700 B.n631 VSUBS 0.00594f
C701 B.n632 VSUBS 0.00594f
C702 B.n633 VSUBS 0.00594f
C703 B.n634 VSUBS 0.00594f
C704 B.n635 VSUBS 0.00594f
C705 B.n636 VSUBS 0.00594f
C706 B.n637 VSUBS 0.00594f
C707 B.n638 VSUBS 0.00594f
C708 B.n639 VSUBS 0.00594f
C709 B.n640 VSUBS 0.00594f
C710 B.n641 VSUBS 0.00594f
C711 B.n642 VSUBS 0.00594f
C712 B.n643 VSUBS 0.00594f
C713 B.n644 VSUBS 0.005591f
C714 B.n645 VSUBS 0.013763f
C715 B.n646 VSUBS 0.00332f
C716 B.n647 VSUBS 0.00594f
C717 B.n648 VSUBS 0.00594f
C718 B.n649 VSUBS 0.00594f
C719 B.n650 VSUBS 0.00594f
C720 B.n651 VSUBS 0.00594f
C721 B.n652 VSUBS 0.00594f
C722 B.n653 VSUBS 0.00594f
C723 B.n654 VSUBS 0.00594f
C724 B.n655 VSUBS 0.00594f
C725 B.n656 VSUBS 0.00594f
C726 B.n657 VSUBS 0.00594f
C727 B.n658 VSUBS 0.00594f
C728 B.n659 VSUBS 0.00332f
C729 B.n660 VSUBS 0.00594f
C730 B.n661 VSUBS 0.00594f
C731 B.n662 VSUBS 0.00594f
C732 B.n663 VSUBS 0.00594f
C733 B.n664 VSUBS 0.00594f
C734 B.n665 VSUBS 0.00594f
C735 B.n666 VSUBS 0.00594f
C736 B.n667 VSUBS 0.00594f
C737 B.n668 VSUBS 0.00594f
C738 B.n669 VSUBS 0.00594f
C739 B.n670 VSUBS 0.00594f
C740 B.n671 VSUBS 0.00594f
C741 B.n672 VSUBS 0.00594f
C742 B.n673 VSUBS 0.00594f
C743 B.n674 VSUBS 0.00594f
C744 B.n675 VSUBS 0.00594f
C745 B.n676 VSUBS 0.00594f
C746 B.n677 VSUBS 0.00594f
C747 B.n678 VSUBS 0.00594f
C748 B.n679 VSUBS 0.00594f
C749 B.n680 VSUBS 0.00594f
C750 B.n681 VSUBS 0.00594f
C751 B.n682 VSUBS 0.00594f
C752 B.n683 VSUBS 0.00594f
C753 B.n684 VSUBS 0.00594f
C754 B.n685 VSUBS 0.00594f
C755 B.n686 VSUBS 0.00594f
C756 B.n687 VSUBS 0.00594f
C757 B.n688 VSUBS 0.00594f
C758 B.n689 VSUBS 0.00594f
C759 B.n690 VSUBS 0.00594f
C760 B.n691 VSUBS 0.00594f
C761 B.n692 VSUBS 0.00594f
C762 B.n693 VSUBS 0.00594f
C763 B.n694 VSUBS 0.00594f
C764 B.n695 VSUBS 0.00594f
C765 B.n696 VSUBS 0.00594f
C766 B.n697 VSUBS 0.00594f
C767 B.n698 VSUBS 0.00594f
C768 B.n699 VSUBS 0.00594f
C769 B.n700 VSUBS 0.00594f
C770 B.n701 VSUBS 0.00594f
C771 B.n702 VSUBS 0.00594f
C772 B.n703 VSUBS 0.00594f
C773 B.n704 VSUBS 0.00594f
C774 B.n705 VSUBS 0.00594f
C775 B.n706 VSUBS 0.00594f
C776 B.n707 VSUBS 0.00594f
C777 B.n708 VSUBS 0.00594f
C778 B.n709 VSUBS 0.00594f
C779 B.n710 VSUBS 0.00594f
C780 B.n711 VSUBS 0.00594f
C781 B.n712 VSUBS 0.00594f
C782 B.n713 VSUBS 0.00594f
C783 B.n714 VSUBS 0.00594f
C784 B.n715 VSUBS 0.00594f
C785 B.n716 VSUBS 0.00594f
C786 B.n717 VSUBS 0.00594f
C787 B.n718 VSUBS 0.00594f
C788 B.n719 VSUBS 0.00594f
C789 B.n720 VSUBS 0.00594f
C790 B.n721 VSUBS 0.00594f
C791 B.n722 VSUBS 0.00594f
C792 B.n723 VSUBS 0.00594f
C793 B.n724 VSUBS 0.00594f
C794 B.n725 VSUBS 0.00594f
C795 B.n726 VSUBS 0.00594f
C796 B.n727 VSUBS 0.00594f
C797 B.n728 VSUBS 0.00594f
C798 B.n729 VSUBS 0.00594f
C799 B.n730 VSUBS 0.00594f
C800 B.n731 VSUBS 0.00594f
C801 B.n732 VSUBS 0.00594f
C802 B.n733 VSUBS 0.00594f
C803 B.n734 VSUBS 0.00594f
C804 B.n735 VSUBS 0.00594f
C805 B.n736 VSUBS 0.00594f
C806 B.n737 VSUBS 0.00594f
C807 B.n738 VSUBS 0.00594f
C808 B.n739 VSUBS 0.00594f
C809 B.n740 VSUBS 0.00594f
C810 B.n741 VSUBS 0.00594f
C811 B.n742 VSUBS 0.00594f
C812 B.n743 VSUBS 0.00594f
C813 B.n744 VSUBS 0.00594f
C814 B.n745 VSUBS 0.013936f
C815 B.n746 VSUBS 0.013319f
C816 B.n747 VSUBS 0.013319f
C817 B.n748 VSUBS 0.00594f
C818 B.n749 VSUBS 0.00594f
C819 B.n750 VSUBS 0.00594f
C820 B.n751 VSUBS 0.00594f
C821 B.n752 VSUBS 0.00594f
C822 B.n753 VSUBS 0.00594f
C823 B.n754 VSUBS 0.00594f
C824 B.n755 VSUBS 0.00594f
C825 B.n756 VSUBS 0.00594f
C826 B.n757 VSUBS 0.00594f
C827 B.n758 VSUBS 0.00594f
C828 B.n759 VSUBS 0.00594f
C829 B.n760 VSUBS 0.00594f
C830 B.n761 VSUBS 0.00594f
C831 B.n762 VSUBS 0.00594f
C832 B.n763 VSUBS 0.00594f
C833 B.n764 VSUBS 0.00594f
C834 B.n765 VSUBS 0.00594f
C835 B.n766 VSUBS 0.00594f
C836 B.n767 VSUBS 0.00594f
C837 B.n768 VSUBS 0.00594f
C838 B.n769 VSUBS 0.00594f
C839 B.n770 VSUBS 0.00594f
C840 B.n771 VSUBS 0.00594f
C841 B.n772 VSUBS 0.00594f
C842 B.n773 VSUBS 0.00594f
C843 B.n774 VSUBS 0.00594f
C844 B.n775 VSUBS 0.00594f
C845 B.n776 VSUBS 0.00594f
C846 B.n777 VSUBS 0.00594f
C847 B.n778 VSUBS 0.00594f
C848 B.n779 VSUBS 0.00594f
C849 B.n780 VSUBS 0.00594f
C850 B.n781 VSUBS 0.00594f
C851 B.n782 VSUBS 0.00594f
C852 B.n783 VSUBS 0.00594f
C853 B.n784 VSUBS 0.00594f
C854 B.n785 VSUBS 0.00594f
C855 B.n786 VSUBS 0.00594f
C856 B.n787 VSUBS 0.00594f
C857 B.n788 VSUBS 0.00594f
C858 B.n789 VSUBS 0.00594f
C859 B.n790 VSUBS 0.00594f
C860 B.n791 VSUBS 0.00594f
C861 B.n792 VSUBS 0.00594f
C862 B.n793 VSUBS 0.00594f
C863 B.n794 VSUBS 0.00594f
C864 B.n795 VSUBS 0.00594f
C865 B.n796 VSUBS 0.00594f
C866 B.n797 VSUBS 0.00594f
C867 B.n798 VSUBS 0.00594f
C868 B.n799 VSUBS 0.007752f
C869 B.n800 VSUBS 0.008258f
C870 B.n801 VSUBS 0.016421f
C871 VDD2.t2 VSUBS 0.361675f
C872 VDD2.t3 VSUBS 0.361675f
C873 VDD2.n0 VSUBS 3.91447f
C874 VDD2.t0 VSUBS 0.361675f
C875 VDD2.t1 VSUBS 0.361675f
C876 VDD2.n1 VSUBS 3.0015f
C877 VDD2.n2 VSUBS 4.895741f
C878 VTAIL.t4 VSUBS 3.17117f
C879 VTAIL.n0 VSUBS 0.766931f
C880 VTAIL.t2 VSUBS 3.17117f
C881 VTAIL.n1 VSUBS 0.863198f
C882 VTAIL.t3 VSUBS 3.17117f
C883 VTAIL.n2 VSUBS 2.41946f
C884 VTAIL.t5 VSUBS 3.1712f
C885 VTAIL.n3 VSUBS 2.41943f
C886 VTAIL.t6 VSUBS 3.1712f
C887 VTAIL.n4 VSUBS 0.863175f
C888 VTAIL.t1 VSUBS 3.1712f
C889 VTAIL.n5 VSUBS 0.863175f
C890 VTAIL.t0 VSUBS 3.17117f
C891 VTAIL.n6 VSUBS 2.41945f
C892 VTAIL.t7 VSUBS 3.17117f
C893 VTAIL.n7 VSUBS 2.31473f
C894 VN.t1 VSUBS 4.15911f
C895 VN.t0 VSUBS 4.15168f
C896 VN.n0 VSUBS 2.61458f
C897 VN.t2 VSUBS 4.15911f
C898 VN.t3 VSUBS 4.15168f
C899 VN.n1 VSUBS 4.41135f
.ends

