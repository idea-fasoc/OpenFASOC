* NGSPICE file created from diff_pair_sample_0919.ext - technology: sky130A

.subckt diff_pair_sample_0919 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t9 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=3.5802 ps=19.14 w=9.18 l=1.63
X1 VDD1.t7 VP.t0 VTAIL.t5 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=3.5802 ps=19.14 w=9.18 l=1.63
X2 B.t11 B.t9 B.t10 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=3.5802 pd=19.14 as=0 ps=0 w=9.18 l=1.63
X3 VDD2.t6 VN.t1 VTAIL.t8 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=1.5147 ps=9.51 w=9.18 l=1.63
X4 VDD1.t6 VP.t1 VTAIL.t1 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=1.5147 ps=9.51 w=9.18 l=1.63
X5 VTAIL.t0 VP.t2 VDD1.t5 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=3.5802 pd=19.14 as=1.5147 ps=9.51 w=9.18 l=1.63
X6 VDD1.t4 VP.t3 VTAIL.t3 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=1.5147 ps=9.51 w=9.18 l=1.63
X7 VDD2.t5 VN.t2 VTAIL.t12 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=3.5802 ps=19.14 w=9.18 l=1.63
X8 VTAIL.t15 VN.t3 VDD2.t4 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=3.5802 pd=19.14 as=1.5147 ps=9.51 w=9.18 l=1.63
X9 B.t8 B.t6 B.t7 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=3.5802 pd=19.14 as=0 ps=0 w=9.18 l=1.63
X10 VTAIL.t4 VP.t4 VDD1.t3 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=1.5147 ps=9.51 w=9.18 l=1.63
X11 B.t5 B.t3 B.t4 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=3.5802 pd=19.14 as=0 ps=0 w=9.18 l=1.63
X12 VDD2.t3 VN.t4 VTAIL.t14 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=1.5147 ps=9.51 w=9.18 l=1.63
X13 VDD1.t2 VP.t5 VTAIL.t7 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=3.5802 ps=19.14 w=9.18 l=1.63
X14 VTAIL.t13 VN.t5 VDD2.t2 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=1.5147 ps=9.51 w=9.18 l=1.63
X15 VTAIL.t10 VN.t6 VDD2.t1 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=3.5802 pd=19.14 as=1.5147 ps=9.51 w=9.18 l=1.63
X16 B.t2 B.t0 B.t1 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=3.5802 pd=19.14 as=0 ps=0 w=9.18 l=1.63
X17 VTAIL.t11 VN.t7 VDD2.t0 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=1.5147 ps=9.51 w=9.18 l=1.63
X18 VTAIL.t6 VP.t6 VDD1.t1 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=3.5802 pd=19.14 as=1.5147 ps=9.51 w=9.18 l=1.63
X19 VTAIL.t2 VP.t7 VDD1.t0 w_n2930_n2804# sky130_fd_pr__pfet_01v8 ad=1.5147 pd=9.51 as=1.5147 ps=9.51 w=9.18 l=1.63
R0 VN.n20 VN.n19 176.548
R1 VN.n41 VN.n40 176.548
R2 VN.n4 VN.t3 169.175
R3 VN.n25 VN.t2 169.175
R4 VN.n39 VN.n21 161.3
R5 VN.n38 VN.n37 161.3
R6 VN.n36 VN.n22 161.3
R7 VN.n35 VN.n34 161.3
R8 VN.n32 VN.n23 161.3
R9 VN.n31 VN.n30 161.3
R10 VN.n29 VN.n24 161.3
R11 VN.n28 VN.n27 161.3
R12 VN.n18 VN.n0 161.3
R13 VN.n17 VN.n16 161.3
R14 VN.n15 VN.n1 161.3
R15 VN.n14 VN.n13 161.3
R16 VN.n11 VN.n2 161.3
R17 VN.n10 VN.n9 161.3
R18 VN.n8 VN.n3 161.3
R19 VN.n7 VN.n6 161.3
R20 VN.n5 VN.t4 135.73
R21 VN.n12 VN.t5 135.73
R22 VN.n19 VN.t0 135.73
R23 VN.n26 VN.t7 135.73
R24 VN.n33 VN.t1 135.73
R25 VN.n40 VN.t6 135.73
R26 VN.n10 VN.n3 56.5617
R27 VN.n17 VN.n1 56.5617
R28 VN.n31 VN.n24 56.5617
R29 VN.n38 VN.n22 56.5617
R30 VN.n5 VN.n4 55.2022
R31 VN.n26 VN.n25 55.2022
R32 VN VN.n41 44.5478
R33 VN.n6 VN.n3 24.5923
R34 VN.n11 VN.n10 24.5923
R35 VN.n13 VN.n1 24.5923
R36 VN.n18 VN.n17 24.5923
R37 VN.n27 VN.n24 24.5923
R38 VN.n34 VN.n22 24.5923
R39 VN.n32 VN.n31 24.5923
R40 VN.n39 VN.n38 24.5923
R41 VN.n28 VN.n25 17.8292
R42 VN.n7 VN.n4 17.8292
R43 VN.n13 VN.n12 13.2801
R44 VN.n34 VN.n33 13.2801
R45 VN.n6 VN.n5 11.3127
R46 VN.n12 VN.n11 11.3127
R47 VN.n27 VN.n26 11.3127
R48 VN.n33 VN.n32 11.3127
R49 VN.n19 VN.n18 9.3454
R50 VN.n40 VN.n39 9.3454
R51 VN.n41 VN.n21 0.189894
R52 VN.n37 VN.n21 0.189894
R53 VN.n37 VN.n36 0.189894
R54 VN.n36 VN.n35 0.189894
R55 VN.n35 VN.n23 0.189894
R56 VN.n30 VN.n23 0.189894
R57 VN.n30 VN.n29 0.189894
R58 VN.n29 VN.n28 0.189894
R59 VN.n8 VN.n7 0.189894
R60 VN.n9 VN.n8 0.189894
R61 VN.n9 VN.n2 0.189894
R62 VN.n14 VN.n2 0.189894
R63 VN.n15 VN.n14 0.189894
R64 VN.n16 VN.n15 0.189894
R65 VN.n16 VN.n0 0.189894
R66 VN.n20 VN.n0 0.189894
R67 VN VN.n20 0.0516364
R68 VTAIL.n14 VTAIL.t5 65.4956
R69 VTAIL.n11 VTAIL.t6 65.4956
R70 VTAIL.n10 VTAIL.t12 65.4956
R71 VTAIL.n7 VTAIL.t10 65.4956
R72 VTAIL.n15 VTAIL.t9 65.4954
R73 VTAIL.n2 VTAIL.t15 65.4954
R74 VTAIL.n3 VTAIL.t7 65.4954
R75 VTAIL.n6 VTAIL.t0 65.4954
R76 VTAIL.n13 VTAIL.n12 61.9548
R77 VTAIL.n9 VTAIL.n8 61.9548
R78 VTAIL.n1 VTAIL.n0 61.9546
R79 VTAIL.n5 VTAIL.n4 61.9546
R80 VTAIL.n15 VTAIL.n14 21.9703
R81 VTAIL.n7 VTAIL.n6 21.9703
R82 VTAIL.n0 VTAIL.t14 3.54135
R83 VTAIL.n0 VTAIL.t13 3.54135
R84 VTAIL.n4 VTAIL.t1 3.54135
R85 VTAIL.n4 VTAIL.t2 3.54135
R86 VTAIL.n12 VTAIL.t3 3.54135
R87 VTAIL.n12 VTAIL.t4 3.54135
R88 VTAIL.n8 VTAIL.t8 3.54135
R89 VTAIL.n8 VTAIL.t11 3.54135
R90 VTAIL.n9 VTAIL.n7 1.69016
R91 VTAIL.n10 VTAIL.n9 1.69016
R92 VTAIL.n13 VTAIL.n11 1.69016
R93 VTAIL.n14 VTAIL.n13 1.69016
R94 VTAIL.n6 VTAIL.n5 1.69016
R95 VTAIL.n5 VTAIL.n3 1.69016
R96 VTAIL.n2 VTAIL.n1 1.69016
R97 VTAIL VTAIL.n15 1.63197
R98 VTAIL.n11 VTAIL.n10 0.470328
R99 VTAIL.n3 VTAIL.n2 0.470328
R100 VTAIL VTAIL.n1 0.0586897
R101 VDD2.n2 VDD2.n1 79.4228
R102 VDD2.n2 VDD2.n0 79.4228
R103 VDD2 VDD2.n5 79.4202
R104 VDD2.n4 VDD2.n3 78.6336
R105 VDD2.n4 VDD2.n2 39.2325
R106 VDD2.n5 VDD2.t0 3.54135
R107 VDD2.n5 VDD2.t5 3.54135
R108 VDD2.n3 VDD2.t1 3.54135
R109 VDD2.n3 VDD2.t6 3.54135
R110 VDD2.n1 VDD2.t2 3.54135
R111 VDD2.n1 VDD2.t7 3.54135
R112 VDD2.n0 VDD2.t4 3.54135
R113 VDD2.n0 VDD2.t3 3.54135
R114 VDD2 VDD2.n4 0.903517
R115 VP.n28 VP.n27 176.548
R116 VP.n50 VP.n49 176.548
R117 VP.n26 VP.n25 176.548
R118 VP.n10 VP.t6 169.175
R119 VP.n13 VP.n12 161.3
R120 VP.n14 VP.n9 161.3
R121 VP.n16 VP.n15 161.3
R122 VP.n17 VP.n8 161.3
R123 VP.n20 VP.n19 161.3
R124 VP.n21 VP.n7 161.3
R125 VP.n23 VP.n22 161.3
R126 VP.n24 VP.n6 161.3
R127 VP.n48 VP.n0 161.3
R128 VP.n47 VP.n46 161.3
R129 VP.n45 VP.n1 161.3
R130 VP.n44 VP.n43 161.3
R131 VP.n41 VP.n2 161.3
R132 VP.n40 VP.n39 161.3
R133 VP.n38 VP.n3 161.3
R134 VP.n37 VP.n36 161.3
R135 VP.n34 VP.n4 161.3
R136 VP.n33 VP.n32 161.3
R137 VP.n31 VP.n5 161.3
R138 VP.n30 VP.n29 161.3
R139 VP.n28 VP.t2 135.73
R140 VP.n35 VP.t1 135.73
R141 VP.n42 VP.t7 135.73
R142 VP.n49 VP.t5 135.73
R143 VP.n25 VP.t0 135.73
R144 VP.n18 VP.t4 135.73
R145 VP.n11 VP.t3 135.73
R146 VP.n33 VP.n5 56.5617
R147 VP.n40 VP.n3 56.5617
R148 VP.n47 VP.n1 56.5617
R149 VP.n23 VP.n7 56.5617
R150 VP.n16 VP.n9 56.5617
R151 VP.n11 VP.n10 55.2022
R152 VP.n27 VP.n26 44.1672
R153 VP.n29 VP.n5 24.5923
R154 VP.n34 VP.n33 24.5923
R155 VP.n36 VP.n3 24.5923
R156 VP.n41 VP.n40 24.5923
R157 VP.n43 VP.n1 24.5923
R158 VP.n48 VP.n47 24.5923
R159 VP.n24 VP.n23 24.5923
R160 VP.n17 VP.n16 24.5923
R161 VP.n19 VP.n7 24.5923
R162 VP.n12 VP.n9 24.5923
R163 VP.n13 VP.n10 17.8292
R164 VP.n35 VP.n34 13.2801
R165 VP.n43 VP.n42 13.2801
R166 VP.n19 VP.n18 13.2801
R167 VP.n36 VP.n35 11.3127
R168 VP.n42 VP.n41 11.3127
R169 VP.n18 VP.n17 11.3127
R170 VP.n12 VP.n11 11.3127
R171 VP.n29 VP.n28 9.3454
R172 VP.n49 VP.n48 9.3454
R173 VP.n25 VP.n24 9.3454
R174 VP.n14 VP.n13 0.189894
R175 VP.n15 VP.n14 0.189894
R176 VP.n15 VP.n8 0.189894
R177 VP.n20 VP.n8 0.189894
R178 VP.n21 VP.n20 0.189894
R179 VP.n22 VP.n21 0.189894
R180 VP.n22 VP.n6 0.189894
R181 VP.n26 VP.n6 0.189894
R182 VP.n30 VP.n27 0.189894
R183 VP.n31 VP.n30 0.189894
R184 VP.n32 VP.n31 0.189894
R185 VP.n32 VP.n4 0.189894
R186 VP.n37 VP.n4 0.189894
R187 VP.n38 VP.n37 0.189894
R188 VP.n39 VP.n38 0.189894
R189 VP.n39 VP.n2 0.189894
R190 VP.n44 VP.n2 0.189894
R191 VP.n45 VP.n44 0.189894
R192 VP.n46 VP.n45 0.189894
R193 VP.n46 VP.n0 0.189894
R194 VP.n50 VP.n0 0.189894
R195 VP VP.n50 0.0516364
R196 VDD1 VDD1.n0 79.5366
R197 VDD1.n3 VDD1.n2 79.4228
R198 VDD1.n3 VDD1.n1 79.4228
R199 VDD1.n5 VDD1.n4 78.6336
R200 VDD1.n5 VDD1.n3 39.8155
R201 VDD1.n4 VDD1.t3 3.54135
R202 VDD1.n4 VDD1.t7 3.54135
R203 VDD1.n0 VDD1.t1 3.54135
R204 VDD1.n0 VDD1.t4 3.54135
R205 VDD1.n2 VDD1.t0 3.54135
R206 VDD1.n2 VDD1.t2 3.54135
R207 VDD1.n1 VDD1.t5 3.54135
R208 VDD1.n1 VDD1.t6 3.54135
R209 VDD1 VDD1.n5 0.787138
R210 B.n444 B.n443 585
R211 B.n445 B.n62 585
R212 B.n447 B.n446 585
R213 B.n448 B.n61 585
R214 B.n450 B.n449 585
R215 B.n451 B.n60 585
R216 B.n453 B.n452 585
R217 B.n454 B.n59 585
R218 B.n456 B.n455 585
R219 B.n457 B.n58 585
R220 B.n459 B.n458 585
R221 B.n460 B.n57 585
R222 B.n462 B.n461 585
R223 B.n463 B.n56 585
R224 B.n465 B.n464 585
R225 B.n466 B.n55 585
R226 B.n468 B.n467 585
R227 B.n469 B.n54 585
R228 B.n471 B.n470 585
R229 B.n472 B.n53 585
R230 B.n474 B.n473 585
R231 B.n475 B.n52 585
R232 B.n477 B.n476 585
R233 B.n478 B.n51 585
R234 B.n480 B.n479 585
R235 B.n481 B.n50 585
R236 B.n483 B.n482 585
R237 B.n484 B.n49 585
R238 B.n486 B.n485 585
R239 B.n487 B.n48 585
R240 B.n489 B.n488 585
R241 B.n490 B.n47 585
R242 B.n492 B.n491 585
R243 B.n494 B.n493 585
R244 B.n495 B.n43 585
R245 B.n497 B.n496 585
R246 B.n498 B.n42 585
R247 B.n500 B.n499 585
R248 B.n501 B.n41 585
R249 B.n503 B.n502 585
R250 B.n504 B.n40 585
R251 B.n506 B.n505 585
R252 B.n507 B.n37 585
R253 B.n510 B.n509 585
R254 B.n511 B.n36 585
R255 B.n513 B.n512 585
R256 B.n514 B.n35 585
R257 B.n516 B.n515 585
R258 B.n517 B.n34 585
R259 B.n519 B.n518 585
R260 B.n520 B.n33 585
R261 B.n522 B.n521 585
R262 B.n523 B.n32 585
R263 B.n525 B.n524 585
R264 B.n526 B.n31 585
R265 B.n528 B.n527 585
R266 B.n529 B.n30 585
R267 B.n531 B.n530 585
R268 B.n532 B.n29 585
R269 B.n534 B.n533 585
R270 B.n535 B.n28 585
R271 B.n537 B.n536 585
R272 B.n538 B.n27 585
R273 B.n540 B.n539 585
R274 B.n541 B.n26 585
R275 B.n543 B.n542 585
R276 B.n544 B.n25 585
R277 B.n546 B.n545 585
R278 B.n547 B.n24 585
R279 B.n549 B.n548 585
R280 B.n550 B.n23 585
R281 B.n552 B.n551 585
R282 B.n553 B.n22 585
R283 B.n555 B.n554 585
R284 B.n556 B.n21 585
R285 B.n558 B.n557 585
R286 B.n442 B.n63 585
R287 B.n441 B.n440 585
R288 B.n439 B.n64 585
R289 B.n438 B.n437 585
R290 B.n436 B.n65 585
R291 B.n435 B.n434 585
R292 B.n433 B.n66 585
R293 B.n432 B.n431 585
R294 B.n430 B.n67 585
R295 B.n429 B.n428 585
R296 B.n427 B.n68 585
R297 B.n426 B.n425 585
R298 B.n424 B.n69 585
R299 B.n423 B.n422 585
R300 B.n421 B.n70 585
R301 B.n420 B.n419 585
R302 B.n418 B.n71 585
R303 B.n417 B.n416 585
R304 B.n415 B.n72 585
R305 B.n414 B.n413 585
R306 B.n412 B.n73 585
R307 B.n411 B.n410 585
R308 B.n409 B.n74 585
R309 B.n408 B.n407 585
R310 B.n406 B.n75 585
R311 B.n405 B.n404 585
R312 B.n403 B.n76 585
R313 B.n402 B.n401 585
R314 B.n400 B.n77 585
R315 B.n399 B.n398 585
R316 B.n397 B.n78 585
R317 B.n396 B.n395 585
R318 B.n394 B.n79 585
R319 B.n393 B.n392 585
R320 B.n391 B.n80 585
R321 B.n390 B.n389 585
R322 B.n388 B.n81 585
R323 B.n387 B.n386 585
R324 B.n385 B.n82 585
R325 B.n384 B.n383 585
R326 B.n382 B.n83 585
R327 B.n381 B.n380 585
R328 B.n379 B.n84 585
R329 B.n378 B.n377 585
R330 B.n376 B.n85 585
R331 B.n375 B.n374 585
R332 B.n373 B.n86 585
R333 B.n372 B.n371 585
R334 B.n370 B.n87 585
R335 B.n369 B.n368 585
R336 B.n367 B.n88 585
R337 B.n366 B.n365 585
R338 B.n364 B.n89 585
R339 B.n363 B.n362 585
R340 B.n361 B.n90 585
R341 B.n360 B.n359 585
R342 B.n358 B.n91 585
R343 B.n357 B.n356 585
R344 B.n355 B.n92 585
R345 B.n354 B.n353 585
R346 B.n352 B.n93 585
R347 B.n351 B.n350 585
R348 B.n349 B.n94 585
R349 B.n348 B.n347 585
R350 B.n346 B.n95 585
R351 B.n345 B.n344 585
R352 B.n343 B.n96 585
R353 B.n342 B.n341 585
R354 B.n340 B.n97 585
R355 B.n339 B.n338 585
R356 B.n337 B.n98 585
R357 B.n336 B.n335 585
R358 B.n334 B.n99 585
R359 B.n333 B.n332 585
R360 B.n331 B.n100 585
R361 B.n216 B.n215 585
R362 B.n217 B.n142 585
R363 B.n219 B.n218 585
R364 B.n220 B.n141 585
R365 B.n222 B.n221 585
R366 B.n223 B.n140 585
R367 B.n225 B.n224 585
R368 B.n226 B.n139 585
R369 B.n228 B.n227 585
R370 B.n229 B.n138 585
R371 B.n231 B.n230 585
R372 B.n232 B.n137 585
R373 B.n234 B.n233 585
R374 B.n235 B.n136 585
R375 B.n237 B.n236 585
R376 B.n238 B.n135 585
R377 B.n240 B.n239 585
R378 B.n241 B.n134 585
R379 B.n243 B.n242 585
R380 B.n244 B.n133 585
R381 B.n246 B.n245 585
R382 B.n247 B.n132 585
R383 B.n249 B.n248 585
R384 B.n250 B.n131 585
R385 B.n252 B.n251 585
R386 B.n253 B.n130 585
R387 B.n255 B.n254 585
R388 B.n256 B.n129 585
R389 B.n258 B.n257 585
R390 B.n259 B.n128 585
R391 B.n261 B.n260 585
R392 B.n262 B.n127 585
R393 B.n264 B.n263 585
R394 B.n266 B.n265 585
R395 B.n267 B.n123 585
R396 B.n269 B.n268 585
R397 B.n270 B.n122 585
R398 B.n272 B.n271 585
R399 B.n273 B.n121 585
R400 B.n275 B.n274 585
R401 B.n276 B.n120 585
R402 B.n278 B.n277 585
R403 B.n279 B.n117 585
R404 B.n282 B.n281 585
R405 B.n283 B.n116 585
R406 B.n285 B.n284 585
R407 B.n286 B.n115 585
R408 B.n288 B.n287 585
R409 B.n289 B.n114 585
R410 B.n291 B.n290 585
R411 B.n292 B.n113 585
R412 B.n294 B.n293 585
R413 B.n295 B.n112 585
R414 B.n297 B.n296 585
R415 B.n298 B.n111 585
R416 B.n300 B.n299 585
R417 B.n301 B.n110 585
R418 B.n303 B.n302 585
R419 B.n304 B.n109 585
R420 B.n306 B.n305 585
R421 B.n307 B.n108 585
R422 B.n309 B.n308 585
R423 B.n310 B.n107 585
R424 B.n312 B.n311 585
R425 B.n313 B.n106 585
R426 B.n315 B.n314 585
R427 B.n316 B.n105 585
R428 B.n318 B.n317 585
R429 B.n319 B.n104 585
R430 B.n321 B.n320 585
R431 B.n322 B.n103 585
R432 B.n324 B.n323 585
R433 B.n325 B.n102 585
R434 B.n327 B.n326 585
R435 B.n328 B.n101 585
R436 B.n330 B.n329 585
R437 B.n214 B.n143 585
R438 B.n213 B.n212 585
R439 B.n211 B.n144 585
R440 B.n210 B.n209 585
R441 B.n208 B.n145 585
R442 B.n207 B.n206 585
R443 B.n205 B.n146 585
R444 B.n204 B.n203 585
R445 B.n202 B.n147 585
R446 B.n201 B.n200 585
R447 B.n199 B.n148 585
R448 B.n198 B.n197 585
R449 B.n196 B.n149 585
R450 B.n195 B.n194 585
R451 B.n193 B.n150 585
R452 B.n192 B.n191 585
R453 B.n190 B.n151 585
R454 B.n189 B.n188 585
R455 B.n187 B.n152 585
R456 B.n186 B.n185 585
R457 B.n184 B.n153 585
R458 B.n183 B.n182 585
R459 B.n181 B.n154 585
R460 B.n180 B.n179 585
R461 B.n178 B.n155 585
R462 B.n177 B.n176 585
R463 B.n175 B.n156 585
R464 B.n174 B.n173 585
R465 B.n172 B.n157 585
R466 B.n171 B.n170 585
R467 B.n169 B.n158 585
R468 B.n168 B.n167 585
R469 B.n166 B.n159 585
R470 B.n165 B.n164 585
R471 B.n163 B.n160 585
R472 B.n162 B.n161 585
R473 B.n2 B.n0 585
R474 B.n613 B.n1 585
R475 B.n612 B.n611 585
R476 B.n610 B.n3 585
R477 B.n609 B.n608 585
R478 B.n607 B.n4 585
R479 B.n606 B.n605 585
R480 B.n604 B.n5 585
R481 B.n603 B.n602 585
R482 B.n601 B.n6 585
R483 B.n600 B.n599 585
R484 B.n598 B.n7 585
R485 B.n597 B.n596 585
R486 B.n595 B.n8 585
R487 B.n594 B.n593 585
R488 B.n592 B.n9 585
R489 B.n591 B.n590 585
R490 B.n589 B.n10 585
R491 B.n588 B.n587 585
R492 B.n586 B.n11 585
R493 B.n585 B.n584 585
R494 B.n583 B.n12 585
R495 B.n582 B.n581 585
R496 B.n580 B.n13 585
R497 B.n579 B.n578 585
R498 B.n577 B.n14 585
R499 B.n576 B.n575 585
R500 B.n574 B.n15 585
R501 B.n573 B.n572 585
R502 B.n571 B.n16 585
R503 B.n570 B.n569 585
R504 B.n568 B.n17 585
R505 B.n567 B.n566 585
R506 B.n565 B.n18 585
R507 B.n564 B.n563 585
R508 B.n562 B.n19 585
R509 B.n561 B.n560 585
R510 B.n559 B.n20 585
R511 B.n615 B.n614 585
R512 B.n216 B.n143 506.916
R513 B.n559 B.n558 506.916
R514 B.n331 B.n330 506.916
R515 B.n444 B.n63 506.916
R516 B.n118 B.t6 341.623
R517 B.n124 B.t3 341.623
R518 B.n38 B.t0 341.623
R519 B.n44 B.t9 341.623
R520 B.n212 B.n143 163.367
R521 B.n212 B.n211 163.367
R522 B.n211 B.n210 163.367
R523 B.n210 B.n145 163.367
R524 B.n206 B.n145 163.367
R525 B.n206 B.n205 163.367
R526 B.n205 B.n204 163.367
R527 B.n204 B.n147 163.367
R528 B.n200 B.n147 163.367
R529 B.n200 B.n199 163.367
R530 B.n199 B.n198 163.367
R531 B.n198 B.n149 163.367
R532 B.n194 B.n149 163.367
R533 B.n194 B.n193 163.367
R534 B.n193 B.n192 163.367
R535 B.n192 B.n151 163.367
R536 B.n188 B.n151 163.367
R537 B.n188 B.n187 163.367
R538 B.n187 B.n186 163.367
R539 B.n186 B.n153 163.367
R540 B.n182 B.n153 163.367
R541 B.n182 B.n181 163.367
R542 B.n181 B.n180 163.367
R543 B.n180 B.n155 163.367
R544 B.n176 B.n155 163.367
R545 B.n176 B.n175 163.367
R546 B.n175 B.n174 163.367
R547 B.n174 B.n157 163.367
R548 B.n170 B.n157 163.367
R549 B.n170 B.n169 163.367
R550 B.n169 B.n168 163.367
R551 B.n168 B.n159 163.367
R552 B.n164 B.n159 163.367
R553 B.n164 B.n163 163.367
R554 B.n163 B.n162 163.367
R555 B.n162 B.n2 163.367
R556 B.n614 B.n2 163.367
R557 B.n614 B.n613 163.367
R558 B.n613 B.n612 163.367
R559 B.n612 B.n3 163.367
R560 B.n608 B.n3 163.367
R561 B.n608 B.n607 163.367
R562 B.n607 B.n606 163.367
R563 B.n606 B.n5 163.367
R564 B.n602 B.n5 163.367
R565 B.n602 B.n601 163.367
R566 B.n601 B.n600 163.367
R567 B.n600 B.n7 163.367
R568 B.n596 B.n7 163.367
R569 B.n596 B.n595 163.367
R570 B.n595 B.n594 163.367
R571 B.n594 B.n9 163.367
R572 B.n590 B.n9 163.367
R573 B.n590 B.n589 163.367
R574 B.n589 B.n588 163.367
R575 B.n588 B.n11 163.367
R576 B.n584 B.n11 163.367
R577 B.n584 B.n583 163.367
R578 B.n583 B.n582 163.367
R579 B.n582 B.n13 163.367
R580 B.n578 B.n13 163.367
R581 B.n578 B.n577 163.367
R582 B.n577 B.n576 163.367
R583 B.n576 B.n15 163.367
R584 B.n572 B.n15 163.367
R585 B.n572 B.n571 163.367
R586 B.n571 B.n570 163.367
R587 B.n570 B.n17 163.367
R588 B.n566 B.n17 163.367
R589 B.n566 B.n565 163.367
R590 B.n565 B.n564 163.367
R591 B.n564 B.n19 163.367
R592 B.n560 B.n19 163.367
R593 B.n560 B.n559 163.367
R594 B.n217 B.n216 163.367
R595 B.n218 B.n217 163.367
R596 B.n218 B.n141 163.367
R597 B.n222 B.n141 163.367
R598 B.n223 B.n222 163.367
R599 B.n224 B.n223 163.367
R600 B.n224 B.n139 163.367
R601 B.n228 B.n139 163.367
R602 B.n229 B.n228 163.367
R603 B.n230 B.n229 163.367
R604 B.n230 B.n137 163.367
R605 B.n234 B.n137 163.367
R606 B.n235 B.n234 163.367
R607 B.n236 B.n235 163.367
R608 B.n236 B.n135 163.367
R609 B.n240 B.n135 163.367
R610 B.n241 B.n240 163.367
R611 B.n242 B.n241 163.367
R612 B.n242 B.n133 163.367
R613 B.n246 B.n133 163.367
R614 B.n247 B.n246 163.367
R615 B.n248 B.n247 163.367
R616 B.n248 B.n131 163.367
R617 B.n252 B.n131 163.367
R618 B.n253 B.n252 163.367
R619 B.n254 B.n253 163.367
R620 B.n254 B.n129 163.367
R621 B.n258 B.n129 163.367
R622 B.n259 B.n258 163.367
R623 B.n260 B.n259 163.367
R624 B.n260 B.n127 163.367
R625 B.n264 B.n127 163.367
R626 B.n265 B.n264 163.367
R627 B.n265 B.n123 163.367
R628 B.n269 B.n123 163.367
R629 B.n270 B.n269 163.367
R630 B.n271 B.n270 163.367
R631 B.n271 B.n121 163.367
R632 B.n275 B.n121 163.367
R633 B.n276 B.n275 163.367
R634 B.n277 B.n276 163.367
R635 B.n277 B.n117 163.367
R636 B.n282 B.n117 163.367
R637 B.n283 B.n282 163.367
R638 B.n284 B.n283 163.367
R639 B.n284 B.n115 163.367
R640 B.n288 B.n115 163.367
R641 B.n289 B.n288 163.367
R642 B.n290 B.n289 163.367
R643 B.n290 B.n113 163.367
R644 B.n294 B.n113 163.367
R645 B.n295 B.n294 163.367
R646 B.n296 B.n295 163.367
R647 B.n296 B.n111 163.367
R648 B.n300 B.n111 163.367
R649 B.n301 B.n300 163.367
R650 B.n302 B.n301 163.367
R651 B.n302 B.n109 163.367
R652 B.n306 B.n109 163.367
R653 B.n307 B.n306 163.367
R654 B.n308 B.n307 163.367
R655 B.n308 B.n107 163.367
R656 B.n312 B.n107 163.367
R657 B.n313 B.n312 163.367
R658 B.n314 B.n313 163.367
R659 B.n314 B.n105 163.367
R660 B.n318 B.n105 163.367
R661 B.n319 B.n318 163.367
R662 B.n320 B.n319 163.367
R663 B.n320 B.n103 163.367
R664 B.n324 B.n103 163.367
R665 B.n325 B.n324 163.367
R666 B.n326 B.n325 163.367
R667 B.n326 B.n101 163.367
R668 B.n330 B.n101 163.367
R669 B.n332 B.n331 163.367
R670 B.n332 B.n99 163.367
R671 B.n336 B.n99 163.367
R672 B.n337 B.n336 163.367
R673 B.n338 B.n337 163.367
R674 B.n338 B.n97 163.367
R675 B.n342 B.n97 163.367
R676 B.n343 B.n342 163.367
R677 B.n344 B.n343 163.367
R678 B.n344 B.n95 163.367
R679 B.n348 B.n95 163.367
R680 B.n349 B.n348 163.367
R681 B.n350 B.n349 163.367
R682 B.n350 B.n93 163.367
R683 B.n354 B.n93 163.367
R684 B.n355 B.n354 163.367
R685 B.n356 B.n355 163.367
R686 B.n356 B.n91 163.367
R687 B.n360 B.n91 163.367
R688 B.n361 B.n360 163.367
R689 B.n362 B.n361 163.367
R690 B.n362 B.n89 163.367
R691 B.n366 B.n89 163.367
R692 B.n367 B.n366 163.367
R693 B.n368 B.n367 163.367
R694 B.n368 B.n87 163.367
R695 B.n372 B.n87 163.367
R696 B.n373 B.n372 163.367
R697 B.n374 B.n373 163.367
R698 B.n374 B.n85 163.367
R699 B.n378 B.n85 163.367
R700 B.n379 B.n378 163.367
R701 B.n380 B.n379 163.367
R702 B.n380 B.n83 163.367
R703 B.n384 B.n83 163.367
R704 B.n385 B.n384 163.367
R705 B.n386 B.n385 163.367
R706 B.n386 B.n81 163.367
R707 B.n390 B.n81 163.367
R708 B.n391 B.n390 163.367
R709 B.n392 B.n391 163.367
R710 B.n392 B.n79 163.367
R711 B.n396 B.n79 163.367
R712 B.n397 B.n396 163.367
R713 B.n398 B.n397 163.367
R714 B.n398 B.n77 163.367
R715 B.n402 B.n77 163.367
R716 B.n403 B.n402 163.367
R717 B.n404 B.n403 163.367
R718 B.n404 B.n75 163.367
R719 B.n408 B.n75 163.367
R720 B.n409 B.n408 163.367
R721 B.n410 B.n409 163.367
R722 B.n410 B.n73 163.367
R723 B.n414 B.n73 163.367
R724 B.n415 B.n414 163.367
R725 B.n416 B.n415 163.367
R726 B.n416 B.n71 163.367
R727 B.n420 B.n71 163.367
R728 B.n421 B.n420 163.367
R729 B.n422 B.n421 163.367
R730 B.n422 B.n69 163.367
R731 B.n426 B.n69 163.367
R732 B.n427 B.n426 163.367
R733 B.n428 B.n427 163.367
R734 B.n428 B.n67 163.367
R735 B.n432 B.n67 163.367
R736 B.n433 B.n432 163.367
R737 B.n434 B.n433 163.367
R738 B.n434 B.n65 163.367
R739 B.n438 B.n65 163.367
R740 B.n439 B.n438 163.367
R741 B.n440 B.n439 163.367
R742 B.n440 B.n63 163.367
R743 B.n558 B.n21 163.367
R744 B.n554 B.n21 163.367
R745 B.n554 B.n553 163.367
R746 B.n553 B.n552 163.367
R747 B.n552 B.n23 163.367
R748 B.n548 B.n23 163.367
R749 B.n548 B.n547 163.367
R750 B.n547 B.n546 163.367
R751 B.n546 B.n25 163.367
R752 B.n542 B.n25 163.367
R753 B.n542 B.n541 163.367
R754 B.n541 B.n540 163.367
R755 B.n540 B.n27 163.367
R756 B.n536 B.n27 163.367
R757 B.n536 B.n535 163.367
R758 B.n535 B.n534 163.367
R759 B.n534 B.n29 163.367
R760 B.n530 B.n29 163.367
R761 B.n530 B.n529 163.367
R762 B.n529 B.n528 163.367
R763 B.n528 B.n31 163.367
R764 B.n524 B.n31 163.367
R765 B.n524 B.n523 163.367
R766 B.n523 B.n522 163.367
R767 B.n522 B.n33 163.367
R768 B.n518 B.n33 163.367
R769 B.n518 B.n517 163.367
R770 B.n517 B.n516 163.367
R771 B.n516 B.n35 163.367
R772 B.n512 B.n35 163.367
R773 B.n512 B.n511 163.367
R774 B.n511 B.n510 163.367
R775 B.n510 B.n37 163.367
R776 B.n505 B.n37 163.367
R777 B.n505 B.n504 163.367
R778 B.n504 B.n503 163.367
R779 B.n503 B.n41 163.367
R780 B.n499 B.n41 163.367
R781 B.n499 B.n498 163.367
R782 B.n498 B.n497 163.367
R783 B.n497 B.n43 163.367
R784 B.n493 B.n43 163.367
R785 B.n493 B.n492 163.367
R786 B.n492 B.n47 163.367
R787 B.n488 B.n47 163.367
R788 B.n488 B.n487 163.367
R789 B.n487 B.n486 163.367
R790 B.n486 B.n49 163.367
R791 B.n482 B.n49 163.367
R792 B.n482 B.n481 163.367
R793 B.n481 B.n480 163.367
R794 B.n480 B.n51 163.367
R795 B.n476 B.n51 163.367
R796 B.n476 B.n475 163.367
R797 B.n475 B.n474 163.367
R798 B.n474 B.n53 163.367
R799 B.n470 B.n53 163.367
R800 B.n470 B.n469 163.367
R801 B.n469 B.n468 163.367
R802 B.n468 B.n55 163.367
R803 B.n464 B.n55 163.367
R804 B.n464 B.n463 163.367
R805 B.n463 B.n462 163.367
R806 B.n462 B.n57 163.367
R807 B.n458 B.n57 163.367
R808 B.n458 B.n457 163.367
R809 B.n457 B.n456 163.367
R810 B.n456 B.n59 163.367
R811 B.n452 B.n59 163.367
R812 B.n452 B.n451 163.367
R813 B.n451 B.n450 163.367
R814 B.n450 B.n61 163.367
R815 B.n446 B.n61 163.367
R816 B.n446 B.n445 163.367
R817 B.n445 B.n444 163.367
R818 B.n118 B.t8 152.63
R819 B.n44 B.t10 152.63
R820 B.n124 B.t5 152.619
R821 B.n38 B.t1 152.619
R822 B.n119 B.t7 114.618
R823 B.n45 B.t11 114.618
R824 B.n125 B.t4 114.608
R825 B.n39 B.t2 114.608
R826 B.n280 B.n119 59.5399
R827 B.n126 B.n125 59.5399
R828 B.n508 B.n39 59.5399
R829 B.n46 B.n45 59.5399
R830 B.n119 B.n118 38.0126
R831 B.n125 B.n124 38.0126
R832 B.n39 B.n38 38.0126
R833 B.n45 B.n44 38.0126
R834 B.n557 B.n20 32.9371
R835 B.n443 B.n442 32.9371
R836 B.n329 B.n100 32.9371
R837 B.n215 B.n214 32.9371
R838 B B.n615 18.0485
R839 B.n557 B.n556 10.6151
R840 B.n556 B.n555 10.6151
R841 B.n555 B.n22 10.6151
R842 B.n551 B.n22 10.6151
R843 B.n551 B.n550 10.6151
R844 B.n550 B.n549 10.6151
R845 B.n549 B.n24 10.6151
R846 B.n545 B.n24 10.6151
R847 B.n545 B.n544 10.6151
R848 B.n544 B.n543 10.6151
R849 B.n543 B.n26 10.6151
R850 B.n539 B.n26 10.6151
R851 B.n539 B.n538 10.6151
R852 B.n538 B.n537 10.6151
R853 B.n537 B.n28 10.6151
R854 B.n533 B.n28 10.6151
R855 B.n533 B.n532 10.6151
R856 B.n532 B.n531 10.6151
R857 B.n531 B.n30 10.6151
R858 B.n527 B.n30 10.6151
R859 B.n527 B.n526 10.6151
R860 B.n526 B.n525 10.6151
R861 B.n525 B.n32 10.6151
R862 B.n521 B.n32 10.6151
R863 B.n521 B.n520 10.6151
R864 B.n520 B.n519 10.6151
R865 B.n519 B.n34 10.6151
R866 B.n515 B.n34 10.6151
R867 B.n515 B.n514 10.6151
R868 B.n514 B.n513 10.6151
R869 B.n513 B.n36 10.6151
R870 B.n509 B.n36 10.6151
R871 B.n507 B.n506 10.6151
R872 B.n506 B.n40 10.6151
R873 B.n502 B.n40 10.6151
R874 B.n502 B.n501 10.6151
R875 B.n501 B.n500 10.6151
R876 B.n500 B.n42 10.6151
R877 B.n496 B.n42 10.6151
R878 B.n496 B.n495 10.6151
R879 B.n495 B.n494 10.6151
R880 B.n491 B.n490 10.6151
R881 B.n490 B.n489 10.6151
R882 B.n489 B.n48 10.6151
R883 B.n485 B.n48 10.6151
R884 B.n485 B.n484 10.6151
R885 B.n484 B.n483 10.6151
R886 B.n483 B.n50 10.6151
R887 B.n479 B.n50 10.6151
R888 B.n479 B.n478 10.6151
R889 B.n478 B.n477 10.6151
R890 B.n477 B.n52 10.6151
R891 B.n473 B.n52 10.6151
R892 B.n473 B.n472 10.6151
R893 B.n472 B.n471 10.6151
R894 B.n471 B.n54 10.6151
R895 B.n467 B.n54 10.6151
R896 B.n467 B.n466 10.6151
R897 B.n466 B.n465 10.6151
R898 B.n465 B.n56 10.6151
R899 B.n461 B.n56 10.6151
R900 B.n461 B.n460 10.6151
R901 B.n460 B.n459 10.6151
R902 B.n459 B.n58 10.6151
R903 B.n455 B.n58 10.6151
R904 B.n455 B.n454 10.6151
R905 B.n454 B.n453 10.6151
R906 B.n453 B.n60 10.6151
R907 B.n449 B.n60 10.6151
R908 B.n449 B.n448 10.6151
R909 B.n448 B.n447 10.6151
R910 B.n447 B.n62 10.6151
R911 B.n443 B.n62 10.6151
R912 B.n333 B.n100 10.6151
R913 B.n334 B.n333 10.6151
R914 B.n335 B.n334 10.6151
R915 B.n335 B.n98 10.6151
R916 B.n339 B.n98 10.6151
R917 B.n340 B.n339 10.6151
R918 B.n341 B.n340 10.6151
R919 B.n341 B.n96 10.6151
R920 B.n345 B.n96 10.6151
R921 B.n346 B.n345 10.6151
R922 B.n347 B.n346 10.6151
R923 B.n347 B.n94 10.6151
R924 B.n351 B.n94 10.6151
R925 B.n352 B.n351 10.6151
R926 B.n353 B.n352 10.6151
R927 B.n353 B.n92 10.6151
R928 B.n357 B.n92 10.6151
R929 B.n358 B.n357 10.6151
R930 B.n359 B.n358 10.6151
R931 B.n359 B.n90 10.6151
R932 B.n363 B.n90 10.6151
R933 B.n364 B.n363 10.6151
R934 B.n365 B.n364 10.6151
R935 B.n365 B.n88 10.6151
R936 B.n369 B.n88 10.6151
R937 B.n370 B.n369 10.6151
R938 B.n371 B.n370 10.6151
R939 B.n371 B.n86 10.6151
R940 B.n375 B.n86 10.6151
R941 B.n376 B.n375 10.6151
R942 B.n377 B.n376 10.6151
R943 B.n377 B.n84 10.6151
R944 B.n381 B.n84 10.6151
R945 B.n382 B.n381 10.6151
R946 B.n383 B.n382 10.6151
R947 B.n383 B.n82 10.6151
R948 B.n387 B.n82 10.6151
R949 B.n388 B.n387 10.6151
R950 B.n389 B.n388 10.6151
R951 B.n389 B.n80 10.6151
R952 B.n393 B.n80 10.6151
R953 B.n394 B.n393 10.6151
R954 B.n395 B.n394 10.6151
R955 B.n395 B.n78 10.6151
R956 B.n399 B.n78 10.6151
R957 B.n400 B.n399 10.6151
R958 B.n401 B.n400 10.6151
R959 B.n401 B.n76 10.6151
R960 B.n405 B.n76 10.6151
R961 B.n406 B.n405 10.6151
R962 B.n407 B.n406 10.6151
R963 B.n407 B.n74 10.6151
R964 B.n411 B.n74 10.6151
R965 B.n412 B.n411 10.6151
R966 B.n413 B.n412 10.6151
R967 B.n413 B.n72 10.6151
R968 B.n417 B.n72 10.6151
R969 B.n418 B.n417 10.6151
R970 B.n419 B.n418 10.6151
R971 B.n419 B.n70 10.6151
R972 B.n423 B.n70 10.6151
R973 B.n424 B.n423 10.6151
R974 B.n425 B.n424 10.6151
R975 B.n425 B.n68 10.6151
R976 B.n429 B.n68 10.6151
R977 B.n430 B.n429 10.6151
R978 B.n431 B.n430 10.6151
R979 B.n431 B.n66 10.6151
R980 B.n435 B.n66 10.6151
R981 B.n436 B.n435 10.6151
R982 B.n437 B.n436 10.6151
R983 B.n437 B.n64 10.6151
R984 B.n441 B.n64 10.6151
R985 B.n442 B.n441 10.6151
R986 B.n215 B.n142 10.6151
R987 B.n219 B.n142 10.6151
R988 B.n220 B.n219 10.6151
R989 B.n221 B.n220 10.6151
R990 B.n221 B.n140 10.6151
R991 B.n225 B.n140 10.6151
R992 B.n226 B.n225 10.6151
R993 B.n227 B.n226 10.6151
R994 B.n227 B.n138 10.6151
R995 B.n231 B.n138 10.6151
R996 B.n232 B.n231 10.6151
R997 B.n233 B.n232 10.6151
R998 B.n233 B.n136 10.6151
R999 B.n237 B.n136 10.6151
R1000 B.n238 B.n237 10.6151
R1001 B.n239 B.n238 10.6151
R1002 B.n239 B.n134 10.6151
R1003 B.n243 B.n134 10.6151
R1004 B.n244 B.n243 10.6151
R1005 B.n245 B.n244 10.6151
R1006 B.n245 B.n132 10.6151
R1007 B.n249 B.n132 10.6151
R1008 B.n250 B.n249 10.6151
R1009 B.n251 B.n250 10.6151
R1010 B.n251 B.n130 10.6151
R1011 B.n255 B.n130 10.6151
R1012 B.n256 B.n255 10.6151
R1013 B.n257 B.n256 10.6151
R1014 B.n257 B.n128 10.6151
R1015 B.n261 B.n128 10.6151
R1016 B.n262 B.n261 10.6151
R1017 B.n263 B.n262 10.6151
R1018 B.n267 B.n266 10.6151
R1019 B.n268 B.n267 10.6151
R1020 B.n268 B.n122 10.6151
R1021 B.n272 B.n122 10.6151
R1022 B.n273 B.n272 10.6151
R1023 B.n274 B.n273 10.6151
R1024 B.n274 B.n120 10.6151
R1025 B.n278 B.n120 10.6151
R1026 B.n279 B.n278 10.6151
R1027 B.n281 B.n116 10.6151
R1028 B.n285 B.n116 10.6151
R1029 B.n286 B.n285 10.6151
R1030 B.n287 B.n286 10.6151
R1031 B.n287 B.n114 10.6151
R1032 B.n291 B.n114 10.6151
R1033 B.n292 B.n291 10.6151
R1034 B.n293 B.n292 10.6151
R1035 B.n293 B.n112 10.6151
R1036 B.n297 B.n112 10.6151
R1037 B.n298 B.n297 10.6151
R1038 B.n299 B.n298 10.6151
R1039 B.n299 B.n110 10.6151
R1040 B.n303 B.n110 10.6151
R1041 B.n304 B.n303 10.6151
R1042 B.n305 B.n304 10.6151
R1043 B.n305 B.n108 10.6151
R1044 B.n309 B.n108 10.6151
R1045 B.n310 B.n309 10.6151
R1046 B.n311 B.n310 10.6151
R1047 B.n311 B.n106 10.6151
R1048 B.n315 B.n106 10.6151
R1049 B.n316 B.n315 10.6151
R1050 B.n317 B.n316 10.6151
R1051 B.n317 B.n104 10.6151
R1052 B.n321 B.n104 10.6151
R1053 B.n322 B.n321 10.6151
R1054 B.n323 B.n322 10.6151
R1055 B.n323 B.n102 10.6151
R1056 B.n327 B.n102 10.6151
R1057 B.n328 B.n327 10.6151
R1058 B.n329 B.n328 10.6151
R1059 B.n214 B.n213 10.6151
R1060 B.n213 B.n144 10.6151
R1061 B.n209 B.n144 10.6151
R1062 B.n209 B.n208 10.6151
R1063 B.n208 B.n207 10.6151
R1064 B.n207 B.n146 10.6151
R1065 B.n203 B.n146 10.6151
R1066 B.n203 B.n202 10.6151
R1067 B.n202 B.n201 10.6151
R1068 B.n201 B.n148 10.6151
R1069 B.n197 B.n148 10.6151
R1070 B.n197 B.n196 10.6151
R1071 B.n196 B.n195 10.6151
R1072 B.n195 B.n150 10.6151
R1073 B.n191 B.n150 10.6151
R1074 B.n191 B.n190 10.6151
R1075 B.n190 B.n189 10.6151
R1076 B.n189 B.n152 10.6151
R1077 B.n185 B.n152 10.6151
R1078 B.n185 B.n184 10.6151
R1079 B.n184 B.n183 10.6151
R1080 B.n183 B.n154 10.6151
R1081 B.n179 B.n154 10.6151
R1082 B.n179 B.n178 10.6151
R1083 B.n178 B.n177 10.6151
R1084 B.n177 B.n156 10.6151
R1085 B.n173 B.n156 10.6151
R1086 B.n173 B.n172 10.6151
R1087 B.n172 B.n171 10.6151
R1088 B.n171 B.n158 10.6151
R1089 B.n167 B.n158 10.6151
R1090 B.n167 B.n166 10.6151
R1091 B.n166 B.n165 10.6151
R1092 B.n165 B.n160 10.6151
R1093 B.n161 B.n160 10.6151
R1094 B.n161 B.n0 10.6151
R1095 B.n611 B.n1 10.6151
R1096 B.n611 B.n610 10.6151
R1097 B.n610 B.n609 10.6151
R1098 B.n609 B.n4 10.6151
R1099 B.n605 B.n4 10.6151
R1100 B.n605 B.n604 10.6151
R1101 B.n604 B.n603 10.6151
R1102 B.n603 B.n6 10.6151
R1103 B.n599 B.n6 10.6151
R1104 B.n599 B.n598 10.6151
R1105 B.n598 B.n597 10.6151
R1106 B.n597 B.n8 10.6151
R1107 B.n593 B.n8 10.6151
R1108 B.n593 B.n592 10.6151
R1109 B.n592 B.n591 10.6151
R1110 B.n591 B.n10 10.6151
R1111 B.n587 B.n10 10.6151
R1112 B.n587 B.n586 10.6151
R1113 B.n586 B.n585 10.6151
R1114 B.n585 B.n12 10.6151
R1115 B.n581 B.n12 10.6151
R1116 B.n581 B.n580 10.6151
R1117 B.n580 B.n579 10.6151
R1118 B.n579 B.n14 10.6151
R1119 B.n575 B.n14 10.6151
R1120 B.n575 B.n574 10.6151
R1121 B.n574 B.n573 10.6151
R1122 B.n573 B.n16 10.6151
R1123 B.n569 B.n16 10.6151
R1124 B.n569 B.n568 10.6151
R1125 B.n568 B.n567 10.6151
R1126 B.n567 B.n18 10.6151
R1127 B.n563 B.n18 10.6151
R1128 B.n563 B.n562 10.6151
R1129 B.n562 B.n561 10.6151
R1130 B.n561 B.n20 10.6151
R1131 B.n509 B.n508 9.36635
R1132 B.n491 B.n46 9.36635
R1133 B.n263 B.n126 9.36635
R1134 B.n281 B.n280 9.36635
R1135 B.n615 B.n0 2.81026
R1136 B.n615 B.n1 2.81026
R1137 B.n508 B.n507 1.24928
R1138 B.n494 B.n46 1.24928
R1139 B.n266 B.n126 1.24928
R1140 B.n280 B.n279 1.24928
C0 B VP 1.59696f
C1 VTAIL w_n2930_n2804# 3.50386f
C2 VDD2 w_n2930_n2804# 1.63643f
C3 VDD2 VTAIL 7.13657f
C4 B VDD1 1.27826f
C5 B VN 0.969288f
C6 VP VDD1 6.29481f
C7 VN VP 5.9477f
C8 B w_n2930_n2804# 7.83924f
C9 B VTAIL 3.62198f
C10 VN VDD1 0.15038f
C11 B VDD2 1.34377f
C12 VP w_n2930_n2804# 6.00101f
C13 VP VTAIL 6.24134f
C14 VP VDD2 0.416858f
C15 VDD1 w_n2930_n2804# 1.56241f
C16 VTAIL VDD1 7.08866f
C17 VN w_n2930_n2804# 5.62349f
C18 VN VTAIL 6.22723f
C19 VDD2 VDD1 1.27335f
C20 VN VDD2 6.02923f
C21 VDD2 VSUBS 1.466897f
C22 VDD1 VSUBS 1.947391f
C23 VTAIL VSUBS 1.010379f
C24 VN VSUBS 5.39767f
C25 VP VSUBS 2.479597f
C26 B VSUBS 3.681748f
C27 w_n2930_n2804# VSUBS 0.101648p
C28 B.n0 VSUBS 0.004875f
C29 B.n1 VSUBS 0.004875f
C30 B.n2 VSUBS 0.00771f
C31 B.n3 VSUBS 0.00771f
C32 B.n4 VSUBS 0.00771f
C33 B.n5 VSUBS 0.00771f
C34 B.n6 VSUBS 0.00771f
C35 B.n7 VSUBS 0.00771f
C36 B.n8 VSUBS 0.00771f
C37 B.n9 VSUBS 0.00771f
C38 B.n10 VSUBS 0.00771f
C39 B.n11 VSUBS 0.00771f
C40 B.n12 VSUBS 0.00771f
C41 B.n13 VSUBS 0.00771f
C42 B.n14 VSUBS 0.00771f
C43 B.n15 VSUBS 0.00771f
C44 B.n16 VSUBS 0.00771f
C45 B.n17 VSUBS 0.00771f
C46 B.n18 VSUBS 0.00771f
C47 B.n19 VSUBS 0.00771f
C48 B.n20 VSUBS 0.017843f
C49 B.n21 VSUBS 0.00771f
C50 B.n22 VSUBS 0.00771f
C51 B.n23 VSUBS 0.00771f
C52 B.n24 VSUBS 0.00771f
C53 B.n25 VSUBS 0.00771f
C54 B.n26 VSUBS 0.00771f
C55 B.n27 VSUBS 0.00771f
C56 B.n28 VSUBS 0.00771f
C57 B.n29 VSUBS 0.00771f
C58 B.n30 VSUBS 0.00771f
C59 B.n31 VSUBS 0.00771f
C60 B.n32 VSUBS 0.00771f
C61 B.n33 VSUBS 0.00771f
C62 B.n34 VSUBS 0.00771f
C63 B.n35 VSUBS 0.00771f
C64 B.n36 VSUBS 0.00771f
C65 B.n37 VSUBS 0.00771f
C66 B.t2 VSUBS 0.318629f
C67 B.t1 VSUBS 0.334431f
C68 B.t0 VSUBS 0.738882f
C69 B.n38 VSUBS 0.16025f
C70 B.n39 VSUBS 0.074441f
C71 B.n40 VSUBS 0.00771f
C72 B.n41 VSUBS 0.00771f
C73 B.n42 VSUBS 0.00771f
C74 B.n43 VSUBS 0.00771f
C75 B.t11 VSUBS 0.318626f
C76 B.t10 VSUBS 0.334428f
C77 B.t9 VSUBS 0.738882f
C78 B.n44 VSUBS 0.160253f
C79 B.n45 VSUBS 0.074445f
C80 B.n46 VSUBS 0.017863f
C81 B.n47 VSUBS 0.00771f
C82 B.n48 VSUBS 0.00771f
C83 B.n49 VSUBS 0.00771f
C84 B.n50 VSUBS 0.00771f
C85 B.n51 VSUBS 0.00771f
C86 B.n52 VSUBS 0.00771f
C87 B.n53 VSUBS 0.00771f
C88 B.n54 VSUBS 0.00771f
C89 B.n55 VSUBS 0.00771f
C90 B.n56 VSUBS 0.00771f
C91 B.n57 VSUBS 0.00771f
C92 B.n58 VSUBS 0.00771f
C93 B.n59 VSUBS 0.00771f
C94 B.n60 VSUBS 0.00771f
C95 B.n61 VSUBS 0.00771f
C96 B.n62 VSUBS 0.00771f
C97 B.n63 VSUBS 0.017843f
C98 B.n64 VSUBS 0.00771f
C99 B.n65 VSUBS 0.00771f
C100 B.n66 VSUBS 0.00771f
C101 B.n67 VSUBS 0.00771f
C102 B.n68 VSUBS 0.00771f
C103 B.n69 VSUBS 0.00771f
C104 B.n70 VSUBS 0.00771f
C105 B.n71 VSUBS 0.00771f
C106 B.n72 VSUBS 0.00771f
C107 B.n73 VSUBS 0.00771f
C108 B.n74 VSUBS 0.00771f
C109 B.n75 VSUBS 0.00771f
C110 B.n76 VSUBS 0.00771f
C111 B.n77 VSUBS 0.00771f
C112 B.n78 VSUBS 0.00771f
C113 B.n79 VSUBS 0.00771f
C114 B.n80 VSUBS 0.00771f
C115 B.n81 VSUBS 0.00771f
C116 B.n82 VSUBS 0.00771f
C117 B.n83 VSUBS 0.00771f
C118 B.n84 VSUBS 0.00771f
C119 B.n85 VSUBS 0.00771f
C120 B.n86 VSUBS 0.00771f
C121 B.n87 VSUBS 0.00771f
C122 B.n88 VSUBS 0.00771f
C123 B.n89 VSUBS 0.00771f
C124 B.n90 VSUBS 0.00771f
C125 B.n91 VSUBS 0.00771f
C126 B.n92 VSUBS 0.00771f
C127 B.n93 VSUBS 0.00771f
C128 B.n94 VSUBS 0.00771f
C129 B.n95 VSUBS 0.00771f
C130 B.n96 VSUBS 0.00771f
C131 B.n97 VSUBS 0.00771f
C132 B.n98 VSUBS 0.00771f
C133 B.n99 VSUBS 0.00771f
C134 B.n100 VSUBS 0.017843f
C135 B.n101 VSUBS 0.00771f
C136 B.n102 VSUBS 0.00771f
C137 B.n103 VSUBS 0.00771f
C138 B.n104 VSUBS 0.00771f
C139 B.n105 VSUBS 0.00771f
C140 B.n106 VSUBS 0.00771f
C141 B.n107 VSUBS 0.00771f
C142 B.n108 VSUBS 0.00771f
C143 B.n109 VSUBS 0.00771f
C144 B.n110 VSUBS 0.00771f
C145 B.n111 VSUBS 0.00771f
C146 B.n112 VSUBS 0.00771f
C147 B.n113 VSUBS 0.00771f
C148 B.n114 VSUBS 0.00771f
C149 B.n115 VSUBS 0.00771f
C150 B.n116 VSUBS 0.00771f
C151 B.n117 VSUBS 0.00771f
C152 B.t7 VSUBS 0.318626f
C153 B.t8 VSUBS 0.334428f
C154 B.t6 VSUBS 0.738882f
C155 B.n118 VSUBS 0.160253f
C156 B.n119 VSUBS 0.074445f
C157 B.n120 VSUBS 0.00771f
C158 B.n121 VSUBS 0.00771f
C159 B.n122 VSUBS 0.00771f
C160 B.n123 VSUBS 0.00771f
C161 B.t4 VSUBS 0.318629f
C162 B.t5 VSUBS 0.334431f
C163 B.t3 VSUBS 0.738882f
C164 B.n124 VSUBS 0.16025f
C165 B.n125 VSUBS 0.074441f
C166 B.n126 VSUBS 0.017863f
C167 B.n127 VSUBS 0.00771f
C168 B.n128 VSUBS 0.00771f
C169 B.n129 VSUBS 0.00771f
C170 B.n130 VSUBS 0.00771f
C171 B.n131 VSUBS 0.00771f
C172 B.n132 VSUBS 0.00771f
C173 B.n133 VSUBS 0.00771f
C174 B.n134 VSUBS 0.00771f
C175 B.n135 VSUBS 0.00771f
C176 B.n136 VSUBS 0.00771f
C177 B.n137 VSUBS 0.00771f
C178 B.n138 VSUBS 0.00771f
C179 B.n139 VSUBS 0.00771f
C180 B.n140 VSUBS 0.00771f
C181 B.n141 VSUBS 0.00771f
C182 B.n142 VSUBS 0.00771f
C183 B.n143 VSUBS 0.017843f
C184 B.n144 VSUBS 0.00771f
C185 B.n145 VSUBS 0.00771f
C186 B.n146 VSUBS 0.00771f
C187 B.n147 VSUBS 0.00771f
C188 B.n148 VSUBS 0.00771f
C189 B.n149 VSUBS 0.00771f
C190 B.n150 VSUBS 0.00771f
C191 B.n151 VSUBS 0.00771f
C192 B.n152 VSUBS 0.00771f
C193 B.n153 VSUBS 0.00771f
C194 B.n154 VSUBS 0.00771f
C195 B.n155 VSUBS 0.00771f
C196 B.n156 VSUBS 0.00771f
C197 B.n157 VSUBS 0.00771f
C198 B.n158 VSUBS 0.00771f
C199 B.n159 VSUBS 0.00771f
C200 B.n160 VSUBS 0.00771f
C201 B.n161 VSUBS 0.00771f
C202 B.n162 VSUBS 0.00771f
C203 B.n163 VSUBS 0.00771f
C204 B.n164 VSUBS 0.00771f
C205 B.n165 VSUBS 0.00771f
C206 B.n166 VSUBS 0.00771f
C207 B.n167 VSUBS 0.00771f
C208 B.n168 VSUBS 0.00771f
C209 B.n169 VSUBS 0.00771f
C210 B.n170 VSUBS 0.00771f
C211 B.n171 VSUBS 0.00771f
C212 B.n172 VSUBS 0.00771f
C213 B.n173 VSUBS 0.00771f
C214 B.n174 VSUBS 0.00771f
C215 B.n175 VSUBS 0.00771f
C216 B.n176 VSUBS 0.00771f
C217 B.n177 VSUBS 0.00771f
C218 B.n178 VSUBS 0.00771f
C219 B.n179 VSUBS 0.00771f
C220 B.n180 VSUBS 0.00771f
C221 B.n181 VSUBS 0.00771f
C222 B.n182 VSUBS 0.00771f
C223 B.n183 VSUBS 0.00771f
C224 B.n184 VSUBS 0.00771f
C225 B.n185 VSUBS 0.00771f
C226 B.n186 VSUBS 0.00771f
C227 B.n187 VSUBS 0.00771f
C228 B.n188 VSUBS 0.00771f
C229 B.n189 VSUBS 0.00771f
C230 B.n190 VSUBS 0.00771f
C231 B.n191 VSUBS 0.00771f
C232 B.n192 VSUBS 0.00771f
C233 B.n193 VSUBS 0.00771f
C234 B.n194 VSUBS 0.00771f
C235 B.n195 VSUBS 0.00771f
C236 B.n196 VSUBS 0.00771f
C237 B.n197 VSUBS 0.00771f
C238 B.n198 VSUBS 0.00771f
C239 B.n199 VSUBS 0.00771f
C240 B.n200 VSUBS 0.00771f
C241 B.n201 VSUBS 0.00771f
C242 B.n202 VSUBS 0.00771f
C243 B.n203 VSUBS 0.00771f
C244 B.n204 VSUBS 0.00771f
C245 B.n205 VSUBS 0.00771f
C246 B.n206 VSUBS 0.00771f
C247 B.n207 VSUBS 0.00771f
C248 B.n208 VSUBS 0.00771f
C249 B.n209 VSUBS 0.00771f
C250 B.n210 VSUBS 0.00771f
C251 B.n211 VSUBS 0.00771f
C252 B.n212 VSUBS 0.00771f
C253 B.n213 VSUBS 0.00771f
C254 B.n214 VSUBS 0.017843f
C255 B.n215 VSUBS 0.018438f
C256 B.n216 VSUBS 0.018438f
C257 B.n217 VSUBS 0.00771f
C258 B.n218 VSUBS 0.00771f
C259 B.n219 VSUBS 0.00771f
C260 B.n220 VSUBS 0.00771f
C261 B.n221 VSUBS 0.00771f
C262 B.n222 VSUBS 0.00771f
C263 B.n223 VSUBS 0.00771f
C264 B.n224 VSUBS 0.00771f
C265 B.n225 VSUBS 0.00771f
C266 B.n226 VSUBS 0.00771f
C267 B.n227 VSUBS 0.00771f
C268 B.n228 VSUBS 0.00771f
C269 B.n229 VSUBS 0.00771f
C270 B.n230 VSUBS 0.00771f
C271 B.n231 VSUBS 0.00771f
C272 B.n232 VSUBS 0.00771f
C273 B.n233 VSUBS 0.00771f
C274 B.n234 VSUBS 0.00771f
C275 B.n235 VSUBS 0.00771f
C276 B.n236 VSUBS 0.00771f
C277 B.n237 VSUBS 0.00771f
C278 B.n238 VSUBS 0.00771f
C279 B.n239 VSUBS 0.00771f
C280 B.n240 VSUBS 0.00771f
C281 B.n241 VSUBS 0.00771f
C282 B.n242 VSUBS 0.00771f
C283 B.n243 VSUBS 0.00771f
C284 B.n244 VSUBS 0.00771f
C285 B.n245 VSUBS 0.00771f
C286 B.n246 VSUBS 0.00771f
C287 B.n247 VSUBS 0.00771f
C288 B.n248 VSUBS 0.00771f
C289 B.n249 VSUBS 0.00771f
C290 B.n250 VSUBS 0.00771f
C291 B.n251 VSUBS 0.00771f
C292 B.n252 VSUBS 0.00771f
C293 B.n253 VSUBS 0.00771f
C294 B.n254 VSUBS 0.00771f
C295 B.n255 VSUBS 0.00771f
C296 B.n256 VSUBS 0.00771f
C297 B.n257 VSUBS 0.00771f
C298 B.n258 VSUBS 0.00771f
C299 B.n259 VSUBS 0.00771f
C300 B.n260 VSUBS 0.00771f
C301 B.n261 VSUBS 0.00771f
C302 B.n262 VSUBS 0.00771f
C303 B.n263 VSUBS 0.007256f
C304 B.n264 VSUBS 0.00771f
C305 B.n265 VSUBS 0.00771f
C306 B.n266 VSUBS 0.004308f
C307 B.n267 VSUBS 0.00771f
C308 B.n268 VSUBS 0.00771f
C309 B.n269 VSUBS 0.00771f
C310 B.n270 VSUBS 0.00771f
C311 B.n271 VSUBS 0.00771f
C312 B.n272 VSUBS 0.00771f
C313 B.n273 VSUBS 0.00771f
C314 B.n274 VSUBS 0.00771f
C315 B.n275 VSUBS 0.00771f
C316 B.n276 VSUBS 0.00771f
C317 B.n277 VSUBS 0.00771f
C318 B.n278 VSUBS 0.00771f
C319 B.n279 VSUBS 0.004308f
C320 B.n280 VSUBS 0.017863f
C321 B.n281 VSUBS 0.007256f
C322 B.n282 VSUBS 0.00771f
C323 B.n283 VSUBS 0.00771f
C324 B.n284 VSUBS 0.00771f
C325 B.n285 VSUBS 0.00771f
C326 B.n286 VSUBS 0.00771f
C327 B.n287 VSUBS 0.00771f
C328 B.n288 VSUBS 0.00771f
C329 B.n289 VSUBS 0.00771f
C330 B.n290 VSUBS 0.00771f
C331 B.n291 VSUBS 0.00771f
C332 B.n292 VSUBS 0.00771f
C333 B.n293 VSUBS 0.00771f
C334 B.n294 VSUBS 0.00771f
C335 B.n295 VSUBS 0.00771f
C336 B.n296 VSUBS 0.00771f
C337 B.n297 VSUBS 0.00771f
C338 B.n298 VSUBS 0.00771f
C339 B.n299 VSUBS 0.00771f
C340 B.n300 VSUBS 0.00771f
C341 B.n301 VSUBS 0.00771f
C342 B.n302 VSUBS 0.00771f
C343 B.n303 VSUBS 0.00771f
C344 B.n304 VSUBS 0.00771f
C345 B.n305 VSUBS 0.00771f
C346 B.n306 VSUBS 0.00771f
C347 B.n307 VSUBS 0.00771f
C348 B.n308 VSUBS 0.00771f
C349 B.n309 VSUBS 0.00771f
C350 B.n310 VSUBS 0.00771f
C351 B.n311 VSUBS 0.00771f
C352 B.n312 VSUBS 0.00771f
C353 B.n313 VSUBS 0.00771f
C354 B.n314 VSUBS 0.00771f
C355 B.n315 VSUBS 0.00771f
C356 B.n316 VSUBS 0.00771f
C357 B.n317 VSUBS 0.00771f
C358 B.n318 VSUBS 0.00771f
C359 B.n319 VSUBS 0.00771f
C360 B.n320 VSUBS 0.00771f
C361 B.n321 VSUBS 0.00771f
C362 B.n322 VSUBS 0.00771f
C363 B.n323 VSUBS 0.00771f
C364 B.n324 VSUBS 0.00771f
C365 B.n325 VSUBS 0.00771f
C366 B.n326 VSUBS 0.00771f
C367 B.n327 VSUBS 0.00771f
C368 B.n328 VSUBS 0.00771f
C369 B.n329 VSUBS 0.018438f
C370 B.n330 VSUBS 0.018438f
C371 B.n331 VSUBS 0.017843f
C372 B.n332 VSUBS 0.00771f
C373 B.n333 VSUBS 0.00771f
C374 B.n334 VSUBS 0.00771f
C375 B.n335 VSUBS 0.00771f
C376 B.n336 VSUBS 0.00771f
C377 B.n337 VSUBS 0.00771f
C378 B.n338 VSUBS 0.00771f
C379 B.n339 VSUBS 0.00771f
C380 B.n340 VSUBS 0.00771f
C381 B.n341 VSUBS 0.00771f
C382 B.n342 VSUBS 0.00771f
C383 B.n343 VSUBS 0.00771f
C384 B.n344 VSUBS 0.00771f
C385 B.n345 VSUBS 0.00771f
C386 B.n346 VSUBS 0.00771f
C387 B.n347 VSUBS 0.00771f
C388 B.n348 VSUBS 0.00771f
C389 B.n349 VSUBS 0.00771f
C390 B.n350 VSUBS 0.00771f
C391 B.n351 VSUBS 0.00771f
C392 B.n352 VSUBS 0.00771f
C393 B.n353 VSUBS 0.00771f
C394 B.n354 VSUBS 0.00771f
C395 B.n355 VSUBS 0.00771f
C396 B.n356 VSUBS 0.00771f
C397 B.n357 VSUBS 0.00771f
C398 B.n358 VSUBS 0.00771f
C399 B.n359 VSUBS 0.00771f
C400 B.n360 VSUBS 0.00771f
C401 B.n361 VSUBS 0.00771f
C402 B.n362 VSUBS 0.00771f
C403 B.n363 VSUBS 0.00771f
C404 B.n364 VSUBS 0.00771f
C405 B.n365 VSUBS 0.00771f
C406 B.n366 VSUBS 0.00771f
C407 B.n367 VSUBS 0.00771f
C408 B.n368 VSUBS 0.00771f
C409 B.n369 VSUBS 0.00771f
C410 B.n370 VSUBS 0.00771f
C411 B.n371 VSUBS 0.00771f
C412 B.n372 VSUBS 0.00771f
C413 B.n373 VSUBS 0.00771f
C414 B.n374 VSUBS 0.00771f
C415 B.n375 VSUBS 0.00771f
C416 B.n376 VSUBS 0.00771f
C417 B.n377 VSUBS 0.00771f
C418 B.n378 VSUBS 0.00771f
C419 B.n379 VSUBS 0.00771f
C420 B.n380 VSUBS 0.00771f
C421 B.n381 VSUBS 0.00771f
C422 B.n382 VSUBS 0.00771f
C423 B.n383 VSUBS 0.00771f
C424 B.n384 VSUBS 0.00771f
C425 B.n385 VSUBS 0.00771f
C426 B.n386 VSUBS 0.00771f
C427 B.n387 VSUBS 0.00771f
C428 B.n388 VSUBS 0.00771f
C429 B.n389 VSUBS 0.00771f
C430 B.n390 VSUBS 0.00771f
C431 B.n391 VSUBS 0.00771f
C432 B.n392 VSUBS 0.00771f
C433 B.n393 VSUBS 0.00771f
C434 B.n394 VSUBS 0.00771f
C435 B.n395 VSUBS 0.00771f
C436 B.n396 VSUBS 0.00771f
C437 B.n397 VSUBS 0.00771f
C438 B.n398 VSUBS 0.00771f
C439 B.n399 VSUBS 0.00771f
C440 B.n400 VSUBS 0.00771f
C441 B.n401 VSUBS 0.00771f
C442 B.n402 VSUBS 0.00771f
C443 B.n403 VSUBS 0.00771f
C444 B.n404 VSUBS 0.00771f
C445 B.n405 VSUBS 0.00771f
C446 B.n406 VSUBS 0.00771f
C447 B.n407 VSUBS 0.00771f
C448 B.n408 VSUBS 0.00771f
C449 B.n409 VSUBS 0.00771f
C450 B.n410 VSUBS 0.00771f
C451 B.n411 VSUBS 0.00771f
C452 B.n412 VSUBS 0.00771f
C453 B.n413 VSUBS 0.00771f
C454 B.n414 VSUBS 0.00771f
C455 B.n415 VSUBS 0.00771f
C456 B.n416 VSUBS 0.00771f
C457 B.n417 VSUBS 0.00771f
C458 B.n418 VSUBS 0.00771f
C459 B.n419 VSUBS 0.00771f
C460 B.n420 VSUBS 0.00771f
C461 B.n421 VSUBS 0.00771f
C462 B.n422 VSUBS 0.00771f
C463 B.n423 VSUBS 0.00771f
C464 B.n424 VSUBS 0.00771f
C465 B.n425 VSUBS 0.00771f
C466 B.n426 VSUBS 0.00771f
C467 B.n427 VSUBS 0.00771f
C468 B.n428 VSUBS 0.00771f
C469 B.n429 VSUBS 0.00771f
C470 B.n430 VSUBS 0.00771f
C471 B.n431 VSUBS 0.00771f
C472 B.n432 VSUBS 0.00771f
C473 B.n433 VSUBS 0.00771f
C474 B.n434 VSUBS 0.00771f
C475 B.n435 VSUBS 0.00771f
C476 B.n436 VSUBS 0.00771f
C477 B.n437 VSUBS 0.00771f
C478 B.n438 VSUBS 0.00771f
C479 B.n439 VSUBS 0.00771f
C480 B.n440 VSUBS 0.00771f
C481 B.n441 VSUBS 0.00771f
C482 B.n442 VSUBS 0.018747f
C483 B.n443 VSUBS 0.017535f
C484 B.n444 VSUBS 0.018438f
C485 B.n445 VSUBS 0.00771f
C486 B.n446 VSUBS 0.00771f
C487 B.n447 VSUBS 0.00771f
C488 B.n448 VSUBS 0.00771f
C489 B.n449 VSUBS 0.00771f
C490 B.n450 VSUBS 0.00771f
C491 B.n451 VSUBS 0.00771f
C492 B.n452 VSUBS 0.00771f
C493 B.n453 VSUBS 0.00771f
C494 B.n454 VSUBS 0.00771f
C495 B.n455 VSUBS 0.00771f
C496 B.n456 VSUBS 0.00771f
C497 B.n457 VSUBS 0.00771f
C498 B.n458 VSUBS 0.00771f
C499 B.n459 VSUBS 0.00771f
C500 B.n460 VSUBS 0.00771f
C501 B.n461 VSUBS 0.00771f
C502 B.n462 VSUBS 0.00771f
C503 B.n463 VSUBS 0.00771f
C504 B.n464 VSUBS 0.00771f
C505 B.n465 VSUBS 0.00771f
C506 B.n466 VSUBS 0.00771f
C507 B.n467 VSUBS 0.00771f
C508 B.n468 VSUBS 0.00771f
C509 B.n469 VSUBS 0.00771f
C510 B.n470 VSUBS 0.00771f
C511 B.n471 VSUBS 0.00771f
C512 B.n472 VSUBS 0.00771f
C513 B.n473 VSUBS 0.00771f
C514 B.n474 VSUBS 0.00771f
C515 B.n475 VSUBS 0.00771f
C516 B.n476 VSUBS 0.00771f
C517 B.n477 VSUBS 0.00771f
C518 B.n478 VSUBS 0.00771f
C519 B.n479 VSUBS 0.00771f
C520 B.n480 VSUBS 0.00771f
C521 B.n481 VSUBS 0.00771f
C522 B.n482 VSUBS 0.00771f
C523 B.n483 VSUBS 0.00771f
C524 B.n484 VSUBS 0.00771f
C525 B.n485 VSUBS 0.00771f
C526 B.n486 VSUBS 0.00771f
C527 B.n487 VSUBS 0.00771f
C528 B.n488 VSUBS 0.00771f
C529 B.n489 VSUBS 0.00771f
C530 B.n490 VSUBS 0.00771f
C531 B.n491 VSUBS 0.007256f
C532 B.n492 VSUBS 0.00771f
C533 B.n493 VSUBS 0.00771f
C534 B.n494 VSUBS 0.004308f
C535 B.n495 VSUBS 0.00771f
C536 B.n496 VSUBS 0.00771f
C537 B.n497 VSUBS 0.00771f
C538 B.n498 VSUBS 0.00771f
C539 B.n499 VSUBS 0.00771f
C540 B.n500 VSUBS 0.00771f
C541 B.n501 VSUBS 0.00771f
C542 B.n502 VSUBS 0.00771f
C543 B.n503 VSUBS 0.00771f
C544 B.n504 VSUBS 0.00771f
C545 B.n505 VSUBS 0.00771f
C546 B.n506 VSUBS 0.00771f
C547 B.n507 VSUBS 0.004308f
C548 B.n508 VSUBS 0.017863f
C549 B.n509 VSUBS 0.007256f
C550 B.n510 VSUBS 0.00771f
C551 B.n511 VSUBS 0.00771f
C552 B.n512 VSUBS 0.00771f
C553 B.n513 VSUBS 0.00771f
C554 B.n514 VSUBS 0.00771f
C555 B.n515 VSUBS 0.00771f
C556 B.n516 VSUBS 0.00771f
C557 B.n517 VSUBS 0.00771f
C558 B.n518 VSUBS 0.00771f
C559 B.n519 VSUBS 0.00771f
C560 B.n520 VSUBS 0.00771f
C561 B.n521 VSUBS 0.00771f
C562 B.n522 VSUBS 0.00771f
C563 B.n523 VSUBS 0.00771f
C564 B.n524 VSUBS 0.00771f
C565 B.n525 VSUBS 0.00771f
C566 B.n526 VSUBS 0.00771f
C567 B.n527 VSUBS 0.00771f
C568 B.n528 VSUBS 0.00771f
C569 B.n529 VSUBS 0.00771f
C570 B.n530 VSUBS 0.00771f
C571 B.n531 VSUBS 0.00771f
C572 B.n532 VSUBS 0.00771f
C573 B.n533 VSUBS 0.00771f
C574 B.n534 VSUBS 0.00771f
C575 B.n535 VSUBS 0.00771f
C576 B.n536 VSUBS 0.00771f
C577 B.n537 VSUBS 0.00771f
C578 B.n538 VSUBS 0.00771f
C579 B.n539 VSUBS 0.00771f
C580 B.n540 VSUBS 0.00771f
C581 B.n541 VSUBS 0.00771f
C582 B.n542 VSUBS 0.00771f
C583 B.n543 VSUBS 0.00771f
C584 B.n544 VSUBS 0.00771f
C585 B.n545 VSUBS 0.00771f
C586 B.n546 VSUBS 0.00771f
C587 B.n547 VSUBS 0.00771f
C588 B.n548 VSUBS 0.00771f
C589 B.n549 VSUBS 0.00771f
C590 B.n550 VSUBS 0.00771f
C591 B.n551 VSUBS 0.00771f
C592 B.n552 VSUBS 0.00771f
C593 B.n553 VSUBS 0.00771f
C594 B.n554 VSUBS 0.00771f
C595 B.n555 VSUBS 0.00771f
C596 B.n556 VSUBS 0.00771f
C597 B.n557 VSUBS 0.018438f
C598 B.n558 VSUBS 0.018438f
C599 B.n559 VSUBS 0.017843f
C600 B.n560 VSUBS 0.00771f
C601 B.n561 VSUBS 0.00771f
C602 B.n562 VSUBS 0.00771f
C603 B.n563 VSUBS 0.00771f
C604 B.n564 VSUBS 0.00771f
C605 B.n565 VSUBS 0.00771f
C606 B.n566 VSUBS 0.00771f
C607 B.n567 VSUBS 0.00771f
C608 B.n568 VSUBS 0.00771f
C609 B.n569 VSUBS 0.00771f
C610 B.n570 VSUBS 0.00771f
C611 B.n571 VSUBS 0.00771f
C612 B.n572 VSUBS 0.00771f
C613 B.n573 VSUBS 0.00771f
C614 B.n574 VSUBS 0.00771f
C615 B.n575 VSUBS 0.00771f
C616 B.n576 VSUBS 0.00771f
C617 B.n577 VSUBS 0.00771f
C618 B.n578 VSUBS 0.00771f
C619 B.n579 VSUBS 0.00771f
C620 B.n580 VSUBS 0.00771f
C621 B.n581 VSUBS 0.00771f
C622 B.n582 VSUBS 0.00771f
C623 B.n583 VSUBS 0.00771f
C624 B.n584 VSUBS 0.00771f
C625 B.n585 VSUBS 0.00771f
C626 B.n586 VSUBS 0.00771f
C627 B.n587 VSUBS 0.00771f
C628 B.n588 VSUBS 0.00771f
C629 B.n589 VSUBS 0.00771f
C630 B.n590 VSUBS 0.00771f
C631 B.n591 VSUBS 0.00771f
C632 B.n592 VSUBS 0.00771f
C633 B.n593 VSUBS 0.00771f
C634 B.n594 VSUBS 0.00771f
C635 B.n595 VSUBS 0.00771f
C636 B.n596 VSUBS 0.00771f
C637 B.n597 VSUBS 0.00771f
C638 B.n598 VSUBS 0.00771f
C639 B.n599 VSUBS 0.00771f
C640 B.n600 VSUBS 0.00771f
C641 B.n601 VSUBS 0.00771f
C642 B.n602 VSUBS 0.00771f
C643 B.n603 VSUBS 0.00771f
C644 B.n604 VSUBS 0.00771f
C645 B.n605 VSUBS 0.00771f
C646 B.n606 VSUBS 0.00771f
C647 B.n607 VSUBS 0.00771f
C648 B.n608 VSUBS 0.00771f
C649 B.n609 VSUBS 0.00771f
C650 B.n610 VSUBS 0.00771f
C651 B.n611 VSUBS 0.00771f
C652 B.n612 VSUBS 0.00771f
C653 B.n613 VSUBS 0.00771f
C654 B.n614 VSUBS 0.00771f
C655 B.n615 VSUBS 0.017458f
C656 VDD1.t1 VSUBS 0.181697f
C657 VDD1.t4 VSUBS 0.181697f
C658 VDD1.n0 VSUBS 1.34103f
C659 VDD1.t5 VSUBS 0.181697f
C660 VDD1.t6 VSUBS 0.181697f
C661 VDD1.n1 VSUBS 1.33998f
C662 VDD1.t0 VSUBS 0.181697f
C663 VDD1.t2 VSUBS 0.181697f
C664 VDD1.n2 VSUBS 1.33998f
C665 VDD1.n3 VSUBS 3.10224f
C666 VDD1.t3 VSUBS 0.181697f
C667 VDD1.t7 VSUBS 0.181697f
C668 VDD1.n4 VSUBS 1.33333f
C669 VDD1.n5 VSUBS 2.68259f
C670 VP.n0 VSUBS 0.04046f
C671 VP.t5 VSUBS 1.63507f
C672 VP.n1 VSUBS 0.054337f
C673 VP.n2 VSUBS 0.04046f
C674 VP.t7 VSUBS 1.63507f
C675 VP.n3 VSUBS 0.058815f
C676 VP.n4 VSUBS 0.04046f
C677 VP.t1 VSUBS 1.63507f
C678 VP.n5 VSUBS 0.063293f
C679 VP.n6 VSUBS 0.04046f
C680 VP.t0 VSUBS 1.63507f
C681 VP.n7 VSUBS 0.054337f
C682 VP.n8 VSUBS 0.04046f
C683 VP.t4 VSUBS 1.63507f
C684 VP.n9 VSUBS 0.058815f
C685 VP.t6 VSUBS 1.78728f
C686 VP.n10 VSUBS 0.694776f
C687 VP.t3 VSUBS 1.63507f
C688 VP.n11 VSUBS 0.680543f
C689 VP.n12 VSUBS 0.055028f
C690 VP.n13 VSUBS 0.259571f
C691 VP.n14 VSUBS 0.04046f
C692 VP.n15 VSUBS 0.04046f
C693 VP.n16 VSUBS 0.058815f
C694 VP.n17 VSUBS 0.055028f
C695 VP.n18 VSUBS 0.602598f
C696 VP.n19 VSUBS 0.057991f
C697 VP.n20 VSUBS 0.04046f
C698 VP.n21 VSUBS 0.04046f
C699 VP.n22 VSUBS 0.04046f
C700 VP.n23 VSUBS 0.063293f
C701 VP.n24 VSUBS 0.052065f
C702 VP.n25 VSUBS 0.692807f
C703 VP.n26 VSUBS 1.82212f
C704 VP.n27 VSUBS 1.85514f
C705 VP.t2 VSUBS 1.63507f
C706 VP.n28 VSUBS 0.692807f
C707 VP.n29 VSUBS 0.052065f
C708 VP.n30 VSUBS 0.04046f
C709 VP.n31 VSUBS 0.04046f
C710 VP.n32 VSUBS 0.04046f
C711 VP.n33 VSUBS 0.054337f
C712 VP.n34 VSUBS 0.057991f
C713 VP.n35 VSUBS 0.602598f
C714 VP.n36 VSUBS 0.055028f
C715 VP.n37 VSUBS 0.04046f
C716 VP.n38 VSUBS 0.04046f
C717 VP.n39 VSUBS 0.04046f
C718 VP.n40 VSUBS 0.058815f
C719 VP.n41 VSUBS 0.055028f
C720 VP.n42 VSUBS 0.602598f
C721 VP.n43 VSUBS 0.057991f
C722 VP.n44 VSUBS 0.04046f
C723 VP.n45 VSUBS 0.04046f
C724 VP.n46 VSUBS 0.04046f
C725 VP.n47 VSUBS 0.063293f
C726 VP.n48 VSUBS 0.052065f
C727 VP.n49 VSUBS 0.692807f
C728 VP.n50 VSUBS 0.039882f
C729 VDD2.t4 VSUBS 0.178864f
C730 VDD2.t3 VSUBS 0.178864f
C731 VDD2.n0 VSUBS 1.31909f
C732 VDD2.t2 VSUBS 0.178864f
C733 VDD2.t7 VSUBS 0.178864f
C734 VDD2.n1 VSUBS 1.31909f
C735 VDD2.n2 VSUBS 3.00181f
C736 VDD2.t1 VSUBS 0.178864f
C737 VDD2.t6 VSUBS 0.178864f
C738 VDD2.n3 VSUBS 1.31254f
C739 VDD2.n4 VSUBS 2.611f
C740 VDD2.t0 VSUBS 0.178864f
C741 VDD2.t5 VSUBS 0.178864f
C742 VDD2.n5 VSUBS 1.31906f
C743 VTAIL.t14 VSUBS 0.183795f
C744 VTAIL.t13 VSUBS 0.183795f
C745 VTAIL.n0 VSUBS 1.22495f
C746 VTAIL.n1 VSUBS 0.696614f
C747 VTAIL.t15 VSUBS 1.64282f
C748 VTAIL.n2 VSUBS 0.813608f
C749 VTAIL.t7 VSUBS 1.64282f
C750 VTAIL.n3 VSUBS 0.813608f
C751 VTAIL.t1 VSUBS 0.183795f
C752 VTAIL.t2 VSUBS 0.183795f
C753 VTAIL.n4 VSUBS 1.22495f
C754 VTAIL.n5 VSUBS 0.829804f
C755 VTAIL.t0 VSUBS 1.64282f
C756 VTAIL.n6 VSUBS 1.90342f
C757 VTAIL.t10 VSUBS 1.64283f
C758 VTAIL.n7 VSUBS 1.90341f
C759 VTAIL.t8 VSUBS 0.183795f
C760 VTAIL.t11 VSUBS 0.183795f
C761 VTAIL.n8 VSUBS 1.22495f
C762 VTAIL.n9 VSUBS 0.829796f
C763 VTAIL.t12 VSUBS 1.64283f
C764 VTAIL.n10 VSUBS 0.813598f
C765 VTAIL.t6 VSUBS 1.64283f
C766 VTAIL.n11 VSUBS 0.813598f
C767 VTAIL.t3 VSUBS 0.183795f
C768 VTAIL.t4 VSUBS 0.183795f
C769 VTAIL.n12 VSUBS 1.22495f
C770 VTAIL.n13 VSUBS 0.829796f
C771 VTAIL.t5 VSUBS 1.64282f
C772 VTAIL.n14 VSUBS 1.90341f
C773 VTAIL.t9 VSUBS 1.64282f
C774 VTAIL.n15 VSUBS 1.89867f
C775 VN.n0 VSUBS 0.039208f
C776 VN.t0 VSUBS 1.58447f
C777 VN.n1 VSUBS 0.052656f
C778 VN.n2 VSUBS 0.039208f
C779 VN.t5 VSUBS 1.58447f
C780 VN.n3 VSUBS 0.056995f
C781 VN.t3 VSUBS 1.73197f
C782 VN.n4 VSUBS 0.673275f
C783 VN.t4 VSUBS 1.58447f
C784 VN.n5 VSUBS 0.659482f
C785 VN.n6 VSUBS 0.053325f
C786 VN.n7 VSUBS 0.251538f
C787 VN.n8 VSUBS 0.039208f
C788 VN.n9 VSUBS 0.039208f
C789 VN.n10 VSUBS 0.056995f
C790 VN.n11 VSUBS 0.053325f
C791 VN.n12 VSUBS 0.58395f
C792 VN.n13 VSUBS 0.056196f
C793 VN.n14 VSUBS 0.039208f
C794 VN.n15 VSUBS 0.039208f
C795 VN.n16 VSUBS 0.039208f
C796 VN.n17 VSUBS 0.061334f
C797 VN.n18 VSUBS 0.050453f
C798 VN.n19 VSUBS 0.671366f
C799 VN.n20 VSUBS 0.038648f
C800 VN.n21 VSUBS 0.039208f
C801 VN.t6 VSUBS 1.58447f
C802 VN.n22 VSUBS 0.052656f
C803 VN.n23 VSUBS 0.039208f
C804 VN.t1 VSUBS 1.58447f
C805 VN.n24 VSUBS 0.056995f
C806 VN.t2 VSUBS 1.73197f
C807 VN.n25 VSUBS 0.673275f
C808 VN.t7 VSUBS 1.58447f
C809 VN.n26 VSUBS 0.659482f
C810 VN.n27 VSUBS 0.053325f
C811 VN.n28 VSUBS 0.251538f
C812 VN.n29 VSUBS 0.039208f
C813 VN.n30 VSUBS 0.039208f
C814 VN.n31 VSUBS 0.056995f
C815 VN.n32 VSUBS 0.053325f
C816 VN.n33 VSUBS 0.58395f
C817 VN.n34 VSUBS 0.056196f
C818 VN.n35 VSUBS 0.039208f
C819 VN.n36 VSUBS 0.039208f
C820 VN.n37 VSUBS 0.039208f
C821 VN.n38 VSUBS 0.061334f
C822 VN.n39 VSUBS 0.050453f
C823 VN.n40 VSUBS 0.671366f
C824 VN.n41 VSUBS 1.79139f
.ends

