* NGSPICE file created from diff_pair_sample_0880.ext - technology: sky130A

.subckt diff_pair_sample_0880 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=2.8587 pd=15.44 as=0 ps=0 w=7.33 l=3.79
X1 VTAIL.t15 VN.t0 VDD2.t0 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=2.8587 pd=15.44 as=1.20945 ps=7.66 w=7.33 l=3.79
X2 VDD2.t1 VN.t1 VTAIL.t14 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=3.79
X3 B.t8 B.t6 B.t7 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=2.8587 pd=15.44 as=0 ps=0 w=7.33 l=3.79
X4 VTAIL.t13 VN.t2 VDD2.t2 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=3.79
X5 VTAIL.t12 VN.t3 VDD2.t3 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=3.79
X6 VDD1.t7 VP.t0 VTAIL.t6 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=3.79
X7 VDD2.t4 VN.t4 VTAIL.t11 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=2.8587 ps=15.44 w=7.33 l=3.79
X8 VDD1.t6 VP.t1 VTAIL.t0 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=2.8587 ps=15.44 w=7.33 l=3.79
X9 VTAIL.t5 VP.t2 VDD1.t5 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=2.8587 pd=15.44 as=1.20945 ps=7.66 w=7.33 l=3.79
X10 VDD2.t5 VN.t5 VTAIL.t10 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=2.8587 ps=15.44 w=7.33 l=3.79
X11 VTAIL.t3 VP.t3 VDD1.t4 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=2.8587 pd=15.44 as=1.20945 ps=7.66 w=7.33 l=3.79
X12 VTAIL.t4 VP.t4 VDD1.t3 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=3.79
X13 VDD2.t6 VN.t6 VTAIL.t9 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=3.79
X14 VDD1.t2 VP.t5 VTAIL.t1 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=3.79
X15 B.t5 B.t3 B.t4 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=2.8587 pd=15.44 as=0 ps=0 w=7.33 l=3.79
X16 VTAIL.t7 VP.t6 VDD1.t1 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=1.20945 ps=7.66 w=7.33 l=3.79
X17 VTAIL.t8 VN.t7 VDD2.t7 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=2.8587 pd=15.44 as=1.20945 ps=7.66 w=7.33 l=3.79
X18 B.t2 B.t0 B.t1 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=2.8587 pd=15.44 as=0 ps=0 w=7.33 l=3.79
X19 VDD1.t0 VP.t7 VTAIL.t2 w_n5090_n2434# sky130_fd_pr__pfet_01v8 ad=1.20945 pd=7.66 as=2.8587 ps=15.44 w=7.33 l=3.79
R0 B.n411 B.n142 585
R1 B.n410 B.n409 585
R2 B.n408 B.n143 585
R3 B.n407 B.n406 585
R4 B.n405 B.n144 585
R5 B.n404 B.n403 585
R6 B.n402 B.n145 585
R7 B.n401 B.n400 585
R8 B.n399 B.n146 585
R9 B.n398 B.n397 585
R10 B.n396 B.n147 585
R11 B.n395 B.n394 585
R12 B.n393 B.n148 585
R13 B.n392 B.n391 585
R14 B.n390 B.n149 585
R15 B.n389 B.n388 585
R16 B.n387 B.n150 585
R17 B.n386 B.n385 585
R18 B.n384 B.n151 585
R19 B.n383 B.n382 585
R20 B.n381 B.n152 585
R21 B.n380 B.n379 585
R22 B.n378 B.n153 585
R23 B.n377 B.n376 585
R24 B.n375 B.n154 585
R25 B.n374 B.n373 585
R26 B.n372 B.n155 585
R27 B.n371 B.n370 585
R28 B.n369 B.n368 585
R29 B.n367 B.n159 585
R30 B.n366 B.n365 585
R31 B.n364 B.n160 585
R32 B.n363 B.n362 585
R33 B.n361 B.n161 585
R34 B.n360 B.n359 585
R35 B.n358 B.n162 585
R36 B.n357 B.n356 585
R37 B.n354 B.n163 585
R38 B.n353 B.n352 585
R39 B.n351 B.n166 585
R40 B.n350 B.n349 585
R41 B.n348 B.n167 585
R42 B.n347 B.n346 585
R43 B.n345 B.n168 585
R44 B.n344 B.n343 585
R45 B.n342 B.n169 585
R46 B.n341 B.n340 585
R47 B.n339 B.n170 585
R48 B.n338 B.n337 585
R49 B.n336 B.n171 585
R50 B.n335 B.n334 585
R51 B.n333 B.n172 585
R52 B.n332 B.n331 585
R53 B.n330 B.n173 585
R54 B.n329 B.n328 585
R55 B.n327 B.n174 585
R56 B.n326 B.n325 585
R57 B.n324 B.n175 585
R58 B.n323 B.n322 585
R59 B.n321 B.n176 585
R60 B.n320 B.n319 585
R61 B.n318 B.n177 585
R62 B.n317 B.n316 585
R63 B.n315 B.n178 585
R64 B.n314 B.n313 585
R65 B.n413 B.n412 585
R66 B.n414 B.n141 585
R67 B.n416 B.n415 585
R68 B.n417 B.n140 585
R69 B.n419 B.n418 585
R70 B.n420 B.n139 585
R71 B.n422 B.n421 585
R72 B.n423 B.n138 585
R73 B.n425 B.n424 585
R74 B.n426 B.n137 585
R75 B.n428 B.n427 585
R76 B.n429 B.n136 585
R77 B.n431 B.n430 585
R78 B.n432 B.n135 585
R79 B.n434 B.n433 585
R80 B.n435 B.n134 585
R81 B.n437 B.n436 585
R82 B.n438 B.n133 585
R83 B.n440 B.n439 585
R84 B.n441 B.n132 585
R85 B.n443 B.n442 585
R86 B.n444 B.n131 585
R87 B.n446 B.n445 585
R88 B.n447 B.n130 585
R89 B.n449 B.n448 585
R90 B.n450 B.n129 585
R91 B.n452 B.n451 585
R92 B.n453 B.n128 585
R93 B.n455 B.n454 585
R94 B.n456 B.n127 585
R95 B.n458 B.n457 585
R96 B.n459 B.n126 585
R97 B.n461 B.n460 585
R98 B.n462 B.n125 585
R99 B.n464 B.n463 585
R100 B.n465 B.n124 585
R101 B.n467 B.n466 585
R102 B.n468 B.n123 585
R103 B.n470 B.n469 585
R104 B.n471 B.n122 585
R105 B.n473 B.n472 585
R106 B.n474 B.n121 585
R107 B.n476 B.n475 585
R108 B.n477 B.n120 585
R109 B.n479 B.n478 585
R110 B.n480 B.n119 585
R111 B.n482 B.n481 585
R112 B.n483 B.n118 585
R113 B.n485 B.n484 585
R114 B.n486 B.n117 585
R115 B.n488 B.n487 585
R116 B.n489 B.n116 585
R117 B.n491 B.n490 585
R118 B.n492 B.n115 585
R119 B.n494 B.n493 585
R120 B.n495 B.n114 585
R121 B.n497 B.n496 585
R122 B.n498 B.n113 585
R123 B.n500 B.n499 585
R124 B.n501 B.n112 585
R125 B.n503 B.n502 585
R126 B.n504 B.n111 585
R127 B.n506 B.n505 585
R128 B.n507 B.n110 585
R129 B.n509 B.n508 585
R130 B.n510 B.n109 585
R131 B.n512 B.n511 585
R132 B.n513 B.n108 585
R133 B.n515 B.n514 585
R134 B.n516 B.n107 585
R135 B.n518 B.n517 585
R136 B.n519 B.n106 585
R137 B.n521 B.n520 585
R138 B.n522 B.n105 585
R139 B.n524 B.n523 585
R140 B.n525 B.n104 585
R141 B.n527 B.n526 585
R142 B.n528 B.n103 585
R143 B.n530 B.n529 585
R144 B.n531 B.n102 585
R145 B.n533 B.n532 585
R146 B.n534 B.n101 585
R147 B.n536 B.n535 585
R148 B.n537 B.n100 585
R149 B.n539 B.n538 585
R150 B.n540 B.n99 585
R151 B.n542 B.n541 585
R152 B.n543 B.n98 585
R153 B.n545 B.n544 585
R154 B.n546 B.n97 585
R155 B.n548 B.n547 585
R156 B.n549 B.n96 585
R157 B.n551 B.n550 585
R158 B.n552 B.n95 585
R159 B.n554 B.n553 585
R160 B.n555 B.n94 585
R161 B.n557 B.n556 585
R162 B.n558 B.n93 585
R163 B.n560 B.n559 585
R164 B.n561 B.n92 585
R165 B.n563 B.n562 585
R166 B.n564 B.n91 585
R167 B.n566 B.n565 585
R168 B.n567 B.n90 585
R169 B.n569 B.n568 585
R170 B.n570 B.n89 585
R171 B.n572 B.n571 585
R172 B.n573 B.n88 585
R173 B.n575 B.n574 585
R174 B.n576 B.n87 585
R175 B.n578 B.n577 585
R176 B.n579 B.n86 585
R177 B.n581 B.n580 585
R178 B.n582 B.n85 585
R179 B.n584 B.n583 585
R180 B.n585 B.n84 585
R181 B.n587 B.n586 585
R182 B.n588 B.n83 585
R183 B.n590 B.n589 585
R184 B.n591 B.n82 585
R185 B.n593 B.n592 585
R186 B.n594 B.n81 585
R187 B.n596 B.n595 585
R188 B.n597 B.n80 585
R189 B.n599 B.n598 585
R190 B.n600 B.n79 585
R191 B.n602 B.n601 585
R192 B.n603 B.n78 585
R193 B.n605 B.n604 585
R194 B.n606 B.n77 585
R195 B.n608 B.n607 585
R196 B.n609 B.n76 585
R197 B.n611 B.n610 585
R198 B.n612 B.n75 585
R199 B.n614 B.n613 585
R200 B.n615 B.n74 585
R201 B.n617 B.n616 585
R202 B.n618 B.n73 585
R203 B.n717 B.n36 585
R204 B.n716 B.n715 585
R205 B.n714 B.n37 585
R206 B.n713 B.n712 585
R207 B.n711 B.n38 585
R208 B.n710 B.n709 585
R209 B.n708 B.n39 585
R210 B.n707 B.n706 585
R211 B.n705 B.n40 585
R212 B.n704 B.n703 585
R213 B.n702 B.n41 585
R214 B.n701 B.n700 585
R215 B.n699 B.n42 585
R216 B.n698 B.n697 585
R217 B.n696 B.n43 585
R218 B.n695 B.n694 585
R219 B.n693 B.n44 585
R220 B.n692 B.n691 585
R221 B.n690 B.n45 585
R222 B.n689 B.n688 585
R223 B.n687 B.n46 585
R224 B.n686 B.n685 585
R225 B.n684 B.n47 585
R226 B.n683 B.n682 585
R227 B.n681 B.n48 585
R228 B.n680 B.n679 585
R229 B.n678 B.n49 585
R230 B.n677 B.n676 585
R231 B.n675 B.n674 585
R232 B.n673 B.n53 585
R233 B.n672 B.n671 585
R234 B.n670 B.n54 585
R235 B.n669 B.n668 585
R236 B.n667 B.n55 585
R237 B.n666 B.n665 585
R238 B.n664 B.n56 585
R239 B.n663 B.n662 585
R240 B.n660 B.n57 585
R241 B.n659 B.n658 585
R242 B.n657 B.n60 585
R243 B.n656 B.n655 585
R244 B.n654 B.n61 585
R245 B.n653 B.n652 585
R246 B.n651 B.n62 585
R247 B.n650 B.n649 585
R248 B.n648 B.n63 585
R249 B.n647 B.n646 585
R250 B.n645 B.n64 585
R251 B.n644 B.n643 585
R252 B.n642 B.n65 585
R253 B.n641 B.n640 585
R254 B.n639 B.n66 585
R255 B.n638 B.n637 585
R256 B.n636 B.n67 585
R257 B.n635 B.n634 585
R258 B.n633 B.n68 585
R259 B.n632 B.n631 585
R260 B.n630 B.n69 585
R261 B.n629 B.n628 585
R262 B.n627 B.n70 585
R263 B.n626 B.n625 585
R264 B.n624 B.n71 585
R265 B.n623 B.n622 585
R266 B.n621 B.n72 585
R267 B.n620 B.n619 585
R268 B.n719 B.n718 585
R269 B.n720 B.n35 585
R270 B.n722 B.n721 585
R271 B.n723 B.n34 585
R272 B.n725 B.n724 585
R273 B.n726 B.n33 585
R274 B.n728 B.n727 585
R275 B.n729 B.n32 585
R276 B.n731 B.n730 585
R277 B.n732 B.n31 585
R278 B.n734 B.n733 585
R279 B.n735 B.n30 585
R280 B.n737 B.n736 585
R281 B.n738 B.n29 585
R282 B.n740 B.n739 585
R283 B.n741 B.n28 585
R284 B.n743 B.n742 585
R285 B.n744 B.n27 585
R286 B.n746 B.n745 585
R287 B.n747 B.n26 585
R288 B.n749 B.n748 585
R289 B.n750 B.n25 585
R290 B.n752 B.n751 585
R291 B.n753 B.n24 585
R292 B.n755 B.n754 585
R293 B.n756 B.n23 585
R294 B.n758 B.n757 585
R295 B.n759 B.n22 585
R296 B.n761 B.n760 585
R297 B.n762 B.n21 585
R298 B.n764 B.n763 585
R299 B.n765 B.n20 585
R300 B.n767 B.n766 585
R301 B.n768 B.n19 585
R302 B.n770 B.n769 585
R303 B.n771 B.n18 585
R304 B.n773 B.n772 585
R305 B.n774 B.n17 585
R306 B.n776 B.n775 585
R307 B.n777 B.n16 585
R308 B.n779 B.n778 585
R309 B.n780 B.n15 585
R310 B.n782 B.n781 585
R311 B.n783 B.n14 585
R312 B.n785 B.n784 585
R313 B.n786 B.n13 585
R314 B.n788 B.n787 585
R315 B.n789 B.n12 585
R316 B.n791 B.n790 585
R317 B.n792 B.n11 585
R318 B.n794 B.n793 585
R319 B.n795 B.n10 585
R320 B.n797 B.n796 585
R321 B.n798 B.n9 585
R322 B.n800 B.n799 585
R323 B.n801 B.n8 585
R324 B.n803 B.n802 585
R325 B.n804 B.n7 585
R326 B.n806 B.n805 585
R327 B.n807 B.n6 585
R328 B.n809 B.n808 585
R329 B.n810 B.n5 585
R330 B.n812 B.n811 585
R331 B.n813 B.n4 585
R332 B.n815 B.n814 585
R333 B.n816 B.n3 585
R334 B.n818 B.n817 585
R335 B.n819 B.n0 585
R336 B.n2 B.n1 585
R337 B.n213 B.n212 585
R338 B.n215 B.n214 585
R339 B.n216 B.n211 585
R340 B.n218 B.n217 585
R341 B.n219 B.n210 585
R342 B.n221 B.n220 585
R343 B.n222 B.n209 585
R344 B.n224 B.n223 585
R345 B.n225 B.n208 585
R346 B.n227 B.n226 585
R347 B.n228 B.n207 585
R348 B.n230 B.n229 585
R349 B.n231 B.n206 585
R350 B.n233 B.n232 585
R351 B.n234 B.n205 585
R352 B.n236 B.n235 585
R353 B.n237 B.n204 585
R354 B.n239 B.n238 585
R355 B.n240 B.n203 585
R356 B.n242 B.n241 585
R357 B.n243 B.n202 585
R358 B.n245 B.n244 585
R359 B.n246 B.n201 585
R360 B.n248 B.n247 585
R361 B.n249 B.n200 585
R362 B.n251 B.n250 585
R363 B.n252 B.n199 585
R364 B.n254 B.n253 585
R365 B.n255 B.n198 585
R366 B.n257 B.n256 585
R367 B.n258 B.n197 585
R368 B.n260 B.n259 585
R369 B.n261 B.n196 585
R370 B.n263 B.n262 585
R371 B.n264 B.n195 585
R372 B.n266 B.n265 585
R373 B.n267 B.n194 585
R374 B.n269 B.n268 585
R375 B.n270 B.n193 585
R376 B.n272 B.n271 585
R377 B.n273 B.n192 585
R378 B.n275 B.n274 585
R379 B.n276 B.n191 585
R380 B.n278 B.n277 585
R381 B.n279 B.n190 585
R382 B.n281 B.n280 585
R383 B.n282 B.n189 585
R384 B.n284 B.n283 585
R385 B.n285 B.n188 585
R386 B.n287 B.n286 585
R387 B.n288 B.n187 585
R388 B.n290 B.n289 585
R389 B.n291 B.n186 585
R390 B.n293 B.n292 585
R391 B.n294 B.n185 585
R392 B.n296 B.n295 585
R393 B.n297 B.n184 585
R394 B.n299 B.n298 585
R395 B.n300 B.n183 585
R396 B.n302 B.n301 585
R397 B.n303 B.n182 585
R398 B.n305 B.n304 585
R399 B.n306 B.n181 585
R400 B.n308 B.n307 585
R401 B.n309 B.n180 585
R402 B.n311 B.n310 585
R403 B.n312 B.n179 585
R404 B.n314 B.n179 559.769
R405 B.n412 B.n411 559.769
R406 B.n620 B.n73 559.769
R407 B.n718 B.n717 559.769
R408 B.n156 B.t7 371.616
R409 B.n58 B.t2 371.616
R410 B.n164 B.t4 371.616
R411 B.n50 B.t11 371.616
R412 B.n157 B.t8 291.714
R413 B.n59 B.t1 291.714
R414 B.n165 B.t5 291.714
R415 B.n51 B.t10 291.714
R416 B.n821 B.n820 256.663
R417 B.n164 B.t3 255.946
R418 B.n156 B.t6 255.946
R419 B.n58 B.t0 255.946
R420 B.n50 B.t9 255.946
R421 B.n820 B.n819 235.042
R422 B.n820 B.n2 235.042
R423 B.n315 B.n314 163.367
R424 B.n316 B.n315 163.367
R425 B.n316 B.n177 163.367
R426 B.n320 B.n177 163.367
R427 B.n321 B.n320 163.367
R428 B.n322 B.n321 163.367
R429 B.n322 B.n175 163.367
R430 B.n326 B.n175 163.367
R431 B.n327 B.n326 163.367
R432 B.n328 B.n327 163.367
R433 B.n328 B.n173 163.367
R434 B.n332 B.n173 163.367
R435 B.n333 B.n332 163.367
R436 B.n334 B.n333 163.367
R437 B.n334 B.n171 163.367
R438 B.n338 B.n171 163.367
R439 B.n339 B.n338 163.367
R440 B.n340 B.n339 163.367
R441 B.n340 B.n169 163.367
R442 B.n344 B.n169 163.367
R443 B.n345 B.n344 163.367
R444 B.n346 B.n345 163.367
R445 B.n346 B.n167 163.367
R446 B.n350 B.n167 163.367
R447 B.n351 B.n350 163.367
R448 B.n352 B.n351 163.367
R449 B.n352 B.n163 163.367
R450 B.n357 B.n163 163.367
R451 B.n358 B.n357 163.367
R452 B.n359 B.n358 163.367
R453 B.n359 B.n161 163.367
R454 B.n363 B.n161 163.367
R455 B.n364 B.n363 163.367
R456 B.n365 B.n364 163.367
R457 B.n365 B.n159 163.367
R458 B.n369 B.n159 163.367
R459 B.n370 B.n369 163.367
R460 B.n370 B.n155 163.367
R461 B.n374 B.n155 163.367
R462 B.n375 B.n374 163.367
R463 B.n376 B.n375 163.367
R464 B.n376 B.n153 163.367
R465 B.n380 B.n153 163.367
R466 B.n381 B.n380 163.367
R467 B.n382 B.n381 163.367
R468 B.n382 B.n151 163.367
R469 B.n386 B.n151 163.367
R470 B.n387 B.n386 163.367
R471 B.n388 B.n387 163.367
R472 B.n388 B.n149 163.367
R473 B.n392 B.n149 163.367
R474 B.n393 B.n392 163.367
R475 B.n394 B.n393 163.367
R476 B.n394 B.n147 163.367
R477 B.n398 B.n147 163.367
R478 B.n399 B.n398 163.367
R479 B.n400 B.n399 163.367
R480 B.n400 B.n145 163.367
R481 B.n404 B.n145 163.367
R482 B.n405 B.n404 163.367
R483 B.n406 B.n405 163.367
R484 B.n406 B.n143 163.367
R485 B.n410 B.n143 163.367
R486 B.n411 B.n410 163.367
R487 B.n616 B.n73 163.367
R488 B.n616 B.n615 163.367
R489 B.n615 B.n614 163.367
R490 B.n614 B.n75 163.367
R491 B.n610 B.n75 163.367
R492 B.n610 B.n609 163.367
R493 B.n609 B.n608 163.367
R494 B.n608 B.n77 163.367
R495 B.n604 B.n77 163.367
R496 B.n604 B.n603 163.367
R497 B.n603 B.n602 163.367
R498 B.n602 B.n79 163.367
R499 B.n598 B.n79 163.367
R500 B.n598 B.n597 163.367
R501 B.n597 B.n596 163.367
R502 B.n596 B.n81 163.367
R503 B.n592 B.n81 163.367
R504 B.n592 B.n591 163.367
R505 B.n591 B.n590 163.367
R506 B.n590 B.n83 163.367
R507 B.n586 B.n83 163.367
R508 B.n586 B.n585 163.367
R509 B.n585 B.n584 163.367
R510 B.n584 B.n85 163.367
R511 B.n580 B.n85 163.367
R512 B.n580 B.n579 163.367
R513 B.n579 B.n578 163.367
R514 B.n578 B.n87 163.367
R515 B.n574 B.n87 163.367
R516 B.n574 B.n573 163.367
R517 B.n573 B.n572 163.367
R518 B.n572 B.n89 163.367
R519 B.n568 B.n89 163.367
R520 B.n568 B.n567 163.367
R521 B.n567 B.n566 163.367
R522 B.n566 B.n91 163.367
R523 B.n562 B.n91 163.367
R524 B.n562 B.n561 163.367
R525 B.n561 B.n560 163.367
R526 B.n560 B.n93 163.367
R527 B.n556 B.n93 163.367
R528 B.n556 B.n555 163.367
R529 B.n555 B.n554 163.367
R530 B.n554 B.n95 163.367
R531 B.n550 B.n95 163.367
R532 B.n550 B.n549 163.367
R533 B.n549 B.n548 163.367
R534 B.n548 B.n97 163.367
R535 B.n544 B.n97 163.367
R536 B.n544 B.n543 163.367
R537 B.n543 B.n542 163.367
R538 B.n542 B.n99 163.367
R539 B.n538 B.n99 163.367
R540 B.n538 B.n537 163.367
R541 B.n537 B.n536 163.367
R542 B.n536 B.n101 163.367
R543 B.n532 B.n101 163.367
R544 B.n532 B.n531 163.367
R545 B.n531 B.n530 163.367
R546 B.n530 B.n103 163.367
R547 B.n526 B.n103 163.367
R548 B.n526 B.n525 163.367
R549 B.n525 B.n524 163.367
R550 B.n524 B.n105 163.367
R551 B.n520 B.n105 163.367
R552 B.n520 B.n519 163.367
R553 B.n519 B.n518 163.367
R554 B.n518 B.n107 163.367
R555 B.n514 B.n107 163.367
R556 B.n514 B.n513 163.367
R557 B.n513 B.n512 163.367
R558 B.n512 B.n109 163.367
R559 B.n508 B.n109 163.367
R560 B.n508 B.n507 163.367
R561 B.n507 B.n506 163.367
R562 B.n506 B.n111 163.367
R563 B.n502 B.n111 163.367
R564 B.n502 B.n501 163.367
R565 B.n501 B.n500 163.367
R566 B.n500 B.n113 163.367
R567 B.n496 B.n113 163.367
R568 B.n496 B.n495 163.367
R569 B.n495 B.n494 163.367
R570 B.n494 B.n115 163.367
R571 B.n490 B.n115 163.367
R572 B.n490 B.n489 163.367
R573 B.n489 B.n488 163.367
R574 B.n488 B.n117 163.367
R575 B.n484 B.n117 163.367
R576 B.n484 B.n483 163.367
R577 B.n483 B.n482 163.367
R578 B.n482 B.n119 163.367
R579 B.n478 B.n119 163.367
R580 B.n478 B.n477 163.367
R581 B.n477 B.n476 163.367
R582 B.n476 B.n121 163.367
R583 B.n472 B.n121 163.367
R584 B.n472 B.n471 163.367
R585 B.n471 B.n470 163.367
R586 B.n470 B.n123 163.367
R587 B.n466 B.n123 163.367
R588 B.n466 B.n465 163.367
R589 B.n465 B.n464 163.367
R590 B.n464 B.n125 163.367
R591 B.n460 B.n125 163.367
R592 B.n460 B.n459 163.367
R593 B.n459 B.n458 163.367
R594 B.n458 B.n127 163.367
R595 B.n454 B.n127 163.367
R596 B.n454 B.n453 163.367
R597 B.n453 B.n452 163.367
R598 B.n452 B.n129 163.367
R599 B.n448 B.n129 163.367
R600 B.n448 B.n447 163.367
R601 B.n447 B.n446 163.367
R602 B.n446 B.n131 163.367
R603 B.n442 B.n131 163.367
R604 B.n442 B.n441 163.367
R605 B.n441 B.n440 163.367
R606 B.n440 B.n133 163.367
R607 B.n436 B.n133 163.367
R608 B.n436 B.n435 163.367
R609 B.n435 B.n434 163.367
R610 B.n434 B.n135 163.367
R611 B.n430 B.n135 163.367
R612 B.n430 B.n429 163.367
R613 B.n429 B.n428 163.367
R614 B.n428 B.n137 163.367
R615 B.n424 B.n137 163.367
R616 B.n424 B.n423 163.367
R617 B.n423 B.n422 163.367
R618 B.n422 B.n139 163.367
R619 B.n418 B.n139 163.367
R620 B.n418 B.n417 163.367
R621 B.n417 B.n416 163.367
R622 B.n416 B.n141 163.367
R623 B.n412 B.n141 163.367
R624 B.n717 B.n716 163.367
R625 B.n716 B.n37 163.367
R626 B.n712 B.n37 163.367
R627 B.n712 B.n711 163.367
R628 B.n711 B.n710 163.367
R629 B.n710 B.n39 163.367
R630 B.n706 B.n39 163.367
R631 B.n706 B.n705 163.367
R632 B.n705 B.n704 163.367
R633 B.n704 B.n41 163.367
R634 B.n700 B.n41 163.367
R635 B.n700 B.n699 163.367
R636 B.n699 B.n698 163.367
R637 B.n698 B.n43 163.367
R638 B.n694 B.n43 163.367
R639 B.n694 B.n693 163.367
R640 B.n693 B.n692 163.367
R641 B.n692 B.n45 163.367
R642 B.n688 B.n45 163.367
R643 B.n688 B.n687 163.367
R644 B.n687 B.n686 163.367
R645 B.n686 B.n47 163.367
R646 B.n682 B.n47 163.367
R647 B.n682 B.n681 163.367
R648 B.n681 B.n680 163.367
R649 B.n680 B.n49 163.367
R650 B.n676 B.n49 163.367
R651 B.n676 B.n675 163.367
R652 B.n675 B.n53 163.367
R653 B.n671 B.n53 163.367
R654 B.n671 B.n670 163.367
R655 B.n670 B.n669 163.367
R656 B.n669 B.n55 163.367
R657 B.n665 B.n55 163.367
R658 B.n665 B.n664 163.367
R659 B.n664 B.n663 163.367
R660 B.n663 B.n57 163.367
R661 B.n658 B.n57 163.367
R662 B.n658 B.n657 163.367
R663 B.n657 B.n656 163.367
R664 B.n656 B.n61 163.367
R665 B.n652 B.n61 163.367
R666 B.n652 B.n651 163.367
R667 B.n651 B.n650 163.367
R668 B.n650 B.n63 163.367
R669 B.n646 B.n63 163.367
R670 B.n646 B.n645 163.367
R671 B.n645 B.n644 163.367
R672 B.n644 B.n65 163.367
R673 B.n640 B.n65 163.367
R674 B.n640 B.n639 163.367
R675 B.n639 B.n638 163.367
R676 B.n638 B.n67 163.367
R677 B.n634 B.n67 163.367
R678 B.n634 B.n633 163.367
R679 B.n633 B.n632 163.367
R680 B.n632 B.n69 163.367
R681 B.n628 B.n69 163.367
R682 B.n628 B.n627 163.367
R683 B.n627 B.n626 163.367
R684 B.n626 B.n71 163.367
R685 B.n622 B.n71 163.367
R686 B.n622 B.n621 163.367
R687 B.n621 B.n620 163.367
R688 B.n718 B.n35 163.367
R689 B.n722 B.n35 163.367
R690 B.n723 B.n722 163.367
R691 B.n724 B.n723 163.367
R692 B.n724 B.n33 163.367
R693 B.n728 B.n33 163.367
R694 B.n729 B.n728 163.367
R695 B.n730 B.n729 163.367
R696 B.n730 B.n31 163.367
R697 B.n734 B.n31 163.367
R698 B.n735 B.n734 163.367
R699 B.n736 B.n735 163.367
R700 B.n736 B.n29 163.367
R701 B.n740 B.n29 163.367
R702 B.n741 B.n740 163.367
R703 B.n742 B.n741 163.367
R704 B.n742 B.n27 163.367
R705 B.n746 B.n27 163.367
R706 B.n747 B.n746 163.367
R707 B.n748 B.n747 163.367
R708 B.n748 B.n25 163.367
R709 B.n752 B.n25 163.367
R710 B.n753 B.n752 163.367
R711 B.n754 B.n753 163.367
R712 B.n754 B.n23 163.367
R713 B.n758 B.n23 163.367
R714 B.n759 B.n758 163.367
R715 B.n760 B.n759 163.367
R716 B.n760 B.n21 163.367
R717 B.n764 B.n21 163.367
R718 B.n765 B.n764 163.367
R719 B.n766 B.n765 163.367
R720 B.n766 B.n19 163.367
R721 B.n770 B.n19 163.367
R722 B.n771 B.n770 163.367
R723 B.n772 B.n771 163.367
R724 B.n772 B.n17 163.367
R725 B.n776 B.n17 163.367
R726 B.n777 B.n776 163.367
R727 B.n778 B.n777 163.367
R728 B.n778 B.n15 163.367
R729 B.n782 B.n15 163.367
R730 B.n783 B.n782 163.367
R731 B.n784 B.n783 163.367
R732 B.n784 B.n13 163.367
R733 B.n788 B.n13 163.367
R734 B.n789 B.n788 163.367
R735 B.n790 B.n789 163.367
R736 B.n790 B.n11 163.367
R737 B.n794 B.n11 163.367
R738 B.n795 B.n794 163.367
R739 B.n796 B.n795 163.367
R740 B.n796 B.n9 163.367
R741 B.n800 B.n9 163.367
R742 B.n801 B.n800 163.367
R743 B.n802 B.n801 163.367
R744 B.n802 B.n7 163.367
R745 B.n806 B.n7 163.367
R746 B.n807 B.n806 163.367
R747 B.n808 B.n807 163.367
R748 B.n808 B.n5 163.367
R749 B.n812 B.n5 163.367
R750 B.n813 B.n812 163.367
R751 B.n814 B.n813 163.367
R752 B.n814 B.n3 163.367
R753 B.n818 B.n3 163.367
R754 B.n819 B.n818 163.367
R755 B.n213 B.n2 163.367
R756 B.n214 B.n213 163.367
R757 B.n214 B.n211 163.367
R758 B.n218 B.n211 163.367
R759 B.n219 B.n218 163.367
R760 B.n220 B.n219 163.367
R761 B.n220 B.n209 163.367
R762 B.n224 B.n209 163.367
R763 B.n225 B.n224 163.367
R764 B.n226 B.n225 163.367
R765 B.n226 B.n207 163.367
R766 B.n230 B.n207 163.367
R767 B.n231 B.n230 163.367
R768 B.n232 B.n231 163.367
R769 B.n232 B.n205 163.367
R770 B.n236 B.n205 163.367
R771 B.n237 B.n236 163.367
R772 B.n238 B.n237 163.367
R773 B.n238 B.n203 163.367
R774 B.n242 B.n203 163.367
R775 B.n243 B.n242 163.367
R776 B.n244 B.n243 163.367
R777 B.n244 B.n201 163.367
R778 B.n248 B.n201 163.367
R779 B.n249 B.n248 163.367
R780 B.n250 B.n249 163.367
R781 B.n250 B.n199 163.367
R782 B.n254 B.n199 163.367
R783 B.n255 B.n254 163.367
R784 B.n256 B.n255 163.367
R785 B.n256 B.n197 163.367
R786 B.n260 B.n197 163.367
R787 B.n261 B.n260 163.367
R788 B.n262 B.n261 163.367
R789 B.n262 B.n195 163.367
R790 B.n266 B.n195 163.367
R791 B.n267 B.n266 163.367
R792 B.n268 B.n267 163.367
R793 B.n268 B.n193 163.367
R794 B.n272 B.n193 163.367
R795 B.n273 B.n272 163.367
R796 B.n274 B.n273 163.367
R797 B.n274 B.n191 163.367
R798 B.n278 B.n191 163.367
R799 B.n279 B.n278 163.367
R800 B.n280 B.n279 163.367
R801 B.n280 B.n189 163.367
R802 B.n284 B.n189 163.367
R803 B.n285 B.n284 163.367
R804 B.n286 B.n285 163.367
R805 B.n286 B.n187 163.367
R806 B.n290 B.n187 163.367
R807 B.n291 B.n290 163.367
R808 B.n292 B.n291 163.367
R809 B.n292 B.n185 163.367
R810 B.n296 B.n185 163.367
R811 B.n297 B.n296 163.367
R812 B.n298 B.n297 163.367
R813 B.n298 B.n183 163.367
R814 B.n302 B.n183 163.367
R815 B.n303 B.n302 163.367
R816 B.n304 B.n303 163.367
R817 B.n304 B.n181 163.367
R818 B.n308 B.n181 163.367
R819 B.n309 B.n308 163.367
R820 B.n310 B.n309 163.367
R821 B.n310 B.n179 163.367
R822 B.n165 B.n164 79.9035
R823 B.n157 B.n156 79.9035
R824 B.n59 B.n58 79.9035
R825 B.n51 B.n50 79.9035
R826 B.n355 B.n165 59.5399
R827 B.n158 B.n157 59.5399
R828 B.n661 B.n59 59.5399
R829 B.n52 B.n51 59.5399
R830 B.n719 B.n36 36.3712
R831 B.n619 B.n618 36.3712
R832 B.n413 B.n142 36.3712
R833 B.n313 B.n312 36.3712
R834 B B.n821 18.0485
R835 B.n720 B.n719 10.6151
R836 B.n721 B.n720 10.6151
R837 B.n721 B.n34 10.6151
R838 B.n725 B.n34 10.6151
R839 B.n726 B.n725 10.6151
R840 B.n727 B.n726 10.6151
R841 B.n727 B.n32 10.6151
R842 B.n731 B.n32 10.6151
R843 B.n732 B.n731 10.6151
R844 B.n733 B.n732 10.6151
R845 B.n733 B.n30 10.6151
R846 B.n737 B.n30 10.6151
R847 B.n738 B.n737 10.6151
R848 B.n739 B.n738 10.6151
R849 B.n739 B.n28 10.6151
R850 B.n743 B.n28 10.6151
R851 B.n744 B.n743 10.6151
R852 B.n745 B.n744 10.6151
R853 B.n745 B.n26 10.6151
R854 B.n749 B.n26 10.6151
R855 B.n750 B.n749 10.6151
R856 B.n751 B.n750 10.6151
R857 B.n751 B.n24 10.6151
R858 B.n755 B.n24 10.6151
R859 B.n756 B.n755 10.6151
R860 B.n757 B.n756 10.6151
R861 B.n757 B.n22 10.6151
R862 B.n761 B.n22 10.6151
R863 B.n762 B.n761 10.6151
R864 B.n763 B.n762 10.6151
R865 B.n763 B.n20 10.6151
R866 B.n767 B.n20 10.6151
R867 B.n768 B.n767 10.6151
R868 B.n769 B.n768 10.6151
R869 B.n769 B.n18 10.6151
R870 B.n773 B.n18 10.6151
R871 B.n774 B.n773 10.6151
R872 B.n775 B.n774 10.6151
R873 B.n775 B.n16 10.6151
R874 B.n779 B.n16 10.6151
R875 B.n780 B.n779 10.6151
R876 B.n781 B.n780 10.6151
R877 B.n781 B.n14 10.6151
R878 B.n785 B.n14 10.6151
R879 B.n786 B.n785 10.6151
R880 B.n787 B.n786 10.6151
R881 B.n787 B.n12 10.6151
R882 B.n791 B.n12 10.6151
R883 B.n792 B.n791 10.6151
R884 B.n793 B.n792 10.6151
R885 B.n793 B.n10 10.6151
R886 B.n797 B.n10 10.6151
R887 B.n798 B.n797 10.6151
R888 B.n799 B.n798 10.6151
R889 B.n799 B.n8 10.6151
R890 B.n803 B.n8 10.6151
R891 B.n804 B.n803 10.6151
R892 B.n805 B.n804 10.6151
R893 B.n805 B.n6 10.6151
R894 B.n809 B.n6 10.6151
R895 B.n810 B.n809 10.6151
R896 B.n811 B.n810 10.6151
R897 B.n811 B.n4 10.6151
R898 B.n815 B.n4 10.6151
R899 B.n816 B.n815 10.6151
R900 B.n817 B.n816 10.6151
R901 B.n817 B.n0 10.6151
R902 B.n715 B.n36 10.6151
R903 B.n715 B.n714 10.6151
R904 B.n714 B.n713 10.6151
R905 B.n713 B.n38 10.6151
R906 B.n709 B.n38 10.6151
R907 B.n709 B.n708 10.6151
R908 B.n708 B.n707 10.6151
R909 B.n707 B.n40 10.6151
R910 B.n703 B.n40 10.6151
R911 B.n703 B.n702 10.6151
R912 B.n702 B.n701 10.6151
R913 B.n701 B.n42 10.6151
R914 B.n697 B.n42 10.6151
R915 B.n697 B.n696 10.6151
R916 B.n696 B.n695 10.6151
R917 B.n695 B.n44 10.6151
R918 B.n691 B.n44 10.6151
R919 B.n691 B.n690 10.6151
R920 B.n690 B.n689 10.6151
R921 B.n689 B.n46 10.6151
R922 B.n685 B.n46 10.6151
R923 B.n685 B.n684 10.6151
R924 B.n684 B.n683 10.6151
R925 B.n683 B.n48 10.6151
R926 B.n679 B.n48 10.6151
R927 B.n679 B.n678 10.6151
R928 B.n678 B.n677 10.6151
R929 B.n674 B.n673 10.6151
R930 B.n673 B.n672 10.6151
R931 B.n672 B.n54 10.6151
R932 B.n668 B.n54 10.6151
R933 B.n668 B.n667 10.6151
R934 B.n667 B.n666 10.6151
R935 B.n666 B.n56 10.6151
R936 B.n662 B.n56 10.6151
R937 B.n660 B.n659 10.6151
R938 B.n659 B.n60 10.6151
R939 B.n655 B.n60 10.6151
R940 B.n655 B.n654 10.6151
R941 B.n654 B.n653 10.6151
R942 B.n653 B.n62 10.6151
R943 B.n649 B.n62 10.6151
R944 B.n649 B.n648 10.6151
R945 B.n648 B.n647 10.6151
R946 B.n647 B.n64 10.6151
R947 B.n643 B.n64 10.6151
R948 B.n643 B.n642 10.6151
R949 B.n642 B.n641 10.6151
R950 B.n641 B.n66 10.6151
R951 B.n637 B.n66 10.6151
R952 B.n637 B.n636 10.6151
R953 B.n636 B.n635 10.6151
R954 B.n635 B.n68 10.6151
R955 B.n631 B.n68 10.6151
R956 B.n631 B.n630 10.6151
R957 B.n630 B.n629 10.6151
R958 B.n629 B.n70 10.6151
R959 B.n625 B.n70 10.6151
R960 B.n625 B.n624 10.6151
R961 B.n624 B.n623 10.6151
R962 B.n623 B.n72 10.6151
R963 B.n619 B.n72 10.6151
R964 B.n618 B.n617 10.6151
R965 B.n617 B.n74 10.6151
R966 B.n613 B.n74 10.6151
R967 B.n613 B.n612 10.6151
R968 B.n612 B.n611 10.6151
R969 B.n611 B.n76 10.6151
R970 B.n607 B.n76 10.6151
R971 B.n607 B.n606 10.6151
R972 B.n606 B.n605 10.6151
R973 B.n605 B.n78 10.6151
R974 B.n601 B.n78 10.6151
R975 B.n601 B.n600 10.6151
R976 B.n600 B.n599 10.6151
R977 B.n599 B.n80 10.6151
R978 B.n595 B.n80 10.6151
R979 B.n595 B.n594 10.6151
R980 B.n594 B.n593 10.6151
R981 B.n593 B.n82 10.6151
R982 B.n589 B.n82 10.6151
R983 B.n589 B.n588 10.6151
R984 B.n588 B.n587 10.6151
R985 B.n587 B.n84 10.6151
R986 B.n583 B.n84 10.6151
R987 B.n583 B.n582 10.6151
R988 B.n582 B.n581 10.6151
R989 B.n581 B.n86 10.6151
R990 B.n577 B.n86 10.6151
R991 B.n577 B.n576 10.6151
R992 B.n576 B.n575 10.6151
R993 B.n575 B.n88 10.6151
R994 B.n571 B.n88 10.6151
R995 B.n571 B.n570 10.6151
R996 B.n570 B.n569 10.6151
R997 B.n569 B.n90 10.6151
R998 B.n565 B.n90 10.6151
R999 B.n565 B.n564 10.6151
R1000 B.n564 B.n563 10.6151
R1001 B.n563 B.n92 10.6151
R1002 B.n559 B.n92 10.6151
R1003 B.n559 B.n558 10.6151
R1004 B.n558 B.n557 10.6151
R1005 B.n557 B.n94 10.6151
R1006 B.n553 B.n94 10.6151
R1007 B.n553 B.n552 10.6151
R1008 B.n552 B.n551 10.6151
R1009 B.n551 B.n96 10.6151
R1010 B.n547 B.n96 10.6151
R1011 B.n547 B.n546 10.6151
R1012 B.n546 B.n545 10.6151
R1013 B.n545 B.n98 10.6151
R1014 B.n541 B.n98 10.6151
R1015 B.n541 B.n540 10.6151
R1016 B.n540 B.n539 10.6151
R1017 B.n539 B.n100 10.6151
R1018 B.n535 B.n100 10.6151
R1019 B.n535 B.n534 10.6151
R1020 B.n534 B.n533 10.6151
R1021 B.n533 B.n102 10.6151
R1022 B.n529 B.n102 10.6151
R1023 B.n529 B.n528 10.6151
R1024 B.n528 B.n527 10.6151
R1025 B.n527 B.n104 10.6151
R1026 B.n523 B.n104 10.6151
R1027 B.n523 B.n522 10.6151
R1028 B.n522 B.n521 10.6151
R1029 B.n521 B.n106 10.6151
R1030 B.n517 B.n106 10.6151
R1031 B.n517 B.n516 10.6151
R1032 B.n516 B.n515 10.6151
R1033 B.n515 B.n108 10.6151
R1034 B.n511 B.n108 10.6151
R1035 B.n511 B.n510 10.6151
R1036 B.n510 B.n509 10.6151
R1037 B.n509 B.n110 10.6151
R1038 B.n505 B.n110 10.6151
R1039 B.n505 B.n504 10.6151
R1040 B.n504 B.n503 10.6151
R1041 B.n503 B.n112 10.6151
R1042 B.n499 B.n112 10.6151
R1043 B.n499 B.n498 10.6151
R1044 B.n498 B.n497 10.6151
R1045 B.n497 B.n114 10.6151
R1046 B.n493 B.n114 10.6151
R1047 B.n493 B.n492 10.6151
R1048 B.n492 B.n491 10.6151
R1049 B.n491 B.n116 10.6151
R1050 B.n487 B.n116 10.6151
R1051 B.n487 B.n486 10.6151
R1052 B.n486 B.n485 10.6151
R1053 B.n485 B.n118 10.6151
R1054 B.n481 B.n118 10.6151
R1055 B.n481 B.n480 10.6151
R1056 B.n480 B.n479 10.6151
R1057 B.n479 B.n120 10.6151
R1058 B.n475 B.n120 10.6151
R1059 B.n475 B.n474 10.6151
R1060 B.n474 B.n473 10.6151
R1061 B.n473 B.n122 10.6151
R1062 B.n469 B.n122 10.6151
R1063 B.n469 B.n468 10.6151
R1064 B.n468 B.n467 10.6151
R1065 B.n467 B.n124 10.6151
R1066 B.n463 B.n124 10.6151
R1067 B.n463 B.n462 10.6151
R1068 B.n462 B.n461 10.6151
R1069 B.n461 B.n126 10.6151
R1070 B.n457 B.n126 10.6151
R1071 B.n457 B.n456 10.6151
R1072 B.n456 B.n455 10.6151
R1073 B.n455 B.n128 10.6151
R1074 B.n451 B.n128 10.6151
R1075 B.n451 B.n450 10.6151
R1076 B.n450 B.n449 10.6151
R1077 B.n449 B.n130 10.6151
R1078 B.n445 B.n130 10.6151
R1079 B.n445 B.n444 10.6151
R1080 B.n444 B.n443 10.6151
R1081 B.n443 B.n132 10.6151
R1082 B.n439 B.n132 10.6151
R1083 B.n439 B.n438 10.6151
R1084 B.n438 B.n437 10.6151
R1085 B.n437 B.n134 10.6151
R1086 B.n433 B.n134 10.6151
R1087 B.n433 B.n432 10.6151
R1088 B.n432 B.n431 10.6151
R1089 B.n431 B.n136 10.6151
R1090 B.n427 B.n136 10.6151
R1091 B.n427 B.n426 10.6151
R1092 B.n426 B.n425 10.6151
R1093 B.n425 B.n138 10.6151
R1094 B.n421 B.n138 10.6151
R1095 B.n421 B.n420 10.6151
R1096 B.n420 B.n419 10.6151
R1097 B.n419 B.n140 10.6151
R1098 B.n415 B.n140 10.6151
R1099 B.n415 B.n414 10.6151
R1100 B.n414 B.n413 10.6151
R1101 B.n212 B.n1 10.6151
R1102 B.n215 B.n212 10.6151
R1103 B.n216 B.n215 10.6151
R1104 B.n217 B.n216 10.6151
R1105 B.n217 B.n210 10.6151
R1106 B.n221 B.n210 10.6151
R1107 B.n222 B.n221 10.6151
R1108 B.n223 B.n222 10.6151
R1109 B.n223 B.n208 10.6151
R1110 B.n227 B.n208 10.6151
R1111 B.n228 B.n227 10.6151
R1112 B.n229 B.n228 10.6151
R1113 B.n229 B.n206 10.6151
R1114 B.n233 B.n206 10.6151
R1115 B.n234 B.n233 10.6151
R1116 B.n235 B.n234 10.6151
R1117 B.n235 B.n204 10.6151
R1118 B.n239 B.n204 10.6151
R1119 B.n240 B.n239 10.6151
R1120 B.n241 B.n240 10.6151
R1121 B.n241 B.n202 10.6151
R1122 B.n245 B.n202 10.6151
R1123 B.n246 B.n245 10.6151
R1124 B.n247 B.n246 10.6151
R1125 B.n247 B.n200 10.6151
R1126 B.n251 B.n200 10.6151
R1127 B.n252 B.n251 10.6151
R1128 B.n253 B.n252 10.6151
R1129 B.n253 B.n198 10.6151
R1130 B.n257 B.n198 10.6151
R1131 B.n258 B.n257 10.6151
R1132 B.n259 B.n258 10.6151
R1133 B.n259 B.n196 10.6151
R1134 B.n263 B.n196 10.6151
R1135 B.n264 B.n263 10.6151
R1136 B.n265 B.n264 10.6151
R1137 B.n265 B.n194 10.6151
R1138 B.n269 B.n194 10.6151
R1139 B.n270 B.n269 10.6151
R1140 B.n271 B.n270 10.6151
R1141 B.n271 B.n192 10.6151
R1142 B.n275 B.n192 10.6151
R1143 B.n276 B.n275 10.6151
R1144 B.n277 B.n276 10.6151
R1145 B.n277 B.n190 10.6151
R1146 B.n281 B.n190 10.6151
R1147 B.n282 B.n281 10.6151
R1148 B.n283 B.n282 10.6151
R1149 B.n283 B.n188 10.6151
R1150 B.n287 B.n188 10.6151
R1151 B.n288 B.n287 10.6151
R1152 B.n289 B.n288 10.6151
R1153 B.n289 B.n186 10.6151
R1154 B.n293 B.n186 10.6151
R1155 B.n294 B.n293 10.6151
R1156 B.n295 B.n294 10.6151
R1157 B.n295 B.n184 10.6151
R1158 B.n299 B.n184 10.6151
R1159 B.n300 B.n299 10.6151
R1160 B.n301 B.n300 10.6151
R1161 B.n301 B.n182 10.6151
R1162 B.n305 B.n182 10.6151
R1163 B.n306 B.n305 10.6151
R1164 B.n307 B.n306 10.6151
R1165 B.n307 B.n180 10.6151
R1166 B.n311 B.n180 10.6151
R1167 B.n312 B.n311 10.6151
R1168 B.n313 B.n178 10.6151
R1169 B.n317 B.n178 10.6151
R1170 B.n318 B.n317 10.6151
R1171 B.n319 B.n318 10.6151
R1172 B.n319 B.n176 10.6151
R1173 B.n323 B.n176 10.6151
R1174 B.n324 B.n323 10.6151
R1175 B.n325 B.n324 10.6151
R1176 B.n325 B.n174 10.6151
R1177 B.n329 B.n174 10.6151
R1178 B.n330 B.n329 10.6151
R1179 B.n331 B.n330 10.6151
R1180 B.n331 B.n172 10.6151
R1181 B.n335 B.n172 10.6151
R1182 B.n336 B.n335 10.6151
R1183 B.n337 B.n336 10.6151
R1184 B.n337 B.n170 10.6151
R1185 B.n341 B.n170 10.6151
R1186 B.n342 B.n341 10.6151
R1187 B.n343 B.n342 10.6151
R1188 B.n343 B.n168 10.6151
R1189 B.n347 B.n168 10.6151
R1190 B.n348 B.n347 10.6151
R1191 B.n349 B.n348 10.6151
R1192 B.n349 B.n166 10.6151
R1193 B.n353 B.n166 10.6151
R1194 B.n354 B.n353 10.6151
R1195 B.n356 B.n162 10.6151
R1196 B.n360 B.n162 10.6151
R1197 B.n361 B.n360 10.6151
R1198 B.n362 B.n361 10.6151
R1199 B.n362 B.n160 10.6151
R1200 B.n366 B.n160 10.6151
R1201 B.n367 B.n366 10.6151
R1202 B.n368 B.n367 10.6151
R1203 B.n372 B.n371 10.6151
R1204 B.n373 B.n372 10.6151
R1205 B.n373 B.n154 10.6151
R1206 B.n377 B.n154 10.6151
R1207 B.n378 B.n377 10.6151
R1208 B.n379 B.n378 10.6151
R1209 B.n379 B.n152 10.6151
R1210 B.n383 B.n152 10.6151
R1211 B.n384 B.n383 10.6151
R1212 B.n385 B.n384 10.6151
R1213 B.n385 B.n150 10.6151
R1214 B.n389 B.n150 10.6151
R1215 B.n390 B.n389 10.6151
R1216 B.n391 B.n390 10.6151
R1217 B.n391 B.n148 10.6151
R1218 B.n395 B.n148 10.6151
R1219 B.n396 B.n395 10.6151
R1220 B.n397 B.n396 10.6151
R1221 B.n397 B.n146 10.6151
R1222 B.n401 B.n146 10.6151
R1223 B.n402 B.n401 10.6151
R1224 B.n403 B.n402 10.6151
R1225 B.n403 B.n144 10.6151
R1226 B.n407 B.n144 10.6151
R1227 B.n408 B.n407 10.6151
R1228 B.n409 B.n408 10.6151
R1229 B.n409 B.n142 10.6151
R1230 B.n821 B.n0 8.11757
R1231 B.n821 B.n1 8.11757
R1232 B.n674 B.n52 6.5566
R1233 B.n662 B.n661 6.5566
R1234 B.n356 B.n355 6.5566
R1235 B.n368 B.n158 6.5566
R1236 B.n677 B.n52 4.05904
R1237 B.n661 B.n660 4.05904
R1238 B.n355 B.n354 4.05904
R1239 B.n371 B.n158 4.05904
R1240 VN.n71 VN.n37 161.3
R1241 VN.n70 VN.n69 161.3
R1242 VN.n68 VN.n38 161.3
R1243 VN.n67 VN.n66 161.3
R1244 VN.n65 VN.n39 161.3
R1245 VN.n64 VN.n63 161.3
R1246 VN.n62 VN.n40 161.3
R1247 VN.n61 VN.n60 161.3
R1248 VN.n58 VN.n41 161.3
R1249 VN.n57 VN.n56 161.3
R1250 VN.n55 VN.n42 161.3
R1251 VN.n54 VN.n53 161.3
R1252 VN.n52 VN.n43 161.3
R1253 VN.n51 VN.n50 161.3
R1254 VN.n49 VN.n44 161.3
R1255 VN.n48 VN.n47 161.3
R1256 VN.n34 VN.n0 161.3
R1257 VN.n33 VN.n32 161.3
R1258 VN.n31 VN.n1 161.3
R1259 VN.n30 VN.n29 161.3
R1260 VN.n28 VN.n2 161.3
R1261 VN.n27 VN.n26 161.3
R1262 VN.n25 VN.n3 161.3
R1263 VN.n24 VN.n23 161.3
R1264 VN.n21 VN.n4 161.3
R1265 VN.n20 VN.n19 161.3
R1266 VN.n18 VN.n5 161.3
R1267 VN.n17 VN.n16 161.3
R1268 VN.n15 VN.n6 161.3
R1269 VN.n14 VN.n13 161.3
R1270 VN.n12 VN.n7 161.3
R1271 VN.n11 VN.n10 161.3
R1272 VN.n8 VN.t0 78.877
R1273 VN.n45 VN.t5 78.877
R1274 VN.n36 VN.n35 61.1402
R1275 VN.n73 VN.n72 61.1402
R1276 VN.n9 VN.n8 59.8758
R1277 VN.n46 VN.n45 59.8758
R1278 VN.n16 VN.n15 56.5193
R1279 VN.n53 VN.n52 56.5193
R1280 VN VN.n73 53.1708
R1281 VN.n29 VN.n28 53.1199
R1282 VN.n66 VN.n65 53.1199
R1283 VN.n9 VN.t6 46.6108
R1284 VN.n22 VN.t2 46.6108
R1285 VN.n35 VN.t4 46.6108
R1286 VN.n46 VN.t3 46.6108
R1287 VN.n59 VN.t1 46.6108
R1288 VN.n72 VN.t7 46.6108
R1289 VN.n29 VN.n1 27.8669
R1290 VN.n66 VN.n38 27.8669
R1291 VN.n10 VN.n7 24.4675
R1292 VN.n14 VN.n7 24.4675
R1293 VN.n15 VN.n14 24.4675
R1294 VN.n16 VN.n5 24.4675
R1295 VN.n20 VN.n5 24.4675
R1296 VN.n21 VN.n20 24.4675
R1297 VN.n23 VN.n3 24.4675
R1298 VN.n27 VN.n3 24.4675
R1299 VN.n28 VN.n27 24.4675
R1300 VN.n33 VN.n1 24.4675
R1301 VN.n34 VN.n33 24.4675
R1302 VN.n52 VN.n51 24.4675
R1303 VN.n51 VN.n44 24.4675
R1304 VN.n47 VN.n44 24.4675
R1305 VN.n65 VN.n64 24.4675
R1306 VN.n64 VN.n40 24.4675
R1307 VN.n60 VN.n40 24.4675
R1308 VN.n58 VN.n57 24.4675
R1309 VN.n57 VN.n42 24.4675
R1310 VN.n53 VN.n42 24.4675
R1311 VN.n71 VN.n70 24.4675
R1312 VN.n70 VN.n38 24.4675
R1313 VN.n35 VN.n34 21.0421
R1314 VN.n72 VN.n71 21.0421
R1315 VN.n10 VN.n9 15.17
R1316 VN.n22 VN.n21 15.17
R1317 VN.n47 VN.n46 15.17
R1318 VN.n59 VN.n58 15.17
R1319 VN.n23 VN.n22 9.29796
R1320 VN.n60 VN.n59 9.29796
R1321 VN.n48 VN.n45 2.65259
R1322 VN.n11 VN.n8 2.65259
R1323 VN.n73 VN.n37 0.417535
R1324 VN.n36 VN.n0 0.417535
R1325 VN VN.n36 0.394291
R1326 VN.n69 VN.n37 0.189894
R1327 VN.n69 VN.n68 0.189894
R1328 VN.n68 VN.n67 0.189894
R1329 VN.n67 VN.n39 0.189894
R1330 VN.n63 VN.n39 0.189894
R1331 VN.n63 VN.n62 0.189894
R1332 VN.n62 VN.n61 0.189894
R1333 VN.n61 VN.n41 0.189894
R1334 VN.n56 VN.n41 0.189894
R1335 VN.n56 VN.n55 0.189894
R1336 VN.n55 VN.n54 0.189894
R1337 VN.n54 VN.n43 0.189894
R1338 VN.n50 VN.n43 0.189894
R1339 VN.n50 VN.n49 0.189894
R1340 VN.n49 VN.n48 0.189894
R1341 VN.n12 VN.n11 0.189894
R1342 VN.n13 VN.n12 0.189894
R1343 VN.n13 VN.n6 0.189894
R1344 VN.n17 VN.n6 0.189894
R1345 VN.n18 VN.n17 0.189894
R1346 VN.n19 VN.n18 0.189894
R1347 VN.n19 VN.n4 0.189894
R1348 VN.n24 VN.n4 0.189894
R1349 VN.n25 VN.n24 0.189894
R1350 VN.n26 VN.n25 0.189894
R1351 VN.n26 VN.n2 0.189894
R1352 VN.n30 VN.n2 0.189894
R1353 VN.n31 VN.n30 0.189894
R1354 VN.n32 VN.n31 0.189894
R1355 VN.n32 VN.n0 0.189894
R1356 VDD2.n2 VDD2.n1 84.8895
R1357 VDD2.n2 VDD2.n0 84.8895
R1358 VDD2 VDD2.n5 84.8867
R1359 VDD2.n4 VDD2.n3 83.1692
R1360 VDD2.n4 VDD2.n2 46.017
R1361 VDD2.n5 VDD2.t3 4.43502
R1362 VDD2.n5 VDD2.t5 4.43502
R1363 VDD2.n3 VDD2.t7 4.43502
R1364 VDD2.n3 VDD2.t1 4.43502
R1365 VDD2.n1 VDD2.t2 4.43502
R1366 VDD2.n1 VDD2.t4 4.43502
R1367 VDD2.n0 VDD2.t0 4.43502
R1368 VDD2.n0 VDD2.t6 4.43502
R1369 VDD2 VDD2.n4 1.83455
R1370 VTAIL.n322 VTAIL.n288 756.745
R1371 VTAIL.n36 VTAIL.n2 756.745
R1372 VTAIL.n76 VTAIL.n42 756.745
R1373 VTAIL.n118 VTAIL.n84 756.745
R1374 VTAIL.n282 VTAIL.n248 756.745
R1375 VTAIL.n240 VTAIL.n206 756.745
R1376 VTAIL.n200 VTAIL.n166 756.745
R1377 VTAIL.n158 VTAIL.n124 756.745
R1378 VTAIL.n300 VTAIL.n299 585
R1379 VTAIL.n305 VTAIL.n304 585
R1380 VTAIL.n307 VTAIL.n306 585
R1381 VTAIL.n296 VTAIL.n295 585
R1382 VTAIL.n313 VTAIL.n312 585
R1383 VTAIL.n315 VTAIL.n314 585
R1384 VTAIL.n292 VTAIL.n291 585
R1385 VTAIL.n321 VTAIL.n320 585
R1386 VTAIL.n323 VTAIL.n322 585
R1387 VTAIL.n14 VTAIL.n13 585
R1388 VTAIL.n19 VTAIL.n18 585
R1389 VTAIL.n21 VTAIL.n20 585
R1390 VTAIL.n10 VTAIL.n9 585
R1391 VTAIL.n27 VTAIL.n26 585
R1392 VTAIL.n29 VTAIL.n28 585
R1393 VTAIL.n6 VTAIL.n5 585
R1394 VTAIL.n35 VTAIL.n34 585
R1395 VTAIL.n37 VTAIL.n36 585
R1396 VTAIL.n54 VTAIL.n53 585
R1397 VTAIL.n59 VTAIL.n58 585
R1398 VTAIL.n61 VTAIL.n60 585
R1399 VTAIL.n50 VTAIL.n49 585
R1400 VTAIL.n67 VTAIL.n66 585
R1401 VTAIL.n69 VTAIL.n68 585
R1402 VTAIL.n46 VTAIL.n45 585
R1403 VTAIL.n75 VTAIL.n74 585
R1404 VTAIL.n77 VTAIL.n76 585
R1405 VTAIL.n96 VTAIL.n95 585
R1406 VTAIL.n101 VTAIL.n100 585
R1407 VTAIL.n103 VTAIL.n102 585
R1408 VTAIL.n92 VTAIL.n91 585
R1409 VTAIL.n109 VTAIL.n108 585
R1410 VTAIL.n111 VTAIL.n110 585
R1411 VTAIL.n88 VTAIL.n87 585
R1412 VTAIL.n117 VTAIL.n116 585
R1413 VTAIL.n119 VTAIL.n118 585
R1414 VTAIL.n283 VTAIL.n282 585
R1415 VTAIL.n281 VTAIL.n280 585
R1416 VTAIL.n252 VTAIL.n251 585
R1417 VTAIL.n275 VTAIL.n274 585
R1418 VTAIL.n273 VTAIL.n272 585
R1419 VTAIL.n256 VTAIL.n255 585
R1420 VTAIL.n267 VTAIL.n266 585
R1421 VTAIL.n265 VTAIL.n264 585
R1422 VTAIL.n260 VTAIL.n259 585
R1423 VTAIL.n241 VTAIL.n240 585
R1424 VTAIL.n239 VTAIL.n238 585
R1425 VTAIL.n210 VTAIL.n209 585
R1426 VTAIL.n233 VTAIL.n232 585
R1427 VTAIL.n231 VTAIL.n230 585
R1428 VTAIL.n214 VTAIL.n213 585
R1429 VTAIL.n225 VTAIL.n224 585
R1430 VTAIL.n223 VTAIL.n222 585
R1431 VTAIL.n218 VTAIL.n217 585
R1432 VTAIL.n201 VTAIL.n200 585
R1433 VTAIL.n199 VTAIL.n198 585
R1434 VTAIL.n170 VTAIL.n169 585
R1435 VTAIL.n193 VTAIL.n192 585
R1436 VTAIL.n191 VTAIL.n190 585
R1437 VTAIL.n174 VTAIL.n173 585
R1438 VTAIL.n185 VTAIL.n184 585
R1439 VTAIL.n183 VTAIL.n182 585
R1440 VTAIL.n178 VTAIL.n177 585
R1441 VTAIL.n159 VTAIL.n158 585
R1442 VTAIL.n157 VTAIL.n156 585
R1443 VTAIL.n128 VTAIL.n127 585
R1444 VTAIL.n151 VTAIL.n150 585
R1445 VTAIL.n149 VTAIL.n148 585
R1446 VTAIL.n132 VTAIL.n131 585
R1447 VTAIL.n143 VTAIL.n142 585
R1448 VTAIL.n141 VTAIL.n140 585
R1449 VTAIL.n136 VTAIL.n135 585
R1450 VTAIL.n301 VTAIL.t11 327.483
R1451 VTAIL.n15 VTAIL.t15 327.483
R1452 VTAIL.n55 VTAIL.t2 327.483
R1453 VTAIL.n97 VTAIL.t3 327.483
R1454 VTAIL.n261 VTAIL.t0 327.483
R1455 VTAIL.n219 VTAIL.t5 327.483
R1456 VTAIL.n179 VTAIL.t10 327.483
R1457 VTAIL.n137 VTAIL.t8 327.483
R1458 VTAIL.n305 VTAIL.n299 171.744
R1459 VTAIL.n306 VTAIL.n305 171.744
R1460 VTAIL.n306 VTAIL.n295 171.744
R1461 VTAIL.n313 VTAIL.n295 171.744
R1462 VTAIL.n314 VTAIL.n313 171.744
R1463 VTAIL.n314 VTAIL.n291 171.744
R1464 VTAIL.n321 VTAIL.n291 171.744
R1465 VTAIL.n322 VTAIL.n321 171.744
R1466 VTAIL.n19 VTAIL.n13 171.744
R1467 VTAIL.n20 VTAIL.n19 171.744
R1468 VTAIL.n20 VTAIL.n9 171.744
R1469 VTAIL.n27 VTAIL.n9 171.744
R1470 VTAIL.n28 VTAIL.n27 171.744
R1471 VTAIL.n28 VTAIL.n5 171.744
R1472 VTAIL.n35 VTAIL.n5 171.744
R1473 VTAIL.n36 VTAIL.n35 171.744
R1474 VTAIL.n59 VTAIL.n53 171.744
R1475 VTAIL.n60 VTAIL.n59 171.744
R1476 VTAIL.n60 VTAIL.n49 171.744
R1477 VTAIL.n67 VTAIL.n49 171.744
R1478 VTAIL.n68 VTAIL.n67 171.744
R1479 VTAIL.n68 VTAIL.n45 171.744
R1480 VTAIL.n75 VTAIL.n45 171.744
R1481 VTAIL.n76 VTAIL.n75 171.744
R1482 VTAIL.n101 VTAIL.n95 171.744
R1483 VTAIL.n102 VTAIL.n101 171.744
R1484 VTAIL.n102 VTAIL.n91 171.744
R1485 VTAIL.n109 VTAIL.n91 171.744
R1486 VTAIL.n110 VTAIL.n109 171.744
R1487 VTAIL.n110 VTAIL.n87 171.744
R1488 VTAIL.n117 VTAIL.n87 171.744
R1489 VTAIL.n118 VTAIL.n117 171.744
R1490 VTAIL.n282 VTAIL.n281 171.744
R1491 VTAIL.n281 VTAIL.n251 171.744
R1492 VTAIL.n274 VTAIL.n251 171.744
R1493 VTAIL.n274 VTAIL.n273 171.744
R1494 VTAIL.n273 VTAIL.n255 171.744
R1495 VTAIL.n266 VTAIL.n255 171.744
R1496 VTAIL.n266 VTAIL.n265 171.744
R1497 VTAIL.n265 VTAIL.n259 171.744
R1498 VTAIL.n240 VTAIL.n239 171.744
R1499 VTAIL.n239 VTAIL.n209 171.744
R1500 VTAIL.n232 VTAIL.n209 171.744
R1501 VTAIL.n232 VTAIL.n231 171.744
R1502 VTAIL.n231 VTAIL.n213 171.744
R1503 VTAIL.n224 VTAIL.n213 171.744
R1504 VTAIL.n224 VTAIL.n223 171.744
R1505 VTAIL.n223 VTAIL.n217 171.744
R1506 VTAIL.n200 VTAIL.n199 171.744
R1507 VTAIL.n199 VTAIL.n169 171.744
R1508 VTAIL.n192 VTAIL.n169 171.744
R1509 VTAIL.n192 VTAIL.n191 171.744
R1510 VTAIL.n191 VTAIL.n173 171.744
R1511 VTAIL.n184 VTAIL.n173 171.744
R1512 VTAIL.n184 VTAIL.n183 171.744
R1513 VTAIL.n183 VTAIL.n177 171.744
R1514 VTAIL.n158 VTAIL.n157 171.744
R1515 VTAIL.n157 VTAIL.n127 171.744
R1516 VTAIL.n150 VTAIL.n127 171.744
R1517 VTAIL.n150 VTAIL.n149 171.744
R1518 VTAIL.n149 VTAIL.n131 171.744
R1519 VTAIL.n142 VTAIL.n131 171.744
R1520 VTAIL.n142 VTAIL.n141 171.744
R1521 VTAIL.n141 VTAIL.n135 171.744
R1522 VTAIL.t11 VTAIL.n299 85.8723
R1523 VTAIL.t15 VTAIL.n13 85.8723
R1524 VTAIL.t2 VTAIL.n53 85.8723
R1525 VTAIL.t3 VTAIL.n95 85.8723
R1526 VTAIL.t0 VTAIL.n259 85.8723
R1527 VTAIL.t5 VTAIL.n217 85.8723
R1528 VTAIL.t10 VTAIL.n177 85.8723
R1529 VTAIL.t8 VTAIL.n135 85.8723
R1530 VTAIL.n247 VTAIL.n246 66.4904
R1531 VTAIL.n165 VTAIL.n164 66.4904
R1532 VTAIL.n1 VTAIL.n0 66.4902
R1533 VTAIL.n83 VTAIL.n82 66.4902
R1534 VTAIL.n327 VTAIL.n326 30.052
R1535 VTAIL.n41 VTAIL.n40 30.052
R1536 VTAIL.n81 VTAIL.n80 30.052
R1537 VTAIL.n123 VTAIL.n122 30.052
R1538 VTAIL.n287 VTAIL.n286 30.052
R1539 VTAIL.n245 VTAIL.n244 30.052
R1540 VTAIL.n205 VTAIL.n204 30.052
R1541 VTAIL.n163 VTAIL.n162 30.052
R1542 VTAIL.n327 VTAIL.n287 22.2376
R1543 VTAIL.n163 VTAIL.n123 22.2376
R1544 VTAIL.n301 VTAIL.n300 16.3891
R1545 VTAIL.n15 VTAIL.n14 16.3891
R1546 VTAIL.n55 VTAIL.n54 16.3891
R1547 VTAIL.n97 VTAIL.n96 16.3891
R1548 VTAIL.n261 VTAIL.n260 16.3891
R1549 VTAIL.n219 VTAIL.n218 16.3891
R1550 VTAIL.n179 VTAIL.n178 16.3891
R1551 VTAIL.n137 VTAIL.n136 16.3891
R1552 VTAIL.n304 VTAIL.n303 12.8005
R1553 VTAIL.n18 VTAIL.n17 12.8005
R1554 VTAIL.n58 VTAIL.n57 12.8005
R1555 VTAIL.n100 VTAIL.n99 12.8005
R1556 VTAIL.n264 VTAIL.n263 12.8005
R1557 VTAIL.n222 VTAIL.n221 12.8005
R1558 VTAIL.n182 VTAIL.n181 12.8005
R1559 VTAIL.n140 VTAIL.n139 12.8005
R1560 VTAIL.n307 VTAIL.n298 12.0247
R1561 VTAIL.n21 VTAIL.n12 12.0247
R1562 VTAIL.n61 VTAIL.n52 12.0247
R1563 VTAIL.n103 VTAIL.n94 12.0247
R1564 VTAIL.n267 VTAIL.n258 12.0247
R1565 VTAIL.n225 VTAIL.n216 12.0247
R1566 VTAIL.n185 VTAIL.n176 12.0247
R1567 VTAIL.n143 VTAIL.n134 12.0247
R1568 VTAIL.n308 VTAIL.n296 11.249
R1569 VTAIL.n22 VTAIL.n10 11.249
R1570 VTAIL.n62 VTAIL.n50 11.249
R1571 VTAIL.n104 VTAIL.n92 11.249
R1572 VTAIL.n268 VTAIL.n256 11.249
R1573 VTAIL.n226 VTAIL.n214 11.249
R1574 VTAIL.n186 VTAIL.n174 11.249
R1575 VTAIL.n144 VTAIL.n132 11.249
R1576 VTAIL.n312 VTAIL.n311 10.4732
R1577 VTAIL.n26 VTAIL.n25 10.4732
R1578 VTAIL.n66 VTAIL.n65 10.4732
R1579 VTAIL.n108 VTAIL.n107 10.4732
R1580 VTAIL.n272 VTAIL.n271 10.4732
R1581 VTAIL.n230 VTAIL.n229 10.4732
R1582 VTAIL.n190 VTAIL.n189 10.4732
R1583 VTAIL.n148 VTAIL.n147 10.4732
R1584 VTAIL.n315 VTAIL.n294 9.69747
R1585 VTAIL.n29 VTAIL.n8 9.69747
R1586 VTAIL.n69 VTAIL.n48 9.69747
R1587 VTAIL.n111 VTAIL.n90 9.69747
R1588 VTAIL.n275 VTAIL.n254 9.69747
R1589 VTAIL.n233 VTAIL.n212 9.69747
R1590 VTAIL.n193 VTAIL.n172 9.69747
R1591 VTAIL.n151 VTAIL.n130 9.69747
R1592 VTAIL.n326 VTAIL.n325 9.45567
R1593 VTAIL.n40 VTAIL.n39 9.45567
R1594 VTAIL.n80 VTAIL.n79 9.45567
R1595 VTAIL.n122 VTAIL.n121 9.45567
R1596 VTAIL.n286 VTAIL.n285 9.45567
R1597 VTAIL.n244 VTAIL.n243 9.45567
R1598 VTAIL.n204 VTAIL.n203 9.45567
R1599 VTAIL.n162 VTAIL.n161 9.45567
R1600 VTAIL.n325 VTAIL.n324 9.3005
R1601 VTAIL.n319 VTAIL.n318 9.3005
R1602 VTAIL.n317 VTAIL.n316 9.3005
R1603 VTAIL.n294 VTAIL.n293 9.3005
R1604 VTAIL.n311 VTAIL.n310 9.3005
R1605 VTAIL.n309 VTAIL.n308 9.3005
R1606 VTAIL.n298 VTAIL.n297 9.3005
R1607 VTAIL.n303 VTAIL.n302 9.3005
R1608 VTAIL.n290 VTAIL.n289 9.3005
R1609 VTAIL.n39 VTAIL.n38 9.3005
R1610 VTAIL.n33 VTAIL.n32 9.3005
R1611 VTAIL.n31 VTAIL.n30 9.3005
R1612 VTAIL.n8 VTAIL.n7 9.3005
R1613 VTAIL.n25 VTAIL.n24 9.3005
R1614 VTAIL.n23 VTAIL.n22 9.3005
R1615 VTAIL.n12 VTAIL.n11 9.3005
R1616 VTAIL.n17 VTAIL.n16 9.3005
R1617 VTAIL.n4 VTAIL.n3 9.3005
R1618 VTAIL.n79 VTAIL.n78 9.3005
R1619 VTAIL.n73 VTAIL.n72 9.3005
R1620 VTAIL.n71 VTAIL.n70 9.3005
R1621 VTAIL.n48 VTAIL.n47 9.3005
R1622 VTAIL.n65 VTAIL.n64 9.3005
R1623 VTAIL.n63 VTAIL.n62 9.3005
R1624 VTAIL.n52 VTAIL.n51 9.3005
R1625 VTAIL.n57 VTAIL.n56 9.3005
R1626 VTAIL.n44 VTAIL.n43 9.3005
R1627 VTAIL.n121 VTAIL.n120 9.3005
R1628 VTAIL.n115 VTAIL.n114 9.3005
R1629 VTAIL.n113 VTAIL.n112 9.3005
R1630 VTAIL.n90 VTAIL.n89 9.3005
R1631 VTAIL.n107 VTAIL.n106 9.3005
R1632 VTAIL.n105 VTAIL.n104 9.3005
R1633 VTAIL.n94 VTAIL.n93 9.3005
R1634 VTAIL.n99 VTAIL.n98 9.3005
R1635 VTAIL.n86 VTAIL.n85 9.3005
R1636 VTAIL.n285 VTAIL.n284 9.3005
R1637 VTAIL.n250 VTAIL.n249 9.3005
R1638 VTAIL.n279 VTAIL.n278 9.3005
R1639 VTAIL.n277 VTAIL.n276 9.3005
R1640 VTAIL.n254 VTAIL.n253 9.3005
R1641 VTAIL.n271 VTAIL.n270 9.3005
R1642 VTAIL.n269 VTAIL.n268 9.3005
R1643 VTAIL.n258 VTAIL.n257 9.3005
R1644 VTAIL.n263 VTAIL.n262 9.3005
R1645 VTAIL.n243 VTAIL.n242 9.3005
R1646 VTAIL.n208 VTAIL.n207 9.3005
R1647 VTAIL.n237 VTAIL.n236 9.3005
R1648 VTAIL.n235 VTAIL.n234 9.3005
R1649 VTAIL.n212 VTAIL.n211 9.3005
R1650 VTAIL.n229 VTAIL.n228 9.3005
R1651 VTAIL.n227 VTAIL.n226 9.3005
R1652 VTAIL.n216 VTAIL.n215 9.3005
R1653 VTAIL.n221 VTAIL.n220 9.3005
R1654 VTAIL.n203 VTAIL.n202 9.3005
R1655 VTAIL.n168 VTAIL.n167 9.3005
R1656 VTAIL.n197 VTAIL.n196 9.3005
R1657 VTAIL.n195 VTAIL.n194 9.3005
R1658 VTAIL.n172 VTAIL.n171 9.3005
R1659 VTAIL.n189 VTAIL.n188 9.3005
R1660 VTAIL.n187 VTAIL.n186 9.3005
R1661 VTAIL.n176 VTAIL.n175 9.3005
R1662 VTAIL.n181 VTAIL.n180 9.3005
R1663 VTAIL.n161 VTAIL.n160 9.3005
R1664 VTAIL.n126 VTAIL.n125 9.3005
R1665 VTAIL.n155 VTAIL.n154 9.3005
R1666 VTAIL.n153 VTAIL.n152 9.3005
R1667 VTAIL.n130 VTAIL.n129 9.3005
R1668 VTAIL.n147 VTAIL.n146 9.3005
R1669 VTAIL.n145 VTAIL.n144 9.3005
R1670 VTAIL.n134 VTAIL.n133 9.3005
R1671 VTAIL.n139 VTAIL.n138 9.3005
R1672 VTAIL.n316 VTAIL.n292 8.92171
R1673 VTAIL.n30 VTAIL.n6 8.92171
R1674 VTAIL.n70 VTAIL.n46 8.92171
R1675 VTAIL.n112 VTAIL.n88 8.92171
R1676 VTAIL.n276 VTAIL.n252 8.92171
R1677 VTAIL.n234 VTAIL.n210 8.92171
R1678 VTAIL.n194 VTAIL.n170 8.92171
R1679 VTAIL.n152 VTAIL.n128 8.92171
R1680 VTAIL.n320 VTAIL.n319 8.14595
R1681 VTAIL.n34 VTAIL.n33 8.14595
R1682 VTAIL.n74 VTAIL.n73 8.14595
R1683 VTAIL.n116 VTAIL.n115 8.14595
R1684 VTAIL.n280 VTAIL.n279 8.14595
R1685 VTAIL.n238 VTAIL.n237 8.14595
R1686 VTAIL.n198 VTAIL.n197 8.14595
R1687 VTAIL.n156 VTAIL.n155 8.14595
R1688 VTAIL.n323 VTAIL.n290 7.3702
R1689 VTAIL.n326 VTAIL.n288 7.3702
R1690 VTAIL.n37 VTAIL.n4 7.3702
R1691 VTAIL.n40 VTAIL.n2 7.3702
R1692 VTAIL.n77 VTAIL.n44 7.3702
R1693 VTAIL.n80 VTAIL.n42 7.3702
R1694 VTAIL.n119 VTAIL.n86 7.3702
R1695 VTAIL.n122 VTAIL.n84 7.3702
R1696 VTAIL.n286 VTAIL.n248 7.3702
R1697 VTAIL.n283 VTAIL.n250 7.3702
R1698 VTAIL.n244 VTAIL.n206 7.3702
R1699 VTAIL.n241 VTAIL.n208 7.3702
R1700 VTAIL.n204 VTAIL.n166 7.3702
R1701 VTAIL.n201 VTAIL.n168 7.3702
R1702 VTAIL.n162 VTAIL.n124 7.3702
R1703 VTAIL.n159 VTAIL.n126 7.3702
R1704 VTAIL.n324 VTAIL.n323 6.59444
R1705 VTAIL.n324 VTAIL.n288 6.59444
R1706 VTAIL.n38 VTAIL.n37 6.59444
R1707 VTAIL.n38 VTAIL.n2 6.59444
R1708 VTAIL.n78 VTAIL.n77 6.59444
R1709 VTAIL.n78 VTAIL.n42 6.59444
R1710 VTAIL.n120 VTAIL.n119 6.59444
R1711 VTAIL.n120 VTAIL.n84 6.59444
R1712 VTAIL.n284 VTAIL.n248 6.59444
R1713 VTAIL.n284 VTAIL.n283 6.59444
R1714 VTAIL.n242 VTAIL.n206 6.59444
R1715 VTAIL.n242 VTAIL.n241 6.59444
R1716 VTAIL.n202 VTAIL.n166 6.59444
R1717 VTAIL.n202 VTAIL.n201 6.59444
R1718 VTAIL.n160 VTAIL.n124 6.59444
R1719 VTAIL.n160 VTAIL.n159 6.59444
R1720 VTAIL.n320 VTAIL.n290 5.81868
R1721 VTAIL.n34 VTAIL.n4 5.81868
R1722 VTAIL.n74 VTAIL.n44 5.81868
R1723 VTAIL.n116 VTAIL.n86 5.81868
R1724 VTAIL.n280 VTAIL.n250 5.81868
R1725 VTAIL.n238 VTAIL.n208 5.81868
R1726 VTAIL.n198 VTAIL.n168 5.81868
R1727 VTAIL.n156 VTAIL.n126 5.81868
R1728 VTAIL.n319 VTAIL.n292 5.04292
R1729 VTAIL.n33 VTAIL.n6 5.04292
R1730 VTAIL.n73 VTAIL.n46 5.04292
R1731 VTAIL.n115 VTAIL.n88 5.04292
R1732 VTAIL.n279 VTAIL.n252 5.04292
R1733 VTAIL.n237 VTAIL.n210 5.04292
R1734 VTAIL.n197 VTAIL.n170 5.04292
R1735 VTAIL.n155 VTAIL.n128 5.04292
R1736 VTAIL.n0 VTAIL.t9 4.43502
R1737 VTAIL.n0 VTAIL.t13 4.43502
R1738 VTAIL.n82 VTAIL.t1 4.43502
R1739 VTAIL.n82 VTAIL.t4 4.43502
R1740 VTAIL.n246 VTAIL.t6 4.43502
R1741 VTAIL.n246 VTAIL.t7 4.43502
R1742 VTAIL.n164 VTAIL.t14 4.43502
R1743 VTAIL.n164 VTAIL.t12 4.43502
R1744 VTAIL.n316 VTAIL.n315 4.26717
R1745 VTAIL.n30 VTAIL.n29 4.26717
R1746 VTAIL.n70 VTAIL.n69 4.26717
R1747 VTAIL.n112 VTAIL.n111 4.26717
R1748 VTAIL.n276 VTAIL.n275 4.26717
R1749 VTAIL.n234 VTAIL.n233 4.26717
R1750 VTAIL.n194 VTAIL.n193 4.26717
R1751 VTAIL.n152 VTAIL.n151 4.26717
R1752 VTAIL.n302 VTAIL.n301 3.71019
R1753 VTAIL.n16 VTAIL.n15 3.71019
R1754 VTAIL.n56 VTAIL.n55 3.71019
R1755 VTAIL.n98 VTAIL.n97 3.71019
R1756 VTAIL.n262 VTAIL.n261 3.71019
R1757 VTAIL.n220 VTAIL.n219 3.71019
R1758 VTAIL.n180 VTAIL.n179 3.71019
R1759 VTAIL.n138 VTAIL.n137 3.71019
R1760 VTAIL.n165 VTAIL.n163 3.55222
R1761 VTAIL.n205 VTAIL.n165 3.55222
R1762 VTAIL.n247 VTAIL.n245 3.55222
R1763 VTAIL.n287 VTAIL.n247 3.55222
R1764 VTAIL.n123 VTAIL.n83 3.55222
R1765 VTAIL.n83 VTAIL.n81 3.55222
R1766 VTAIL.n41 VTAIL.n1 3.55222
R1767 VTAIL VTAIL.n327 3.49403
R1768 VTAIL.n312 VTAIL.n294 3.49141
R1769 VTAIL.n26 VTAIL.n8 3.49141
R1770 VTAIL.n66 VTAIL.n48 3.49141
R1771 VTAIL.n108 VTAIL.n90 3.49141
R1772 VTAIL.n272 VTAIL.n254 3.49141
R1773 VTAIL.n230 VTAIL.n212 3.49141
R1774 VTAIL.n190 VTAIL.n172 3.49141
R1775 VTAIL.n148 VTAIL.n130 3.49141
R1776 VTAIL.n311 VTAIL.n296 2.71565
R1777 VTAIL.n25 VTAIL.n10 2.71565
R1778 VTAIL.n65 VTAIL.n50 2.71565
R1779 VTAIL.n107 VTAIL.n92 2.71565
R1780 VTAIL.n271 VTAIL.n256 2.71565
R1781 VTAIL.n229 VTAIL.n214 2.71565
R1782 VTAIL.n189 VTAIL.n174 2.71565
R1783 VTAIL.n147 VTAIL.n132 2.71565
R1784 VTAIL.n308 VTAIL.n307 1.93989
R1785 VTAIL.n22 VTAIL.n21 1.93989
R1786 VTAIL.n62 VTAIL.n61 1.93989
R1787 VTAIL.n104 VTAIL.n103 1.93989
R1788 VTAIL.n268 VTAIL.n267 1.93989
R1789 VTAIL.n226 VTAIL.n225 1.93989
R1790 VTAIL.n186 VTAIL.n185 1.93989
R1791 VTAIL.n144 VTAIL.n143 1.93989
R1792 VTAIL.n304 VTAIL.n298 1.16414
R1793 VTAIL.n18 VTAIL.n12 1.16414
R1794 VTAIL.n58 VTAIL.n52 1.16414
R1795 VTAIL.n100 VTAIL.n94 1.16414
R1796 VTAIL.n264 VTAIL.n258 1.16414
R1797 VTAIL.n222 VTAIL.n216 1.16414
R1798 VTAIL.n182 VTAIL.n176 1.16414
R1799 VTAIL.n140 VTAIL.n134 1.16414
R1800 VTAIL.n245 VTAIL.n205 0.470328
R1801 VTAIL.n81 VTAIL.n41 0.470328
R1802 VTAIL.n303 VTAIL.n300 0.388379
R1803 VTAIL.n17 VTAIL.n14 0.388379
R1804 VTAIL.n57 VTAIL.n54 0.388379
R1805 VTAIL.n99 VTAIL.n96 0.388379
R1806 VTAIL.n263 VTAIL.n260 0.388379
R1807 VTAIL.n221 VTAIL.n218 0.388379
R1808 VTAIL.n181 VTAIL.n178 0.388379
R1809 VTAIL.n139 VTAIL.n136 0.388379
R1810 VTAIL.n302 VTAIL.n297 0.155672
R1811 VTAIL.n309 VTAIL.n297 0.155672
R1812 VTAIL.n310 VTAIL.n309 0.155672
R1813 VTAIL.n310 VTAIL.n293 0.155672
R1814 VTAIL.n317 VTAIL.n293 0.155672
R1815 VTAIL.n318 VTAIL.n317 0.155672
R1816 VTAIL.n318 VTAIL.n289 0.155672
R1817 VTAIL.n325 VTAIL.n289 0.155672
R1818 VTAIL.n16 VTAIL.n11 0.155672
R1819 VTAIL.n23 VTAIL.n11 0.155672
R1820 VTAIL.n24 VTAIL.n23 0.155672
R1821 VTAIL.n24 VTAIL.n7 0.155672
R1822 VTAIL.n31 VTAIL.n7 0.155672
R1823 VTAIL.n32 VTAIL.n31 0.155672
R1824 VTAIL.n32 VTAIL.n3 0.155672
R1825 VTAIL.n39 VTAIL.n3 0.155672
R1826 VTAIL.n56 VTAIL.n51 0.155672
R1827 VTAIL.n63 VTAIL.n51 0.155672
R1828 VTAIL.n64 VTAIL.n63 0.155672
R1829 VTAIL.n64 VTAIL.n47 0.155672
R1830 VTAIL.n71 VTAIL.n47 0.155672
R1831 VTAIL.n72 VTAIL.n71 0.155672
R1832 VTAIL.n72 VTAIL.n43 0.155672
R1833 VTAIL.n79 VTAIL.n43 0.155672
R1834 VTAIL.n98 VTAIL.n93 0.155672
R1835 VTAIL.n105 VTAIL.n93 0.155672
R1836 VTAIL.n106 VTAIL.n105 0.155672
R1837 VTAIL.n106 VTAIL.n89 0.155672
R1838 VTAIL.n113 VTAIL.n89 0.155672
R1839 VTAIL.n114 VTAIL.n113 0.155672
R1840 VTAIL.n114 VTAIL.n85 0.155672
R1841 VTAIL.n121 VTAIL.n85 0.155672
R1842 VTAIL.n285 VTAIL.n249 0.155672
R1843 VTAIL.n278 VTAIL.n249 0.155672
R1844 VTAIL.n278 VTAIL.n277 0.155672
R1845 VTAIL.n277 VTAIL.n253 0.155672
R1846 VTAIL.n270 VTAIL.n253 0.155672
R1847 VTAIL.n270 VTAIL.n269 0.155672
R1848 VTAIL.n269 VTAIL.n257 0.155672
R1849 VTAIL.n262 VTAIL.n257 0.155672
R1850 VTAIL.n243 VTAIL.n207 0.155672
R1851 VTAIL.n236 VTAIL.n207 0.155672
R1852 VTAIL.n236 VTAIL.n235 0.155672
R1853 VTAIL.n235 VTAIL.n211 0.155672
R1854 VTAIL.n228 VTAIL.n211 0.155672
R1855 VTAIL.n228 VTAIL.n227 0.155672
R1856 VTAIL.n227 VTAIL.n215 0.155672
R1857 VTAIL.n220 VTAIL.n215 0.155672
R1858 VTAIL.n203 VTAIL.n167 0.155672
R1859 VTAIL.n196 VTAIL.n167 0.155672
R1860 VTAIL.n196 VTAIL.n195 0.155672
R1861 VTAIL.n195 VTAIL.n171 0.155672
R1862 VTAIL.n188 VTAIL.n171 0.155672
R1863 VTAIL.n188 VTAIL.n187 0.155672
R1864 VTAIL.n187 VTAIL.n175 0.155672
R1865 VTAIL.n180 VTAIL.n175 0.155672
R1866 VTAIL.n161 VTAIL.n125 0.155672
R1867 VTAIL.n154 VTAIL.n125 0.155672
R1868 VTAIL.n154 VTAIL.n153 0.155672
R1869 VTAIL.n153 VTAIL.n129 0.155672
R1870 VTAIL.n146 VTAIL.n129 0.155672
R1871 VTAIL.n146 VTAIL.n145 0.155672
R1872 VTAIL.n145 VTAIL.n133 0.155672
R1873 VTAIL.n138 VTAIL.n133 0.155672
R1874 VTAIL VTAIL.n1 0.0586897
R1875 VP.n23 VP.n22 161.3
R1876 VP.n24 VP.n19 161.3
R1877 VP.n26 VP.n25 161.3
R1878 VP.n27 VP.n18 161.3
R1879 VP.n29 VP.n28 161.3
R1880 VP.n30 VP.n17 161.3
R1881 VP.n32 VP.n31 161.3
R1882 VP.n33 VP.n16 161.3
R1883 VP.n36 VP.n35 161.3
R1884 VP.n37 VP.n15 161.3
R1885 VP.n39 VP.n38 161.3
R1886 VP.n40 VP.n14 161.3
R1887 VP.n42 VP.n41 161.3
R1888 VP.n43 VP.n13 161.3
R1889 VP.n45 VP.n44 161.3
R1890 VP.n46 VP.n12 161.3
R1891 VP.n88 VP.n0 161.3
R1892 VP.n87 VP.n86 161.3
R1893 VP.n85 VP.n1 161.3
R1894 VP.n84 VP.n83 161.3
R1895 VP.n82 VP.n2 161.3
R1896 VP.n81 VP.n80 161.3
R1897 VP.n79 VP.n3 161.3
R1898 VP.n78 VP.n77 161.3
R1899 VP.n75 VP.n4 161.3
R1900 VP.n74 VP.n73 161.3
R1901 VP.n72 VP.n5 161.3
R1902 VP.n71 VP.n70 161.3
R1903 VP.n69 VP.n6 161.3
R1904 VP.n68 VP.n67 161.3
R1905 VP.n66 VP.n7 161.3
R1906 VP.n65 VP.n64 161.3
R1907 VP.n62 VP.n8 161.3
R1908 VP.n61 VP.n60 161.3
R1909 VP.n59 VP.n9 161.3
R1910 VP.n58 VP.n57 161.3
R1911 VP.n56 VP.n10 161.3
R1912 VP.n55 VP.n54 161.3
R1913 VP.n53 VP.n11 161.3
R1914 VP.n52 VP.n51 161.3
R1915 VP.n20 VP.t2 78.8767
R1916 VP.n50 VP.n49 61.1402
R1917 VP.n90 VP.n89 61.1402
R1918 VP.n48 VP.n47 61.1402
R1919 VP.n21 VP.n20 59.8759
R1920 VP.n70 VP.n69 56.5193
R1921 VP.n28 VP.n27 56.5193
R1922 VP.n49 VP.n48 53.1328
R1923 VP.n57 VP.n56 53.1199
R1924 VP.n83 VP.n82 53.1199
R1925 VP.n41 VP.n40 53.1199
R1926 VP.n50 VP.t3 46.6108
R1927 VP.n63 VP.t5 46.6108
R1928 VP.n76 VP.t4 46.6108
R1929 VP.n89 VP.t7 46.6108
R1930 VP.n47 VP.t1 46.6108
R1931 VP.n34 VP.t6 46.6108
R1932 VP.n21 VP.t0 46.6108
R1933 VP.n56 VP.n55 27.8669
R1934 VP.n83 VP.n1 27.8669
R1935 VP.n41 VP.n13 27.8669
R1936 VP.n51 VP.n11 24.4675
R1937 VP.n55 VP.n11 24.4675
R1938 VP.n57 VP.n9 24.4675
R1939 VP.n61 VP.n9 24.4675
R1940 VP.n62 VP.n61 24.4675
R1941 VP.n64 VP.n7 24.4675
R1942 VP.n68 VP.n7 24.4675
R1943 VP.n69 VP.n68 24.4675
R1944 VP.n70 VP.n5 24.4675
R1945 VP.n74 VP.n5 24.4675
R1946 VP.n75 VP.n74 24.4675
R1947 VP.n77 VP.n3 24.4675
R1948 VP.n81 VP.n3 24.4675
R1949 VP.n82 VP.n81 24.4675
R1950 VP.n87 VP.n1 24.4675
R1951 VP.n88 VP.n87 24.4675
R1952 VP.n45 VP.n13 24.4675
R1953 VP.n46 VP.n45 24.4675
R1954 VP.n28 VP.n17 24.4675
R1955 VP.n32 VP.n17 24.4675
R1956 VP.n33 VP.n32 24.4675
R1957 VP.n35 VP.n15 24.4675
R1958 VP.n39 VP.n15 24.4675
R1959 VP.n40 VP.n39 24.4675
R1960 VP.n22 VP.n19 24.4675
R1961 VP.n26 VP.n19 24.4675
R1962 VP.n27 VP.n26 24.4675
R1963 VP.n51 VP.n50 21.0421
R1964 VP.n89 VP.n88 21.0421
R1965 VP.n47 VP.n46 21.0421
R1966 VP.n64 VP.n63 15.17
R1967 VP.n76 VP.n75 15.17
R1968 VP.n34 VP.n33 15.17
R1969 VP.n22 VP.n21 15.17
R1970 VP.n63 VP.n62 9.29796
R1971 VP.n77 VP.n76 9.29796
R1972 VP.n35 VP.n34 9.29796
R1973 VP.n23 VP.n20 2.65257
R1974 VP.n48 VP.n12 0.417535
R1975 VP.n52 VP.n49 0.417535
R1976 VP.n90 VP.n0 0.417535
R1977 VP VP.n90 0.394291
R1978 VP.n24 VP.n23 0.189894
R1979 VP.n25 VP.n24 0.189894
R1980 VP.n25 VP.n18 0.189894
R1981 VP.n29 VP.n18 0.189894
R1982 VP.n30 VP.n29 0.189894
R1983 VP.n31 VP.n30 0.189894
R1984 VP.n31 VP.n16 0.189894
R1985 VP.n36 VP.n16 0.189894
R1986 VP.n37 VP.n36 0.189894
R1987 VP.n38 VP.n37 0.189894
R1988 VP.n38 VP.n14 0.189894
R1989 VP.n42 VP.n14 0.189894
R1990 VP.n43 VP.n42 0.189894
R1991 VP.n44 VP.n43 0.189894
R1992 VP.n44 VP.n12 0.189894
R1993 VP.n53 VP.n52 0.189894
R1994 VP.n54 VP.n53 0.189894
R1995 VP.n54 VP.n10 0.189894
R1996 VP.n58 VP.n10 0.189894
R1997 VP.n59 VP.n58 0.189894
R1998 VP.n60 VP.n59 0.189894
R1999 VP.n60 VP.n8 0.189894
R2000 VP.n65 VP.n8 0.189894
R2001 VP.n66 VP.n65 0.189894
R2002 VP.n67 VP.n66 0.189894
R2003 VP.n67 VP.n6 0.189894
R2004 VP.n71 VP.n6 0.189894
R2005 VP.n72 VP.n71 0.189894
R2006 VP.n73 VP.n72 0.189894
R2007 VP.n73 VP.n4 0.189894
R2008 VP.n78 VP.n4 0.189894
R2009 VP.n79 VP.n78 0.189894
R2010 VP.n80 VP.n79 0.189894
R2011 VP.n80 VP.n2 0.189894
R2012 VP.n84 VP.n2 0.189894
R2013 VP.n85 VP.n84 0.189894
R2014 VP.n86 VP.n85 0.189894
R2015 VP.n86 VP.n0 0.189894
R2016 VDD1 VDD1.n0 85.0032
R2017 VDD1.n3 VDD1.n2 84.8895
R2018 VDD1.n3 VDD1.n1 84.8895
R2019 VDD1.n5 VDD1.n4 83.169
R2020 VDD1.n5 VDD1.n3 46.6
R2021 VDD1.n4 VDD1.t1 4.43502
R2022 VDD1.n4 VDD1.t6 4.43502
R2023 VDD1.n0 VDD1.t5 4.43502
R2024 VDD1.n0 VDD1.t7 4.43502
R2025 VDD1.n2 VDD1.t3 4.43502
R2026 VDD1.n2 VDD1.t0 4.43502
R2027 VDD1.n1 VDD1.t4 4.43502
R2028 VDD1.n1 VDD1.t2 4.43502
R2029 VDD1 VDD1.n5 1.71817
C0 VP B 2.56727f
C1 VDD1 VDD2 2.3951f
C2 VN VDD2 5.83545f
C3 VTAIL VDD2 7.3646f
C4 B VDD2 2.02058f
C5 VP w_n5090_n2434# 11.2775f
C6 VN VDD1 0.153885f
C7 w_n5090_n2434# VDD2 2.37637f
C8 VDD1 VTAIL 7.30221f
C9 VN VTAIL 6.85636f
C10 B VDD1 1.88712f
C11 VN B 1.44734f
C12 B VTAIL 3.85047f
C13 VDD1 w_n5090_n2434# 2.21174f
C14 VN w_n5090_n2434# 10.6132f
C15 w_n5090_n2434# VTAIL 3.30493f
C16 B w_n5090_n2434# 10.629f
C17 VP VDD2 0.646305f
C18 VP VDD1 6.325871f
C19 VN VP 8.25861f
C20 VP VTAIL 6.87047f
C21 VDD2 VSUBS 2.50476f
C22 VDD1 VSUBS 3.19701f
C23 VTAIL VSUBS 1.371791f
C24 VN VSUBS 8.351609f
C25 VP VSUBS 4.662338f
C26 B VSUBS 5.936588f
C27 w_n5090_n2434# VSUBS 0.153983p
C28 VDD1.t5 VSUBS 0.190503f
C29 VDD1.t7 VSUBS 0.190503f
C30 VDD1.n0 VSUBS 1.34921f
C31 VDD1.t4 VSUBS 0.190503f
C32 VDD1.t2 VSUBS 0.190503f
C33 VDD1.n1 VSUBS 1.34746f
C34 VDD1.t3 VSUBS 0.190503f
C35 VDD1.t0 VSUBS 0.190503f
C36 VDD1.n2 VSUBS 1.34746f
C37 VDD1.n3 VSUBS 5.50158f
C38 VDD1.t1 VSUBS 0.190503f
C39 VDD1.t6 VSUBS 0.190503f
C40 VDD1.n4 VSUBS 1.32426f
C41 VDD1.n5 VSUBS 4.29849f
C42 VP.n0 VSUBS 0.060685f
C43 VP.t7 VSUBS 2.39752f
C44 VP.n1 VSUBS 0.063241f
C45 VP.n2 VSUBS 0.032262f
C46 VP.n3 VSUBS 0.060128f
C47 VP.n4 VSUBS 0.032262f
C48 VP.t4 VSUBS 2.39752f
C49 VP.n5 VSUBS 0.060128f
C50 VP.n6 VSUBS 0.032262f
C51 VP.n7 VSUBS 0.060128f
C52 VP.n8 VSUBS 0.032262f
C53 VP.t5 VSUBS 2.39752f
C54 VP.n9 VSUBS 0.060128f
C55 VP.n10 VSUBS 0.032262f
C56 VP.n11 VSUBS 0.060128f
C57 VP.n12 VSUBS 0.060685f
C58 VP.t1 VSUBS 2.39752f
C59 VP.n13 VSUBS 0.063241f
C60 VP.n14 VSUBS 0.032262f
C61 VP.n15 VSUBS 0.060128f
C62 VP.n16 VSUBS 0.032262f
C63 VP.t6 VSUBS 2.39752f
C64 VP.n17 VSUBS 0.060128f
C65 VP.n18 VSUBS 0.032262f
C66 VP.n19 VSUBS 0.060128f
C67 VP.t2 VSUBS 2.85439f
C68 VP.n20 VSUBS 0.947954f
C69 VP.t0 VSUBS 2.39752f
C70 VP.n21 VSUBS 0.986188f
C71 VP.n22 VSUBS 0.048848f
C72 VP.n23 VSUBS 0.421534f
C73 VP.n24 VSUBS 0.032262f
C74 VP.n25 VSUBS 0.032262f
C75 VP.n26 VSUBS 0.060128f
C76 VP.n27 VSUBS 0.047097f
C77 VP.n28 VSUBS 0.047097f
C78 VP.n29 VSUBS 0.032262f
C79 VP.n30 VSUBS 0.032262f
C80 VP.n31 VSUBS 0.032262f
C81 VP.n32 VSUBS 0.060128f
C82 VP.n33 VSUBS 0.048848f
C83 VP.n34 VSUBS 0.866933f
C84 VP.n35 VSUBS 0.041723f
C85 VP.n36 VSUBS 0.032262f
C86 VP.n37 VSUBS 0.032262f
C87 VP.n38 VSUBS 0.032262f
C88 VP.n39 VSUBS 0.060128f
C89 VP.n40 VSUBS 0.057243f
C90 VP.n41 VSUBS 0.033838f
C91 VP.n42 VSUBS 0.032262f
C92 VP.n43 VSUBS 0.032262f
C93 VP.n44 VSUBS 0.032262f
C94 VP.n45 VSUBS 0.060128f
C95 VP.n46 VSUBS 0.055972f
C96 VP.n47 VSUBS 1.00525f
C97 VP.n48 VSUBS 2.03712f
C98 VP.n49 VSUBS 2.05895f
C99 VP.t3 VSUBS 2.39752f
C100 VP.n50 VSUBS 1.00525f
C101 VP.n51 VSUBS 0.055972f
C102 VP.n52 VSUBS 0.060685f
C103 VP.n53 VSUBS 0.032262f
C104 VP.n54 VSUBS 0.032262f
C105 VP.n55 VSUBS 0.063241f
C106 VP.n56 VSUBS 0.033838f
C107 VP.n57 VSUBS 0.057243f
C108 VP.n58 VSUBS 0.032262f
C109 VP.n59 VSUBS 0.032262f
C110 VP.n60 VSUBS 0.032262f
C111 VP.n61 VSUBS 0.060128f
C112 VP.n62 VSUBS 0.041723f
C113 VP.n63 VSUBS 0.866933f
C114 VP.n64 VSUBS 0.048848f
C115 VP.n65 VSUBS 0.032262f
C116 VP.n66 VSUBS 0.032262f
C117 VP.n67 VSUBS 0.032262f
C118 VP.n68 VSUBS 0.060128f
C119 VP.n69 VSUBS 0.047097f
C120 VP.n70 VSUBS 0.047097f
C121 VP.n71 VSUBS 0.032262f
C122 VP.n72 VSUBS 0.032262f
C123 VP.n73 VSUBS 0.032262f
C124 VP.n74 VSUBS 0.060128f
C125 VP.n75 VSUBS 0.048848f
C126 VP.n76 VSUBS 0.866933f
C127 VP.n77 VSUBS 0.041723f
C128 VP.n78 VSUBS 0.032262f
C129 VP.n79 VSUBS 0.032262f
C130 VP.n80 VSUBS 0.032262f
C131 VP.n81 VSUBS 0.060128f
C132 VP.n82 VSUBS 0.057243f
C133 VP.n83 VSUBS 0.033838f
C134 VP.n84 VSUBS 0.032262f
C135 VP.n85 VSUBS 0.032262f
C136 VP.n86 VSUBS 0.032262f
C137 VP.n87 VSUBS 0.060128f
C138 VP.n88 VSUBS 0.055972f
C139 VP.n89 VSUBS 1.00525f
C140 VP.n90 VSUBS 0.098753f
C141 VTAIL.t9 VSUBS 0.16963f
C142 VTAIL.t13 VSUBS 0.16963f
C143 VTAIL.n0 VSUBS 1.05278f
C144 VTAIL.n1 VSUBS 0.936631f
C145 VTAIL.n2 VSUBS 0.031683f
C146 VTAIL.n3 VSUBS 0.029285f
C147 VTAIL.n4 VSUBS 0.015736f
C148 VTAIL.n5 VSUBS 0.037195f
C149 VTAIL.n6 VSUBS 0.016662f
C150 VTAIL.n7 VSUBS 0.029285f
C151 VTAIL.n8 VSUBS 0.015736f
C152 VTAIL.n9 VSUBS 0.037195f
C153 VTAIL.n10 VSUBS 0.016662f
C154 VTAIL.n11 VSUBS 0.029285f
C155 VTAIL.n12 VSUBS 0.015736f
C156 VTAIL.n13 VSUBS 0.027897f
C157 VTAIL.n14 VSUBS 0.02366f
C158 VTAIL.t15 VSUBS 0.07935f
C159 VTAIL.n15 VSUBS 0.140456f
C160 VTAIL.n16 VSUBS 0.84966f
C161 VTAIL.n17 VSUBS 0.015736f
C162 VTAIL.n18 VSUBS 0.016662f
C163 VTAIL.n19 VSUBS 0.037195f
C164 VTAIL.n20 VSUBS 0.037195f
C165 VTAIL.n21 VSUBS 0.016662f
C166 VTAIL.n22 VSUBS 0.015736f
C167 VTAIL.n23 VSUBS 0.029285f
C168 VTAIL.n24 VSUBS 0.029285f
C169 VTAIL.n25 VSUBS 0.015736f
C170 VTAIL.n26 VSUBS 0.016662f
C171 VTAIL.n27 VSUBS 0.037195f
C172 VTAIL.n28 VSUBS 0.037195f
C173 VTAIL.n29 VSUBS 0.016662f
C174 VTAIL.n30 VSUBS 0.015736f
C175 VTAIL.n31 VSUBS 0.029285f
C176 VTAIL.n32 VSUBS 0.029285f
C177 VTAIL.n33 VSUBS 0.015736f
C178 VTAIL.n34 VSUBS 0.016662f
C179 VTAIL.n35 VSUBS 0.037195f
C180 VTAIL.n36 VSUBS 0.08836f
C181 VTAIL.n37 VSUBS 0.016662f
C182 VTAIL.n38 VSUBS 0.015736f
C183 VTAIL.n39 VSUBS 0.06329f
C184 VTAIL.n40 VSUBS 0.044221f
C185 VTAIL.n41 VSUBS 0.402018f
C186 VTAIL.n42 VSUBS 0.031683f
C187 VTAIL.n43 VSUBS 0.029285f
C188 VTAIL.n44 VSUBS 0.015736f
C189 VTAIL.n45 VSUBS 0.037195f
C190 VTAIL.n46 VSUBS 0.016662f
C191 VTAIL.n47 VSUBS 0.029285f
C192 VTAIL.n48 VSUBS 0.015736f
C193 VTAIL.n49 VSUBS 0.037195f
C194 VTAIL.n50 VSUBS 0.016662f
C195 VTAIL.n51 VSUBS 0.029285f
C196 VTAIL.n52 VSUBS 0.015736f
C197 VTAIL.n53 VSUBS 0.027897f
C198 VTAIL.n54 VSUBS 0.02366f
C199 VTAIL.t2 VSUBS 0.07935f
C200 VTAIL.n55 VSUBS 0.140456f
C201 VTAIL.n56 VSUBS 0.84966f
C202 VTAIL.n57 VSUBS 0.015736f
C203 VTAIL.n58 VSUBS 0.016662f
C204 VTAIL.n59 VSUBS 0.037195f
C205 VTAIL.n60 VSUBS 0.037195f
C206 VTAIL.n61 VSUBS 0.016662f
C207 VTAIL.n62 VSUBS 0.015736f
C208 VTAIL.n63 VSUBS 0.029285f
C209 VTAIL.n64 VSUBS 0.029285f
C210 VTAIL.n65 VSUBS 0.015736f
C211 VTAIL.n66 VSUBS 0.016662f
C212 VTAIL.n67 VSUBS 0.037195f
C213 VTAIL.n68 VSUBS 0.037195f
C214 VTAIL.n69 VSUBS 0.016662f
C215 VTAIL.n70 VSUBS 0.015736f
C216 VTAIL.n71 VSUBS 0.029285f
C217 VTAIL.n72 VSUBS 0.029285f
C218 VTAIL.n73 VSUBS 0.015736f
C219 VTAIL.n74 VSUBS 0.016662f
C220 VTAIL.n75 VSUBS 0.037195f
C221 VTAIL.n76 VSUBS 0.08836f
C222 VTAIL.n77 VSUBS 0.016662f
C223 VTAIL.n78 VSUBS 0.015736f
C224 VTAIL.n79 VSUBS 0.06329f
C225 VTAIL.n80 VSUBS 0.044221f
C226 VTAIL.n81 VSUBS 0.402018f
C227 VTAIL.t1 VSUBS 0.16963f
C228 VTAIL.t4 VSUBS 0.16963f
C229 VTAIL.n82 VSUBS 1.05278f
C230 VTAIL.n83 VSUBS 1.26629f
C231 VTAIL.n84 VSUBS 0.031683f
C232 VTAIL.n85 VSUBS 0.029285f
C233 VTAIL.n86 VSUBS 0.015736f
C234 VTAIL.n87 VSUBS 0.037195f
C235 VTAIL.n88 VSUBS 0.016662f
C236 VTAIL.n89 VSUBS 0.029285f
C237 VTAIL.n90 VSUBS 0.015736f
C238 VTAIL.n91 VSUBS 0.037195f
C239 VTAIL.n92 VSUBS 0.016662f
C240 VTAIL.n93 VSUBS 0.029285f
C241 VTAIL.n94 VSUBS 0.015736f
C242 VTAIL.n95 VSUBS 0.027897f
C243 VTAIL.n96 VSUBS 0.02366f
C244 VTAIL.t3 VSUBS 0.07935f
C245 VTAIL.n97 VSUBS 0.140456f
C246 VTAIL.n98 VSUBS 0.84966f
C247 VTAIL.n99 VSUBS 0.015736f
C248 VTAIL.n100 VSUBS 0.016662f
C249 VTAIL.n101 VSUBS 0.037195f
C250 VTAIL.n102 VSUBS 0.037195f
C251 VTAIL.n103 VSUBS 0.016662f
C252 VTAIL.n104 VSUBS 0.015736f
C253 VTAIL.n105 VSUBS 0.029285f
C254 VTAIL.n106 VSUBS 0.029285f
C255 VTAIL.n107 VSUBS 0.015736f
C256 VTAIL.n108 VSUBS 0.016662f
C257 VTAIL.n109 VSUBS 0.037195f
C258 VTAIL.n110 VSUBS 0.037195f
C259 VTAIL.n111 VSUBS 0.016662f
C260 VTAIL.n112 VSUBS 0.015736f
C261 VTAIL.n113 VSUBS 0.029285f
C262 VTAIL.n114 VSUBS 0.029285f
C263 VTAIL.n115 VSUBS 0.015736f
C264 VTAIL.n116 VSUBS 0.016662f
C265 VTAIL.n117 VSUBS 0.037195f
C266 VTAIL.n118 VSUBS 0.08836f
C267 VTAIL.n119 VSUBS 0.016662f
C268 VTAIL.n120 VSUBS 0.015736f
C269 VTAIL.n121 VSUBS 0.06329f
C270 VTAIL.n122 VSUBS 0.044221f
C271 VTAIL.n123 VSUBS 1.68691f
C272 VTAIL.n124 VSUBS 0.031683f
C273 VTAIL.n125 VSUBS 0.029285f
C274 VTAIL.n126 VSUBS 0.015736f
C275 VTAIL.n127 VSUBS 0.037195f
C276 VTAIL.n128 VSUBS 0.016662f
C277 VTAIL.n129 VSUBS 0.029285f
C278 VTAIL.n130 VSUBS 0.015736f
C279 VTAIL.n131 VSUBS 0.037195f
C280 VTAIL.n132 VSUBS 0.016662f
C281 VTAIL.n133 VSUBS 0.029285f
C282 VTAIL.n134 VSUBS 0.015736f
C283 VTAIL.n135 VSUBS 0.027897f
C284 VTAIL.n136 VSUBS 0.02366f
C285 VTAIL.t8 VSUBS 0.07935f
C286 VTAIL.n137 VSUBS 0.140456f
C287 VTAIL.n138 VSUBS 0.84966f
C288 VTAIL.n139 VSUBS 0.015736f
C289 VTAIL.n140 VSUBS 0.016662f
C290 VTAIL.n141 VSUBS 0.037195f
C291 VTAIL.n142 VSUBS 0.037195f
C292 VTAIL.n143 VSUBS 0.016662f
C293 VTAIL.n144 VSUBS 0.015736f
C294 VTAIL.n145 VSUBS 0.029285f
C295 VTAIL.n146 VSUBS 0.029285f
C296 VTAIL.n147 VSUBS 0.015736f
C297 VTAIL.n148 VSUBS 0.016662f
C298 VTAIL.n149 VSUBS 0.037195f
C299 VTAIL.n150 VSUBS 0.037195f
C300 VTAIL.n151 VSUBS 0.016662f
C301 VTAIL.n152 VSUBS 0.015736f
C302 VTAIL.n153 VSUBS 0.029285f
C303 VTAIL.n154 VSUBS 0.029285f
C304 VTAIL.n155 VSUBS 0.015736f
C305 VTAIL.n156 VSUBS 0.016662f
C306 VTAIL.n157 VSUBS 0.037195f
C307 VTAIL.n158 VSUBS 0.08836f
C308 VTAIL.n159 VSUBS 0.016662f
C309 VTAIL.n160 VSUBS 0.015736f
C310 VTAIL.n161 VSUBS 0.06329f
C311 VTAIL.n162 VSUBS 0.044221f
C312 VTAIL.n163 VSUBS 1.68691f
C313 VTAIL.t14 VSUBS 0.16963f
C314 VTAIL.t12 VSUBS 0.16963f
C315 VTAIL.n164 VSUBS 1.05279f
C316 VTAIL.n165 VSUBS 1.26628f
C317 VTAIL.n166 VSUBS 0.031683f
C318 VTAIL.n167 VSUBS 0.029285f
C319 VTAIL.n168 VSUBS 0.015736f
C320 VTAIL.n169 VSUBS 0.037195f
C321 VTAIL.n170 VSUBS 0.016662f
C322 VTAIL.n171 VSUBS 0.029285f
C323 VTAIL.n172 VSUBS 0.015736f
C324 VTAIL.n173 VSUBS 0.037195f
C325 VTAIL.n174 VSUBS 0.016662f
C326 VTAIL.n175 VSUBS 0.029285f
C327 VTAIL.n176 VSUBS 0.015736f
C328 VTAIL.n177 VSUBS 0.027897f
C329 VTAIL.n178 VSUBS 0.02366f
C330 VTAIL.t10 VSUBS 0.07935f
C331 VTAIL.n179 VSUBS 0.140456f
C332 VTAIL.n180 VSUBS 0.84966f
C333 VTAIL.n181 VSUBS 0.015736f
C334 VTAIL.n182 VSUBS 0.016662f
C335 VTAIL.n183 VSUBS 0.037195f
C336 VTAIL.n184 VSUBS 0.037195f
C337 VTAIL.n185 VSUBS 0.016662f
C338 VTAIL.n186 VSUBS 0.015736f
C339 VTAIL.n187 VSUBS 0.029285f
C340 VTAIL.n188 VSUBS 0.029285f
C341 VTAIL.n189 VSUBS 0.015736f
C342 VTAIL.n190 VSUBS 0.016662f
C343 VTAIL.n191 VSUBS 0.037195f
C344 VTAIL.n192 VSUBS 0.037195f
C345 VTAIL.n193 VSUBS 0.016662f
C346 VTAIL.n194 VSUBS 0.015736f
C347 VTAIL.n195 VSUBS 0.029285f
C348 VTAIL.n196 VSUBS 0.029285f
C349 VTAIL.n197 VSUBS 0.015736f
C350 VTAIL.n198 VSUBS 0.016662f
C351 VTAIL.n199 VSUBS 0.037195f
C352 VTAIL.n200 VSUBS 0.08836f
C353 VTAIL.n201 VSUBS 0.016662f
C354 VTAIL.n202 VSUBS 0.015736f
C355 VTAIL.n203 VSUBS 0.06329f
C356 VTAIL.n204 VSUBS 0.044221f
C357 VTAIL.n205 VSUBS 0.402018f
C358 VTAIL.n206 VSUBS 0.031683f
C359 VTAIL.n207 VSUBS 0.029285f
C360 VTAIL.n208 VSUBS 0.015736f
C361 VTAIL.n209 VSUBS 0.037195f
C362 VTAIL.n210 VSUBS 0.016662f
C363 VTAIL.n211 VSUBS 0.029285f
C364 VTAIL.n212 VSUBS 0.015736f
C365 VTAIL.n213 VSUBS 0.037195f
C366 VTAIL.n214 VSUBS 0.016662f
C367 VTAIL.n215 VSUBS 0.029285f
C368 VTAIL.n216 VSUBS 0.015736f
C369 VTAIL.n217 VSUBS 0.027897f
C370 VTAIL.n218 VSUBS 0.02366f
C371 VTAIL.t5 VSUBS 0.07935f
C372 VTAIL.n219 VSUBS 0.140456f
C373 VTAIL.n220 VSUBS 0.84966f
C374 VTAIL.n221 VSUBS 0.015736f
C375 VTAIL.n222 VSUBS 0.016662f
C376 VTAIL.n223 VSUBS 0.037195f
C377 VTAIL.n224 VSUBS 0.037195f
C378 VTAIL.n225 VSUBS 0.016662f
C379 VTAIL.n226 VSUBS 0.015736f
C380 VTAIL.n227 VSUBS 0.029285f
C381 VTAIL.n228 VSUBS 0.029285f
C382 VTAIL.n229 VSUBS 0.015736f
C383 VTAIL.n230 VSUBS 0.016662f
C384 VTAIL.n231 VSUBS 0.037195f
C385 VTAIL.n232 VSUBS 0.037195f
C386 VTAIL.n233 VSUBS 0.016662f
C387 VTAIL.n234 VSUBS 0.015736f
C388 VTAIL.n235 VSUBS 0.029285f
C389 VTAIL.n236 VSUBS 0.029285f
C390 VTAIL.n237 VSUBS 0.015736f
C391 VTAIL.n238 VSUBS 0.016662f
C392 VTAIL.n239 VSUBS 0.037195f
C393 VTAIL.n240 VSUBS 0.08836f
C394 VTAIL.n241 VSUBS 0.016662f
C395 VTAIL.n242 VSUBS 0.015736f
C396 VTAIL.n243 VSUBS 0.06329f
C397 VTAIL.n244 VSUBS 0.044221f
C398 VTAIL.n245 VSUBS 0.402018f
C399 VTAIL.t6 VSUBS 0.16963f
C400 VTAIL.t7 VSUBS 0.16963f
C401 VTAIL.n246 VSUBS 1.05279f
C402 VTAIL.n247 VSUBS 1.26628f
C403 VTAIL.n248 VSUBS 0.031683f
C404 VTAIL.n249 VSUBS 0.029285f
C405 VTAIL.n250 VSUBS 0.015736f
C406 VTAIL.n251 VSUBS 0.037195f
C407 VTAIL.n252 VSUBS 0.016662f
C408 VTAIL.n253 VSUBS 0.029285f
C409 VTAIL.n254 VSUBS 0.015736f
C410 VTAIL.n255 VSUBS 0.037195f
C411 VTAIL.n256 VSUBS 0.016662f
C412 VTAIL.n257 VSUBS 0.029285f
C413 VTAIL.n258 VSUBS 0.015736f
C414 VTAIL.n259 VSUBS 0.027897f
C415 VTAIL.n260 VSUBS 0.02366f
C416 VTAIL.t0 VSUBS 0.07935f
C417 VTAIL.n261 VSUBS 0.140456f
C418 VTAIL.n262 VSUBS 0.84966f
C419 VTAIL.n263 VSUBS 0.015736f
C420 VTAIL.n264 VSUBS 0.016662f
C421 VTAIL.n265 VSUBS 0.037195f
C422 VTAIL.n266 VSUBS 0.037195f
C423 VTAIL.n267 VSUBS 0.016662f
C424 VTAIL.n268 VSUBS 0.015736f
C425 VTAIL.n269 VSUBS 0.029285f
C426 VTAIL.n270 VSUBS 0.029285f
C427 VTAIL.n271 VSUBS 0.015736f
C428 VTAIL.n272 VSUBS 0.016662f
C429 VTAIL.n273 VSUBS 0.037195f
C430 VTAIL.n274 VSUBS 0.037195f
C431 VTAIL.n275 VSUBS 0.016662f
C432 VTAIL.n276 VSUBS 0.015736f
C433 VTAIL.n277 VSUBS 0.029285f
C434 VTAIL.n278 VSUBS 0.029285f
C435 VTAIL.n279 VSUBS 0.015736f
C436 VTAIL.n280 VSUBS 0.016662f
C437 VTAIL.n281 VSUBS 0.037195f
C438 VTAIL.n282 VSUBS 0.08836f
C439 VTAIL.n283 VSUBS 0.016662f
C440 VTAIL.n284 VSUBS 0.015736f
C441 VTAIL.n285 VSUBS 0.06329f
C442 VTAIL.n286 VSUBS 0.044221f
C443 VTAIL.n287 VSUBS 1.68691f
C444 VTAIL.n288 VSUBS 0.031683f
C445 VTAIL.n289 VSUBS 0.029285f
C446 VTAIL.n290 VSUBS 0.015736f
C447 VTAIL.n291 VSUBS 0.037195f
C448 VTAIL.n292 VSUBS 0.016662f
C449 VTAIL.n293 VSUBS 0.029285f
C450 VTAIL.n294 VSUBS 0.015736f
C451 VTAIL.n295 VSUBS 0.037195f
C452 VTAIL.n296 VSUBS 0.016662f
C453 VTAIL.n297 VSUBS 0.029285f
C454 VTAIL.n298 VSUBS 0.015736f
C455 VTAIL.n299 VSUBS 0.027897f
C456 VTAIL.n300 VSUBS 0.02366f
C457 VTAIL.t11 VSUBS 0.07935f
C458 VTAIL.n301 VSUBS 0.140456f
C459 VTAIL.n302 VSUBS 0.84966f
C460 VTAIL.n303 VSUBS 0.015736f
C461 VTAIL.n304 VSUBS 0.016662f
C462 VTAIL.n305 VSUBS 0.037195f
C463 VTAIL.n306 VSUBS 0.037195f
C464 VTAIL.n307 VSUBS 0.016662f
C465 VTAIL.n308 VSUBS 0.015736f
C466 VTAIL.n309 VSUBS 0.029285f
C467 VTAIL.n310 VSUBS 0.029285f
C468 VTAIL.n311 VSUBS 0.015736f
C469 VTAIL.n312 VSUBS 0.016662f
C470 VTAIL.n313 VSUBS 0.037195f
C471 VTAIL.n314 VSUBS 0.037195f
C472 VTAIL.n315 VSUBS 0.016662f
C473 VTAIL.n316 VSUBS 0.015736f
C474 VTAIL.n317 VSUBS 0.029285f
C475 VTAIL.n318 VSUBS 0.029285f
C476 VTAIL.n319 VSUBS 0.015736f
C477 VTAIL.n320 VSUBS 0.016662f
C478 VTAIL.n321 VSUBS 0.037195f
C479 VTAIL.n322 VSUBS 0.08836f
C480 VTAIL.n323 VSUBS 0.016662f
C481 VTAIL.n324 VSUBS 0.015736f
C482 VTAIL.n325 VSUBS 0.06329f
C483 VTAIL.n326 VSUBS 0.044221f
C484 VTAIL.n327 VSUBS 1.68142f
C485 VDD2.t0 VSUBS 0.21075f
C486 VDD2.t6 VSUBS 0.21075f
C487 VDD2.n0 VSUBS 1.49067f
C488 VDD2.t2 VSUBS 0.21075f
C489 VDD2.t4 VSUBS 0.21075f
C490 VDD2.n1 VSUBS 1.49067f
C491 VDD2.n2 VSUBS 6.01124f
C492 VDD2.t7 VSUBS 0.21075f
C493 VDD2.t1 VSUBS 0.21075f
C494 VDD2.n3 VSUBS 1.46502f
C495 VDD2.n4 VSUBS 4.70968f
C496 VDD2.t3 VSUBS 0.21075f
C497 VDD2.t5 VSUBS 0.21075f
C498 VDD2.n5 VSUBS 1.49061f
C499 VN.n0 VSUBS 0.054101f
C500 VN.t4 VSUBS 2.13742f
C501 VN.n1 VSUBS 0.05638f
C502 VN.n2 VSUBS 0.028762f
C503 VN.n3 VSUBS 0.053605f
C504 VN.n4 VSUBS 0.028762f
C505 VN.t2 VSUBS 2.13742f
C506 VN.n5 VSUBS 0.053605f
C507 VN.n6 VSUBS 0.028762f
C508 VN.n7 VSUBS 0.053605f
C509 VN.t0 VSUBS 2.54473f
C510 VN.n8 VSUBS 0.845111f
C511 VN.t6 VSUBS 2.13742f
C512 VN.n9 VSUBS 0.8792f
C513 VN.n10 VSUBS 0.043548f
C514 VN.n11 VSUBS 0.375802f
C515 VN.n12 VSUBS 0.028762f
C516 VN.n13 VSUBS 0.028762f
C517 VN.n14 VSUBS 0.053605f
C518 VN.n15 VSUBS 0.041987f
C519 VN.n16 VSUBS 0.041987f
C520 VN.n17 VSUBS 0.028762f
C521 VN.n18 VSUBS 0.028762f
C522 VN.n19 VSUBS 0.028762f
C523 VN.n20 VSUBS 0.053605f
C524 VN.n21 VSUBS 0.043548f
C525 VN.n22 VSUBS 0.772882f
C526 VN.n23 VSUBS 0.037197f
C527 VN.n24 VSUBS 0.028762f
C528 VN.n25 VSUBS 0.028762f
C529 VN.n26 VSUBS 0.028762f
C530 VN.n27 VSUBS 0.053605f
C531 VN.n28 VSUBS 0.051033f
C532 VN.n29 VSUBS 0.030167f
C533 VN.n30 VSUBS 0.028762f
C534 VN.n31 VSUBS 0.028762f
C535 VN.n32 VSUBS 0.028762f
C536 VN.n33 VSUBS 0.053605f
C537 VN.n34 VSUBS 0.0499f
C538 VN.n35 VSUBS 0.896194f
C539 VN.n36 VSUBS 0.088039f
C540 VN.n37 VSUBS 0.054101f
C541 VN.t7 VSUBS 2.13742f
C542 VN.n38 VSUBS 0.05638f
C543 VN.n39 VSUBS 0.028762f
C544 VN.n40 VSUBS 0.053605f
C545 VN.n41 VSUBS 0.028762f
C546 VN.t1 VSUBS 2.13742f
C547 VN.n42 VSUBS 0.053605f
C548 VN.n43 VSUBS 0.028762f
C549 VN.n44 VSUBS 0.053605f
C550 VN.t5 VSUBS 2.54473f
C551 VN.n45 VSUBS 0.845111f
C552 VN.t3 VSUBS 2.13742f
C553 VN.n46 VSUBS 0.8792f
C554 VN.n47 VSUBS 0.043548f
C555 VN.n48 VSUBS 0.375802f
C556 VN.n49 VSUBS 0.028762f
C557 VN.n50 VSUBS 0.028762f
C558 VN.n51 VSUBS 0.053605f
C559 VN.n52 VSUBS 0.041987f
C560 VN.n53 VSUBS 0.041987f
C561 VN.n54 VSUBS 0.028762f
C562 VN.n55 VSUBS 0.028762f
C563 VN.n56 VSUBS 0.028762f
C564 VN.n57 VSUBS 0.053605f
C565 VN.n58 VSUBS 0.043548f
C566 VN.n59 VSUBS 0.772882f
C567 VN.n60 VSUBS 0.037197f
C568 VN.n61 VSUBS 0.028762f
C569 VN.n62 VSUBS 0.028762f
C570 VN.n63 VSUBS 0.028762f
C571 VN.n64 VSUBS 0.053605f
C572 VN.n65 VSUBS 0.051033f
C573 VN.n66 VSUBS 0.030167f
C574 VN.n67 VSUBS 0.028762f
C575 VN.n68 VSUBS 0.028762f
C576 VN.n69 VSUBS 0.028762f
C577 VN.n70 VSUBS 0.053605f
C578 VN.n71 VSUBS 0.0499f
C579 VN.n72 VSUBS 0.896194f
C580 VN.n73 VSUBS 1.82332f
C581 B.n0 VSUBS 0.008422f
C582 B.n1 VSUBS 0.008422f
C583 B.n2 VSUBS 0.012456f
C584 B.n3 VSUBS 0.009545f
C585 B.n4 VSUBS 0.009545f
C586 B.n5 VSUBS 0.009545f
C587 B.n6 VSUBS 0.009545f
C588 B.n7 VSUBS 0.009545f
C589 B.n8 VSUBS 0.009545f
C590 B.n9 VSUBS 0.009545f
C591 B.n10 VSUBS 0.009545f
C592 B.n11 VSUBS 0.009545f
C593 B.n12 VSUBS 0.009545f
C594 B.n13 VSUBS 0.009545f
C595 B.n14 VSUBS 0.009545f
C596 B.n15 VSUBS 0.009545f
C597 B.n16 VSUBS 0.009545f
C598 B.n17 VSUBS 0.009545f
C599 B.n18 VSUBS 0.009545f
C600 B.n19 VSUBS 0.009545f
C601 B.n20 VSUBS 0.009545f
C602 B.n21 VSUBS 0.009545f
C603 B.n22 VSUBS 0.009545f
C604 B.n23 VSUBS 0.009545f
C605 B.n24 VSUBS 0.009545f
C606 B.n25 VSUBS 0.009545f
C607 B.n26 VSUBS 0.009545f
C608 B.n27 VSUBS 0.009545f
C609 B.n28 VSUBS 0.009545f
C610 B.n29 VSUBS 0.009545f
C611 B.n30 VSUBS 0.009545f
C612 B.n31 VSUBS 0.009545f
C613 B.n32 VSUBS 0.009545f
C614 B.n33 VSUBS 0.009545f
C615 B.n34 VSUBS 0.009545f
C616 B.n35 VSUBS 0.009545f
C617 B.n36 VSUBS 0.02451f
C618 B.n37 VSUBS 0.009545f
C619 B.n38 VSUBS 0.009545f
C620 B.n39 VSUBS 0.009545f
C621 B.n40 VSUBS 0.009545f
C622 B.n41 VSUBS 0.009545f
C623 B.n42 VSUBS 0.009545f
C624 B.n43 VSUBS 0.009545f
C625 B.n44 VSUBS 0.009545f
C626 B.n45 VSUBS 0.009545f
C627 B.n46 VSUBS 0.009545f
C628 B.n47 VSUBS 0.009545f
C629 B.n48 VSUBS 0.009545f
C630 B.n49 VSUBS 0.009545f
C631 B.t10 VSUBS 0.155049f
C632 B.t11 VSUBS 0.206432f
C633 B.t9 VSUBS 1.80719f
C634 B.n50 VSUBS 0.336625f
C635 B.n51 VSUBS 0.252588f
C636 B.n52 VSUBS 0.022115f
C637 B.n53 VSUBS 0.009545f
C638 B.n54 VSUBS 0.009545f
C639 B.n55 VSUBS 0.009545f
C640 B.n56 VSUBS 0.009545f
C641 B.n57 VSUBS 0.009545f
C642 B.t1 VSUBS 0.155052f
C643 B.t2 VSUBS 0.206435f
C644 B.t0 VSUBS 1.80719f
C645 B.n58 VSUBS 0.336623f
C646 B.n59 VSUBS 0.252585f
C647 B.n60 VSUBS 0.009545f
C648 B.n61 VSUBS 0.009545f
C649 B.n62 VSUBS 0.009545f
C650 B.n63 VSUBS 0.009545f
C651 B.n64 VSUBS 0.009545f
C652 B.n65 VSUBS 0.009545f
C653 B.n66 VSUBS 0.009545f
C654 B.n67 VSUBS 0.009545f
C655 B.n68 VSUBS 0.009545f
C656 B.n69 VSUBS 0.009545f
C657 B.n70 VSUBS 0.009545f
C658 B.n71 VSUBS 0.009545f
C659 B.n72 VSUBS 0.009545f
C660 B.n73 VSUBS 0.023497f
C661 B.n74 VSUBS 0.009545f
C662 B.n75 VSUBS 0.009545f
C663 B.n76 VSUBS 0.009545f
C664 B.n77 VSUBS 0.009545f
C665 B.n78 VSUBS 0.009545f
C666 B.n79 VSUBS 0.009545f
C667 B.n80 VSUBS 0.009545f
C668 B.n81 VSUBS 0.009545f
C669 B.n82 VSUBS 0.009545f
C670 B.n83 VSUBS 0.009545f
C671 B.n84 VSUBS 0.009545f
C672 B.n85 VSUBS 0.009545f
C673 B.n86 VSUBS 0.009545f
C674 B.n87 VSUBS 0.009545f
C675 B.n88 VSUBS 0.009545f
C676 B.n89 VSUBS 0.009545f
C677 B.n90 VSUBS 0.009545f
C678 B.n91 VSUBS 0.009545f
C679 B.n92 VSUBS 0.009545f
C680 B.n93 VSUBS 0.009545f
C681 B.n94 VSUBS 0.009545f
C682 B.n95 VSUBS 0.009545f
C683 B.n96 VSUBS 0.009545f
C684 B.n97 VSUBS 0.009545f
C685 B.n98 VSUBS 0.009545f
C686 B.n99 VSUBS 0.009545f
C687 B.n100 VSUBS 0.009545f
C688 B.n101 VSUBS 0.009545f
C689 B.n102 VSUBS 0.009545f
C690 B.n103 VSUBS 0.009545f
C691 B.n104 VSUBS 0.009545f
C692 B.n105 VSUBS 0.009545f
C693 B.n106 VSUBS 0.009545f
C694 B.n107 VSUBS 0.009545f
C695 B.n108 VSUBS 0.009545f
C696 B.n109 VSUBS 0.009545f
C697 B.n110 VSUBS 0.009545f
C698 B.n111 VSUBS 0.009545f
C699 B.n112 VSUBS 0.009545f
C700 B.n113 VSUBS 0.009545f
C701 B.n114 VSUBS 0.009545f
C702 B.n115 VSUBS 0.009545f
C703 B.n116 VSUBS 0.009545f
C704 B.n117 VSUBS 0.009545f
C705 B.n118 VSUBS 0.009545f
C706 B.n119 VSUBS 0.009545f
C707 B.n120 VSUBS 0.009545f
C708 B.n121 VSUBS 0.009545f
C709 B.n122 VSUBS 0.009545f
C710 B.n123 VSUBS 0.009545f
C711 B.n124 VSUBS 0.009545f
C712 B.n125 VSUBS 0.009545f
C713 B.n126 VSUBS 0.009545f
C714 B.n127 VSUBS 0.009545f
C715 B.n128 VSUBS 0.009545f
C716 B.n129 VSUBS 0.009545f
C717 B.n130 VSUBS 0.009545f
C718 B.n131 VSUBS 0.009545f
C719 B.n132 VSUBS 0.009545f
C720 B.n133 VSUBS 0.009545f
C721 B.n134 VSUBS 0.009545f
C722 B.n135 VSUBS 0.009545f
C723 B.n136 VSUBS 0.009545f
C724 B.n137 VSUBS 0.009545f
C725 B.n138 VSUBS 0.009545f
C726 B.n139 VSUBS 0.009545f
C727 B.n140 VSUBS 0.009545f
C728 B.n141 VSUBS 0.009545f
C729 B.n142 VSUBS 0.023497f
C730 B.n143 VSUBS 0.009545f
C731 B.n144 VSUBS 0.009545f
C732 B.n145 VSUBS 0.009545f
C733 B.n146 VSUBS 0.009545f
C734 B.n147 VSUBS 0.009545f
C735 B.n148 VSUBS 0.009545f
C736 B.n149 VSUBS 0.009545f
C737 B.n150 VSUBS 0.009545f
C738 B.n151 VSUBS 0.009545f
C739 B.n152 VSUBS 0.009545f
C740 B.n153 VSUBS 0.009545f
C741 B.n154 VSUBS 0.009545f
C742 B.n155 VSUBS 0.009545f
C743 B.t8 VSUBS 0.155052f
C744 B.t7 VSUBS 0.206435f
C745 B.t6 VSUBS 1.80719f
C746 B.n156 VSUBS 0.336623f
C747 B.n157 VSUBS 0.252585f
C748 B.n158 VSUBS 0.022115f
C749 B.n159 VSUBS 0.009545f
C750 B.n160 VSUBS 0.009545f
C751 B.n161 VSUBS 0.009545f
C752 B.n162 VSUBS 0.009545f
C753 B.n163 VSUBS 0.009545f
C754 B.t5 VSUBS 0.155049f
C755 B.t4 VSUBS 0.206432f
C756 B.t3 VSUBS 1.80719f
C757 B.n164 VSUBS 0.336625f
C758 B.n165 VSUBS 0.252588f
C759 B.n166 VSUBS 0.009545f
C760 B.n167 VSUBS 0.009545f
C761 B.n168 VSUBS 0.009545f
C762 B.n169 VSUBS 0.009545f
C763 B.n170 VSUBS 0.009545f
C764 B.n171 VSUBS 0.009545f
C765 B.n172 VSUBS 0.009545f
C766 B.n173 VSUBS 0.009545f
C767 B.n174 VSUBS 0.009545f
C768 B.n175 VSUBS 0.009545f
C769 B.n176 VSUBS 0.009545f
C770 B.n177 VSUBS 0.009545f
C771 B.n178 VSUBS 0.009545f
C772 B.n179 VSUBS 0.023497f
C773 B.n180 VSUBS 0.009545f
C774 B.n181 VSUBS 0.009545f
C775 B.n182 VSUBS 0.009545f
C776 B.n183 VSUBS 0.009545f
C777 B.n184 VSUBS 0.009545f
C778 B.n185 VSUBS 0.009545f
C779 B.n186 VSUBS 0.009545f
C780 B.n187 VSUBS 0.009545f
C781 B.n188 VSUBS 0.009545f
C782 B.n189 VSUBS 0.009545f
C783 B.n190 VSUBS 0.009545f
C784 B.n191 VSUBS 0.009545f
C785 B.n192 VSUBS 0.009545f
C786 B.n193 VSUBS 0.009545f
C787 B.n194 VSUBS 0.009545f
C788 B.n195 VSUBS 0.009545f
C789 B.n196 VSUBS 0.009545f
C790 B.n197 VSUBS 0.009545f
C791 B.n198 VSUBS 0.009545f
C792 B.n199 VSUBS 0.009545f
C793 B.n200 VSUBS 0.009545f
C794 B.n201 VSUBS 0.009545f
C795 B.n202 VSUBS 0.009545f
C796 B.n203 VSUBS 0.009545f
C797 B.n204 VSUBS 0.009545f
C798 B.n205 VSUBS 0.009545f
C799 B.n206 VSUBS 0.009545f
C800 B.n207 VSUBS 0.009545f
C801 B.n208 VSUBS 0.009545f
C802 B.n209 VSUBS 0.009545f
C803 B.n210 VSUBS 0.009545f
C804 B.n211 VSUBS 0.009545f
C805 B.n212 VSUBS 0.009545f
C806 B.n213 VSUBS 0.009545f
C807 B.n214 VSUBS 0.009545f
C808 B.n215 VSUBS 0.009545f
C809 B.n216 VSUBS 0.009545f
C810 B.n217 VSUBS 0.009545f
C811 B.n218 VSUBS 0.009545f
C812 B.n219 VSUBS 0.009545f
C813 B.n220 VSUBS 0.009545f
C814 B.n221 VSUBS 0.009545f
C815 B.n222 VSUBS 0.009545f
C816 B.n223 VSUBS 0.009545f
C817 B.n224 VSUBS 0.009545f
C818 B.n225 VSUBS 0.009545f
C819 B.n226 VSUBS 0.009545f
C820 B.n227 VSUBS 0.009545f
C821 B.n228 VSUBS 0.009545f
C822 B.n229 VSUBS 0.009545f
C823 B.n230 VSUBS 0.009545f
C824 B.n231 VSUBS 0.009545f
C825 B.n232 VSUBS 0.009545f
C826 B.n233 VSUBS 0.009545f
C827 B.n234 VSUBS 0.009545f
C828 B.n235 VSUBS 0.009545f
C829 B.n236 VSUBS 0.009545f
C830 B.n237 VSUBS 0.009545f
C831 B.n238 VSUBS 0.009545f
C832 B.n239 VSUBS 0.009545f
C833 B.n240 VSUBS 0.009545f
C834 B.n241 VSUBS 0.009545f
C835 B.n242 VSUBS 0.009545f
C836 B.n243 VSUBS 0.009545f
C837 B.n244 VSUBS 0.009545f
C838 B.n245 VSUBS 0.009545f
C839 B.n246 VSUBS 0.009545f
C840 B.n247 VSUBS 0.009545f
C841 B.n248 VSUBS 0.009545f
C842 B.n249 VSUBS 0.009545f
C843 B.n250 VSUBS 0.009545f
C844 B.n251 VSUBS 0.009545f
C845 B.n252 VSUBS 0.009545f
C846 B.n253 VSUBS 0.009545f
C847 B.n254 VSUBS 0.009545f
C848 B.n255 VSUBS 0.009545f
C849 B.n256 VSUBS 0.009545f
C850 B.n257 VSUBS 0.009545f
C851 B.n258 VSUBS 0.009545f
C852 B.n259 VSUBS 0.009545f
C853 B.n260 VSUBS 0.009545f
C854 B.n261 VSUBS 0.009545f
C855 B.n262 VSUBS 0.009545f
C856 B.n263 VSUBS 0.009545f
C857 B.n264 VSUBS 0.009545f
C858 B.n265 VSUBS 0.009545f
C859 B.n266 VSUBS 0.009545f
C860 B.n267 VSUBS 0.009545f
C861 B.n268 VSUBS 0.009545f
C862 B.n269 VSUBS 0.009545f
C863 B.n270 VSUBS 0.009545f
C864 B.n271 VSUBS 0.009545f
C865 B.n272 VSUBS 0.009545f
C866 B.n273 VSUBS 0.009545f
C867 B.n274 VSUBS 0.009545f
C868 B.n275 VSUBS 0.009545f
C869 B.n276 VSUBS 0.009545f
C870 B.n277 VSUBS 0.009545f
C871 B.n278 VSUBS 0.009545f
C872 B.n279 VSUBS 0.009545f
C873 B.n280 VSUBS 0.009545f
C874 B.n281 VSUBS 0.009545f
C875 B.n282 VSUBS 0.009545f
C876 B.n283 VSUBS 0.009545f
C877 B.n284 VSUBS 0.009545f
C878 B.n285 VSUBS 0.009545f
C879 B.n286 VSUBS 0.009545f
C880 B.n287 VSUBS 0.009545f
C881 B.n288 VSUBS 0.009545f
C882 B.n289 VSUBS 0.009545f
C883 B.n290 VSUBS 0.009545f
C884 B.n291 VSUBS 0.009545f
C885 B.n292 VSUBS 0.009545f
C886 B.n293 VSUBS 0.009545f
C887 B.n294 VSUBS 0.009545f
C888 B.n295 VSUBS 0.009545f
C889 B.n296 VSUBS 0.009545f
C890 B.n297 VSUBS 0.009545f
C891 B.n298 VSUBS 0.009545f
C892 B.n299 VSUBS 0.009545f
C893 B.n300 VSUBS 0.009545f
C894 B.n301 VSUBS 0.009545f
C895 B.n302 VSUBS 0.009545f
C896 B.n303 VSUBS 0.009545f
C897 B.n304 VSUBS 0.009545f
C898 B.n305 VSUBS 0.009545f
C899 B.n306 VSUBS 0.009545f
C900 B.n307 VSUBS 0.009545f
C901 B.n308 VSUBS 0.009545f
C902 B.n309 VSUBS 0.009545f
C903 B.n310 VSUBS 0.009545f
C904 B.n311 VSUBS 0.009545f
C905 B.n312 VSUBS 0.023497f
C906 B.n313 VSUBS 0.02451f
C907 B.n314 VSUBS 0.02451f
C908 B.n315 VSUBS 0.009545f
C909 B.n316 VSUBS 0.009545f
C910 B.n317 VSUBS 0.009545f
C911 B.n318 VSUBS 0.009545f
C912 B.n319 VSUBS 0.009545f
C913 B.n320 VSUBS 0.009545f
C914 B.n321 VSUBS 0.009545f
C915 B.n322 VSUBS 0.009545f
C916 B.n323 VSUBS 0.009545f
C917 B.n324 VSUBS 0.009545f
C918 B.n325 VSUBS 0.009545f
C919 B.n326 VSUBS 0.009545f
C920 B.n327 VSUBS 0.009545f
C921 B.n328 VSUBS 0.009545f
C922 B.n329 VSUBS 0.009545f
C923 B.n330 VSUBS 0.009545f
C924 B.n331 VSUBS 0.009545f
C925 B.n332 VSUBS 0.009545f
C926 B.n333 VSUBS 0.009545f
C927 B.n334 VSUBS 0.009545f
C928 B.n335 VSUBS 0.009545f
C929 B.n336 VSUBS 0.009545f
C930 B.n337 VSUBS 0.009545f
C931 B.n338 VSUBS 0.009545f
C932 B.n339 VSUBS 0.009545f
C933 B.n340 VSUBS 0.009545f
C934 B.n341 VSUBS 0.009545f
C935 B.n342 VSUBS 0.009545f
C936 B.n343 VSUBS 0.009545f
C937 B.n344 VSUBS 0.009545f
C938 B.n345 VSUBS 0.009545f
C939 B.n346 VSUBS 0.009545f
C940 B.n347 VSUBS 0.009545f
C941 B.n348 VSUBS 0.009545f
C942 B.n349 VSUBS 0.009545f
C943 B.n350 VSUBS 0.009545f
C944 B.n351 VSUBS 0.009545f
C945 B.n352 VSUBS 0.009545f
C946 B.n353 VSUBS 0.009545f
C947 B.n354 VSUBS 0.006597f
C948 B.n355 VSUBS 0.022115f
C949 B.n356 VSUBS 0.00772f
C950 B.n357 VSUBS 0.009545f
C951 B.n358 VSUBS 0.009545f
C952 B.n359 VSUBS 0.009545f
C953 B.n360 VSUBS 0.009545f
C954 B.n361 VSUBS 0.009545f
C955 B.n362 VSUBS 0.009545f
C956 B.n363 VSUBS 0.009545f
C957 B.n364 VSUBS 0.009545f
C958 B.n365 VSUBS 0.009545f
C959 B.n366 VSUBS 0.009545f
C960 B.n367 VSUBS 0.009545f
C961 B.n368 VSUBS 0.00772f
C962 B.n369 VSUBS 0.009545f
C963 B.n370 VSUBS 0.009545f
C964 B.n371 VSUBS 0.006597f
C965 B.n372 VSUBS 0.009545f
C966 B.n373 VSUBS 0.009545f
C967 B.n374 VSUBS 0.009545f
C968 B.n375 VSUBS 0.009545f
C969 B.n376 VSUBS 0.009545f
C970 B.n377 VSUBS 0.009545f
C971 B.n378 VSUBS 0.009545f
C972 B.n379 VSUBS 0.009545f
C973 B.n380 VSUBS 0.009545f
C974 B.n381 VSUBS 0.009545f
C975 B.n382 VSUBS 0.009545f
C976 B.n383 VSUBS 0.009545f
C977 B.n384 VSUBS 0.009545f
C978 B.n385 VSUBS 0.009545f
C979 B.n386 VSUBS 0.009545f
C980 B.n387 VSUBS 0.009545f
C981 B.n388 VSUBS 0.009545f
C982 B.n389 VSUBS 0.009545f
C983 B.n390 VSUBS 0.009545f
C984 B.n391 VSUBS 0.009545f
C985 B.n392 VSUBS 0.009545f
C986 B.n393 VSUBS 0.009545f
C987 B.n394 VSUBS 0.009545f
C988 B.n395 VSUBS 0.009545f
C989 B.n396 VSUBS 0.009545f
C990 B.n397 VSUBS 0.009545f
C991 B.n398 VSUBS 0.009545f
C992 B.n399 VSUBS 0.009545f
C993 B.n400 VSUBS 0.009545f
C994 B.n401 VSUBS 0.009545f
C995 B.n402 VSUBS 0.009545f
C996 B.n403 VSUBS 0.009545f
C997 B.n404 VSUBS 0.009545f
C998 B.n405 VSUBS 0.009545f
C999 B.n406 VSUBS 0.009545f
C1000 B.n407 VSUBS 0.009545f
C1001 B.n408 VSUBS 0.009545f
C1002 B.n409 VSUBS 0.009545f
C1003 B.n410 VSUBS 0.009545f
C1004 B.n411 VSUBS 0.02451f
C1005 B.n412 VSUBS 0.023497f
C1006 B.n413 VSUBS 0.02451f
C1007 B.n414 VSUBS 0.009545f
C1008 B.n415 VSUBS 0.009545f
C1009 B.n416 VSUBS 0.009545f
C1010 B.n417 VSUBS 0.009545f
C1011 B.n418 VSUBS 0.009545f
C1012 B.n419 VSUBS 0.009545f
C1013 B.n420 VSUBS 0.009545f
C1014 B.n421 VSUBS 0.009545f
C1015 B.n422 VSUBS 0.009545f
C1016 B.n423 VSUBS 0.009545f
C1017 B.n424 VSUBS 0.009545f
C1018 B.n425 VSUBS 0.009545f
C1019 B.n426 VSUBS 0.009545f
C1020 B.n427 VSUBS 0.009545f
C1021 B.n428 VSUBS 0.009545f
C1022 B.n429 VSUBS 0.009545f
C1023 B.n430 VSUBS 0.009545f
C1024 B.n431 VSUBS 0.009545f
C1025 B.n432 VSUBS 0.009545f
C1026 B.n433 VSUBS 0.009545f
C1027 B.n434 VSUBS 0.009545f
C1028 B.n435 VSUBS 0.009545f
C1029 B.n436 VSUBS 0.009545f
C1030 B.n437 VSUBS 0.009545f
C1031 B.n438 VSUBS 0.009545f
C1032 B.n439 VSUBS 0.009545f
C1033 B.n440 VSUBS 0.009545f
C1034 B.n441 VSUBS 0.009545f
C1035 B.n442 VSUBS 0.009545f
C1036 B.n443 VSUBS 0.009545f
C1037 B.n444 VSUBS 0.009545f
C1038 B.n445 VSUBS 0.009545f
C1039 B.n446 VSUBS 0.009545f
C1040 B.n447 VSUBS 0.009545f
C1041 B.n448 VSUBS 0.009545f
C1042 B.n449 VSUBS 0.009545f
C1043 B.n450 VSUBS 0.009545f
C1044 B.n451 VSUBS 0.009545f
C1045 B.n452 VSUBS 0.009545f
C1046 B.n453 VSUBS 0.009545f
C1047 B.n454 VSUBS 0.009545f
C1048 B.n455 VSUBS 0.009545f
C1049 B.n456 VSUBS 0.009545f
C1050 B.n457 VSUBS 0.009545f
C1051 B.n458 VSUBS 0.009545f
C1052 B.n459 VSUBS 0.009545f
C1053 B.n460 VSUBS 0.009545f
C1054 B.n461 VSUBS 0.009545f
C1055 B.n462 VSUBS 0.009545f
C1056 B.n463 VSUBS 0.009545f
C1057 B.n464 VSUBS 0.009545f
C1058 B.n465 VSUBS 0.009545f
C1059 B.n466 VSUBS 0.009545f
C1060 B.n467 VSUBS 0.009545f
C1061 B.n468 VSUBS 0.009545f
C1062 B.n469 VSUBS 0.009545f
C1063 B.n470 VSUBS 0.009545f
C1064 B.n471 VSUBS 0.009545f
C1065 B.n472 VSUBS 0.009545f
C1066 B.n473 VSUBS 0.009545f
C1067 B.n474 VSUBS 0.009545f
C1068 B.n475 VSUBS 0.009545f
C1069 B.n476 VSUBS 0.009545f
C1070 B.n477 VSUBS 0.009545f
C1071 B.n478 VSUBS 0.009545f
C1072 B.n479 VSUBS 0.009545f
C1073 B.n480 VSUBS 0.009545f
C1074 B.n481 VSUBS 0.009545f
C1075 B.n482 VSUBS 0.009545f
C1076 B.n483 VSUBS 0.009545f
C1077 B.n484 VSUBS 0.009545f
C1078 B.n485 VSUBS 0.009545f
C1079 B.n486 VSUBS 0.009545f
C1080 B.n487 VSUBS 0.009545f
C1081 B.n488 VSUBS 0.009545f
C1082 B.n489 VSUBS 0.009545f
C1083 B.n490 VSUBS 0.009545f
C1084 B.n491 VSUBS 0.009545f
C1085 B.n492 VSUBS 0.009545f
C1086 B.n493 VSUBS 0.009545f
C1087 B.n494 VSUBS 0.009545f
C1088 B.n495 VSUBS 0.009545f
C1089 B.n496 VSUBS 0.009545f
C1090 B.n497 VSUBS 0.009545f
C1091 B.n498 VSUBS 0.009545f
C1092 B.n499 VSUBS 0.009545f
C1093 B.n500 VSUBS 0.009545f
C1094 B.n501 VSUBS 0.009545f
C1095 B.n502 VSUBS 0.009545f
C1096 B.n503 VSUBS 0.009545f
C1097 B.n504 VSUBS 0.009545f
C1098 B.n505 VSUBS 0.009545f
C1099 B.n506 VSUBS 0.009545f
C1100 B.n507 VSUBS 0.009545f
C1101 B.n508 VSUBS 0.009545f
C1102 B.n509 VSUBS 0.009545f
C1103 B.n510 VSUBS 0.009545f
C1104 B.n511 VSUBS 0.009545f
C1105 B.n512 VSUBS 0.009545f
C1106 B.n513 VSUBS 0.009545f
C1107 B.n514 VSUBS 0.009545f
C1108 B.n515 VSUBS 0.009545f
C1109 B.n516 VSUBS 0.009545f
C1110 B.n517 VSUBS 0.009545f
C1111 B.n518 VSUBS 0.009545f
C1112 B.n519 VSUBS 0.009545f
C1113 B.n520 VSUBS 0.009545f
C1114 B.n521 VSUBS 0.009545f
C1115 B.n522 VSUBS 0.009545f
C1116 B.n523 VSUBS 0.009545f
C1117 B.n524 VSUBS 0.009545f
C1118 B.n525 VSUBS 0.009545f
C1119 B.n526 VSUBS 0.009545f
C1120 B.n527 VSUBS 0.009545f
C1121 B.n528 VSUBS 0.009545f
C1122 B.n529 VSUBS 0.009545f
C1123 B.n530 VSUBS 0.009545f
C1124 B.n531 VSUBS 0.009545f
C1125 B.n532 VSUBS 0.009545f
C1126 B.n533 VSUBS 0.009545f
C1127 B.n534 VSUBS 0.009545f
C1128 B.n535 VSUBS 0.009545f
C1129 B.n536 VSUBS 0.009545f
C1130 B.n537 VSUBS 0.009545f
C1131 B.n538 VSUBS 0.009545f
C1132 B.n539 VSUBS 0.009545f
C1133 B.n540 VSUBS 0.009545f
C1134 B.n541 VSUBS 0.009545f
C1135 B.n542 VSUBS 0.009545f
C1136 B.n543 VSUBS 0.009545f
C1137 B.n544 VSUBS 0.009545f
C1138 B.n545 VSUBS 0.009545f
C1139 B.n546 VSUBS 0.009545f
C1140 B.n547 VSUBS 0.009545f
C1141 B.n548 VSUBS 0.009545f
C1142 B.n549 VSUBS 0.009545f
C1143 B.n550 VSUBS 0.009545f
C1144 B.n551 VSUBS 0.009545f
C1145 B.n552 VSUBS 0.009545f
C1146 B.n553 VSUBS 0.009545f
C1147 B.n554 VSUBS 0.009545f
C1148 B.n555 VSUBS 0.009545f
C1149 B.n556 VSUBS 0.009545f
C1150 B.n557 VSUBS 0.009545f
C1151 B.n558 VSUBS 0.009545f
C1152 B.n559 VSUBS 0.009545f
C1153 B.n560 VSUBS 0.009545f
C1154 B.n561 VSUBS 0.009545f
C1155 B.n562 VSUBS 0.009545f
C1156 B.n563 VSUBS 0.009545f
C1157 B.n564 VSUBS 0.009545f
C1158 B.n565 VSUBS 0.009545f
C1159 B.n566 VSUBS 0.009545f
C1160 B.n567 VSUBS 0.009545f
C1161 B.n568 VSUBS 0.009545f
C1162 B.n569 VSUBS 0.009545f
C1163 B.n570 VSUBS 0.009545f
C1164 B.n571 VSUBS 0.009545f
C1165 B.n572 VSUBS 0.009545f
C1166 B.n573 VSUBS 0.009545f
C1167 B.n574 VSUBS 0.009545f
C1168 B.n575 VSUBS 0.009545f
C1169 B.n576 VSUBS 0.009545f
C1170 B.n577 VSUBS 0.009545f
C1171 B.n578 VSUBS 0.009545f
C1172 B.n579 VSUBS 0.009545f
C1173 B.n580 VSUBS 0.009545f
C1174 B.n581 VSUBS 0.009545f
C1175 B.n582 VSUBS 0.009545f
C1176 B.n583 VSUBS 0.009545f
C1177 B.n584 VSUBS 0.009545f
C1178 B.n585 VSUBS 0.009545f
C1179 B.n586 VSUBS 0.009545f
C1180 B.n587 VSUBS 0.009545f
C1181 B.n588 VSUBS 0.009545f
C1182 B.n589 VSUBS 0.009545f
C1183 B.n590 VSUBS 0.009545f
C1184 B.n591 VSUBS 0.009545f
C1185 B.n592 VSUBS 0.009545f
C1186 B.n593 VSUBS 0.009545f
C1187 B.n594 VSUBS 0.009545f
C1188 B.n595 VSUBS 0.009545f
C1189 B.n596 VSUBS 0.009545f
C1190 B.n597 VSUBS 0.009545f
C1191 B.n598 VSUBS 0.009545f
C1192 B.n599 VSUBS 0.009545f
C1193 B.n600 VSUBS 0.009545f
C1194 B.n601 VSUBS 0.009545f
C1195 B.n602 VSUBS 0.009545f
C1196 B.n603 VSUBS 0.009545f
C1197 B.n604 VSUBS 0.009545f
C1198 B.n605 VSUBS 0.009545f
C1199 B.n606 VSUBS 0.009545f
C1200 B.n607 VSUBS 0.009545f
C1201 B.n608 VSUBS 0.009545f
C1202 B.n609 VSUBS 0.009545f
C1203 B.n610 VSUBS 0.009545f
C1204 B.n611 VSUBS 0.009545f
C1205 B.n612 VSUBS 0.009545f
C1206 B.n613 VSUBS 0.009545f
C1207 B.n614 VSUBS 0.009545f
C1208 B.n615 VSUBS 0.009545f
C1209 B.n616 VSUBS 0.009545f
C1210 B.n617 VSUBS 0.009545f
C1211 B.n618 VSUBS 0.023497f
C1212 B.n619 VSUBS 0.02451f
C1213 B.n620 VSUBS 0.02451f
C1214 B.n621 VSUBS 0.009545f
C1215 B.n622 VSUBS 0.009545f
C1216 B.n623 VSUBS 0.009545f
C1217 B.n624 VSUBS 0.009545f
C1218 B.n625 VSUBS 0.009545f
C1219 B.n626 VSUBS 0.009545f
C1220 B.n627 VSUBS 0.009545f
C1221 B.n628 VSUBS 0.009545f
C1222 B.n629 VSUBS 0.009545f
C1223 B.n630 VSUBS 0.009545f
C1224 B.n631 VSUBS 0.009545f
C1225 B.n632 VSUBS 0.009545f
C1226 B.n633 VSUBS 0.009545f
C1227 B.n634 VSUBS 0.009545f
C1228 B.n635 VSUBS 0.009545f
C1229 B.n636 VSUBS 0.009545f
C1230 B.n637 VSUBS 0.009545f
C1231 B.n638 VSUBS 0.009545f
C1232 B.n639 VSUBS 0.009545f
C1233 B.n640 VSUBS 0.009545f
C1234 B.n641 VSUBS 0.009545f
C1235 B.n642 VSUBS 0.009545f
C1236 B.n643 VSUBS 0.009545f
C1237 B.n644 VSUBS 0.009545f
C1238 B.n645 VSUBS 0.009545f
C1239 B.n646 VSUBS 0.009545f
C1240 B.n647 VSUBS 0.009545f
C1241 B.n648 VSUBS 0.009545f
C1242 B.n649 VSUBS 0.009545f
C1243 B.n650 VSUBS 0.009545f
C1244 B.n651 VSUBS 0.009545f
C1245 B.n652 VSUBS 0.009545f
C1246 B.n653 VSUBS 0.009545f
C1247 B.n654 VSUBS 0.009545f
C1248 B.n655 VSUBS 0.009545f
C1249 B.n656 VSUBS 0.009545f
C1250 B.n657 VSUBS 0.009545f
C1251 B.n658 VSUBS 0.009545f
C1252 B.n659 VSUBS 0.009545f
C1253 B.n660 VSUBS 0.006597f
C1254 B.n661 VSUBS 0.022115f
C1255 B.n662 VSUBS 0.00772f
C1256 B.n663 VSUBS 0.009545f
C1257 B.n664 VSUBS 0.009545f
C1258 B.n665 VSUBS 0.009545f
C1259 B.n666 VSUBS 0.009545f
C1260 B.n667 VSUBS 0.009545f
C1261 B.n668 VSUBS 0.009545f
C1262 B.n669 VSUBS 0.009545f
C1263 B.n670 VSUBS 0.009545f
C1264 B.n671 VSUBS 0.009545f
C1265 B.n672 VSUBS 0.009545f
C1266 B.n673 VSUBS 0.009545f
C1267 B.n674 VSUBS 0.00772f
C1268 B.n675 VSUBS 0.009545f
C1269 B.n676 VSUBS 0.009545f
C1270 B.n677 VSUBS 0.006597f
C1271 B.n678 VSUBS 0.009545f
C1272 B.n679 VSUBS 0.009545f
C1273 B.n680 VSUBS 0.009545f
C1274 B.n681 VSUBS 0.009545f
C1275 B.n682 VSUBS 0.009545f
C1276 B.n683 VSUBS 0.009545f
C1277 B.n684 VSUBS 0.009545f
C1278 B.n685 VSUBS 0.009545f
C1279 B.n686 VSUBS 0.009545f
C1280 B.n687 VSUBS 0.009545f
C1281 B.n688 VSUBS 0.009545f
C1282 B.n689 VSUBS 0.009545f
C1283 B.n690 VSUBS 0.009545f
C1284 B.n691 VSUBS 0.009545f
C1285 B.n692 VSUBS 0.009545f
C1286 B.n693 VSUBS 0.009545f
C1287 B.n694 VSUBS 0.009545f
C1288 B.n695 VSUBS 0.009545f
C1289 B.n696 VSUBS 0.009545f
C1290 B.n697 VSUBS 0.009545f
C1291 B.n698 VSUBS 0.009545f
C1292 B.n699 VSUBS 0.009545f
C1293 B.n700 VSUBS 0.009545f
C1294 B.n701 VSUBS 0.009545f
C1295 B.n702 VSUBS 0.009545f
C1296 B.n703 VSUBS 0.009545f
C1297 B.n704 VSUBS 0.009545f
C1298 B.n705 VSUBS 0.009545f
C1299 B.n706 VSUBS 0.009545f
C1300 B.n707 VSUBS 0.009545f
C1301 B.n708 VSUBS 0.009545f
C1302 B.n709 VSUBS 0.009545f
C1303 B.n710 VSUBS 0.009545f
C1304 B.n711 VSUBS 0.009545f
C1305 B.n712 VSUBS 0.009545f
C1306 B.n713 VSUBS 0.009545f
C1307 B.n714 VSUBS 0.009545f
C1308 B.n715 VSUBS 0.009545f
C1309 B.n716 VSUBS 0.009545f
C1310 B.n717 VSUBS 0.02451f
C1311 B.n718 VSUBS 0.023497f
C1312 B.n719 VSUBS 0.023497f
C1313 B.n720 VSUBS 0.009545f
C1314 B.n721 VSUBS 0.009545f
C1315 B.n722 VSUBS 0.009545f
C1316 B.n723 VSUBS 0.009545f
C1317 B.n724 VSUBS 0.009545f
C1318 B.n725 VSUBS 0.009545f
C1319 B.n726 VSUBS 0.009545f
C1320 B.n727 VSUBS 0.009545f
C1321 B.n728 VSUBS 0.009545f
C1322 B.n729 VSUBS 0.009545f
C1323 B.n730 VSUBS 0.009545f
C1324 B.n731 VSUBS 0.009545f
C1325 B.n732 VSUBS 0.009545f
C1326 B.n733 VSUBS 0.009545f
C1327 B.n734 VSUBS 0.009545f
C1328 B.n735 VSUBS 0.009545f
C1329 B.n736 VSUBS 0.009545f
C1330 B.n737 VSUBS 0.009545f
C1331 B.n738 VSUBS 0.009545f
C1332 B.n739 VSUBS 0.009545f
C1333 B.n740 VSUBS 0.009545f
C1334 B.n741 VSUBS 0.009545f
C1335 B.n742 VSUBS 0.009545f
C1336 B.n743 VSUBS 0.009545f
C1337 B.n744 VSUBS 0.009545f
C1338 B.n745 VSUBS 0.009545f
C1339 B.n746 VSUBS 0.009545f
C1340 B.n747 VSUBS 0.009545f
C1341 B.n748 VSUBS 0.009545f
C1342 B.n749 VSUBS 0.009545f
C1343 B.n750 VSUBS 0.009545f
C1344 B.n751 VSUBS 0.009545f
C1345 B.n752 VSUBS 0.009545f
C1346 B.n753 VSUBS 0.009545f
C1347 B.n754 VSUBS 0.009545f
C1348 B.n755 VSUBS 0.009545f
C1349 B.n756 VSUBS 0.009545f
C1350 B.n757 VSUBS 0.009545f
C1351 B.n758 VSUBS 0.009545f
C1352 B.n759 VSUBS 0.009545f
C1353 B.n760 VSUBS 0.009545f
C1354 B.n761 VSUBS 0.009545f
C1355 B.n762 VSUBS 0.009545f
C1356 B.n763 VSUBS 0.009545f
C1357 B.n764 VSUBS 0.009545f
C1358 B.n765 VSUBS 0.009545f
C1359 B.n766 VSUBS 0.009545f
C1360 B.n767 VSUBS 0.009545f
C1361 B.n768 VSUBS 0.009545f
C1362 B.n769 VSUBS 0.009545f
C1363 B.n770 VSUBS 0.009545f
C1364 B.n771 VSUBS 0.009545f
C1365 B.n772 VSUBS 0.009545f
C1366 B.n773 VSUBS 0.009545f
C1367 B.n774 VSUBS 0.009545f
C1368 B.n775 VSUBS 0.009545f
C1369 B.n776 VSUBS 0.009545f
C1370 B.n777 VSUBS 0.009545f
C1371 B.n778 VSUBS 0.009545f
C1372 B.n779 VSUBS 0.009545f
C1373 B.n780 VSUBS 0.009545f
C1374 B.n781 VSUBS 0.009545f
C1375 B.n782 VSUBS 0.009545f
C1376 B.n783 VSUBS 0.009545f
C1377 B.n784 VSUBS 0.009545f
C1378 B.n785 VSUBS 0.009545f
C1379 B.n786 VSUBS 0.009545f
C1380 B.n787 VSUBS 0.009545f
C1381 B.n788 VSUBS 0.009545f
C1382 B.n789 VSUBS 0.009545f
C1383 B.n790 VSUBS 0.009545f
C1384 B.n791 VSUBS 0.009545f
C1385 B.n792 VSUBS 0.009545f
C1386 B.n793 VSUBS 0.009545f
C1387 B.n794 VSUBS 0.009545f
C1388 B.n795 VSUBS 0.009545f
C1389 B.n796 VSUBS 0.009545f
C1390 B.n797 VSUBS 0.009545f
C1391 B.n798 VSUBS 0.009545f
C1392 B.n799 VSUBS 0.009545f
C1393 B.n800 VSUBS 0.009545f
C1394 B.n801 VSUBS 0.009545f
C1395 B.n802 VSUBS 0.009545f
C1396 B.n803 VSUBS 0.009545f
C1397 B.n804 VSUBS 0.009545f
C1398 B.n805 VSUBS 0.009545f
C1399 B.n806 VSUBS 0.009545f
C1400 B.n807 VSUBS 0.009545f
C1401 B.n808 VSUBS 0.009545f
C1402 B.n809 VSUBS 0.009545f
C1403 B.n810 VSUBS 0.009545f
C1404 B.n811 VSUBS 0.009545f
C1405 B.n812 VSUBS 0.009545f
C1406 B.n813 VSUBS 0.009545f
C1407 B.n814 VSUBS 0.009545f
C1408 B.n815 VSUBS 0.009545f
C1409 B.n816 VSUBS 0.009545f
C1410 B.n817 VSUBS 0.009545f
C1411 B.n818 VSUBS 0.009545f
C1412 B.n819 VSUBS 0.012456f
C1413 B.n820 VSUBS 0.013269f
C1414 B.n821 VSUBS 0.026386f
.ends

