* NGSPICE file created from diff_pair_sample_1332.ext - technology: sky130A

.subckt diff_pair_sample_1332 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3946 pd=13.06 as=1.0131 ps=6.47 w=6.14 l=3.32
X1 VDD1.t9 VP.t0 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X2 VDD2.t8 VN.t1 VTAIL.t16 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3946 pd=13.06 as=1.0131 ps=6.47 w=6.14 l=3.32
X3 VDD1.t8 VP.t1 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X4 VTAIL.t14 VN.t2 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X5 VDD1.t7 VP.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.3946 pd=13.06 as=1.0131 ps=6.47 w=6.14 l=3.32
X6 VDD1.t6 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.3946 pd=13.06 as=1.0131 ps=6.47 w=6.14 l=3.32
X7 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=2.3946 pd=13.06 as=0 ps=0 w=6.14 l=3.32
X8 VTAIL.t2 VP.t4 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X9 VTAIL.t3 VP.t5 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X10 VDD2.t6 VN.t3 VTAIL.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X11 VDD2.t5 VN.t4 VTAIL.t19 B.t8 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X12 VTAIL.t7 VP.t6 VDD1.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X13 VDD1.t2 VP.t7 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=2.3946 ps=13.06 w=6.14 l=3.32
X14 VTAIL.t1 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X15 VDD2.t4 VN.t5 VTAIL.t18 B.t6 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=2.3946 ps=13.06 w=6.14 l=3.32
X16 VDD1.t0 VP.t9 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=2.3946 ps=13.06 w=6.14 l=3.32
X17 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=2.3946 pd=13.06 as=0 ps=0 w=6.14 l=3.32
X18 VDD2.t3 VN.t6 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=2.3946 ps=13.06 w=6.14 l=3.32
X19 VTAIL.t17 VN.t7 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X20 VTAIL.t10 VN.t8 VDD2.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X21 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.3946 pd=13.06 as=0 ps=0 w=6.14 l=3.32
X22 VTAIL.t15 VN.t9 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=1.0131 pd=6.47 as=1.0131 ps=6.47 w=6.14 l=3.32
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.3946 pd=13.06 as=0 ps=0 w=6.14 l=3.32
R0 VN.n96 VN.n95 161.3
R1 VN.n94 VN.n50 161.3
R2 VN.n93 VN.n92 161.3
R3 VN.n91 VN.n51 161.3
R4 VN.n90 VN.n89 161.3
R5 VN.n88 VN.n52 161.3
R6 VN.n87 VN.n86 161.3
R7 VN.n85 VN.n84 161.3
R8 VN.n83 VN.n54 161.3
R9 VN.n82 VN.n81 161.3
R10 VN.n80 VN.n55 161.3
R11 VN.n79 VN.n78 161.3
R12 VN.n77 VN.n56 161.3
R13 VN.n76 VN.n75 161.3
R14 VN.n74 VN.n57 161.3
R15 VN.n73 VN.n72 161.3
R16 VN.n71 VN.n58 161.3
R17 VN.n70 VN.n69 161.3
R18 VN.n68 VN.n59 161.3
R19 VN.n67 VN.n66 161.3
R20 VN.n65 VN.n60 161.3
R21 VN.n64 VN.n63 161.3
R22 VN.n47 VN.n46 161.3
R23 VN.n45 VN.n1 161.3
R24 VN.n44 VN.n43 161.3
R25 VN.n42 VN.n2 161.3
R26 VN.n41 VN.n40 161.3
R27 VN.n39 VN.n3 161.3
R28 VN.n38 VN.n37 161.3
R29 VN.n36 VN.n35 161.3
R30 VN.n34 VN.n5 161.3
R31 VN.n33 VN.n32 161.3
R32 VN.n31 VN.n6 161.3
R33 VN.n30 VN.n29 161.3
R34 VN.n28 VN.n7 161.3
R35 VN.n27 VN.n26 161.3
R36 VN.n25 VN.n8 161.3
R37 VN.n24 VN.n23 161.3
R38 VN.n22 VN.n9 161.3
R39 VN.n21 VN.n20 161.3
R40 VN.n19 VN.n10 161.3
R41 VN.n18 VN.n17 161.3
R42 VN.n16 VN.n11 161.3
R43 VN.n15 VN.n14 161.3
R44 VN.n62 VN.t5 77.5432
R45 VN.n13 VN.t1 77.5432
R46 VN.n48 VN.n0 75.4905
R47 VN.n97 VN.n49 75.4905
R48 VN.n62 VN.n61 67.3352
R49 VN.n13 VN.n12 67.3352
R50 VN.n21 VN.n10 56.5617
R51 VN.n29 VN.n6 56.5617
R52 VN.n70 VN.n59 56.5617
R53 VN.n78 VN.n55 56.5617
R54 VN VN.n97 52.8731
R55 VN.n8 VN.t3 44.571
R56 VN.n12 VN.t7 44.571
R57 VN.n4 VN.t9 44.571
R58 VN.n0 VN.t6 44.571
R59 VN.n57 VN.t4 44.571
R60 VN.n61 VN.t8 44.571
R61 VN.n53 VN.t2 44.571
R62 VN.n49 VN.t0 44.571
R63 VN.n40 VN.n2 42.999
R64 VN.n89 VN.n51 42.999
R65 VN.n44 VN.n2 38.1551
R66 VN.n93 VN.n51 38.1551
R67 VN.n16 VN.n15 24.5923
R68 VN.n17 VN.n16 24.5923
R69 VN.n17 VN.n10 24.5923
R70 VN.n22 VN.n21 24.5923
R71 VN.n23 VN.n22 24.5923
R72 VN.n23 VN.n8 24.5923
R73 VN.n27 VN.n8 24.5923
R74 VN.n28 VN.n27 24.5923
R75 VN.n29 VN.n28 24.5923
R76 VN.n33 VN.n6 24.5923
R77 VN.n34 VN.n33 24.5923
R78 VN.n35 VN.n34 24.5923
R79 VN.n39 VN.n38 24.5923
R80 VN.n40 VN.n39 24.5923
R81 VN.n45 VN.n44 24.5923
R82 VN.n46 VN.n45 24.5923
R83 VN.n66 VN.n59 24.5923
R84 VN.n66 VN.n65 24.5923
R85 VN.n65 VN.n64 24.5923
R86 VN.n78 VN.n77 24.5923
R87 VN.n77 VN.n76 24.5923
R88 VN.n76 VN.n57 24.5923
R89 VN.n72 VN.n57 24.5923
R90 VN.n72 VN.n71 24.5923
R91 VN.n71 VN.n70 24.5923
R92 VN.n89 VN.n88 24.5923
R93 VN.n88 VN.n87 24.5923
R94 VN.n84 VN.n83 24.5923
R95 VN.n83 VN.n82 24.5923
R96 VN.n82 VN.n55 24.5923
R97 VN.n95 VN.n94 24.5923
R98 VN.n94 VN.n93 24.5923
R99 VN.n38 VN.n4 17.2148
R100 VN.n87 VN.n53 17.2148
R101 VN.n46 VN.n0 14.7556
R102 VN.n95 VN.n49 14.7556
R103 VN.n15 VN.n12 7.37805
R104 VN.n35 VN.n4 7.37805
R105 VN.n64 VN.n61 7.37805
R106 VN.n84 VN.n53 7.37805
R107 VN.n63 VN.n62 4.1475
R108 VN.n14 VN.n13 4.1475
R109 VN.n97 VN.n96 0.354861
R110 VN.n48 VN.n47 0.354861
R111 VN VN.n48 0.267071
R112 VN.n96 VN.n50 0.189894
R113 VN.n92 VN.n50 0.189894
R114 VN.n92 VN.n91 0.189894
R115 VN.n91 VN.n90 0.189894
R116 VN.n90 VN.n52 0.189894
R117 VN.n86 VN.n52 0.189894
R118 VN.n86 VN.n85 0.189894
R119 VN.n85 VN.n54 0.189894
R120 VN.n81 VN.n54 0.189894
R121 VN.n81 VN.n80 0.189894
R122 VN.n80 VN.n79 0.189894
R123 VN.n79 VN.n56 0.189894
R124 VN.n75 VN.n56 0.189894
R125 VN.n75 VN.n74 0.189894
R126 VN.n74 VN.n73 0.189894
R127 VN.n73 VN.n58 0.189894
R128 VN.n69 VN.n58 0.189894
R129 VN.n69 VN.n68 0.189894
R130 VN.n68 VN.n67 0.189894
R131 VN.n67 VN.n60 0.189894
R132 VN.n63 VN.n60 0.189894
R133 VN.n14 VN.n11 0.189894
R134 VN.n18 VN.n11 0.189894
R135 VN.n19 VN.n18 0.189894
R136 VN.n20 VN.n19 0.189894
R137 VN.n20 VN.n9 0.189894
R138 VN.n24 VN.n9 0.189894
R139 VN.n25 VN.n24 0.189894
R140 VN.n26 VN.n25 0.189894
R141 VN.n26 VN.n7 0.189894
R142 VN.n30 VN.n7 0.189894
R143 VN.n31 VN.n30 0.189894
R144 VN.n32 VN.n31 0.189894
R145 VN.n32 VN.n5 0.189894
R146 VN.n36 VN.n5 0.189894
R147 VN.n37 VN.n36 0.189894
R148 VN.n37 VN.n3 0.189894
R149 VN.n41 VN.n3 0.189894
R150 VN.n42 VN.n41 0.189894
R151 VN.n43 VN.n42 0.189894
R152 VN.n43 VN.n1 0.189894
R153 VN.n47 VN.n1 0.189894
R154 VTAIL.n11 VTAIL.t18 55.1232
R155 VTAIL.n16 VTAIL.t5 55.1222
R156 VTAIL.n17 VTAIL.t11 55.1222
R157 VTAIL.n2 VTAIL.t6 55.1222
R158 VTAIL.n15 VTAIL.n14 51.8984
R159 VTAIL.n13 VTAIL.n12 51.8984
R160 VTAIL.n10 VTAIL.n9 51.8984
R161 VTAIL.n8 VTAIL.n7 51.8984
R162 VTAIL.n19 VTAIL.n18 51.8983
R163 VTAIL.n1 VTAIL.n0 51.8983
R164 VTAIL.n4 VTAIL.n3 51.8983
R165 VTAIL.n6 VTAIL.n5 51.8983
R166 VTAIL.n8 VTAIL.n6 23.9531
R167 VTAIL.n17 VTAIL.n16 20.8065
R168 VTAIL.n18 VTAIL.t13 3.22526
R169 VTAIL.n18 VTAIL.t15 3.22526
R170 VTAIL.n0 VTAIL.t16 3.22526
R171 VTAIL.n0 VTAIL.t17 3.22526
R172 VTAIL.n3 VTAIL.t8 3.22526
R173 VTAIL.n3 VTAIL.t7 3.22526
R174 VTAIL.n5 VTAIL.t0 3.22526
R175 VTAIL.n5 VTAIL.t1 3.22526
R176 VTAIL.n14 VTAIL.t9 3.22526
R177 VTAIL.n14 VTAIL.t2 3.22526
R178 VTAIL.n12 VTAIL.t4 3.22526
R179 VTAIL.n12 VTAIL.t3 3.22526
R180 VTAIL.n9 VTAIL.t19 3.22526
R181 VTAIL.n9 VTAIL.t10 3.22526
R182 VTAIL.n7 VTAIL.t12 3.22526
R183 VTAIL.n7 VTAIL.t14 3.22526
R184 VTAIL.n10 VTAIL.n8 3.14705
R185 VTAIL.n11 VTAIL.n10 3.14705
R186 VTAIL.n15 VTAIL.n13 3.14705
R187 VTAIL.n16 VTAIL.n15 3.14705
R188 VTAIL.n6 VTAIL.n4 3.14705
R189 VTAIL.n4 VTAIL.n2 3.14705
R190 VTAIL.n19 VTAIL.n17 3.14705
R191 VTAIL VTAIL.n1 2.4186
R192 VTAIL.n13 VTAIL.n11 2.0436
R193 VTAIL.n2 VTAIL.n1 2.0436
R194 VTAIL VTAIL.n19 0.728948
R195 VDD2.n1 VDD2.t8 74.9475
R196 VDD2.n4 VDD2.t9 71.802
R197 VDD2.n3 VDD2.n2 70.8816
R198 VDD2 VDD2.n7 70.878
R199 VDD2.n6 VDD2.n5 68.5772
R200 VDD2.n1 VDD2.n0 68.5771
R201 VDD2.n4 VDD2.n3 43.9545
R202 VDD2.n7 VDD2.t1 3.22526
R203 VDD2.n7 VDD2.t4 3.22526
R204 VDD2.n5 VDD2.t7 3.22526
R205 VDD2.n5 VDD2.t5 3.22526
R206 VDD2.n2 VDD2.t0 3.22526
R207 VDD2.n2 VDD2.t3 3.22526
R208 VDD2.n0 VDD2.t2 3.22526
R209 VDD2.n0 VDD2.t6 3.22526
R210 VDD2.n6 VDD2.n4 3.14705
R211 VDD2 VDD2.n6 0.845328
R212 VDD2.n3 VDD2.n1 0.731792
R213 B.n881 B.n880 585
R214 B.n278 B.n161 585
R215 B.n277 B.n276 585
R216 B.n275 B.n274 585
R217 B.n273 B.n272 585
R218 B.n271 B.n270 585
R219 B.n269 B.n268 585
R220 B.n267 B.n266 585
R221 B.n265 B.n264 585
R222 B.n263 B.n262 585
R223 B.n261 B.n260 585
R224 B.n259 B.n258 585
R225 B.n257 B.n256 585
R226 B.n255 B.n254 585
R227 B.n253 B.n252 585
R228 B.n251 B.n250 585
R229 B.n249 B.n248 585
R230 B.n247 B.n246 585
R231 B.n245 B.n244 585
R232 B.n243 B.n242 585
R233 B.n241 B.n240 585
R234 B.n239 B.n238 585
R235 B.n237 B.n236 585
R236 B.n235 B.n234 585
R237 B.n233 B.n232 585
R238 B.n231 B.n230 585
R239 B.n229 B.n228 585
R240 B.n227 B.n226 585
R241 B.n225 B.n224 585
R242 B.n223 B.n222 585
R243 B.n221 B.n220 585
R244 B.n219 B.n218 585
R245 B.n217 B.n216 585
R246 B.n215 B.n214 585
R247 B.n213 B.n212 585
R248 B.n211 B.n210 585
R249 B.n209 B.n208 585
R250 B.n207 B.n206 585
R251 B.n205 B.n204 585
R252 B.n203 B.n202 585
R253 B.n201 B.n200 585
R254 B.n199 B.n198 585
R255 B.n197 B.n196 585
R256 B.n195 B.n194 585
R257 B.n193 B.n192 585
R258 B.n191 B.n190 585
R259 B.n189 B.n188 585
R260 B.n187 B.n186 585
R261 B.n185 B.n184 585
R262 B.n183 B.n182 585
R263 B.n181 B.n180 585
R264 B.n179 B.n178 585
R265 B.n177 B.n176 585
R266 B.n175 B.n174 585
R267 B.n173 B.n172 585
R268 B.n171 B.n170 585
R269 B.n169 B.n168 585
R270 B.n131 B.n130 585
R271 B.n879 B.n132 585
R272 B.n884 B.n132 585
R273 B.n878 B.n877 585
R274 B.n877 B.n128 585
R275 B.n876 B.n127 585
R276 B.n890 B.n127 585
R277 B.n875 B.n126 585
R278 B.n891 B.n126 585
R279 B.n874 B.n125 585
R280 B.n892 B.n125 585
R281 B.n873 B.n872 585
R282 B.n872 B.n121 585
R283 B.n871 B.n120 585
R284 B.n898 B.n120 585
R285 B.n870 B.n119 585
R286 B.n899 B.n119 585
R287 B.n869 B.n118 585
R288 B.n900 B.n118 585
R289 B.n868 B.n867 585
R290 B.n867 B.n114 585
R291 B.n866 B.n113 585
R292 B.n906 B.n113 585
R293 B.n865 B.n112 585
R294 B.n907 B.n112 585
R295 B.n864 B.n111 585
R296 B.n908 B.n111 585
R297 B.n863 B.n862 585
R298 B.n862 B.n107 585
R299 B.n861 B.n106 585
R300 B.n914 B.n106 585
R301 B.n860 B.n105 585
R302 B.n915 B.n105 585
R303 B.n859 B.n104 585
R304 B.n916 B.n104 585
R305 B.n858 B.n857 585
R306 B.n857 B.n100 585
R307 B.n856 B.n99 585
R308 B.n922 B.n99 585
R309 B.n855 B.n98 585
R310 B.n923 B.n98 585
R311 B.n854 B.n97 585
R312 B.n924 B.n97 585
R313 B.n853 B.n852 585
R314 B.n852 B.n93 585
R315 B.n851 B.n92 585
R316 B.n930 B.n92 585
R317 B.n850 B.n91 585
R318 B.n931 B.n91 585
R319 B.n849 B.n90 585
R320 B.n932 B.n90 585
R321 B.n848 B.n847 585
R322 B.n847 B.n86 585
R323 B.n846 B.n85 585
R324 B.n938 B.n85 585
R325 B.n845 B.n84 585
R326 B.n939 B.n84 585
R327 B.n844 B.n83 585
R328 B.n940 B.n83 585
R329 B.n843 B.n842 585
R330 B.n842 B.n79 585
R331 B.n841 B.n78 585
R332 B.n946 B.n78 585
R333 B.n840 B.n77 585
R334 B.n947 B.n77 585
R335 B.n839 B.n76 585
R336 B.n948 B.n76 585
R337 B.n838 B.n837 585
R338 B.n837 B.n75 585
R339 B.n836 B.n71 585
R340 B.n954 B.n71 585
R341 B.n835 B.n70 585
R342 B.n955 B.n70 585
R343 B.n834 B.n69 585
R344 B.n956 B.n69 585
R345 B.n833 B.n832 585
R346 B.n832 B.n65 585
R347 B.n831 B.n64 585
R348 B.n962 B.n64 585
R349 B.n830 B.n63 585
R350 B.n963 B.n63 585
R351 B.n829 B.n62 585
R352 B.n964 B.n62 585
R353 B.n828 B.n827 585
R354 B.n827 B.n58 585
R355 B.n826 B.n57 585
R356 B.n970 B.n57 585
R357 B.n825 B.n56 585
R358 B.n971 B.n56 585
R359 B.n824 B.n55 585
R360 B.n972 B.n55 585
R361 B.n823 B.n822 585
R362 B.n822 B.n51 585
R363 B.n821 B.n50 585
R364 B.n978 B.n50 585
R365 B.n820 B.n49 585
R366 B.n979 B.n49 585
R367 B.n819 B.n48 585
R368 B.n980 B.n48 585
R369 B.n818 B.n817 585
R370 B.n817 B.n44 585
R371 B.n816 B.n43 585
R372 B.n986 B.n43 585
R373 B.n815 B.n42 585
R374 B.n987 B.n42 585
R375 B.n814 B.n41 585
R376 B.n988 B.n41 585
R377 B.n813 B.n812 585
R378 B.n812 B.n37 585
R379 B.n811 B.n36 585
R380 B.n994 B.n36 585
R381 B.n810 B.n35 585
R382 B.n995 B.n35 585
R383 B.n809 B.n34 585
R384 B.n996 B.n34 585
R385 B.n808 B.n807 585
R386 B.n807 B.n30 585
R387 B.n806 B.n29 585
R388 B.n1002 B.n29 585
R389 B.n805 B.n28 585
R390 B.n1003 B.n28 585
R391 B.n804 B.n27 585
R392 B.n1004 B.n27 585
R393 B.n803 B.n802 585
R394 B.n802 B.n23 585
R395 B.n801 B.n22 585
R396 B.n1010 B.n22 585
R397 B.n800 B.n21 585
R398 B.n1011 B.n21 585
R399 B.n799 B.n20 585
R400 B.n1012 B.n20 585
R401 B.n798 B.n797 585
R402 B.n797 B.n19 585
R403 B.n796 B.n15 585
R404 B.n1018 B.n15 585
R405 B.n795 B.n14 585
R406 B.n1019 B.n14 585
R407 B.n794 B.n13 585
R408 B.n1020 B.n13 585
R409 B.n793 B.n792 585
R410 B.n792 B.n12 585
R411 B.n791 B.n790 585
R412 B.n791 B.n8 585
R413 B.n789 B.n7 585
R414 B.n1027 B.n7 585
R415 B.n788 B.n6 585
R416 B.n1028 B.n6 585
R417 B.n787 B.n5 585
R418 B.n1029 B.n5 585
R419 B.n786 B.n785 585
R420 B.n785 B.n4 585
R421 B.n784 B.n279 585
R422 B.n784 B.n783 585
R423 B.n774 B.n280 585
R424 B.n281 B.n280 585
R425 B.n776 B.n775 585
R426 B.n777 B.n776 585
R427 B.n773 B.n286 585
R428 B.n286 B.n285 585
R429 B.n772 B.n771 585
R430 B.n771 B.n770 585
R431 B.n288 B.n287 585
R432 B.n763 B.n288 585
R433 B.n762 B.n761 585
R434 B.n764 B.n762 585
R435 B.n760 B.n293 585
R436 B.n293 B.n292 585
R437 B.n759 B.n758 585
R438 B.n758 B.n757 585
R439 B.n295 B.n294 585
R440 B.n296 B.n295 585
R441 B.n750 B.n749 585
R442 B.n751 B.n750 585
R443 B.n748 B.n301 585
R444 B.n301 B.n300 585
R445 B.n747 B.n746 585
R446 B.n746 B.n745 585
R447 B.n303 B.n302 585
R448 B.n304 B.n303 585
R449 B.n738 B.n737 585
R450 B.n739 B.n738 585
R451 B.n736 B.n309 585
R452 B.n309 B.n308 585
R453 B.n735 B.n734 585
R454 B.n734 B.n733 585
R455 B.n311 B.n310 585
R456 B.n312 B.n311 585
R457 B.n726 B.n725 585
R458 B.n727 B.n726 585
R459 B.n724 B.n317 585
R460 B.n317 B.n316 585
R461 B.n723 B.n722 585
R462 B.n722 B.n721 585
R463 B.n319 B.n318 585
R464 B.n320 B.n319 585
R465 B.n714 B.n713 585
R466 B.n715 B.n714 585
R467 B.n712 B.n325 585
R468 B.n325 B.n324 585
R469 B.n711 B.n710 585
R470 B.n710 B.n709 585
R471 B.n327 B.n326 585
R472 B.n328 B.n327 585
R473 B.n702 B.n701 585
R474 B.n703 B.n702 585
R475 B.n700 B.n333 585
R476 B.n333 B.n332 585
R477 B.n699 B.n698 585
R478 B.n698 B.n697 585
R479 B.n335 B.n334 585
R480 B.n336 B.n335 585
R481 B.n690 B.n689 585
R482 B.n691 B.n690 585
R483 B.n688 B.n341 585
R484 B.n341 B.n340 585
R485 B.n687 B.n686 585
R486 B.n686 B.n685 585
R487 B.n343 B.n342 585
R488 B.n344 B.n343 585
R489 B.n678 B.n677 585
R490 B.n679 B.n678 585
R491 B.n676 B.n349 585
R492 B.n349 B.n348 585
R493 B.n675 B.n674 585
R494 B.n674 B.n673 585
R495 B.n351 B.n350 585
R496 B.n666 B.n351 585
R497 B.n665 B.n664 585
R498 B.n667 B.n665 585
R499 B.n663 B.n356 585
R500 B.n356 B.n355 585
R501 B.n662 B.n661 585
R502 B.n661 B.n660 585
R503 B.n358 B.n357 585
R504 B.n359 B.n358 585
R505 B.n653 B.n652 585
R506 B.n654 B.n653 585
R507 B.n651 B.n364 585
R508 B.n364 B.n363 585
R509 B.n650 B.n649 585
R510 B.n649 B.n648 585
R511 B.n366 B.n365 585
R512 B.n367 B.n366 585
R513 B.n641 B.n640 585
R514 B.n642 B.n641 585
R515 B.n639 B.n372 585
R516 B.n372 B.n371 585
R517 B.n638 B.n637 585
R518 B.n637 B.n636 585
R519 B.n374 B.n373 585
R520 B.n375 B.n374 585
R521 B.n629 B.n628 585
R522 B.n630 B.n629 585
R523 B.n627 B.n380 585
R524 B.n380 B.n379 585
R525 B.n626 B.n625 585
R526 B.n625 B.n624 585
R527 B.n382 B.n381 585
R528 B.n383 B.n382 585
R529 B.n617 B.n616 585
R530 B.n618 B.n617 585
R531 B.n615 B.n388 585
R532 B.n388 B.n387 585
R533 B.n614 B.n613 585
R534 B.n613 B.n612 585
R535 B.n390 B.n389 585
R536 B.n391 B.n390 585
R537 B.n605 B.n604 585
R538 B.n606 B.n605 585
R539 B.n603 B.n396 585
R540 B.n396 B.n395 585
R541 B.n602 B.n601 585
R542 B.n601 B.n600 585
R543 B.n398 B.n397 585
R544 B.n399 B.n398 585
R545 B.n593 B.n592 585
R546 B.n594 B.n593 585
R547 B.n591 B.n404 585
R548 B.n404 B.n403 585
R549 B.n590 B.n589 585
R550 B.n589 B.n588 585
R551 B.n406 B.n405 585
R552 B.n407 B.n406 585
R553 B.n581 B.n580 585
R554 B.n582 B.n581 585
R555 B.n579 B.n412 585
R556 B.n412 B.n411 585
R557 B.n578 B.n577 585
R558 B.n577 B.n576 585
R559 B.n414 B.n413 585
R560 B.n415 B.n414 585
R561 B.n569 B.n568 585
R562 B.n570 B.n569 585
R563 B.n418 B.n417 585
R564 B.n453 B.n451 585
R565 B.n454 B.n450 585
R566 B.n454 B.n419 585
R567 B.n457 B.n456 585
R568 B.n458 B.n449 585
R569 B.n460 B.n459 585
R570 B.n462 B.n448 585
R571 B.n465 B.n464 585
R572 B.n466 B.n447 585
R573 B.n468 B.n467 585
R574 B.n470 B.n446 585
R575 B.n473 B.n472 585
R576 B.n474 B.n445 585
R577 B.n476 B.n475 585
R578 B.n478 B.n444 585
R579 B.n481 B.n480 585
R580 B.n482 B.n443 585
R581 B.n484 B.n483 585
R582 B.n486 B.n442 585
R583 B.n489 B.n488 585
R584 B.n490 B.n441 585
R585 B.n492 B.n491 585
R586 B.n494 B.n440 585
R587 B.n497 B.n496 585
R588 B.n499 B.n437 585
R589 B.n501 B.n500 585
R590 B.n503 B.n436 585
R591 B.n506 B.n505 585
R592 B.n507 B.n435 585
R593 B.n509 B.n508 585
R594 B.n511 B.n434 585
R595 B.n514 B.n513 585
R596 B.n515 B.n433 585
R597 B.n520 B.n519 585
R598 B.n522 B.n432 585
R599 B.n525 B.n524 585
R600 B.n526 B.n431 585
R601 B.n528 B.n527 585
R602 B.n530 B.n430 585
R603 B.n533 B.n532 585
R604 B.n534 B.n429 585
R605 B.n536 B.n535 585
R606 B.n538 B.n428 585
R607 B.n541 B.n540 585
R608 B.n542 B.n427 585
R609 B.n544 B.n543 585
R610 B.n546 B.n426 585
R611 B.n549 B.n548 585
R612 B.n550 B.n425 585
R613 B.n552 B.n551 585
R614 B.n554 B.n424 585
R615 B.n557 B.n556 585
R616 B.n558 B.n423 585
R617 B.n560 B.n559 585
R618 B.n562 B.n422 585
R619 B.n563 B.n421 585
R620 B.n566 B.n565 585
R621 B.n567 B.n420 585
R622 B.n420 B.n419 585
R623 B.n572 B.n571 585
R624 B.n571 B.n570 585
R625 B.n573 B.n416 585
R626 B.n416 B.n415 585
R627 B.n575 B.n574 585
R628 B.n576 B.n575 585
R629 B.n410 B.n409 585
R630 B.n411 B.n410 585
R631 B.n584 B.n583 585
R632 B.n583 B.n582 585
R633 B.n585 B.n408 585
R634 B.n408 B.n407 585
R635 B.n587 B.n586 585
R636 B.n588 B.n587 585
R637 B.n402 B.n401 585
R638 B.n403 B.n402 585
R639 B.n596 B.n595 585
R640 B.n595 B.n594 585
R641 B.n597 B.n400 585
R642 B.n400 B.n399 585
R643 B.n599 B.n598 585
R644 B.n600 B.n599 585
R645 B.n394 B.n393 585
R646 B.n395 B.n394 585
R647 B.n608 B.n607 585
R648 B.n607 B.n606 585
R649 B.n609 B.n392 585
R650 B.n392 B.n391 585
R651 B.n611 B.n610 585
R652 B.n612 B.n611 585
R653 B.n386 B.n385 585
R654 B.n387 B.n386 585
R655 B.n620 B.n619 585
R656 B.n619 B.n618 585
R657 B.n621 B.n384 585
R658 B.n384 B.n383 585
R659 B.n623 B.n622 585
R660 B.n624 B.n623 585
R661 B.n378 B.n377 585
R662 B.n379 B.n378 585
R663 B.n632 B.n631 585
R664 B.n631 B.n630 585
R665 B.n633 B.n376 585
R666 B.n376 B.n375 585
R667 B.n635 B.n634 585
R668 B.n636 B.n635 585
R669 B.n370 B.n369 585
R670 B.n371 B.n370 585
R671 B.n644 B.n643 585
R672 B.n643 B.n642 585
R673 B.n645 B.n368 585
R674 B.n368 B.n367 585
R675 B.n647 B.n646 585
R676 B.n648 B.n647 585
R677 B.n362 B.n361 585
R678 B.n363 B.n362 585
R679 B.n656 B.n655 585
R680 B.n655 B.n654 585
R681 B.n657 B.n360 585
R682 B.n360 B.n359 585
R683 B.n659 B.n658 585
R684 B.n660 B.n659 585
R685 B.n354 B.n353 585
R686 B.n355 B.n354 585
R687 B.n669 B.n668 585
R688 B.n668 B.n667 585
R689 B.n670 B.n352 585
R690 B.n666 B.n352 585
R691 B.n672 B.n671 585
R692 B.n673 B.n672 585
R693 B.n347 B.n346 585
R694 B.n348 B.n347 585
R695 B.n681 B.n680 585
R696 B.n680 B.n679 585
R697 B.n682 B.n345 585
R698 B.n345 B.n344 585
R699 B.n684 B.n683 585
R700 B.n685 B.n684 585
R701 B.n339 B.n338 585
R702 B.n340 B.n339 585
R703 B.n693 B.n692 585
R704 B.n692 B.n691 585
R705 B.n694 B.n337 585
R706 B.n337 B.n336 585
R707 B.n696 B.n695 585
R708 B.n697 B.n696 585
R709 B.n331 B.n330 585
R710 B.n332 B.n331 585
R711 B.n705 B.n704 585
R712 B.n704 B.n703 585
R713 B.n706 B.n329 585
R714 B.n329 B.n328 585
R715 B.n708 B.n707 585
R716 B.n709 B.n708 585
R717 B.n323 B.n322 585
R718 B.n324 B.n323 585
R719 B.n717 B.n716 585
R720 B.n716 B.n715 585
R721 B.n718 B.n321 585
R722 B.n321 B.n320 585
R723 B.n720 B.n719 585
R724 B.n721 B.n720 585
R725 B.n315 B.n314 585
R726 B.n316 B.n315 585
R727 B.n729 B.n728 585
R728 B.n728 B.n727 585
R729 B.n730 B.n313 585
R730 B.n313 B.n312 585
R731 B.n732 B.n731 585
R732 B.n733 B.n732 585
R733 B.n307 B.n306 585
R734 B.n308 B.n307 585
R735 B.n741 B.n740 585
R736 B.n740 B.n739 585
R737 B.n742 B.n305 585
R738 B.n305 B.n304 585
R739 B.n744 B.n743 585
R740 B.n745 B.n744 585
R741 B.n299 B.n298 585
R742 B.n300 B.n299 585
R743 B.n753 B.n752 585
R744 B.n752 B.n751 585
R745 B.n754 B.n297 585
R746 B.n297 B.n296 585
R747 B.n756 B.n755 585
R748 B.n757 B.n756 585
R749 B.n291 B.n290 585
R750 B.n292 B.n291 585
R751 B.n766 B.n765 585
R752 B.n765 B.n764 585
R753 B.n767 B.n289 585
R754 B.n763 B.n289 585
R755 B.n769 B.n768 585
R756 B.n770 B.n769 585
R757 B.n284 B.n283 585
R758 B.n285 B.n284 585
R759 B.n779 B.n778 585
R760 B.n778 B.n777 585
R761 B.n780 B.n282 585
R762 B.n282 B.n281 585
R763 B.n782 B.n781 585
R764 B.n783 B.n782 585
R765 B.n3 B.n0 585
R766 B.n4 B.n3 585
R767 B.n1026 B.n1 585
R768 B.n1027 B.n1026 585
R769 B.n1025 B.n1024 585
R770 B.n1025 B.n8 585
R771 B.n1023 B.n9 585
R772 B.n12 B.n9 585
R773 B.n1022 B.n1021 585
R774 B.n1021 B.n1020 585
R775 B.n11 B.n10 585
R776 B.n1019 B.n11 585
R777 B.n1017 B.n1016 585
R778 B.n1018 B.n1017 585
R779 B.n1015 B.n16 585
R780 B.n19 B.n16 585
R781 B.n1014 B.n1013 585
R782 B.n1013 B.n1012 585
R783 B.n18 B.n17 585
R784 B.n1011 B.n18 585
R785 B.n1009 B.n1008 585
R786 B.n1010 B.n1009 585
R787 B.n1007 B.n24 585
R788 B.n24 B.n23 585
R789 B.n1006 B.n1005 585
R790 B.n1005 B.n1004 585
R791 B.n26 B.n25 585
R792 B.n1003 B.n26 585
R793 B.n1001 B.n1000 585
R794 B.n1002 B.n1001 585
R795 B.n999 B.n31 585
R796 B.n31 B.n30 585
R797 B.n998 B.n997 585
R798 B.n997 B.n996 585
R799 B.n33 B.n32 585
R800 B.n995 B.n33 585
R801 B.n993 B.n992 585
R802 B.n994 B.n993 585
R803 B.n991 B.n38 585
R804 B.n38 B.n37 585
R805 B.n990 B.n989 585
R806 B.n989 B.n988 585
R807 B.n40 B.n39 585
R808 B.n987 B.n40 585
R809 B.n985 B.n984 585
R810 B.n986 B.n985 585
R811 B.n983 B.n45 585
R812 B.n45 B.n44 585
R813 B.n982 B.n981 585
R814 B.n981 B.n980 585
R815 B.n47 B.n46 585
R816 B.n979 B.n47 585
R817 B.n977 B.n976 585
R818 B.n978 B.n977 585
R819 B.n975 B.n52 585
R820 B.n52 B.n51 585
R821 B.n974 B.n973 585
R822 B.n973 B.n972 585
R823 B.n54 B.n53 585
R824 B.n971 B.n54 585
R825 B.n969 B.n968 585
R826 B.n970 B.n969 585
R827 B.n967 B.n59 585
R828 B.n59 B.n58 585
R829 B.n966 B.n965 585
R830 B.n965 B.n964 585
R831 B.n61 B.n60 585
R832 B.n963 B.n61 585
R833 B.n961 B.n960 585
R834 B.n962 B.n961 585
R835 B.n959 B.n66 585
R836 B.n66 B.n65 585
R837 B.n958 B.n957 585
R838 B.n957 B.n956 585
R839 B.n68 B.n67 585
R840 B.n955 B.n68 585
R841 B.n953 B.n952 585
R842 B.n954 B.n953 585
R843 B.n951 B.n72 585
R844 B.n75 B.n72 585
R845 B.n950 B.n949 585
R846 B.n949 B.n948 585
R847 B.n74 B.n73 585
R848 B.n947 B.n74 585
R849 B.n945 B.n944 585
R850 B.n946 B.n945 585
R851 B.n943 B.n80 585
R852 B.n80 B.n79 585
R853 B.n942 B.n941 585
R854 B.n941 B.n940 585
R855 B.n82 B.n81 585
R856 B.n939 B.n82 585
R857 B.n937 B.n936 585
R858 B.n938 B.n937 585
R859 B.n935 B.n87 585
R860 B.n87 B.n86 585
R861 B.n934 B.n933 585
R862 B.n933 B.n932 585
R863 B.n89 B.n88 585
R864 B.n931 B.n89 585
R865 B.n929 B.n928 585
R866 B.n930 B.n929 585
R867 B.n927 B.n94 585
R868 B.n94 B.n93 585
R869 B.n926 B.n925 585
R870 B.n925 B.n924 585
R871 B.n96 B.n95 585
R872 B.n923 B.n96 585
R873 B.n921 B.n920 585
R874 B.n922 B.n921 585
R875 B.n919 B.n101 585
R876 B.n101 B.n100 585
R877 B.n918 B.n917 585
R878 B.n917 B.n916 585
R879 B.n103 B.n102 585
R880 B.n915 B.n103 585
R881 B.n913 B.n912 585
R882 B.n914 B.n913 585
R883 B.n911 B.n108 585
R884 B.n108 B.n107 585
R885 B.n910 B.n909 585
R886 B.n909 B.n908 585
R887 B.n110 B.n109 585
R888 B.n907 B.n110 585
R889 B.n905 B.n904 585
R890 B.n906 B.n905 585
R891 B.n903 B.n115 585
R892 B.n115 B.n114 585
R893 B.n902 B.n901 585
R894 B.n901 B.n900 585
R895 B.n117 B.n116 585
R896 B.n899 B.n117 585
R897 B.n897 B.n896 585
R898 B.n898 B.n897 585
R899 B.n895 B.n122 585
R900 B.n122 B.n121 585
R901 B.n894 B.n893 585
R902 B.n893 B.n892 585
R903 B.n124 B.n123 585
R904 B.n891 B.n124 585
R905 B.n889 B.n888 585
R906 B.n890 B.n889 585
R907 B.n887 B.n129 585
R908 B.n129 B.n128 585
R909 B.n886 B.n885 585
R910 B.n885 B.n884 585
R911 B.n1030 B.n1029 585
R912 B.n1028 B.n2 585
R913 B.n885 B.n131 530.939
R914 B.n881 B.n132 530.939
R915 B.n569 B.n420 530.939
R916 B.n571 B.n418 530.939
R917 B.n883 B.n882 256.663
R918 B.n883 B.n160 256.663
R919 B.n883 B.n159 256.663
R920 B.n883 B.n158 256.663
R921 B.n883 B.n157 256.663
R922 B.n883 B.n156 256.663
R923 B.n883 B.n155 256.663
R924 B.n883 B.n154 256.663
R925 B.n883 B.n153 256.663
R926 B.n883 B.n152 256.663
R927 B.n883 B.n151 256.663
R928 B.n883 B.n150 256.663
R929 B.n883 B.n149 256.663
R930 B.n883 B.n148 256.663
R931 B.n883 B.n147 256.663
R932 B.n883 B.n146 256.663
R933 B.n883 B.n145 256.663
R934 B.n883 B.n144 256.663
R935 B.n883 B.n143 256.663
R936 B.n883 B.n142 256.663
R937 B.n883 B.n141 256.663
R938 B.n883 B.n140 256.663
R939 B.n883 B.n139 256.663
R940 B.n883 B.n138 256.663
R941 B.n883 B.n137 256.663
R942 B.n883 B.n136 256.663
R943 B.n883 B.n135 256.663
R944 B.n883 B.n134 256.663
R945 B.n883 B.n133 256.663
R946 B.n452 B.n419 256.663
R947 B.n455 B.n419 256.663
R948 B.n461 B.n419 256.663
R949 B.n463 B.n419 256.663
R950 B.n469 B.n419 256.663
R951 B.n471 B.n419 256.663
R952 B.n477 B.n419 256.663
R953 B.n479 B.n419 256.663
R954 B.n485 B.n419 256.663
R955 B.n487 B.n419 256.663
R956 B.n493 B.n419 256.663
R957 B.n495 B.n419 256.663
R958 B.n502 B.n419 256.663
R959 B.n504 B.n419 256.663
R960 B.n510 B.n419 256.663
R961 B.n512 B.n419 256.663
R962 B.n521 B.n419 256.663
R963 B.n523 B.n419 256.663
R964 B.n529 B.n419 256.663
R965 B.n531 B.n419 256.663
R966 B.n537 B.n419 256.663
R967 B.n539 B.n419 256.663
R968 B.n545 B.n419 256.663
R969 B.n547 B.n419 256.663
R970 B.n553 B.n419 256.663
R971 B.n555 B.n419 256.663
R972 B.n561 B.n419 256.663
R973 B.n564 B.n419 256.663
R974 B.n1032 B.n1031 256.663
R975 B.n165 B.t14 253.495
R976 B.n162 B.t21 253.495
R977 B.n516 B.t10 253.495
R978 B.n438 B.t18 253.495
R979 B.n170 B.n169 163.367
R980 B.n174 B.n173 163.367
R981 B.n178 B.n177 163.367
R982 B.n182 B.n181 163.367
R983 B.n186 B.n185 163.367
R984 B.n190 B.n189 163.367
R985 B.n194 B.n193 163.367
R986 B.n198 B.n197 163.367
R987 B.n202 B.n201 163.367
R988 B.n206 B.n205 163.367
R989 B.n210 B.n209 163.367
R990 B.n214 B.n213 163.367
R991 B.n218 B.n217 163.367
R992 B.n222 B.n221 163.367
R993 B.n226 B.n225 163.367
R994 B.n230 B.n229 163.367
R995 B.n234 B.n233 163.367
R996 B.n238 B.n237 163.367
R997 B.n242 B.n241 163.367
R998 B.n246 B.n245 163.367
R999 B.n250 B.n249 163.367
R1000 B.n254 B.n253 163.367
R1001 B.n258 B.n257 163.367
R1002 B.n262 B.n261 163.367
R1003 B.n266 B.n265 163.367
R1004 B.n270 B.n269 163.367
R1005 B.n274 B.n273 163.367
R1006 B.n276 B.n161 163.367
R1007 B.n569 B.n414 163.367
R1008 B.n577 B.n414 163.367
R1009 B.n577 B.n412 163.367
R1010 B.n581 B.n412 163.367
R1011 B.n581 B.n406 163.367
R1012 B.n589 B.n406 163.367
R1013 B.n589 B.n404 163.367
R1014 B.n593 B.n404 163.367
R1015 B.n593 B.n398 163.367
R1016 B.n601 B.n398 163.367
R1017 B.n601 B.n396 163.367
R1018 B.n605 B.n396 163.367
R1019 B.n605 B.n390 163.367
R1020 B.n613 B.n390 163.367
R1021 B.n613 B.n388 163.367
R1022 B.n617 B.n388 163.367
R1023 B.n617 B.n382 163.367
R1024 B.n625 B.n382 163.367
R1025 B.n625 B.n380 163.367
R1026 B.n629 B.n380 163.367
R1027 B.n629 B.n374 163.367
R1028 B.n637 B.n374 163.367
R1029 B.n637 B.n372 163.367
R1030 B.n641 B.n372 163.367
R1031 B.n641 B.n366 163.367
R1032 B.n649 B.n366 163.367
R1033 B.n649 B.n364 163.367
R1034 B.n653 B.n364 163.367
R1035 B.n653 B.n358 163.367
R1036 B.n661 B.n358 163.367
R1037 B.n661 B.n356 163.367
R1038 B.n665 B.n356 163.367
R1039 B.n665 B.n351 163.367
R1040 B.n674 B.n351 163.367
R1041 B.n674 B.n349 163.367
R1042 B.n678 B.n349 163.367
R1043 B.n678 B.n343 163.367
R1044 B.n686 B.n343 163.367
R1045 B.n686 B.n341 163.367
R1046 B.n690 B.n341 163.367
R1047 B.n690 B.n335 163.367
R1048 B.n698 B.n335 163.367
R1049 B.n698 B.n333 163.367
R1050 B.n702 B.n333 163.367
R1051 B.n702 B.n327 163.367
R1052 B.n710 B.n327 163.367
R1053 B.n710 B.n325 163.367
R1054 B.n714 B.n325 163.367
R1055 B.n714 B.n319 163.367
R1056 B.n722 B.n319 163.367
R1057 B.n722 B.n317 163.367
R1058 B.n726 B.n317 163.367
R1059 B.n726 B.n311 163.367
R1060 B.n734 B.n311 163.367
R1061 B.n734 B.n309 163.367
R1062 B.n738 B.n309 163.367
R1063 B.n738 B.n303 163.367
R1064 B.n746 B.n303 163.367
R1065 B.n746 B.n301 163.367
R1066 B.n750 B.n301 163.367
R1067 B.n750 B.n295 163.367
R1068 B.n758 B.n295 163.367
R1069 B.n758 B.n293 163.367
R1070 B.n762 B.n293 163.367
R1071 B.n762 B.n288 163.367
R1072 B.n771 B.n288 163.367
R1073 B.n771 B.n286 163.367
R1074 B.n776 B.n286 163.367
R1075 B.n776 B.n280 163.367
R1076 B.n784 B.n280 163.367
R1077 B.n785 B.n784 163.367
R1078 B.n785 B.n5 163.367
R1079 B.n6 B.n5 163.367
R1080 B.n7 B.n6 163.367
R1081 B.n791 B.n7 163.367
R1082 B.n792 B.n791 163.367
R1083 B.n792 B.n13 163.367
R1084 B.n14 B.n13 163.367
R1085 B.n15 B.n14 163.367
R1086 B.n797 B.n15 163.367
R1087 B.n797 B.n20 163.367
R1088 B.n21 B.n20 163.367
R1089 B.n22 B.n21 163.367
R1090 B.n802 B.n22 163.367
R1091 B.n802 B.n27 163.367
R1092 B.n28 B.n27 163.367
R1093 B.n29 B.n28 163.367
R1094 B.n807 B.n29 163.367
R1095 B.n807 B.n34 163.367
R1096 B.n35 B.n34 163.367
R1097 B.n36 B.n35 163.367
R1098 B.n812 B.n36 163.367
R1099 B.n812 B.n41 163.367
R1100 B.n42 B.n41 163.367
R1101 B.n43 B.n42 163.367
R1102 B.n817 B.n43 163.367
R1103 B.n817 B.n48 163.367
R1104 B.n49 B.n48 163.367
R1105 B.n50 B.n49 163.367
R1106 B.n822 B.n50 163.367
R1107 B.n822 B.n55 163.367
R1108 B.n56 B.n55 163.367
R1109 B.n57 B.n56 163.367
R1110 B.n827 B.n57 163.367
R1111 B.n827 B.n62 163.367
R1112 B.n63 B.n62 163.367
R1113 B.n64 B.n63 163.367
R1114 B.n832 B.n64 163.367
R1115 B.n832 B.n69 163.367
R1116 B.n70 B.n69 163.367
R1117 B.n71 B.n70 163.367
R1118 B.n837 B.n71 163.367
R1119 B.n837 B.n76 163.367
R1120 B.n77 B.n76 163.367
R1121 B.n78 B.n77 163.367
R1122 B.n842 B.n78 163.367
R1123 B.n842 B.n83 163.367
R1124 B.n84 B.n83 163.367
R1125 B.n85 B.n84 163.367
R1126 B.n847 B.n85 163.367
R1127 B.n847 B.n90 163.367
R1128 B.n91 B.n90 163.367
R1129 B.n92 B.n91 163.367
R1130 B.n852 B.n92 163.367
R1131 B.n852 B.n97 163.367
R1132 B.n98 B.n97 163.367
R1133 B.n99 B.n98 163.367
R1134 B.n857 B.n99 163.367
R1135 B.n857 B.n104 163.367
R1136 B.n105 B.n104 163.367
R1137 B.n106 B.n105 163.367
R1138 B.n862 B.n106 163.367
R1139 B.n862 B.n111 163.367
R1140 B.n112 B.n111 163.367
R1141 B.n113 B.n112 163.367
R1142 B.n867 B.n113 163.367
R1143 B.n867 B.n118 163.367
R1144 B.n119 B.n118 163.367
R1145 B.n120 B.n119 163.367
R1146 B.n872 B.n120 163.367
R1147 B.n872 B.n125 163.367
R1148 B.n126 B.n125 163.367
R1149 B.n127 B.n126 163.367
R1150 B.n877 B.n127 163.367
R1151 B.n877 B.n132 163.367
R1152 B.n454 B.n453 163.367
R1153 B.n456 B.n454 163.367
R1154 B.n460 B.n449 163.367
R1155 B.n464 B.n462 163.367
R1156 B.n468 B.n447 163.367
R1157 B.n472 B.n470 163.367
R1158 B.n476 B.n445 163.367
R1159 B.n480 B.n478 163.367
R1160 B.n484 B.n443 163.367
R1161 B.n488 B.n486 163.367
R1162 B.n492 B.n441 163.367
R1163 B.n496 B.n494 163.367
R1164 B.n501 B.n437 163.367
R1165 B.n505 B.n503 163.367
R1166 B.n509 B.n435 163.367
R1167 B.n513 B.n511 163.367
R1168 B.n520 B.n433 163.367
R1169 B.n524 B.n522 163.367
R1170 B.n528 B.n431 163.367
R1171 B.n532 B.n530 163.367
R1172 B.n536 B.n429 163.367
R1173 B.n540 B.n538 163.367
R1174 B.n544 B.n427 163.367
R1175 B.n548 B.n546 163.367
R1176 B.n552 B.n425 163.367
R1177 B.n556 B.n554 163.367
R1178 B.n560 B.n423 163.367
R1179 B.n563 B.n562 163.367
R1180 B.n565 B.n420 163.367
R1181 B.n571 B.n416 163.367
R1182 B.n575 B.n416 163.367
R1183 B.n575 B.n410 163.367
R1184 B.n583 B.n410 163.367
R1185 B.n583 B.n408 163.367
R1186 B.n587 B.n408 163.367
R1187 B.n587 B.n402 163.367
R1188 B.n595 B.n402 163.367
R1189 B.n595 B.n400 163.367
R1190 B.n599 B.n400 163.367
R1191 B.n599 B.n394 163.367
R1192 B.n607 B.n394 163.367
R1193 B.n607 B.n392 163.367
R1194 B.n611 B.n392 163.367
R1195 B.n611 B.n386 163.367
R1196 B.n619 B.n386 163.367
R1197 B.n619 B.n384 163.367
R1198 B.n623 B.n384 163.367
R1199 B.n623 B.n378 163.367
R1200 B.n631 B.n378 163.367
R1201 B.n631 B.n376 163.367
R1202 B.n635 B.n376 163.367
R1203 B.n635 B.n370 163.367
R1204 B.n643 B.n370 163.367
R1205 B.n643 B.n368 163.367
R1206 B.n647 B.n368 163.367
R1207 B.n647 B.n362 163.367
R1208 B.n655 B.n362 163.367
R1209 B.n655 B.n360 163.367
R1210 B.n659 B.n360 163.367
R1211 B.n659 B.n354 163.367
R1212 B.n668 B.n354 163.367
R1213 B.n668 B.n352 163.367
R1214 B.n672 B.n352 163.367
R1215 B.n672 B.n347 163.367
R1216 B.n680 B.n347 163.367
R1217 B.n680 B.n345 163.367
R1218 B.n684 B.n345 163.367
R1219 B.n684 B.n339 163.367
R1220 B.n692 B.n339 163.367
R1221 B.n692 B.n337 163.367
R1222 B.n696 B.n337 163.367
R1223 B.n696 B.n331 163.367
R1224 B.n704 B.n331 163.367
R1225 B.n704 B.n329 163.367
R1226 B.n708 B.n329 163.367
R1227 B.n708 B.n323 163.367
R1228 B.n716 B.n323 163.367
R1229 B.n716 B.n321 163.367
R1230 B.n720 B.n321 163.367
R1231 B.n720 B.n315 163.367
R1232 B.n728 B.n315 163.367
R1233 B.n728 B.n313 163.367
R1234 B.n732 B.n313 163.367
R1235 B.n732 B.n307 163.367
R1236 B.n740 B.n307 163.367
R1237 B.n740 B.n305 163.367
R1238 B.n744 B.n305 163.367
R1239 B.n744 B.n299 163.367
R1240 B.n752 B.n299 163.367
R1241 B.n752 B.n297 163.367
R1242 B.n756 B.n297 163.367
R1243 B.n756 B.n291 163.367
R1244 B.n765 B.n291 163.367
R1245 B.n765 B.n289 163.367
R1246 B.n769 B.n289 163.367
R1247 B.n769 B.n284 163.367
R1248 B.n778 B.n284 163.367
R1249 B.n778 B.n282 163.367
R1250 B.n782 B.n282 163.367
R1251 B.n782 B.n3 163.367
R1252 B.n1030 B.n3 163.367
R1253 B.n1026 B.n2 163.367
R1254 B.n1026 B.n1025 163.367
R1255 B.n1025 B.n9 163.367
R1256 B.n1021 B.n9 163.367
R1257 B.n1021 B.n11 163.367
R1258 B.n1017 B.n11 163.367
R1259 B.n1017 B.n16 163.367
R1260 B.n1013 B.n16 163.367
R1261 B.n1013 B.n18 163.367
R1262 B.n1009 B.n18 163.367
R1263 B.n1009 B.n24 163.367
R1264 B.n1005 B.n24 163.367
R1265 B.n1005 B.n26 163.367
R1266 B.n1001 B.n26 163.367
R1267 B.n1001 B.n31 163.367
R1268 B.n997 B.n31 163.367
R1269 B.n997 B.n33 163.367
R1270 B.n993 B.n33 163.367
R1271 B.n993 B.n38 163.367
R1272 B.n989 B.n38 163.367
R1273 B.n989 B.n40 163.367
R1274 B.n985 B.n40 163.367
R1275 B.n985 B.n45 163.367
R1276 B.n981 B.n45 163.367
R1277 B.n981 B.n47 163.367
R1278 B.n977 B.n47 163.367
R1279 B.n977 B.n52 163.367
R1280 B.n973 B.n52 163.367
R1281 B.n973 B.n54 163.367
R1282 B.n969 B.n54 163.367
R1283 B.n969 B.n59 163.367
R1284 B.n965 B.n59 163.367
R1285 B.n965 B.n61 163.367
R1286 B.n961 B.n61 163.367
R1287 B.n961 B.n66 163.367
R1288 B.n957 B.n66 163.367
R1289 B.n957 B.n68 163.367
R1290 B.n953 B.n68 163.367
R1291 B.n953 B.n72 163.367
R1292 B.n949 B.n72 163.367
R1293 B.n949 B.n74 163.367
R1294 B.n945 B.n74 163.367
R1295 B.n945 B.n80 163.367
R1296 B.n941 B.n80 163.367
R1297 B.n941 B.n82 163.367
R1298 B.n937 B.n82 163.367
R1299 B.n937 B.n87 163.367
R1300 B.n933 B.n87 163.367
R1301 B.n933 B.n89 163.367
R1302 B.n929 B.n89 163.367
R1303 B.n929 B.n94 163.367
R1304 B.n925 B.n94 163.367
R1305 B.n925 B.n96 163.367
R1306 B.n921 B.n96 163.367
R1307 B.n921 B.n101 163.367
R1308 B.n917 B.n101 163.367
R1309 B.n917 B.n103 163.367
R1310 B.n913 B.n103 163.367
R1311 B.n913 B.n108 163.367
R1312 B.n909 B.n108 163.367
R1313 B.n909 B.n110 163.367
R1314 B.n905 B.n110 163.367
R1315 B.n905 B.n115 163.367
R1316 B.n901 B.n115 163.367
R1317 B.n901 B.n117 163.367
R1318 B.n897 B.n117 163.367
R1319 B.n897 B.n122 163.367
R1320 B.n893 B.n122 163.367
R1321 B.n893 B.n124 163.367
R1322 B.n889 B.n124 163.367
R1323 B.n889 B.n129 163.367
R1324 B.n885 B.n129 163.367
R1325 B.n162 B.t22 140.543
R1326 B.n516 B.t13 140.543
R1327 B.n165 B.t16 140.536
R1328 B.n438 B.t20 140.536
R1329 B.n570 B.n419 120.457
R1330 B.n884 B.n883 120.457
R1331 B.n133 B.n131 71.676
R1332 B.n170 B.n134 71.676
R1333 B.n174 B.n135 71.676
R1334 B.n178 B.n136 71.676
R1335 B.n182 B.n137 71.676
R1336 B.n186 B.n138 71.676
R1337 B.n190 B.n139 71.676
R1338 B.n194 B.n140 71.676
R1339 B.n198 B.n141 71.676
R1340 B.n202 B.n142 71.676
R1341 B.n206 B.n143 71.676
R1342 B.n210 B.n144 71.676
R1343 B.n214 B.n145 71.676
R1344 B.n218 B.n146 71.676
R1345 B.n222 B.n147 71.676
R1346 B.n226 B.n148 71.676
R1347 B.n230 B.n149 71.676
R1348 B.n234 B.n150 71.676
R1349 B.n238 B.n151 71.676
R1350 B.n242 B.n152 71.676
R1351 B.n246 B.n153 71.676
R1352 B.n250 B.n154 71.676
R1353 B.n254 B.n155 71.676
R1354 B.n258 B.n156 71.676
R1355 B.n262 B.n157 71.676
R1356 B.n266 B.n158 71.676
R1357 B.n270 B.n159 71.676
R1358 B.n274 B.n160 71.676
R1359 B.n882 B.n161 71.676
R1360 B.n882 B.n881 71.676
R1361 B.n276 B.n160 71.676
R1362 B.n273 B.n159 71.676
R1363 B.n269 B.n158 71.676
R1364 B.n265 B.n157 71.676
R1365 B.n261 B.n156 71.676
R1366 B.n257 B.n155 71.676
R1367 B.n253 B.n154 71.676
R1368 B.n249 B.n153 71.676
R1369 B.n245 B.n152 71.676
R1370 B.n241 B.n151 71.676
R1371 B.n237 B.n150 71.676
R1372 B.n233 B.n149 71.676
R1373 B.n229 B.n148 71.676
R1374 B.n225 B.n147 71.676
R1375 B.n221 B.n146 71.676
R1376 B.n217 B.n145 71.676
R1377 B.n213 B.n144 71.676
R1378 B.n209 B.n143 71.676
R1379 B.n205 B.n142 71.676
R1380 B.n201 B.n141 71.676
R1381 B.n197 B.n140 71.676
R1382 B.n193 B.n139 71.676
R1383 B.n189 B.n138 71.676
R1384 B.n185 B.n137 71.676
R1385 B.n181 B.n136 71.676
R1386 B.n177 B.n135 71.676
R1387 B.n173 B.n134 71.676
R1388 B.n169 B.n133 71.676
R1389 B.n452 B.n418 71.676
R1390 B.n456 B.n455 71.676
R1391 B.n461 B.n460 71.676
R1392 B.n464 B.n463 71.676
R1393 B.n469 B.n468 71.676
R1394 B.n472 B.n471 71.676
R1395 B.n477 B.n476 71.676
R1396 B.n480 B.n479 71.676
R1397 B.n485 B.n484 71.676
R1398 B.n488 B.n487 71.676
R1399 B.n493 B.n492 71.676
R1400 B.n496 B.n495 71.676
R1401 B.n502 B.n501 71.676
R1402 B.n505 B.n504 71.676
R1403 B.n510 B.n509 71.676
R1404 B.n513 B.n512 71.676
R1405 B.n521 B.n520 71.676
R1406 B.n524 B.n523 71.676
R1407 B.n529 B.n528 71.676
R1408 B.n532 B.n531 71.676
R1409 B.n537 B.n536 71.676
R1410 B.n540 B.n539 71.676
R1411 B.n545 B.n544 71.676
R1412 B.n548 B.n547 71.676
R1413 B.n553 B.n552 71.676
R1414 B.n556 B.n555 71.676
R1415 B.n561 B.n560 71.676
R1416 B.n564 B.n563 71.676
R1417 B.n453 B.n452 71.676
R1418 B.n455 B.n449 71.676
R1419 B.n462 B.n461 71.676
R1420 B.n463 B.n447 71.676
R1421 B.n470 B.n469 71.676
R1422 B.n471 B.n445 71.676
R1423 B.n478 B.n477 71.676
R1424 B.n479 B.n443 71.676
R1425 B.n486 B.n485 71.676
R1426 B.n487 B.n441 71.676
R1427 B.n494 B.n493 71.676
R1428 B.n495 B.n437 71.676
R1429 B.n503 B.n502 71.676
R1430 B.n504 B.n435 71.676
R1431 B.n511 B.n510 71.676
R1432 B.n512 B.n433 71.676
R1433 B.n522 B.n521 71.676
R1434 B.n523 B.n431 71.676
R1435 B.n530 B.n529 71.676
R1436 B.n531 B.n429 71.676
R1437 B.n538 B.n537 71.676
R1438 B.n539 B.n427 71.676
R1439 B.n546 B.n545 71.676
R1440 B.n547 B.n425 71.676
R1441 B.n554 B.n553 71.676
R1442 B.n555 B.n423 71.676
R1443 B.n562 B.n561 71.676
R1444 B.n565 B.n564 71.676
R1445 B.n1031 B.n1030 71.676
R1446 B.n1031 B.n2 71.676
R1447 B.n166 B.n165 70.7884
R1448 B.n163 B.n162 70.7884
R1449 B.n517 B.n516 70.7884
R1450 B.n439 B.n438 70.7884
R1451 B.n163 B.t23 69.7558
R1452 B.n517 B.t12 69.7558
R1453 B.n166 B.t17 69.749
R1454 B.n439 B.t19 69.749
R1455 B.n570 B.n415 65.5283
R1456 B.n576 B.n415 65.5283
R1457 B.n576 B.n411 65.5283
R1458 B.n582 B.n411 65.5283
R1459 B.n582 B.n407 65.5283
R1460 B.n588 B.n407 65.5283
R1461 B.n588 B.n403 65.5283
R1462 B.n594 B.n403 65.5283
R1463 B.n600 B.n399 65.5283
R1464 B.n600 B.n395 65.5283
R1465 B.n606 B.n395 65.5283
R1466 B.n606 B.n391 65.5283
R1467 B.n612 B.n391 65.5283
R1468 B.n612 B.n387 65.5283
R1469 B.n618 B.n387 65.5283
R1470 B.n618 B.n383 65.5283
R1471 B.n624 B.n383 65.5283
R1472 B.n624 B.n379 65.5283
R1473 B.n630 B.n379 65.5283
R1474 B.n630 B.n375 65.5283
R1475 B.n636 B.n375 65.5283
R1476 B.n642 B.n371 65.5283
R1477 B.n642 B.n367 65.5283
R1478 B.n648 B.n367 65.5283
R1479 B.n648 B.n363 65.5283
R1480 B.n654 B.n363 65.5283
R1481 B.n654 B.n359 65.5283
R1482 B.n660 B.n359 65.5283
R1483 B.n660 B.n355 65.5283
R1484 B.n667 B.n355 65.5283
R1485 B.n667 B.n666 65.5283
R1486 B.n673 B.n348 65.5283
R1487 B.n679 B.n348 65.5283
R1488 B.n679 B.n344 65.5283
R1489 B.n685 B.n344 65.5283
R1490 B.n685 B.n340 65.5283
R1491 B.n691 B.n340 65.5283
R1492 B.n691 B.n336 65.5283
R1493 B.n697 B.n336 65.5283
R1494 B.n697 B.n332 65.5283
R1495 B.n703 B.n332 65.5283
R1496 B.n709 B.n328 65.5283
R1497 B.n709 B.n324 65.5283
R1498 B.n715 B.n324 65.5283
R1499 B.n715 B.n320 65.5283
R1500 B.n721 B.n320 65.5283
R1501 B.n721 B.n316 65.5283
R1502 B.n727 B.n316 65.5283
R1503 B.n727 B.n312 65.5283
R1504 B.n733 B.n312 65.5283
R1505 B.n739 B.n308 65.5283
R1506 B.n739 B.n304 65.5283
R1507 B.n745 B.n304 65.5283
R1508 B.n745 B.n300 65.5283
R1509 B.n751 B.n300 65.5283
R1510 B.n751 B.n296 65.5283
R1511 B.n757 B.n296 65.5283
R1512 B.n757 B.n292 65.5283
R1513 B.n764 B.n292 65.5283
R1514 B.n764 B.n763 65.5283
R1515 B.n770 B.n285 65.5283
R1516 B.n777 B.n285 65.5283
R1517 B.n777 B.n281 65.5283
R1518 B.n783 B.n281 65.5283
R1519 B.n783 B.n4 65.5283
R1520 B.n1029 B.n4 65.5283
R1521 B.n1029 B.n1028 65.5283
R1522 B.n1028 B.n1027 65.5283
R1523 B.n1027 B.n8 65.5283
R1524 B.n12 B.n8 65.5283
R1525 B.n1020 B.n12 65.5283
R1526 B.n1020 B.n1019 65.5283
R1527 B.n1019 B.n1018 65.5283
R1528 B.n1012 B.n19 65.5283
R1529 B.n1012 B.n1011 65.5283
R1530 B.n1011 B.n1010 65.5283
R1531 B.n1010 B.n23 65.5283
R1532 B.n1004 B.n23 65.5283
R1533 B.n1004 B.n1003 65.5283
R1534 B.n1003 B.n1002 65.5283
R1535 B.n1002 B.n30 65.5283
R1536 B.n996 B.n30 65.5283
R1537 B.n996 B.n995 65.5283
R1538 B.n994 B.n37 65.5283
R1539 B.n988 B.n37 65.5283
R1540 B.n988 B.n987 65.5283
R1541 B.n987 B.n986 65.5283
R1542 B.n986 B.n44 65.5283
R1543 B.n980 B.n44 65.5283
R1544 B.n980 B.n979 65.5283
R1545 B.n979 B.n978 65.5283
R1546 B.n978 B.n51 65.5283
R1547 B.n972 B.n971 65.5283
R1548 B.n971 B.n970 65.5283
R1549 B.n970 B.n58 65.5283
R1550 B.n964 B.n58 65.5283
R1551 B.n964 B.n963 65.5283
R1552 B.n963 B.n962 65.5283
R1553 B.n962 B.n65 65.5283
R1554 B.n956 B.n65 65.5283
R1555 B.n956 B.n955 65.5283
R1556 B.n955 B.n954 65.5283
R1557 B.n948 B.n75 65.5283
R1558 B.n948 B.n947 65.5283
R1559 B.n947 B.n946 65.5283
R1560 B.n946 B.n79 65.5283
R1561 B.n940 B.n79 65.5283
R1562 B.n940 B.n939 65.5283
R1563 B.n939 B.n938 65.5283
R1564 B.n938 B.n86 65.5283
R1565 B.n932 B.n86 65.5283
R1566 B.n932 B.n931 65.5283
R1567 B.n930 B.n93 65.5283
R1568 B.n924 B.n93 65.5283
R1569 B.n924 B.n923 65.5283
R1570 B.n923 B.n922 65.5283
R1571 B.n922 B.n100 65.5283
R1572 B.n916 B.n100 65.5283
R1573 B.n916 B.n915 65.5283
R1574 B.n915 B.n914 65.5283
R1575 B.n914 B.n107 65.5283
R1576 B.n908 B.n107 65.5283
R1577 B.n908 B.n907 65.5283
R1578 B.n907 B.n906 65.5283
R1579 B.n906 B.n114 65.5283
R1580 B.n900 B.n899 65.5283
R1581 B.n899 B.n898 65.5283
R1582 B.n898 B.n121 65.5283
R1583 B.n892 B.n121 65.5283
R1584 B.n892 B.n891 65.5283
R1585 B.n891 B.n890 65.5283
R1586 B.n890 B.n128 65.5283
R1587 B.n884 B.n128 65.5283
R1588 B.t8 B.n328 61.6737
R1589 B.t9 B.n51 61.6737
R1590 B.n167 B.n166 59.5399
R1591 B.n164 B.n163 59.5399
R1592 B.n518 B.n517 59.5399
R1593 B.n498 B.n439 59.5399
R1594 B.n733 B.t7 52.0373
R1595 B.t3 B.n994 52.0373
R1596 B.n673 B.t1 44.3281
R1597 B.n954 B.t2 44.3281
R1598 B.n594 B.t11 42.4009
R1599 B.n900 B.t15 42.4009
R1600 B.n636 B.t0 38.5463
R1601 B.t5 B.n930 38.5463
R1602 B.n763 B.t6 34.6917
R1603 B.n19 B.t4 34.6917
R1604 B.n572 B.n417 34.4981
R1605 B.n568 B.n567 34.4981
R1606 B.n880 B.n879 34.4981
R1607 B.n886 B.n130 34.4981
R1608 B.n770 B.t6 30.8371
R1609 B.n1018 B.t4 30.8371
R1610 B.t0 B.n371 26.9825
R1611 B.n931 B.t5 26.9825
R1612 B.t11 B.n399 23.128
R1613 B.t15 B.n114 23.128
R1614 B.n666 B.t1 21.2007
R1615 B.n75 B.t2 21.2007
R1616 B B.n1032 18.0485
R1617 B.t7 B.n308 13.4915
R1618 B.n995 B.t3 13.4915
R1619 B.n573 B.n572 10.6151
R1620 B.n574 B.n573 10.6151
R1621 B.n574 B.n409 10.6151
R1622 B.n584 B.n409 10.6151
R1623 B.n585 B.n584 10.6151
R1624 B.n586 B.n585 10.6151
R1625 B.n586 B.n401 10.6151
R1626 B.n596 B.n401 10.6151
R1627 B.n597 B.n596 10.6151
R1628 B.n598 B.n597 10.6151
R1629 B.n598 B.n393 10.6151
R1630 B.n608 B.n393 10.6151
R1631 B.n609 B.n608 10.6151
R1632 B.n610 B.n609 10.6151
R1633 B.n610 B.n385 10.6151
R1634 B.n620 B.n385 10.6151
R1635 B.n621 B.n620 10.6151
R1636 B.n622 B.n621 10.6151
R1637 B.n622 B.n377 10.6151
R1638 B.n632 B.n377 10.6151
R1639 B.n633 B.n632 10.6151
R1640 B.n634 B.n633 10.6151
R1641 B.n634 B.n369 10.6151
R1642 B.n644 B.n369 10.6151
R1643 B.n645 B.n644 10.6151
R1644 B.n646 B.n645 10.6151
R1645 B.n646 B.n361 10.6151
R1646 B.n656 B.n361 10.6151
R1647 B.n657 B.n656 10.6151
R1648 B.n658 B.n657 10.6151
R1649 B.n658 B.n353 10.6151
R1650 B.n669 B.n353 10.6151
R1651 B.n670 B.n669 10.6151
R1652 B.n671 B.n670 10.6151
R1653 B.n671 B.n346 10.6151
R1654 B.n681 B.n346 10.6151
R1655 B.n682 B.n681 10.6151
R1656 B.n683 B.n682 10.6151
R1657 B.n683 B.n338 10.6151
R1658 B.n693 B.n338 10.6151
R1659 B.n694 B.n693 10.6151
R1660 B.n695 B.n694 10.6151
R1661 B.n695 B.n330 10.6151
R1662 B.n705 B.n330 10.6151
R1663 B.n706 B.n705 10.6151
R1664 B.n707 B.n706 10.6151
R1665 B.n707 B.n322 10.6151
R1666 B.n717 B.n322 10.6151
R1667 B.n718 B.n717 10.6151
R1668 B.n719 B.n718 10.6151
R1669 B.n719 B.n314 10.6151
R1670 B.n729 B.n314 10.6151
R1671 B.n730 B.n729 10.6151
R1672 B.n731 B.n730 10.6151
R1673 B.n731 B.n306 10.6151
R1674 B.n741 B.n306 10.6151
R1675 B.n742 B.n741 10.6151
R1676 B.n743 B.n742 10.6151
R1677 B.n743 B.n298 10.6151
R1678 B.n753 B.n298 10.6151
R1679 B.n754 B.n753 10.6151
R1680 B.n755 B.n754 10.6151
R1681 B.n755 B.n290 10.6151
R1682 B.n766 B.n290 10.6151
R1683 B.n767 B.n766 10.6151
R1684 B.n768 B.n767 10.6151
R1685 B.n768 B.n283 10.6151
R1686 B.n779 B.n283 10.6151
R1687 B.n780 B.n779 10.6151
R1688 B.n781 B.n780 10.6151
R1689 B.n781 B.n0 10.6151
R1690 B.n451 B.n417 10.6151
R1691 B.n451 B.n450 10.6151
R1692 B.n457 B.n450 10.6151
R1693 B.n458 B.n457 10.6151
R1694 B.n459 B.n458 10.6151
R1695 B.n459 B.n448 10.6151
R1696 B.n465 B.n448 10.6151
R1697 B.n466 B.n465 10.6151
R1698 B.n467 B.n466 10.6151
R1699 B.n467 B.n446 10.6151
R1700 B.n473 B.n446 10.6151
R1701 B.n474 B.n473 10.6151
R1702 B.n475 B.n474 10.6151
R1703 B.n475 B.n444 10.6151
R1704 B.n481 B.n444 10.6151
R1705 B.n482 B.n481 10.6151
R1706 B.n483 B.n482 10.6151
R1707 B.n483 B.n442 10.6151
R1708 B.n489 B.n442 10.6151
R1709 B.n490 B.n489 10.6151
R1710 B.n491 B.n490 10.6151
R1711 B.n491 B.n440 10.6151
R1712 B.n497 B.n440 10.6151
R1713 B.n500 B.n499 10.6151
R1714 B.n500 B.n436 10.6151
R1715 B.n506 B.n436 10.6151
R1716 B.n507 B.n506 10.6151
R1717 B.n508 B.n507 10.6151
R1718 B.n508 B.n434 10.6151
R1719 B.n514 B.n434 10.6151
R1720 B.n515 B.n514 10.6151
R1721 B.n519 B.n515 10.6151
R1722 B.n525 B.n432 10.6151
R1723 B.n526 B.n525 10.6151
R1724 B.n527 B.n526 10.6151
R1725 B.n527 B.n430 10.6151
R1726 B.n533 B.n430 10.6151
R1727 B.n534 B.n533 10.6151
R1728 B.n535 B.n534 10.6151
R1729 B.n535 B.n428 10.6151
R1730 B.n541 B.n428 10.6151
R1731 B.n542 B.n541 10.6151
R1732 B.n543 B.n542 10.6151
R1733 B.n543 B.n426 10.6151
R1734 B.n549 B.n426 10.6151
R1735 B.n550 B.n549 10.6151
R1736 B.n551 B.n550 10.6151
R1737 B.n551 B.n424 10.6151
R1738 B.n557 B.n424 10.6151
R1739 B.n558 B.n557 10.6151
R1740 B.n559 B.n558 10.6151
R1741 B.n559 B.n422 10.6151
R1742 B.n422 B.n421 10.6151
R1743 B.n566 B.n421 10.6151
R1744 B.n567 B.n566 10.6151
R1745 B.n568 B.n413 10.6151
R1746 B.n578 B.n413 10.6151
R1747 B.n579 B.n578 10.6151
R1748 B.n580 B.n579 10.6151
R1749 B.n580 B.n405 10.6151
R1750 B.n590 B.n405 10.6151
R1751 B.n591 B.n590 10.6151
R1752 B.n592 B.n591 10.6151
R1753 B.n592 B.n397 10.6151
R1754 B.n602 B.n397 10.6151
R1755 B.n603 B.n602 10.6151
R1756 B.n604 B.n603 10.6151
R1757 B.n604 B.n389 10.6151
R1758 B.n614 B.n389 10.6151
R1759 B.n615 B.n614 10.6151
R1760 B.n616 B.n615 10.6151
R1761 B.n616 B.n381 10.6151
R1762 B.n626 B.n381 10.6151
R1763 B.n627 B.n626 10.6151
R1764 B.n628 B.n627 10.6151
R1765 B.n628 B.n373 10.6151
R1766 B.n638 B.n373 10.6151
R1767 B.n639 B.n638 10.6151
R1768 B.n640 B.n639 10.6151
R1769 B.n640 B.n365 10.6151
R1770 B.n650 B.n365 10.6151
R1771 B.n651 B.n650 10.6151
R1772 B.n652 B.n651 10.6151
R1773 B.n652 B.n357 10.6151
R1774 B.n662 B.n357 10.6151
R1775 B.n663 B.n662 10.6151
R1776 B.n664 B.n663 10.6151
R1777 B.n664 B.n350 10.6151
R1778 B.n675 B.n350 10.6151
R1779 B.n676 B.n675 10.6151
R1780 B.n677 B.n676 10.6151
R1781 B.n677 B.n342 10.6151
R1782 B.n687 B.n342 10.6151
R1783 B.n688 B.n687 10.6151
R1784 B.n689 B.n688 10.6151
R1785 B.n689 B.n334 10.6151
R1786 B.n699 B.n334 10.6151
R1787 B.n700 B.n699 10.6151
R1788 B.n701 B.n700 10.6151
R1789 B.n701 B.n326 10.6151
R1790 B.n711 B.n326 10.6151
R1791 B.n712 B.n711 10.6151
R1792 B.n713 B.n712 10.6151
R1793 B.n713 B.n318 10.6151
R1794 B.n723 B.n318 10.6151
R1795 B.n724 B.n723 10.6151
R1796 B.n725 B.n724 10.6151
R1797 B.n725 B.n310 10.6151
R1798 B.n735 B.n310 10.6151
R1799 B.n736 B.n735 10.6151
R1800 B.n737 B.n736 10.6151
R1801 B.n737 B.n302 10.6151
R1802 B.n747 B.n302 10.6151
R1803 B.n748 B.n747 10.6151
R1804 B.n749 B.n748 10.6151
R1805 B.n749 B.n294 10.6151
R1806 B.n759 B.n294 10.6151
R1807 B.n760 B.n759 10.6151
R1808 B.n761 B.n760 10.6151
R1809 B.n761 B.n287 10.6151
R1810 B.n772 B.n287 10.6151
R1811 B.n773 B.n772 10.6151
R1812 B.n775 B.n773 10.6151
R1813 B.n775 B.n774 10.6151
R1814 B.n774 B.n279 10.6151
R1815 B.n786 B.n279 10.6151
R1816 B.n787 B.n786 10.6151
R1817 B.n788 B.n787 10.6151
R1818 B.n789 B.n788 10.6151
R1819 B.n790 B.n789 10.6151
R1820 B.n793 B.n790 10.6151
R1821 B.n794 B.n793 10.6151
R1822 B.n795 B.n794 10.6151
R1823 B.n796 B.n795 10.6151
R1824 B.n798 B.n796 10.6151
R1825 B.n799 B.n798 10.6151
R1826 B.n800 B.n799 10.6151
R1827 B.n801 B.n800 10.6151
R1828 B.n803 B.n801 10.6151
R1829 B.n804 B.n803 10.6151
R1830 B.n805 B.n804 10.6151
R1831 B.n806 B.n805 10.6151
R1832 B.n808 B.n806 10.6151
R1833 B.n809 B.n808 10.6151
R1834 B.n810 B.n809 10.6151
R1835 B.n811 B.n810 10.6151
R1836 B.n813 B.n811 10.6151
R1837 B.n814 B.n813 10.6151
R1838 B.n815 B.n814 10.6151
R1839 B.n816 B.n815 10.6151
R1840 B.n818 B.n816 10.6151
R1841 B.n819 B.n818 10.6151
R1842 B.n820 B.n819 10.6151
R1843 B.n821 B.n820 10.6151
R1844 B.n823 B.n821 10.6151
R1845 B.n824 B.n823 10.6151
R1846 B.n825 B.n824 10.6151
R1847 B.n826 B.n825 10.6151
R1848 B.n828 B.n826 10.6151
R1849 B.n829 B.n828 10.6151
R1850 B.n830 B.n829 10.6151
R1851 B.n831 B.n830 10.6151
R1852 B.n833 B.n831 10.6151
R1853 B.n834 B.n833 10.6151
R1854 B.n835 B.n834 10.6151
R1855 B.n836 B.n835 10.6151
R1856 B.n838 B.n836 10.6151
R1857 B.n839 B.n838 10.6151
R1858 B.n840 B.n839 10.6151
R1859 B.n841 B.n840 10.6151
R1860 B.n843 B.n841 10.6151
R1861 B.n844 B.n843 10.6151
R1862 B.n845 B.n844 10.6151
R1863 B.n846 B.n845 10.6151
R1864 B.n848 B.n846 10.6151
R1865 B.n849 B.n848 10.6151
R1866 B.n850 B.n849 10.6151
R1867 B.n851 B.n850 10.6151
R1868 B.n853 B.n851 10.6151
R1869 B.n854 B.n853 10.6151
R1870 B.n855 B.n854 10.6151
R1871 B.n856 B.n855 10.6151
R1872 B.n858 B.n856 10.6151
R1873 B.n859 B.n858 10.6151
R1874 B.n860 B.n859 10.6151
R1875 B.n861 B.n860 10.6151
R1876 B.n863 B.n861 10.6151
R1877 B.n864 B.n863 10.6151
R1878 B.n865 B.n864 10.6151
R1879 B.n866 B.n865 10.6151
R1880 B.n868 B.n866 10.6151
R1881 B.n869 B.n868 10.6151
R1882 B.n870 B.n869 10.6151
R1883 B.n871 B.n870 10.6151
R1884 B.n873 B.n871 10.6151
R1885 B.n874 B.n873 10.6151
R1886 B.n875 B.n874 10.6151
R1887 B.n876 B.n875 10.6151
R1888 B.n878 B.n876 10.6151
R1889 B.n879 B.n878 10.6151
R1890 B.n1024 B.n1 10.6151
R1891 B.n1024 B.n1023 10.6151
R1892 B.n1023 B.n1022 10.6151
R1893 B.n1022 B.n10 10.6151
R1894 B.n1016 B.n10 10.6151
R1895 B.n1016 B.n1015 10.6151
R1896 B.n1015 B.n1014 10.6151
R1897 B.n1014 B.n17 10.6151
R1898 B.n1008 B.n17 10.6151
R1899 B.n1008 B.n1007 10.6151
R1900 B.n1007 B.n1006 10.6151
R1901 B.n1006 B.n25 10.6151
R1902 B.n1000 B.n25 10.6151
R1903 B.n1000 B.n999 10.6151
R1904 B.n999 B.n998 10.6151
R1905 B.n998 B.n32 10.6151
R1906 B.n992 B.n32 10.6151
R1907 B.n992 B.n991 10.6151
R1908 B.n991 B.n990 10.6151
R1909 B.n990 B.n39 10.6151
R1910 B.n984 B.n39 10.6151
R1911 B.n984 B.n983 10.6151
R1912 B.n983 B.n982 10.6151
R1913 B.n982 B.n46 10.6151
R1914 B.n976 B.n46 10.6151
R1915 B.n976 B.n975 10.6151
R1916 B.n975 B.n974 10.6151
R1917 B.n974 B.n53 10.6151
R1918 B.n968 B.n53 10.6151
R1919 B.n968 B.n967 10.6151
R1920 B.n967 B.n966 10.6151
R1921 B.n966 B.n60 10.6151
R1922 B.n960 B.n60 10.6151
R1923 B.n960 B.n959 10.6151
R1924 B.n959 B.n958 10.6151
R1925 B.n958 B.n67 10.6151
R1926 B.n952 B.n67 10.6151
R1927 B.n952 B.n951 10.6151
R1928 B.n951 B.n950 10.6151
R1929 B.n950 B.n73 10.6151
R1930 B.n944 B.n73 10.6151
R1931 B.n944 B.n943 10.6151
R1932 B.n943 B.n942 10.6151
R1933 B.n942 B.n81 10.6151
R1934 B.n936 B.n81 10.6151
R1935 B.n936 B.n935 10.6151
R1936 B.n935 B.n934 10.6151
R1937 B.n934 B.n88 10.6151
R1938 B.n928 B.n88 10.6151
R1939 B.n928 B.n927 10.6151
R1940 B.n927 B.n926 10.6151
R1941 B.n926 B.n95 10.6151
R1942 B.n920 B.n95 10.6151
R1943 B.n920 B.n919 10.6151
R1944 B.n919 B.n918 10.6151
R1945 B.n918 B.n102 10.6151
R1946 B.n912 B.n102 10.6151
R1947 B.n912 B.n911 10.6151
R1948 B.n911 B.n910 10.6151
R1949 B.n910 B.n109 10.6151
R1950 B.n904 B.n109 10.6151
R1951 B.n904 B.n903 10.6151
R1952 B.n903 B.n902 10.6151
R1953 B.n902 B.n116 10.6151
R1954 B.n896 B.n116 10.6151
R1955 B.n896 B.n895 10.6151
R1956 B.n895 B.n894 10.6151
R1957 B.n894 B.n123 10.6151
R1958 B.n888 B.n123 10.6151
R1959 B.n888 B.n887 10.6151
R1960 B.n887 B.n886 10.6151
R1961 B.n168 B.n130 10.6151
R1962 B.n171 B.n168 10.6151
R1963 B.n172 B.n171 10.6151
R1964 B.n175 B.n172 10.6151
R1965 B.n176 B.n175 10.6151
R1966 B.n179 B.n176 10.6151
R1967 B.n180 B.n179 10.6151
R1968 B.n183 B.n180 10.6151
R1969 B.n184 B.n183 10.6151
R1970 B.n187 B.n184 10.6151
R1971 B.n188 B.n187 10.6151
R1972 B.n191 B.n188 10.6151
R1973 B.n192 B.n191 10.6151
R1974 B.n195 B.n192 10.6151
R1975 B.n196 B.n195 10.6151
R1976 B.n199 B.n196 10.6151
R1977 B.n200 B.n199 10.6151
R1978 B.n203 B.n200 10.6151
R1979 B.n204 B.n203 10.6151
R1980 B.n207 B.n204 10.6151
R1981 B.n208 B.n207 10.6151
R1982 B.n211 B.n208 10.6151
R1983 B.n212 B.n211 10.6151
R1984 B.n216 B.n215 10.6151
R1985 B.n219 B.n216 10.6151
R1986 B.n220 B.n219 10.6151
R1987 B.n223 B.n220 10.6151
R1988 B.n224 B.n223 10.6151
R1989 B.n227 B.n224 10.6151
R1990 B.n228 B.n227 10.6151
R1991 B.n231 B.n228 10.6151
R1992 B.n232 B.n231 10.6151
R1993 B.n236 B.n235 10.6151
R1994 B.n239 B.n236 10.6151
R1995 B.n240 B.n239 10.6151
R1996 B.n243 B.n240 10.6151
R1997 B.n244 B.n243 10.6151
R1998 B.n247 B.n244 10.6151
R1999 B.n248 B.n247 10.6151
R2000 B.n251 B.n248 10.6151
R2001 B.n252 B.n251 10.6151
R2002 B.n255 B.n252 10.6151
R2003 B.n256 B.n255 10.6151
R2004 B.n259 B.n256 10.6151
R2005 B.n260 B.n259 10.6151
R2006 B.n263 B.n260 10.6151
R2007 B.n264 B.n263 10.6151
R2008 B.n267 B.n264 10.6151
R2009 B.n268 B.n267 10.6151
R2010 B.n271 B.n268 10.6151
R2011 B.n272 B.n271 10.6151
R2012 B.n275 B.n272 10.6151
R2013 B.n277 B.n275 10.6151
R2014 B.n278 B.n277 10.6151
R2015 B.n880 B.n278 10.6151
R2016 B.n498 B.n497 9.36635
R2017 B.n518 B.n432 9.36635
R2018 B.n212 B.n167 9.36635
R2019 B.n235 B.n164 9.36635
R2020 B.n1032 B.n0 8.11757
R2021 B.n1032 B.n1 8.11757
R2022 B.n703 B.t8 3.85508
R2023 B.n972 B.t9 3.85508
R2024 B.n499 B.n498 1.24928
R2025 B.n519 B.n518 1.24928
R2026 B.n215 B.n167 1.24928
R2027 B.n232 B.n164 1.24928
R2028 VP.n32 VP.n31 161.3
R2029 VP.n33 VP.n28 161.3
R2030 VP.n35 VP.n34 161.3
R2031 VP.n36 VP.n27 161.3
R2032 VP.n38 VP.n37 161.3
R2033 VP.n39 VP.n26 161.3
R2034 VP.n41 VP.n40 161.3
R2035 VP.n42 VP.n25 161.3
R2036 VP.n44 VP.n43 161.3
R2037 VP.n45 VP.n24 161.3
R2038 VP.n47 VP.n46 161.3
R2039 VP.n48 VP.n23 161.3
R2040 VP.n50 VP.n49 161.3
R2041 VP.n51 VP.n22 161.3
R2042 VP.n53 VP.n52 161.3
R2043 VP.n55 VP.n54 161.3
R2044 VP.n56 VP.n20 161.3
R2045 VP.n58 VP.n57 161.3
R2046 VP.n59 VP.n19 161.3
R2047 VP.n61 VP.n60 161.3
R2048 VP.n62 VP.n18 161.3
R2049 VP.n64 VP.n63 161.3
R2050 VP.n111 VP.n110 161.3
R2051 VP.n109 VP.n1 161.3
R2052 VP.n108 VP.n107 161.3
R2053 VP.n106 VP.n2 161.3
R2054 VP.n105 VP.n104 161.3
R2055 VP.n103 VP.n3 161.3
R2056 VP.n102 VP.n101 161.3
R2057 VP.n100 VP.n99 161.3
R2058 VP.n98 VP.n5 161.3
R2059 VP.n97 VP.n96 161.3
R2060 VP.n95 VP.n6 161.3
R2061 VP.n94 VP.n93 161.3
R2062 VP.n92 VP.n7 161.3
R2063 VP.n91 VP.n90 161.3
R2064 VP.n89 VP.n8 161.3
R2065 VP.n88 VP.n87 161.3
R2066 VP.n86 VP.n9 161.3
R2067 VP.n85 VP.n84 161.3
R2068 VP.n83 VP.n10 161.3
R2069 VP.n82 VP.n81 161.3
R2070 VP.n80 VP.n11 161.3
R2071 VP.n79 VP.n78 161.3
R2072 VP.n77 VP.n76 161.3
R2073 VP.n75 VP.n13 161.3
R2074 VP.n74 VP.n73 161.3
R2075 VP.n72 VP.n14 161.3
R2076 VP.n71 VP.n70 161.3
R2077 VP.n69 VP.n15 161.3
R2078 VP.n68 VP.n67 161.3
R2079 VP.n30 VP.t3 77.543
R2080 VP.n66 VP.n16 75.4905
R2081 VP.n112 VP.n0 75.4905
R2082 VP.n65 VP.n17 75.4905
R2083 VP.n30 VP.n29 67.3352
R2084 VP.n85 VP.n10 56.5617
R2085 VP.n93 VP.n6 56.5617
R2086 VP.n46 VP.n23 56.5617
R2087 VP.n38 VP.n27 56.5617
R2088 VP.n66 VP.n65 52.7079
R2089 VP.n8 VP.t1 44.571
R2090 VP.n16 VP.t2 44.571
R2091 VP.n12 VP.t8 44.571
R2092 VP.n4 VP.t6 44.571
R2093 VP.n0 VP.t9 44.571
R2094 VP.n25 VP.t0 44.571
R2095 VP.n17 VP.t7 44.571
R2096 VP.n21 VP.t4 44.571
R2097 VP.n29 VP.t5 44.571
R2098 VP.n74 VP.n14 42.999
R2099 VP.n104 VP.n2 42.999
R2100 VP.n57 VP.n19 42.999
R2101 VP.n70 VP.n14 38.1551
R2102 VP.n108 VP.n2 38.1551
R2103 VP.n61 VP.n19 38.1551
R2104 VP.n69 VP.n68 24.5923
R2105 VP.n70 VP.n69 24.5923
R2106 VP.n75 VP.n74 24.5923
R2107 VP.n76 VP.n75 24.5923
R2108 VP.n80 VP.n79 24.5923
R2109 VP.n81 VP.n80 24.5923
R2110 VP.n81 VP.n10 24.5923
R2111 VP.n86 VP.n85 24.5923
R2112 VP.n87 VP.n86 24.5923
R2113 VP.n87 VP.n8 24.5923
R2114 VP.n91 VP.n8 24.5923
R2115 VP.n92 VP.n91 24.5923
R2116 VP.n93 VP.n92 24.5923
R2117 VP.n97 VP.n6 24.5923
R2118 VP.n98 VP.n97 24.5923
R2119 VP.n99 VP.n98 24.5923
R2120 VP.n103 VP.n102 24.5923
R2121 VP.n104 VP.n103 24.5923
R2122 VP.n109 VP.n108 24.5923
R2123 VP.n110 VP.n109 24.5923
R2124 VP.n62 VP.n61 24.5923
R2125 VP.n63 VP.n62 24.5923
R2126 VP.n50 VP.n23 24.5923
R2127 VP.n51 VP.n50 24.5923
R2128 VP.n52 VP.n51 24.5923
R2129 VP.n56 VP.n55 24.5923
R2130 VP.n57 VP.n56 24.5923
R2131 VP.n39 VP.n38 24.5923
R2132 VP.n40 VP.n39 24.5923
R2133 VP.n40 VP.n25 24.5923
R2134 VP.n44 VP.n25 24.5923
R2135 VP.n45 VP.n44 24.5923
R2136 VP.n46 VP.n45 24.5923
R2137 VP.n33 VP.n32 24.5923
R2138 VP.n34 VP.n33 24.5923
R2139 VP.n34 VP.n27 24.5923
R2140 VP.n76 VP.n12 17.2148
R2141 VP.n102 VP.n4 17.2148
R2142 VP.n55 VP.n21 17.2148
R2143 VP.n68 VP.n16 14.7556
R2144 VP.n110 VP.n0 14.7556
R2145 VP.n63 VP.n17 14.7556
R2146 VP.n79 VP.n12 7.37805
R2147 VP.n99 VP.n4 7.37805
R2148 VP.n52 VP.n21 7.37805
R2149 VP.n32 VP.n29 7.37805
R2150 VP.n31 VP.n30 4.14747
R2151 VP.n65 VP.n64 0.354861
R2152 VP.n67 VP.n66 0.354861
R2153 VP.n112 VP.n111 0.354861
R2154 VP VP.n112 0.267071
R2155 VP.n31 VP.n28 0.189894
R2156 VP.n35 VP.n28 0.189894
R2157 VP.n36 VP.n35 0.189894
R2158 VP.n37 VP.n36 0.189894
R2159 VP.n37 VP.n26 0.189894
R2160 VP.n41 VP.n26 0.189894
R2161 VP.n42 VP.n41 0.189894
R2162 VP.n43 VP.n42 0.189894
R2163 VP.n43 VP.n24 0.189894
R2164 VP.n47 VP.n24 0.189894
R2165 VP.n48 VP.n47 0.189894
R2166 VP.n49 VP.n48 0.189894
R2167 VP.n49 VP.n22 0.189894
R2168 VP.n53 VP.n22 0.189894
R2169 VP.n54 VP.n53 0.189894
R2170 VP.n54 VP.n20 0.189894
R2171 VP.n58 VP.n20 0.189894
R2172 VP.n59 VP.n58 0.189894
R2173 VP.n60 VP.n59 0.189894
R2174 VP.n60 VP.n18 0.189894
R2175 VP.n64 VP.n18 0.189894
R2176 VP.n67 VP.n15 0.189894
R2177 VP.n71 VP.n15 0.189894
R2178 VP.n72 VP.n71 0.189894
R2179 VP.n73 VP.n72 0.189894
R2180 VP.n73 VP.n13 0.189894
R2181 VP.n77 VP.n13 0.189894
R2182 VP.n78 VP.n77 0.189894
R2183 VP.n78 VP.n11 0.189894
R2184 VP.n82 VP.n11 0.189894
R2185 VP.n83 VP.n82 0.189894
R2186 VP.n84 VP.n83 0.189894
R2187 VP.n84 VP.n9 0.189894
R2188 VP.n88 VP.n9 0.189894
R2189 VP.n89 VP.n88 0.189894
R2190 VP.n90 VP.n89 0.189894
R2191 VP.n90 VP.n7 0.189894
R2192 VP.n94 VP.n7 0.189894
R2193 VP.n95 VP.n94 0.189894
R2194 VP.n96 VP.n95 0.189894
R2195 VP.n96 VP.n5 0.189894
R2196 VP.n100 VP.n5 0.189894
R2197 VP.n101 VP.n100 0.189894
R2198 VP.n101 VP.n3 0.189894
R2199 VP.n105 VP.n3 0.189894
R2200 VP.n106 VP.n105 0.189894
R2201 VP.n107 VP.n106 0.189894
R2202 VP.n107 VP.n1 0.189894
R2203 VP.n111 VP.n1 0.189894
R2204 VDD1.n1 VDD1.t6 74.9485
R2205 VDD1.n3 VDD1.t7 74.9475
R2206 VDD1.n5 VDD1.n4 70.8816
R2207 VDD1.n1 VDD1.n0 68.5772
R2208 VDD1.n3 VDD1.n2 68.5771
R2209 VDD1.n7 VDD1.n6 68.5763
R2210 VDD1.n7 VDD1.n5 46.1108
R2211 VDD1.n6 VDD1.t5 3.22526
R2212 VDD1.n6 VDD1.t2 3.22526
R2213 VDD1.n0 VDD1.t4 3.22526
R2214 VDD1.n0 VDD1.t9 3.22526
R2215 VDD1.n4 VDD1.t3 3.22526
R2216 VDD1.n4 VDD1.t0 3.22526
R2217 VDD1.n2 VDD1.t1 3.22526
R2218 VDD1.n2 VDD1.t8 3.22526
R2219 VDD1 VDD1.n7 2.30222
R2220 VDD1 VDD1.n1 0.845328
R2221 VDD1.n5 VDD1.n3 0.731792
C0 VTAIL VDD2 8.34105f
C1 VDD1 VP 6.48716f
C2 VDD1 VDD2 2.64226f
C3 VP VDD2 0.675307f
C4 VTAIL VN 7.44331f
C5 VDD1 VN 0.155254f
C6 VP VN 8.367339f
C7 VDD2 VN 5.97019f
C8 VDD1 VTAIL 8.28358f
C9 VTAIL VP 7.457479f
C10 VDD2 B 7.063401f
C11 VDD1 B 6.997525f
C12 VTAIL B 5.848364f
C13 VN B 20.91988f
C14 VP B 19.475908f
C15 VDD1.t6 B 1.43305f
C16 VDD1.t4 B 0.131514f
C17 VDD1.t9 B 0.131514f
C18 VDD1.n0 B 1.11119f
C19 VDD1.n1 B 1.08946f
C20 VDD1.t7 B 1.43306f
C21 VDD1.t1 B 0.131514f
C22 VDD1.t8 B 0.131514f
C23 VDD1.n2 B 1.11118f
C24 VDD1.n3 B 1.0804f
C25 VDD1.t3 B 0.131514f
C26 VDD1.t0 B 0.131514f
C27 VDD1.n4 B 1.13383f
C28 VDD1.n5 B 3.3066f
C29 VDD1.t5 B 0.131514f
C30 VDD1.t2 B 0.131514f
C31 VDD1.n6 B 1.11118f
C32 VDD1.n7 B 3.26312f
C33 VP.t9 B 1.1608f
C34 VP.n0 B 0.513277f
C35 VP.n1 B 0.021486f
C36 VP.n2 B 0.017525f
C37 VP.n3 B 0.021486f
C38 VP.t6 B 1.1608f
C39 VP.n4 B 0.428816f
C40 VP.n5 B 0.021486f
C41 VP.n6 B 0.026775f
C42 VP.n7 B 0.021486f
C43 VP.t1 B 1.1608f
C44 VP.n8 B 0.44899f
C45 VP.n9 B 0.021486f
C46 VP.n10 B 0.026775f
C47 VP.n11 B 0.021486f
C48 VP.t8 B 1.1608f
C49 VP.n12 B 0.428816f
C50 VP.n13 B 0.021486f
C51 VP.n14 B 0.017525f
C52 VP.n15 B 0.021486f
C53 VP.t2 B 1.1608f
C54 VP.n16 B 0.513277f
C55 VP.t7 B 1.1608f
C56 VP.n17 B 0.513277f
C57 VP.n18 B 0.021486f
C58 VP.n19 B 0.017525f
C59 VP.n20 B 0.021486f
C60 VP.t4 B 1.1608f
C61 VP.n21 B 0.428816f
C62 VP.n22 B 0.021486f
C63 VP.n23 B 0.026775f
C64 VP.n24 B 0.021486f
C65 VP.t0 B 1.1608f
C66 VP.n25 B 0.44899f
C67 VP.n26 B 0.021486f
C68 VP.n27 B 0.026775f
C69 VP.n28 B 0.021486f
C70 VP.t5 B 1.1608f
C71 VP.n29 B 0.496766f
C72 VP.t3 B 1.40828f
C73 VP.n30 B 0.474531f
C74 VP.n31 B 0.252938f
C75 VP.n32 B 0.026075f
C76 VP.n33 B 0.039844f
C77 VP.n34 B 0.039844f
C78 VP.n35 B 0.021486f
C79 VP.n36 B 0.021486f
C80 VP.n37 B 0.021486f
C81 VP.n38 B 0.035691f
C82 VP.n39 B 0.039844f
C83 VP.n40 B 0.039844f
C84 VP.n41 B 0.021486f
C85 VP.n42 B 0.021486f
C86 VP.n43 B 0.021486f
C87 VP.n44 B 0.039844f
C88 VP.n45 B 0.039844f
C89 VP.n46 B 0.035691f
C90 VP.n47 B 0.021486f
C91 VP.n48 B 0.021486f
C92 VP.n49 B 0.021486f
C93 VP.n50 B 0.039844f
C94 VP.n51 B 0.039844f
C95 VP.n52 B 0.026075f
C96 VP.n53 B 0.021486f
C97 VP.n54 B 0.021486f
C98 VP.n55 B 0.033943f
C99 VP.n56 B 0.039844f
C100 VP.n57 B 0.041864f
C101 VP.n58 B 0.021486f
C102 VP.n59 B 0.021486f
C103 VP.n60 B 0.021486f
C104 VP.n61 B 0.04292f
C105 VP.n62 B 0.039844f
C106 VP.n63 B 0.031976f
C107 VP.n64 B 0.034672f
C108 VP.n65 B 1.3177f
C109 VP.n66 B 1.3324f
C110 VP.n67 B 0.034672f
C111 VP.n68 B 0.031976f
C112 VP.n69 B 0.039844f
C113 VP.n70 B 0.04292f
C114 VP.n71 B 0.021486f
C115 VP.n72 B 0.021486f
C116 VP.n73 B 0.021486f
C117 VP.n74 B 0.041864f
C118 VP.n75 B 0.039844f
C119 VP.n76 B 0.033943f
C120 VP.n77 B 0.021486f
C121 VP.n78 B 0.021486f
C122 VP.n79 B 0.026075f
C123 VP.n80 B 0.039844f
C124 VP.n81 B 0.039844f
C125 VP.n82 B 0.021486f
C126 VP.n83 B 0.021486f
C127 VP.n84 B 0.021486f
C128 VP.n85 B 0.035691f
C129 VP.n86 B 0.039844f
C130 VP.n87 B 0.039844f
C131 VP.n88 B 0.021486f
C132 VP.n89 B 0.021486f
C133 VP.n90 B 0.021486f
C134 VP.n91 B 0.039844f
C135 VP.n92 B 0.039844f
C136 VP.n93 B 0.035691f
C137 VP.n94 B 0.021486f
C138 VP.n95 B 0.021486f
C139 VP.n96 B 0.021486f
C140 VP.n97 B 0.039844f
C141 VP.n98 B 0.039844f
C142 VP.n99 B 0.026075f
C143 VP.n100 B 0.021486f
C144 VP.n101 B 0.021486f
C145 VP.n102 B 0.033943f
C146 VP.n103 B 0.039844f
C147 VP.n104 B 0.041864f
C148 VP.n105 B 0.021486f
C149 VP.n106 B 0.021486f
C150 VP.n107 B 0.021486f
C151 VP.n108 B 0.04292f
C152 VP.n109 B 0.039844f
C153 VP.n110 B 0.031976f
C154 VP.n111 B 0.034672f
C155 VP.n112 B 0.052118f
C156 VDD2.t8 B 1.39993f
C157 VDD2.t2 B 0.128474f
C158 VDD2.t6 B 0.128474f
C159 VDD2.n0 B 1.0855f
C160 VDD2.n1 B 1.05543f
C161 VDD2.t0 B 0.128474f
C162 VDD2.t3 B 0.128474f
C163 VDD2.n2 B 1.10762f
C164 VDD2.n3 B 3.08238f
C165 VDD2.t9 B 1.37717f
C166 VDD2.n4 B 3.10002f
C167 VDD2.t7 B 0.128474f
C168 VDD2.t5 B 0.128474f
C169 VDD2.n5 B 1.0855f
C170 VDD2.n6 B 0.544866f
C171 VDD2.t1 B 0.128474f
C172 VDD2.t4 B 0.128474f
C173 VDD2.n7 B 1.10758f
C174 VTAIL.t16 B 0.14274f
C175 VTAIL.t17 B 0.14274f
C176 VTAIL.n0 B 1.13488f
C177 VTAIL.n1 B 0.681082f
C178 VTAIL.t6 B 1.44336f
C179 VTAIL.n2 B 0.830946f
C180 VTAIL.t8 B 0.14274f
C181 VTAIL.t7 B 0.14274f
C182 VTAIL.n3 B 1.13488f
C183 VTAIL.n4 B 0.854735f
C184 VTAIL.t0 B 0.14274f
C185 VTAIL.t1 B 0.14274f
C186 VTAIL.n5 B 1.13488f
C187 VTAIL.n6 B 2.05438f
C188 VTAIL.t12 B 0.14274f
C189 VTAIL.t14 B 0.14274f
C190 VTAIL.n7 B 1.13488f
C191 VTAIL.n8 B 2.05438f
C192 VTAIL.t19 B 0.14274f
C193 VTAIL.t10 B 0.14274f
C194 VTAIL.n9 B 1.13488f
C195 VTAIL.n10 B 0.854729f
C196 VTAIL.t18 B 1.44336f
C197 VTAIL.n11 B 0.830945f
C198 VTAIL.t4 B 0.14274f
C199 VTAIL.t3 B 0.14274f
C200 VTAIL.n12 B 1.13488f
C201 VTAIL.n13 B 0.750129f
C202 VTAIL.t9 B 0.14274f
C203 VTAIL.t2 B 0.14274f
C204 VTAIL.n14 B 1.13488f
C205 VTAIL.n15 B 0.854729f
C206 VTAIL.t5 B 1.44335f
C207 VTAIL.n16 B 1.83692f
C208 VTAIL.t11 B 1.44336f
C209 VTAIL.n17 B 1.83692f
C210 VTAIL.t13 B 0.14274f
C211 VTAIL.t15 B 0.14274f
C212 VTAIL.n18 B 1.13488f
C213 VTAIL.n19 B 0.625514f
C214 VN.t6 B 1.12819f
C215 VN.n0 B 0.498856f
C216 VN.n1 B 0.020882f
C217 VN.n2 B 0.017033f
C218 VN.n3 B 0.020882f
C219 VN.t9 B 1.12819f
C220 VN.n4 B 0.416768f
C221 VN.n5 B 0.020882f
C222 VN.n6 B 0.026022f
C223 VN.n7 B 0.020882f
C224 VN.t3 B 1.12819f
C225 VN.n8 B 0.436375f
C226 VN.n9 B 0.020882f
C227 VN.n10 B 0.026022f
C228 VN.n11 B 0.020882f
C229 VN.t7 B 1.12819f
C230 VN.n12 B 0.482809f
C231 VN.t1 B 1.36871f
C232 VN.n13 B 0.461198f
C233 VN.n14 B 0.245831f
C234 VN.n15 B 0.025342f
C235 VN.n16 B 0.038724f
C236 VN.n17 B 0.038724f
C237 VN.n18 B 0.020882f
C238 VN.n19 B 0.020882f
C239 VN.n20 B 0.020882f
C240 VN.n21 B 0.034689f
C241 VN.n22 B 0.038724f
C242 VN.n23 B 0.038724f
C243 VN.n24 B 0.020882f
C244 VN.n25 B 0.020882f
C245 VN.n26 B 0.020882f
C246 VN.n27 B 0.038724f
C247 VN.n28 B 0.038724f
C248 VN.n29 B 0.034689f
C249 VN.n30 B 0.020882f
C250 VN.n31 B 0.020882f
C251 VN.n32 B 0.020882f
C252 VN.n33 B 0.038724f
C253 VN.n34 B 0.038724f
C254 VN.n35 B 0.025342f
C255 VN.n36 B 0.020882f
C256 VN.n37 B 0.020882f
C257 VN.n38 B 0.032989f
C258 VN.n39 B 0.038724f
C259 VN.n40 B 0.040688f
C260 VN.n41 B 0.020882f
C261 VN.n42 B 0.020882f
C262 VN.n43 B 0.020882f
C263 VN.n44 B 0.041714f
C264 VN.n45 B 0.038724f
C265 VN.n46 B 0.031077f
C266 VN.n47 B 0.033698f
C267 VN.n48 B 0.050653f
C268 VN.t0 B 1.12819f
C269 VN.n49 B 0.498856f
C270 VN.n50 B 0.020882f
C271 VN.n51 B 0.017033f
C272 VN.n52 B 0.020882f
C273 VN.t2 B 1.12819f
C274 VN.n53 B 0.416768f
C275 VN.n54 B 0.020882f
C276 VN.n55 B 0.026022f
C277 VN.n56 B 0.020882f
C278 VN.t4 B 1.12819f
C279 VN.n57 B 0.436375f
C280 VN.n58 B 0.020882f
C281 VN.n59 B 0.026022f
C282 VN.n60 B 0.020882f
C283 VN.t8 B 1.12819f
C284 VN.n61 B 0.482809f
C285 VN.t5 B 1.36871f
C286 VN.n62 B 0.461198f
C287 VN.n63 B 0.245831f
C288 VN.n64 B 0.025342f
C289 VN.n65 B 0.038724f
C290 VN.n66 B 0.038724f
C291 VN.n67 B 0.020882f
C292 VN.n68 B 0.020882f
C293 VN.n69 B 0.020882f
C294 VN.n70 B 0.034689f
C295 VN.n71 B 0.038724f
C296 VN.n72 B 0.038724f
C297 VN.n73 B 0.020882f
C298 VN.n74 B 0.020882f
C299 VN.n75 B 0.020882f
C300 VN.n76 B 0.038724f
C301 VN.n77 B 0.038724f
C302 VN.n78 B 0.034689f
C303 VN.n79 B 0.020882f
C304 VN.n80 B 0.020882f
C305 VN.n81 B 0.020882f
C306 VN.n82 B 0.038724f
C307 VN.n83 B 0.038724f
C308 VN.n84 B 0.025342f
C309 VN.n85 B 0.020882f
C310 VN.n86 B 0.020882f
C311 VN.n87 B 0.032989f
C312 VN.n88 B 0.038724f
C313 VN.n89 B 0.040688f
C314 VN.n90 B 0.020882f
C315 VN.n91 B 0.020882f
C316 VN.n92 B 0.020882f
C317 VN.n93 B 0.041714f
C318 VN.n94 B 0.038724f
C319 VN.n95 B 0.031077f
C320 VN.n96 B 0.033698f
C321 VN.n97 B 1.28907f
.ends

