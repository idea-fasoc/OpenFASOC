* NGSPICE file created from diff_pair_sample_0471.ext - technology: sky130A

.subckt diff_pair_sample_0471 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0 ps=0 w=2.12 l=3.62
X1 B.t8 B.t6 B.t7 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0 ps=0 w=2.12 l=3.62
X2 VDD2.t7 VN.t0 VTAIL.t6 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.8268 ps=5.02 w=2.12 l=3.62
X3 VDD1.t7 VP.t0 VTAIL.t14 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=3.62
X4 VDD1.t6 VP.t1 VTAIL.t13 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=3.62
X5 VDD2.t6 VN.t1 VTAIL.t1 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=3.62
X6 VTAIL.t2 VN.t2 VDD2.t5 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=3.62
X7 B.t5 B.t3 B.t4 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0 ps=0 w=2.12 l=3.62
X8 VTAIL.t5 VN.t3 VDD2.t4 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0.3498 ps=2.45 w=2.12 l=3.62
X9 VTAIL.t11 VP.t2 VDD1.t5 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0.3498 ps=2.45 w=2.12 l=3.62
X10 VDD2.t3 VN.t4 VTAIL.t4 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.8268 ps=5.02 w=2.12 l=3.62
X11 VDD1.t4 VP.t3 VTAIL.t8 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.8268 ps=5.02 w=2.12 l=3.62
X12 VTAIL.t3 VN.t5 VDD2.t2 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=3.62
X13 VDD1.t3 VP.t4 VTAIL.t9 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.8268 ps=5.02 w=2.12 l=3.62
X14 B.t2 B.t0 B.t1 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0 ps=0 w=2.12 l=3.62
X15 VDD2.t1 VN.t6 VTAIL.t0 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=3.62
X16 VTAIL.t10 VP.t5 VDD1.t2 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=3.62
X17 VTAIL.t7 VN.t7 VDD2.t0 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0.3498 ps=2.45 w=2.12 l=3.62
X18 VTAIL.t15 VP.t6 VDD1.t1 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.3498 pd=2.45 as=0.3498 ps=2.45 w=2.12 l=3.62
X19 VTAIL.t12 VP.t7 VDD1.t0 w_n4920_n1392# sky130_fd_pr__pfet_01v8 ad=0.8268 pd=5.02 as=0.3498 ps=2.45 w=2.12 l=3.62
R0 B.n530 B.n529 585
R1 B.n531 B.n56 585
R2 B.n533 B.n532 585
R3 B.n534 B.n55 585
R4 B.n536 B.n535 585
R5 B.n537 B.n54 585
R6 B.n539 B.n538 585
R7 B.n540 B.n53 585
R8 B.n542 B.n541 585
R9 B.n543 B.n52 585
R10 B.n545 B.n544 585
R11 B.n546 B.n51 585
R12 B.n548 B.n547 585
R13 B.n550 B.n549 585
R14 B.n551 B.n47 585
R15 B.n553 B.n552 585
R16 B.n554 B.n46 585
R17 B.n556 B.n555 585
R18 B.n557 B.n45 585
R19 B.n559 B.n558 585
R20 B.n560 B.n44 585
R21 B.n562 B.n561 585
R22 B.n564 B.n41 585
R23 B.n566 B.n565 585
R24 B.n567 B.n40 585
R25 B.n569 B.n568 585
R26 B.n570 B.n39 585
R27 B.n572 B.n571 585
R28 B.n573 B.n38 585
R29 B.n575 B.n574 585
R30 B.n576 B.n37 585
R31 B.n578 B.n577 585
R32 B.n579 B.n36 585
R33 B.n581 B.n580 585
R34 B.n582 B.n35 585
R35 B.n528 B.n57 585
R36 B.n527 B.n526 585
R37 B.n525 B.n58 585
R38 B.n524 B.n523 585
R39 B.n522 B.n59 585
R40 B.n521 B.n520 585
R41 B.n519 B.n60 585
R42 B.n518 B.n517 585
R43 B.n516 B.n61 585
R44 B.n515 B.n514 585
R45 B.n513 B.n62 585
R46 B.n512 B.n511 585
R47 B.n510 B.n63 585
R48 B.n509 B.n508 585
R49 B.n507 B.n64 585
R50 B.n506 B.n505 585
R51 B.n504 B.n65 585
R52 B.n503 B.n502 585
R53 B.n501 B.n66 585
R54 B.n500 B.n499 585
R55 B.n498 B.n67 585
R56 B.n497 B.n496 585
R57 B.n495 B.n68 585
R58 B.n494 B.n493 585
R59 B.n492 B.n69 585
R60 B.n491 B.n490 585
R61 B.n489 B.n70 585
R62 B.n488 B.n487 585
R63 B.n486 B.n71 585
R64 B.n485 B.n484 585
R65 B.n483 B.n72 585
R66 B.n482 B.n481 585
R67 B.n480 B.n73 585
R68 B.n479 B.n478 585
R69 B.n477 B.n74 585
R70 B.n476 B.n475 585
R71 B.n474 B.n75 585
R72 B.n473 B.n472 585
R73 B.n471 B.n76 585
R74 B.n470 B.n469 585
R75 B.n468 B.n77 585
R76 B.n467 B.n466 585
R77 B.n465 B.n78 585
R78 B.n464 B.n463 585
R79 B.n462 B.n79 585
R80 B.n461 B.n460 585
R81 B.n459 B.n80 585
R82 B.n458 B.n457 585
R83 B.n456 B.n81 585
R84 B.n455 B.n454 585
R85 B.n453 B.n82 585
R86 B.n452 B.n451 585
R87 B.n450 B.n83 585
R88 B.n449 B.n448 585
R89 B.n447 B.n84 585
R90 B.n446 B.n445 585
R91 B.n444 B.n85 585
R92 B.n443 B.n442 585
R93 B.n441 B.n86 585
R94 B.n440 B.n439 585
R95 B.n438 B.n87 585
R96 B.n437 B.n436 585
R97 B.n435 B.n88 585
R98 B.n434 B.n433 585
R99 B.n432 B.n89 585
R100 B.n431 B.n430 585
R101 B.n429 B.n90 585
R102 B.n428 B.n427 585
R103 B.n426 B.n91 585
R104 B.n425 B.n424 585
R105 B.n423 B.n92 585
R106 B.n422 B.n421 585
R107 B.n420 B.n93 585
R108 B.n419 B.n418 585
R109 B.n417 B.n94 585
R110 B.n416 B.n415 585
R111 B.n414 B.n95 585
R112 B.n413 B.n412 585
R113 B.n411 B.n96 585
R114 B.n410 B.n409 585
R115 B.n408 B.n97 585
R116 B.n407 B.n406 585
R117 B.n405 B.n98 585
R118 B.n404 B.n403 585
R119 B.n402 B.n99 585
R120 B.n401 B.n400 585
R121 B.n399 B.n100 585
R122 B.n398 B.n397 585
R123 B.n396 B.n101 585
R124 B.n395 B.n394 585
R125 B.n393 B.n102 585
R126 B.n392 B.n391 585
R127 B.n390 B.n103 585
R128 B.n389 B.n388 585
R129 B.n387 B.n104 585
R130 B.n386 B.n385 585
R131 B.n384 B.n105 585
R132 B.n383 B.n382 585
R133 B.n381 B.n106 585
R134 B.n380 B.n379 585
R135 B.n378 B.n107 585
R136 B.n377 B.n376 585
R137 B.n375 B.n108 585
R138 B.n374 B.n373 585
R139 B.n372 B.n109 585
R140 B.n371 B.n370 585
R141 B.n369 B.n110 585
R142 B.n368 B.n367 585
R143 B.n366 B.n111 585
R144 B.n365 B.n364 585
R145 B.n363 B.n112 585
R146 B.n362 B.n361 585
R147 B.n360 B.n113 585
R148 B.n359 B.n358 585
R149 B.n357 B.n114 585
R150 B.n356 B.n355 585
R151 B.n354 B.n115 585
R152 B.n353 B.n352 585
R153 B.n351 B.n116 585
R154 B.n350 B.n349 585
R155 B.n348 B.n117 585
R156 B.n347 B.n346 585
R157 B.n345 B.n118 585
R158 B.n344 B.n343 585
R159 B.n342 B.n119 585
R160 B.n341 B.n340 585
R161 B.n339 B.n120 585
R162 B.n338 B.n337 585
R163 B.n336 B.n121 585
R164 B.n335 B.n334 585
R165 B.n333 B.n122 585
R166 B.n332 B.n331 585
R167 B.n330 B.n123 585
R168 B.n276 B.n145 585
R169 B.n278 B.n277 585
R170 B.n279 B.n144 585
R171 B.n281 B.n280 585
R172 B.n282 B.n143 585
R173 B.n284 B.n283 585
R174 B.n285 B.n142 585
R175 B.n287 B.n286 585
R176 B.n288 B.n141 585
R177 B.n290 B.n289 585
R178 B.n291 B.n140 585
R179 B.n293 B.n292 585
R180 B.n294 B.n137 585
R181 B.n297 B.n296 585
R182 B.n298 B.n136 585
R183 B.n300 B.n299 585
R184 B.n301 B.n135 585
R185 B.n303 B.n302 585
R186 B.n304 B.n134 585
R187 B.n306 B.n305 585
R188 B.n307 B.n133 585
R189 B.n309 B.n308 585
R190 B.n311 B.n310 585
R191 B.n312 B.n129 585
R192 B.n314 B.n313 585
R193 B.n315 B.n128 585
R194 B.n317 B.n316 585
R195 B.n318 B.n127 585
R196 B.n320 B.n319 585
R197 B.n321 B.n126 585
R198 B.n323 B.n322 585
R199 B.n324 B.n125 585
R200 B.n326 B.n325 585
R201 B.n327 B.n124 585
R202 B.n329 B.n328 585
R203 B.n275 B.n274 585
R204 B.n273 B.n146 585
R205 B.n272 B.n271 585
R206 B.n270 B.n147 585
R207 B.n269 B.n268 585
R208 B.n267 B.n148 585
R209 B.n266 B.n265 585
R210 B.n264 B.n149 585
R211 B.n263 B.n262 585
R212 B.n261 B.n150 585
R213 B.n260 B.n259 585
R214 B.n258 B.n151 585
R215 B.n257 B.n256 585
R216 B.n255 B.n152 585
R217 B.n254 B.n253 585
R218 B.n252 B.n153 585
R219 B.n251 B.n250 585
R220 B.n249 B.n154 585
R221 B.n248 B.n247 585
R222 B.n246 B.n155 585
R223 B.n245 B.n244 585
R224 B.n243 B.n156 585
R225 B.n242 B.n241 585
R226 B.n240 B.n157 585
R227 B.n239 B.n238 585
R228 B.n237 B.n158 585
R229 B.n236 B.n235 585
R230 B.n234 B.n159 585
R231 B.n233 B.n232 585
R232 B.n231 B.n160 585
R233 B.n230 B.n229 585
R234 B.n228 B.n161 585
R235 B.n227 B.n226 585
R236 B.n225 B.n162 585
R237 B.n224 B.n223 585
R238 B.n222 B.n163 585
R239 B.n221 B.n220 585
R240 B.n219 B.n164 585
R241 B.n218 B.n217 585
R242 B.n216 B.n165 585
R243 B.n215 B.n214 585
R244 B.n213 B.n166 585
R245 B.n212 B.n211 585
R246 B.n210 B.n167 585
R247 B.n209 B.n208 585
R248 B.n207 B.n168 585
R249 B.n206 B.n205 585
R250 B.n204 B.n169 585
R251 B.n203 B.n202 585
R252 B.n201 B.n170 585
R253 B.n200 B.n199 585
R254 B.n198 B.n171 585
R255 B.n197 B.n196 585
R256 B.n195 B.n172 585
R257 B.n194 B.n193 585
R258 B.n192 B.n173 585
R259 B.n191 B.n190 585
R260 B.n189 B.n174 585
R261 B.n188 B.n187 585
R262 B.n186 B.n175 585
R263 B.n185 B.n184 585
R264 B.n183 B.n176 585
R265 B.n182 B.n181 585
R266 B.n180 B.n177 585
R267 B.n179 B.n178 585
R268 B.n2 B.n0 585
R269 B.n681 B.n1 585
R270 B.n680 B.n679 585
R271 B.n678 B.n3 585
R272 B.n677 B.n676 585
R273 B.n675 B.n4 585
R274 B.n674 B.n673 585
R275 B.n672 B.n5 585
R276 B.n671 B.n670 585
R277 B.n669 B.n6 585
R278 B.n668 B.n667 585
R279 B.n666 B.n7 585
R280 B.n665 B.n664 585
R281 B.n663 B.n8 585
R282 B.n662 B.n661 585
R283 B.n660 B.n9 585
R284 B.n659 B.n658 585
R285 B.n657 B.n10 585
R286 B.n656 B.n655 585
R287 B.n654 B.n11 585
R288 B.n653 B.n652 585
R289 B.n651 B.n12 585
R290 B.n650 B.n649 585
R291 B.n648 B.n13 585
R292 B.n647 B.n646 585
R293 B.n645 B.n14 585
R294 B.n644 B.n643 585
R295 B.n642 B.n15 585
R296 B.n641 B.n640 585
R297 B.n639 B.n16 585
R298 B.n638 B.n637 585
R299 B.n636 B.n17 585
R300 B.n635 B.n634 585
R301 B.n633 B.n18 585
R302 B.n632 B.n631 585
R303 B.n630 B.n19 585
R304 B.n629 B.n628 585
R305 B.n627 B.n20 585
R306 B.n626 B.n625 585
R307 B.n624 B.n21 585
R308 B.n623 B.n622 585
R309 B.n621 B.n22 585
R310 B.n620 B.n619 585
R311 B.n618 B.n23 585
R312 B.n617 B.n616 585
R313 B.n615 B.n24 585
R314 B.n614 B.n613 585
R315 B.n612 B.n25 585
R316 B.n611 B.n610 585
R317 B.n609 B.n26 585
R318 B.n608 B.n607 585
R319 B.n606 B.n27 585
R320 B.n605 B.n604 585
R321 B.n603 B.n28 585
R322 B.n602 B.n601 585
R323 B.n600 B.n29 585
R324 B.n599 B.n598 585
R325 B.n597 B.n30 585
R326 B.n596 B.n595 585
R327 B.n594 B.n31 585
R328 B.n593 B.n592 585
R329 B.n591 B.n32 585
R330 B.n590 B.n589 585
R331 B.n588 B.n33 585
R332 B.n587 B.n586 585
R333 B.n585 B.n34 585
R334 B.n584 B.n583 585
R335 B.n683 B.n682 585
R336 B.n274 B.n145 506.916
R337 B.n584 B.n35 506.916
R338 B.n328 B.n123 506.916
R339 B.n530 B.n57 506.916
R340 B.n130 B.t8 248.46
R341 B.n48 B.t4 248.46
R342 B.n138 B.t11 248.459
R343 B.n42 B.t1 248.459
R344 B.n130 B.t6 223.312
R345 B.n138 B.t9 223.312
R346 B.n42 B.t0 223.312
R347 B.n48 B.t3 223.312
R348 B.n131 B.t7 171.855
R349 B.n49 B.t5 171.855
R350 B.n139 B.t10 171.853
R351 B.n43 B.t2 171.853
R352 B.n274 B.n273 163.367
R353 B.n273 B.n272 163.367
R354 B.n272 B.n147 163.367
R355 B.n268 B.n147 163.367
R356 B.n268 B.n267 163.367
R357 B.n267 B.n266 163.367
R358 B.n266 B.n149 163.367
R359 B.n262 B.n149 163.367
R360 B.n262 B.n261 163.367
R361 B.n261 B.n260 163.367
R362 B.n260 B.n151 163.367
R363 B.n256 B.n151 163.367
R364 B.n256 B.n255 163.367
R365 B.n255 B.n254 163.367
R366 B.n254 B.n153 163.367
R367 B.n250 B.n153 163.367
R368 B.n250 B.n249 163.367
R369 B.n249 B.n248 163.367
R370 B.n248 B.n155 163.367
R371 B.n244 B.n155 163.367
R372 B.n244 B.n243 163.367
R373 B.n243 B.n242 163.367
R374 B.n242 B.n157 163.367
R375 B.n238 B.n157 163.367
R376 B.n238 B.n237 163.367
R377 B.n237 B.n236 163.367
R378 B.n236 B.n159 163.367
R379 B.n232 B.n159 163.367
R380 B.n232 B.n231 163.367
R381 B.n231 B.n230 163.367
R382 B.n230 B.n161 163.367
R383 B.n226 B.n161 163.367
R384 B.n226 B.n225 163.367
R385 B.n225 B.n224 163.367
R386 B.n224 B.n163 163.367
R387 B.n220 B.n163 163.367
R388 B.n220 B.n219 163.367
R389 B.n219 B.n218 163.367
R390 B.n218 B.n165 163.367
R391 B.n214 B.n165 163.367
R392 B.n214 B.n213 163.367
R393 B.n213 B.n212 163.367
R394 B.n212 B.n167 163.367
R395 B.n208 B.n167 163.367
R396 B.n208 B.n207 163.367
R397 B.n207 B.n206 163.367
R398 B.n206 B.n169 163.367
R399 B.n202 B.n169 163.367
R400 B.n202 B.n201 163.367
R401 B.n201 B.n200 163.367
R402 B.n200 B.n171 163.367
R403 B.n196 B.n171 163.367
R404 B.n196 B.n195 163.367
R405 B.n195 B.n194 163.367
R406 B.n194 B.n173 163.367
R407 B.n190 B.n173 163.367
R408 B.n190 B.n189 163.367
R409 B.n189 B.n188 163.367
R410 B.n188 B.n175 163.367
R411 B.n184 B.n175 163.367
R412 B.n184 B.n183 163.367
R413 B.n183 B.n182 163.367
R414 B.n182 B.n177 163.367
R415 B.n178 B.n177 163.367
R416 B.n178 B.n2 163.367
R417 B.n682 B.n2 163.367
R418 B.n682 B.n681 163.367
R419 B.n681 B.n680 163.367
R420 B.n680 B.n3 163.367
R421 B.n676 B.n3 163.367
R422 B.n676 B.n675 163.367
R423 B.n675 B.n674 163.367
R424 B.n674 B.n5 163.367
R425 B.n670 B.n5 163.367
R426 B.n670 B.n669 163.367
R427 B.n669 B.n668 163.367
R428 B.n668 B.n7 163.367
R429 B.n664 B.n7 163.367
R430 B.n664 B.n663 163.367
R431 B.n663 B.n662 163.367
R432 B.n662 B.n9 163.367
R433 B.n658 B.n9 163.367
R434 B.n658 B.n657 163.367
R435 B.n657 B.n656 163.367
R436 B.n656 B.n11 163.367
R437 B.n652 B.n11 163.367
R438 B.n652 B.n651 163.367
R439 B.n651 B.n650 163.367
R440 B.n650 B.n13 163.367
R441 B.n646 B.n13 163.367
R442 B.n646 B.n645 163.367
R443 B.n645 B.n644 163.367
R444 B.n644 B.n15 163.367
R445 B.n640 B.n15 163.367
R446 B.n640 B.n639 163.367
R447 B.n639 B.n638 163.367
R448 B.n638 B.n17 163.367
R449 B.n634 B.n17 163.367
R450 B.n634 B.n633 163.367
R451 B.n633 B.n632 163.367
R452 B.n632 B.n19 163.367
R453 B.n628 B.n19 163.367
R454 B.n628 B.n627 163.367
R455 B.n627 B.n626 163.367
R456 B.n626 B.n21 163.367
R457 B.n622 B.n21 163.367
R458 B.n622 B.n621 163.367
R459 B.n621 B.n620 163.367
R460 B.n620 B.n23 163.367
R461 B.n616 B.n23 163.367
R462 B.n616 B.n615 163.367
R463 B.n615 B.n614 163.367
R464 B.n614 B.n25 163.367
R465 B.n610 B.n25 163.367
R466 B.n610 B.n609 163.367
R467 B.n609 B.n608 163.367
R468 B.n608 B.n27 163.367
R469 B.n604 B.n27 163.367
R470 B.n604 B.n603 163.367
R471 B.n603 B.n602 163.367
R472 B.n602 B.n29 163.367
R473 B.n598 B.n29 163.367
R474 B.n598 B.n597 163.367
R475 B.n597 B.n596 163.367
R476 B.n596 B.n31 163.367
R477 B.n592 B.n31 163.367
R478 B.n592 B.n591 163.367
R479 B.n591 B.n590 163.367
R480 B.n590 B.n33 163.367
R481 B.n586 B.n33 163.367
R482 B.n586 B.n585 163.367
R483 B.n585 B.n584 163.367
R484 B.n278 B.n145 163.367
R485 B.n279 B.n278 163.367
R486 B.n280 B.n279 163.367
R487 B.n280 B.n143 163.367
R488 B.n284 B.n143 163.367
R489 B.n285 B.n284 163.367
R490 B.n286 B.n285 163.367
R491 B.n286 B.n141 163.367
R492 B.n290 B.n141 163.367
R493 B.n291 B.n290 163.367
R494 B.n292 B.n291 163.367
R495 B.n292 B.n137 163.367
R496 B.n297 B.n137 163.367
R497 B.n298 B.n297 163.367
R498 B.n299 B.n298 163.367
R499 B.n299 B.n135 163.367
R500 B.n303 B.n135 163.367
R501 B.n304 B.n303 163.367
R502 B.n305 B.n304 163.367
R503 B.n305 B.n133 163.367
R504 B.n309 B.n133 163.367
R505 B.n310 B.n309 163.367
R506 B.n310 B.n129 163.367
R507 B.n314 B.n129 163.367
R508 B.n315 B.n314 163.367
R509 B.n316 B.n315 163.367
R510 B.n316 B.n127 163.367
R511 B.n320 B.n127 163.367
R512 B.n321 B.n320 163.367
R513 B.n322 B.n321 163.367
R514 B.n322 B.n125 163.367
R515 B.n326 B.n125 163.367
R516 B.n327 B.n326 163.367
R517 B.n328 B.n327 163.367
R518 B.n332 B.n123 163.367
R519 B.n333 B.n332 163.367
R520 B.n334 B.n333 163.367
R521 B.n334 B.n121 163.367
R522 B.n338 B.n121 163.367
R523 B.n339 B.n338 163.367
R524 B.n340 B.n339 163.367
R525 B.n340 B.n119 163.367
R526 B.n344 B.n119 163.367
R527 B.n345 B.n344 163.367
R528 B.n346 B.n345 163.367
R529 B.n346 B.n117 163.367
R530 B.n350 B.n117 163.367
R531 B.n351 B.n350 163.367
R532 B.n352 B.n351 163.367
R533 B.n352 B.n115 163.367
R534 B.n356 B.n115 163.367
R535 B.n357 B.n356 163.367
R536 B.n358 B.n357 163.367
R537 B.n358 B.n113 163.367
R538 B.n362 B.n113 163.367
R539 B.n363 B.n362 163.367
R540 B.n364 B.n363 163.367
R541 B.n364 B.n111 163.367
R542 B.n368 B.n111 163.367
R543 B.n369 B.n368 163.367
R544 B.n370 B.n369 163.367
R545 B.n370 B.n109 163.367
R546 B.n374 B.n109 163.367
R547 B.n375 B.n374 163.367
R548 B.n376 B.n375 163.367
R549 B.n376 B.n107 163.367
R550 B.n380 B.n107 163.367
R551 B.n381 B.n380 163.367
R552 B.n382 B.n381 163.367
R553 B.n382 B.n105 163.367
R554 B.n386 B.n105 163.367
R555 B.n387 B.n386 163.367
R556 B.n388 B.n387 163.367
R557 B.n388 B.n103 163.367
R558 B.n392 B.n103 163.367
R559 B.n393 B.n392 163.367
R560 B.n394 B.n393 163.367
R561 B.n394 B.n101 163.367
R562 B.n398 B.n101 163.367
R563 B.n399 B.n398 163.367
R564 B.n400 B.n399 163.367
R565 B.n400 B.n99 163.367
R566 B.n404 B.n99 163.367
R567 B.n405 B.n404 163.367
R568 B.n406 B.n405 163.367
R569 B.n406 B.n97 163.367
R570 B.n410 B.n97 163.367
R571 B.n411 B.n410 163.367
R572 B.n412 B.n411 163.367
R573 B.n412 B.n95 163.367
R574 B.n416 B.n95 163.367
R575 B.n417 B.n416 163.367
R576 B.n418 B.n417 163.367
R577 B.n418 B.n93 163.367
R578 B.n422 B.n93 163.367
R579 B.n423 B.n422 163.367
R580 B.n424 B.n423 163.367
R581 B.n424 B.n91 163.367
R582 B.n428 B.n91 163.367
R583 B.n429 B.n428 163.367
R584 B.n430 B.n429 163.367
R585 B.n430 B.n89 163.367
R586 B.n434 B.n89 163.367
R587 B.n435 B.n434 163.367
R588 B.n436 B.n435 163.367
R589 B.n436 B.n87 163.367
R590 B.n440 B.n87 163.367
R591 B.n441 B.n440 163.367
R592 B.n442 B.n441 163.367
R593 B.n442 B.n85 163.367
R594 B.n446 B.n85 163.367
R595 B.n447 B.n446 163.367
R596 B.n448 B.n447 163.367
R597 B.n448 B.n83 163.367
R598 B.n452 B.n83 163.367
R599 B.n453 B.n452 163.367
R600 B.n454 B.n453 163.367
R601 B.n454 B.n81 163.367
R602 B.n458 B.n81 163.367
R603 B.n459 B.n458 163.367
R604 B.n460 B.n459 163.367
R605 B.n460 B.n79 163.367
R606 B.n464 B.n79 163.367
R607 B.n465 B.n464 163.367
R608 B.n466 B.n465 163.367
R609 B.n466 B.n77 163.367
R610 B.n470 B.n77 163.367
R611 B.n471 B.n470 163.367
R612 B.n472 B.n471 163.367
R613 B.n472 B.n75 163.367
R614 B.n476 B.n75 163.367
R615 B.n477 B.n476 163.367
R616 B.n478 B.n477 163.367
R617 B.n478 B.n73 163.367
R618 B.n482 B.n73 163.367
R619 B.n483 B.n482 163.367
R620 B.n484 B.n483 163.367
R621 B.n484 B.n71 163.367
R622 B.n488 B.n71 163.367
R623 B.n489 B.n488 163.367
R624 B.n490 B.n489 163.367
R625 B.n490 B.n69 163.367
R626 B.n494 B.n69 163.367
R627 B.n495 B.n494 163.367
R628 B.n496 B.n495 163.367
R629 B.n496 B.n67 163.367
R630 B.n500 B.n67 163.367
R631 B.n501 B.n500 163.367
R632 B.n502 B.n501 163.367
R633 B.n502 B.n65 163.367
R634 B.n506 B.n65 163.367
R635 B.n507 B.n506 163.367
R636 B.n508 B.n507 163.367
R637 B.n508 B.n63 163.367
R638 B.n512 B.n63 163.367
R639 B.n513 B.n512 163.367
R640 B.n514 B.n513 163.367
R641 B.n514 B.n61 163.367
R642 B.n518 B.n61 163.367
R643 B.n519 B.n518 163.367
R644 B.n520 B.n519 163.367
R645 B.n520 B.n59 163.367
R646 B.n524 B.n59 163.367
R647 B.n525 B.n524 163.367
R648 B.n526 B.n525 163.367
R649 B.n526 B.n57 163.367
R650 B.n580 B.n35 163.367
R651 B.n580 B.n579 163.367
R652 B.n579 B.n578 163.367
R653 B.n578 B.n37 163.367
R654 B.n574 B.n37 163.367
R655 B.n574 B.n573 163.367
R656 B.n573 B.n572 163.367
R657 B.n572 B.n39 163.367
R658 B.n568 B.n39 163.367
R659 B.n568 B.n567 163.367
R660 B.n567 B.n566 163.367
R661 B.n566 B.n41 163.367
R662 B.n561 B.n41 163.367
R663 B.n561 B.n560 163.367
R664 B.n560 B.n559 163.367
R665 B.n559 B.n45 163.367
R666 B.n555 B.n45 163.367
R667 B.n555 B.n554 163.367
R668 B.n554 B.n553 163.367
R669 B.n553 B.n47 163.367
R670 B.n549 B.n47 163.367
R671 B.n549 B.n548 163.367
R672 B.n548 B.n51 163.367
R673 B.n544 B.n51 163.367
R674 B.n544 B.n543 163.367
R675 B.n543 B.n542 163.367
R676 B.n542 B.n53 163.367
R677 B.n538 B.n53 163.367
R678 B.n538 B.n537 163.367
R679 B.n537 B.n536 163.367
R680 B.n536 B.n55 163.367
R681 B.n532 B.n55 163.367
R682 B.n532 B.n531 163.367
R683 B.n531 B.n530 163.367
R684 B.n131 B.n130 76.6066
R685 B.n139 B.n138 76.6066
R686 B.n43 B.n42 76.6066
R687 B.n49 B.n48 76.6066
R688 B.n132 B.n131 59.5399
R689 B.n295 B.n139 59.5399
R690 B.n563 B.n43 59.5399
R691 B.n50 B.n49 59.5399
R692 B.n583 B.n582 32.9371
R693 B.n529 B.n528 32.9371
R694 B.n330 B.n329 32.9371
R695 B.n276 B.n275 32.9371
R696 B B.n683 18.0485
R697 B.n582 B.n581 10.6151
R698 B.n581 B.n36 10.6151
R699 B.n577 B.n36 10.6151
R700 B.n577 B.n576 10.6151
R701 B.n576 B.n575 10.6151
R702 B.n575 B.n38 10.6151
R703 B.n571 B.n38 10.6151
R704 B.n571 B.n570 10.6151
R705 B.n570 B.n569 10.6151
R706 B.n569 B.n40 10.6151
R707 B.n565 B.n40 10.6151
R708 B.n565 B.n564 10.6151
R709 B.n562 B.n44 10.6151
R710 B.n558 B.n44 10.6151
R711 B.n558 B.n557 10.6151
R712 B.n557 B.n556 10.6151
R713 B.n556 B.n46 10.6151
R714 B.n552 B.n46 10.6151
R715 B.n552 B.n551 10.6151
R716 B.n551 B.n550 10.6151
R717 B.n547 B.n546 10.6151
R718 B.n546 B.n545 10.6151
R719 B.n545 B.n52 10.6151
R720 B.n541 B.n52 10.6151
R721 B.n541 B.n540 10.6151
R722 B.n540 B.n539 10.6151
R723 B.n539 B.n54 10.6151
R724 B.n535 B.n54 10.6151
R725 B.n535 B.n534 10.6151
R726 B.n534 B.n533 10.6151
R727 B.n533 B.n56 10.6151
R728 B.n529 B.n56 10.6151
R729 B.n331 B.n330 10.6151
R730 B.n331 B.n122 10.6151
R731 B.n335 B.n122 10.6151
R732 B.n336 B.n335 10.6151
R733 B.n337 B.n336 10.6151
R734 B.n337 B.n120 10.6151
R735 B.n341 B.n120 10.6151
R736 B.n342 B.n341 10.6151
R737 B.n343 B.n342 10.6151
R738 B.n343 B.n118 10.6151
R739 B.n347 B.n118 10.6151
R740 B.n348 B.n347 10.6151
R741 B.n349 B.n348 10.6151
R742 B.n349 B.n116 10.6151
R743 B.n353 B.n116 10.6151
R744 B.n354 B.n353 10.6151
R745 B.n355 B.n354 10.6151
R746 B.n355 B.n114 10.6151
R747 B.n359 B.n114 10.6151
R748 B.n360 B.n359 10.6151
R749 B.n361 B.n360 10.6151
R750 B.n361 B.n112 10.6151
R751 B.n365 B.n112 10.6151
R752 B.n366 B.n365 10.6151
R753 B.n367 B.n366 10.6151
R754 B.n367 B.n110 10.6151
R755 B.n371 B.n110 10.6151
R756 B.n372 B.n371 10.6151
R757 B.n373 B.n372 10.6151
R758 B.n373 B.n108 10.6151
R759 B.n377 B.n108 10.6151
R760 B.n378 B.n377 10.6151
R761 B.n379 B.n378 10.6151
R762 B.n379 B.n106 10.6151
R763 B.n383 B.n106 10.6151
R764 B.n384 B.n383 10.6151
R765 B.n385 B.n384 10.6151
R766 B.n385 B.n104 10.6151
R767 B.n389 B.n104 10.6151
R768 B.n390 B.n389 10.6151
R769 B.n391 B.n390 10.6151
R770 B.n391 B.n102 10.6151
R771 B.n395 B.n102 10.6151
R772 B.n396 B.n395 10.6151
R773 B.n397 B.n396 10.6151
R774 B.n397 B.n100 10.6151
R775 B.n401 B.n100 10.6151
R776 B.n402 B.n401 10.6151
R777 B.n403 B.n402 10.6151
R778 B.n403 B.n98 10.6151
R779 B.n407 B.n98 10.6151
R780 B.n408 B.n407 10.6151
R781 B.n409 B.n408 10.6151
R782 B.n409 B.n96 10.6151
R783 B.n413 B.n96 10.6151
R784 B.n414 B.n413 10.6151
R785 B.n415 B.n414 10.6151
R786 B.n415 B.n94 10.6151
R787 B.n419 B.n94 10.6151
R788 B.n420 B.n419 10.6151
R789 B.n421 B.n420 10.6151
R790 B.n421 B.n92 10.6151
R791 B.n425 B.n92 10.6151
R792 B.n426 B.n425 10.6151
R793 B.n427 B.n426 10.6151
R794 B.n427 B.n90 10.6151
R795 B.n431 B.n90 10.6151
R796 B.n432 B.n431 10.6151
R797 B.n433 B.n432 10.6151
R798 B.n433 B.n88 10.6151
R799 B.n437 B.n88 10.6151
R800 B.n438 B.n437 10.6151
R801 B.n439 B.n438 10.6151
R802 B.n439 B.n86 10.6151
R803 B.n443 B.n86 10.6151
R804 B.n444 B.n443 10.6151
R805 B.n445 B.n444 10.6151
R806 B.n445 B.n84 10.6151
R807 B.n449 B.n84 10.6151
R808 B.n450 B.n449 10.6151
R809 B.n451 B.n450 10.6151
R810 B.n451 B.n82 10.6151
R811 B.n455 B.n82 10.6151
R812 B.n456 B.n455 10.6151
R813 B.n457 B.n456 10.6151
R814 B.n457 B.n80 10.6151
R815 B.n461 B.n80 10.6151
R816 B.n462 B.n461 10.6151
R817 B.n463 B.n462 10.6151
R818 B.n463 B.n78 10.6151
R819 B.n467 B.n78 10.6151
R820 B.n468 B.n467 10.6151
R821 B.n469 B.n468 10.6151
R822 B.n469 B.n76 10.6151
R823 B.n473 B.n76 10.6151
R824 B.n474 B.n473 10.6151
R825 B.n475 B.n474 10.6151
R826 B.n475 B.n74 10.6151
R827 B.n479 B.n74 10.6151
R828 B.n480 B.n479 10.6151
R829 B.n481 B.n480 10.6151
R830 B.n481 B.n72 10.6151
R831 B.n485 B.n72 10.6151
R832 B.n486 B.n485 10.6151
R833 B.n487 B.n486 10.6151
R834 B.n487 B.n70 10.6151
R835 B.n491 B.n70 10.6151
R836 B.n492 B.n491 10.6151
R837 B.n493 B.n492 10.6151
R838 B.n493 B.n68 10.6151
R839 B.n497 B.n68 10.6151
R840 B.n498 B.n497 10.6151
R841 B.n499 B.n498 10.6151
R842 B.n499 B.n66 10.6151
R843 B.n503 B.n66 10.6151
R844 B.n504 B.n503 10.6151
R845 B.n505 B.n504 10.6151
R846 B.n505 B.n64 10.6151
R847 B.n509 B.n64 10.6151
R848 B.n510 B.n509 10.6151
R849 B.n511 B.n510 10.6151
R850 B.n511 B.n62 10.6151
R851 B.n515 B.n62 10.6151
R852 B.n516 B.n515 10.6151
R853 B.n517 B.n516 10.6151
R854 B.n517 B.n60 10.6151
R855 B.n521 B.n60 10.6151
R856 B.n522 B.n521 10.6151
R857 B.n523 B.n522 10.6151
R858 B.n523 B.n58 10.6151
R859 B.n527 B.n58 10.6151
R860 B.n528 B.n527 10.6151
R861 B.n277 B.n276 10.6151
R862 B.n277 B.n144 10.6151
R863 B.n281 B.n144 10.6151
R864 B.n282 B.n281 10.6151
R865 B.n283 B.n282 10.6151
R866 B.n283 B.n142 10.6151
R867 B.n287 B.n142 10.6151
R868 B.n288 B.n287 10.6151
R869 B.n289 B.n288 10.6151
R870 B.n289 B.n140 10.6151
R871 B.n293 B.n140 10.6151
R872 B.n294 B.n293 10.6151
R873 B.n296 B.n136 10.6151
R874 B.n300 B.n136 10.6151
R875 B.n301 B.n300 10.6151
R876 B.n302 B.n301 10.6151
R877 B.n302 B.n134 10.6151
R878 B.n306 B.n134 10.6151
R879 B.n307 B.n306 10.6151
R880 B.n308 B.n307 10.6151
R881 B.n312 B.n311 10.6151
R882 B.n313 B.n312 10.6151
R883 B.n313 B.n128 10.6151
R884 B.n317 B.n128 10.6151
R885 B.n318 B.n317 10.6151
R886 B.n319 B.n318 10.6151
R887 B.n319 B.n126 10.6151
R888 B.n323 B.n126 10.6151
R889 B.n324 B.n323 10.6151
R890 B.n325 B.n324 10.6151
R891 B.n325 B.n124 10.6151
R892 B.n329 B.n124 10.6151
R893 B.n275 B.n146 10.6151
R894 B.n271 B.n146 10.6151
R895 B.n271 B.n270 10.6151
R896 B.n270 B.n269 10.6151
R897 B.n269 B.n148 10.6151
R898 B.n265 B.n148 10.6151
R899 B.n265 B.n264 10.6151
R900 B.n264 B.n263 10.6151
R901 B.n263 B.n150 10.6151
R902 B.n259 B.n150 10.6151
R903 B.n259 B.n258 10.6151
R904 B.n258 B.n257 10.6151
R905 B.n257 B.n152 10.6151
R906 B.n253 B.n152 10.6151
R907 B.n253 B.n252 10.6151
R908 B.n252 B.n251 10.6151
R909 B.n251 B.n154 10.6151
R910 B.n247 B.n154 10.6151
R911 B.n247 B.n246 10.6151
R912 B.n246 B.n245 10.6151
R913 B.n245 B.n156 10.6151
R914 B.n241 B.n156 10.6151
R915 B.n241 B.n240 10.6151
R916 B.n240 B.n239 10.6151
R917 B.n239 B.n158 10.6151
R918 B.n235 B.n158 10.6151
R919 B.n235 B.n234 10.6151
R920 B.n234 B.n233 10.6151
R921 B.n233 B.n160 10.6151
R922 B.n229 B.n160 10.6151
R923 B.n229 B.n228 10.6151
R924 B.n228 B.n227 10.6151
R925 B.n227 B.n162 10.6151
R926 B.n223 B.n162 10.6151
R927 B.n223 B.n222 10.6151
R928 B.n222 B.n221 10.6151
R929 B.n221 B.n164 10.6151
R930 B.n217 B.n164 10.6151
R931 B.n217 B.n216 10.6151
R932 B.n216 B.n215 10.6151
R933 B.n215 B.n166 10.6151
R934 B.n211 B.n166 10.6151
R935 B.n211 B.n210 10.6151
R936 B.n210 B.n209 10.6151
R937 B.n209 B.n168 10.6151
R938 B.n205 B.n168 10.6151
R939 B.n205 B.n204 10.6151
R940 B.n204 B.n203 10.6151
R941 B.n203 B.n170 10.6151
R942 B.n199 B.n170 10.6151
R943 B.n199 B.n198 10.6151
R944 B.n198 B.n197 10.6151
R945 B.n197 B.n172 10.6151
R946 B.n193 B.n172 10.6151
R947 B.n193 B.n192 10.6151
R948 B.n192 B.n191 10.6151
R949 B.n191 B.n174 10.6151
R950 B.n187 B.n174 10.6151
R951 B.n187 B.n186 10.6151
R952 B.n186 B.n185 10.6151
R953 B.n185 B.n176 10.6151
R954 B.n181 B.n176 10.6151
R955 B.n181 B.n180 10.6151
R956 B.n180 B.n179 10.6151
R957 B.n179 B.n0 10.6151
R958 B.n679 B.n1 10.6151
R959 B.n679 B.n678 10.6151
R960 B.n678 B.n677 10.6151
R961 B.n677 B.n4 10.6151
R962 B.n673 B.n4 10.6151
R963 B.n673 B.n672 10.6151
R964 B.n672 B.n671 10.6151
R965 B.n671 B.n6 10.6151
R966 B.n667 B.n6 10.6151
R967 B.n667 B.n666 10.6151
R968 B.n666 B.n665 10.6151
R969 B.n665 B.n8 10.6151
R970 B.n661 B.n8 10.6151
R971 B.n661 B.n660 10.6151
R972 B.n660 B.n659 10.6151
R973 B.n659 B.n10 10.6151
R974 B.n655 B.n10 10.6151
R975 B.n655 B.n654 10.6151
R976 B.n654 B.n653 10.6151
R977 B.n653 B.n12 10.6151
R978 B.n649 B.n12 10.6151
R979 B.n649 B.n648 10.6151
R980 B.n648 B.n647 10.6151
R981 B.n647 B.n14 10.6151
R982 B.n643 B.n14 10.6151
R983 B.n643 B.n642 10.6151
R984 B.n642 B.n641 10.6151
R985 B.n641 B.n16 10.6151
R986 B.n637 B.n16 10.6151
R987 B.n637 B.n636 10.6151
R988 B.n636 B.n635 10.6151
R989 B.n635 B.n18 10.6151
R990 B.n631 B.n18 10.6151
R991 B.n631 B.n630 10.6151
R992 B.n630 B.n629 10.6151
R993 B.n629 B.n20 10.6151
R994 B.n625 B.n20 10.6151
R995 B.n625 B.n624 10.6151
R996 B.n624 B.n623 10.6151
R997 B.n623 B.n22 10.6151
R998 B.n619 B.n22 10.6151
R999 B.n619 B.n618 10.6151
R1000 B.n618 B.n617 10.6151
R1001 B.n617 B.n24 10.6151
R1002 B.n613 B.n24 10.6151
R1003 B.n613 B.n612 10.6151
R1004 B.n612 B.n611 10.6151
R1005 B.n611 B.n26 10.6151
R1006 B.n607 B.n26 10.6151
R1007 B.n607 B.n606 10.6151
R1008 B.n606 B.n605 10.6151
R1009 B.n605 B.n28 10.6151
R1010 B.n601 B.n28 10.6151
R1011 B.n601 B.n600 10.6151
R1012 B.n600 B.n599 10.6151
R1013 B.n599 B.n30 10.6151
R1014 B.n595 B.n30 10.6151
R1015 B.n595 B.n594 10.6151
R1016 B.n594 B.n593 10.6151
R1017 B.n593 B.n32 10.6151
R1018 B.n589 B.n32 10.6151
R1019 B.n589 B.n588 10.6151
R1020 B.n588 B.n587 10.6151
R1021 B.n587 B.n34 10.6151
R1022 B.n583 B.n34 10.6151
R1023 B.n563 B.n562 6.5566
R1024 B.n550 B.n50 6.5566
R1025 B.n296 B.n295 6.5566
R1026 B.n308 B.n132 6.5566
R1027 B.n564 B.n563 4.05904
R1028 B.n547 B.n50 4.05904
R1029 B.n295 B.n294 4.05904
R1030 B.n311 B.n132 4.05904
R1031 B.n683 B.n0 2.81026
R1032 B.n683 B.n1 2.81026
R1033 VN.n72 VN.n71 161.3
R1034 VN.n70 VN.n38 161.3
R1035 VN.n69 VN.n68 161.3
R1036 VN.n67 VN.n39 161.3
R1037 VN.n66 VN.n65 161.3
R1038 VN.n64 VN.n40 161.3
R1039 VN.n63 VN.n62 161.3
R1040 VN.n61 VN.n41 161.3
R1041 VN.n60 VN.n59 161.3
R1042 VN.n58 VN.n42 161.3
R1043 VN.n57 VN.n56 161.3
R1044 VN.n55 VN.n44 161.3
R1045 VN.n54 VN.n53 161.3
R1046 VN.n52 VN.n45 161.3
R1047 VN.n51 VN.n50 161.3
R1048 VN.n49 VN.n46 161.3
R1049 VN.n35 VN.n34 161.3
R1050 VN.n33 VN.n1 161.3
R1051 VN.n32 VN.n31 161.3
R1052 VN.n30 VN.n2 161.3
R1053 VN.n29 VN.n28 161.3
R1054 VN.n27 VN.n3 161.3
R1055 VN.n26 VN.n25 161.3
R1056 VN.n24 VN.n4 161.3
R1057 VN.n23 VN.n22 161.3
R1058 VN.n20 VN.n5 161.3
R1059 VN.n19 VN.n18 161.3
R1060 VN.n17 VN.n6 161.3
R1061 VN.n16 VN.n15 161.3
R1062 VN.n14 VN.n7 161.3
R1063 VN.n13 VN.n12 161.3
R1064 VN.n11 VN.n8 161.3
R1065 VN.n36 VN.n0 81.6384
R1066 VN.n73 VN.n37 81.6384
R1067 VN.n10 VN.n9 63.7241
R1068 VN.n48 VN.n47 63.7241
R1069 VN.n15 VN.n6 56.5617
R1070 VN.n28 VN.n2 56.5617
R1071 VN.n53 VN.n44 56.5617
R1072 VN.n65 VN.n39 56.5617
R1073 VN VN.n73 48.4451
R1074 VN.n48 VN.t4 47.3529
R1075 VN.n10 VN.t3 47.3529
R1076 VN.n13 VN.n8 24.5923
R1077 VN.n14 VN.n13 24.5923
R1078 VN.n15 VN.n14 24.5923
R1079 VN.n19 VN.n6 24.5923
R1080 VN.n20 VN.n19 24.5923
R1081 VN.n22 VN.n20 24.5923
R1082 VN.n26 VN.n4 24.5923
R1083 VN.n27 VN.n26 24.5923
R1084 VN.n28 VN.n27 24.5923
R1085 VN.n32 VN.n2 24.5923
R1086 VN.n33 VN.n32 24.5923
R1087 VN.n34 VN.n33 24.5923
R1088 VN.n53 VN.n52 24.5923
R1089 VN.n52 VN.n51 24.5923
R1090 VN.n51 VN.n46 24.5923
R1091 VN.n65 VN.n64 24.5923
R1092 VN.n64 VN.n63 24.5923
R1093 VN.n63 VN.n41 24.5923
R1094 VN.n59 VN.n58 24.5923
R1095 VN.n58 VN.n57 24.5923
R1096 VN.n57 VN.n44 24.5923
R1097 VN.n71 VN.n70 24.5923
R1098 VN.n70 VN.n69 24.5923
R1099 VN.n69 VN.n39 24.5923
R1100 VN.n9 VN.t6 14.1143
R1101 VN.n21 VN.t5 14.1143
R1102 VN.n0 VN.t0 14.1143
R1103 VN.n47 VN.t2 14.1143
R1104 VN.n43 VN.t1 14.1143
R1105 VN.n37 VN.t7 14.1143
R1106 VN.n21 VN.n4 13.526
R1107 VN.n43 VN.n41 13.526
R1108 VN.n9 VN.n8 11.0668
R1109 VN.n22 VN.n21 11.0668
R1110 VN.n47 VN.n46 11.0668
R1111 VN.n59 VN.n43 11.0668
R1112 VN.n34 VN.n0 8.60764
R1113 VN.n71 VN.n37 8.60764
R1114 VN.n49 VN.n48 3.19096
R1115 VN.n11 VN.n10 3.19096
R1116 VN.n73 VN.n72 0.354861
R1117 VN.n36 VN.n35 0.354861
R1118 VN VN.n36 0.267071
R1119 VN.n72 VN.n38 0.189894
R1120 VN.n68 VN.n38 0.189894
R1121 VN.n68 VN.n67 0.189894
R1122 VN.n67 VN.n66 0.189894
R1123 VN.n66 VN.n40 0.189894
R1124 VN.n62 VN.n40 0.189894
R1125 VN.n62 VN.n61 0.189894
R1126 VN.n61 VN.n60 0.189894
R1127 VN.n60 VN.n42 0.189894
R1128 VN.n56 VN.n42 0.189894
R1129 VN.n56 VN.n55 0.189894
R1130 VN.n55 VN.n54 0.189894
R1131 VN.n54 VN.n45 0.189894
R1132 VN.n50 VN.n45 0.189894
R1133 VN.n50 VN.n49 0.189894
R1134 VN.n12 VN.n11 0.189894
R1135 VN.n12 VN.n7 0.189894
R1136 VN.n16 VN.n7 0.189894
R1137 VN.n17 VN.n16 0.189894
R1138 VN.n18 VN.n17 0.189894
R1139 VN.n18 VN.n5 0.189894
R1140 VN.n23 VN.n5 0.189894
R1141 VN.n24 VN.n23 0.189894
R1142 VN.n25 VN.n24 0.189894
R1143 VN.n25 VN.n3 0.189894
R1144 VN.n29 VN.n3 0.189894
R1145 VN.n30 VN.n29 0.189894
R1146 VN.n31 VN.n30 0.189894
R1147 VN.n31 VN.n1 0.189894
R1148 VN.n35 VN.n1 0.189894
R1149 VTAIL.n15 VTAIL.t6 171.044
R1150 VTAIL.n2 VTAIL.t5 171.044
R1151 VTAIL.n3 VTAIL.t9 171.044
R1152 VTAIL.n6 VTAIL.t12 171.044
R1153 VTAIL.n14 VTAIL.t8 171.044
R1154 VTAIL.n11 VTAIL.t11 171.044
R1155 VTAIL.n10 VTAIL.t4 171.044
R1156 VTAIL.n7 VTAIL.t7 171.044
R1157 VTAIL.n13 VTAIL.n12 155.713
R1158 VTAIL.n9 VTAIL.n8 155.713
R1159 VTAIL.n1 VTAIL.n0 155.712
R1160 VTAIL.n5 VTAIL.n4 155.712
R1161 VTAIL.n15 VTAIL.n14 17.5996
R1162 VTAIL.n7 VTAIL.n6 17.5996
R1163 VTAIL.n0 VTAIL.t0 15.333
R1164 VTAIL.n0 VTAIL.t3 15.333
R1165 VTAIL.n4 VTAIL.t14 15.333
R1166 VTAIL.n4 VTAIL.t15 15.333
R1167 VTAIL.n12 VTAIL.t13 15.333
R1168 VTAIL.n12 VTAIL.t10 15.333
R1169 VTAIL.n8 VTAIL.t1 15.333
R1170 VTAIL.n8 VTAIL.t2 15.333
R1171 VTAIL.n9 VTAIL.n7 3.40567
R1172 VTAIL.n10 VTAIL.n9 3.40567
R1173 VTAIL.n13 VTAIL.n11 3.40567
R1174 VTAIL.n14 VTAIL.n13 3.40567
R1175 VTAIL.n6 VTAIL.n5 3.40567
R1176 VTAIL.n5 VTAIL.n3 3.40567
R1177 VTAIL.n2 VTAIL.n1 3.40567
R1178 VTAIL VTAIL.n15 3.34748
R1179 VTAIL.n11 VTAIL.n10 0.470328
R1180 VTAIL.n3 VTAIL.n2 0.470328
R1181 VTAIL VTAIL.n1 0.0586897
R1182 VDD2.n2 VDD2.n1 174.037
R1183 VDD2.n2 VDD2.n0 174.037
R1184 VDD2 VDD2.n5 174.036
R1185 VDD2.n4 VDD2.n3 172.391
R1186 VDD2.n4 VDD2.n2 40.8662
R1187 VDD2.n5 VDD2.t5 15.333
R1188 VDD2.n5 VDD2.t3 15.333
R1189 VDD2.n3 VDD2.t0 15.333
R1190 VDD2.n3 VDD2.t6 15.333
R1191 VDD2.n1 VDD2.t2 15.333
R1192 VDD2.n1 VDD2.t7 15.333
R1193 VDD2.n0 VDD2.t4 15.333
R1194 VDD2.n0 VDD2.t1 15.333
R1195 VDD2 VDD2.n4 1.76128
R1196 VP.n24 VP.n21 161.3
R1197 VP.n26 VP.n25 161.3
R1198 VP.n27 VP.n20 161.3
R1199 VP.n29 VP.n28 161.3
R1200 VP.n30 VP.n19 161.3
R1201 VP.n32 VP.n31 161.3
R1202 VP.n33 VP.n18 161.3
R1203 VP.n36 VP.n35 161.3
R1204 VP.n37 VP.n17 161.3
R1205 VP.n39 VP.n38 161.3
R1206 VP.n40 VP.n16 161.3
R1207 VP.n42 VP.n41 161.3
R1208 VP.n43 VP.n15 161.3
R1209 VP.n45 VP.n44 161.3
R1210 VP.n46 VP.n14 161.3
R1211 VP.n48 VP.n47 161.3
R1212 VP.n89 VP.n88 161.3
R1213 VP.n87 VP.n1 161.3
R1214 VP.n86 VP.n85 161.3
R1215 VP.n84 VP.n2 161.3
R1216 VP.n83 VP.n82 161.3
R1217 VP.n81 VP.n3 161.3
R1218 VP.n80 VP.n79 161.3
R1219 VP.n78 VP.n4 161.3
R1220 VP.n77 VP.n76 161.3
R1221 VP.n74 VP.n5 161.3
R1222 VP.n73 VP.n72 161.3
R1223 VP.n71 VP.n6 161.3
R1224 VP.n70 VP.n69 161.3
R1225 VP.n68 VP.n7 161.3
R1226 VP.n67 VP.n66 161.3
R1227 VP.n65 VP.n8 161.3
R1228 VP.n64 VP.n63 161.3
R1229 VP.n61 VP.n9 161.3
R1230 VP.n60 VP.n59 161.3
R1231 VP.n58 VP.n10 161.3
R1232 VP.n57 VP.n56 161.3
R1233 VP.n55 VP.n11 161.3
R1234 VP.n54 VP.n53 161.3
R1235 VP.n52 VP.n12 161.3
R1236 VP.n51 VP.n50 81.6384
R1237 VP.n90 VP.n0 81.6384
R1238 VP.n49 VP.n13 81.6384
R1239 VP.n23 VP.n22 63.7241
R1240 VP.n56 VP.n10 56.5617
R1241 VP.n69 VP.n6 56.5617
R1242 VP.n82 VP.n2 56.5617
R1243 VP.n41 VP.n15 56.5617
R1244 VP.n28 VP.n19 56.5617
R1245 VP.n51 VP.n49 48.2799
R1246 VP.n23 VP.t2 47.3528
R1247 VP.n54 VP.n12 24.5923
R1248 VP.n55 VP.n54 24.5923
R1249 VP.n56 VP.n55 24.5923
R1250 VP.n60 VP.n10 24.5923
R1251 VP.n61 VP.n60 24.5923
R1252 VP.n63 VP.n61 24.5923
R1253 VP.n67 VP.n8 24.5923
R1254 VP.n68 VP.n67 24.5923
R1255 VP.n69 VP.n68 24.5923
R1256 VP.n73 VP.n6 24.5923
R1257 VP.n74 VP.n73 24.5923
R1258 VP.n76 VP.n74 24.5923
R1259 VP.n80 VP.n4 24.5923
R1260 VP.n81 VP.n80 24.5923
R1261 VP.n82 VP.n81 24.5923
R1262 VP.n86 VP.n2 24.5923
R1263 VP.n87 VP.n86 24.5923
R1264 VP.n88 VP.n87 24.5923
R1265 VP.n45 VP.n15 24.5923
R1266 VP.n46 VP.n45 24.5923
R1267 VP.n47 VP.n46 24.5923
R1268 VP.n32 VP.n19 24.5923
R1269 VP.n33 VP.n32 24.5923
R1270 VP.n35 VP.n33 24.5923
R1271 VP.n39 VP.n17 24.5923
R1272 VP.n40 VP.n39 24.5923
R1273 VP.n41 VP.n40 24.5923
R1274 VP.n26 VP.n21 24.5923
R1275 VP.n27 VP.n26 24.5923
R1276 VP.n28 VP.n27 24.5923
R1277 VP.n50 VP.t7 14.1143
R1278 VP.n62 VP.t0 14.1143
R1279 VP.n75 VP.t6 14.1143
R1280 VP.n0 VP.t4 14.1143
R1281 VP.n13 VP.t3 14.1143
R1282 VP.n34 VP.t5 14.1143
R1283 VP.n22 VP.t1 14.1143
R1284 VP.n63 VP.n62 13.526
R1285 VP.n75 VP.n4 13.526
R1286 VP.n34 VP.n17 13.526
R1287 VP.n62 VP.n8 11.0668
R1288 VP.n76 VP.n75 11.0668
R1289 VP.n35 VP.n34 11.0668
R1290 VP.n22 VP.n21 11.0668
R1291 VP.n50 VP.n12 8.60764
R1292 VP.n88 VP.n0 8.60764
R1293 VP.n47 VP.n13 8.60764
R1294 VP.n24 VP.n23 3.19095
R1295 VP.n49 VP.n48 0.354861
R1296 VP.n52 VP.n51 0.354861
R1297 VP.n90 VP.n89 0.354861
R1298 VP VP.n90 0.267071
R1299 VP.n25 VP.n24 0.189894
R1300 VP.n25 VP.n20 0.189894
R1301 VP.n29 VP.n20 0.189894
R1302 VP.n30 VP.n29 0.189894
R1303 VP.n31 VP.n30 0.189894
R1304 VP.n31 VP.n18 0.189894
R1305 VP.n36 VP.n18 0.189894
R1306 VP.n37 VP.n36 0.189894
R1307 VP.n38 VP.n37 0.189894
R1308 VP.n38 VP.n16 0.189894
R1309 VP.n42 VP.n16 0.189894
R1310 VP.n43 VP.n42 0.189894
R1311 VP.n44 VP.n43 0.189894
R1312 VP.n44 VP.n14 0.189894
R1313 VP.n48 VP.n14 0.189894
R1314 VP.n53 VP.n52 0.189894
R1315 VP.n53 VP.n11 0.189894
R1316 VP.n57 VP.n11 0.189894
R1317 VP.n58 VP.n57 0.189894
R1318 VP.n59 VP.n58 0.189894
R1319 VP.n59 VP.n9 0.189894
R1320 VP.n64 VP.n9 0.189894
R1321 VP.n65 VP.n64 0.189894
R1322 VP.n66 VP.n65 0.189894
R1323 VP.n66 VP.n7 0.189894
R1324 VP.n70 VP.n7 0.189894
R1325 VP.n71 VP.n70 0.189894
R1326 VP.n72 VP.n71 0.189894
R1327 VP.n72 VP.n5 0.189894
R1328 VP.n77 VP.n5 0.189894
R1329 VP.n78 VP.n77 0.189894
R1330 VP.n79 VP.n78 0.189894
R1331 VP.n79 VP.n3 0.189894
R1332 VP.n83 VP.n3 0.189894
R1333 VP.n84 VP.n83 0.189894
R1334 VP.n85 VP.n84 0.189894
R1335 VP.n85 VP.n1 0.189894
R1336 VP.n89 VP.n1 0.189894
R1337 VDD1 VDD1.n0 174.151
R1338 VDD1.n3 VDD1.n2 174.037
R1339 VDD1.n3 VDD1.n1 174.037
R1340 VDD1.n5 VDD1.n4 172.391
R1341 VDD1.n5 VDD1.n3 41.4492
R1342 VDD1.n4 VDD1.t2 15.333
R1343 VDD1.n4 VDD1.t4 15.333
R1344 VDD1.n0 VDD1.t5 15.333
R1345 VDD1.n0 VDD1.t6 15.333
R1346 VDD1.n2 VDD1.t1 15.333
R1347 VDD1.n2 VDD1.t3 15.333
R1348 VDD1.n1 VDD1.t0 15.333
R1349 VDD1.n1 VDD1.t7 15.333
R1350 VDD1 VDD1.n5 1.6449
C0 VTAIL VDD2 5.75303f
C1 VDD1 VN 0.159754f
C2 VDD1 VP 2.48939f
C3 VN VTAIL 3.5893f
C4 VP VTAIL 3.6034f
C5 w_n4920_n1392# B 8.97971f
C6 VDD1 w_n4920_n1392# 2.01518f
C7 VDD1 B 1.69406f
C8 VTAIL w_n4920_n1392# 2.10526f
C9 VN VDD2 2.01705f
C10 VP VDD2 0.635754f
C11 VTAIL B 1.88059f
C12 VDD1 VTAIL 5.69177f
C13 VP VN 7.08054f
C14 w_n4920_n1392# VDD2 2.17197f
C15 VDD2 B 1.82261f
C16 VDD1 VDD2 2.30735f
C17 VN w_n4920_n1392# 10.1268f
C18 VP w_n4920_n1392# 10.764299f
C19 VN B 1.35695f
C20 VP B 2.43743f
C21 VDD2 VSUBS 2.155366f
C22 VDD1 VSUBS 2.98664f
C23 VTAIL VSUBS 0.695596f
C24 VN VSUBS 8.36443f
C25 VP VSUBS 3.964023f
C26 B VSUBS 4.971448f
C27 w_n4920_n1392# VSUBS 87.320206f
C28 VDD1.t5 VSUBS 0.063991f
C29 VDD1.t6 VSUBS 0.063991f
C30 VDD1.n0 VSUBS 0.30296f
C31 VDD1.t0 VSUBS 0.063991f
C32 VDD1.t7 VSUBS 0.063991f
C33 VDD1.n1 VSUBS 0.302145f
C34 VDD1.t1 VSUBS 0.063991f
C35 VDD1.t3 VSUBS 0.063991f
C36 VDD1.n2 VSUBS 0.302145f
C37 VDD1.n3 VSUBS 5.28405f
C38 VDD1.t2 VSUBS 0.063991f
C39 VDD1.t4 VSUBS 0.063991f
C40 VDD1.n4 VSUBS 0.29219f
C41 VDD1.n5 VSUBS 4.03114f
C42 VP.t4 VSUBS 1.01105f
C43 VP.n0 VSUBS 0.666758f
C44 VP.n1 VSUBS 0.05578f
C45 VP.n2 VSUBS 0.088802f
C46 VP.n3 VSUBS 0.05578f
C47 VP.n4 VSUBS 0.08046f
C48 VP.n5 VSUBS 0.05578f
C49 VP.n6 VSUBS 0.081085f
C50 VP.n7 VSUBS 0.05578f
C51 VP.n8 VSUBS 0.075354f
C52 VP.n9 VSUBS 0.05578f
C53 VP.n10 VSUBS 0.073369f
C54 VP.n11 VSUBS 0.05578f
C55 VP.n12 VSUBS 0.070247f
C56 VP.t3 VSUBS 1.01105f
C57 VP.n13 VSUBS 0.666758f
C58 VP.n14 VSUBS 0.05578f
C59 VP.n15 VSUBS 0.088802f
C60 VP.n16 VSUBS 0.05578f
C61 VP.n17 VSUBS 0.08046f
C62 VP.n18 VSUBS 0.05578f
C63 VP.n19 VSUBS 0.081085f
C64 VP.n20 VSUBS 0.05578f
C65 VP.n21 VSUBS 0.075354f
C66 VP.t2 VSUBS 1.6238f
C67 VP.t1 VSUBS 1.01105f
C68 VP.n22 VSUBS 0.64129f
C69 VP.n23 VSUBS 0.702309f
C70 VP.n24 VSUBS 0.69818f
C71 VP.n25 VSUBS 0.05578f
C72 VP.n26 VSUBS 0.103439f
C73 VP.n27 VSUBS 0.103439f
C74 VP.n28 VSUBS 0.081085f
C75 VP.n29 VSUBS 0.05578f
C76 VP.n30 VSUBS 0.05578f
C77 VP.n31 VSUBS 0.05578f
C78 VP.n32 VSUBS 0.103439f
C79 VP.n33 VSUBS 0.103439f
C80 VP.t5 VSUBS 1.01105f
C81 VP.n34 VSUBS 0.45096f
C82 VP.n35 VSUBS 0.075354f
C83 VP.n36 VSUBS 0.05578f
C84 VP.n37 VSUBS 0.05578f
C85 VP.n38 VSUBS 0.05578f
C86 VP.n39 VSUBS 0.103439f
C87 VP.n40 VSUBS 0.103439f
C88 VP.n41 VSUBS 0.073369f
C89 VP.n42 VSUBS 0.05578f
C90 VP.n43 VSUBS 0.05578f
C91 VP.n44 VSUBS 0.05578f
C92 VP.n45 VSUBS 0.103439f
C93 VP.n46 VSUBS 0.103439f
C94 VP.n47 VSUBS 0.070247f
C95 VP.n48 VSUBS 0.090014f
C96 VP.n49 VSUBS 3.0385f
C97 VP.t7 VSUBS 1.01105f
C98 VP.n50 VSUBS 0.666758f
C99 VP.n51 VSUBS 3.08015f
C100 VP.n52 VSUBS 0.090014f
C101 VP.n53 VSUBS 0.05578f
C102 VP.n54 VSUBS 0.103439f
C103 VP.n55 VSUBS 0.103439f
C104 VP.n56 VSUBS 0.088802f
C105 VP.n57 VSUBS 0.05578f
C106 VP.n58 VSUBS 0.05578f
C107 VP.n59 VSUBS 0.05578f
C108 VP.n60 VSUBS 0.103439f
C109 VP.n61 VSUBS 0.103439f
C110 VP.t0 VSUBS 1.01105f
C111 VP.n62 VSUBS 0.45096f
C112 VP.n63 VSUBS 0.08046f
C113 VP.n64 VSUBS 0.05578f
C114 VP.n65 VSUBS 0.05578f
C115 VP.n66 VSUBS 0.05578f
C116 VP.n67 VSUBS 0.103439f
C117 VP.n68 VSUBS 0.103439f
C118 VP.n69 VSUBS 0.081085f
C119 VP.n70 VSUBS 0.05578f
C120 VP.n71 VSUBS 0.05578f
C121 VP.n72 VSUBS 0.05578f
C122 VP.n73 VSUBS 0.103439f
C123 VP.n74 VSUBS 0.103439f
C124 VP.t6 VSUBS 1.01105f
C125 VP.n75 VSUBS 0.45096f
C126 VP.n76 VSUBS 0.075354f
C127 VP.n77 VSUBS 0.05578f
C128 VP.n78 VSUBS 0.05578f
C129 VP.n79 VSUBS 0.05578f
C130 VP.n80 VSUBS 0.103439f
C131 VP.n81 VSUBS 0.103439f
C132 VP.n82 VSUBS 0.073369f
C133 VP.n83 VSUBS 0.05578f
C134 VP.n84 VSUBS 0.05578f
C135 VP.n85 VSUBS 0.05578f
C136 VP.n86 VSUBS 0.103439f
C137 VP.n87 VSUBS 0.103439f
C138 VP.n88 VSUBS 0.070247f
C139 VP.n89 VSUBS 0.090014f
C140 VP.n90 VSUBS 0.155686f
C141 VDD2.t4 VSUBS 0.063686f
C142 VDD2.t1 VSUBS 0.063686f
C143 VDD2.n0 VSUBS 0.300704f
C144 VDD2.t2 VSUBS 0.063686f
C145 VDD2.t7 VSUBS 0.063686f
C146 VDD2.n1 VSUBS 0.300704f
C147 VDD2.n2 VSUBS 5.180181f
C148 VDD2.t0 VSUBS 0.063686f
C149 VDD2.t6 VSUBS 0.063686f
C150 VDD2.n3 VSUBS 0.290799f
C151 VDD2.n4 VSUBS 3.96445f
C152 VDD2.t5 VSUBS 0.063686f
C153 VDD2.t3 VSUBS 0.063686f
C154 VDD2.n5 VSUBS 0.300679f
C155 VTAIL.t0 VSUBS 0.062352f
C156 VTAIL.t3 VSUBS 0.062352f
C157 VTAIL.n0 VSUBS 0.242268f
C158 VTAIL.n1 VSUBS 0.810493f
C159 VTAIL.t5 VSUBS 0.380948f
C160 VTAIL.n2 VSUBS 0.891231f
C161 VTAIL.t9 VSUBS 0.380948f
C162 VTAIL.n3 VSUBS 0.891231f
C163 VTAIL.t14 VSUBS 0.062352f
C164 VTAIL.t15 VSUBS 0.062352f
C165 VTAIL.n4 VSUBS 0.242268f
C166 VTAIL.n5 VSUBS 1.21189f
C167 VTAIL.t12 VSUBS 0.380948f
C168 VTAIL.n6 VSUBS 1.96801f
C169 VTAIL.t7 VSUBS 0.38095f
C170 VTAIL.n7 VSUBS 1.96801f
C171 VTAIL.t1 VSUBS 0.062352f
C172 VTAIL.t2 VSUBS 0.062352f
C173 VTAIL.n8 VSUBS 0.242269f
C174 VTAIL.n9 VSUBS 1.21189f
C175 VTAIL.t4 VSUBS 0.38095f
C176 VTAIL.n10 VSUBS 0.89123f
C177 VTAIL.t11 VSUBS 0.38095f
C178 VTAIL.n11 VSUBS 0.89123f
C179 VTAIL.t13 VSUBS 0.062352f
C180 VTAIL.t10 VSUBS 0.062352f
C181 VTAIL.n12 VSUBS 0.242269f
C182 VTAIL.n13 VSUBS 1.21189f
C183 VTAIL.t8 VSUBS 0.380948f
C184 VTAIL.n14 VSUBS 1.96801f
C185 VTAIL.t6 VSUBS 0.380948f
C186 VTAIL.n15 VSUBS 1.96103f
C187 VN.t0 VSUBS 0.870597f
C188 VN.n0 VSUBS 0.574132f
C189 VN.n1 VSUBS 0.048031f
C190 VN.n2 VSUBS 0.076465f
C191 VN.n3 VSUBS 0.048031f
C192 VN.n4 VSUBS 0.069283f
C193 VN.n5 VSUBS 0.048031f
C194 VN.n6 VSUBS 0.069821f
C195 VN.n7 VSUBS 0.048031f
C196 VN.n8 VSUBS 0.064885f
C197 VN.t6 VSUBS 0.870597f
C198 VN.n9 VSUBS 0.552201f
C199 VN.t3 VSUBS 1.39823f
C200 VN.n10 VSUBS 0.604743f
C201 VN.n11 VSUBS 0.601187f
C202 VN.n12 VSUBS 0.048031f
C203 VN.n13 VSUBS 0.08907f
C204 VN.n14 VSUBS 0.08907f
C205 VN.n15 VSUBS 0.069821f
C206 VN.n16 VSUBS 0.048031f
C207 VN.n17 VSUBS 0.048031f
C208 VN.n18 VSUBS 0.048031f
C209 VN.n19 VSUBS 0.08907f
C210 VN.n20 VSUBS 0.08907f
C211 VN.t5 VSUBS 0.870597f
C212 VN.n21 VSUBS 0.388312f
C213 VN.n22 VSUBS 0.064885f
C214 VN.n23 VSUBS 0.048031f
C215 VN.n24 VSUBS 0.048031f
C216 VN.n25 VSUBS 0.048031f
C217 VN.n26 VSUBS 0.08907f
C218 VN.n27 VSUBS 0.08907f
C219 VN.n28 VSUBS 0.063176f
C220 VN.n29 VSUBS 0.048031f
C221 VN.n30 VSUBS 0.048031f
C222 VN.n31 VSUBS 0.048031f
C223 VN.n32 VSUBS 0.08907f
C224 VN.n33 VSUBS 0.08907f
C225 VN.n34 VSUBS 0.060488f
C226 VN.n35 VSUBS 0.077509f
C227 VN.n36 VSUBS 0.134058f
C228 VN.t7 VSUBS 0.870597f
C229 VN.n37 VSUBS 0.574132f
C230 VN.n38 VSUBS 0.048031f
C231 VN.n39 VSUBS 0.076465f
C232 VN.n40 VSUBS 0.048031f
C233 VN.n41 VSUBS 0.069283f
C234 VN.n42 VSUBS 0.048031f
C235 VN.t1 VSUBS 0.870597f
C236 VN.n43 VSUBS 0.388312f
C237 VN.n44 VSUBS 0.069821f
C238 VN.n45 VSUBS 0.048031f
C239 VN.n46 VSUBS 0.064885f
C240 VN.t4 VSUBS 1.39823f
C241 VN.t2 VSUBS 0.870597f
C242 VN.n47 VSUBS 0.552201f
C243 VN.n48 VSUBS 0.604743f
C244 VN.n49 VSUBS 0.601187f
C245 VN.n50 VSUBS 0.048031f
C246 VN.n51 VSUBS 0.08907f
C247 VN.n52 VSUBS 0.08907f
C248 VN.n53 VSUBS 0.069821f
C249 VN.n54 VSUBS 0.048031f
C250 VN.n55 VSUBS 0.048031f
C251 VN.n56 VSUBS 0.048031f
C252 VN.n57 VSUBS 0.08907f
C253 VN.n58 VSUBS 0.08907f
C254 VN.n59 VSUBS 0.064885f
C255 VN.n60 VSUBS 0.048031f
C256 VN.n61 VSUBS 0.048031f
C257 VN.n62 VSUBS 0.048031f
C258 VN.n63 VSUBS 0.08907f
C259 VN.n64 VSUBS 0.08907f
C260 VN.n65 VSUBS 0.063176f
C261 VN.n66 VSUBS 0.048031f
C262 VN.n67 VSUBS 0.048031f
C263 VN.n68 VSUBS 0.048031f
C264 VN.n69 VSUBS 0.08907f
C265 VN.n70 VSUBS 0.08907f
C266 VN.n71 VSUBS 0.060488f
C267 VN.n72 VSUBS 0.077509f
C268 VN.n73 VSUBS 2.63627f
C269 B.n0 VSUBS 0.006771f
C270 B.n1 VSUBS 0.006771f
C271 B.n2 VSUBS 0.010708f
C272 B.n3 VSUBS 0.010708f
C273 B.n4 VSUBS 0.010708f
C274 B.n5 VSUBS 0.010708f
C275 B.n6 VSUBS 0.010708f
C276 B.n7 VSUBS 0.010708f
C277 B.n8 VSUBS 0.010708f
C278 B.n9 VSUBS 0.010708f
C279 B.n10 VSUBS 0.010708f
C280 B.n11 VSUBS 0.010708f
C281 B.n12 VSUBS 0.010708f
C282 B.n13 VSUBS 0.010708f
C283 B.n14 VSUBS 0.010708f
C284 B.n15 VSUBS 0.010708f
C285 B.n16 VSUBS 0.010708f
C286 B.n17 VSUBS 0.010708f
C287 B.n18 VSUBS 0.010708f
C288 B.n19 VSUBS 0.010708f
C289 B.n20 VSUBS 0.010708f
C290 B.n21 VSUBS 0.010708f
C291 B.n22 VSUBS 0.010708f
C292 B.n23 VSUBS 0.010708f
C293 B.n24 VSUBS 0.010708f
C294 B.n25 VSUBS 0.010708f
C295 B.n26 VSUBS 0.010708f
C296 B.n27 VSUBS 0.010708f
C297 B.n28 VSUBS 0.010708f
C298 B.n29 VSUBS 0.010708f
C299 B.n30 VSUBS 0.010708f
C300 B.n31 VSUBS 0.010708f
C301 B.n32 VSUBS 0.010708f
C302 B.n33 VSUBS 0.010708f
C303 B.n34 VSUBS 0.010708f
C304 B.n35 VSUBS 0.02616f
C305 B.n36 VSUBS 0.010708f
C306 B.n37 VSUBS 0.010708f
C307 B.n38 VSUBS 0.010708f
C308 B.n39 VSUBS 0.010708f
C309 B.n40 VSUBS 0.010708f
C310 B.n41 VSUBS 0.010708f
C311 B.t2 VSUBS 0.071007f
C312 B.t1 VSUBS 0.096227f
C313 B.t0 VSUBS 0.580232f
C314 B.n42 VSUBS 0.124291f
C315 B.n43 VSUBS 0.09707f
C316 B.n44 VSUBS 0.010708f
C317 B.n45 VSUBS 0.010708f
C318 B.n46 VSUBS 0.010708f
C319 B.n47 VSUBS 0.010708f
C320 B.t5 VSUBS 0.071007f
C321 B.t4 VSUBS 0.096227f
C322 B.t3 VSUBS 0.580232f
C323 B.n48 VSUBS 0.124291f
C324 B.n49 VSUBS 0.09707f
C325 B.n50 VSUBS 0.02481f
C326 B.n51 VSUBS 0.010708f
C327 B.n52 VSUBS 0.010708f
C328 B.n53 VSUBS 0.010708f
C329 B.n54 VSUBS 0.010708f
C330 B.n55 VSUBS 0.010708f
C331 B.n56 VSUBS 0.010708f
C332 B.n57 VSUBS 0.024232f
C333 B.n58 VSUBS 0.010708f
C334 B.n59 VSUBS 0.010708f
C335 B.n60 VSUBS 0.010708f
C336 B.n61 VSUBS 0.010708f
C337 B.n62 VSUBS 0.010708f
C338 B.n63 VSUBS 0.010708f
C339 B.n64 VSUBS 0.010708f
C340 B.n65 VSUBS 0.010708f
C341 B.n66 VSUBS 0.010708f
C342 B.n67 VSUBS 0.010708f
C343 B.n68 VSUBS 0.010708f
C344 B.n69 VSUBS 0.010708f
C345 B.n70 VSUBS 0.010708f
C346 B.n71 VSUBS 0.010708f
C347 B.n72 VSUBS 0.010708f
C348 B.n73 VSUBS 0.010708f
C349 B.n74 VSUBS 0.010708f
C350 B.n75 VSUBS 0.010708f
C351 B.n76 VSUBS 0.010708f
C352 B.n77 VSUBS 0.010708f
C353 B.n78 VSUBS 0.010708f
C354 B.n79 VSUBS 0.010708f
C355 B.n80 VSUBS 0.010708f
C356 B.n81 VSUBS 0.010708f
C357 B.n82 VSUBS 0.010708f
C358 B.n83 VSUBS 0.010708f
C359 B.n84 VSUBS 0.010708f
C360 B.n85 VSUBS 0.010708f
C361 B.n86 VSUBS 0.010708f
C362 B.n87 VSUBS 0.010708f
C363 B.n88 VSUBS 0.010708f
C364 B.n89 VSUBS 0.010708f
C365 B.n90 VSUBS 0.010708f
C366 B.n91 VSUBS 0.010708f
C367 B.n92 VSUBS 0.010708f
C368 B.n93 VSUBS 0.010708f
C369 B.n94 VSUBS 0.010708f
C370 B.n95 VSUBS 0.010708f
C371 B.n96 VSUBS 0.010708f
C372 B.n97 VSUBS 0.010708f
C373 B.n98 VSUBS 0.010708f
C374 B.n99 VSUBS 0.010708f
C375 B.n100 VSUBS 0.010708f
C376 B.n101 VSUBS 0.010708f
C377 B.n102 VSUBS 0.010708f
C378 B.n103 VSUBS 0.010708f
C379 B.n104 VSUBS 0.010708f
C380 B.n105 VSUBS 0.010708f
C381 B.n106 VSUBS 0.010708f
C382 B.n107 VSUBS 0.010708f
C383 B.n108 VSUBS 0.010708f
C384 B.n109 VSUBS 0.010708f
C385 B.n110 VSUBS 0.010708f
C386 B.n111 VSUBS 0.010708f
C387 B.n112 VSUBS 0.010708f
C388 B.n113 VSUBS 0.010708f
C389 B.n114 VSUBS 0.010708f
C390 B.n115 VSUBS 0.010708f
C391 B.n116 VSUBS 0.010708f
C392 B.n117 VSUBS 0.010708f
C393 B.n118 VSUBS 0.010708f
C394 B.n119 VSUBS 0.010708f
C395 B.n120 VSUBS 0.010708f
C396 B.n121 VSUBS 0.010708f
C397 B.n122 VSUBS 0.010708f
C398 B.n123 VSUBS 0.024232f
C399 B.n124 VSUBS 0.010708f
C400 B.n125 VSUBS 0.010708f
C401 B.n126 VSUBS 0.010708f
C402 B.n127 VSUBS 0.010708f
C403 B.n128 VSUBS 0.010708f
C404 B.n129 VSUBS 0.010708f
C405 B.t7 VSUBS 0.071007f
C406 B.t8 VSUBS 0.096227f
C407 B.t6 VSUBS 0.580232f
C408 B.n130 VSUBS 0.124291f
C409 B.n131 VSUBS 0.09707f
C410 B.n132 VSUBS 0.02481f
C411 B.n133 VSUBS 0.010708f
C412 B.n134 VSUBS 0.010708f
C413 B.n135 VSUBS 0.010708f
C414 B.n136 VSUBS 0.010708f
C415 B.n137 VSUBS 0.010708f
C416 B.t10 VSUBS 0.071007f
C417 B.t11 VSUBS 0.096227f
C418 B.t9 VSUBS 0.580232f
C419 B.n138 VSUBS 0.124291f
C420 B.n139 VSUBS 0.09707f
C421 B.n140 VSUBS 0.010708f
C422 B.n141 VSUBS 0.010708f
C423 B.n142 VSUBS 0.010708f
C424 B.n143 VSUBS 0.010708f
C425 B.n144 VSUBS 0.010708f
C426 B.n145 VSUBS 0.02616f
C427 B.n146 VSUBS 0.010708f
C428 B.n147 VSUBS 0.010708f
C429 B.n148 VSUBS 0.010708f
C430 B.n149 VSUBS 0.010708f
C431 B.n150 VSUBS 0.010708f
C432 B.n151 VSUBS 0.010708f
C433 B.n152 VSUBS 0.010708f
C434 B.n153 VSUBS 0.010708f
C435 B.n154 VSUBS 0.010708f
C436 B.n155 VSUBS 0.010708f
C437 B.n156 VSUBS 0.010708f
C438 B.n157 VSUBS 0.010708f
C439 B.n158 VSUBS 0.010708f
C440 B.n159 VSUBS 0.010708f
C441 B.n160 VSUBS 0.010708f
C442 B.n161 VSUBS 0.010708f
C443 B.n162 VSUBS 0.010708f
C444 B.n163 VSUBS 0.010708f
C445 B.n164 VSUBS 0.010708f
C446 B.n165 VSUBS 0.010708f
C447 B.n166 VSUBS 0.010708f
C448 B.n167 VSUBS 0.010708f
C449 B.n168 VSUBS 0.010708f
C450 B.n169 VSUBS 0.010708f
C451 B.n170 VSUBS 0.010708f
C452 B.n171 VSUBS 0.010708f
C453 B.n172 VSUBS 0.010708f
C454 B.n173 VSUBS 0.010708f
C455 B.n174 VSUBS 0.010708f
C456 B.n175 VSUBS 0.010708f
C457 B.n176 VSUBS 0.010708f
C458 B.n177 VSUBS 0.010708f
C459 B.n178 VSUBS 0.010708f
C460 B.n179 VSUBS 0.010708f
C461 B.n180 VSUBS 0.010708f
C462 B.n181 VSUBS 0.010708f
C463 B.n182 VSUBS 0.010708f
C464 B.n183 VSUBS 0.010708f
C465 B.n184 VSUBS 0.010708f
C466 B.n185 VSUBS 0.010708f
C467 B.n186 VSUBS 0.010708f
C468 B.n187 VSUBS 0.010708f
C469 B.n188 VSUBS 0.010708f
C470 B.n189 VSUBS 0.010708f
C471 B.n190 VSUBS 0.010708f
C472 B.n191 VSUBS 0.010708f
C473 B.n192 VSUBS 0.010708f
C474 B.n193 VSUBS 0.010708f
C475 B.n194 VSUBS 0.010708f
C476 B.n195 VSUBS 0.010708f
C477 B.n196 VSUBS 0.010708f
C478 B.n197 VSUBS 0.010708f
C479 B.n198 VSUBS 0.010708f
C480 B.n199 VSUBS 0.010708f
C481 B.n200 VSUBS 0.010708f
C482 B.n201 VSUBS 0.010708f
C483 B.n202 VSUBS 0.010708f
C484 B.n203 VSUBS 0.010708f
C485 B.n204 VSUBS 0.010708f
C486 B.n205 VSUBS 0.010708f
C487 B.n206 VSUBS 0.010708f
C488 B.n207 VSUBS 0.010708f
C489 B.n208 VSUBS 0.010708f
C490 B.n209 VSUBS 0.010708f
C491 B.n210 VSUBS 0.010708f
C492 B.n211 VSUBS 0.010708f
C493 B.n212 VSUBS 0.010708f
C494 B.n213 VSUBS 0.010708f
C495 B.n214 VSUBS 0.010708f
C496 B.n215 VSUBS 0.010708f
C497 B.n216 VSUBS 0.010708f
C498 B.n217 VSUBS 0.010708f
C499 B.n218 VSUBS 0.010708f
C500 B.n219 VSUBS 0.010708f
C501 B.n220 VSUBS 0.010708f
C502 B.n221 VSUBS 0.010708f
C503 B.n222 VSUBS 0.010708f
C504 B.n223 VSUBS 0.010708f
C505 B.n224 VSUBS 0.010708f
C506 B.n225 VSUBS 0.010708f
C507 B.n226 VSUBS 0.010708f
C508 B.n227 VSUBS 0.010708f
C509 B.n228 VSUBS 0.010708f
C510 B.n229 VSUBS 0.010708f
C511 B.n230 VSUBS 0.010708f
C512 B.n231 VSUBS 0.010708f
C513 B.n232 VSUBS 0.010708f
C514 B.n233 VSUBS 0.010708f
C515 B.n234 VSUBS 0.010708f
C516 B.n235 VSUBS 0.010708f
C517 B.n236 VSUBS 0.010708f
C518 B.n237 VSUBS 0.010708f
C519 B.n238 VSUBS 0.010708f
C520 B.n239 VSUBS 0.010708f
C521 B.n240 VSUBS 0.010708f
C522 B.n241 VSUBS 0.010708f
C523 B.n242 VSUBS 0.010708f
C524 B.n243 VSUBS 0.010708f
C525 B.n244 VSUBS 0.010708f
C526 B.n245 VSUBS 0.010708f
C527 B.n246 VSUBS 0.010708f
C528 B.n247 VSUBS 0.010708f
C529 B.n248 VSUBS 0.010708f
C530 B.n249 VSUBS 0.010708f
C531 B.n250 VSUBS 0.010708f
C532 B.n251 VSUBS 0.010708f
C533 B.n252 VSUBS 0.010708f
C534 B.n253 VSUBS 0.010708f
C535 B.n254 VSUBS 0.010708f
C536 B.n255 VSUBS 0.010708f
C537 B.n256 VSUBS 0.010708f
C538 B.n257 VSUBS 0.010708f
C539 B.n258 VSUBS 0.010708f
C540 B.n259 VSUBS 0.010708f
C541 B.n260 VSUBS 0.010708f
C542 B.n261 VSUBS 0.010708f
C543 B.n262 VSUBS 0.010708f
C544 B.n263 VSUBS 0.010708f
C545 B.n264 VSUBS 0.010708f
C546 B.n265 VSUBS 0.010708f
C547 B.n266 VSUBS 0.010708f
C548 B.n267 VSUBS 0.010708f
C549 B.n268 VSUBS 0.010708f
C550 B.n269 VSUBS 0.010708f
C551 B.n270 VSUBS 0.010708f
C552 B.n271 VSUBS 0.010708f
C553 B.n272 VSUBS 0.010708f
C554 B.n273 VSUBS 0.010708f
C555 B.n274 VSUBS 0.024232f
C556 B.n275 VSUBS 0.024232f
C557 B.n276 VSUBS 0.02616f
C558 B.n277 VSUBS 0.010708f
C559 B.n278 VSUBS 0.010708f
C560 B.n279 VSUBS 0.010708f
C561 B.n280 VSUBS 0.010708f
C562 B.n281 VSUBS 0.010708f
C563 B.n282 VSUBS 0.010708f
C564 B.n283 VSUBS 0.010708f
C565 B.n284 VSUBS 0.010708f
C566 B.n285 VSUBS 0.010708f
C567 B.n286 VSUBS 0.010708f
C568 B.n287 VSUBS 0.010708f
C569 B.n288 VSUBS 0.010708f
C570 B.n289 VSUBS 0.010708f
C571 B.n290 VSUBS 0.010708f
C572 B.n291 VSUBS 0.010708f
C573 B.n292 VSUBS 0.010708f
C574 B.n293 VSUBS 0.010708f
C575 B.n294 VSUBS 0.007401f
C576 B.n295 VSUBS 0.02481f
C577 B.n296 VSUBS 0.008661f
C578 B.n297 VSUBS 0.010708f
C579 B.n298 VSUBS 0.010708f
C580 B.n299 VSUBS 0.010708f
C581 B.n300 VSUBS 0.010708f
C582 B.n301 VSUBS 0.010708f
C583 B.n302 VSUBS 0.010708f
C584 B.n303 VSUBS 0.010708f
C585 B.n304 VSUBS 0.010708f
C586 B.n305 VSUBS 0.010708f
C587 B.n306 VSUBS 0.010708f
C588 B.n307 VSUBS 0.010708f
C589 B.n308 VSUBS 0.008661f
C590 B.n309 VSUBS 0.010708f
C591 B.n310 VSUBS 0.010708f
C592 B.n311 VSUBS 0.007401f
C593 B.n312 VSUBS 0.010708f
C594 B.n313 VSUBS 0.010708f
C595 B.n314 VSUBS 0.010708f
C596 B.n315 VSUBS 0.010708f
C597 B.n316 VSUBS 0.010708f
C598 B.n317 VSUBS 0.010708f
C599 B.n318 VSUBS 0.010708f
C600 B.n319 VSUBS 0.010708f
C601 B.n320 VSUBS 0.010708f
C602 B.n321 VSUBS 0.010708f
C603 B.n322 VSUBS 0.010708f
C604 B.n323 VSUBS 0.010708f
C605 B.n324 VSUBS 0.010708f
C606 B.n325 VSUBS 0.010708f
C607 B.n326 VSUBS 0.010708f
C608 B.n327 VSUBS 0.010708f
C609 B.n328 VSUBS 0.02616f
C610 B.n329 VSUBS 0.02616f
C611 B.n330 VSUBS 0.024232f
C612 B.n331 VSUBS 0.010708f
C613 B.n332 VSUBS 0.010708f
C614 B.n333 VSUBS 0.010708f
C615 B.n334 VSUBS 0.010708f
C616 B.n335 VSUBS 0.010708f
C617 B.n336 VSUBS 0.010708f
C618 B.n337 VSUBS 0.010708f
C619 B.n338 VSUBS 0.010708f
C620 B.n339 VSUBS 0.010708f
C621 B.n340 VSUBS 0.010708f
C622 B.n341 VSUBS 0.010708f
C623 B.n342 VSUBS 0.010708f
C624 B.n343 VSUBS 0.010708f
C625 B.n344 VSUBS 0.010708f
C626 B.n345 VSUBS 0.010708f
C627 B.n346 VSUBS 0.010708f
C628 B.n347 VSUBS 0.010708f
C629 B.n348 VSUBS 0.010708f
C630 B.n349 VSUBS 0.010708f
C631 B.n350 VSUBS 0.010708f
C632 B.n351 VSUBS 0.010708f
C633 B.n352 VSUBS 0.010708f
C634 B.n353 VSUBS 0.010708f
C635 B.n354 VSUBS 0.010708f
C636 B.n355 VSUBS 0.010708f
C637 B.n356 VSUBS 0.010708f
C638 B.n357 VSUBS 0.010708f
C639 B.n358 VSUBS 0.010708f
C640 B.n359 VSUBS 0.010708f
C641 B.n360 VSUBS 0.010708f
C642 B.n361 VSUBS 0.010708f
C643 B.n362 VSUBS 0.010708f
C644 B.n363 VSUBS 0.010708f
C645 B.n364 VSUBS 0.010708f
C646 B.n365 VSUBS 0.010708f
C647 B.n366 VSUBS 0.010708f
C648 B.n367 VSUBS 0.010708f
C649 B.n368 VSUBS 0.010708f
C650 B.n369 VSUBS 0.010708f
C651 B.n370 VSUBS 0.010708f
C652 B.n371 VSUBS 0.010708f
C653 B.n372 VSUBS 0.010708f
C654 B.n373 VSUBS 0.010708f
C655 B.n374 VSUBS 0.010708f
C656 B.n375 VSUBS 0.010708f
C657 B.n376 VSUBS 0.010708f
C658 B.n377 VSUBS 0.010708f
C659 B.n378 VSUBS 0.010708f
C660 B.n379 VSUBS 0.010708f
C661 B.n380 VSUBS 0.010708f
C662 B.n381 VSUBS 0.010708f
C663 B.n382 VSUBS 0.010708f
C664 B.n383 VSUBS 0.010708f
C665 B.n384 VSUBS 0.010708f
C666 B.n385 VSUBS 0.010708f
C667 B.n386 VSUBS 0.010708f
C668 B.n387 VSUBS 0.010708f
C669 B.n388 VSUBS 0.010708f
C670 B.n389 VSUBS 0.010708f
C671 B.n390 VSUBS 0.010708f
C672 B.n391 VSUBS 0.010708f
C673 B.n392 VSUBS 0.010708f
C674 B.n393 VSUBS 0.010708f
C675 B.n394 VSUBS 0.010708f
C676 B.n395 VSUBS 0.010708f
C677 B.n396 VSUBS 0.010708f
C678 B.n397 VSUBS 0.010708f
C679 B.n398 VSUBS 0.010708f
C680 B.n399 VSUBS 0.010708f
C681 B.n400 VSUBS 0.010708f
C682 B.n401 VSUBS 0.010708f
C683 B.n402 VSUBS 0.010708f
C684 B.n403 VSUBS 0.010708f
C685 B.n404 VSUBS 0.010708f
C686 B.n405 VSUBS 0.010708f
C687 B.n406 VSUBS 0.010708f
C688 B.n407 VSUBS 0.010708f
C689 B.n408 VSUBS 0.010708f
C690 B.n409 VSUBS 0.010708f
C691 B.n410 VSUBS 0.010708f
C692 B.n411 VSUBS 0.010708f
C693 B.n412 VSUBS 0.010708f
C694 B.n413 VSUBS 0.010708f
C695 B.n414 VSUBS 0.010708f
C696 B.n415 VSUBS 0.010708f
C697 B.n416 VSUBS 0.010708f
C698 B.n417 VSUBS 0.010708f
C699 B.n418 VSUBS 0.010708f
C700 B.n419 VSUBS 0.010708f
C701 B.n420 VSUBS 0.010708f
C702 B.n421 VSUBS 0.010708f
C703 B.n422 VSUBS 0.010708f
C704 B.n423 VSUBS 0.010708f
C705 B.n424 VSUBS 0.010708f
C706 B.n425 VSUBS 0.010708f
C707 B.n426 VSUBS 0.010708f
C708 B.n427 VSUBS 0.010708f
C709 B.n428 VSUBS 0.010708f
C710 B.n429 VSUBS 0.010708f
C711 B.n430 VSUBS 0.010708f
C712 B.n431 VSUBS 0.010708f
C713 B.n432 VSUBS 0.010708f
C714 B.n433 VSUBS 0.010708f
C715 B.n434 VSUBS 0.010708f
C716 B.n435 VSUBS 0.010708f
C717 B.n436 VSUBS 0.010708f
C718 B.n437 VSUBS 0.010708f
C719 B.n438 VSUBS 0.010708f
C720 B.n439 VSUBS 0.010708f
C721 B.n440 VSUBS 0.010708f
C722 B.n441 VSUBS 0.010708f
C723 B.n442 VSUBS 0.010708f
C724 B.n443 VSUBS 0.010708f
C725 B.n444 VSUBS 0.010708f
C726 B.n445 VSUBS 0.010708f
C727 B.n446 VSUBS 0.010708f
C728 B.n447 VSUBS 0.010708f
C729 B.n448 VSUBS 0.010708f
C730 B.n449 VSUBS 0.010708f
C731 B.n450 VSUBS 0.010708f
C732 B.n451 VSUBS 0.010708f
C733 B.n452 VSUBS 0.010708f
C734 B.n453 VSUBS 0.010708f
C735 B.n454 VSUBS 0.010708f
C736 B.n455 VSUBS 0.010708f
C737 B.n456 VSUBS 0.010708f
C738 B.n457 VSUBS 0.010708f
C739 B.n458 VSUBS 0.010708f
C740 B.n459 VSUBS 0.010708f
C741 B.n460 VSUBS 0.010708f
C742 B.n461 VSUBS 0.010708f
C743 B.n462 VSUBS 0.010708f
C744 B.n463 VSUBS 0.010708f
C745 B.n464 VSUBS 0.010708f
C746 B.n465 VSUBS 0.010708f
C747 B.n466 VSUBS 0.010708f
C748 B.n467 VSUBS 0.010708f
C749 B.n468 VSUBS 0.010708f
C750 B.n469 VSUBS 0.010708f
C751 B.n470 VSUBS 0.010708f
C752 B.n471 VSUBS 0.010708f
C753 B.n472 VSUBS 0.010708f
C754 B.n473 VSUBS 0.010708f
C755 B.n474 VSUBS 0.010708f
C756 B.n475 VSUBS 0.010708f
C757 B.n476 VSUBS 0.010708f
C758 B.n477 VSUBS 0.010708f
C759 B.n478 VSUBS 0.010708f
C760 B.n479 VSUBS 0.010708f
C761 B.n480 VSUBS 0.010708f
C762 B.n481 VSUBS 0.010708f
C763 B.n482 VSUBS 0.010708f
C764 B.n483 VSUBS 0.010708f
C765 B.n484 VSUBS 0.010708f
C766 B.n485 VSUBS 0.010708f
C767 B.n486 VSUBS 0.010708f
C768 B.n487 VSUBS 0.010708f
C769 B.n488 VSUBS 0.010708f
C770 B.n489 VSUBS 0.010708f
C771 B.n490 VSUBS 0.010708f
C772 B.n491 VSUBS 0.010708f
C773 B.n492 VSUBS 0.010708f
C774 B.n493 VSUBS 0.010708f
C775 B.n494 VSUBS 0.010708f
C776 B.n495 VSUBS 0.010708f
C777 B.n496 VSUBS 0.010708f
C778 B.n497 VSUBS 0.010708f
C779 B.n498 VSUBS 0.010708f
C780 B.n499 VSUBS 0.010708f
C781 B.n500 VSUBS 0.010708f
C782 B.n501 VSUBS 0.010708f
C783 B.n502 VSUBS 0.010708f
C784 B.n503 VSUBS 0.010708f
C785 B.n504 VSUBS 0.010708f
C786 B.n505 VSUBS 0.010708f
C787 B.n506 VSUBS 0.010708f
C788 B.n507 VSUBS 0.010708f
C789 B.n508 VSUBS 0.010708f
C790 B.n509 VSUBS 0.010708f
C791 B.n510 VSUBS 0.010708f
C792 B.n511 VSUBS 0.010708f
C793 B.n512 VSUBS 0.010708f
C794 B.n513 VSUBS 0.010708f
C795 B.n514 VSUBS 0.010708f
C796 B.n515 VSUBS 0.010708f
C797 B.n516 VSUBS 0.010708f
C798 B.n517 VSUBS 0.010708f
C799 B.n518 VSUBS 0.010708f
C800 B.n519 VSUBS 0.010708f
C801 B.n520 VSUBS 0.010708f
C802 B.n521 VSUBS 0.010708f
C803 B.n522 VSUBS 0.010708f
C804 B.n523 VSUBS 0.010708f
C805 B.n524 VSUBS 0.010708f
C806 B.n525 VSUBS 0.010708f
C807 B.n526 VSUBS 0.010708f
C808 B.n527 VSUBS 0.010708f
C809 B.n528 VSUBS 0.025486f
C810 B.n529 VSUBS 0.024905f
C811 B.n530 VSUBS 0.02616f
C812 B.n531 VSUBS 0.010708f
C813 B.n532 VSUBS 0.010708f
C814 B.n533 VSUBS 0.010708f
C815 B.n534 VSUBS 0.010708f
C816 B.n535 VSUBS 0.010708f
C817 B.n536 VSUBS 0.010708f
C818 B.n537 VSUBS 0.010708f
C819 B.n538 VSUBS 0.010708f
C820 B.n539 VSUBS 0.010708f
C821 B.n540 VSUBS 0.010708f
C822 B.n541 VSUBS 0.010708f
C823 B.n542 VSUBS 0.010708f
C824 B.n543 VSUBS 0.010708f
C825 B.n544 VSUBS 0.010708f
C826 B.n545 VSUBS 0.010708f
C827 B.n546 VSUBS 0.010708f
C828 B.n547 VSUBS 0.007401f
C829 B.n548 VSUBS 0.010708f
C830 B.n549 VSUBS 0.010708f
C831 B.n550 VSUBS 0.008661f
C832 B.n551 VSUBS 0.010708f
C833 B.n552 VSUBS 0.010708f
C834 B.n553 VSUBS 0.010708f
C835 B.n554 VSUBS 0.010708f
C836 B.n555 VSUBS 0.010708f
C837 B.n556 VSUBS 0.010708f
C838 B.n557 VSUBS 0.010708f
C839 B.n558 VSUBS 0.010708f
C840 B.n559 VSUBS 0.010708f
C841 B.n560 VSUBS 0.010708f
C842 B.n561 VSUBS 0.010708f
C843 B.n562 VSUBS 0.008661f
C844 B.n563 VSUBS 0.02481f
C845 B.n564 VSUBS 0.007401f
C846 B.n565 VSUBS 0.010708f
C847 B.n566 VSUBS 0.010708f
C848 B.n567 VSUBS 0.010708f
C849 B.n568 VSUBS 0.010708f
C850 B.n569 VSUBS 0.010708f
C851 B.n570 VSUBS 0.010708f
C852 B.n571 VSUBS 0.010708f
C853 B.n572 VSUBS 0.010708f
C854 B.n573 VSUBS 0.010708f
C855 B.n574 VSUBS 0.010708f
C856 B.n575 VSUBS 0.010708f
C857 B.n576 VSUBS 0.010708f
C858 B.n577 VSUBS 0.010708f
C859 B.n578 VSUBS 0.010708f
C860 B.n579 VSUBS 0.010708f
C861 B.n580 VSUBS 0.010708f
C862 B.n581 VSUBS 0.010708f
C863 B.n582 VSUBS 0.02616f
C864 B.n583 VSUBS 0.024232f
C865 B.n584 VSUBS 0.024232f
C866 B.n585 VSUBS 0.010708f
C867 B.n586 VSUBS 0.010708f
C868 B.n587 VSUBS 0.010708f
C869 B.n588 VSUBS 0.010708f
C870 B.n589 VSUBS 0.010708f
C871 B.n590 VSUBS 0.010708f
C872 B.n591 VSUBS 0.010708f
C873 B.n592 VSUBS 0.010708f
C874 B.n593 VSUBS 0.010708f
C875 B.n594 VSUBS 0.010708f
C876 B.n595 VSUBS 0.010708f
C877 B.n596 VSUBS 0.010708f
C878 B.n597 VSUBS 0.010708f
C879 B.n598 VSUBS 0.010708f
C880 B.n599 VSUBS 0.010708f
C881 B.n600 VSUBS 0.010708f
C882 B.n601 VSUBS 0.010708f
C883 B.n602 VSUBS 0.010708f
C884 B.n603 VSUBS 0.010708f
C885 B.n604 VSUBS 0.010708f
C886 B.n605 VSUBS 0.010708f
C887 B.n606 VSUBS 0.010708f
C888 B.n607 VSUBS 0.010708f
C889 B.n608 VSUBS 0.010708f
C890 B.n609 VSUBS 0.010708f
C891 B.n610 VSUBS 0.010708f
C892 B.n611 VSUBS 0.010708f
C893 B.n612 VSUBS 0.010708f
C894 B.n613 VSUBS 0.010708f
C895 B.n614 VSUBS 0.010708f
C896 B.n615 VSUBS 0.010708f
C897 B.n616 VSUBS 0.010708f
C898 B.n617 VSUBS 0.010708f
C899 B.n618 VSUBS 0.010708f
C900 B.n619 VSUBS 0.010708f
C901 B.n620 VSUBS 0.010708f
C902 B.n621 VSUBS 0.010708f
C903 B.n622 VSUBS 0.010708f
C904 B.n623 VSUBS 0.010708f
C905 B.n624 VSUBS 0.010708f
C906 B.n625 VSUBS 0.010708f
C907 B.n626 VSUBS 0.010708f
C908 B.n627 VSUBS 0.010708f
C909 B.n628 VSUBS 0.010708f
C910 B.n629 VSUBS 0.010708f
C911 B.n630 VSUBS 0.010708f
C912 B.n631 VSUBS 0.010708f
C913 B.n632 VSUBS 0.010708f
C914 B.n633 VSUBS 0.010708f
C915 B.n634 VSUBS 0.010708f
C916 B.n635 VSUBS 0.010708f
C917 B.n636 VSUBS 0.010708f
C918 B.n637 VSUBS 0.010708f
C919 B.n638 VSUBS 0.010708f
C920 B.n639 VSUBS 0.010708f
C921 B.n640 VSUBS 0.010708f
C922 B.n641 VSUBS 0.010708f
C923 B.n642 VSUBS 0.010708f
C924 B.n643 VSUBS 0.010708f
C925 B.n644 VSUBS 0.010708f
C926 B.n645 VSUBS 0.010708f
C927 B.n646 VSUBS 0.010708f
C928 B.n647 VSUBS 0.010708f
C929 B.n648 VSUBS 0.010708f
C930 B.n649 VSUBS 0.010708f
C931 B.n650 VSUBS 0.010708f
C932 B.n651 VSUBS 0.010708f
C933 B.n652 VSUBS 0.010708f
C934 B.n653 VSUBS 0.010708f
C935 B.n654 VSUBS 0.010708f
C936 B.n655 VSUBS 0.010708f
C937 B.n656 VSUBS 0.010708f
C938 B.n657 VSUBS 0.010708f
C939 B.n658 VSUBS 0.010708f
C940 B.n659 VSUBS 0.010708f
C941 B.n660 VSUBS 0.010708f
C942 B.n661 VSUBS 0.010708f
C943 B.n662 VSUBS 0.010708f
C944 B.n663 VSUBS 0.010708f
C945 B.n664 VSUBS 0.010708f
C946 B.n665 VSUBS 0.010708f
C947 B.n666 VSUBS 0.010708f
C948 B.n667 VSUBS 0.010708f
C949 B.n668 VSUBS 0.010708f
C950 B.n669 VSUBS 0.010708f
C951 B.n670 VSUBS 0.010708f
C952 B.n671 VSUBS 0.010708f
C953 B.n672 VSUBS 0.010708f
C954 B.n673 VSUBS 0.010708f
C955 B.n674 VSUBS 0.010708f
C956 B.n675 VSUBS 0.010708f
C957 B.n676 VSUBS 0.010708f
C958 B.n677 VSUBS 0.010708f
C959 B.n678 VSUBS 0.010708f
C960 B.n679 VSUBS 0.010708f
C961 B.n680 VSUBS 0.010708f
C962 B.n681 VSUBS 0.010708f
C963 B.n682 VSUBS 0.010708f
C964 B.n683 VSUBS 0.024247f
.ends

