* NGSPICE file created from diff_pair_sample_0132.ext - technology: sky130A

.subckt diff_pair_sample_0132 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t2 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=1.3464 ps=8.49 w=8.16 l=2.17
X1 VTAIL.t4 VN.t0 VDD2.t7 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=3.1824 pd=17.1 as=1.3464 ps=8.49 w=8.16 l=2.17
X2 VTAIL.t14 VP.t1 VDD1.t3 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=3.1824 pd=17.1 as=1.3464 ps=8.49 w=8.16 l=2.17
X3 VTAIL.t13 VP.t2 VDD1.t1 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=3.1824 pd=17.1 as=1.3464 ps=8.49 w=8.16 l=2.17
X4 VDD2.t6 VN.t1 VTAIL.t5 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=3.1824 ps=17.1 w=8.16 l=2.17
X5 VDD2.t5 VN.t2 VTAIL.t0 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=1.3464 ps=8.49 w=8.16 l=2.17
X6 VTAIL.t12 VP.t3 VDD1.t0 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=1.3464 ps=8.49 w=8.16 l=2.17
X7 VDD1.t6 VP.t4 VTAIL.t11 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=3.1824 ps=17.1 w=8.16 l=2.17
X8 B.t11 B.t9 B.t10 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=3.1824 pd=17.1 as=0 ps=0 w=8.16 l=2.17
X9 VDD2.t4 VN.t3 VTAIL.t1 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=3.1824 ps=17.1 w=8.16 l=2.17
X10 B.t8 B.t6 B.t7 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=3.1824 pd=17.1 as=0 ps=0 w=8.16 l=2.17
X11 VDD1.t5 VP.t5 VTAIL.t10 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=1.3464 ps=8.49 w=8.16 l=2.17
X12 VDD2.t3 VN.t4 VTAIL.t2 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=1.3464 ps=8.49 w=8.16 l=2.17
X13 VDD1.t4 VP.t6 VTAIL.t9 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=1.3464 ps=8.49 w=8.16 l=2.17
X14 B.t5 B.t3 B.t4 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=3.1824 pd=17.1 as=0 ps=0 w=8.16 l=2.17
X15 VTAIL.t3 VN.t5 VDD2.t2 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=3.1824 pd=17.1 as=1.3464 ps=8.49 w=8.16 l=2.17
X16 VDD1.t7 VP.t7 VTAIL.t8 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=3.1824 ps=17.1 w=8.16 l=2.17
X17 VTAIL.t6 VN.t6 VDD2.t1 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=1.3464 ps=8.49 w=8.16 l=2.17
X18 B.t2 B.t0 B.t1 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=3.1824 pd=17.1 as=0 ps=0 w=8.16 l=2.17
X19 VTAIL.t7 VN.t7 VDD2.t0 w_n3470_n2600# sky130_fd_pr__pfet_01v8 ad=1.3464 pd=8.49 as=1.3464 ps=8.49 w=8.16 l=2.17
R0 VP.n16 VP.n15 161.3
R1 VP.n17 VP.n12 161.3
R2 VP.n19 VP.n18 161.3
R3 VP.n20 VP.n11 161.3
R4 VP.n22 VP.n21 161.3
R5 VP.n24 VP.n10 161.3
R6 VP.n26 VP.n25 161.3
R7 VP.n27 VP.n9 161.3
R8 VP.n29 VP.n28 161.3
R9 VP.n30 VP.n8 161.3
R10 VP.n58 VP.n0 161.3
R11 VP.n57 VP.n56 161.3
R12 VP.n55 VP.n1 161.3
R13 VP.n54 VP.n53 161.3
R14 VP.n52 VP.n2 161.3
R15 VP.n50 VP.n49 161.3
R16 VP.n48 VP.n3 161.3
R17 VP.n47 VP.n46 161.3
R18 VP.n45 VP.n4 161.3
R19 VP.n44 VP.n43 161.3
R20 VP.n42 VP.n41 161.3
R21 VP.n40 VP.n6 161.3
R22 VP.n39 VP.n38 161.3
R23 VP.n37 VP.n7 161.3
R24 VP.n36 VP.n35 161.3
R25 VP.n14 VP.t1 122.703
R26 VP.n34 VP.n33 98.6123
R27 VP.n60 VP.n59 98.6123
R28 VP.n32 VP.n31 98.6123
R29 VP.n34 VP.t2 90.6254
R30 VP.n5 VP.t6 90.6254
R31 VP.n51 VP.t3 90.6254
R32 VP.n59 VP.t7 90.6254
R33 VP.n31 VP.t4 90.6254
R34 VP.n23 VP.t0 90.6254
R35 VP.n13 VP.t5 90.6254
R36 VP.n14 VP.n13 59.4159
R37 VP.n33 VP.n32 45.9239
R38 VP.n39 VP.n7 40.577
R39 VP.n40 VP.n39 40.577
R40 VP.n46 VP.n45 40.577
R41 VP.n46 VP.n3 40.577
R42 VP.n53 VP.n1 40.577
R43 VP.n57 VP.n1 40.577
R44 VP.n29 VP.n9 40.577
R45 VP.n25 VP.n9 40.577
R46 VP.n18 VP.n11 40.577
R47 VP.n18 VP.n17 40.577
R48 VP.n35 VP.n7 24.5923
R49 VP.n41 VP.n40 24.5923
R50 VP.n45 VP.n44 24.5923
R51 VP.n50 VP.n3 24.5923
R52 VP.n53 VP.n52 24.5923
R53 VP.n58 VP.n57 24.5923
R54 VP.n30 VP.n29 24.5923
R55 VP.n22 VP.n11 24.5923
R56 VP.n25 VP.n24 24.5923
R57 VP.n17 VP.n16 24.5923
R58 VP.n35 VP.n34 12.2964
R59 VP.n41 VP.n5 12.2964
R60 VP.n44 VP.n5 12.2964
R61 VP.n51 VP.n50 12.2964
R62 VP.n52 VP.n51 12.2964
R63 VP.n59 VP.n58 12.2964
R64 VP.n31 VP.n30 12.2964
R65 VP.n23 VP.n22 12.2964
R66 VP.n24 VP.n23 12.2964
R67 VP.n16 VP.n13 12.2964
R68 VP.n15 VP.n14 9.706
R69 VP.n32 VP.n8 0.278335
R70 VP.n36 VP.n33 0.278335
R71 VP.n60 VP.n0 0.278335
R72 VP.n15 VP.n12 0.189894
R73 VP.n19 VP.n12 0.189894
R74 VP.n20 VP.n19 0.189894
R75 VP.n21 VP.n20 0.189894
R76 VP.n21 VP.n10 0.189894
R77 VP.n26 VP.n10 0.189894
R78 VP.n27 VP.n26 0.189894
R79 VP.n28 VP.n27 0.189894
R80 VP.n28 VP.n8 0.189894
R81 VP.n37 VP.n36 0.189894
R82 VP.n38 VP.n37 0.189894
R83 VP.n38 VP.n6 0.189894
R84 VP.n42 VP.n6 0.189894
R85 VP.n43 VP.n42 0.189894
R86 VP.n43 VP.n4 0.189894
R87 VP.n47 VP.n4 0.189894
R88 VP.n48 VP.n47 0.189894
R89 VP.n49 VP.n48 0.189894
R90 VP.n49 VP.n2 0.189894
R91 VP.n54 VP.n2 0.189894
R92 VP.n55 VP.n54 0.189894
R93 VP.n56 VP.n55 0.189894
R94 VP.n56 VP.n0 0.189894
R95 VP VP.n60 0.153485
R96 VDD1 VDD1.n0 82.4206
R97 VDD1.n3 VDD1.n2 82.3068
R98 VDD1.n3 VDD1.n1 82.3068
R99 VDD1.n5 VDD1.n4 81.2847
R100 VDD1.n5 VDD1.n3 41.0311
R101 VDD1.n4 VDD1.t2 3.98396
R102 VDD1.n4 VDD1.t6 3.98396
R103 VDD1.n0 VDD1.t3 3.98396
R104 VDD1.n0 VDD1.t5 3.98396
R105 VDD1.n2 VDD1.t0 3.98396
R106 VDD1.n2 VDD1.t7 3.98396
R107 VDD1.n1 VDD1.t1 3.98396
R108 VDD1.n1 VDD1.t4 3.98396
R109 VDD1 VDD1.n5 1.0199
R110 VTAIL.n11 VTAIL.t14 68.5894
R111 VTAIL.n10 VTAIL.t1 68.5894
R112 VTAIL.n7 VTAIL.t4 68.5894
R113 VTAIL.n15 VTAIL.t5 68.5893
R114 VTAIL.n2 VTAIL.t3 68.5893
R115 VTAIL.n3 VTAIL.t8 68.5893
R116 VTAIL.n6 VTAIL.t13 68.5893
R117 VTAIL.n14 VTAIL.t11 68.5893
R118 VTAIL.n13 VTAIL.n12 64.6061
R119 VTAIL.n9 VTAIL.n8 64.6061
R120 VTAIL.n1 VTAIL.n0 64.6058
R121 VTAIL.n5 VTAIL.n4 64.6058
R122 VTAIL.n15 VTAIL.n14 21.5565
R123 VTAIL.n7 VTAIL.n6 21.5565
R124 VTAIL.n0 VTAIL.t0 3.98396
R125 VTAIL.n0 VTAIL.t6 3.98396
R126 VTAIL.n4 VTAIL.t9 3.98396
R127 VTAIL.n4 VTAIL.t12 3.98396
R128 VTAIL.n12 VTAIL.t10 3.98396
R129 VTAIL.n12 VTAIL.t15 3.98396
R130 VTAIL.n8 VTAIL.t2 3.98396
R131 VTAIL.n8 VTAIL.t7 3.98396
R132 VTAIL.n9 VTAIL.n7 2.15567
R133 VTAIL.n10 VTAIL.n9 2.15567
R134 VTAIL.n13 VTAIL.n11 2.15567
R135 VTAIL.n14 VTAIL.n13 2.15567
R136 VTAIL.n6 VTAIL.n5 2.15567
R137 VTAIL.n5 VTAIL.n3 2.15567
R138 VTAIL.n2 VTAIL.n1 2.15567
R139 VTAIL VTAIL.n15 2.09748
R140 VTAIL.n11 VTAIL.n10 0.470328
R141 VTAIL.n3 VTAIL.n2 0.470328
R142 VTAIL VTAIL.n1 0.0586897
R143 VN.n47 VN.n25 161.3
R144 VN.n46 VN.n45 161.3
R145 VN.n44 VN.n26 161.3
R146 VN.n43 VN.n42 161.3
R147 VN.n41 VN.n27 161.3
R148 VN.n39 VN.n38 161.3
R149 VN.n37 VN.n28 161.3
R150 VN.n36 VN.n35 161.3
R151 VN.n34 VN.n29 161.3
R152 VN.n33 VN.n32 161.3
R153 VN.n22 VN.n0 161.3
R154 VN.n21 VN.n20 161.3
R155 VN.n19 VN.n1 161.3
R156 VN.n18 VN.n17 161.3
R157 VN.n16 VN.n2 161.3
R158 VN.n14 VN.n13 161.3
R159 VN.n12 VN.n3 161.3
R160 VN.n11 VN.n10 161.3
R161 VN.n9 VN.n4 161.3
R162 VN.n8 VN.n7 161.3
R163 VN.n6 VN.t5 122.703
R164 VN.n31 VN.t3 122.703
R165 VN.n24 VN.n23 98.6123
R166 VN.n49 VN.n48 98.6123
R167 VN.n5 VN.t2 90.6254
R168 VN.n15 VN.t6 90.6254
R169 VN.n23 VN.t1 90.6254
R170 VN.n30 VN.t7 90.6254
R171 VN.n40 VN.t4 90.6254
R172 VN.n48 VN.t0 90.6254
R173 VN.n6 VN.n5 59.4159
R174 VN.n31 VN.n30 59.4159
R175 VN VN.n49 46.2027
R176 VN.n10 VN.n9 40.577
R177 VN.n10 VN.n3 40.577
R178 VN.n17 VN.n1 40.577
R179 VN.n21 VN.n1 40.577
R180 VN.n35 VN.n34 40.577
R181 VN.n35 VN.n28 40.577
R182 VN.n42 VN.n26 40.577
R183 VN.n46 VN.n26 40.577
R184 VN.n9 VN.n8 24.5923
R185 VN.n14 VN.n3 24.5923
R186 VN.n17 VN.n16 24.5923
R187 VN.n22 VN.n21 24.5923
R188 VN.n34 VN.n33 24.5923
R189 VN.n42 VN.n41 24.5923
R190 VN.n39 VN.n28 24.5923
R191 VN.n47 VN.n46 24.5923
R192 VN.n8 VN.n5 12.2964
R193 VN.n15 VN.n14 12.2964
R194 VN.n16 VN.n15 12.2964
R195 VN.n23 VN.n22 12.2964
R196 VN.n33 VN.n30 12.2964
R197 VN.n41 VN.n40 12.2964
R198 VN.n40 VN.n39 12.2964
R199 VN.n48 VN.n47 12.2964
R200 VN.n32 VN.n31 9.706
R201 VN.n7 VN.n6 9.706
R202 VN.n49 VN.n25 0.278335
R203 VN.n24 VN.n0 0.278335
R204 VN.n45 VN.n25 0.189894
R205 VN.n45 VN.n44 0.189894
R206 VN.n44 VN.n43 0.189894
R207 VN.n43 VN.n27 0.189894
R208 VN.n38 VN.n27 0.189894
R209 VN.n38 VN.n37 0.189894
R210 VN.n37 VN.n36 0.189894
R211 VN.n36 VN.n29 0.189894
R212 VN.n32 VN.n29 0.189894
R213 VN.n7 VN.n4 0.189894
R214 VN.n11 VN.n4 0.189894
R215 VN.n12 VN.n11 0.189894
R216 VN.n13 VN.n12 0.189894
R217 VN.n13 VN.n2 0.189894
R218 VN.n18 VN.n2 0.189894
R219 VN.n19 VN.n18 0.189894
R220 VN.n20 VN.n19 0.189894
R221 VN.n20 VN.n0 0.189894
R222 VN VN.n24 0.153485
R223 VDD2.n2 VDD2.n1 82.3068
R224 VDD2.n2 VDD2.n0 82.3068
R225 VDD2 VDD2.n5 82.3041
R226 VDD2.n4 VDD2.n3 81.2849
R227 VDD2.n4 VDD2.n2 40.4481
R228 VDD2.n5 VDD2.t0 3.98396
R229 VDD2.n5 VDD2.t4 3.98396
R230 VDD2.n3 VDD2.t7 3.98396
R231 VDD2.n3 VDD2.t3 3.98396
R232 VDD2.n1 VDD2.t1 3.98396
R233 VDD2.n1 VDD2.t6 3.98396
R234 VDD2.n0 VDD2.t2 3.98396
R235 VDD2.n0 VDD2.t5 3.98396
R236 VDD2 VDD2.n4 1.13628
R237 B.n481 B.n64 585
R238 B.n483 B.n482 585
R239 B.n484 B.n63 585
R240 B.n486 B.n485 585
R241 B.n487 B.n62 585
R242 B.n489 B.n488 585
R243 B.n490 B.n61 585
R244 B.n492 B.n491 585
R245 B.n493 B.n60 585
R246 B.n495 B.n494 585
R247 B.n496 B.n59 585
R248 B.n498 B.n497 585
R249 B.n499 B.n58 585
R250 B.n501 B.n500 585
R251 B.n502 B.n57 585
R252 B.n504 B.n503 585
R253 B.n505 B.n56 585
R254 B.n507 B.n506 585
R255 B.n508 B.n55 585
R256 B.n510 B.n509 585
R257 B.n511 B.n54 585
R258 B.n513 B.n512 585
R259 B.n514 B.n53 585
R260 B.n516 B.n515 585
R261 B.n517 B.n52 585
R262 B.n519 B.n518 585
R263 B.n520 B.n51 585
R264 B.n522 B.n521 585
R265 B.n523 B.n47 585
R266 B.n525 B.n524 585
R267 B.n526 B.n46 585
R268 B.n528 B.n527 585
R269 B.n529 B.n45 585
R270 B.n531 B.n530 585
R271 B.n532 B.n44 585
R272 B.n534 B.n533 585
R273 B.n535 B.n43 585
R274 B.n537 B.n536 585
R275 B.n538 B.n42 585
R276 B.n540 B.n539 585
R277 B.n542 B.n39 585
R278 B.n544 B.n543 585
R279 B.n545 B.n38 585
R280 B.n547 B.n546 585
R281 B.n548 B.n37 585
R282 B.n550 B.n549 585
R283 B.n551 B.n36 585
R284 B.n553 B.n552 585
R285 B.n554 B.n35 585
R286 B.n556 B.n555 585
R287 B.n557 B.n34 585
R288 B.n559 B.n558 585
R289 B.n560 B.n33 585
R290 B.n562 B.n561 585
R291 B.n563 B.n32 585
R292 B.n565 B.n564 585
R293 B.n566 B.n31 585
R294 B.n568 B.n567 585
R295 B.n569 B.n30 585
R296 B.n571 B.n570 585
R297 B.n572 B.n29 585
R298 B.n574 B.n573 585
R299 B.n575 B.n28 585
R300 B.n577 B.n576 585
R301 B.n578 B.n27 585
R302 B.n580 B.n579 585
R303 B.n581 B.n26 585
R304 B.n583 B.n582 585
R305 B.n584 B.n25 585
R306 B.n586 B.n585 585
R307 B.n480 B.n479 585
R308 B.n478 B.n65 585
R309 B.n477 B.n476 585
R310 B.n475 B.n66 585
R311 B.n474 B.n473 585
R312 B.n472 B.n67 585
R313 B.n471 B.n470 585
R314 B.n469 B.n68 585
R315 B.n468 B.n467 585
R316 B.n466 B.n69 585
R317 B.n465 B.n464 585
R318 B.n463 B.n70 585
R319 B.n462 B.n461 585
R320 B.n460 B.n71 585
R321 B.n459 B.n458 585
R322 B.n457 B.n72 585
R323 B.n456 B.n455 585
R324 B.n454 B.n73 585
R325 B.n453 B.n452 585
R326 B.n451 B.n74 585
R327 B.n450 B.n449 585
R328 B.n448 B.n75 585
R329 B.n447 B.n446 585
R330 B.n445 B.n76 585
R331 B.n444 B.n443 585
R332 B.n442 B.n77 585
R333 B.n441 B.n440 585
R334 B.n439 B.n78 585
R335 B.n438 B.n437 585
R336 B.n436 B.n79 585
R337 B.n435 B.n434 585
R338 B.n433 B.n80 585
R339 B.n432 B.n431 585
R340 B.n430 B.n81 585
R341 B.n429 B.n428 585
R342 B.n427 B.n82 585
R343 B.n426 B.n425 585
R344 B.n424 B.n83 585
R345 B.n423 B.n422 585
R346 B.n421 B.n84 585
R347 B.n420 B.n419 585
R348 B.n418 B.n85 585
R349 B.n417 B.n416 585
R350 B.n415 B.n86 585
R351 B.n414 B.n413 585
R352 B.n412 B.n87 585
R353 B.n411 B.n410 585
R354 B.n409 B.n88 585
R355 B.n408 B.n407 585
R356 B.n406 B.n89 585
R357 B.n405 B.n404 585
R358 B.n403 B.n90 585
R359 B.n402 B.n401 585
R360 B.n400 B.n91 585
R361 B.n399 B.n398 585
R362 B.n397 B.n92 585
R363 B.n396 B.n395 585
R364 B.n394 B.n93 585
R365 B.n393 B.n392 585
R366 B.n391 B.n94 585
R367 B.n390 B.n389 585
R368 B.n388 B.n95 585
R369 B.n387 B.n386 585
R370 B.n385 B.n96 585
R371 B.n384 B.n383 585
R372 B.n382 B.n97 585
R373 B.n381 B.n380 585
R374 B.n379 B.n98 585
R375 B.n378 B.n377 585
R376 B.n376 B.n99 585
R377 B.n375 B.n374 585
R378 B.n373 B.n100 585
R379 B.n372 B.n371 585
R380 B.n370 B.n101 585
R381 B.n369 B.n368 585
R382 B.n367 B.n102 585
R383 B.n366 B.n365 585
R384 B.n364 B.n103 585
R385 B.n363 B.n362 585
R386 B.n361 B.n104 585
R387 B.n360 B.n359 585
R388 B.n358 B.n105 585
R389 B.n357 B.n356 585
R390 B.n355 B.n106 585
R391 B.n354 B.n353 585
R392 B.n352 B.n107 585
R393 B.n351 B.n350 585
R394 B.n349 B.n108 585
R395 B.n348 B.n347 585
R396 B.n346 B.n109 585
R397 B.n345 B.n344 585
R398 B.n238 B.n149 585
R399 B.n240 B.n239 585
R400 B.n241 B.n148 585
R401 B.n243 B.n242 585
R402 B.n244 B.n147 585
R403 B.n246 B.n245 585
R404 B.n247 B.n146 585
R405 B.n249 B.n248 585
R406 B.n250 B.n145 585
R407 B.n252 B.n251 585
R408 B.n253 B.n144 585
R409 B.n255 B.n254 585
R410 B.n256 B.n143 585
R411 B.n258 B.n257 585
R412 B.n259 B.n142 585
R413 B.n261 B.n260 585
R414 B.n262 B.n141 585
R415 B.n264 B.n263 585
R416 B.n265 B.n140 585
R417 B.n267 B.n266 585
R418 B.n268 B.n139 585
R419 B.n270 B.n269 585
R420 B.n271 B.n138 585
R421 B.n273 B.n272 585
R422 B.n274 B.n137 585
R423 B.n276 B.n275 585
R424 B.n277 B.n136 585
R425 B.n279 B.n278 585
R426 B.n280 B.n135 585
R427 B.n282 B.n281 585
R428 B.n284 B.n132 585
R429 B.n286 B.n285 585
R430 B.n287 B.n131 585
R431 B.n289 B.n288 585
R432 B.n290 B.n130 585
R433 B.n292 B.n291 585
R434 B.n293 B.n129 585
R435 B.n295 B.n294 585
R436 B.n296 B.n128 585
R437 B.n298 B.n297 585
R438 B.n300 B.n299 585
R439 B.n301 B.n124 585
R440 B.n303 B.n302 585
R441 B.n304 B.n123 585
R442 B.n306 B.n305 585
R443 B.n307 B.n122 585
R444 B.n309 B.n308 585
R445 B.n310 B.n121 585
R446 B.n312 B.n311 585
R447 B.n313 B.n120 585
R448 B.n315 B.n314 585
R449 B.n316 B.n119 585
R450 B.n318 B.n317 585
R451 B.n319 B.n118 585
R452 B.n321 B.n320 585
R453 B.n322 B.n117 585
R454 B.n324 B.n323 585
R455 B.n325 B.n116 585
R456 B.n327 B.n326 585
R457 B.n328 B.n115 585
R458 B.n330 B.n329 585
R459 B.n331 B.n114 585
R460 B.n333 B.n332 585
R461 B.n334 B.n113 585
R462 B.n336 B.n335 585
R463 B.n337 B.n112 585
R464 B.n339 B.n338 585
R465 B.n340 B.n111 585
R466 B.n342 B.n341 585
R467 B.n343 B.n110 585
R468 B.n237 B.n236 585
R469 B.n235 B.n150 585
R470 B.n234 B.n233 585
R471 B.n232 B.n151 585
R472 B.n231 B.n230 585
R473 B.n229 B.n152 585
R474 B.n228 B.n227 585
R475 B.n226 B.n153 585
R476 B.n225 B.n224 585
R477 B.n223 B.n154 585
R478 B.n222 B.n221 585
R479 B.n220 B.n155 585
R480 B.n219 B.n218 585
R481 B.n217 B.n156 585
R482 B.n216 B.n215 585
R483 B.n214 B.n157 585
R484 B.n213 B.n212 585
R485 B.n211 B.n158 585
R486 B.n210 B.n209 585
R487 B.n208 B.n159 585
R488 B.n207 B.n206 585
R489 B.n205 B.n160 585
R490 B.n204 B.n203 585
R491 B.n202 B.n161 585
R492 B.n201 B.n200 585
R493 B.n199 B.n162 585
R494 B.n198 B.n197 585
R495 B.n196 B.n163 585
R496 B.n195 B.n194 585
R497 B.n193 B.n164 585
R498 B.n192 B.n191 585
R499 B.n190 B.n165 585
R500 B.n189 B.n188 585
R501 B.n187 B.n166 585
R502 B.n186 B.n185 585
R503 B.n184 B.n167 585
R504 B.n183 B.n182 585
R505 B.n181 B.n168 585
R506 B.n180 B.n179 585
R507 B.n178 B.n169 585
R508 B.n177 B.n176 585
R509 B.n175 B.n170 585
R510 B.n174 B.n173 585
R511 B.n172 B.n171 585
R512 B.n2 B.n0 585
R513 B.n653 B.n1 585
R514 B.n652 B.n651 585
R515 B.n650 B.n3 585
R516 B.n649 B.n648 585
R517 B.n647 B.n4 585
R518 B.n646 B.n645 585
R519 B.n644 B.n5 585
R520 B.n643 B.n642 585
R521 B.n641 B.n6 585
R522 B.n640 B.n639 585
R523 B.n638 B.n7 585
R524 B.n637 B.n636 585
R525 B.n635 B.n8 585
R526 B.n634 B.n633 585
R527 B.n632 B.n9 585
R528 B.n631 B.n630 585
R529 B.n629 B.n10 585
R530 B.n628 B.n627 585
R531 B.n626 B.n11 585
R532 B.n625 B.n624 585
R533 B.n623 B.n12 585
R534 B.n622 B.n621 585
R535 B.n620 B.n13 585
R536 B.n619 B.n618 585
R537 B.n617 B.n14 585
R538 B.n616 B.n615 585
R539 B.n614 B.n15 585
R540 B.n613 B.n612 585
R541 B.n611 B.n16 585
R542 B.n610 B.n609 585
R543 B.n608 B.n17 585
R544 B.n607 B.n606 585
R545 B.n605 B.n18 585
R546 B.n604 B.n603 585
R547 B.n602 B.n19 585
R548 B.n601 B.n600 585
R549 B.n599 B.n20 585
R550 B.n598 B.n597 585
R551 B.n596 B.n21 585
R552 B.n595 B.n594 585
R553 B.n593 B.n22 585
R554 B.n592 B.n591 585
R555 B.n590 B.n23 585
R556 B.n589 B.n588 585
R557 B.n587 B.n24 585
R558 B.n655 B.n654 585
R559 B.n238 B.n237 497.305
R560 B.n587 B.n586 497.305
R561 B.n345 B.n110 497.305
R562 B.n479 B.n64 497.305
R563 B.n125 B.t6 297.916
R564 B.n133 B.t0 297.916
R565 B.n40 B.t9 297.916
R566 B.n48 B.t3 297.916
R567 B.n237 B.n150 163.367
R568 B.n233 B.n150 163.367
R569 B.n233 B.n232 163.367
R570 B.n232 B.n231 163.367
R571 B.n231 B.n152 163.367
R572 B.n227 B.n152 163.367
R573 B.n227 B.n226 163.367
R574 B.n226 B.n225 163.367
R575 B.n225 B.n154 163.367
R576 B.n221 B.n154 163.367
R577 B.n221 B.n220 163.367
R578 B.n220 B.n219 163.367
R579 B.n219 B.n156 163.367
R580 B.n215 B.n156 163.367
R581 B.n215 B.n214 163.367
R582 B.n214 B.n213 163.367
R583 B.n213 B.n158 163.367
R584 B.n209 B.n158 163.367
R585 B.n209 B.n208 163.367
R586 B.n208 B.n207 163.367
R587 B.n207 B.n160 163.367
R588 B.n203 B.n160 163.367
R589 B.n203 B.n202 163.367
R590 B.n202 B.n201 163.367
R591 B.n201 B.n162 163.367
R592 B.n197 B.n162 163.367
R593 B.n197 B.n196 163.367
R594 B.n196 B.n195 163.367
R595 B.n195 B.n164 163.367
R596 B.n191 B.n164 163.367
R597 B.n191 B.n190 163.367
R598 B.n190 B.n189 163.367
R599 B.n189 B.n166 163.367
R600 B.n185 B.n166 163.367
R601 B.n185 B.n184 163.367
R602 B.n184 B.n183 163.367
R603 B.n183 B.n168 163.367
R604 B.n179 B.n168 163.367
R605 B.n179 B.n178 163.367
R606 B.n178 B.n177 163.367
R607 B.n177 B.n170 163.367
R608 B.n173 B.n170 163.367
R609 B.n173 B.n172 163.367
R610 B.n172 B.n2 163.367
R611 B.n654 B.n2 163.367
R612 B.n654 B.n653 163.367
R613 B.n653 B.n652 163.367
R614 B.n652 B.n3 163.367
R615 B.n648 B.n3 163.367
R616 B.n648 B.n647 163.367
R617 B.n647 B.n646 163.367
R618 B.n646 B.n5 163.367
R619 B.n642 B.n5 163.367
R620 B.n642 B.n641 163.367
R621 B.n641 B.n640 163.367
R622 B.n640 B.n7 163.367
R623 B.n636 B.n7 163.367
R624 B.n636 B.n635 163.367
R625 B.n635 B.n634 163.367
R626 B.n634 B.n9 163.367
R627 B.n630 B.n9 163.367
R628 B.n630 B.n629 163.367
R629 B.n629 B.n628 163.367
R630 B.n628 B.n11 163.367
R631 B.n624 B.n11 163.367
R632 B.n624 B.n623 163.367
R633 B.n623 B.n622 163.367
R634 B.n622 B.n13 163.367
R635 B.n618 B.n13 163.367
R636 B.n618 B.n617 163.367
R637 B.n617 B.n616 163.367
R638 B.n616 B.n15 163.367
R639 B.n612 B.n15 163.367
R640 B.n612 B.n611 163.367
R641 B.n611 B.n610 163.367
R642 B.n610 B.n17 163.367
R643 B.n606 B.n17 163.367
R644 B.n606 B.n605 163.367
R645 B.n605 B.n604 163.367
R646 B.n604 B.n19 163.367
R647 B.n600 B.n19 163.367
R648 B.n600 B.n599 163.367
R649 B.n599 B.n598 163.367
R650 B.n598 B.n21 163.367
R651 B.n594 B.n21 163.367
R652 B.n594 B.n593 163.367
R653 B.n593 B.n592 163.367
R654 B.n592 B.n23 163.367
R655 B.n588 B.n23 163.367
R656 B.n588 B.n587 163.367
R657 B.n239 B.n238 163.367
R658 B.n239 B.n148 163.367
R659 B.n243 B.n148 163.367
R660 B.n244 B.n243 163.367
R661 B.n245 B.n244 163.367
R662 B.n245 B.n146 163.367
R663 B.n249 B.n146 163.367
R664 B.n250 B.n249 163.367
R665 B.n251 B.n250 163.367
R666 B.n251 B.n144 163.367
R667 B.n255 B.n144 163.367
R668 B.n256 B.n255 163.367
R669 B.n257 B.n256 163.367
R670 B.n257 B.n142 163.367
R671 B.n261 B.n142 163.367
R672 B.n262 B.n261 163.367
R673 B.n263 B.n262 163.367
R674 B.n263 B.n140 163.367
R675 B.n267 B.n140 163.367
R676 B.n268 B.n267 163.367
R677 B.n269 B.n268 163.367
R678 B.n269 B.n138 163.367
R679 B.n273 B.n138 163.367
R680 B.n274 B.n273 163.367
R681 B.n275 B.n274 163.367
R682 B.n275 B.n136 163.367
R683 B.n279 B.n136 163.367
R684 B.n280 B.n279 163.367
R685 B.n281 B.n280 163.367
R686 B.n281 B.n132 163.367
R687 B.n286 B.n132 163.367
R688 B.n287 B.n286 163.367
R689 B.n288 B.n287 163.367
R690 B.n288 B.n130 163.367
R691 B.n292 B.n130 163.367
R692 B.n293 B.n292 163.367
R693 B.n294 B.n293 163.367
R694 B.n294 B.n128 163.367
R695 B.n298 B.n128 163.367
R696 B.n299 B.n298 163.367
R697 B.n299 B.n124 163.367
R698 B.n303 B.n124 163.367
R699 B.n304 B.n303 163.367
R700 B.n305 B.n304 163.367
R701 B.n305 B.n122 163.367
R702 B.n309 B.n122 163.367
R703 B.n310 B.n309 163.367
R704 B.n311 B.n310 163.367
R705 B.n311 B.n120 163.367
R706 B.n315 B.n120 163.367
R707 B.n316 B.n315 163.367
R708 B.n317 B.n316 163.367
R709 B.n317 B.n118 163.367
R710 B.n321 B.n118 163.367
R711 B.n322 B.n321 163.367
R712 B.n323 B.n322 163.367
R713 B.n323 B.n116 163.367
R714 B.n327 B.n116 163.367
R715 B.n328 B.n327 163.367
R716 B.n329 B.n328 163.367
R717 B.n329 B.n114 163.367
R718 B.n333 B.n114 163.367
R719 B.n334 B.n333 163.367
R720 B.n335 B.n334 163.367
R721 B.n335 B.n112 163.367
R722 B.n339 B.n112 163.367
R723 B.n340 B.n339 163.367
R724 B.n341 B.n340 163.367
R725 B.n341 B.n110 163.367
R726 B.n346 B.n345 163.367
R727 B.n347 B.n346 163.367
R728 B.n347 B.n108 163.367
R729 B.n351 B.n108 163.367
R730 B.n352 B.n351 163.367
R731 B.n353 B.n352 163.367
R732 B.n353 B.n106 163.367
R733 B.n357 B.n106 163.367
R734 B.n358 B.n357 163.367
R735 B.n359 B.n358 163.367
R736 B.n359 B.n104 163.367
R737 B.n363 B.n104 163.367
R738 B.n364 B.n363 163.367
R739 B.n365 B.n364 163.367
R740 B.n365 B.n102 163.367
R741 B.n369 B.n102 163.367
R742 B.n370 B.n369 163.367
R743 B.n371 B.n370 163.367
R744 B.n371 B.n100 163.367
R745 B.n375 B.n100 163.367
R746 B.n376 B.n375 163.367
R747 B.n377 B.n376 163.367
R748 B.n377 B.n98 163.367
R749 B.n381 B.n98 163.367
R750 B.n382 B.n381 163.367
R751 B.n383 B.n382 163.367
R752 B.n383 B.n96 163.367
R753 B.n387 B.n96 163.367
R754 B.n388 B.n387 163.367
R755 B.n389 B.n388 163.367
R756 B.n389 B.n94 163.367
R757 B.n393 B.n94 163.367
R758 B.n394 B.n393 163.367
R759 B.n395 B.n394 163.367
R760 B.n395 B.n92 163.367
R761 B.n399 B.n92 163.367
R762 B.n400 B.n399 163.367
R763 B.n401 B.n400 163.367
R764 B.n401 B.n90 163.367
R765 B.n405 B.n90 163.367
R766 B.n406 B.n405 163.367
R767 B.n407 B.n406 163.367
R768 B.n407 B.n88 163.367
R769 B.n411 B.n88 163.367
R770 B.n412 B.n411 163.367
R771 B.n413 B.n412 163.367
R772 B.n413 B.n86 163.367
R773 B.n417 B.n86 163.367
R774 B.n418 B.n417 163.367
R775 B.n419 B.n418 163.367
R776 B.n419 B.n84 163.367
R777 B.n423 B.n84 163.367
R778 B.n424 B.n423 163.367
R779 B.n425 B.n424 163.367
R780 B.n425 B.n82 163.367
R781 B.n429 B.n82 163.367
R782 B.n430 B.n429 163.367
R783 B.n431 B.n430 163.367
R784 B.n431 B.n80 163.367
R785 B.n435 B.n80 163.367
R786 B.n436 B.n435 163.367
R787 B.n437 B.n436 163.367
R788 B.n437 B.n78 163.367
R789 B.n441 B.n78 163.367
R790 B.n442 B.n441 163.367
R791 B.n443 B.n442 163.367
R792 B.n443 B.n76 163.367
R793 B.n447 B.n76 163.367
R794 B.n448 B.n447 163.367
R795 B.n449 B.n448 163.367
R796 B.n449 B.n74 163.367
R797 B.n453 B.n74 163.367
R798 B.n454 B.n453 163.367
R799 B.n455 B.n454 163.367
R800 B.n455 B.n72 163.367
R801 B.n459 B.n72 163.367
R802 B.n460 B.n459 163.367
R803 B.n461 B.n460 163.367
R804 B.n461 B.n70 163.367
R805 B.n465 B.n70 163.367
R806 B.n466 B.n465 163.367
R807 B.n467 B.n466 163.367
R808 B.n467 B.n68 163.367
R809 B.n471 B.n68 163.367
R810 B.n472 B.n471 163.367
R811 B.n473 B.n472 163.367
R812 B.n473 B.n66 163.367
R813 B.n477 B.n66 163.367
R814 B.n478 B.n477 163.367
R815 B.n479 B.n478 163.367
R816 B.n586 B.n25 163.367
R817 B.n582 B.n25 163.367
R818 B.n582 B.n581 163.367
R819 B.n581 B.n580 163.367
R820 B.n580 B.n27 163.367
R821 B.n576 B.n27 163.367
R822 B.n576 B.n575 163.367
R823 B.n575 B.n574 163.367
R824 B.n574 B.n29 163.367
R825 B.n570 B.n29 163.367
R826 B.n570 B.n569 163.367
R827 B.n569 B.n568 163.367
R828 B.n568 B.n31 163.367
R829 B.n564 B.n31 163.367
R830 B.n564 B.n563 163.367
R831 B.n563 B.n562 163.367
R832 B.n562 B.n33 163.367
R833 B.n558 B.n33 163.367
R834 B.n558 B.n557 163.367
R835 B.n557 B.n556 163.367
R836 B.n556 B.n35 163.367
R837 B.n552 B.n35 163.367
R838 B.n552 B.n551 163.367
R839 B.n551 B.n550 163.367
R840 B.n550 B.n37 163.367
R841 B.n546 B.n37 163.367
R842 B.n546 B.n545 163.367
R843 B.n545 B.n544 163.367
R844 B.n544 B.n39 163.367
R845 B.n539 B.n39 163.367
R846 B.n539 B.n538 163.367
R847 B.n538 B.n537 163.367
R848 B.n537 B.n43 163.367
R849 B.n533 B.n43 163.367
R850 B.n533 B.n532 163.367
R851 B.n532 B.n531 163.367
R852 B.n531 B.n45 163.367
R853 B.n527 B.n45 163.367
R854 B.n527 B.n526 163.367
R855 B.n526 B.n525 163.367
R856 B.n525 B.n47 163.367
R857 B.n521 B.n47 163.367
R858 B.n521 B.n520 163.367
R859 B.n520 B.n519 163.367
R860 B.n519 B.n52 163.367
R861 B.n515 B.n52 163.367
R862 B.n515 B.n514 163.367
R863 B.n514 B.n513 163.367
R864 B.n513 B.n54 163.367
R865 B.n509 B.n54 163.367
R866 B.n509 B.n508 163.367
R867 B.n508 B.n507 163.367
R868 B.n507 B.n56 163.367
R869 B.n503 B.n56 163.367
R870 B.n503 B.n502 163.367
R871 B.n502 B.n501 163.367
R872 B.n501 B.n58 163.367
R873 B.n497 B.n58 163.367
R874 B.n497 B.n496 163.367
R875 B.n496 B.n495 163.367
R876 B.n495 B.n60 163.367
R877 B.n491 B.n60 163.367
R878 B.n491 B.n490 163.367
R879 B.n490 B.n489 163.367
R880 B.n489 B.n62 163.367
R881 B.n485 B.n62 163.367
R882 B.n485 B.n484 163.367
R883 B.n484 B.n483 163.367
R884 B.n483 B.n64 163.367
R885 B.n125 B.t8 157.03
R886 B.n48 B.t4 157.03
R887 B.n133 B.t2 157.02
R888 B.n40 B.t10 157.02
R889 B.n126 B.t7 108.546
R890 B.n49 B.t5 108.546
R891 B.n134 B.t1 108.537
R892 B.n41 B.t11 108.537
R893 B.n127 B.n126 59.5399
R894 B.n283 B.n134 59.5399
R895 B.n541 B.n41 59.5399
R896 B.n50 B.n49 59.5399
R897 B.n126 B.n125 48.4853
R898 B.n134 B.n133 48.4853
R899 B.n41 B.n40 48.4853
R900 B.n49 B.n48 48.4853
R901 B.n585 B.n24 32.3127
R902 B.n481 B.n480 32.3127
R903 B.n344 B.n343 32.3127
R904 B.n236 B.n149 32.3127
R905 B B.n655 18.0485
R906 B.n585 B.n584 10.6151
R907 B.n584 B.n583 10.6151
R908 B.n583 B.n26 10.6151
R909 B.n579 B.n26 10.6151
R910 B.n579 B.n578 10.6151
R911 B.n578 B.n577 10.6151
R912 B.n577 B.n28 10.6151
R913 B.n573 B.n28 10.6151
R914 B.n573 B.n572 10.6151
R915 B.n572 B.n571 10.6151
R916 B.n571 B.n30 10.6151
R917 B.n567 B.n30 10.6151
R918 B.n567 B.n566 10.6151
R919 B.n566 B.n565 10.6151
R920 B.n565 B.n32 10.6151
R921 B.n561 B.n32 10.6151
R922 B.n561 B.n560 10.6151
R923 B.n560 B.n559 10.6151
R924 B.n559 B.n34 10.6151
R925 B.n555 B.n34 10.6151
R926 B.n555 B.n554 10.6151
R927 B.n554 B.n553 10.6151
R928 B.n553 B.n36 10.6151
R929 B.n549 B.n36 10.6151
R930 B.n549 B.n548 10.6151
R931 B.n548 B.n547 10.6151
R932 B.n547 B.n38 10.6151
R933 B.n543 B.n38 10.6151
R934 B.n543 B.n542 10.6151
R935 B.n540 B.n42 10.6151
R936 B.n536 B.n42 10.6151
R937 B.n536 B.n535 10.6151
R938 B.n535 B.n534 10.6151
R939 B.n534 B.n44 10.6151
R940 B.n530 B.n44 10.6151
R941 B.n530 B.n529 10.6151
R942 B.n529 B.n528 10.6151
R943 B.n528 B.n46 10.6151
R944 B.n524 B.n523 10.6151
R945 B.n523 B.n522 10.6151
R946 B.n522 B.n51 10.6151
R947 B.n518 B.n51 10.6151
R948 B.n518 B.n517 10.6151
R949 B.n517 B.n516 10.6151
R950 B.n516 B.n53 10.6151
R951 B.n512 B.n53 10.6151
R952 B.n512 B.n511 10.6151
R953 B.n511 B.n510 10.6151
R954 B.n510 B.n55 10.6151
R955 B.n506 B.n55 10.6151
R956 B.n506 B.n505 10.6151
R957 B.n505 B.n504 10.6151
R958 B.n504 B.n57 10.6151
R959 B.n500 B.n57 10.6151
R960 B.n500 B.n499 10.6151
R961 B.n499 B.n498 10.6151
R962 B.n498 B.n59 10.6151
R963 B.n494 B.n59 10.6151
R964 B.n494 B.n493 10.6151
R965 B.n493 B.n492 10.6151
R966 B.n492 B.n61 10.6151
R967 B.n488 B.n61 10.6151
R968 B.n488 B.n487 10.6151
R969 B.n487 B.n486 10.6151
R970 B.n486 B.n63 10.6151
R971 B.n482 B.n63 10.6151
R972 B.n482 B.n481 10.6151
R973 B.n344 B.n109 10.6151
R974 B.n348 B.n109 10.6151
R975 B.n349 B.n348 10.6151
R976 B.n350 B.n349 10.6151
R977 B.n350 B.n107 10.6151
R978 B.n354 B.n107 10.6151
R979 B.n355 B.n354 10.6151
R980 B.n356 B.n355 10.6151
R981 B.n356 B.n105 10.6151
R982 B.n360 B.n105 10.6151
R983 B.n361 B.n360 10.6151
R984 B.n362 B.n361 10.6151
R985 B.n362 B.n103 10.6151
R986 B.n366 B.n103 10.6151
R987 B.n367 B.n366 10.6151
R988 B.n368 B.n367 10.6151
R989 B.n368 B.n101 10.6151
R990 B.n372 B.n101 10.6151
R991 B.n373 B.n372 10.6151
R992 B.n374 B.n373 10.6151
R993 B.n374 B.n99 10.6151
R994 B.n378 B.n99 10.6151
R995 B.n379 B.n378 10.6151
R996 B.n380 B.n379 10.6151
R997 B.n380 B.n97 10.6151
R998 B.n384 B.n97 10.6151
R999 B.n385 B.n384 10.6151
R1000 B.n386 B.n385 10.6151
R1001 B.n386 B.n95 10.6151
R1002 B.n390 B.n95 10.6151
R1003 B.n391 B.n390 10.6151
R1004 B.n392 B.n391 10.6151
R1005 B.n392 B.n93 10.6151
R1006 B.n396 B.n93 10.6151
R1007 B.n397 B.n396 10.6151
R1008 B.n398 B.n397 10.6151
R1009 B.n398 B.n91 10.6151
R1010 B.n402 B.n91 10.6151
R1011 B.n403 B.n402 10.6151
R1012 B.n404 B.n403 10.6151
R1013 B.n404 B.n89 10.6151
R1014 B.n408 B.n89 10.6151
R1015 B.n409 B.n408 10.6151
R1016 B.n410 B.n409 10.6151
R1017 B.n410 B.n87 10.6151
R1018 B.n414 B.n87 10.6151
R1019 B.n415 B.n414 10.6151
R1020 B.n416 B.n415 10.6151
R1021 B.n416 B.n85 10.6151
R1022 B.n420 B.n85 10.6151
R1023 B.n421 B.n420 10.6151
R1024 B.n422 B.n421 10.6151
R1025 B.n422 B.n83 10.6151
R1026 B.n426 B.n83 10.6151
R1027 B.n427 B.n426 10.6151
R1028 B.n428 B.n427 10.6151
R1029 B.n428 B.n81 10.6151
R1030 B.n432 B.n81 10.6151
R1031 B.n433 B.n432 10.6151
R1032 B.n434 B.n433 10.6151
R1033 B.n434 B.n79 10.6151
R1034 B.n438 B.n79 10.6151
R1035 B.n439 B.n438 10.6151
R1036 B.n440 B.n439 10.6151
R1037 B.n440 B.n77 10.6151
R1038 B.n444 B.n77 10.6151
R1039 B.n445 B.n444 10.6151
R1040 B.n446 B.n445 10.6151
R1041 B.n446 B.n75 10.6151
R1042 B.n450 B.n75 10.6151
R1043 B.n451 B.n450 10.6151
R1044 B.n452 B.n451 10.6151
R1045 B.n452 B.n73 10.6151
R1046 B.n456 B.n73 10.6151
R1047 B.n457 B.n456 10.6151
R1048 B.n458 B.n457 10.6151
R1049 B.n458 B.n71 10.6151
R1050 B.n462 B.n71 10.6151
R1051 B.n463 B.n462 10.6151
R1052 B.n464 B.n463 10.6151
R1053 B.n464 B.n69 10.6151
R1054 B.n468 B.n69 10.6151
R1055 B.n469 B.n468 10.6151
R1056 B.n470 B.n469 10.6151
R1057 B.n470 B.n67 10.6151
R1058 B.n474 B.n67 10.6151
R1059 B.n475 B.n474 10.6151
R1060 B.n476 B.n475 10.6151
R1061 B.n476 B.n65 10.6151
R1062 B.n480 B.n65 10.6151
R1063 B.n240 B.n149 10.6151
R1064 B.n241 B.n240 10.6151
R1065 B.n242 B.n241 10.6151
R1066 B.n242 B.n147 10.6151
R1067 B.n246 B.n147 10.6151
R1068 B.n247 B.n246 10.6151
R1069 B.n248 B.n247 10.6151
R1070 B.n248 B.n145 10.6151
R1071 B.n252 B.n145 10.6151
R1072 B.n253 B.n252 10.6151
R1073 B.n254 B.n253 10.6151
R1074 B.n254 B.n143 10.6151
R1075 B.n258 B.n143 10.6151
R1076 B.n259 B.n258 10.6151
R1077 B.n260 B.n259 10.6151
R1078 B.n260 B.n141 10.6151
R1079 B.n264 B.n141 10.6151
R1080 B.n265 B.n264 10.6151
R1081 B.n266 B.n265 10.6151
R1082 B.n266 B.n139 10.6151
R1083 B.n270 B.n139 10.6151
R1084 B.n271 B.n270 10.6151
R1085 B.n272 B.n271 10.6151
R1086 B.n272 B.n137 10.6151
R1087 B.n276 B.n137 10.6151
R1088 B.n277 B.n276 10.6151
R1089 B.n278 B.n277 10.6151
R1090 B.n278 B.n135 10.6151
R1091 B.n282 B.n135 10.6151
R1092 B.n285 B.n284 10.6151
R1093 B.n285 B.n131 10.6151
R1094 B.n289 B.n131 10.6151
R1095 B.n290 B.n289 10.6151
R1096 B.n291 B.n290 10.6151
R1097 B.n291 B.n129 10.6151
R1098 B.n295 B.n129 10.6151
R1099 B.n296 B.n295 10.6151
R1100 B.n297 B.n296 10.6151
R1101 B.n301 B.n300 10.6151
R1102 B.n302 B.n301 10.6151
R1103 B.n302 B.n123 10.6151
R1104 B.n306 B.n123 10.6151
R1105 B.n307 B.n306 10.6151
R1106 B.n308 B.n307 10.6151
R1107 B.n308 B.n121 10.6151
R1108 B.n312 B.n121 10.6151
R1109 B.n313 B.n312 10.6151
R1110 B.n314 B.n313 10.6151
R1111 B.n314 B.n119 10.6151
R1112 B.n318 B.n119 10.6151
R1113 B.n319 B.n318 10.6151
R1114 B.n320 B.n319 10.6151
R1115 B.n320 B.n117 10.6151
R1116 B.n324 B.n117 10.6151
R1117 B.n325 B.n324 10.6151
R1118 B.n326 B.n325 10.6151
R1119 B.n326 B.n115 10.6151
R1120 B.n330 B.n115 10.6151
R1121 B.n331 B.n330 10.6151
R1122 B.n332 B.n331 10.6151
R1123 B.n332 B.n113 10.6151
R1124 B.n336 B.n113 10.6151
R1125 B.n337 B.n336 10.6151
R1126 B.n338 B.n337 10.6151
R1127 B.n338 B.n111 10.6151
R1128 B.n342 B.n111 10.6151
R1129 B.n343 B.n342 10.6151
R1130 B.n236 B.n235 10.6151
R1131 B.n235 B.n234 10.6151
R1132 B.n234 B.n151 10.6151
R1133 B.n230 B.n151 10.6151
R1134 B.n230 B.n229 10.6151
R1135 B.n229 B.n228 10.6151
R1136 B.n228 B.n153 10.6151
R1137 B.n224 B.n153 10.6151
R1138 B.n224 B.n223 10.6151
R1139 B.n223 B.n222 10.6151
R1140 B.n222 B.n155 10.6151
R1141 B.n218 B.n155 10.6151
R1142 B.n218 B.n217 10.6151
R1143 B.n217 B.n216 10.6151
R1144 B.n216 B.n157 10.6151
R1145 B.n212 B.n157 10.6151
R1146 B.n212 B.n211 10.6151
R1147 B.n211 B.n210 10.6151
R1148 B.n210 B.n159 10.6151
R1149 B.n206 B.n159 10.6151
R1150 B.n206 B.n205 10.6151
R1151 B.n205 B.n204 10.6151
R1152 B.n204 B.n161 10.6151
R1153 B.n200 B.n161 10.6151
R1154 B.n200 B.n199 10.6151
R1155 B.n199 B.n198 10.6151
R1156 B.n198 B.n163 10.6151
R1157 B.n194 B.n163 10.6151
R1158 B.n194 B.n193 10.6151
R1159 B.n193 B.n192 10.6151
R1160 B.n192 B.n165 10.6151
R1161 B.n188 B.n165 10.6151
R1162 B.n188 B.n187 10.6151
R1163 B.n187 B.n186 10.6151
R1164 B.n186 B.n167 10.6151
R1165 B.n182 B.n167 10.6151
R1166 B.n182 B.n181 10.6151
R1167 B.n181 B.n180 10.6151
R1168 B.n180 B.n169 10.6151
R1169 B.n176 B.n169 10.6151
R1170 B.n176 B.n175 10.6151
R1171 B.n175 B.n174 10.6151
R1172 B.n174 B.n171 10.6151
R1173 B.n171 B.n0 10.6151
R1174 B.n651 B.n1 10.6151
R1175 B.n651 B.n650 10.6151
R1176 B.n650 B.n649 10.6151
R1177 B.n649 B.n4 10.6151
R1178 B.n645 B.n4 10.6151
R1179 B.n645 B.n644 10.6151
R1180 B.n644 B.n643 10.6151
R1181 B.n643 B.n6 10.6151
R1182 B.n639 B.n6 10.6151
R1183 B.n639 B.n638 10.6151
R1184 B.n638 B.n637 10.6151
R1185 B.n637 B.n8 10.6151
R1186 B.n633 B.n8 10.6151
R1187 B.n633 B.n632 10.6151
R1188 B.n632 B.n631 10.6151
R1189 B.n631 B.n10 10.6151
R1190 B.n627 B.n10 10.6151
R1191 B.n627 B.n626 10.6151
R1192 B.n626 B.n625 10.6151
R1193 B.n625 B.n12 10.6151
R1194 B.n621 B.n12 10.6151
R1195 B.n621 B.n620 10.6151
R1196 B.n620 B.n619 10.6151
R1197 B.n619 B.n14 10.6151
R1198 B.n615 B.n14 10.6151
R1199 B.n615 B.n614 10.6151
R1200 B.n614 B.n613 10.6151
R1201 B.n613 B.n16 10.6151
R1202 B.n609 B.n16 10.6151
R1203 B.n609 B.n608 10.6151
R1204 B.n608 B.n607 10.6151
R1205 B.n607 B.n18 10.6151
R1206 B.n603 B.n18 10.6151
R1207 B.n603 B.n602 10.6151
R1208 B.n602 B.n601 10.6151
R1209 B.n601 B.n20 10.6151
R1210 B.n597 B.n20 10.6151
R1211 B.n597 B.n596 10.6151
R1212 B.n596 B.n595 10.6151
R1213 B.n595 B.n22 10.6151
R1214 B.n591 B.n22 10.6151
R1215 B.n591 B.n590 10.6151
R1216 B.n590 B.n589 10.6151
R1217 B.n589 B.n24 10.6151
R1218 B.n542 B.n541 9.36635
R1219 B.n524 B.n50 9.36635
R1220 B.n283 B.n282 9.36635
R1221 B.n300 B.n127 9.36635
R1222 B.n655 B.n0 2.81026
R1223 B.n655 B.n1 2.81026
R1224 B.n541 B.n540 1.24928
R1225 B.n50 B.n46 1.24928
R1226 B.n284 B.n283 1.24928
R1227 B.n297 B.n127 1.24928
C0 VN VDD2 5.8371f
C1 VDD1 B 1.41586f
C2 VDD2 w_n3470_n2600# 1.80052f
C3 VP VDD2 0.473738f
C4 VN VDD1 0.150774f
C5 w_n3470_n2600# VDD1 1.70385f
C6 VP VDD1 6.15889f
C7 VN B 1.08352f
C8 w_n3470_n2600# B 8.380651f
C9 VP B 1.83426f
C10 VN w_n3470_n2600# 6.87944f
C11 VN VP 6.42438f
C12 VP w_n3470_n2600# 7.32865f
C13 VDD2 VTAIL 6.68707f
C14 VDD1 VTAIL 6.63554f
C15 B VTAIL 3.55134f
C16 VN VTAIL 6.25216f
C17 w_n3470_n2600# VTAIL 3.29894f
C18 VP VTAIL 6.26626f
C19 VDD2 VDD1 1.55004f
C20 VDD2 B 1.49836f
C21 VDD2 VSUBS 1.547147f
C22 VDD1 VSUBS 2.124348f
C23 VTAIL VSUBS 1.088265f
C24 VN VSUBS 6.07049f
C25 VP VSUBS 3.002135f
C26 B VSUBS 4.195756f
C27 w_n3470_n2600# VSUBS 0.111887p
C28 B.n0 VSUBS 0.004865f
C29 B.n1 VSUBS 0.004865f
C30 B.n2 VSUBS 0.007693f
C31 B.n3 VSUBS 0.007693f
C32 B.n4 VSUBS 0.007693f
C33 B.n5 VSUBS 0.007693f
C34 B.n6 VSUBS 0.007693f
C35 B.n7 VSUBS 0.007693f
C36 B.n8 VSUBS 0.007693f
C37 B.n9 VSUBS 0.007693f
C38 B.n10 VSUBS 0.007693f
C39 B.n11 VSUBS 0.007693f
C40 B.n12 VSUBS 0.007693f
C41 B.n13 VSUBS 0.007693f
C42 B.n14 VSUBS 0.007693f
C43 B.n15 VSUBS 0.007693f
C44 B.n16 VSUBS 0.007693f
C45 B.n17 VSUBS 0.007693f
C46 B.n18 VSUBS 0.007693f
C47 B.n19 VSUBS 0.007693f
C48 B.n20 VSUBS 0.007693f
C49 B.n21 VSUBS 0.007693f
C50 B.n22 VSUBS 0.007693f
C51 B.n23 VSUBS 0.007693f
C52 B.n24 VSUBS 0.017617f
C53 B.n25 VSUBS 0.007693f
C54 B.n26 VSUBS 0.007693f
C55 B.n27 VSUBS 0.007693f
C56 B.n28 VSUBS 0.007693f
C57 B.n29 VSUBS 0.007693f
C58 B.n30 VSUBS 0.007693f
C59 B.n31 VSUBS 0.007693f
C60 B.n32 VSUBS 0.007693f
C61 B.n33 VSUBS 0.007693f
C62 B.n34 VSUBS 0.007693f
C63 B.n35 VSUBS 0.007693f
C64 B.n36 VSUBS 0.007693f
C65 B.n37 VSUBS 0.007693f
C66 B.n38 VSUBS 0.007693f
C67 B.n39 VSUBS 0.007693f
C68 B.t11 VSUBS 0.277658f
C69 B.t10 VSUBS 0.297887f
C70 B.t9 VSUBS 0.896466f
C71 B.n40 VSUBS 0.154785f
C72 B.n41 VSUBS 0.076485f
C73 B.n42 VSUBS 0.007693f
C74 B.n43 VSUBS 0.007693f
C75 B.n44 VSUBS 0.007693f
C76 B.n45 VSUBS 0.007693f
C77 B.n46 VSUBS 0.004299f
C78 B.n47 VSUBS 0.007693f
C79 B.t5 VSUBS 0.277655f
C80 B.t4 VSUBS 0.297884f
C81 B.t3 VSUBS 0.896466f
C82 B.n48 VSUBS 0.154788f
C83 B.n49 VSUBS 0.076487f
C84 B.n50 VSUBS 0.017824f
C85 B.n51 VSUBS 0.007693f
C86 B.n52 VSUBS 0.007693f
C87 B.n53 VSUBS 0.007693f
C88 B.n54 VSUBS 0.007693f
C89 B.n55 VSUBS 0.007693f
C90 B.n56 VSUBS 0.007693f
C91 B.n57 VSUBS 0.007693f
C92 B.n58 VSUBS 0.007693f
C93 B.n59 VSUBS 0.007693f
C94 B.n60 VSUBS 0.007693f
C95 B.n61 VSUBS 0.007693f
C96 B.n62 VSUBS 0.007693f
C97 B.n63 VSUBS 0.007693f
C98 B.n64 VSUBS 0.018133f
C99 B.n65 VSUBS 0.007693f
C100 B.n66 VSUBS 0.007693f
C101 B.n67 VSUBS 0.007693f
C102 B.n68 VSUBS 0.007693f
C103 B.n69 VSUBS 0.007693f
C104 B.n70 VSUBS 0.007693f
C105 B.n71 VSUBS 0.007693f
C106 B.n72 VSUBS 0.007693f
C107 B.n73 VSUBS 0.007693f
C108 B.n74 VSUBS 0.007693f
C109 B.n75 VSUBS 0.007693f
C110 B.n76 VSUBS 0.007693f
C111 B.n77 VSUBS 0.007693f
C112 B.n78 VSUBS 0.007693f
C113 B.n79 VSUBS 0.007693f
C114 B.n80 VSUBS 0.007693f
C115 B.n81 VSUBS 0.007693f
C116 B.n82 VSUBS 0.007693f
C117 B.n83 VSUBS 0.007693f
C118 B.n84 VSUBS 0.007693f
C119 B.n85 VSUBS 0.007693f
C120 B.n86 VSUBS 0.007693f
C121 B.n87 VSUBS 0.007693f
C122 B.n88 VSUBS 0.007693f
C123 B.n89 VSUBS 0.007693f
C124 B.n90 VSUBS 0.007693f
C125 B.n91 VSUBS 0.007693f
C126 B.n92 VSUBS 0.007693f
C127 B.n93 VSUBS 0.007693f
C128 B.n94 VSUBS 0.007693f
C129 B.n95 VSUBS 0.007693f
C130 B.n96 VSUBS 0.007693f
C131 B.n97 VSUBS 0.007693f
C132 B.n98 VSUBS 0.007693f
C133 B.n99 VSUBS 0.007693f
C134 B.n100 VSUBS 0.007693f
C135 B.n101 VSUBS 0.007693f
C136 B.n102 VSUBS 0.007693f
C137 B.n103 VSUBS 0.007693f
C138 B.n104 VSUBS 0.007693f
C139 B.n105 VSUBS 0.007693f
C140 B.n106 VSUBS 0.007693f
C141 B.n107 VSUBS 0.007693f
C142 B.n108 VSUBS 0.007693f
C143 B.n109 VSUBS 0.007693f
C144 B.n110 VSUBS 0.018133f
C145 B.n111 VSUBS 0.007693f
C146 B.n112 VSUBS 0.007693f
C147 B.n113 VSUBS 0.007693f
C148 B.n114 VSUBS 0.007693f
C149 B.n115 VSUBS 0.007693f
C150 B.n116 VSUBS 0.007693f
C151 B.n117 VSUBS 0.007693f
C152 B.n118 VSUBS 0.007693f
C153 B.n119 VSUBS 0.007693f
C154 B.n120 VSUBS 0.007693f
C155 B.n121 VSUBS 0.007693f
C156 B.n122 VSUBS 0.007693f
C157 B.n123 VSUBS 0.007693f
C158 B.n124 VSUBS 0.007693f
C159 B.t7 VSUBS 0.277655f
C160 B.t8 VSUBS 0.297884f
C161 B.t6 VSUBS 0.896466f
C162 B.n125 VSUBS 0.154788f
C163 B.n126 VSUBS 0.076487f
C164 B.n127 VSUBS 0.017824f
C165 B.n128 VSUBS 0.007693f
C166 B.n129 VSUBS 0.007693f
C167 B.n130 VSUBS 0.007693f
C168 B.n131 VSUBS 0.007693f
C169 B.n132 VSUBS 0.007693f
C170 B.t1 VSUBS 0.277658f
C171 B.t2 VSUBS 0.297887f
C172 B.t0 VSUBS 0.896466f
C173 B.n133 VSUBS 0.154785f
C174 B.n134 VSUBS 0.076485f
C175 B.n135 VSUBS 0.007693f
C176 B.n136 VSUBS 0.007693f
C177 B.n137 VSUBS 0.007693f
C178 B.n138 VSUBS 0.007693f
C179 B.n139 VSUBS 0.007693f
C180 B.n140 VSUBS 0.007693f
C181 B.n141 VSUBS 0.007693f
C182 B.n142 VSUBS 0.007693f
C183 B.n143 VSUBS 0.007693f
C184 B.n144 VSUBS 0.007693f
C185 B.n145 VSUBS 0.007693f
C186 B.n146 VSUBS 0.007693f
C187 B.n147 VSUBS 0.007693f
C188 B.n148 VSUBS 0.007693f
C189 B.n149 VSUBS 0.018133f
C190 B.n150 VSUBS 0.007693f
C191 B.n151 VSUBS 0.007693f
C192 B.n152 VSUBS 0.007693f
C193 B.n153 VSUBS 0.007693f
C194 B.n154 VSUBS 0.007693f
C195 B.n155 VSUBS 0.007693f
C196 B.n156 VSUBS 0.007693f
C197 B.n157 VSUBS 0.007693f
C198 B.n158 VSUBS 0.007693f
C199 B.n159 VSUBS 0.007693f
C200 B.n160 VSUBS 0.007693f
C201 B.n161 VSUBS 0.007693f
C202 B.n162 VSUBS 0.007693f
C203 B.n163 VSUBS 0.007693f
C204 B.n164 VSUBS 0.007693f
C205 B.n165 VSUBS 0.007693f
C206 B.n166 VSUBS 0.007693f
C207 B.n167 VSUBS 0.007693f
C208 B.n168 VSUBS 0.007693f
C209 B.n169 VSUBS 0.007693f
C210 B.n170 VSUBS 0.007693f
C211 B.n171 VSUBS 0.007693f
C212 B.n172 VSUBS 0.007693f
C213 B.n173 VSUBS 0.007693f
C214 B.n174 VSUBS 0.007693f
C215 B.n175 VSUBS 0.007693f
C216 B.n176 VSUBS 0.007693f
C217 B.n177 VSUBS 0.007693f
C218 B.n178 VSUBS 0.007693f
C219 B.n179 VSUBS 0.007693f
C220 B.n180 VSUBS 0.007693f
C221 B.n181 VSUBS 0.007693f
C222 B.n182 VSUBS 0.007693f
C223 B.n183 VSUBS 0.007693f
C224 B.n184 VSUBS 0.007693f
C225 B.n185 VSUBS 0.007693f
C226 B.n186 VSUBS 0.007693f
C227 B.n187 VSUBS 0.007693f
C228 B.n188 VSUBS 0.007693f
C229 B.n189 VSUBS 0.007693f
C230 B.n190 VSUBS 0.007693f
C231 B.n191 VSUBS 0.007693f
C232 B.n192 VSUBS 0.007693f
C233 B.n193 VSUBS 0.007693f
C234 B.n194 VSUBS 0.007693f
C235 B.n195 VSUBS 0.007693f
C236 B.n196 VSUBS 0.007693f
C237 B.n197 VSUBS 0.007693f
C238 B.n198 VSUBS 0.007693f
C239 B.n199 VSUBS 0.007693f
C240 B.n200 VSUBS 0.007693f
C241 B.n201 VSUBS 0.007693f
C242 B.n202 VSUBS 0.007693f
C243 B.n203 VSUBS 0.007693f
C244 B.n204 VSUBS 0.007693f
C245 B.n205 VSUBS 0.007693f
C246 B.n206 VSUBS 0.007693f
C247 B.n207 VSUBS 0.007693f
C248 B.n208 VSUBS 0.007693f
C249 B.n209 VSUBS 0.007693f
C250 B.n210 VSUBS 0.007693f
C251 B.n211 VSUBS 0.007693f
C252 B.n212 VSUBS 0.007693f
C253 B.n213 VSUBS 0.007693f
C254 B.n214 VSUBS 0.007693f
C255 B.n215 VSUBS 0.007693f
C256 B.n216 VSUBS 0.007693f
C257 B.n217 VSUBS 0.007693f
C258 B.n218 VSUBS 0.007693f
C259 B.n219 VSUBS 0.007693f
C260 B.n220 VSUBS 0.007693f
C261 B.n221 VSUBS 0.007693f
C262 B.n222 VSUBS 0.007693f
C263 B.n223 VSUBS 0.007693f
C264 B.n224 VSUBS 0.007693f
C265 B.n225 VSUBS 0.007693f
C266 B.n226 VSUBS 0.007693f
C267 B.n227 VSUBS 0.007693f
C268 B.n228 VSUBS 0.007693f
C269 B.n229 VSUBS 0.007693f
C270 B.n230 VSUBS 0.007693f
C271 B.n231 VSUBS 0.007693f
C272 B.n232 VSUBS 0.007693f
C273 B.n233 VSUBS 0.007693f
C274 B.n234 VSUBS 0.007693f
C275 B.n235 VSUBS 0.007693f
C276 B.n236 VSUBS 0.017617f
C277 B.n237 VSUBS 0.017617f
C278 B.n238 VSUBS 0.018133f
C279 B.n239 VSUBS 0.007693f
C280 B.n240 VSUBS 0.007693f
C281 B.n241 VSUBS 0.007693f
C282 B.n242 VSUBS 0.007693f
C283 B.n243 VSUBS 0.007693f
C284 B.n244 VSUBS 0.007693f
C285 B.n245 VSUBS 0.007693f
C286 B.n246 VSUBS 0.007693f
C287 B.n247 VSUBS 0.007693f
C288 B.n248 VSUBS 0.007693f
C289 B.n249 VSUBS 0.007693f
C290 B.n250 VSUBS 0.007693f
C291 B.n251 VSUBS 0.007693f
C292 B.n252 VSUBS 0.007693f
C293 B.n253 VSUBS 0.007693f
C294 B.n254 VSUBS 0.007693f
C295 B.n255 VSUBS 0.007693f
C296 B.n256 VSUBS 0.007693f
C297 B.n257 VSUBS 0.007693f
C298 B.n258 VSUBS 0.007693f
C299 B.n259 VSUBS 0.007693f
C300 B.n260 VSUBS 0.007693f
C301 B.n261 VSUBS 0.007693f
C302 B.n262 VSUBS 0.007693f
C303 B.n263 VSUBS 0.007693f
C304 B.n264 VSUBS 0.007693f
C305 B.n265 VSUBS 0.007693f
C306 B.n266 VSUBS 0.007693f
C307 B.n267 VSUBS 0.007693f
C308 B.n268 VSUBS 0.007693f
C309 B.n269 VSUBS 0.007693f
C310 B.n270 VSUBS 0.007693f
C311 B.n271 VSUBS 0.007693f
C312 B.n272 VSUBS 0.007693f
C313 B.n273 VSUBS 0.007693f
C314 B.n274 VSUBS 0.007693f
C315 B.n275 VSUBS 0.007693f
C316 B.n276 VSUBS 0.007693f
C317 B.n277 VSUBS 0.007693f
C318 B.n278 VSUBS 0.007693f
C319 B.n279 VSUBS 0.007693f
C320 B.n280 VSUBS 0.007693f
C321 B.n281 VSUBS 0.007693f
C322 B.n282 VSUBS 0.00724f
C323 B.n283 VSUBS 0.017824f
C324 B.n284 VSUBS 0.004299f
C325 B.n285 VSUBS 0.007693f
C326 B.n286 VSUBS 0.007693f
C327 B.n287 VSUBS 0.007693f
C328 B.n288 VSUBS 0.007693f
C329 B.n289 VSUBS 0.007693f
C330 B.n290 VSUBS 0.007693f
C331 B.n291 VSUBS 0.007693f
C332 B.n292 VSUBS 0.007693f
C333 B.n293 VSUBS 0.007693f
C334 B.n294 VSUBS 0.007693f
C335 B.n295 VSUBS 0.007693f
C336 B.n296 VSUBS 0.007693f
C337 B.n297 VSUBS 0.004299f
C338 B.n298 VSUBS 0.007693f
C339 B.n299 VSUBS 0.007693f
C340 B.n300 VSUBS 0.00724f
C341 B.n301 VSUBS 0.007693f
C342 B.n302 VSUBS 0.007693f
C343 B.n303 VSUBS 0.007693f
C344 B.n304 VSUBS 0.007693f
C345 B.n305 VSUBS 0.007693f
C346 B.n306 VSUBS 0.007693f
C347 B.n307 VSUBS 0.007693f
C348 B.n308 VSUBS 0.007693f
C349 B.n309 VSUBS 0.007693f
C350 B.n310 VSUBS 0.007693f
C351 B.n311 VSUBS 0.007693f
C352 B.n312 VSUBS 0.007693f
C353 B.n313 VSUBS 0.007693f
C354 B.n314 VSUBS 0.007693f
C355 B.n315 VSUBS 0.007693f
C356 B.n316 VSUBS 0.007693f
C357 B.n317 VSUBS 0.007693f
C358 B.n318 VSUBS 0.007693f
C359 B.n319 VSUBS 0.007693f
C360 B.n320 VSUBS 0.007693f
C361 B.n321 VSUBS 0.007693f
C362 B.n322 VSUBS 0.007693f
C363 B.n323 VSUBS 0.007693f
C364 B.n324 VSUBS 0.007693f
C365 B.n325 VSUBS 0.007693f
C366 B.n326 VSUBS 0.007693f
C367 B.n327 VSUBS 0.007693f
C368 B.n328 VSUBS 0.007693f
C369 B.n329 VSUBS 0.007693f
C370 B.n330 VSUBS 0.007693f
C371 B.n331 VSUBS 0.007693f
C372 B.n332 VSUBS 0.007693f
C373 B.n333 VSUBS 0.007693f
C374 B.n334 VSUBS 0.007693f
C375 B.n335 VSUBS 0.007693f
C376 B.n336 VSUBS 0.007693f
C377 B.n337 VSUBS 0.007693f
C378 B.n338 VSUBS 0.007693f
C379 B.n339 VSUBS 0.007693f
C380 B.n340 VSUBS 0.007693f
C381 B.n341 VSUBS 0.007693f
C382 B.n342 VSUBS 0.007693f
C383 B.n343 VSUBS 0.018133f
C384 B.n344 VSUBS 0.017617f
C385 B.n345 VSUBS 0.017617f
C386 B.n346 VSUBS 0.007693f
C387 B.n347 VSUBS 0.007693f
C388 B.n348 VSUBS 0.007693f
C389 B.n349 VSUBS 0.007693f
C390 B.n350 VSUBS 0.007693f
C391 B.n351 VSUBS 0.007693f
C392 B.n352 VSUBS 0.007693f
C393 B.n353 VSUBS 0.007693f
C394 B.n354 VSUBS 0.007693f
C395 B.n355 VSUBS 0.007693f
C396 B.n356 VSUBS 0.007693f
C397 B.n357 VSUBS 0.007693f
C398 B.n358 VSUBS 0.007693f
C399 B.n359 VSUBS 0.007693f
C400 B.n360 VSUBS 0.007693f
C401 B.n361 VSUBS 0.007693f
C402 B.n362 VSUBS 0.007693f
C403 B.n363 VSUBS 0.007693f
C404 B.n364 VSUBS 0.007693f
C405 B.n365 VSUBS 0.007693f
C406 B.n366 VSUBS 0.007693f
C407 B.n367 VSUBS 0.007693f
C408 B.n368 VSUBS 0.007693f
C409 B.n369 VSUBS 0.007693f
C410 B.n370 VSUBS 0.007693f
C411 B.n371 VSUBS 0.007693f
C412 B.n372 VSUBS 0.007693f
C413 B.n373 VSUBS 0.007693f
C414 B.n374 VSUBS 0.007693f
C415 B.n375 VSUBS 0.007693f
C416 B.n376 VSUBS 0.007693f
C417 B.n377 VSUBS 0.007693f
C418 B.n378 VSUBS 0.007693f
C419 B.n379 VSUBS 0.007693f
C420 B.n380 VSUBS 0.007693f
C421 B.n381 VSUBS 0.007693f
C422 B.n382 VSUBS 0.007693f
C423 B.n383 VSUBS 0.007693f
C424 B.n384 VSUBS 0.007693f
C425 B.n385 VSUBS 0.007693f
C426 B.n386 VSUBS 0.007693f
C427 B.n387 VSUBS 0.007693f
C428 B.n388 VSUBS 0.007693f
C429 B.n389 VSUBS 0.007693f
C430 B.n390 VSUBS 0.007693f
C431 B.n391 VSUBS 0.007693f
C432 B.n392 VSUBS 0.007693f
C433 B.n393 VSUBS 0.007693f
C434 B.n394 VSUBS 0.007693f
C435 B.n395 VSUBS 0.007693f
C436 B.n396 VSUBS 0.007693f
C437 B.n397 VSUBS 0.007693f
C438 B.n398 VSUBS 0.007693f
C439 B.n399 VSUBS 0.007693f
C440 B.n400 VSUBS 0.007693f
C441 B.n401 VSUBS 0.007693f
C442 B.n402 VSUBS 0.007693f
C443 B.n403 VSUBS 0.007693f
C444 B.n404 VSUBS 0.007693f
C445 B.n405 VSUBS 0.007693f
C446 B.n406 VSUBS 0.007693f
C447 B.n407 VSUBS 0.007693f
C448 B.n408 VSUBS 0.007693f
C449 B.n409 VSUBS 0.007693f
C450 B.n410 VSUBS 0.007693f
C451 B.n411 VSUBS 0.007693f
C452 B.n412 VSUBS 0.007693f
C453 B.n413 VSUBS 0.007693f
C454 B.n414 VSUBS 0.007693f
C455 B.n415 VSUBS 0.007693f
C456 B.n416 VSUBS 0.007693f
C457 B.n417 VSUBS 0.007693f
C458 B.n418 VSUBS 0.007693f
C459 B.n419 VSUBS 0.007693f
C460 B.n420 VSUBS 0.007693f
C461 B.n421 VSUBS 0.007693f
C462 B.n422 VSUBS 0.007693f
C463 B.n423 VSUBS 0.007693f
C464 B.n424 VSUBS 0.007693f
C465 B.n425 VSUBS 0.007693f
C466 B.n426 VSUBS 0.007693f
C467 B.n427 VSUBS 0.007693f
C468 B.n428 VSUBS 0.007693f
C469 B.n429 VSUBS 0.007693f
C470 B.n430 VSUBS 0.007693f
C471 B.n431 VSUBS 0.007693f
C472 B.n432 VSUBS 0.007693f
C473 B.n433 VSUBS 0.007693f
C474 B.n434 VSUBS 0.007693f
C475 B.n435 VSUBS 0.007693f
C476 B.n436 VSUBS 0.007693f
C477 B.n437 VSUBS 0.007693f
C478 B.n438 VSUBS 0.007693f
C479 B.n439 VSUBS 0.007693f
C480 B.n440 VSUBS 0.007693f
C481 B.n441 VSUBS 0.007693f
C482 B.n442 VSUBS 0.007693f
C483 B.n443 VSUBS 0.007693f
C484 B.n444 VSUBS 0.007693f
C485 B.n445 VSUBS 0.007693f
C486 B.n446 VSUBS 0.007693f
C487 B.n447 VSUBS 0.007693f
C488 B.n448 VSUBS 0.007693f
C489 B.n449 VSUBS 0.007693f
C490 B.n450 VSUBS 0.007693f
C491 B.n451 VSUBS 0.007693f
C492 B.n452 VSUBS 0.007693f
C493 B.n453 VSUBS 0.007693f
C494 B.n454 VSUBS 0.007693f
C495 B.n455 VSUBS 0.007693f
C496 B.n456 VSUBS 0.007693f
C497 B.n457 VSUBS 0.007693f
C498 B.n458 VSUBS 0.007693f
C499 B.n459 VSUBS 0.007693f
C500 B.n460 VSUBS 0.007693f
C501 B.n461 VSUBS 0.007693f
C502 B.n462 VSUBS 0.007693f
C503 B.n463 VSUBS 0.007693f
C504 B.n464 VSUBS 0.007693f
C505 B.n465 VSUBS 0.007693f
C506 B.n466 VSUBS 0.007693f
C507 B.n467 VSUBS 0.007693f
C508 B.n468 VSUBS 0.007693f
C509 B.n469 VSUBS 0.007693f
C510 B.n470 VSUBS 0.007693f
C511 B.n471 VSUBS 0.007693f
C512 B.n472 VSUBS 0.007693f
C513 B.n473 VSUBS 0.007693f
C514 B.n474 VSUBS 0.007693f
C515 B.n475 VSUBS 0.007693f
C516 B.n476 VSUBS 0.007693f
C517 B.n477 VSUBS 0.007693f
C518 B.n478 VSUBS 0.007693f
C519 B.n479 VSUBS 0.017617f
C520 B.n480 VSUBS 0.018536f
C521 B.n481 VSUBS 0.017214f
C522 B.n482 VSUBS 0.007693f
C523 B.n483 VSUBS 0.007693f
C524 B.n484 VSUBS 0.007693f
C525 B.n485 VSUBS 0.007693f
C526 B.n486 VSUBS 0.007693f
C527 B.n487 VSUBS 0.007693f
C528 B.n488 VSUBS 0.007693f
C529 B.n489 VSUBS 0.007693f
C530 B.n490 VSUBS 0.007693f
C531 B.n491 VSUBS 0.007693f
C532 B.n492 VSUBS 0.007693f
C533 B.n493 VSUBS 0.007693f
C534 B.n494 VSUBS 0.007693f
C535 B.n495 VSUBS 0.007693f
C536 B.n496 VSUBS 0.007693f
C537 B.n497 VSUBS 0.007693f
C538 B.n498 VSUBS 0.007693f
C539 B.n499 VSUBS 0.007693f
C540 B.n500 VSUBS 0.007693f
C541 B.n501 VSUBS 0.007693f
C542 B.n502 VSUBS 0.007693f
C543 B.n503 VSUBS 0.007693f
C544 B.n504 VSUBS 0.007693f
C545 B.n505 VSUBS 0.007693f
C546 B.n506 VSUBS 0.007693f
C547 B.n507 VSUBS 0.007693f
C548 B.n508 VSUBS 0.007693f
C549 B.n509 VSUBS 0.007693f
C550 B.n510 VSUBS 0.007693f
C551 B.n511 VSUBS 0.007693f
C552 B.n512 VSUBS 0.007693f
C553 B.n513 VSUBS 0.007693f
C554 B.n514 VSUBS 0.007693f
C555 B.n515 VSUBS 0.007693f
C556 B.n516 VSUBS 0.007693f
C557 B.n517 VSUBS 0.007693f
C558 B.n518 VSUBS 0.007693f
C559 B.n519 VSUBS 0.007693f
C560 B.n520 VSUBS 0.007693f
C561 B.n521 VSUBS 0.007693f
C562 B.n522 VSUBS 0.007693f
C563 B.n523 VSUBS 0.007693f
C564 B.n524 VSUBS 0.00724f
C565 B.n525 VSUBS 0.007693f
C566 B.n526 VSUBS 0.007693f
C567 B.n527 VSUBS 0.007693f
C568 B.n528 VSUBS 0.007693f
C569 B.n529 VSUBS 0.007693f
C570 B.n530 VSUBS 0.007693f
C571 B.n531 VSUBS 0.007693f
C572 B.n532 VSUBS 0.007693f
C573 B.n533 VSUBS 0.007693f
C574 B.n534 VSUBS 0.007693f
C575 B.n535 VSUBS 0.007693f
C576 B.n536 VSUBS 0.007693f
C577 B.n537 VSUBS 0.007693f
C578 B.n538 VSUBS 0.007693f
C579 B.n539 VSUBS 0.007693f
C580 B.n540 VSUBS 0.004299f
C581 B.n541 VSUBS 0.017824f
C582 B.n542 VSUBS 0.00724f
C583 B.n543 VSUBS 0.007693f
C584 B.n544 VSUBS 0.007693f
C585 B.n545 VSUBS 0.007693f
C586 B.n546 VSUBS 0.007693f
C587 B.n547 VSUBS 0.007693f
C588 B.n548 VSUBS 0.007693f
C589 B.n549 VSUBS 0.007693f
C590 B.n550 VSUBS 0.007693f
C591 B.n551 VSUBS 0.007693f
C592 B.n552 VSUBS 0.007693f
C593 B.n553 VSUBS 0.007693f
C594 B.n554 VSUBS 0.007693f
C595 B.n555 VSUBS 0.007693f
C596 B.n556 VSUBS 0.007693f
C597 B.n557 VSUBS 0.007693f
C598 B.n558 VSUBS 0.007693f
C599 B.n559 VSUBS 0.007693f
C600 B.n560 VSUBS 0.007693f
C601 B.n561 VSUBS 0.007693f
C602 B.n562 VSUBS 0.007693f
C603 B.n563 VSUBS 0.007693f
C604 B.n564 VSUBS 0.007693f
C605 B.n565 VSUBS 0.007693f
C606 B.n566 VSUBS 0.007693f
C607 B.n567 VSUBS 0.007693f
C608 B.n568 VSUBS 0.007693f
C609 B.n569 VSUBS 0.007693f
C610 B.n570 VSUBS 0.007693f
C611 B.n571 VSUBS 0.007693f
C612 B.n572 VSUBS 0.007693f
C613 B.n573 VSUBS 0.007693f
C614 B.n574 VSUBS 0.007693f
C615 B.n575 VSUBS 0.007693f
C616 B.n576 VSUBS 0.007693f
C617 B.n577 VSUBS 0.007693f
C618 B.n578 VSUBS 0.007693f
C619 B.n579 VSUBS 0.007693f
C620 B.n580 VSUBS 0.007693f
C621 B.n581 VSUBS 0.007693f
C622 B.n582 VSUBS 0.007693f
C623 B.n583 VSUBS 0.007693f
C624 B.n584 VSUBS 0.007693f
C625 B.n585 VSUBS 0.018133f
C626 B.n586 VSUBS 0.018133f
C627 B.n587 VSUBS 0.017617f
C628 B.n588 VSUBS 0.007693f
C629 B.n589 VSUBS 0.007693f
C630 B.n590 VSUBS 0.007693f
C631 B.n591 VSUBS 0.007693f
C632 B.n592 VSUBS 0.007693f
C633 B.n593 VSUBS 0.007693f
C634 B.n594 VSUBS 0.007693f
C635 B.n595 VSUBS 0.007693f
C636 B.n596 VSUBS 0.007693f
C637 B.n597 VSUBS 0.007693f
C638 B.n598 VSUBS 0.007693f
C639 B.n599 VSUBS 0.007693f
C640 B.n600 VSUBS 0.007693f
C641 B.n601 VSUBS 0.007693f
C642 B.n602 VSUBS 0.007693f
C643 B.n603 VSUBS 0.007693f
C644 B.n604 VSUBS 0.007693f
C645 B.n605 VSUBS 0.007693f
C646 B.n606 VSUBS 0.007693f
C647 B.n607 VSUBS 0.007693f
C648 B.n608 VSUBS 0.007693f
C649 B.n609 VSUBS 0.007693f
C650 B.n610 VSUBS 0.007693f
C651 B.n611 VSUBS 0.007693f
C652 B.n612 VSUBS 0.007693f
C653 B.n613 VSUBS 0.007693f
C654 B.n614 VSUBS 0.007693f
C655 B.n615 VSUBS 0.007693f
C656 B.n616 VSUBS 0.007693f
C657 B.n617 VSUBS 0.007693f
C658 B.n618 VSUBS 0.007693f
C659 B.n619 VSUBS 0.007693f
C660 B.n620 VSUBS 0.007693f
C661 B.n621 VSUBS 0.007693f
C662 B.n622 VSUBS 0.007693f
C663 B.n623 VSUBS 0.007693f
C664 B.n624 VSUBS 0.007693f
C665 B.n625 VSUBS 0.007693f
C666 B.n626 VSUBS 0.007693f
C667 B.n627 VSUBS 0.007693f
C668 B.n628 VSUBS 0.007693f
C669 B.n629 VSUBS 0.007693f
C670 B.n630 VSUBS 0.007693f
C671 B.n631 VSUBS 0.007693f
C672 B.n632 VSUBS 0.007693f
C673 B.n633 VSUBS 0.007693f
C674 B.n634 VSUBS 0.007693f
C675 B.n635 VSUBS 0.007693f
C676 B.n636 VSUBS 0.007693f
C677 B.n637 VSUBS 0.007693f
C678 B.n638 VSUBS 0.007693f
C679 B.n639 VSUBS 0.007693f
C680 B.n640 VSUBS 0.007693f
C681 B.n641 VSUBS 0.007693f
C682 B.n642 VSUBS 0.007693f
C683 B.n643 VSUBS 0.007693f
C684 B.n644 VSUBS 0.007693f
C685 B.n645 VSUBS 0.007693f
C686 B.n646 VSUBS 0.007693f
C687 B.n647 VSUBS 0.007693f
C688 B.n648 VSUBS 0.007693f
C689 B.n649 VSUBS 0.007693f
C690 B.n650 VSUBS 0.007693f
C691 B.n651 VSUBS 0.007693f
C692 B.n652 VSUBS 0.007693f
C693 B.n653 VSUBS 0.007693f
C694 B.n654 VSUBS 0.007693f
C695 B.n655 VSUBS 0.01742f
C696 VDD2.t2 VSUBS 0.157271f
C697 VDD2.t5 VSUBS 0.157271f
C698 VDD2.n0 VSUBS 1.14762f
C699 VDD2.t1 VSUBS 0.157271f
C700 VDD2.t6 VSUBS 0.157271f
C701 VDD2.n1 VSUBS 1.14762f
C702 VDD2.n2 VSUBS 3.1586f
C703 VDD2.t7 VSUBS 0.157271f
C704 VDD2.t3 VSUBS 0.157271f
C705 VDD2.n3 VSUBS 1.13918f
C706 VDD2.n4 VSUBS 2.66162f
C707 VDD2.t0 VSUBS 0.157271f
C708 VDD2.t4 VSUBS 0.157271f
C709 VDD2.n5 VSUBS 1.14758f
C710 VN.n0 VSUBS 0.046955f
C711 VN.t1 VSUBS 1.69525f
C712 VN.n1 VSUBS 0.028767f
C713 VN.n2 VSUBS 0.035617f
C714 VN.t6 VSUBS 1.69525f
C715 VN.n3 VSUBS 0.070416f
C716 VN.n4 VSUBS 0.035617f
C717 VN.t2 VSUBS 1.69525f
C718 VN.n5 VSUBS 0.712342f
C719 VN.t5 VSUBS 1.90647f
C720 VN.n6 VSUBS 0.702729f
C721 VN.n7 VSUBS 0.301855f
C722 VN.n8 VSUBS 0.049745f
C723 VN.n9 VSUBS 0.070416f
C724 VN.n10 VSUBS 0.028767f
C725 VN.n11 VSUBS 0.035617f
C726 VN.n12 VSUBS 0.035617f
C727 VN.n13 VSUBS 0.035617f
C728 VN.n14 VSUBS 0.049745f
C729 VN.n15 VSUBS 0.621757f
C730 VN.n16 VSUBS 0.049745f
C731 VN.n17 VSUBS 0.070416f
C732 VN.n18 VSUBS 0.035617f
C733 VN.n19 VSUBS 0.035617f
C734 VN.n20 VSUBS 0.035617f
C735 VN.n21 VSUBS 0.070416f
C736 VN.n22 VSUBS 0.049745f
C737 VN.n23 VSUBS 0.723884f
C738 VN.n24 VSUBS 0.051464f
C739 VN.n25 VSUBS 0.046955f
C740 VN.t0 VSUBS 1.69525f
C741 VN.n26 VSUBS 0.028767f
C742 VN.n27 VSUBS 0.035617f
C743 VN.t4 VSUBS 1.69525f
C744 VN.n28 VSUBS 0.070416f
C745 VN.n29 VSUBS 0.035617f
C746 VN.t7 VSUBS 1.69525f
C747 VN.n30 VSUBS 0.712342f
C748 VN.t3 VSUBS 1.90647f
C749 VN.n31 VSUBS 0.702729f
C750 VN.n32 VSUBS 0.301855f
C751 VN.n33 VSUBS 0.049745f
C752 VN.n34 VSUBS 0.070416f
C753 VN.n35 VSUBS 0.028767f
C754 VN.n36 VSUBS 0.035617f
C755 VN.n37 VSUBS 0.035617f
C756 VN.n38 VSUBS 0.035617f
C757 VN.n39 VSUBS 0.049745f
C758 VN.n40 VSUBS 0.621757f
C759 VN.n41 VSUBS 0.049745f
C760 VN.n42 VSUBS 0.070416f
C761 VN.n43 VSUBS 0.035617f
C762 VN.n44 VSUBS 0.035617f
C763 VN.n45 VSUBS 0.035617f
C764 VN.n46 VSUBS 0.070416f
C765 VN.n47 VSUBS 0.049745f
C766 VN.n48 VSUBS 0.723884f
C767 VN.n49 VSUBS 1.75553f
C768 VTAIL.t0 VSUBS 0.171574f
C769 VTAIL.t6 VSUBS 0.171574f
C770 VTAIL.n0 VSUBS 1.12599f
C771 VTAIL.n1 VSUBS 0.727872f
C772 VTAIL.t3 VSUBS 1.51131f
C773 VTAIL.n2 VSUBS 0.845774f
C774 VTAIL.t8 VSUBS 1.51131f
C775 VTAIL.n3 VSUBS 0.845774f
C776 VTAIL.t9 VSUBS 0.171574f
C777 VTAIL.t12 VSUBS 0.171574f
C778 VTAIL.n4 VSUBS 1.12599f
C779 VTAIL.n5 VSUBS 0.90766f
C780 VTAIL.t13 VSUBS 1.51131f
C781 VTAIL.n6 VSUBS 1.95481f
C782 VTAIL.t4 VSUBS 1.51132f
C783 VTAIL.n7 VSUBS 1.9548f
C784 VTAIL.t2 VSUBS 0.171574f
C785 VTAIL.t7 VSUBS 0.171574f
C786 VTAIL.n8 VSUBS 1.12599f
C787 VTAIL.n9 VSUBS 0.907655f
C788 VTAIL.t1 VSUBS 1.51132f
C789 VTAIL.n10 VSUBS 0.845763f
C790 VTAIL.t14 VSUBS 1.51132f
C791 VTAIL.n11 VSUBS 0.845763f
C792 VTAIL.t10 VSUBS 0.171574f
C793 VTAIL.t15 VSUBS 0.171574f
C794 VTAIL.n12 VSUBS 1.12599f
C795 VTAIL.n13 VSUBS 0.907655f
C796 VTAIL.t11 VSUBS 1.51131f
C797 VTAIL.n14 VSUBS 1.95481f
C798 VTAIL.t5 VSUBS 1.51131f
C799 VTAIL.n15 VSUBS 1.94982f
C800 VDD1.t3 VSUBS 0.159893f
C801 VDD1.t5 VSUBS 0.159893f
C802 VDD1.n0 VSUBS 1.16781f
C803 VDD1.t1 VSUBS 0.159893f
C804 VDD1.t4 VSUBS 0.159893f
C805 VDD1.n1 VSUBS 1.16675f
C806 VDD1.t0 VSUBS 0.159893f
C807 VDD1.t7 VSUBS 0.159893f
C808 VDD1.n2 VSUBS 1.16675f
C809 VDD1.n3 VSUBS 3.26329f
C810 VDD1.t2 VSUBS 0.159893f
C811 VDD1.t6 VSUBS 0.159893f
C812 VDD1.n4 VSUBS 1.15817f
C813 VDD1.n5 VSUBS 2.73626f
C814 VP.n0 VSUBS 0.048529f
C815 VP.t7 VSUBS 1.7521f
C816 VP.n1 VSUBS 0.029731f
C817 VP.n2 VSUBS 0.036811f
C818 VP.t3 VSUBS 1.7521f
C819 VP.n3 VSUBS 0.072777f
C820 VP.n4 VSUBS 0.036811f
C821 VP.t6 VSUBS 1.7521f
C822 VP.n5 VSUBS 0.642606f
C823 VP.n6 VSUBS 0.036811f
C824 VP.n7 VSUBS 0.072777f
C825 VP.n8 VSUBS 0.048529f
C826 VP.t4 VSUBS 1.7521f
C827 VP.n9 VSUBS 0.029731f
C828 VP.n10 VSUBS 0.036811f
C829 VP.t0 VSUBS 1.7521f
C830 VP.n11 VSUBS 0.072777f
C831 VP.n12 VSUBS 0.036811f
C832 VP.t5 VSUBS 1.7521f
C833 VP.n13 VSUBS 0.736229f
C834 VP.t1 VSUBS 1.97041f
C835 VP.n14 VSUBS 0.726294f
C836 VP.n15 VSUBS 0.311977f
C837 VP.n16 VSUBS 0.051413f
C838 VP.n17 VSUBS 0.072777f
C839 VP.n18 VSUBS 0.029731f
C840 VP.n19 VSUBS 0.036811f
C841 VP.n20 VSUBS 0.036811f
C842 VP.n21 VSUBS 0.036811f
C843 VP.n22 VSUBS 0.051413f
C844 VP.n23 VSUBS 0.642606f
C845 VP.n24 VSUBS 0.051413f
C846 VP.n25 VSUBS 0.072777f
C847 VP.n26 VSUBS 0.036811f
C848 VP.n27 VSUBS 0.036811f
C849 VP.n28 VSUBS 0.036811f
C850 VP.n29 VSUBS 0.072777f
C851 VP.n30 VSUBS 0.051413f
C852 VP.n31 VSUBS 0.748158f
C853 VP.n32 VSUBS 1.79434f
C854 VP.n33 VSUBS 1.82324f
C855 VP.t2 VSUBS 1.7521f
C856 VP.n34 VSUBS 0.748158f
C857 VP.n35 VSUBS 0.051413f
C858 VP.n36 VSUBS 0.048529f
C859 VP.n37 VSUBS 0.036811f
C860 VP.n38 VSUBS 0.036811f
C861 VP.n39 VSUBS 0.029731f
C862 VP.n40 VSUBS 0.072777f
C863 VP.n41 VSUBS 0.051413f
C864 VP.n42 VSUBS 0.036811f
C865 VP.n43 VSUBS 0.036811f
C866 VP.n44 VSUBS 0.051413f
C867 VP.n45 VSUBS 0.072777f
C868 VP.n46 VSUBS 0.029731f
C869 VP.n47 VSUBS 0.036811f
C870 VP.n48 VSUBS 0.036811f
C871 VP.n49 VSUBS 0.036811f
C872 VP.n50 VSUBS 0.051413f
C873 VP.n51 VSUBS 0.642606f
C874 VP.n52 VSUBS 0.051413f
C875 VP.n53 VSUBS 0.072777f
C876 VP.n54 VSUBS 0.036811f
C877 VP.n55 VSUBS 0.036811f
C878 VP.n56 VSUBS 0.036811f
C879 VP.n57 VSUBS 0.072777f
C880 VP.n58 VSUBS 0.051413f
C881 VP.n59 VSUBS 0.748158f
C882 VP.n60 VSUBS 0.05319f
.ends

