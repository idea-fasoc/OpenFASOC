* NGSPICE file created from diff_pair_sample_1092.ext - technology: sky130A

.subckt diff_pair_sample_1092 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2478_n1074# sky130_fd_pr__pfet_01v8 ad=0.2067 pd=1.84 as=0 ps=0 w=0.53 l=3.44
X1 B.t8 B.t6 B.t7 w_n2478_n1074# sky130_fd_pr__pfet_01v8 ad=0.2067 pd=1.84 as=0 ps=0 w=0.53 l=3.44
X2 VDD1.t1 VP.t0 VTAIL.t3 w_n2478_n1074# sky130_fd_pr__pfet_01v8 ad=0.2067 pd=1.84 as=0.2067 ps=1.84 w=0.53 l=3.44
X3 VDD2.t1 VN.t0 VTAIL.t0 w_n2478_n1074# sky130_fd_pr__pfet_01v8 ad=0.2067 pd=1.84 as=0.2067 ps=1.84 w=0.53 l=3.44
X4 B.t5 B.t3 B.t4 w_n2478_n1074# sky130_fd_pr__pfet_01v8 ad=0.2067 pd=1.84 as=0 ps=0 w=0.53 l=3.44
X5 B.t2 B.t0 B.t1 w_n2478_n1074# sky130_fd_pr__pfet_01v8 ad=0.2067 pd=1.84 as=0 ps=0 w=0.53 l=3.44
X6 VDD1.t0 VP.t1 VTAIL.t2 w_n2478_n1074# sky130_fd_pr__pfet_01v8 ad=0.2067 pd=1.84 as=0.2067 ps=1.84 w=0.53 l=3.44
X7 VDD2.t0 VN.t1 VTAIL.t1 w_n2478_n1074# sky130_fd_pr__pfet_01v8 ad=0.2067 pd=1.84 as=0.2067 ps=1.84 w=0.53 l=3.44
R0 B.n74 B.t7 739.422
R1 B.n162 B.t10 739.422
R2 B.n28 B.t2 739.422
R3 B.n22 B.t5 739.422
R4 B.n75 B.t8 666.307
R5 B.n163 B.t11 666.307
R6 B.n29 B.t1 666.307
R7 B.n23 B.t4 666.307
R8 B.n178 B.n177 585
R9 B.n176 B.n65 585
R10 B.n175 B.n174 585
R11 B.n173 B.n66 585
R12 B.n172 B.n171 585
R13 B.n170 B.n67 585
R14 B.n169 B.n168 585
R15 B.n167 B.n68 585
R16 B.n166 B.n165 585
R17 B.n161 B.n69 585
R18 B.n160 B.n159 585
R19 B.n158 B.n70 585
R20 B.n157 B.n156 585
R21 B.n155 B.n71 585
R22 B.n154 B.n153 585
R23 B.n152 B.n72 585
R24 B.n151 B.n150 585
R25 B.n148 B.n73 585
R26 B.n147 B.n146 585
R27 B.n145 B.n76 585
R28 B.n144 B.n143 585
R29 B.n142 B.n77 585
R30 B.n141 B.n140 585
R31 B.n139 B.n78 585
R32 B.n138 B.n137 585
R33 B.n179 B.n64 585
R34 B.n181 B.n180 585
R35 B.n182 B.n63 585
R36 B.n184 B.n183 585
R37 B.n185 B.n62 585
R38 B.n187 B.n186 585
R39 B.n188 B.n61 585
R40 B.n190 B.n189 585
R41 B.n191 B.n60 585
R42 B.n193 B.n192 585
R43 B.n194 B.n59 585
R44 B.n196 B.n195 585
R45 B.n197 B.n58 585
R46 B.n199 B.n198 585
R47 B.n200 B.n57 585
R48 B.n202 B.n201 585
R49 B.n203 B.n56 585
R50 B.n205 B.n204 585
R51 B.n206 B.n55 585
R52 B.n208 B.n207 585
R53 B.n209 B.n54 585
R54 B.n211 B.n210 585
R55 B.n212 B.n53 585
R56 B.n214 B.n213 585
R57 B.n215 B.n52 585
R58 B.n217 B.n216 585
R59 B.n218 B.n51 585
R60 B.n220 B.n219 585
R61 B.n221 B.n50 585
R62 B.n223 B.n222 585
R63 B.n224 B.n49 585
R64 B.n226 B.n225 585
R65 B.n227 B.n48 585
R66 B.n229 B.n228 585
R67 B.n230 B.n47 585
R68 B.n232 B.n231 585
R69 B.n233 B.n46 585
R70 B.n235 B.n234 585
R71 B.n236 B.n45 585
R72 B.n238 B.n237 585
R73 B.n239 B.n44 585
R74 B.n241 B.n240 585
R75 B.n242 B.n43 585
R76 B.n244 B.n243 585
R77 B.n245 B.n42 585
R78 B.n247 B.n246 585
R79 B.n248 B.n41 585
R80 B.n250 B.n249 585
R81 B.n251 B.n40 585
R82 B.n253 B.n252 585
R83 B.n254 B.n39 585
R84 B.n256 B.n255 585
R85 B.n257 B.n38 585
R86 B.n259 B.n258 585
R87 B.n260 B.n37 585
R88 B.n262 B.n261 585
R89 B.n263 B.n36 585
R90 B.n265 B.n264 585
R91 B.n266 B.n35 585
R92 B.n268 B.n267 585
R93 B.n269 B.n34 585
R94 B.n271 B.n270 585
R95 B.n310 B.n17 585
R96 B.n309 B.n308 585
R97 B.n307 B.n18 585
R98 B.n306 B.n305 585
R99 B.n304 B.n19 585
R100 B.n303 B.n302 585
R101 B.n301 B.n20 585
R102 B.n300 B.n299 585
R103 B.n297 B.n21 585
R104 B.n296 B.n295 585
R105 B.n294 B.n24 585
R106 B.n293 B.n292 585
R107 B.n291 B.n25 585
R108 B.n290 B.n289 585
R109 B.n288 B.n26 585
R110 B.n287 B.n286 585
R111 B.n285 B.n27 585
R112 B.n283 B.n282 585
R113 B.n281 B.n30 585
R114 B.n280 B.n279 585
R115 B.n278 B.n31 585
R116 B.n277 B.n276 585
R117 B.n275 B.n32 585
R118 B.n274 B.n273 585
R119 B.n272 B.n33 585
R120 B.n312 B.n311 585
R121 B.n313 B.n16 585
R122 B.n315 B.n314 585
R123 B.n316 B.n15 585
R124 B.n318 B.n317 585
R125 B.n319 B.n14 585
R126 B.n321 B.n320 585
R127 B.n322 B.n13 585
R128 B.n324 B.n323 585
R129 B.n325 B.n12 585
R130 B.n327 B.n326 585
R131 B.n328 B.n11 585
R132 B.n330 B.n329 585
R133 B.n331 B.n10 585
R134 B.n333 B.n332 585
R135 B.n334 B.n9 585
R136 B.n336 B.n335 585
R137 B.n337 B.n8 585
R138 B.n339 B.n338 585
R139 B.n340 B.n7 585
R140 B.n342 B.n341 585
R141 B.n343 B.n6 585
R142 B.n345 B.n344 585
R143 B.n346 B.n5 585
R144 B.n348 B.n347 585
R145 B.n349 B.n4 585
R146 B.n351 B.n350 585
R147 B.n352 B.n3 585
R148 B.n354 B.n353 585
R149 B.n355 B.n0 585
R150 B.n2 B.n1 585
R151 B.n94 B.n93 585
R152 B.n96 B.n95 585
R153 B.n97 B.n92 585
R154 B.n99 B.n98 585
R155 B.n100 B.n91 585
R156 B.n102 B.n101 585
R157 B.n103 B.n90 585
R158 B.n105 B.n104 585
R159 B.n106 B.n89 585
R160 B.n108 B.n107 585
R161 B.n109 B.n88 585
R162 B.n111 B.n110 585
R163 B.n112 B.n87 585
R164 B.n114 B.n113 585
R165 B.n115 B.n86 585
R166 B.n117 B.n116 585
R167 B.n118 B.n85 585
R168 B.n120 B.n119 585
R169 B.n121 B.n84 585
R170 B.n123 B.n122 585
R171 B.n124 B.n83 585
R172 B.n126 B.n125 585
R173 B.n127 B.n82 585
R174 B.n129 B.n128 585
R175 B.n130 B.n81 585
R176 B.n132 B.n131 585
R177 B.n133 B.n80 585
R178 B.n135 B.n134 585
R179 B.n136 B.n79 585
R180 B.n138 B.n79 492.5
R181 B.n179 B.n178 492.5
R182 B.n270 B.n33 492.5
R183 B.n312 B.n17 492.5
R184 B.n357 B.n356 256.663
R185 B.n356 B.n355 235.042
R186 B.n356 B.n2 235.042
R187 B.n74 B.t6 210.166
R188 B.n162 B.t9 210.166
R189 B.n28 B.t0 210.166
R190 B.n22 B.t3 210.166
R191 B.n139 B.n138 163.367
R192 B.n140 B.n139 163.367
R193 B.n140 B.n77 163.367
R194 B.n144 B.n77 163.367
R195 B.n145 B.n144 163.367
R196 B.n146 B.n145 163.367
R197 B.n146 B.n73 163.367
R198 B.n151 B.n73 163.367
R199 B.n152 B.n151 163.367
R200 B.n153 B.n152 163.367
R201 B.n153 B.n71 163.367
R202 B.n157 B.n71 163.367
R203 B.n158 B.n157 163.367
R204 B.n159 B.n158 163.367
R205 B.n159 B.n69 163.367
R206 B.n166 B.n69 163.367
R207 B.n167 B.n166 163.367
R208 B.n168 B.n167 163.367
R209 B.n168 B.n67 163.367
R210 B.n172 B.n67 163.367
R211 B.n173 B.n172 163.367
R212 B.n174 B.n173 163.367
R213 B.n174 B.n65 163.367
R214 B.n178 B.n65 163.367
R215 B.n270 B.n269 163.367
R216 B.n269 B.n268 163.367
R217 B.n268 B.n35 163.367
R218 B.n264 B.n35 163.367
R219 B.n264 B.n263 163.367
R220 B.n263 B.n262 163.367
R221 B.n262 B.n37 163.367
R222 B.n258 B.n37 163.367
R223 B.n258 B.n257 163.367
R224 B.n257 B.n256 163.367
R225 B.n256 B.n39 163.367
R226 B.n252 B.n39 163.367
R227 B.n252 B.n251 163.367
R228 B.n251 B.n250 163.367
R229 B.n250 B.n41 163.367
R230 B.n246 B.n41 163.367
R231 B.n246 B.n245 163.367
R232 B.n245 B.n244 163.367
R233 B.n244 B.n43 163.367
R234 B.n240 B.n43 163.367
R235 B.n240 B.n239 163.367
R236 B.n239 B.n238 163.367
R237 B.n238 B.n45 163.367
R238 B.n234 B.n45 163.367
R239 B.n234 B.n233 163.367
R240 B.n233 B.n232 163.367
R241 B.n232 B.n47 163.367
R242 B.n228 B.n47 163.367
R243 B.n228 B.n227 163.367
R244 B.n227 B.n226 163.367
R245 B.n226 B.n49 163.367
R246 B.n222 B.n49 163.367
R247 B.n222 B.n221 163.367
R248 B.n221 B.n220 163.367
R249 B.n220 B.n51 163.367
R250 B.n216 B.n51 163.367
R251 B.n216 B.n215 163.367
R252 B.n215 B.n214 163.367
R253 B.n214 B.n53 163.367
R254 B.n210 B.n53 163.367
R255 B.n210 B.n209 163.367
R256 B.n209 B.n208 163.367
R257 B.n208 B.n55 163.367
R258 B.n204 B.n55 163.367
R259 B.n204 B.n203 163.367
R260 B.n203 B.n202 163.367
R261 B.n202 B.n57 163.367
R262 B.n198 B.n57 163.367
R263 B.n198 B.n197 163.367
R264 B.n197 B.n196 163.367
R265 B.n196 B.n59 163.367
R266 B.n192 B.n59 163.367
R267 B.n192 B.n191 163.367
R268 B.n191 B.n190 163.367
R269 B.n190 B.n61 163.367
R270 B.n186 B.n61 163.367
R271 B.n186 B.n185 163.367
R272 B.n185 B.n184 163.367
R273 B.n184 B.n63 163.367
R274 B.n180 B.n63 163.367
R275 B.n180 B.n179 163.367
R276 B.n308 B.n17 163.367
R277 B.n308 B.n307 163.367
R278 B.n307 B.n306 163.367
R279 B.n306 B.n19 163.367
R280 B.n302 B.n19 163.367
R281 B.n302 B.n301 163.367
R282 B.n301 B.n300 163.367
R283 B.n300 B.n21 163.367
R284 B.n295 B.n21 163.367
R285 B.n295 B.n294 163.367
R286 B.n294 B.n293 163.367
R287 B.n293 B.n25 163.367
R288 B.n289 B.n25 163.367
R289 B.n289 B.n288 163.367
R290 B.n288 B.n287 163.367
R291 B.n287 B.n27 163.367
R292 B.n282 B.n27 163.367
R293 B.n282 B.n281 163.367
R294 B.n281 B.n280 163.367
R295 B.n280 B.n31 163.367
R296 B.n276 B.n31 163.367
R297 B.n276 B.n275 163.367
R298 B.n275 B.n274 163.367
R299 B.n274 B.n33 163.367
R300 B.n313 B.n312 163.367
R301 B.n314 B.n313 163.367
R302 B.n314 B.n15 163.367
R303 B.n318 B.n15 163.367
R304 B.n319 B.n318 163.367
R305 B.n320 B.n319 163.367
R306 B.n320 B.n13 163.367
R307 B.n324 B.n13 163.367
R308 B.n325 B.n324 163.367
R309 B.n326 B.n325 163.367
R310 B.n326 B.n11 163.367
R311 B.n330 B.n11 163.367
R312 B.n331 B.n330 163.367
R313 B.n332 B.n331 163.367
R314 B.n332 B.n9 163.367
R315 B.n336 B.n9 163.367
R316 B.n337 B.n336 163.367
R317 B.n338 B.n337 163.367
R318 B.n338 B.n7 163.367
R319 B.n342 B.n7 163.367
R320 B.n343 B.n342 163.367
R321 B.n344 B.n343 163.367
R322 B.n344 B.n5 163.367
R323 B.n348 B.n5 163.367
R324 B.n349 B.n348 163.367
R325 B.n350 B.n349 163.367
R326 B.n350 B.n3 163.367
R327 B.n354 B.n3 163.367
R328 B.n355 B.n354 163.367
R329 B.n93 B.n2 163.367
R330 B.n96 B.n93 163.367
R331 B.n97 B.n96 163.367
R332 B.n98 B.n97 163.367
R333 B.n98 B.n91 163.367
R334 B.n102 B.n91 163.367
R335 B.n103 B.n102 163.367
R336 B.n104 B.n103 163.367
R337 B.n104 B.n89 163.367
R338 B.n108 B.n89 163.367
R339 B.n109 B.n108 163.367
R340 B.n110 B.n109 163.367
R341 B.n110 B.n87 163.367
R342 B.n114 B.n87 163.367
R343 B.n115 B.n114 163.367
R344 B.n116 B.n115 163.367
R345 B.n116 B.n85 163.367
R346 B.n120 B.n85 163.367
R347 B.n121 B.n120 163.367
R348 B.n122 B.n121 163.367
R349 B.n122 B.n83 163.367
R350 B.n126 B.n83 163.367
R351 B.n127 B.n126 163.367
R352 B.n128 B.n127 163.367
R353 B.n128 B.n81 163.367
R354 B.n132 B.n81 163.367
R355 B.n133 B.n132 163.367
R356 B.n134 B.n133 163.367
R357 B.n134 B.n79 163.367
R358 B.n75 B.n74 73.1157
R359 B.n163 B.n162 73.1157
R360 B.n29 B.n28 73.1157
R361 B.n23 B.n22 73.1157
R362 B.n149 B.n75 59.5399
R363 B.n164 B.n163 59.5399
R364 B.n284 B.n29 59.5399
R365 B.n298 B.n23 59.5399
R366 B.n311 B.n310 32.0005
R367 B.n272 B.n271 32.0005
R368 B.n177 B.n64 32.0005
R369 B.n137 B.n136 32.0005
R370 B B.n357 18.0485
R371 B.n311 B.n16 10.6151
R372 B.n315 B.n16 10.6151
R373 B.n316 B.n315 10.6151
R374 B.n317 B.n316 10.6151
R375 B.n317 B.n14 10.6151
R376 B.n321 B.n14 10.6151
R377 B.n322 B.n321 10.6151
R378 B.n323 B.n322 10.6151
R379 B.n323 B.n12 10.6151
R380 B.n327 B.n12 10.6151
R381 B.n328 B.n327 10.6151
R382 B.n329 B.n328 10.6151
R383 B.n329 B.n10 10.6151
R384 B.n333 B.n10 10.6151
R385 B.n334 B.n333 10.6151
R386 B.n335 B.n334 10.6151
R387 B.n335 B.n8 10.6151
R388 B.n339 B.n8 10.6151
R389 B.n340 B.n339 10.6151
R390 B.n341 B.n340 10.6151
R391 B.n341 B.n6 10.6151
R392 B.n345 B.n6 10.6151
R393 B.n346 B.n345 10.6151
R394 B.n347 B.n346 10.6151
R395 B.n347 B.n4 10.6151
R396 B.n351 B.n4 10.6151
R397 B.n352 B.n351 10.6151
R398 B.n353 B.n352 10.6151
R399 B.n353 B.n0 10.6151
R400 B.n310 B.n309 10.6151
R401 B.n309 B.n18 10.6151
R402 B.n305 B.n18 10.6151
R403 B.n305 B.n304 10.6151
R404 B.n304 B.n303 10.6151
R405 B.n303 B.n20 10.6151
R406 B.n299 B.n20 10.6151
R407 B.n297 B.n296 10.6151
R408 B.n296 B.n24 10.6151
R409 B.n292 B.n24 10.6151
R410 B.n292 B.n291 10.6151
R411 B.n291 B.n290 10.6151
R412 B.n290 B.n26 10.6151
R413 B.n286 B.n26 10.6151
R414 B.n286 B.n285 10.6151
R415 B.n283 B.n30 10.6151
R416 B.n279 B.n30 10.6151
R417 B.n279 B.n278 10.6151
R418 B.n278 B.n277 10.6151
R419 B.n277 B.n32 10.6151
R420 B.n273 B.n32 10.6151
R421 B.n273 B.n272 10.6151
R422 B.n271 B.n34 10.6151
R423 B.n267 B.n34 10.6151
R424 B.n267 B.n266 10.6151
R425 B.n266 B.n265 10.6151
R426 B.n265 B.n36 10.6151
R427 B.n261 B.n36 10.6151
R428 B.n261 B.n260 10.6151
R429 B.n260 B.n259 10.6151
R430 B.n259 B.n38 10.6151
R431 B.n255 B.n38 10.6151
R432 B.n255 B.n254 10.6151
R433 B.n254 B.n253 10.6151
R434 B.n253 B.n40 10.6151
R435 B.n249 B.n40 10.6151
R436 B.n249 B.n248 10.6151
R437 B.n248 B.n247 10.6151
R438 B.n247 B.n42 10.6151
R439 B.n243 B.n42 10.6151
R440 B.n243 B.n242 10.6151
R441 B.n242 B.n241 10.6151
R442 B.n241 B.n44 10.6151
R443 B.n237 B.n44 10.6151
R444 B.n237 B.n236 10.6151
R445 B.n236 B.n235 10.6151
R446 B.n235 B.n46 10.6151
R447 B.n231 B.n46 10.6151
R448 B.n231 B.n230 10.6151
R449 B.n230 B.n229 10.6151
R450 B.n229 B.n48 10.6151
R451 B.n225 B.n48 10.6151
R452 B.n225 B.n224 10.6151
R453 B.n224 B.n223 10.6151
R454 B.n223 B.n50 10.6151
R455 B.n219 B.n50 10.6151
R456 B.n219 B.n218 10.6151
R457 B.n218 B.n217 10.6151
R458 B.n217 B.n52 10.6151
R459 B.n213 B.n52 10.6151
R460 B.n213 B.n212 10.6151
R461 B.n212 B.n211 10.6151
R462 B.n211 B.n54 10.6151
R463 B.n207 B.n54 10.6151
R464 B.n207 B.n206 10.6151
R465 B.n206 B.n205 10.6151
R466 B.n205 B.n56 10.6151
R467 B.n201 B.n56 10.6151
R468 B.n201 B.n200 10.6151
R469 B.n200 B.n199 10.6151
R470 B.n199 B.n58 10.6151
R471 B.n195 B.n58 10.6151
R472 B.n195 B.n194 10.6151
R473 B.n194 B.n193 10.6151
R474 B.n193 B.n60 10.6151
R475 B.n189 B.n60 10.6151
R476 B.n189 B.n188 10.6151
R477 B.n188 B.n187 10.6151
R478 B.n187 B.n62 10.6151
R479 B.n183 B.n62 10.6151
R480 B.n183 B.n182 10.6151
R481 B.n182 B.n181 10.6151
R482 B.n181 B.n64 10.6151
R483 B.n94 B.n1 10.6151
R484 B.n95 B.n94 10.6151
R485 B.n95 B.n92 10.6151
R486 B.n99 B.n92 10.6151
R487 B.n100 B.n99 10.6151
R488 B.n101 B.n100 10.6151
R489 B.n101 B.n90 10.6151
R490 B.n105 B.n90 10.6151
R491 B.n106 B.n105 10.6151
R492 B.n107 B.n106 10.6151
R493 B.n107 B.n88 10.6151
R494 B.n111 B.n88 10.6151
R495 B.n112 B.n111 10.6151
R496 B.n113 B.n112 10.6151
R497 B.n113 B.n86 10.6151
R498 B.n117 B.n86 10.6151
R499 B.n118 B.n117 10.6151
R500 B.n119 B.n118 10.6151
R501 B.n119 B.n84 10.6151
R502 B.n123 B.n84 10.6151
R503 B.n124 B.n123 10.6151
R504 B.n125 B.n124 10.6151
R505 B.n125 B.n82 10.6151
R506 B.n129 B.n82 10.6151
R507 B.n130 B.n129 10.6151
R508 B.n131 B.n130 10.6151
R509 B.n131 B.n80 10.6151
R510 B.n135 B.n80 10.6151
R511 B.n136 B.n135 10.6151
R512 B.n137 B.n78 10.6151
R513 B.n141 B.n78 10.6151
R514 B.n142 B.n141 10.6151
R515 B.n143 B.n142 10.6151
R516 B.n143 B.n76 10.6151
R517 B.n147 B.n76 10.6151
R518 B.n148 B.n147 10.6151
R519 B.n150 B.n72 10.6151
R520 B.n154 B.n72 10.6151
R521 B.n155 B.n154 10.6151
R522 B.n156 B.n155 10.6151
R523 B.n156 B.n70 10.6151
R524 B.n160 B.n70 10.6151
R525 B.n161 B.n160 10.6151
R526 B.n165 B.n161 10.6151
R527 B.n169 B.n68 10.6151
R528 B.n170 B.n169 10.6151
R529 B.n171 B.n170 10.6151
R530 B.n171 B.n66 10.6151
R531 B.n175 B.n66 10.6151
R532 B.n176 B.n175 10.6151
R533 B.n177 B.n176 10.6151
R534 B.n357 B.n0 8.11757
R535 B.n357 B.n1 8.11757
R536 B.n298 B.n297 6.5566
R537 B.n285 B.n284 6.5566
R538 B.n150 B.n149 6.5566
R539 B.n165 B.n164 6.5566
R540 B.n299 B.n298 4.05904
R541 B.n284 B.n283 4.05904
R542 B.n149 B.n148 4.05904
R543 B.n164 B.n68 4.05904
R544 VP.n0 VP.t0 80.6958
R545 VP.n0 VP.t1 42.5013
R546 VP VP.n0 0.52637
R547 VTAIL.n3 VTAIL.t1 677.158
R548 VTAIL.n0 VTAIL.t2 677.158
R549 VTAIL.n2 VTAIL.t3 677.158
R550 VTAIL.n1 VTAIL.t0 677.158
R551 VTAIL.n1 VTAIL.n0 19.3238
R552 VTAIL.n3 VTAIL.n2 16.0738
R553 VTAIL.n2 VTAIL.n1 2.09533
R554 VTAIL VTAIL.n0 1.34102
R555 VTAIL VTAIL.n3 0.75481
R556 VDD1 VDD1.t0 725.79
R557 VDD1 VDD1.t1 694.707
R558 VN VN.t0 80.6029
R559 VN VN.t1 43.0272
R560 VDD2.n0 VDD2.t0 724.453
R561 VDD2.n0 VDD2.t1 693.837
R562 VDD2 VDD2.n0 0.87119
C0 VDD1 VP 0.599638f
C1 VDD2 B 0.934935f
C2 B VP 1.45687f
C3 VDD2 VTAIL 2.38438f
C4 VN VDD1 0.15698f
C5 w_n2478_n1074# VDD2 1.11263f
C6 VTAIL VP 1.03852f
C7 B VN 0.933169f
C8 w_n2478_n1074# VP 3.55132f
C9 B VDD1 0.896357f
C10 VTAIL VN 1.02441f
C11 w_n2478_n1074# VN 3.24338f
C12 VTAIL VDD1 2.32541f
C13 w_n2478_n1074# VDD1 1.07772f
C14 VTAIL B 1.02189f
C15 w_n2478_n1074# B 6.62432f
C16 VDD2 VP 0.377719f
C17 w_n2478_n1074# VTAIL 1.10516f
C18 VDD2 VN 0.38134f
C19 VN VP 3.73531f
C20 VDD2 VDD1 0.776245f
C21 VDD2 VSUBS 0.607997f
C22 VDD1 VSUBS 2.915478f
C23 VTAIL VSUBS 0.37448f
C24 VN VSUBS 6.43066f
C25 VP VSUBS 1.465638f
C26 B VSUBS 3.361667f
C27 w_n2478_n1074# VSUBS 34.523502f
C28 VDD2.t0 VSUBS 0.079163f
C29 VDD2.t1 VSUBS 0.042565f
C30 VDD2.n0 VSUBS 2.10026f
C31 VN.t1 VSUBS 0.7079f
C32 VN.t0 VSUBS 1.97258f
C33 VDD1.t1 VSUBS 0.039607f
C34 VDD1.t0 VSUBS 0.077874f
C35 VTAIL.t2 VSUBS 0.05361f
C36 VTAIL.n0 VSUBS 1.20202f
C37 VTAIL.t0 VSUBS 0.05361f
C38 VTAIL.n1 VSUBS 1.27188f
C39 VTAIL.t3 VSUBS 0.05361f
C40 VTAIL.n2 VSUBS 0.9709f
C41 VTAIL.t1 VSUBS 0.05361f
C42 VTAIL.n3 VSUBS 0.846756f
C43 VP.t0 VSUBS 2.10917f
C44 VP.t1 VSUBS 0.752134f
C45 VP.n0 VSUBS 4.19829f
C46 B.n0 VSUBS 0.011541f
C47 B.n1 VSUBS 0.011541f
C48 B.n2 VSUBS 0.017068f
C49 B.n3 VSUBS 0.013079f
C50 B.n4 VSUBS 0.013079f
C51 B.n5 VSUBS 0.013079f
C52 B.n6 VSUBS 0.013079f
C53 B.n7 VSUBS 0.013079f
C54 B.n8 VSUBS 0.013079f
C55 B.n9 VSUBS 0.013079f
C56 B.n10 VSUBS 0.013079f
C57 B.n11 VSUBS 0.013079f
C58 B.n12 VSUBS 0.013079f
C59 B.n13 VSUBS 0.013079f
C60 B.n14 VSUBS 0.013079f
C61 B.n15 VSUBS 0.013079f
C62 B.n16 VSUBS 0.013079f
C63 B.n17 VSUBS 0.030448f
C64 B.n18 VSUBS 0.013079f
C65 B.n19 VSUBS 0.013079f
C66 B.n20 VSUBS 0.013079f
C67 B.n21 VSUBS 0.013079f
C68 B.t4 VSUBS 0.018472f
C69 B.t5 VSUBS 0.024342f
C70 B.t3 VSUBS 0.171877f
C71 B.n22 VSUBS 0.121267f
C72 B.n23 VSUBS 0.07802f
C73 B.n24 VSUBS 0.013079f
C74 B.n25 VSUBS 0.013079f
C75 B.n26 VSUBS 0.013079f
C76 B.n27 VSUBS 0.013079f
C77 B.t1 VSUBS 0.018472f
C78 B.t2 VSUBS 0.024342f
C79 B.t0 VSUBS 0.171877f
C80 B.n28 VSUBS 0.121267f
C81 B.n29 VSUBS 0.07802f
C82 B.n30 VSUBS 0.013079f
C83 B.n31 VSUBS 0.013079f
C84 B.n32 VSUBS 0.013079f
C85 B.n33 VSUBS 0.030448f
C86 B.n34 VSUBS 0.013079f
C87 B.n35 VSUBS 0.013079f
C88 B.n36 VSUBS 0.013079f
C89 B.n37 VSUBS 0.013079f
C90 B.n38 VSUBS 0.013079f
C91 B.n39 VSUBS 0.013079f
C92 B.n40 VSUBS 0.013079f
C93 B.n41 VSUBS 0.013079f
C94 B.n42 VSUBS 0.013079f
C95 B.n43 VSUBS 0.013079f
C96 B.n44 VSUBS 0.013079f
C97 B.n45 VSUBS 0.013079f
C98 B.n46 VSUBS 0.013079f
C99 B.n47 VSUBS 0.013079f
C100 B.n48 VSUBS 0.013079f
C101 B.n49 VSUBS 0.013079f
C102 B.n50 VSUBS 0.013079f
C103 B.n51 VSUBS 0.013079f
C104 B.n52 VSUBS 0.013079f
C105 B.n53 VSUBS 0.013079f
C106 B.n54 VSUBS 0.013079f
C107 B.n55 VSUBS 0.013079f
C108 B.n56 VSUBS 0.013079f
C109 B.n57 VSUBS 0.013079f
C110 B.n58 VSUBS 0.013079f
C111 B.n59 VSUBS 0.013079f
C112 B.n60 VSUBS 0.013079f
C113 B.n61 VSUBS 0.013079f
C114 B.n62 VSUBS 0.013079f
C115 B.n63 VSUBS 0.013079f
C116 B.n64 VSUBS 0.031526f
C117 B.n65 VSUBS 0.013079f
C118 B.n66 VSUBS 0.013079f
C119 B.n67 VSUBS 0.013079f
C120 B.n68 VSUBS 0.00904f
C121 B.n69 VSUBS 0.013079f
C122 B.n70 VSUBS 0.013079f
C123 B.n71 VSUBS 0.013079f
C124 B.n72 VSUBS 0.013079f
C125 B.n73 VSUBS 0.013079f
C126 B.t8 VSUBS 0.018472f
C127 B.t7 VSUBS 0.024342f
C128 B.t6 VSUBS 0.171877f
C129 B.n74 VSUBS 0.121267f
C130 B.n75 VSUBS 0.07802f
C131 B.n76 VSUBS 0.013079f
C132 B.n77 VSUBS 0.013079f
C133 B.n78 VSUBS 0.013079f
C134 B.n79 VSUBS 0.029948f
C135 B.n80 VSUBS 0.013079f
C136 B.n81 VSUBS 0.013079f
C137 B.n82 VSUBS 0.013079f
C138 B.n83 VSUBS 0.013079f
C139 B.n84 VSUBS 0.013079f
C140 B.n85 VSUBS 0.013079f
C141 B.n86 VSUBS 0.013079f
C142 B.n87 VSUBS 0.013079f
C143 B.n88 VSUBS 0.013079f
C144 B.n89 VSUBS 0.013079f
C145 B.n90 VSUBS 0.013079f
C146 B.n91 VSUBS 0.013079f
C147 B.n92 VSUBS 0.013079f
C148 B.n93 VSUBS 0.013079f
C149 B.n94 VSUBS 0.013079f
C150 B.n95 VSUBS 0.013079f
C151 B.n96 VSUBS 0.013079f
C152 B.n97 VSUBS 0.013079f
C153 B.n98 VSUBS 0.013079f
C154 B.n99 VSUBS 0.013079f
C155 B.n100 VSUBS 0.013079f
C156 B.n101 VSUBS 0.013079f
C157 B.n102 VSUBS 0.013079f
C158 B.n103 VSUBS 0.013079f
C159 B.n104 VSUBS 0.013079f
C160 B.n105 VSUBS 0.013079f
C161 B.n106 VSUBS 0.013079f
C162 B.n107 VSUBS 0.013079f
C163 B.n108 VSUBS 0.013079f
C164 B.n109 VSUBS 0.013079f
C165 B.n110 VSUBS 0.013079f
C166 B.n111 VSUBS 0.013079f
C167 B.n112 VSUBS 0.013079f
C168 B.n113 VSUBS 0.013079f
C169 B.n114 VSUBS 0.013079f
C170 B.n115 VSUBS 0.013079f
C171 B.n116 VSUBS 0.013079f
C172 B.n117 VSUBS 0.013079f
C173 B.n118 VSUBS 0.013079f
C174 B.n119 VSUBS 0.013079f
C175 B.n120 VSUBS 0.013079f
C176 B.n121 VSUBS 0.013079f
C177 B.n122 VSUBS 0.013079f
C178 B.n123 VSUBS 0.013079f
C179 B.n124 VSUBS 0.013079f
C180 B.n125 VSUBS 0.013079f
C181 B.n126 VSUBS 0.013079f
C182 B.n127 VSUBS 0.013079f
C183 B.n128 VSUBS 0.013079f
C184 B.n129 VSUBS 0.013079f
C185 B.n130 VSUBS 0.013079f
C186 B.n131 VSUBS 0.013079f
C187 B.n132 VSUBS 0.013079f
C188 B.n133 VSUBS 0.013079f
C189 B.n134 VSUBS 0.013079f
C190 B.n135 VSUBS 0.013079f
C191 B.n136 VSUBS 0.029948f
C192 B.n137 VSUBS 0.030448f
C193 B.n138 VSUBS 0.030448f
C194 B.n139 VSUBS 0.013079f
C195 B.n140 VSUBS 0.013079f
C196 B.n141 VSUBS 0.013079f
C197 B.n142 VSUBS 0.013079f
C198 B.n143 VSUBS 0.013079f
C199 B.n144 VSUBS 0.013079f
C200 B.n145 VSUBS 0.013079f
C201 B.n146 VSUBS 0.013079f
C202 B.n147 VSUBS 0.013079f
C203 B.n148 VSUBS 0.00904f
C204 B.n149 VSUBS 0.030304f
C205 B.n150 VSUBS 0.010579f
C206 B.n151 VSUBS 0.013079f
C207 B.n152 VSUBS 0.013079f
C208 B.n153 VSUBS 0.013079f
C209 B.n154 VSUBS 0.013079f
C210 B.n155 VSUBS 0.013079f
C211 B.n156 VSUBS 0.013079f
C212 B.n157 VSUBS 0.013079f
C213 B.n158 VSUBS 0.013079f
C214 B.n159 VSUBS 0.013079f
C215 B.n160 VSUBS 0.013079f
C216 B.n161 VSUBS 0.013079f
C217 B.t11 VSUBS 0.018472f
C218 B.t10 VSUBS 0.024342f
C219 B.t9 VSUBS 0.171877f
C220 B.n162 VSUBS 0.121267f
C221 B.n163 VSUBS 0.07802f
C222 B.n164 VSUBS 0.030304f
C223 B.n165 VSUBS 0.010579f
C224 B.n166 VSUBS 0.013079f
C225 B.n167 VSUBS 0.013079f
C226 B.n168 VSUBS 0.013079f
C227 B.n169 VSUBS 0.013079f
C228 B.n170 VSUBS 0.013079f
C229 B.n171 VSUBS 0.013079f
C230 B.n172 VSUBS 0.013079f
C231 B.n173 VSUBS 0.013079f
C232 B.n174 VSUBS 0.013079f
C233 B.n175 VSUBS 0.013079f
C234 B.n176 VSUBS 0.013079f
C235 B.n177 VSUBS 0.028871f
C236 B.n178 VSUBS 0.030448f
C237 B.n179 VSUBS 0.029948f
C238 B.n180 VSUBS 0.013079f
C239 B.n181 VSUBS 0.013079f
C240 B.n182 VSUBS 0.013079f
C241 B.n183 VSUBS 0.013079f
C242 B.n184 VSUBS 0.013079f
C243 B.n185 VSUBS 0.013079f
C244 B.n186 VSUBS 0.013079f
C245 B.n187 VSUBS 0.013079f
C246 B.n188 VSUBS 0.013079f
C247 B.n189 VSUBS 0.013079f
C248 B.n190 VSUBS 0.013079f
C249 B.n191 VSUBS 0.013079f
C250 B.n192 VSUBS 0.013079f
C251 B.n193 VSUBS 0.013079f
C252 B.n194 VSUBS 0.013079f
C253 B.n195 VSUBS 0.013079f
C254 B.n196 VSUBS 0.013079f
C255 B.n197 VSUBS 0.013079f
C256 B.n198 VSUBS 0.013079f
C257 B.n199 VSUBS 0.013079f
C258 B.n200 VSUBS 0.013079f
C259 B.n201 VSUBS 0.013079f
C260 B.n202 VSUBS 0.013079f
C261 B.n203 VSUBS 0.013079f
C262 B.n204 VSUBS 0.013079f
C263 B.n205 VSUBS 0.013079f
C264 B.n206 VSUBS 0.013079f
C265 B.n207 VSUBS 0.013079f
C266 B.n208 VSUBS 0.013079f
C267 B.n209 VSUBS 0.013079f
C268 B.n210 VSUBS 0.013079f
C269 B.n211 VSUBS 0.013079f
C270 B.n212 VSUBS 0.013079f
C271 B.n213 VSUBS 0.013079f
C272 B.n214 VSUBS 0.013079f
C273 B.n215 VSUBS 0.013079f
C274 B.n216 VSUBS 0.013079f
C275 B.n217 VSUBS 0.013079f
C276 B.n218 VSUBS 0.013079f
C277 B.n219 VSUBS 0.013079f
C278 B.n220 VSUBS 0.013079f
C279 B.n221 VSUBS 0.013079f
C280 B.n222 VSUBS 0.013079f
C281 B.n223 VSUBS 0.013079f
C282 B.n224 VSUBS 0.013079f
C283 B.n225 VSUBS 0.013079f
C284 B.n226 VSUBS 0.013079f
C285 B.n227 VSUBS 0.013079f
C286 B.n228 VSUBS 0.013079f
C287 B.n229 VSUBS 0.013079f
C288 B.n230 VSUBS 0.013079f
C289 B.n231 VSUBS 0.013079f
C290 B.n232 VSUBS 0.013079f
C291 B.n233 VSUBS 0.013079f
C292 B.n234 VSUBS 0.013079f
C293 B.n235 VSUBS 0.013079f
C294 B.n236 VSUBS 0.013079f
C295 B.n237 VSUBS 0.013079f
C296 B.n238 VSUBS 0.013079f
C297 B.n239 VSUBS 0.013079f
C298 B.n240 VSUBS 0.013079f
C299 B.n241 VSUBS 0.013079f
C300 B.n242 VSUBS 0.013079f
C301 B.n243 VSUBS 0.013079f
C302 B.n244 VSUBS 0.013079f
C303 B.n245 VSUBS 0.013079f
C304 B.n246 VSUBS 0.013079f
C305 B.n247 VSUBS 0.013079f
C306 B.n248 VSUBS 0.013079f
C307 B.n249 VSUBS 0.013079f
C308 B.n250 VSUBS 0.013079f
C309 B.n251 VSUBS 0.013079f
C310 B.n252 VSUBS 0.013079f
C311 B.n253 VSUBS 0.013079f
C312 B.n254 VSUBS 0.013079f
C313 B.n255 VSUBS 0.013079f
C314 B.n256 VSUBS 0.013079f
C315 B.n257 VSUBS 0.013079f
C316 B.n258 VSUBS 0.013079f
C317 B.n259 VSUBS 0.013079f
C318 B.n260 VSUBS 0.013079f
C319 B.n261 VSUBS 0.013079f
C320 B.n262 VSUBS 0.013079f
C321 B.n263 VSUBS 0.013079f
C322 B.n264 VSUBS 0.013079f
C323 B.n265 VSUBS 0.013079f
C324 B.n266 VSUBS 0.013079f
C325 B.n267 VSUBS 0.013079f
C326 B.n268 VSUBS 0.013079f
C327 B.n269 VSUBS 0.013079f
C328 B.n270 VSUBS 0.029948f
C329 B.n271 VSUBS 0.029948f
C330 B.n272 VSUBS 0.030448f
C331 B.n273 VSUBS 0.013079f
C332 B.n274 VSUBS 0.013079f
C333 B.n275 VSUBS 0.013079f
C334 B.n276 VSUBS 0.013079f
C335 B.n277 VSUBS 0.013079f
C336 B.n278 VSUBS 0.013079f
C337 B.n279 VSUBS 0.013079f
C338 B.n280 VSUBS 0.013079f
C339 B.n281 VSUBS 0.013079f
C340 B.n282 VSUBS 0.013079f
C341 B.n283 VSUBS 0.00904f
C342 B.n284 VSUBS 0.030304f
C343 B.n285 VSUBS 0.010579f
C344 B.n286 VSUBS 0.013079f
C345 B.n287 VSUBS 0.013079f
C346 B.n288 VSUBS 0.013079f
C347 B.n289 VSUBS 0.013079f
C348 B.n290 VSUBS 0.013079f
C349 B.n291 VSUBS 0.013079f
C350 B.n292 VSUBS 0.013079f
C351 B.n293 VSUBS 0.013079f
C352 B.n294 VSUBS 0.013079f
C353 B.n295 VSUBS 0.013079f
C354 B.n296 VSUBS 0.013079f
C355 B.n297 VSUBS 0.010579f
C356 B.n298 VSUBS 0.030304f
C357 B.n299 VSUBS 0.00904f
C358 B.n300 VSUBS 0.013079f
C359 B.n301 VSUBS 0.013079f
C360 B.n302 VSUBS 0.013079f
C361 B.n303 VSUBS 0.013079f
C362 B.n304 VSUBS 0.013079f
C363 B.n305 VSUBS 0.013079f
C364 B.n306 VSUBS 0.013079f
C365 B.n307 VSUBS 0.013079f
C366 B.n308 VSUBS 0.013079f
C367 B.n309 VSUBS 0.013079f
C368 B.n310 VSUBS 0.030448f
C369 B.n311 VSUBS 0.029948f
C370 B.n312 VSUBS 0.029948f
C371 B.n313 VSUBS 0.013079f
C372 B.n314 VSUBS 0.013079f
C373 B.n315 VSUBS 0.013079f
C374 B.n316 VSUBS 0.013079f
C375 B.n317 VSUBS 0.013079f
C376 B.n318 VSUBS 0.013079f
C377 B.n319 VSUBS 0.013079f
C378 B.n320 VSUBS 0.013079f
C379 B.n321 VSUBS 0.013079f
C380 B.n322 VSUBS 0.013079f
C381 B.n323 VSUBS 0.013079f
C382 B.n324 VSUBS 0.013079f
C383 B.n325 VSUBS 0.013079f
C384 B.n326 VSUBS 0.013079f
C385 B.n327 VSUBS 0.013079f
C386 B.n328 VSUBS 0.013079f
C387 B.n329 VSUBS 0.013079f
C388 B.n330 VSUBS 0.013079f
C389 B.n331 VSUBS 0.013079f
C390 B.n332 VSUBS 0.013079f
C391 B.n333 VSUBS 0.013079f
C392 B.n334 VSUBS 0.013079f
C393 B.n335 VSUBS 0.013079f
C394 B.n336 VSUBS 0.013079f
C395 B.n337 VSUBS 0.013079f
C396 B.n338 VSUBS 0.013079f
C397 B.n339 VSUBS 0.013079f
C398 B.n340 VSUBS 0.013079f
C399 B.n341 VSUBS 0.013079f
C400 B.n342 VSUBS 0.013079f
C401 B.n343 VSUBS 0.013079f
C402 B.n344 VSUBS 0.013079f
C403 B.n345 VSUBS 0.013079f
C404 B.n346 VSUBS 0.013079f
C405 B.n347 VSUBS 0.013079f
C406 B.n348 VSUBS 0.013079f
C407 B.n349 VSUBS 0.013079f
C408 B.n350 VSUBS 0.013079f
C409 B.n351 VSUBS 0.013079f
C410 B.n352 VSUBS 0.013079f
C411 B.n353 VSUBS 0.013079f
C412 B.n354 VSUBS 0.013079f
C413 B.n355 VSUBS 0.017068f
C414 B.n356 VSUBS 0.018182f
C415 B.n357 VSUBS 0.036156f
.ends

