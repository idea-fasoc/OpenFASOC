* NGSPICE file created from diff_pair_sample_0639.ext - technology: sky130A

.subckt diff_pair_sample_0639 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0.6162 ps=3.94 w=1.58 l=0.93
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0 ps=0 w=1.58 l=0.93
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0 ps=0 w=1.58 l=0.93
X3 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0.6162 ps=3.94 w=1.58 l=0.93
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0 ps=0 w=1.58 l=0.93
X5 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0.6162 ps=3.94 w=1.58 l=0.93
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0 ps=0 w=1.58 l=0.93
X7 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.6162 pd=3.94 as=0.6162 ps=3.94 w=1.58 l=0.93
R0 VN VN.t0 277.214
R1 VN VN.t1 244.536
R2 VTAIL.n3 VTAIL.t3 110.665
R3 VTAIL.n0 VTAIL.t1 110.665
R4 VTAIL.n2 VTAIL.t0 110.665
R5 VTAIL.n1 VTAIL.t2 110.665
R6 VTAIL.n1 VTAIL.n0 15.9186
R7 VTAIL.n3 VTAIL.n2 14.8324
R8 VTAIL.n2 VTAIL.n1 1.01343
R9 VTAIL VTAIL.n0 0.800069
R10 VTAIL VTAIL.n3 0.213862
R11 VDD2.n0 VDD2.t0 154.555
R12 VDD2.n0 VDD2.t1 127.344
R13 VDD2 VDD2.n0 0.330241
R14 B.n293 B.n292 585
R15 B.n112 B.n48 585
R16 B.n111 B.n110 585
R17 B.n109 B.n108 585
R18 B.n107 B.n106 585
R19 B.n105 B.n104 585
R20 B.n103 B.n102 585
R21 B.n101 B.n100 585
R22 B.n99 B.n98 585
R23 B.n97 B.n96 585
R24 B.n95 B.n94 585
R25 B.n92 B.n91 585
R26 B.n90 B.n89 585
R27 B.n88 B.n87 585
R28 B.n86 B.n85 585
R29 B.n84 B.n83 585
R30 B.n82 B.n81 585
R31 B.n80 B.n79 585
R32 B.n78 B.n77 585
R33 B.n76 B.n75 585
R34 B.n74 B.n73 585
R35 B.n71 B.n70 585
R36 B.n69 B.n68 585
R37 B.n67 B.n66 585
R38 B.n65 B.n64 585
R39 B.n63 B.n62 585
R40 B.n61 B.n60 585
R41 B.n59 B.n58 585
R42 B.n57 B.n56 585
R43 B.n55 B.n54 585
R44 B.n33 B.n32 585
R45 B.n298 B.n297 585
R46 B.n291 B.n49 585
R47 B.n49 B.n30 585
R48 B.n290 B.n29 585
R49 B.n302 B.n29 585
R50 B.n289 B.n28 585
R51 B.n303 B.n28 585
R52 B.n288 B.n27 585
R53 B.n304 B.n27 585
R54 B.n287 B.n286 585
R55 B.n286 B.n23 585
R56 B.n285 B.n22 585
R57 B.n310 B.n22 585
R58 B.n284 B.n21 585
R59 B.n311 B.n21 585
R60 B.n283 B.n20 585
R61 B.n312 B.n20 585
R62 B.n282 B.n281 585
R63 B.n281 B.n16 585
R64 B.n280 B.n15 585
R65 B.n318 B.n15 585
R66 B.n279 B.n14 585
R67 B.n319 B.n14 585
R68 B.n278 B.n13 585
R69 B.n320 B.n13 585
R70 B.n277 B.n276 585
R71 B.n276 B.n12 585
R72 B.n275 B.n274 585
R73 B.n275 B.n8 585
R74 B.n273 B.n7 585
R75 B.n327 B.n7 585
R76 B.n272 B.n6 585
R77 B.n328 B.n6 585
R78 B.n271 B.n5 585
R79 B.n329 B.n5 585
R80 B.n270 B.n269 585
R81 B.n269 B.n4 585
R82 B.n268 B.n113 585
R83 B.n268 B.n267 585
R84 B.n257 B.n114 585
R85 B.n260 B.n114 585
R86 B.n259 B.n258 585
R87 B.n261 B.n259 585
R88 B.n256 B.n119 585
R89 B.n119 B.n118 585
R90 B.n255 B.n254 585
R91 B.n254 B.n253 585
R92 B.n121 B.n120 585
R93 B.n122 B.n121 585
R94 B.n246 B.n245 585
R95 B.n247 B.n246 585
R96 B.n244 B.n127 585
R97 B.n127 B.n126 585
R98 B.n243 B.n242 585
R99 B.n242 B.n241 585
R100 B.n129 B.n128 585
R101 B.n130 B.n129 585
R102 B.n234 B.n233 585
R103 B.n235 B.n234 585
R104 B.n232 B.n135 585
R105 B.n135 B.n134 585
R106 B.n231 B.n230 585
R107 B.n230 B.n229 585
R108 B.n137 B.n136 585
R109 B.n138 B.n137 585
R110 B.n225 B.n224 585
R111 B.n141 B.n140 585
R112 B.n221 B.n220 585
R113 B.n222 B.n221 585
R114 B.n219 B.n157 585
R115 B.n218 B.n217 585
R116 B.n216 B.n215 585
R117 B.n214 B.n213 585
R118 B.n212 B.n211 585
R119 B.n210 B.n209 585
R120 B.n208 B.n207 585
R121 B.n206 B.n205 585
R122 B.n204 B.n203 585
R123 B.n202 B.n201 585
R124 B.n200 B.n199 585
R125 B.n198 B.n197 585
R126 B.n196 B.n195 585
R127 B.n194 B.n193 585
R128 B.n192 B.n191 585
R129 B.n190 B.n189 585
R130 B.n188 B.n187 585
R131 B.n186 B.n185 585
R132 B.n184 B.n183 585
R133 B.n182 B.n181 585
R134 B.n180 B.n179 585
R135 B.n178 B.n177 585
R136 B.n176 B.n175 585
R137 B.n174 B.n173 585
R138 B.n172 B.n171 585
R139 B.n170 B.n169 585
R140 B.n168 B.n167 585
R141 B.n166 B.n165 585
R142 B.n164 B.n156 585
R143 B.n222 B.n156 585
R144 B.n226 B.n139 585
R145 B.n139 B.n138 585
R146 B.n228 B.n227 585
R147 B.n229 B.n228 585
R148 B.n133 B.n132 585
R149 B.n134 B.n133 585
R150 B.n237 B.n236 585
R151 B.n236 B.n235 585
R152 B.n238 B.n131 585
R153 B.n131 B.n130 585
R154 B.n240 B.n239 585
R155 B.n241 B.n240 585
R156 B.n125 B.n124 585
R157 B.n126 B.n125 585
R158 B.n249 B.n248 585
R159 B.n248 B.n247 585
R160 B.n250 B.n123 585
R161 B.n123 B.n122 585
R162 B.n252 B.n251 585
R163 B.n253 B.n252 585
R164 B.n117 B.n116 585
R165 B.n118 B.n117 585
R166 B.n263 B.n262 585
R167 B.n262 B.n261 585
R168 B.n264 B.n115 585
R169 B.n260 B.n115 585
R170 B.n266 B.n265 585
R171 B.n267 B.n266 585
R172 B.n3 B.n0 585
R173 B.n4 B.n3 585
R174 B.n326 B.n1 585
R175 B.n327 B.n326 585
R176 B.n325 B.n324 585
R177 B.n325 B.n8 585
R178 B.n323 B.n9 585
R179 B.n12 B.n9 585
R180 B.n322 B.n321 585
R181 B.n321 B.n320 585
R182 B.n11 B.n10 585
R183 B.n319 B.n11 585
R184 B.n317 B.n316 585
R185 B.n318 B.n317 585
R186 B.n315 B.n17 585
R187 B.n17 B.n16 585
R188 B.n314 B.n313 585
R189 B.n313 B.n312 585
R190 B.n19 B.n18 585
R191 B.n311 B.n19 585
R192 B.n309 B.n308 585
R193 B.n310 B.n309 585
R194 B.n307 B.n24 585
R195 B.n24 B.n23 585
R196 B.n306 B.n305 585
R197 B.n305 B.n304 585
R198 B.n26 B.n25 585
R199 B.n303 B.n26 585
R200 B.n301 B.n300 585
R201 B.n302 B.n301 585
R202 B.n299 B.n31 585
R203 B.n31 B.n30 585
R204 B.n330 B.n329 585
R205 B.n328 B.n2 585
R206 B.n297 B.n31 473.281
R207 B.n293 B.n49 473.281
R208 B.n156 B.n137 473.281
R209 B.n224 B.n139 473.281
R210 B.n295 B.n294 256.663
R211 B.n295 B.n47 256.663
R212 B.n295 B.n46 256.663
R213 B.n295 B.n45 256.663
R214 B.n295 B.n44 256.663
R215 B.n295 B.n43 256.663
R216 B.n295 B.n42 256.663
R217 B.n295 B.n41 256.663
R218 B.n295 B.n40 256.663
R219 B.n295 B.n39 256.663
R220 B.n295 B.n38 256.663
R221 B.n295 B.n37 256.663
R222 B.n295 B.n36 256.663
R223 B.n295 B.n35 256.663
R224 B.n295 B.n34 256.663
R225 B.n296 B.n295 256.663
R226 B.n223 B.n222 256.663
R227 B.n222 B.n142 256.663
R228 B.n222 B.n143 256.663
R229 B.n222 B.n144 256.663
R230 B.n222 B.n145 256.663
R231 B.n222 B.n146 256.663
R232 B.n222 B.n147 256.663
R233 B.n222 B.n148 256.663
R234 B.n222 B.n149 256.663
R235 B.n222 B.n150 256.663
R236 B.n222 B.n151 256.663
R237 B.n222 B.n152 256.663
R238 B.n222 B.n153 256.663
R239 B.n222 B.n154 256.663
R240 B.n222 B.n155 256.663
R241 B.n332 B.n331 256.663
R242 B.n52 B.t2 243.371
R243 B.n50 B.t13 243.371
R244 B.n161 B.t10 243.371
R245 B.n158 B.t6 243.371
R246 B.n222 B.n138 200
R247 B.n295 B.n30 200
R248 B.n54 B.n33 163.367
R249 B.n58 B.n57 163.367
R250 B.n62 B.n61 163.367
R251 B.n66 B.n65 163.367
R252 B.n70 B.n69 163.367
R253 B.n75 B.n74 163.367
R254 B.n79 B.n78 163.367
R255 B.n83 B.n82 163.367
R256 B.n87 B.n86 163.367
R257 B.n91 B.n90 163.367
R258 B.n96 B.n95 163.367
R259 B.n100 B.n99 163.367
R260 B.n104 B.n103 163.367
R261 B.n108 B.n107 163.367
R262 B.n110 B.n48 163.367
R263 B.n230 B.n137 163.367
R264 B.n230 B.n135 163.367
R265 B.n234 B.n135 163.367
R266 B.n234 B.n129 163.367
R267 B.n242 B.n129 163.367
R268 B.n242 B.n127 163.367
R269 B.n246 B.n127 163.367
R270 B.n246 B.n121 163.367
R271 B.n254 B.n121 163.367
R272 B.n254 B.n119 163.367
R273 B.n259 B.n119 163.367
R274 B.n259 B.n114 163.367
R275 B.n268 B.n114 163.367
R276 B.n269 B.n268 163.367
R277 B.n269 B.n5 163.367
R278 B.n6 B.n5 163.367
R279 B.n7 B.n6 163.367
R280 B.n275 B.n7 163.367
R281 B.n276 B.n275 163.367
R282 B.n276 B.n13 163.367
R283 B.n14 B.n13 163.367
R284 B.n15 B.n14 163.367
R285 B.n281 B.n15 163.367
R286 B.n281 B.n20 163.367
R287 B.n21 B.n20 163.367
R288 B.n22 B.n21 163.367
R289 B.n286 B.n22 163.367
R290 B.n286 B.n27 163.367
R291 B.n28 B.n27 163.367
R292 B.n29 B.n28 163.367
R293 B.n49 B.n29 163.367
R294 B.n221 B.n141 163.367
R295 B.n221 B.n157 163.367
R296 B.n217 B.n216 163.367
R297 B.n213 B.n212 163.367
R298 B.n209 B.n208 163.367
R299 B.n205 B.n204 163.367
R300 B.n201 B.n200 163.367
R301 B.n197 B.n196 163.367
R302 B.n193 B.n192 163.367
R303 B.n189 B.n188 163.367
R304 B.n185 B.n184 163.367
R305 B.n181 B.n180 163.367
R306 B.n177 B.n176 163.367
R307 B.n173 B.n172 163.367
R308 B.n169 B.n168 163.367
R309 B.n165 B.n156 163.367
R310 B.n228 B.n139 163.367
R311 B.n228 B.n133 163.367
R312 B.n236 B.n133 163.367
R313 B.n236 B.n131 163.367
R314 B.n240 B.n131 163.367
R315 B.n240 B.n125 163.367
R316 B.n248 B.n125 163.367
R317 B.n248 B.n123 163.367
R318 B.n252 B.n123 163.367
R319 B.n252 B.n117 163.367
R320 B.n262 B.n117 163.367
R321 B.n262 B.n115 163.367
R322 B.n266 B.n115 163.367
R323 B.n266 B.n3 163.367
R324 B.n330 B.n3 163.367
R325 B.n326 B.n2 163.367
R326 B.n326 B.n325 163.367
R327 B.n325 B.n9 163.367
R328 B.n321 B.n9 163.367
R329 B.n321 B.n11 163.367
R330 B.n317 B.n11 163.367
R331 B.n317 B.n17 163.367
R332 B.n313 B.n17 163.367
R333 B.n313 B.n19 163.367
R334 B.n309 B.n19 163.367
R335 B.n309 B.n24 163.367
R336 B.n305 B.n24 163.367
R337 B.n305 B.n26 163.367
R338 B.n301 B.n26 163.367
R339 B.n301 B.n31 163.367
R340 B.n50 B.t14 132.659
R341 B.n161 B.t12 132.659
R342 B.n52 B.t4 132.659
R343 B.n158 B.t9 132.659
R344 B.n229 B.n138 108.8
R345 B.n229 B.n134 108.8
R346 B.n235 B.n134 108.8
R347 B.n235 B.n130 108.8
R348 B.n241 B.n130 108.8
R349 B.n247 B.n126 108.8
R350 B.n247 B.n122 108.8
R351 B.n253 B.n122 108.8
R352 B.n253 B.n118 108.8
R353 B.n261 B.n118 108.8
R354 B.n261 B.n260 108.8
R355 B.n267 B.n4 108.8
R356 B.n329 B.n4 108.8
R357 B.n329 B.n328 108.8
R358 B.n328 B.n327 108.8
R359 B.n327 B.n8 108.8
R360 B.n320 B.n12 108.8
R361 B.n320 B.n319 108.8
R362 B.n319 B.n318 108.8
R363 B.n318 B.n16 108.8
R364 B.n312 B.n16 108.8
R365 B.n312 B.n311 108.8
R366 B.n310 B.n23 108.8
R367 B.n304 B.n23 108.8
R368 B.n304 B.n303 108.8
R369 B.n303 B.n302 108.8
R370 B.n302 B.n30 108.8
R371 B.n51 B.t15 108.222
R372 B.n162 B.t11 108.222
R373 B.n53 B.t5 108.222
R374 B.n159 B.t8 108.222
R375 B.n267 B.t1 104.001
R376 B.t0 B.n8 104.001
R377 B.t7 B.n126 94.4005
R378 B.n311 B.t3 94.4005
R379 B.n297 B.n296 71.676
R380 B.n54 B.n34 71.676
R381 B.n58 B.n35 71.676
R382 B.n62 B.n36 71.676
R383 B.n66 B.n37 71.676
R384 B.n70 B.n38 71.676
R385 B.n75 B.n39 71.676
R386 B.n79 B.n40 71.676
R387 B.n83 B.n41 71.676
R388 B.n87 B.n42 71.676
R389 B.n91 B.n43 71.676
R390 B.n96 B.n44 71.676
R391 B.n100 B.n45 71.676
R392 B.n104 B.n46 71.676
R393 B.n108 B.n47 71.676
R394 B.n294 B.n48 71.676
R395 B.n294 B.n293 71.676
R396 B.n110 B.n47 71.676
R397 B.n107 B.n46 71.676
R398 B.n103 B.n45 71.676
R399 B.n99 B.n44 71.676
R400 B.n95 B.n43 71.676
R401 B.n90 B.n42 71.676
R402 B.n86 B.n41 71.676
R403 B.n82 B.n40 71.676
R404 B.n78 B.n39 71.676
R405 B.n74 B.n38 71.676
R406 B.n69 B.n37 71.676
R407 B.n65 B.n36 71.676
R408 B.n61 B.n35 71.676
R409 B.n57 B.n34 71.676
R410 B.n296 B.n33 71.676
R411 B.n224 B.n223 71.676
R412 B.n157 B.n142 71.676
R413 B.n216 B.n143 71.676
R414 B.n212 B.n144 71.676
R415 B.n208 B.n145 71.676
R416 B.n204 B.n146 71.676
R417 B.n200 B.n147 71.676
R418 B.n196 B.n148 71.676
R419 B.n192 B.n149 71.676
R420 B.n188 B.n150 71.676
R421 B.n184 B.n151 71.676
R422 B.n180 B.n152 71.676
R423 B.n176 B.n153 71.676
R424 B.n172 B.n154 71.676
R425 B.n168 B.n155 71.676
R426 B.n223 B.n141 71.676
R427 B.n217 B.n142 71.676
R428 B.n213 B.n143 71.676
R429 B.n209 B.n144 71.676
R430 B.n205 B.n145 71.676
R431 B.n201 B.n146 71.676
R432 B.n197 B.n147 71.676
R433 B.n193 B.n148 71.676
R434 B.n189 B.n149 71.676
R435 B.n185 B.n150 71.676
R436 B.n181 B.n151 71.676
R437 B.n177 B.n152 71.676
R438 B.n173 B.n153 71.676
R439 B.n169 B.n154 71.676
R440 B.n165 B.n155 71.676
R441 B.n331 B.n330 71.676
R442 B.n331 B.n2 71.676
R443 B.n72 B.n53 59.5399
R444 B.n93 B.n51 59.5399
R445 B.n163 B.n162 59.5399
R446 B.n160 B.n159 59.5399
R447 B.n226 B.n225 30.7517
R448 B.n164 B.n136 30.7517
R449 B.n292 B.n291 30.7517
R450 B.n299 B.n298 30.7517
R451 B.n53 B.n52 24.4369
R452 B.n51 B.n50 24.4369
R453 B.n162 B.n161 24.4369
R454 B.n159 B.n158 24.4369
R455 B B.n332 18.0485
R456 B.n241 B.t7 14.4005
R457 B.t3 B.n310 14.4005
R458 B.n227 B.n226 10.6151
R459 B.n227 B.n132 10.6151
R460 B.n237 B.n132 10.6151
R461 B.n238 B.n237 10.6151
R462 B.n239 B.n238 10.6151
R463 B.n239 B.n124 10.6151
R464 B.n249 B.n124 10.6151
R465 B.n250 B.n249 10.6151
R466 B.n251 B.n250 10.6151
R467 B.n251 B.n116 10.6151
R468 B.n263 B.n116 10.6151
R469 B.n264 B.n263 10.6151
R470 B.n265 B.n264 10.6151
R471 B.n265 B.n0 10.6151
R472 B.n225 B.n140 10.6151
R473 B.n220 B.n140 10.6151
R474 B.n220 B.n219 10.6151
R475 B.n219 B.n218 10.6151
R476 B.n218 B.n215 10.6151
R477 B.n215 B.n214 10.6151
R478 B.n214 B.n211 10.6151
R479 B.n211 B.n210 10.6151
R480 B.n210 B.n207 10.6151
R481 B.n207 B.n206 10.6151
R482 B.n203 B.n202 10.6151
R483 B.n202 B.n199 10.6151
R484 B.n199 B.n198 10.6151
R485 B.n198 B.n195 10.6151
R486 B.n195 B.n194 10.6151
R487 B.n194 B.n191 10.6151
R488 B.n191 B.n190 10.6151
R489 B.n190 B.n187 10.6151
R490 B.n187 B.n186 10.6151
R491 B.n183 B.n182 10.6151
R492 B.n182 B.n179 10.6151
R493 B.n179 B.n178 10.6151
R494 B.n178 B.n175 10.6151
R495 B.n175 B.n174 10.6151
R496 B.n174 B.n171 10.6151
R497 B.n171 B.n170 10.6151
R498 B.n170 B.n167 10.6151
R499 B.n167 B.n166 10.6151
R500 B.n166 B.n164 10.6151
R501 B.n231 B.n136 10.6151
R502 B.n232 B.n231 10.6151
R503 B.n233 B.n232 10.6151
R504 B.n233 B.n128 10.6151
R505 B.n243 B.n128 10.6151
R506 B.n244 B.n243 10.6151
R507 B.n245 B.n244 10.6151
R508 B.n245 B.n120 10.6151
R509 B.n255 B.n120 10.6151
R510 B.n256 B.n255 10.6151
R511 B.n258 B.n256 10.6151
R512 B.n258 B.n257 10.6151
R513 B.n257 B.n113 10.6151
R514 B.n270 B.n113 10.6151
R515 B.n271 B.n270 10.6151
R516 B.n272 B.n271 10.6151
R517 B.n273 B.n272 10.6151
R518 B.n274 B.n273 10.6151
R519 B.n277 B.n274 10.6151
R520 B.n278 B.n277 10.6151
R521 B.n279 B.n278 10.6151
R522 B.n280 B.n279 10.6151
R523 B.n282 B.n280 10.6151
R524 B.n283 B.n282 10.6151
R525 B.n284 B.n283 10.6151
R526 B.n285 B.n284 10.6151
R527 B.n287 B.n285 10.6151
R528 B.n288 B.n287 10.6151
R529 B.n289 B.n288 10.6151
R530 B.n290 B.n289 10.6151
R531 B.n291 B.n290 10.6151
R532 B.n324 B.n1 10.6151
R533 B.n324 B.n323 10.6151
R534 B.n323 B.n322 10.6151
R535 B.n322 B.n10 10.6151
R536 B.n316 B.n10 10.6151
R537 B.n316 B.n315 10.6151
R538 B.n315 B.n314 10.6151
R539 B.n314 B.n18 10.6151
R540 B.n308 B.n18 10.6151
R541 B.n308 B.n307 10.6151
R542 B.n307 B.n306 10.6151
R543 B.n306 B.n25 10.6151
R544 B.n300 B.n25 10.6151
R545 B.n300 B.n299 10.6151
R546 B.n298 B.n32 10.6151
R547 B.n55 B.n32 10.6151
R548 B.n56 B.n55 10.6151
R549 B.n59 B.n56 10.6151
R550 B.n60 B.n59 10.6151
R551 B.n63 B.n60 10.6151
R552 B.n64 B.n63 10.6151
R553 B.n67 B.n64 10.6151
R554 B.n68 B.n67 10.6151
R555 B.n71 B.n68 10.6151
R556 B.n76 B.n73 10.6151
R557 B.n77 B.n76 10.6151
R558 B.n80 B.n77 10.6151
R559 B.n81 B.n80 10.6151
R560 B.n84 B.n81 10.6151
R561 B.n85 B.n84 10.6151
R562 B.n88 B.n85 10.6151
R563 B.n89 B.n88 10.6151
R564 B.n92 B.n89 10.6151
R565 B.n97 B.n94 10.6151
R566 B.n98 B.n97 10.6151
R567 B.n101 B.n98 10.6151
R568 B.n102 B.n101 10.6151
R569 B.n105 B.n102 10.6151
R570 B.n106 B.n105 10.6151
R571 B.n109 B.n106 10.6151
R572 B.n111 B.n109 10.6151
R573 B.n112 B.n111 10.6151
R574 B.n292 B.n112 10.6151
R575 B.n206 B.n160 8.74196
R576 B.n183 B.n163 8.74196
R577 B.n72 B.n71 8.74196
R578 B.n94 B.n93 8.74196
R579 B.n332 B.n0 8.11757
R580 B.n332 B.n1 8.11757
R581 B.n260 B.t1 4.8005
R582 B.n12 B.t0 4.8005
R583 B.n203 B.n160 1.87367
R584 B.n186 B.n163 1.87367
R585 B.n73 B.n72 1.87367
R586 B.n93 B.n92 1.87367
R587 VP.n0 VP.t1 276.832
R588 VP.n0 VP.t0 244.484
R589 VP VP.n0 0.0516364
R590 VDD1 VDD1.t1 155.351
R591 VDD1 VDD1.t0 127.674
C0 VTAIL VP 0.608832f
C1 VTAIL VDD1 1.8409f
C2 VDD2 VP 0.271149f
C3 VDD2 VDD1 0.482356f
C4 VTAIL VN 0.594668f
C5 VDD2 VN 0.497797f
C6 VTAIL VDD2 1.88223f
C7 VP VDD1 0.611495f
C8 VN VP 2.74176f
C9 VN VDD1 0.155951f
C10 VDD2 B 1.88508f
C11 VDD1 B 2.02422f
C12 VTAIL B 2.19261f
C13 VN B 5.58028f
C14 VP B 3.438225f
C15 VP.t1 B 0.394878f
C16 VP.t0 B 0.271436f
C17 VP.n0 B 2.0144f
C18 VN.t1 B 0.266005f
C19 VN.t0 B 0.391252f
.ends

