* NGSPICE file created from diff_pair_sample_1611.ext - technology: sky130A

.subckt diff_pair_sample_1611 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 w_n1914_n3500# sky130_fd_pr__pfet_01v8 ad=4.9374 pd=26.1 as=4.9374 ps=26.1 w=12.66 l=2.03
X1 VDD1.t1 VP.t0 VTAIL.t0 w_n1914_n3500# sky130_fd_pr__pfet_01v8 ad=4.9374 pd=26.1 as=4.9374 ps=26.1 w=12.66 l=2.03
X2 B.t11 B.t9 B.t10 w_n1914_n3500# sky130_fd_pr__pfet_01v8 ad=4.9374 pd=26.1 as=0 ps=0 w=12.66 l=2.03
X3 VDD2.t0 VN.t1 VTAIL.t3 w_n1914_n3500# sky130_fd_pr__pfet_01v8 ad=4.9374 pd=26.1 as=4.9374 ps=26.1 w=12.66 l=2.03
X4 B.t8 B.t6 B.t7 w_n1914_n3500# sky130_fd_pr__pfet_01v8 ad=4.9374 pd=26.1 as=0 ps=0 w=12.66 l=2.03
X5 B.t5 B.t3 B.t4 w_n1914_n3500# sky130_fd_pr__pfet_01v8 ad=4.9374 pd=26.1 as=0 ps=0 w=12.66 l=2.03
X6 B.t2 B.t0 B.t1 w_n1914_n3500# sky130_fd_pr__pfet_01v8 ad=4.9374 pd=26.1 as=0 ps=0 w=12.66 l=2.03
X7 VDD1.t0 VP.t1 VTAIL.t1 w_n1914_n3500# sky130_fd_pr__pfet_01v8 ad=4.9374 pd=26.1 as=4.9374 ps=26.1 w=12.66 l=2.03
R0 VN VN.t1 253.02
R1 VN VN.t0 209.427
R2 VTAIL.n278 VTAIL.n277 756.745
R3 VTAIL.n68 VTAIL.n67 756.745
R4 VTAIL.n208 VTAIL.n207 756.745
R5 VTAIL.n138 VTAIL.n137 756.745
R6 VTAIL.n232 VTAIL.n231 585
R7 VTAIL.n237 VTAIL.n236 585
R8 VTAIL.n239 VTAIL.n238 585
R9 VTAIL.n228 VTAIL.n227 585
R10 VTAIL.n245 VTAIL.n244 585
R11 VTAIL.n247 VTAIL.n246 585
R12 VTAIL.n224 VTAIL.n223 585
R13 VTAIL.n253 VTAIL.n252 585
R14 VTAIL.n255 VTAIL.n254 585
R15 VTAIL.n220 VTAIL.n219 585
R16 VTAIL.n261 VTAIL.n260 585
R17 VTAIL.n263 VTAIL.n262 585
R18 VTAIL.n216 VTAIL.n215 585
R19 VTAIL.n269 VTAIL.n268 585
R20 VTAIL.n271 VTAIL.n270 585
R21 VTAIL.n212 VTAIL.n211 585
R22 VTAIL.n277 VTAIL.n276 585
R23 VTAIL.n22 VTAIL.n21 585
R24 VTAIL.n27 VTAIL.n26 585
R25 VTAIL.n29 VTAIL.n28 585
R26 VTAIL.n18 VTAIL.n17 585
R27 VTAIL.n35 VTAIL.n34 585
R28 VTAIL.n37 VTAIL.n36 585
R29 VTAIL.n14 VTAIL.n13 585
R30 VTAIL.n43 VTAIL.n42 585
R31 VTAIL.n45 VTAIL.n44 585
R32 VTAIL.n10 VTAIL.n9 585
R33 VTAIL.n51 VTAIL.n50 585
R34 VTAIL.n53 VTAIL.n52 585
R35 VTAIL.n6 VTAIL.n5 585
R36 VTAIL.n59 VTAIL.n58 585
R37 VTAIL.n61 VTAIL.n60 585
R38 VTAIL.n2 VTAIL.n1 585
R39 VTAIL.n67 VTAIL.n66 585
R40 VTAIL.n207 VTAIL.n206 585
R41 VTAIL.n142 VTAIL.n141 585
R42 VTAIL.n201 VTAIL.n200 585
R43 VTAIL.n199 VTAIL.n198 585
R44 VTAIL.n146 VTAIL.n145 585
R45 VTAIL.n193 VTAIL.n192 585
R46 VTAIL.n191 VTAIL.n190 585
R47 VTAIL.n150 VTAIL.n149 585
R48 VTAIL.n185 VTAIL.n184 585
R49 VTAIL.n183 VTAIL.n182 585
R50 VTAIL.n154 VTAIL.n153 585
R51 VTAIL.n177 VTAIL.n176 585
R52 VTAIL.n175 VTAIL.n174 585
R53 VTAIL.n158 VTAIL.n157 585
R54 VTAIL.n169 VTAIL.n168 585
R55 VTAIL.n167 VTAIL.n166 585
R56 VTAIL.n162 VTAIL.n161 585
R57 VTAIL.n137 VTAIL.n136 585
R58 VTAIL.n72 VTAIL.n71 585
R59 VTAIL.n131 VTAIL.n130 585
R60 VTAIL.n129 VTAIL.n128 585
R61 VTAIL.n76 VTAIL.n75 585
R62 VTAIL.n123 VTAIL.n122 585
R63 VTAIL.n121 VTAIL.n120 585
R64 VTAIL.n80 VTAIL.n79 585
R65 VTAIL.n115 VTAIL.n114 585
R66 VTAIL.n113 VTAIL.n112 585
R67 VTAIL.n84 VTAIL.n83 585
R68 VTAIL.n107 VTAIL.n106 585
R69 VTAIL.n105 VTAIL.n104 585
R70 VTAIL.n88 VTAIL.n87 585
R71 VTAIL.n99 VTAIL.n98 585
R72 VTAIL.n97 VTAIL.n96 585
R73 VTAIL.n92 VTAIL.n91 585
R74 VTAIL.n233 VTAIL.t2 327.466
R75 VTAIL.n23 VTAIL.t1 327.466
R76 VTAIL.n163 VTAIL.t0 327.466
R77 VTAIL.n93 VTAIL.t3 327.466
R78 VTAIL.n237 VTAIL.n231 171.744
R79 VTAIL.n238 VTAIL.n237 171.744
R80 VTAIL.n238 VTAIL.n227 171.744
R81 VTAIL.n245 VTAIL.n227 171.744
R82 VTAIL.n246 VTAIL.n245 171.744
R83 VTAIL.n246 VTAIL.n223 171.744
R84 VTAIL.n253 VTAIL.n223 171.744
R85 VTAIL.n254 VTAIL.n253 171.744
R86 VTAIL.n254 VTAIL.n219 171.744
R87 VTAIL.n261 VTAIL.n219 171.744
R88 VTAIL.n262 VTAIL.n261 171.744
R89 VTAIL.n262 VTAIL.n215 171.744
R90 VTAIL.n269 VTAIL.n215 171.744
R91 VTAIL.n270 VTAIL.n269 171.744
R92 VTAIL.n270 VTAIL.n211 171.744
R93 VTAIL.n277 VTAIL.n211 171.744
R94 VTAIL.n27 VTAIL.n21 171.744
R95 VTAIL.n28 VTAIL.n27 171.744
R96 VTAIL.n28 VTAIL.n17 171.744
R97 VTAIL.n35 VTAIL.n17 171.744
R98 VTAIL.n36 VTAIL.n35 171.744
R99 VTAIL.n36 VTAIL.n13 171.744
R100 VTAIL.n43 VTAIL.n13 171.744
R101 VTAIL.n44 VTAIL.n43 171.744
R102 VTAIL.n44 VTAIL.n9 171.744
R103 VTAIL.n51 VTAIL.n9 171.744
R104 VTAIL.n52 VTAIL.n51 171.744
R105 VTAIL.n52 VTAIL.n5 171.744
R106 VTAIL.n59 VTAIL.n5 171.744
R107 VTAIL.n60 VTAIL.n59 171.744
R108 VTAIL.n60 VTAIL.n1 171.744
R109 VTAIL.n67 VTAIL.n1 171.744
R110 VTAIL.n207 VTAIL.n141 171.744
R111 VTAIL.n200 VTAIL.n141 171.744
R112 VTAIL.n200 VTAIL.n199 171.744
R113 VTAIL.n199 VTAIL.n145 171.744
R114 VTAIL.n192 VTAIL.n145 171.744
R115 VTAIL.n192 VTAIL.n191 171.744
R116 VTAIL.n191 VTAIL.n149 171.744
R117 VTAIL.n184 VTAIL.n149 171.744
R118 VTAIL.n184 VTAIL.n183 171.744
R119 VTAIL.n183 VTAIL.n153 171.744
R120 VTAIL.n176 VTAIL.n153 171.744
R121 VTAIL.n176 VTAIL.n175 171.744
R122 VTAIL.n175 VTAIL.n157 171.744
R123 VTAIL.n168 VTAIL.n157 171.744
R124 VTAIL.n168 VTAIL.n167 171.744
R125 VTAIL.n167 VTAIL.n161 171.744
R126 VTAIL.n137 VTAIL.n71 171.744
R127 VTAIL.n130 VTAIL.n71 171.744
R128 VTAIL.n130 VTAIL.n129 171.744
R129 VTAIL.n129 VTAIL.n75 171.744
R130 VTAIL.n122 VTAIL.n75 171.744
R131 VTAIL.n122 VTAIL.n121 171.744
R132 VTAIL.n121 VTAIL.n79 171.744
R133 VTAIL.n114 VTAIL.n79 171.744
R134 VTAIL.n114 VTAIL.n113 171.744
R135 VTAIL.n113 VTAIL.n83 171.744
R136 VTAIL.n106 VTAIL.n83 171.744
R137 VTAIL.n106 VTAIL.n105 171.744
R138 VTAIL.n105 VTAIL.n87 171.744
R139 VTAIL.n98 VTAIL.n87 171.744
R140 VTAIL.n98 VTAIL.n97 171.744
R141 VTAIL.n97 VTAIL.n91 171.744
R142 VTAIL.t2 VTAIL.n231 85.8723
R143 VTAIL.t1 VTAIL.n21 85.8723
R144 VTAIL.t0 VTAIL.n161 85.8723
R145 VTAIL.t3 VTAIL.n91 85.8723
R146 VTAIL.n279 VTAIL.n278 35.2884
R147 VTAIL.n69 VTAIL.n68 35.2884
R148 VTAIL.n209 VTAIL.n208 35.2884
R149 VTAIL.n139 VTAIL.n138 35.2884
R150 VTAIL.n139 VTAIL.n69 27.3496
R151 VTAIL.n279 VTAIL.n209 25.3152
R152 VTAIL.n233 VTAIL.n232 16.3895
R153 VTAIL.n23 VTAIL.n22 16.3895
R154 VTAIL.n163 VTAIL.n162 16.3895
R155 VTAIL.n93 VTAIL.n92 16.3895
R156 VTAIL.n236 VTAIL.n235 12.8005
R157 VTAIL.n276 VTAIL.n210 12.8005
R158 VTAIL.n26 VTAIL.n25 12.8005
R159 VTAIL.n66 VTAIL.n0 12.8005
R160 VTAIL.n206 VTAIL.n140 12.8005
R161 VTAIL.n166 VTAIL.n165 12.8005
R162 VTAIL.n136 VTAIL.n70 12.8005
R163 VTAIL.n96 VTAIL.n95 12.8005
R164 VTAIL.n239 VTAIL.n230 12.0247
R165 VTAIL.n275 VTAIL.n212 12.0247
R166 VTAIL.n29 VTAIL.n20 12.0247
R167 VTAIL.n65 VTAIL.n2 12.0247
R168 VTAIL.n205 VTAIL.n142 12.0247
R169 VTAIL.n169 VTAIL.n160 12.0247
R170 VTAIL.n135 VTAIL.n72 12.0247
R171 VTAIL.n99 VTAIL.n90 12.0247
R172 VTAIL.n240 VTAIL.n228 11.249
R173 VTAIL.n272 VTAIL.n271 11.249
R174 VTAIL.n30 VTAIL.n18 11.249
R175 VTAIL.n62 VTAIL.n61 11.249
R176 VTAIL.n202 VTAIL.n201 11.249
R177 VTAIL.n170 VTAIL.n158 11.249
R178 VTAIL.n132 VTAIL.n131 11.249
R179 VTAIL.n100 VTAIL.n88 11.249
R180 VTAIL.n244 VTAIL.n243 10.4732
R181 VTAIL.n268 VTAIL.n214 10.4732
R182 VTAIL.n34 VTAIL.n33 10.4732
R183 VTAIL.n58 VTAIL.n4 10.4732
R184 VTAIL.n198 VTAIL.n144 10.4732
R185 VTAIL.n174 VTAIL.n173 10.4732
R186 VTAIL.n128 VTAIL.n74 10.4732
R187 VTAIL.n104 VTAIL.n103 10.4732
R188 VTAIL.n247 VTAIL.n226 9.69747
R189 VTAIL.n267 VTAIL.n216 9.69747
R190 VTAIL.n37 VTAIL.n16 9.69747
R191 VTAIL.n57 VTAIL.n6 9.69747
R192 VTAIL.n197 VTAIL.n146 9.69747
R193 VTAIL.n177 VTAIL.n156 9.69747
R194 VTAIL.n127 VTAIL.n76 9.69747
R195 VTAIL.n107 VTAIL.n86 9.69747
R196 VTAIL.n274 VTAIL.n210 9.45567
R197 VTAIL.n64 VTAIL.n0 9.45567
R198 VTAIL.n204 VTAIL.n140 9.45567
R199 VTAIL.n134 VTAIL.n70 9.45567
R200 VTAIL.n257 VTAIL.n256 9.3005
R201 VTAIL.n259 VTAIL.n258 9.3005
R202 VTAIL.n218 VTAIL.n217 9.3005
R203 VTAIL.n265 VTAIL.n264 9.3005
R204 VTAIL.n267 VTAIL.n266 9.3005
R205 VTAIL.n214 VTAIL.n213 9.3005
R206 VTAIL.n273 VTAIL.n272 9.3005
R207 VTAIL.n275 VTAIL.n274 9.3005
R208 VTAIL.n251 VTAIL.n250 9.3005
R209 VTAIL.n249 VTAIL.n248 9.3005
R210 VTAIL.n226 VTAIL.n225 9.3005
R211 VTAIL.n243 VTAIL.n242 9.3005
R212 VTAIL.n241 VTAIL.n240 9.3005
R213 VTAIL.n230 VTAIL.n229 9.3005
R214 VTAIL.n235 VTAIL.n234 9.3005
R215 VTAIL.n222 VTAIL.n221 9.3005
R216 VTAIL.n47 VTAIL.n46 9.3005
R217 VTAIL.n49 VTAIL.n48 9.3005
R218 VTAIL.n8 VTAIL.n7 9.3005
R219 VTAIL.n55 VTAIL.n54 9.3005
R220 VTAIL.n57 VTAIL.n56 9.3005
R221 VTAIL.n4 VTAIL.n3 9.3005
R222 VTAIL.n63 VTAIL.n62 9.3005
R223 VTAIL.n65 VTAIL.n64 9.3005
R224 VTAIL.n41 VTAIL.n40 9.3005
R225 VTAIL.n39 VTAIL.n38 9.3005
R226 VTAIL.n16 VTAIL.n15 9.3005
R227 VTAIL.n33 VTAIL.n32 9.3005
R228 VTAIL.n31 VTAIL.n30 9.3005
R229 VTAIL.n20 VTAIL.n19 9.3005
R230 VTAIL.n25 VTAIL.n24 9.3005
R231 VTAIL.n12 VTAIL.n11 9.3005
R232 VTAIL.n205 VTAIL.n204 9.3005
R233 VTAIL.n203 VTAIL.n202 9.3005
R234 VTAIL.n144 VTAIL.n143 9.3005
R235 VTAIL.n197 VTAIL.n196 9.3005
R236 VTAIL.n195 VTAIL.n194 9.3005
R237 VTAIL.n148 VTAIL.n147 9.3005
R238 VTAIL.n189 VTAIL.n188 9.3005
R239 VTAIL.n187 VTAIL.n186 9.3005
R240 VTAIL.n152 VTAIL.n151 9.3005
R241 VTAIL.n181 VTAIL.n180 9.3005
R242 VTAIL.n179 VTAIL.n178 9.3005
R243 VTAIL.n156 VTAIL.n155 9.3005
R244 VTAIL.n173 VTAIL.n172 9.3005
R245 VTAIL.n171 VTAIL.n170 9.3005
R246 VTAIL.n160 VTAIL.n159 9.3005
R247 VTAIL.n165 VTAIL.n164 9.3005
R248 VTAIL.n119 VTAIL.n118 9.3005
R249 VTAIL.n78 VTAIL.n77 9.3005
R250 VTAIL.n125 VTAIL.n124 9.3005
R251 VTAIL.n127 VTAIL.n126 9.3005
R252 VTAIL.n74 VTAIL.n73 9.3005
R253 VTAIL.n133 VTAIL.n132 9.3005
R254 VTAIL.n135 VTAIL.n134 9.3005
R255 VTAIL.n117 VTAIL.n116 9.3005
R256 VTAIL.n82 VTAIL.n81 9.3005
R257 VTAIL.n111 VTAIL.n110 9.3005
R258 VTAIL.n109 VTAIL.n108 9.3005
R259 VTAIL.n86 VTAIL.n85 9.3005
R260 VTAIL.n103 VTAIL.n102 9.3005
R261 VTAIL.n101 VTAIL.n100 9.3005
R262 VTAIL.n90 VTAIL.n89 9.3005
R263 VTAIL.n95 VTAIL.n94 9.3005
R264 VTAIL.n248 VTAIL.n224 8.92171
R265 VTAIL.n264 VTAIL.n263 8.92171
R266 VTAIL.n38 VTAIL.n14 8.92171
R267 VTAIL.n54 VTAIL.n53 8.92171
R268 VTAIL.n194 VTAIL.n193 8.92171
R269 VTAIL.n178 VTAIL.n154 8.92171
R270 VTAIL.n124 VTAIL.n123 8.92171
R271 VTAIL.n108 VTAIL.n84 8.92171
R272 VTAIL.n252 VTAIL.n251 8.14595
R273 VTAIL.n260 VTAIL.n218 8.14595
R274 VTAIL.n42 VTAIL.n41 8.14595
R275 VTAIL.n50 VTAIL.n8 8.14595
R276 VTAIL.n190 VTAIL.n148 8.14595
R277 VTAIL.n182 VTAIL.n181 8.14595
R278 VTAIL.n120 VTAIL.n78 8.14595
R279 VTAIL.n112 VTAIL.n111 8.14595
R280 VTAIL.n255 VTAIL.n222 7.3702
R281 VTAIL.n259 VTAIL.n220 7.3702
R282 VTAIL.n45 VTAIL.n12 7.3702
R283 VTAIL.n49 VTAIL.n10 7.3702
R284 VTAIL.n189 VTAIL.n150 7.3702
R285 VTAIL.n185 VTAIL.n152 7.3702
R286 VTAIL.n119 VTAIL.n80 7.3702
R287 VTAIL.n115 VTAIL.n82 7.3702
R288 VTAIL.n256 VTAIL.n255 6.59444
R289 VTAIL.n256 VTAIL.n220 6.59444
R290 VTAIL.n46 VTAIL.n45 6.59444
R291 VTAIL.n46 VTAIL.n10 6.59444
R292 VTAIL.n186 VTAIL.n150 6.59444
R293 VTAIL.n186 VTAIL.n185 6.59444
R294 VTAIL.n116 VTAIL.n80 6.59444
R295 VTAIL.n116 VTAIL.n115 6.59444
R296 VTAIL.n252 VTAIL.n222 5.81868
R297 VTAIL.n260 VTAIL.n259 5.81868
R298 VTAIL.n42 VTAIL.n12 5.81868
R299 VTAIL.n50 VTAIL.n49 5.81868
R300 VTAIL.n190 VTAIL.n189 5.81868
R301 VTAIL.n182 VTAIL.n152 5.81868
R302 VTAIL.n120 VTAIL.n119 5.81868
R303 VTAIL.n112 VTAIL.n82 5.81868
R304 VTAIL.n251 VTAIL.n224 5.04292
R305 VTAIL.n263 VTAIL.n218 5.04292
R306 VTAIL.n41 VTAIL.n14 5.04292
R307 VTAIL.n53 VTAIL.n8 5.04292
R308 VTAIL.n193 VTAIL.n148 5.04292
R309 VTAIL.n181 VTAIL.n154 5.04292
R310 VTAIL.n123 VTAIL.n78 5.04292
R311 VTAIL.n111 VTAIL.n84 5.04292
R312 VTAIL.n248 VTAIL.n247 4.26717
R313 VTAIL.n264 VTAIL.n216 4.26717
R314 VTAIL.n38 VTAIL.n37 4.26717
R315 VTAIL.n54 VTAIL.n6 4.26717
R316 VTAIL.n194 VTAIL.n146 4.26717
R317 VTAIL.n178 VTAIL.n177 4.26717
R318 VTAIL.n124 VTAIL.n76 4.26717
R319 VTAIL.n108 VTAIL.n107 4.26717
R320 VTAIL.n234 VTAIL.n233 3.70982
R321 VTAIL.n24 VTAIL.n23 3.70982
R322 VTAIL.n164 VTAIL.n163 3.70982
R323 VTAIL.n94 VTAIL.n93 3.70982
R324 VTAIL.n244 VTAIL.n226 3.49141
R325 VTAIL.n268 VTAIL.n267 3.49141
R326 VTAIL.n34 VTAIL.n16 3.49141
R327 VTAIL.n58 VTAIL.n57 3.49141
R328 VTAIL.n198 VTAIL.n197 3.49141
R329 VTAIL.n174 VTAIL.n156 3.49141
R330 VTAIL.n128 VTAIL.n127 3.49141
R331 VTAIL.n104 VTAIL.n86 3.49141
R332 VTAIL.n243 VTAIL.n228 2.71565
R333 VTAIL.n271 VTAIL.n214 2.71565
R334 VTAIL.n33 VTAIL.n18 2.71565
R335 VTAIL.n61 VTAIL.n4 2.71565
R336 VTAIL.n201 VTAIL.n144 2.71565
R337 VTAIL.n173 VTAIL.n158 2.71565
R338 VTAIL.n131 VTAIL.n74 2.71565
R339 VTAIL.n103 VTAIL.n88 2.71565
R340 VTAIL.n240 VTAIL.n239 1.93989
R341 VTAIL.n272 VTAIL.n212 1.93989
R342 VTAIL.n30 VTAIL.n29 1.93989
R343 VTAIL.n62 VTAIL.n2 1.93989
R344 VTAIL.n202 VTAIL.n142 1.93989
R345 VTAIL.n170 VTAIL.n169 1.93989
R346 VTAIL.n132 VTAIL.n72 1.93989
R347 VTAIL.n100 VTAIL.n99 1.93989
R348 VTAIL.n209 VTAIL.n139 1.48757
R349 VTAIL.n236 VTAIL.n230 1.16414
R350 VTAIL.n276 VTAIL.n275 1.16414
R351 VTAIL.n26 VTAIL.n20 1.16414
R352 VTAIL.n66 VTAIL.n65 1.16414
R353 VTAIL.n206 VTAIL.n205 1.16414
R354 VTAIL.n166 VTAIL.n160 1.16414
R355 VTAIL.n136 VTAIL.n135 1.16414
R356 VTAIL.n96 VTAIL.n90 1.16414
R357 VTAIL VTAIL.n69 1.03714
R358 VTAIL VTAIL.n279 0.450931
R359 VTAIL.n235 VTAIL.n232 0.388379
R360 VTAIL.n278 VTAIL.n210 0.388379
R361 VTAIL.n25 VTAIL.n22 0.388379
R362 VTAIL.n68 VTAIL.n0 0.388379
R363 VTAIL.n208 VTAIL.n140 0.388379
R364 VTAIL.n165 VTAIL.n162 0.388379
R365 VTAIL.n138 VTAIL.n70 0.388379
R366 VTAIL.n95 VTAIL.n92 0.388379
R367 VTAIL.n234 VTAIL.n229 0.155672
R368 VTAIL.n241 VTAIL.n229 0.155672
R369 VTAIL.n242 VTAIL.n241 0.155672
R370 VTAIL.n242 VTAIL.n225 0.155672
R371 VTAIL.n249 VTAIL.n225 0.155672
R372 VTAIL.n250 VTAIL.n249 0.155672
R373 VTAIL.n250 VTAIL.n221 0.155672
R374 VTAIL.n257 VTAIL.n221 0.155672
R375 VTAIL.n258 VTAIL.n257 0.155672
R376 VTAIL.n258 VTAIL.n217 0.155672
R377 VTAIL.n265 VTAIL.n217 0.155672
R378 VTAIL.n266 VTAIL.n265 0.155672
R379 VTAIL.n266 VTAIL.n213 0.155672
R380 VTAIL.n273 VTAIL.n213 0.155672
R381 VTAIL.n274 VTAIL.n273 0.155672
R382 VTAIL.n24 VTAIL.n19 0.155672
R383 VTAIL.n31 VTAIL.n19 0.155672
R384 VTAIL.n32 VTAIL.n31 0.155672
R385 VTAIL.n32 VTAIL.n15 0.155672
R386 VTAIL.n39 VTAIL.n15 0.155672
R387 VTAIL.n40 VTAIL.n39 0.155672
R388 VTAIL.n40 VTAIL.n11 0.155672
R389 VTAIL.n47 VTAIL.n11 0.155672
R390 VTAIL.n48 VTAIL.n47 0.155672
R391 VTAIL.n48 VTAIL.n7 0.155672
R392 VTAIL.n55 VTAIL.n7 0.155672
R393 VTAIL.n56 VTAIL.n55 0.155672
R394 VTAIL.n56 VTAIL.n3 0.155672
R395 VTAIL.n63 VTAIL.n3 0.155672
R396 VTAIL.n64 VTAIL.n63 0.155672
R397 VTAIL.n204 VTAIL.n203 0.155672
R398 VTAIL.n203 VTAIL.n143 0.155672
R399 VTAIL.n196 VTAIL.n143 0.155672
R400 VTAIL.n196 VTAIL.n195 0.155672
R401 VTAIL.n195 VTAIL.n147 0.155672
R402 VTAIL.n188 VTAIL.n147 0.155672
R403 VTAIL.n188 VTAIL.n187 0.155672
R404 VTAIL.n187 VTAIL.n151 0.155672
R405 VTAIL.n180 VTAIL.n151 0.155672
R406 VTAIL.n180 VTAIL.n179 0.155672
R407 VTAIL.n179 VTAIL.n155 0.155672
R408 VTAIL.n172 VTAIL.n155 0.155672
R409 VTAIL.n172 VTAIL.n171 0.155672
R410 VTAIL.n171 VTAIL.n159 0.155672
R411 VTAIL.n164 VTAIL.n159 0.155672
R412 VTAIL.n134 VTAIL.n133 0.155672
R413 VTAIL.n133 VTAIL.n73 0.155672
R414 VTAIL.n126 VTAIL.n73 0.155672
R415 VTAIL.n126 VTAIL.n125 0.155672
R416 VTAIL.n125 VTAIL.n77 0.155672
R417 VTAIL.n118 VTAIL.n77 0.155672
R418 VTAIL.n118 VTAIL.n117 0.155672
R419 VTAIL.n117 VTAIL.n81 0.155672
R420 VTAIL.n110 VTAIL.n81 0.155672
R421 VTAIL.n110 VTAIL.n109 0.155672
R422 VTAIL.n109 VTAIL.n85 0.155672
R423 VTAIL.n102 VTAIL.n85 0.155672
R424 VTAIL.n102 VTAIL.n101 0.155672
R425 VTAIL.n101 VTAIL.n89 0.155672
R426 VTAIL.n94 VTAIL.n89 0.155672
R427 VDD2.n137 VDD2.n136 756.745
R428 VDD2.n68 VDD2.n67 756.745
R429 VDD2.n136 VDD2.n135 585
R430 VDD2.n71 VDD2.n70 585
R431 VDD2.n130 VDD2.n129 585
R432 VDD2.n128 VDD2.n127 585
R433 VDD2.n75 VDD2.n74 585
R434 VDD2.n122 VDD2.n121 585
R435 VDD2.n120 VDD2.n119 585
R436 VDD2.n79 VDD2.n78 585
R437 VDD2.n114 VDD2.n113 585
R438 VDD2.n112 VDD2.n111 585
R439 VDD2.n83 VDD2.n82 585
R440 VDD2.n106 VDD2.n105 585
R441 VDD2.n104 VDD2.n103 585
R442 VDD2.n87 VDD2.n86 585
R443 VDD2.n98 VDD2.n97 585
R444 VDD2.n96 VDD2.n95 585
R445 VDD2.n91 VDD2.n90 585
R446 VDD2.n22 VDD2.n21 585
R447 VDD2.n27 VDD2.n26 585
R448 VDD2.n29 VDD2.n28 585
R449 VDD2.n18 VDD2.n17 585
R450 VDD2.n35 VDD2.n34 585
R451 VDD2.n37 VDD2.n36 585
R452 VDD2.n14 VDD2.n13 585
R453 VDD2.n43 VDD2.n42 585
R454 VDD2.n45 VDD2.n44 585
R455 VDD2.n10 VDD2.n9 585
R456 VDD2.n51 VDD2.n50 585
R457 VDD2.n53 VDD2.n52 585
R458 VDD2.n6 VDD2.n5 585
R459 VDD2.n59 VDD2.n58 585
R460 VDD2.n61 VDD2.n60 585
R461 VDD2.n2 VDD2.n1 585
R462 VDD2.n67 VDD2.n66 585
R463 VDD2.n92 VDD2.t0 327.466
R464 VDD2.n23 VDD2.t1 327.466
R465 VDD2.n136 VDD2.n70 171.744
R466 VDD2.n129 VDD2.n70 171.744
R467 VDD2.n129 VDD2.n128 171.744
R468 VDD2.n128 VDD2.n74 171.744
R469 VDD2.n121 VDD2.n74 171.744
R470 VDD2.n121 VDD2.n120 171.744
R471 VDD2.n120 VDD2.n78 171.744
R472 VDD2.n113 VDD2.n78 171.744
R473 VDD2.n113 VDD2.n112 171.744
R474 VDD2.n112 VDD2.n82 171.744
R475 VDD2.n105 VDD2.n82 171.744
R476 VDD2.n105 VDD2.n104 171.744
R477 VDD2.n104 VDD2.n86 171.744
R478 VDD2.n97 VDD2.n86 171.744
R479 VDD2.n97 VDD2.n96 171.744
R480 VDD2.n96 VDD2.n90 171.744
R481 VDD2.n27 VDD2.n21 171.744
R482 VDD2.n28 VDD2.n27 171.744
R483 VDD2.n28 VDD2.n17 171.744
R484 VDD2.n35 VDD2.n17 171.744
R485 VDD2.n36 VDD2.n35 171.744
R486 VDD2.n36 VDD2.n13 171.744
R487 VDD2.n43 VDD2.n13 171.744
R488 VDD2.n44 VDD2.n43 171.744
R489 VDD2.n44 VDD2.n9 171.744
R490 VDD2.n51 VDD2.n9 171.744
R491 VDD2.n52 VDD2.n51 171.744
R492 VDD2.n52 VDD2.n5 171.744
R493 VDD2.n59 VDD2.n5 171.744
R494 VDD2.n60 VDD2.n59 171.744
R495 VDD2.n60 VDD2.n1 171.744
R496 VDD2.n67 VDD2.n1 171.744
R497 VDD2.n138 VDD2.n68 90.6094
R498 VDD2.t0 VDD2.n90 85.8723
R499 VDD2.t1 VDD2.n21 85.8723
R500 VDD2.n138 VDD2.n137 51.9672
R501 VDD2.n92 VDD2.n91 16.3895
R502 VDD2.n23 VDD2.n22 16.3895
R503 VDD2.n135 VDD2.n69 12.8005
R504 VDD2.n95 VDD2.n94 12.8005
R505 VDD2.n26 VDD2.n25 12.8005
R506 VDD2.n66 VDD2.n0 12.8005
R507 VDD2.n134 VDD2.n71 12.0247
R508 VDD2.n98 VDD2.n89 12.0247
R509 VDD2.n29 VDD2.n20 12.0247
R510 VDD2.n65 VDD2.n2 12.0247
R511 VDD2.n131 VDD2.n130 11.249
R512 VDD2.n99 VDD2.n87 11.249
R513 VDD2.n30 VDD2.n18 11.249
R514 VDD2.n62 VDD2.n61 11.249
R515 VDD2.n127 VDD2.n73 10.4732
R516 VDD2.n103 VDD2.n102 10.4732
R517 VDD2.n34 VDD2.n33 10.4732
R518 VDD2.n58 VDD2.n4 10.4732
R519 VDD2.n126 VDD2.n75 9.69747
R520 VDD2.n106 VDD2.n85 9.69747
R521 VDD2.n37 VDD2.n16 9.69747
R522 VDD2.n57 VDD2.n6 9.69747
R523 VDD2.n133 VDD2.n69 9.45567
R524 VDD2.n64 VDD2.n0 9.45567
R525 VDD2.n134 VDD2.n133 9.3005
R526 VDD2.n132 VDD2.n131 9.3005
R527 VDD2.n73 VDD2.n72 9.3005
R528 VDD2.n126 VDD2.n125 9.3005
R529 VDD2.n124 VDD2.n123 9.3005
R530 VDD2.n77 VDD2.n76 9.3005
R531 VDD2.n118 VDD2.n117 9.3005
R532 VDD2.n116 VDD2.n115 9.3005
R533 VDD2.n81 VDD2.n80 9.3005
R534 VDD2.n110 VDD2.n109 9.3005
R535 VDD2.n108 VDD2.n107 9.3005
R536 VDD2.n85 VDD2.n84 9.3005
R537 VDD2.n102 VDD2.n101 9.3005
R538 VDD2.n100 VDD2.n99 9.3005
R539 VDD2.n89 VDD2.n88 9.3005
R540 VDD2.n94 VDD2.n93 9.3005
R541 VDD2.n47 VDD2.n46 9.3005
R542 VDD2.n49 VDD2.n48 9.3005
R543 VDD2.n8 VDD2.n7 9.3005
R544 VDD2.n55 VDD2.n54 9.3005
R545 VDD2.n57 VDD2.n56 9.3005
R546 VDD2.n4 VDD2.n3 9.3005
R547 VDD2.n63 VDD2.n62 9.3005
R548 VDD2.n65 VDD2.n64 9.3005
R549 VDD2.n41 VDD2.n40 9.3005
R550 VDD2.n39 VDD2.n38 9.3005
R551 VDD2.n16 VDD2.n15 9.3005
R552 VDD2.n33 VDD2.n32 9.3005
R553 VDD2.n31 VDD2.n30 9.3005
R554 VDD2.n20 VDD2.n19 9.3005
R555 VDD2.n25 VDD2.n24 9.3005
R556 VDD2.n12 VDD2.n11 9.3005
R557 VDD2.n123 VDD2.n122 8.92171
R558 VDD2.n107 VDD2.n83 8.92171
R559 VDD2.n38 VDD2.n14 8.92171
R560 VDD2.n54 VDD2.n53 8.92171
R561 VDD2.n119 VDD2.n77 8.14595
R562 VDD2.n111 VDD2.n110 8.14595
R563 VDD2.n42 VDD2.n41 8.14595
R564 VDD2.n50 VDD2.n8 8.14595
R565 VDD2.n118 VDD2.n79 7.3702
R566 VDD2.n114 VDD2.n81 7.3702
R567 VDD2.n45 VDD2.n12 7.3702
R568 VDD2.n49 VDD2.n10 7.3702
R569 VDD2.n115 VDD2.n79 6.59444
R570 VDD2.n115 VDD2.n114 6.59444
R571 VDD2.n46 VDD2.n45 6.59444
R572 VDD2.n46 VDD2.n10 6.59444
R573 VDD2.n119 VDD2.n118 5.81868
R574 VDD2.n111 VDD2.n81 5.81868
R575 VDD2.n42 VDD2.n12 5.81868
R576 VDD2.n50 VDD2.n49 5.81868
R577 VDD2.n122 VDD2.n77 5.04292
R578 VDD2.n110 VDD2.n83 5.04292
R579 VDD2.n41 VDD2.n14 5.04292
R580 VDD2.n53 VDD2.n8 5.04292
R581 VDD2.n123 VDD2.n75 4.26717
R582 VDD2.n107 VDD2.n106 4.26717
R583 VDD2.n38 VDD2.n37 4.26717
R584 VDD2.n54 VDD2.n6 4.26717
R585 VDD2.n93 VDD2.n92 3.70982
R586 VDD2.n24 VDD2.n23 3.70982
R587 VDD2.n127 VDD2.n126 3.49141
R588 VDD2.n103 VDD2.n85 3.49141
R589 VDD2.n34 VDD2.n16 3.49141
R590 VDD2.n58 VDD2.n57 3.49141
R591 VDD2.n130 VDD2.n73 2.71565
R592 VDD2.n102 VDD2.n87 2.71565
R593 VDD2.n33 VDD2.n18 2.71565
R594 VDD2.n61 VDD2.n4 2.71565
R595 VDD2.n131 VDD2.n71 1.93989
R596 VDD2.n99 VDD2.n98 1.93989
R597 VDD2.n30 VDD2.n29 1.93989
R598 VDD2.n62 VDD2.n2 1.93989
R599 VDD2.n135 VDD2.n134 1.16414
R600 VDD2.n95 VDD2.n89 1.16414
R601 VDD2.n26 VDD2.n20 1.16414
R602 VDD2.n66 VDD2.n65 1.16414
R603 VDD2 VDD2.n138 0.56731
R604 VDD2.n137 VDD2.n69 0.388379
R605 VDD2.n94 VDD2.n91 0.388379
R606 VDD2.n25 VDD2.n22 0.388379
R607 VDD2.n68 VDD2.n0 0.388379
R608 VDD2.n133 VDD2.n132 0.155672
R609 VDD2.n132 VDD2.n72 0.155672
R610 VDD2.n125 VDD2.n72 0.155672
R611 VDD2.n125 VDD2.n124 0.155672
R612 VDD2.n124 VDD2.n76 0.155672
R613 VDD2.n117 VDD2.n76 0.155672
R614 VDD2.n117 VDD2.n116 0.155672
R615 VDD2.n116 VDD2.n80 0.155672
R616 VDD2.n109 VDD2.n80 0.155672
R617 VDD2.n109 VDD2.n108 0.155672
R618 VDD2.n108 VDD2.n84 0.155672
R619 VDD2.n101 VDD2.n84 0.155672
R620 VDD2.n101 VDD2.n100 0.155672
R621 VDD2.n100 VDD2.n88 0.155672
R622 VDD2.n93 VDD2.n88 0.155672
R623 VDD2.n24 VDD2.n19 0.155672
R624 VDD2.n31 VDD2.n19 0.155672
R625 VDD2.n32 VDD2.n31 0.155672
R626 VDD2.n32 VDD2.n15 0.155672
R627 VDD2.n39 VDD2.n15 0.155672
R628 VDD2.n40 VDD2.n39 0.155672
R629 VDD2.n40 VDD2.n11 0.155672
R630 VDD2.n47 VDD2.n11 0.155672
R631 VDD2.n48 VDD2.n47 0.155672
R632 VDD2.n48 VDD2.n7 0.155672
R633 VDD2.n55 VDD2.n7 0.155672
R634 VDD2.n56 VDD2.n55 0.155672
R635 VDD2.n56 VDD2.n3 0.155672
R636 VDD2.n63 VDD2.n3 0.155672
R637 VDD2.n64 VDD2.n63 0.155672
R638 VP.n0 VP.t0 252.829
R639 VP.n0 VP.t1 209.185
R640 VP VP.n0 0.241678
R641 VDD1.n68 VDD1.n67 756.745
R642 VDD1.n137 VDD1.n136 756.745
R643 VDD1.n67 VDD1.n66 585
R644 VDD1.n2 VDD1.n1 585
R645 VDD1.n61 VDD1.n60 585
R646 VDD1.n59 VDD1.n58 585
R647 VDD1.n6 VDD1.n5 585
R648 VDD1.n53 VDD1.n52 585
R649 VDD1.n51 VDD1.n50 585
R650 VDD1.n10 VDD1.n9 585
R651 VDD1.n45 VDD1.n44 585
R652 VDD1.n43 VDD1.n42 585
R653 VDD1.n14 VDD1.n13 585
R654 VDD1.n37 VDD1.n36 585
R655 VDD1.n35 VDD1.n34 585
R656 VDD1.n18 VDD1.n17 585
R657 VDD1.n29 VDD1.n28 585
R658 VDD1.n27 VDD1.n26 585
R659 VDD1.n22 VDD1.n21 585
R660 VDD1.n91 VDD1.n90 585
R661 VDD1.n96 VDD1.n95 585
R662 VDD1.n98 VDD1.n97 585
R663 VDD1.n87 VDD1.n86 585
R664 VDD1.n104 VDD1.n103 585
R665 VDD1.n106 VDD1.n105 585
R666 VDD1.n83 VDD1.n82 585
R667 VDD1.n112 VDD1.n111 585
R668 VDD1.n114 VDD1.n113 585
R669 VDD1.n79 VDD1.n78 585
R670 VDD1.n120 VDD1.n119 585
R671 VDD1.n122 VDD1.n121 585
R672 VDD1.n75 VDD1.n74 585
R673 VDD1.n128 VDD1.n127 585
R674 VDD1.n130 VDD1.n129 585
R675 VDD1.n71 VDD1.n70 585
R676 VDD1.n136 VDD1.n135 585
R677 VDD1.n23 VDD1.t1 327.466
R678 VDD1.n92 VDD1.t0 327.466
R679 VDD1.n67 VDD1.n1 171.744
R680 VDD1.n60 VDD1.n1 171.744
R681 VDD1.n60 VDD1.n59 171.744
R682 VDD1.n59 VDD1.n5 171.744
R683 VDD1.n52 VDD1.n5 171.744
R684 VDD1.n52 VDD1.n51 171.744
R685 VDD1.n51 VDD1.n9 171.744
R686 VDD1.n44 VDD1.n9 171.744
R687 VDD1.n44 VDD1.n43 171.744
R688 VDD1.n43 VDD1.n13 171.744
R689 VDD1.n36 VDD1.n13 171.744
R690 VDD1.n36 VDD1.n35 171.744
R691 VDD1.n35 VDD1.n17 171.744
R692 VDD1.n28 VDD1.n17 171.744
R693 VDD1.n28 VDD1.n27 171.744
R694 VDD1.n27 VDD1.n21 171.744
R695 VDD1.n96 VDD1.n90 171.744
R696 VDD1.n97 VDD1.n96 171.744
R697 VDD1.n97 VDD1.n86 171.744
R698 VDD1.n104 VDD1.n86 171.744
R699 VDD1.n105 VDD1.n104 171.744
R700 VDD1.n105 VDD1.n82 171.744
R701 VDD1.n112 VDD1.n82 171.744
R702 VDD1.n113 VDD1.n112 171.744
R703 VDD1.n113 VDD1.n78 171.744
R704 VDD1.n120 VDD1.n78 171.744
R705 VDD1.n121 VDD1.n120 171.744
R706 VDD1.n121 VDD1.n74 171.744
R707 VDD1.n128 VDD1.n74 171.744
R708 VDD1.n129 VDD1.n128 171.744
R709 VDD1.n129 VDD1.n70 171.744
R710 VDD1.n136 VDD1.n70 171.744
R711 VDD1 VDD1.n137 91.6428
R712 VDD1.t1 VDD1.n21 85.8723
R713 VDD1.t0 VDD1.n90 85.8723
R714 VDD1 VDD1.n68 52.534
R715 VDD1.n23 VDD1.n22 16.3895
R716 VDD1.n92 VDD1.n91 16.3895
R717 VDD1.n66 VDD1.n0 12.8005
R718 VDD1.n26 VDD1.n25 12.8005
R719 VDD1.n95 VDD1.n94 12.8005
R720 VDD1.n135 VDD1.n69 12.8005
R721 VDD1.n65 VDD1.n2 12.0247
R722 VDD1.n29 VDD1.n20 12.0247
R723 VDD1.n98 VDD1.n89 12.0247
R724 VDD1.n134 VDD1.n71 12.0247
R725 VDD1.n62 VDD1.n61 11.249
R726 VDD1.n30 VDD1.n18 11.249
R727 VDD1.n99 VDD1.n87 11.249
R728 VDD1.n131 VDD1.n130 11.249
R729 VDD1.n58 VDD1.n4 10.4732
R730 VDD1.n34 VDD1.n33 10.4732
R731 VDD1.n103 VDD1.n102 10.4732
R732 VDD1.n127 VDD1.n73 10.4732
R733 VDD1.n57 VDD1.n6 9.69747
R734 VDD1.n37 VDD1.n16 9.69747
R735 VDD1.n106 VDD1.n85 9.69747
R736 VDD1.n126 VDD1.n75 9.69747
R737 VDD1.n64 VDD1.n0 9.45567
R738 VDD1.n133 VDD1.n69 9.45567
R739 VDD1.n65 VDD1.n64 9.3005
R740 VDD1.n63 VDD1.n62 9.3005
R741 VDD1.n4 VDD1.n3 9.3005
R742 VDD1.n57 VDD1.n56 9.3005
R743 VDD1.n55 VDD1.n54 9.3005
R744 VDD1.n8 VDD1.n7 9.3005
R745 VDD1.n49 VDD1.n48 9.3005
R746 VDD1.n47 VDD1.n46 9.3005
R747 VDD1.n12 VDD1.n11 9.3005
R748 VDD1.n41 VDD1.n40 9.3005
R749 VDD1.n39 VDD1.n38 9.3005
R750 VDD1.n16 VDD1.n15 9.3005
R751 VDD1.n33 VDD1.n32 9.3005
R752 VDD1.n31 VDD1.n30 9.3005
R753 VDD1.n20 VDD1.n19 9.3005
R754 VDD1.n25 VDD1.n24 9.3005
R755 VDD1.n116 VDD1.n115 9.3005
R756 VDD1.n118 VDD1.n117 9.3005
R757 VDD1.n77 VDD1.n76 9.3005
R758 VDD1.n124 VDD1.n123 9.3005
R759 VDD1.n126 VDD1.n125 9.3005
R760 VDD1.n73 VDD1.n72 9.3005
R761 VDD1.n132 VDD1.n131 9.3005
R762 VDD1.n134 VDD1.n133 9.3005
R763 VDD1.n110 VDD1.n109 9.3005
R764 VDD1.n108 VDD1.n107 9.3005
R765 VDD1.n85 VDD1.n84 9.3005
R766 VDD1.n102 VDD1.n101 9.3005
R767 VDD1.n100 VDD1.n99 9.3005
R768 VDD1.n89 VDD1.n88 9.3005
R769 VDD1.n94 VDD1.n93 9.3005
R770 VDD1.n81 VDD1.n80 9.3005
R771 VDD1.n54 VDD1.n53 8.92171
R772 VDD1.n38 VDD1.n14 8.92171
R773 VDD1.n107 VDD1.n83 8.92171
R774 VDD1.n123 VDD1.n122 8.92171
R775 VDD1.n50 VDD1.n8 8.14595
R776 VDD1.n42 VDD1.n41 8.14595
R777 VDD1.n111 VDD1.n110 8.14595
R778 VDD1.n119 VDD1.n77 8.14595
R779 VDD1.n49 VDD1.n10 7.3702
R780 VDD1.n45 VDD1.n12 7.3702
R781 VDD1.n114 VDD1.n81 7.3702
R782 VDD1.n118 VDD1.n79 7.3702
R783 VDD1.n46 VDD1.n10 6.59444
R784 VDD1.n46 VDD1.n45 6.59444
R785 VDD1.n115 VDD1.n114 6.59444
R786 VDD1.n115 VDD1.n79 6.59444
R787 VDD1.n50 VDD1.n49 5.81868
R788 VDD1.n42 VDD1.n12 5.81868
R789 VDD1.n111 VDD1.n81 5.81868
R790 VDD1.n119 VDD1.n118 5.81868
R791 VDD1.n53 VDD1.n8 5.04292
R792 VDD1.n41 VDD1.n14 5.04292
R793 VDD1.n110 VDD1.n83 5.04292
R794 VDD1.n122 VDD1.n77 5.04292
R795 VDD1.n54 VDD1.n6 4.26717
R796 VDD1.n38 VDD1.n37 4.26717
R797 VDD1.n107 VDD1.n106 4.26717
R798 VDD1.n123 VDD1.n75 4.26717
R799 VDD1.n24 VDD1.n23 3.70982
R800 VDD1.n93 VDD1.n92 3.70982
R801 VDD1.n58 VDD1.n57 3.49141
R802 VDD1.n34 VDD1.n16 3.49141
R803 VDD1.n103 VDD1.n85 3.49141
R804 VDD1.n127 VDD1.n126 3.49141
R805 VDD1.n61 VDD1.n4 2.71565
R806 VDD1.n33 VDD1.n18 2.71565
R807 VDD1.n102 VDD1.n87 2.71565
R808 VDD1.n130 VDD1.n73 2.71565
R809 VDD1.n62 VDD1.n2 1.93989
R810 VDD1.n30 VDD1.n29 1.93989
R811 VDD1.n99 VDD1.n98 1.93989
R812 VDD1.n131 VDD1.n71 1.93989
R813 VDD1.n66 VDD1.n65 1.16414
R814 VDD1.n26 VDD1.n20 1.16414
R815 VDD1.n95 VDD1.n89 1.16414
R816 VDD1.n135 VDD1.n134 1.16414
R817 VDD1.n68 VDD1.n0 0.388379
R818 VDD1.n25 VDD1.n22 0.388379
R819 VDD1.n94 VDD1.n91 0.388379
R820 VDD1.n137 VDD1.n69 0.388379
R821 VDD1.n64 VDD1.n63 0.155672
R822 VDD1.n63 VDD1.n3 0.155672
R823 VDD1.n56 VDD1.n3 0.155672
R824 VDD1.n56 VDD1.n55 0.155672
R825 VDD1.n55 VDD1.n7 0.155672
R826 VDD1.n48 VDD1.n7 0.155672
R827 VDD1.n48 VDD1.n47 0.155672
R828 VDD1.n47 VDD1.n11 0.155672
R829 VDD1.n40 VDD1.n11 0.155672
R830 VDD1.n40 VDD1.n39 0.155672
R831 VDD1.n39 VDD1.n15 0.155672
R832 VDD1.n32 VDD1.n15 0.155672
R833 VDD1.n32 VDD1.n31 0.155672
R834 VDD1.n31 VDD1.n19 0.155672
R835 VDD1.n24 VDD1.n19 0.155672
R836 VDD1.n93 VDD1.n88 0.155672
R837 VDD1.n100 VDD1.n88 0.155672
R838 VDD1.n101 VDD1.n100 0.155672
R839 VDD1.n101 VDD1.n84 0.155672
R840 VDD1.n108 VDD1.n84 0.155672
R841 VDD1.n109 VDD1.n108 0.155672
R842 VDD1.n109 VDD1.n80 0.155672
R843 VDD1.n116 VDD1.n80 0.155672
R844 VDD1.n117 VDD1.n116 0.155672
R845 VDD1.n117 VDD1.n76 0.155672
R846 VDD1.n124 VDD1.n76 0.155672
R847 VDD1.n125 VDD1.n124 0.155672
R848 VDD1.n125 VDD1.n72 0.155672
R849 VDD1.n132 VDD1.n72 0.155672
R850 VDD1.n133 VDD1.n132 0.155672
R851 B.n398 B.n65 585
R852 B.n400 B.n399 585
R853 B.n401 B.n64 585
R854 B.n403 B.n402 585
R855 B.n404 B.n63 585
R856 B.n406 B.n405 585
R857 B.n407 B.n62 585
R858 B.n409 B.n408 585
R859 B.n410 B.n61 585
R860 B.n412 B.n411 585
R861 B.n413 B.n60 585
R862 B.n415 B.n414 585
R863 B.n416 B.n59 585
R864 B.n418 B.n417 585
R865 B.n419 B.n58 585
R866 B.n421 B.n420 585
R867 B.n422 B.n57 585
R868 B.n424 B.n423 585
R869 B.n425 B.n56 585
R870 B.n427 B.n426 585
R871 B.n428 B.n55 585
R872 B.n430 B.n429 585
R873 B.n431 B.n54 585
R874 B.n433 B.n432 585
R875 B.n434 B.n53 585
R876 B.n436 B.n435 585
R877 B.n437 B.n52 585
R878 B.n439 B.n438 585
R879 B.n440 B.n51 585
R880 B.n442 B.n441 585
R881 B.n443 B.n50 585
R882 B.n445 B.n444 585
R883 B.n446 B.n49 585
R884 B.n448 B.n447 585
R885 B.n449 B.n48 585
R886 B.n451 B.n450 585
R887 B.n452 B.n47 585
R888 B.n454 B.n453 585
R889 B.n455 B.n46 585
R890 B.n457 B.n456 585
R891 B.n458 B.n45 585
R892 B.n460 B.n459 585
R893 B.n461 B.n44 585
R894 B.n463 B.n462 585
R895 B.n465 B.n41 585
R896 B.n467 B.n466 585
R897 B.n468 B.n40 585
R898 B.n470 B.n469 585
R899 B.n471 B.n39 585
R900 B.n473 B.n472 585
R901 B.n474 B.n38 585
R902 B.n476 B.n475 585
R903 B.n477 B.n35 585
R904 B.n480 B.n479 585
R905 B.n481 B.n34 585
R906 B.n483 B.n482 585
R907 B.n484 B.n33 585
R908 B.n486 B.n485 585
R909 B.n487 B.n32 585
R910 B.n489 B.n488 585
R911 B.n490 B.n31 585
R912 B.n492 B.n491 585
R913 B.n493 B.n30 585
R914 B.n495 B.n494 585
R915 B.n496 B.n29 585
R916 B.n498 B.n497 585
R917 B.n499 B.n28 585
R918 B.n501 B.n500 585
R919 B.n502 B.n27 585
R920 B.n504 B.n503 585
R921 B.n505 B.n26 585
R922 B.n507 B.n506 585
R923 B.n508 B.n25 585
R924 B.n510 B.n509 585
R925 B.n511 B.n24 585
R926 B.n513 B.n512 585
R927 B.n514 B.n23 585
R928 B.n516 B.n515 585
R929 B.n517 B.n22 585
R930 B.n519 B.n518 585
R931 B.n520 B.n21 585
R932 B.n522 B.n521 585
R933 B.n523 B.n20 585
R934 B.n525 B.n524 585
R935 B.n526 B.n19 585
R936 B.n528 B.n527 585
R937 B.n529 B.n18 585
R938 B.n531 B.n530 585
R939 B.n532 B.n17 585
R940 B.n534 B.n533 585
R941 B.n535 B.n16 585
R942 B.n537 B.n536 585
R943 B.n538 B.n15 585
R944 B.n540 B.n539 585
R945 B.n541 B.n14 585
R946 B.n543 B.n542 585
R947 B.n544 B.n13 585
R948 B.n397 B.n396 585
R949 B.n395 B.n66 585
R950 B.n394 B.n393 585
R951 B.n392 B.n67 585
R952 B.n391 B.n390 585
R953 B.n389 B.n68 585
R954 B.n388 B.n387 585
R955 B.n386 B.n69 585
R956 B.n385 B.n384 585
R957 B.n383 B.n70 585
R958 B.n382 B.n381 585
R959 B.n380 B.n71 585
R960 B.n379 B.n378 585
R961 B.n377 B.n72 585
R962 B.n376 B.n375 585
R963 B.n374 B.n73 585
R964 B.n373 B.n372 585
R965 B.n371 B.n74 585
R966 B.n370 B.n369 585
R967 B.n368 B.n75 585
R968 B.n367 B.n366 585
R969 B.n365 B.n76 585
R970 B.n364 B.n363 585
R971 B.n362 B.n77 585
R972 B.n361 B.n360 585
R973 B.n359 B.n78 585
R974 B.n358 B.n357 585
R975 B.n356 B.n79 585
R976 B.n355 B.n354 585
R977 B.n353 B.n80 585
R978 B.n352 B.n351 585
R979 B.n350 B.n81 585
R980 B.n349 B.n348 585
R981 B.n347 B.n82 585
R982 B.n346 B.n345 585
R983 B.n344 B.n83 585
R984 B.n343 B.n342 585
R985 B.n341 B.n84 585
R986 B.n340 B.n339 585
R987 B.n338 B.n85 585
R988 B.n337 B.n336 585
R989 B.n335 B.n86 585
R990 B.n334 B.n333 585
R991 B.n332 B.n87 585
R992 B.n331 B.n330 585
R993 B.n184 B.n183 585
R994 B.n185 B.n140 585
R995 B.n187 B.n186 585
R996 B.n188 B.n139 585
R997 B.n190 B.n189 585
R998 B.n191 B.n138 585
R999 B.n193 B.n192 585
R1000 B.n194 B.n137 585
R1001 B.n196 B.n195 585
R1002 B.n197 B.n136 585
R1003 B.n199 B.n198 585
R1004 B.n200 B.n135 585
R1005 B.n202 B.n201 585
R1006 B.n203 B.n134 585
R1007 B.n205 B.n204 585
R1008 B.n206 B.n133 585
R1009 B.n208 B.n207 585
R1010 B.n209 B.n132 585
R1011 B.n211 B.n210 585
R1012 B.n212 B.n131 585
R1013 B.n214 B.n213 585
R1014 B.n215 B.n130 585
R1015 B.n217 B.n216 585
R1016 B.n218 B.n129 585
R1017 B.n220 B.n219 585
R1018 B.n221 B.n128 585
R1019 B.n223 B.n222 585
R1020 B.n224 B.n127 585
R1021 B.n226 B.n225 585
R1022 B.n227 B.n126 585
R1023 B.n229 B.n228 585
R1024 B.n230 B.n125 585
R1025 B.n232 B.n231 585
R1026 B.n233 B.n124 585
R1027 B.n235 B.n234 585
R1028 B.n236 B.n123 585
R1029 B.n238 B.n237 585
R1030 B.n239 B.n122 585
R1031 B.n241 B.n240 585
R1032 B.n242 B.n121 585
R1033 B.n244 B.n243 585
R1034 B.n245 B.n120 585
R1035 B.n247 B.n246 585
R1036 B.n248 B.n117 585
R1037 B.n251 B.n250 585
R1038 B.n252 B.n116 585
R1039 B.n254 B.n253 585
R1040 B.n255 B.n115 585
R1041 B.n257 B.n256 585
R1042 B.n258 B.n114 585
R1043 B.n260 B.n259 585
R1044 B.n261 B.n113 585
R1045 B.n263 B.n262 585
R1046 B.n265 B.n264 585
R1047 B.n266 B.n109 585
R1048 B.n268 B.n267 585
R1049 B.n269 B.n108 585
R1050 B.n271 B.n270 585
R1051 B.n272 B.n107 585
R1052 B.n274 B.n273 585
R1053 B.n275 B.n106 585
R1054 B.n277 B.n276 585
R1055 B.n278 B.n105 585
R1056 B.n280 B.n279 585
R1057 B.n281 B.n104 585
R1058 B.n283 B.n282 585
R1059 B.n284 B.n103 585
R1060 B.n286 B.n285 585
R1061 B.n287 B.n102 585
R1062 B.n289 B.n288 585
R1063 B.n290 B.n101 585
R1064 B.n292 B.n291 585
R1065 B.n293 B.n100 585
R1066 B.n295 B.n294 585
R1067 B.n296 B.n99 585
R1068 B.n298 B.n297 585
R1069 B.n299 B.n98 585
R1070 B.n301 B.n300 585
R1071 B.n302 B.n97 585
R1072 B.n304 B.n303 585
R1073 B.n305 B.n96 585
R1074 B.n307 B.n306 585
R1075 B.n308 B.n95 585
R1076 B.n310 B.n309 585
R1077 B.n311 B.n94 585
R1078 B.n313 B.n312 585
R1079 B.n314 B.n93 585
R1080 B.n316 B.n315 585
R1081 B.n317 B.n92 585
R1082 B.n319 B.n318 585
R1083 B.n320 B.n91 585
R1084 B.n322 B.n321 585
R1085 B.n323 B.n90 585
R1086 B.n325 B.n324 585
R1087 B.n326 B.n89 585
R1088 B.n328 B.n327 585
R1089 B.n329 B.n88 585
R1090 B.n182 B.n141 585
R1091 B.n181 B.n180 585
R1092 B.n179 B.n142 585
R1093 B.n178 B.n177 585
R1094 B.n176 B.n143 585
R1095 B.n175 B.n174 585
R1096 B.n173 B.n144 585
R1097 B.n172 B.n171 585
R1098 B.n170 B.n145 585
R1099 B.n169 B.n168 585
R1100 B.n167 B.n146 585
R1101 B.n166 B.n165 585
R1102 B.n164 B.n147 585
R1103 B.n163 B.n162 585
R1104 B.n161 B.n148 585
R1105 B.n160 B.n159 585
R1106 B.n158 B.n149 585
R1107 B.n157 B.n156 585
R1108 B.n155 B.n150 585
R1109 B.n154 B.n153 585
R1110 B.n152 B.n151 585
R1111 B.n2 B.n0 585
R1112 B.n577 B.n1 585
R1113 B.n576 B.n575 585
R1114 B.n574 B.n3 585
R1115 B.n573 B.n572 585
R1116 B.n571 B.n4 585
R1117 B.n570 B.n569 585
R1118 B.n568 B.n5 585
R1119 B.n567 B.n566 585
R1120 B.n565 B.n6 585
R1121 B.n564 B.n563 585
R1122 B.n562 B.n7 585
R1123 B.n561 B.n560 585
R1124 B.n559 B.n8 585
R1125 B.n558 B.n557 585
R1126 B.n556 B.n9 585
R1127 B.n555 B.n554 585
R1128 B.n553 B.n10 585
R1129 B.n552 B.n551 585
R1130 B.n550 B.n11 585
R1131 B.n549 B.n548 585
R1132 B.n547 B.n12 585
R1133 B.n546 B.n545 585
R1134 B.n579 B.n578 585
R1135 B.n184 B.n141 473.281
R1136 B.n546 B.n13 473.281
R1137 B.n330 B.n329 473.281
R1138 B.n396 B.n65 473.281
R1139 B.n110 B.t8 433.159
R1140 B.n42 B.t1 433.159
R1141 B.n118 B.t5 433.159
R1142 B.n36 B.t10 433.159
R1143 B.n111 B.t7 387.389
R1144 B.n43 B.t2 387.389
R1145 B.n119 B.t4 387.389
R1146 B.n37 B.t11 387.389
R1147 B.n110 B.t6 357.286
R1148 B.n118 B.t3 357.286
R1149 B.n36 B.t9 357.286
R1150 B.n42 B.t0 357.286
R1151 B.n180 B.n141 163.367
R1152 B.n180 B.n179 163.367
R1153 B.n179 B.n178 163.367
R1154 B.n178 B.n143 163.367
R1155 B.n174 B.n143 163.367
R1156 B.n174 B.n173 163.367
R1157 B.n173 B.n172 163.367
R1158 B.n172 B.n145 163.367
R1159 B.n168 B.n145 163.367
R1160 B.n168 B.n167 163.367
R1161 B.n167 B.n166 163.367
R1162 B.n166 B.n147 163.367
R1163 B.n162 B.n147 163.367
R1164 B.n162 B.n161 163.367
R1165 B.n161 B.n160 163.367
R1166 B.n160 B.n149 163.367
R1167 B.n156 B.n149 163.367
R1168 B.n156 B.n155 163.367
R1169 B.n155 B.n154 163.367
R1170 B.n154 B.n151 163.367
R1171 B.n151 B.n2 163.367
R1172 B.n578 B.n2 163.367
R1173 B.n578 B.n577 163.367
R1174 B.n577 B.n576 163.367
R1175 B.n576 B.n3 163.367
R1176 B.n572 B.n3 163.367
R1177 B.n572 B.n571 163.367
R1178 B.n571 B.n570 163.367
R1179 B.n570 B.n5 163.367
R1180 B.n566 B.n5 163.367
R1181 B.n566 B.n565 163.367
R1182 B.n565 B.n564 163.367
R1183 B.n564 B.n7 163.367
R1184 B.n560 B.n7 163.367
R1185 B.n560 B.n559 163.367
R1186 B.n559 B.n558 163.367
R1187 B.n558 B.n9 163.367
R1188 B.n554 B.n9 163.367
R1189 B.n554 B.n553 163.367
R1190 B.n553 B.n552 163.367
R1191 B.n552 B.n11 163.367
R1192 B.n548 B.n11 163.367
R1193 B.n548 B.n547 163.367
R1194 B.n547 B.n546 163.367
R1195 B.n185 B.n184 163.367
R1196 B.n186 B.n185 163.367
R1197 B.n186 B.n139 163.367
R1198 B.n190 B.n139 163.367
R1199 B.n191 B.n190 163.367
R1200 B.n192 B.n191 163.367
R1201 B.n192 B.n137 163.367
R1202 B.n196 B.n137 163.367
R1203 B.n197 B.n196 163.367
R1204 B.n198 B.n197 163.367
R1205 B.n198 B.n135 163.367
R1206 B.n202 B.n135 163.367
R1207 B.n203 B.n202 163.367
R1208 B.n204 B.n203 163.367
R1209 B.n204 B.n133 163.367
R1210 B.n208 B.n133 163.367
R1211 B.n209 B.n208 163.367
R1212 B.n210 B.n209 163.367
R1213 B.n210 B.n131 163.367
R1214 B.n214 B.n131 163.367
R1215 B.n215 B.n214 163.367
R1216 B.n216 B.n215 163.367
R1217 B.n216 B.n129 163.367
R1218 B.n220 B.n129 163.367
R1219 B.n221 B.n220 163.367
R1220 B.n222 B.n221 163.367
R1221 B.n222 B.n127 163.367
R1222 B.n226 B.n127 163.367
R1223 B.n227 B.n226 163.367
R1224 B.n228 B.n227 163.367
R1225 B.n228 B.n125 163.367
R1226 B.n232 B.n125 163.367
R1227 B.n233 B.n232 163.367
R1228 B.n234 B.n233 163.367
R1229 B.n234 B.n123 163.367
R1230 B.n238 B.n123 163.367
R1231 B.n239 B.n238 163.367
R1232 B.n240 B.n239 163.367
R1233 B.n240 B.n121 163.367
R1234 B.n244 B.n121 163.367
R1235 B.n245 B.n244 163.367
R1236 B.n246 B.n245 163.367
R1237 B.n246 B.n117 163.367
R1238 B.n251 B.n117 163.367
R1239 B.n252 B.n251 163.367
R1240 B.n253 B.n252 163.367
R1241 B.n253 B.n115 163.367
R1242 B.n257 B.n115 163.367
R1243 B.n258 B.n257 163.367
R1244 B.n259 B.n258 163.367
R1245 B.n259 B.n113 163.367
R1246 B.n263 B.n113 163.367
R1247 B.n264 B.n263 163.367
R1248 B.n264 B.n109 163.367
R1249 B.n268 B.n109 163.367
R1250 B.n269 B.n268 163.367
R1251 B.n270 B.n269 163.367
R1252 B.n270 B.n107 163.367
R1253 B.n274 B.n107 163.367
R1254 B.n275 B.n274 163.367
R1255 B.n276 B.n275 163.367
R1256 B.n276 B.n105 163.367
R1257 B.n280 B.n105 163.367
R1258 B.n281 B.n280 163.367
R1259 B.n282 B.n281 163.367
R1260 B.n282 B.n103 163.367
R1261 B.n286 B.n103 163.367
R1262 B.n287 B.n286 163.367
R1263 B.n288 B.n287 163.367
R1264 B.n288 B.n101 163.367
R1265 B.n292 B.n101 163.367
R1266 B.n293 B.n292 163.367
R1267 B.n294 B.n293 163.367
R1268 B.n294 B.n99 163.367
R1269 B.n298 B.n99 163.367
R1270 B.n299 B.n298 163.367
R1271 B.n300 B.n299 163.367
R1272 B.n300 B.n97 163.367
R1273 B.n304 B.n97 163.367
R1274 B.n305 B.n304 163.367
R1275 B.n306 B.n305 163.367
R1276 B.n306 B.n95 163.367
R1277 B.n310 B.n95 163.367
R1278 B.n311 B.n310 163.367
R1279 B.n312 B.n311 163.367
R1280 B.n312 B.n93 163.367
R1281 B.n316 B.n93 163.367
R1282 B.n317 B.n316 163.367
R1283 B.n318 B.n317 163.367
R1284 B.n318 B.n91 163.367
R1285 B.n322 B.n91 163.367
R1286 B.n323 B.n322 163.367
R1287 B.n324 B.n323 163.367
R1288 B.n324 B.n89 163.367
R1289 B.n328 B.n89 163.367
R1290 B.n329 B.n328 163.367
R1291 B.n330 B.n87 163.367
R1292 B.n334 B.n87 163.367
R1293 B.n335 B.n334 163.367
R1294 B.n336 B.n335 163.367
R1295 B.n336 B.n85 163.367
R1296 B.n340 B.n85 163.367
R1297 B.n341 B.n340 163.367
R1298 B.n342 B.n341 163.367
R1299 B.n342 B.n83 163.367
R1300 B.n346 B.n83 163.367
R1301 B.n347 B.n346 163.367
R1302 B.n348 B.n347 163.367
R1303 B.n348 B.n81 163.367
R1304 B.n352 B.n81 163.367
R1305 B.n353 B.n352 163.367
R1306 B.n354 B.n353 163.367
R1307 B.n354 B.n79 163.367
R1308 B.n358 B.n79 163.367
R1309 B.n359 B.n358 163.367
R1310 B.n360 B.n359 163.367
R1311 B.n360 B.n77 163.367
R1312 B.n364 B.n77 163.367
R1313 B.n365 B.n364 163.367
R1314 B.n366 B.n365 163.367
R1315 B.n366 B.n75 163.367
R1316 B.n370 B.n75 163.367
R1317 B.n371 B.n370 163.367
R1318 B.n372 B.n371 163.367
R1319 B.n372 B.n73 163.367
R1320 B.n376 B.n73 163.367
R1321 B.n377 B.n376 163.367
R1322 B.n378 B.n377 163.367
R1323 B.n378 B.n71 163.367
R1324 B.n382 B.n71 163.367
R1325 B.n383 B.n382 163.367
R1326 B.n384 B.n383 163.367
R1327 B.n384 B.n69 163.367
R1328 B.n388 B.n69 163.367
R1329 B.n389 B.n388 163.367
R1330 B.n390 B.n389 163.367
R1331 B.n390 B.n67 163.367
R1332 B.n394 B.n67 163.367
R1333 B.n395 B.n394 163.367
R1334 B.n396 B.n395 163.367
R1335 B.n542 B.n13 163.367
R1336 B.n542 B.n541 163.367
R1337 B.n541 B.n540 163.367
R1338 B.n540 B.n15 163.367
R1339 B.n536 B.n15 163.367
R1340 B.n536 B.n535 163.367
R1341 B.n535 B.n534 163.367
R1342 B.n534 B.n17 163.367
R1343 B.n530 B.n17 163.367
R1344 B.n530 B.n529 163.367
R1345 B.n529 B.n528 163.367
R1346 B.n528 B.n19 163.367
R1347 B.n524 B.n19 163.367
R1348 B.n524 B.n523 163.367
R1349 B.n523 B.n522 163.367
R1350 B.n522 B.n21 163.367
R1351 B.n518 B.n21 163.367
R1352 B.n518 B.n517 163.367
R1353 B.n517 B.n516 163.367
R1354 B.n516 B.n23 163.367
R1355 B.n512 B.n23 163.367
R1356 B.n512 B.n511 163.367
R1357 B.n511 B.n510 163.367
R1358 B.n510 B.n25 163.367
R1359 B.n506 B.n25 163.367
R1360 B.n506 B.n505 163.367
R1361 B.n505 B.n504 163.367
R1362 B.n504 B.n27 163.367
R1363 B.n500 B.n27 163.367
R1364 B.n500 B.n499 163.367
R1365 B.n499 B.n498 163.367
R1366 B.n498 B.n29 163.367
R1367 B.n494 B.n29 163.367
R1368 B.n494 B.n493 163.367
R1369 B.n493 B.n492 163.367
R1370 B.n492 B.n31 163.367
R1371 B.n488 B.n31 163.367
R1372 B.n488 B.n487 163.367
R1373 B.n487 B.n486 163.367
R1374 B.n486 B.n33 163.367
R1375 B.n482 B.n33 163.367
R1376 B.n482 B.n481 163.367
R1377 B.n481 B.n480 163.367
R1378 B.n480 B.n35 163.367
R1379 B.n475 B.n35 163.367
R1380 B.n475 B.n474 163.367
R1381 B.n474 B.n473 163.367
R1382 B.n473 B.n39 163.367
R1383 B.n469 B.n39 163.367
R1384 B.n469 B.n468 163.367
R1385 B.n468 B.n467 163.367
R1386 B.n467 B.n41 163.367
R1387 B.n462 B.n41 163.367
R1388 B.n462 B.n461 163.367
R1389 B.n461 B.n460 163.367
R1390 B.n460 B.n45 163.367
R1391 B.n456 B.n45 163.367
R1392 B.n456 B.n455 163.367
R1393 B.n455 B.n454 163.367
R1394 B.n454 B.n47 163.367
R1395 B.n450 B.n47 163.367
R1396 B.n450 B.n449 163.367
R1397 B.n449 B.n448 163.367
R1398 B.n448 B.n49 163.367
R1399 B.n444 B.n49 163.367
R1400 B.n444 B.n443 163.367
R1401 B.n443 B.n442 163.367
R1402 B.n442 B.n51 163.367
R1403 B.n438 B.n51 163.367
R1404 B.n438 B.n437 163.367
R1405 B.n437 B.n436 163.367
R1406 B.n436 B.n53 163.367
R1407 B.n432 B.n53 163.367
R1408 B.n432 B.n431 163.367
R1409 B.n431 B.n430 163.367
R1410 B.n430 B.n55 163.367
R1411 B.n426 B.n55 163.367
R1412 B.n426 B.n425 163.367
R1413 B.n425 B.n424 163.367
R1414 B.n424 B.n57 163.367
R1415 B.n420 B.n57 163.367
R1416 B.n420 B.n419 163.367
R1417 B.n419 B.n418 163.367
R1418 B.n418 B.n59 163.367
R1419 B.n414 B.n59 163.367
R1420 B.n414 B.n413 163.367
R1421 B.n413 B.n412 163.367
R1422 B.n412 B.n61 163.367
R1423 B.n408 B.n61 163.367
R1424 B.n408 B.n407 163.367
R1425 B.n407 B.n406 163.367
R1426 B.n406 B.n63 163.367
R1427 B.n402 B.n63 163.367
R1428 B.n402 B.n401 163.367
R1429 B.n401 B.n400 163.367
R1430 B.n400 B.n65 163.367
R1431 B.n112 B.n111 59.5399
R1432 B.n249 B.n119 59.5399
R1433 B.n478 B.n37 59.5399
R1434 B.n464 B.n43 59.5399
R1435 B.n111 B.n110 45.7702
R1436 B.n119 B.n118 45.7702
R1437 B.n37 B.n36 45.7702
R1438 B.n43 B.n42 45.7702
R1439 B.n545 B.n544 30.7517
R1440 B.n398 B.n397 30.7517
R1441 B.n331 B.n88 30.7517
R1442 B.n183 B.n182 30.7517
R1443 B B.n579 18.0485
R1444 B.n544 B.n543 10.6151
R1445 B.n543 B.n14 10.6151
R1446 B.n539 B.n14 10.6151
R1447 B.n539 B.n538 10.6151
R1448 B.n538 B.n537 10.6151
R1449 B.n537 B.n16 10.6151
R1450 B.n533 B.n16 10.6151
R1451 B.n533 B.n532 10.6151
R1452 B.n532 B.n531 10.6151
R1453 B.n531 B.n18 10.6151
R1454 B.n527 B.n18 10.6151
R1455 B.n527 B.n526 10.6151
R1456 B.n526 B.n525 10.6151
R1457 B.n525 B.n20 10.6151
R1458 B.n521 B.n20 10.6151
R1459 B.n521 B.n520 10.6151
R1460 B.n520 B.n519 10.6151
R1461 B.n519 B.n22 10.6151
R1462 B.n515 B.n22 10.6151
R1463 B.n515 B.n514 10.6151
R1464 B.n514 B.n513 10.6151
R1465 B.n513 B.n24 10.6151
R1466 B.n509 B.n24 10.6151
R1467 B.n509 B.n508 10.6151
R1468 B.n508 B.n507 10.6151
R1469 B.n507 B.n26 10.6151
R1470 B.n503 B.n26 10.6151
R1471 B.n503 B.n502 10.6151
R1472 B.n502 B.n501 10.6151
R1473 B.n501 B.n28 10.6151
R1474 B.n497 B.n28 10.6151
R1475 B.n497 B.n496 10.6151
R1476 B.n496 B.n495 10.6151
R1477 B.n495 B.n30 10.6151
R1478 B.n491 B.n30 10.6151
R1479 B.n491 B.n490 10.6151
R1480 B.n490 B.n489 10.6151
R1481 B.n489 B.n32 10.6151
R1482 B.n485 B.n32 10.6151
R1483 B.n485 B.n484 10.6151
R1484 B.n484 B.n483 10.6151
R1485 B.n483 B.n34 10.6151
R1486 B.n479 B.n34 10.6151
R1487 B.n477 B.n476 10.6151
R1488 B.n476 B.n38 10.6151
R1489 B.n472 B.n38 10.6151
R1490 B.n472 B.n471 10.6151
R1491 B.n471 B.n470 10.6151
R1492 B.n470 B.n40 10.6151
R1493 B.n466 B.n40 10.6151
R1494 B.n466 B.n465 10.6151
R1495 B.n463 B.n44 10.6151
R1496 B.n459 B.n44 10.6151
R1497 B.n459 B.n458 10.6151
R1498 B.n458 B.n457 10.6151
R1499 B.n457 B.n46 10.6151
R1500 B.n453 B.n46 10.6151
R1501 B.n453 B.n452 10.6151
R1502 B.n452 B.n451 10.6151
R1503 B.n451 B.n48 10.6151
R1504 B.n447 B.n48 10.6151
R1505 B.n447 B.n446 10.6151
R1506 B.n446 B.n445 10.6151
R1507 B.n445 B.n50 10.6151
R1508 B.n441 B.n50 10.6151
R1509 B.n441 B.n440 10.6151
R1510 B.n440 B.n439 10.6151
R1511 B.n439 B.n52 10.6151
R1512 B.n435 B.n52 10.6151
R1513 B.n435 B.n434 10.6151
R1514 B.n434 B.n433 10.6151
R1515 B.n433 B.n54 10.6151
R1516 B.n429 B.n54 10.6151
R1517 B.n429 B.n428 10.6151
R1518 B.n428 B.n427 10.6151
R1519 B.n427 B.n56 10.6151
R1520 B.n423 B.n56 10.6151
R1521 B.n423 B.n422 10.6151
R1522 B.n422 B.n421 10.6151
R1523 B.n421 B.n58 10.6151
R1524 B.n417 B.n58 10.6151
R1525 B.n417 B.n416 10.6151
R1526 B.n416 B.n415 10.6151
R1527 B.n415 B.n60 10.6151
R1528 B.n411 B.n60 10.6151
R1529 B.n411 B.n410 10.6151
R1530 B.n410 B.n409 10.6151
R1531 B.n409 B.n62 10.6151
R1532 B.n405 B.n62 10.6151
R1533 B.n405 B.n404 10.6151
R1534 B.n404 B.n403 10.6151
R1535 B.n403 B.n64 10.6151
R1536 B.n399 B.n64 10.6151
R1537 B.n399 B.n398 10.6151
R1538 B.n332 B.n331 10.6151
R1539 B.n333 B.n332 10.6151
R1540 B.n333 B.n86 10.6151
R1541 B.n337 B.n86 10.6151
R1542 B.n338 B.n337 10.6151
R1543 B.n339 B.n338 10.6151
R1544 B.n339 B.n84 10.6151
R1545 B.n343 B.n84 10.6151
R1546 B.n344 B.n343 10.6151
R1547 B.n345 B.n344 10.6151
R1548 B.n345 B.n82 10.6151
R1549 B.n349 B.n82 10.6151
R1550 B.n350 B.n349 10.6151
R1551 B.n351 B.n350 10.6151
R1552 B.n351 B.n80 10.6151
R1553 B.n355 B.n80 10.6151
R1554 B.n356 B.n355 10.6151
R1555 B.n357 B.n356 10.6151
R1556 B.n357 B.n78 10.6151
R1557 B.n361 B.n78 10.6151
R1558 B.n362 B.n361 10.6151
R1559 B.n363 B.n362 10.6151
R1560 B.n363 B.n76 10.6151
R1561 B.n367 B.n76 10.6151
R1562 B.n368 B.n367 10.6151
R1563 B.n369 B.n368 10.6151
R1564 B.n369 B.n74 10.6151
R1565 B.n373 B.n74 10.6151
R1566 B.n374 B.n373 10.6151
R1567 B.n375 B.n374 10.6151
R1568 B.n375 B.n72 10.6151
R1569 B.n379 B.n72 10.6151
R1570 B.n380 B.n379 10.6151
R1571 B.n381 B.n380 10.6151
R1572 B.n381 B.n70 10.6151
R1573 B.n385 B.n70 10.6151
R1574 B.n386 B.n385 10.6151
R1575 B.n387 B.n386 10.6151
R1576 B.n387 B.n68 10.6151
R1577 B.n391 B.n68 10.6151
R1578 B.n392 B.n391 10.6151
R1579 B.n393 B.n392 10.6151
R1580 B.n393 B.n66 10.6151
R1581 B.n397 B.n66 10.6151
R1582 B.n183 B.n140 10.6151
R1583 B.n187 B.n140 10.6151
R1584 B.n188 B.n187 10.6151
R1585 B.n189 B.n188 10.6151
R1586 B.n189 B.n138 10.6151
R1587 B.n193 B.n138 10.6151
R1588 B.n194 B.n193 10.6151
R1589 B.n195 B.n194 10.6151
R1590 B.n195 B.n136 10.6151
R1591 B.n199 B.n136 10.6151
R1592 B.n200 B.n199 10.6151
R1593 B.n201 B.n200 10.6151
R1594 B.n201 B.n134 10.6151
R1595 B.n205 B.n134 10.6151
R1596 B.n206 B.n205 10.6151
R1597 B.n207 B.n206 10.6151
R1598 B.n207 B.n132 10.6151
R1599 B.n211 B.n132 10.6151
R1600 B.n212 B.n211 10.6151
R1601 B.n213 B.n212 10.6151
R1602 B.n213 B.n130 10.6151
R1603 B.n217 B.n130 10.6151
R1604 B.n218 B.n217 10.6151
R1605 B.n219 B.n218 10.6151
R1606 B.n219 B.n128 10.6151
R1607 B.n223 B.n128 10.6151
R1608 B.n224 B.n223 10.6151
R1609 B.n225 B.n224 10.6151
R1610 B.n225 B.n126 10.6151
R1611 B.n229 B.n126 10.6151
R1612 B.n230 B.n229 10.6151
R1613 B.n231 B.n230 10.6151
R1614 B.n231 B.n124 10.6151
R1615 B.n235 B.n124 10.6151
R1616 B.n236 B.n235 10.6151
R1617 B.n237 B.n236 10.6151
R1618 B.n237 B.n122 10.6151
R1619 B.n241 B.n122 10.6151
R1620 B.n242 B.n241 10.6151
R1621 B.n243 B.n242 10.6151
R1622 B.n243 B.n120 10.6151
R1623 B.n247 B.n120 10.6151
R1624 B.n248 B.n247 10.6151
R1625 B.n250 B.n116 10.6151
R1626 B.n254 B.n116 10.6151
R1627 B.n255 B.n254 10.6151
R1628 B.n256 B.n255 10.6151
R1629 B.n256 B.n114 10.6151
R1630 B.n260 B.n114 10.6151
R1631 B.n261 B.n260 10.6151
R1632 B.n262 B.n261 10.6151
R1633 B.n266 B.n265 10.6151
R1634 B.n267 B.n266 10.6151
R1635 B.n267 B.n108 10.6151
R1636 B.n271 B.n108 10.6151
R1637 B.n272 B.n271 10.6151
R1638 B.n273 B.n272 10.6151
R1639 B.n273 B.n106 10.6151
R1640 B.n277 B.n106 10.6151
R1641 B.n278 B.n277 10.6151
R1642 B.n279 B.n278 10.6151
R1643 B.n279 B.n104 10.6151
R1644 B.n283 B.n104 10.6151
R1645 B.n284 B.n283 10.6151
R1646 B.n285 B.n284 10.6151
R1647 B.n285 B.n102 10.6151
R1648 B.n289 B.n102 10.6151
R1649 B.n290 B.n289 10.6151
R1650 B.n291 B.n290 10.6151
R1651 B.n291 B.n100 10.6151
R1652 B.n295 B.n100 10.6151
R1653 B.n296 B.n295 10.6151
R1654 B.n297 B.n296 10.6151
R1655 B.n297 B.n98 10.6151
R1656 B.n301 B.n98 10.6151
R1657 B.n302 B.n301 10.6151
R1658 B.n303 B.n302 10.6151
R1659 B.n303 B.n96 10.6151
R1660 B.n307 B.n96 10.6151
R1661 B.n308 B.n307 10.6151
R1662 B.n309 B.n308 10.6151
R1663 B.n309 B.n94 10.6151
R1664 B.n313 B.n94 10.6151
R1665 B.n314 B.n313 10.6151
R1666 B.n315 B.n314 10.6151
R1667 B.n315 B.n92 10.6151
R1668 B.n319 B.n92 10.6151
R1669 B.n320 B.n319 10.6151
R1670 B.n321 B.n320 10.6151
R1671 B.n321 B.n90 10.6151
R1672 B.n325 B.n90 10.6151
R1673 B.n326 B.n325 10.6151
R1674 B.n327 B.n326 10.6151
R1675 B.n327 B.n88 10.6151
R1676 B.n182 B.n181 10.6151
R1677 B.n181 B.n142 10.6151
R1678 B.n177 B.n142 10.6151
R1679 B.n177 B.n176 10.6151
R1680 B.n176 B.n175 10.6151
R1681 B.n175 B.n144 10.6151
R1682 B.n171 B.n144 10.6151
R1683 B.n171 B.n170 10.6151
R1684 B.n170 B.n169 10.6151
R1685 B.n169 B.n146 10.6151
R1686 B.n165 B.n146 10.6151
R1687 B.n165 B.n164 10.6151
R1688 B.n164 B.n163 10.6151
R1689 B.n163 B.n148 10.6151
R1690 B.n159 B.n148 10.6151
R1691 B.n159 B.n158 10.6151
R1692 B.n158 B.n157 10.6151
R1693 B.n157 B.n150 10.6151
R1694 B.n153 B.n150 10.6151
R1695 B.n153 B.n152 10.6151
R1696 B.n152 B.n0 10.6151
R1697 B.n575 B.n1 10.6151
R1698 B.n575 B.n574 10.6151
R1699 B.n574 B.n573 10.6151
R1700 B.n573 B.n4 10.6151
R1701 B.n569 B.n4 10.6151
R1702 B.n569 B.n568 10.6151
R1703 B.n568 B.n567 10.6151
R1704 B.n567 B.n6 10.6151
R1705 B.n563 B.n6 10.6151
R1706 B.n563 B.n562 10.6151
R1707 B.n562 B.n561 10.6151
R1708 B.n561 B.n8 10.6151
R1709 B.n557 B.n8 10.6151
R1710 B.n557 B.n556 10.6151
R1711 B.n556 B.n555 10.6151
R1712 B.n555 B.n10 10.6151
R1713 B.n551 B.n10 10.6151
R1714 B.n551 B.n550 10.6151
R1715 B.n550 B.n549 10.6151
R1716 B.n549 B.n12 10.6151
R1717 B.n545 B.n12 10.6151
R1718 B.n478 B.n477 6.5566
R1719 B.n465 B.n464 6.5566
R1720 B.n250 B.n249 6.5566
R1721 B.n262 B.n112 6.5566
R1722 B.n479 B.n478 4.05904
R1723 B.n464 B.n463 4.05904
R1724 B.n249 B.n248 4.05904
R1725 B.n265 B.n112 4.05904
R1726 B.n579 B.n0 2.81026
R1727 B.n579 B.n1 2.81026
C0 VN w_n1914_n3500# 2.59909f
C1 VDD1 w_n1914_n3500# 1.76393f
C2 VN VTAIL 2.38923f
C3 VDD1 VTAIL 5.20227f
C4 VN B 0.964661f
C5 VN VP 5.30496f
C6 VDD1 B 1.67845f
C7 w_n1914_n3500# VDD2 1.78299f
C8 VDD1 VP 2.95627f
C9 VDD2 VTAIL 5.24814f
C10 VDD2 B 1.70349f
C11 VP VDD2 0.309561f
C12 w_n1914_n3500# VTAIL 2.87122f
C13 w_n1914_n3500# B 8.37875f
C14 VP w_n1914_n3500# 2.84167f
C15 B VTAIL 3.55544f
C16 VP VTAIL 2.40359f
C17 VP B 1.36118f
C18 VDD1 VN 0.148194f
C19 VN VDD2 2.79792f
C20 VDD1 VDD2 0.60695f
C21 VDD2 VSUBS 0.862594f
C22 VDD1 VSUBS 3.607516f
C23 VTAIL VSUBS 0.960722f
C24 VN VSUBS 7.83285f
C25 VP VSUBS 1.54024f
C26 B VSUBS 3.524449f
C27 w_n1914_n3500# VSUBS 82.38621f
C28 B.n0 VSUBS 0.004001f
C29 B.n1 VSUBS 0.004001f
C30 B.n2 VSUBS 0.006327f
C31 B.n3 VSUBS 0.006327f
C32 B.n4 VSUBS 0.006327f
C33 B.n5 VSUBS 0.006327f
C34 B.n6 VSUBS 0.006327f
C35 B.n7 VSUBS 0.006327f
C36 B.n8 VSUBS 0.006327f
C37 B.n9 VSUBS 0.006327f
C38 B.n10 VSUBS 0.006327f
C39 B.n11 VSUBS 0.006327f
C40 B.n12 VSUBS 0.006327f
C41 B.n13 VSUBS 0.01471f
C42 B.n14 VSUBS 0.006327f
C43 B.n15 VSUBS 0.006327f
C44 B.n16 VSUBS 0.006327f
C45 B.n17 VSUBS 0.006327f
C46 B.n18 VSUBS 0.006327f
C47 B.n19 VSUBS 0.006327f
C48 B.n20 VSUBS 0.006327f
C49 B.n21 VSUBS 0.006327f
C50 B.n22 VSUBS 0.006327f
C51 B.n23 VSUBS 0.006327f
C52 B.n24 VSUBS 0.006327f
C53 B.n25 VSUBS 0.006327f
C54 B.n26 VSUBS 0.006327f
C55 B.n27 VSUBS 0.006327f
C56 B.n28 VSUBS 0.006327f
C57 B.n29 VSUBS 0.006327f
C58 B.n30 VSUBS 0.006327f
C59 B.n31 VSUBS 0.006327f
C60 B.n32 VSUBS 0.006327f
C61 B.n33 VSUBS 0.006327f
C62 B.n34 VSUBS 0.006327f
C63 B.n35 VSUBS 0.006327f
C64 B.t11 VSUBS 0.203965f
C65 B.t10 VSUBS 0.227719f
C66 B.t9 VSUBS 1.03595f
C67 B.n36 VSUBS 0.354154f
C68 B.n37 VSUBS 0.233823f
C69 B.n38 VSUBS 0.006327f
C70 B.n39 VSUBS 0.006327f
C71 B.n40 VSUBS 0.006327f
C72 B.n41 VSUBS 0.006327f
C73 B.t2 VSUBS 0.203968f
C74 B.t1 VSUBS 0.227721f
C75 B.t0 VSUBS 1.03595f
C76 B.n42 VSUBS 0.354151f
C77 B.n43 VSUBS 0.23382f
C78 B.n44 VSUBS 0.006327f
C79 B.n45 VSUBS 0.006327f
C80 B.n46 VSUBS 0.006327f
C81 B.n47 VSUBS 0.006327f
C82 B.n48 VSUBS 0.006327f
C83 B.n49 VSUBS 0.006327f
C84 B.n50 VSUBS 0.006327f
C85 B.n51 VSUBS 0.006327f
C86 B.n52 VSUBS 0.006327f
C87 B.n53 VSUBS 0.006327f
C88 B.n54 VSUBS 0.006327f
C89 B.n55 VSUBS 0.006327f
C90 B.n56 VSUBS 0.006327f
C91 B.n57 VSUBS 0.006327f
C92 B.n58 VSUBS 0.006327f
C93 B.n59 VSUBS 0.006327f
C94 B.n60 VSUBS 0.006327f
C95 B.n61 VSUBS 0.006327f
C96 B.n62 VSUBS 0.006327f
C97 B.n63 VSUBS 0.006327f
C98 B.n64 VSUBS 0.006327f
C99 B.n65 VSUBS 0.01471f
C100 B.n66 VSUBS 0.006327f
C101 B.n67 VSUBS 0.006327f
C102 B.n68 VSUBS 0.006327f
C103 B.n69 VSUBS 0.006327f
C104 B.n70 VSUBS 0.006327f
C105 B.n71 VSUBS 0.006327f
C106 B.n72 VSUBS 0.006327f
C107 B.n73 VSUBS 0.006327f
C108 B.n74 VSUBS 0.006327f
C109 B.n75 VSUBS 0.006327f
C110 B.n76 VSUBS 0.006327f
C111 B.n77 VSUBS 0.006327f
C112 B.n78 VSUBS 0.006327f
C113 B.n79 VSUBS 0.006327f
C114 B.n80 VSUBS 0.006327f
C115 B.n81 VSUBS 0.006327f
C116 B.n82 VSUBS 0.006327f
C117 B.n83 VSUBS 0.006327f
C118 B.n84 VSUBS 0.006327f
C119 B.n85 VSUBS 0.006327f
C120 B.n86 VSUBS 0.006327f
C121 B.n87 VSUBS 0.006327f
C122 B.n88 VSUBS 0.01471f
C123 B.n89 VSUBS 0.006327f
C124 B.n90 VSUBS 0.006327f
C125 B.n91 VSUBS 0.006327f
C126 B.n92 VSUBS 0.006327f
C127 B.n93 VSUBS 0.006327f
C128 B.n94 VSUBS 0.006327f
C129 B.n95 VSUBS 0.006327f
C130 B.n96 VSUBS 0.006327f
C131 B.n97 VSUBS 0.006327f
C132 B.n98 VSUBS 0.006327f
C133 B.n99 VSUBS 0.006327f
C134 B.n100 VSUBS 0.006327f
C135 B.n101 VSUBS 0.006327f
C136 B.n102 VSUBS 0.006327f
C137 B.n103 VSUBS 0.006327f
C138 B.n104 VSUBS 0.006327f
C139 B.n105 VSUBS 0.006327f
C140 B.n106 VSUBS 0.006327f
C141 B.n107 VSUBS 0.006327f
C142 B.n108 VSUBS 0.006327f
C143 B.n109 VSUBS 0.006327f
C144 B.t7 VSUBS 0.203968f
C145 B.t8 VSUBS 0.227721f
C146 B.t6 VSUBS 1.03595f
C147 B.n110 VSUBS 0.354151f
C148 B.n111 VSUBS 0.23382f
C149 B.n112 VSUBS 0.014659f
C150 B.n113 VSUBS 0.006327f
C151 B.n114 VSUBS 0.006327f
C152 B.n115 VSUBS 0.006327f
C153 B.n116 VSUBS 0.006327f
C154 B.n117 VSUBS 0.006327f
C155 B.t4 VSUBS 0.203965f
C156 B.t5 VSUBS 0.227719f
C157 B.t3 VSUBS 1.03595f
C158 B.n118 VSUBS 0.354154f
C159 B.n119 VSUBS 0.233823f
C160 B.n120 VSUBS 0.006327f
C161 B.n121 VSUBS 0.006327f
C162 B.n122 VSUBS 0.006327f
C163 B.n123 VSUBS 0.006327f
C164 B.n124 VSUBS 0.006327f
C165 B.n125 VSUBS 0.006327f
C166 B.n126 VSUBS 0.006327f
C167 B.n127 VSUBS 0.006327f
C168 B.n128 VSUBS 0.006327f
C169 B.n129 VSUBS 0.006327f
C170 B.n130 VSUBS 0.006327f
C171 B.n131 VSUBS 0.006327f
C172 B.n132 VSUBS 0.006327f
C173 B.n133 VSUBS 0.006327f
C174 B.n134 VSUBS 0.006327f
C175 B.n135 VSUBS 0.006327f
C176 B.n136 VSUBS 0.006327f
C177 B.n137 VSUBS 0.006327f
C178 B.n138 VSUBS 0.006327f
C179 B.n139 VSUBS 0.006327f
C180 B.n140 VSUBS 0.006327f
C181 B.n141 VSUBS 0.013761f
C182 B.n142 VSUBS 0.006327f
C183 B.n143 VSUBS 0.006327f
C184 B.n144 VSUBS 0.006327f
C185 B.n145 VSUBS 0.006327f
C186 B.n146 VSUBS 0.006327f
C187 B.n147 VSUBS 0.006327f
C188 B.n148 VSUBS 0.006327f
C189 B.n149 VSUBS 0.006327f
C190 B.n150 VSUBS 0.006327f
C191 B.n151 VSUBS 0.006327f
C192 B.n152 VSUBS 0.006327f
C193 B.n153 VSUBS 0.006327f
C194 B.n154 VSUBS 0.006327f
C195 B.n155 VSUBS 0.006327f
C196 B.n156 VSUBS 0.006327f
C197 B.n157 VSUBS 0.006327f
C198 B.n158 VSUBS 0.006327f
C199 B.n159 VSUBS 0.006327f
C200 B.n160 VSUBS 0.006327f
C201 B.n161 VSUBS 0.006327f
C202 B.n162 VSUBS 0.006327f
C203 B.n163 VSUBS 0.006327f
C204 B.n164 VSUBS 0.006327f
C205 B.n165 VSUBS 0.006327f
C206 B.n166 VSUBS 0.006327f
C207 B.n167 VSUBS 0.006327f
C208 B.n168 VSUBS 0.006327f
C209 B.n169 VSUBS 0.006327f
C210 B.n170 VSUBS 0.006327f
C211 B.n171 VSUBS 0.006327f
C212 B.n172 VSUBS 0.006327f
C213 B.n173 VSUBS 0.006327f
C214 B.n174 VSUBS 0.006327f
C215 B.n175 VSUBS 0.006327f
C216 B.n176 VSUBS 0.006327f
C217 B.n177 VSUBS 0.006327f
C218 B.n178 VSUBS 0.006327f
C219 B.n179 VSUBS 0.006327f
C220 B.n180 VSUBS 0.006327f
C221 B.n181 VSUBS 0.006327f
C222 B.n182 VSUBS 0.013761f
C223 B.n183 VSUBS 0.01471f
C224 B.n184 VSUBS 0.01471f
C225 B.n185 VSUBS 0.006327f
C226 B.n186 VSUBS 0.006327f
C227 B.n187 VSUBS 0.006327f
C228 B.n188 VSUBS 0.006327f
C229 B.n189 VSUBS 0.006327f
C230 B.n190 VSUBS 0.006327f
C231 B.n191 VSUBS 0.006327f
C232 B.n192 VSUBS 0.006327f
C233 B.n193 VSUBS 0.006327f
C234 B.n194 VSUBS 0.006327f
C235 B.n195 VSUBS 0.006327f
C236 B.n196 VSUBS 0.006327f
C237 B.n197 VSUBS 0.006327f
C238 B.n198 VSUBS 0.006327f
C239 B.n199 VSUBS 0.006327f
C240 B.n200 VSUBS 0.006327f
C241 B.n201 VSUBS 0.006327f
C242 B.n202 VSUBS 0.006327f
C243 B.n203 VSUBS 0.006327f
C244 B.n204 VSUBS 0.006327f
C245 B.n205 VSUBS 0.006327f
C246 B.n206 VSUBS 0.006327f
C247 B.n207 VSUBS 0.006327f
C248 B.n208 VSUBS 0.006327f
C249 B.n209 VSUBS 0.006327f
C250 B.n210 VSUBS 0.006327f
C251 B.n211 VSUBS 0.006327f
C252 B.n212 VSUBS 0.006327f
C253 B.n213 VSUBS 0.006327f
C254 B.n214 VSUBS 0.006327f
C255 B.n215 VSUBS 0.006327f
C256 B.n216 VSUBS 0.006327f
C257 B.n217 VSUBS 0.006327f
C258 B.n218 VSUBS 0.006327f
C259 B.n219 VSUBS 0.006327f
C260 B.n220 VSUBS 0.006327f
C261 B.n221 VSUBS 0.006327f
C262 B.n222 VSUBS 0.006327f
C263 B.n223 VSUBS 0.006327f
C264 B.n224 VSUBS 0.006327f
C265 B.n225 VSUBS 0.006327f
C266 B.n226 VSUBS 0.006327f
C267 B.n227 VSUBS 0.006327f
C268 B.n228 VSUBS 0.006327f
C269 B.n229 VSUBS 0.006327f
C270 B.n230 VSUBS 0.006327f
C271 B.n231 VSUBS 0.006327f
C272 B.n232 VSUBS 0.006327f
C273 B.n233 VSUBS 0.006327f
C274 B.n234 VSUBS 0.006327f
C275 B.n235 VSUBS 0.006327f
C276 B.n236 VSUBS 0.006327f
C277 B.n237 VSUBS 0.006327f
C278 B.n238 VSUBS 0.006327f
C279 B.n239 VSUBS 0.006327f
C280 B.n240 VSUBS 0.006327f
C281 B.n241 VSUBS 0.006327f
C282 B.n242 VSUBS 0.006327f
C283 B.n243 VSUBS 0.006327f
C284 B.n244 VSUBS 0.006327f
C285 B.n245 VSUBS 0.006327f
C286 B.n246 VSUBS 0.006327f
C287 B.n247 VSUBS 0.006327f
C288 B.n248 VSUBS 0.004373f
C289 B.n249 VSUBS 0.014659f
C290 B.n250 VSUBS 0.005117f
C291 B.n251 VSUBS 0.006327f
C292 B.n252 VSUBS 0.006327f
C293 B.n253 VSUBS 0.006327f
C294 B.n254 VSUBS 0.006327f
C295 B.n255 VSUBS 0.006327f
C296 B.n256 VSUBS 0.006327f
C297 B.n257 VSUBS 0.006327f
C298 B.n258 VSUBS 0.006327f
C299 B.n259 VSUBS 0.006327f
C300 B.n260 VSUBS 0.006327f
C301 B.n261 VSUBS 0.006327f
C302 B.n262 VSUBS 0.005117f
C303 B.n263 VSUBS 0.006327f
C304 B.n264 VSUBS 0.006327f
C305 B.n265 VSUBS 0.004373f
C306 B.n266 VSUBS 0.006327f
C307 B.n267 VSUBS 0.006327f
C308 B.n268 VSUBS 0.006327f
C309 B.n269 VSUBS 0.006327f
C310 B.n270 VSUBS 0.006327f
C311 B.n271 VSUBS 0.006327f
C312 B.n272 VSUBS 0.006327f
C313 B.n273 VSUBS 0.006327f
C314 B.n274 VSUBS 0.006327f
C315 B.n275 VSUBS 0.006327f
C316 B.n276 VSUBS 0.006327f
C317 B.n277 VSUBS 0.006327f
C318 B.n278 VSUBS 0.006327f
C319 B.n279 VSUBS 0.006327f
C320 B.n280 VSUBS 0.006327f
C321 B.n281 VSUBS 0.006327f
C322 B.n282 VSUBS 0.006327f
C323 B.n283 VSUBS 0.006327f
C324 B.n284 VSUBS 0.006327f
C325 B.n285 VSUBS 0.006327f
C326 B.n286 VSUBS 0.006327f
C327 B.n287 VSUBS 0.006327f
C328 B.n288 VSUBS 0.006327f
C329 B.n289 VSUBS 0.006327f
C330 B.n290 VSUBS 0.006327f
C331 B.n291 VSUBS 0.006327f
C332 B.n292 VSUBS 0.006327f
C333 B.n293 VSUBS 0.006327f
C334 B.n294 VSUBS 0.006327f
C335 B.n295 VSUBS 0.006327f
C336 B.n296 VSUBS 0.006327f
C337 B.n297 VSUBS 0.006327f
C338 B.n298 VSUBS 0.006327f
C339 B.n299 VSUBS 0.006327f
C340 B.n300 VSUBS 0.006327f
C341 B.n301 VSUBS 0.006327f
C342 B.n302 VSUBS 0.006327f
C343 B.n303 VSUBS 0.006327f
C344 B.n304 VSUBS 0.006327f
C345 B.n305 VSUBS 0.006327f
C346 B.n306 VSUBS 0.006327f
C347 B.n307 VSUBS 0.006327f
C348 B.n308 VSUBS 0.006327f
C349 B.n309 VSUBS 0.006327f
C350 B.n310 VSUBS 0.006327f
C351 B.n311 VSUBS 0.006327f
C352 B.n312 VSUBS 0.006327f
C353 B.n313 VSUBS 0.006327f
C354 B.n314 VSUBS 0.006327f
C355 B.n315 VSUBS 0.006327f
C356 B.n316 VSUBS 0.006327f
C357 B.n317 VSUBS 0.006327f
C358 B.n318 VSUBS 0.006327f
C359 B.n319 VSUBS 0.006327f
C360 B.n320 VSUBS 0.006327f
C361 B.n321 VSUBS 0.006327f
C362 B.n322 VSUBS 0.006327f
C363 B.n323 VSUBS 0.006327f
C364 B.n324 VSUBS 0.006327f
C365 B.n325 VSUBS 0.006327f
C366 B.n326 VSUBS 0.006327f
C367 B.n327 VSUBS 0.006327f
C368 B.n328 VSUBS 0.006327f
C369 B.n329 VSUBS 0.01471f
C370 B.n330 VSUBS 0.013761f
C371 B.n331 VSUBS 0.013761f
C372 B.n332 VSUBS 0.006327f
C373 B.n333 VSUBS 0.006327f
C374 B.n334 VSUBS 0.006327f
C375 B.n335 VSUBS 0.006327f
C376 B.n336 VSUBS 0.006327f
C377 B.n337 VSUBS 0.006327f
C378 B.n338 VSUBS 0.006327f
C379 B.n339 VSUBS 0.006327f
C380 B.n340 VSUBS 0.006327f
C381 B.n341 VSUBS 0.006327f
C382 B.n342 VSUBS 0.006327f
C383 B.n343 VSUBS 0.006327f
C384 B.n344 VSUBS 0.006327f
C385 B.n345 VSUBS 0.006327f
C386 B.n346 VSUBS 0.006327f
C387 B.n347 VSUBS 0.006327f
C388 B.n348 VSUBS 0.006327f
C389 B.n349 VSUBS 0.006327f
C390 B.n350 VSUBS 0.006327f
C391 B.n351 VSUBS 0.006327f
C392 B.n352 VSUBS 0.006327f
C393 B.n353 VSUBS 0.006327f
C394 B.n354 VSUBS 0.006327f
C395 B.n355 VSUBS 0.006327f
C396 B.n356 VSUBS 0.006327f
C397 B.n357 VSUBS 0.006327f
C398 B.n358 VSUBS 0.006327f
C399 B.n359 VSUBS 0.006327f
C400 B.n360 VSUBS 0.006327f
C401 B.n361 VSUBS 0.006327f
C402 B.n362 VSUBS 0.006327f
C403 B.n363 VSUBS 0.006327f
C404 B.n364 VSUBS 0.006327f
C405 B.n365 VSUBS 0.006327f
C406 B.n366 VSUBS 0.006327f
C407 B.n367 VSUBS 0.006327f
C408 B.n368 VSUBS 0.006327f
C409 B.n369 VSUBS 0.006327f
C410 B.n370 VSUBS 0.006327f
C411 B.n371 VSUBS 0.006327f
C412 B.n372 VSUBS 0.006327f
C413 B.n373 VSUBS 0.006327f
C414 B.n374 VSUBS 0.006327f
C415 B.n375 VSUBS 0.006327f
C416 B.n376 VSUBS 0.006327f
C417 B.n377 VSUBS 0.006327f
C418 B.n378 VSUBS 0.006327f
C419 B.n379 VSUBS 0.006327f
C420 B.n380 VSUBS 0.006327f
C421 B.n381 VSUBS 0.006327f
C422 B.n382 VSUBS 0.006327f
C423 B.n383 VSUBS 0.006327f
C424 B.n384 VSUBS 0.006327f
C425 B.n385 VSUBS 0.006327f
C426 B.n386 VSUBS 0.006327f
C427 B.n387 VSUBS 0.006327f
C428 B.n388 VSUBS 0.006327f
C429 B.n389 VSUBS 0.006327f
C430 B.n390 VSUBS 0.006327f
C431 B.n391 VSUBS 0.006327f
C432 B.n392 VSUBS 0.006327f
C433 B.n393 VSUBS 0.006327f
C434 B.n394 VSUBS 0.006327f
C435 B.n395 VSUBS 0.006327f
C436 B.n396 VSUBS 0.013761f
C437 B.n397 VSUBS 0.014555f
C438 B.n398 VSUBS 0.013916f
C439 B.n399 VSUBS 0.006327f
C440 B.n400 VSUBS 0.006327f
C441 B.n401 VSUBS 0.006327f
C442 B.n402 VSUBS 0.006327f
C443 B.n403 VSUBS 0.006327f
C444 B.n404 VSUBS 0.006327f
C445 B.n405 VSUBS 0.006327f
C446 B.n406 VSUBS 0.006327f
C447 B.n407 VSUBS 0.006327f
C448 B.n408 VSUBS 0.006327f
C449 B.n409 VSUBS 0.006327f
C450 B.n410 VSUBS 0.006327f
C451 B.n411 VSUBS 0.006327f
C452 B.n412 VSUBS 0.006327f
C453 B.n413 VSUBS 0.006327f
C454 B.n414 VSUBS 0.006327f
C455 B.n415 VSUBS 0.006327f
C456 B.n416 VSUBS 0.006327f
C457 B.n417 VSUBS 0.006327f
C458 B.n418 VSUBS 0.006327f
C459 B.n419 VSUBS 0.006327f
C460 B.n420 VSUBS 0.006327f
C461 B.n421 VSUBS 0.006327f
C462 B.n422 VSUBS 0.006327f
C463 B.n423 VSUBS 0.006327f
C464 B.n424 VSUBS 0.006327f
C465 B.n425 VSUBS 0.006327f
C466 B.n426 VSUBS 0.006327f
C467 B.n427 VSUBS 0.006327f
C468 B.n428 VSUBS 0.006327f
C469 B.n429 VSUBS 0.006327f
C470 B.n430 VSUBS 0.006327f
C471 B.n431 VSUBS 0.006327f
C472 B.n432 VSUBS 0.006327f
C473 B.n433 VSUBS 0.006327f
C474 B.n434 VSUBS 0.006327f
C475 B.n435 VSUBS 0.006327f
C476 B.n436 VSUBS 0.006327f
C477 B.n437 VSUBS 0.006327f
C478 B.n438 VSUBS 0.006327f
C479 B.n439 VSUBS 0.006327f
C480 B.n440 VSUBS 0.006327f
C481 B.n441 VSUBS 0.006327f
C482 B.n442 VSUBS 0.006327f
C483 B.n443 VSUBS 0.006327f
C484 B.n444 VSUBS 0.006327f
C485 B.n445 VSUBS 0.006327f
C486 B.n446 VSUBS 0.006327f
C487 B.n447 VSUBS 0.006327f
C488 B.n448 VSUBS 0.006327f
C489 B.n449 VSUBS 0.006327f
C490 B.n450 VSUBS 0.006327f
C491 B.n451 VSUBS 0.006327f
C492 B.n452 VSUBS 0.006327f
C493 B.n453 VSUBS 0.006327f
C494 B.n454 VSUBS 0.006327f
C495 B.n455 VSUBS 0.006327f
C496 B.n456 VSUBS 0.006327f
C497 B.n457 VSUBS 0.006327f
C498 B.n458 VSUBS 0.006327f
C499 B.n459 VSUBS 0.006327f
C500 B.n460 VSUBS 0.006327f
C501 B.n461 VSUBS 0.006327f
C502 B.n462 VSUBS 0.006327f
C503 B.n463 VSUBS 0.004373f
C504 B.n464 VSUBS 0.014659f
C505 B.n465 VSUBS 0.005117f
C506 B.n466 VSUBS 0.006327f
C507 B.n467 VSUBS 0.006327f
C508 B.n468 VSUBS 0.006327f
C509 B.n469 VSUBS 0.006327f
C510 B.n470 VSUBS 0.006327f
C511 B.n471 VSUBS 0.006327f
C512 B.n472 VSUBS 0.006327f
C513 B.n473 VSUBS 0.006327f
C514 B.n474 VSUBS 0.006327f
C515 B.n475 VSUBS 0.006327f
C516 B.n476 VSUBS 0.006327f
C517 B.n477 VSUBS 0.005117f
C518 B.n478 VSUBS 0.014659f
C519 B.n479 VSUBS 0.004373f
C520 B.n480 VSUBS 0.006327f
C521 B.n481 VSUBS 0.006327f
C522 B.n482 VSUBS 0.006327f
C523 B.n483 VSUBS 0.006327f
C524 B.n484 VSUBS 0.006327f
C525 B.n485 VSUBS 0.006327f
C526 B.n486 VSUBS 0.006327f
C527 B.n487 VSUBS 0.006327f
C528 B.n488 VSUBS 0.006327f
C529 B.n489 VSUBS 0.006327f
C530 B.n490 VSUBS 0.006327f
C531 B.n491 VSUBS 0.006327f
C532 B.n492 VSUBS 0.006327f
C533 B.n493 VSUBS 0.006327f
C534 B.n494 VSUBS 0.006327f
C535 B.n495 VSUBS 0.006327f
C536 B.n496 VSUBS 0.006327f
C537 B.n497 VSUBS 0.006327f
C538 B.n498 VSUBS 0.006327f
C539 B.n499 VSUBS 0.006327f
C540 B.n500 VSUBS 0.006327f
C541 B.n501 VSUBS 0.006327f
C542 B.n502 VSUBS 0.006327f
C543 B.n503 VSUBS 0.006327f
C544 B.n504 VSUBS 0.006327f
C545 B.n505 VSUBS 0.006327f
C546 B.n506 VSUBS 0.006327f
C547 B.n507 VSUBS 0.006327f
C548 B.n508 VSUBS 0.006327f
C549 B.n509 VSUBS 0.006327f
C550 B.n510 VSUBS 0.006327f
C551 B.n511 VSUBS 0.006327f
C552 B.n512 VSUBS 0.006327f
C553 B.n513 VSUBS 0.006327f
C554 B.n514 VSUBS 0.006327f
C555 B.n515 VSUBS 0.006327f
C556 B.n516 VSUBS 0.006327f
C557 B.n517 VSUBS 0.006327f
C558 B.n518 VSUBS 0.006327f
C559 B.n519 VSUBS 0.006327f
C560 B.n520 VSUBS 0.006327f
C561 B.n521 VSUBS 0.006327f
C562 B.n522 VSUBS 0.006327f
C563 B.n523 VSUBS 0.006327f
C564 B.n524 VSUBS 0.006327f
C565 B.n525 VSUBS 0.006327f
C566 B.n526 VSUBS 0.006327f
C567 B.n527 VSUBS 0.006327f
C568 B.n528 VSUBS 0.006327f
C569 B.n529 VSUBS 0.006327f
C570 B.n530 VSUBS 0.006327f
C571 B.n531 VSUBS 0.006327f
C572 B.n532 VSUBS 0.006327f
C573 B.n533 VSUBS 0.006327f
C574 B.n534 VSUBS 0.006327f
C575 B.n535 VSUBS 0.006327f
C576 B.n536 VSUBS 0.006327f
C577 B.n537 VSUBS 0.006327f
C578 B.n538 VSUBS 0.006327f
C579 B.n539 VSUBS 0.006327f
C580 B.n540 VSUBS 0.006327f
C581 B.n541 VSUBS 0.006327f
C582 B.n542 VSUBS 0.006327f
C583 B.n543 VSUBS 0.006327f
C584 B.n544 VSUBS 0.01471f
C585 B.n545 VSUBS 0.013761f
C586 B.n546 VSUBS 0.013761f
C587 B.n547 VSUBS 0.006327f
C588 B.n548 VSUBS 0.006327f
C589 B.n549 VSUBS 0.006327f
C590 B.n550 VSUBS 0.006327f
C591 B.n551 VSUBS 0.006327f
C592 B.n552 VSUBS 0.006327f
C593 B.n553 VSUBS 0.006327f
C594 B.n554 VSUBS 0.006327f
C595 B.n555 VSUBS 0.006327f
C596 B.n556 VSUBS 0.006327f
C597 B.n557 VSUBS 0.006327f
C598 B.n558 VSUBS 0.006327f
C599 B.n559 VSUBS 0.006327f
C600 B.n560 VSUBS 0.006327f
C601 B.n561 VSUBS 0.006327f
C602 B.n562 VSUBS 0.006327f
C603 B.n563 VSUBS 0.006327f
C604 B.n564 VSUBS 0.006327f
C605 B.n565 VSUBS 0.006327f
C606 B.n566 VSUBS 0.006327f
C607 B.n567 VSUBS 0.006327f
C608 B.n568 VSUBS 0.006327f
C609 B.n569 VSUBS 0.006327f
C610 B.n570 VSUBS 0.006327f
C611 B.n571 VSUBS 0.006327f
C612 B.n572 VSUBS 0.006327f
C613 B.n573 VSUBS 0.006327f
C614 B.n574 VSUBS 0.006327f
C615 B.n575 VSUBS 0.006327f
C616 B.n576 VSUBS 0.006327f
C617 B.n577 VSUBS 0.006327f
C618 B.n578 VSUBS 0.006327f
C619 B.n579 VSUBS 0.014326f
C620 VDD1.n0 VSUBS 0.011467f
C621 VDD1.n1 VSUBS 0.025854f
C622 VDD1.n2 VSUBS 0.011582f
C623 VDD1.n3 VSUBS 0.020356f
C624 VDD1.n4 VSUBS 0.010938f
C625 VDD1.n5 VSUBS 0.025854f
C626 VDD1.n6 VSUBS 0.011582f
C627 VDD1.n7 VSUBS 0.020356f
C628 VDD1.n8 VSUBS 0.010938f
C629 VDD1.n9 VSUBS 0.025854f
C630 VDD1.n10 VSUBS 0.011582f
C631 VDD1.n11 VSUBS 0.020356f
C632 VDD1.n12 VSUBS 0.010938f
C633 VDD1.n13 VSUBS 0.025854f
C634 VDD1.n14 VSUBS 0.011582f
C635 VDD1.n15 VSUBS 0.020356f
C636 VDD1.n16 VSUBS 0.010938f
C637 VDD1.n17 VSUBS 0.025854f
C638 VDD1.n18 VSUBS 0.011582f
C639 VDD1.n19 VSUBS 0.020356f
C640 VDD1.n20 VSUBS 0.010938f
C641 VDD1.n21 VSUBS 0.01939f
C642 VDD1.n22 VSUBS 0.016447f
C643 VDD1.t1 VSUBS 0.055231f
C644 VDD1.n23 VSUBS 0.129441f
C645 VDD1.n24 VSUBS 1.0835f
C646 VDD1.n25 VSUBS 0.010938f
C647 VDD1.n26 VSUBS 0.011582f
C648 VDD1.n27 VSUBS 0.025854f
C649 VDD1.n28 VSUBS 0.025854f
C650 VDD1.n29 VSUBS 0.011582f
C651 VDD1.n30 VSUBS 0.010938f
C652 VDD1.n31 VSUBS 0.020356f
C653 VDD1.n32 VSUBS 0.020356f
C654 VDD1.n33 VSUBS 0.010938f
C655 VDD1.n34 VSUBS 0.011582f
C656 VDD1.n35 VSUBS 0.025854f
C657 VDD1.n36 VSUBS 0.025854f
C658 VDD1.n37 VSUBS 0.011582f
C659 VDD1.n38 VSUBS 0.010938f
C660 VDD1.n39 VSUBS 0.020356f
C661 VDD1.n40 VSUBS 0.020356f
C662 VDD1.n41 VSUBS 0.010938f
C663 VDD1.n42 VSUBS 0.011582f
C664 VDD1.n43 VSUBS 0.025854f
C665 VDD1.n44 VSUBS 0.025854f
C666 VDD1.n45 VSUBS 0.011582f
C667 VDD1.n46 VSUBS 0.010938f
C668 VDD1.n47 VSUBS 0.020356f
C669 VDD1.n48 VSUBS 0.020356f
C670 VDD1.n49 VSUBS 0.010938f
C671 VDD1.n50 VSUBS 0.011582f
C672 VDD1.n51 VSUBS 0.025854f
C673 VDD1.n52 VSUBS 0.025854f
C674 VDD1.n53 VSUBS 0.011582f
C675 VDD1.n54 VSUBS 0.010938f
C676 VDD1.n55 VSUBS 0.020356f
C677 VDD1.n56 VSUBS 0.020356f
C678 VDD1.n57 VSUBS 0.010938f
C679 VDD1.n58 VSUBS 0.011582f
C680 VDD1.n59 VSUBS 0.025854f
C681 VDD1.n60 VSUBS 0.025854f
C682 VDD1.n61 VSUBS 0.011582f
C683 VDD1.n62 VSUBS 0.010938f
C684 VDD1.n63 VSUBS 0.020356f
C685 VDD1.n64 VSUBS 0.052056f
C686 VDD1.n65 VSUBS 0.010938f
C687 VDD1.n66 VSUBS 0.011582f
C688 VDD1.n67 VSUBS 0.058185f
C689 VDD1.n68 VSUBS 0.053365f
C690 VDD1.n69 VSUBS 0.011467f
C691 VDD1.n70 VSUBS 0.025854f
C692 VDD1.n71 VSUBS 0.011582f
C693 VDD1.n72 VSUBS 0.020356f
C694 VDD1.n73 VSUBS 0.010938f
C695 VDD1.n74 VSUBS 0.025854f
C696 VDD1.n75 VSUBS 0.011582f
C697 VDD1.n76 VSUBS 0.020356f
C698 VDD1.n77 VSUBS 0.010938f
C699 VDD1.n78 VSUBS 0.025854f
C700 VDD1.n79 VSUBS 0.011582f
C701 VDD1.n80 VSUBS 0.020356f
C702 VDD1.n81 VSUBS 0.010938f
C703 VDD1.n82 VSUBS 0.025854f
C704 VDD1.n83 VSUBS 0.011582f
C705 VDD1.n84 VSUBS 0.020356f
C706 VDD1.n85 VSUBS 0.010938f
C707 VDD1.n86 VSUBS 0.025854f
C708 VDD1.n87 VSUBS 0.011582f
C709 VDD1.n88 VSUBS 0.020356f
C710 VDD1.n89 VSUBS 0.010938f
C711 VDD1.n90 VSUBS 0.01939f
C712 VDD1.n91 VSUBS 0.016447f
C713 VDD1.t0 VSUBS 0.055231f
C714 VDD1.n92 VSUBS 0.129441f
C715 VDD1.n93 VSUBS 1.0835f
C716 VDD1.n94 VSUBS 0.010938f
C717 VDD1.n95 VSUBS 0.011582f
C718 VDD1.n96 VSUBS 0.025854f
C719 VDD1.n97 VSUBS 0.025854f
C720 VDD1.n98 VSUBS 0.011582f
C721 VDD1.n99 VSUBS 0.010938f
C722 VDD1.n100 VSUBS 0.020356f
C723 VDD1.n101 VSUBS 0.020356f
C724 VDD1.n102 VSUBS 0.010938f
C725 VDD1.n103 VSUBS 0.011582f
C726 VDD1.n104 VSUBS 0.025854f
C727 VDD1.n105 VSUBS 0.025854f
C728 VDD1.n106 VSUBS 0.011582f
C729 VDD1.n107 VSUBS 0.010938f
C730 VDD1.n108 VSUBS 0.020356f
C731 VDD1.n109 VSUBS 0.020356f
C732 VDD1.n110 VSUBS 0.010938f
C733 VDD1.n111 VSUBS 0.011582f
C734 VDD1.n112 VSUBS 0.025854f
C735 VDD1.n113 VSUBS 0.025854f
C736 VDD1.n114 VSUBS 0.011582f
C737 VDD1.n115 VSUBS 0.010938f
C738 VDD1.n116 VSUBS 0.020356f
C739 VDD1.n117 VSUBS 0.020356f
C740 VDD1.n118 VSUBS 0.010938f
C741 VDD1.n119 VSUBS 0.011582f
C742 VDD1.n120 VSUBS 0.025854f
C743 VDD1.n121 VSUBS 0.025854f
C744 VDD1.n122 VSUBS 0.011582f
C745 VDD1.n123 VSUBS 0.010938f
C746 VDD1.n124 VSUBS 0.020356f
C747 VDD1.n125 VSUBS 0.020356f
C748 VDD1.n126 VSUBS 0.010938f
C749 VDD1.n127 VSUBS 0.011582f
C750 VDD1.n128 VSUBS 0.025854f
C751 VDD1.n129 VSUBS 0.025854f
C752 VDD1.n130 VSUBS 0.011582f
C753 VDD1.n131 VSUBS 0.010938f
C754 VDD1.n132 VSUBS 0.020356f
C755 VDD1.n133 VSUBS 0.052056f
C756 VDD1.n134 VSUBS 0.010938f
C757 VDD1.n135 VSUBS 0.011582f
C758 VDD1.n136 VSUBS 0.058185f
C759 VDD1.n137 VSUBS 0.612149f
C760 VP.t0 VSUBS 4.14043f
C761 VP.t1 VSUBS 3.59989f
C762 VP.n0 VSUBS 5.68166f
C763 VDD2.n0 VSUBS 0.011291f
C764 VDD2.n1 VSUBS 0.025457f
C765 VDD2.n2 VSUBS 0.011404f
C766 VDD2.n3 VSUBS 0.020043f
C767 VDD2.n4 VSUBS 0.01077f
C768 VDD2.n5 VSUBS 0.025457f
C769 VDD2.n6 VSUBS 0.011404f
C770 VDD2.n7 VSUBS 0.020043f
C771 VDD2.n8 VSUBS 0.01077f
C772 VDD2.n9 VSUBS 0.025457f
C773 VDD2.n10 VSUBS 0.011404f
C774 VDD2.n11 VSUBS 0.020043f
C775 VDD2.n12 VSUBS 0.01077f
C776 VDD2.n13 VSUBS 0.025457f
C777 VDD2.n14 VSUBS 0.011404f
C778 VDD2.n15 VSUBS 0.020043f
C779 VDD2.n16 VSUBS 0.01077f
C780 VDD2.n17 VSUBS 0.025457f
C781 VDD2.n18 VSUBS 0.011404f
C782 VDD2.n19 VSUBS 0.020043f
C783 VDD2.n20 VSUBS 0.01077f
C784 VDD2.n21 VSUBS 0.019093f
C785 VDD2.n22 VSUBS 0.016194f
C786 VDD2.t1 VSUBS 0.054383f
C787 VDD2.n23 VSUBS 0.127453f
C788 VDD2.n24 VSUBS 1.06686f
C789 VDD2.n25 VSUBS 0.01077f
C790 VDD2.n26 VSUBS 0.011404f
C791 VDD2.n27 VSUBS 0.025457f
C792 VDD2.n28 VSUBS 0.025457f
C793 VDD2.n29 VSUBS 0.011404f
C794 VDD2.n30 VSUBS 0.01077f
C795 VDD2.n31 VSUBS 0.020043f
C796 VDD2.n32 VSUBS 0.020043f
C797 VDD2.n33 VSUBS 0.01077f
C798 VDD2.n34 VSUBS 0.011404f
C799 VDD2.n35 VSUBS 0.025457f
C800 VDD2.n36 VSUBS 0.025457f
C801 VDD2.n37 VSUBS 0.011404f
C802 VDD2.n38 VSUBS 0.01077f
C803 VDD2.n39 VSUBS 0.020043f
C804 VDD2.n40 VSUBS 0.020043f
C805 VDD2.n41 VSUBS 0.01077f
C806 VDD2.n42 VSUBS 0.011404f
C807 VDD2.n43 VSUBS 0.025457f
C808 VDD2.n44 VSUBS 0.025457f
C809 VDD2.n45 VSUBS 0.011404f
C810 VDD2.n46 VSUBS 0.01077f
C811 VDD2.n47 VSUBS 0.020043f
C812 VDD2.n48 VSUBS 0.020043f
C813 VDD2.n49 VSUBS 0.01077f
C814 VDD2.n50 VSUBS 0.011404f
C815 VDD2.n51 VSUBS 0.025457f
C816 VDD2.n52 VSUBS 0.025457f
C817 VDD2.n53 VSUBS 0.011404f
C818 VDD2.n54 VSUBS 0.01077f
C819 VDD2.n55 VSUBS 0.020043f
C820 VDD2.n56 VSUBS 0.020043f
C821 VDD2.n57 VSUBS 0.01077f
C822 VDD2.n58 VSUBS 0.011404f
C823 VDD2.n59 VSUBS 0.025457f
C824 VDD2.n60 VSUBS 0.025457f
C825 VDD2.n61 VSUBS 0.011404f
C826 VDD2.n62 VSUBS 0.01077f
C827 VDD2.n63 VSUBS 0.020043f
C828 VDD2.n64 VSUBS 0.051257f
C829 VDD2.n65 VSUBS 0.01077f
C830 VDD2.n66 VSUBS 0.011404f
C831 VDD2.n67 VSUBS 0.057291f
C832 VDD2.n68 VSUBS 0.567954f
C833 VDD2.n69 VSUBS 0.011291f
C834 VDD2.n70 VSUBS 0.025457f
C835 VDD2.n71 VSUBS 0.011404f
C836 VDD2.n72 VSUBS 0.020043f
C837 VDD2.n73 VSUBS 0.01077f
C838 VDD2.n74 VSUBS 0.025457f
C839 VDD2.n75 VSUBS 0.011404f
C840 VDD2.n76 VSUBS 0.020043f
C841 VDD2.n77 VSUBS 0.01077f
C842 VDD2.n78 VSUBS 0.025457f
C843 VDD2.n79 VSUBS 0.011404f
C844 VDD2.n80 VSUBS 0.020043f
C845 VDD2.n81 VSUBS 0.01077f
C846 VDD2.n82 VSUBS 0.025457f
C847 VDD2.n83 VSUBS 0.011404f
C848 VDD2.n84 VSUBS 0.020043f
C849 VDD2.n85 VSUBS 0.01077f
C850 VDD2.n86 VSUBS 0.025457f
C851 VDD2.n87 VSUBS 0.011404f
C852 VDD2.n88 VSUBS 0.020043f
C853 VDD2.n89 VSUBS 0.01077f
C854 VDD2.n90 VSUBS 0.019093f
C855 VDD2.n91 VSUBS 0.016194f
C856 VDD2.t0 VSUBS 0.054383f
C857 VDD2.n92 VSUBS 0.127453f
C858 VDD2.n93 VSUBS 1.06686f
C859 VDD2.n94 VSUBS 0.01077f
C860 VDD2.n95 VSUBS 0.011404f
C861 VDD2.n96 VSUBS 0.025457f
C862 VDD2.n97 VSUBS 0.025457f
C863 VDD2.n98 VSUBS 0.011404f
C864 VDD2.n99 VSUBS 0.01077f
C865 VDD2.n100 VSUBS 0.020043f
C866 VDD2.n101 VSUBS 0.020043f
C867 VDD2.n102 VSUBS 0.01077f
C868 VDD2.n103 VSUBS 0.011404f
C869 VDD2.n104 VSUBS 0.025457f
C870 VDD2.n105 VSUBS 0.025457f
C871 VDD2.n106 VSUBS 0.011404f
C872 VDD2.n107 VSUBS 0.01077f
C873 VDD2.n108 VSUBS 0.020043f
C874 VDD2.n109 VSUBS 0.020043f
C875 VDD2.n110 VSUBS 0.01077f
C876 VDD2.n111 VSUBS 0.011404f
C877 VDD2.n112 VSUBS 0.025457f
C878 VDD2.n113 VSUBS 0.025457f
C879 VDD2.n114 VSUBS 0.011404f
C880 VDD2.n115 VSUBS 0.01077f
C881 VDD2.n116 VSUBS 0.020043f
C882 VDD2.n117 VSUBS 0.020043f
C883 VDD2.n118 VSUBS 0.01077f
C884 VDD2.n119 VSUBS 0.011404f
C885 VDD2.n120 VSUBS 0.025457f
C886 VDD2.n121 VSUBS 0.025457f
C887 VDD2.n122 VSUBS 0.011404f
C888 VDD2.n123 VSUBS 0.01077f
C889 VDD2.n124 VSUBS 0.020043f
C890 VDD2.n125 VSUBS 0.020043f
C891 VDD2.n126 VSUBS 0.01077f
C892 VDD2.n127 VSUBS 0.011404f
C893 VDD2.n128 VSUBS 0.025457f
C894 VDD2.n129 VSUBS 0.025457f
C895 VDD2.n130 VSUBS 0.011404f
C896 VDD2.n131 VSUBS 0.01077f
C897 VDD2.n132 VSUBS 0.020043f
C898 VDD2.n133 VSUBS 0.051257f
C899 VDD2.n134 VSUBS 0.01077f
C900 VDD2.n135 VSUBS 0.011404f
C901 VDD2.n136 VSUBS 0.057291f
C902 VDD2.n137 VSUBS 0.051707f
C903 VDD2.n138 VSUBS 2.43538f
C904 VTAIL.n0 VSUBS 0.01634f
C905 VTAIL.n1 VSUBS 0.03684f
C906 VTAIL.n2 VSUBS 0.016503f
C907 VTAIL.n3 VSUBS 0.029005f
C908 VTAIL.n4 VSUBS 0.015586f
C909 VTAIL.n5 VSUBS 0.03684f
C910 VTAIL.n6 VSUBS 0.016503f
C911 VTAIL.n7 VSUBS 0.029005f
C912 VTAIL.n8 VSUBS 0.015586f
C913 VTAIL.n9 VSUBS 0.03684f
C914 VTAIL.n10 VSUBS 0.016503f
C915 VTAIL.n11 VSUBS 0.029005f
C916 VTAIL.n12 VSUBS 0.015586f
C917 VTAIL.n13 VSUBS 0.03684f
C918 VTAIL.n14 VSUBS 0.016503f
C919 VTAIL.n15 VSUBS 0.029005f
C920 VTAIL.n16 VSUBS 0.015586f
C921 VTAIL.n17 VSUBS 0.03684f
C922 VTAIL.n18 VSUBS 0.016503f
C923 VTAIL.n19 VSUBS 0.029005f
C924 VTAIL.n20 VSUBS 0.015586f
C925 VTAIL.n21 VSUBS 0.02763f
C926 VTAIL.n22 VSUBS 0.023436f
C927 VTAIL.t1 VSUBS 0.0787f
C928 VTAIL.n23 VSUBS 0.184442f
C929 VTAIL.n24 VSUBS 1.54389f
C930 VTAIL.n25 VSUBS 0.015586f
C931 VTAIL.n26 VSUBS 0.016503f
C932 VTAIL.n27 VSUBS 0.03684f
C933 VTAIL.n28 VSUBS 0.03684f
C934 VTAIL.n29 VSUBS 0.016503f
C935 VTAIL.n30 VSUBS 0.015586f
C936 VTAIL.n31 VSUBS 0.029005f
C937 VTAIL.n32 VSUBS 0.029005f
C938 VTAIL.n33 VSUBS 0.015586f
C939 VTAIL.n34 VSUBS 0.016503f
C940 VTAIL.n35 VSUBS 0.03684f
C941 VTAIL.n36 VSUBS 0.03684f
C942 VTAIL.n37 VSUBS 0.016503f
C943 VTAIL.n38 VSUBS 0.015586f
C944 VTAIL.n39 VSUBS 0.029005f
C945 VTAIL.n40 VSUBS 0.029005f
C946 VTAIL.n41 VSUBS 0.015586f
C947 VTAIL.n42 VSUBS 0.016503f
C948 VTAIL.n43 VSUBS 0.03684f
C949 VTAIL.n44 VSUBS 0.03684f
C950 VTAIL.n45 VSUBS 0.016503f
C951 VTAIL.n46 VSUBS 0.015586f
C952 VTAIL.n47 VSUBS 0.029005f
C953 VTAIL.n48 VSUBS 0.029005f
C954 VTAIL.n49 VSUBS 0.015586f
C955 VTAIL.n50 VSUBS 0.016503f
C956 VTAIL.n51 VSUBS 0.03684f
C957 VTAIL.n52 VSUBS 0.03684f
C958 VTAIL.n53 VSUBS 0.016503f
C959 VTAIL.n54 VSUBS 0.015586f
C960 VTAIL.n55 VSUBS 0.029005f
C961 VTAIL.n56 VSUBS 0.029005f
C962 VTAIL.n57 VSUBS 0.015586f
C963 VTAIL.n58 VSUBS 0.016503f
C964 VTAIL.n59 VSUBS 0.03684f
C965 VTAIL.n60 VSUBS 0.03684f
C966 VTAIL.n61 VSUBS 0.016503f
C967 VTAIL.n62 VSUBS 0.015586f
C968 VTAIL.n63 VSUBS 0.029005f
C969 VTAIL.n64 VSUBS 0.074175f
C970 VTAIL.n65 VSUBS 0.015586f
C971 VTAIL.n66 VSUBS 0.016503f
C972 VTAIL.n67 VSUBS 0.082908f
C973 VTAIL.n68 VSUBS 0.054845f
C974 VTAIL.n69 VSUBS 1.91953f
C975 VTAIL.n70 VSUBS 0.01634f
C976 VTAIL.n71 VSUBS 0.03684f
C977 VTAIL.n72 VSUBS 0.016503f
C978 VTAIL.n73 VSUBS 0.029005f
C979 VTAIL.n74 VSUBS 0.015586f
C980 VTAIL.n75 VSUBS 0.03684f
C981 VTAIL.n76 VSUBS 0.016503f
C982 VTAIL.n77 VSUBS 0.029005f
C983 VTAIL.n78 VSUBS 0.015586f
C984 VTAIL.n79 VSUBS 0.03684f
C985 VTAIL.n80 VSUBS 0.016503f
C986 VTAIL.n81 VSUBS 0.029005f
C987 VTAIL.n82 VSUBS 0.015586f
C988 VTAIL.n83 VSUBS 0.03684f
C989 VTAIL.n84 VSUBS 0.016503f
C990 VTAIL.n85 VSUBS 0.029005f
C991 VTAIL.n86 VSUBS 0.015586f
C992 VTAIL.n87 VSUBS 0.03684f
C993 VTAIL.n88 VSUBS 0.016503f
C994 VTAIL.n89 VSUBS 0.029005f
C995 VTAIL.n90 VSUBS 0.015586f
C996 VTAIL.n91 VSUBS 0.02763f
C997 VTAIL.n92 VSUBS 0.023436f
C998 VTAIL.t3 VSUBS 0.0787f
C999 VTAIL.n93 VSUBS 0.184442f
C1000 VTAIL.n94 VSUBS 1.54389f
C1001 VTAIL.n95 VSUBS 0.015586f
C1002 VTAIL.n96 VSUBS 0.016503f
C1003 VTAIL.n97 VSUBS 0.03684f
C1004 VTAIL.n98 VSUBS 0.03684f
C1005 VTAIL.n99 VSUBS 0.016503f
C1006 VTAIL.n100 VSUBS 0.015586f
C1007 VTAIL.n101 VSUBS 0.029005f
C1008 VTAIL.n102 VSUBS 0.029005f
C1009 VTAIL.n103 VSUBS 0.015586f
C1010 VTAIL.n104 VSUBS 0.016503f
C1011 VTAIL.n105 VSUBS 0.03684f
C1012 VTAIL.n106 VSUBS 0.03684f
C1013 VTAIL.n107 VSUBS 0.016503f
C1014 VTAIL.n108 VSUBS 0.015586f
C1015 VTAIL.n109 VSUBS 0.029005f
C1016 VTAIL.n110 VSUBS 0.029005f
C1017 VTAIL.n111 VSUBS 0.015586f
C1018 VTAIL.n112 VSUBS 0.016503f
C1019 VTAIL.n113 VSUBS 0.03684f
C1020 VTAIL.n114 VSUBS 0.03684f
C1021 VTAIL.n115 VSUBS 0.016503f
C1022 VTAIL.n116 VSUBS 0.015586f
C1023 VTAIL.n117 VSUBS 0.029005f
C1024 VTAIL.n118 VSUBS 0.029005f
C1025 VTAIL.n119 VSUBS 0.015586f
C1026 VTAIL.n120 VSUBS 0.016503f
C1027 VTAIL.n121 VSUBS 0.03684f
C1028 VTAIL.n122 VSUBS 0.03684f
C1029 VTAIL.n123 VSUBS 0.016503f
C1030 VTAIL.n124 VSUBS 0.015586f
C1031 VTAIL.n125 VSUBS 0.029005f
C1032 VTAIL.n126 VSUBS 0.029005f
C1033 VTAIL.n127 VSUBS 0.015586f
C1034 VTAIL.n128 VSUBS 0.016503f
C1035 VTAIL.n129 VSUBS 0.03684f
C1036 VTAIL.n130 VSUBS 0.03684f
C1037 VTAIL.n131 VSUBS 0.016503f
C1038 VTAIL.n132 VSUBS 0.015586f
C1039 VTAIL.n133 VSUBS 0.029005f
C1040 VTAIL.n134 VSUBS 0.074175f
C1041 VTAIL.n135 VSUBS 0.015586f
C1042 VTAIL.n136 VSUBS 0.016503f
C1043 VTAIL.n137 VSUBS 0.082908f
C1044 VTAIL.n138 VSUBS 0.054845f
C1045 VTAIL.n139 VSUBS 1.96162f
C1046 VTAIL.n140 VSUBS 0.01634f
C1047 VTAIL.n141 VSUBS 0.03684f
C1048 VTAIL.n142 VSUBS 0.016503f
C1049 VTAIL.n143 VSUBS 0.029005f
C1050 VTAIL.n144 VSUBS 0.015586f
C1051 VTAIL.n145 VSUBS 0.03684f
C1052 VTAIL.n146 VSUBS 0.016503f
C1053 VTAIL.n147 VSUBS 0.029005f
C1054 VTAIL.n148 VSUBS 0.015586f
C1055 VTAIL.n149 VSUBS 0.03684f
C1056 VTAIL.n150 VSUBS 0.016503f
C1057 VTAIL.n151 VSUBS 0.029005f
C1058 VTAIL.n152 VSUBS 0.015586f
C1059 VTAIL.n153 VSUBS 0.03684f
C1060 VTAIL.n154 VSUBS 0.016503f
C1061 VTAIL.n155 VSUBS 0.029005f
C1062 VTAIL.n156 VSUBS 0.015586f
C1063 VTAIL.n157 VSUBS 0.03684f
C1064 VTAIL.n158 VSUBS 0.016503f
C1065 VTAIL.n159 VSUBS 0.029005f
C1066 VTAIL.n160 VSUBS 0.015586f
C1067 VTAIL.n161 VSUBS 0.02763f
C1068 VTAIL.n162 VSUBS 0.023436f
C1069 VTAIL.t0 VSUBS 0.0787f
C1070 VTAIL.n163 VSUBS 0.184442f
C1071 VTAIL.n164 VSUBS 1.54389f
C1072 VTAIL.n165 VSUBS 0.015586f
C1073 VTAIL.n166 VSUBS 0.016503f
C1074 VTAIL.n167 VSUBS 0.03684f
C1075 VTAIL.n168 VSUBS 0.03684f
C1076 VTAIL.n169 VSUBS 0.016503f
C1077 VTAIL.n170 VSUBS 0.015586f
C1078 VTAIL.n171 VSUBS 0.029005f
C1079 VTAIL.n172 VSUBS 0.029005f
C1080 VTAIL.n173 VSUBS 0.015586f
C1081 VTAIL.n174 VSUBS 0.016503f
C1082 VTAIL.n175 VSUBS 0.03684f
C1083 VTAIL.n176 VSUBS 0.03684f
C1084 VTAIL.n177 VSUBS 0.016503f
C1085 VTAIL.n178 VSUBS 0.015586f
C1086 VTAIL.n179 VSUBS 0.029005f
C1087 VTAIL.n180 VSUBS 0.029005f
C1088 VTAIL.n181 VSUBS 0.015586f
C1089 VTAIL.n182 VSUBS 0.016503f
C1090 VTAIL.n183 VSUBS 0.03684f
C1091 VTAIL.n184 VSUBS 0.03684f
C1092 VTAIL.n185 VSUBS 0.016503f
C1093 VTAIL.n186 VSUBS 0.015586f
C1094 VTAIL.n187 VSUBS 0.029005f
C1095 VTAIL.n188 VSUBS 0.029005f
C1096 VTAIL.n189 VSUBS 0.015586f
C1097 VTAIL.n190 VSUBS 0.016503f
C1098 VTAIL.n191 VSUBS 0.03684f
C1099 VTAIL.n192 VSUBS 0.03684f
C1100 VTAIL.n193 VSUBS 0.016503f
C1101 VTAIL.n194 VSUBS 0.015586f
C1102 VTAIL.n195 VSUBS 0.029005f
C1103 VTAIL.n196 VSUBS 0.029005f
C1104 VTAIL.n197 VSUBS 0.015586f
C1105 VTAIL.n198 VSUBS 0.016503f
C1106 VTAIL.n199 VSUBS 0.03684f
C1107 VTAIL.n200 VSUBS 0.03684f
C1108 VTAIL.n201 VSUBS 0.016503f
C1109 VTAIL.n202 VSUBS 0.015586f
C1110 VTAIL.n203 VSUBS 0.029005f
C1111 VTAIL.n204 VSUBS 0.074175f
C1112 VTAIL.n205 VSUBS 0.015586f
C1113 VTAIL.n206 VSUBS 0.016503f
C1114 VTAIL.n207 VSUBS 0.082908f
C1115 VTAIL.n208 VSUBS 0.054845f
C1116 VTAIL.n209 VSUBS 1.77148f
C1117 VTAIL.n210 VSUBS 0.01634f
C1118 VTAIL.n211 VSUBS 0.03684f
C1119 VTAIL.n212 VSUBS 0.016503f
C1120 VTAIL.n213 VSUBS 0.029005f
C1121 VTAIL.n214 VSUBS 0.015586f
C1122 VTAIL.n215 VSUBS 0.03684f
C1123 VTAIL.n216 VSUBS 0.016503f
C1124 VTAIL.n217 VSUBS 0.029005f
C1125 VTAIL.n218 VSUBS 0.015586f
C1126 VTAIL.n219 VSUBS 0.03684f
C1127 VTAIL.n220 VSUBS 0.016503f
C1128 VTAIL.n221 VSUBS 0.029005f
C1129 VTAIL.n222 VSUBS 0.015586f
C1130 VTAIL.n223 VSUBS 0.03684f
C1131 VTAIL.n224 VSUBS 0.016503f
C1132 VTAIL.n225 VSUBS 0.029005f
C1133 VTAIL.n226 VSUBS 0.015586f
C1134 VTAIL.n227 VSUBS 0.03684f
C1135 VTAIL.n228 VSUBS 0.016503f
C1136 VTAIL.n229 VSUBS 0.029005f
C1137 VTAIL.n230 VSUBS 0.015586f
C1138 VTAIL.n231 VSUBS 0.02763f
C1139 VTAIL.n232 VSUBS 0.023436f
C1140 VTAIL.t2 VSUBS 0.0787f
C1141 VTAIL.n233 VSUBS 0.184442f
C1142 VTAIL.n234 VSUBS 1.54389f
C1143 VTAIL.n235 VSUBS 0.015586f
C1144 VTAIL.n236 VSUBS 0.016503f
C1145 VTAIL.n237 VSUBS 0.03684f
C1146 VTAIL.n238 VSUBS 0.03684f
C1147 VTAIL.n239 VSUBS 0.016503f
C1148 VTAIL.n240 VSUBS 0.015586f
C1149 VTAIL.n241 VSUBS 0.029005f
C1150 VTAIL.n242 VSUBS 0.029005f
C1151 VTAIL.n243 VSUBS 0.015586f
C1152 VTAIL.n244 VSUBS 0.016503f
C1153 VTAIL.n245 VSUBS 0.03684f
C1154 VTAIL.n246 VSUBS 0.03684f
C1155 VTAIL.n247 VSUBS 0.016503f
C1156 VTAIL.n248 VSUBS 0.015586f
C1157 VTAIL.n249 VSUBS 0.029005f
C1158 VTAIL.n250 VSUBS 0.029005f
C1159 VTAIL.n251 VSUBS 0.015586f
C1160 VTAIL.n252 VSUBS 0.016503f
C1161 VTAIL.n253 VSUBS 0.03684f
C1162 VTAIL.n254 VSUBS 0.03684f
C1163 VTAIL.n255 VSUBS 0.016503f
C1164 VTAIL.n256 VSUBS 0.015586f
C1165 VTAIL.n257 VSUBS 0.029005f
C1166 VTAIL.n258 VSUBS 0.029005f
C1167 VTAIL.n259 VSUBS 0.015586f
C1168 VTAIL.n260 VSUBS 0.016503f
C1169 VTAIL.n261 VSUBS 0.03684f
C1170 VTAIL.n262 VSUBS 0.03684f
C1171 VTAIL.n263 VSUBS 0.016503f
C1172 VTAIL.n264 VSUBS 0.015586f
C1173 VTAIL.n265 VSUBS 0.029005f
C1174 VTAIL.n266 VSUBS 0.029005f
C1175 VTAIL.n267 VSUBS 0.015586f
C1176 VTAIL.n268 VSUBS 0.016503f
C1177 VTAIL.n269 VSUBS 0.03684f
C1178 VTAIL.n270 VSUBS 0.03684f
C1179 VTAIL.n271 VSUBS 0.016503f
C1180 VTAIL.n272 VSUBS 0.015586f
C1181 VTAIL.n273 VSUBS 0.029005f
C1182 VTAIL.n274 VSUBS 0.074175f
C1183 VTAIL.n275 VSUBS 0.015586f
C1184 VTAIL.n276 VSUBS 0.016503f
C1185 VTAIL.n277 VSUBS 0.082908f
C1186 VTAIL.n278 VSUBS 0.054845f
C1187 VTAIL.n279 VSUBS 1.6746f
C1188 VN.t0 VSUBS 3.47794f
C1189 VN.t1 VSUBS 4.0041f
.ends

