* NGSPICE file created from diff_pair_sample_0989.ext - technology: sky130A

.subckt diff_pair_sample_0989 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t3 w_n2534_n4764# sky130_fd_pr__pfet_01v8 ad=7.4022 pd=38.74 as=7.4022 ps=38.74 w=18.98 l=3.58
X1 VDD1.t0 VP.t1 VTAIL.t2 w_n2534_n4764# sky130_fd_pr__pfet_01v8 ad=7.4022 pd=38.74 as=7.4022 ps=38.74 w=18.98 l=3.58
X2 VDD2.t1 VN.t0 VTAIL.t1 w_n2534_n4764# sky130_fd_pr__pfet_01v8 ad=7.4022 pd=38.74 as=7.4022 ps=38.74 w=18.98 l=3.58
X3 B.t11 B.t9 B.t10 w_n2534_n4764# sky130_fd_pr__pfet_01v8 ad=7.4022 pd=38.74 as=0 ps=0 w=18.98 l=3.58
X4 VDD2.t0 VN.t1 VTAIL.t0 w_n2534_n4764# sky130_fd_pr__pfet_01v8 ad=7.4022 pd=38.74 as=7.4022 ps=38.74 w=18.98 l=3.58
X5 B.t8 B.t6 B.t7 w_n2534_n4764# sky130_fd_pr__pfet_01v8 ad=7.4022 pd=38.74 as=0 ps=0 w=18.98 l=3.58
X6 B.t5 B.t3 B.t4 w_n2534_n4764# sky130_fd_pr__pfet_01v8 ad=7.4022 pd=38.74 as=0 ps=0 w=18.98 l=3.58
X7 B.t2 B.t0 B.t1 w_n2534_n4764# sky130_fd_pr__pfet_01v8 ad=7.4022 pd=38.74 as=0 ps=0 w=18.98 l=3.58
R0 VP.n0 VP.t0 219.16
R1 VP.n0 VP.t1 166.617
R2 VP VP.n0 0.526373
R3 VTAIL.n418 VTAIL.n318 756.745
R4 VTAIL.n100 VTAIL.n0 756.745
R5 VTAIL.n312 VTAIL.n212 756.745
R6 VTAIL.n206 VTAIL.n106 756.745
R7 VTAIL.n353 VTAIL.n352 585
R8 VTAIL.n350 VTAIL.n349 585
R9 VTAIL.n359 VTAIL.n358 585
R10 VTAIL.n361 VTAIL.n360 585
R11 VTAIL.n346 VTAIL.n345 585
R12 VTAIL.n367 VTAIL.n366 585
R13 VTAIL.n369 VTAIL.n368 585
R14 VTAIL.n342 VTAIL.n341 585
R15 VTAIL.n375 VTAIL.n374 585
R16 VTAIL.n377 VTAIL.n376 585
R17 VTAIL.n338 VTAIL.n337 585
R18 VTAIL.n383 VTAIL.n382 585
R19 VTAIL.n385 VTAIL.n384 585
R20 VTAIL.n334 VTAIL.n333 585
R21 VTAIL.n391 VTAIL.n390 585
R22 VTAIL.n394 VTAIL.n393 585
R23 VTAIL.n392 VTAIL.n330 585
R24 VTAIL.n399 VTAIL.n329 585
R25 VTAIL.n401 VTAIL.n400 585
R26 VTAIL.n403 VTAIL.n402 585
R27 VTAIL.n326 VTAIL.n325 585
R28 VTAIL.n409 VTAIL.n408 585
R29 VTAIL.n411 VTAIL.n410 585
R30 VTAIL.n322 VTAIL.n321 585
R31 VTAIL.n417 VTAIL.n416 585
R32 VTAIL.n419 VTAIL.n418 585
R33 VTAIL.n35 VTAIL.n34 585
R34 VTAIL.n32 VTAIL.n31 585
R35 VTAIL.n41 VTAIL.n40 585
R36 VTAIL.n43 VTAIL.n42 585
R37 VTAIL.n28 VTAIL.n27 585
R38 VTAIL.n49 VTAIL.n48 585
R39 VTAIL.n51 VTAIL.n50 585
R40 VTAIL.n24 VTAIL.n23 585
R41 VTAIL.n57 VTAIL.n56 585
R42 VTAIL.n59 VTAIL.n58 585
R43 VTAIL.n20 VTAIL.n19 585
R44 VTAIL.n65 VTAIL.n64 585
R45 VTAIL.n67 VTAIL.n66 585
R46 VTAIL.n16 VTAIL.n15 585
R47 VTAIL.n73 VTAIL.n72 585
R48 VTAIL.n76 VTAIL.n75 585
R49 VTAIL.n74 VTAIL.n12 585
R50 VTAIL.n81 VTAIL.n11 585
R51 VTAIL.n83 VTAIL.n82 585
R52 VTAIL.n85 VTAIL.n84 585
R53 VTAIL.n8 VTAIL.n7 585
R54 VTAIL.n91 VTAIL.n90 585
R55 VTAIL.n93 VTAIL.n92 585
R56 VTAIL.n4 VTAIL.n3 585
R57 VTAIL.n99 VTAIL.n98 585
R58 VTAIL.n101 VTAIL.n100 585
R59 VTAIL.n313 VTAIL.n312 585
R60 VTAIL.n311 VTAIL.n310 585
R61 VTAIL.n216 VTAIL.n215 585
R62 VTAIL.n305 VTAIL.n304 585
R63 VTAIL.n303 VTAIL.n302 585
R64 VTAIL.n220 VTAIL.n219 585
R65 VTAIL.n297 VTAIL.n296 585
R66 VTAIL.n295 VTAIL.n294 585
R67 VTAIL.n293 VTAIL.n223 585
R68 VTAIL.n227 VTAIL.n224 585
R69 VTAIL.n288 VTAIL.n287 585
R70 VTAIL.n286 VTAIL.n285 585
R71 VTAIL.n229 VTAIL.n228 585
R72 VTAIL.n280 VTAIL.n279 585
R73 VTAIL.n278 VTAIL.n277 585
R74 VTAIL.n233 VTAIL.n232 585
R75 VTAIL.n272 VTAIL.n271 585
R76 VTAIL.n270 VTAIL.n269 585
R77 VTAIL.n237 VTAIL.n236 585
R78 VTAIL.n264 VTAIL.n263 585
R79 VTAIL.n262 VTAIL.n261 585
R80 VTAIL.n241 VTAIL.n240 585
R81 VTAIL.n256 VTAIL.n255 585
R82 VTAIL.n254 VTAIL.n253 585
R83 VTAIL.n245 VTAIL.n244 585
R84 VTAIL.n248 VTAIL.n247 585
R85 VTAIL.n207 VTAIL.n206 585
R86 VTAIL.n205 VTAIL.n204 585
R87 VTAIL.n110 VTAIL.n109 585
R88 VTAIL.n199 VTAIL.n198 585
R89 VTAIL.n197 VTAIL.n196 585
R90 VTAIL.n114 VTAIL.n113 585
R91 VTAIL.n191 VTAIL.n190 585
R92 VTAIL.n189 VTAIL.n188 585
R93 VTAIL.n187 VTAIL.n117 585
R94 VTAIL.n121 VTAIL.n118 585
R95 VTAIL.n182 VTAIL.n181 585
R96 VTAIL.n180 VTAIL.n179 585
R97 VTAIL.n123 VTAIL.n122 585
R98 VTAIL.n174 VTAIL.n173 585
R99 VTAIL.n172 VTAIL.n171 585
R100 VTAIL.n127 VTAIL.n126 585
R101 VTAIL.n166 VTAIL.n165 585
R102 VTAIL.n164 VTAIL.n163 585
R103 VTAIL.n131 VTAIL.n130 585
R104 VTAIL.n158 VTAIL.n157 585
R105 VTAIL.n156 VTAIL.n155 585
R106 VTAIL.n135 VTAIL.n134 585
R107 VTAIL.n150 VTAIL.n149 585
R108 VTAIL.n148 VTAIL.n147 585
R109 VTAIL.n139 VTAIL.n138 585
R110 VTAIL.n142 VTAIL.n141 585
R111 VTAIL.t3 VTAIL.n246 327.466
R112 VTAIL.t1 VTAIL.n140 327.466
R113 VTAIL.t0 VTAIL.n351 327.466
R114 VTAIL.t2 VTAIL.n33 327.466
R115 VTAIL.n352 VTAIL.n349 171.744
R116 VTAIL.n359 VTAIL.n349 171.744
R117 VTAIL.n360 VTAIL.n359 171.744
R118 VTAIL.n360 VTAIL.n345 171.744
R119 VTAIL.n367 VTAIL.n345 171.744
R120 VTAIL.n368 VTAIL.n367 171.744
R121 VTAIL.n368 VTAIL.n341 171.744
R122 VTAIL.n375 VTAIL.n341 171.744
R123 VTAIL.n376 VTAIL.n375 171.744
R124 VTAIL.n376 VTAIL.n337 171.744
R125 VTAIL.n383 VTAIL.n337 171.744
R126 VTAIL.n384 VTAIL.n383 171.744
R127 VTAIL.n384 VTAIL.n333 171.744
R128 VTAIL.n391 VTAIL.n333 171.744
R129 VTAIL.n393 VTAIL.n391 171.744
R130 VTAIL.n393 VTAIL.n392 171.744
R131 VTAIL.n392 VTAIL.n329 171.744
R132 VTAIL.n401 VTAIL.n329 171.744
R133 VTAIL.n402 VTAIL.n401 171.744
R134 VTAIL.n402 VTAIL.n325 171.744
R135 VTAIL.n409 VTAIL.n325 171.744
R136 VTAIL.n410 VTAIL.n409 171.744
R137 VTAIL.n410 VTAIL.n321 171.744
R138 VTAIL.n417 VTAIL.n321 171.744
R139 VTAIL.n418 VTAIL.n417 171.744
R140 VTAIL.n34 VTAIL.n31 171.744
R141 VTAIL.n41 VTAIL.n31 171.744
R142 VTAIL.n42 VTAIL.n41 171.744
R143 VTAIL.n42 VTAIL.n27 171.744
R144 VTAIL.n49 VTAIL.n27 171.744
R145 VTAIL.n50 VTAIL.n49 171.744
R146 VTAIL.n50 VTAIL.n23 171.744
R147 VTAIL.n57 VTAIL.n23 171.744
R148 VTAIL.n58 VTAIL.n57 171.744
R149 VTAIL.n58 VTAIL.n19 171.744
R150 VTAIL.n65 VTAIL.n19 171.744
R151 VTAIL.n66 VTAIL.n65 171.744
R152 VTAIL.n66 VTAIL.n15 171.744
R153 VTAIL.n73 VTAIL.n15 171.744
R154 VTAIL.n75 VTAIL.n73 171.744
R155 VTAIL.n75 VTAIL.n74 171.744
R156 VTAIL.n74 VTAIL.n11 171.744
R157 VTAIL.n83 VTAIL.n11 171.744
R158 VTAIL.n84 VTAIL.n83 171.744
R159 VTAIL.n84 VTAIL.n7 171.744
R160 VTAIL.n91 VTAIL.n7 171.744
R161 VTAIL.n92 VTAIL.n91 171.744
R162 VTAIL.n92 VTAIL.n3 171.744
R163 VTAIL.n99 VTAIL.n3 171.744
R164 VTAIL.n100 VTAIL.n99 171.744
R165 VTAIL.n312 VTAIL.n311 171.744
R166 VTAIL.n311 VTAIL.n215 171.744
R167 VTAIL.n304 VTAIL.n215 171.744
R168 VTAIL.n304 VTAIL.n303 171.744
R169 VTAIL.n303 VTAIL.n219 171.744
R170 VTAIL.n296 VTAIL.n219 171.744
R171 VTAIL.n296 VTAIL.n295 171.744
R172 VTAIL.n295 VTAIL.n223 171.744
R173 VTAIL.n227 VTAIL.n223 171.744
R174 VTAIL.n287 VTAIL.n227 171.744
R175 VTAIL.n287 VTAIL.n286 171.744
R176 VTAIL.n286 VTAIL.n228 171.744
R177 VTAIL.n279 VTAIL.n228 171.744
R178 VTAIL.n279 VTAIL.n278 171.744
R179 VTAIL.n278 VTAIL.n232 171.744
R180 VTAIL.n271 VTAIL.n232 171.744
R181 VTAIL.n271 VTAIL.n270 171.744
R182 VTAIL.n270 VTAIL.n236 171.744
R183 VTAIL.n263 VTAIL.n236 171.744
R184 VTAIL.n263 VTAIL.n262 171.744
R185 VTAIL.n262 VTAIL.n240 171.744
R186 VTAIL.n255 VTAIL.n240 171.744
R187 VTAIL.n255 VTAIL.n254 171.744
R188 VTAIL.n254 VTAIL.n244 171.744
R189 VTAIL.n247 VTAIL.n244 171.744
R190 VTAIL.n206 VTAIL.n205 171.744
R191 VTAIL.n205 VTAIL.n109 171.744
R192 VTAIL.n198 VTAIL.n109 171.744
R193 VTAIL.n198 VTAIL.n197 171.744
R194 VTAIL.n197 VTAIL.n113 171.744
R195 VTAIL.n190 VTAIL.n113 171.744
R196 VTAIL.n190 VTAIL.n189 171.744
R197 VTAIL.n189 VTAIL.n117 171.744
R198 VTAIL.n121 VTAIL.n117 171.744
R199 VTAIL.n181 VTAIL.n121 171.744
R200 VTAIL.n181 VTAIL.n180 171.744
R201 VTAIL.n180 VTAIL.n122 171.744
R202 VTAIL.n173 VTAIL.n122 171.744
R203 VTAIL.n173 VTAIL.n172 171.744
R204 VTAIL.n172 VTAIL.n126 171.744
R205 VTAIL.n165 VTAIL.n126 171.744
R206 VTAIL.n165 VTAIL.n164 171.744
R207 VTAIL.n164 VTAIL.n130 171.744
R208 VTAIL.n157 VTAIL.n130 171.744
R209 VTAIL.n157 VTAIL.n156 171.744
R210 VTAIL.n156 VTAIL.n134 171.744
R211 VTAIL.n149 VTAIL.n134 171.744
R212 VTAIL.n149 VTAIL.n148 171.744
R213 VTAIL.n148 VTAIL.n138 171.744
R214 VTAIL.n141 VTAIL.n138 171.744
R215 VTAIL.n352 VTAIL.t0 85.8723
R216 VTAIL.n34 VTAIL.t2 85.8723
R217 VTAIL.n247 VTAIL.t3 85.8723
R218 VTAIL.n141 VTAIL.t1 85.8723
R219 VTAIL.n211 VTAIL.n105 35.4703
R220 VTAIL.n423 VTAIL.n422 32.5732
R221 VTAIL.n105 VTAIL.n104 32.5732
R222 VTAIL.n317 VTAIL.n316 32.5732
R223 VTAIL.n211 VTAIL.n210 32.5732
R224 VTAIL.n423 VTAIL.n317 32.0996
R225 VTAIL.n353 VTAIL.n351 16.3895
R226 VTAIL.n35 VTAIL.n33 16.3895
R227 VTAIL.n248 VTAIL.n246 16.3895
R228 VTAIL.n142 VTAIL.n140 16.3895
R229 VTAIL.n400 VTAIL.n399 13.1884
R230 VTAIL.n82 VTAIL.n81 13.1884
R231 VTAIL.n294 VTAIL.n293 13.1884
R232 VTAIL.n188 VTAIL.n187 13.1884
R233 VTAIL.n354 VTAIL.n350 12.8005
R234 VTAIL.n398 VTAIL.n330 12.8005
R235 VTAIL.n403 VTAIL.n328 12.8005
R236 VTAIL.n36 VTAIL.n32 12.8005
R237 VTAIL.n80 VTAIL.n12 12.8005
R238 VTAIL.n85 VTAIL.n10 12.8005
R239 VTAIL.n297 VTAIL.n222 12.8005
R240 VTAIL.n292 VTAIL.n224 12.8005
R241 VTAIL.n249 VTAIL.n245 12.8005
R242 VTAIL.n191 VTAIL.n116 12.8005
R243 VTAIL.n186 VTAIL.n118 12.8005
R244 VTAIL.n143 VTAIL.n139 12.8005
R245 VTAIL.n358 VTAIL.n357 12.0247
R246 VTAIL.n395 VTAIL.n394 12.0247
R247 VTAIL.n404 VTAIL.n326 12.0247
R248 VTAIL.n40 VTAIL.n39 12.0247
R249 VTAIL.n77 VTAIL.n76 12.0247
R250 VTAIL.n86 VTAIL.n8 12.0247
R251 VTAIL.n298 VTAIL.n220 12.0247
R252 VTAIL.n289 VTAIL.n288 12.0247
R253 VTAIL.n253 VTAIL.n252 12.0247
R254 VTAIL.n192 VTAIL.n114 12.0247
R255 VTAIL.n183 VTAIL.n182 12.0247
R256 VTAIL.n147 VTAIL.n146 12.0247
R257 VTAIL.n361 VTAIL.n348 11.249
R258 VTAIL.n390 VTAIL.n332 11.249
R259 VTAIL.n408 VTAIL.n407 11.249
R260 VTAIL.n43 VTAIL.n30 11.249
R261 VTAIL.n72 VTAIL.n14 11.249
R262 VTAIL.n90 VTAIL.n89 11.249
R263 VTAIL.n302 VTAIL.n301 11.249
R264 VTAIL.n285 VTAIL.n226 11.249
R265 VTAIL.n256 VTAIL.n243 11.249
R266 VTAIL.n196 VTAIL.n195 11.249
R267 VTAIL.n179 VTAIL.n120 11.249
R268 VTAIL.n150 VTAIL.n137 11.249
R269 VTAIL.n362 VTAIL.n346 10.4732
R270 VTAIL.n389 VTAIL.n334 10.4732
R271 VTAIL.n411 VTAIL.n324 10.4732
R272 VTAIL.n44 VTAIL.n28 10.4732
R273 VTAIL.n71 VTAIL.n16 10.4732
R274 VTAIL.n93 VTAIL.n6 10.4732
R275 VTAIL.n305 VTAIL.n218 10.4732
R276 VTAIL.n284 VTAIL.n229 10.4732
R277 VTAIL.n257 VTAIL.n241 10.4732
R278 VTAIL.n199 VTAIL.n112 10.4732
R279 VTAIL.n178 VTAIL.n123 10.4732
R280 VTAIL.n151 VTAIL.n135 10.4732
R281 VTAIL.n366 VTAIL.n365 9.69747
R282 VTAIL.n386 VTAIL.n385 9.69747
R283 VTAIL.n412 VTAIL.n322 9.69747
R284 VTAIL.n48 VTAIL.n47 9.69747
R285 VTAIL.n68 VTAIL.n67 9.69747
R286 VTAIL.n94 VTAIL.n4 9.69747
R287 VTAIL.n306 VTAIL.n216 9.69747
R288 VTAIL.n281 VTAIL.n280 9.69747
R289 VTAIL.n261 VTAIL.n260 9.69747
R290 VTAIL.n200 VTAIL.n110 9.69747
R291 VTAIL.n175 VTAIL.n174 9.69747
R292 VTAIL.n155 VTAIL.n154 9.69747
R293 VTAIL.n422 VTAIL.n421 9.45567
R294 VTAIL.n104 VTAIL.n103 9.45567
R295 VTAIL.n316 VTAIL.n315 9.45567
R296 VTAIL.n210 VTAIL.n209 9.45567
R297 VTAIL.n320 VTAIL.n319 9.3005
R298 VTAIL.n415 VTAIL.n414 9.3005
R299 VTAIL.n413 VTAIL.n412 9.3005
R300 VTAIL.n324 VTAIL.n323 9.3005
R301 VTAIL.n407 VTAIL.n406 9.3005
R302 VTAIL.n405 VTAIL.n404 9.3005
R303 VTAIL.n328 VTAIL.n327 9.3005
R304 VTAIL.n373 VTAIL.n372 9.3005
R305 VTAIL.n371 VTAIL.n370 9.3005
R306 VTAIL.n344 VTAIL.n343 9.3005
R307 VTAIL.n365 VTAIL.n364 9.3005
R308 VTAIL.n363 VTAIL.n362 9.3005
R309 VTAIL.n348 VTAIL.n347 9.3005
R310 VTAIL.n357 VTAIL.n356 9.3005
R311 VTAIL.n355 VTAIL.n354 9.3005
R312 VTAIL.n340 VTAIL.n339 9.3005
R313 VTAIL.n379 VTAIL.n378 9.3005
R314 VTAIL.n381 VTAIL.n380 9.3005
R315 VTAIL.n336 VTAIL.n335 9.3005
R316 VTAIL.n387 VTAIL.n386 9.3005
R317 VTAIL.n389 VTAIL.n388 9.3005
R318 VTAIL.n332 VTAIL.n331 9.3005
R319 VTAIL.n396 VTAIL.n395 9.3005
R320 VTAIL.n398 VTAIL.n397 9.3005
R321 VTAIL.n421 VTAIL.n420 9.3005
R322 VTAIL.n2 VTAIL.n1 9.3005
R323 VTAIL.n97 VTAIL.n96 9.3005
R324 VTAIL.n95 VTAIL.n94 9.3005
R325 VTAIL.n6 VTAIL.n5 9.3005
R326 VTAIL.n89 VTAIL.n88 9.3005
R327 VTAIL.n87 VTAIL.n86 9.3005
R328 VTAIL.n10 VTAIL.n9 9.3005
R329 VTAIL.n55 VTAIL.n54 9.3005
R330 VTAIL.n53 VTAIL.n52 9.3005
R331 VTAIL.n26 VTAIL.n25 9.3005
R332 VTAIL.n47 VTAIL.n46 9.3005
R333 VTAIL.n45 VTAIL.n44 9.3005
R334 VTAIL.n30 VTAIL.n29 9.3005
R335 VTAIL.n39 VTAIL.n38 9.3005
R336 VTAIL.n37 VTAIL.n36 9.3005
R337 VTAIL.n22 VTAIL.n21 9.3005
R338 VTAIL.n61 VTAIL.n60 9.3005
R339 VTAIL.n63 VTAIL.n62 9.3005
R340 VTAIL.n18 VTAIL.n17 9.3005
R341 VTAIL.n69 VTAIL.n68 9.3005
R342 VTAIL.n71 VTAIL.n70 9.3005
R343 VTAIL.n14 VTAIL.n13 9.3005
R344 VTAIL.n78 VTAIL.n77 9.3005
R345 VTAIL.n80 VTAIL.n79 9.3005
R346 VTAIL.n103 VTAIL.n102 9.3005
R347 VTAIL.n274 VTAIL.n273 9.3005
R348 VTAIL.n276 VTAIL.n275 9.3005
R349 VTAIL.n231 VTAIL.n230 9.3005
R350 VTAIL.n282 VTAIL.n281 9.3005
R351 VTAIL.n284 VTAIL.n283 9.3005
R352 VTAIL.n226 VTAIL.n225 9.3005
R353 VTAIL.n290 VTAIL.n289 9.3005
R354 VTAIL.n292 VTAIL.n291 9.3005
R355 VTAIL.n315 VTAIL.n314 9.3005
R356 VTAIL.n214 VTAIL.n213 9.3005
R357 VTAIL.n309 VTAIL.n308 9.3005
R358 VTAIL.n307 VTAIL.n306 9.3005
R359 VTAIL.n218 VTAIL.n217 9.3005
R360 VTAIL.n301 VTAIL.n300 9.3005
R361 VTAIL.n299 VTAIL.n298 9.3005
R362 VTAIL.n222 VTAIL.n221 9.3005
R363 VTAIL.n235 VTAIL.n234 9.3005
R364 VTAIL.n268 VTAIL.n267 9.3005
R365 VTAIL.n266 VTAIL.n265 9.3005
R366 VTAIL.n239 VTAIL.n238 9.3005
R367 VTAIL.n260 VTAIL.n259 9.3005
R368 VTAIL.n258 VTAIL.n257 9.3005
R369 VTAIL.n243 VTAIL.n242 9.3005
R370 VTAIL.n252 VTAIL.n251 9.3005
R371 VTAIL.n250 VTAIL.n249 9.3005
R372 VTAIL.n168 VTAIL.n167 9.3005
R373 VTAIL.n170 VTAIL.n169 9.3005
R374 VTAIL.n125 VTAIL.n124 9.3005
R375 VTAIL.n176 VTAIL.n175 9.3005
R376 VTAIL.n178 VTAIL.n177 9.3005
R377 VTAIL.n120 VTAIL.n119 9.3005
R378 VTAIL.n184 VTAIL.n183 9.3005
R379 VTAIL.n186 VTAIL.n185 9.3005
R380 VTAIL.n209 VTAIL.n208 9.3005
R381 VTAIL.n108 VTAIL.n107 9.3005
R382 VTAIL.n203 VTAIL.n202 9.3005
R383 VTAIL.n201 VTAIL.n200 9.3005
R384 VTAIL.n112 VTAIL.n111 9.3005
R385 VTAIL.n195 VTAIL.n194 9.3005
R386 VTAIL.n193 VTAIL.n192 9.3005
R387 VTAIL.n116 VTAIL.n115 9.3005
R388 VTAIL.n129 VTAIL.n128 9.3005
R389 VTAIL.n162 VTAIL.n161 9.3005
R390 VTAIL.n160 VTAIL.n159 9.3005
R391 VTAIL.n133 VTAIL.n132 9.3005
R392 VTAIL.n154 VTAIL.n153 9.3005
R393 VTAIL.n152 VTAIL.n151 9.3005
R394 VTAIL.n137 VTAIL.n136 9.3005
R395 VTAIL.n146 VTAIL.n145 9.3005
R396 VTAIL.n144 VTAIL.n143 9.3005
R397 VTAIL.n369 VTAIL.n344 8.92171
R398 VTAIL.n382 VTAIL.n336 8.92171
R399 VTAIL.n416 VTAIL.n415 8.92171
R400 VTAIL.n51 VTAIL.n26 8.92171
R401 VTAIL.n64 VTAIL.n18 8.92171
R402 VTAIL.n98 VTAIL.n97 8.92171
R403 VTAIL.n310 VTAIL.n309 8.92171
R404 VTAIL.n277 VTAIL.n231 8.92171
R405 VTAIL.n264 VTAIL.n239 8.92171
R406 VTAIL.n204 VTAIL.n203 8.92171
R407 VTAIL.n171 VTAIL.n125 8.92171
R408 VTAIL.n158 VTAIL.n133 8.92171
R409 VTAIL.n370 VTAIL.n342 8.14595
R410 VTAIL.n381 VTAIL.n338 8.14595
R411 VTAIL.n419 VTAIL.n320 8.14595
R412 VTAIL.n52 VTAIL.n24 8.14595
R413 VTAIL.n63 VTAIL.n20 8.14595
R414 VTAIL.n101 VTAIL.n2 8.14595
R415 VTAIL.n313 VTAIL.n214 8.14595
R416 VTAIL.n276 VTAIL.n233 8.14595
R417 VTAIL.n265 VTAIL.n237 8.14595
R418 VTAIL.n207 VTAIL.n108 8.14595
R419 VTAIL.n170 VTAIL.n127 8.14595
R420 VTAIL.n159 VTAIL.n131 8.14595
R421 VTAIL.n374 VTAIL.n373 7.3702
R422 VTAIL.n378 VTAIL.n377 7.3702
R423 VTAIL.n420 VTAIL.n318 7.3702
R424 VTAIL.n56 VTAIL.n55 7.3702
R425 VTAIL.n60 VTAIL.n59 7.3702
R426 VTAIL.n102 VTAIL.n0 7.3702
R427 VTAIL.n314 VTAIL.n212 7.3702
R428 VTAIL.n273 VTAIL.n272 7.3702
R429 VTAIL.n269 VTAIL.n268 7.3702
R430 VTAIL.n208 VTAIL.n106 7.3702
R431 VTAIL.n167 VTAIL.n166 7.3702
R432 VTAIL.n163 VTAIL.n162 7.3702
R433 VTAIL.n374 VTAIL.n340 6.59444
R434 VTAIL.n377 VTAIL.n340 6.59444
R435 VTAIL.n422 VTAIL.n318 6.59444
R436 VTAIL.n56 VTAIL.n22 6.59444
R437 VTAIL.n59 VTAIL.n22 6.59444
R438 VTAIL.n104 VTAIL.n0 6.59444
R439 VTAIL.n316 VTAIL.n212 6.59444
R440 VTAIL.n272 VTAIL.n235 6.59444
R441 VTAIL.n269 VTAIL.n235 6.59444
R442 VTAIL.n210 VTAIL.n106 6.59444
R443 VTAIL.n166 VTAIL.n129 6.59444
R444 VTAIL.n163 VTAIL.n129 6.59444
R445 VTAIL.n373 VTAIL.n342 5.81868
R446 VTAIL.n378 VTAIL.n338 5.81868
R447 VTAIL.n420 VTAIL.n419 5.81868
R448 VTAIL.n55 VTAIL.n24 5.81868
R449 VTAIL.n60 VTAIL.n20 5.81868
R450 VTAIL.n102 VTAIL.n101 5.81868
R451 VTAIL.n314 VTAIL.n313 5.81868
R452 VTAIL.n273 VTAIL.n233 5.81868
R453 VTAIL.n268 VTAIL.n237 5.81868
R454 VTAIL.n208 VTAIL.n207 5.81868
R455 VTAIL.n167 VTAIL.n127 5.81868
R456 VTAIL.n162 VTAIL.n131 5.81868
R457 VTAIL.n370 VTAIL.n369 5.04292
R458 VTAIL.n382 VTAIL.n381 5.04292
R459 VTAIL.n416 VTAIL.n320 5.04292
R460 VTAIL.n52 VTAIL.n51 5.04292
R461 VTAIL.n64 VTAIL.n63 5.04292
R462 VTAIL.n98 VTAIL.n2 5.04292
R463 VTAIL.n310 VTAIL.n214 5.04292
R464 VTAIL.n277 VTAIL.n276 5.04292
R465 VTAIL.n265 VTAIL.n264 5.04292
R466 VTAIL.n204 VTAIL.n108 5.04292
R467 VTAIL.n171 VTAIL.n170 5.04292
R468 VTAIL.n159 VTAIL.n158 5.04292
R469 VTAIL.n366 VTAIL.n344 4.26717
R470 VTAIL.n385 VTAIL.n336 4.26717
R471 VTAIL.n415 VTAIL.n322 4.26717
R472 VTAIL.n48 VTAIL.n26 4.26717
R473 VTAIL.n67 VTAIL.n18 4.26717
R474 VTAIL.n97 VTAIL.n4 4.26717
R475 VTAIL.n309 VTAIL.n216 4.26717
R476 VTAIL.n280 VTAIL.n231 4.26717
R477 VTAIL.n261 VTAIL.n239 4.26717
R478 VTAIL.n203 VTAIL.n110 4.26717
R479 VTAIL.n174 VTAIL.n125 4.26717
R480 VTAIL.n155 VTAIL.n133 4.26717
R481 VTAIL.n355 VTAIL.n351 3.70982
R482 VTAIL.n37 VTAIL.n33 3.70982
R483 VTAIL.n250 VTAIL.n246 3.70982
R484 VTAIL.n144 VTAIL.n140 3.70982
R485 VTAIL.n365 VTAIL.n346 3.49141
R486 VTAIL.n386 VTAIL.n334 3.49141
R487 VTAIL.n412 VTAIL.n411 3.49141
R488 VTAIL.n47 VTAIL.n28 3.49141
R489 VTAIL.n68 VTAIL.n16 3.49141
R490 VTAIL.n94 VTAIL.n93 3.49141
R491 VTAIL.n306 VTAIL.n305 3.49141
R492 VTAIL.n281 VTAIL.n229 3.49141
R493 VTAIL.n260 VTAIL.n241 3.49141
R494 VTAIL.n200 VTAIL.n199 3.49141
R495 VTAIL.n175 VTAIL.n123 3.49141
R496 VTAIL.n154 VTAIL.n135 3.49141
R497 VTAIL.n362 VTAIL.n361 2.71565
R498 VTAIL.n390 VTAIL.n389 2.71565
R499 VTAIL.n408 VTAIL.n324 2.71565
R500 VTAIL.n44 VTAIL.n43 2.71565
R501 VTAIL.n72 VTAIL.n71 2.71565
R502 VTAIL.n90 VTAIL.n6 2.71565
R503 VTAIL.n302 VTAIL.n218 2.71565
R504 VTAIL.n285 VTAIL.n284 2.71565
R505 VTAIL.n257 VTAIL.n256 2.71565
R506 VTAIL.n196 VTAIL.n112 2.71565
R507 VTAIL.n179 VTAIL.n178 2.71565
R508 VTAIL.n151 VTAIL.n150 2.71565
R509 VTAIL.n317 VTAIL.n211 2.15567
R510 VTAIL.n358 VTAIL.n348 1.93989
R511 VTAIL.n394 VTAIL.n332 1.93989
R512 VTAIL.n407 VTAIL.n326 1.93989
R513 VTAIL.n40 VTAIL.n30 1.93989
R514 VTAIL.n76 VTAIL.n14 1.93989
R515 VTAIL.n89 VTAIL.n8 1.93989
R516 VTAIL.n301 VTAIL.n220 1.93989
R517 VTAIL.n288 VTAIL.n226 1.93989
R518 VTAIL.n253 VTAIL.n243 1.93989
R519 VTAIL.n195 VTAIL.n114 1.93989
R520 VTAIL.n182 VTAIL.n120 1.93989
R521 VTAIL.n147 VTAIL.n137 1.93989
R522 VTAIL VTAIL.n105 1.37119
R523 VTAIL.n357 VTAIL.n350 1.16414
R524 VTAIL.n395 VTAIL.n330 1.16414
R525 VTAIL.n404 VTAIL.n403 1.16414
R526 VTAIL.n39 VTAIL.n32 1.16414
R527 VTAIL.n77 VTAIL.n12 1.16414
R528 VTAIL.n86 VTAIL.n85 1.16414
R529 VTAIL.n298 VTAIL.n297 1.16414
R530 VTAIL.n289 VTAIL.n224 1.16414
R531 VTAIL.n252 VTAIL.n245 1.16414
R532 VTAIL.n192 VTAIL.n191 1.16414
R533 VTAIL.n183 VTAIL.n118 1.16414
R534 VTAIL.n146 VTAIL.n139 1.16414
R535 VTAIL VTAIL.n423 0.784983
R536 VTAIL.n354 VTAIL.n353 0.388379
R537 VTAIL.n399 VTAIL.n398 0.388379
R538 VTAIL.n400 VTAIL.n328 0.388379
R539 VTAIL.n36 VTAIL.n35 0.388379
R540 VTAIL.n81 VTAIL.n80 0.388379
R541 VTAIL.n82 VTAIL.n10 0.388379
R542 VTAIL.n294 VTAIL.n222 0.388379
R543 VTAIL.n293 VTAIL.n292 0.388379
R544 VTAIL.n249 VTAIL.n248 0.388379
R545 VTAIL.n188 VTAIL.n116 0.388379
R546 VTAIL.n187 VTAIL.n186 0.388379
R547 VTAIL.n143 VTAIL.n142 0.388379
R548 VTAIL.n356 VTAIL.n355 0.155672
R549 VTAIL.n356 VTAIL.n347 0.155672
R550 VTAIL.n363 VTAIL.n347 0.155672
R551 VTAIL.n364 VTAIL.n363 0.155672
R552 VTAIL.n364 VTAIL.n343 0.155672
R553 VTAIL.n371 VTAIL.n343 0.155672
R554 VTAIL.n372 VTAIL.n371 0.155672
R555 VTAIL.n372 VTAIL.n339 0.155672
R556 VTAIL.n379 VTAIL.n339 0.155672
R557 VTAIL.n380 VTAIL.n379 0.155672
R558 VTAIL.n380 VTAIL.n335 0.155672
R559 VTAIL.n387 VTAIL.n335 0.155672
R560 VTAIL.n388 VTAIL.n387 0.155672
R561 VTAIL.n388 VTAIL.n331 0.155672
R562 VTAIL.n396 VTAIL.n331 0.155672
R563 VTAIL.n397 VTAIL.n396 0.155672
R564 VTAIL.n397 VTAIL.n327 0.155672
R565 VTAIL.n405 VTAIL.n327 0.155672
R566 VTAIL.n406 VTAIL.n405 0.155672
R567 VTAIL.n406 VTAIL.n323 0.155672
R568 VTAIL.n413 VTAIL.n323 0.155672
R569 VTAIL.n414 VTAIL.n413 0.155672
R570 VTAIL.n414 VTAIL.n319 0.155672
R571 VTAIL.n421 VTAIL.n319 0.155672
R572 VTAIL.n38 VTAIL.n37 0.155672
R573 VTAIL.n38 VTAIL.n29 0.155672
R574 VTAIL.n45 VTAIL.n29 0.155672
R575 VTAIL.n46 VTAIL.n45 0.155672
R576 VTAIL.n46 VTAIL.n25 0.155672
R577 VTAIL.n53 VTAIL.n25 0.155672
R578 VTAIL.n54 VTAIL.n53 0.155672
R579 VTAIL.n54 VTAIL.n21 0.155672
R580 VTAIL.n61 VTAIL.n21 0.155672
R581 VTAIL.n62 VTAIL.n61 0.155672
R582 VTAIL.n62 VTAIL.n17 0.155672
R583 VTAIL.n69 VTAIL.n17 0.155672
R584 VTAIL.n70 VTAIL.n69 0.155672
R585 VTAIL.n70 VTAIL.n13 0.155672
R586 VTAIL.n78 VTAIL.n13 0.155672
R587 VTAIL.n79 VTAIL.n78 0.155672
R588 VTAIL.n79 VTAIL.n9 0.155672
R589 VTAIL.n87 VTAIL.n9 0.155672
R590 VTAIL.n88 VTAIL.n87 0.155672
R591 VTAIL.n88 VTAIL.n5 0.155672
R592 VTAIL.n95 VTAIL.n5 0.155672
R593 VTAIL.n96 VTAIL.n95 0.155672
R594 VTAIL.n96 VTAIL.n1 0.155672
R595 VTAIL.n103 VTAIL.n1 0.155672
R596 VTAIL.n315 VTAIL.n213 0.155672
R597 VTAIL.n308 VTAIL.n213 0.155672
R598 VTAIL.n308 VTAIL.n307 0.155672
R599 VTAIL.n307 VTAIL.n217 0.155672
R600 VTAIL.n300 VTAIL.n217 0.155672
R601 VTAIL.n300 VTAIL.n299 0.155672
R602 VTAIL.n299 VTAIL.n221 0.155672
R603 VTAIL.n291 VTAIL.n221 0.155672
R604 VTAIL.n291 VTAIL.n290 0.155672
R605 VTAIL.n290 VTAIL.n225 0.155672
R606 VTAIL.n283 VTAIL.n225 0.155672
R607 VTAIL.n283 VTAIL.n282 0.155672
R608 VTAIL.n282 VTAIL.n230 0.155672
R609 VTAIL.n275 VTAIL.n230 0.155672
R610 VTAIL.n275 VTAIL.n274 0.155672
R611 VTAIL.n274 VTAIL.n234 0.155672
R612 VTAIL.n267 VTAIL.n234 0.155672
R613 VTAIL.n267 VTAIL.n266 0.155672
R614 VTAIL.n266 VTAIL.n238 0.155672
R615 VTAIL.n259 VTAIL.n238 0.155672
R616 VTAIL.n259 VTAIL.n258 0.155672
R617 VTAIL.n258 VTAIL.n242 0.155672
R618 VTAIL.n251 VTAIL.n242 0.155672
R619 VTAIL.n251 VTAIL.n250 0.155672
R620 VTAIL.n209 VTAIL.n107 0.155672
R621 VTAIL.n202 VTAIL.n107 0.155672
R622 VTAIL.n202 VTAIL.n201 0.155672
R623 VTAIL.n201 VTAIL.n111 0.155672
R624 VTAIL.n194 VTAIL.n111 0.155672
R625 VTAIL.n194 VTAIL.n193 0.155672
R626 VTAIL.n193 VTAIL.n115 0.155672
R627 VTAIL.n185 VTAIL.n115 0.155672
R628 VTAIL.n185 VTAIL.n184 0.155672
R629 VTAIL.n184 VTAIL.n119 0.155672
R630 VTAIL.n177 VTAIL.n119 0.155672
R631 VTAIL.n177 VTAIL.n176 0.155672
R632 VTAIL.n176 VTAIL.n124 0.155672
R633 VTAIL.n169 VTAIL.n124 0.155672
R634 VTAIL.n169 VTAIL.n168 0.155672
R635 VTAIL.n168 VTAIL.n128 0.155672
R636 VTAIL.n161 VTAIL.n128 0.155672
R637 VTAIL.n161 VTAIL.n160 0.155672
R638 VTAIL.n160 VTAIL.n132 0.155672
R639 VTAIL.n153 VTAIL.n132 0.155672
R640 VTAIL.n153 VTAIL.n152 0.155672
R641 VTAIL.n152 VTAIL.n136 0.155672
R642 VTAIL.n145 VTAIL.n136 0.155672
R643 VTAIL.n145 VTAIL.n144 0.155672
R644 VDD1.n100 VDD1.n0 756.745
R645 VDD1.n205 VDD1.n105 756.745
R646 VDD1.n101 VDD1.n100 585
R647 VDD1.n99 VDD1.n98 585
R648 VDD1.n4 VDD1.n3 585
R649 VDD1.n93 VDD1.n92 585
R650 VDD1.n91 VDD1.n90 585
R651 VDD1.n8 VDD1.n7 585
R652 VDD1.n85 VDD1.n84 585
R653 VDD1.n83 VDD1.n82 585
R654 VDD1.n81 VDD1.n11 585
R655 VDD1.n15 VDD1.n12 585
R656 VDD1.n76 VDD1.n75 585
R657 VDD1.n74 VDD1.n73 585
R658 VDD1.n17 VDD1.n16 585
R659 VDD1.n68 VDD1.n67 585
R660 VDD1.n66 VDD1.n65 585
R661 VDD1.n21 VDD1.n20 585
R662 VDD1.n60 VDD1.n59 585
R663 VDD1.n58 VDD1.n57 585
R664 VDD1.n25 VDD1.n24 585
R665 VDD1.n52 VDD1.n51 585
R666 VDD1.n50 VDD1.n49 585
R667 VDD1.n29 VDD1.n28 585
R668 VDD1.n44 VDD1.n43 585
R669 VDD1.n42 VDD1.n41 585
R670 VDD1.n33 VDD1.n32 585
R671 VDD1.n36 VDD1.n35 585
R672 VDD1.n140 VDD1.n139 585
R673 VDD1.n137 VDD1.n136 585
R674 VDD1.n146 VDD1.n145 585
R675 VDD1.n148 VDD1.n147 585
R676 VDD1.n133 VDD1.n132 585
R677 VDD1.n154 VDD1.n153 585
R678 VDD1.n156 VDD1.n155 585
R679 VDD1.n129 VDD1.n128 585
R680 VDD1.n162 VDD1.n161 585
R681 VDD1.n164 VDD1.n163 585
R682 VDD1.n125 VDD1.n124 585
R683 VDD1.n170 VDD1.n169 585
R684 VDD1.n172 VDD1.n171 585
R685 VDD1.n121 VDD1.n120 585
R686 VDD1.n178 VDD1.n177 585
R687 VDD1.n181 VDD1.n180 585
R688 VDD1.n179 VDD1.n117 585
R689 VDD1.n186 VDD1.n116 585
R690 VDD1.n188 VDD1.n187 585
R691 VDD1.n190 VDD1.n189 585
R692 VDD1.n113 VDD1.n112 585
R693 VDD1.n196 VDD1.n195 585
R694 VDD1.n198 VDD1.n197 585
R695 VDD1.n109 VDD1.n108 585
R696 VDD1.n204 VDD1.n203 585
R697 VDD1.n206 VDD1.n205 585
R698 VDD1.t1 VDD1.n34 327.466
R699 VDD1.t0 VDD1.n138 327.466
R700 VDD1.n100 VDD1.n99 171.744
R701 VDD1.n99 VDD1.n3 171.744
R702 VDD1.n92 VDD1.n3 171.744
R703 VDD1.n92 VDD1.n91 171.744
R704 VDD1.n91 VDD1.n7 171.744
R705 VDD1.n84 VDD1.n7 171.744
R706 VDD1.n84 VDD1.n83 171.744
R707 VDD1.n83 VDD1.n11 171.744
R708 VDD1.n15 VDD1.n11 171.744
R709 VDD1.n75 VDD1.n15 171.744
R710 VDD1.n75 VDD1.n74 171.744
R711 VDD1.n74 VDD1.n16 171.744
R712 VDD1.n67 VDD1.n16 171.744
R713 VDD1.n67 VDD1.n66 171.744
R714 VDD1.n66 VDD1.n20 171.744
R715 VDD1.n59 VDD1.n20 171.744
R716 VDD1.n59 VDD1.n58 171.744
R717 VDD1.n58 VDD1.n24 171.744
R718 VDD1.n51 VDD1.n24 171.744
R719 VDD1.n51 VDD1.n50 171.744
R720 VDD1.n50 VDD1.n28 171.744
R721 VDD1.n43 VDD1.n28 171.744
R722 VDD1.n43 VDD1.n42 171.744
R723 VDD1.n42 VDD1.n32 171.744
R724 VDD1.n35 VDD1.n32 171.744
R725 VDD1.n139 VDD1.n136 171.744
R726 VDD1.n146 VDD1.n136 171.744
R727 VDD1.n147 VDD1.n146 171.744
R728 VDD1.n147 VDD1.n132 171.744
R729 VDD1.n154 VDD1.n132 171.744
R730 VDD1.n155 VDD1.n154 171.744
R731 VDD1.n155 VDD1.n128 171.744
R732 VDD1.n162 VDD1.n128 171.744
R733 VDD1.n163 VDD1.n162 171.744
R734 VDD1.n163 VDD1.n124 171.744
R735 VDD1.n170 VDD1.n124 171.744
R736 VDD1.n171 VDD1.n170 171.744
R737 VDD1.n171 VDD1.n120 171.744
R738 VDD1.n178 VDD1.n120 171.744
R739 VDD1.n180 VDD1.n178 171.744
R740 VDD1.n180 VDD1.n179 171.744
R741 VDD1.n179 VDD1.n116 171.744
R742 VDD1.n188 VDD1.n116 171.744
R743 VDD1.n189 VDD1.n188 171.744
R744 VDD1.n189 VDD1.n112 171.744
R745 VDD1.n196 VDD1.n112 171.744
R746 VDD1.n197 VDD1.n196 171.744
R747 VDD1.n197 VDD1.n108 171.744
R748 VDD1.n204 VDD1.n108 171.744
R749 VDD1.n205 VDD1.n204 171.744
R750 VDD1 VDD1.n209 97.3824
R751 VDD1.n35 VDD1.t1 85.8723
R752 VDD1.n139 VDD1.t0 85.8723
R753 VDD1 VDD1.n104 50.1529
R754 VDD1.n36 VDD1.n34 16.3895
R755 VDD1.n140 VDD1.n138 16.3895
R756 VDD1.n82 VDD1.n81 13.1884
R757 VDD1.n187 VDD1.n186 13.1884
R758 VDD1.n85 VDD1.n10 12.8005
R759 VDD1.n80 VDD1.n12 12.8005
R760 VDD1.n37 VDD1.n33 12.8005
R761 VDD1.n141 VDD1.n137 12.8005
R762 VDD1.n185 VDD1.n117 12.8005
R763 VDD1.n190 VDD1.n115 12.8005
R764 VDD1.n86 VDD1.n8 12.0247
R765 VDD1.n77 VDD1.n76 12.0247
R766 VDD1.n41 VDD1.n40 12.0247
R767 VDD1.n145 VDD1.n144 12.0247
R768 VDD1.n182 VDD1.n181 12.0247
R769 VDD1.n191 VDD1.n113 12.0247
R770 VDD1.n90 VDD1.n89 11.249
R771 VDD1.n73 VDD1.n14 11.249
R772 VDD1.n44 VDD1.n31 11.249
R773 VDD1.n148 VDD1.n135 11.249
R774 VDD1.n177 VDD1.n119 11.249
R775 VDD1.n195 VDD1.n194 11.249
R776 VDD1.n93 VDD1.n6 10.4732
R777 VDD1.n72 VDD1.n17 10.4732
R778 VDD1.n45 VDD1.n29 10.4732
R779 VDD1.n149 VDD1.n133 10.4732
R780 VDD1.n176 VDD1.n121 10.4732
R781 VDD1.n198 VDD1.n111 10.4732
R782 VDD1.n94 VDD1.n4 9.69747
R783 VDD1.n69 VDD1.n68 9.69747
R784 VDD1.n49 VDD1.n48 9.69747
R785 VDD1.n153 VDD1.n152 9.69747
R786 VDD1.n173 VDD1.n172 9.69747
R787 VDD1.n199 VDD1.n109 9.69747
R788 VDD1.n104 VDD1.n103 9.45567
R789 VDD1.n209 VDD1.n208 9.45567
R790 VDD1.n62 VDD1.n61 9.3005
R791 VDD1.n64 VDD1.n63 9.3005
R792 VDD1.n19 VDD1.n18 9.3005
R793 VDD1.n70 VDD1.n69 9.3005
R794 VDD1.n72 VDD1.n71 9.3005
R795 VDD1.n14 VDD1.n13 9.3005
R796 VDD1.n78 VDD1.n77 9.3005
R797 VDD1.n80 VDD1.n79 9.3005
R798 VDD1.n103 VDD1.n102 9.3005
R799 VDD1.n2 VDD1.n1 9.3005
R800 VDD1.n97 VDD1.n96 9.3005
R801 VDD1.n95 VDD1.n94 9.3005
R802 VDD1.n6 VDD1.n5 9.3005
R803 VDD1.n89 VDD1.n88 9.3005
R804 VDD1.n87 VDD1.n86 9.3005
R805 VDD1.n10 VDD1.n9 9.3005
R806 VDD1.n23 VDD1.n22 9.3005
R807 VDD1.n56 VDD1.n55 9.3005
R808 VDD1.n54 VDD1.n53 9.3005
R809 VDD1.n27 VDD1.n26 9.3005
R810 VDD1.n48 VDD1.n47 9.3005
R811 VDD1.n46 VDD1.n45 9.3005
R812 VDD1.n31 VDD1.n30 9.3005
R813 VDD1.n40 VDD1.n39 9.3005
R814 VDD1.n38 VDD1.n37 9.3005
R815 VDD1.n107 VDD1.n106 9.3005
R816 VDD1.n202 VDD1.n201 9.3005
R817 VDD1.n200 VDD1.n199 9.3005
R818 VDD1.n111 VDD1.n110 9.3005
R819 VDD1.n194 VDD1.n193 9.3005
R820 VDD1.n192 VDD1.n191 9.3005
R821 VDD1.n115 VDD1.n114 9.3005
R822 VDD1.n160 VDD1.n159 9.3005
R823 VDD1.n158 VDD1.n157 9.3005
R824 VDD1.n131 VDD1.n130 9.3005
R825 VDD1.n152 VDD1.n151 9.3005
R826 VDD1.n150 VDD1.n149 9.3005
R827 VDD1.n135 VDD1.n134 9.3005
R828 VDD1.n144 VDD1.n143 9.3005
R829 VDD1.n142 VDD1.n141 9.3005
R830 VDD1.n127 VDD1.n126 9.3005
R831 VDD1.n166 VDD1.n165 9.3005
R832 VDD1.n168 VDD1.n167 9.3005
R833 VDD1.n123 VDD1.n122 9.3005
R834 VDD1.n174 VDD1.n173 9.3005
R835 VDD1.n176 VDD1.n175 9.3005
R836 VDD1.n119 VDD1.n118 9.3005
R837 VDD1.n183 VDD1.n182 9.3005
R838 VDD1.n185 VDD1.n184 9.3005
R839 VDD1.n208 VDD1.n207 9.3005
R840 VDD1.n98 VDD1.n97 8.92171
R841 VDD1.n65 VDD1.n19 8.92171
R842 VDD1.n52 VDD1.n27 8.92171
R843 VDD1.n156 VDD1.n131 8.92171
R844 VDD1.n169 VDD1.n123 8.92171
R845 VDD1.n203 VDD1.n202 8.92171
R846 VDD1.n101 VDD1.n2 8.14595
R847 VDD1.n64 VDD1.n21 8.14595
R848 VDD1.n53 VDD1.n25 8.14595
R849 VDD1.n157 VDD1.n129 8.14595
R850 VDD1.n168 VDD1.n125 8.14595
R851 VDD1.n206 VDD1.n107 8.14595
R852 VDD1.n102 VDD1.n0 7.3702
R853 VDD1.n61 VDD1.n60 7.3702
R854 VDD1.n57 VDD1.n56 7.3702
R855 VDD1.n161 VDD1.n160 7.3702
R856 VDD1.n165 VDD1.n164 7.3702
R857 VDD1.n207 VDD1.n105 7.3702
R858 VDD1.n104 VDD1.n0 6.59444
R859 VDD1.n60 VDD1.n23 6.59444
R860 VDD1.n57 VDD1.n23 6.59444
R861 VDD1.n161 VDD1.n127 6.59444
R862 VDD1.n164 VDD1.n127 6.59444
R863 VDD1.n209 VDD1.n105 6.59444
R864 VDD1.n102 VDD1.n101 5.81868
R865 VDD1.n61 VDD1.n21 5.81868
R866 VDD1.n56 VDD1.n25 5.81868
R867 VDD1.n160 VDD1.n129 5.81868
R868 VDD1.n165 VDD1.n125 5.81868
R869 VDD1.n207 VDD1.n206 5.81868
R870 VDD1.n98 VDD1.n2 5.04292
R871 VDD1.n65 VDD1.n64 5.04292
R872 VDD1.n53 VDD1.n52 5.04292
R873 VDD1.n157 VDD1.n156 5.04292
R874 VDD1.n169 VDD1.n168 5.04292
R875 VDD1.n203 VDD1.n107 5.04292
R876 VDD1.n97 VDD1.n4 4.26717
R877 VDD1.n68 VDD1.n19 4.26717
R878 VDD1.n49 VDD1.n27 4.26717
R879 VDD1.n153 VDD1.n131 4.26717
R880 VDD1.n172 VDD1.n123 4.26717
R881 VDD1.n202 VDD1.n109 4.26717
R882 VDD1.n38 VDD1.n34 3.70982
R883 VDD1.n142 VDD1.n138 3.70982
R884 VDD1.n94 VDD1.n93 3.49141
R885 VDD1.n69 VDD1.n17 3.49141
R886 VDD1.n48 VDD1.n29 3.49141
R887 VDD1.n152 VDD1.n133 3.49141
R888 VDD1.n173 VDD1.n121 3.49141
R889 VDD1.n199 VDD1.n198 3.49141
R890 VDD1.n90 VDD1.n6 2.71565
R891 VDD1.n73 VDD1.n72 2.71565
R892 VDD1.n45 VDD1.n44 2.71565
R893 VDD1.n149 VDD1.n148 2.71565
R894 VDD1.n177 VDD1.n176 2.71565
R895 VDD1.n195 VDD1.n111 2.71565
R896 VDD1.n89 VDD1.n8 1.93989
R897 VDD1.n76 VDD1.n14 1.93989
R898 VDD1.n41 VDD1.n31 1.93989
R899 VDD1.n145 VDD1.n135 1.93989
R900 VDD1.n181 VDD1.n119 1.93989
R901 VDD1.n194 VDD1.n113 1.93989
R902 VDD1.n86 VDD1.n85 1.16414
R903 VDD1.n77 VDD1.n12 1.16414
R904 VDD1.n40 VDD1.n33 1.16414
R905 VDD1.n144 VDD1.n137 1.16414
R906 VDD1.n182 VDD1.n117 1.16414
R907 VDD1.n191 VDD1.n190 1.16414
R908 VDD1.n82 VDD1.n10 0.388379
R909 VDD1.n81 VDD1.n80 0.388379
R910 VDD1.n37 VDD1.n36 0.388379
R911 VDD1.n141 VDD1.n140 0.388379
R912 VDD1.n186 VDD1.n185 0.388379
R913 VDD1.n187 VDD1.n115 0.388379
R914 VDD1.n103 VDD1.n1 0.155672
R915 VDD1.n96 VDD1.n1 0.155672
R916 VDD1.n96 VDD1.n95 0.155672
R917 VDD1.n95 VDD1.n5 0.155672
R918 VDD1.n88 VDD1.n5 0.155672
R919 VDD1.n88 VDD1.n87 0.155672
R920 VDD1.n87 VDD1.n9 0.155672
R921 VDD1.n79 VDD1.n9 0.155672
R922 VDD1.n79 VDD1.n78 0.155672
R923 VDD1.n78 VDD1.n13 0.155672
R924 VDD1.n71 VDD1.n13 0.155672
R925 VDD1.n71 VDD1.n70 0.155672
R926 VDD1.n70 VDD1.n18 0.155672
R927 VDD1.n63 VDD1.n18 0.155672
R928 VDD1.n63 VDD1.n62 0.155672
R929 VDD1.n62 VDD1.n22 0.155672
R930 VDD1.n55 VDD1.n22 0.155672
R931 VDD1.n55 VDD1.n54 0.155672
R932 VDD1.n54 VDD1.n26 0.155672
R933 VDD1.n47 VDD1.n26 0.155672
R934 VDD1.n47 VDD1.n46 0.155672
R935 VDD1.n46 VDD1.n30 0.155672
R936 VDD1.n39 VDD1.n30 0.155672
R937 VDD1.n39 VDD1.n38 0.155672
R938 VDD1.n143 VDD1.n142 0.155672
R939 VDD1.n143 VDD1.n134 0.155672
R940 VDD1.n150 VDD1.n134 0.155672
R941 VDD1.n151 VDD1.n150 0.155672
R942 VDD1.n151 VDD1.n130 0.155672
R943 VDD1.n158 VDD1.n130 0.155672
R944 VDD1.n159 VDD1.n158 0.155672
R945 VDD1.n159 VDD1.n126 0.155672
R946 VDD1.n166 VDD1.n126 0.155672
R947 VDD1.n167 VDD1.n166 0.155672
R948 VDD1.n167 VDD1.n122 0.155672
R949 VDD1.n174 VDD1.n122 0.155672
R950 VDD1.n175 VDD1.n174 0.155672
R951 VDD1.n175 VDD1.n118 0.155672
R952 VDD1.n183 VDD1.n118 0.155672
R953 VDD1.n184 VDD1.n183 0.155672
R954 VDD1.n184 VDD1.n114 0.155672
R955 VDD1.n192 VDD1.n114 0.155672
R956 VDD1.n193 VDD1.n192 0.155672
R957 VDD1.n193 VDD1.n110 0.155672
R958 VDD1.n200 VDD1.n110 0.155672
R959 VDD1.n201 VDD1.n200 0.155672
R960 VDD1.n201 VDD1.n106 0.155672
R961 VDD1.n208 VDD1.n106 0.155672
R962 VN VN.t0 219.066
R963 VN VN.t1 167.143
R964 VDD2.n205 VDD2.n105 756.745
R965 VDD2.n100 VDD2.n0 756.745
R966 VDD2.n206 VDD2.n205 585
R967 VDD2.n204 VDD2.n203 585
R968 VDD2.n109 VDD2.n108 585
R969 VDD2.n198 VDD2.n197 585
R970 VDD2.n196 VDD2.n195 585
R971 VDD2.n113 VDD2.n112 585
R972 VDD2.n190 VDD2.n189 585
R973 VDD2.n188 VDD2.n187 585
R974 VDD2.n186 VDD2.n116 585
R975 VDD2.n120 VDD2.n117 585
R976 VDD2.n181 VDD2.n180 585
R977 VDD2.n179 VDD2.n178 585
R978 VDD2.n122 VDD2.n121 585
R979 VDD2.n173 VDD2.n172 585
R980 VDD2.n171 VDD2.n170 585
R981 VDD2.n126 VDD2.n125 585
R982 VDD2.n165 VDD2.n164 585
R983 VDD2.n163 VDD2.n162 585
R984 VDD2.n130 VDD2.n129 585
R985 VDD2.n157 VDD2.n156 585
R986 VDD2.n155 VDD2.n154 585
R987 VDD2.n134 VDD2.n133 585
R988 VDD2.n149 VDD2.n148 585
R989 VDD2.n147 VDD2.n146 585
R990 VDD2.n138 VDD2.n137 585
R991 VDD2.n141 VDD2.n140 585
R992 VDD2.n35 VDD2.n34 585
R993 VDD2.n32 VDD2.n31 585
R994 VDD2.n41 VDD2.n40 585
R995 VDD2.n43 VDD2.n42 585
R996 VDD2.n28 VDD2.n27 585
R997 VDD2.n49 VDD2.n48 585
R998 VDD2.n51 VDD2.n50 585
R999 VDD2.n24 VDD2.n23 585
R1000 VDD2.n57 VDD2.n56 585
R1001 VDD2.n59 VDD2.n58 585
R1002 VDD2.n20 VDD2.n19 585
R1003 VDD2.n65 VDD2.n64 585
R1004 VDD2.n67 VDD2.n66 585
R1005 VDD2.n16 VDD2.n15 585
R1006 VDD2.n73 VDD2.n72 585
R1007 VDD2.n76 VDD2.n75 585
R1008 VDD2.n74 VDD2.n12 585
R1009 VDD2.n81 VDD2.n11 585
R1010 VDD2.n83 VDD2.n82 585
R1011 VDD2.n85 VDD2.n84 585
R1012 VDD2.n8 VDD2.n7 585
R1013 VDD2.n91 VDD2.n90 585
R1014 VDD2.n93 VDD2.n92 585
R1015 VDD2.n4 VDD2.n3 585
R1016 VDD2.n99 VDD2.n98 585
R1017 VDD2.n101 VDD2.n100 585
R1018 VDD2.t1 VDD2.n139 327.466
R1019 VDD2.t0 VDD2.n33 327.466
R1020 VDD2.n205 VDD2.n204 171.744
R1021 VDD2.n204 VDD2.n108 171.744
R1022 VDD2.n197 VDD2.n108 171.744
R1023 VDD2.n197 VDD2.n196 171.744
R1024 VDD2.n196 VDD2.n112 171.744
R1025 VDD2.n189 VDD2.n112 171.744
R1026 VDD2.n189 VDD2.n188 171.744
R1027 VDD2.n188 VDD2.n116 171.744
R1028 VDD2.n120 VDD2.n116 171.744
R1029 VDD2.n180 VDD2.n120 171.744
R1030 VDD2.n180 VDD2.n179 171.744
R1031 VDD2.n179 VDD2.n121 171.744
R1032 VDD2.n172 VDD2.n121 171.744
R1033 VDD2.n172 VDD2.n171 171.744
R1034 VDD2.n171 VDD2.n125 171.744
R1035 VDD2.n164 VDD2.n125 171.744
R1036 VDD2.n164 VDD2.n163 171.744
R1037 VDD2.n163 VDD2.n129 171.744
R1038 VDD2.n156 VDD2.n129 171.744
R1039 VDD2.n156 VDD2.n155 171.744
R1040 VDD2.n155 VDD2.n133 171.744
R1041 VDD2.n148 VDD2.n133 171.744
R1042 VDD2.n148 VDD2.n147 171.744
R1043 VDD2.n147 VDD2.n137 171.744
R1044 VDD2.n140 VDD2.n137 171.744
R1045 VDD2.n34 VDD2.n31 171.744
R1046 VDD2.n41 VDD2.n31 171.744
R1047 VDD2.n42 VDD2.n41 171.744
R1048 VDD2.n42 VDD2.n27 171.744
R1049 VDD2.n49 VDD2.n27 171.744
R1050 VDD2.n50 VDD2.n49 171.744
R1051 VDD2.n50 VDD2.n23 171.744
R1052 VDD2.n57 VDD2.n23 171.744
R1053 VDD2.n58 VDD2.n57 171.744
R1054 VDD2.n58 VDD2.n19 171.744
R1055 VDD2.n65 VDD2.n19 171.744
R1056 VDD2.n66 VDD2.n65 171.744
R1057 VDD2.n66 VDD2.n15 171.744
R1058 VDD2.n73 VDD2.n15 171.744
R1059 VDD2.n75 VDD2.n73 171.744
R1060 VDD2.n75 VDD2.n74 171.744
R1061 VDD2.n74 VDD2.n11 171.744
R1062 VDD2.n83 VDD2.n11 171.744
R1063 VDD2.n84 VDD2.n83 171.744
R1064 VDD2.n84 VDD2.n7 171.744
R1065 VDD2.n91 VDD2.n7 171.744
R1066 VDD2.n92 VDD2.n91 171.744
R1067 VDD2.n92 VDD2.n3 171.744
R1068 VDD2.n99 VDD2.n3 171.744
R1069 VDD2.n100 VDD2.n99 171.744
R1070 VDD2.n210 VDD2.n104 96.0149
R1071 VDD2.n140 VDD2.t1 85.8723
R1072 VDD2.n34 VDD2.t0 85.8723
R1073 VDD2.n210 VDD2.n209 49.252
R1074 VDD2.n141 VDD2.n139 16.3895
R1075 VDD2.n35 VDD2.n33 16.3895
R1076 VDD2.n187 VDD2.n186 13.1884
R1077 VDD2.n82 VDD2.n81 13.1884
R1078 VDD2.n190 VDD2.n115 12.8005
R1079 VDD2.n185 VDD2.n117 12.8005
R1080 VDD2.n142 VDD2.n138 12.8005
R1081 VDD2.n36 VDD2.n32 12.8005
R1082 VDD2.n80 VDD2.n12 12.8005
R1083 VDD2.n85 VDD2.n10 12.8005
R1084 VDD2.n191 VDD2.n113 12.0247
R1085 VDD2.n182 VDD2.n181 12.0247
R1086 VDD2.n146 VDD2.n145 12.0247
R1087 VDD2.n40 VDD2.n39 12.0247
R1088 VDD2.n77 VDD2.n76 12.0247
R1089 VDD2.n86 VDD2.n8 12.0247
R1090 VDD2.n195 VDD2.n194 11.249
R1091 VDD2.n178 VDD2.n119 11.249
R1092 VDD2.n149 VDD2.n136 11.249
R1093 VDD2.n43 VDD2.n30 11.249
R1094 VDD2.n72 VDD2.n14 11.249
R1095 VDD2.n90 VDD2.n89 11.249
R1096 VDD2.n198 VDD2.n111 10.4732
R1097 VDD2.n177 VDD2.n122 10.4732
R1098 VDD2.n150 VDD2.n134 10.4732
R1099 VDD2.n44 VDD2.n28 10.4732
R1100 VDD2.n71 VDD2.n16 10.4732
R1101 VDD2.n93 VDD2.n6 10.4732
R1102 VDD2.n199 VDD2.n109 9.69747
R1103 VDD2.n174 VDD2.n173 9.69747
R1104 VDD2.n154 VDD2.n153 9.69747
R1105 VDD2.n48 VDD2.n47 9.69747
R1106 VDD2.n68 VDD2.n67 9.69747
R1107 VDD2.n94 VDD2.n4 9.69747
R1108 VDD2.n209 VDD2.n208 9.45567
R1109 VDD2.n104 VDD2.n103 9.45567
R1110 VDD2.n167 VDD2.n166 9.3005
R1111 VDD2.n169 VDD2.n168 9.3005
R1112 VDD2.n124 VDD2.n123 9.3005
R1113 VDD2.n175 VDD2.n174 9.3005
R1114 VDD2.n177 VDD2.n176 9.3005
R1115 VDD2.n119 VDD2.n118 9.3005
R1116 VDD2.n183 VDD2.n182 9.3005
R1117 VDD2.n185 VDD2.n184 9.3005
R1118 VDD2.n208 VDD2.n207 9.3005
R1119 VDD2.n107 VDD2.n106 9.3005
R1120 VDD2.n202 VDD2.n201 9.3005
R1121 VDD2.n200 VDD2.n199 9.3005
R1122 VDD2.n111 VDD2.n110 9.3005
R1123 VDD2.n194 VDD2.n193 9.3005
R1124 VDD2.n192 VDD2.n191 9.3005
R1125 VDD2.n115 VDD2.n114 9.3005
R1126 VDD2.n128 VDD2.n127 9.3005
R1127 VDD2.n161 VDD2.n160 9.3005
R1128 VDD2.n159 VDD2.n158 9.3005
R1129 VDD2.n132 VDD2.n131 9.3005
R1130 VDD2.n153 VDD2.n152 9.3005
R1131 VDD2.n151 VDD2.n150 9.3005
R1132 VDD2.n136 VDD2.n135 9.3005
R1133 VDD2.n145 VDD2.n144 9.3005
R1134 VDD2.n143 VDD2.n142 9.3005
R1135 VDD2.n2 VDD2.n1 9.3005
R1136 VDD2.n97 VDD2.n96 9.3005
R1137 VDD2.n95 VDD2.n94 9.3005
R1138 VDD2.n6 VDD2.n5 9.3005
R1139 VDD2.n89 VDD2.n88 9.3005
R1140 VDD2.n87 VDD2.n86 9.3005
R1141 VDD2.n10 VDD2.n9 9.3005
R1142 VDD2.n55 VDD2.n54 9.3005
R1143 VDD2.n53 VDD2.n52 9.3005
R1144 VDD2.n26 VDD2.n25 9.3005
R1145 VDD2.n47 VDD2.n46 9.3005
R1146 VDD2.n45 VDD2.n44 9.3005
R1147 VDD2.n30 VDD2.n29 9.3005
R1148 VDD2.n39 VDD2.n38 9.3005
R1149 VDD2.n37 VDD2.n36 9.3005
R1150 VDD2.n22 VDD2.n21 9.3005
R1151 VDD2.n61 VDD2.n60 9.3005
R1152 VDD2.n63 VDD2.n62 9.3005
R1153 VDD2.n18 VDD2.n17 9.3005
R1154 VDD2.n69 VDD2.n68 9.3005
R1155 VDD2.n71 VDD2.n70 9.3005
R1156 VDD2.n14 VDD2.n13 9.3005
R1157 VDD2.n78 VDD2.n77 9.3005
R1158 VDD2.n80 VDD2.n79 9.3005
R1159 VDD2.n103 VDD2.n102 9.3005
R1160 VDD2.n203 VDD2.n202 8.92171
R1161 VDD2.n170 VDD2.n124 8.92171
R1162 VDD2.n157 VDD2.n132 8.92171
R1163 VDD2.n51 VDD2.n26 8.92171
R1164 VDD2.n64 VDD2.n18 8.92171
R1165 VDD2.n98 VDD2.n97 8.92171
R1166 VDD2.n206 VDD2.n107 8.14595
R1167 VDD2.n169 VDD2.n126 8.14595
R1168 VDD2.n158 VDD2.n130 8.14595
R1169 VDD2.n52 VDD2.n24 8.14595
R1170 VDD2.n63 VDD2.n20 8.14595
R1171 VDD2.n101 VDD2.n2 8.14595
R1172 VDD2.n207 VDD2.n105 7.3702
R1173 VDD2.n166 VDD2.n165 7.3702
R1174 VDD2.n162 VDD2.n161 7.3702
R1175 VDD2.n56 VDD2.n55 7.3702
R1176 VDD2.n60 VDD2.n59 7.3702
R1177 VDD2.n102 VDD2.n0 7.3702
R1178 VDD2.n209 VDD2.n105 6.59444
R1179 VDD2.n165 VDD2.n128 6.59444
R1180 VDD2.n162 VDD2.n128 6.59444
R1181 VDD2.n56 VDD2.n22 6.59444
R1182 VDD2.n59 VDD2.n22 6.59444
R1183 VDD2.n104 VDD2.n0 6.59444
R1184 VDD2.n207 VDD2.n206 5.81868
R1185 VDD2.n166 VDD2.n126 5.81868
R1186 VDD2.n161 VDD2.n130 5.81868
R1187 VDD2.n55 VDD2.n24 5.81868
R1188 VDD2.n60 VDD2.n20 5.81868
R1189 VDD2.n102 VDD2.n101 5.81868
R1190 VDD2.n203 VDD2.n107 5.04292
R1191 VDD2.n170 VDD2.n169 5.04292
R1192 VDD2.n158 VDD2.n157 5.04292
R1193 VDD2.n52 VDD2.n51 5.04292
R1194 VDD2.n64 VDD2.n63 5.04292
R1195 VDD2.n98 VDD2.n2 5.04292
R1196 VDD2.n202 VDD2.n109 4.26717
R1197 VDD2.n173 VDD2.n124 4.26717
R1198 VDD2.n154 VDD2.n132 4.26717
R1199 VDD2.n48 VDD2.n26 4.26717
R1200 VDD2.n67 VDD2.n18 4.26717
R1201 VDD2.n97 VDD2.n4 4.26717
R1202 VDD2.n143 VDD2.n139 3.70982
R1203 VDD2.n37 VDD2.n33 3.70982
R1204 VDD2.n199 VDD2.n198 3.49141
R1205 VDD2.n174 VDD2.n122 3.49141
R1206 VDD2.n153 VDD2.n134 3.49141
R1207 VDD2.n47 VDD2.n28 3.49141
R1208 VDD2.n68 VDD2.n16 3.49141
R1209 VDD2.n94 VDD2.n93 3.49141
R1210 VDD2.n195 VDD2.n111 2.71565
R1211 VDD2.n178 VDD2.n177 2.71565
R1212 VDD2.n150 VDD2.n149 2.71565
R1213 VDD2.n44 VDD2.n43 2.71565
R1214 VDD2.n72 VDD2.n71 2.71565
R1215 VDD2.n90 VDD2.n6 2.71565
R1216 VDD2.n194 VDD2.n113 1.93989
R1217 VDD2.n181 VDD2.n119 1.93989
R1218 VDD2.n146 VDD2.n136 1.93989
R1219 VDD2.n40 VDD2.n30 1.93989
R1220 VDD2.n76 VDD2.n14 1.93989
R1221 VDD2.n89 VDD2.n8 1.93989
R1222 VDD2.n191 VDD2.n190 1.16414
R1223 VDD2.n182 VDD2.n117 1.16414
R1224 VDD2.n145 VDD2.n138 1.16414
R1225 VDD2.n39 VDD2.n32 1.16414
R1226 VDD2.n77 VDD2.n12 1.16414
R1227 VDD2.n86 VDD2.n85 1.16414
R1228 VDD2 VDD2.n210 0.901362
R1229 VDD2.n187 VDD2.n115 0.388379
R1230 VDD2.n186 VDD2.n185 0.388379
R1231 VDD2.n142 VDD2.n141 0.388379
R1232 VDD2.n36 VDD2.n35 0.388379
R1233 VDD2.n81 VDD2.n80 0.388379
R1234 VDD2.n82 VDD2.n10 0.388379
R1235 VDD2.n208 VDD2.n106 0.155672
R1236 VDD2.n201 VDD2.n106 0.155672
R1237 VDD2.n201 VDD2.n200 0.155672
R1238 VDD2.n200 VDD2.n110 0.155672
R1239 VDD2.n193 VDD2.n110 0.155672
R1240 VDD2.n193 VDD2.n192 0.155672
R1241 VDD2.n192 VDD2.n114 0.155672
R1242 VDD2.n184 VDD2.n114 0.155672
R1243 VDD2.n184 VDD2.n183 0.155672
R1244 VDD2.n183 VDD2.n118 0.155672
R1245 VDD2.n176 VDD2.n118 0.155672
R1246 VDD2.n176 VDD2.n175 0.155672
R1247 VDD2.n175 VDD2.n123 0.155672
R1248 VDD2.n168 VDD2.n123 0.155672
R1249 VDD2.n168 VDD2.n167 0.155672
R1250 VDD2.n167 VDD2.n127 0.155672
R1251 VDD2.n160 VDD2.n127 0.155672
R1252 VDD2.n160 VDD2.n159 0.155672
R1253 VDD2.n159 VDD2.n131 0.155672
R1254 VDD2.n152 VDD2.n131 0.155672
R1255 VDD2.n152 VDD2.n151 0.155672
R1256 VDD2.n151 VDD2.n135 0.155672
R1257 VDD2.n144 VDD2.n135 0.155672
R1258 VDD2.n144 VDD2.n143 0.155672
R1259 VDD2.n38 VDD2.n37 0.155672
R1260 VDD2.n38 VDD2.n29 0.155672
R1261 VDD2.n45 VDD2.n29 0.155672
R1262 VDD2.n46 VDD2.n45 0.155672
R1263 VDD2.n46 VDD2.n25 0.155672
R1264 VDD2.n53 VDD2.n25 0.155672
R1265 VDD2.n54 VDD2.n53 0.155672
R1266 VDD2.n54 VDD2.n21 0.155672
R1267 VDD2.n61 VDD2.n21 0.155672
R1268 VDD2.n62 VDD2.n61 0.155672
R1269 VDD2.n62 VDD2.n17 0.155672
R1270 VDD2.n69 VDD2.n17 0.155672
R1271 VDD2.n70 VDD2.n69 0.155672
R1272 VDD2.n70 VDD2.n13 0.155672
R1273 VDD2.n78 VDD2.n13 0.155672
R1274 VDD2.n79 VDD2.n78 0.155672
R1275 VDD2.n79 VDD2.n9 0.155672
R1276 VDD2.n87 VDD2.n9 0.155672
R1277 VDD2.n88 VDD2.n87 0.155672
R1278 VDD2.n88 VDD2.n5 0.155672
R1279 VDD2.n95 VDD2.n5 0.155672
R1280 VDD2.n96 VDD2.n95 0.155672
R1281 VDD2.n96 VDD2.n1 0.155672
R1282 VDD2.n103 VDD2.n1 0.155672
R1283 B.n550 B.n89 585
R1284 B.n552 B.n551 585
R1285 B.n553 B.n88 585
R1286 B.n555 B.n554 585
R1287 B.n556 B.n87 585
R1288 B.n558 B.n557 585
R1289 B.n559 B.n86 585
R1290 B.n561 B.n560 585
R1291 B.n562 B.n85 585
R1292 B.n564 B.n563 585
R1293 B.n565 B.n84 585
R1294 B.n567 B.n566 585
R1295 B.n568 B.n83 585
R1296 B.n570 B.n569 585
R1297 B.n571 B.n82 585
R1298 B.n573 B.n572 585
R1299 B.n574 B.n81 585
R1300 B.n576 B.n575 585
R1301 B.n577 B.n80 585
R1302 B.n579 B.n578 585
R1303 B.n580 B.n79 585
R1304 B.n582 B.n581 585
R1305 B.n583 B.n78 585
R1306 B.n585 B.n584 585
R1307 B.n586 B.n77 585
R1308 B.n588 B.n587 585
R1309 B.n589 B.n76 585
R1310 B.n591 B.n590 585
R1311 B.n592 B.n75 585
R1312 B.n594 B.n593 585
R1313 B.n595 B.n74 585
R1314 B.n597 B.n596 585
R1315 B.n598 B.n73 585
R1316 B.n600 B.n599 585
R1317 B.n601 B.n72 585
R1318 B.n603 B.n602 585
R1319 B.n604 B.n71 585
R1320 B.n606 B.n605 585
R1321 B.n607 B.n70 585
R1322 B.n609 B.n608 585
R1323 B.n610 B.n69 585
R1324 B.n612 B.n611 585
R1325 B.n613 B.n68 585
R1326 B.n615 B.n614 585
R1327 B.n616 B.n67 585
R1328 B.n618 B.n617 585
R1329 B.n619 B.n66 585
R1330 B.n621 B.n620 585
R1331 B.n622 B.n65 585
R1332 B.n624 B.n623 585
R1333 B.n625 B.n64 585
R1334 B.n627 B.n626 585
R1335 B.n628 B.n63 585
R1336 B.n630 B.n629 585
R1337 B.n631 B.n62 585
R1338 B.n633 B.n632 585
R1339 B.n634 B.n61 585
R1340 B.n636 B.n635 585
R1341 B.n637 B.n60 585
R1342 B.n639 B.n638 585
R1343 B.n640 B.n59 585
R1344 B.n642 B.n641 585
R1345 B.n644 B.n56 585
R1346 B.n646 B.n645 585
R1347 B.n647 B.n55 585
R1348 B.n649 B.n648 585
R1349 B.n650 B.n54 585
R1350 B.n652 B.n651 585
R1351 B.n653 B.n53 585
R1352 B.n655 B.n654 585
R1353 B.n656 B.n49 585
R1354 B.n658 B.n657 585
R1355 B.n659 B.n48 585
R1356 B.n661 B.n660 585
R1357 B.n662 B.n47 585
R1358 B.n664 B.n663 585
R1359 B.n665 B.n46 585
R1360 B.n667 B.n666 585
R1361 B.n668 B.n45 585
R1362 B.n670 B.n669 585
R1363 B.n671 B.n44 585
R1364 B.n673 B.n672 585
R1365 B.n674 B.n43 585
R1366 B.n676 B.n675 585
R1367 B.n677 B.n42 585
R1368 B.n679 B.n678 585
R1369 B.n680 B.n41 585
R1370 B.n682 B.n681 585
R1371 B.n683 B.n40 585
R1372 B.n685 B.n684 585
R1373 B.n686 B.n39 585
R1374 B.n688 B.n687 585
R1375 B.n689 B.n38 585
R1376 B.n691 B.n690 585
R1377 B.n692 B.n37 585
R1378 B.n694 B.n693 585
R1379 B.n695 B.n36 585
R1380 B.n697 B.n696 585
R1381 B.n698 B.n35 585
R1382 B.n700 B.n699 585
R1383 B.n701 B.n34 585
R1384 B.n703 B.n702 585
R1385 B.n704 B.n33 585
R1386 B.n706 B.n705 585
R1387 B.n707 B.n32 585
R1388 B.n709 B.n708 585
R1389 B.n710 B.n31 585
R1390 B.n712 B.n711 585
R1391 B.n713 B.n30 585
R1392 B.n715 B.n714 585
R1393 B.n716 B.n29 585
R1394 B.n718 B.n717 585
R1395 B.n719 B.n28 585
R1396 B.n721 B.n720 585
R1397 B.n722 B.n27 585
R1398 B.n724 B.n723 585
R1399 B.n725 B.n26 585
R1400 B.n727 B.n726 585
R1401 B.n728 B.n25 585
R1402 B.n730 B.n729 585
R1403 B.n731 B.n24 585
R1404 B.n733 B.n732 585
R1405 B.n734 B.n23 585
R1406 B.n736 B.n735 585
R1407 B.n737 B.n22 585
R1408 B.n739 B.n738 585
R1409 B.n740 B.n21 585
R1410 B.n742 B.n741 585
R1411 B.n743 B.n20 585
R1412 B.n745 B.n744 585
R1413 B.n746 B.n19 585
R1414 B.n748 B.n747 585
R1415 B.n749 B.n18 585
R1416 B.n751 B.n750 585
R1417 B.n549 B.n548 585
R1418 B.n547 B.n90 585
R1419 B.n546 B.n545 585
R1420 B.n544 B.n91 585
R1421 B.n543 B.n542 585
R1422 B.n541 B.n92 585
R1423 B.n540 B.n539 585
R1424 B.n538 B.n93 585
R1425 B.n537 B.n536 585
R1426 B.n535 B.n94 585
R1427 B.n534 B.n533 585
R1428 B.n532 B.n95 585
R1429 B.n531 B.n530 585
R1430 B.n529 B.n96 585
R1431 B.n528 B.n527 585
R1432 B.n526 B.n97 585
R1433 B.n525 B.n524 585
R1434 B.n523 B.n98 585
R1435 B.n522 B.n521 585
R1436 B.n520 B.n99 585
R1437 B.n519 B.n518 585
R1438 B.n517 B.n100 585
R1439 B.n516 B.n515 585
R1440 B.n514 B.n101 585
R1441 B.n513 B.n512 585
R1442 B.n511 B.n102 585
R1443 B.n510 B.n509 585
R1444 B.n508 B.n103 585
R1445 B.n507 B.n506 585
R1446 B.n505 B.n104 585
R1447 B.n504 B.n503 585
R1448 B.n502 B.n105 585
R1449 B.n501 B.n500 585
R1450 B.n499 B.n106 585
R1451 B.n498 B.n497 585
R1452 B.n496 B.n107 585
R1453 B.n495 B.n494 585
R1454 B.n493 B.n108 585
R1455 B.n492 B.n491 585
R1456 B.n490 B.n109 585
R1457 B.n489 B.n488 585
R1458 B.n487 B.n110 585
R1459 B.n486 B.n485 585
R1460 B.n484 B.n111 585
R1461 B.n483 B.n482 585
R1462 B.n481 B.n112 585
R1463 B.n480 B.n479 585
R1464 B.n478 B.n113 585
R1465 B.n477 B.n476 585
R1466 B.n475 B.n114 585
R1467 B.n474 B.n473 585
R1468 B.n472 B.n115 585
R1469 B.n471 B.n470 585
R1470 B.n469 B.n116 585
R1471 B.n468 B.n467 585
R1472 B.n466 B.n117 585
R1473 B.n465 B.n464 585
R1474 B.n463 B.n118 585
R1475 B.n462 B.n461 585
R1476 B.n460 B.n119 585
R1477 B.n459 B.n458 585
R1478 B.n457 B.n120 585
R1479 B.n456 B.n455 585
R1480 B.n253 B.n192 585
R1481 B.n255 B.n254 585
R1482 B.n256 B.n191 585
R1483 B.n258 B.n257 585
R1484 B.n259 B.n190 585
R1485 B.n261 B.n260 585
R1486 B.n262 B.n189 585
R1487 B.n264 B.n263 585
R1488 B.n265 B.n188 585
R1489 B.n267 B.n266 585
R1490 B.n268 B.n187 585
R1491 B.n270 B.n269 585
R1492 B.n271 B.n186 585
R1493 B.n273 B.n272 585
R1494 B.n274 B.n185 585
R1495 B.n276 B.n275 585
R1496 B.n277 B.n184 585
R1497 B.n279 B.n278 585
R1498 B.n280 B.n183 585
R1499 B.n282 B.n281 585
R1500 B.n283 B.n182 585
R1501 B.n285 B.n284 585
R1502 B.n286 B.n181 585
R1503 B.n288 B.n287 585
R1504 B.n289 B.n180 585
R1505 B.n291 B.n290 585
R1506 B.n292 B.n179 585
R1507 B.n294 B.n293 585
R1508 B.n295 B.n178 585
R1509 B.n297 B.n296 585
R1510 B.n298 B.n177 585
R1511 B.n300 B.n299 585
R1512 B.n301 B.n176 585
R1513 B.n303 B.n302 585
R1514 B.n304 B.n175 585
R1515 B.n306 B.n305 585
R1516 B.n307 B.n174 585
R1517 B.n309 B.n308 585
R1518 B.n310 B.n173 585
R1519 B.n312 B.n311 585
R1520 B.n313 B.n172 585
R1521 B.n315 B.n314 585
R1522 B.n316 B.n171 585
R1523 B.n318 B.n317 585
R1524 B.n319 B.n170 585
R1525 B.n321 B.n320 585
R1526 B.n322 B.n169 585
R1527 B.n324 B.n323 585
R1528 B.n325 B.n168 585
R1529 B.n327 B.n326 585
R1530 B.n328 B.n167 585
R1531 B.n330 B.n329 585
R1532 B.n331 B.n166 585
R1533 B.n333 B.n332 585
R1534 B.n334 B.n165 585
R1535 B.n336 B.n335 585
R1536 B.n337 B.n164 585
R1537 B.n339 B.n338 585
R1538 B.n340 B.n163 585
R1539 B.n342 B.n341 585
R1540 B.n343 B.n162 585
R1541 B.n345 B.n344 585
R1542 B.n347 B.n346 585
R1543 B.n348 B.n158 585
R1544 B.n350 B.n349 585
R1545 B.n351 B.n157 585
R1546 B.n353 B.n352 585
R1547 B.n354 B.n156 585
R1548 B.n356 B.n355 585
R1549 B.n357 B.n155 585
R1550 B.n359 B.n358 585
R1551 B.n360 B.n152 585
R1552 B.n363 B.n362 585
R1553 B.n364 B.n151 585
R1554 B.n366 B.n365 585
R1555 B.n367 B.n150 585
R1556 B.n369 B.n368 585
R1557 B.n370 B.n149 585
R1558 B.n372 B.n371 585
R1559 B.n373 B.n148 585
R1560 B.n375 B.n374 585
R1561 B.n376 B.n147 585
R1562 B.n378 B.n377 585
R1563 B.n379 B.n146 585
R1564 B.n381 B.n380 585
R1565 B.n382 B.n145 585
R1566 B.n384 B.n383 585
R1567 B.n385 B.n144 585
R1568 B.n387 B.n386 585
R1569 B.n388 B.n143 585
R1570 B.n390 B.n389 585
R1571 B.n391 B.n142 585
R1572 B.n393 B.n392 585
R1573 B.n394 B.n141 585
R1574 B.n396 B.n395 585
R1575 B.n397 B.n140 585
R1576 B.n399 B.n398 585
R1577 B.n400 B.n139 585
R1578 B.n402 B.n401 585
R1579 B.n403 B.n138 585
R1580 B.n405 B.n404 585
R1581 B.n406 B.n137 585
R1582 B.n408 B.n407 585
R1583 B.n409 B.n136 585
R1584 B.n411 B.n410 585
R1585 B.n412 B.n135 585
R1586 B.n414 B.n413 585
R1587 B.n415 B.n134 585
R1588 B.n417 B.n416 585
R1589 B.n418 B.n133 585
R1590 B.n420 B.n419 585
R1591 B.n421 B.n132 585
R1592 B.n423 B.n422 585
R1593 B.n424 B.n131 585
R1594 B.n426 B.n425 585
R1595 B.n427 B.n130 585
R1596 B.n429 B.n428 585
R1597 B.n430 B.n129 585
R1598 B.n432 B.n431 585
R1599 B.n433 B.n128 585
R1600 B.n435 B.n434 585
R1601 B.n436 B.n127 585
R1602 B.n438 B.n437 585
R1603 B.n439 B.n126 585
R1604 B.n441 B.n440 585
R1605 B.n442 B.n125 585
R1606 B.n444 B.n443 585
R1607 B.n445 B.n124 585
R1608 B.n447 B.n446 585
R1609 B.n448 B.n123 585
R1610 B.n450 B.n449 585
R1611 B.n451 B.n122 585
R1612 B.n453 B.n452 585
R1613 B.n454 B.n121 585
R1614 B.n252 B.n251 585
R1615 B.n250 B.n193 585
R1616 B.n249 B.n248 585
R1617 B.n247 B.n194 585
R1618 B.n246 B.n245 585
R1619 B.n244 B.n195 585
R1620 B.n243 B.n242 585
R1621 B.n241 B.n196 585
R1622 B.n240 B.n239 585
R1623 B.n238 B.n197 585
R1624 B.n237 B.n236 585
R1625 B.n235 B.n198 585
R1626 B.n234 B.n233 585
R1627 B.n232 B.n199 585
R1628 B.n231 B.n230 585
R1629 B.n229 B.n200 585
R1630 B.n228 B.n227 585
R1631 B.n226 B.n201 585
R1632 B.n225 B.n224 585
R1633 B.n223 B.n202 585
R1634 B.n222 B.n221 585
R1635 B.n220 B.n203 585
R1636 B.n219 B.n218 585
R1637 B.n217 B.n204 585
R1638 B.n216 B.n215 585
R1639 B.n214 B.n205 585
R1640 B.n213 B.n212 585
R1641 B.n211 B.n206 585
R1642 B.n210 B.n209 585
R1643 B.n208 B.n207 585
R1644 B.n2 B.n0 585
R1645 B.n797 B.n1 585
R1646 B.n796 B.n795 585
R1647 B.n794 B.n3 585
R1648 B.n793 B.n792 585
R1649 B.n791 B.n4 585
R1650 B.n790 B.n789 585
R1651 B.n788 B.n5 585
R1652 B.n787 B.n786 585
R1653 B.n785 B.n6 585
R1654 B.n784 B.n783 585
R1655 B.n782 B.n7 585
R1656 B.n781 B.n780 585
R1657 B.n779 B.n8 585
R1658 B.n778 B.n777 585
R1659 B.n776 B.n9 585
R1660 B.n775 B.n774 585
R1661 B.n773 B.n10 585
R1662 B.n772 B.n771 585
R1663 B.n770 B.n11 585
R1664 B.n769 B.n768 585
R1665 B.n767 B.n12 585
R1666 B.n766 B.n765 585
R1667 B.n764 B.n13 585
R1668 B.n763 B.n762 585
R1669 B.n761 B.n14 585
R1670 B.n760 B.n759 585
R1671 B.n758 B.n15 585
R1672 B.n757 B.n756 585
R1673 B.n755 B.n16 585
R1674 B.n754 B.n753 585
R1675 B.n752 B.n17 585
R1676 B.n799 B.n798 585
R1677 B.n153 B.t2 577.332
R1678 B.n57 B.t7 577.332
R1679 B.n159 B.t11 577.332
R1680 B.n50 B.t4 577.332
R1681 B.n251 B.n192 506.916
R1682 B.n750 B.n17 506.916
R1683 B.n455 B.n454 506.916
R1684 B.n550 B.n549 506.916
R1685 B.n154 B.t1 501.5
R1686 B.n58 B.t8 501.5
R1687 B.n160 B.t10 501.5
R1688 B.n51 B.t5 501.5
R1689 B.n153 B.t0 336.935
R1690 B.n159 B.t9 336.935
R1691 B.n50 B.t3 336.935
R1692 B.n57 B.t6 336.935
R1693 B.n251 B.n250 163.367
R1694 B.n250 B.n249 163.367
R1695 B.n249 B.n194 163.367
R1696 B.n245 B.n194 163.367
R1697 B.n245 B.n244 163.367
R1698 B.n244 B.n243 163.367
R1699 B.n243 B.n196 163.367
R1700 B.n239 B.n196 163.367
R1701 B.n239 B.n238 163.367
R1702 B.n238 B.n237 163.367
R1703 B.n237 B.n198 163.367
R1704 B.n233 B.n198 163.367
R1705 B.n233 B.n232 163.367
R1706 B.n232 B.n231 163.367
R1707 B.n231 B.n200 163.367
R1708 B.n227 B.n200 163.367
R1709 B.n227 B.n226 163.367
R1710 B.n226 B.n225 163.367
R1711 B.n225 B.n202 163.367
R1712 B.n221 B.n202 163.367
R1713 B.n221 B.n220 163.367
R1714 B.n220 B.n219 163.367
R1715 B.n219 B.n204 163.367
R1716 B.n215 B.n204 163.367
R1717 B.n215 B.n214 163.367
R1718 B.n214 B.n213 163.367
R1719 B.n213 B.n206 163.367
R1720 B.n209 B.n206 163.367
R1721 B.n209 B.n208 163.367
R1722 B.n208 B.n2 163.367
R1723 B.n798 B.n2 163.367
R1724 B.n798 B.n797 163.367
R1725 B.n797 B.n796 163.367
R1726 B.n796 B.n3 163.367
R1727 B.n792 B.n3 163.367
R1728 B.n792 B.n791 163.367
R1729 B.n791 B.n790 163.367
R1730 B.n790 B.n5 163.367
R1731 B.n786 B.n5 163.367
R1732 B.n786 B.n785 163.367
R1733 B.n785 B.n784 163.367
R1734 B.n784 B.n7 163.367
R1735 B.n780 B.n7 163.367
R1736 B.n780 B.n779 163.367
R1737 B.n779 B.n778 163.367
R1738 B.n778 B.n9 163.367
R1739 B.n774 B.n9 163.367
R1740 B.n774 B.n773 163.367
R1741 B.n773 B.n772 163.367
R1742 B.n772 B.n11 163.367
R1743 B.n768 B.n11 163.367
R1744 B.n768 B.n767 163.367
R1745 B.n767 B.n766 163.367
R1746 B.n766 B.n13 163.367
R1747 B.n762 B.n13 163.367
R1748 B.n762 B.n761 163.367
R1749 B.n761 B.n760 163.367
R1750 B.n760 B.n15 163.367
R1751 B.n756 B.n15 163.367
R1752 B.n756 B.n755 163.367
R1753 B.n755 B.n754 163.367
R1754 B.n754 B.n17 163.367
R1755 B.n255 B.n192 163.367
R1756 B.n256 B.n255 163.367
R1757 B.n257 B.n256 163.367
R1758 B.n257 B.n190 163.367
R1759 B.n261 B.n190 163.367
R1760 B.n262 B.n261 163.367
R1761 B.n263 B.n262 163.367
R1762 B.n263 B.n188 163.367
R1763 B.n267 B.n188 163.367
R1764 B.n268 B.n267 163.367
R1765 B.n269 B.n268 163.367
R1766 B.n269 B.n186 163.367
R1767 B.n273 B.n186 163.367
R1768 B.n274 B.n273 163.367
R1769 B.n275 B.n274 163.367
R1770 B.n275 B.n184 163.367
R1771 B.n279 B.n184 163.367
R1772 B.n280 B.n279 163.367
R1773 B.n281 B.n280 163.367
R1774 B.n281 B.n182 163.367
R1775 B.n285 B.n182 163.367
R1776 B.n286 B.n285 163.367
R1777 B.n287 B.n286 163.367
R1778 B.n287 B.n180 163.367
R1779 B.n291 B.n180 163.367
R1780 B.n292 B.n291 163.367
R1781 B.n293 B.n292 163.367
R1782 B.n293 B.n178 163.367
R1783 B.n297 B.n178 163.367
R1784 B.n298 B.n297 163.367
R1785 B.n299 B.n298 163.367
R1786 B.n299 B.n176 163.367
R1787 B.n303 B.n176 163.367
R1788 B.n304 B.n303 163.367
R1789 B.n305 B.n304 163.367
R1790 B.n305 B.n174 163.367
R1791 B.n309 B.n174 163.367
R1792 B.n310 B.n309 163.367
R1793 B.n311 B.n310 163.367
R1794 B.n311 B.n172 163.367
R1795 B.n315 B.n172 163.367
R1796 B.n316 B.n315 163.367
R1797 B.n317 B.n316 163.367
R1798 B.n317 B.n170 163.367
R1799 B.n321 B.n170 163.367
R1800 B.n322 B.n321 163.367
R1801 B.n323 B.n322 163.367
R1802 B.n323 B.n168 163.367
R1803 B.n327 B.n168 163.367
R1804 B.n328 B.n327 163.367
R1805 B.n329 B.n328 163.367
R1806 B.n329 B.n166 163.367
R1807 B.n333 B.n166 163.367
R1808 B.n334 B.n333 163.367
R1809 B.n335 B.n334 163.367
R1810 B.n335 B.n164 163.367
R1811 B.n339 B.n164 163.367
R1812 B.n340 B.n339 163.367
R1813 B.n341 B.n340 163.367
R1814 B.n341 B.n162 163.367
R1815 B.n345 B.n162 163.367
R1816 B.n346 B.n345 163.367
R1817 B.n346 B.n158 163.367
R1818 B.n350 B.n158 163.367
R1819 B.n351 B.n350 163.367
R1820 B.n352 B.n351 163.367
R1821 B.n352 B.n156 163.367
R1822 B.n356 B.n156 163.367
R1823 B.n357 B.n356 163.367
R1824 B.n358 B.n357 163.367
R1825 B.n358 B.n152 163.367
R1826 B.n363 B.n152 163.367
R1827 B.n364 B.n363 163.367
R1828 B.n365 B.n364 163.367
R1829 B.n365 B.n150 163.367
R1830 B.n369 B.n150 163.367
R1831 B.n370 B.n369 163.367
R1832 B.n371 B.n370 163.367
R1833 B.n371 B.n148 163.367
R1834 B.n375 B.n148 163.367
R1835 B.n376 B.n375 163.367
R1836 B.n377 B.n376 163.367
R1837 B.n377 B.n146 163.367
R1838 B.n381 B.n146 163.367
R1839 B.n382 B.n381 163.367
R1840 B.n383 B.n382 163.367
R1841 B.n383 B.n144 163.367
R1842 B.n387 B.n144 163.367
R1843 B.n388 B.n387 163.367
R1844 B.n389 B.n388 163.367
R1845 B.n389 B.n142 163.367
R1846 B.n393 B.n142 163.367
R1847 B.n394 B.n393 163.367
R1848 B.n395 B.n394 163.367
R1849 B.n395 B.n140 163.367
R1850 B.n399 B.n140 163.367
R1851 B.n400 B.n399 163.367
R1852 B.n401 B.n400 163.367
R1853 B.n401 B.n138 163.367
R1854 B.n405 B.n138 163.367
R1855 B.n406 B.n405 163.367
R1856 B.n407 B.n406 163.367
R1857 B.n407 B.n136 163.367
R1858 B.n411 B.n136 163.367
R1859 B.n412 B.n411 163.367
R1860 B.n413 B.n412 163.367
R1861 B.n413 B.n134 163.367
R1862 B.n417 B.n134 163.367
R1863 B.n418 B.n417 163.367
R1864 B.n419 B.n418 163.367
R1865 B.n419 B.n132 163.367
R1866 B.n423 B.n132 163.367
R1867 B.n424 B.n423 163.367
R1868 B.n425 B.n424 163.367
R1869 B.n425 B.n130 163.367
R1870 B.n429 B.n130 163.367
R1871 B.n430 B.n429 163.367
R1872 B.n431 B.n430 163.367
R1873 B.n431 B.n128 163.367
R1874 B.n435 B.n128 163.367
R1875 B.n436 B.n435 163.367
R1876 B.n437 B.n436 163.367
R1877 B.n437 B.n126 163.367
R1878 B.n441 B.n126 163.367
R1879 B.n442 B.n441 163.367
R1880 B.n443 B.n442 163.367
R1881 B.n443 B.n124 163.367
R1882 B.n447 B.n124 163.367
R1883 B.n448 B.n447 163.367
R1884 B.n449 B.n448 163.367
R1885 B.n449 B.n122 163.367
R1886 B.n453 B.n122 163.367
R1887 B.n454 B.n453 163.367
R1888 B.n455 B.n120 163.367
R1889 B.n459 B.n120 163.367
R1890 B.n460 B.n459 163.367
R1891 B.n461 B.n460 163.367
R1892 B.n461 B.n118 163.367
R1893 B.n465 B.n118 163.367
R1894 B.n466 B.n465 163.367
R1895 B.n467 B.n466 163.367
R1896 B.n467 B.n116 163.367
R1897 B.n471 B.n116 163.367
R1898 B.n472 B.n471 163.367
R1899 B.n473 B.n472 163.367
R1900 B.n473 B.n114 163.367
R1901 B.n477 B.n114 163.367
R1902 B.n478 B.n477 163.367
R1903 B.n479 B.n478 163.367
R1904 B.n479 B.n112 163.367
R1905 B.n483 B.n112 163.367
R1906 B.n484 B.n483 163.367
R1907 B.n485 B.n484 163.367
R1908 B.n485 B.n110 163.367
R1909 B.n489 B.n110 163.367
R1910 B.n490 B.n489 163.367
R1911 B.n491 B.n490 163.367
R1912 B.n491 B.n108 163.367
R1913 B.n495 B.n108 163.367
R1914 B.n496 B.n495 163.367
R1915 B.n497 B.n496 163.367
R1916 B.n497 B.n106 163.367
R1917 B.n501 B.n106 163.367
R1918 B.n502 B.n501 163.367
R1919 B.n503 B.n502 163.367
R1920 B.n503 B.n104 163.367
R1921 B.n507 B.n104 163.367
R1922 B.n508 B.n507 163.367
R1923 B.n509 B.n508 163.367
R1924 B.n509 B.n102 163.367
R1925 B.n513 B.n102 163.367
R1926 B.n514 B.n513 163.367
R1927 B.n515 B.n514 163.367
R1928 B.n515 B.n100 163.367
R1929 B.n519 B.n100 163.367
R1930 B.n520 B.n519 163.367
R1931 B.n521 B.n520 163.367
R1932 B.n521 B.n98 163.367
R1933 B.n525 B.n98 163.367
R1934 B.n526 B.n525 163.367
R1935 B.n527 B.n526 163.367
R1936 B.n527 B.n96 163.367
R1937 B.n531 B.n96 163.367
R1938 B.n532 B.n531 163.367
R1939 B.n533 B.n532 163.367
R1940 B.n533 B.n94 163.367
R1941 B.n537 B.n94 163.367
R1942 B.n538 B.n537 163.367
R1943 B.n539 B.n538 163.367
R1944 B.n539 B.n92 163.367
R1945 B.n543 B.n92 163.367
R1946 B.n544 B.n543 163.367
R1947 B.n545 B.n544 163.367
R1948 B.n545 B.n90 163.367
R1949 B.n549 B.n90 163.367
R1950 B.n750 B.n749 163.367
R1951 B.n749 B.n748 163.367
R1952 B.n748 B.n19 163.367
R1953 B.n744 B.n19 163.367
R1954 B.n744 B.n743 163.367
R1955 B.n743 B.n742 163.367
R1956 B.n742 B.n21 163.367
R1957 B.n738 B.n21 163.367
R1958 B.n738 B.n737 163.367
R1959 B.n737 B.n736 163.367
R1960 B.n736 B.n23 163.367
R1961 B.n732 B.n23 163.367
R1962 B.n732 B.n731 163.367
R1963 B.n731 B.n730 163.367
R1964 B.n730 B.n25 163.367
R1965 B.n726 B.n25 163.367
R1966 B.n726 B.n725 163.367
R1967 B.n725 B.n724 163.367
R1968 B.n724 B.n27 163.367
R1969 B.n720 B.n27 163.367
R1970 B.n720 B.n719 163.367
R1971 B.n719 B.n718 163.367
R1972 B.n718 B.n29 163.367
R1973 B.n714 B.n29 163.367
R1974 B.n714 B.n713 163.367
R1975 B.n713 B.n712 163.367
R1976 B.n712 B.n31 163.367
R1977 B.n708 B.n31 163.367
R1978 B.n708 B.n707 163.367
R1979 B.n707 B.n706 163.367
R1980 B.n706 B.n33 163.367
R1981 B.n702 B.n33 163.367
R1982 B.n702 B.n701 163.367
R1983 B.n701 B.n700 163.367
R1984 B.n700 B.n35 163.367
R1985 B.n696 B.n35 163.367
R1986 B.n696 B.n695 163.367
R1987 B.n695 B.n694 163.367
R1988 B.n694 B.n37 163.367
R1989 B.n690 B.n37 163.367
R1990 B.n690 B.n689 163.367
R1991 B.n689 B.n688 163.367
R1992 B.n688 B.n39 163.367
R1993 B.n684 B.n39 163.367
R1994 B.n684 B.n683 163.367
R1995 B.n683 B.n682 163.367
R1996 B.n682 B.n41 163.367
R1997 B.n678 B.n41 163.367
R1998 B.n678 B.n677 163.367
R1999 B.n677 B.n676 163.367
R2000 B.n676 B.n43 163.367
R2001 B.n672 B.n43 163.367
R2002 B.n672 B.n671 163.367
R2003 B.n671 B.n670 163.367
R2004 B.n670 B.n45 163.367
R2005 B.n666 B.n45 163.367
R2006 B.n666 B.n665 163.367
R2007 B.n665 B.n664 163.367
R2008 B.n664 B.n47 163.367
R2009 B.n660 B.n47 163.367
R2010 B.n660 B.n659 163.367
R2011 B.n659 B.n658 163.367
R2012 B.n658 B.n49 163.367
R2013 B.n654 B.n49 163.367
R2014 B.n654 B.n653 163.367
R2015 B.n653 B.n652 163.367
R2016 B.n652 B.n54 163.367
R2017 B.n648 B.n54 163.367
R2018 B.n648 B.n647 163.367
R2019 B.n647 B.n646 163.367
R2020 B.n646 B.n56 163.367
R2021 B.n641 B.n56 163.367
R2022 B.n641 B.n640 163.367
R2023 B.n640 B.n639 163.367
R2024 B.n639 B.n60 163.367
R2025 B.n635 B.n60 163.367
R2026 B.n635 B.n634 163.367
R2027 B.n634 B.n633 163.367
R2028 B.n633 B.n62 163.367
R2029 B.n629 B.n62 163.367
R2030 B.n629 B.n628 163.367
R2031 B.n628 B.n627 163.367
R2032 B.n627 B.n64 163.367
R2033 B.n623 B.n64 163.367
R2034 B.n623 B.n622 163.367
R2035 B.n622 B.n621 163.367
R2036 B.n621 B.n66 163.367
R2037 B.n617 B.n66 163.367
R2038 B.n617 B.n616 163.367
R2039 B.n616 B.n615 163.367
R2040 B.n615 B.n68 163.367
R2041 B.n611 B.n68 163.367
R2042 B.n611 B.n610 163.367
R2043 B.n610 B.n609 163.367
R2044 B.n609 B.n70 163.367
R2045 B.n605 B.n70 163.367
R2046 B.n605 B.n604 163.367
R2047 B.n604 B.n603 163.367
R2048 B.n603 B.n72 163.367
R2049 B.n599 B.n72 163.367
R2050 B.n599 B.n598 163.367
R2051 B.n598 B.n597 163.367
R2052 B.n597 B.n74 163.367
R2053 B.n593 B.n74 163.367
R2054 B.n593 B.n592 163.367
R2055 B.n592 B.n591 163.367
R2056 B.n591 B.n76 163.367
R2057 B.n587 B.n76 163.367
R2058 B.n587 B.n586 163.367
R2059 B.n586 B.n585 163.367
R2060 B.n585 B.n78 163.367
R2061 B.n581 B.n78 163.367
R2062 B.n581 B.n580 163.367
R2063 B.n580 B.n579 163.367
R2064 B.n579 B.n80 163.367
R2065 B.n575 B.n80 163.367
R2066 B.n575 B.n574 163.367
R2067 B.n574 B.n573 163.367
R2068 B.n573 B.n82 163.367
R2069 B.n569 B.n82 163.367
R2070 B.n569 B.n568 163.367
R2071 B.n568 B.n567 163.367
R2072 B.n567 B.n84 163.367
R2073 B.n563 B.n84 163.367
R2074 B.n563 B.n562 163.367
R2075 B.n562 B.n561 163.367
R2076 B.n561 B.n86 163.367
R2077 B.n557 B.n86 163.367
R2078 B.n557 B.n556 163.367
R2079 B.n556 B.n555 163.367
R2080 B.n555 B.n88 163.367
R2081 B.n551 B.n88 163.367
R2082 B.n551 B.n550 163.367
R2083 B.n154 B.n153 75.8308
R2084 B.n160 B.n159 75.8308
R2085 B.n51 B.n50 75.8308
R2086 B.n58 B.n57 75.8308
R2087 B.n361 B.n154 59.5399
R2088 B.n161 B.n160 59.5399
R2089 B.n52 B.n51 59.5399
R2090 B.n643 B.n58 59.5399
R2091 B.n752 B.n751 32.9371
R2092 B.n548 B.n89 32.9371
R2093 B.n456 B.n121 32.9371
R2094 B.n253 B.n252 32.9371
R2095 B B.n799 18.0485
R2096 B.n751 B.n18 10.6151
R2097 B.n747 B.n18 10.6151
R2098 B.n747 B.n746 10.6151
R2099 B.n746 B.n745 10.6151
R2100 B.n745 B.n20 10.6151
R2101 B.n741 B.n20 10.6151
R2102 B.n741 B.n740 10.6151
R2103 B.n740 B.n739 10.6151
R2104 B.n739 B.n22 10.6151
R2105 B.n735 B.n22 10.6151
R2106 B.n735 B.n734 10.6151
R2107 B.n734 B.n733 10.6151
R2108 B.n733 B.n24 10.6151
R2109 B.n729 B.n24 10.6151
R2110 B.n729 B.n728 10.6151
R2111 B.n728 B.n727 10.6151
R2112 B.n727 B.n26 10.6151
R2113 B.n723 B.n26 10.6151
R2114 B.n723 B.n722 10.6151
R2115 B.n722 B.n721 10.6151
R2116 B.n721 B.n28 10.6151
R2117 B.n717 B.n28 10.6151
R2118 B.n717 B.n716 10.6151
R2119 B.n716 B.n715 10.6151
R2120 B.n715 B.n30 10.6151
R2121 B.n711 B.n30 10.6151
R2122 B.n711 B.n710 10.6151
R2123 B.n710 B.n709 10.6151
R2124 B.n709 B.n32 10.6151
R2125 B.n705 B.n32 10.6151
R2126 B.n705 B.n704 10.6151
R2127 B.n704 B.n703 10.6151
R2128 B.n703 B.n34 10.6151
R2129 B.n699 B.n34 10.6151
R2130 B.n699 B.n698 10.6151
R2131 B.n698 B.n697 10.6151
R2132 B.n697 B.n36 10.6151
R2133 B.n693 B.n36 10.6151
R2134 B.n693 B.n692 10.6151
R2135 B.n692 B.n691 10.6151
R2136 B.n691 B.n38 10.6151
R2137 B.n687 B.n38 10.6151
R2138 B.n687 B.n686 10.6151
R2139 B.n686 B.n685 10.6151
R2140 B.n685 B.n40 10.6151
R2141 B.n681 B.n40 10.6151
R2142 B.n681 B.n680 10.6151
R2143 B.n680 B.n679 10.6151
R2144 B.n679 B.n42 10.6151
R2145 B.n675 B.n42 10.6151
R2146 B.n675 B.n674 10.6151
R2147 B.n674 B.n673 10.6151
R2148 B.n673 B.n44 10.6151
R2149 B.n669 B.n44 10.6151
R2150 B.n669 B.n668 10.6151
R2151 B.n668 B.n667 10.6151
R2152 B.n667 B.n46 10.6151
R2153 B.n663 B.n46 10.6151
R2154 B.n663 B.n662 10.6151
R2155 B.n662 B.n661 10.6151
R2156 B.n661 B.n48 10.6151
R2157 B.n657 B.n656 10.6151
R2158 B.n656 B.n655 10.6151
R2159 B.n655 B.n53 10.6151
R2160 B.n651 B.n53 10.6151
R2161 B.n651 B.n650 10.6151
R2162 B.n650 B.n649 10.6151
R2163 B.n649 B.n55 10.6151
R2164 B.n645 B.n55 10.6151
R2165 B.n645 B.n644 10.6151
R2166 B.n642 B.n59 10.6151
R2167 B.n638 B.n59 10.6151
R2168 B.n638 B.n637 10.6151
R2169 B.n637 B.n636 10.6151
R2170 B.n636 B.n61 10.6151
R2171 B.n632 B.n61 10.6151
R2172 B.n632 B.n631 10.6151
R2173 B.n631 B.n630 10.6151
R2174 B.n630 B.n63 10.6151
R2175 B.n626 B.n63 10.6151
R2176 B.n626 B.n625 10.6151
R2177 B.n625 B.n624 10.6151
R2178 B.n624 B.n65 10.6151
R2179 B.n620 B.n65 10.6151
R2180 B.n620 B.n619 10.6151
R2181 B.n619 B.n618 10.6151
R2182 B.n618 B.n67 10.6151
R2183 B.n614 B.n67 10.6151
R2184 B.n614 B.n613 10.6151
R2185 B.n613 B.n612 10.6151
R2186 B.n612 B.n69 10.6151
R2187 B.n608 B.n69 10.6151
R2188 B.n608 B.n607 10.6151
R2189 B.n607 B.n606 10.6151
R2190 B.n606 B.n71 10.6151
R2191 B.n602 B.n71 10.6151
R2192 B.n602 B.n601 10.6151
R2193 B.n601 B.n600 10.6151
R2194 B.n600 B.n73 10.6151
R2195 B.n596 B.n73 10.6151
R2196 B.n596 B.n595 10.6151
R2197 B.n595 B.n594 10.6151
R2198 B.n594 B.n75 10.6151
R2199 B.n590 B.n75 10.6151
R2200 B.n590 B.n589 10.6151
R2201 B.n589 B.n588 10.6151
R2202 B.n588 B.n77 10.6151
R2203 B.n584 B.n77 10.6151
R2204 B.n584 B.n583 10.6151
R2205 B.n583 B.n582 10.6151
R2206 B.n582 B.n79 10.6151
R2207 B.n578 B.n79 10.6151
R2208 B.n578 B.n577 10.6151
R2209 B.n577 B.n576 10.6151
R2210 B.n576 B.n81 10.6151
R2211 B.n572 B.n81 10.6151
R2212 B.n572 B.n571 10.6151
R2213 B.n571 B.n570 10.6151
R2214 B.n570 B.n83 10.6151
R2215 B.n566 B.n83 10.6151
R2216 B.n566 B.n565 10.6151
R2217 B.n565 B.n564 10.6151
R2218 B.n564 B.n85 10.6151
R2219 B.n560 B.n85 10.6151
R2220 B.n560 B.n559 10.6151
R2221 B.n559 B.n558 10.6151
R2222 B.n558 B.n87 10.6151
R2223 B.n554 B.n87 10.6151
R2224 B.n554 B.n553 10.6151
R2225 B.n553 B.n552 10.6151
R2226 B.n552 B.n89 10.6151
R2227 B.n457 B.n456 10.6151
R2228 B.n458 B.n457 10.6151
R2229 B.n458 B.n119 10.6151
R2230 B.n462 B.n119 10.6151
R2231 B.n463 B.n462 10.6151
R2232 B.n464 B.n463 10.6151
R2233 B.n464 B.n117 10.6151
R2234 B.n468 B.n117 10.6151
R2235 B.n469 B.n468 10.6151
R2236 B.n470 B.n469 10.6151
R2237 B.n470 B.n115 10.6151
R2238 B.n474 B.n115 10.6151
R2239 B.n475 B.n474 10.6151
R2240 B.n476 B.n475 10.6151
R2241 B.n476 B.n113 10.6151
R2242 B.n480 B.n113 10.6151
R2243 B.n481 B.n480 10.6151
R2244 B.n482 B.n481 10.6151
R2245 B.n482 B.n111 10.6151
R2246 B.n486 B.n111 10.6151
R2247 B.n487 B.n486 10.6151
R2248 B.n488 B.n487 10.6151
R2249 B.n488 B.n109 10.6151
R2250 B.n492 B.n109 10.6151
R2251 B.n493 B.n492 10.6151
R2252 B.n494 B.n493 10.6151
R2253 B.n494 B.n107 10.6151
R2254 B.n498 B.n107 10.6151
R2255 B.n499 B.n498 10.6151
R2256 B.n500 B.n499 10.6151
R2257 B.n500 B.n105 10.6151
R2258 B.n504 B.n105 10.6151
R2259 B.n505 B.n504 10.6151
R2260 B.n506 B.n505 10.6151
R2261 B.n506 B.n103 10.6151
R2262 B.n510 B.n103 10.6151
R2263 B.n511 B.n510 10.6151
R2264 B.n512 B.n511 10.6151
R2265 B.n512 B.n101 10.6151
R2266 B.n516 B.n101 10.6151
R2267 B.n517 B.n516 10.6151
R2268 B.n518 B.n517 10.6151
R2269 B.n518 B.n99 10.6151
R2270 B.n522 B.n99 10.6151
R2271 B.n523 B.n522 10.6151
R2272 B.n524 B.n523 10.6151
R2273 B.n524 B.n97 10.6151
R2274 B.n528 B.n97 10.6151
R2275 B.n529 B.n528 10.6151
R2276 B.n530 B.n529 10.6151
R2277 B.n530 B.n95 10.6151
R2278 B.n534 B.n95 10.6151
R2279 B.n535 B.n534 10.6151
R2280 B.n536 B.n535 10.6151
R2281 B.n536 B.n93 10.6151
R2282 B.n540 B.n93 10.6151
R2283 B.n541 B.n540 10.6151
R2284 B.n542 B.n541 10.6151
R2285 B.n542 B.n91 10.6151
R2286 B.n546 B.n91 10.6151
R2287 B.n547 B.n546 10.6151
R2288 B.n548 B.n547 10.6151
R2289 B.n254 B.n253 10.6151
R2290 B.n254 B.n191 10.6151
R2291 B.n258 B.n191 10.6151
R2292 B.n259 B.n258 10.6151
R2293 B.n260 B.n259 10.6151
R2294 B.n260 B.n189 10.6151
R2295 B.n264 B.n189 10.6151
R2296 B.n265 B.n264 10.6151
R2297 B.n266 B.n265 10.6151
R2298 B.n266 B.n187 10.6151
R2299 B.n270 B.n187 10.6151
R2300 B.n271 B.n270 10.6151
R2301 B.n272 B.n271 10.6151
R2302 B.n272 B.n185 10.6151
R2303 B.n276 B.n185 10.6151
R2304 B.n277 B.n276 10.6151
R2305 B.n278 B.n277 10.6151
R2306 B.n278 B.n183 10.6151
R2307 B.n282 B.n183 10.6151
R2308 B.n283 B.n282 10.6151
R2309 B.n284 B.n283 10.6151
R2310 B.n284 B.n181 10.6151
R2311 B.n288 B.n181 10.6151
R2312 B.n289 B.n288 10.6151
R2313 B.n290 B.n289 10.6151
R2314 B.n290 B.n179 10.6151
R2315 B.n294 B.n179 10.6151
R2316 B.n295 B.n294 10.6151
R2317 B.n296 B.n295 10.6151
R2318 B.n296 B.n177 10.6151
R2319 B.n300 B.n177 10.6151
R2320 B.n301 B.n300 10.6151
R2321 B.n302 B.n301 10.6151
R2322 B.n302 B.n175 10.6151
R2323 B.n306 B.n175 10.6151
R2324 B.n307 B.n306 10.6151
R2325 B.n308 B.n307 10.6151
R2326 B.n308 B.n173 10.6151
R2327 B.n312 B.n173 10.6151
R2328 B.n313 B.n312 10.6151
R2329 B.n314 B.n313 10.6151
R2330 B.n314 B.n171 10.6151
R2331 B.n318 B.n171 10.6151
R2332 B.n319 B.n318 10.6151
R2333 B.n320 B.n319 10.6151
R2334 B.n320 B.n169 10.6151
R2335 B.n324 B.n169 10.6151
R2336 B.n325 B.n324 10.6151
R2337 B.n326 B.n325 10.6151
R2338 B.n326 B.n167 10.6151
R2339 B.n330 B.n167 10.6151
R2340 B.n331 B.n330 10.6151
R2341 B.n332 B.n331 10.6151
R2342 B.n332 B.n165 10.6151
R2343 B.n336 B.n165 10.6151
R2344 B.n337 B.n336 10.6151
R2345 B.n338 B.n337 10.6151
R2346 B.n338 B.n163 10.6151
R2347 B.n342 B.n163 10.6151
R2348 B.n343 B.n342 10.6151
R2349 B.n344 B.n343 10.6151
R2350 B.n348 B.n347 10.6151
R2351 B.n349 B.n348 10.6151
R2352 B.n349 B.n157 10.6151
R2353 B.n353 B.n157 10.6151
R2354 B.n354 B.n353 10.6151
R2355 B.n355 B.n354 10.6151
R2356 B.n355 B.n155 10.6151
R2357 B.n359 B.n155 10.6151
R2358 B.n360 B.n359 10.6151
R2359 B.n362 B.n151 10.6151
R2360 B.n366 B.n151 10.6151
R2361 B.n367 B.n366 10.6151
R2362 B.n368 B.n367 10.6151
R2363 B.n368 B.n149 10.6151
R2364 B.n372 B.n149 10.6151
R2365 B.n373 B.n372 10.6151
R2366 B.n374 B.n373 10.6151
R2367 B.n374 B.n147 10.6151
R2368 B.n378 B.n147 10.6151
R2369 B.n379 B.n378 10.6151
R2370 B.n380 B.n379 10.6151
R2371 B.n380 B.n145 10.6151
R2372 B.n384 B.n145 10.6151
R2373 B.n385 B.n384 10.6151
R2374 B.n386 B.n385 10.6151
R2375 B.n386 B.n143 10.6151
R2376 B.n390 B.n143 10.6151
R2377 B.n391 B.n390 10.6151
R2378 B.n392 B.n391 10.6151
R2379 B.n392 B.n141 10.6151
R2380 B.n396 B.n141 10.6151
R2381 B.n397 B.n396 10.6151
R2382 B.n398 B.n397 10.6151
R2383 B.n398 B.n139 10.6151
R2384 B.n402 B.n139 10.6151
R2385 B.n403 B.n402 10.6151
R2386 B.n404 B.n403 10.6151
R2387 B.n404 B.n137 10.6151
R2388 B.n408 B.n137 10.6151
R2389 B.n409 B.n408 10.6151
R2390 B.n410 B.n409 10.6151
R2391 B.n410 B.n135 10.6151
R2392 B.n414 B.n135 10.6151
R2393 B.n415 B.n414 10.6151
R2394 B.n416 B.n415 10.6151
R2395 B.n416 B.n133 10.6151
R2396 B.n420 B.n133 10.6151
R2397 B.n421 B.n420 10.6151
R2398 B.n422 B.n421 10.6151
R2399 B.n422 B.n131 10.6151
R2400 B.n426 B.n131 10.6151
R2401 B.n427 B.n426 10.6151
R2402 B.n428 B.n427 10.6151
R2403 B.n428 B.n129 10.6151
R2404 B.n432 B.n129 10.6151
R2405 B.n433 B.n432 10.6151
R2406 B.n434 B.n433 10.6151
R2407 B.n434 B.n127 10.6151
R2408 B.n438 B.n127 10.6151
R2409 B.n439 B.n438 10.6151
R2410 B.n440 B.n439 10.6151
R2411 B.n440 B.n125 10.6151
R2412 B.n444 B.n125 10.6151
R2413 B.n445 B.n444 10.6151
R2414 B.n446 B.n445 10.6151
R2415 B.n446 B.n123 10.6151
R2416 B.n450 B.n123 10.6151
R2417 B.n451 B.n450 10.6151
R2418 B.n452 B.n451 10.6151
R2419 B.n452 B.n121 10.6151
R2420 B.n252 B.n193 10.6151
R2421 B.n248 B.n193 10.6151
R2422 B.n248 B.n247 10.6151
R2423 B.n247 B.n246 10.6151
R2424 B.n246 B.n195 10.6151
R2425 B.n242 B.n195 10.6151
R2426 B.n242 B.n241 10.6151
R2427 B.n241 B.n240 10.6151
R2428 B.n240 B.n197 10.6151
R2429 B.n236 B.n197 10.6151
R2430 B.n236 B.n235 10.6151
R2431 B.n235 B.n234 10.6151
R2432 B.n234 B.n199 10.6151
R2433 B.n230 B.n199 10.6151
R2434 B.n230 B.n229 10.6151
R2435 B.n229 B.n228 10.6151
R2436 B.n228 B.n201 10.6151
R2437 B.n224 B.n201 10.6151
R2438 B.n224 B.n223 10.6151
R2439 B.n223 B.n222 10.6151
R2440 B.n222 B.n203 10.6151
R2441 B.n218 B.n203 10.6151
R2442 B.n218 B.n217 10.6151
R2443 B.n217 B.n216 10.6151
R2444 B.n216 B.n205 10.6151
R2445 B.n212 B.n205 10.6151
R2446 B.n212 B.n211 10.6151
R2447 B.n211 B.n210 10.6151
R2448 B.n210 B.n207 10.6151
R2449 B.n207 B.n0 10.6151
R2450 B.n795 B.n1 10.6151
R2451 B.n795 B.n794 10.6151
R2452 B.n794 B.n793 10.6151
R2453 B.n793 B.n4 10.6151
R2454 B.n789 B.n4 10.6151
R2455 B.n789 B.n788 10.6151
R2456 B.n788 B.n787 10.6151
R2457 B.n787 B.n6 10.6151
R2458 B.n783 B.n6 10.6151
R2459 B.n783 B.n782 10.6151
R2460 B.n782 B.n781 10.6151
R2461 B.n781 B.n8 10.6151
R2462 B.n777 B.n8 10.6151
R2463 B.n777 B.n776 10.6151
R2464 B.n776 B.n775 10.6151
R2465 B.n775 B.n10 10.6151
R2466 B.n771 B.n10 10.6151
R2467 B.n771 B.n770 10.6151
R2468 B.n770 B.n769 10.6151
R2469 B.n769 B.n12 10.6151
R2470 B.n765 B.n12 10.6151
R2471 B.n765 B.n764 10.6151
R2472 B.n764 B.n763 10.6151
R2473 B.n763 B.n14 10.6151
R2474 B.n759 B.n14 10.6151
R2475 B.n759 B.n758 10.6151
R2476 B.n758 B.n757 10.6151
R2477 B.n757 B.n16 10.6151
R2478 B.n753 B.n16 10.6151
R2479 B.n753 B.n752 10.6151
R2480 B.n52 B.n48 9.36635
R2481 B.n643 B.n642 9.36635
R2482 B.n344 B.n161 9.36635
R2483 B.n362 B.n361 9.36635
R2484 B.n799 B.n0 2.81026
R2485 B.n799 B.n1 2.81026
R2486 B.n657 B.n52 1.24928
R2487 B.n644 B.n643 1.24928
R2488 B.n347 B.n161 1.24928
R2489 B.n361 B.n360 1.24928
C0 VP VTAIL 3.85296f
C1 B VN 1.30118f
C2 VDD1 w_n2534_n4764# 2.36848f
C3 VP VN 7.20207f
C4 VN VTAIL 3.83859f
C5 VDD2 w_n2534_n4764# 2.40646f
C6 VDD1 VDD2 0.780666f
C7 B w_n2534_n4764# 11.824599f
C8 B VDD1 2.39715f
C9 VP w_n2534_n4764# 4.03794f
C10 VTAIL w_n2534_n4764# 3.71469f
C11 VP VDD1 4.664f
C12 B VDD2 2.43598f
C13 VDD1 VTAIL 7.01185f
C14 VP VDD2 0.374941f
C15 VN w_n2534_n4764# 3.71304f
C16 VDD2 VTAIL 7.0687f
C17 VDD1 VN 0.148906f
C18 VDD2 VN 4.44097f
C19 B VP 1.83925f
C20 B VTAIL 5.66991f
C21 VDD2 VSUBS 1.266783f
C22 VDD1 VSUBS 6.10145f
C23 VTAIL VSUBS 1.376629f
C24 VN VSUBS 9.43259f
C25 VP VSUBS 2.22044f
C26 B VSUBS 5.218378f
C27 w_n2534_n4764# VSUBS 0.147509p
C28 B.n0 VSUBS 0.00391f
C29 B.n1 VSUBS 0.00391f
C30 B.n2 VSUBS 0.006183f
C31 B.n3 VSUBS 0.006183f
C32 B.n4 VSUBS 0.006183f
C33 B.n5 VSUBS 0.006183f
C34 B.n6 VSUBS 0.006183f
C35 B.n7 VSUBS 0.006183f
C36 B.n8 VSUBS 0.006183f
C37 B.n9 VSUBS 0.006183f
C38 B.n10 VSUBS 0.006183f
C39 B.n11 VSUBS 0.006183f
C40 B.n12 VSUBS 0.006183f
C41 B.n13 VSUBS 0.006183f
C42 B.n14 VSUBS 0.006183f
C43 B.n15 VSUBS 0.006183f
C44 B.n16 VSUBS 0.006183f
C45 B.n17 VSUBS 0.014099f
C46 B.n18 VSUBS 0.006183f
C47 B.n19 VSUBS 0.006183f
C48 B.n20 VSUBS 0.006183f
C49 B.n21 VSUBS 0.006183f
C50 B.n22 VSUBS 0.006183f
C51 B.n23 VSUBS 0.006183f
C52 B.n24 VSUBS 0.006183f
C53 B.n25 VSUBS 0.006183f
C54 B.n26 VSUBS 0.006183f
C55 B.n27 VSUBS 0.006183f
C56 B.n28 VSUBS 0.006183f
C57 B.n29 VSUBS 0.006183f
C58 B.n30 VSUBS 0.006183f
C59 B.n31 VSUBS 0.006183f
C60 B.n32 VSUBS 0.006183f
C61 B.n33 VSUBS 0.006183f
C62 B.n34 VSUBS 0.006183f
C63 B.n35 VSUBS 0.006183f
C64 B.n36 VSUBS 0.006183f
C65 B.n37 VSUBS 0.006183f
C66 B.n38 VSUBS 0.006183f
C67 B.n39 VSUBS 0.006183f
C68 B.n40 VSUBS 0.006183f
C69 B.n41 VSUBS 0.006183f
C70 B.n42 VSUBS 0.006183f
C71 B.n43 VSUBS 0.006183f
C72 B.n44 VSUBS 0.006183f
C73 B.n45 VSUBS 0.006183f
C74 B.n46 VSUBS 0.006183f
C75 B.n47 VSUBS 0.006183f
C76 B.n48 VSUBS 0.00582f
C77 B.n49 VSUBS 0.006183f
C78 B.t5 VSUBS 0.331284f
C79 B.t4 VSUBS 0.370067f
C80 B.t3 VSUBS 2.71492f
C81 B.n50 VSUBS 0.589031f
C82 B.n51 VSUBS 0.30409f
C83 B.n52 VSUBS 0.014326f
C84 B.n53 VSUBS 0.006183f
C85 B.n54 VSUBS 0.006183f
C86 B.n55 VSUBS 0.006183f
C87 B.n56 VSUBS 0.006183f
C88 B.t8 VSUBS 0.331288f
C89 B.t7 VSUBS 0.37007f
C90 B.t6 VSUBS 2.71492f
C91 B.n57 VSUBS 0.589028f
C92 B.n58 VSUBS 0.304086f
C93 B.n59 VSUBS 0.006183f
C94 B.n60 VSUBS 0.006183f
C95 B.n61 VSUBS 0.006183f
C96 B.n62 VSUBS 0.006183f
C97 B.n63 VSUBS 0.006183f
C98 B.n64 VSUBS 0.006183f
C99 B.n65 VSUBS 0.006183f
C100 B.n66 VSUBS 0.006183f
C101 B.n67 VSUBS 0.006183f
C102 B.n68 VSUBS 0.006183f
C103 B.n69 VSUBS 0.006183f
C104 B.n70 VSUBS 0.006183f
C105 B.n71 VSUBS 0.006183f
C106 B.n72 VSUBS 0.006183f
C107 B.n73 VSUBS 0.006183f
C108 B.n74 VSUBS 0.006183f
C109 B.n75 VSUBS 0.006183f
C110 B.n76 VSUBS 0.006183f
C111 B.n77 VSUBS 0.006183f
C112 B.n78 VSUBS 0.006183f
C113 B.n79 VSUBS 0.006183f
C114 B.n80 VSUBS 0.006183f
C115 B.n81 VSUBS 0.006183f
C116 B.n82 VSUBS 0.006183f
C117 B.n83 VSUBS 0.006183f
C118 B.n84 VSUBS 0.006183f
C119 B.n85 VSUBS 0.006183f
C120 B.n86 VSUBS 0.006183f
C121 B.n87 VSUBS 0.006183f
C122 B.n88 VSUBS 0.006183f
C123 B.n89 VSUBS 0.014275f
C124 B.n90 VSUBS 0.006183f
C125 B.n91 VSUBS 0.006183f
C126 B.n92 VSUBS 0.006183f
C127 B.n93 VSUBS 0.006183f
C128 B.n94 VSUBS 0.006183f
C129 B.n95 VSUBS 0.006183f
C130 B.n96 VSUBS 0.006183f
C131 B.n97 VSUBS 0.006183f
C132 B.n98 VSUBS 0.006183f
C133 B.n99 VSUBS 0.006183f
C134 B.n100 VSUBS 0.006183f
C135 B.n101 VSUBS 0.006183f
C136 B.n102 VSUBS 0.006183f
C137 B.n103 VSUBS 0.006183f
C138 B.n104 VSUBS 0.006183f
C139 B.n105 VSUBS 0.006183f
C140 B.n106 VSUBS 0.006183f
C141 B.n107 VSUBS 0.006183f
C142 B.n108 VSUBS 0.006183f
C143 B.n109 VSUBS 0.006183f
C144 B.n110 VSUBS 0.006183f
C145 B.n111 VSUBS 0.006183f
C146 B.n112 VSUBS 0.006183f
C147 B.n113 VSUBS 0.006183f
C148 B.n114 VSUBS 0.006183f
C149 B.n115 VSUBS 0.006183f
C150 B.n116 VSUBS 0.006183f
C151 B.n117 VSUBS 0.006183f
C152 B.n118 VSUBS 0.006183f
C153 B.n119 VSUBS 0.006183f
C154 B.n120 VSUBS 0.006183f
C155 B.n121 VSUBS 0.015f
C156 B.n122 VSUBS 0.006183f
C157 B.n123 VSUBS 0.006183f
C158 B.n124 VSUBS 0.006183f
C159 B.n125 VSUBS 0.006183f
C160 B.n126 VSUBS 0.006183f
C161 B.n127 VSUBS 0.006183f
C162 B.n128 VSUBS 0.006183f
C163 B.n129 VSUBS 0.006183f
C164 B.n130 VSUBS 0.006183f
C165 B.n131 VSUBS 0.006183f
C166 B.n132 VSUBS 0.006183f
C167 B.n133 VSUBS 0.006183f
C168 B.n134 VSUBS 0.006183f
C169 B.n135 VSUBS 0.006183f
C170 B.n136 VSUBS 0.006183f
C171 B.n137 VSUBS 0.006183f
C172 B.n138 VSUBS 0.006183f
C173 B.n139 VSUBS 0.006183f
C174 B.n140 VSUBS 0.006183f
C175 B.n141 VSUBS 0.006183f
C176 B.n142 VSUBS 0.006183f
C177 B.n143 VSUBS 0.006183f
C178 B.n144 VSUBS 0.006183f
C179 B.n145 VSUBS 0.006183f
C180 B.n146 VSUBS 0.006183f
C181 B.n147 VSUBS 0.006183f
C182 B.n148 VSUBS 0.006183f
C183 B.n149 VSUBS 0.006183f
C184 B.n150 VSUBS 0.006183f
C185 B.n151 VSUBS 0.006183f
C186 B.n152 VSUBS 0.006183f
C187 B.t1 VSUBS 0.331288f
C188 B.t2 VSUBS 0.37007f
C189 B.t0 VSUBS 2.71492f
C190 B.n153 VSUBS 0.589028f
C191 B.n154 VSUBS 0.304086f
C192 B.n155 VSUBS 0.006183f
C193 B.n156 VSUBS 0.006183f
C194 B.n157 VSUBS 0.006183f
C195 B.n158 VSUBS 0.006183f
C196 B.t10 VSUBS 0.331284f
C197 B.t11 VSUBS 0.370067f
C198 B.t9 VSUBS 2.71492f
C199 B.n159 VSUBS 0.589031f
C200 B.n160 VSUBS 0.30409f
C201 B.n161 VSUBS 0.014326f
C202 B.n162 VSUBS 0.006183f
C203 B.n163 VSUBS 0.006183f
C204 B.n164 VSUBS 0.006183f
C205 B.n165 VSUBS 0.006183f
C206 B.n166 VSUBS 0.006183f
C207 B.n167 VSUBS 0.006183f
C208 B.n168 VSUBS 0.006183f
C209 B.n169 VSUBS 0.006183f
C210 B.n170 VSUBS 0.006183f
C211 B.n171 VSUBS 0.006183f
C212 B.n172 VSUBS 0.006183f
C213 B.n173 VSUBS 0.006183f
C214 B.n174 VSUBS 0.006183f
C215 B.n175 VSUBS 0.006183f
C216 B.n176 VSUBS 0.006183f
C217 B.n177 VSUBS 0.006183f
C218 B.n178 VSUBS 0.006183f
C219 B.n179 VSUBS 0.006183f
C220 B.n180 VSUBS 0.006183f
C221 B.n181 VSUBS 0.006183f
C222 B.n182 VSUBS 0.006183f
C223 B.n183 VSUBS 0.006183f
C224 B.n184 VSUBS 0.006183f
C225 B.n185 VSUBS 0.006183f
C226 B.n186 VSUBS 0.006183f
C227 B.n187 VSUBS 0.006183f
C228 B.n188 VSUBS 0.006183f
C229 B.n189 VSUBS 0.006183f
C230 B.n190 VSUBS 0.006183f
C231 B.n191 VSUBS 0.006183f
C232 B.n192 VSUBS 0.015f
C233 B.n193 VSUBS 0.006183f
C234 B.n194 VSUBS 0.006183f
C235 B.n195 VSUBS 0.006183f
C236 B.n196 VSUBS 0.006183f
C237 B.n197 VSUBS 0.006183f
C238 B.n198 VSUBS 0.006183f
C239 B.n199 VSUBS 0.006183f
C240 B.n200 VSUBS 0.006183f
C241 B.n201 VSUBS 0.006183f
C242 B.n202 VSUBS 0.006183f
C243 B.n203 VSUBS 0.006183f
C244 B.n204 VSUBS 0.006183f
C245 B.n205 VSUBS 0.006183f
C246 B.n206 VSUBS 0.006183f
C247 B.n207 VSUBS 0.006183f
C248 B.n208 VSUBS 0.006183f
C249 B.n209 VSUBS 0.006183f
C250 B.n210 VSUBS 0.006183f
C251 B.n211 VSUBS 0.006183f
C252 B.n212 VSUBS 0.006183f
C253 B.n213 VSUBS 0.006183f
C254 B.n214 VSUBS 0.006183f
C255 B.n215 VSUBS 0.006183f
C256 B.n216 VSUBS 0.006183f
C257 B.n217 VSUBS 0.006183f
C258 B.n218 VSUBS 0.006183f
C259 B.n219 VSUBS 0.006183f
C260 B.n220 VSUBS 0.006183f
C261 B.n221 VSUBS 0.006183f
C262 B.n222 VSUBS 0.006183f
C263 B.n223 VSUBS 0.006183f
C264 B.n224 VSUBS 0.006183f
C265 B.n225 VSUBS 0.006183f
C266 B.n226 VSUBS 0.006183f
C267 B.n227 VSUBS 0.006183f
C268 B.n228 VSUBS 0.006183f
C269 B.n229 VSUBS 0.006183f
C270 B.n230 VSUBS 0.006183f
C271 B.n231 VSUBS 0.006183f
C272 B.n232 VSUBS 0.006183f
C273 B.n233 VSUBS 0.006183f
C274 B.n234 VSUBS 0.006183f
C275 B.n235 VSUBS 0.006183f
C276 B.n236 VSUBS 0.006183f
C277 B.n237 VSUBS 0.006183f
C278 B.n238 VSUBS 0.006183f
C279 B.n239 VSUBS 0.006183f
C280 B.n240 VSUBS 0.006183f
C281 B.n241 VSUBS 0.006183f
C282 B.n242 VSUBS 0.006183f
C283 B.n243 VSUBS 0.006183f
C284 B.n244 VSUBS 0.006183f
C285 B.n245 VSUBS 0.006183f
C286 B.n246 VSUBS 0.006183f
C287 B.n247 VSUBS 0.006183f
C288 B.n248 VSUBS 0.006183f
C289 B.n249 VSUBS 0.006183f
C290 B.n250 VSUBS 0.006183f
C291 B.n251 VSUBS 0.014099f
C292 B.n252 VSUBS 0.014099f
C293 B.n253 VSUBS 0.015f
C294 B.n254 VSUBS 0.006183f
C295 B.n255 VSUBS 0.006183f
C296 B.n256 VSUBS 0.006183f
C297 B.n257 VSUBS 0.006183f
C298 B.n258 VSUBS 0.006183f
C299 B.n259 VSUBS 0.006183f
C300 B.n260 VSUBS 0.006183f
C301 B.n261 VSUBS 0.006183f
C302 B.n262 VSUBS 0.006183f
C303 B.n263 VSUBS 0.006183f
C304 B.n264 VSUBS 0.006183f
C305 B.n265 VSUBS 0.006183f
C306 B.n266 VSUBS 0.006183f
C307 B.n267 VSUBS 0.006183f
C308 B.n268 VSUBS 0.006183f
C309 B.n269 VSUBS 0.006183f
C310 B.n270 VSUBS 0.006183f
C311 B.n271 VSUBS 0.006183f
C312 B.n272 VSUBS 0.006183f
C313 B.n273 VSUBS 0.006183f
C314 B.n274 VSUBS 0.006183f
C315 B.n275 VSUBS 0.006183f
C316 B.n276 VSUBS 0.006183f
C317 B.n277 VSUBS 0.006183f
C318 B.n278 VSUBS 0.006183f
C319 B.n279 VSUBS 0.006183f
C320 B.n280 VSUBS 0.006183f
C321 B.n281 VSUBS 0.006183f
C322 B.n282 VSUBS 0.006183f
C323 B.n283 VSUBS 0.006183f
C324 B.n284 VSUBS 0.006183f
C325 B.n285 VSUBS 0.006183f
C326 B.n286 VSUBS 0.006183f
C327 B.n287 VSUBS 0.006183f
C328 B.n288 VSUBS 0.006183f
C329 B.n289 VSUBS 0.006183f
C330 B.n290 VSUBS 0.006183f
C331 B.n291 VSUBS 0.006183f
C332 B.n292 VSUBS 0.006183f
C333 B.n293 VSUBS 0.006183f
C334 B.n294 VSUBS 0.006183f
C335 B.n295 VSUBS 0.006183f
C336 B.n296 VSUBS 0.006183f
C337 B.n297 VSUBS 0.006183f
C338 B.n298 VSUBS 0.006183f
C339 B.n299 VSUBS 0.006183f
C340 B.n300 VSUBS 0.006183f
C341 B.n301 VSUBS 0.006183f
C342 B.n302 VSUBS 0.006183f
C343 B.n303 VSUBS 0.006183f
C344 B.n304 VSUBS 0.006183f
C345 B.n305 VSUBS 0.006183f
C346 B.n306 VSUBS 0.006183f
C347 B.n307 VSUBS 0.006183f
C348 B.n308 VSUBS 0.006183f
C349 B.n309 VSUBS 0.006183f
C350 B.n310 VSUBS 0.006183f
C351 B.n311 VSUBS 0.006183f
C352 B.n312 VSUBS 0.006183f
C353 B.n313 VSUBS 0.006183f
C354 B.n314 VSUBS 0.006183f
C355 B.n315 VSUBS 0.006183f
C356 B.n316 VSUBS 0.006183f
C357 B.n317 VSUBS 0.006183f
C358 B.n318 VSUBS 0.006183f
C359 B.n319 VSUBS 0.006183f
C360 B.n320 VSUBS 0.006183f
C361 B.n321 VSUBS 0.006183f
C362 B.n322 VSUBS 0.006183f
C363 B.n323 VSUBS 0.006183f
C364 B.n324 VSUBS 0.006183f
C365 B.n325 VSUBS 0.006183f
C366 B.n326 VSUBS 0.006183f
C367 B.n327 VSUBS 0.006183f
C368 B.n328 VSUBS 0.006183f
C369 B.n329 VSUBS 0.006183f
C370 B.n330 VSUBS 0.006183f
C371 B.n331 VSUBS 0.006183f
C372 B.n332 VSUBS 0.006183f
C373 B.n333 VSUBS 0.006183f
C374 B.n334 VSUBS 0.006183f
C375 B.n335 VSUBS 0.006183f
C376 B.n336 VSUBS 0.006183f
C377 B.n337 VSUBS 0.006183f
C378 B.n338 VSUBS 0.006183f
C379 B.n339 VSUBS 0.006183f
C380 B.n340 VSUBS 0.006183f
C381 B.n341 VSUBS 0.006183f
C382 B.n342 VSUBS 0.006183f
C383 B.n343 VSUBS 0.006183f
C384 B.n344 VSUBS 0.00582f
C385 B.n345 VSUBS 0.006183f
C386 B.n346 VSUBS 0.006183f
C387 B.n347 VSUBS 0.003455f
C388 B.n348 VSUBS 0.006183f
C389 B.n349 VSUBS 0.006183f
C390 B.n350 VSUBS 0.006183f
C391 B.n351 VSUBS 0.006183f
C392 B.n352 VSUBS 0.006183f
C393 B.n353 VSUBS 0.006183f
C394 B.n354 VSUBS 0.006183f
C395 B.n355 VSUBS 0.006183f
C396 B.n356 VSUBS 0.006183f
C397 B.n357 VSUBS 0.006183f
C398 B.n358 VSUBS 0.006183f
C399 B.n359 VSUBS 0.006183f
C400 B.n360 VSUBS 0.003455f
C401 B.n361 VSUBS 0.014326f
C402 B.n362 VSUBS 0.00582f
C403 B.n363 VSUBS 0.006183f
C404 B.n364 VSUBS 0.006183f
C405 B.n365 VSUBS 0.006183f
C406 B.n366 VSUBS 0.006183f
C407 B.n367 VSUBS 0.006183f
C408 B.n368 VSUBS 0.006183f
C409 B.n369 VSUBS 0.006183f
C410 B.n370 VSUBS 0.006183f
C411 B.n371 VSUBS 0.006183f
C412 B.n372 VSUBS 0.006183f
C413 B.n373 VSUBS 0.006183f
C414 B.n374 VSUBS 0.006183f
C415 B.n375 VSUBS 0.006183f
C416 B.n376 VSUBS 0.006183f
C417 B.n377 VSUBS 0.006183f
C418 B.n378 VSUBS 0.006183f
C419 B.n379 VSUBS 0.006183f
C420 B.n380 VSUBS 0.006183f
C421 B.n381 VSUBS 0.006183f
C422 B.n382 VSUBS 0.006183f
C423 B.n383 VSUBS 0.006183f
C424 B.n384 VSUBS 0.006183f
C425 B.n385 VSUBS 0.006183f
C426 B.n386 VSUBS 0.006183f
C427 B.n387 VSUBS 0.006183f
C428 B.n388 VSUBS 0.006183f
C429 B.n389 VSUBS 0.006183f
C430 B.n390 VSUBS 0.006183f
C431 B.n391 VSUBS 0.006183f
C432 B.n392 VSUBS 0.006183f
C433 B.n393 VSUBS 0.006183f
C434 B.n394 VSUBS 0.006183f
C435 B.n395 VSUBS 0.006183f
C436 B.n396 VSUBS 0.006183f
C437 B.n397 VSUBS 0.006183f
C438 B.n398 VSUBS 0.006183f
C439 B.n399 VSUBS 0.006183f
C440 B.n400 VSUBS 0.006183f
C441 B.n401 VSUBS 0.006183f
C442 B.n402 VSUBS 0.006183f
C443 B.n403 VSUBS 0.006183f
C444 B.n404 VSUBS 0.006183f
C445 B.n405 VSUBS 0.006183f
C446 B.n406 VSUBS 0.006183f
C447 B.n407 VSUBS 0.006183f
C448 B.n408 VSUBS 0.006183f
C449 B.n409 VSUBS 0.006183f
C450 B.n410 VSUBS 0.006183f
C451 B.n411 VSUBS 0.006183f
C452 B.n412 VSUBS 0.006183f
C453 B.n413 VSUBS 0.006183f
C454 B.n414 VSUBS 0.006183f
C455 B.n415 VSUBS 0.006183f
C456 B.n416 VSUBS 0.006183f
C457 B.n417 VSUBS 0.006183f
C458 B.n418 VSUBS 0.006183f
C459 B.n419 VSUBS 0.006183f
C460 B.n420 VSUBS 0.006183f
C461 B.n421 VSUBS 0.006183f
C462 B.n422 VSUBS 0.006183f
C463 B.n423 VSUBS 0.006183f
C464 B.n424 VSUBS 0.006183f
C465 B.n425 VSUBS 0.006183f
C466 B.n426 VSUBS 0.006183f
C467 B.n427 VSUBS 0.006183f
C468 B.n428 VSUBS 0.006183f
C469 B.n429 VSUBS 0.006183f
C470 B.n430 VSUBS 0.006183f
C471 B.n431 VSUBS 0.006183f
C472 B.n432 VSUBS 0.006183f
C473 B.n433 VSUBS 0.006183f
C474 B.n434 VSUBS 0.006183f
C475 B.n435 VSUBS 0.006183f
C476 B.n436 VSUBS 0.006183f
C477 B.n437 VSUBS 0.006183f
C478 B.n438 VSUBS 0.006183f
C479 B.n439 VSUBS 0.006183f
C480 B.n440 VSUBS 0.006183f
C481 B.n441 VSUBS 0.006183f
C482 B.n442 VSUBS 0.006183f
C483 B.n443 VSUBS 0.006183f
C484 B.n444 VSUBS 0.006183f
C485 B.n445 VSUBS 0.006183f
C486 B.n446 VSUBS 0.006183f
C487 B.n447 VSUBS 0.006183f
C488 B.n448 VSUBS 0.006183f
C489 B.n449 VSUBS 0.006183f
C490 B.n450 VSUBS 0.006183f
C491 B.n451 VSUBS 0.006183f
C492 B.n452 VSUBS 0.006183f
C493 B.n453 VSUBS 0.006183f
C494 B.n454 VSUBS 0.015f
C495 B.n455 VSUBS 0.014099f
C496 B.n456 VSUBS 0.014099f
C497 B.n457 VSUBS 0.006183f
C498 B.n458 VSUBS 0.006183f
C499 B.n459 VSUBS 0.006183f
C500 B.n460 VSUBS 0.006183f
C501 B.n461 VSUBS 0.006183f
C502 B.n462 VSUBS 0.006183f
C503 B.n463 VSUBS 0.006183f
C504 B.n464 VSUBS 0.006183f
C505 B.n465 VSUBS 0.006183f
C506 B.n466 VSUBS 0.006183f
C507 B.n467 VSUBS 0.006183f
C508 B.n468 VSUBS 0.006183f
C509 B.n469 VSUBS 0.006183f
C510 B.n470 VSUBS 0.006183f
C511 B.n471 VSUBS 0.006183f
C512 B.n472 VSUBS 0.006183f
C513 B.n473 VSUBS 0.006183f
C514 B.n474 VSUBS 0.006183f
C515 B.n475 VSUBS 0.006183f
C516 B.n476 VSUBS 0.006183f
C517 B.n477 VSUBS 0.006183f
C518 B.n478 VSUBS 0.006183f
C519 B.n479 VSUBS 0.006183f
C520 B.n480 VSUBS 0.006183f
C521 B.n481 VSUBS 0.006183f
C522 B.n482 VSUBS 0.006183f
C523 B.n483 VSUBS 0.006183f
C524 B.n484 VSUBS 0.006183f
C525 B.n485 VSUBS 0.006183f
C526 B.n486 VSUBS 0.006183f
C527 B.n487 VSUBS 0.006183f
C528 B.n488 VSUBS 0.006183f
C529 B.n489 VSUBS 0.006183f
C530 B.n490 VSUBS 0.006183f
C531 B.n491 VSUBS 0.006183f
C532 B.n492 VSUBS 0.006183f
C533 B.n493 VSUBS 0.006183f
C534 B.n494 VSUBS 0.006183f
C535 B.n495 VSUBS 0.006183f
C536 B.n496 VSUBS 0.006183f
C537 B.n497 VSUBS 0.006183f
C538 B.n498 VSUBS 0.006183f
C539 B.n499 VSUBS 0.006183f
C540 B.n500 VSUBS 0.006183f
C541 B.n501 VSUBS 0.006183f
C542 B.n502 VSUBS 0.006183f
C543 B.n503 VSUBS 0.006183f
C544 B.n504 VSUBS 0.006183f
C545 B.n505 VSUBS 0.006183f
C546 B.n506 VSUBS 0.006183f
C547 B.n507 VSUBS 0.006183f
C548 B.n508 VSUBS 0.006183f
C549 B.n509 VSUBS 0.006183f
C550 B.n510 VSUBS 0.006183f
C551 B.n511 VSUBS 0.006183f
C552 B.n512 VSUBS 0.006183f
C553 B.n513 VSUBS 0.006183f
C554 B.n514 VSUBS 0.006183f
C555 B.n515 VSUBS 0.006183f
C556 B.n516 VSUBS 0.006183f
C557 B.n517 VSUBS 0.006183f
C558 B.n518 VSUBS 0.006183f
C559 B.n519 VSUBS 0.006183f
C560 B.n520 VSUBS 0.006183f
C561 B.n521 VSUBS 0.006183f
C562 B.n522 VSUBS 0.006183f
C563 B.n523 VSUBS 0.006183f
C564 B.n524 VSUBS 0.006183f
C565 B.n525 VSUBS 0.006183f
C566 B.n526 VSUBS 0.006183f
C567 B.n527 VSUBS 0.006183f
C568 B.n528 VSUBS 0.006183f
C569 B.n529 VSUBS 0.006183f
C570 B.n530 VSUBS 0.006183f
C571 B.n531 VSUBS 0.006183f
C572 B.n532 VSUBS 0.006183f
C573 B.n533 VSUBS 0.006183f
C574 B.n534 VSUBS 0.006183f
C575 B.n535 VSUBS 0.006183f
C576 B.n536 VSUBS 0.006183f
C577 B.n537 VSUBS 0.006183f
C578 B.n538 VSUBS 0.006183f
C579 B.n539 VSUBS 0.006183f
C580 B.n540 VSUBS 0.006183f
C581 B.n541 VSUBS 0.006183f
C582 B.n542 VSUBS 0.006183f
C583 B.n543 VSUBS 0.006183f
C584 B.n544 VSUBS 0.006183f
C585 B.n545 VSUBS 0.006183f
C586 B.n546 VSUBS 0.006183f
C587 B.n547 VSUBS 0.006183f
C588 B.n548 VSUBS 0.014823f
C589 B.n549 VSUBS 0.014099f
C590 B.n550 VSUBS 0.015f
C591 B.n551 VSUBS 0.006183f
C592 B.n552 VSUBS 0.006183f
C593 B.n553 VSUBS 0.006183f
C594 B.n554 VSUBS 0.006183f
C595 B.n555 VSUBS 0.006183f
C596 B.n556 VSUBS 0.006183f
C597 B.n557 VSUBS 0.006183f
C598 B.n558 VSUBS 0.006183f
C599 B.n559 VSUBS 0.006183f
C600 B.n560 VSUBS 0.006183f
C601 B.n561 VSUBS 0.006183f
C602 B.n562 VSUBS 0.006183f
C603 B.n563 VSUBS 0.006183f
C604 B.n564 VSUBS 0.006183f
C605 B.n565 VSUBS 0.006183f
C606 B.n566 VSUBS 0.006183f
C607 B.n567 VSUBS 0.006183f
C608 B.n568 VSUBS 0.006183f
C609 B.n569 VSUBS 0.006183f
C610 B.n570 VSUBS 0.006183f
C611 B.n571 VSUBS 0.006183f
C612 B.n572 VSUBS 0.006183f
C613 B.n573 VSUBS 0.006183f
C614 B.n574 VSUBS 0.006183f
C615 B.n575 VSUBS 0.006183f
C616 B.n576 VSUBS 0.006183f
C617 B.n577 VSUBS 0.006183f
C618 B.n578 VSUBS 0.006183f
C619 B.n579 VSUBS 0.006183f
C620 B.n580 VSUBS 0.006183f
C621 B.n581 VSUBS 0.006183f
C622 B.n582 VSUBS 0.006183f
C623 B.n583 VSUBS 0.006183f
C624 B.n584 VSUBS 0.006183f
C625 B.n585 VSUBS 0.006183f
C626 B.n586 VSUBS 0.006183f
C627 B.n587 VSUBS 0.006183f
C628 B.n588 VSUBS 0.006183f
C629 B.n589 VSUBS 0.006183f
C630 B.n590 VSUBS 0.006183f
C631 B.n591 VSUBS 0.006183f
C632 B.n592 VSUBS 0.006183f
C633 B.n593 VSUBS 0.006183f
C634 B.n594 VSUBS 0.006183f
C635 B.n595 VSUBS 0.006183f
C636 B.n596 VSUBS 0.006183f
C637 B.n597 VSUBS 0.006183f
C638 B.n598 VSUBS 0.006183f
C639 B.n599 VSUBS 0.006183f
C640 B.n600 VSUBS 0.006183f
C641 B.n601 VSUBS 0.006183f
C642 B.n602 VSUBS 0.006183f
C643 B.n603 VSUBS 0.006183f
C644 B.n604 VSUBS 0.006183f
C645 B.n605 VSUBS 0.006183f
C646 B.n606 VSUBS 0.006183f
C647 B.n607 VSUBS 0.006183f
C648 B.n608 VSUBS 0.006183f
C649 B.n609 VSUBS 0.006183f
C650 B.n610 VSUBS 0.006183f
C651 B.n611 VSUBS 0.006183f
C652 B.n612 VSUBS 0.006183f
C653 B.n613 VSUBS 0.006183f
C654 B.n614 VSUBS 0.006183f
C655 B.n615 VSUBS 0.006183f
C656 B.n616 VSUBS 0.006183f
C657 B.n617 VSUBS 0.006183f
C658 B.n618 VSUBS 0.006183f
C659 B.n619 VSUBS 0.006183f
C660 B.n620 VSUBS 0.006183f
C661 B.n621 VSUBS 0.006183f
C662 B.n622 VSUBS 0.006183f
C663 B.n623 VSUBS 0.006183f
C664 B.n624 VSUBS 0.006183f
C665 B.n625 VSUBS 0.006183f
C666 B.n626 VSUBS 0.006183f
C667 B.n627 VSUBS 0.006183f
C668 B.n628 VSUBS 0.006183f
C669 B.n629 VSUBS 0.006183f
C670 B.n630 VSUBS 0.006183f
C671 B.n631 VSUBS 0.006183f
C672 B.n632 VSUBS 0.006183f
C673 B.n633 VSUBS 0.006183f
C674 B.n634 VSUBS 0.006183f
C675 B.n635 VSUBS 0.006183f
C676 B.n636 VSUBS 0.006183f
C677 B.n637 VSUBS 0.006183f
C678 B.n638 VSUBS 0.006183f
C679 B.n639 VSUBS 0.006183f
C680 B.n640 VSUBS 0.006183f
C681 B.n641 VSUBS 0.006183f
C682 B.n642 VSUBS 0.00582f
C683 B.n643 VSUBS 0.014326f
C684 B.n644 VSUBS 0.003455f
C685 B.n645 VSUBS 0.006183f
C686 B.n646 VSUBS 0.006183f
C687 B.n647 VSUBS 0.006183f
C688 B.n648 VSUBS 0.006183f
C689 B.n649 VSUBS 0.006183f
C690 B.n650 VSUBS 0.006183f
C691 B.n651 VSUBS 0.006183f
C692 B.n652 VSUBS 0.006183f
C693 B.n653 VSUBS 0.006183f
C694 B.n654 VSUBS 0.006183f
C695 B.n655 VSUBS 0.006183f
C696 B.n656 VSUBS 0.006183f
C697 B.n657 VSUBS 0.003455f
C698 B.n658 VSUBS 0.006183f
C699 B.n659 VSUBS 0.006183f
C700 B.n660 VSUBS 0.006183f
C701 B.n661 VSUBS 0.006183f
C702 B.n662 VSUBS 0.006183f
C703 B.n663 VSUBS 0.006183f
C704 B.n664 VSUBS 0.006183f
C705 B.n665 VSUBS 0.006183f
C706 B.n666 VSUBS 0.006183f
C707 B.n667 VSUBS 0.006183f
C708 B.n668 VSUBS 0.006183f
C709 B.n669 VSUBS 0.006183f
C710 B.n670 VSUBS 0.006183f
C711 B.n671 VSUBS 0.006183f
C712 B.n672 VSUBS 0.006183f
C713 B.n673 VSUBS 0.006183f
C714 B.n674 VSUBS 0.006183f
C715 B.n675 VSUBS 0.006183f
C716 B.n676 VSUBS 0.006183f
C717 B.n677 VSUBS 0.006183f
C718 B.n678 VSUBS 0.006183f
C719 B.n679 VSUBS 0.006183f
C720 B.n680 VSUBS 0.006183f
C721 B.n681 VSUBS 0.006183f
C722 B.n682 VSUBS 0.006183f
C723 B.n683 VSUBS 0.006183f
C724 B.n684 VSUBS 0.006183f
C725 B.n685 VSUBS 0.006183f
C726 B.n686 VSUBS 0.006183f
C727 B.n687 VSUBS 0.006183f
C728 B.n688 VSUBS 0.006183f
C729 B.n689 VSUBS 0.006183f
C730 B.n690 VSUBS 0.006183f
C731 B.n691 VSUBS 0.006183f
C732 B.n692 VSUBS 0.006183f
C733 B.n693 VSUBS 0.006183f
C734 B.n694 VSUBS 0.006183f
C735 B.n695 VSUBS 0.006183f
C736 B.n696 VSUBS 0.006183f
C737 B.n697 VSUBS 0.006183f
C738 B.n698 VSUBS 0.006183f
C739 B.n699 VSUBS 0.006183f
C740 B.n700 VSUBS 0.006183f
C741 B.n701 VSUBS 0.006183f
C742 B.n702 VSUBS 0.006183f
C743 B.n703 VSUBS 0.006183f
C744 B.n704 VSUBS 0.006183f
C745 B.n705 VSUBS 0.006183f
C746 B.n706 VSUBS 0.006183f
C747 B.n707 VSUBS 0.006183f
C748 B.n708 VSUBS 0.006183f
C749 B.n709 VSUBS 0.006183f
C750 B.n710 VSUBS 0.006183f
C751 B.n711 VSUBS 0.006183f
C752 B.n712 VSUBS 0.006183f
C753 B.n713 VSUBS 0.006183f
C754 B.n714 VSUBS 0.006183f
C755 B.n715 VSUBS 0.006183f
C756 B.n716 VSUBS 0.006183f
C757 B.n717 VSUBS 0.006183f
C758 B.n718 VSUBS 0.006183f
C759 B.n719 VSUBS 0.006183f
C760 B.n720 VSUBS 0.006183f
C761 B.n721 VSUBS 0.006183f
C762 B.n722 VSUBS 0.006183f
C763 B.n723 VSUBS 0.006183f
C764 B.n724 VSUBS 0.006183f
C765 B.n725 VSUBS 0.006183f
C766 B.n726 VSUBS 0.006183f
C767 B.n727 VSUBS 0.006183f
C768 B.n728 VSUBS 0.006183f
C769 B.n729 VSUBS 0.006183f
C770 B.n730 VSUBS 0.006183f
C771 B.n731 VSUBS 0.006183f
C772 B.n732 VSUBS 0.006183f
C773 B.n733 VSUBS 0.006183f
C774 B.n734 VSUBS 0.006183f
C775 B.n735 VSUBS 0.006183f
C776 B.n736 VSUBS 0.006183f
C777 B.n737 VSUBS 0.006183f
C778 B.n738 VSUBS 0.006183f
C779 B.n739 VSUBS 0.006183f
C780 B.n740 VSUBS 0.006183f
C781 B.n741 VSUBS 0.006183f
C782 B.n742 VSUBS 0.006183f
C783 B.n743 VSUBS 0.006183f
C784 B.n744 VSUBS 0.006183f
C785 B.n745 VSUBS 0.006183f
C786 B.n746 VSUBS 0.006183f
C787 B.n747 VSUBS 0.006183f
C788 B.n748 VSUBS 0.006183f
C789 B.n749 VSUBS 0.006183f
C790 B.n750 VSUBS 0.015f
C791 B.n751 VSUBS 0.015f
C792 B.n752 VSUBS 0.014099f
C793 B.n753 VSUBS 0.006183f
C794 B.n754 VSUBS 0.006183f
C795 B.n755 VSUBS 0.006183f
C796 B.n756 VSUBS 0.006183f
C797 B.n757 VSUBS 0.006183f
C798 B.n758 VSUBS 0.006183f
C799 B.n759 VSUBS 0.006183f
C800 B.n760 VSUBS 0.006183f
C801 B.n761 VSUBS 0.006183f
C802 B.n762 VSUBS 0.006183f
C803 B.n763 VSUBS 0.006183f
C804 B.n764 VSUBS 0.006183f
C805 B.n765 VSUBS 0.006183f
C806 B.n766 VSUBS 0.006183f
C807 B.n767 VSUBS 0.006183f
C808 B.n768 VSUBS 0.006183f
C809 B.n769 VSUBS 0.006183f
C810 B.n770 VSUBS 0.006183f
C811 B.n771 VSUBS 0.006183f
C812 B.n772 VSUBS 0.006183f
C813 B.n773 VSUBS 0.006183f
C814 B.n774 VSUBS 0.006183f
C815 B.n775 VSUBS 0.006183f
C816 B.n776 VSUBS 0.006183f
C817 B.n777 VSUBS 0.006183f
C818 B.n778 VSUBS 0.006183f
C819 B.n779 VSUBS 0.006183f
C820 B.n780 VSUBS 0.006183f
C821 B.n781 VSUBS 0.006183f
C822 B.n782 VSUBS 0.006183f
C823 B.n783 VSUBS 0.006183f
C824 B.n784 VSUBS 0.006183f
C825 B.n785 VSUBS 0.006183f
C826 B.n786 VSUBS 0.006183f
C827 B.n787 VSUBS 0.006183f
C828 B.n788 VSUBS 0.006183f
C829 B.n789 VSUBS 0.006183f
C830 B.n790 VSUBS 0.006183f
C831 B.n791 VSUBS 0.006183f
C832 B.n792 VSUBS 0.006183f
C833 B.n793 VSUBS 0.006183f
C834 B.n794 VSUBS 0.006183f
C835 B.n795 VSUBS 0.006183f
C836 B.n796 VSUBS 0.006183f
C837 B.n797 VSUBS 0.006183f
C838 B.n798 VSUBS 0.006183f
C839 B.n799 VSUBS 0.014001f
C840 VDD2.n0 VSUBS 0.0317f
C841 VDD2.n1 VSUBS 0.028303f
C842 VDD2.n2 VSUBS 0.015209f
C843 VDD2.n3 VSUBS 0.035948f
C844 VDD2.n4 VSUBS 0.016103f
C845 VDD2.n5 VSUBS 0.028303f
C846 VDD2.n6 VSUBS 0.015209f
C847 VDD2.n7 VSUBS 0.035948f
C848 VDD2.n8 VSUBS 0.016103f
C849 VDD2.n9 VSUBS 0.028303f
C850 VDD2.n10 VSUBS 0.015209f
C851 VDD2.n11 VSUBS 0.035948f
C852 VDD2.n12 VSUBS 0.016103f
C853 VDD2.n13 VSUBS 0.028303f
C854 VDD2.n14 VSUBS 0.015209f
C855 VDD2.n15 VSUBS 0.035948f
C856 VDD2.n16 VSUBS 0.016103f
C857 VDD2.n17 VSUBS 0.028303f
C858 VDD2.n18 VSUBS 0.015209f
C859 VDD2.n19 VSUBS 0.035948f
C860 VDD2.n20 VSUBS 0.016103f
C861 VDD2.n21 VSUBS 0.028303f
C862 VDD2.n22 VSUBS 0.015209f
C863 VDD2.n23 VSUBS 0.035948f
C864 VDD2.n24 VSUBS 0.016103f
C865 VDD2.n25 VSUBS 0.028303f
C866 VDD2.n26 VSUBS 0.015209f
C867 VDD2.n27 VSUBS 0.035948f
C868 VDD2.n28 VSUBS 0.016103f
C869 VDD2.n29 VSUBS 0.028303f
C870 VDD2.n30 VSUBS 0.015209f
C871 VDD2.n31 VSUBS 0.035948f
C872 VDD2.n32 VSUBS 0.016103f
C873 VDD2.n33 VSUBS 0.232736f
C874 VDD2.t0 VSUBS 0.077237f
C875 VDD2.n34 VSUBS 0.026961f
C876 VDD2.n35 VSUBS 0.022868f
C877 VDD2.n36 VSUBS 0.015209f
C878 VDD2.n37 VSUBS 2.31857f
C879 VDD2.n38 VSUBS 0.028303f
C880 VDD2.n39 VSUBS 0.015209f
C881 VDD2.n40 VSUBS 0.016103f
C882 VDD2.n41 VSUBS 0.035948f
C883 VDD2.n42 VSUBS 0.035948f
C884 VDD2.n43 VSUBS 0.016103f
C885 VDD2.n44 VSUBS 0.015209f
C886 VDD2.n45 VSUBS 0.028303f
C887 VDD2.n46 VSUBS 0.028303f
C888 VDD2.n47 VSUBS 0.015209f
C889 VDD2.n48 VSUBS 0.016103f
C890 VDD2.n49 VSUBS 0.035948f
C891 VDD2.n50 VSUBS 0.035948f
C892 VDD2.n51 VSUBS 0.016103f
C893 VDD2.n52 VSUBS 0.015209f
C894 VDD2.n53 VSUBS 0.028303f
C895 VDD2.n54 VSUBS 0.028303f
C896 VDD2.n55 VSUBS 0.015209f
C897 VDD2.n56 VSUBS 0.016103f
C898 VDD2.n57 VSUBS 0.035948f
C899 VDD2.n58 VSUBS 0.035948f
C900 VDD2.n59 VSUBS 0.016103f
C901 VDD2.n60 VSUBS 0.015209f
C902 VDD2.n61 VSUBS 0.028303f
C903 VDD2.n62 VSUBS 0.028303f
C904 VDD2.n63 VSUBS 0.015209f
C905 VDD2.n64 VSUBS 0.016103f
C906 VDD2.n65 VSUBS 0.035948f
C907 VDD2.n66 VSUBS 0.035948f
C908 VDD2.n67 VSUBS 0.016103f
C909 VDD2.n68 VSUBS 0.015209f
C910 VDD2.n69 VSUBS 0.028303f
C911 VDD2.n70 VSUBS 0.028303f
C912 VDD2.n71 VSUBS 0.015209f
C913 VDD2.n72 VSUBS 0.016103f
C914 VDD2.n73 VSUBS 0.035948f
C915 VDD2.n74 VSUBS 0.035948f
C916 VDD2.n75 VSUBS 0.035948f
C917 VDD2.n76 VSUBS 0.016103f
C918 VDD2.n77 VSUBS 0.015209f
C919 VDD2.n78 VSUBS 0.028303f
C920 VDD2.n79 VSUBS 0.028303f
C921 VDD2.n80 VSUBS 0.015209f
C922 VDD2.n81 VSUBS 0.015656f
C923 VDD2.n82 VSUBS 0.015656f
C924 VDD2.n83 VSUBS 0.035948f
C925 VDD2.n84 VSUBS 0.035948f
C926 VDD2.n85 VSUBS 0.016103f
C927 VDD2.n86 VSUBS 0.015209f
C928 VDD2.n87 VSUBS 0.028303f
C929 VDD2.n88 VSUBS 0.028303f
C930 VDD2.n89 VSUBS 0.015209f
C931 VDD2.n90 VSUBS 0.016103f
C932 VDD2.n91 VSUBS 0.035948f
C933 VDD2.n92 VSUBS 0.035948f
C934 VDD2.n93 VSUBS 0.016103f
C935 VDD2.n94 VSUBS 0.015209f
C936 VDD2.n95 VSUBS 0.028303f
C937 VDD2.n96 VSUBS 0.028303f
C938 VDD2.n97 VSUBS 0.015209f
C939 VDD2.n98 VSUBS 0.016103f
C940 VDD2.n99 VSUBS 0.035948f
C941 VDD2.n100 VSUBS 0.089075f
C942 VDD2.n101 VSUBS 0.016103f
C943 VDD2.n102 VSUBS 0.015209f
C944 VDD2.n103 VSUBS 0.066194f
C945 VDD2.n104 VSUBS 1.20717f
C946 VDD2.n105 VSUBS 0.0317f
C947 VDD2.n106 VSUBS 0.028303f
C948 VDD2.n107 VSUBS 0.015209f
C949 VDD2.n108 VSUBS 0.035948f
C950 VDD2.n109 VSUBS 0.016103f
C951 VDD2.n110 VSUBS 0.028303f
C952 VDD2.n111 VSUBS 0.015209f
C953 VDD2.n112 VSUBS 0.035948f
C954 VDD2.n113 VSUBS 0.016103f
C955 VDD2.n114 VSUBS 0.028303f
C956 VDD2.n115 VSUBS 0.015209f
C957 VDD2.n116 VSUBS 0.035948f
C958 VDD2.n117 VSUBS 0.016103f
C959 VDD2.n118 VSUBS 0.028303f
C960 VDD2.n119 VSUBS 0.015209f
C961 VDD2.n120 VSUBS 0.035948f
C962 VDD2.n121 VSUBS 0.035948f
C963 VDD2.n122 VSUBS 0.016103f
C964 VDD2.n123 VSUBS 0.028303f
C965 VDD2.n124 VSUBS 0.015209f
C966 VDD2.n125 VSUBS 0.035948f
C967 VDD2.n126 VSUBS 0.016103f
C968 VDD2.n127 VSUBS 0.028303f
C969 VDD2.n128 VSUBS 0.015209f
C970 VDD2.n129 VSUBS 0.035948f
C971 VDD2.n130 VSUBS 0.016103f
C972 VDD2.n131 VSUBS 0.028303f
C973 VDD2.n132 VSUBS 0.015209f
C974 VDD2.n133 VSUBS 0.035948f
C975 VDD2.n134 VSUBS 0.016103f
C976 VDD2.n135 VSUBS 0.028303f
C977 VDD2.n136 VSUBS 0.015209f
C978 VDD2.n137 VSUBS 0.035948f
C979 VDD2.n138 VSUBS 0.016103f
C980 VDD2.n139 VSUBS 0.232736f
C981 VDD2.t1 VSUBS 0.077237f
C982 VDD2.n140 VSUBS 0.026961f
C983 VDD2.n141 VSUBS 0.022868f
C984 VDD2.n142 VSUBS 0.015209f
C985 VDD2.n143 VSUBS 2.31857f
C986 VDD2.n144 VSUBS 0.028303f
C987 VDD2.n145 VSUBS 0.015209f
C988 VDD2.n146 VSUBS 0.016103f
C989 VDD2.n147 VSUBS 0.035948f
C990 VDD2.n148 VSUBS 0.035948f
C991 VDD2.n149 VSUBS 0.016103f
C992 VDD2.n150 VSUBS 0.015209f
C993 VDD2.n151 VSUBS 0.028303f
C994 VDD2.n152 VSUBS 0.028303f
C995 VDD2.n153 VSUBS 0.015209f
C996 VDD2.n154 VSUBS 0.016103f
C997 VDD2.n155 VSUBS 0.035948f
C998 VDD2.n156 VSUBS 0.035948f
C999 VDD2.n157 VSUBS 0.016103f
C1000 VDD2.n158 VSUBS 0.015209f
C1001 VDD2.n159 VSUBS 0.028303f
C1002 VDD2.n160 VSUBS 0.028303f
C1003 VDD2.n161 VSUBS 0.015209f
C1004 VDD2.n162 VSUBS 0.016103f
C1005 VDD2.n163 VSUBS 0.035948f
C1006 VDD2.n164 VSUBS 0.035948f
C1007 VDD2.n165 VSUBS 0.016103f
C1008 VDD2.n166 VSUBS 0.015209f
C1009 VDD2.n167 VSUBS 0.028303f
C1010 VDD2.n168 VSUBS 0.028303f
C1011 VDD2.n169 VSUBS 0.015209f
C1012 VDD2.n170 VSUBS 0.016103f
C1013 VDD2.n171 VSUBS 0.035948f
C1014 VDD2.n172 VSUBS 0.035948f
C1015 VDD2.n173 VSUBS 0.016103f
C1016 VDD2.n174 VSUBS 0.015209f
C1017 VDD2.n175 VSUBS 0.028303f
C1018 VDD2.n176 VSUBS 0.028303f
C1019 VDD2.n177 VSUBS 0.015209f
C1020 VDD2.n178 VSUBS 0.016103f
C1021 VDD2.n179 VSUBS 0.035948f
C1022 VDD2.n180 VSUBS 0.035948f
C1023 VDD2.n181 VSUBS 0.016103f
C1024 VDD2.n182 VSUBS 0.015209f
C1025 VDD2.n183 VSUBS 0.028303f
C1026 VDD2.n184 VSUBS 0.028303f
C1027 VDD2.n185 VSUBS 0.015209f
C1028 VDD2.n186 VSUBS 0.015656f
C1029 VDD2.n187 VSUBS 0.015656f
C1030 VDD2.n188 VSUBS 0.035948f
C1031 VDD2.n189 VSUBS 0.035948f
C1032 VDD2.n190 VSUBS 0.016103f
C1033 VDD2.n191 VSUBS 0.015209f
C1034 VDD2.n192 VSUBS 0.028303f
C1035 VDD2.n193 VSUBS 0.028303f
C1036 VDD2.n194 VSUBS 0.015209f
C1037 VDD2.n195 VSUBS 0.016103f
C1038 VDD2.n196 VSUBS 0.035948f
C1039 VDD2.n197 VSUBS 0.035948f
C1040 VDD2.n198 VSUBS 0.016103f
C1041 VDD2.n199 VSUBS 0.015209f
C1042 VDD2.n200 VSUBS 0.028303f
C1043 VDD2.n201 VSUBS 0.028303f
C1044 VDD2.n202 VSUBS 0.015209f
C1045 VDD2.n203 VSUBS 0.016103f
C1046 VDD2.n204 VSUBS 0.035948f
C1047 VDD2.n205 VSUBS 0.089075f
C1048 VDD2.n206 VSUBS 0.016103f
C1049 VDD2.n207 VSUBS 0.015209f
C1050 VDD2.n208 VSUBS 0.066194f
C1051 VDD2.n209 VSUBS 0.064446f
C1052 VDD2.n210 VSUBS 4.46982f
C1053 VN.t1 VSUBS 5.959569f
C1054 VN.t0 VSUBS 6.80819f
C1055 VDD1.n0 VSUBS 0.031885f
C1056 VDD1.n1 VSUBS 0.028468f
C1057 VDD1.n2 VSUBS 0.015297f
C1058 VDD1.n3 VSUBS 0.036157f
C1059 VDD1.n4 VSUBS 0.016197f
C1060 VDD1.n5 VSUBS 0.028468f
C1061 VDD1.n6 VSUBS 0.015297f
C1062 VDD1.n7 VSUBS 0.036157f
C1063 VDD1.n8 VSUBS 0.016197f
C1064 VDD1.n9 VSUBS 0.028468f
C1065 VDD1.n10 VSUBS 0.015297f
C1066 VDD1.n11 VSUBS 0.036157f
C1067 VDD1.n12 VSUBS 0.016197f
C1068 VDD1.n13 VSUBS 0.028468f
C1069 VDD1.n14 VSUBS 0.015297f
C1070 VDD1.n15 VSUBS 0.036157f
C1071 VDD1.n16 VSUBS 0.036157f
C1072 VDD1.n17 VSUBS 0.016197f
C1073 VDD1.n18 VSUBS 0.028468f
C1074 VDD1.n19 VSUBS 0.015297f
C1075 VDD1.n20 VSUBS 0.036157f
C1076 VDD1.n21 VSUBS 0.016197f
C1077 VDD1.n22 VSUBS 0.028468f
C1078 VDD1.n23 VSUBS 0.015297f
C1079 VDD1.n24 VSUBS 0.036157f
C1080 VDD1.n25 VSUBS 0.016197f
C1081 VDD1.n26 VSUBS 0.028468f
C1082 VDD1.n27 VSUBS 0.015297f
C1083 VDD1.n28 VSUBS 0.036157f
C1084 VDD1.n29 VSUBS 0.016197f
C1085 VDD1.n30 VSUBS 0.028468f
C1086 VDD1.n31 VSUBS 0.015297f
C1087 VDD1.n32 VSUBS 0.036157f
C1088 VDD1.n33 VSUBS 0.016197f
C1089 VDD1.n34 VSUBS 0.23409f
C1090 VDD1.t1 VSUBS 0.077687f
C1091 VDD1.n35 VSUBS 0.027118f
C1092 VDD1.n36 VSUBS 0.023001f
C1093 VDD1.n37 VSUBS 0.015297f
C1094 VDD1.n38 VSUBS 2.33206f
C1095 VDD1.n39 VSUBS 0.028468f
C1096 VDD1.n40 VSUBS 0.015297f
C1097 VDD1.n41 VSUBS 0.016197f
C1098 VDD1.n42 VSUBS 0.036157f
C1099 VDD1.n43 VSUBS 0.036157f
C1100 VDD1.n44 VSUBS 0.016197f
C1101 VDD1.n45 VSUBS 0.015297f
C1102 VDD1.n46 VSUBS 0.028468f
C1103 VDD1.n47 VSUBS 0.028468f
C1104 VDD1.n48 VSUBS 0.015297f
C1105 VDD1.n49 VSUBS 0.016197f
C1106 VDD1.n50 VSUBS 0.036157f
C1107 VDD1.n51 VSUBS 0.036157f
C1108 VDD1.n52 VSUBS 0.016197f
C1109 VDD1.n53 VSUBS 0.015297f
C1110 VDD1.n54 VSUBS 0.028468f
C1111 VDD1.n55 VSUBS 0.028468f
C1112 VDD1.n56 VSUBS 0.015297f
C1113 VDD1.n57 VSUBS 0.016197f
C1114 VDD1.n58 VSUBS 0.036157f
C1115 VDD1.n59 VSUBS 0.036157f
C1116 VDD1.n60 VSUBS 0.016197f
C1117 VDD1.n61 VSUBS 0.015297f
C1118 VDD1.n62 VSUBS 0.028468f
C1119 VDD1.n63 VSUBS 0.028468f
C1120 VDD1.n64 VSUBS 0.015297f
C1121 VDD1.n65 VSUBS 0.016197f
C1122 VDD1.n66 VSUBS 0.036157f
C1123 VDD1.n67 VSUBS 0.036157f
C1124 VDD1.n68 VSUBS 0.016197f
C1125 VDD1.n69 VSUBS 0.015297f
C1126 VDD1.n70 VSUBS 0.028468f
C1127 VDD1.n71 VSUBS 0.028468f
C1128 VDD1.n72 VSUBS 0.015297f
C1129 VDD1.n73 VSUBS 0.016197f
C1130 VDD1.n74 VSUBS 0.036157f
C1131 VDD1.n75 VSUBS 0.036157f
C1132 VDD1.n76 VSUBS 0.016197f
C1133 VDD1.n77 VSUBS 0.015297f
C1134 VDD1.n78 VSUBS 0.028468f
C1135 VDD1.n79 VSUBS 0.028468f
C1136 VDD1.n80 VSUBS 0.015297f
C1137 VDD1.n81 VSUBS 0.015747f
C1138 VDD1.n82 VSUBS 0.015747f
C1139 VDD1.n83 VSUBS 0.036157f
C1140 VDD1.n84 VSUBS 0.036157f
C1141 VDD1.n85 VSUBS 0.016197f
C1142 VDD1.n86 VSUBS 0.015297f
C1143 VDD1.n87 VSUBS 0.028468f
C1144 VDD1.n88 VSUBS 0.028468f
C1145 VDD1.n89 VSUBS 0.015297f
C1146 VDD1.n90 VSUBS 0.016197f
C1147 VDD1.n91 VSUBS 0.036157f
C1148 VDD1.n92 VSUBS 0.036157f
C1149 VDD1.n93 VSUBS 0.016197f
C1150 VDD1.n94 VSUBS 0.015297f
C1151 VDD1.n95 VSUBS 0.028468f
C1152 VDD1.n96 VSUBS 0.028468f
C1153 VDD1.n97 VSUBS 0.015297f
C1154 VDD1.n98 VSUBS 0.016197f
C1155 VDD1.n99 VSUBS 0.036157f
C1156 VDD1.n100 VSUBS 0.089593f
C1157 VDD1.n101 VSUBS 0.016197f
C1158 VDD1.n102 VSUBS 0.015297f
C1159 VDD1.n103 VSUBS 0.066579f
C1160 VDD1.n104 VSUBS 0.067298f
C1161 VDD1.n105 VSUBS 0.031885f
C1162 VDD1.n106 VSUBS 0.028468f
C1163 VDD1.n107 VSUBS 0.015297f
C1164 VDD1.n108 VSUBS 0.036157f
C1165 VDD1.n109 VSUBS 0.016197f
C1166 VDD1.n110 VSUBS 0.028468f
C1167 VDD1.n111 VSUBS 0.015297f
C1168 VDD1.n112 VSUBS 0.036157f
C1169 VDD1.n113 VSUBS 0.016197f
C1170 VDD1.n114 VSUBS 0.028468f
C1171 VDD1.n115 VSUBS 0.015297f
C1172 VDD1.n116 VSUBS 0.036157f
C1173 VDD1.n117 VSUBS 0.016197f
C1174 VDD1.n118 VSUBS 0.028468f
C1175 VDD1.n119 VSUBS 0.015297f
C1176 VDD1.n120 VSUBS 0.036157f
C1177 VDD1.n121 VSUBS 0.016197f
C1178 VDD1.n122 VSUBS 0.028468f
C1179 VDD1.n123 VSUBS 0.015297f
C1180 VDD1.n124 VSUBS 0.036157f
C1181 VDD1.n125 VSUBS 0.016197f
C1182 VDD1.n126 VSUBS 0.028468f
C1183 VDD1.n127 VSUBS 0.015297f
C1184 VDD1.n128 VSUBS 0.036157f
C1185 VDD1.n129 VSUBS 0.016197f
C1186 VDD1.n130 VSUBS 0.028468f
C1187 VDD1.n131 VSUBS 0.015297f
C1188 VDD1.n132 VSUBS 0.036157f
C1189 VDD1.n133 VSUBS 0.016197f
C1190 VDD1.n134 VSUBS 0.028468f
C1191 VDD1.n135 VSUBS 0.015297f
C1192 VDD1.n136 VSUBS 0.036157f
C1193 VDD1.n137 VSUBS 0.016197f
C1194 VDD1.n138 VSUBS 0.23409f
C1195 VDD1.t0 VSUBS 0.077687f
C1196 VDD1.n139 VSUBS 0.027118f
C1197 VDD1.n140 VSUBS 0.023001f
C1198 VDD1.n141 VSUBS 0.015297f
C1199 VDD1.n142 VSUBS 2.33206f
C1200 VDD1.n143 VSUBS 0.028468f
C1201 VDD1.n144 VSUBS 0.015297f
C1202 VDD1.n145 VSUBS 0.016197f
C1203 VDD1.n146 VSUBS 0.036157f
C1204 VDD1.n147 VSUBS 0.036157f
C1205 VDD1.n148 VSUBS 0.016197f
C1206 VDD1.n149 VSUBS 0.015297f
C1207 VDD1.n150 VSUBS 0.028468f
C1208 VDD1.n151 VSUBS 0.028468f
C1209 VDD1.n152 VSUBS 0.015297f
C1210 VDD1.n153 VSUBS 0.016197f
C1211 VDD1.n154 VSUBS 0.036157f
C1212 VDD1.n155 VSUBS 0.036157f
C1213 VDD1.n156 VSUBS 0.016197f
C1214 VDD1.n157 VSUBS 0.015297f
C1215 VDD1.n158 VSUBS 0.028468f
C1216 VDD1.n159 VSUBS 0.028468f
C1217 VDD1.n160 VSUBS 0.015297f
C1218 VDD1.n161 VSUBS 0.016197f
C1219 VDD1.n162 VSUBS 0.036157f
C1220 VDD1.n163 VSUBS 0.036157f
C1221 VDD1.n164 VSUBS 0.016197f
C1222 VDD1.n165 VSUBS 0.015297f
C1223 VDD1.n166 VSUBS 0.028468f
C1224 VDD1.n167 VSUBS 0.028468f
C1225 VDD1.n168 VSUBS 0.015297f
C1226 VDD1.n169 VSUBS 0.016197f
C1227 VDD1.n170 VSUBS 0.036157f
C1228 VDD1.n171 VSUBS 0.036157f
C1229 VDD1.n172 VSUBS 0.016197f
C1230 VDD1.n173 VSUBS 0.015297f
C1231 VDD1.n174 VSUBS 0.028468f
C1232 VDD1.n175 VSUBS 0.028468f
C1233 VDD1.n176 VSUBS 0.015297f
C1234 VDD1.n177 VSUBS 0.016197f
C1235 VDD1.n178 VSUBS 0.036157f
C1236 VDD1.n179 VSUBS 0.036157f
C1237 VDD1.n180 VSUBS 0.036157f
C1238 VDD1.n181 VSUBS 0.016197f
C1239 VDD1.n182 VSUBS 0.015297f
C1240 VDD1.n183 VSUBS 0.028468f
C1241 VDD1.n184 VSUBS 0.028468f
C1242 VDD1.n185 VSUBS 0.015297f
C1243 VDD1.n186 VSUBS 0.015747f
C1244 VDD1.n187 VSUBS 0.015747f
C1245 VDD1.n188 VSUBS 0.036157f
C1246 VDD1.n189 VSUBS 0.036157f
C1247 VDD1.n190 VSUBS 0.016197f
C1248 VDD1.n191 VSUBS 0.015297f
C1249 VDD1.n192 VSUBS 0.028468f
C1250 VDD1.n193 VSUBS 0.028468f
C1251 VDD1.n194 VSUBS 0.015297f
C1252 VDD1.n195 VSUBS 0.016197f
C1253 VDD1.n196 VSUBS 0.036157f
C1254 VDD1.n197 VSUBS 0.036157f
C1255 VDD1.n198 VSUBS 0.016197f
C1256 VDD1.n199 VSUBS 0.015297f
C1257 VDD1.n200 VSUBS 0.028468f
C1258 VDD1.n201 VSUBS 0.028468f
C1259 VDD1.n202 VSUBS 0.015297f
C1260 VDD1.n203 VSUBS 0.016197f
C1261 VDD1.n204 VSUBS 0.036157f
C1262 VDD1.n205 VSUBS 0.089593f
C1263 VDD1.n206 VSUBS 0.016197f
C1264 VDD1.n207 VSUBS 0.015297f
C1265 VDD1.n208 VSUBS 0.066579f
C1266 VDD1.n209 VSUBS 1.287f
C1267 VTAIL.n0 VSUBS 0.031844f
C1268 VTAIL.n1 VSUBS 0.028431f
C1269 VTAIL.n2 VSUBS 0.015278f
C1270 VTAIL.n3 VSUBS 0.036111f
C1271 VTAIL.n4 VSUBS 0.016176f
C1272 VTAIL.n5 VSUBS 0.028431f
C1273 VTAIL.n6 VSUBS 0.015278f
C1274 VTAIL.n7 VSUBS 0.036111f
C1275 VTAIL.n8 VSUBS 0.016176f
C1276 VTAIL.n9 VSUBS 0.028431f
C1277 VTAIL.n10 VSUBS 0.015278f
C1278 VTAIL.n11 VSUBS 0.036111f
C1279 VTAIL.n12 VSUBS 0.016176f
C1280 VTAIL.n13 VSUBS 0.028431f
C1281 VTAIL.n14 VSUBS 0.015278f
C1282 VTAIL.n15 VSUBS 0.036111f
C1283 VTAIL.n16 VSUBS 0.016176f
C1284 VTAIL.n17 VSUBS 0.028431f
C1285 VTAIL.n18 VSUBS 0.015278f
C1286 VTAIL.n19 VSUBS 0.036111f
C1287 VTAIL.n20 VSUBS 0.016176f
C1288 VTAIL.n21 VSUBS 0.028431f
C1289 VTAIL.n22 VSUBS 0.015278f
C1290 VTAIL.n23 VSUBS 0.036111f
C1291 VTAIL.n24 VSUBS 0.016176f
C1292 VTAIL.n25 VSUBS 0.028431f
C1293 VTAIL.n26 VSUBS 0.015278f
C1294 VTAIL.n27 VSUBS 0.036111f
C1295 VTAIL.n28 VSUBS 0.016176f
C1296 VTAIL.n29 VSUBS 0.028431f
C1297 VTAIL.n30 VSUBS 0.015278f
C1298 VTAIL.n31 VSUBS 0.036111f
C1299 VTAIL.n32 VSUBS 0.016176f
C1300 VTAIL.n33 VSUBS 0.233792f
C1301 VTAIL.t2 VSUBS 0.077588f
C1302 VTAIL.n34 VSUBS 0.027083f
C1303 VTAIL.n35 VSUBS 0.022972f
C1304 VTAIL.n36 VSUBS 0.015278f
C1305 VTAIL.n37 VSUBS 2.32909f
C1306 VTAIL.n38 VSUBS 0.028431f
C1307 VTAIL.n39 VSUBS 0.015278f
C1308 VTAIL.n40 VSUBS 0.016176f
C1309 VTAIL.n41 VSUBS 0.036111f
C1310 VTAIL.n42 VSUBS 0.036111f
C1311 VTAIL.n43 VSUBS 0.016176f
C1312 VTAIL.n44 VSUBS 0.015278f
C1313 VTAIL.n45 VSUBS 0.028431f
C1314 VTAIL.n46 VSUBS 0.028431f
C1315 VTAIL.n47 VSUBS 0.015278f
C1316 VTAIL.n48 VSUBS 0.016176f
C1317 VTAIL.n49 VSUBS 0.036111f
C1318 VTAIL.n50 VSUBS 0.036111f
C1319 VTAIL.n51 VSUBS 0.016176f
C1320 VTAIL.n52 VSUBS 0.015278f
C1321 VTAIL.n53 VSUBS 0.028431f
C1322 VTAIL.n54 VSUBS 0.028431f
C1323 VTAIL.n55 VSUBS 0.015278f
C1324 VTAIL.n56 VSUBS 0.016176f
C1325 VTAIL.n57 VSUBS 0.036111f
C1326 VTAIL.n58 VSUBS 0.036111f
C1327 VTAIL.n59 VSUBS 0.016176f
C1328 VTAIL.n60 VSUBS 0.015278f
C1329 VTAIL.n61 VSUBS 0.028431f
C1330 VTAIL.n62 VSUBS 0.028431f
C1331 VTAIL.n63 VSUBS 0.015278f
C1332 VTAIL.n64 VSUBS 0.016176f
C1333 VTAIL.n65 VSUBS 0.036111f
C1334 VTAIL.n66 VSUBS 0.036111f
C1335 VTAIL.n67 VSUBS 0.016176f
C1336 VTAIL.n68 VSUBS 0.015278f
C1337 VTAIL.n69 VSUBS 0.028431f
C1338 VTAIL.n70 VSUBS 0.028431f
C1339 VTAIL.n71 VSUBS 0.015278f
C1340 VTAIL.n72 VSUBS 0.016176f
C1341 VTAIL.n73 VSUBS 0.036111f
C1342 VTAIL.n74 VSUBS 0.036111f
C1343 VTAIL.n75 VSUBS 0.036111f
C1344 VTAIL.n76 VSUBS 0.016176f
C1345 VTAIL.n77 VSUBS 0.015278f
C1346 VTAIL.n78 VSUBS 0.028431f
C1347 VTAIL.n79 VSUBS 0.028431f
C1348 VTAIL.n80 VSUBS 0.015278f
C1349 VTAIL.n81 VSUBS 0.015727f
C1350 VTAIL.n82 VSUBS 0.015727f
C1351 VTAIL.n83 VSUBS 0.036111f
C1352 VTAIL.n84 VSUBS 0.036111f
C1353 VTAIL.n85 VSUBS 0.016176f
C1354 VTAIL.n86 VSUBS 0.015278f
C1355 VTAIL.n87 VSUBS 0.028431f
C1356 VTAIL.n88 VSUBS 0.028431f
C1357 VTAIL.n89 VSUBS 0.015278f
C1358 VTAIL.n90 VSUBS 0.016176f
C1359 VTAIL.n91 VSUBS 0.036111f
C1360 VTAIL.n92 VSUBS 0.036111f
C1361 VTAIL.n93 VSUBS 0.016176f
C1362 VTAIL.n94 VSUBS 0.015278f
C1363 VTAIL.n95 VSUBS 0.028431f
C1364 VTAIL.n96 VSUBS 0.028431f
C1365 VTAIL.n97 VSUBS 0.015278f
C1366 VTAIL.n98 VSUBS 0.016176f
C1367 VTAIL.n99 VSUBS 0.036111f
C1368 VTAIL.n100 VSUBS 0.089479f
C1369 VTAIL.n101 VSUBS 0.016176f
C1370 VTAIL.n102 VSUBS 0.015278f
C1371 VTAIL.n103 VSUBS 0.066494f
C1372 VTAIL.n104 VSUBS 0.045113f
C1373 VTAIL.n105 VSUBS 2.65304f
C1374 VTAIL.n106 VSUBS 0.031844f
C1375 VTAIL.n107 VSUBS 0.028431f
C1376 VTAIL.n108 VSUBS 0.015278f
C1377 VTAIL.n109 VSUBS 0.036111f
C1378 VTAIL.n110 VSUBS 0.016176f
C1379 VTAIL.n111 VSUBS 0.028431f
C1380 VTAIL.n112 VSUBS 0.015278f
C1381 VTAIL.n113 VSUBS 0.036111f
C1382 VTAIL.n114 VSUBS 0.016176f
C1383 VTAIL.n115 VSUBS 0.028431f
C1384 VTAIL.n116 VSUBS 0.015278f
C1385 VTAIL.n117 VSUBS 0.036111f
C1386 VTAIL.n118 VSUBS 0.016176f
C1387 VTAIL.n119 VSUBS 0.028431f
C1388 VTAIL.n120 VSUBS 0.015278f
C1389 VTAIL.n121 VSUBS 0.036111f
C1390 VTAIL.n122 VSUBS 0.036111f
C1391 VTAIL.n123 VSUBS 0.016176f
C1392 VTAIL.n124 VSUBS 0.028431f
C1393 VTAIL.n125 VSUBS 0.015278f
C1394 VTAIL.n126 VSUBS 0.036111f
C1395 VTAIL.n127 VSUBS 0.016176f
C1396 VTAIL.n128 VSUBS 0.028431f
C1397 VTAIL.n129 VSUBS 0.015278f
C1398 VTAIL.n130 VSUBS 0.036111f
C1399 VTAIL.n131 VSUBS 0.016176f
C1400 VTAIL.n132 VSUBS 0.028431f
C1401 VTAIL.n133 VSUBS 0.015278f
C1402 VTAIL.n134 VSUBS 0.036111f
C1403 VTAIL.n135 VSUBS 0.016176f
C1404 VTAIL.n136 VSUBS 0.028431f
C1405 VTAIL.n137 VSUBS 0.015278f
C1406 VTAIL.n138 VSUBS 0.036111f
C1407 VTAIL.n139 VSUBS 0.016176f
C1408 VTAIL.n140 VSUBS 0.233792f
C1409 VTAIL.t1 VSUBS 0.077588f
C1410 VTAIL.n141 VSUBS 0.027083f
C1411 VTAIL.n142 VSUBS 0.022972f
C1412 VTAIL.n143 VSUBS 0.015278f
C1413 VTAIL.n144 VSUBS 2.32909f
C1414 VTAIL.n145 VSUBS 0.028431f
C1415 VTAIL.n146 VSUBS 0.015278f
C1416 VTAIL.n147 VSUBS 0.016176f
C1417 VTAIL.n148 VSUBS 0.036111f
C1418 VTAIL.n149 VSUBS 0.036111f
C1419 VTAIL.n150 VSUBS 0.016176f
C1420 VTAIL.n151 VSUBS 0.015278f
C1421 VTAIL.n152 VSUBS 0.028431f
C1422 VTAIL.n153 VSUBS 0.028431f
C1423 VTAIL.n154 VSUBS 0.015278f
C1424 VTAIL.n155 VSUBS 0.016176f
C1425 VTAIL.n156 VSUBS 0.036111f
C1426 VTAIL.n157 VSUBS 0.036111f
C1427 VTAIL.n158 VSUBS 0.016176f
C1428 VTAIL.n159 VSUBS 0.015278f
C1429 VTAIL.n160 VSUBS 0.028431f
C1430 VTAIL.n161 VSUBS 0.028431f
C1431 VTAIL.n162 VSUBS 0.015278f
C1432 VTAIL.n163 VSUBS 0.016176f
C1433 VTAIL.n164 VSUBS 0.036111f
C1434 VTAIL.n165 VSUBS 0.036111f
C1435 VTAIL.n166 VSUBS 0.016176f
C1436 VTAIL.n167 VSUBS 0.015278f
C1437 VTAIL.n168 VSUBS 0.028431f
C1438 VTAIL.n169 VSUBS 0.028431f
C1439 VTAIL.n170 VSUBS 0.015278f
C1440 VTAIL.n171 VSUBS 0.016176f
C1441 VTAIL.n172 VSUBS 0.036111f
C1442 VTAIL.n173 VSUBS 0.036111f
C1443 VTAIL.n174 VSUBS 0.016176f
C1444 VTAIL.n175 VSUBS 0.015278f
C1445 VTAIL.n176 VSUBS 0.028431f
C1446 VTAIL.n177 VSUBS 0.028431f
C1447 VTAIL.n178 VSUBS 0.015278f
C1448 VTAIL.n179 VSUBS 0.016176f
C1449 VTAIL.n180 VSUBS 0.036111f
C1450 VTAIL.n181 VSUBS 0.036111f
C1451 VTAIL.n182 VSUBS 0.016176f
C1452 VTAIL.n183 VSUBS 0.015278f
C1453 VTAIL.n184 VSUBS 0.028431f
C1454 VTAIL.n185 VSUBS 0.028431f
C1455 VTAIL.n186 VSUBS 0.015278f
C1456 VTAIL.n187 VSUBS 0.015727f
C1457 VTAIL.n188 VSUBS 0.015727f
C1458 VTAIL.n189 VSUBS 0.036111f
C1459 VTAIL.n190 VSUBS 0.036111f
C1460 VTAIL.n191 VSUBS 0.016176f
C1461 VTAIL.n192 VSUBS 0.015278f
C1462 VTAIL.n193 VSUBS 0.028431f
C1463 VTAIL.n194 VSUBS 0.028431f
C1464 VTAIL.n195 VSUBS 0.015278f
C1465 VTAIL.n196 VSUBS 0.016176f
C1466 VTAIL.n197 VSUBS 0.036111f
C1467 VTAIL.n198 VSUBS 0.036111f
C1468 VTAIL.n199 VSUBS 0.016176f
C1469 VTAIL.n200 VSUBS 0.015278f
C1470 VTAIL.n201 VSUBS 0.028431f
C1471 VTAIL.n202 VSUBS 0.028431f
C1472 VTAIL.n203 VSUBS 0.015278f
C1473 VTAIL.n204 VSUBS 0.016176f
C1474 VTAIL.n205 VSUBS 0.036111f
C1475 VTAIL.n206 VSUBS 0.089479f
C1476 VTAIL.n207 VSUBS 0.016176f
C1477 VTAIL.n208 VSUBS 0.015278f
C1478 VTAIL.n209 VSUBS 0.066494f
C1479 VTAIL.n210 VSUBS 0.045113f
C1480 VTAIL.n211 VSUBS 2.72491f
C1481 VTAIL.n212 VSUBS 0.031844f
C1482 VTAIL.n213 VSUBS 0.028431f
C1483 VTAIL.n214 VSUBS 0.015278f
C1484 VTAIL.n215 VSUBS 0.036111f
C1485 VTAIL.n216 VSUBS 0.016176f
C1486 VTAIL.n217 VSUBS 0.028431f
C1487 VTAIL.n218 VSUBS 0.015278f
C1488 VTAIL.n219 VSUBS 0.036111f
C1489 VTAIL.n220 VSUBS 0.016176f
C1490 VTAIL.n221 VSUBS 0.028431f
C1491 VTAIL.n222 VSUBS 0.015278f
C1492 VTAIL.n223 VSUBS 0.036111f
C1493 VTAIL.n224 VSUBS 0.016176f
C1494 VTAIL.n225 VSUBS 0.028431f
C1495 VTAIL.n226 VSUBS 0.015278f
C1496 VTAIL.n227 VSUBS 0.036111f
C1497 VTAIL.n228 VSUBS 0.036111f
C1498 VTAIL.n229 VSUBS 0.016176f
C1499 VTAIL.n230 VSUBS 0.028431f
C1500 VTAIL.n231 VSUBS 0.015278f
C1501 VTAIL.n232 VSUBS 0.036111f
C1502 VTAIL.n233 VSUBS 0.016176f
C1503 VTAIL.n234 VSUBS 0.028431f
C1504 VTAIL.n235 VSUBS 0.015278f
C1505 VTAIL.n236 VSUBS 0.036111f
C1506 VTAIL.n237 VSUBS 0.016176f
C1507 VTAIL.n238 VSUBS 0.028431f
C1508 VTAIL.n239 VSUBS 0.015278f
C1509 VTAIL.n240 VSUBS 0.036111f
C1510 VTAIL.n241 VSUBS 0.016176f
C1511 VTAIL.n242 VSUBS 0.028431f
C1512 VTAIL.n243 VSUBS 0.015278f
C1513 VTAIL.n244 VSUBS 0.036111f
C1514 VTAIL.n245 VSUBS 0.016176f
C1515 VTAIL.n246 VSUBS 0.233792f
C1516 VTAIL.t3 VSUBS 0.077588f
C1517 VTAIL.n247 VSUBS 0.027083f
C1518 VTAIL.n248 VSUBS 0.022972f
C1519 VTAIL.n249 VSUBS 0.015278f
C1520 VTAIL.n250 VSUBS 2.32909f
C1521 VTAIL.n251 VSUBS 0.028431f
C1522 VTAIL.n252 VSUBS 0.015278f
C1523 VTAIL.n253 VSUBS 0.016176f
C1524 VTAIL.n254 VSUBS 0.036111f
C1525 VTAIL.n255 VSUBS 0.036111f
C1526 VTAIL.n256 VSUBS 0.016176f
C1527 VTAIL.n257 VSUBS 0.015278f
C1528 VTAIL.n258 VSUBS 0.028431f
C1529 VTAIL.n259 VSUBS 0.028431f
C1530 VTAIL.n260 VSUBS 0.015278f
C1531 VTAIL.n261 VSUBS 0.016176f
C1532 VTAIL.n262 VSUBS 0.036111f
C1533 VTAIL.n263 VSUBS 0.036111f
C1534 VTAIL.n264 VSUBS 0.016176f
C1535 VTAIL.n265 VSUBS 0.015278f
C1536 VTAIL.n266 VSUBS 0.028431f
C1537 VTAIL.n267 VSUBS 0.028431f
C1538 VTAIL.n268 VSUBS 0.015278f
C1539 VTAIL.n269 VSUBS 0.016176f
C1540 VTAIL.n270 VSUBS 0.036111f
C1541 VTAIL.n271 VSUBS 0.036111f
C1542 VTAIL.n272 VSUBS 0.016176f
C1543 VTAIL.n273 VSUBS 0.015278f
C1544 VTAIL.n274 VSUBS 0.028431f
C1545 VTAIL.n275 VSUBS 0.028431f
C1546 VTAIL.n276 VSUBS 0.015278f
C1547 VTAIL.n277 VSUBS 0.016176f
C1548 VTAIL.n278 VSUBS 0.036111f
C1549 VTAIL.n279 VSUBS 0.036111f
C1550 VTAIL.n280 VSUBS 0.016176f
C1551 VTAIL.n281 VSUBS 0.015278f
C1552 VTAIL.n282 VSUBS 0.028431f
C1553 VTAIL.n283 VSUBS 0.028431f
C1554 VTAIL.n284 VSUBS 0.015278f
C1555 VTAIL.n285 VSUBS 0.016176f
C1556 VTAIL.n286 VSUBS 0.036111f
C1557 VTAIL.n287 VSUBS 0.036111f
C1558 VTAIL.n288 VSUBS 0.016176f
C1559 VTAIL.n289 VSUBS 0.015278f
C1560 VTAIL.n290 VSUBS 0.028431f
C1561 VTAIL.n291 VSUBS 0.028431f
C1562 VTAIL.n292 VSUBS 0.015278f
C1563 VTAIL.n293 VSUBS 0.015727f
C1564 VTAIL.n294 VSUBS 0.015727f
C1565 VTAIL.n295 VSUBS 0.036111f
C1566 VTAIL.n296 VSUBS 0.036111f
C1567 VTAIL.n297 VSUBS 0.016176f
C1568 VTAIL.n298 VSUBS 0.015278f
C1569 VTAIL.n299 VSUBS 0.028431f
C1570 VTAIL.n300 VSUBS 0.028431f
C1571 VTAIL.n301 VSUBS 0.015278f
C1572 VTAIL.n302 VSUBS 0.016176f
C1573 VTAIL.n303 VSUBS 0.036111f
C1574 VTAIL.n304 VSUBS 0.036111f
C1575 VTAIL.n305 VSUBS 0.016176f
C1576 VTAIL.n306 VSUBS 0.015278f
C1577 VTAIL.n307 VSUBS 0.028431f
C1578 VTAIL.n308 VSUBS 0.028431f
C1579 VTAIL.n309 VSUBS 0.015278f
C1580 VTAIL.n310 VSUBS 0.016176f
C1581 VTAIL.n311 VSUBS 0.036111f
C1582 VTAIL.n312 VSUBS 0.089479f
C1583 VTAIL.n313 VSUBS 0.016176f
C1584 VTAIL.n314 VSUBS 0.015278f
C1585 VTAIL.n315 VSUBS 0.066494f
C1586 VTAIL.n316 VSUBS 0.045113f
C1587 VTAIL.n317 VSUBS 2.41612f
C1588 VTAIL.n318 VSUBS 0.031844f
C1589 VTAIL.n319 VSUBS 0.028431f
C1590 VTAIL.n320 VSUBS 0.015278f
C1591 VTAIL.n321 VSUBS 0.036111f
C1592 VTAIL.n322 VSUBS 0.016176f
C1593 VTAIL.n323 VSUBS 0.028431f
C1594 VTAIL.n324 VSUBS 0.015278f
C1595 VTAIL.n325 VSUBS 0.036111f
C1596 VTAIL.n326 VSUBS 0.016176f
C1597 VTAIL.n327 VSUBS 0.028431f
C1598 VTAIL.n328 VSUBS 0.015278f
C1599 VTAIL.n329 VSUBS 0.036111f
C1600 VTAIL.n330 VSUBS 0.016176f
C1601 VTAIL.n331 VSUBS 0.028431f
C1602 VTAIL.n332 VSUBS 0.015278f
C1603 VTAIL.n333 VSUBS 0.036111f
C1604 VTAIL.n334 VSUBS 0.016176f
C1605 VTAIL.n335 VSUBS 0.028431f
C1606 VTAIL.n336 VSUBS 0.015278f
C1607 VTAIL.n337 VSUBS 0.036111f
C1608 VTAIL.n338 VSUBS 0.016176f
C1609 VTAIL.n339 VSUBS 0.028431f
C1610 VTAIL.n340 VSUBS 0.015278f
C1611 VTAIL.n341 VSUBS 0.036111f
C1612 VTAIL.n342 VSUBS 0.016176f
C1613 VTAIL.n343 VSUBS 0.028431f
C1614 VTAIL.n344 VSUBS 0.015278f
C1615 VTAIL.n345 VSUBS 0.036111f
C1616 VTAIL.n346 VSUBS 0.016176f
C1617 VTAIL.n347 VSUBS 0.028431f
C1618 VTAIL.n348 VSUBS 0.015278f
C1619 VTAIL.n349 VSUBS 0.036111f
C1620 VTAIL.n350 VSUBS 0.016176f
C1621 VTAIL.n351 VSUBS 0.233792f
C1622 VTAIL.t0 VSUBS 0.077588f
C1623 VTAIL.n352 VSUBS 0.027083f
C1624 VTAIL.n353 VSUBS 0.022972f
C1625 VTAIL.n354 VSUBS 0.015278f
C1626 VTAIL.n355 VSUBS 2.32909f
C1627 VTAIL.n356 VSUBS 0.028431f
C1628 VTAIL.n357 VSUBS 0.015278f
C1629 VTAIL.n358 VSUBS 0.016176f
C1630 VTAIL.n359 VSUBS 0.036111f
C1631 VTAIL.n360 VSUBS 0.036111f
C1632 VTAIL.n361 VSUBS 0.016176f
C1633 VTAIL.n362 VSUBS 0.015278f
C1634 VTAIL.n363 VSUBS 0.028431f
C1635 VTAIL.n364 VSUBS 0.028431f
C1636 VTAIL.n365 VSUBS 0.015278f
C1637 VTAIL.n366 VSUBS 0.016176f
C1638 VTAIL.n367 VSUBS 0.036111f
C1639 VTAIL.n368 VSUBS 0.036111f
C1640 VTAIL.n369 VSUBS 0.016176f
C1641 VTAIL.n370 VSUBS 0.015278f
C1642 VTAIL.n371 VSUBS 0.028431f
C1643 VTAIL.n372 VSUBS 0.028431f
C1644 VTAIL.n373 VSUBS 0.015278f
C1645 VTAIL.n374 VSUBS 0.016176f
C1646 VTAIL.n375 VSUBS 0.036111f
C1647 VTAIL.n376 VSUBS 0.036111f
C1648 VTAIL.n377 VSUBS 0.016176f
C1649 VTAIL.n378 VSUBS 0.015278f
C1650 VTAIL.n379 VSUBS 0.028431f
C1651 VTAIL.n380 VSUBS 0.028431f
C1652 VTAIL.n381 VSUBS 0.015278f
C1653 VTAIL.n382 VSUBS 0.016176f
C1654 VTAIL.n383 VSUBS 0.036111f
C1655 VTAIL.n384 VSUBS 0.036111f
C1656 VTAIL.n385 VSUBS 0.016176f
C1657 VTAIL.n386 VSUBS 0.015278f
C1658 VTAIL.n387 VSUBS 0.028431f
C1659 VTAIL.n388 VSUBS 0.028431f
C1660 VTAIL.n389 VSUBS 0.015278f
C1661 VTAIL.n390 VSUBS 0.016176f
C1662 VTAIL.n391 VSUBS 0.036111f
C1663 VTAIL.n392 VSUBS 0.036111f
C1664 VTAIL.n393 VSUBS 0.036111f
C1665 VTAIL.n394 VSUBS 0.016176f
C1666 VTAIL.n395 VSUBS 0.015278f
C1667 VTAIL.n396 VSUBS 0.028431f
C1668 VTAIL.n397 VSUBS 0.028431f
C1669 VTAIL.n398 VSUBS 0.015278f
C1670 VTAIL.n399 VSUBS 0.015727f
C1671 VTAIL.n400 VSUBS 0.015727f
C1672 VTAIL.n401 VSUBS 0.036111f
C1673 VTAIL.n402 VSUBS 0.036111f
C1674 VTAIL.n403 VSUBS 0.016176f
C1675 VTAIL.n404 VSUBS 0.015278f
C1676 VTAIL.n405 VSUBS 0.028431f
C1677 VTAIL.n406 VSUBS 0.028431f
C1678 VTAIL.n407 VSUBS 0.015278f
C1679 VTAIL.n408 VSUBS 0.016176f
C1680 VTAIL.n409 VSUBS 0.036111f
C1681 VTAIL.n410 VSUBS 0.036111f
C1682 VTAIL.n411 VSUBS 0.016176f
C1683 VTAIL.n412 VSUBS 0.015278f
C1684 VTAIL.n413 VSUBS 0.028431f
C1685 VTAIL.n414 VSUBS 0.028431f
C1686 VTAIL.n415 VSUBS 0.015278f
C1687 VTAIL.n416 VSUBS 0.016176f
C1688 VTAIL.n417 VSUBS 0.036111f
C1689 VTAIL.n418 VSUBS 0.089479f
C1690 VTAIL.n419 VSUBS 0.016176f
C1691 VTAIL.n420 VSUBS 0.015278f
C1692 VTAIL.n421 VSUBS 0.066494f
C1693 VTAIL.n422 VSUBS 0.045113f
C1694 VTAIL.n423 VSUBS 2.29054f
C1695 VP.t0 VSUBS 7.073411f
C1696 VP.t1 VSUBS 6.1853f
C1697 VP.n0 VSUBS 6.42523f
.ends

