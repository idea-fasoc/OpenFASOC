* NGSPICE file created from diff_pair_sample_1286.ext - technology: sky130A

.subckt diff_pair_sample_1286 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=6.1425 ps=32.28 w=15.75 l=2.48
X1 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=0 ps=0 w=15.75 l=2.48
X2 VDD1.t7 VP.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=2.59875 ps=16.08 w=15.75 l=2.48
X3 VTAIL.t7 VP.t1 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=2.59875 ps=16.08 w=15.75 l=2.48
X4 VTAIL.t12 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=2.59875 ps=16.08 w=15.75 l=2.48
X5 VTAIL.t14 VN.t2 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=2.59875 ps=16.08 w=15.75 l=2.48
X6 VTAIL.t9 VN.t3 VDD2.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=2.59875 ps=16.08 w=15.75 l=2.48
X7 VTAIL.t8 VN.t4 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=2.59875 ps=16.08 w=15.75 l=2.48
X8 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=0 ps=0 w=15.75 l=2.48
X9 VTAIL.t5 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=2.59875 ps=16.08 w=15.75 l=2.48
X10 VDD1.t4 VP.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=6.1425 ps=32.28 w=15.75 l=2.48
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=0 ps=0 w=15.75 l=2.48
X12 VDD1.t3 VP.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=2.59875 ps=16.08 w=15.75 l=2.48
X13 VDD2.t2 VN.t5 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=6.1425 ps=32.28 w=15.75 l=2.48
X14 VDD2.t1 VN.t6 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=2.59875 ps=16.08 w=15.75 l=2.48
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=0 ps=0 w=15.75 l=2.48
X16 VDD2.t0 VN.t7 VTAIL.t13 B.t3 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=2.59875 ps=16.08 w=15.75 l=2.48
X17 VTAIL.t0 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=2.59875 ps=16.08 w=15.75 l=2.48
X18 VTAIL.t1 VP.t6 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=6.1425 pd=32.28 as=2.59875 ps=16.08 w=15.75 l=2.48
X19 VDD1.t0 VP.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.59875 pd=16.08 as=6.1425 ps=32.28 w=15.75 l=2.48
R0 VN.n6 VN.t3 186.806
R1 VN.n33 VN.t5 186.806
R2 VN.n51 VN.n27 161.3
R3 VN.n50 VN.n49 161.3
R4 VN.n48 VN.n28 161.3
R5 VN.n47 VN.n46 161.3
R6 VN.n45 VN.n29 161.3
R7 VN.n44 VN.n43 161.3
R8 VN.n42 VN.n41 161.3
R9 VN.n40 VN.n31 161.3
R10 VN.n39 VN.n38 161.3
R11 VN.n37 VN.n32 161.3
R12 VN.n36 VN.n35 161.3
R13 VN.n24 VN.n0 161.3
R14 VN.n23 VN.n22 161.3
R15 VN.n21 VN.n1 161.3
R16 VN.n20 VN.n19 161.3
R17 VN.n18 VN.n2 161.3
R18 VN.n17 VN.n16 161.3
R19 VN.n15 VN.n14 161.3
R20 VN.n13 VN.n4 161.3
R21 VN.n12 VN.n11 161.3
R22 VN.n10 VN.n5 161.3
R23 VN.n9 VN.n8 161.3
R24 VN.n7 VN.t7 153.054
R25 VN.n3 VN.t4 153.054
R26 VN.n25 VN.t0 153.054
R27 VN.n34 VN.t1 153.054
R28 VN.n30 VN.t6 153.054
R29 VN.n52 VN.t2 153.054
R30 VN.n26 VN.n25 100.236
R31 VN.n53 VN.n52 100.236
R32 VN.n19 VN.n1 56.5193
R33 VN.n46 VN.n28 56.5193
R34 VN VN.n53 53.4527
R35 VN.n7 VN.n6 52.6675
R36 VN.n34 VN.n33 52.6675
R37 VN.n12 VN.n5 40.4934
R38 VN.n13 VN.n12 40.4934
R39 VN.n39 VN.n32 40.4934
R40 VN.n40 VN.n39 40.4934
R41 VN.n8 VN.n5 24.4675
R42 VN.n14 VN.n13 24.4675
R43 VN.n18 VN.n17 24.4675
R44 VN.n19 VN.n18 24.4675
R45 VN.n23 VN.n1 24.4675
R46 VN.n24 VN.n23 24.4675
R47 VN.n35 VN.n32 24.4675
R48 VN.n46 VN.n45 24.4675
R49 VN.n45 VN.n44 24.4675
R50 VN.n41 VN.n40 24.4675
R51 VN.n51 VN.n50 24.4675
R52 VN.n50 VN.n28 24.4675
R53 VN.n8 VN.n7 19.8188
R54 VN.n14 VN.n3 19.8188
R55 VN.n35 VN.n34 19.8188
R56 VN.n41 VN.n30 19.8188
R57 VN.n25 VN.n24 10.5213
R58 VN.n52 VN.n51 10.5213
R59 VN.n36 VN.n33 6.81722
R60 VN.n9 VN.n6 6.81722
R61 VN.n17 VN.n3 4.64923
R62 VN.n44 VN.n30 4.64923
R63 VN.n53 VN.n27 0.278367
R64 VN.n26 VN.n0 0.278367
R65 VN.n49 VN.n27 0.189894
R66 VN.n49 VN.n48 0.189894
R67 VN.n48 VN.n47 0.189894
R68 VN.n47 VN.n29 0.189894
R69 VN.n43 VN.n29 0.189894
R70 VN.n43 VN.n42 0.189894
R71 VN.n42 VN.n31 0.189894
R72 VN.n38 VN.n31 0.189894
R73 VN.n38 VN.n37 0.189894
R74 VN.n37 VN.n36 0.189894
R75 VN.n10 VN.n9 0.189894
R76 VN.n11 VN.n10 0.189894
R77 VN.n11 VN.n4 0.189894
R78 VN.n15 VN.n4 0.189894
R79 VN.n16 VN.n15 0.189894
R80 VN.n16 VN.n2 0.189894
R81 VN.n20 VN.n2 0.189894
R82 VN.n21 VN.n20 0.189894
R83 VN.n22 VN.n21 0.189894
R84 VN.n22 VN.n0 0.189894
R85 VN VN.n26 0.153454
R86 VTAIL.n11 VTAIL.t5 45.9684
R87 VTAIL.n10 VTAIL.t15 45.9684
R88 VTAIL.n7 VTAIL.t14 45.9684
R89 VTAIL.n15 VTAIL.t11 45.9683
R90 VTAIL.n2 VTAIL.t9 45.9683
R91 VTAIL.n3 VTAIL.t2 45.9683
R92 VTAIL.n6 VTAIL.t1 45.9683
R93 VTAIL.n14 VTAIL.t6 45.9683
R94 VTAIL.n13 VTAIL.n12 44.7113
R95 VTAIL.n9 VTAIL.n8 44.7113
R96 VTAIL.n1 VTAIL.n0 44.7111
R97 VTAIL.n5 VTAIL.n4 44.7111
R98 VTAIL.n15 VTAIL.n14 28.3669
R99 VTAIL.n7 VTAIL.n6 28.3669
R100 VTAIL.n9 VTAIL.n7 2.42291
R101 VTAIL.n10 VTAIL.n9 2.42291
R102 VTAIL.n13 VTAIL.n11 2.42291
R103 VTAIL.n14 VTAIL.n13 2.42291
R104 VTAIL.n6 VTAIL.n5 2.42291
R105 VTAIL.n5 VTAIL.n3 2.42291
R106 VTAIL.n2 VTAIL.n1 2.42291
R107 VTAIL VTAIL.n15 2.36472
R108 VTAIL.n0 VTAIL.t13 1.25764
R109 VTAIL.n0 VTAIL.t8 1.25764
R110 VTAIL.n4 VTAIL.t4 1.25764
R111 VTAIL.n4 VTAIL.t0 1.25764
R112 VTAIL.n12 VTAIL.t3 1.25764
R113 VTAIL.n12 VTAIL.t7 1.25764
R114 VTAIL.n8 VTAIL.t10 1.25764
R115 VTAIL.n8 VTAIL.t12 1.25764
R116 VTAIL.n11 VTAIL.n10 0.470328
R117 VTAIL.n3 VTAIL.n2 0.470328
R118 VTAIL VTAIL.n1 0.0586897
R119 VDD2.n2 VDD2.n1 62.5457
R120 VDD2.n2 VDD2.n0 62.5457
R121 VDD2 VDD2.n5 62.543
R122 VDD2.n4 VDD2.n3 61.3901
R123 VDD2.n4 VDD2.n2 48.1937
R124 VDD2 VDD2.n4 1.2699
R125 VDD2.n5 VDD2.t6 1.25764
R126 VDD2.n5 VDD2.t2 1.25764
R127 VDD2.n3 VDD2.t5 1.25764
R128 VDD2.n3 VDD2.t1 1.25764
R129 VDD2.n1 VDD2.t3 1.25764
R130 VDD2.n1 VDD2.t7 1.25764
R131 VDD2.n0 VDD2.t4 1.25764
R132 VDD2.n0 VDD2.t0 1.25764
R133 B.n984 B.n983 585
R134 B.n985 B.n984 585
R135 B.n382 B.n149 585
R136 B.n381 B.n380 585
R137 B.n379 B.n378 585
R138 B.n377 B.n376 585
R139 B.n375 B.n374 585
R140 B.n373 B.n372 585
R141 B.n371 B.n370 585
R142 B.n369 B.n368 585
R143 B.n367 B.n366 585
R144 B.n365 B.n364 585
R145 B.n363 B.n362 585
R146 B.n361 B.n360 585
R147 B.n359 B.n358 585
R148 B.n357 B.n356 585
R149 B.n355 B.n354 585
R150 B.n353 B.n352 585
R151 B.n351 B.n350 585
R152 B.n349 B.n348 585
R153 B.n347 B.n346 585
R154 B.n345 B.n344 585
R155 B.n343 B.n342 585
R156 B.n341 B.n340 585
R157 B.n339 B.n338 585
R158 B.n337 B.n336 585
R159 B.n335 B.n334 585
R160 B.n333 B.n332 585
R161 B.n331 B.n330 585
R162 B.n329 B.n328 585
R163 B.n327 B.n326 585
R164 B.n325 B.n324 585
R165 B.n323 B.n322 585
R166 B.n321 B.n320 585
R167 B.n319 B.n318 585
R168 B.n317 B.n316 585
R169 B.n315 B.n314 585
R170 B.n313 B.n312 585
R171 B.n311 B.n310 585
R172 B.n309 B.n308 585
R173 B.n307 B.n306 585
R174 B.n305 B.n304 585
R175 B.n303 B.n302 585
R176 B.n301 B.n300 585
R177 B.n299 B.n298 585
R178 B.n297 B.n296 585
R179 B.n295 B.n294 585
R180 B.n293 B.n292 585
R181 B.n291 B.n290 585
R182 B.n289 B.n288 585
R183 B.n287 B.n286 585
R184 B.n285 B.n284 585
R185 B.n283 B.n282 585
R186 B.n281 B.n280 585
R187 B.n279 B.n278 585
R188 B.n277 B.n276 585
R189 B.n275 B.n274 585
R190 B.n273 B.n272 585
R191 B.n271 B.n270 585
R192 B.n269 B.n268 585
R193 B.n267 B.n266 585
R194 B.n265 B.n264 585
R195 B.n263 B.n262 585
R196 B.n260 B.n259 585
R197 B.n258 B.n257 585
R198 B.n256 B.n255 585
R199 B.n254 B.n253 585
R200 B.n252 B.n251 585
R201 B.n250 B.n249 585
R202 B.n248 B.n247 585
R203 B.n246 B.n245 585
R204 B.n244 B.n243 585
R205 B.n242 B.n241 585
R206 B.n240 B.n239 585
R207 B.n238 B.n237 585
R208 B.n236 B.n235 585
R209 B.n234 B.n233 585
R210 B.n232 B.n231 585
R211 B.n230 B.n229 585
R212 B.n228 B.n227 585
R213 B.n226 B.n225 585
R214 B.n224 B.n223 585
R215 B.n222 B.n221 585
R216 B.n220 B.n219 585
R217 B.n218 B.n217 585
R218 B.n216 B.n215 585
R219 B.n214 B.n213 585
R220 B.n212 B.n211 585
R221 B.n210 B.n209 585
R222 B.n208 B.n207 585
R223 B.n206 B.n205 585
R224 B.n204 B.n203 585
R225 B.n202 B.n201 585
R226 B.n200 B.n199 585
R227 B.n198 B.n197 585
R228 B.n196 B.n195 585
R229 B.n194 B.n193 585
R230 B.n192 B.n191 585
R231 B.n190 B.n189 585
R232 B.n188 B.n187 585
R233 B.n186 B.n185 585
R234 B.n184 B.n183 585
R235 B.n182 B.n181 585
R236 B.n180 B.n179 585
R237 B.n178 B.n177 585
R238 B.n176 B.n175 585
R239 B.n174 B.n173 585
R240 B.n172 B.n171 585
R241 B.n170 B.n169 585
R242 B.n168 B.n167 585
R243 B.n166 B.n165 585
R244 B.n164 B.n163 585
R245 B.n162 B.n161 585
R246 B.n160 B.n159 585
R247 B.n158 B.n157 585
R248 B.n156 B.n155 585
R249 B.n982 B.n91 585
R250 B.n986 B.n91 585
R251 B.n981 B.n90 585
R252 B.n987 B.n90 585
R253 B.n980 B.n979 585
R254 B.n979 B.n86 585
R255 B.n978 B.n85 585
R256 B.n993 B.n85 585
R257 B.n977 B.n84 585
R258 B.n994 B.n84 585
R259 B.n976 B.n83 585
R260 B.n995 B.n83 585
R261 B.n975 B.n974 585
R262 B.n974 B.n79 585
R263 B.n973 B.n78 585
R264 B.n1001 B.n78 585
R265 B.n972 B.n77 585
R266 B.n1002 B.n77 585
R267 B.n971 B.n76 585
R268 B.n1003 B.n76 585
R269 B.n970 B.n969 585
R270 B.n969 B.n72 585
R271 B.n968 B.n71 585
R272 B.n1009 B.n71 585
R273 B.n967 B.n70 585
R274 B.n1010 B.n70 585
R275 B.n966 B.n69 585
R276 B.n1011 B.n69 585
R277 B.n965 B.n964 585
R278 B.n964 B.n65 585
R279 B.n963 B.n64 585
R280 B.n1017 B.n64 585
R281 B.n962 B.n63 585
R282 B.n1018 B.n63 585
R283 B.n961 B.n62 585
R284 B.n1019 B.n62 585
R285 B.n960 B.n959 585
R286 B.n959 B.n61 585
R287 B.n958 B.n57 585
R288 B.n1025 B.n57 585
R289 B.n957 B.n56 585
R290 B.n1026 B.n56 585
R291 B.n956 B.n55 585
R292 B.n1027 B.n55 585
R293 B.n955 B.n954 585
R294 B.n954 B.n51 585
R295 B.n953 B.n50 585
R296 B.n1033 B.n50 585
R297 B.n952 B.n49 585
R298 B.n1034 B.n49 585
R299 B.n951 B.n48 585
R300 B.n1035 B.n48 585
R301 B.n950 B.n949 585
R302 B.n949 B.n44 585
R303 B.n948 B.n43 585
R304 B.n1041 B.n43 585
R305 B.n947 B.n42 585
R306 B.n1042 B.n42 585
R307 B.n946 B.n41 585
R308 B.n1043 B.n41 585
R309 B.n945 B.n944 585
R310 B.n944 B.n37 585
R311 B.n943 B.n36 585
R312 B.n1049 B.n36 585
R313 B.n942 B.n35 585
R314 B.n1050 B.n35 585
R315 B.n941 B.n34 585
R316 B.n1051 B.n34 585
R317 B.n940 B.n939 585
R318 B.n939 B.n30 585
R319 B.n938 B.n29 585
R320 B.n1057 B.n29 585
R321 B.n937 B.n28 585
R322 B.n1058 B.n28 585
R323 B.n936 B.n27 585
R324 B.n1059 B.n27 585
R325 B.n935 B.n934 585
R326 B.n934 B.n23 585
R327 B.n933 B.n22 585
R328 B.n1065 B.n22 585
R329 B.n932 B.n21 585
R330 B.n1066 B.n21 585
R331 B.n931 B.n20 585
R332 B.n1067 B.n20 585
R333 B.n930 B.n929 585
R334 B.n929 B.n16 585
R335 B.n928 B.n15 585
R336 B.n1073 B.n15 585
R337 B.n927 B.n14 585
R338 B.n1074 B.n14 585
R339 B.n926 B.n13 585
R340 B.n1075 B.n13 585
R341 B.n925 B.n924 585
R342 B.n924 B.n12 585
R343 B.n923 B.n922 585
R344 B.n923 B.n8 585
R345 B.n921 B.n7 585
R346 B.n1082 B.n7 585
R347 B.n920 B.n6 585
R348 B.n1083 B.n6 585
R349 B.n919 B.n5 585
R350 B.n1084 B.n5 585
R351 B.n918 B.n917 585
R352 B.n917 B.n4 585
R353 B.n916 B.n383 585
R354 B.n916 B.n915 585
R355 B.n906 B.n384 585
R356 B.n385 B.n384 585
R357 B.n908 B.n907 585
R358 B.n909 B.n908 585
R359 B.n905 B.n390 585
R360 B.n390 B.n389 585
R361 B.n904 B.n903 585
R362 B.n903 B.n902 585
R363 B.n392 B.n391 585
R364 B.n393 B.n392 585
R365 B.n895 B.n894 585
R366 B.n896 B.n895 585
R367 B.n893 B.n398 585
R368 B.n398 B.n397 585
R369 B.n892 B.n891 585
R370 B.n891 B.n890 585
R371 B.n400 B.n399 585
R372 B.n401 B.n400 585
R373 B.n883 B.n882 585
R374 B.n884 B.n883 585
R375 B.n881 B.n406 585
R376 B.n406 B.n405 585
R377 B.n880 B.n879 585
R378 B.n879 B.n878 585
R379 B.n408 B.n407 585
R380 B.n409 B.n408 585
R381 B.n871 B.n870 585
R382 B.n872 B.n871 585
R383 B.n869 B.n414 585
R384 B.n414 B.n413 585
R385 B.n868 B.n867 585
R386 B.n867 B.n866 585
R387 B.n416 B.n415 585
R388 B.n417 B.n416 585
R389 B.n859 B.n858 585
R390 B.n860 B.n859 585
R391 B.n857 B.n422 585
R392 B.n422 B.n421 585
R393 B.n856 B.n855 585
R394 B.n855 B.n854 585
R395 B.n424 B.n423 585
R396 B.n425 B.n424 585
R397 B.n847 B.n846 585
R398 B.n848 B.n847 585
R399 B.n845 B.n430 585
R400 B.n430 B.n429 585
R401 B.n844 B.n843 585
R402 B.n843 B.n842 585
R403 B.n432 B.n431 585
R404 B.n433 B.n432 585
R405 B.n835 B.n834 585
R406 B.n836 B.n835 585
R407 B.n833 B.n438 585
R408 B.n438 B.n437 585
R409 B.n832 B.n831 585
R410 B.n831 B.n830 585
R411 B.n440 B.n439 585
R412 B.n823 B.n440 585
R413 B.n822 B.n821 585
R414 B.n824 B.n822 585
R415 B.n820 B.n445 585
R416 B.n445 B.n444 585
R417 B.n819 B.n818 585
R418 B.n818 B.n817 585
R419 B.n447 B.n446 585
R420 B.n448 B.n447 585
R421 B.n810 B.n809 585
R422 B.n811 B.n810 585
R423 B.n808 B.n453 585
R424 B.n453 B.n452 585
R425 B.n807 B.n806 585
R426 B.n806 B.n805 585
R427 B.n455 B.n454 585
R428 B.n456 B.n455 585
R429 B.n798 B.n797 585
R430 B.n799 B.n798 585
R431 B.n796 B.n461 585
R432 B.n461 B.n460 585
R433 B.n795 B.n794 585
R434 B.n794 B.n793 585
R435 B.n463 B.n462 585
R436 B.n464 B.n463 585
R437 B.n786 B.n785 585
R438 B.n787 B.n786 585
R439 B.n784 B.n469 585
R440 B.n469 B.n468 585
R441 B.n783 B.n782 585
R442 B.n782 B.n781 585
R443 B.n471 B.n470 585
R444 B.n472 B.n471 585
R445 B.n774 B.n773 585
R446 B.n775 B.n774 585
R447 B.n772 B.n477 585
R448 B.n477 B.n476 585
R449 B.n766 B.n765 585
R450 B.n764 B.n536 585
R451 B.n763 B.n535 585
R452 B.n768 B.n535 585
R453 B.n762 B.n761 585
R454 B.n760 B.n759 585
R455 B.n758 B.n757 585
R456 B.n756 B.n755 585
R457 B.n754 B.n753 585
R458 B.n752 B.n751 585
R459 B.n750 B.n749 585
R460 B.n748 B.n747 585
R461 B.n746 B.n745 585
R462 B.n744 B.n743 585
R463 B.n742 B.n741 585
R464 B.n740 B.n739 585
R465 B.n738 B.n737 585
R466 B.n736 B.n735 585
R467 B.n734 B.n733 585
R468 B.n732 B.n731 585
R469 B.n730 B.n729 585
R470 B.n728 B.n727 585
R471 B.n726 B.n725 585
R472 B.n724 B.n723 585
R473 B.n722 B.n721 585
R474 B.n720 B.n719 585
R475 B.n718 B.n717 585
R476 B.n716 B.n715 585
R477 B.n714 B.n713 585
R478 B.n712 B.n711 585
R479 B.n710 B.n709 585
R480 B.n708 B.n707 585
R481 B.n706 B.n705 585
R482 B.n704 B.n703 585
R483 B.n702 B.n701 585
R484 B.n700 B.n699 585
R485 B.n698 B.n697 585
R486 B.n696 B.n695 585
R487 B.n694 B.n693 585
R488 B.n692 B.n691 585
R489 B.n690 B.n689 585
R490 B.n688 B.n687 585
R491 B.n686 B.n685 585
R492 B.n684 B.n683 585
R493 B.n682 B.n681 585
R494 B.n680 B.n679 585
R495 B.n678 B.n677 585
R496 B.n676 B.n675 585
R497 B.n674 B.n673 585
R498 B.n672 B.n671 585
R499 B.n670 B.n669 585
R500 B.n668 B.n667 585
R501 B.n666 B.n665 585
R502 B.n664 B.n663 585
R503 B.n662 B.n661 585
R504 B.n660 B.n659 585
R505 B.n658 B.n657 585
R506 B.n656 B.n655 585
R507 B.n654 B.n653 585
R508 B.n652 B.n651 585
R509 B.n650 B.n649 585
R510 B.n648 B.n647 585
R511 B.n646 B.n645 585
R512 B.n643 B.n642 585
R513 B.n641 B.n640 585
R514 B.n639 B.n638 585
R515 B.n637 B.n636 585
R516 B.n635 B.n634 585
R517 B.n633 B.n632 585
R518 B.n631 B.n630 585
R519 B.n629 B.n628 585
R520 B.n627 B.n626 585
R521 B.n625 B.n624 585
R522 B.n623 B.n622 585
R523 B.n621 B.n620 585
R524 B.n619 B.n618 585
R525 B.n617 B.n616 585
R526 B.n615 B.n614 585
R527 B.n613 B.n612 585
R528 B.n611 B.n610 585
R529 B.n609 B.n608 585
R530 B.n607 B.n606 585
R531 B.n605 B.n604 585
R532 B.n603 B.n602 585
R533 B.n601 B.n600 585
R534 B.n599 B.n598 585
R535 B.n597 B.n596 585
R536 B.n595 B.n594 585
R537 B.n593 B.n592 585
R538 B.n591 B.n590 585
R539 B.n589 B.n588 585
R540 B.n587 B.n586 585
R541 B.n585 B.n584 585
R542 B.n583 B.n582 585
R543 B.n581 B.n580 585
R544 B.n579 B.n578 585
R545 B.n577 B.n576 585
R546 B.n575 B.n574 585
R547 B.n573 B.n572 585
R548 B.n571 B.n570 585
R549 B.n569 B.n568 585
R550 B.n567 B.n566 585
R551 B.n565 B.n564 585
R552 B.n563 B.n562 585
R553 B.n561 B.n560 585
R554 B.n559 B.n558 585
R555 B.n557 B.n556 585
R556 B.n555 B.n554 585
R557 B.n553 B.n552 585
R558 B.n551 B.n550 585
R559 B.n549 B.n548 585
R560 B.n547 B.n546 585
R561 B.n545 B.n544 585
R562 B.n543 B.n542 585
R563 B.n479 B.n478 585
R564 B.n771 B.n770 585
R565 B.n475 B.n474 585
R566 B.n476 B.n475 585
R567 B.n777 B.n776 585
R568 B.n776 B.n775 585
R569 B.n778 B.n473 585
R570 B.n473 B.n472 585
R571 B.n780 B.n779 585
R572 B.n781 B.n780 585
R573 B.n467 B.n466 585
R574 B.n468 B.n467 585
R575 B.n789 B.n788 585
R576 B.n788 B.n787 585
R577 B.n790 B.n465 585
R578 B.n465 B.n464 585
R579 B.n792 B.n791 585
R580 B.n793 B.n792 585
R581 B.n459 B.n458 585
R582 B.n460 B.n459 585
R583 B.n801 B.n800 585
R584 B.n800 B.n799 585
R585 B.n802 B.n457 585
R586 B.n457 B.n456 585
R587 B.n804 B.n803 585
R588 B.n805 B.n804 585
R589 B.n451 B.n450 585
R590 B.n452 B.n451 585
R591 B.n813 B.n812 585
R592 B.n812 B.n811 585
R593 B.n814 B.n449 585
R594 B.n449 B.n448 585
R595 B.n816 B.n815 585
R596 B.n817 B.n816 585
R597 B.n443 B.n442 585
R598 B.n444 B.n443 585
R599 B.n826 B.n825 585
R600 B.n825 B.n824 585
R601 B.n827 B.n441 585
R602 B.n823 B.n441 585
R603 B.n829 B.n828 585
R604 B.n830 B.n829 585
R605 B.n436 B.n435 585
R606 B.n437 B.n436 585
R607 B.n838 B.n837 585
R608 B.n837 B.n836 585
R609 B.n839 B.n434 585
R610 B.n434 B.n433 585
R611 B.n841 B.n840 585
R612 B.n842 B.n841 585
R613 B.n428 B.n427 585
R614 B.n429 B.n428 585
R615 B.n850 B.n849 585
R616 B.n849 B.n848 585
R617 B.n851 B.n426 585
R618 B.n426 B.n425 585
R619 B.n853 B.n852 585
R620 B.n854 B.n853 585
R621 B.n420 B.n419 585
R622 B.n421 B.n420 585
R623 B.n862 B.n861 585
R624 B.n861 B.n860 585
R625 B.n863 B.n418 585
R626 B.n418 B.n417 585
R627 B.n865 B.n864 585
R628 B.n866 B.n865 585
R629 B.n412 B.n411 585
R630 B.n413 B.n412 585
R631 B.n874 B.n873 585
R632 B.n873 B.n872 585
R633 B.n875 B.n410 585
R634 B.n410 B.n409 585
R635 B.n877 B.n876 585
R636 B.n878 B.n877 585
R637 B.n404 B.n403 585
R638 B.n405 B.n404 585
R639 B.n886 B.n885 585
R640 B.n885 B.n884 585
R641 B.n887 B.n402 585
R642 B.n402 B.n401 585
R643 B.n889 B.n888 585
R644 B.n890 B.n889 585
R645 B.n396 B.n395 585
R646 B.n397 B.n396 585
R647 B.n898 B.n897 585
R648 B.n897 B.n896 585
R649 B.n899 B.n394 585
R650 B.n394 B.n393 585
R651 B.n901 B.n900 585
R652 B.n902 B.n901 585
R653 B.n388 B.n387 585
R654 B.n389 B.n388 585
R655 B.n911 B.n910 585
R656 B.n910 B.n909 585
R657 B.n912 B.n386 585
R658 B.n386 B.n385 585
R659 B.n914 B.n913 585
R660 B.n915 B.n914 585
R661 B.n3 B.n0 585
R662 B.n4 B.n3 585
R663 B.n1081 B.n1 585
R664 B.n1082 B.n1081 585
R665 B.n1080 B.n1079 585
R666 B.n1080 B.n8 585
R667 B.n1078 B.n9 585
R668 B.n12 B.n9 585
R669 B.n1077 B.n1076 585
R670 B.n1076 B.n1075 585
R671 B.n11 B.n10 585
R672 B.n1074 B.n11 585
R673 B.n1072 B.n1071 585
R674 B.n1073 B.n1072 585
R675 B.n1070 B.n17 585
R676 B.n17 B.n16 585
R677 B.n1069 B.n1068 585
R678 B.n1068 B.n1067 585
R679 B.n19 B.n18 585
R680 B.n1066 B.n19 585
R681 B.n1064 B.n1063 585
R682 B.n1065 B.n1064 585
R683 B.n1062 B.n24 585
R684 B.n24 B.n23 585
R685 B.n1061 B.n1060 585
R686 B.n1060 B.n1059 585
R687 B.n26 B.n25 585
R688 B.n1058 B.n26 585
R689 B.n1056 B.n1055 585
R690 B.n1057 B.n1056 585
R691 B.n1054 B.n31 585
R692 B.n31 B.n30 585
R693 B.n1053 B.n1052 585
R694 B.n1052 B.n1051 585
R695 B.n33 B.n32 585
R696 B.n1050 B.n33 585
R697 B.n1048 B.n1047 585
R698 B.n1049 B.n1048 585
R699 B.n1046 B.n38 585
R700 B.n38 B.n37 585
R701 B.n1045 B.n1044 585
R702 B.n1044 B.n1043 585
R703 B.n40 B.n39 585
R704 B.n1042 B.n40 585
R705 B.n1040 B.n1039 585
R706 B.n1041 B.n1040 585
R707 B.n1038 B.n45 585
R708 B.n45 B.n44 585
R709 B.n1037 B.n1036 585
R710 B.n1036 B.n1035 585
R711 B.n47 B.n46 585
R712 B.n1034 B.n47 585
R713 B.n1032 B.n1031 585
R714 B.n1033 B.n1032 585
R715 B.n1030 B.n52 585
R716 B.n52 B.n51 585
R717 B.n1029 B.n1028 585
R718 B.n1028 B.n1027 585
R719 B.n54 B.n53 585
R720 B.n1026 B.n54 585
R721 B.n1024 B.n1023 585
R722 B.n1025 B.n1024 585
R723 B.n1022 B.n58 585
R724 B.n61 B.n58 585
R725 B.n1021 B.n1020 585
R726 B.n1020 B.n1019 585
R727 B.n60 B.n59 585
R728 B.n1018 B.n60 585
R729 B.n1016 B.n1015 585
R730 B.n1017 B.n1016 585
R731 B.n1014 B.n66 585
R732 B.n66 B.n65 585
R733 B.n1013 B.n1012 585
R734 B.n1012 B.n1011 585
R735 B.n68 B.n67 585
R736 B.n1010 B.n68 585
R737 B.n1008 B.n1007 585
R738 B.n1009 B.n1008 585
R739 B.n1006 B.n73 585
R740 B.n73 B.n72 585
R741 B.n1005 B.n1004 585
R742 B.n1004 B.n1003 585
R743 B.n75 B.n74 585
R744 B.n1002 B.n75 585
R745 B.n1000 B.n999 585
R746 B.n1001 B.n1000 585
R747 B.n998 B.n80 585
R748 B.n80 B.n79 585
R749 B.n997 B.n996 585
R750 B.n996 B.n995 585
R751 B.n82 B.n81 585
R752 B.n994 B.n82 585
R753 B.n992 B.n991 585
R754 B.n993 B.n992 585
R755 B.n990 B.n87 585
R756 B.n87 B.n86 585
R757 B.n989 B.n988 585
R758 B.n988 B.n987 585
R759 B.n89 B.n88 585
R760 B.n986 B.n89 585
R761 B.n1085 B.n1084 585
R762 B.n1083 B.n2 585
R763 B.n155 B.n89 478.086
R764 B.n984 B.n91 478.086
R765 B.n770 B.n477 478.086
R766 B.n766 B.n475 478.086
R767 B.n153 B.t16 360.913
R768 B.n150 B.t8 360.913
R769 B.n540 B.t12 360.913
R770 B.n537 B.t19 360.913
R771 B.n985 B.n148 256.663
R772 B.n985 B.n147 256.663
R773 B.n985 B.n146 256.663
R774 B.n985 B.n145 256.663
R775 B.n985 B.n144 256.663
R776 B.n985 B.n143 256.663
R777 B.n985 B.n142 256.663
R778 B.n985 B.n141 256.663
R779 B.n985 B.n140 256.663
R780 B.n985 B.n139 256.663
R781 B.n985 B.n138 256.663
R782 B.n985 B.n137 256.663
R783 B.n985 B.n136 256.663
R784 B.n985 B.n135 256.663
R785 B.n985 B.n134 256.663
R786 B.n985 B.n133 256.663
R787 B.n985 B.n132 256.663
R788 B.n985 B.n131 256.663
R789 B.n985 B.n130 256.663
R790 B.n985 B.n129 256.663
R791 B.n985 B.n128 256.663
R792 B.n985 B.n127 256.663
R793 B.n985 B.n126 256.663
R794 B.n985 B.n125 256.663
R795 B.n985 B.n124 256.663
R796 B.n985 B.n123 256.663
R797 B.n985 B.n122 256.663
R798 B.n985 B.n121 256.663
R799 B.n985 B.n120 256.663
R800 B.n985 B.n119 256.663
R801 B.n985 B.n118 256.663
R802 B.n985 B.n117 256.663
R803 B.n985 B.n116 256.663
R804 B.n985 B.n115 256.663
R805 B.n985 B.n114 256.663
R806 B.n985 B.n113 256.663
R807 B.n985 B.n112 256.663
R808 B.n985 B.n111 256.663
R809 B.n985 B.n110 256.663
R810 B.n985 B.n109 256.663
R811 B.n985 B.n108 256.663
R812 B.n985 B.n107 256.663
R813 B.n985 B.n106 256.663
R814 B.n985 B.n105 256.663
R815 B.n985 B.n104 256.663
R816 B.n985 B.n103 256.663
R817 B.n985 B.n102 256.663
R818 B.n985 B.n101 256.663
R819 B.n985 B.n100 256.663
R820 B.n985 B.n99 256.663
R821 B.n985 B.n98 256.663
R822 B.n985 B.n97 256.663
R823 B.n985 B.n96 256.663
R824 B.n985 B.n95 256.663
R825 B.n985 B.n94 256.663
R826 B.n985 B.n93 256.663
R827 B.n985 B.n92 256.663
R828 B.n768 B.n767 256.663
R829 B.n768 B.n480 256.663
R830 B.n768 B.n481 256.663
R831 B.n768 B.n482 256.663
R832 B.n768 B.n483 256.663
R833 B.n768 B.n484 256.663
R834 B.n768 B.n485 256.663
R835 B.n768 B.n486 256.663
R836 B.n768 B.n487 256.663
R837 B.n768 B.n488 256.663
R838 B.n768 B.n489 256.663
R839 B.n768 B.n490 256.663
R840 B.n768 B.n491 256.663
R841 B.n768 B.n492 256.663
R842 B.n768 B.n493 256.663
R843 B.n768 B.n494 256.663
R844 B.n768 B.n495 256.663
R845 B.n768 B.n496 256.663
R846 B.n768 B.n497 256.663
R847 B.n768 B.n498 256.663
R848 B.n768 B.n499 256.663
R849 B.n768 B.n500 256.663
R850 B.n768 B.n501 256.663
R851 B.n768 B.n502 256.663
R852 B.n768 B.n503 256.663
R853 B.n768 B.n504 256.663
R854 B.n768 B.n505 256.663
R855 B.n768 B.n506 256.663
R856 B.n768 B.n507 256.663
R857 B.n768 B.n508 256.663
R858 B.n768 B.n509 256.663
R859 B.n768 B.n510 256.663
R860 B.n768 B.n511 256.663
R861 B.n768 B.n512 256.663
R862 B.n768 B.n513 256.663
R863 B.n768 B.n514 256.663
R864 B.n768 B.n515 256.663
R865 B.n768 B.n516 256.663
R866 B.n768 B.n517 256.663
R867 B.n768 B.n518 256.663
R868 B.n768 B.n519 256.663
R869 B.n768 B.n520 256.663
R870 B.n768 B.n521 256.663
R871 B.n768 B.n522 256.663
R872 B.n768 B.n523 256.663
R873 B.n768 B.n524 256.663
R874 B.n768 B.n525 256.663
R875 B.n768 B.n526 256.663
R876 B.n768 B.n527 256.663
R877 B.n768 B.n528 256.663
R878 B.n768 B.n529 256.663
R879 B.n768 B.n530 256.663
R880 B.n768 B.n531 256.663
R881 B.n768 B.n532 256.663
R882 B.n768 B.n533 256.663
R883 B.n768 B.n534 256.663
R884 B.n769 B.n768 256.663
R885 B.n1087 B.n1086 256.663
R886 B.n159 B.n158 163.367
R887 B.n163 B.n162 163.367
R888 B.n167 B.n166 163.367
R889 B.n171 B.n170 163.367
R890 B.n175 B.n174 163.367
R891 B.n179 B.n178 163.367
R892 B.n183 B.n182 163.367
R893 B.n187 B.n186 163.367
R894 B.n191 B.n190 163.367
R895 B.n195 B.n194 163.367
R896 B.n199 B.n198 163.367
R897 B.n203 B.n202 163.367
R898 B.n207 B.n206 163.367
R899 B.n211 B.n210 163.367
R900 B.n215 B.n214 163.367
R901 B.n219 B.n218 163.367
R902 B.n223 B.n222 163.367
R903 B.n227 B.n226 163.367
R904 B.n231 B.n230 163.367
R905 B.n235 B.n234 163.367
R906 B.n239 B.n238 163.367
R907 B.n243 B.n242 163.367
R908 B.n247 B.n246 163.367
R909 B.n251 B.n250 163.367
R910 B.n255 B.n254 163.367
R911 B.n259 B.n258 163.367
R912 B.n264 B.n263 163.367
R913 B.n268 B.n267 163.367
R914 B.n272 B.n271 163.367
R915 B.n276 B.n275 163.367
R916 B.n280 B.n279 163.367
R917 B.n284 B.n283 163.367
R918 B.n288 B.n287 163.367
R919 B.n292 B.n291 163.367
R920 B.n296 B.n295 163.367
R921 B.n300 B.n299 163.367
R922 B.n304 B.n303 163.367
R923 B.n308 B.n307 163.367
R924 B.n312 B.n311 163.367
R925 B.n316 B.n315 163.367
R926 B.n320 B.n319 163.367
R927 B.n324 B.n323 163.367
R928 B.n328 B.n327 163.367
R929 B.n332 B.n331 163.367
R930 B.n336 B.n335 163.367
R931 B.n340 B.n339 163.367
R932 B.n344 B.n343 163.367
R933 B.n348 B.n347 163.367
R934 B.n352 B.n351 163.367
R935 B.n356 B.n355 163.367
R936 B.n360 B.n359 163.367
R937 B.n364 B.n363 163.367
R938 B.n368 B.n367 163.367
R939 B.n372 B.n371 163.367
R940 B.n376 B.n375 163.367
R941 B.n380 B.n379 163.367
R942 B.n984 B.n149 163.367
R943 B.n774 B.n477 163.367
R944 B.n774 B.n471 163.367
R945 B.n782 B.n471 163.367
R946 B.n782 B.n469 163.367
R947 B.n786 B.n469 163.367
R948 B.n786 B.n463 163.367
R949 B.n794 B.n463 163.367
R950 B.n794 B.n461 163.367
R951 B.n798 B.n461 163.367
R952 B.n798 B.n455 163.367
R953 B.n806 B.n455 163.367
R954 B.n806 B.n453 163.367
R955 B.n810 B.n453 163.367
R956 B.n810 B.n447 163.367
R957 B.n818 B.n447 163.367
R958 B.n818 B.n445 163.367
R959 B.n822 B.n445 163.367
R960 B.n822 B.n440 163.367
R961 B.n831 B.n440 163.367
R962 B.n831 B.n438 163.367
R963 B.n835 B.n438 163.367
R964 B.n835 B.n432 163.367
R965 B.n843 B.n432 163.367
R966 B.n843 B.n430 163.367
R967 B.n847 B.n430 163.367
R968 B.n847 B.n424 163.367
R969 B.n855 B.n424 163.367
R970 B.n855 B.n422 163.367
R971 B.n859 B.n422 163.367
R972 B.n859 B.n416 163.367
R973 B.n867 B.n416 163.367
R974 B.n867 B.n414 163.367
R975 B.n871 B.n414 163.367
R976 B.n871 B.n408 163.367
R977 B.n879 B.n408 163.367
R978 B.n879 B.n406 163.367
R979 B.n883 B.n406 163.367
R980 B.n883 B.n400 163.367
R981 B.n891 B.n400 163.367
R982 B.n891 B.n398 163.367
R983 B.n895 B.n398 163.367
R984 B.n895 B.n392 163.367
R985 B.n903 B.n392 163.367
R986 B.n903 B.n390 163.367
R987 B.n908 B.n390 163.367
R988 B.n908 B.n384 163.367
R989 B.n916 B.n384 163.367
R990 B.n917 B.n916 163.367
R991 B.n917 B.n5 163.367
R992 B.n6 B.n5 163.367
R993 B.n7 B.n6 163.367
R994 B.n923 B.n7 163.367
R995 B.n924 B.n923 163.367
R996 B.n924 B.n13 163.367
R997 B.n14 B.n13 163.367
R998 B.n15 B.n14 163.367
R999 B.n929 B.n15 163.367
R1000 B.n929 B.n20 163.367
R1001 B.n21 B.n20 163.367
R1002 B.n22 B.n21 163.367
R1003 B.n934 B.n22 163.367
R1004 B.n934 B.n27 163.367
R1005 B.n28 B.n27 163.367
R1006 B.n29 B.n28 163.367
R1007 B.n939 B.n29 163.367
R1008 B.n939 B.n34 163.367
R1009 B.n35 B.n34 163.367
R1010 B.n36 B.n35 163.367
R1011 B.n944 B.n36 163.367
R1012 B.n944 B.n41 163.367
R1013 B.n42 B.n41 163.367
R1014 B.n43 B.n42 163.367
R1015 B.n949 B.n43 163.367
R1016 B.n949 B.n48 163.367
R1017 B.n49 B.n48 163.367
R1018 B.n50 B.n49 163.367
R1019 B.n954 B.n50 163.367
R1020 B.n954 B.n55 163.367
R1021 B.n56 B.n55 163.367
R1022 B.n57 B.n56 163.367
R1023 B.n959 B.n57 163.367
R1024 B.n959 B.n62 163.367
R1025 B.n63 B.n62 163.367
R1026 B.n64 B.n63 163.367
R1027 B.n964 B.n64 163.367
R1028 B.n964 B.n69 163.367
R1029 B.n70 B.n69 163.367
R1030 B.n71 B.n70 163.367
R1031 B.n969 B.n71 163.367
R1032 B.n969 B.n76 163.367
R1033 B.n77 B.n76 163.367
R1034 B.n78 B.n77 163.367
R1035 B.n974 B.n78 163.367
R1036 B.n974 B.n83 163.367
R1037 B.n84 B.n83 163.367
R1038 B.n85 B.n84 163.367
R1039 B.n979 B.n85 163.367
R1040 B.n979 B.n90 163.367
R1041 B.n91 B.n90 163.367
R1042 B.n536 B.n535 163.367
R1043 B.n761 B.n535 163.367
R1044 B.n759 B.n758 163.367
R1045 B.n755 B.n754 163.367
R1046 B.n751 B.n750 163.367
R1047 B.n747 B.n746 163.367
R1048 B.n743 B.n742 163.367
R1049 B.n739 B.n738 163.367
R1050 B.n735 B.n734 163.367
R1051 B.n731 B.n730 163.367
R1052 B.n727 B.n726 163.367
R1053 B.n723 B.n722 163.367
R1054 B.n719 B.n718 163.367
R1055 B.n715 B.n714 163.367
R1056 B.n711 B.n710 163.367
R1057 B.n707 B.n706 163.367
R1058 B.n703 B.n702 163.367
R1059 B.n699 B.n698 163.367
R1060 B.n695 B.n694 163.367
R1061 B.n691 B.n690 163.367
R1062 B.n687 B.n686 163.367
R1063 B.n683 B.n682 163.367
R1064 B.n679 B.n678 163.367
R1065 B.n675 B.n674 163.367
R1066 B.n671 B.n670 163.367
R1067 B.n667 B.n666 163.367
R1068 B.n663 B.n662 163.367
R1069 B.n659 B.n658 163.367
R1070 B.n655 B.n654 163.367
R1071 B.n651 B.n650 163.367
R1072 B.n647 B.n646 163.367
R1073 B.n642 B.n641 163.367
R1074 B.n638 B.n637 163.367
R1075 B.n634 B.n633 163.367
R1076 B.n630 B.n629 163.367
R1077 B.n626 B.n625 163.367
R1078 B.n622 B.n621 163.367
R1079 B.n618 B.n617 163.367
R1080 B.n614 B.n613 163.367
R1081 B.n610 B.n609 163.367
R1082 B.n606 B.n605 163.367
R1083 B.n602 B.n601 163.367
R1084 B.n598 B.n597 163.367
R1085 B.n594 B.n593 163.367
R1086 B.n590 B.n589 163.367
R1087 B.n586 B.n585 163.367
R1088 B.n582 B.n581 163.367
R1089 B.n578 B.n577 163.367
R1090 B.n574 B.n573 163.367
R1091 B.n570 B.n569 163.367
R1092 B.n566 B.n565 163.367
R1093 B.n562 B.n561 163.367
R1094 B.n558 B.n557 163.367
R1095 B.n554 B.n553 163.367
R1096 B.n550 B.n549 163.367
R1097 B.n546 B.n545 163.367
R1098 B.n542 B.n479 163.367
R1099 B.n776 B.n475 163.367
R1100 B.n776 B.n473 163.367
R1101 B.n780 B.n473 163.367
R1102 B.n780 B.n467 163.367
R1103 B.n788 B.n467 163.367
R1104 B.n788 B.n465 163.367
R1105 B.n792 B.n465 163.367
R1106 B.n792 B.n459 163.367
R1107 B.n800 B.n459 163.367
R1108 B.n800 B.n457 163.367
R1109 B.n804 B.n457 163.367
R1110 B.n804 B.n451 163.367
R1111 B.n812 B.n451 163.367
R1112 B.n812 B.n449 163.367
R1113 B.n816 B.n449 163.367
R1114 B.n816 B.n443 163.367
R1115 B.n825 B.n443 163.367
R1116 B.n825 B.n441 163.367
R1117 B.n829 B.n441 163.367
R1118 B.n829 B.n436 163.367
R1119 B.n837 B.n436 163.367
R1120 B.n837 B.n434 163.367
R1121 B.n841 B.n434 163.367
R1122 B.n841 B.n428 163.367
R1123 B.n849 B.n428 163.367
R1124 B.n849 B.n426 163.367
R1125 B.n853 B.n426 163.367
R1126 B.n853 B.n420 163.367
R1127 B.n861 B.n420 163.367
R1128 B.n861 B.n418 163.367
R1129 B.n865 B.n418 163.367
R1130 B.n865 B.n412 163.367
R1131 B.n873 B.n412 163.367
R1132 B.n873 B.n410 163.367
R1133 B.n877 B.n410 163.367
R1134 B.n877 B.n404 163.367
R1135 B.n885 B.n404 163.367
R1136 B.n885 B.n402 163.367
R1137 B.n889 B.n402 163.367
R1138 B.n889 B.n396 163.367
R1139 B.n897 B.n396 163.367
R1140 B.n897 B.n394 163.367
R1141 B.n901 B.n394 163.367
R1142 B.n901 B.n388 163.367
R1143 B.n910 B.n388 163.367
R1144 B.n910 B.n386 163.367
R1145 B.n914 B.n386 163.367
R1146 B.n914 B.n3 163.367
R1147 B.n1085 B.n3 163.367
R1148 B.n1081 B.n2 163.367
R1149 B.n1081 B.n1080 163.367
R1150 B.n1080 B.n9 163.367
R1151 B.n1076 B.n9 163.367
R1152 B.n1076 B.n11 163.367
R1153 B.n1072 B.n11 163.367
R1154 B.n1072 B.n17 163.367
R1155 B.n1068 B.n17 163.367
R1156 B.n1068 B.n19 163.367
R1157 B.n1064 B.n19 163.367
R1158 B.n1064 B.n24 163.367
R1159 B.n1060 B.n24 163.367
R1160 B.n1060 B.n26 163.367
R1161 B.n1056 B.n26 163.367
R1162 B.n1056 B.n31 163.367
R1163 B.n1052 B.n31 163.367
R1164 B.n1052 B.n33 163.367
R1165 B.n1048 B.n33 163.367
R1166 B.n1048 B.n38 163.367
R1167 B.n1044 B.n38 163.367
R1168 B.n1044 B.n40 163.367
R1169 B.n1040 B.n40 163.367
R1170 B.n1040 B.n45 163.367
R1171 B.n1036 B.n45 163.367
R1172 B.n1036 B.n47 163.367
R1173 B.n1032 B.n47 163.367
R1174 B.n1032 B.n52 163.367
R1175 B.n1028 B.n52 163.367
R1176 B.n1028 B.n54 163.367
R1177 B.n1024 B.n54 163.367
R1178 B.n1024 B.n58 163.367
R1179 B.n1020 B.n58 163.367
R1180 B.n1020 B.n60 163.367
R1181 B.n1016 B.n60 163.367
R1182 B.n1016 B.n66 163.367
R1183 B.n1012 B.n66 163.367
R1184 B.n1012 B.n68 163.367
R1185 B.n1008 B.n68 163.367
R1186 B.n1008 B.n73 163.367
R1187 B.n1004 B.n73 163.367
R1188 B.n1004 B.n75 163.367
R1189 B.n1000 B.n75 163.367
R1190 B.n1000 B.n80 163.367
R1191 B.n996 B.n80 163.367
R1192 B.n996 B.n82 163.367
R1193 B.n992 B.n82 163.367
R1194 B.n992 B.n87 163.367
R1195 B.n988 B.n87 163.367
R1196 B.n988 B.n89 163.367
R1197 B.n150 B.t10 124.032
R1198 B.n540 B.t15 124.032
R1199 B.n153 B.t17 124.013
R1200 B.n537 B.t21 124.013
R1201 B.n155 B.n92 71.676
R1202 B.n159 B.n93 71.676
R1203 B.n163 B.n94 71.676
R1204 B.n167 B.n95 71.676
R1205 B.n171 B.n96 71.676
R1206 B.n175 B.n97 71.676
R1207 B.n179 B.n98 71.676
R1208 B.n183 B.n99 71.676
R1209 B.n187 B.n100 71.676
R1210 B.n191 B.n101 71.676
R1211 B.n195 B.n102 71.676
R1212 B.n199 B.n103 71.676
R1213 B.n203 B.n104 71.676
R1214 B.n207 B.n105 71.676
R1215 B.n211 B.n106 71.676
R1216 B.n215 B.n107 71.676
R1217 B.n219 B.n108 71.676
R1218 B.n223 B.n109 71.676
R1219 B.n227 B.n110 71.676
R1220 B.n231 B.n111 71.676
R1221 B.n235 B.n112 71.676
R1222 B.n239 B.n113 71.676
R1223 B.n243 B.n114 71.676
R1224 B.n247 B.n115 71.676
R1225 B.n251 B.n116 71.676
R1226 B.n255 B.n117 71.676
R1227 B.n259 B.n118 71.676
R1228 B.n264 B.n119 71.676
R1229 B.n268 B.n120 71.676
R1230 B.n272 B.n121 71.676
R1231 B.n276 B.n122 71.676
R1232 B.n280 B.n123 71.676
R1233 B.n284 B.n124 71.676
R1234 B.n288 B.n125 71.676
R1235 B.n292 B.n126 71.676
R1236 B.n296 B.n127 71.676
R1237 B.n300 B.n128 71.676
R1238 B.n304 B.n129 71.676
R1239 B.n308 B.n130 71.676
R1240 B.n312 B.n131 71.676
R1241 B.n316 B.n132 71.676
R1242 B.n320 B.n133 71.676
R1243 B.n324 B.n134 71.676
R1244 B.n328 B.n135 71.676
R1245 B.n332 B.n136 71.676
R1246 B.n336 B.n137 71.676
R1247 B.n340 B.n138 71.676
R1248 B.n344 B.n139 71.676
R1249 B.n348 B.n140 71.676
R1250 B.n352 B.n141 71.676
R1251 B.n356 B.n142 71.676
R1252 B.n360 B.n143 71.676
R1253 B.n364 B.n144 71.676
R1254 B.n368 B.n145 71.676
R1255 B.n372 B.n146 71.676
R1256 B.n376 B.n147 71.676
R1257 B.n380 B.n148 71.676
R1258 B.n149 B.n148 71.676
R1259 B.n379 B.n147 71.676
R1260 B.n375 B.n146 71.676
R1261 B.n371 B.n145 71.676
R1262 B.n367 B.n144 71.676
R1263 B.n363 B.n143 71.676
R1264 B.n359 B.n142 71.676
R1265 B.n355 B.n141 71.676
R1266 B.n351 B.n140 71.676
R1267 B.n347 B.n139 71.676
R1268 B.n343 B.n138 71.676
R1269 B.n339 B.n137 71.676
R1270 B.n335 B.n136 71.676
R1271 B.n331 B.n135 71.676
R1272 B.n327 B.n134 71.676
R1273 B.n323 B.n133 71.676
R1274 B.n319 B.n132 71.676
R1275 B.n315 B.n131 71.676
R1276 B.n311 B.n130 71.676
R1277 B.n307 B.n129 71.676
R1278 B.n303 B.n128 71.676
R1279 B.n299 B.n127 71.676
R1280 B.n295 B.n126 71.676
R1281 B.n291 B.n125 71.676
R1282 B.n287 B.n124 71.676
R1283 B.n283 B.n123 71.676
R1284 B.n279 B.n122 71.676
R1285 B.n275 B.n121 71.676
R1286 B.n271 B.n120 71.676
R1287 B.n267 B.n119 71.676
R1288 B.n263 B.n118 71.676
R1289 B.n258 B.n117 71.676
R1290 B.n254 B.n116 71.676
R1291 B.n250 B.n115 71.676
R1292 B.n246 B.n114 71.676
R1293 B.n242 B.n113 71.676
R1294 B.n238 B.n112 71.676
R1295 B.n234 B.n111 71.676
R1296 B.n230 B.n110 71.676
R1297 B.n226 B.n109 71.676
R1298 B.n222 B.n108 71.676
R1299 B.n218 B.n107 71.676
R1300 B.n214 B.n106 71.676
R1301 B.n210 B.n105 71.676
R1302 B.n206 B.n104 71.676
R1303 B.n202 B.n103 71.676
R1304 B.n198 B.n102 71.676
R1305 B.n194 B.n101 71.676
R1306 B.n190 B.n100 71.676
R1307 B.n186 B.n99 71.676
R1308 B.n182 B.n98 71.676
R1309 B.n178 B.n97 71.676
R1310 B.n174 B.n96 71.676
R1311 B.n170 B.n95 71.676
R1312 B.n166 B.n94 71.676
R1313 B.n162 B.n93 71.676
R1314 B.n158 B.n92 71.676
R1315 B.n767 B.n766 71.676
R1316 B.n761 B.n480 71.676
R1317 B.n758 B.n481 71.676
R1318 B.n754 B.n482 71.676
R1319 B.n750 B.n483 71.676
R1320 B.n746 B.n484 71.676
R1321 B.n742 B.n485 71.676
R1322 B.n738 B.n486 71.676
R1323 B.n734 B.n487 71.676
R1324 B.n730 B.n488 71.676
R1325 B.n726 B.n489 71.676
R1326 B.n722 B.n490 71.676
R1327 B.n718 B.n491 71.676
R1328 B.n714 B.n492 71.676
R1329 B.n710 B.n493 71.676
R1330 B.n706 B.n494 71.676
R1331 B.n702 B.n495 71.676
R1332 B.n698 B.n496 71.676
R1333 B.n694 B.n497 71.676
R1334 B.n690 B.n498 71.676
R1335 B.n686 B.n499 71.676
R1336 B.n682 B.n500 71.676
R1337 B.n678 B.n501 71.676
R1338 B.n674 B.n502 71.676
R1339 B.n670 B.n503 71.676
R1340 B.n666 B.n504 71.676
R1341 B.n662 B.n505 71.676
R1342 B.n658 B.n506 71.676
R1343 B.n654 B.n507 71.676
R1344 B.n650 B.n508 71.676
R1345 B.n646 B.n509 71.676
R1346 B.n641 B.n510 71.676
R1347 B.n637 B.n511 71.676
R1348 B.n633 B.n512 71.676
R1349 B.n629 B.n513 71.676
R1350 B.n625 B.n514 71.676
R1351 B.n621 B.n515 71.676
R1352 B.n617 B.n516 71.676
R1353 B.n613 B.n517 71.676
R1354 B.n609 B.n518 71.676
R1355 B.n605 B.n519 71.676
R1356 B.n601 B.n520 71.676
R1357 B.n597 B.n521 71.676
R1358 B.n593 B.n522 71.676
R1359 B.n589 B.n523 71.676
R1360 B.n585 B.n524 71.676
R1361 B.n581 B.n525 71.676
R1362 B.n577 B.n526 71.676
R1363 B.n573 B.n527 71.676
R1364 B.n569 B.n528 71.676
R1365 B.n565 B.n529 71.676
R1366 B.n561 B.n530 71.676
R1367 B.n557 B.n531 71.676
R1368 B.n553 B.n532 71.676
R1369 B.n549 B.n533 71.676
R1370 B.n545 B.n534 71.676
R1371 B.n769 B.n479 71.676
R1372 B.n767 B.n536 71.676
R1373 B.n759 B.n480 71.676
R1374 B.n755 B.n481 71.676
R1375 B.n751 B.n482 71.676
R1376 B.n747 B.n483 71.676
R1377 B.n743 B.n484 71.676
R1378 B.n739 B.n485 71.676
R1379 B.n735 B.n486 71.676
R1380 B.n731 B.n487 71.676
R1381 B.n727 B.n488 71.676
R1382 B.n723 B.n489 71.676
R1383 B.n719 B.n490 71.676
R1384 B.n715 B.n491 71.676
R1385 B.n711 B.n492 71.676
R1386 B.n707 B.n493 71.676
R1387 B.n703 B.n494 71.676
R1388 B.n699 B.n495 71.676
R1389 B.n695 B.n496 71.676
R1390 B.n691 B.n497 71.676
R1391 B.n687 B.n498 71.676
R1392 B.n683 B.n499 71.676
R1393 B.n679 B.n500 71.676
R1394 B.n675 B.n501 71.676
R1395 B.n671 B.n502 71.676
R1396 B.n667 B.n503 71.676
R1397 B.n663 B.n504 71.676
R1398 B.n659 B.n505 71.676
R1399 B.n655 B.n506 71.676
R1400 B.n651 B.n507 71.676
R1401 B.n647 B.n508 71.676
R1402 B.n642 B.n509 71.676
R1403 B.n638 B.n510 71.676
R1404 B.n634 B.n511 71.676
R1405 B.n630 B.n512 71.676
R1406 B.n626 B.n513 71.676
R1407 B.n622 B.n514 71.676
R1408 B.n618 B.n515 71.676
R1409 B.n614 B.n516 71.676
R1410 B.n610 B.n517 71.676
R1411 B.n606 B.n518 71.676
R1412 B.n602 B.n519 71.676
R1413 B.n598 B.n520 71.676
R1414 B.n594 B.n521 71.676
R1415 B.n590 B.n522 71.676
R1416 B.n586 B.n523 71.676
R1417 B.n582 B.n524 71.676
R1418 B.n578 B.n525 71.676
R1419 B.n574 B.n526 71.676
R1420 B.n570 B.n527 71.676
R1421 B.n566 B.n528 71.676
R1422 B.n562 B.n529 71.676
R1423 B.n558 B.n530 71.676
R1424 B.n554 B.n531 71.676
R1425 B.n550 B.n532 71.676
R1426 B.n546 B.n533 71.676
R1427 B.n542 B.n534 71.676
R1428 B.n770 B.n769 71.676
R1429 B.n1086 B.n1085 71.676
R1430 B.n1086 B.n2 71.676
R1431 B.n151 B.t11 69.5359
R1432 B.n541 B.t14 69.5359
R1433 B.n154 B.t18 69.5151
R1434 B.n538 B.t20 69.5151
R1435 B.n768 B.n476 62.2597
R1436 B.n986 B.n985 62.2597
R1437 B.n261 B.n154 59.5399
R1438 B.n152 B.n151 59.5399
R1439 B.n644 B.n541 59.5399
R1440 B.n539 B.n538 59.5399
R1441 B.n154 B.n153 54.4975
R1442 B.n151 B.n150 54.4975
R1443 B.n541 B.n540 54.4975
R1444 B.n538 B.n537 54.4975
R1445 B.n775 B.n476 35.5772
R1446 B.n775 B.n472 35.5772
R1447 B.n781 B.n472 35.5772
R1448 B.n781 B.n468 35.5772
R1449 B.n787 B.n468 35.5772
R1450 B.n787 B.n464 35.5772
R1451 B.n793 B.n464 35.5772
R1452 B.n799 B.n460 35.5772
R1453 B.n799 B.n456 35.5772
R1454 B.n805 B.n456 35.5772
R1455 B.n805 B.n452 35.5772
R1456 B.n811 B.n452 35.5772
R1457 B.n811 B.n448 35.5772
R1458 B.n817 B.n448 35.5772
R1459 B.n817 B.n444 35.5772
R1460 B.n824 B.n444 35.5772
R1461 B.n824 B.n823 35.5772
R1462 B.n830 B.n437 35.5772
R1463 B.n836 B.n437 35.5772
R1464 B.n836 B.n433 35.5772
R1465 B.n842 B.n433 35.5772
R1466 B.n842 B.n429 35.5772
R1467 B.n848 B.n429 35.5772
R1468 B.n848 B.n425 35.5772
R1469 B.n854 B.n425 35.5772
R1470 B.n860 B.n421 35.5772
R1471 B.n860 B.n417 35.5772
R1472 B.n866 B.n417 35.5772
R1473 B.n866 B.n413 35.5772
R1474 B.n872 B.n413 35.5772
R1475 B.n872 B.n409 35.5772
R1476 B.n878 B.n409 35.5772
R1477 B.n884 B.n405 35.5772
R1478 B.n884 B.n401 35.5772
R1479 B.n890 B.n401 35.5772
R1480 B.n890 B.n397 35.5772
R1481 B.n896 B.n397 35.5772
R1482 B.n896 B.n393 35.5772
R1483 B.n902 B.n393 35.5772
R1484 B.n909 B.n389 35.5772
R1485 B.n909 B.n385 35.5772
R1486 B.n915 B.n385 35.5772
R1487 B.n915 B.n4 35.5772
R1488 B.n1084 B.n4 35.5772
R1489 B.n1084 B.n1083 35.5772
R1490 B.n1083 B.n1082 35.5772
R1491 B.n1082 B.n8 35.5772
R1492 B.n12 B.n8 35.5772
R1493 B.n1075 B.n12 35.5772
R1494 B.n1075 B.n1074 35.5772
R1495 B.n1073 B.n16 35.5772
R1496 B.n1067 B.n16 35.5772
R1497 B.n1067 B.n1066 35.5772
R1498 B.n1066 B.n1065 35.5772
R1499 B.n1065 B.n23 35.5772
R1500 B.n1059 B.n23 35.5772
R1501 B.n1059 B.n1058 35.5772
R1502 B.n1057 B.n30 35.5772
R1503 B.n1051 B.n30 35.5772
R1504 B.n1051 B.n1050 35.5772
R1505 B.n1050 B.n1049 35.5772
R1506 B.n1049 B.n37 35.5772
R1507 B.n1043 B.n37 35.5772
R1508 B.n1043 B.n1042 35.5772
R1509 B.n1041 B.n44 35.5772
R1510 B.n1035 B.n44 35.5772
R1511 B.n1035 B.n1034 35.5772
R1512 B.n1034 B.n1033 35.5772
R1513 B.n1033 B.n51 35.5772
R1514 B.n1027 B.n51 35.5772
R1515 B.n1027 B.n1026 35.5772
R1516 B.n1026 B.n1025 35.5772
R1517 B.n1019 B.n61 35.5772
R1518 B.n1019 B.n1018 35.5772
R1519 B.n1018 B.n1017 35.5772
R1520 B.n1017 B.n65 35.5772
R1521 B.n1011 B.n65 35.5772
R1522 B.n1011 B.n1010 35.5772
R1523 B.n1010 B.n1009 35.5772
R1524 B.n1009 B.n72 35.5772
R1525 B.n1003 B.n72 35.5772
R1526 B.n1003 B.n1002 35.5772
R1527 B.n1001 B.n79 35.5772
R1528 B.n995 B.n79 35.5772
R1529 B.n995 B.n994 35.5772
R1530 B.n994 B.n993 35.5772
R1531 B.n993 B.n86 35.5772
R1532 B.n987 B.n86 35.5772
R1533 B.n987 B.n986 35.5772
R1534 B.n823 B.t1 34.5308
R1535 B.n61 B.t6 34.5308
R1536 B.n765 B.n474 31.0639
R1537 B.n772 B.n771 31.0639
R1538 B.n983 B.n982 31.0639
R1539 B.n156 B.n88 31.0639
R1540 B.t4 B.n421 27.2062
R1541 B.n902 B.t2 27.2062
R1542 B.t5 B.n1073 27.2062
R1543 B.n1042 B.t7 27.2062
R1544 B B.n1087 18.0485
R1545 B.n793 B.t13 17.7888
R1546 B.t13 B.n460 17.7888
R1547 B.n878 B.t0 17.7888
R1548 B.t0 B.n405 17.7888
R1549 B.n1058 B.t3 17.7888
R1550 B.t3 B.n1057 17.7888
R1551 B.n1002 B.t9 17.7888
R1552 B.t9 B.n1001 17.7888
R1553 B.n777 B.n474 10.6151
R1554 B.n778 B.n777 10.6151
R1555 B.n779 B.n778 10.6151
R1556 B.n779 B.n466 10.6151
R1557 B.n789 B.n466 10.6151
R1558 B.n790 B.n789 10.6151
R1559 B.n791 B.n790 10.6151
R1560 B.n791 B.n458 10.6151
R1561 B.n801 B.n458 10.6151
R1562 B.n802 B.n801 10.6151
R1563 B.n803 B.n802 10.6151
R1564 B.n803 B.n450 10.6151
R1565 B.n813 B.n450 10.6151
R1566 B.n814 B.n813 10.6151
R1567 B.n815 B.n814 10.6151
R1568 B.n815 B.n442 10.6151
R1569 B.n826 B.n442 10.6151
R1570 B.n827 B.n826 10.6151
R1571 B.n828 B.n827 10.6151
R1572 B.n828 B.n435 10.6151
R1573 B.n838 B.n435 10.6151
R1574 B.n839 B.n838 10.6151
R1575 B.n840 B.n839 10.6151
R1576 B.n840 B.n427 10.6151
R1577 B.n850 B.n427 10.6151
R1578 B.n851 B.n850 10.6151
R1579 B.n852 B.n851 10.6151
R1580 B.n852 B.n419 10.6151
R1581 B.n862 B.n419 10.6151
R1582 B.n863 B.n862 10.6151
R1583 B.n864 B.n863 10.6151
R1584 B.n864 B.n411 10.6151
R1585 B.n874 B.n411 10.6151
R1586 B.n875 B.n874 10.6151
R1587 B.n876 B.n875 10.6151
R1588 B.n876 B.n403 10.6151
R1589 B.n886 B.n403 10.6151
R1590 B.n887 B.n886 10.6151
R1591 B.n888 B.n887 10.6151
R1592 B.n888 B.n395 10.6151
R1593 B.n898 B.n395 10.6151
R1594 B.n899 B.n898 10.6151
R1595 B.n900 B.n899 10.6151
R1596 B.n900 B.n387 10.6151
R1597 B.n911 B.n387 10.6151
R1598 B.n912 B.n911 10.6151
R1599 B.n913 B.n912 10.6151
R1600 B.n913 B.n0 10.6151
R1601 B.n765 B.n764 10.6151
R1602 B.n764 B.n763 10.6151
R1603 B.n763 B.n762 10.6151
R1604 B.n762 B.n760 10.6151
R1605 B.n760 B.n757 10.6151
R1606 B.n757 B.n756 10.6151
R1607 B.n756 B.n753 10.6151
R1608 B.n753 B.n752 10.6151
R1609 B.n752 B.n749 10.6151
R1610 B.n749 B.n748 10.6151
R1611 B.n748 B.n745 10.6151
R1612 B.n745 B.n744 10.6151
R1613 B.n744 B.n741 10.6151
R1614 B.n741 B.n740 10.6151
R1615 B.n740 B.n737 10.6151
R1616 B.n737 B.n736 10.6151
R1617 B.n736 B.n733 10.6151
R1618 B.n733 B.n732 10.6151
R1619 B.n732 B.n729 10.6151
R1620 B.n729 B.n728 10.6151
R1621 B.n728 B.n725 10.6151
R1622 B.n725 B.n724 10.6151
R1623 B.n724 B.n721 10.6151
R1624 B.n721 B.n720 10.6151
R1625 B.n720 B.n717 10.6151
R1626 B.n717 B.n716 10.6151
R1627 B.n716 B.n713 10.6151
R1628 B.n713 B.n712 10.6151
R1629 B.n712 B.n709 10.6151
R1630 B.n709 B.n708 10.6151
R1631 B.n708 B.n705 10.6151
R1632 B.n705 B.n704 10.6151
R1633 B.n704 B.n701 10.6151
R1634 B.n701 B.n700 10.6151
R1635 B.n700 B.n697 10.6151
R1636 B.n697 B.n696 10.6151
R1637 B.n696 B.n693 10.6151
R1638 B.n693 B.n692 10.6151
R1639 B.n692 B.n689 10.6151
R1640 B.n689 B.n688 10.6151
R1641 B.n688 B.n685 10.6151
R1642 B.n685 B.n684 10.6151
R1643 B.n684 B.n681 10.6151
R1644 B.n681 B.n680 10.6151
R1645 B.n680 B.n677 10.6151
R1646 B.n677 B.n676 10.6151
R1647 B.n676 B.n673 10.6151
R1648 B.n673 B.n672 10.6151
R1649 B.n672 B.n669 10.6151
R1650 B.n669 B.n668 10.6151
R1651 B.n668 B.n665 10.6151
R1652 B.n665 B.n664 10.6151
R1653 B.n661 B.n660 10.6151
R1654 B.n660 B.n657 10.6151
R1655 B.n657 B.n656 10.6151
R1656 B.n656 B.n653 10.6151
R1657 B.n653 B.n652 10.6151
R1658 B.n652 B.n649 10.6151
R1659 B.n649 B.n648 10.6151
R1660 B.n648 B.n645 10.6151
R1661 B.n643 B.n640 10.6151
R1662 B.n640 B.n639 10.6151
R1663 B.n639 B.n636 10.6151
R1664 B.n636 B.n635 10.6151
R1665 B.n635 B.n632 10.6151
R1666 B.n632 B.n631 10.6151
R1667 B.n631 B.n628 10.6151
R1668 B.n628 B.n627 10.6151
R1669 B.n627 B.n624 10.6151
R1670 B.n624 B.n623 10.6151
R1671 B.n623 B.n620 10.6151
R1672 B.n620 B.n619 10.6151
R1673 B.n619 B.n616 10.6151
R1674 B.n616 B.n615 10.6151
R1675 B.n615 B.n612 10.6151
R1676 B.n612 B.n611 10.6151
R1677 B.n611 B.n608 10.6151
R1678 B.n608 B.n607 10.6151
R1679 B.n607 B.n604 10.6151
R1680 B.n604 B.n603 10.6151
R1681 B.n603 B.n600 10.6151
R1682 B.n600 B.n599 10.6151
R1683 B.n599 B.n596 10.6151
R1684 B.n596 B.n595 10.6151
R1685 B.n595 B.n592 10.6151
R1686 B.n592 B.n591 10.6151
R1687 B.n591 B.n588 10.6151
R1688 B.n588 B.n587 10.6151
R1689 B.n587 B.n584 10.6151
R1690 B.n584 B.n583 10.6151
R1691 B.n583 B.n580 10.6151
R1692 B.n580 B.n579 10.6151
R1693 B.n579 B.n576 10.6151
R1694 B.n576 B.n575 10.6151
R1695 B.n575 B.n572 10.6151
R1696 B.n572 B.n571 10.6151
R1697 B.n571 B.n568 10.6151
R1698 B.n568 B.n567 10.6151
R1699 B.n567 B.n564 10.6151
R1700 B.n564 B.n563 10.6151
R1701 B.n563 B.n560 10.6151
R1702 B.n560 B.n559 10.6151
R1703 B.n559 B.n556 10.6151
R1704 B.n556 B.n555 10.6151
R1705 B.n555 B.n552 10.6151
R1706 B.n552 B.n551 10.6151
R1707 B.n551 B.n548 10.6151
R1708 B.n548 B.n547 10.6151
R1709 B.n547 B.n544 10.6151
R1710 B.n544 B.n543 10.6151
R1711 B.n543 B.n478 10.6151
R1712 B.n771 B.n478 10.6151
R1713 B.n773 B.n772 10.6151
R1714 B.n773 B.n470 10.6151
R1715 B.n783 B.n470 10.6151
R1716 B.n784 B.n783 10.6151
R1717 B.n785 B.n784 10.6151
R1718 B.n785 B.n462 10.6151
R1719 B.n795 B.n462 10.6151
R1720 B.n796 B.n795 10.6151
R1721 B.n797 B.n796 10.6151
R1722 B.n797 B.n454 10.6151
R1723 B.n807 B.n454 10.6151
R1724 B.n808 B.n807 10.6151
R1725 B.n809 B.n808 10.6151
R1726 B.n809 B.n446 10.6151
R1727 B.n819 B.n446 10.6151
R1728 B.n820 B.n819 10.6151
R1729 B.n821 B.n820 10.6151
R1730 B.n821 B.n439 10.6151
R1731 B.n832 B.n439 10.6151
R1732 B.n833 B.n832 10.6151
R1733 B.n834 B.n833 10.6151
R1734 B.n834 B.n431 10.6151
R1735 B.n844 B.n431 10.6151
R1736 B.n845 B.n844 10.6151
R1737 B.n846 B.n845 10.6151
R1738 B.n846 B.n423 10.6151
R1739 B.n856 B.n423 10.6151
R1740 B.n857 B.n856 10.6151
R1741 B.n858 B.n857 10.6151
R1742 B.n858 B.n415 10.6151
R1743 B.n868 B.n415 10.6151
R1744 B.n869 B.n868 10.6151
R1745 B.n870 B.n869 10.6151
R1746 B.n870 B.n407 10.6151
R1747 B.n880 B.n407 10.6151
R1748 B.n881 B.n880 10.6151
R1749 B.n882 B.n881 10.6151
R1750 B.n882 B.n399 10.6151
R1751 B.n892 B.n399 10.6151
R1752 B.n893 B.n892 10.6151
R1753 B.n894 B.n893 10.6151
R1754 B.n894 B.n391 10.6151
R1755 B.n904 B.n391 10.6151
R1756 B.n905 B.n904 10.6151
R1757 B.n907 B.n905 10.6151
R1758 B.n907 B.n906 10.6151
R1759 B.n906 B.n383 10.6151
R1760 B.n918 B.n383 10.6151
R1761 B.n919 B.n918 10.6151
R1762 B.n920 B.n919 10.6151
R1763 B.n921 B.n920 10.6151
R1764 B.n922 B.n921 10.6151
R1765 B.n925 B.n922 10.6151
R1766 B.n926 B.n925 10.6151
R1767 B.n927 B.n926 10.6151
R1768 B.n928 B.n927 10.6151
R1769 B.n930 B.n928 10.6151
R1770 B.n931 B.n930 10.6151
R1771 B.n932 B.n931 10.6151
R1772 B.n933 B.n932 10.6151
R1773 B.n935 B.n933 10.6151
R1774 B.n936 B.n935 10.6151
R1775 B.n937 B.n936 10.6151
R1776 B.n938 B.n937 10.6151
R1777 B.n940 B.n938 10.6151
R1778 B.n941 B.n940 10.6151
R1779 B.n942 B.n941 10.6151
R1780 B.n943 B.n942 10.6151
R1781 B.n945 B.n943 10.6151
R1782 B.n946 B.n945 10.6151
R1783 B.n947 B.n946 10.6151
R1784 B.n948 B.n947 10.6151
R1785 B.n950 B.n948 10.6151
R1786 B.n951 B.n950 10.6151
R1787 B.n952 B.n951 10.6151
R1788 B.n953 B.n952 10.6151
R1789 B.n955 B.n953 10.6151
R1790 B.n956 B.n955 10.6151
R1791 B.n957 B.n956 10.6151
R1792 B.n958 B.n957 10.6151
R1793 B.n960 B.n958 10.6151
R1794 B.n961 B.n960 10.6151
R1795 B.n962 B.n961 10.6151
R1796 B.n963 B.n962 10.6151
R1797 B.n965 B.n963 10.6151
R1798 B.n966 B.n965 10.6151
R1799 B.n967 B.n966 10.6151
R1800 B.n968 B.n967 10.6151
R1801 B.n970 B.n968 10.6151
R1802 B.n971 B.n970 10.6151
R1803 B.n972 B.n971 10.6151
R1804 B.n973 B.n972 10.6151
R1805 B.n975 B.n973 10.6151
R1806 B.n976 B.n975 10.6151
R1807 B.n977 B.n976 10.6151
R1808 B.n978 B.n977 10.6151
R1809 B.n980 B.n978 10.6151
R1810 B.n981 B.n980 10.6151
R1811 B.n982 B.n981 10.6151
R1812 B.n1079 B.n1 10.6151
R1813 B.n1079 B.n1078 10.6151
R1814 B.n1078 B.n1077 10.6151
R1815 B.n1077 B.n10 10.6151
R1816 B.n1071 B.n10 10.6151
R1817 B.n1071 B.n1070 10.6151
R1818 B.n1070 B.n1069 10.6151
R1819 B.n1069 B.n18 10.6151
R1820 B.n1063 B.n18 10.6151
R1821 B.n1063 B.n1062 10.6151
R1822 B.n1062 B.n1061 10.6151
R1823 B.n1061 B.n25 10.6151
R1824 B.n1055 B.n25 10.6151
R1825 B.n1055 B.n1054 10.6151
R1826 B.n1054 B.n1053 10.6151
R1827 B.n1053 B.n32 10.6151
R1828 B.n1047 B.n32 10.6151
R1829 B.n1047 B.n1046 10.6151
R1830 B.n1046 B.n1045 10.6151
R1831 B.n1045 B.n39 10.6151
R1832 B.n1039 B.n39 10.6151
R1833 B.n1039 B.n1038 10.6151
R1834 B.n1038 B.n1037 10.6151
R1835 B.n1037 B.n46 10.6151
R1836 B.n1031 B.n46 10.6151
R1837 B.n1031 B.n1030 10.6151
R1838 B.n1030 B.n1029 10.6151
R1839 B.n1029 B.n53 10.6151
R1840 B.n1023 B.n53 10.6151
R1841 B.n1023 B.n1022 10.6151
R1842 B.n1022 B.n1021 10.6151
R1843 B.n1021 B.n59 10.6151
R1844 B.n1015 B.n59 10.6151
R1845 B.n1015 B.n1014 10.6151
R1846 B.n1014 B.n1013 10.6151
R1847 B.n1013 B.n67 10.6151
R1848 B.n1007 B.n67 10.6151
R1849 B.n1007 B.n1006 10.6151
R1850 B.n1006 B.n1005 10.6151
R1851 B.n1005 B.n74 10.6151
R1852 B.n999 B.n74 10.6151
R1853 B.n999 B.n998 10.6151
R1854 B.n998 B.n997 10.6151
R1855 B.n997 B.n81 10.6151
R1856 B.n991 B.n81 10.6151
R1857 B.n991 B.n990 10.6151
R1858 B.n990 B.n989 10.6151
R1859 B.n989 B.n88 10.6151
R1860 B.n157 B.n156 10.6151
R1861 B.n160 B.n157 10.6151
R1862 B.n161 B.n160 10.6151
R1863 B.n164 B.n161 10.6151
R1864 B.n165 B.n164 10.6151
R1865 B.n168 B.n165 10.6151
R1866 B.n169 B.n168 10.6151
R1867 B.n172 B.n169 10.6151
R1868 B.n173 B.n172 10.6151
R1869 B.n176 B.n173 10.6151
R1870 B.n177 B.n176 10.6151
R1871 B.n180 B.n177 10.6151
R1872 B.n181 B.n180 10.6151
R1873 B.n184 B.n181 10.6151
R1874 B.n185 B.n184 10.6151
R1875 B.n188 B.n185 10.6151
R1876 B.n189 B.n188 10.6151
R1877 B.n192 B.n189 10.6151
R1878 B.n193 B.n192 10.6151
R1879 B.n196 B.n193 10.6151
R1880 B.n197 B.n196 10.6151
R1881 B.n200 B.n197 10.6151
R1882 B.n201 B.n200 10.6151
R1883 B.n204 B.n201 10.6151
R1884 B.n205 B.n204 10.6151
R1885 B.n208 B.n205 10.6151
R1886 B.n209 B.n208 10.6151
R1887 B.n212 B.n209 10.6151
R1888 B.n213 B.n212 10.6151
R1889 B.n216 B.n213 10.6151
R1890 B.n217 B.n216 10.6151
R1891 B.n220 B.n217 10.6151
R1892 B.n221 B.n220 10.6151
R1893 B.n224 B.n221 10.6151
R1894 B.n225 B.n224 10.6151
R1895 B.n228 B.n225 10.6151
R1896 B.n229 B.n228 10.6151
R1897 B.n232 B.n229 10.6151
R1898 B.n233 B.n232 10.6151
R1899 B.n236 B.n233 10.6151
R1900 B.n237 B.n236 10.6151
R1901 B.n240 B.n237 10.6151
R1902 B.n241 B.n240 10.6151
R1903 B.n244 B.n241 10.6151
R1904 B.n245 B.n244 10.6151
R1905 B.n248 B.n245 10.6151
R1906 B.n249 B.n248 10.6151
R1907 B.n252 B.n249 10.6151
R1908 B.n253 B.n252 10.6151
R1909 B.n256 B.n253 10.6151
R1910 B.n257 B.n256 10.6151
R1911 B.n260 B.n257 10.6151
R1912 B.n265 B.n262 10.6151
R1913 B.n266 B.n265 10.6151
R1914 B.n269 B.n266 10.6151
R1915 B.n270 B.n269 10.6151
R1916 B.n273 B.n270 10.6151
R1917 B.n274 B.n273 10.6151
R1918 B.n277 B.n274 10.6151
R1919 B.n278 B.n277 10.6151
R1920 B.n282 B.n281 10.6151
R1921 B.n285 B.n282 10.6151
R1922 B.n286 B.n285 10.6151
R1923 B.n289 B.n286 10.6151
R1924 B.n290 B.n289 10.6151
R1925 B.n293 B.n290 10.6151
R1926 B.n294 B.n293 10.6151
R1927 B.n297 B.n294 10.6151
R1928 B.n298 B.n297 10.6151
R1929 B.n301 B.n298 10.6151
R1930 B.n302 B.n301 10.6151
R1931 B.n305 B.n302 10.6151
R1932 B.n306 B.n305 10.6151
R1933 B.n309 B.n306 10.6151
R1934 B.n310 B.n309 10.6151
R1935 B.n313 B.n310 10.6151
R1936 B.n314 B.n313 10.6151
R1937 B.n317 B.n314 10.6151
R1938 B.n318 B.n317 10.6151
R1939 B.n321 B.n318 10.6151
R1940 B.n322 B.n321 10.6151
R1941 B.n325 B.n322 10.6151
R1942 B.n326 B.n325 10.6151
R1943 B.n329 B.n326 10.6151
R1944 B.n330 B.n329 10.6151
R1945 B.n333 B.n330 10.6151
R1946 B.n334 B.n333 10.6151
R1947 B.n337 B.n334 10.6151
R1948 B.n338 B.n337 10.6151
R1949 B.n341 B.n338 10.6151
R1950 B.n342 B.n341 10.6151
R1951 B.n345 B.n342 10.6151
R1952 B.n346 B.n345 10.6151
R1953 B.n349 B.n346 10.6151
R1954 B.n350 B.n349 10.6151
R1955 B.n353 B.n350 10.6151
R1956 B.n354 B.n353 10.6151
R1957 B.n357 B.n354 10.6151
R1958 B.n358 B.n357 10.6151
R1959 B.n361 B.n358 10.6151
R1960 B.n362 B.n361 10.6151
R1961 B.n365 B.n362 10.6151
R1962 B.n366 B.n365 10.6151
R1963 B.n369 B.n366 10.6151
R1964 B.n370 B.n369 10.6151
R1965 B.n373 B.n370 10.6151
R1966 B.n374 B.n373 10.6151
R1967 B.n377 B.n374 10.6151
R1968 B.n378 B.n377 10.6151
R1969 B.n381 B.n378 10.6151
R1970 B.n382 B.n381 10.6151
R1971 B.n983 B.n382 10.6151
R1972 B.n854 B.t4 8.37149
R1973 B.t2 B.n389 8.37149
R1974 B.n1074 B.t5 8.37149
R1975 B.t7 B.n1041 8.37149
R1976 B.n1087 B.n0 8.11757
R1977 B.n1087 B.n1 8.11757
R1978 B.n661 B.n539 6.5566
R1979 B.n645 B.n644 6.5566
R1980 B.n262 B.n261 6.5566
R1981 B.n278 B.n152 6.5566
R1982 B.n664 B.n539 4.05904
R1983 B.n644 B.n643 4.05904
R1984 B.n261 B.n260 4.05904
R1985 B.n281 B.n152 4.05904
R1986 B.n830 B.t1 1.04687
R1987 B.n1025 B.t6 1.04687
R1988 VP.n16 VP.t2 186.806
R1989 VP.n19 VP.n18 161.3
R1990 VP.n20 VP.n15 161.3
R1991 VP.n22 VP.n21 161.3
R1992 VP.n23 VP.n14 161.3
R1993 VP.n25 VP.n24 161.3
R1994 VP.n27 VP.n26 161.3
R1995 VP.n28 VP.n12 161.3
R1996 VP.n30 VP.n29 161.3
R1997 VP.n31 VP.n11 161.3
R1998 VP.n33 VP.n32 161.3
R1999 VP.n34 VP.n10 161.3
R2000 VP.n64 VP.n0 161.3
R2001 VP.n63 VP.n62 161.3
R2002 VP.n61 VP.n1 161.3
R2003 VP.n60 VP.n59 161.3
R2004 VP.n58 VP.n2 161.3
R2005 VP.n57 VP.n56 161.3
R2006 VP.n55 VP.n54 161.3
R2007 VP.n53 VP.n4 161.3
R2008 VP.n52 VP.n51 161.3
R2009 VP.n50 VP.n5 161.3
R2010 VP.n49 VP.n48 161.3
R2011 VP.n46 VP.n6 161.3
R2012 VP.n45 VP.n44 161.3
R2013 VP.n43 VP.n7 161.3
R2014 VP.n42 VP.n41 161.3
R2015 VP.n40 VP.n8 161.3
R2016 VP.n39 VP.n38 161.3
R2017 VP.n9 VP.t6 153.054
R2018 VP.n47 VP.t0 153.054
R2019 VP.n3 VP.t5 153.054
R2020 VP.n65 VP.t7 153.054
R2021 VP.n35 VP.t3 153.054
R2022 VP.n13 VP.t1 153.054
R2023 VP.n17 VP.t4 153.054
R2024 VP.n37 VP.n9 100.236
R2025 VP.n66 VP.n65 100.236
R2026 VP.n36 VP.n35 100.236
R2027 VP.n41 VP.n7 56.5193
R2028 VP.n59 VP.n1 56.5193
R2029 VP.n29 VP.n11 56.5193
R2030 VP.n37 VP.n36 53.1738
R2031 VP.n17 VP.n16 52.6675
R2032 VP.n52 VP.n5 40.4934
R2033 VP.n53 VP.n52 40.4934
R2034 VP.n23 VP.n22 40.4934
R2035 VP.n22 VP.n15 40.4934
R2036 VP.n40 VP.n39 24.4675
R2037 VP.n41 VP.n40 24.4675
R2038 VP.n45 VP.n7 24.4675
R2039 VP.n46 VP.n45 24.4675
R2040 VP.n48 VP.n5 24.4675
R2041 VP.n54 VP.n53 24.4675
R2042 VP.n58 VP.n57 24.4675
R2043 VP.n59 VP.n58 24.4675
R2044 VP.n63 VP.n1 24.4675
R2045 VP.n64 VP.n63 24.4675
R2046 VP.n33 VP.n11 24.4675
R2047 VP.n34 VP.n33 24.4675
R2048 VP.n24 VP.n23 24.4675
R2049 VP.n28 VP.n27 24.4675
R2050 VP.n29 VP.n28 24.4675
R2051 VP.n18 VP.n15 24.4675
R2052 VP.n48 VP.n47 19.8188
R2053 VP.n54 VP.n3 19.8188
R2054 VP.n24 VP.n13 19.8188
R2055 VP.n18 VP.n17 19.8188
R2056 VP.n39 VP.n9 10.5213
R2057 VP.n65 VP.n64 10.5213
R2058 VP.n35 VP.n34 10.5213
R2059 VP.n19 VP.n16 6.81722
R2060 VP.n47 VP.n46 4.64923
R2061 VP.n57 VP.n3 4.64923
R2062 VP.n27 VP.n13 4.64923
R2063 VP.n36 VP.n10 0.278367
R2064 VP.n38 VP.n37 0.278367
R2065 VP.n66 VP.n0 0.278367
R2066 VP.n20 VP.n19 0.189894
R2067 VP.n21 VP.n20 0.189894
R2068 VP.n21 VP.n14 0.189894
R2069 VP.n25 VP.n14 0.189894
R2070 VP.n26 VP.n25 0.189894
R2071 VP.n26 VP.n12 0.189894
R2072 VP.n30 VP.n12 0.189894
R2073 VP.n31 VP.n30 0.189894
R2074 VP.n32 VP.n31 0.189894
R2075 VP.n32 VP.n10 0.189894
R2076 VP.n38 VP.n8 0.189894
R2077 VP.n42 VP.n8 0.189894
R2078 VP.n43 VP.n42 0.189894
R2079 VP.n44 VP.n43 0.189894
R2080 VP.n44 VP.n6 0.189894
R2081 VP.n49 VP.n6 0.189894
R2082 VP.n50 VP.n49 0.189894
R2083 VP.n51 VP.n50 0.189894
R2084 VP.n51 VP.n4 0.189894
R2085 VP.n55 VP.n4 0.189894
R2086 VP.n56 VP.n55 0.189894
R2087 VP.n56 VP.n2 0.189894
R2088 VP.n60 VP.n2 0.189894
R2089 VP.n61 VP.n60 0.189894
R2090 VP.n62 VP.n61 0.189894
R2091 VP.n62 VP.n0 0.189894
R2092 VP VP.n66 0.153454
R2093 VDD1 VDD1.n0 62.6595
R2094 VDD1.n3 VDD1.n2 62.5457
R2095 VDD1.n3 VDD1.n1 62.5457
R2096 VDD1.n5 VDD1.n4 61.3899
R2097 VDD1.n5 VDD1.n3 48.7768
R2098 VDD1.n4 VDD1.t6 1.25764
R2099 VDD1.n4 VDD1.t4 1.25764
R2100 VDD1.n0 VDD1.t5 1.25764
R2101 VDD1.n0 VDD1.t3 1.25764
R2102 VDD1.n2 VDD1.t2 1.25764
R2103 VDD1.n2 VDD1.t0 1.25764
R2104 VDD1.n1 VDD1.t1 1.25764
R2105 VDD1.n1 VDD1.t7 1.25764
R2106 VDD1 VDD1.n5 1.15352
C0 VDD2 VDD1 1.71564f
C1 VN VP 8.210639f
C2 VDD1 VN 0.151613f
C3 VDD2 VTAIL 9.4081f
C4 VN VTAIL 11.3593f
C5 VDD1 VP 11.5133f
C6 VDD2 VN 11.1592f
C7 VTAIL VP 11.373401f
C8 VDD1 VTAIL 9.35448f
C9 VDD2 VP 0.507003f
C10 VDD2 B 5.522882f
C11 VDD1 B 5.945598f
C12 VTAIL B 12.638032f
C13 VN B 15.36759f
C14 VP B 13.872665f
C15 VDD1.t5 B 0.3066f
C16 VDD1.t3 B 0.3066f
C17 VDD1.n0 B 2.78832f
C18 VDD1.t1 B 0.3066f
C19 VDD1.t7 B 0.3066f
C20 VDD1.n1 B 2.78727f
C21 VDD1.t2 B 0.3066f
C22 VDD1.t0 B 0.3066f
C23 VDD1.n2 B 2.78727f
C24 VDD1.n3 B 3.44309f
C25 VDD1.t6 B 0.3066f
C26 VDD1.t4 B 0.3066f
C27 VDD1.n4 B 2.77809f
C28 VDD1.n5 B 3.17622f
C29 VP.n0 B 0.029601f
C30 VP.t7 B 2.40571f
C31 VP.n1 B 0.029022f
C32 VP.n2 B 0.022452f
C33 VP.t5 B 2.40571f
C34 VP.n3 B 0.839899f
C35 VP.n4 B 0.022452f
C36 VP.n5 B 0.044624f
C37 VP.n6 B 0.022452f
C38 VP.t0 B 2.40571f
C39 VP.n7 B 0.03653f
C40 VP.n8 B 0.022452f
C41 VP.t6 B 2.40571f
C42 VP.n9 B 0.912215f
C43 VP.n10 B 0.029601f
C44 VP.t3 B 2.40571f
C45 VP.n11 B 0.029022f
C46 VP.n12 B 0.022452f
C47 VP.t1 B 2.40571f
C48 VP.n13 B 0.839899f
C49 VP.n14 B 0.022452f
C50 VP.n15 B 0.044624f
C51 VP.t2 B 2.58184f
C52 VP.n16 B 0.883256f
C53 VP.t4 B 2.40571f
C54 VP.n17 B 0.909986f
C55 VP.n18 B 0.037919f
C56 VP.n19 B 0.214339f
C57 VP.n20 B 0.022452f
C58 VP.n21 B 0.022452f
C59 VP.n22 B 0.018151f
C60 VP.n23 B 0.044624f
C61 VP.n24 B 0.037919f
C62 VP.n25 B 0.022452f
C63 VP.n26 B 0.022452f
C64 VP.n27 B 0.02511f
C65 VP.n28 B 0.041845f
C66 VP.n29 B 0.03653f
C67 VP.n30 B 0.022452f
C68 VP.n31 B 0.022452f
C69 VP.n32 B 0.022452f
C70 VP.n33 B 0.041845f
C71 VP.n34 B 0.030069f
C72 VP.n35 B 0.912215f
C73 VP.n36 B 1.36442f
C74 VP.n37 B 1.3796f
C75 VP.n38 B 0.029601f
C76 VP.n39 B 0.030069f
C77 VP.n40 B 0.041845f
C78 VP.n41 B 0.029022f
C79 VP.n42 B 0.022452f
C80 VP.n43 B 0.022452f
C81 VP.n44 B 0.022452f
C82 VP.n45 B 0.041845f
C83 VP.n46 B 0.02511f
C84 VP.n47 B 0.839899f
C85 VP.n48 B 0.037919f
C86 VP.n49 B 0.022452f
C87 VP.n50 B 0.022452f
C88 VP.n51 B 0.022452f
C89 VP.n52 B 0.018151f
C90 VP.n53 B 0.044624f
C91 VP.n54 B 0.037919f
C92 VP.n55 B 0.022452f
C93 VP.n56 B 0.022452f
C94 VP.n57 B 0.02511f
C95 VP.n58 B 0.041845f
C96 VP.n59 B 0.03653f
C97 VP.n60 B 0.022452f
C98 VP.n61 B 0.022452f
C99 VP.n62 B 0.022452f
C100 VP.n63 B 0.041845f
C101 VP.n64 B 0.030069f
C102 VP.n65 B 0.912215f
C103 VP.n66 B 0.035397f
C104 VDD2.t4 B 0.30352f
C105 VDD2.t0 B 0.30352f
C106 VDD2.n0 B 2.75927f
C107 VDD2.t3 B 0.30352f
C108 VDD2.t7 B 0.30352f
C109 VDD2.n1 B 2.75927f
C110 VDD2.n2 B 3.3578f
C111 VDD2.t5 B 0.30352f
C112 VDD2.t1 B 0.30352f
C113 VDD2.n3 B 2.75019f
C114 VDD2.n4 B 3.11409f
C115 VDD2.t6 B 0.30352f
C116 VDD2.t2 B 0.30352f
C117 VDD2.n5 B 2.75923f
C118 VTAIL.t13 B 0.235562f
C119 VTAIL.t8 B 0.235562f
C120 VTAIL.n0 B 2.0779f
C121 VTAIL.n1 B 0.337231f
C122 VTAIL.t9 B 2.65238f
C123 VTAIL.n2 B 0.430297f
C124 VTAIL.t2 B 2.65238f
C125 VTAIL.n3 B 0.430297f
C126 VTAIL.t4 B 0.235562f
C127 VTAIL.t0 B 0.235562f
C128 VTAIL.n4 B 2.0779f
C129 VTAIL.n5 B 0.481415f
C130 VTAIL.t1 B 2.65238f
C131 VTAIL.n6 B 1.63451f
C132 VTAIL.t14 B 2.6524f
C133 VTAIL.n7 B 1.63449f
C134 VTAIL.t10 B 0.235562f
C135 VTAIL.t12 B 0.235562f
C136 VTAIL.n8 B 2.0779f
C137 VTAIL.n9 B 0.481412f
C138 VTAIL.t15 B 2.6524f
C139 VTAIL.n10 B 0.430279f
C140 VTAIL.t5 B 2.6524f
C141 VTAIL.n11 B 0.430279f
C142 VTAIL.t3 B 0.235562f
C143 VTAIL.t7 B 0.235562f
C144 VTAIL.n12 B 2.0779f
C145 VTAIL.n13 B 0.481412f
C146 VTAIL.t6 B 2.65238f
C147 VTAIL.n14 B 1.63451f
C148 VTAIL.t11 B 2.65238f
C149 VTAIL.n15 B 1.63096f
C150 VN.n0 B 0.029286f
C151 VN.t0 B 2.38009f
C152 VN.n1 B 0.028713f
C153 VN.n2 B 0.022213f
C154 VN.t4 B 2.38009f
C155 VN.n3 B 0.830953f
C156 VN.n4 B 0.022213f
C157 VN.n5 B 0.044148f
C158 VN.t3 B 2.55434f
C159 VN.n6 B 0.873849f
C160 VN.t7 B 2.38009f
C161 VN.n7 B 0.900294f
C162 VN.n8 B 0.037515f
C163 VN.n9 B 0.212056f
C164 VN.n10 B 0.022213f
C165 VN.n11 B 0.022213f
C166 VN.n12 B 0.017957f
C167 VN.n13 B 0.044148f
C168 VN.n14 B 0.037515f
C169 VN.n15 B 0.022213f
C170 VN.n16 B 0.022213f
C171 VN.n17 B 0.024843f
C172 VN.n18 B 0.0414f
C173 VN.n19 B 0.036141f
C174 VN.n20 B 0.022213f
C175 VN.n21 B 0.022213f
C176 VN.n22 B 0.022213f
C177 VN.n23 B 0.0414f
C178 VN.n24 B 0.029748f
C179 VN.n25 B 0.9025f
C180 VN.n26 B 0.03502f
C181 VN.n27 B 0.029286f
C182 VN.t2 B 2.38009f
C183 VN.n28 B 0.028713f
C184 VN.n29 B 0.022213f
C185 VN.t6 B 2.38009f
C186 VN.n30 B 0.830953f
C187 VN.n31 B 0.022213f
C188 VN.n32 B 0.044148f
C189 VN.t5 B 2.55434f
C190 VN.n33 B 0.873849f
C191 VN.t1 B 2.38009f
C192 VN.n34 B 0.900294f
C193 VN.n35 B 0.037515f
C194 VN.n36 B 0.212056f
C195 VN.n37 B 0.022213f
C196 VN.n38 B 0.022213f
C197 VN.n39 B 0.017957f
C198 VN.n40 B 0.044148f
C199 VN.n41 B 0.037515f
C200 VN.n42 B 0.022213f
C201 VN.n43 B 0.022213f
C202 VN.n44 B 0.024843f
C203 VN.n45 B 0.0414f
C204 VN.n46 B 0.036141f
C205 VN.n47 B 0.022213f
C206 VN.n48 B 0.022213f
C207 VN.n49 B 0.022213f
C208 VN.n50 B 0.0414f
C209 VN.n51 B 0.029748f
C210 VN.n52 B 0.9025f
C211 VN.n53 B 1.36171f
.ends

