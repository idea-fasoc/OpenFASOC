* NGSPICE file created from diff_pair_sample_1607.ext - technology: sky130A

.subckt diff_pair_sample_1607 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=6.8874 pd=36.1 as=0 ps=0 w=17.66 l=3.06
X1 VTAIL.t11 VN.t0 VDD2.t1 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=2.9139 pd=17.99 as=2.9139 ps=17.99 w=17.66 l=3.06
X2 VTAIL.t3 VP.t0 VDD1.t5 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=2.9139 pd=17.99 as=2.9139 ps=17.99 w=17.66 l=3.06
X3 VDD2.t0 VN.t1 VTAIL.t10 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=2.9139 pd=17.99 as=6.8874 ps=36.1 w=17.66 l=3.06
X4 VDD2.t4 VN.t2 VTAIL.t9 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=6.8874 pd=36.1 as=2.9139 ps=17.99 w=17.66 l=3.06
X5 VDD1.t4 VP.t1 VTAIL.t0 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=2.9139 pd=17.99 as=6.8874 ps=36.1 w=17.66 l=3.06
X6 VDD1.t3 VP.t2 VTAIL.t1 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=6.8874 pd=36.1 as=2.9139 ps=17.99 w=17.66 l=3.06
X7 VTAIL.t8 VN.t3 VDD2.t3 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=2.9139 pd=17.99 as=2.9139 ps=17.99 w=17.66 l=3.06
X8 VTAIL.t5 VP.t3 VDD1.t2 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=2.9139 pd=17.99 as=2.9139 ps=17.99 w=17.66 l=3.06
X9 VDD1.t1 VP.t4 VTAIL.t4 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=6.8874 pd=36.1 as=2.9139 ps=17.99 w=17.66 l=3.06
X10 VDD2.t2 VN.t4 VTAIL.t7 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=6.8874 pd=36.1 as=2.9139 ps=17.99 w=17.66 l=3.06
X11 B.t8 B.t6 B.t7 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=6.8874 pd=36.1 as=0 ps=0 w=17.66 l=3.06
X12 B.t5 B.t3 B.t4 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=6.8874 pd=36.1 as=0 ps=0 w=17.66 l=3.06
X13 VDD2.t5 VN.t5 VTAIL.t6 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=2.9139 pd=17.99 as=6.8874 ps=36.1 w=17.66 l=3.06
X14 B.t2 B.t0 B.t1 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=6.8874 pd=36.1 as=0 ps=0 w=17.66 l=3.06
X15 VDD1.t0 VP.t5 VTAIL.t2 w_n3682_n4500# sky130_fd_pr__pfet_01v8 ad=2.9139 pd=17.99 as=6.8874 ps=36.1 w=17.66 l=3.06
R0 B.n640 B.n93 585
R1 B.n642 B.n641 585
R2 B.n643 B.n92 585
R3 B.n645 B.n644 585
R4 B.n646 B.n91 585
R5 B.n648 B.n647 585
R6 B.n649 B.n90 585
R7 B.n651 B.n650 585
R8 B.n652 B.n89 585
R9 B.n654 B.n653 585
R10 B.n655 B.n88 585
R11 B.n657 B.n656 585
R12 B.n658 B.n87 585
R13 B.n660 B.n659 585
R14 B.n661 B.n86 585
R15 B.n663 B.n662 585
R16 B.n664 B.n85 585
R17 B.n666 B.n665 585
R18 B.n667 B.n84 585
R19 B.n669 B.n668 585
R20 B.n670 B.n83 585
R21 B.n672 B.n671 585
R22 B.n673 B.n82 585
R23 B.n675 B.n674 585
R24 B.n676 B.n81 585
R25 B.n678 B.n677 585
R26 B.n679 B.n80 585
R27 B.n681 B.n680 585
R28 B.n682 B.n79 585
R29 B.n684 B.n683 585
R30 B.n685 B.n78 585
R31 B.n687 B.n686 585
R32 B.n688 B.n77 585
R33 B.n690 B.n689 585
R34 B.n691 B.n76 585
R35 B.n693 B.n692 585
R36 B.n694 B.n75 585
R37 B.n696 B.n695 585
R38 B.n697 B.n74 585
R39 B.n699 B.n698 585
R40 B.n700 B.n73 585
R41 B.n702 B.n701 585
R42 B.n703 B.n72 585
R43 B.n705 B.n704 585
R44 B.n706 B.n71 585
R45 B.n708 B.n707 585
R46 B.n709 B.n70 585
R47 B.n711 B.n710 585
R48 B.n712 B.n69 585
R49 B.n714 B.n713 585
R50 B.n715 B.n68 585
R51 B.n717 B.n716 585
R52 B.n718 B.n67 585
R53 B.n720 B.n719 585
R54 B.n721 B.n66 585
R55 B.n723 B.n722 585
R56 B.n724 B.n65 585
R57 B.n726 B.n725 585
R58 B.n728 B.n727 585
R59 B.n729 B.n61 585
R60 B.n731 B.n730 585
R61 B.n732 B.n60 585
R62 B.n734 B.n733 585
R63 B.n735 B.n59 585
R64 B.n737 B.n736 585
R65 B.n738 B.n58 585
R66 B.n740 B.n739 585
R67 B.n741 B.n55 585
R68 B.n744 B.n743 585
R69 B.n745 B.n54 585
R70 B.n747 B.n746 585
R71 B.n748 B.n53 585
R72 B.n750 B.n749 585
R73 B.n751 B.n52 585
R74 B.n753 B.n752 585
R75 B.n754 B.n51 585
R76 B.n756 B.n755 585
R77 B.n757 B.n50 585
R78 B.n759 B.n758 585
R79 B.n760 B.n49 585
R80 B.n762 B.n761 585
R81 B.n763 B.n48 585
R82 B.n765 B.n764 585
R83 B.n766 B.n47 585
R84 B.n768 B.n767 585
R85 B.n769 B.n46 585
R86 B.n771 B.n770 585
R87 B.n772 B.n45 585
R88 B.n774 B.n773 585
R89 B.n775 B.n44 585
R90 B.n777 B.n776 585
R91 B.n778 B.n43 585
R92 B.n780 B.n779 585
R93 B.n781 B.n42 585
R94 B.n783 B.n782 585
R95 B.n784 B.n41 585
R96 B.n786 B.n785 585
R97 B.n787 B.n40 585
R98 B.n789 B.n788 585
R99 B.n790 B.n39 585
R100 B.n792 B.n791 585
R101 B.n793 B.n38 585
R102 B.n795 B.n794 585
R103 B.n796 B.n37 585
R104 B.n798 B.n797 585
R105 B.n799 B.n36 585
R106 B.n801 B.n800 585
R107 B.n802 B.n35 585
R108 B.n804 B.n803 585
R109 B.n805 B.n34 585
R110 B.n807 B.n806 585
R111 B.n808 B.n33 585
R112 B.n810 B.n809 585
R113 B.n811 B.n32 585
R114 B.n813 B.n812 585
R115 B.n814 B.n31 585
R116 B.n816 B.n815 585
R117 B.n817 B.n30 585
R118 B.n819 B.n818 585
R119 B.n820 B.n29 585
R120 B.n822 B.n821 585
R121 B.n823 B.n28 585
R122 B.n825 B.n824 585
R123 B.n826 B.n27 585
R124 B.n828 B.n827 585
R125 B.n829 B.n26 585
R126 B.n639 B.n638 585
R127 B.n637 B.n94 585
R128 B.n636 B.n635 585
R129 B.n634 B.n95 585
R130 B.n633 B.n632 585
R131 B.n631 B.n96 585
R132 B.n630 B.n629 585
R133 B.n628 B.n97 585
R134 B.n627 B.n626 585
R135 B.n625 B.n98 585
R136 B.n624 B.n623 585
R137 B.n622 B.n99 585
R138 B.n621 B.n620 585
R139 B.n619 B.n100 585
R140 B.n618 B.n617 585
R141 B.n616 B.n101 585
R142 B.n615 B.n614 585
R143 B.n613 B.n102 585
R144 B.n612 B.n611 585
R145 B.n610 B.n103 585
R146 B.n609 B.n608 585
R147 B.n607 B.n104 585
R148 B.n606 B.n605 585
R149 B.n604 B.n105 585
R150 B.n603 B.n602 585
R151 B.n601 B.n106 585
R152 B.n600 B.n599 585
R153 B.n598 B.n107 585
R154 B.n597 B.n596 585
R155 B.n595 B.n108 585
R156 B.n594 B.n593 585
R157 B.n592 B.n109 585
R158 B.n591 B.n590 585
R159 B.n589 B.n110 585
R160 B.n588 B.n587 585
R161 B.n586 B.n111 585
R162 B.n585 B.n584 585
R163 B.n583 B.n112 585
R164 B.n582 B.n581 585
R165 B.n580 B.n113 585
R166 B.n579 B.n578 585
R167 B.n577 B.n114 585
R168 B.n576 B.n575 585
R169 B.n574 B.n115 585
R170 B.n573 B.n572 585
R171 B.n571 B.n116 585
R172 B.n570 B.n569 585
R173 B.n568 B.n117 585
R174 B.n567 B.n566 585
R175 B.n565 B.n118 585
R176 B.n564 B.n563 585
R177 B.n562 B.n119 585
R178 B.n561 B.n560 585
R179 B.n559 B.n120 585
R180 B.n558 B.n557 585
R181 B.n556 B.n121 585
R182 B.n555 B.n554 585
R183 B.n553 B.n122 585
R184 B.n552 B.n551 585
R185 B.n550 B.n123 585
R186 B.n549 B.n548 585
R187 B.n547 B.n124 585
R188 B.n546 B.n545 585
R189 B.n544 B.n125 585
R190 B.n543 B.n542 585
R191 B.n541 B.n126 585
R192 B.n540 B.n539 585
R193 B.n538 B.n127 585
R194 B.n537 B.n536 585
R195 B.n535 B.n128 585
R196 B.n534 B.n533 585
R197 B.n532 B.n129 585
R198 B.n531 B.n530 585
R199 B.n529 B.n130 585
R200 B.n528 B.n527 585
R201 B.n526 B.n131 585
R202 B.n525 B.n524 585
R203 B.n523 B.n132 585
R204 B.n522 B.n521 585
R205 B.n520 B.n133 585
R206 B.n519 B.n518 585
R207 B.n517 B.n134 585
R208 B.n516 B.n515 585
R209 B.n514 B.n135 585
R210 B.n513 B.n512 585
R211 B.n511 B.n136 585
R212 B.n510 B.n509 585
R213 B.n508 B.n137 585
R214 B.n507 B.n506 585
R215 B.n505 B.n138 585
R216 B.n504 B.n503 585
R217 B.n502 B.n139 585
R218 B.n501 B.n500 585
R219 B.n499 B.n140 585
R220 B.n498 B.n497 585
R221 B.n496 B.n141 585
R222 B.n495 B.n494 585
R223 B.n304 B.n209 585
R224 B.n306 B.n305 585
R225 B.n307 B.n208 585
R226 B.n309 B.n308 585
R227 B.n310 B.n207 585
R228 B.n312 B.n311 585
R229 B.n313 B.n206 585
R230 B.n315 B.n314 585
R231 B.n316 B.n205 585
R232 B.n318 B.n317 585
R233 B.n319 B.n204 585
R234 B.n321 B.n320 585
R235 B.n322 B.n203 585
R236 B.n324 B.n323 585
R237 B.n325 B.n202 585
R238 B.n327 B.n326 585
R239 B.n328 B.n201 585
R240 B.n330 B.n329 585
R241 B.n331 B.n200 585
R242 B.n333 B.n332 585
R243 B.n334 B.n199 585
R244 B.n336 B.n335 585
R245 B.n337 B.n198 585
R246 B.n339 B.n338 585
R247 B.n340 B.n197 585
R248 B.n342 B.n341 585
R249 B.n343 B.n196 585
R250 B.n345 B.n344 585
R251 B.n346 B.n195 585
R252 B.n348 B.n347 585
R253 B.n349 B.n194 585
R254 B.n351 B.n350 585
R255 B.n352 B.n193 585
R256 B.n354 B.n353 585
R257 B.n355 B.n192 585
R258 B.n357 B.n356 585
R259 B.n358 B.n191 585
R260 B.n360 B.n359 585
R261 B.n361 B.n190 585
R262 B.n363 B.n362 585
R263 B.n364 B.n189 585
R264 B.n366 B.n365 585
R265 B.n367 B.n188 585
R266 B.n369 B.n368 585
R267 B.n370 B.n187 585
R268 B.n372 B.n371 585
R269 B.n373 B.n186 585
R270 B.n375 B.n374 585
R271 B.n376 B.n185 585
R272 B.n378 B.n377 585
R273 B.n379 B.n184 585
R274 B.n381 B.n380 585
R275 B.n382 B.n183 585
R276 B.n384 B.n383 585
R277 B.n385 B.n182 585
R278 B.n387 B.n386 585
R279 B.n388 B.n181 585
R280 B.n390 B.n389 585
R281 B.n392 B.n391 585
R282 B.n393 B.n177 585
R283 B.n395 B.n394 585
R284 B.n396 B.n176 585
R285 B.n398 B.n397 585
R286 B.n399 B.n175 585
R287 B.n401 B.n400 585
R288 B.n402 B.n174 585
R289 B.n404 B.n403 585
R290 B.n405 B.n171 585
R291 B.n408 B.n407 585
R292 B.n409 B.n170 585
R293 B.n411 B.n410 585
R294 B.n412 B.n169 585
R295 B.n414 B.n413 585
R296 B.n415 B.n168 585
R297 B.n417 B.n416 585
R298 B.n418 B.n167 585
R299 B.n420 B.n419 585
R300 B.n421 B.n166 585
R301 B.n423 B.n422 585
R302 B.n424 B.n165 585
R303 B.n426 B.n425 585
R304 B.n427 B.n164 585
R305 B.n429 B.n428 585
R306 B.n430 B.n163 585
R307 B.n432 B.n431 585
R308 B.n433 B.n162 585
R309 B.n435 B.n434 585
R310 B.n436 B.n161 585
R311 B.n438 B.n437 585
R312 B.n439 B.n160 585
R313 B.n441 B.n440 585
R314 B.n442 B.n159 585
R315 B.n444 B.n443 585
R316 B.n445 B.n158 585
R317 B.n447 B.n446 585
R318 B.n448 B.n157 585
R319 B.n450 B.n449 585
R320 B.n451 B.n156 585
R321 B.n453 B.n452 585
R322 B.n454 B.n155 585
R323 B.n456 B.n455 585
R324 B.n457 B.n154 585
R325 B.n459 B.n458 585
R326 B.n460 B.n153 585
R327 B.n462 B.n461 585
R328 B.n463 B.n152 585
R329 B.n465 B.n464 585
R330 B.n466 B.n151 585
R331 B.n468 B.n467 585
R332 B.n469 B.n150 585
R333 B.n471 B.n470 585
R334 B.n472 B.n149 585
R335 B.n474 B.n473 585
R336 B.n475 B.n148 585
R337 B.n477 B.n476 585
R338 B.n478 B.n147 585
R339 B.n480 B.n479 585
R340 B.n481 B.n146 585
R341 B.n483 B.n482 585
R342 B.n484 B.n145 585
R343 B.n486 B.n485 585
R344 B.n487 B.n144 585
R345 B.n489 B.n488 585
R346 B.n490 B.n143 585
R347 B.n492 B.n491 585
R348 B.n493 B.n142 585
R349 B.n303 B.n302 585
R350 B.n301 B.n210 585
R351 B.n300 B.n299 585
R352 B.n298 B.n211 585
R353 B.n297 B.n296 585
R354 B.n295 B.n212 585
R355 B.n294 B.n293 585
R356 B.n292 B.n213 585
R357 B.n291 B.n290 585
R358 B.n289 B.n214 585
R359 B.n288 B.n287 585
R360 B.n286 B.n215 585
R361 B.n285 B.n284 585
R362 B.n283 B.n216 585
R363 B.n282 B.n281 585
R364 B.n280 B.n217 585
R365 B.n279 B.n278 585
R366 B.n277 B.n218 585
R367 B.n276 B.n275 585
R368 B.n274 B.n219 585
R369 B.n273 B.n272 585
R370 B.n271 B.n220 585
R371 B.n270 B.n269 585
R372 B.n268 B.n221 585
R373 B.n267 B.n266 585
R374 B.n265 B.n222 585
R375 B.n264 B.n263 585
R376 B.n262 B.n223 585
R377 B.n261 B.n260 585
R378 B.n259 B.n224 585
R379 B.n258 B.n257 585
R380 B.n256 B.n225 585
R381 B.n255 B.n254 585
R382 B.n253 B.n226 585
R383 B.n252 B.n251 585
R384 B.n250 B.n227 585
R385 B.n249 B.n248 585
R386 B.n247 B.n228 585
R387 B.n246 B.n245 585
R388 B.n244 B.n229 585
R389 B.n243 B.n242 585
R390 B.n241 B.n230 585
R391 B.n240 B.n239 585
R392 B.n238 B.n231 585
R393 B.n237 B.n236 585
R394 B.n235 B.n232 585
R395 B.n234 B.n233 585
R396 B.n2 B.n0 585
R397 B.n901 B.n1 585
R398 B.n900 B.n899 585
R399 B.n898 B.n3 585
R400 B.n897 B.n896 585
R401 B.n895 B.n4 585
R402 B.n894 B.n893 585
R403 B.n892 B.n5 585
R404 B.n891 B.n890 585
R405 B.n889 B.n6 585
R406 B.n888 B.n887 585
R407 B.n886 B.n7 585
R408 B.n885 B.n884 585
R409 B.n883 B.n8 585
R410 B.n882 B.n881 585
R411 B.n880 B.n9 585
R412 B.n879 B.n878 585
R413 B.n877 B.n10 585
R414 B.n876 B.n875 585
R415 B.n874 B.n11 585
R416 B.n873 B.n872 585
R417 B.n871 B.n12 585
R418 B.n870 B.n869 585
R419 B.n868 B.n13 585
R420 B.n867 B.n866 585
R421 B.n865 B.n14 585
R422 B.n864 B.n863 585
R423 B.n862 B.n15 585
R424 B.n861 B.n860 585
R425 B.n859 B.n16 585
R426 B.n858 B.n857 585
R427 B.n856 B.n17 585
R428 B.n855 B.n854 585
R429 B.n853 B.n18 585
R430 B.n852 B.n851 585
R431 B.n850 B.n19 585
R432 B.n849 B.n848 585
R433 B.n847 B.n20 585
R434 B.n846 B.n845 585
R435 B.n844 B.n21 585
R436 B.n843 B.n842 585
R437 B.n841 B.n22 585
R438 B.n840 B.n839 585
R439 B.n838 B.n23 585
R440 B.n837 B.n836 585
R441 B.n835 B.n24 585
R442 B.n834 B.n833 585
R443 B.n832 B.n25 585
R444 B.n831 B.n830 585
R445 B.n903 B.n902 585
R446 B.n172 B.t8 543.525
R447 B.n62 B.t10 543.525
R448 B.n178 B.t5 543.525
R449 B.n56 B.t1 543.525
R450 B.n302 B.n209 506.916
R451 B.n830 B.n829 506.916
R452 B.n494 B.n493 506.916
R453 B.n638 B.n93 506.916
R454 B.n173 B.t7 477.781
R455 B.n63 B.t11 477.781
R456 B.n179 B.t4 477.779
R457 B.n57 B.t2 477.779
R458 B.n172 B.t6 347.736
R459 B.n178 B.t3 347.736
R460 B.n56 B.t0 347.736
R461 B.n62 B.t9 347.736
R462 B.n302 B.n301 163.367
R463 B.n301 B.n300 163.367
R464 B.n300 B.n211 163.367
R465 B.n296 B.n211 163.367
R466 B.n296 B.n295 163.367
R467 B.n295 B.n294 163.367
R468 B.n294 B.n213 163.367
R469 B.n290 B.n213 163.367
R470 B.n290 B.n289 163.367
R471 B.n289 B.n288 163.367
R472 B.n288 B.n215 163.367
R473 B.n284 B.n215 163.367
R474 B.n284 B.n283 163.367
R475 B.n283 B.n282 163.367
R476 B.n282 B.n217 163.367
R477 B.n278 B.n217 163.367
R478 B.n278 B.n277 163.367
R479 B.n277 B.n276 163.367
R480 B.n276 B.n219 163.367
R481 B.n272 B.n219 163.367
R482 B.n272 B.n271 163.367
R483 B.n271 B.n270 163.367
R484 B.n270 B.n221 163.367
R485 B.n266 B.n221 163.367
R486 B.n266 B.n265 163.367
R487 B.n265 B.n264 163.367
R488 B.n264 B.n223 163.367
R489 B.n260 B.n223 163.367
R490 B.n260 B.n259 163.367
R491 B.n259 B.n258 163.367
R492 B.n258 B.n225 163.367
R493 B.n254 B.n225 163.367
R494 B.n254 B.n253 163.367
R495 B.n253 B.n252 163.367
R496 B.n252 B.n227 163.367
R497 B.n248 B.n227 163.367
R498 B.n248 B.n247 163.367
R499 B.n247 B.n246 163.367
R500 B.n246 B.n229 163.367
R501 B.n242 B.n229 163.367
R502 B.n242 B.n241 163.367
R503 B.n241 B.n240 163.367
R504 B.n240 B.n231 163.367
R505 B.n236 B.n231 163.367
R506 B.n236 B.n235 163.367
R507 B.n235 B.n234 163.367
R508 B.n234 B.n2 163.367
R509 B.n902 B.n2 163.367
R510 B.n902 B.n901 163.367
R511 B.n901 B.n900 163.367
R512 B.n900 B.n3 163.367
R513 B.n896 B.n3 163.367
R514 B.n896 B.n895 163.367
R515 B.n895 B.n894 163.367
R516 B.n894 B.n5 163.367
R517 B.n890 B.n5 163.367
R518 B.n890 B.n889 163.367
R519 B.n889 B.n888 163.367
R520 B.n888 B.n7 163.367
R521 B.n884 B.n7 163.367
R522 B.n884 B.n883 163.367
R523 B.n883 B.n882 163.367
R524 B.n882 B.n9 163.367
R525 B.n878 B.n9 163.367
R526 B.n878 B.n877 163.367
R527 B.n877 B.n876 163.367
R528 B.n876 B.n11 163.367
R529 B.n872 B.n11 163.367
R530 B.n872 B.n871 163.367
R531 B.n871 B.n870 163.367
R532 B.n870 B.n13 163.367
R533 B.n866 B.n13 163.367
R534 B.n866 B.n865 163.367
R535 B.n865 B.n864 163.367
R536 B.n864 B.n15 163.367
R537 B.n860 B.n15 163.367
R538 B.n860 B.n859 163.367
R539 B.n859 B.n858 163.367
R540 B.n858 B.n17 163.367
R541 B.n854 B.n17 163.367
R542 B.n854 B.n853 163.367
R543 B.n853 B.n852 163.367
R544 B.n852 B.n19 163.367
R545 B.n848 B.n19 163.367
R546 B.n848 B.n847 163.367
R547 B.n847 B.n846 163.367
R548 B.n846 B.n21 163.367
R549 B.n842 B.n21 163.367
R550 B.n842 B.n841 163.367
R551 B.n841 B.n840 163.367
R552 B.n840 B.n23 163.367
R553 B.n836 B.n23 163.367
R554 B.n836 B.n835 163.367
R555 B.n835 B.n834 163.367
R556 B.n834 B.n25 163.367
R557 B.n830 B.n25 163.367
R558 B.n306 B.n209 163.367
R559 B.n307 B.n306 163.367
R560 B.n308 B.n307 163.367
R561 B.n308 B.n207 163.367
R562 B.n312 B.n207 163.367
R563 B.n313 B.n312 163.367
R564 B.n314 B.n313 163.367
R565 B.n314 B.n205 163.367
R566 B.n318 B.n205 163.367
R567 B.n319 B.n318 163.367
R568 B.n320 B.n319 163.367
R569 B.n320 B.n203 163.367
R570 B.n324 B.n203 163.367
R571 B.n325 B.n324 163.367
R572 B.n326 B.n325 163.367
R573 B.n326 B.n201 163.367
R574 B.n330 B.n201 163.367
R575 B.n331 B.n330 163.367
R576 B.n332 B.n331 163.367
R577 B.n332 B.n199 163.367
R578 B.n336 B.n199 163.367
R579 B.n337 B.n336 163.367
R580 B.n338 B.n337 163.367
R581 B.n338 B.n197 163.367
R582 B.n342 B.n197 163.367
R583 B.n343 B.n342 163.367
R584 B.n344 B.n343 163.367
R585 B.n344 B.n195 163.367
R586 B.n348 B.n195 163.367
R587 B.n349 B.n348 163.367
R588 B.n350 B.n349 163.367
R589 B.n350 B.n193 163.367
R590 B.n354 B.n193 163.367
R591 B.n355 B.n354 163.367
R592 B.n356 B.n355 163.367
R593 B.n356 B.n191 163.367
R594 B.n360 B.n191 163.367
R595 B.n361 B.n360 163.367
R596 B.n362 B.n361 163.367
R597 B.n362 B.n189 163.367
R598 B.n366 B.n189 163.367
R599 B.n367 B.n366 163.367
R600 B.n368 B.n367 163.367
R601 B.n368 B.n187 163.367
R602 B.n372 B.n187 163.367
R603 B.n373 B.n372 163.367
R604 B.n374 B.n373 163.367
R605 B.n374 B.n185 163.367
R606 B.n378 B.n185 163.367
R607 B.n379 B.n378 163.367
R608 B.n380 B.n379 163.367
R609 B.n380 B.n183 163.367
R610 B.n384 B.n183 163.367
R611 B.n385 B.n384 163.367
R612 B.n386 B.n385 163.367
R613 B.n386 B.n181 163.367
R614 B.n390 B.n181 163.367
R615 B.n391 B.n390 163.367
R616 B.n391 B.n177 163.367
R617 B.n395 B.n177 163.367
R618 B.n396 B.n395 163.367
R619 B.n397 B.n396 163.367
R620 B.n397 B.n175 163.367
R621 B.n401 B.n175 163.367
R622 B.n402 B.n401 163.367
R623 B.n403 B.n402 163.367
R624 B.n403 B.n171 163.367
R625 B.n408 B.n171 163.367
R626 B.n409 B.n408 163.367
R627 B.n410 B.n409 163.367
R628 B.n410 B.n169 163.367
R629 B.n414 B.n169 163.367
R630 B.n415 B.n414 163.367
R631 B.n416 B.n415 163.367
R632 B.n416 B.n167 163.367
R633 B.n420 B.n167 163.367
R634 B.n421 B.n420 163.367
R635 B.n422 B.n421 163.367
R636 B.n422 B.n165 163.367
R637 B.n426 B.n165 163.367
R638 B.n427 B.n426 163.367
R639 B.n428 B.n427 163.367
R640 B.n428 B.n163 163.367
R641 B.n432 B.n163 163.367
R642 B.n433 B.n432 163.367
R643 B.n434 B.n433 163.367
R644 B.n434 B.n161 163.367
R645 B.n438 B.n161 163.367
R646 B.n439 B.n438 163.367
R647 B.n440 B.n439 163.367
R648 B.n440 B.n159 163.367
R649 B.n444 B.n159 163.367
R650 B.n445 B.n444 163.367
R651 B.n446 B.n445 163.367
R652 B.n446 B.n157 163.367
R653 B.n450 B.n157 163.367
R654 B.n451 B.n450 163.367
R655 B.n452 B.n451 163.367
R656 B.n452 B.n155 163.367
R657 B.n456 B.n155 163.367
R658 B.n457 B.n456 163.367
R659 B.n458 B.n457 163.367
R660 B.n458 B.n153 163.367
R661 B.n462 B.n153 163.367
R662 B.n463 B.n462 163.367
R663 B.n464 B.n463 163.367
R664 B.n464 B.n151 163.367
R665 B.n468 B.n151 163.367
R666 B.n469 B.n468 163.367
R667 B.n470 B.n469 163.367
R668 B.n470 B.n149 163.367
R669 B.n474 B.n149 163.367
R670 B.n475 B.n474 163.367
R671 B.n476 B.n475 163.367
R672 B.n476 B.n147 163.367
R673 B.n480 B.n147 163.367
R674 B.n481 B.n480 163.367
R675 B.n482 B.n481 163.367
R676 B.n482 B.n145 163.367
R677 B.n486 B.n145 163.367
R678 B.n487 B.n486 163.367
R679 B.n488 B.n487 163.367
R680 B.n488 B.n143 163.367
R681 B.n492 B.n143 163.367
R682 B.n493 B.n492 163.367
R683 B.n494 B.n141 163.367
R684 B.n498 B.n141 163.367
R685 B.n499 B.n498 163.367
R686 B.n500 B.n499 163.367
R687 B.n500 B.n139 163.367
R688 B.n504 B.n139 163.367
R689 B.n505 B.n504 163.367
R690 B.n506 B.n505 163.367
R691 B.n506 B.n137 163.367
R692 B.n510 B.n137 163.367
R693 B.n511 B.n510 163.367
R694 B.n512 B.n511 163.367
R695 B.n512 B.n135 163.367
R696 B.n516 B.n135 163.367
R697 B.n517 B.n516 163.367
R698 B.n518 B.n517 163.367
R699 B.n518 B.n133 163.367
R700 B.n522 B.n133 163.367
R701 B.n523 B.n522 163.367
R702 B.n524 B.n523 163.367
R703 B.n524 B.n131 163.367
R704 B.n528 B.n131 163.367
R705 B.n529 B.n528 163.367
R706 B.n530 B.n529 163.367
R707 B.n530 B.n129 163.367
R708 B.n534 B.n129 163.367
R709 B.n535 B.n534 163.367
R710 B.n536 B.n535 163.367
R711 B.n536 B.n127 163.367
R712 B.n540 B.n127 163.367
R713 B.n541 B.n540 163.367
R714 B.n542 B.n541 163.367
R715 B.n542 B.n125 163.367
R716 B.n546 B.n125 163.367
R717 B.n547 B.n546 163.367
R718 B.n548 B.n547 163.367
R719 B.n548 B.n123 163.367
R720 B.n552 B.n123 163.367
R721 B.n553 B.n552 163.367
R722 B.n554 B.n553 163.367
R723 B.n554 B.n121 163.367
R724 B.n558 B.n121 163.367
R725 B.n559 B.n558 163.367
R726 B.n560 B.n559 163.367
R727 B.n560 B.n119 163.367
R728 B.n564 B.n119 163.367
R729 B.n565 B.n564 163.367
R730 B.n566 B.n565 163.367
R731 B.n566 B.n117 163.367
R732 B.n570 B.n117 163.367
R733 B.n571 B.n570 163.367
R734 B.n572 B.n571 163.367
R735 B.n572 B.n115 163.367
R736 B.n576 B.n115 163.367
R737 B.n577 B.n576 163.367
R738 B.n578 B.n577 163.367
R739 B.n578 B.n113 163.367
R740 B.n582 B.n113 163.367
R741 B.n583 B.n582 163.367
R742 B.n584 B.n583 163.367
R743 B.n584 B.n111 163.367
R744 B.n588 B.n111 163.367
R745 B.n589 B.n588 163.367
R746 B.n590 B.n589 163.367
R747 B.n590 B.n109 163.367
R748 B.n594 B.n109 163.367
R749 B.n595 B.n594 163.367
R750 B.n596 B.n595 163.367
R751 B.n596 B.n107 163.367
R752 B.n600 B.n107 163.367
R753 B.n601 B.n600 163.367
R754 B.n602 B.n601 163.367
R755 B.n602 B.n105 163.367
R756 B.n606 B.n105 163.367
R757 B.n607 B.n606 163.367
R758 B.n608 B.n607 163.367
R759 B.n608 B.n103 163.367
R760 B.n612 B.n103 163.367
R761 B.n613 B.n612 163.367
R762 B.n614 B.n613 163.367
R763 B.n614 B.n101 163.367
R764 B.n618 B.n101 163.367
R765 B.n619 B.n618 163.367
R766 B.n620 B.n619 163.367
R767 B.n620 B.n99 163.367
R768 B.n624 B.n99 163.367
R769 B.n625 B.n624 163.367
R770 B.n626 B.n625 163.367
R771 B.n626 B.n97 163.367
R772 B.n630 B.n97 163.367
R773 B.n631 B.n630 163.367
R774 B.n632 B.n631 163.367
R775 B.n632 B.n95 163.367
R776 B.n636 B.n95 163.367
R777 B.n637 B.n636 163.367
R778 B.n638 B.n637 163.367
R779 B.n829 B.n828 163.367
R780 B.n828 B.n27 163.367
R781 B.n824 B.n27 163.367
R782 B.n824 B.n823 163.367
R783 B.n823 B.n822 163.367
R784 B.n822 B.n29 163.367
R785 B.n818 B.n29 163.367
R786 B.n818 B.n817 163.367
R787 B.n817 B.n816 163.367
R788 B.n816 B.n31 163.367
R789 B.n812 B.n31 163.367
R790 B.n812 B.n811 163.367
R791 B.n811 B.n810 163.367
R792 B.n810 B.n33 163.367
R793 B.n806 B.n33 163.367
R794 B.n806 B.n805 163.367
R795 B.n805 B.n804 163.367
R796 B.n804 B.n35 163.367
R797 B.n800 B.n35 163.367
R798 B.n800 B.n799 163.367
R799 B.n799 B.n798 163.367
R800 B.n798 B.n37 163.367
R801 B.n794 B.n37 163.367
R802 B.n794 B.n793 163.367
R803 B.n793 B.n792 163.367
R804 B.n792 B.n39 163.367
R805 B.n788 B.n39 163.367
R806 B.n788 B.n787 163.367
R807 B.n787 B.n786 163.367
R808 B.n786 B.n41 163.367
R809 B.n782 B.n41 163.367
R810 B.n782 B.n781 163.367
R811 B.n781 B.n780 163.367
R812 B.n780 B.n43 163.367
R813 B.n776 B.n43 163.367
R814 B.n776 B.n775 163.367
R815 B.n775 B.n774 163.367
R816 B.n774 B.n45 163.367
R817 B.n770 B.n45 163.367
R818 B.n770 B.n769 163.367
R819 B.n769 B.n768 163.367
R820 B.n768 B.n47 163.367
R821 B.n764 B.n47 163.367
R822 B.n764 B.n763 163.367
R823 B.n763 B.n762 163.367
R824 B.n762 B.n49 163.367
R825 B.n758 B.n49 163.367
R826 B.n758 B.n757 163.367
R827 B.n757 B.n756 163.367
R828 B.n756 B.n51 163.367
R829 B.n752 B.n51 163.367
R830 B.n752 B.n751 163.367
R831 B.n751 B.n750 163.367
R832 B.n750 B.n53 163.367
R833 B.n746 B.n53 163.367
R834 B.n746 B.n745 163.367
R835 B.n745 B.n744 163.367
R836 B.n744 B.n55 163.367
R837 B.n739 B.n55 163.367
R838 B.n739 B.n738 163.367
R839 B.n738 B.n737 163.367
R840 B.n737 B.n59 163.367
R841 B.n733 B.n59 163.367
R842 B.n733 B.n732 163.367
R843 B.n732 B.n731 163.367
R844 B.n731 B.n61 163.367
R845 B.n727 B.n61 163.367
R846 B.n727 B.n726 163.367
R847 B.n726 B.n65 163.367
R848 B.n722 B.n65 163.367
R849 B.n722 B.n721 163.367
R850 B.n721 B.n720 163.367
R851 B.n720 B.n67 163.367
R852 B.n716 B.n67 163.367
R853 B.n716 B.n715 163.367
R854 B.n715 B.n714 163.367
R855 B.n714 B.n69 163.367
R856 B.n710 B.n69 163.367
R857 B.n710 B.n709 163.367
R858 B.n709 B.n708 163.367
R859 B.n708 B.n71 163.367
R860 B.n704 B.n71 163.367
R861 B.n704 B.n703 163.367
R862 B.n703 B.n702 163.367
R863 B.n702 B.n73 163.367
R864 B.n698 B.n73 163.367
R865 B.n698 B.n697 163.367
R866 B.n697 B.n696 163.367
R867 B.n696 B.n75 163.367
R868 B.n692 B.n75 163.367
R869 B.n692 B.n691 163.367
R870 B.n691 B.n690 163.367
R871 B.n690 B.n77 163.367
R872 B.n686 B.n77 163.367
R873 B.n686 B.n685 163.367
R874 B.n685 B.n684 163.367
R875 B.n684 B.n79 163.367
R876 B.n680 B.n79 163.367
R877 B.n680 B.n679 163.367
R878 B.n679 B.n678 163.367
R879 B.n678 B.n81 163.367
R880 B.n674 B.n81 163.367
R881 B.n674 B.n673 163.367
R882 B.n673 B.n672 163.367
R883 B.n672 B.n83 163.367
R884 B.n668 B.n83 163.367
R885 B.n668 B.n667 163.367
R886 B.n667 B.n666 163.367
R887 B.n666 B.n85 163.367
R888 B.n662 B.n85 163.367
R889 B.n662 B.n661 163.367
R890 B.n661 B.n660 163.367
R891 B.n660 B.n87 163.367
R892 B.n656 B.n87 163.367
R893 B.n656 B.n655 163.367
R894 B.n655 B.n654 163.367
R895 B.n654 B.n89 163.367
R896 B.n650 B.n89 163.367
R897 B.n650 B.n649 163.367
R898 B.n649 B.n648 163.367
R899 B.n648 B.n91 163.367
R900 B.n644 B.n91 163.367
R901 B.n644 B.n643 163.367
R902 B.n643 B.n642 163.367
R903 B.n642 B.n93 163.367
R904 B.n173 B.n172 65.746
R905 B.n179 B.n178 65.746
R906 B.n57 B.n56 65.746
R907 B.n63 B.n62 65.746
R908 B.n406 B.n173 59.5399
R909 B.n180 B.n179 59.5399
R910 B.n742 B.n57 59.5399
R911 B.n64 B.n63 59.5399
R912 B.n831 B.n26 32.9371
R913 B.n640 B.n639 32.9371
R914 B.n495 B.n142 32.9371
R915 B.n304 B.n303 32.9371
R916 B B.n903 18.0485
R917 B.n827 B.n26 10.6151
R918 B.n827 B.n826 10.6151
R919 B.n826 B.n825 10.6151
R920 B.n825 B.n28 10.6151
R921 B.n821 B.n28 10.6151
R922 B.n821 B.n820 10.6151
R923 B.n820 B.n819 10.6151
R924 B.n819 B.n30 10.6151
R925 B.n815 B.n30 10.6151
R926 B.n815 B.n814 10.6151
R927 B.n814 B.n813 10.6151
R928 B.n813 B.n32 10.6151
R929 B.n809 B.n32 10.6151
R930 B.n809 B.n808 10.6151
R931 B.n808 B.n807 10.6151
R932 B.n807 B.n34 10.6151
R933 B.n803 B.n34 10.6151
R934 B.n803 B.n802 10.6151
R935 B.n802 B.n801 10.6151
R936 B.n801 B.n36 10.6151
R937 B.n797 B.n36 10.6151
R938 B.n797 B.n796 10.6151
R939 B.n796 B.n795 10.6151
R940 B.n795 B.n38 10.6151
R941 B.n791 B.n38 10.6151
R942 B.n791 B.n790 10.6151
R943 B.n790 B.n789 10.6151
R944 B.n789 B.n40 10.6151
R945 B.n785 B.n40 10.6151
R946 B.n785 B.n784 10.6151
R947 B.n784 B.n783 10.6151
R948 B.n783 B.n42 10.6151
R949 B.n779 B.n42 10.6151
R950 B.n779 B.n778 10.6151
R951 B.n778 B.n777 10.6151
R952 B.n777 B.n44 10.6151
R953 B.n773 B.n44 10.6151
R954 B.n773 B.n772 10.6151
R955 B.n772 B.n771 10.6151
R956 B.n771 B.n46 10.6151
R957 B.n767 B.n46 10.6151
R958 B.n767 B.n766 10.6151
R959 B.n766 B.n765 10.6151
R960 B.n765 B.n48 10.6151
R961 B.n761 B.n48 10.6151
R962 B.n761 B.n760 10.6151
R963 B.n760 B.n759 10.6151
R964 B.n759 B.n50 10.6151
R965 B.n755 B.n50 10.6151
R966 B.n755 B.n754 10.6151
R967 B.n754 B.n753 10.6151
R968 B.n753 B.n52 10.6151
R969 B.n749 B.n52 10.6151
R970 B.n749 B.n748 10.6151
R971 B.n748 B.n747 10.6151
R972 B.n747 B.n54 10.6151
R973 B.n743 B.n54 10.6151
R974 B.n741 B.n740 10.6151
R975 B.n740 B.n58 10.6151
R976 B.n736 B.n58 10.6151
R977 B.n736 B.n735 10.6151
R978 B.n735 B.n734 10.6151
R979 B.n734 B.n60 10.6151
R980 B.n730 B.n60 10.6151
R981 B.n730 B.n729 10.6151
R982 B.n729 B.n728 10.6151
R983 B.n725 B.n724 10.6151
R984 B.n724 B.n723 10.6151
R985 B.n723 B.n66 10.6151
R986 B.n719 B.n66 10.6151
R987 B.n719 B.n718 10.6151
R988 B.n718 B.n717 10.6151
R989 B.n717 B.n68 10.6151
R990 B.n713 B.n68 10.6151
R991 B.n713 B.n712 10.6151
R992 B.n712 B.n711 10.6151
R993 B.n711 B.n70 10.6151
R994 B.n707 B.n70 10.6151
R995 B.n707 B.n706 10.6151
R996 B.n706 B.n705 10.6151
R997 B.n705 B.n72 10.6151
R998 B.n701 B.n72 10.6151
R999 B.n701 B.n700 10.6151
R1000 B.n700 B.n699 10.6151
R1001 B.n699 B.n74 10.6151
R1002 B.n695 B.n74 10.6151
R1003 B.n695 B.n694 10.6151
R1004 B.n694 B.n693 10.6151
R1005 B.n693 B.n76 10.6151
R1006 B.n689 B.n76 10.6151
R1007 B.n689 B.n688 10.6151
R1008 B.n688 B.n687 10.6151
R1009 B.n687 B.n78 10.6151
R1010 B.n683 B.n78 10.6151
R1011 B.n683 B.n682 10.6151
R1012 B.n682 B.n681 10.6151
R1013 B.n681 B.n80 10.6151
R1014 B.n677 B.n80 10.6151
R1015 B.n677 B.n676 10.6151
R1016 B.n676 B.n675 10.6151
R1017 B.n675 B.n82 10.6151
R1018 B.n671 B.n82 10.6151
R1019 B.n671 B.n670 10.6151
R1020 B.n670 B.n669 10.6151
R1021 B.n669 B.n84 10.6151
R1022 B.n665 B.n84 10.6151
R1023 B.n665 B.n664 10.6151
R1024 B.n664 B.n663 10.6151
R1025 B.n663 B.n86 10.6151
R1026 B.n659 B.n86 10.6151
R1027 B.n659 B.n658 10.6151
R1028 B.n658 B.n657 10.6151
R1029 B.n657 B.n88 10.6151
R1030 B.n653 B.n88 10.6151
R1031 B.n653 B.n652 10.6151
R1032 B.n652 B.n651 10.6151
R1033 B.n651 B.n90 10.6151
R1034 B.n647 B.n90 10.6151
R1035 B.n647 B.n646 10.6151
R1036 B.n646 B.n645 10.6151
R1037 B.n645 B.n92 10.6151
R1038 B.n641 B.n92 10.6151
R1039 B.n641 B.n640 10.6151
R1040 B.n496 B.n495 10.6151
R1041 B.n497 B.n496 10.6151
R1042 B.n497 B.n140 10.6151
R1043 B.n501 B.n140 10.6151
R1044 B.n502 B.n501 10.6151
R1045 B.n503 B.n502 10.6151
R1046 B.n503 B.n138 10.6151
R1047 B.n507 B.n138 10.6151
R1048 B.n508 B.n507 10.6151
R1049 B.n509 B.n508 10.6151
R1050 B.n509 B.n136 10.6151
R1051 B.n513 B.n136 10.6151
R1052 B.n514 B.n513 10.6151
R1053 B.n515 B.n514 10.6151
R1054 B.n515 B.n134 10.6151
R1055 B.n519 B.n134 10.6151
R1056 B.n520 B.n519 10.6151
R1057 B.n521 B.n520 10.6151
R1058 B.n521 B.n132 10.6151
R1059 B.n525 B.n132 10.6151
R1060 B.n526 B.n525 10.6151
R1061 B.n527 B.n526 10.6151
R1062 B.n527 B.n130 10.6151
R1063 B.n531 B.n130 10.6151
R1064 B.n532 B.n531 10.6151
R1065 B.n533 B.n532 10.6151
R1066 B.n533 B.n128 10.6151
R1067 B.n537 B.n128 10.6151
R1068 B.n538 B.n537 10.6151
R1069 B.n539 B.n538 10.6151
R1070 B.n539 B.n126 10.6151
R1071 B.n543 B.n126 10.6151
R1072 B.n544 B.n543 10.6151
R1073 B.n545 B.n544 10.6151
R1074 B.n545 B.n124 10.6151
R1075 B.n549 B.n124 10.6151
R1076 B.n550 B.n549 10.6151
R1077 B.n551 B.n550 10.6151
R1078 B.n551 B.n122 10.6151
R1079 B.n555 B.n122 10.6151
R1080 B.n556 B.n555 10.6151
R1081 B.n557 B.n556 10.6151
R1082 B.n557 B.n120 10.6151
R1083 B.n561 B.n120 10.6151
R1084 B.n562 B.n561 10.6151
R1085 B.n563 B.n562 10.6151
R1086 B.n563 B.n118 10.6151
R1087 B.n567 B.n118 10.6151
R1088 B.n568 B.n567 10.6151
R1089 B.n569 B.n568 10.6151
R1090 B.n569 B.n116 10.6151
R1091 B.n573 B.n116 10.6151
R1092 B.n574 B.n573 10.6151
R1093 B.n575 B.n574 10.6151
R1094 B.n575 B.n114 10.6151
R1095 B.n579 B.n114 10.6151
R1096 B.n580 B.n579 10.6151
R1097 B.n581 B.n580 10.6151
R1098 B.n581 B.n112 10.6151
R1099 B.n585 B.n112 10.6151
R1100 B.n586 B.n585 10.6151
R1101 B.n587 B.n586 10.6151
R1102 B.n587 B.n110 10.6151
R1103 B.n591 B.n110 10.6151
R1104 B.n592 B.n591 10.6151
R1105 B.n593 B.n592 10.6151
R1106 B.n593 B.n108 10.6151
R1107 B.n597 B.n108 10.6151
R1108 B.n598 B.n597 10.6151
R1109 B.n599 B.n598 10.6151
R1110 B.n599 B.n106 10.6151
R1111 B.n603 B.n106 10.6151
R1112 B.n604 B.n603 10.6151
R1113 B.n605 B.n604 10.6151
R1114 B.n605 B.n104 10.6151
R1115 B.n609 B.n104 10.6151
R1116 B.n610 B.n609 10.6151
R1117 B.n611 B.n610 10.6151
R1118 B.n611 B.n102 10.6151
R1119 B.n615 B.n102 10.6151
R1120 B.n616 B.n615 10.6151
R1121 B.n617 B.n616 10.6151
R1122 B.n617 B.n100 10.6151
R1123 B.n621 B.n100 10.6151
R1124 B.n622 B.n621 10.6151
R1125 B.n623 B.n622 10.6151
R1126 B.n623 B.n98 10.6151
R1127 B.n627 B.n98 10.6151
R1128 B.n628 B.n627 10.6151
R1129 B.n629 B.n628 10.6151
R1130 B.n629 B.n96 10.6151
R1131 B.n633 B.n96 10.6151
R1132 B.n634 B.n633 10.6151
R1133 B.n635 B.n634 10.6151
R1134 B.n635 B.n94 10.6151
R1135 B.n639 B.n94 10.6151
R1136 B.n305 B.n304 10.6151
R1137 B.n305 B.n208 10.6151
R1138 B.n309 B.n208 10.6151
R1139 B.n310 B.n309 10.6151
R1140 B.n311 B.n310 10.6151
R1141 B.n311 B.n206 10.6151
R1142 B.n315 B.n206 10.6151
R1143 B.n316 B.n315 10.6151
R1144 B.n317 B.n316 10.6151
R1145 B.n317 B.n204 10.6151
R1146 B.n321 B.n204 10.6151
R1147 B.n322 B.n321 10.6151
R1148 B.n323 B.n322 10.6151
R1149 B.n323 B.n202 10.6151
R1150 B.n327 B.n202 10.6151
R1151 B.n328 B.n327 10.6151
R1152 B.n329 B.n328 10.6151
R1153 B.n329 B.n200 10.6151
R1154 B.n333 B.n200 10.6151
R1155 B.n334 B.n333 10.6151
R1156 B.n335 B.n334 10.6151
R1157 B.n335 B.n198 10.6151
R1158 B.n339 B.n198 10.6151
R1159 B.n340 B.n339 10.6151
R1160 B.n341 B.n340 10.6151
R1161 B.n341 B.n196 10.6151
R1162 B.n345 B.n196 10.6151
R1163 B.n346 B.n345 10.6151
R1164 B.n347 B.n346 10.6151
R1165 B.n347 B.n194 10.6151
R1166 B.n351 B.n194 10.6151
R1167 B.n352 B.n351 10.6151
R1168 B.n353 B.n352 10.6151
R1169 B.n353 B.n192 10.6151
R1170 B.n357 B.n192 10.6151
R1171 B.n358 B.n357 10.6151
R1172 B.n359 B.n358 10.6151
R1173 B.n359 B.n190 10.6151
R1174 B.n363 B.n190 10.6151
R1175 B.n364 B.n363 10.6151
R1176 B.n365 B.n364 10.6151
R1177 B.n365 B.n188 10.6151
R1178 B.n369 B.n188 10.6151
R1179 B.n370 B.n369 10.6151
R1180 B.n371 B.n370 10.6151
R1181 B.n371 B.n186 10.6151
R1182 B.n375 B.n186 10.6151
R1183 B.n376 B.n375 10.6151
R1184 B.n377 B.n376 10.6151
R1185 B.n377 B.n184 10.6151
R1186 B.n381 B.n184 10.6151
R1187 B.n382 B.n381 10.6151
R1188 B.n383 B.n382 10.6151
R1189 B.n383 B.n182 10.6151
R1190 B.n387 B.n182 10.6151
R1191 B.n388 B.n387 10.6151
R1192 B.n389 B.n388 10.6151
R1193 B.n393 B.n392 10.6151
R1194 B.n394 B.n393 10.6151
R1195 B.n394 B.n176 10.6151
R1196 B.n398 B.n176 10.6151
R1197 B.n399 B.n398 10.6151
R1198 B.n400 B.n399 10.6151
R1199 B.n400 B.n174 10.6151
R1200 B.n404 B.n174 10.6151
R1201 B.n405 B.n404 10.6151
R1202 B.n407 B.n170 10.6151
R1203 B.n411 B.n170 10.6151
R1204 B.n412 B.n411 10.6151
R1205 B.n413 B.n412 10.6151
R1206 B.n413 B.n168 10.6151
R1207 B.n417 B.n168 10.6151
R1208 B.n418 B.n417 10.6151
R1209 B.n419 B.n418 10.6151
R1210 B.n419 B.n166 10.6151
R1211 B.n423 B.n166 10.6151
R1212 B.n424 B.n423 10.6151
R1213 B.n425 B.n424 10.6151
R1214 B.n425 B.n164 10.6151
R1215 B.n429 B.n164 10.6151
R1216 B.n430 B.n429 10.6151
R1217 B.n431 B.n430 10.6151
R1218 B.n431 B.n162 10.6151
R1219 B.n435 B.n162 10.6151
R1220 B.n436 B.n435 10.6151
R1221 B.n437 B.n436 10.6151
R1222 B.n437 B.n160 10.6151
R1223 B.n441 B.n160 10.6151
R1224 B.n442 B.n441 10.6151
R1225 B.n443 B.n442 10.6151
R1226 B.n443 B.n158 10.6151
R1227 B.n447 B.n158 10.6151
R1228 B.n448 B.n447 10.6151
R1229 B.n449 B.n448 10.6151
R1230 B.n449 B.n156 10.6151
R1231 B.n453 B.n156 10.6151
R1232 B.n454 B.n453 10.6151
R1233 B.n455 B.n454 10.6151
R1234 B.n455 B.n154 10.6151
R1235 B.n459 B.n154 10.6151
R1236 B.n460 B.n459 10.6151
R1237 B.n461 B.n460 10.6151
R1238 B.n461 B.n152 10.6151
R1239 B.n465 B.n152 10.6151
R1240 B.n466 B.n465 10.6151
R1241 B.n467 B.n466 10.6151
R1242 B.n467 B.n150 10.6151
R1243 B.n471 B.n150 10.6151
R1244 B.n472 B.n471 10.6151
R1245 B.n473 B.n472 10.6151
R1246 B.n473 B.n148 10.6151
R1247 B.n477 B.n148 10.6151
R1248 B.n478 B.n477 10.6151
R1249 B.n479 B.n478 10.6151
R1250 B.n479 B.n146 10.6151
R1251 B.n483 B.n146 10.6151
R1252 B.n484 B.n483 10.6151
R1253 B.n485 B.n484 10.6151
R1254 B.n485 B.n144 10.6151
R1255 B.n489 B.n144 10.6151
R1256 B.n490 B.n489 10.6151
R1257 B.n491 B.n490 10.6151
R1258 B.n491 B.n142 10.6151
R1259 B.n303 B.n210 10.6151
R1260 B.n299 B.n210 10.6151
R1261 B.n299 B.n298 10.6151
R1262 B.n298 B.n297 10.6151
R1263 B.n297 B.n212 10.6151
R1264 B.n293 B.n212 10.6151
R1265 B.n293 B.n292 10.6151
R1266 B.n292 B.n291 10.6151
R1267 B.n291 B.n214 10.6151
R1268 B.n287 B.n214 10.6151
R1269 B.n287 B.n286 10.6151
R1270 B.n286 B.n285 10.6151
R1271 B.n285 B.n216 10.6151
R1272 B.n281 B.n216 10.6151
R1273 B.n281 B.n280 10.6151
R1274 B.n280 B.n279 10.6151
R1275 B.n279 B.n218 10.6151
R1276 B.n275 B.n218 10.6151
R1277 B.n275 B.n274 10.6151
R1278 B.n274 B.n273 10.6151
R1279 B.n273 B.n220 10.6151
R1280 B.n269 B.n220 10.6151
R1281 B.n269 B.n268 10.6151
R1282 B.n268 B.n267 10.6151
R1283 B.n267 B.n222 10.6151
R1284 B.n263 B.n222 10.6151
R1285 B.n263 B.n262 10.6151
R1286 B.n262 B.n261 10.6151
R1287 B.n261 B.n224 10.6151
R1288 B.n257 B.n224 10.6151
R1289 B.n257 B.n256 10.6151
R1290 B.n256 B.n255 10.6151
R1291 B.n255 B.n226 10.6151
R1292 B.n251 B.n226 10.6151
R1293 B.n251 B.n250 10.6151
R1294 B.n250 B.n249 10.6151
R1295 B.n249 B.n228 10.6151
R1296 B.n245 B.n228 10.6151
R1297 B.n245 B.n244 10.6151
R1298 B.n244 B.n243 10.6151
R1299 B.n243 B.n230 10.6151
R1300 B.n239 B.n230 10.6151
R1301 B.n239 B.n238 10.6151
R1302 B.n238 B.n237 10.6151
R1303 B.n237 B.n232 10.6151
R1304 B.n233 B.n232 10.6151
R1305 B.n233 B.n0 10.6151
R1306 B.n899 B.n1 10.6151
R1307 B.n899 B.n898 10.6151
R1308 B.n898 B.n897 10.6151
R1309 B.n897 B.n4 10.6151
R1310 B.n893 B.n4 10.6151
R1311 B.n893 B.n892 10.6151
R1312 B.n892 B.n891 10.6151
R1313 B.n891 B.n6 10.6151
R1314 B.n887 B.n6 10.6151
R1315 B.n887 B.n886 10.6151
R1316 B.n886 B.n885 10.6151
R1317 B.n885 B.n8 10.6151
R1318 B.n881 B.n8 10.6151
R1319 B.n881 B.n880 10.6151
R1320 B.n880 B.n879 10.6151
R1321 B.n879 B.n10 10.6151
R1322 B.n875 B.n10 10.6151
R1323 B.n875 B.n874 10.6151
R1324 B.n874 B.n873 10.6151
R1325 B.n873 B.n12 10.6151
R1326 B.n869 B.n12 10.6151
R1327 B.n869 B.n868 10.6151
R1328 B.n868 B.n867 10.6151
R1329 B.n867 B.n14 10.6151
R1330 B.n863 B.n14 10.6151
R1331 B.n863 B.n862 10.6151
R1332 B.n862 B.n861 10.6151
R1333 B.n861 B.n16 10.6151
R1334 B.n857 B.n16 10.6151
R1335 B.n857 B.n856 10.6151
R1336 B.n856 B.n855 10.6151
R1337 B.n855 B.n18 10.6151
R1338 B.n851 B.n18 10.6151
R1339 B.n851 B.n850 10.6151
R1340 B.n850 B.n849 10.6151
R1341 B.n849 B.n20 10.6151
R1342 B.n845 B.n20 10.6151
R1343 B.n845 B.n844 10.6151
R1344 B.n844 B.n843 10.6151
R1345 B.n843 B.n22 10.6151
R1346 B.n839 B.n22 10.6151
R1347 B.n839 B.n838 10.6151
R1348 B.n838 B.n837 10.6151
R1349 B.n837 B.n24 10.6151
R1350 B.n833 B.n24 10.6151
R1351 B.n833 B.n832 10.6151
R1352 B.n832 B.n831 10.6151
R1353 B.n743 B.n742 9.36635
R1354 B.n725 B.n64 9.36635
R1355 B.n389 B.n180 9.36635
R1356 B.n407 B.n406 9.36635
R1357 B.n903 B.n0 2.81026
R1358 B.n903 B.n1 2.81026
R1359 B.n742 B.n741 1.24928
R1360 B.n728 B.n64 1.24928
R1361 B.n392 B.n180 1.24928
R1362 B.n406 B.n405 1.24928
R1363 VN.n20 VN.t1 172.542
R1364 VN.n4 VN.t4 172.542
R1365 VN.n30 VN.n29 161.3
R1366 VN.n28 VN.n17 161.3
R1367 VN.n27 VN.n26 161.3
R1368 VN.n25 VN.n18 161.3
R1369 VN.n24 VN.n23 161.3
R1370 VN.n22 VN.n19 161.3
R1371 VN.n14 VN.n13 161.3
R1372 VN.n12 VN.n1 161.3
R1373 VN.n11 VN.n10 161.3
R1374 VN.n9 VN.n2 161.3
R1375 VN.n8 VN.n7 161.3
R1376 VN.n6 VN.n3 161.3
R1377 VN.n5 VN.t0 139.088
R1378 VN.n0 VN.t5 139.088
R1379 VN.n21 VN.t3 139.088
R1380 VN.n16 VN.t2 139.088
R1381 VN.n15 VN.n0 71.0639
R1382 VN.n31 VN.n16 71.0639
R1383 VN.n11 VN.n2 56.5617
R1384 VN.n27 VN.n18 56.5617
R1385 VN VN.n31 55.055
R1386 VN.n5 VN.n4 49.4645
R1387 VN.n21 VN.n20 49.4645
R1388 VN.n6 VN.n5 24.5923
R1389 VN.n7 VN.n6 24.5923
R1390 VN.n7 VN.n2 24.5923
R1391 VN.n12 VN.n11 24.5923
R1392 VN.n13 VN.n12 24.5923
R1393 VN.n23 VN.n18 24.5923
R1394 VN.n23 VN.n22 24.5923
R1395 VN.n22 VN.n21 24.5923
R1396 VN.n29 VN.n28 24.5923
R1397 VN.n28 VN.n27 24.5923
R1398 VN.n13 VN.n0 19.1821
R1399 VN.n29 VN.n16 19.1821
R1400 VN.n4 VN.n3 3.94397
R1401 VN.n20 VN.n19 3.94397
R1402 VN.n31 VN.n30 0.354861
R1403 VN.n15 VN.n14 0.354861
R1404 VN VN.n15 0.267071
R1405 VN.n30 VN.n17 0.189894
R1406 VN.n26 VN.n17 0.189894
R1407 VN.n26 VN.n25 0.189894
R1408 VN.n25 VN.n24 0.189894
R1409 VN.n24 VN.n19 0.189894
R1410 VN.n8 VN.n3 0.189894
R1411 VN.n9 VN.n8 0.189894
R1412 VN.n10 VN.n9 0.189894
R1413 VN.n10 VN.n1 0.189894
R1414 VN.n14 VN.n1 0.189894
R1415 VDD2.n191 VDD2.n99 756.745
R1416 VDD2.n92 VDD2.n0 756.745
R1417 VDD2.n192 VDD2.n191 585
R1418 VDD2.n190 VDD2.n189 585
R1419 VDD2.n103 VDD2.n102 585
R1420 VDD2.n184 VDD2.n183 585
R1421 VDD2.n182 VDD2.n181 585
R1422 VDD2.n107 VDD2.n106 585
R1423 VDD2.n111 VDD2.n109 585
R1424 VDD2.n176 VDD2.n175 585
R1425 VDD2.n174 VDD2.n173 585
R1426 VDD2.n113 VDD2.n112 585
R1427 VDD2.n168 VDD2.n167 585
R1428 VDD2.n166 VDD2.n165 585
R1429 VDD2.n117 VDD2.n116 585
R1430 VDD2.n160 VDD2.n159 585
R1431 VDD2.n158 VDD2.n157 585
R1432 VDD2.n121 VDD2.n120 585
R1433 VDD2.n152 VDD2.n151 585
R1434 VDD2.n150 VDD2.n149 585
R1435 VDD2.n125 VDD2.n124 585
R1436 VDD2.n144 VDD2.n143 585
R1437 VDD2.n142 VDD2.n141 585
R1438 VDD2.n129 VDD2.n128 585
R1439 VDD2.n136 VDD2.n135 585
R1440 VDD2.n134 VDD2.n133 585
R1441 VDD2.n33 VDD2.n32 585
R1442 VDD2.n35 VDD2.n34 585
R1443 VDD2.n28 VDD2.n27 585
R1444 VDD2.n41 VDD2.n40 585
R1445 VDD2.n43 VDD2.n42 585
R1446 VDD2.n24 VDD2.n23 585
R1447 VDD2.n49 VDD2.n48 585
R1448 VDD2.n51 VDD2.n50 585
R1449 VDD2.n20 VDD2.n19 585
R1450 VDD2.n57 VDD2.n56 585
R1451 VDD2.n59 VDD2.n58 585
R1452 VDD2.n16 VDD2.n15 585
R1453 VDD2.n65 VDD2.n64 585
R1454 VDD2.n67 VDD2.n66 585
R1455 VDD2.n12 VDD2.n11 585
R1456 VDD2.n74 VDD2.n73 585
R1457 VDD2.n75 VDD2.n10 585
R1458 VDD2.n77 VDD2.n76 585
R1459 VDD2.n8 VDD2.n7 585
R1460 VDD2.n83 VDD2.n82 585
R1461 VDD2.n85 VDD2.n84 585
R1462 VDD2.n4 VDD2.n3 585
R1463 VDD2.n91 VDD2.n90 585
R1464 VDD2.n93 VDD2.n92 585
R1465 VDD2.n132 VDD2.t4 327.466
R1466 VDD2.n31 VDD2.t2 327.466
R1467 VDD2.n191 VDD2.n190 171.744
R1468 VDD2.n190 VDD2.n102 171.744
R1469 VDD2.n183 VDD2.n102 171.744
R1470 VDD2.n183 VDD2.n182 171.744
R1471 VDD2.n182 VDD2.n106 171.744
R1472 VDD2.n111 VDD2.n106 171.744
R1473 VDD2.n175 VDD2.n111 171.744
R1474 VDD2.n175 VDD2.n174 171.744
R1475 VDD2.n174 VDD2.n112 171.744
R1476 VDD2.n167 VDD2.n112 171.744
R1477 VDD2.n167 VDD2.n166 171.744
R1478 VDD2.n166 VDD2.n116 171.744
R1479 VDD2.n159 VDD2.n116 171.744
R1480 VDD2.n159 VDD2.n158 171.744
R1481 VDD2.n158 VDD2.n120 171.744
R1482 VDD2.n151 VDD2.n120 171.744
R1483 VDD2.n151 VDD2.n150 171.744
R1484 VDD2.n150 VDD2.n124 171.744
R1485 VDD2.n143 VDD2.n124 171.744
R1486 VDD2.n143 VDD2.n142 171.744
R1487 VDD2.n142 VDD2.n128 171.744
R1488 VDD2.n135 VDD2.n128 171.744
R1489 VDD2.n135 VDD2.n134 171.744
R1490 VDD2.n34 VDD2.n33 171.744
R1491 VDD2.n34 VDD2.n27 171.744
R1492 VDD2.n41 VDD2.n27 171.744
R1493 VDD2.n42 VDD2.n41 171.744
R1494 VDD2.n42 VDD2.n23 171.744
R1495 VDD2.n49 VDD2.n23 171.744
R1496 VDD2.n50 VDD2.n49 171.744
R1497 VDD2.n50 VDD2.n19 171.744
R1498 VDD2.n57 VDD2.n19 171.744
R1499 VDD2.n58 VDD2.n57 171.744
R1500 VDD2.n58 VDD2.n15 171.744
R1501 VDD2.n65 VDD2.n15 171.744
R1502 VDD2.n66 VDD2.n65 171.744
R1503 VDD2.n66 VDD2.n11 171.744
R1504 VDD2.n74 VDD2.n11 171.744
R1505 VDD2.n75 VDD2.n74 171.744
R1506 VDD2.n76 VDD2.n75 171.744
R1507 VDD2.n76 VDD2.n7 171.744
R1508 VDD2.n83 VDD2.n7 171.744
R1509 VDD2.n84 VDD2.n83 171.744
R1510 VDD2.n84 VDD2.n3 171.744
R1511 VDD2.n91 VDD2.n3 171.744
R1512 VDD2.n92 VDD2.n91 171.744
R1513 VDD2.n134 VDD2.t4 85.8723
R1514 VDD2.n33 VDD2.t2 85.8723
R1515 VDD2.n98 VDD2.n97 72.4125
R1516 VDD2 VDD2.n197 72.4096
R1517 VDD2.n98 VDD2.n96 53.7158
R1518 VDD2.n196 VDD2.n195 51.5793
R1519 VDD2.n196 VDD2.n98 48.4373
R1520 VDD2.n133 VDD2.n132 16.3895
R1521 VDD2.n32 VDD2.n31 16.3895
R1522 VDD2.n109 VDD2.n107 13.1884
R1523 VDD2.n77 VDD2.n8 13.1884
R1524 VDD2.n181 VDD2.n180 12.8005
R1525 VDD2.n177 VDD2.n176 12.8005
R1526 VDD2.n136 VDD2.n131 12.8005
R1527 VDD2.n35 VDD2.n30 12.8005
R1528 VDD2.n78 VDD2.n10 12.8005
R1529 VDD2.n82 VDD2.n81 12.8005
R1530 VDD2.n184 VDD2.n105 12.0247
R1531 VDD2.n173 VDD2.n110 12.0247
R1532 VDD2.n137 VDD2.n129 12.0247
R1533 VDD2.n36 VDD2.n28 12.0247
R1534 VDD2.n73 VDD2.n72 12.0247
R1535 VDD2.n85 VDD2.n6 12.0247
R1536 VDD2.n185 VDD2.n103 11.249
R1537 VDD2.n172 VDD2.n113 11.249
R1538 VDD2.n141 VDD2.n140 11.249
R1539 VDD2.n40 VDD2.n39 11.249
R1540 VDD2.n71 VDD2.n12 11.249
R1541 VDD2.n86 VDD2.n4 11.249
R1542 VDD2.n189 VDD2.n188 10.4732
R1543 VDD2.n169 VDD2.n168 10.4732
R1544 VDD2.n144 VDD2.n127 10.4732
R1545 VDD2.n43 VDD2.n26 10.4732
R1546 VDD2.n68 VDD2.n67 10.4732
R1547 VDD2.n90 VDD2.n89 10.4732
R1548 VDD2.n192 VDD2.n101 9.69747
R1549 VDD2.n165 VDD2.n115 9.69747
R1550 VDD2.n145 VDD2.n125 9.69747
R1551 VDD2.n44 VDD2.n24 9.69747
R1552 VDD2.n64 VDD2.n14 9.69747
R1553 VDD2.n93 VDD2.n2 9.69747
R1554 VDD2.n195 VDD2.n194 9.45567
R1555 VDD2.n96 VDD2.n95 9.45567
R1556 VDD2.n119 VDD2.n118 9.3005
R1557 VDD2.n162 VDD2.n161 9.3005
R1558 VDD2.n164 VDD2.n163 9.3005
R1559 VDD2.n115 VDD2.n114 9.3005
R1560 VDD2.n170 VDD2.n169 9.3005
R1561 VDD2.n172 VDD2.n171 9.3005
R1562 VDD2.n110 VDD2.n108 9.3005
R1563 VDD2.n178 VDD2.n177 9.3005
R1564 VDD2.n194 VDD2.n193 9.3005
R1565 VDD2.n101 VDD2.n100 9.3005
R1566 VDD2.n188 VDD2.n187 9.3005
R1567 VDD2.n186 VDD2.n185 9.3005
R1568 VDD2.n105 VDD2.n104 9.3005
R1569 VDD2.n180 VDD2.n179 9.3005
R1570 VDD2.n156 VDD2.n155 9.3005
R1571 VDD2.n154 VDD2.n153 9.3005
R1572 VDD2.n123 VDD2.n122 9.3005
R1573 VDD2.n148 VDD2.n147 9.3005
R1574 VDD2.n146 VDD2.n145 9.3005
R1575 VDD2.n127 VDD2.n126 9.3005
R1576 VDD2.n140 VDD2.n139 9.3005
R1577 VDD2.n138 VDD2.n137 9.3005
R1578 VDD2.n131 VDD2.n130 9.3005
R1579 VDD2.n95 VDD2.n94 9.3005
R1580 VDD2.n2 VDD2.n1 9.3005
R1581 VDD2.n89 VDD2.n88 9.3005
R1582 VDD2.n87 VDD2.n86 9.3005
R1583 VDD2.n6 VDD2.n5 9.3005
R1584 VDD2.n81 VDD2.n80 9.3005
R1585 VDD2.n53 VDD2.n52 9.3005
R1586 VDD2.n22 VDD2.n21 9.3005
R1587 VDD2.n47 VDD2.n46 9.3005
R1588 VDD2.n45 VDD2.n44 9.3005
R1589 VDD2.n26 VDD2.n25 9.3005
R1590 VDD2.n39 VDD2.n38 9.3005
R1591 VDD2.n37 VDD2.n36 9.3005
R1592 VDD2.n30 VDD2.n29 9.3005
R1593 VDD2.n55 VDD2.n54 9.3005
R1594 VDD2.n18 VDD2.n17 9.3005
R1595 VDD2.n61 VDD2.n60 9.3005
R1596 VDD2.n63 VDD2.n62 9.3005
R1597 VDD2.n14 VDD2.n13 9.3005
R1598 VDD2.n69 VDD2.n68 9.3005
R1599 VDD2.n71 VDD2.n70 9.3005
R1600 VDD2.n72 VDD2.n9 9.3005
R1601 VDD2.n79 VDD2.n78 9.3005
R1602 VDD2.n193 VDD2.n99 8.92171
R1603 VDD2.n164 VDD2.n117 8.92171
R1604 VDD2.n149 VDD2.n148 8.92171
R1605 VDD2.n48 VDD2.n47 8.92171
R1606 VDD2.n63 VDD2.n16 8.92171
R1607 VDD2.n94 VDD2.n0 8.92171
R1608 VDD2.n161 VDD2.n160 8.14595
R1609 VDD2.n152 VDD2.n123 8.14595
R1610 VDD2.n51 VDD2.n22 8.14595
R1611 VDD2.n60 VDD2.n59 8.14595
R1612 VDD2.n157 VDD2.n119 7.3702
R1613 VDD2.n153 VDD2.n121 7.3702
R1614 VDD2.n52 VDD2.n20 7.3702
R1615 VDD2.n56 VDD2.n18 7.3702
R1616 VDD2.n157 VDD2.n156 6.59444
R1617 VDD2.n156 VDD2.n121 6.59444
R1618 VDD2.n55 VDD2.n20 6.59444
R1619 VDD2.n56 VDD2.n55 6.59444
R1620 VDD2.n160 VDD2.n119 5.81868
R1621 VDD2.n153 VDD2.n152 5.81868
R1622 VDD2.n52 VDD2.n51 5.81868
R1623 VDD2.n59 VDD2.n18 5.81868
R1624 VDD2.n195 VDD2.n99 5.04292
R1625 VDD2.n161 VDD2.n117 5.04292
R1626 VDD2.n149 VDD2.n123 5.04292
R1627 VDD2.n48 VDD2.n22 5.04292
R1628 VDD2.n60 VDD2.n16 5.04292
R1629 VDD2.n96 VDD2.n0 5.04292
R1630 VDD2.n193 VDD2.n192 4.26717
R1631 VDD2.n165 VDD2.n164 4.26717
R1632 VDD2.n148 VDD2.n125 4.26717
R1633 VDD2.n47 VDD2.n24 4.26717
R1634 VDD2.n64 VDD2.n63 4.26717
R1635 VDD2.n94 VDD2.n93 4.26717
R1636 VDD2.n132 VDD2.n130 3.70982
R1637 VDD2.n31 VDD2.n29 3.70982
R1638 VDD2.n189 VDD2.n101 3.49141
R1639 VDD2.n168 VDD2.n115 3.49141
R1640 VDD2.n145 VDD2.n144 3.49141
R1641 VDD2.n44 VDD2.n43 3.49141
R1642 VDD2.n67 VDD2.n14 3.49141
R1643 VDD2.n90 VDD2.n2 3.49141
R1644 VDD2.n188 VDD2.n103 2.71565
R1645 VDD2.n169 VDD2.n113 2.71565
R1646 VDD2.n141 VDD2.n127 2.71565
R1647 VDD2.n40 VDD2.n26 2.71565
R1648 VDD2.n68 VDD2.n12 2.71565
R1649 VDD2.n89 VDD2.n4 2.71565
R1650 VDD2 VDD2.n196 2.2505
R1651 VDD2.n185 VDD2.n184 1.93989
R1652 VDD2.n173 VDD2.n172 1.93989
R1653 VDD2.n140 VDD2.n129 1.93989
R1654 VDD2.n39 VDD2.n28 1.93989
R1655 VDD2.n73 VDD2.n71 1.93989
R1656 VDD2.n86 VDD2.n85 1.93989
R1657 VDD2.n197 VDD2.t3 1.8411
R1658 VDD2.n197 VDD2.t0 1.8411
R1659 VDD2.n97 VDD2.t1 1.8411
R1660 VDD2.n97 VDD2.t5 1.8411
R1661 VDD2.n181 VDD2.n105 1.16414
R1662 VDD2.n176 VDD2.n110 1.16414
R1663 VDD2.n137 VDD2.n136 1.16414
R1664 VDD2.n36 VDD2.n35 1.16414
R1665 VDD2.n72 VDD2.n10 1.16414
R1666 VDD2.n82 VDD2.n6 1.16414
R1667 VDD2.n180 VDD2.n107 0.388379
R1668 VDD2.n177 VDD2.n109 0.388379
R1669 VDD2.n133 VDD2.n131 0.388379
R1670 VDD2.n32 VDD2.n30 0.388379
R1671 VDD2.n78 VDD2.n77 0.388379
R1672 VDD2.n81 VDD2.n8 0.388379
R1673 VDD2.n194 VDD2.n100 0.155672
R1674 VDD2.n187 VDD2.n100 0.155672
R1675 VDD2.n187 VDD2.n186 0.155672
R1676 VDD2.n186 VDD2.n104 0.155672
R1677 VDD2.n179 VDD2.n104 0.155672
R1678 VDD2.n179 VDD2.n178 0.155672
R1679 VDD2.n178 VDD2.n108 0.155672
R1680 VDD2.n171 VDD2.n108 0.155672
R1681 VDD2.n171 VDD2.n170 0.155672
R1682 VDD2.n170 VDD2.n114 0.155672
R1683 VDD2.n163 VDD2.n114 0.155672
R1684 VDD2.n163 VDD2.n162 0.155672
R1685 VDD2.n162 VDD2.n118 0.155672
R1686 VDD2.n155 VDD2.n118 0.155672
R1687 VDD2.n155 VDD2.n154 0.155672
R1688 VDD2.n154 VDD2.n122 0.155672
R1689 VDD2.n147 VDD2.n122 0.155672
R1690 VDD2.n147 VDD2.n146 0.155672
R1691 VDD2.n146 VDD2.n126 0.155672
R1692 VDD2.n139 VDD2.n126 0.155672
R1693 VDD2.n139 VDD2.n138 0.155672
R1694 VDD2.n138 VDD2.n130 0.155672
R1695 VDD2.n37 VDD2.n29 0.155672
R1696 VDD2.n38 VDD2.n37 0.155672
R1697 VDD2.n38 VDD2.n25 0.155672
R1698 VDD2.n45 VDD2.n25 0.155672
R1699 VDD2.n46 VDD2.n45 0.155672
R1700 VDD2.n46 VDD2.n21 0.155672
R1701 VDD2.n53 VDD2.n21 0.155672
R1702 VDD2.n54 VDD2.n53 0.155672
R1703 VDD2.n54 VDD2.n17 0.155672
R1704 VDD2.n61 VDD2.n17 0.155672
R1705 VDD2.n62 VDD2.n61 0.155672
R1706 VDD2.n62 VDD2.n13 0.155672
R1707 VDD2.n69 VDD2.n13 0.155672
R1708 VDD2.n70 VDD2.n69 0.155672
R1709 VDD2.n70 VDD2.n9 0.155672
R1710 VDD2.n79 VDD2.n9 0.155672
R1711 VDD2.n80 VDD2.n79 0.155672
R1712 VDD2.n80 VDD2.n5 0.155672
R1713 VDD2.n87 VDD2.n5 0.155672
R1714 VDD2.n88 VDD2.n87 0.155672
R1715 VDD2.n88 VDD2.n1 0.155672
R1716 VDD2.n95 VDD2.n1 0.155672
R1717 VTAIL.n394 VTAIL.n302 756.745
R1718 VTAIL.n94 VTAIL.n2 756.745
R1719 VTAIL.n296 VTAIL.n204 756.745
R1720 VTAIL.n196 VTAIL.n104 756.745
R1721 VTAIL.n335 VTAIL.n334 585
R1722 VTAIL.n337 VTAIL.n336 585
R1723 VTAIL.n330 VTAIL.n329 585
R1724 VTAIL.n343 VTAIL.n342 585
R1725 VTAIL.n345 VTAIL.n344 585
R1726 VTAIL.n326 VTAIL.n325 585
R1727 VTAIL.n351 VTAIL.n350 585
R1728 VTAIL.n353 VTAIL.n352 585
R1729 VTAIL.n322 VTAIL.n321 585
R1730 VTAIL.n359 VTAIL.n358 585
R1731 VTAIL.n361 VTAIL.n360 585
R1732 VTAIL.n318 VTAIL.n317 585
R1733 VTAIL.n367 VTAIL.n366 585
R1734 VTAIL.n369 VTAIL.n368 585
R1735 VTAIL.n314 VTAIL.n313 585
R1736 VTAIL.n376 VTAIL.n375 585
R1737 VTAIL.n377 VTAIL.n312 585
R1738 VTAIL.n379 VTAIL.n378 585
R1739 VTAIL.n310 VTAIL.n309 585
R1740 VTAIL.n385 VTAIL.n384 585
R1741 VTAIL.n387 VTAIL.n386 585
R1742 VTAIL.n306 VTAIL.n305 585
R1743 VTAIL.n393 VTAIL.n392 585
R1744 VTAIL.n395 VTAIL.n394 585
R1745 VTAIL.n35 VTAIL.n34 585
R1746 VTAIL.n37 VTAIL.n36 585
R1747 VTAIL.n30 VTAIL.n29 585
R1748 VTAIL.n43 VTAIL.n42 585
R1749 VTAIL.n45 VTAIL.n44 585
R1750 VTAIL.n26 VTAIL.n25 585
R1751 VTAIL.n51 VTAIL.n50 585
R1752 VTAIL.n53 VTAIL.n52 585
R1753 VTAIL.n22 VTAIL.n21 585
R1754 VTAIL.n59 VTAIL.n58 585
R1755 VTAIL.n61 VTAIL.n60 585
R1756 VTAIL.n18 VTAIL.n17 585
R1757 VTAIL.n67 VTAIL.n66 585
R1758 VTAIL.n69 VTAIL.n68 585
R1759 VTAIL.n14 VTAIL.n13 585
R1760 VTAIL.n76 VTAIL.n75 585
R1761 VTAIL.n77 VTAIL.n12 585
R1762 VTAIL.n79 VTAIL.n78 585
R1763 VTAIL.n10 VTAIL.n9 585
R1764 VTAIL.n85 VTAIL.n84 585
R1765 VTAIL.n87 VTAIL.n86 585
R1766 VTAIL.n6 VTAIL.n5 585
R1767 VTAIL.n93 VTAIL.n92 585
R1768 VTAIL.n95 VTAIL.n94 585
R1769 VTAIL.n297 VTAIL.n296 585
R1770 VTAIL.n295 VTAIL.n294 585
R1771 VTAIL.n208 VTAIL.n207 585
R1772 VTAIL.n289 VTAIL.n288 585
R1773 VTAIL.n287 VTAIL.n286 585
R1774 VTAIL.n212 VTAIL.n211 585
R1775 VTAIL.n216 VTAIL.n214 585
R1776 VTAIL.n281 VTAIL.n280 585
R1777 VTAIL.n279 VTAIL.n278 585
R1778 VTAIL.n218 VTAIL.n217 585
R1779 VTAIL.n273 VTAIL.n272 585
R1780 VTAIL.n271 VTAIL.n270 585
R1781 VTAIL.n222 VTAIL.n221 585
R1782 VTAIL.n265 VTAIL.n264 585
R1783 VTAIL.n263 VTAIL.n262 585
R1784 VTAIL.n226 VTAIL.n225 585
R1785 VTAIL.n257 VTAIL.n256 585
R1786 VTAIL.n255 VTAIL.n254 585
R1787 VTAIL.n230 VTAIL.n229 585
R1788 VTAIL.n249 VTAIL.n248 585
R1789 VTAIL.n247 VTAIL.n246 585
R1790 VTAIL.n234 VTAIL.n233 585
R1791 VTAIL.n241 VTAIL.n240 585
R1792 VTAIL.n239 VTAIL.n238 585
R1793 VTAIL.n197 VTAIL.n196 585
R1794 VTAIL.n195 VTAIL.n194 585
R1795 VTAIL.n108 VTAIL.n107 585
R1796 VTAIL.n189 VTAIL.n188 585
R1797 VTAIL.n187 VTAIL.n186 585
R1798 VTAIL.n112 VTAIL.n111 585
R1799 VTAIL.n116 VTAIL.n114 585
R1800 VTAIL.n181 VTAIL.n180 585
R1801 VTAIL.n179 VTAIL.n178 585
R1802 VTAIL.n118 VTAIL.n117 585
R1803 VTAIL.n173 VTAIL.n172 585
R1804 VTAIL.n171 VTAIL.n170 585
R1805 VTAIL.n122 VTAIL.n121 585
R1806 VTAIL.n165 VTAIL.n164 585
R1807 VTAIL.n163 VTAIL.n162 585
R1808 VTAIL.n126 VTAIL.n125 585
R1809 VTAIL.n157 VTAIL.n156 585
R1810 VTAIL.n155 VTAIL.n154 585
R1811 VTAIL.n130 VTAIL.n129 585
R1812 VTAIL.n149 VTAIL.n148 585
R1813 VTAIL.n147 VTAIL.n146 585
R1814 VTAIL.n134 VTAIL.n133 585
R1815 VTAIL.n141 VTAIL.n140 585
R1816 VTAIL.n139 VTAIL.n138 585
R1817 VTAIL.n333 VTAIL.t6 327.466
R1818 VTAIL.n33 VTAIL.t2 327.466
R1819 VTAIL.n237 VTAIL.t0 327.466
R1820 VTAIL.n137 VTAIL.t10 327.466
R1821 VTAIL.n336 VTAIL.n335 171.744
R1822 VTAIL.n336 VTAIL.n329 171.744
R1823 VTAIL.n343 VTAIL.n329 171.744
R1824 VTAIL.n344 VTAIL.n343 171.744
R1825 VTAIL.n344 VTAIL.n325 171.744
R1826 VTAIL.n351 VTAIL.n325 171.744
R1827 VTAIL.n352 VTAIL.n351 171.744
R1828 VTAIL.n352 VTAIL.n321 171.744
R1829 VTAIL.n359 VTAIL.n321 171.744
R1830 VTAIL.n360 VTAIL.n359 171.744
R1831 VTAIL.n360 VTAIL.n317 171.744
R1832 VTAIL.n367 VTAIL.n317 171.744
R1833 VTAIL.n368 VTAIL.n367 171.744
R1834 VTAIL.n368 VTAIL.n313 171.744
R1835 VTAIL.n376 VTAIL.n313 171.744
R1836 VTAIL.n377 VTAIL.n376 171.744
R1837 VTAIL.n378 VTAIL.n377 171.744
R1838 VTAIL.n378 VTAIL.n309 171.744
R1839 VTAIL.n385 VTAIL.n309 171.744
R1840 VTAIL.n386 VTAIL.n385 171.744
R1841 VTAIL.n386 VTAIL.n305 171.744
R1842 VTAIL.n393 VTAIL.n305 171.744
R1843 VTAIL.n394 VTAIL.n393 171.744
R1844 VTAIL.n36 VTAIL.n35 171.744
R1845 VTAIL.n36 VTAIL.n29 171.744
R1846 VTAIL.n43 VTAIL.n29 171.744
R1847 VTAIL.n44 VTAIL.n43 171.744
R1848 VTAIL.n44 VTAIL.n25 171.744
R1849 VTAIL.n51 VTAIL.n25 171.744
R1850 VTAIL.n52 VTAIL.n51 171.744
R1851 VTAIL.n52 VTAIL.n21 171.744
R1852 VTAIL.n59 VTAIL.n21 171.744
R1853 VTAIL.n60 VTAIL.n59 171.744
R1854 VTAIL.n60 VTAIL.n17 171.744
R1855 VTAIL.n67 VTAIL.n17 171.744
R1856 VTAIL.n68 VTAIL.n67 171.744
R1857 VTAIL.n68 VTAIL.n13 171.744
R1858 VTAIL.n76 VTAIL.n13 171.744
R1859 VTAIL.n77 VTAIL.n76 171.744
R1860 VTAIL.n78 VTAIL.n77 171.744
R1861 VTAIL.n78 VTAIL.n9 171.744
R1862 VTAIL.n85 VTAIL.n9 171.744
R1863 VTAIL.n86 VTAIL.n85 171.744
R1864 VTAIL.n86 VTAIL.n5 171.744
R1865 VTAIL.n93 VTAIL.n5 171.744
R1866 VTAIL.n94 VTAIL.n93 171.744
R1867 VTAIL.n296 VTAIL.n295 171.744
R1868 VTAIL.n295 VTAIL.n207 171.744
R1869 VTAIL.n288 VTAIL.n207 171.744
R1870 VTAIL.n288 VTAIL.n287 171.744
R1871 VTAIL.n287 VTAIL.n211 171.744
R1872 VTAIL.n216 VTAIL.n211 171.744
R1873 VTAIL.n280 VTAIL.n216 171.744
R1874 VTAIL.n280 VTAIL.n279 171.744
R1875 VTAIL.n279 VTAIL.n217 171.744
R1876 VTAIL.n272 VTAIL.n217 171.744
R1877 VTAIL.n272 VTAIL.n271 171.744
R1878 VTAIL.n271 VTAIL.n221 171.744
R1879 VTAIL.n264 VTAIL.n221 171.744
R1880 VTAIL.n264 VTAIL.n263 171.744
R1881 VTAIL.n263 VTAIL.n225 171.744
R1882 VTAIL.n256 VTAIL.n225 171.744
R1883 VTAIL.n256 VTAIL.n255 171.744
R1884 VTAIL.n255 VTAIL.n229 171.744
R1885 VTAIL.n248 VTAIL.n229 171.744
R1886 VTAIL.n248 VTAIL.n247 171.744
R1887 VTAIL.n247 VTAIL.n233 171.744
R1888 VTAIL.n240 VTAIL.n233 171.744
R1889 VTAIL.n240 VTAIL.n239 171.744
R1890 VTAIL.n196 VTAIL.n195 171.744
R1891 VTAIL.n195 VTAIL.n107 171.744
R1892 VTAIL.n188 VTAIL.n107 171.744
R1893 VTAIL.n188 VTAIL.n187 171.744
R1894 VTAIL.n187 VTAIL.n111 171.744
R1895 VTAIL.n116 VTAIL.n111 171.744
R1896 VTAIL.n180 VTAIL.n116 171.744
R1897 VTAIL.n180 VTAIL.n179 171.744
R1898 VTAIL.n179 VTAIL.n117 171.744
R1899 VTAIL.n172 VTAIL.n117 171.744
R1900 VTAIL.n172 VTAIL.n171 171.744
R1901 VTAIL.n171 VTAIL.n121 171.744
R1902 VTAIL.n164 VTAIL.n121 171.744
R1903 VTAIL.n164 VTAIL.n163 171.744
R1904 VTAIL.n163 VTAIL.n125 171.744
R1905 VTAIL.n156 VTAIL.n125 171.744
R1906 VTAIL.n156 VTAIL.n155 171.744
R1907 VTAIL.n155 VTAIL.n129 171.744
R1908 VTAIL.n148 VTAIL.n129 171.744
R1909 VTAIL.n148 VTAIL.n147 171.744
R1910 VTAIL.n147 VTAIL.n133 171.744
R1911 VTAIL.n140 VTAIL.n133 171.744
R1912 VTAIL.n140 VTAIL.n139 171.744
R1913 VTAIL.n335 VTAIL.t6 85.8723
R1914 VTAIL.n35 VTAIL.t2 85.8723
R1915 VTAIL.n239 VTAIL.t0 85.8723
R1916 VTAIL.n139 VTAIL.t10 85.8723
R1917 VTAIL.n203 VTAIL.n202 55.0586
R1918 VTAIL.n103 VTAIL.n102 55.0586
R1919 VTAIL.n1 VTAIL.n0 55.0584
R1920 VTAIL.n101 VTAIL.n100 55.0584
R1921 VTAIL.n399 VTAIL.n398 34.9005
R1922 VTAIL.n99 VTAIL.n98 34.9005
R1923 VTAIL.n301 VTAIL.n300 34.9005
R1924 VTAIL.n201 VTAIL.n200 34.9005
R1925 VTAIL.n103 VTAIL.n101 33.4358
R1926 VTAIL.n399 VTAIL.n301 30.5134
R1927 VTAIL.n334 VTAIL.n333 16.3895
R1928 VTAIL.n34 VTAIL.n33 16.3895
R1929 VTAIL.n238 VTAIL.n237 16.3895
R1930 VTAIL.n138 VTAIL.n137 16.3895
R1931 VTAIL.n379 VTAIL.n310 13.1884
R1932 VTAIL.n79 VTAIL.n10 13.1884
R1933 VTAIL.n214 VTAIL.n212 13.1884
R1934 VTAIL.n114 VTAIL.n112 13.1884
R1935 VTAIL.n337 VTAIL.n332 12.8005
R1936 VTAIL.n380 VTAIL.n312 12.8005
R1937 VTAIL.n384 VTAIL.n383 12.8005
R1938 VTAIL.n37 VTAIL.n32 12.8005
R1939 VTAIL.n80 VTAIL.n12 12.8005
R1940 VTAIL.n84 VTAIL.n83 12.8005
R1941 VTAIL.n286 VTAIL.n285 12.8005
R1942 VTAIL.n282 VTAIL.n281 12.8005
R1943 VTAIL.n241 VTAIL.n236 12.8005
R1944 VTAIL.n186 VTAIL.n185 12.8005
R1945 VTAIL.n182 VTAIL.n181 12.8005
R1946 VTAIL.n141 VTAIL.n136 12.8005
R1947 VTAIL.n338 VTAIL.n330 12.0247
R1948 VTAIL.n375 VTAIL.n374 12.0247
R1949 VTAIL.n387 VTAIL.n308 12.0247
R1950 VTAIL.n38 VTAIL.n30 12.0247
R1951 VTAIL.n75 VTAIL.n74 12.0247
R1952 VTAIL.n87 VTAIL.n8 12.0247
R1953 VTAIL.n289 VTAIL.n210 12.0247
R1954 VTAIL.n278 VTAIL.n215 12.0247
R1955 VTAIL.n242 VTAIL.n234 12.0247
R1956 VTAIL.n189 VTAIL.n110 12.0247
R1957 VTAIL.n178 VTAIL.n115 12.0247
R1958 VTAIL.n142 VTAIL.n134 12.0247
R1959 VTAIL.n342 VTAIL.n341 11.249
R1960 VTAIL.n373 VTAIL.n314 11.249
R1961 VTAIL.n388 VTAIL.n306 11.249
R1962 VTAIL.n42 VTAIL.n41 11.249
R1963 VTAIL.n73 VTAIL.n14 11.249
R1964 VTAIL.n88 VTAIL.n6 11.249
R1965 VTAIL.n290 VTAIL.n208 11.249
R1966 VTAIL.n277 VTAIL.n218 11.249
R1967 VTAIL.n246 VTAIL.n245 11.249
R1968 VTAIL.n190 VTAIL.n108 11.249
R1969 VTAIL.n177 VTAIL.n118 11.249
R1970 VTAIL.n146 VTAIL.n145 11.249
R1971 VTAIL.n345 VTAIL.n328 10.4732
R1972 VTAIL.n370 VTAIL.n369 10.4732
R1973 VTAIL.n392 VTAIL.n391 10.4732
R1974 VTAIL.n45 VTAIL.n28 10.4732
R1975 VTAIL.n70 VTAIL.n69 10.4732
R1976 VTAIL.n92 VTAIL.n91 10.4732
R1977 VTAIL.n294 VTAIL.n293 10.4732
R1978 VTAIL.n274 VTAIL.n273 10.4732
R1979 VTAIL.n249 VTAIL.n232 10.4732
R1980 VTAIL.n194 VTAIL.n193 10.4732
R1981 VTAIL.n174 VTAIL.n173 10.4732
R1982 VTAIL.n149 VTAIL.n132 10.4732
R1983 VTAIL.n346 VTAIL.n326 9.69747
R1984 VTAIL.n366 VTAIL.n316 9.69747
R1985 VTAIL.n395 VTAIL.n304 9.69747
R1986 VTAIL.n46 VTAIL.n26 9.69747
R1987 VTAIL.n66 VTAIL.n16 9.69747
R1988 VTAIL.n95 VTAIL.n4 9.69747
R1989 VTAIL.n297 VTAIL.n206 9.69747
R1990 VTAIL.n270 VTAIL.n220 9.69747
R1991 VTAIL.n250 VTAIL.n230 9.69747
R1992 VTAIL.n197 VTAIL.n106 9.69747
R1993 VTAIL.n170 VTAIL.n120 9.69747
R1994 VTAIL.n150 VTAIL.n130 9.69747
R1995 VTAIL.n398 VTAIL.n397 9.45567
R1996 VTAIL.n98 VTAIL.n97 9.45567
R1997 VTAIL.n300 VTAIL.n299 9.45567
R1998 VTAIL.n200 VTAIL.n199 9.45567
R1999 VTAIL.n397 VTAIL.n396 9.3005
R2000 VTAIL.n304 VTAIL.n303 9.3005
R2001 VTAIL.n391 VTAIL.n390 9.3005
R2002 VTAIL.n389 VTAIL.n388 9.3005
R2003 VTAIL.n308 VTAIL.n307 9.3005
R2004 VTAIL.n383 VTAIL.n382 9.3005
R2005 VTAIL.n355 VTAIL.n354 9.3005
R2006 VTAIL.n324 VTAIL.n323 9.3005
R2007 VTAIL.n349 VTAIL.n348 9.3005
R2008 VTAIL.n347 VTAIL.n346 9.3005
R2009 VTAIL.n328 VTAIL.n327 9.3005
R2010 VTAIL.n341 VTAIL.n340 9.3005
R2011 VTAIL.n339 VTAIL.n338 9.3005
R2012 VTAIL.n332 VTAIL.n331 9.3005
R2013 VTAIL.n357 VTAIL.n356 9.3005
R2014 VTAIL.n320 VTAIL.n319 9.3005
R2015 VTAIL.n363 VTAIL.n362 9.3005
R2016 VTAIL.n365 VTAIL.n364 9.3005
R2017 VTAIL.n316 VTAIL.n315 9.3005
R2018 VTAIL.n371 VTAIL.n370 9.3005
R2019 VTAIL.n373 VTAIL.n372 9.3005
R2020 VTAIL.n374 VTAIL.n311 9.3005
R2021 VTAIL.n381 VTAIL.n380 9.3005
R2022 VTAIL.n97 VTAIL.n96 9.3005
R2023 VTAIL.n4 VTAIL.n3 9.3005
R2024 VTAIL.n91 VTAIL.n90 9.3005
R2025 VTAIL.n89 VTAIL.n88 9.3005
R2026 VTAIL.n8 VTAIL.n7 9.3005
R2027 VTAIL.n83 VTAIL.n82 9.3005
R2028 VTAIL.n55 VTAIL.n54 9.3005
R2029 VTAIL.n24 VTAIL.n23 9.3005
R2030 VTAIL.n49 VTAIL.n48 9.3005
R2031 VTAIL.n47 VTAIL.n46 9.3005
R2032 VTAIL.n28 VTAIL.n27 9.3005
R2033 VTAIL.n41 VTAIL.n40 9.3005
R2034 VTAIL.n39 VTAIL.n38 9.3005
R2035 VTAIL.n32 VTAIL.n31 9.3005
R2036 VTAIL.n57 VTAIL.n56 9.3005
R2037 VTAIL.n20 VTAIL.n19 9.3005
R2038 VTAIL.n63 VTAIL.n62 9.3005
R2039 VTAIL.n65 VTAIL.n64 9.3005
R2040 VTAIL.n16 VTAIL.n15 9.3005
R2041 VTAIL.n71 VTAIL.n70 9.3005
R2042 VTAIL.n73 VTAIL.n72 9.3005
R2043 VTAIL.n74 VTAIL.n11 9.3005
R2044 VTAIL.n81 VTAIL.n80 9.3005
R2045 VTAIL.n224 VTAIL.n223 9.3005
R2046 VTAIL.n267 VTAIL.n266 9.3005
R2047 VTAIL.n269 VTAIL.n268 9.3005
R2048 VTAIL.n220 VTAIL.n219 9.3005
R2049 VTAIL.n275 VTAIL.n274 9.3005
R2050 VTAIL.n277 VTAIL.n276 9.3005
R2051 VTAIL.n215 VTAIL.n213 9.3005
R2052 VTAIL.n283 VTAIL.n282 9.3005
R2053 VTAIL.n299 VTAIL.n298 9.3005
R2054 VTAIL.n206 VTAIL.n205 9.3005
R2055 VTAIL.n293 VTAIL.n292 9.3005
R2056 VTAIL.n291 VTAIL.n290 9.3005
R2057 VTAIL.n210 VTAIL.n209 9.3005
R2058 VTAIL.n285 VTAIL.n284 9.3005
R2059 VTAIL.n261 VTAIL.n260 9.3005
R2060 VTAIL.n259 VTAIL.n258 9.3005
R2061 VTAIL.n228 VTAIL.n227 9.3005
R2062 VTAIL.n253 VTAIL.n252 9.3005
R2063 VTAIL.n251 VTAIL.n250 9.3005
R2064 VTAIL.n232 VTAIL.n231 9.3005
R2065 VTAIL.n245 VTAIL.n244 9.3005
R2066 VTAIL.n243 VTAIL.n242 9.3005
R2067 VTAIL.n236 VTAIL.n235 9.3005
R2068 VTAIL.n124 VTAIL.n123 9.3005
R2069 VTAIL.n167 VTAIL.n166 9.3005
R2070 VTAIL.n169 VTAIL.n168 9.3005
R2071 VTAIL.n120 VTAIL.n119 9.3005
R2072 VTAIL.n175 VTAIL.n174 9.3005
R2073 VTAIL.n177 VTAIL.n176 9.3005
R2074 VTAIL.n115 VTAIL.n113 9.3005
R2075 VTAIL.n183 VTAIL.n182 9.3005
R2076 VTAIL.n199 VTAIL.n198 9.3005
R2077 VTAIL.n106 VTAIL.n105 9.3005
R2078 VTAIL.n193 VTAIL.n192 9.3005
R2079 VTAIL.n191 VTAIL.n190 9.3005
R2080 VTAIL.n110 VTAIL.n109 9.3005
R2081 VTAIL.n185 VTAIL.n184 9.3005
R2082 VTAIL.n161 VTAIL.n160 9.3005
R2083 VTAIL.n159 VTAIL.n158 9.3005
R2084 VTAIL.n128 VTAIL.n127 9.3005
R2085 VTAIL.n153 VTAIL.n152 9.3005
R2086 VTAIL.n151 VTAIL.n150 9.3005
R2087 VTAIL.n132 VTAIL.n131 9.3005
R2088 VTAIL.n145 VTAIL.n144 9.3005
R2089 VTAIL.n143 VTAIL.n142 9.3005
R2090 VTAIL.n136 VTAIL.n135 9.3005
R2091 VTAIL.n350 VTAIL.n349 8.92171
R2092 VTAIL.n365 VTAIL.n318 8.92171
R2093 VTAIL.n396 VTAIL.n302 8.92171
R2094 VTAIL.n50 VTAIL.n49 8.92171
R2095 VTAIL.n65 VTAIL.n18 8.92171
R2096 VTAIL.n96 VTAIL.n2 8.92171
R2097 VTAIL.n298 VTAIL.n204 8.92171
R2098 VTAIL.n269 VTAIL.n222 8.92171
R2099 VTAIL.n254 VTAIL.n253 8.92171
R2100 VTAIL.n198 VTAIL.n104 8.92171
R2101 VTAIL.n169 VTAIL.n122 8.92171
R2102 VTAIL.n154 VTAIL.n153 8.92171
R2103 VTAIL.n353 VTAIL.n324 8.14595
R2104 VTAIL.n362 VTAIL.n361 8.14595
R2105 VTAIL.n53 VTAIL.n24 8.14595
R2106 VTAIL.n62 VTAIL.n61 8.14595
R2107 VTAIL.n266 VTAIL.n265 8.14595
R2108 VTAIL.n257 VTAIL.n228 8.14595
R2109 VTAIL.n166 VTAIL.n165 8.14595
R2110 VTAIL.n157 VTAIL.n128 8.14595
R2111 VTAIL.n354 VTAIL.n322 7.3702
R2112 VTAIL.n358 VTAIL.n320 7.3702
R2113 VTAIL.n54 VTAIL.n22 7.3702
R2114 VTAIL.n58 VTAIL.n20 7.3702
R2115 VTAIL.n262 VTAIL.n224 7.3702
R2116 VTAIL.n258 VTAIL.n226 7.3702
R2117 VTAIL.n162 VTAIL.n124 7.3702
R2118 VTAIL.n158 VTAIL.n126 7.3702
R2119 VTAIL.n357 VTAIL.n322 6.59444
R2120 VTAIL.n358 VTAIL.n357 6.59444
R2121 VTAIL.n57 VTAIL.n22 6.59444
R2122 VTAIL.n58 VTAIL.n57 6.59444
R2123 VTAIL.n262 VTAIL.n261 6.59444
R2124 VTAIL.n261 VTAIL.n226 6.59444
R2125 VTAIL.n162 VTAIL.n161 6.59444
R2126 VTAIL.n161 VTAIL.n126 6.59444
R2127 VTAIL.n354 VTAIL.n353 5.81868
R2128 VTAIL.n361 VTAIL.n320 5.81868
R2129 VTAIL.n54 VTAIL.n53 5.81868
R2130 VTAIL.n61 VTAIL.n20 5.81868
R2131 VTAIL.n265 VTAIL.n224 5.81868
R2132 VTAIL.n258 VTAIL.n257 5.81868
R2133 VTAIL.n165 VTAIL.n124 5.81868
R2134 VTAIL.n158 VTAIL.n157 5.81868
R2135 VTAIL.n350 VTAIL.n324 5.04292
R2136 VTAIL.n362 VTAIL.n318 5.04292
R2137 VTAIL.n398 VTAIL.n302 5.04292
R2138 VTAIL.n50 VTAIL.n24 5.04292
R2139 VTAIL.n62 VTAIL.n18 5.04292
R2140 VTAIL.n98 VTAIL.n2 5.04292
R2141 VTAIL.n300 VTAIL.n204 5.04292
R2142 VTAIL.n266 VTAIL.n222 5.04292
R2143 VTAIL.n254 VTAIL.n228 5.04292
R2144 VTAIL.n200 VTAIL.n104 5.04292
R2145 VTAIL.n166 VTAIL.n122 5.04292
R2146 VTAIL.n154 VTAIL.n128 5.04292
R2147 VTAIL.n349 VTAIL.n326 4.26717
R2148 VTAIL.n366 VTAIL.n365 4.26717
R2149 VTAIL.n396 VTAIL.n395 4.26717
R2150 VTAIL.n49 VTAIL.n26 4.26717
R2151 VTAIL.n66 VTAIL.n65 4.26717
R2152 VTAIL.n96 VTAIL.n95 4.26717
R2153 VTAIL.n298 VTAIL.n297 4.26717
R2154 VTAIL.n270 VTAIL.n269 4.26717
R2155 VTAIL.n253 VTAIL.n230 4.26717
R2156 VTAIL.n198 VTAIL.n197 4.26717
R2157 VTAIL.n170 VTAIL.n169 4.26717
R2158 VTAIL.n153 VTAIL.n130 4.26717
R2159 VTAIL.n333 VTAIL.n331 3.70982
R2160 VTAIL.n33 VTAIL.n31 3.70982
R2161 VTAIL.n237 VTAIL.n235 3.70982
R2162 VTAIL.n137 VTAIL.n135 3.70982
R2163 VTAIL.n346 VTAIL.n345 3.49141
R2164 VTAIL.n369 VTAIL.n316 3.49141
R2165 VTAIL.n392 VTAIL.n304 3.49141
R2166 VTAIL.n46 VTAIL.n45 3.49141
R2167 VTAIL.n69 VTAIL.n16 3.49141
R2168 VTAIL.n92 VTAIL.n4 3.49141
R2169 VTAIL.n294 VTAIL.n206 3.49141
R2170 VTAIL.n273 VTAIL.n220 3.49141
R2171 VTAIL.n250 VTAIL.n249 3.49141
R2172 VTAIL.n194 VTAIL.n106 3.49141
R2173 VTAIL.n173 VTAIL.n120 3.49141
R2174 VTAIL.n150 VTAIL.n149 3.49141
R2175 VTAIL.n201 VTAIL.n103 2.92291
R2176 VTAIL.n301 VTAIL.n203 2.92291
R2177 VTAIL.n101 VTAIL.n99 2.92291
R2178 VTAIL.n342 VTAIL.n328 2.71565
R2179 VTAIL.n370 VTAIL.n314 2.71565
R2180 VTAIL.n391 VTAIL.n306 2.71565
R2181 VTAIL.n42 VTAIL.n28 2.71565
R2182 VTAIL.n70 VTAIL.n14 2.71565
R2183 VTAIL.n91 VTAIL.n6 2.71565
R2184 VTAIL.n293 VTAIL.n208 2.71565
R2185 VTAIL.n274 VTAIL.n218 2.71565
R2186 VTAIL.n246 VTAIL.n232 2.71565
R2187 VTAIL.n193 VTAIL.n108 2.71565
R2188 VTAIL.n174 VTAIL.n118 2.71565
R2189 VTAIL.n146 VTAIL.n132 2.71565
R2190 VTAIL VTAIL.n399 2.13412
R2191 VTAIL.n341 VTAIL.n330 1.93989
R2192 VTAIL.n375 VTAIL.n373 1.93989
R2193 VTAIL.n388 VTAIL.n387 1.93989
R2194 VTAIL.n41 VTAIL.n30 1.93989
R2195 VTAIL.n75 VTAIL.n73 1.93989
R2196 VTAIL.n88 VTAIL.n87 1.93989
R2197 VTAIL.n290 VTAIL.n289 1.93989
R2198 VTAIL.n278 VTAIL.n277 1.93989
R2199 VTAIL.n245 VTAIL.n234 1.93989
R2200 VTAIL.n190 VTAIL.n189 1.93989
R2201 VTAIL.n178 VTAIL.n177 1.93989
R2202 VTAIL.n145 VTAIL.n134 1.93989
R2203 VTAIL.n203 VTAIL.n201 1.93153
R2204 VTAIL.n99 VTAIL.n1 1.93153
R2205 VTAIL.n0 VTAIL.t7 1.8411
R2206 VTAIL.n0 VTAIL.t11 1.8411
R2207 VTAIL.n100 VTAIL.t1 1.8411
R2208 VTAIL.n100 VTAIL.t3 1.8411
R2209 VTAIL.n202 VTAIL.t4 1.8411
R2210 VTAIL.n202 VTAIL.t5 1.8411
R2211 VTAIL.n102 VTAIL.t9 1.8411
R2212 VTAIL.n102 VTAIL.t8 1.8411
R2213 VTAIL.n338 VTAIL.n337 1.16414
R2214 VTAIL.n374 VTAIL.n312 1.16414
R2215 VTAIL.n384 VTAIL.n308 1.16414
R2216 VTAIL.n38 VTAIL.n37 1.16414
R2217 VTAIL.n74 VTAIL.n12 1.16414
R2218 VTAIL.n84 VTAIL.n8 1.16414
R2219 VTAIL.n286 VTAIL.n210 1.16414
R2220 VTAIL.n281 VTAIL.n215 1.16414
R2221 VTAIL.n242 VTAIL.n241 1.16414
R2222 VTAIL.n186 VTAIL.n110 1.16414
R2223 VTAIL.n181 VTAIL.n115 1.16414
R2224 VTAIL.n142 VTAIL.n141 1.16414
R2225 VTAIL VTAIL.n1 0.789293
R2226 VTAIL.n334 VTAIL.n332 0.388379
R2227 VTAIL.n380 VTAIL.n379 0.388379
R2228 VTAIL.n383 VTAIL.n310 0.388379
R2229 VTAIL.n34 VTAIL.n32 0.388379
R2230 VTAIL.n80 VTAIL.n79 0.388379
R2231 VTAIL.n83 VTAIL.n10 0.388379
R2232 VTAIL.n285 VTAIL.n212 0.388379
R2233 VTAIL.n282 VTAIL.n214 0.388379
R2234 VTAIL.n238 VTAIL.n236 0.388379
R2235 VTAIL.n185 VTAIL.n112 0.388379
R2236 VTAIL.n182 VTAIL.n114 0.388379
R2237 VTAIL.n138 VTAIL.n136 0.388379
R2238 VTAIL.n339 VTAIL.n331 0.155672
R2239 VTAIL.n340 VTAIL.n339 0.155672
R2240 VTAIL.n340 VTAIL.n327 0.155672
R2241 VTAIL.n347 VTAIL.n327 0.155672
R2242 VTAIL.n348 VTAIL.n347 0.155672
R2243 VTAIL.n348 VTAIL.n323 0.155672
R2244 VTAIL.n355 VTAIL.n323 0.155672
R2245 VTAIL.n356 VTAIL.n355 0.155672
R2246 VTAIL.n356 VTAIL.n319 0.155672
R2247 VTAIL.n363 VTAIL.n319 0.155672
R2248 VTAIL.n364 VTAIL.n363 0.155672
R2249 VTAIL.n364 VTAIL.n315 0.155672
R2250 VTAIL.n371 VTAIL.n315 0.155672
R2251 VTAIL.n372 VTAIL.n371 0.155672
R2252 VTAIL.n372 VTAIL.n311 0.155672
R2253 VTAIL.n381 VTAIL.n311 0.155672
R2254 VTAIL.n382 VTAIL.n381 0.155672
R2255 VTAIL.n382 VTAIL.n307 0.155672
R2256 VTAIL.n389 VTAIL.n307 0.155672
R2257 VTAIL.n390 VTAIL.n389 0.155672
R2258 VTAIL.n390 VTAIL.n303 0.155672
R2259 VTAIL.n397 VTAIL.n303 0.155672
R2260 VTAIL.n39 VTAIL.n31 0.155672
R2261 VTAIL.n40 VTAIL.n39 0.155672
R2262 VTAIL.n40 VTAIL.n27 0.155672
R2263 VTAIL.n47 VTAIL.n27 0.155672
R2264 VTAIL.n48 VTAIL.n47 0.155672
R2265 VTAIL.n48 VTAIL.n23 0.155672
R2266 VTAIL.n55 VTAIL.n23 0.155672
R2267 VTAIL.n56 VTAIL.n55 0.155672
R2268 VTAIL.n56 VTAIL.n19 0.155672
R2269 VTAIL.n63 VTAIL.n19 0.155672
R2270 VTAIL.n64 VTAIL.n63 0.155672
R2271 VTAIL.n64 VTAIL.n15 0.155672
R2272 VTAIL.n71 VTAIL.n15 0.155672
R2273 VTAIL.n72 VTAIL.n71 0.155672
R2274 VTAIL.n72 VTAIL.n11 0.155672
R2275 VTAIL.n81 VTAIL.n11 0.155672
R2276 VTAIL.n82 VTAIL.n81 0.155672
R2277 VTAIL.n82 VTAIL.n7 0.155672
R2278 VTAIL.n89 VTAIL.n7 0.155672
R2279 VTAIL.n90 VTAIL.n89 0.155672
R2280 VTAIL.n90 VTAIL.n3 0.155672
R2281 VTAIL.n97 VTAIL.n3 0.155672
R2282 VTAIL.n299 VTAIL.n205 0.155672
R2283 VTAIL.n292 VTAIL.n205 0.155672
R2284 VTAIL.n292 VTAIL.n291 0.155672
R2285 VTAIL.n291 VTAIL.n209 0.155672
R2286 VTAIL.n284 VTAIL.n209 0.155672
R2287 VTAIL.n284 VTAIL.n283 0.155672
R2288 VTAIL.n283 VTAIL.n213 0.155672
R2289 VTAIL.n276 VTAIL.n213 0.155672
R2290 VTAIL.n276 VTAIL.n275 0.155672
R2291 VTAIL.n275 VTAIL.n219 0.155672
R2292 VTAIL.n268 VTAIL.n219 0.155672
R2293 VTAIL.n268 VTAIL.n267 0.155672
R2294 VTAIL.n267 VTAIL.n223 0.155672
R2295 VTAIL.n260 VTAIL.n223 0.155672
R2296 VTAIL.n260 VTAIL.n259 0.155672
R2297 VTAIL.n259 VTAIL.n227 0.155672
R2298 VTAIL.n252 VTAIL.n227 0.155672
R2299 VTAIL.n252 VTAIL.n251 0.155672
R2300 VTAIL.n251 VTAIL.n231 0.155672
R2301 VTAIL.n244 VTAIL.n231 0.155672
R2302 VTAIL.n244 VTAIL.n243 0.155672
R2303 VTAIL.n243 VTAIL.n235 0.155672
R2304 VTAIL.n199 VTAIL.n105 0.155672
R2305 VTAIL.n192 VTAIL.n105 0.155672
R2306 VTAIL.n192 VTAIL.n191 0.155672
R2307 VTAIL.n191 VTAIL.n109 0.155672
R2308 VTAIL.n184 VTAIL.n109 0.155672
R2309 VTAIL.n184 VTAIL.n183 0.155672
R2310 VTAIL.n183 VTAIL.n113 0.155672
R2311 VTAIL.n176 VTAIL.n113 0.155672
R2312 VTAIL.n176 VTAIL.n175 0.155672
R2313 VTAIL.n175 VTAIL.n119 0.155672
R2314 VTAIL.n168 VTAIL.n119 0.155672
R2315 VTAIL.n168 VTAIL.n167 0.155672
R2316 VTAIL.n167 VTAIL.n123 0.155672
R2317 VTAIL.n160 VTAIL.n123 0.155672
R2318 VTAIL.n160 VTAIL.n159 0.155672
R2319 VTAIL.n159 VTAIL.n127 0.155672
R2320 VTAIL.n152 VTAIL.n127 0.155672
R2321 VTAIL.n152 VTAIL.n151 0.155672
R2322 VTAIL.n151 VTAIL.n131 0.155672
R2323 VTAIL.n144 VTAIL.n131 0.155672
R2324 VTAIL.n144 VTAIL.n143 0.155672
R2325 VTAIL.n143 VTAIL.n135 0.155672
R2326 VP.n11 VP.t4 172.542
R2327 VP.n13 VP.n10 161.3
R2328 VP.n15 VP.n14 161.3
R2329 VP.n16 VP.n9 161.3
R2330 VP.n18 VP.n17 161.3
R2331 VP.n19 VP.n8 161.3
R2332 VP.n21 VP.n20 161.3
R2333 VP.n44 VP.n43 161.3
R2334 VP.n42 VP.n1 161.3
R2335 VP.n41 VP.n40 161.3
R2336 VP.n39 VP.n2 161.3
R2337 VP.n38 VP.n37 161.3
R2338 VP.n36 VP.n3 161.3
R2339 VP.n35 VP.n34 161.3
R2340 VP.n33 VP.n4 161.3
R2341 VP.n32 VP.n31 161.3
R2342 VP.n30 VP.n5 161.3
R2343 VP.n29 VP.n28 161.3
R2344 VP.n27 VP.n6 161.3
R2345 VP.n26 VP.n25 161.3
R2346 VP.n35 VP.t0 139.088
R2347 VP.n24 VP.t2 139.088
R2348 VP.n0 VP.t5 139.088
R2349 VP.n12 VP.t3 139.088
R2350 VP.n7 VP.t1 139.088
R2351 VP.n24 VP.n23 71.0639
R2352 VP.n45 VP.n0 71.0639
R2353 VP.n22 VP.n7 71.0639
R2354 VP.n30 VP.n29 56.5617
R2355 VP.n41 VP.n2 56.5617
R2356 VP.n18 VP.n9 56.5617
R2357 VP.n23 VP.n22 54.8897
R2358 VP.n12 VP.n11 49.4645
R2359 VP.n25 VP.n6 24.5923
R2360 VP.n29 VP.n6 24.5923
R2361 VP.n31 VP.n30 24.5923
R2362 VP.n31 VP.n4 24.5923
R2363 VP.n35 VP.n4 24.5923
R2364 VP.n36 VP.n35 24.5923
R2365 VP.n37 VP.n36 24.5923
R2366 VP.n37 VP.n2 24.5923
R2367 VP.n42 VP.n41 24.5923
R2368 VP.n43 VP.n42 24.5923
R2369 VP.n19 VP.n18 24.5923
R2370 VP.n20 VP.n19 24.5923
R2371 VP.n13 VP.n12 24.5923
R2372 VP.n14 VP.n13 24.5923
R2373 VP.n14 VP.n9 24.5923
R2374 VP.n25 VP.n24 19.1821
R2375 VP.n43 VP.n0 19.1821
R2376 VP.n20 VP.n7 19.1821
R2377 VP.n11 VP.n10 3.94395
R2378 VP.n22 VP.n21 0.354861
R2379 VP.n26 VP.n23 0.354861
R2380 VP.n45 VP.n44 0.354861
R2381 VP VP.n45 0.267071
R2382 VP.n15 VP.n10 0.189894
R2383 VP.n16 VP.n15 0.189894
R2384 VP.n17 VP.n16 0.189894
R2385 VP.n17 VP.n8 0.189894
R2386 VP.n21 VP.n8 0.189894
R2387 VP.n27 VP.n26 0.189894
R2388 VP.n28 VP.n27 0.189894
R2389 VP.n28 VP.n5 0.189894
R2390 VP.n32 VP.n5 0.189894
R2391 VP.n33 VP.n32 0.189894
R2392 VP.n34 VP.n33 0.189894
R2393 VP.n34 VP.n3 0.189894
R2394 VP.n38 VP.n3 0.189894
R2395 VP.n39 VP.n38 0.189894
R2396 VP.n40 VP.n39 0.189894
R2397 VP.n40 VP.n1 0.189894
R2398 VP.n44 VP.n1 0.189894
R2399 VDD1.n92 VDD1.n0 756.745
R2400 VDD1.n189 VDD1.n97 756.745
R2401 VDD1.n93 VDD1.n92 585
R2402 VDD1.n91 VDD1.n90 585
R2403 VDD1.n4 VDD1.n3 585
R2404 VDD1.n85 VDD1.n84 585
R2405 VDD1.n83 VDD1.n82 585
R2406 VDD1.n8 VDD1.n7 585
R2407 VDD1.n12 VDD1.n10 585
R2408 VDD1.n77 VDD1.n76 585
R2409 VDD1.n75 VDD1.n74 585
R2410 VDD1.n14 VDD1.n13 585
R2411 VDD1.n69 VDD1.n68 585
R2412 VDD1.n67 VDD1.n66 585
R2413 VDD1.n18 VDD1.n17 585
R2414 VDD1.n61 VDD1.n60 585
R2415 VDD1.n59 VDD1.n58 585
R2416 VDD1.n22 VDD1.n21 585
R2417 VDD1.n53 VDD1.n52 585
R2418 VDD1.n51 VDD1.n50 585
R2419 VDD1.n26 VDD1.n25 585
R2420 VDD1.n45 VDD1.n44 585
R2421 VDD1.n43 VDD1.n42 585
R2422 VDD1.n30 VDD1.n29 585
R2423 VDD1.n37 VDD1.n36 585
R2424 VDD1.n35 VDD1.n34 585
R2425 VDD1.n130 VDD1.n129 585
R2426 VDD1.n132 VDD1.n131 585
R2427 VDD1.n125 VDD1.n124 585
R2428 VDD1.n138 VDD1.n137 585
R2429 VDD1.n140 VDD1.n139 585
R2430 VDD1.n121 VDD1.n120 585
R2431 VDD1.n146 VDD1.n145 585
R2432 VDD1.n148 VDD1.n147 585
R2433 VDD1.n117 VDD1.n116 585
R2434 VDD1.n154 VDD1.n153 585
R2435 VDD1.n156 VDD1.n155 585
R2436 VDD1.n113 VDD1.n112 585
R2437 VDD1.n162 VDD1.n161 585
R2438 VDD1.n164 VDD1.n163 585
R2439 VDD1.n109 VDD1.n108 585
R2440 VDD1.n171 VDD1.n170 585
R2441 VDD1.n172 VDD1.n107 585
R2442 VDD1.n174 VDD1.n173 585
R2443 VDD1.n105 VDD1.n104 585
R2444 VDD1.n180 VDD1.n179 585
R2445 VDD1.n182 VDD1.n181 585
R2446 VDD1.n101 VDD1.n100 585
R2447 VDD1.n188 VDD1.n187 585
R2448 VDD1.n190 VDD1.n189 585
R2449 VDD1.n33 VDD1.t1 327.466
R2450 VDD1.n128 VDD1.t3 327.466
R2451 VDD1.n92 VDD1.n91 171.744
R2452 VDD1.n91 VDD1.n3 171.744
R2453 VDD1.n84 VDD1.n3 171.744
R2454 VDD1.n84 VDD1.n83 171.744
R2455 VDD1.n83 VDD1.n7 171.744
R2456 VDD1.n12 VDD1.n7 171.744
R2457 VDD1.n76 VDD1.n12 171.744
R2458 VDD1.n76 VDD1.n75 171.744
R2459 VDD1.n75 VDD1.n13 171.744
R2460 VDD1.n68 VDD1.n13 171.744
R2461 VDD1.n68 VDD1.n67 171.744
R2462 VDD1.n67 VDD1.n17 171.744
R2463 VDD1.n60 VDD1.n17 171.744
R2464 VDD1.n60 VDD1.n59 171.744
R2465 VDD1.n59 VDD1.n21 171.744
R2466 VDD1.n52 VDD1.n21 171.744
R2467 VDD1.n52 VDD1.n51 171.744
R2468 VDD1.n51 VDD1.n25 171.744
R2469 VDD1.n44 VDD1.n25 171.744
R2470 VDD1.n44 VDD1.n43 171.744
R2471 VDD1.n43 VDD1.n29 171.744
R2472 VDD1.n36 VDD1.n29 171.744
R2473 VDD1.n36 VDD1.n35 171.744
R2474 VDD1.n131 VDD1.n130 171.744
R2475 VDD1.n131 VDD1.n124 171.744
R2476 VDD1.n138 VDD1.n124 171.744
R2477 VDD1.n139 VDD1.n138 171.744
R2478 VDD1.n139 VDD1.n120 171.744
R2479 VDD1.n146 VDD1.n120 171.744
R2480 VDD1.n147 VDD1.n146 171.744
R2481 VDD1.n147 VDD1.n116 171.744
R2482 VDD1.n154 VDD1.n116 171.744
R2483 VDD1.n155 VDD1.n154 171.744
R2484 VDD1.n155 VDD1.n112 171.744
R2485 VDD1.n162 VDD1.n112 171.744
R2486 VDD1.n163 VDD1.n162 171.744
R2487 VDD1.n163 VDD1.n108 171.744
R2488 VDD1.n171 VDD1.n108 171.744
R2489 VDD1.n172 VDD1.n171 171.744
R2490 VDD1.n173 VDD1.n172 171.744
R2491 VDD1.n173 VDD1.n104 171.744
R2492 VDD1.n180 VDD1.n104 171.744
R2493 VDD1.n181 VDD1.n180 171.744
R2494 VDD1.n181 VDD1.n100 171.744
R2495 VDD1.n188 VDD1.n100 171.744
R2496 VDD1.n189 VDD1.n188 171.744
R2497 VDD1.n35 VDD1.t1 85.8723
R2498 VDD1.n130 VDD1.t3 85.8723
R2499 VDD1.n195 VDD1.n194 72.4125
R2500 VDD1.n197 VDD1.n196 71.7372
R2501 VDD1 VDD1.n96 53.8293
R2502 VDD1.n195 VDD1.n193 53.7158
R2503 VDD1.n197 VDD1.n195 50.4815
R2504 VDD1.n34 VDD1.n33 16.3895
R2505 VDD1.n129 VDD1.n128 16.3895
R2506 VDD1.n10 VDD1.n8 13.1884
R2507 VDD1.n174 VDD1.n105 13.1884
R2508 VDD1.n82 VDD1.n81 12.8005
R2509 VDD1.n78 VDD1.n77 12.8005
R2510 VDD1.n37 VDD1.n32 12.8005
R2511 VDD1.n132 VDD1.n127 12.8005
R2512 VDD1.n175 VDD1.n107 12.8005
R2513 VDD1.n179 VDD1.n178 12.8005
R2514 VDD1.n85 VDD1.n6 12.0247
R2515 VDD1.n74 VDD1.n11 12.0247
R2516 VDD1.n38 VDD1.n30 12.0247
R2517 VDD1.n133 VDD1.n125 12.0247
R2518 VDD1.n170 VDD1.n169 12.0247
R2519 VDD1.n182 VDD1.n103 12.0247
R2520 VDD1.n86 VDD1.n4 11.249
R2521 VDD1.n73 VDD1.n14 11.249
R2522 VDD1.n42 VDD1.n41 11.249
R2523 VDD1.n137 VDD1.n136 11.249
R2524 VDD1.n168 VDD1.n109 11.249
R2525 VDD1.n183 VDD1.n101 11.249
R2526 VDD1.n90 VDD1.n89 10.4732
R2527 VDD1.n70 VDD1.n69 10.4732
R2528 VDD1.n45 VDD1.n28 10.4732
R2529 VDD1.n140 VDD1.n123 10.4732
R2530 VDD1.n165 VDD1.n164 10.4732
R2531 VDD1.n187 VDD1.n186 10.4732
R2532 VDD1.n93 VDD1.n2 9.69747
R2533 VDD1.n66 VDD1.n16 9.69747
R2534 VDD1.n46 VDD1.n26 9.69747
R2535 VDD1.n141 VDD1.n121 9.69747
R2536 VDD1.n161 VDD1.n111 9.69747
R2537 VDD1.n190 VDD1.n99 9.69747
R2538 VDD1.n96 VDD1.n95 9.45567
R2539 VDD1.n193 VDD1.n192 9.45567
R2540 VDD1.n20 VDD1.n19 9.3005
R2541 VDD1.n63 VDD1.n62 9.3005
R2542 VDD1.n65 VDD1.n64 9.3005
R2543 VDD1.n16 VDD1.n15 9.3005
R2544 VDD1.n71 VDD1.n70 9.3005
R2545 VDD1.n73 VDD1.n72 9.3005
R2546 VDD1.n11 VDD1.n9 9.3005
R2547 VDD1.n79 VDD1.n78 9.3005
R2548 VDD1.n95 VDD1.n94 9.3005
R2549 VDD1.n2 VDD1.n1 9.3005
R2550 VDD1.n89 VDD1.n88 9.3005
R2551 VDD1.n87 VDD1.n86 9.3005
R2552 VDD1.n6 VDD1.n5 9.3005
R2553 VDD1.n81 VDD1.n80 9.3005
R2554 VDD1.n57 VDD1.n56 9.3005
R2555 VDD1.n55 VDD1.n54 9.3005
R2556 VDD1.n24 VDD1.n23 9.3005
R2557 VDD1.n49 VDD1.n48 9.3005
R2558 VDD1.n47 VDD1.n46 9.3005
R2559 VDD1.n28 VDD1.n27 9.3005
R2560 VDD1.n41 VDD1.n40 9.3005
R2561 VDD1.n39 VDD1.n38 9.3005
R2562 VDD1.n32 VDD1.n31 9.3005
R2563 VDD1.n192 VDD1.n191 9.3005
R2564 VDD1.n99 VDD1.n98 9.3005
R2565 VDD1.n186 VDD1.n185 9.3005
R2566 VDD1.n184 VDD1.n183 9.3005
R2567 VDD1.n103 VDD1.n102 9.3005
R2568 VDD1.n178 VDD1.n177 9.3005
R2569 VDD1.n150 VDD1.n149 9.3005
R2570 VDD1.n119 VDD1.n118 9.3005
R2571 VDD1.n144 VDD1.n143 9.3005
R2572 VDD1.n142 VDD1.n141 9.3005
R2573 VDD1.n123 VDD1.n122 9.3005
R2574 VDD1.n136 VDD1.n135 9.3005
R2575 VDD1.n134 VDD1.n133 9.3005
R2576 VDD1.n127 VDD1.n126 9.3005
R2577 VDD1.n152 VDD1.n151 9.3005
R2578 VDD1.n115 VDD1.n114 9.3005
R2579 VDD1.n158 VDD1.n157 9.3005
R2580 VDD1.n160 VDD1.n159 9.3005
R2581 VDD1.n111 VDD1.n110 9.3005
R2582 VDD1.n166 VDD1.n165 9.3005
R2583 VDD1.n168 VDD1.n167 9.3005
R2584 VDD1.n169 VDD1.n106 9.3005
R2585 VDD1.n176 VDD1.n175 9.3005
R2586 VDD1.n94 VDD1.n0 8.92171
R2587 VDD1.n65 VDD1.n18 8.92171
R2588 VDD1.n50 VDD1.n49 8.92171
R2589 VDD1.n145 VDD1.n144 8.92171
R2590 VDD1.n160 VDD1.n113 8.92171
R2591 VDD1.n191 VDD1.n97 8.92171
R2592 VDD1.n62 VDD1.n61 8.14595
R2593 VDD1.n53 VDD1.n24 8.14595
R2594 VDD1.n148 VDD1.n119 8.14595
R2595 VDD1.n157 VDD1.n156 8.14595
R2596 VDD1.n58 VDD1.n20 7.3702
R2597 VDD1.n54 VDD1.n22 7.3702
R2598 VDD1.n149 VDD1.n117 7.3702
R2599 VDD1.n153 VDD1.n115 7.3702
R2600 VDD1.n58 VDD1.n57 6.59444
R2601 VDD1.n57 VDD1.n22 6.59444
R2602 VDD1.n152 VDD1.n117 6.59444
R2603 VDD1.n153 VDD1.n152 6.59444
R2604 VDD1.n61 VDD1.n20 5.81868
R2605 VDD1.n54 VDD1.n53 5.81868
R2606 VDD1.n149 VDD1.n148 5.81868
R2607 VDD1.n156 VDD1.n115 5.81868
R2608 VDD1.n96 VDD1.n0 5.04292
R2609 VDD1.n62 VDD1.n18 5.04292
R2610 VDD1.n50 VDD1.n24 5.04292
R2611 VDD1.n145 VDD1.n119 5.04292
R2612 VDD1.n157 VDD1.n113 5.04292
R2613 VDD1.n193 VDD1.n97 5.04292
R2614 VDD1.n94 VDD1.n93 4.26717
R2615 VDD1.n66 VDD1.n65 4.26717
R2616 VDD1.n49 VDD1.n26 4.26717
R2617 VDD1.n144 VDD1.n121 4.26717
R2618 VDD1.n161 VDD1.n160 4.26717
R2619 VDD1.n191 VDD1.n190 4.26717
R2620 VDD1.n33 VDD1.n31 3.70982
R2621 VDD1.n128 VDD1.n126 3.70982
R2622 VDD1.n90 VDD1.n2 3.49141
R2623 VDD1.n69 VDD1.n16 3.49141
R2624 VDD1.n46 VDD1.n45 3.49141
R2625 VDD1.n141 VDD1.n140 3.49141
R2626 VDD1.n164 VDD1.n111 3.49141
R2627 VDD1.n187 VDD1.n99 3.49141
R2628 VDD1.n89 VDD1.n4 2.71565
R2629 VDD1.n70 VDD1.n14 2.71565
R2630 VDD1.n42 VDD1.n28 2.71565
R2631 VDD1.n137 VDD1.n123 2.71565
R2632 VDD1.n165 VDD1.n109 2.71565
R2633 VDD1.n186 VDD1.n101 2.71565
R2634 VDD1.n86 VDD1.n85 1.93989
R2635 VDD1.n74 VDD1.n73 1.93989
R2636 VDD1.n41 VDD1.n30 1.93989
R2637 VDD1.n136 VDD1.n125 1.93989
R2638 VDD1.n170 VDD1.n168 1.93989
R2639 VDD1.n183 VDD1.n182 1.93989
R2640 VDD1.n196 VDD1.t2 1.8411
R2641 VDD1.n196 VDD1.t4 1.8411
R2642 VDD1.n194 VDD1.t5 1.8411
R2643 VDD1.n194 VDD1.t0 1.8411
R2644 VDD1.n82 VDD1.n6 1.16414
R2645 VDD1.n77 VDD1.n11 1.16414
R2646 VDD1.n38 VDD1.n37 1.16414
R2647 VDD1.n133 VDD1.n132 1.16414
R2648 VDD1.n169 VDD1.n107 1.16414
R2649 VDD1.n179 VDD1.n103 1.16414
R2650 VDD1 VDD1.n197 0.672914
R2651 VDD1.n81 VDD1.n8 0.388379
R2652 VDD1.n78 VDD1.n10 0.388379
R2653 VDD1.n34 VDD1.n32 0.388379
R2654 VDD1.n129 VDD1.n127 0.388379
R2655 VDD1.n175 VDD1.n174 0.388379
R2656 VDD1.n178 VDD1.n105 0.388379
R2657 VDD1.n95 VDD1.n1 0.155672
R2658 VDD1.n88 VDD1.n1 0.155672
R2659 VDD1.n88 VDD1.n87 0.155672
R2660 VDD1.n87 VDD1.n5 0.155672
R2661 VDD1.n80 VDD1.n5 0.155672
R2662 VDD1.n80 VDD1.n79 0.155672
R2663 VDD1.n79 VDD1.n9 0.155672
R2664 VDD1.n72 VDD1.n9 0.155672
R2665 VDD1.n72 VDD1.n71 0.155672
R2666 VDD1.n71 VDD1.n15 0.155672
R2667 VDD1.n64 VDD1.n15 0.155672
R2668 VDD1.n64 VDD1.n63 0.155672
R2669 VDD1.n63 VDD1.n19 0.155672
R2670 VDD1.n56 VDD1.n19 0.155672
R2671 VDD1.n56 VDD1.n55 0.155672
R2672 VDD1.n55 VDD1.n23 0.155672
R2673 VDD1.n48 VDD1.n23 0.155672
R2674 VDD1.n48 VDD1.n47 0.155672
R2675 VDD1.n47 VDD1.n27 0.155672
R2676 VDD1.n40 VDD1.n27 0.155672
R2677 VDD1.n40 VDD1.n39 0.155672
R2678 VDD1.n39 VDD1.n31 0.155672
R2679 VDD1.n134 VDD1.n126 0.155672
R2680 VDD1.n135 VDD1.n134 0.155672
R2681 VDD1.n135 VDD1.n122 0.155672
R2682 VDD1.n142 VDD1.n122 0.155672
R2683 VDD1.n143 VDD1.n142 0.155672
R2684 VDD1.n143 VDD1.n118 0.155672
R2685 VDD1.n150 VDD1.n118 0.155672
R2686 VDD1.n151 VDD1.n150 0.155672
R2687 VDD1.n151 VDD1.n114 0.155672
R2688 VDD1.n158 VDD1.n114 0.155672
R2689 VDD1.n159 VDD1.n158 0.155672
R2690 VDD1.n159 VDD1.n110 0.155672
R2691 VDD1.n166 VDD1.n110 0.155672
R2692 VDD1.n167 VDD1.n166 0.155672
R2693 VDD1.n167 VDD1.n106 0.155672
R2694 VDD1.n176 VDD1.n106 0.155672
R2695 VDD1.n177 VDD1.n176 0.155672
R2696 VDD1.n177 VDD1.n102 0.155672
R2697 VDD1.n184 VDD1.n102 0.155672
R2698 VDD1.n185 VDD1.n184 0.155672
R2699 VDD1.n185 VDD1.n98 0.155672
R2700 VDD1.n192 VDD1.n98 0.155672
C0 VDD2 VN 9.99884f
C1 VDD1 B 2.66521f
C2 VDD1 VP 10.3412f
C3 VDD2 B 2.75033f
C4 VTAIL w_n3682_n4500# 3.7933f
C5 VDD2 VP 0.498138f
C6 VN w_n3682_n4500# 7.18485f
C7 VDD1 VDD2 1.58755f
C8 w_n3682_n4500# B 11.8986f
C9 w_n3682_n4500# VP 7.66217f
C10 VN VTAIL 10.0109f
C11 VDD1 w_n3682_n4500# 2.79433f
C12 VTAIL B 5.17917f
C13 VDD2 w_n3682_n4500# 2.89409f
C14 VTAIL VP 10.0252f
C15 VN B 1.33481f
C16 VDD1 VTAIL 9.78217f
C17 VN VP 8.418281f
C18 VDD2 VTAIL 9.83541f
C19 VDD1 VN 0.151789f
C20 B VP 2.13405f
C21 VDD2 VSUBS 2.17259f
C22 VDD1 VSUBS 2.142432f
C23 VTAIL VSUBS 1.490361f
C24 VN VSUBS 6.50248f
C25 VP VSUBS 3.509484f
C26 B VSUBS 5.570963f
C27 w_n3682_n4500# VSUBS 0.202672p
C28 VDD1.n0 VSUBS 0.03091f
C29 VDD1.n1 VSUBS 0.027186f
C30 VDD1.n2 VSUBS 0.014608f
C31 VDD1.n3 VSUBS 0.034529f
C32 VDD1.n4 VSUBS 0.015468f
C33 VDD1.n5 VSUBS 0.027186f
C34 VDD1.n6 VSUBS 0.014608f
C35 VDD1.n7 VSUBS 0.034529f
C36 VDD1.n8 VSUBS 0.015038f
C37 VDD1.n9 VSUBS 0.027186f
C38 VDD1.n10 VSUBS 0.015038f
C39 VDD1.n11 VSUBS 0.014608f
C40 VDD1.n12 VSUBS 0.034529f
C41 VDD1.n13 VSUBS 0.034529f
C42 VDD1.n14 VSUBS 0.015468f
C43 VDD1.n15 VSUBS 0.027186f
C44 VDD1.n16 VSUBS 0.014608f
C45 VDD1.n17 VSUBS 0.034529f
C46 VDD1.n18 VSUBS 0.015468f
C47 VDD1.n19 VSUBS 0.027186f
C48 VDD1.n20 VSUBS 0.014608f
C49 VDD1.n21 VSUBS 0.034529f
C50 VDD1.n22 VSUBS 0.015468f
C51 VDD1.n23 VSUBS 0.027186f
C52 VDD1.n24 VSUBS 0.014608f
C53 VDD1.n25 VSUBS 0.034529f
C54 VDD1.n26 VSUBS 0.015468f
C55 VDD1.n27 VSUBS 0.027186f
C56 VDD1.n28 VSUBS 0.014608f
C57 VDD1.n29 VSUBS 0.034529f
C58 VDD1.n30 VSUBS 0.015468f
C59 VDD1.n31 VSUBS 2.06416f
C60 VDD1.n32 VSUBS 0.014608f
C61 VDD1.t1 VSUBS 0.0741f
C62 VDD1.n33 VSUBS 0.212966f
C63 VDD1.n34 VSUBS 0.021966f
C64 VDD1.n35 VSUBS 0.025897f
C65 VDD1.n36 VSUBS 0.034529f
C66 VDD1.n37 VSUBS 0.015468f
C67 VDD1.n38 VSUBS 0.014608f
C68 VDD1.n39 VSUBS 0.027186f
C69 VDD1.n40 VSUBS 0.027186f
C70 VDD1.n41 VSUBS 0.014608f
C71 VDD1.n42 VSUBS 0.015468f
C72 VDD1.n43 VSUBS 0.034529f
C73 VDD1.n44 VSUBS 0.034529f
C74 VDD1.n45 VSUBS 0.015468f
C75 VDD1.n46 VSUBS 0.014608f
C76 VDD1.n47 VSUBS 0.027186f
C77 VDD1.n48 VSUBS 0.027186f
C78 VDD1.n49 VSUBS 0.014608f
C79 VDD1.n50 VSUBS 0.015468f
C80 VDD1.n51 VSUBS 0.034529f
C81 VDD1.n52 VSUBS 0.034529f
C82 VDD1.n53 VSUBS 0.015468f
C83 VDD1.n54 VSUBS 0.014608f
C84 VDD1.n55 VSUBS 0.027186f
C85 VDD1.n56 VSUBS 0.027186f
C86 VDD1.n57 VSUBS 0.014608f
C87 VDD1.n58 VSUBS 0.015468f
C88 VDD1.n59 VSUBS 0.034529f
C89 VDD1.n60 VSUBS 0.034529f
C90 VDD1.n61 VSUBS 0.015468f
C91 VDD1.n62 VSUBS 0.014608f
C92 VDD1.n63 VSUBS 0.027186f
C93 VDD1.n64 VSUBS 0.027186f
C94 VDD1.n65 VSUBS 0.014608f
C95 VDD1.n66 VSUBS 0.015468f
C96 VDD1.n67 VSUBS 0.034529f
C97 VDD1.n68 VSUBS 0.034529f
C98 VDD1.n69 VSUBS 0.015468f
C99 VDD1.n70 VSUBS 0.014608f
C100 VDD1.n71 VSUBS 0.027186f
C101 VDD1.n72 VSUBS 0.027186f
C102 VDD1.n73 VSUBS 0.014608f
C103 VDD1.n74 VSUBS 0.015468f
C104 VDD1.n75 VSUBS 0.034529f
C105 VDD1.n76 VSUBS 0.034529f
C106 VDD1.n77 VSUBS 0.015468f
C107 VDD1.n78 VSUBS 0.014608f
C108 VDD1.n79 VSUBS 0.027186f
C109 VDD1.n80 VSUBS 0.027186f
C110 VDD1.n81 VSUBS 0.014608f
C111 VDD1.n82 VSUBS 0.015468f
C112 VDD1.n83 VSUBS 0.034529f
C113 VDD1.n84 VSUBS 0.034529f
C114 VDD1.n85 VSUBS 0.015468f
C115 VDD1.n86 VSUBS 0.014608f
C116 VDD1.n87 VSUBS 0.027186f
C117 VDD1.n88 VSUBS 0.027186f
C118 VDD1.n89 VSUBS 0.014608f
C119 VDD1.n90 VSUBS 0.015468f
C120 VDD1.n91 VSUBS 0.034529f
C121 VDD1.n92 VSUBS 0.08713f
C122 VDD1.n93 VSUBS 0.015468f
C123 VDD1.n94 VSUBS 0.014608f
C124 VDD1.n95 VSUBS 0.068038f
C125 VDD1.n96 VSUBS 0.073413f
C126 VDD1.n97 VSUBS 0.03091f
C127 VDD1.n98 VSUBS 0.027186f
C128 VDD1.n99 VSUBS 0.014608f
C129 VDD1.n100 VSUBS 0.034529f
C130 VDD1.n101 VSUBS 0.015468f
C131 VDD1.n102 VSUBS 0.027186f
C132 VDD1.n103 VSUBS 0.014608f
C133 VDD1.n104 VSUBS 0.034529f
C134 VDD1.n105 VSUBS 0.015038f
C135 VDD1.n106 VSUBS 0.027186f
C136 VDD1.n107 VSUBS 0.015468f
C137 VDD1.n108 VSUBS 0.034529f
C138 VDD1.n109 VSUBS 0.015468f
C139 VDD1.n110 VSUBS 0.027186f
C140 VDD1.n111 VSUBS 0.014608f
C141 VDD1.n112 VSUBS 0.034529f
C142 VDD1.n113 VSUBS 0.015468f
C143 VDD1.n114 VSUBS 0.027186f
C144 VDD1.n115 VSUBS 0.014608f
C145 VDD1.n116 VSUBS 0.034529f
C146 VDD1.n117 VSUBS 0.015468f
C147 VDD1.n118 VSUBS 0.027186f
C148 VDD1.n119 VSUBS 0.014608f
C149 VDD1.n120 VSUBS 0.034529f
C150 VDD1.n121 VSUBS 0.015468f
C151 VDD1.n122 VSUBS 0.027186f
C152 VDD1.n123 VSUBS 0.014608f
C153 VDD1.n124 VSUBS 0.034529f
C154 VDD1.n125 VSUBS 0.015468f
C155 VDD1.n126 VSUBS 2.06416f
C156 VDD1.n127 VSUBS 0.014608f
C157 VDD1.t3 VSUBS 0.0741f
C158 VDD1.n128 VSUBS 0.212966f
C159 VDD1.n129 VSUBS 0.021966f
C160 VDD1.n130 VSUBS 0.025897f
C161 VDD1.n131 VSUBS 0.034529f
C162 VDD1.n132 VSUBS 0.015468f
C163 VDD1.n133 VSUBS 0.014608f
C164 VDD1.n134 VSUBS 0.027186f
C165 VDD1.n135 VSUBS 0.027186f
C166 VDD1.n136 VSUBS 0.014608f
C167 VDD1.n137 VSUBS 0.015468f
C168 VDD1.n138 VSUBS 0.034529f
C169 VDD1.n139 VSUBS 0.034529f
C170 VDD1.n140 VSUBS 0.015468f
C171 VDD1.n141 VSUBS 0.014608f
C172 VDD1.n142 VSUBS 0.027186f
C173 VDD1.n143 VSUBS 0.027186f
C174 VDD1.n144 VSUBS 0.014608f
C175 VDD1.n145 VSUBS 0.015468f
C176 VDD1.n146 VSUBS 0.034529f
C177 VDD1.n147 VSUBS 0.034529f
C178 VDD1.n148 VSUBS 0.015468f
C179 VDD1.n149 VSUBS 0.014608f
C180 VDD1.n150 VSUBS 0.027186f
C181 VDD1.n151 VSUBS 0.027186f
C182 VDD1.n152 VSUBS 0.014608f
C183 VDD1.n153 VSUBS 0.015468f
C184 VDD1.n154 VSUBS 0.034529f
C185 VDD1.n155 VSUBS 0.034529f
C186 VDD1.n156 VSUBS 0.015468f
C187 VDD1.n157 VSUBS 0.014608f
C188 VDD1.n158 VSUBS 0.027186f
C189 VDD1.n159 VSUBS 0.027186f
C190 VDD1.n160 VSUBS 0.014608f
C191 VDD1.n161 VSUBS 0.015468f
C192 VDD1.n162 VSUBS 0.034529f
C193 VDD1.n163 VSUBS 0.034529f
C194 VDD1.n164 VSUBS 0.015468f
C195 VDD1.n165 VSUBS 0.014608f
C196 VDD1.n166 VSUBS 0.027186f
C197 VDD1.n167 VSUBS 0.027186f
C198 VDD1.n168 VSUBS 0.014608f
C199 VDD1.n169 VSUBS 0.014608f
C200 VDD1.n170 VSUBS 0.015468f
C201 VDD1.n171 VSUBS 0.034529f
C202 VDD1.n172 VSUBS 0.034529f
C203 VDD1.n173 VSUBS 0.034529f
C204 VDD1.n174 VSUBS 0.015038f
C205 VDD1.n175 VSUBS 0.014608f
C206 VDD1.n176 VSUBS 0.027186f
C207 VDD1.n177 VSUBS 0.027186f
C208 VDD1.n178 VSUBS 0.014608f
C209 VDD1.n179 VSUBS 0.015468f
C210 VDD1.n180 VSUBS 0.034529f
C211 VDD1.n181 VSUBS 0.034529f
C212 VDD1.n182 VSUBS 0.015468f
C213 VDD1.n183 VSUBS 0.014608f
C214 VDD1.n184 VSUBS 0.027186f
C215 VDD1.n185 VSUBS 0.027186f
C216 VDD1.n186 VSUBS 0.014608f
C217 VDD1.n187 VSUBS 0.015468f
C218 VDD1.n188 VSUBS 0.034529f
C219 VDD1.n189 VSUBS 0.08713f
C220 VDD1.n190 VSUBS 0.015468f
C221 VDD1.n191 VSUBS 0.014608f
C222 VDD1.n192 VSUBS 0.068038f
C223 VDD1.n193 VSUBS 0.072518f
C224 VDD1.t5 VSUBS 0.379391f
C225 VDD1.t0 VSUBS 0.379391f
C226 VDD1.n194 VSUBS 3.16431f
C227 VDD1.n195 VSUBS 3.96631f
C228 VDD1.t2 VSUBS 0.379391f
C229 VDD1.t4 VSUBS 0.379391f
C230 VDD1.n196 VSUBS 3.15638f
C231 VDD1.n197 VSUBS 3.93842f
C232 VP.t5 VSUBS 4.01571f
C233 VP.n0 VSUBS 1.49534f
C234 VP.n1 VSUBS 0.027026f
C235 VP.n2 VSUBS 0.035174f
C236 VP.n3 VSUBS 0.027026f
C237 VP.t0 VSUBS 4.01571f
C238 VP.n4 VSUBS 0.050118f
C239 VP.n5 VSUBS 0.027026f
C240 VP.n6 VSUBS 0.050118f
C241 VP.t1 VSUBS 4.01571f
C242 VP.n7 VSUBS 1.49534f
C243 VP.n8 VSUBS 0.027026f
C244 VP.n9 VSUBS 0.035174f
C245 VP.n10 VSUBS 0.307391f
C246 VP.t3 VSUBS 4.01571f
C247 VP.t4 VSUBS 4.32158f
C248 VP.n11 VSUBS 1.42522f
C249 VP.n12 VSUBS 1.48947f
C250 VP.n13 VSUBS 0.050118f
C251 VP.n14 VSUBS 0.050118f
C252 VP.n15 VSUBS 0.027026f
C253 VP.n16 VSUBS 0.027026f
C254 VP.n17 VSUBS 0.027026f
C255 VP.n18 VSUBS 0.043399f
C256 VP.n19 VSUBS 0.050118f
C257 VP.n20 VSUBS 0.044675f
C258 VP.n21 VSUBS 0.043613f
C259 VP.n22 VSUBS 1.74538f
C260 VP.n23 VSUBS 1.76314f
C261 VP.t2 VSUBS 4.01571f
C262 VP.n24 VSUBS 1.49534f
C263 VP.n25 VSUBS 0.044675f
C264 VP.n26 VSUBS 0.043613f
C265 VP.n27 VSUBS 0.027026f
C266 VP.n28 VSUBS 0.027026f
C267 VP.n29 VSUBS 0.043399f
C268 VP.n30 VSUBS 0.035174f
C269 VP.n31 VSUBS 0.050118f
C270 VP.n32 VSUBS 0.027026f
C271 VP.n33 VSUBS 0.027026f
C272 VP.n34 VSUBS 0.027026f
C273 VP.n35 VSUBS 1.41444f
C274 VP.n36 VSUBS 0.050118f
C275 VP.n37 VSUBS 0.050118f
C276 VP.n38 VSUBS 0.027026f
C277 VP.n39 VSUBS 0.027026f
C278 VP.n40 VSUBS 0.027026f
C279 VP.n41 VSUBS 0.043399f
C280 VP.n42 VSUBS 0.050118f
C281 VP.n43 VSUBS 0.044675f
C282 VP.n44 VSUBS 0.043613f
C283 VP.n45 VSUBS 0.057859f
C284 VTAIL.t7 VSUBS 0.38913f
C285 VTAIL.t11 VSUBS 0.38913f
C286 VTAIL.n0 VSUBS 3.07659f
C287 VTAIL.n1 VSUBS 0.903464f
C288 VTAIL.n2 VSUBS 0.031704f
C289 VTAIL.n3 VSUBS 0.027884f
C290 VTAIL.n4 VSUBS 0.014984f
C291 VTAIL.n5 VSUBS 0.035416f
C292 VTAIL.n6 VSUBS 0.015865f
C293 VTAIL.n7 VSUBS 0.027884f
C294 VTAIL.n8 VSUBS 0.014984f
C295 VTAIL.n9 VSUBS 0.035416f
C296 VTAIL.n10 VSUBS 0.015424f
C297 VTAIL.n11 VSUBS 0.027884f
C298 VTAIL.n12 VSUBS 0.015865f
C299 VTAIL.n13 VSUBS 0.035416f
C300 VTAIL.n14 VSUBS 0.015865f
C301 VTAIL.n15 VSUBS 0.027884f
C302 VTAIL.n16 VSUBS 0.014984f
C303 VTAIL.n17 VSUBS 0.035416f
C304 VTAIL.n18 VSUBS 0.015865f
C305 VTAIL.n19 VSUBS 0.027884f
C306 VTAIL.n20 VSUBS 0.014984f
C307 VTAIL.n21 VSUBS 0.035416f
C308 VTAIL.n22 VSUBS 0.015865f
C309 VTAIL.n23 VSUBS 0.027884f
C310 VTAIL.n24 VSUBS 0.014984f
C311 VTAIL.n25 VSUBS 0.035416f
C312 VTAIL.n26 VSUBS 0.015865f
C313 VTAIL.n27 VSUBS 0.027884f
C314 VTAIL.n28 VSUBS 0.014984f
C315 VTAIL.n29 VSUBS 0.035416f
C316 VTAIL.n30 VSUBS 0.015865f
C317 VTAIL.n31 VSUBS 2.11714f
C318 VTAIL.n32 VSUBS 0.014984f
C319 VTAIL.t2 VSUBS 0.076002f
C320 VTAIL.n33 VSUBS 0.218433f
C321 VTAIL.n34 VSUBS 0.02253f
C322 VTAIL.n35 VSUBS 0.026562f
C323 VTAIL.n36 VSUBS 0.035416f
C324 VTAIL.n37 VSUBS 0.015865f
C325 VTAIL.n38 VSUBS 0.014984f
C326 VTAIL.n39 VSUBS 0.027884f
C327 VTAIL.n40 VSUBS 0.027884f
C328 VTAIL.n41 VSUBS 0.014984f
C329 VTAIL.n42 VSUBS 0.015865f
C330 VTAIL.n43 VSUBS 0.035416f
C331 VTAIL.n44 VSUBS 0.035416f
C332 VTAIL.n45 VSUBS 0.015865f
C333 VTAIL.n46 VSUBS 0.014984f
C334 VTAIL.n47 VSUBS 0.027884f
C335 VTAIL.n48 VSUBS 0.027884f
C336 VTAIL.n49 VSUBS 0.014984f
C337 VTAIL.n50 VSUBS 0.015865f
C338 VTAIL.n51 VSUBS 0.035416f
C339 VTAIL.n52 VSUBS 0.035416f
C340 VTAIL.n53 VSUBS 0.015865f
C341 VTAIL.n54 VSUBS 0.014984f
C342 VTAIL.n55 VSUBS 0.027884f
C343 VTAIL.n56 VSUBS 0.027884f
C344 VTAIL.n57 VSUBS 0.014984f
C345 VTAIL.n58 VSUBS 0.015865f
C346 VTAIL.n59 VSUBS 0.035416f
C347 VTAIL.n60 VSUBS 0.035416f
C348 VTAIL.n61 VSUBS 0.015865f
C349 VTAIL.n62 VSUBS 0.014984f
C350 VTAIL.n63 VSUBS 0.027884f
C351 VTAIL.n64 VSUBS 0.027884f
C352 VTAIL.n65 VSUBS 0.014984f
C353 VTAIL.n66 VSUBS 0.015865f
C354 VTAIL.n67 VSUBS 0.035416f
C355 VTAIL.n68 VSUBS 0.035416f
C356 VTAIL.n69 VSUBS 0.015865f
C357 VTAIL.n70 VSUBS 0.014984f
C358 VTAIL.n71 VSUBS 0.027884f
C359 VTAIL.n72 VSUBS 0.027884f
C360 VTAIL.n73 VSUBS 0.014984f
C361 VTAIL.n74 VSUBS 0.014984f
C362 VTAIL.n75 VSUBS 0.015865f
C363 VTAIL.n76 VSUBS 0.035416f
C364 VTAIL.n77 VSUBS 0.035416f
C365 VTAIL.n78 VSUBS 0.035416f
C366 VTAIL.n79 VSUBS 0.015424f
C367 VTAIL.n80 VSUBS 0.014984f
C368 VTAIL.n81 VSUBS 0.027884f
C369 VTAIL.n82 VSUBS 0.027884f
C370 VTAIL.n83 VSUBS 0.014984f
C371 VTAIL.n84 VSUBS 0.015865f
C372 VTAIL.n85 VSUBS 0.035416f
C373 VTAIL.n86 VSUBS 0.035416f
C374 VTAIL.n87 VSUBS 0.015865f
C375 VTAIL.n88 VSUBS 0.014984f
C376 VTAIL.n89 VSUBS 0.027884f
C377 VTAIL.n90 VSUBS 0.027884f
C378 VTAIL.n91 VSUBS 0.014984f
C379 VTAIL.n92 VSUBS 0.015865f
C380 VTAIL.n93 VSUBS 0.035416f
C381 VTAIL.n94 VSUBS 0.089366f
C382 VTAIL.n95 VSUBS 0.015865f
C383 VTAIL.n96 VSUBS 0.014984f
C384 VTAIL.n97 VSUBS 0.069785f
C385 VTAIL.n98 VSUBS 0.045261f
C386 VTAIL.n99 VSUBS 0.4629f
C387 VTAIL.t1 VSUBS 0.38913f
C388 VTAIL.t3 VSUBS 0.38913f
C389 VTAIL.n100 VSUBS 3.07659f
C390 VTAIL.n101 VSUBS 3.19343f
C391 VTAIL.t9 VSUBS 0.38913f
C392 VTAIL.t8 VSUBS 0.38913f
C393 VTAIL.n102 VSUBS 3.0766f
C394 VTAIL.n103 VSUBS 3.19341f
C395 VTAIL.n104 VSUBS 0.031704f
C396 VTAIL.n105 VSUBS 0.027884f
C397 VTAIL.n106 VSUBS 0.014984f
C398 VTAIL.n107 VSUBS 0.035416f
C399 VTAIL.n108 VSUBS 0.015865f
C400 VTAIL.n109 VSUBS 0.027884f
C401 VTAIL.n110 VSUBS 0.014984f
C402 VTAIL.n111 VSUBS 0.035416f
C403 VTAIL.n112 VSUBS 0.015424f
C404 VTAIL.n113 VSUBS 0.027884f
C405 VTAIL.n114 VSUBS 0.015424f
C406 VTAIL.n115 VSUBS 0.014984f
C407 VTAIL.n116 VSUBS 0.035416f
C408 VTAIL.n117 VSUBS 0.035416f
C409 VTAIL.n118 VSUBS 0.015865f
C410 VTAIL.n119 VSUBS 0.027884f
C411 VTAIL.n120 VSUBS 0.014984f
C412 VTAIL.n121 VSUBS 0.035416f
C413 VTAIL.n122 VSUBS 0.015865f
C414 VTAIL.n123 VSUBS 0.027884f
C415 VTAIL.n124 VSUBS 0.014984f
C416 VTAIL.n125 VSUBS 0.035416f
C417 VTAIL.n126 VSUBS 0.015865f
C418 VTAIL.n127 VSUBS 0.027884f
C419 VTAIL.n128 VSUBS 0.014984f
C420 VTAIL.n129 VSUBS 0.035416f
C421 VTAIL.n130 VSUBS 0.015865f
C422 VTAIL.n131 VSUBS 0.027884f
C423 VTAIL.n132 VSUBS 0.014984f
C424 VTAIL.n133 VSUBS 0.035416f
C425 VTAIL.n134 VSUBS 0.015865f
C426 VTAIL.n135 VSUBS 2.11714f
C427 VTAIL.n136 VSUBS 0.014984f
C428 VTAIL.t10 VSUBS 0.076002f
C429 VTAIL.n137 VSUBS 0.218433f
C430 VTAIL.n138 VSUBS 0.02253f
C431 VTAIL.n139 VSUBS 0.026562f
C432 VTAIL.n140 VSUBS 0.035416f
C433 VTAIL.n141 VSUBS 0.015865f
C434 VTAIL.n142 VSUBS 0.014984f
C435 VTAIL.n143 VSUBS 0.027884f
C436 VTAIL.n144 VSUBS 0.027884f
C437 VTAIL.n145 VSUBS 0.014984f
C438 VTAIL.n146 VSUBS 0.015865f
C439 VTAIL.n147 VSUBS 0.035416f
C440 VTAIL.n148 VSUBS 0.035416f
C441 VTAIL.n149 VSUBS 0.015865f
C442 VTAIL.n150 VSUBS 0.014984f
C443 VTAIL.n151 VSUBS 0.027884f
C444 VTAIL.n152 VSUBS 0.027884f
C445 VTAIL.n153 VSUBS 0.014984f
C446 VTAIL.n154 VSUBS 0.015865f
C447 VTAIL.n155 VSUBS 0.035416f
C448 VTAIL.n156 VSUBS 0.035416f
C449 VTAIL.n157 VSUBS 0.015865f
C450 VTAIL.n158 VSUBS 0.014984f
C451 VTAIL.n159 VSUBS 0.027884f
C452 VTAIL.n160 VSUBS 0.027884f
C453 VTAIL.n161 VSUBS 0.014984f
C454 VTAIL.n162 VSUBS 0.015865f
C455 VTAIL.n163 VSUBS 0.035416f
C456 VTAIL.n164 VSUBS 0.035416f
C457 VTAIL.n165 VSUBS 0.015865f
C458 VTAIL.n166 VSUBS 0.014984f
C459 VTAIL.n167 VSUBS 0.027884f
C460 VTAIL.n168 VSUBS 0.027884f
C461 VTAIL.n169 VSUBS 0.014984f
C462 VTAIL.n170 VSUBS 0.015865f
C463 VTAIL.n171 VSUBS 0.035416f
C464 VTAIL.n172 VSUBS 0.035416f
C465 VTAIL.n173 VSUBS 0.015865f
C466 VTAIL.n174 VSUBS 0.014984f
C467 VTAIL.n175 VSUBS 0.027884f
C468 VTAIL.n176 VSUBS 0.027884f
C469 VTAIL.n177 VSUBS 0.014984f
C470 VTAIL.n178 VSUBS 0.015865f
C471 VTAIL.n179 VSUBS 0.035416f
C472 VTAIL.n180 VSUBS 0.035416f
C473 VTAIL.n181 VSUBS 0.015865f
C474 VTAIL.n182 VSUBS 0.014984f
C475 VTAIL.n183 VSUBS 0.027884f
C476 VTAIL.n184 VSUBS 0.027884f
C477 VTAIL.n185 VSUBS 0.014984f
C478 VTAIL.n186 VSUBS 0.015865f
C479 VTAIL.n187 VSUBS 0.035416f
C480 VTAIL.n188 VSUBS 0.035416f
C481 VTAIL.n189 VSUBS 0.015865f
C482 VTAIL.n190 VSUBS 0.014984f
C483 VTAIL.n191 VSUBS 0.027884f
C484 VTAIL.n192 VSUBS 0.027884f
C485 VTAIL.n193 VSUBS 0.014984f
C486 VTAIL.n194 VSUBS 0.015865f
C487 VTAIL.n195 VSUBS 0.035416f
C488 VTAIL.n196 VSUBS 0.089366f
C489 VTAIL.n197 VSUBS 0.015865f
C490 VTAIL.n198 VSUBS 0.014984f
C491 VTAIL.n199 VSUBS 0.069785f
C492 VTAIL.n200 VSUBS 0.045261f
C493 VTAIL.n201 VSUBS 0.4629f
C494 VTAIL.t4 VSUBS 0.38913f
C495 VTAIL.t5 VSUBS 0.38913f
C496 VTAIL.n202 VSUBS 3.0766f
C497 VTAIL.n203 VSUBS 1.09515f
C498 VTAIL.n204 VSUBS 0.031704f
C499 VTAIL.n205 VSUBS 0.027884f
C500 VTAIL.n206 VSUBS 0.014984f
C501 VTAIL.n207 VSUBS 0.035416f
C502 VTAIL.n208 VSUBS 0.015865f
C503 VTAIL.n209 VSUBS 0.027884f
C504 VTAIL.n210 VSUBS 0.014984f
C505 VTAIL.n211 VSUBS 0.035416f
C506 VTAIL.n212 VSUBS 0.015424f
C507 VTAIL.n213 VSUBS 0.027884f
C508 VTAIL.n214 VSUBS 0.015424f
C509 VTAIL.n215 VSUBS 0.014984f
C510 VTAIL.n216 VSUBS 0.035416f
C511 VTAIL.n217 VSUBS 0.035416f
C512 VTAIL.n218 VSUBS 0.015865f
C513 VTAIL.n219 VSUBS 0.027884f
C514 VTAIL.n220 VSUBS 0.014984f
C515 VTAIL.n221 VSUBS 0.035416f
C516 VTAIL.n222 VSUBS 0.015865f
C517 VTAIL.n223 VSUBS 0.027884f
C518 VTAIL.n224 VSUBS 0.014984f
C519 VTAIL.n225 VSUBS 0.035416f
C520 VTAIL.n226 VSUBS 0.015865f
C521 VTAIL.n227 VSUBS 0.027884f
C522 VTAIL.n228 VSUBS 0.014984f
C523 VTAIL.n229 VSUBS 0.035416f
C524 VTAIL.n230 VSUBS 0.015865f
C525 VTAIL.n231 VSUBS 0.027884f
C526 VTAIL.n232 VSUBS 0.014984f
C527 VTAIL.n233 VSUBS 0.035416f
C528 VTAIL.n234 VSUBS 0.015865f
C529 VTAIL.n235 VSUBS 2.11714f
C530 VTAIL.n236 VSUBS 0.014984f
C531 VTAIL.t0 VSUBS 0.076002f
C532 VTAIL.n237 VSUBS 0.218433f
C533 VTAIL.n238 VSUBS 0.02253f
C534 VTAIL.n239 VSUBS 0.026562f
C535 VTAIL.n240 VSUBS 0.035416f
C536 VTAIL.n241 VSUBS 0.015865f
C537 VTAIL.n242 VSUBS 0.014984f
C538 VTAIL.n243 VSUBS 0.027884f
C539 VTAIL.n244 VSUBS 0.027884f
C540 VTAIL.n245 VSUBS 0.014984f
C541 VTAIL.n246 VSUBS 0.015865f
C542 VTAIL.n247 VSUBS 0.035416f
C543 VTAIL.n248 VSUBS 0.035416f
C544 VTAIL.n249 VSUBS 0.015865f
C545 VTAIL.n250 VSUBS 0.014984f
C546 VTAIL.n251 VSUBS 0.027884f
C547 VTAIL.n252 VSUBS 0.027884f
C548 VTAIL.n253 VSUBS 0.014984f
C549 VTAIL.n254 VSUBS 0.015865f
C550 VTAIL.n255 VSUBS 0.035416f
C551 VTAIL.n256 VSUBS 0.035416f
C552 VTAIL.n257 VSUBS 0.015865f
C553 VTAIL.n258 VSUBS 0.014984f
C554 VTAIL.n259 VSUBS 0.027884f
C555 VTAIL.n260 VSUBS 0.027884f
C556 VTAIL.n261 VSUBS 0.014984f
C557 VTAIL.n262 VSUBS 0.015865f
C558 VTAIL.n263 VSUBS 0.035416f
C559 VTAIL.n264 VSUBS 0.035416f
C560 VTAIL.n265 VSUBS 0.015865f
C561 VTAIL.n266 VSUBS 0.014984f
C562 VTAIL.n267 VSUBS 0.027884f
C563 VTAIL.n268 VSUBS 0.027884f
C564 VTAIL.n269 VSUBS 0.014984f
C565 VTAIL.n270 VSUBS 0.015865f
C566 VTAIL.n271 VSUBS 0.035416f
C567 VTAIL.n272 VSUBS 0.035416f
C568 VTAIL.n273 VSUBS 0.015865f
C569 VTAIL.n274 VSUBS 0.014984f
C570 VTAIL.n275 VSUBS 0.027884f
C571 VTAIL.n276 VSUBS 0.027884f
C572 VTAIL.n277 VSUBS 0.014984f
C573 VTAIL.n278 VSUBS 0.015865f
C574 VTAIL.n279 VSUBS 0.035416f
C575 VTAIL.n280 VSUBS 0.035416f
C576 VTAIL.n281 VSUBS 0.015865f
C577 VTAIL.n282 VSUBS 0.014984f
C578 VTAIL.n283 VSUBS 0.027884f
C579 VTAIL.n284 VSUBS 0.027884f
C580 VTAIL.n285 VSUBS 0.014984f
C581 VTAIL.n286 VSUBS 0.015865f
C582 VTAIL.n287 VSUBS 0.035416f
C583 VTAIL.n288 VSUBS 0.035416f
C584 VTAIL.n289 VSUBS 0.015865f
C585 VTAIL.n290 VSUBS 0.014984f
C586 VTAIL.n291 VSUBS 0.027884f
C587 VTAIL.n292 VSUBS 0.027884f
C588 VTAIL.n293 VSUBS 0.014984f
C589 VTAIL.n294 VSUBS 0.015865f
C590 VTAIL.n295 VSUBS 0.035416f
C591 VTAIL.n296 VSUBS 0.089366f
C592 VTAIL.n297 VSUBS 0.015865f
C593 VTAIL.n298 VSUBS 0.014984f
C594 VTAIL.n299 VSUBS 0.069785f
C595 VTAIL.n300 VSUBS 0.045261f
C596 VTAIL.n301 VSUBS 2.29859f
C597 VTAIL.n302 VSUBS 0.031704f
C598 VTAIL.n303 VSUBS 0.027884f
C599 VTAIL.n304 VSUBS 0.014984f
C600 VTAIL.n305 VSUBS 0.035416f
C601 VTAIL.n306 VSUBS 0.015865f
C602 VTAIL.n307 VSUBS 0.027884f
C603 VTAIL.n308 VSUBS 0.014984f
C604 VTAIL.n309 VSUBS 0.035416f
C605 VTAIL.n310 VSUBS 0.015424f
C606 VTAIL.n311 VSUBS 0.027884f
C607 VTAIL.n312 VSUBS 0.015865f
C608 VTAIL.n313 VSUBS 0.035416f
C609 VTAIL.n314 VSUBS 0.015865f
C610 VTAIL.n315 VSUBS 0.027884f
C611 VTAIL.n316 VSUBS 0.014984f
C612 VTAIL.n317 VSUBS 0.035416f
C613 VTAIL.n318 VSUBS 0.015865f
C614 VTAIL.n319 VSUBS 0.027884f
C615 VTAIL.n320 VSUBS 0.014984f
C616 VTAIL.n321 VSUBS 0.035416f
C617 VTAIL.n322 VSUBS 0.015865f
C618 VTAIL.n323 VSUBS 0.027884f
C619 VTAIL.n324 VSUBS 0.014984f
C620 VTAIL.n325 VSUBS 0.035416f
C621 VTAIL.n326 VSUBS 0.015865f
C622 VTAIL.n327 VSUBS 0.027884f
C623 VTAIL.n328 VSUBS 0.014984f
C624 VTAIL.n329 VSUBS 0.035416f
C625 VTAIL.n330 VSUBS 0.015865f
C626 VTAIL.n331 VSUBS 2.11714f
C627 VTAIL.n332 VSUBS 0.014984f
C628 VTAIL.t6 VSUBS 0.076002f
C629 VTAIL.n333 VSUBS 0.218433f
C630 VTAIL.n334 VSUBS 0.02253f
C631 VTAIL.n335 VSUBS 0.026562f
C632 VTAIL.n336 VSUBS 0.035416f
C633 VTAIL.n337 VSUBS 0.015865f
C634 VTAIL.n338 VSUBS 0.014984f
C635 VTAIL.n339 VSUBS 0.027884f
C636 VTAIL.n340 VSUBS 0.027884f
C637 VTAIL.n341 VSUBS 0.014984f
C638 VTAIL.n342 VSUBS 0.015865f
C639 VTAIL.n343 VSUBS 0.035416f
C640 VTAIL.n344 VSUBS 0.035416f
C641 VTAIL.n345 VSUBS 0.015865f
C642 VTAIL.n346 VSUBS 0.014984f
C643 VTAIL.n347 VSUBS 0.027884f
C644 VTAIL.n348 VSUBS 0.027884f
C645 VTAIL.n349 VSUBS 0.014984f
C646 VTAIL.n350 VSUBS 0.015865f
C647 VTAIL.n351 VSUBS 0.035416f
C648 VTAIL.n352 VSUBS 0.035416f
C649 VTAIL.n353 VSUBS 0.015865f
C650 VTAIL.n354 VSUBS 0.014984f
C651 VTAIL.n355 VSUBS 0.027884f
C652 VTAIL.n356 VSUBS 0.027884f
C653 VTAIL.n357 VSUBS 0.014984f
C654 VTAIL.n358 VSUBS 0.015865f
C655 VTAIL.n359 VSUBS 0.035416f
C656 VTAIL.n360 VSUBS 0.035416f
C657 VTAIL.n361 VSUBS 0.015865f
C658 VTAIL.n362 VSUBS 0.014984f
C659 VTAIL.n363 VSUBS 0.027884f
C660 VTAIL.n364 VSUBS 0.027884f
C661 VTAIL.n365 VSUBS 0.014984f
C662 VTAIL.n366 VSUBS 0.015865f
C663 VTAIL.n367 VSUBS 0.035416f
C664 VTAIL.n368 VSUBS 0.035416f
C665 VTAIL.n369 VSUBS 0.015865f
C666 VTAIL.n370 VSUBS 0.014984f
C667 VTAIL.n371 VSUBS 0.027884f
C668 VTAIL.n372 VSUBS 0.027884f
C669 VTAIL.n373 VSUBS 0.014984f
C670 VTAIL.n374 VSUBS 0.014984f
C671 VTAIL.n375 VSUBS 0.015865f
C672 VTAIL.n376 VSUBS 0.035416f
C673 VTAIL.n377 VSUBS 0.035416f
C674 VTAIL.n378 VSUBS 0.035416f
C675 VTAIL.n379 VSUBS 0.015424f
C676 VTAIL.n380 VSUBS 0.014984f
C677 VTAIL.n381 VSUBS 0.027884f
C678 VTAIL.n382 VSUBS 0.027884f
C679 VTAIL.n383 VSUBS 0.014984f
C680 VTAIL.n384 VSUBS 0.015865f
C681 VTAIL.n385 VSUBS 0.035416f
C682 VTAIL.n386 VSUBS 0.035416f
C683 VTAIL.n387 VSUBS 0.015865f
C684 VTAIL.n388 VSUBS 0.014984f
C685 VTAIL.n389 VSUBS 0.027884f
C686 VTAIL.n390 VSUBS 0.027884f
C687 VTAIL.n391 VSUBS 0.014984f
C688 VTAIL.n392 VSUBS 0.015865f
C689 VTAIL.n393 VSUBS 0.035416f
C690 VTAIL.n394 VSUBS 0.089366f
C691 VTAIL.n395 VSUBS 0.015865f
C692 VTAIL.n396 VSUBS 0.014984f
C693 VTAIL.n397 VSUBS 0.069785f
C694 VTAIL.n398 VSUBS 0.045261f
C695 VTAIL.n399 VSUBS 2.22772f
C696 VDD2.n0 VSUBS 0.030911f
C697 VDD2.n1 VSUBS 0.027186f
C698 VDD2.n2 VSUBS 0.014609f
C699 VDD2.n3 VSUBS 0.03453f
C700 VDD2.n4 VSUBS 0.015468f
C701 VDD2.n5 VSUBS 0.027186f
C702 VDD2.n6 VSUBS 0.014609f
C703 VDD2.n7 VSUBS 0.03453f
C704 VDD2.n8 VSUBS 0.015038f
C705 VDD2.n9 VSUBS 0.027186f
C706 VDD2.n10 VSUBS 0.015468f
C707 VDD2.n11 VSUBS 0.03453f
C708 VDD2.n12 VSUBS 0.015468f
C709 VDD2.n13 VSUBS 0.027186f
C710 VDD2.n14 VSUBS 0.014609f
C711 VDD2.n15 VSUBS 0.03453f
C712 VDD2.n16 VSUBS 0.015468f
C713 VDD2.n17 VSUBS 0.027186f
C714 VDD2.n18 VSUBS 0.014609f
C715 VDD2.n19 VSUBS 0.03453f
C716 VDD2.n20 VSUBS 0.015468f
C717 VDD2.n21 VSUBS 0.027186f
C718 VDD2.n22 VSUBS 0.014609f
C719 VDD2.n23 VSUBS 0.03453f
C720 VDD2.n24 VSUBS 0.015468f
C721 VDD2.n25 VSUBS 0.027186f
C722 VDD2.n26 VSUBS 0.014609f
C723 VDD2.n27 VSUBS 0.03453f
C724 VDD2.n28 VSUBS 0.015468f
C725 VDD2.n29 VSUBS 2.06419f
C726 VDD2.n30 VSUBS 0.014609f
C727 VDD2.t2 VSUBS 0.074101f
C728 VDD2.n31 VSUBS 0.21297f
C729 VDD2.n32 VSUBS 0.021966f
C730 VDD2.n33 VSUBS 0.025897f
C731 VDD2.n34 VSUBS 0.03453f
C732 VDD2.n35 VSUBS 0.015468f
C733 VDD2.n36 VSUBS 0.014609f
C734 VDD2.n37 VSUBS 0.027186f
C735 VDD2.n38 VSUBS 0.027186f
C736 VDD2.n39 VSUBS 0.014609f
C737 VDD2.n40 VSUBS 0.015468f
C738 VDD2.n41 VSUBS 0.03453f
C739 VDD2.n42 VSUBS 0.03453f
C740 VDD2.n43 VSUBS 0.015468f
C741 VDD2.n44 VSUBS 0.014609f
C742 VDD2.n45 VSUBS 0.027186f
C743 VDD2.n46 VSUBS 0.027186f
C744 VDD2.n47 VSUBS 0.014609f
C745 VDD2.n48 VSUBS 0.015468f
C746 VDD2.n49 VSUBS 0.03453f
C747 VDD2.n50 VSUBS 0.03453f
C748 VDD2.n51 VSUBS 0.015468f
C749 VDD2.n52 VSUBS 0.014609f
C750 VDD2.n53 VSUBS 0.027186f
C751 VDD2.n54 VSUBS 0.027186f
C752 VDD2.n55 VSUBS 0.014609f
C753 VDD2.n56 VSUBS 0.015468f
C754 VDD2.n57 VSUBS 0.03453f
C755 VDD2.n58 VSUBS 0.03453f
C756 VDD2.n59 VSUBS 0.015468f
C757 VDD2.n60 VSUBS 0.014609f
C758 VDD2.n61 VSUBS 0.027186f
C759 VDD2.n62 VSUBS 0.027186f
C760 VDD2.n63 VSUBS 0.014609f
C761 VDD2.n64 VSUBS 0.015468f
C762 VDD2.n65 VSUBS 0.03453f
C763 VDD2.n66 VSUBS 0.03453f
C764 VDD2.n67 VSUBS 0.015468f
C765 VDD2.n68 VSUBS 0.014609f
C766 VDD2.n69 VSUBS 0.027186f
C767 VDD2.n70 VSUBS 0.027186f
C768 VDD2.n71 VSUBS 0.014609f
C769 VDD2.n72 VSUBS 0.014609f
C770 VDD2.n73 VSUBS 0.015468f
C771 VDD2.n74 VSUBS 0.03453f
C772 VDD2.n75 VSUBS 0.03453f
C773 VDD2.n76 VSUBS 0.03453f
C774 VDD2.n77 VSUBS 0.015038f
C775 VDD2.n78 VSUBS 0.014609f
C776 VDD2.n79 VSUBS 0.027186f
C777 VDD2.n80 VSUBS 0.027186f
C778 VDD2.n81 VSUBS 0.014609f
C779 VDD2.n82 VSUBS 0.015468f
C780 VDD2.n83 VSUBS 0.03453f
C781 VDD2.n84 VSUBS 0.03453f
C782 VDD2.n85 VSUBS 0.015468f
C783 VDD2.n86 VSUBS 0.014609f
C784 VDD2.n87 VSUBS 0.027186f
C785 VDD2.n88 VSUBS 0.027186f
C786 VDD2.n89 VSUBS 0.014609f
C787 VDD2.n90 VSUBS 0.015468f
C788 VDD2.n91 VSUBS 0.03453f
C789 VDD2.n92 VSUBS 0.087131f
C790 VDD2.n93 VSUBS 0.015468f
C791 VDD2.n94 VSUBS 0.014609f
C792 VDD2.n95 VSUBS 0.068039f
C793 VDD2.n96 VSUBS 0.072519f
C794 VDD2.t1 VSUBS 0.379397f
C795 VDD2.t5 VSUBS 0.379397f
C796 VDD2.n97 VSUBS 3.16436f
C797 VDD2.n98 VSUBS 3.81371f
C798 VDD2.n99 VSUBS 0.030911f
C799 VDD2.n100 VSUBS 0.027186f
C800 VDD2.n101 VSUBS 0.014609f
C801 VDD2.n102 VSUBS 0.03453f
C802 VDD2.n103 VSUBS 0.015468f
C803 VDD2.n104 VSUBS 0.027186f
C804 VDD2.n105 VSUBS 0.014609f
C805 VDD2.n106 VSUBS 0.03453f
C806 VDD2.n107 VSUBS 0.015038f
C807 VDD2.n108 VSUBS 0.027186f
C808 VDD2.n109 VSUBS 0.015038f
C809 VDD2.n110 VSUBS 0.014609f
C810 VDD2.n111 VSUBS 0.03453f
C811 VDD2.n112 VSUBS 0.03453f
C812 VDD2.n113 VSUBS 0.015468f
C813 VDD2.n114 VSUBS 0.027186f
C814 VDD2.n115 VSUBS 0.014609f
C815 VDD2.n116 VSUBS 0.03453f
C816 VDD2.n117 VSUBS 0.015468f
C817 VDD2.n118 VSUBS 0.027186f
C818 VDD2.n119 VSUBS 0.014609f
C819 VDD2.n120 VSUBS 0.03453f
C820 VDD2.n121 VSUBS 0.015468f
C821 VDD2.n122 VSUBS 0.027186f
C822 VDD2.n123 VSUBS 0.014609f
C823 VDD2.n124 VSUBS 0.03453f
C824 VDD2.n125 VSUBS 0.015468f
C825 VDD2.n126 VSUBS 0.027186f
C826 VDD2.n127 VSUBS 0.014609f
C827 VDD2.n128 VSUBS 0.03453f
C828 VDD2.n129 VSUBS 0.015468f
C829 VDD2.n130 VSUBS 2.06419f
C830 VDD2.n131 VSUBS 0.014609f
C831 VDD2.t4 VSUBS 0.074101f
C832 VDD2.n132 VSUBS 0.21297f
C833 VDD2.n133 VSUBS 0.021966f
C834 VDD2.n134 VSUBS 0.025897f
C835 VDD2.n135 VSUBS 0.03453f
C836 VDD2.n136 VSUBS 0.015468f
C837 VDD2.n137 VSUBS 0.014609f
C838 VDD2.n138 VSUBS 0.027186f
C839 VDD2.n139 VSUBS 0.027186f
C840 VDD2.n140 VSUBS 0.014609f
C841 VDD2.n141 VSUBS 0.015468f
C842 VDD2.n142 VSUBS 0.03453f
C843 VDD2.n143 VSUBS 0.03453f
C844 VDD2.n144 VSUBS 0.015468f
C845 VDD2.n145 VSUBS 0.014609f
C846 VDD2.n146 VSUBS 0.027186f
C847 VDD2.n147 VSUBS 0.027186f
C848 VDD2.n148 VSUBS 0.014609f
C849 VDD2.n149 VSUBS 0.015468f
C850 VDD2.n150 VSUBS 0.03453f
C851 VDD2.n151 VSUBS 0.03453f
C852 VDD2.n152 VSUBS 0.015468f
C853 VDD2.n153 VSUBS 0.014609f
C854 VDD2.n154 VSUBS 0.027186f
C855 VDD2.n155 VSUBS 0.027186f
C856 VDD2.n156 VSUBS 0.014609f
C857 VDD2.n157 VSUBS 0.015468f
C858 VDD2.n158 VSUBS 0.03453f
C859 VDD2.n159 VSUBS 0.03453f
C860 VDD2.n160 VSUBS 0.015468f
C861 VDD2.n161 VSUBS 0.014609f
C862 VDD2.n162 VSUBS 0.027186f
C863 VDD2.n163 VSUBS 0.027186f
C864 VDD2.n164 VSUBS 0.014609f
C865 VDD2.n165 VSUBS 0.015468f
C866 VDD2.n166 VSUBS 0.03453f
C867 VDD2.n167 VSUBS 0.03453f
C868 VDD2.n168 VSUBS 0.015468f
C869 VDD2.n169 VSUBS 0.014609f
C870 VDD2.n170 VSUBS 0.027186f
C871 VDD2.n171 VSUBS 0.027186f
C872 VDD2.n172 VSUBS 0.014609f
C873 VDD2.n173 VSUBS 0.015468f
C874 VDD2.n174 VSUBS 0.03453f
C875 VDD2.n175 VSUBS 0.03453f
C876 VDD2.n176 VSUBS 0.015468f
C877 VDD2.n177 VSUBS 0.014609f
C878 VDD2.n178 VSUBS 0.027186f
C879 VDD2.n179 VSUBS 0.027186f
C880 VDD2.n180 VSUBS 0.014609f
C881 VDD2.n181 VSUBS 0.015468f
C882 VDD2.n182 VSUBS 0.03453f
C883 VDD2.n183 VSUBS 0.03453f
C884 VDD2.n184 VSUBS 0.015468f
C885 VDD2.n185 VSUBS 0.014609f
C886 VDD2.n186 VSUBS 0.027186f
C887 VDD2.n187 VSUBS 0.027186f
C888 VDD2.n188 VSUBS 0.014609f
C889 VDD2.n189 VSUBS 0.015468f
C890 VDD2.n190 VSUBS 0.03453f
C891 VDD2.n191 VSUBS 0.087131f
C892 VDD2.n192 VSUBS 0.015468f
C893 VDD2.n193 VSUBS 0.014609f
C894 VDD2.n194 VSUBS 0.068039f
C895 VDD2.n195 VSUBS 0.062863f
C896 VDD2.n196 VSUBS 3.39455f
C897 VDD2.t3 VSUBS 0.379397f
C898 VDD2.t0 VSUBS 0.379397f
C899 VDD2.n197 VSUBS 3.16431f
C900 VN.t5 VSUBS 3.70957f
C901 VN.n0 VSUBS 1.38134f
C902 VN.n1 VSUBS 0.024966f
C903 VN.n2 VSUBS 0.032493f
C904 VN.n3 VSUBS 0.283957f
C905 VN.t0 VSUBS 3.70957f
C906 VN.t4 VSUBS 3.99212f
C907 VN.n4 VSUBS 1.31657f
C908 VN.n5 VSUBS 1.37592f
C909 VN.n6 VSUBS 0.046297f
C910 VN.n7 VSUBS 0.046297f
C911 VN.n8 VSUBS 0.024966f
C912 VN.n9 VSUBS 0.024966f
C913 VN.n10 VSUBS 0.024966f
C914 VN.n11 VSUBS 0.040091f
C915 VN.n12 VSUBS 0.046297f
C916 VN.n13 VSUBS 0.041269f
C917 VN.n14 VSUBS 0.040288f
C918 VN.n15 VSUBS 0.053448f
C919 VN.t2 VSUBS 3.70957f
C920 VN.n16 VSUBS 1.38134f
C921 VN.n17 VSUBS 0.024966f
C922 VN.n18 VSUBS 0.032493f
C923 VN.n19 VSUBS 0.283957f
C924 VN.t3 VSUBS 3.70957f
C925 VN.t1 VSUBS 3.99212f
C926 VN.n20 VSUBS 1.31657f
C927 VN.n21 VSUBS 1.37592f
C928 VN.n22 VSUBS 0.046297f
C929 VN.n23 VSUBS 0.046297f
C930 VN.n24 VSUBS 0.024966f
C931 VN.n25 VSUBS 0.024966f
C932 VN.n26 VSUBS 0.024966f
C933 VN.n27 VSUBS 0.040091f
C934 VN.n28 VSUBS 0.046297f
C935 VN.n29 VSUBS 0.041269f
C936 VN.n30 VSUBS 0.040288f
C937 VN.n31 VSUBS 1.62222f
C938 B.n0 VSUBS 0.004803f
C939 B.n1 VSUBS 0.004803f
C940 B.n2 VSUBS 0.007596f
C941 B.n3 VSUBS 0.007596f
C942 B.n4 VSUBS 0.007596f
C943 B.n5 VSUBS 0.007596f
C944 B.n6 VSUBS 0.007596f
C945 B.n7 VSUBS 0.007596f
C946 B.n8 VSUBS 0.007596f
C947 B.n9 VSUBS 0.007596f
C948 B.n10 VSUBS 0.007596f
C949 B.n11 VSUBS 0.007596f
C950 B.n12 VSUBS 0.007596f
C951 B.n13 VSUBS 0.007596f
C952 B.n14 VSUBS 0.007596f
C953 B.n15 VSUBS 0.007596f
C954 B.n16 VSUBS 0.007596f
C955 B.n17 VSUBS 0.007596f
C956 B.n18 VSUBS 0.007596f
C957 B.n19 VSUBS 0.007596f
C958 B.n20 VSUBS 0.007596f
C959 B.n21 VSUBS 0.007596f
C960 B.n22 VSUBS 0.007596f
C961 B.n23 VSUBS 0.007596f
C962 B.n24 VSUBS 0.007596f
C963 B.n25 VSUBS 0.007596f
C964 B.n26 VSUBS 0.018252f
C965 B.n27 VSUBS 0.007596f
C966 B.n28 VSUBS 0.007596f
C967 B.n29 VSUBS 0.007596f
C968 B.n30 VSUBS 0.007596f
C969 B.n31 VSUBS 0.007596f
C970 B.n32 VSUBS 0.007596f
C971 B.n33 VSUBS 0.007596f
C972 B.n34 VSUBS 0.007596f
C973 B.n35 VSUBS 0.007596f
C974 B.n36 VSUBS 0.007596f
C975 B.n37 VSUBS 0.007596f
C976 B.n38 VSUBS 0.007596f
C977 B.n39 VSUBS 0.007596f
C978 B.n40 VSUBS 0.007596f
C979 B.n41 VSUBS 0.007596f
C980 B.n42 VSUBS 0.007596f
C981 B.n43 VSUBS 0.007596f
C982 B.n44 VSUBS 0.007596f
C983 B.n45 VSUBS 0.007596f
C984 B.n46 VSUBS 0.007596f
C985 B.n47 VSUBS 0.007596f
C986 B.n48 VSUBS 0.007596f
C987 B.n49 VSUBS 0.007596f
C988 B.n50 VSUBS 0.007596f
C989 B.n51 VSUBS 0.007596f
C990 B.n52 VSUBS 0.007596f
C991 B.n53 VSUBS 0.007596f
C992 B.n54 VSUBS 0.007596f
C993 B.n55 VSUBS 0.007596f
C994 B.t2 VSUBS 0.372279f
C995 B.t1 VSUBS 0.4138f
C996 B.t0 VSUBS 2.63554f
C997 B.n56 VSUBS 0.647139f
C998 B.n57 VSUBS 0.354088f
C999 B.n58 VSUBS 0.007596f
C1000 B.n59 VSUBS 0.007596f
C1001 B.n60 VSUBS 0.007596f
C1002 B.n61 VSUBS 0.007596f
C1003 B.t11 VSUBS 0.372283f
C1004 B.t10 VSUBS 0.413803f
C1005 B.t9 VSUBS 2.63554f
C1006 B.n62 VSUBS 0.647136f
C1007 B.n63 VSUBS 0.354084f
C1008 B.n64 VSUBS 0.017598f
C1009 B.n65 VSUBS 0.007596f
C1010 B.n66 VSUBS 0.007596f
C1011 B.n67 VSUBS 0.007596f
C1012 B.n68 VSUBS 0.007596f
C1013 B.n69 VSUBS 0.007596f
C1014 B.n70 VSUBS 0.007596f
C1015 B.n71 VSUBS 0.007596f
C1016 B.n72 VSUBS 0.007596f
C1017 B.n73 VSUBS 0.007596f
C1018 B.n74 VSUBS 0.007596f
C1019 B.n75 VSUBS 0.007596f
C1020 B.n76 VSUBS 0.007596f
C1021 B.n77 VSUBS 0.007596f
C1022 B.n78 VSUBS 0.007596f
C1023 B.n79 VSUBS 0.007596f
C1024 B.n80 VSUBS 0.007596f
C1025 B.n81 VSUBS 0.007596f
C1026 B.n82 VSUBS 0.007596f
C1027 B.n83 VSUBS 0.007596f
C1028 B.n84 VSUBS 0.007596f
C1029 B.n85 VSUBS 0.007596f
C1030 B.n86 VSUBS 0.007596f
C1031 B.n87 VSUBS 0.007596f
C1032 B.n88 VSUBS 0.007596f
C1033 B.n89 VSUBS 0.007596f
C1034 B.n90 VSUBS 0.007596f
C1035 B.n91 VSUBS 0.007596f
C1036 B.n92 VSUBS 0.007596f
C1037 B.n93 VSUBS 0.018252f
C1038 B.n94 VSUBS 0.007596f
C1039 B.n95 VSUBS 0.007596f
C1040 B.n96 VSUBS 0.007596f
C1041 B.n97 VSUBS 0.007596f
C1042 B.n98 VSUBS 0.007596f
C1043 B.n99 VSUBS 0.007596f
C1044 B.n100 VSUBS 0.007596f
C1045 B.n101 VSUBS 0.007596f
C1046 B.n102 VSUBS 0.007596f
C1047 B.n103 VSUBS 0.007596f
C1048 B.n104 VSUBS 0.007596f
C1049 B.n105 VSUBS 0.007596f
C1050 B.n106 VSUBS 0.007596f
C1051 B.n107 VSUBS 0.007596f
C1052 B.n108 VSUBS 0.007596f
C1053 B.n109 VSUBS 0.007596f
C1054 B.n110 VSUBS 0.007596f
C1055 B.n111 VSUBS 0.007596f
C1056 B.n112 VSUBS 0.007596f
C1057 B.n113 VSUBS 0.007596f
C1058 B.n114 VSUBS 0.007596f
C1059 B.n115 VSUBS 0.007596f
C1060 B.n116 VSUBS 0.007596f
C1061 B.n117 VSUBS 0.007596f
C1062 B.n118 VSUBS 0.007596f
C1063 B.n119 VSUBS 0.007596f
C1064 B.n120 VSUBS 0.007596f
C1065 B.n121 VSUBS 0.007596f
C1066 B.n122 VSUBS 0.007596f
C1067 B.n123 VSUBS 0.007596f
C1068 B.n124 VSUBS 0.007596f
C1069 B.n125 VSUBS 0.007596f
C1070 B.n126 VSUBS 0.007596f
C1071 B.n127 VSUBS 0.007596f
C1072 B.n128 VSUBS 0.007596f
C1073 B.n129 VSUBS 0.007596f
C1074 B.n130 VSUBS 0.007596f
C1075 B.n131 VSUBS 0.007596f
C1076 B.n132 VSUBS 0.007596f
C1077 B.n133 VSUBS 0.007596f
C1078 B.n134 VSUBS 0.007596f
C1079 B.n135 VSUBS 0.007596f
C1080 B.n136 VSUBS 0.007596f
C1081 B.n137 VSUBS 0.007596f
C1082 B.n138 VSUBS 0.007596f
C1083 B.n139 VSUBS 0.007596f
C1084 B.n140 VSUBS 0.007596f
C1085 B.n141 VSUBS 0.007596f
C1086 B.n142 VSUBS 0.018252f
C1087 B.n143 VSUBS 0.007596f
C1088 B.n144 VSUBS 0.007596f
C1089 B.n145 VSUBS 0.007596f
C1090 B.n146 VSUBS 0.007596f
C1091 B.n147 VSUBS 0.007596f
C1092 B.n148 VSUBS 0.007596f
C1093 B.n149 VSUBS 0.007596f
C1094 B.n150 VSUBS 0.007596f
C1095 B.n151 VSUBS 0.007596f
C1096 B.n152 VSUBS 0.007596f
C1097 B.n153 VSUBS 0.007596f
C1098 B.n154 VSUBS 0.007596f
C1099 B.n155 VSUBS 0.007596f
C1100 B.n156 VSUBS 0.007596f
C1101 B.n157 VSUBS 0.007596f
C1102 B.n158 VSUBS 0.007596f
C1103 B.n159 VSUBS 0.007596f
C1104 B.n160 VSUBS 0.007596f
C1105 B.n161 VSUBS 0.007596f
C1106 B.n162 VSUBS 0.007596f
C1107 B.n163 VSUBS 0.007596f
C1108 B.n164 VSUBS 0.007596f
C1109 B.n165 VSUBS 0.007596f
C1110 B.n166 VSUBS 0.007596f
C1111 B.n167 VSUBS 0.007596f
C1112 B.n168 VSUBS 0.007596f
C1113 B.n169 VSUBS 0.007596f
C1114 B.n170 VSUBS 0.007596f
C1115 B.n171 VSUBS 0.007596f
C1116 B.t7 VSUBS 0.372283f
C1117 B.t8 VSUBS 0.413803f
C1118 B.t6 VSUBS 2.63554f
C1119 B.n172 VSUBS 0.647136f
C1120 B.n173 VSUBS 0.354084f
C1121 B.n174 VSUBS 0.007596f
C1122 B.n175 VSUBS 0.007596f
C1123 B.n176 VSUBS 0.007596f
C1124 B.n177 VSUBS 0.007596f
C1125 B.t4 VSUBS 0.372279f
C1126 B.t5 VSUBS 0.4138f
C1127 B.t3 VSUBS 2.63554f
C1128 B.n178 VSUBS 0.647139f
C1129 B.n179 VSUBS 0.354088f
C1130 B.n180 VSUBS 0.017598f
C1131 B.n181 VSUBS 0.007596f
C1132 B.n182 VSUBS 0.007596f
C1133 B.n183 VSUBS 0.007596f
C1134 B.n184 VSUBS 0.007596f
C1135 B.n185 VSUBS 0.007596f
C1136 B.n186 VSUBS 0.007596f
C1137 B.n187 VSUBS 0.007596f
C1138 B.n188 VSUBS 0.007596f
C1139 B.n189 VSUBS 0.007596f
C1140 B.n190 VSUBS 0.007596f
C1141 B.n191 VSUBS 0.007596f
C1142 B.n192 VSUBS 0.007596f
C1143 B.n193 VSUBS 0.007596f
C1144 B.n194 VSUBS 0.007596f
C1145 B.n195 VSUBS 0.007596f
C1146 B.n196 VSUBS 0.007596f
C1147 B.n197 VSUBS 0.007596f
C1148 B.n198 VSUBS 0.007596f
C1149 B.n199 VSUBS 0.007596f
C1150 B.n200 VSUBS 0.007596f
C1151 B.n201 VSUBS 0.007596f
C1152 B.n202 VSUBS 0.007596f
C1153 B.n203 VSUBS 0.007596f
C1154 B.n204 VSUBS 0.007596f
C1155 B.n205 VSUBS 0.007596f
C1156 B.n206 VSUBS 0.007596f
C1157 B.n207 VSUBS 0.007596f
C1158 B.n208 VSUBS 0.007596f
C1159 B.n209 VSUBS 0.018252f
C1160 B.n210 VSUBS 0.007596f
C1161 B.n211 VSUBS 0.007596f
C1162 B.n212 VSUBS 0.007596f
C1163 B.n213 VSUBS 0.007596f
C1164 B.n214 VSUBS 0.007596f
C1165 B.n215 VSUBS 0.007596f
C1166 B.n216 VSUBS 0.007596f
C1167 B.n217 VSUBS 0.007596f
C1168 B.n218 VSUBS 0.007596f
C1169 B.n219 VSUBS 0.007596f
C1170 B.n220 VSUBS 0.007596f
C1171 B.n221 VSUBS 0.007596f
C1172 B.n222 VSUBS 0.007596f
C1173 B.n223 VSUBS 0.007596f
C1174 B.n224 VSUBS 0.007596f
C1175 B.n225 VSUBS 0.007596f
C1176 B.n226 VSUBS 0.007596f
C1177 B.n227 VSUBS 0.007596f
C1178 B.n228 VSUBS 0.007596f
C1179 B.n229 VSUBS 0.007596f
C1180 B.n230 VSUBS 0.007596f
C1181 B.n231 VSUBS 0.007596f
C1182 B.n232 VSUBS 0.007596f
C1183 B.n233 VSUBS 0.007596f
C1184 B.n234 VSUBS 0.007596f
C1185 B.n235 VSUBS 0.007596f
C1186 B.n236 VSUBS 0.007596f
C1187 B.n237 VSUBS 0.007596f
C1188 B.n238 VSUBS 0.007596f
C1189 B.n239 VSUBS 0.007596f
C1190 B.n240 VSUBS 0.007596f
C1191 B.n241 VSUBS 0.007596f
C1192 B.n242 VSUBS 0.007596f
C1193 B.n243 VSUBS 0.007596f
C1194 B.n244 VSUBS 0.007596f
C1195 B.n245 VSUBS 0.007596f
C1196 B.n246 VSUBS 0.007596f
C1197 B.n247 VSUBS 0.007596f
C1198 B.n248 VSUBS 0.007596f
C1199 B.n249 VSUBS 0.007596f
C1200 B.n250 VSUBS 0.007596f
C1201 B.n251 VSUBS 0.007596f
C1202 B.n252 VSUBS 0.007596f
C1203 B.n253 VSUBS 0.007596f
C1204 B.n254 VSUBS 0.007596f
C1205 B.n255 VSUBS 0.007596f
C1206 B.n256 VSUBS 0.007596f
C1207 B.n257 VSUBS 0.007596f
C1208 B.n258 VSUBS 0.007596f
C1209 B.n259 VSUBS 0.007596f
C1210 B.n260 VSUBS 0.007596f
C1211 B.n261 VSUBS 0.007596f
C1212 B.n262 VSUBS 0.007596f
C1213 B.n263 VSUBS 0.007596f
C1214 B.n264 VSUBS 0.007596f
C1215 B.n265 VSUBS 0.007596f
C1216 B.n266 VSUBS 0.007596f
C1217 B.n267 VSUBS 0.007596f
C1218 B.n268 VSUBS 0.007596f
C1219 B.n269 VSUBS 0.007596f
C1220 B.n270 VSUBS 0.007596f
C1221 B.n271 VSUBS 0.007596f
C1222 B.n272 VSUBS 0.007596f
C1223 B.n273 VSUBS 0.007596f
C1224 B.n274 VSUBS 0.007596f
C1225 B.n275 VSUBS 0.007596f
C1226 B.n276 VSUBS 0.007596f
C1227 B.n277 VSUBS 0.007596f
C1228 B.n278 VSUBS 0.007596f
C1229 B.n279 VSUBS 0.007596f
C1230 B.n280 VSUBS 0.007596f
C1231 B.n281 VSUBS 0.007596f
C1232 B.n282 VSUBS 0.007596f
C1233 B.n283 VSUBS 0.007596f
C1234 B.n284 VSUBS 0.007596f
C1235 B.n285 VSUBS 0.007596f
C1236 B.n286 VSUBS 0.007596f
C1237 B.n287 VSUBS 0.007596f
C1238 B.n288 VSUBS 0.007596f
C1239 B.n289 VSUBS 0.007596f
C1240 B.n290 VSUBS 0.007596f
C1241 B.n291 VSUBS 0.007596f
C1242 B.n292 VSUBS 0.007596f
C1243 B.n293 VSUBS 0.007596f
C1244 B.n294 VSUBS 0.007596f
C1245 B.n295 VSUBS 0.007596f
C1246 B.n296 VSUBS 0.007596f
C1247 B.n297 VSUBS 0.007596f
C1248 B.n298 VSUBS 0.007596f
C1249 B.n299 VSUBS 0.007596f
C1250 B.n300 VSUBS 0.007596f
C1251 B.n301 VSUBS 0.007596f
C1252 B.n302 VSUBS 0.017492f
C1253 B.n303 VSUBS 0.017492f
C1254 B.n304 VSUBS 0.018252f
C1255 B.n305 VSUBS 0.007596f
C1256 B.n306 VSUBS 0.007596f
C1257 B.n307 VSUBS 0.007596f
C1258 B.n308 VSUBS 0.007596f
C1259 B.n309 VSUBS 0.007596f
C1260 B.n310 VSUBS 0.007596f
C1261 B.n311 VSUBS 0.007596f
C1262 B.n312 VSUBS 0.007596f
C1263 B.n313 VSUBS 0.007596f
C1264 B.n314 VSUBS 0.007596f
C1265 B.n315 VSUBS 0.007596f
C1266 B.n316 VSUBS 0.007596f
C1267 B.n317 VSUBS 0.007596f
C1268 B.n318 VSUBS 0.007596f
C1269 B.n319 VSUBS 0.007596f
C1270 B.n320 VSUBS 0.007596f
C1271 B.n321 VSUBS 0.007596f
C1272 B.n322 VSUBS 0.007596f
C1273 B.n323 VSUBS 0.007596f
C1274 B.n324 VSUBS 0.007596f
C1275 B.n325 VSUBS 0.007596f
C1276 B.n326 VSUBS 0.007596f
C1277 B.n327 VSUBS 0.007596f
C1278 B.n328 VSUBS 0.007596f
C1279 B.n329 VSUBS 0.007596f
C1280 B.n330 VSUBS 0.007596f
C1281 B.n331 VSUBS 0.007596f
C1282 B.n332 VSUBS 0.007596f
C1283 B.n333 VSUBS 0.007596f
C1284 B.n334 VSUBS 0.007596f
C1285 B.n335 VSUBS 0.007596f
C1286 B.n336 VSUBS 0.007596f
C1287 B.n337 VSUBS 0.007596f
C1288 B.n338 VSUBS 0.007596f
C1289 B.n339 VSUBS 0.007596f
C1290 B.n340 VSUBS 0.007596f
C1291 B.n341 VSUBS 0.007596f
C1292 B.n342 VSUBS 0.007596f
C1293 B.n343 VSUBS 0.007596f
C1294 B.n344 VSUBS 0.007596f
C1295 B.n345 VSUBS 0.007596f
C1296 B.n346 VSUBS 0.007596f
C1297 B.n347 VSUBS 0.007596f
C1298 B.n348 VSUBS 0.007596f
C1299 B.n349 VSUBS 0.007596f
C1300 B.n350 VSUBS 0.007596f
C1301 B.n351 VSUBS 0.007596f
C1302 B.n352 VSUBS 0.007596f
C1303 B.n353 VSUBS 0.007596f
C1304 B.n354 VSUBS 0.007596f
C1305 B.n355 VSUBS 0.007596f
C1306 B.n356 VSUBS 0.007596f
C1307 B.n357 VSUBS 0.007596f
C1308 B.n358 VSUBS 0.007596f
C1309 B.n359 VSUBS 0.007596f
C1310 B.n360 VSUBS 0.007596f
C1311 B.n361 VSUBS 0.007596f
C1312 B.n362 VSUBS 0.007596f
C1313 B.n363 VSUBS 0.007596f
C1314 B.n364 VSUBS 0.007596f
C1315 B.n365 VSUBS 0.007596f
C1316 B.n366 VSUBS 0.007596f
C1317 B.n367 VSUBS 0.007596f
C1318 B.n368 VSUBS 0.007596f
C1319 B.n369 VSUBS 0.007596f
C1320 B.n370 VSUBS 0.007596f
C1321 B.n371 VSUBS 0.007596f
C1322 B.n372 VSUBS 0.007596f
C1323 B.n373 VSUBS 0.007596f
C1324 B.n374 VSUBS 0.007596f
C1325 B.n375 VSUBS 0.007596f
C1326 B.n376 VSUBS 0.007596f
C1327 B.n377 VSUBS 0.007596f
C1328 B.n378 VSUBS 0.007596f
C1329 B.n379 VSUBS 0.007596f
C1330 B.n380 VSUBS 0.007596f
C1331 B.n381 VSUBS 0.007596f
C1332 B.n382 VSUBS 0.007596f
C1333 B.n383 VSUBS 0.007596f
C1334 B.n384 VSUBS 0.007596f
C1335 B.n385 VSUBS 0.007596f
C1336 B.n386 VSUBS 0.007596f
C1337 B.n387 VSUBS 0.007596f
C1338 B.n388 VSUBS 0.007596f
C1339 B.n389 VSUBS 0.007149f
C1340 B.n390 VSUBS 0.007596f
C1341 B.n391 VSUBS 0.007596f
C1342 B.n392 VSUBS 0.004245f
C1343 B.n393 VSUBS 0.007596f
C1344 B.n394 VSUBS 0.007596f
C1345 B.n395 VSUBS 0.007596f
C1346 B.n396 VSUBS 0.007596f
C1347 B.n397 VSUBS 0.007596f
C1348 B.n398 VSUBS 0.007596f
C1349 B.n399 VSUBS 0.007596f
C1350 B.n400 VSUBS 0.007596f
C1351 B.n401 VSUBS 0.007596f
C1352 B.n402 VSUBS 0.007596f
C1353 B.n403 VSUBS 0.007596f
C1354 B.n404 VSUBS 0.007596f
C1355 B.n405 VSUBS 0.004245f
C1356 B.n406 VSUBS 0.017598f
C1357 B.n407 VSUBS 0.007149f
C1358 B.n408 VSUBS 0.007596f
C1359 B.n409 VSUBS 0.007596f
C1360 B.n410 VSUBS 0.007596f
C1361 B.n411 VSUBS 0.007596f
C1362 B.n412 VSUBS 0.007596f
C1363 B.n413 VSUBS 0.007596f
C1364 B.n414 VSUBS 0.007596f
C1365 B.n415 VSUBS 0.007596f
C1366 B.n416 VSUBS 0.007596f
C1367 B.n417 VSUBS 0.007596f
C1368 B.n418 VSUBS 0.007596f
C1369 B.n419 VSUBS 0.007596f
C1370 B.n420 VSUBS 0.007596f
C1371 B.n421 VSUBS 0.007596f
C1372 B.n422 VSUBS 0.007596f
C1373 B.n423 VSUBS 0.007596f
C1374 B.n424 VSUBS 0.007596f
C1375 B.n425 VSUBS 0.007596f
C1376 B.n426 VSUBS 0.007596f
C1377 B.n427 VSUBS 0.007596f
C1378 B.n428 VSUBS 0.007596f
C1379 B.n429 VSUBS 0.007596f
C1380 B.n430 VSUBS 0.007596f
C1381 B.n431 VSUBS 0.007596f
C1382 B.n432 VSUBS 0.007596f
C1383 B.n433 VSUBS 0.007596f
C1384 B.n434 VSUBS 0.007596f
C1385 B.n435 VSUBS 0.007596f
C1386 B.n436 VSUBS 0.007596f
C1387 B.n437 VSUBS 0.007596f
C1388 B.n438 VSUBS 0.007596f
C1389 B.n439 VSUBS 0.007596f
C1390 B.n440 VSUBS 0.007596f
C1391 B.n441 VSUBS 0.007596f
C1392 B.n442 VSUBS 0.007596f
C1393 B.n443 VSUBS 0.007596f
C1394 B.n444 VSUBS 0.007596f
C1395 B.n445 VSUBS 0.007596f
C1396 B.n446 VSUBS 0.007596f
C1397 B.n447 VSUBS 0.007596f
C1398 B.n448 VSUBS 0.007596f
C1399 B.n449 VSUBS 0.007596f
C1400 B.n450 VSUBS 0.007596f
C1401 B.n451 VSUBS 0.007596f
C1402 B.n452 VSUBS 0.007596f
C1403 B.n453 VSUBS 0.007596f
C1404 B.n454 VSUBS 0.007596f
C1405 B.n455 VSUBS 0.007596f
C1406 B.n456 VSUBS 0.007596f
C1407 B.n457 VSUBS 0.007596f
C1408 B.n458 VSUBS 0.007596f
C1409 B.n459 VSUBS 0.007596f
C1410 B.n460 VSUBS 0.007596f
C1411 B.n461 VSUBS 0.007596f
C1412 B.n462 VSUBS 0.007596f
C1413 B.n463 VSUBS 0.007596f
C1414 B.n464 VSUBS 0.007596f
C1415 B.n465 VSUBS 0.007596f
C1416 B.n466 VSUBS 0.007596f
C1417 B.n467 VSUBS 0.007596f
C1418 B.n468 VSUBS 0.007596f
C1419 B.n469 VSUBS 0.007596f
C1420 B.n470 VSUBS 0.007596f
C1421 B.n471 VSUBS 0.007596f
C1422 B.n472 VSUBS 0.007596f
C1423 B.n473 VSUBS 0.007596f
C1424 B.n474 VSUBS 0.007596f
C1425 B.n475 VSUBS 0.007596f
C1426 B.n476 VSUBS 0.007596f
C1427 B.n477 VSUBS 0.007596f
C1428 B.n478 VSUBS 0.007596f
C1429 B.n479 VSUBS 0.007596f
C1430 B.n480 VSUBS 0.007596f
C1431 B.n481 VSUBS 0.007596f
C1432 B.n482 VSUBS 0.007596f
C1433 B.n483 VSUBS 0.007596f
C1434 B.n484 VSUBS 0.007596f
C1435 B.n485 VSUBS 0.007596f
C1436 B.n486 VSUBS 0.007596f
C1437 B.n487 VSUBS 0.007596f
C1438 B.n488 VSUBS 0.007596f
C1439 B.n489 VSUBS 0.007596f
C1440 B.n490 VSUBS 0.007596f
C1441 B.n491 VSUBS 0.007596f
C1442 B.n492 VSUBS 0.007596f
C1443 B.n493 VSUBS 0.018252f
C1444 B.n494 VSUBS 0.017492f
C1445 B.n495 VSUBS 0.017492f
C1446 B.n496 VSUBS 0.007596f
C1447 B.n497 VSUBS 0.007596f
C1448 B.n498 VSUBS 0.007596f
C1449 B.n499 VSUBS 0.007596f
C1450 B.n500 VSUBS 0.007596f
C1451 B.n501 VSUBS 0.007596f
C1452 B.n502 VSUBS 0.007596f
C1453 B.n503 VSUBS 0.007596f
C1454 B.n504 VSUBS 0.007596f
C1455 B.n505 VSUBS 0.007596f
C1456 B.n506 VSUBS 0.007596f
C1457 B.n507 VSUBS 0.007596f
C1458 B.n508 VSUBS 0.007596f
C1459 B.n509 VSUBS 0.007596f
C1460 B.n510 VSUBS 0.007596f
C1461 B.n511 VSUBS 0.007596f
C1462 B.n512 VSUBS 0.007596f
C1463 B.n513 VSUBS 0.007596f
C1464 B.n514 VSUBS 0.007596f
C1465 B.n515 VSUBS 0.007596f
C1466 B.n516 VSUBS 0.007596f
C1467 B.n517 VSUBS 0.007596f
C1468 B.n518 VSUBS 0.007596f
C1469 B.n519 VSUBS 0.007596f
C1470 B.n520 VSUBS 0.007596f
C1471 B.n521 VSUBS 0.007596f
C1472 B.n522 VSUBS 0.007596f
C1473 B.n523 VSUBS 0.007596f
C1474 B.n524 VSUBS 0.007596f
C1475 B.n525 VSUBS 0.007596f
C1476 B.n526 VSUBS 0.007596f
C1477 B.n527 VSUBS 0.007596f
C1478 B.n528 VSUBS 0.007596f
C1479 B.n529 VSUBS 0.007596f
C1480 B.n530 VSUBS 0.007596f
C1481 B.n531 VSUBS 0.007596f
C1482 B.n532 VSUBS 0.007596f
C1483 B.n533 VSUBS 0.007596f
C1484 B.n534 VSUBS 0.007596f
C1485 B.n535 VSUBS 0.007596f
C1486 B.n536 VSUBS 0.007596f
C1487 B.n537 VSUBS 0.007596f
C1488 B.n538 VSUBS 0.007596f
C1489 B.n539 VSUBS 0.007596f
C1490 B.n540 VSUBS 0.007596f
C1491 B.n541 VSUBS 0.007596f
C1492 B.n542 VSUBS 0.007596f
C1493 B.n543 VSUBS 0.007596f
C1494 B.n544 VSUBS 0.007596f
C1495 B.n545 VSUBS 0.007596f
C1496 B.n546 VSUBS 0.007596f
C1497 B.n547 VSUBS 0.007596f
C1498 B.n548 VSUBS 0.007596f
C1499 B.n549 VSUBS 0.007596f
C1500 B.n550 VSUBS 0.007596f
C1501 B.n551 VSUBS 0.007596f
C1502 B.n552 VSUBS 0.007596f
C1503 B.n553 VSUBS 0.007596f
C1504 B.n554 VSUBS 0.007596f
C1505 B.n555 VSUBS 0.007596f
C1506 B.n556 VSUBS 0.007596f
C1507 B.n557 VSUBS 0.007596f
C1508 B.n558 VSUBS 0.007596f
C1509 B.n559 VSUBS 0.007596f
C1510 B.n560 VSUBS 0.007596f
C1511 B.n561 VSUBS 0.007596f
C1512 B.n562 VSUBS 0.007596f
C1513 B.n563 VSUBS 0.007596f
C1514 B.n564 VSUBS 0.007596f
C1515 B.n565 VSUBS 0.007596f
C1516 B.n566 VSUBS 0.007596f
C1517 B.n567 VSUBS 0.007596f
C1518 B.n568 VSUBS 0.007596f
C1519 B.n569 VSUBS 0.007596f
C1520 B.n570 VSUBS 0.007596f
C1521 B.n571 VSUBS 0.007596f
C1522 B.n572 VSUBS 0.007596f
C1523 B.n573 VSUBS 0.007596f
C1524 B.n574 VSUBS 0.007596f
C1525 B.n575 VSUBS 0.007596f
C1526 B.n576 VSUBS 0.007596f
C1527 B.n577 VSUBS 0.007596f
C1528 B.n578 VSUBS 0.007596f
C1529 B.n579 VSUBS 0.007596f
C1530 B.n580 VSUBS 0.007596f
C1531 B.n581 VSUBS 0.007596f
C1532 B.n582 VSUBS 0.007596f
C1533 B.n583 VSUBS 0.007596f
C1534 B.n584 VSUBS 0.007596f
C1535 B.n585 VSUBS 0.007596f
C1536 B.n586 VSUBS 0.007596f
C1537 B.n587 VSUBS 0.007596f
C1538 B.n588 VSUBS 0.007596f
C1539 B.n589 VSUBS 0.007596f
C1540 B.n590 VSUBS 0.007596f
C1541 B.n591 VSUBS 0.007596f
C1542 B.n592 VSUBS 0.007596f
C1543 B.n593 VSUBS 0.007596f
C1544 B.n594 VSUBS 0.007596f
C1545 B.n595 VSUBS 0.007596f
C1546 B.n596 VSUBS 0.007596f
C1547 B.n597 VSUBS 0.007596f
C1548 B.n598 VSUBS 0.007596f
C1549 B.n599 VSUBS 0.007596f
C1550 B.n600 VSUBS 0.007596f
C1551 B.n601 VSUBS 0.007596f
C1552 B.n602 VSUBS 0.007596f
C1553 B.n603 VSUBS 0.007596f
C1554 B.n604 VSUBS 0.007596f
C1555 B.n605 VSUBS 0.007596f
C1556 B.n606 VSUBS 0.007596f
C1557 B.n607 VSUBS 0.007596f
C1558 B.n608 VSUBS 0.007596f
C1559 B.n609 VSUBS 0.007596f
C1560 B.n610 VSUBS 0.007596f
C1561 B.n611 VSUBS 0.007596f
C1562 B.n612 VSUBS 0.007596f
C1563 B.n613 VSUBS 0.007596f
C1564 B.n614 VSUBS 0.007596f
C1565 B.n615 VSUBS 0.007596f
C1566 B.n616 VSUBS 0.007596f
C1567 B.n617 VSUBS 0.007596f
C1568 B.n618 VSUBS 0.007596f
C1569 B.n619 VSUBS 0.007596f
C1570 B.n620 VSUBS 0.007596f
C1571 B.n621 VSUBS 0.007596f
C1572 B.n622 VSUBS 0.007596f
C1573 B.n623 VSUBS 0.007596f
C1574 B.n624 VSUBS 0.007596f
C1575 B.n625 VSUBS 0.007596f
C1576 B.n626 VSUBS 0.007596f
C1577 B.n627 VSUBS 0.007596f
C1578 B.n628 VSUBS 0.007596f
C1579 B.n629 VSUBS 0.007596f
C1580 B.n630 VSUBS 0.007596f
C1581 B.n631 VSUBS 0.007596f
C1582 B.n632 VSUBS 0.007596f
C1583 B.n633 VSUBS 0.007596f
C1584 B.n634 VSUBS 0.007596f
C1585 B.n635 VSUBS 0.007596f
C1586 B.n636 VSUBS 0.007596f
C1587 B.n637 VSUBS 0.007596f
C1588 B.n638 VSUBS 0.017492f
C1589 B.n639 VSUBS 0.018382f
C1590 B.n640 VSUBS 0.017362f
C1591 B.n641 VSUBS 0.007596f
C1592 B.n642 VSUBS 0.007596f
C1593 B.n643 VSUBS 0.007596f
C1594 B.n644 VSUBS 0.007596f
C1595 B.n645 VSUBS 0.007596f
C1596 B.n646 VSUBS 0.007596f
C1597 B.n647 VSUBS 0.007596f
C1598 B.n648 VSUBS 0.007596f
C1599 B.n649 VSUBS 0.007596f
C1600 B.n650 VSUBS 0.007596f
C1601 B.n651 VSUBS 0.007596f
C1602 B.n652 VSUBS 0.007596f
C1603 B.n653 VSUBS 0.007596f
C1604 B.n654 VSUBS 0.007596f
C1605 B.n655 VSUBS 0.007596f
C1606 B.n656 VSUBS 0.007596f
C1607 B.n657 VSUBS 0.007596f
C1608 B.n658 VSUBS 0.007596f
C1609 B.n659 VSUBS 0.007596f
C1610 B.n660 VSUBS 0.007596f
C1611 B.n661 VSUBS 0.007596f
C1612 B.n662 VSUBS 0.007596f
C1613 B.n663 VSUBS 0.007596f
C1614 B.n664 VSUBS 0.007596f
C1615 B.n665 VSUBS 0.007596f
C1616 B.n666 VSUBS 0.007596f
C1617 B.n667 VSUBS 0.007596f
C1618 B.n668 VSUBS 0.007596f
C1619 B.n669 VSUBS 0.007596f
C1620 B.n670 VSUBS 0.007596f
C1621 B.n671 VSUBS 0.007596f
C1622 B.n672 VSUBS 0.007596f
C1623 B.n673 VSUBS 0.007596f
C1624 B.n674 VSUBS 0.007596f
C1625 B.n675 VSUBS 0.007596f
C1626 B.n676 VSUBS 0.007596f
C1627 B.n677 VSUBS 0.007596f
C1628 B.n678 VSUBS 0.007596f
C1629 B.n679 VSUBS 0.007596f
C1630 B.n680 VSUBS 0.007596f
C1631 B.n681 VSUBS 0.007596f
C1632 B.n682 VSUBS 0.007596f
C1633 B.n683 VSUBS 0.007596f
C1634 B.n684 VSUBS 0.007596f
C1635 B.n685 VSUBS 0.007596f
C1636 B.n686 VSUBS 0.007596f
C1637 B.n687 VSUBS 0.007596f
C1638 B.n688 VSUBS 0.007596f
C1639 B.n689 VSUBS 0.007596f
C1640 B.n690 VSUBS 0.007596f
C1641 B.n691 VSUBS 0.007596f
C1642 B.n692 VSUBS 0.007596f
C1643 B.n693 VSUBS 0.007596f
C1644 B.n694 VSUBS 0.007596f
C1645 B.n695 VSUBS 0.007596f
C1646 B.n696 VSUBS 0.007596f
C1647 B.n697 VSUBS 0.007596f
C1648 B.n698 VSUBS 0.007596f
C1649 B.n699 VSUBS 0.007596f
C1650 B.n700 VSUBS 0.007596f
C1651 B.n701 VSUBS 0.007596f
C1652 B.n702 VSUBS 0.007596f
C1653 B.n703 VSUBS 0.007596f
C1654 B.n704 VSUBS 0.007596f
C1655 B.n705 VSUBS 0.007596f
C1656 B.n706 VSUBS 0.007596f
C1657 B.n707 VSUBS 0.007596f
C1658 B.n708 VSUBS 0.007596f
C1659 B.n709 VSUBS 0.007596f
C1660 B.n710 VSUBS 0.007596f
C1661 B.n711 VSUBS 0.007596f
C1662 B.n712 VSUBS 0.007596f
C1663 B.n713 VSUBS 0.007596f
C1664 B.n714 VSUBS 0.007596f
C1665 B.n715 VSUBS 0.007596f
C1666 B.n716 VSUBS 0.007596f
C1667 B.n717 VSUBS 0.007596f
C1668 B.n718 VSUBS 0.007596f
C1669 B.n719 VSUBS 0.007596f
C1670 B.n720 VSUBS 0.007596f
C1671 B.n721 VSUBS 0.007596f
C1672 B.n722 VSUBS 0.007596f
C1673 B.n723 VSUBS 0.007596f
C1674 B.n724 VSUBS 0.007596f
C1675 B.n725 VSUBS 0.007149f
C1676 B.n726 VSUBS 0.007596f
C1677 B.n727 VSUBS 0.007596f
C1678 B.n728 VSUBS 0.004245f
C1679 B.n729 VSUBS 0.007596f
C1680 B.n730 VSUBS 0.007596f
C1681 B.n731 VSUBS 0.007596f
C1682 B.n732 VSUBS 0.007596f
C1683 B.n733 VSUBS 0.007596f
C1684 B.n734 VSUBS 0.007596f
C1685 B.n735 VSUBS 0.007596f
C1686 B.n736 VSUBS 0.007596f
C1687 B.n737 VSUBS 0.007596f
C1688 B.n738 VSUBS 0.007596f
C1689 B.n739 VSUBS 0.007596f
C1690 B.n740 VSUBS 0.007596f
C1691 B.n741 VSUBS 0.004245f
C1692 B.n742 VSUBS 0.017598f
C1693 B.n743 VSUBS 0.007149f
C1694 B.n744 VSUBS 0.007596f
C1695 B.n745 VSUBS 0.007596f
C1696 B.n746 VSUBS 0.007596f
C1697 B.n747 VSUBS 0.007596f
C1698 B.n748 VSUBS 0.007596f
C1699 B.n749 VSUBS 0.007596f
C1700 B.n750 VSUBS 0.007596f
C1701 B.n751 VSUBS 0.007596f
C1702 B.n752 VSUBS 0.007596f
C1703 B.n753 VSUBS 0.007596f
C1704 B.n754 VSUBS 0.007596f
C1705 B.n755 VSUBS 0.007596f
C1706 B.n756 VSUBS 0.007596f
C1707 B.n757 VSUBS 0.007596f
C1708 B.n758 VSUBS 0.007596f
C1709 B.n759 VSUBS 0.007596f
C1710 B.n760 VSUBS 0.007596f
C1711 B.n761 VSUBS 0.007596f
C1712 B.n762 VSUBS 0.007596f
C1713 B.n763 VSUBS 0.007596f
C1714 B.n764 VSUBS 0.007596f
C1715 B.n765 VSUBS 0.007596f
C1716 B.n766 VSUBS 0.007596f
C1717 B.n767 VSUBS 0.007596f
C1718 B.n768 VSUBS 0.007596f
C1719 B.n769 VSUBS 0.007596f
C1720 B.n770 VSUBS 0.007596f
C1721 B.n771 VSUBS 0.007596f
C1722 B.n772 VSUBS 0.007596f
C1723 B.n773 VSUBS 0.007596f
C1724 B.n774 VSUBS 0.007596f
C1725 B.n775 VSUBS 0.007596f
C1726 B.n776 VSUBS 0.007596f
C1727 B.n777 VSUBS 0.007596f
C1728 B.n778 VSUBS 0.007596f
C1729 B.n779 VSUBS 0.007596f
C1730 B.n780 VSUBS 0.007596f
C1731 B.n781 VSUBS 0.007596f
C1732 B.n782 VSUBS 0.007596f
C1733 B.n783 VSUBS 0.007596f
C1734 B.n784 VSUBS 0.007596f
C1735 B.n785 VSUBS 0.007596f
C1736 B.n786 VSUBS 0.007596f
C1737 B.n787 VSUBS 0.007596f
C1738 B.n788 VSUBS 0.007596f
C1739 B.n789 VSUBS 0.007596f
C1740 B.n790 VSUBS 0.007596f
C1741 B.n791 VSUBS 0.007596f
C1742 B.n792 VSUBS 0.007596f
C1743 B.n793 VSUBS 0.007596f
C1744 B.n794 VSUBS 0.007596f
C1745 B.n795 VSUBS 0.007596f
C1746 B.n796 VSUBS 0.007596f
C1747 B.n797 VSUBS 0.007596f
C1748 B.n798 VSUBS 0.007596f
C1749 B.n799 VSUBS 0.007596f
C1750 B.n800 VSUBS 0.007596f
C1751 B.n801 VSUBS 0.007596f
C1752 B.n802 VSUBS 0.007596f
C1753 B.n803 VSUBS 0.007596f
C1754 B.n804 VSUBS 0.007596f
C1755 B.n805 VSUBS 0.007596f
C1756 B.n806 VSUBS 0.007596f
C1757 B.n807 VSUBS 0.007596f
C1758 B.n808 VSUBS 0.007596f
C1759 B.n809 VSUBS 0.007596f
C1760 B.n810 VSUBS 0.007596f
C1761 B.n811 VSUBS 0.007596f
C1762 B.n812 VSUBS 0.007596f
C1763 B.n813 VSUBS 0.007596f
C1764 B.n814 VSUBS 0.007596f
C1765 B.n815 VSUBS 0.007596f
C1766 B.n816 VSUBS 0.007596f
C1767 B.n817 VSUBS 0.007596f
C1768 B.n818 VSUBS 0.007596f
C1769 B.n819 VSUBS 0.007596f
C1770 B.n820 VSUBS 0.007596f
C1771 B.n821 VSUBS 0.007596f
C1772 B.n822 VSUBS 0.007596f
C1773 B.n823 VSUBS 0.007596f
C1774 B.n824 VSUBS 0.007596f
C1775 B.n825 VSUBS 0.007596f
C1776 B.n826 VSUBS 0.007596f
C1777 B.n827 VSUBS 0.007596f
C1778 B.n828 VSUBS 0.007596f
C1779 B.n829 VSUBS 0.018252f
C1780 B.n830 VSUBS 0.017492f
C1781 B.n831 VSUBS 0.017492f
C1782 B.n832 VSUBS 0.007596f
C1783 B.n833 VSUBS 0.007596f
C1784 B.n834 VSUBS 0.007596f
C1785 B.n835 VSUBS 0.007596f
C1786 B.n836 VSUBS 0.007596f
C1787 B.n837 VSUBS 0.007596f
C1788 B.n838 VSUBS 0.007596f
C1789 B.n839 VSUBS 0.007596f
C1790 B.n840 VSUBS 0.007596f
C1791 B.n841 VSUBS 0.007596f
C1792 B.n842 VSUBS 0.007596f
C1793 B.n843 VSUBS 0.007596f
C1794 B.n844 VSUBS 0.007596f
C1795 B.n845 VSUBS 0.007596f
C1796 B.n846 VSUBS 0.007596f
C1797 B.n847 VSUBS 0.007596f
C1798 B.n848 VSUBS 0.007596f
C1799 B.n849 VSUBS 0.007596f
C1800 B.n850 VSUBS 0.007596f
C1801 B.n851 VSUBS 0.007596f
C1802 B.n852 VSUBS 0.007596f
C1803 B.n853 VSUBS 0.007596f
C1804 B.n854 VSUBS 0.007596f
C1805 B.n855 VSUBS 0.007596f
C1806 B.n856 VSUBS 0.007596f
C1807 B.n857 VSUBS 0.007596f
C1808 B.n858 VSUBS 0.007596f
C1809 B.n859 VSUBS 0.007596f
C1810 B.n860 VSUBS 0.007596f
C1811 B.n861 VSUBS 0.007596f
C1812 B.n862 VSUBS 0.007596f
C1813 B.n863 VSUBS 0.007596f
C1814 B.n864 VSUBS 0.007596f
C1815 B.n865 VSUBS 0.007596f
C1816 B.n866 VSUBS 0.007596f
C1817 B.n867 VSUBS 0.007596f
C1818 B.n868 VSUBS 0.007596f
C1819 B.n869 VSUBS 0.007596f
C1820 B.n870 VSUBS 0.007596f
C1821 B.n871 VSUBS 0.007596f
C1822 B.n872 VSUBS 0.007596f
C1823 B.n873 VSUBS 0.007596f
C1824 B.n874 VSUBS 0.007596f
C1825 B.n875 VSUBS 0.007596f
C1826 B.n876 VSUBS 0.007596f
C1827 B.n877 VSUBS 0.007596f
C1828 B.n878 VSUBS 0.007596f
C1829 B.n879 VSUBS 0.007596f
C1830 B.n880 VSUBS 0.007596f
C1831 B.n881 VSUBS 0.007596f
C1832 B.n882 VSUBS 0.007596f
C1833 B.n883 VSUBS 0.007596f
C1834 B.n884 VSUBS 0.007596f
C1835 B.n885 VSUBS 0.007596f
C1836 B.n886 VSUBS 0.007596f
C1837 B.n887 VSUBS 0.007596f
C1838 B.n888 VSUBS 0.007596f
C1839 B.n889 VSUBS 0.007596f
C1840 B.n890 VSUBS 0.007596f
C1841 B.n891 VSUBS 0.007596f
C1842 B.n892 VSUBS 0.007596f
C1843 B.n893 VSUBS 0.007596f
C1844 B.n894 VSUBS 0.007596f
C1845 B.n895 VSUBS 0.007596f
C1846 B.n896 VSUBS 0.007596f
C1847 B.n897 VSUBS 0.007596f
C1848 B.n898 VSUBS 0.007596f
C1849 B.n899 VSUBS 0.007596f
C1850 B.n900 VSUBS 0.007596f
C1851 B.n901 VSUBS 0.007596f
C1852 B.n902 VSUBS 0.007596f
C1853 B.n903 VSUBS 0.017199f
.ends

