* NGSPICE file created from diff_pair_sample_0872.ext - technology: sky130A

.subckt diff_pair_sample_0872 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VP.t0 VDD1.t0 B.t8 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X1 VDD1.t8 VP.t1 VTAIL.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=2.6754 pd=14.5 as=1.1319 ps=7.19 w=6.86 l=3.74
X2 B.t22 B.t20 B.t21 B.t17 sky130_fd_pr__nfet_01v8 ad=2.6754 pd=14.5 as=0 ps=0 w=6.86 l=3.74
X3 VTAIL.t16 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X4 VDD1.t6 VP.t3 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=2.6754 ps=14.5 w=6.86 l=3.74
X5 VDD2.t9 VN.t0 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.6754 pd=14.5 as=1.1319 ps=7.19 w=6.86 l=3.74
X6 VDD2.t8 VN.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X7 VTAIL.t14 VP.t4 VDD1.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X8 VDD1.t5 VP.t5 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=2.6754 ps=14.5 w=6.86 l=3.74
X9 VTAIL.t12 VP.t6 VDD1.t3 B.t23 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X10 VTAIL.t4 VN.t2 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X11 VDD2.t6 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=2.6754 ps=14.5 w=6.86 l=3.74
X12 VDD2.t5 VN.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=2.6754 ps=14.5 w=6.86 l=3.74
X13 VTAIL.t8 VN.t5 VDD2.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X14 VTAIL.t2 VN.t6 VDD2.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X15 VDD1.t2 VP.t7 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X16 B.t19 B.t16 B.t18 B.t17 sky130_fd_pr__nfet_01v8 ad=2.6754 pd=14.5 as=0 ps=0 w=6.86 l=3.74
X17 VDD2.t2 VN.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X18 VDD2.t1 VN.t8 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6754 pd=14.5 as=1.1319 ps=7.19 w=6.86 l=3.74
X19 VDD1.t7 VP.t8 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6754 pd=14.5 as=1.1319 ps=7.19 w=6.86 l=3.74
X20 VDD1.t9 VP.t9 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X21 VTAIL.t19 VN.t9 VDD2.t0 B.t23 sky130_fd_pr__nfet_01v8 ad=1.1319 pd=7.19 as=1.1319 ps=7.19 w=6.86 l=3.74
X22 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.6754 pd=14.5 as=0 ps=0 w=6.86 l=3.74
X23 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.6754 pd=14.5 as=0 ps=0 w=6.86 l=3.74
R0 VP.n33 VP.n32 161.3
R1 VP.n34 VP.n29 161.3
R2 VP.n36 VP.n35 161.3
R3 VP.n37 VP.n28 161.3
R4 VP.n39 VP.n38 161.3
R5 VP.n40 VP.n27 161.3
R6 VP.n42 VP.n41 161.3
R7 VP.n43 VP.n26 161.3
R8 VP.n45 VP.n44 161.3
R9 VP.n46 VP.n25 161.3
R10 VP.n48 VP.n47 161.3
R11 VP.n49 VP.n24 161.3
R12 VP.n51 VP.n50 161.3
R13 VP.n52 VP.n23 161.3
R14 VP.n54 VP.n53 161.3
R15 VP.n55 VP.n22 161.3
R16 VP.n58 VP.n57 161.3
R17 VP.n59 VP.n21 161.3
R18 VP.n61 VP.n60 161.3
R19 VP.n62 VP.n20 161.3
R20 VP.n64 VP.n63 161.3
R21 VP.n65 VP.n19 161.3
R22 VP.n67 VP.n66 161.3
R23 VP.n68 VP.n18 161.3
R24 VP.n70 VP.n69 161.3
R25 VP.n125 VP.n124 161.3
R26 VP.n123 VP.n1 161.3
R27 VP.n122 VP.n121 161.3
R28 VP.n120 VP.n2 161.3
R29 VP.n119 VP.n118 161.3
R30 VP.n117 VP.n3 161.3
R31 VP.n116 VP.n115 161.3
R32 VP.n114 VP.n4 161.3
R33 VP.n113 VP.n112 161.3
R34 VP.n110 VP.n5 161.3
R35 VP.n109 VP.n108 161.3
R36 VP.n107 VP.n6 161.3
R37 VP.n106 VP.n105 161.3
R38 VP.n104 VP.n7 161.3
R39 VP.n103 VP.n102 161.3
R40 VP.n101 VP.n8 161.3
R41 VP.n100 VP.n99 161.3
R42 VP.n98 VP.n9 161.3
R43 VP.n97 VP.n96 161.3
R44 VP.n95 VP.n10 161.3
R45 VP.n94 VP.n93 161.3
R46 VP.n92 VP.n11 161.3
R47 VP.n91 VP.n90 161.3
R48 VP.n89 VP.n12 161.3
R49 VP.n88 VP.n87 161.3
R50 VP.n85 VP.n13 161.3
R51 VP.n84 VP.n83 161.3
R52 VP.n82 VP.n14 161.3
R53 VP.n81 VP.n80 161.3
R54 VP.n79 VP.n15 161.3
R55 VP.n78 VP.n77 161.3
R56 VP.n76 VP.n16 161.3
R57 VP.n75 VP.n74 161.3
R58 VP.n73 VP.n72 83.3598
R59 VP.n126 VP.n0 83.3598
R60 VP.n71 VP.n17 83.3598
R61 VP.n30 VP.t8 77.0929
R62 VP.n31 VP.n30 71.5921
R63 VP.n72 VP.n71 55.5185
R64 VP.n80 VP.n79 50.7491
R65 VP.n118 VP.n2 50.7491
R66 VP.n63 VP.n19 50.7491
R67 VP.n99 VP.t7 44.2053
R68 VP.n73 VP.t1 44.2053
R69 VP.n86 VP.t4 44.2053
R70 VP.n111 VP.t2 44.2053
R71 VP.n0 VP.t5 44.2053
R72 VP.n44 VP.t9 44.2053
R73 VP.n17 VP.t3 44.2053
R74 VP.n56 VP.t6 44.2053
R75 VP.n31 VP.t0 44.2053
R76 VP.n93 VP.n92 43.9677
R77 VP.n105 VP.n6 43.9677
R78 VP.n50 VP.n23 43.9677
R79 VP.n38 VP.n37 43.9677
R80 VP.n93 VP.n10 37.1863
R81 VP.n105 VP.n104 37.1863
R82 VP.n50 VP.n49 37.1863
R83 VP.n38 VP.n27 37.1863
R84 VP.n80 VP.n14 30.405
R85 VP.n118 VP.n117 30.405
R86 VP.n63 VP.n62 30.405
R87 VP.n74 VP.n16 24.5923
R88 VP.n78 VP.n16 24.5923
R89 VP.n79 VP.n78 24.5923
R90 VP.n84 VP.n14 24.5923
R91 VP.n85 VP.n84 24.5923
R92 VP.n87 VP.n12 24.5923
R93 VP.n91 VP.n12 24.5923
R94 VP.n92 VP.n91 24.5923
R95 VP.n97 VP.n10 24.5923
R96 VP.n98 VP.n97 24.5923
R97 VP.n99 VP.n98 24.5923
R98 VP.n99 VP.n8 24.5923
R99 VP.n103 VP.n8 24.5923
R100 VP.n104 VP.n103 24.5923
R101 VP.n109 VP.n6 24.5923
R102 VP.n110 VP.n109 24.5923
R103 VP.n112 VP.n110 24.5923
R104 VP.n116 VP.n4 24.5923
R105 VP.n117 VP.n116 24.5923
R106 VP.n122 VP.n2 24.5923
R107 VP.n123 VP.n122 24.5923
R108 VP.n124 VP.n123 24.5923
R109 VP.n67 VP.n19 24.5923
R110 VP.n68 VP.n67 24.5923
R111 VP.n69 VP.n68 24.5923
R112 VP.n54 VP.n23 24.5923
R113 VP.n55 VP.n54 24.5923
R114 VP.n57 VP.n55 24.5923
R115 VP.n61 VP.n21 24.5923
R116 VP.n62 VP.n61 24.5923
R117 VP.n42 VP.n27 24.5923
R118 VP.n43 VP.n42 24.5923
R119 VP.n44 VP.n43 24.5923
R120 VP.n44 VP.n25 24.5923
R121 VP.n48 VP.n25 24.5923
R122 VP.n49 VP.n48 24.5923
R123 VP.n32 VP.n29 24.5923
R124 VP.n36 VP.n29 24.5923
R125 VP.n37 VP.n36 24.5923
R126 VP.n86 VP.n85 21.1495
R127 VP.n111 VP.n4 21.1495
R128 VP.n56 VP.n21 21.1495
R129 VP.n74 VP.n73 6.88621
R130 VP.n124 VP.n0 6.88621
R131 VP.n69 VP.n17 6.88621
R132 VP.n87 VP.n86 3.44336
R133 VP.n112 VP.n111 3.44336
R134 VP.n57 VP.n56 3.44336
R135 VP.n32 VP.n31 3.44336
R136 VP.n33 VP.n30 3.23942
R137 VP.n71 VP.n70 0.354861
R138 VP.n75 VP.n72 0.354861
R139 VP.n126 VP.n125 0.354861
R140 VP VP.n126 0.267071
R141 VP.n34 VP.n33 0.189894
R142 VP.n35 VP.n34 0.189894
R143 VP.n35 VP.n28 0.189894
R144 VP.n39 VP.n28 0.189894
R145 VP.n40 VP.n39 0.189894
R146 VP.n41 VP.n40 0.189894
R147 VP.n41 VP.n26 0.189894
R148 VP.n45 VP.n26 0.189894
R149 VP.n46 VP.n45 0.189894
R150 VP.n47 VP.n46 0.189894
R151 VP.n47 VP.n24 0.189894
R152 VP.n51 VP.n24 0.189894
R153 VP.n52 VP.n51 0.189894
R154 VP.n53 VP.n52 0.189894
R155 VP.n53 VP.n22 0.189894
R156 VP.n58 VP.n22 0.189894
R157 VP.n59 VP.n58 0.189894
R158 VP.n60 VP.n59 0.189894
R159 VP.n60 VP.n20 0.189894
R160 VP.n64 VP.n20 0.189894
R161 VP.n65 VP.n64 0.189894
R162 VP.n66 VP.n65 0.189894
R163 VP.n66 VP.n18 0.189894
R164 VP.n70 VP.n18 0.189894
R165 VP.n76 VP.n75 0.189894
R166 VP.n77 VP.n76 0.189894
R167 VP.n77 VP.n15 0.189894
R168 VP.n81 VP.n15 0.189894
R169 VP.n82 VP.n81 0.189894
R170 VP.n83 VP.n82 0.189894
R171 VP.n83 VP.n13 0.189894
R172 VP.n88 VP.n13 0.189894
R173 VP.n89 VP.n88 0.189894
R174 VP.n90 VP.n89 0.189894
R175 VP.n90 VP.n11 0.189894
R176 VP.n94 VP.n11 0.189894
R177 VP.n95 VP.n94 0.189894
R178 VP.n96 VP.n95 0.189894
R179 VP.n96 VP.n9 0.189894
R180 VP.n100 VP.n9 0.189894
R181 VP.n101 VP.n100 0.189894
R182 VP.n102 VP.n101 0.189894
R183 VP.n102 VP.n7 0.189894
R184 VP.n106 VP.n7 0.189894
R185 VP.n107 VP.n106 0.189894
R186 VP.n108 VP.n107 0.189894
R187 VP.n108 VP.n5 0.189894
R188 VP.n113 VP.n5 0.189894
R189 VP.n114 VP.n113 0.189894
R190 VP.n115 VP.n114 0.189894
R191 VP.n115 VP.n3 0.189894
R192 VP.n119 VP.n3 0.189894
R193 VP.n120 VP.n119 0.189894
R194 VP.n121 VP.n120 0.189894
R195 VP.n121 VP.n1 0.189894
R196 VP.n125 VP.n1 0.189894
R197 VDD1.n1 VDD1.t7 74.13
R198 VDD1.n3 VDD1.t8 74.1299
R199 VDD1.n5 VDD1.n4 70.3101
R200 VDD1.n1 VDD1.n0 67.7351
R201 VDD1.n7 VDD1.n6 67.735
R202 VDD1.n3 VDD1.n2 67.734
R203 VDD1.n7 VDD1.n5 48.6324
R204 VDD1.n6 VDD1.t3 2.8868
R205 VDD1.n6 VDD1.t6 2.8868
R206 VDD1.n0 VDD1.t0 2.8868
R207 VDD1.n0 VDD1.t9 2.8868
R208 VDD1.n4 VDD1.t1 2.8868
R209 VDD1.n4 VDD1.t5 2.8868
R210 VDD1.n2 VDD1.t4 2.8868
R211 VDD1.n2 VDD1.t2 2.8868
R212 VDD1 VDD1.n7 2.57378
R213 VDD1 VDD1.n1 0.935845
R214 VDD1.n5 VDD1.n3 0.822309
R215 VTAIL.n11 VTAIL.t0 53.9426
R216 VTAIL.n17 VTAIL.t3 53.9425
R217 VTAIL.n2 VTAIL.t13 53.9425
R218 VTAIL.n16 VTAIL.t15 53.9425
R219 VTAIL.n15 VTAIL.n14 51.0563
R220 VTAIL.n13 VTAIL.n12 51.0563
R221 VTAIL.n10 VTAIL.n9 51.0563
R222 VTAIL.n8 VTAIL.n7 51.0563
R223 VTAIL.n19 VTAIL.n18 51.0552
R224 VTAIL.n1 VTAIL.n0 51.0552
R225 VTAIL.n4 VTAIL.n3 51.0552
R226 VTAIL.n6 VTAIL.n5 51.0552
R227 VTAIL.n8 VTAIL.n6 25.2979
R228 VTAIL.n17 VTAIL.n16 21.7893
R229 VTAIL.n10 VTAIL.n8 3.50912
R230 VTAIL.n11 VTAIL.n10 3.50912
R231 VTAIL.n15 VTAIL.n13 3.50912
R232 VTAIL.n16 VTAIL.n15 3.50912
R233 VTAIL.n6 VTAIL.n4 3.50912
R234 VTAIL.n4 VTAIL.n2 3.50912
R235 VTAIL.n19 VTAIL.n17 3.50912
R236 VTAIL.n18 VTAIL.t5 2.8868
R237 VTAIL.n18 VTAIL.t19 2.8868
R238 VTAIL.n0 VTAIL.t1 2.8868
R239 VTAIL.n0 VTAIL.t8 2.8868
R240 VTAIL.n3 VTAIL.t11 2.8868
R241 VTAIL.n3 VTAIL.t16 2.8868
R242 VTAIL.n5 VTAIL.t17 2.8868
R243 VTAIL.n5 VTAIL.t14 2.8868
R244 VTAIL.n14 VTAIL.t9 2.8868
R245 VTAIL.n14 VTAIL.t12 2.8868
R246 VTAIL.n12 VTAIL.t10 2.8868
R247 VTAIL.n12 VTAIL.t18 2.8868
R248 VTAIL.n9 VTAIL.t7 2.8868
R249 VTAIL.n9 VTAIL.t2 2.8868
R250 VTAIL.n7 VTAIL.t6 2.8868
R251 VTAIL.n7 VTAIL.t4 2.8868
R252 VTAIL VTAIL.n1 2.69016
R253 VTAIL.n13 VTAIL.n11 2.22464
R254 VTAIL.n2 VTAIL.n1 2.22464
R255 VTAIL VTAIL.n19 0.819465
R256 B.n968 B.n967 585
R257 B.n969 B.n968 585
R258 B.n304 B.n177 585
R259 B.n303 B.n302 585
R260 B.n301 B.n300 585
R261 B.n299 B.n298 585
R262 B.n297 B.n296 585
R263 B.n295 B.n294 585
R264 B.n293 B.n292 585
R265 B.n291 B.n290 585
R266 B.n289 B.n288 585
R267 B.n287 B.n286 585
R268 B.n285 B.n284 585
R269 B.n283 B.n282 585
R270 B.n281 B.n280 585
R271 B.n279 B.n278 585
R272 B.n277 B.n276 585
R273 B.n275 B.n274 585
R274 B.n273 B.n272 585
R275 B.n271 B.n270 585
R276 B.n269 B.n268 585
R277 B.n267 B.n266 585
R278 B.n265 B.n264 585
R279 B.n263 B.n262 585
R280 B.n261 B.n260 585
R281 B.n259 B.n258 585
R282 B.n257 B.n256 585
R283 B.n255 B.n254 585
R284 B.n253 B.n252 585
R285 B.n251 B.n250 585
R286 B.n249 B.n248 585
R287 B.n247 B.n246 585
R288 B.n245 B.n244 585
R289 B.n243 B.n242 585
R290 B.n241 B.n240 585
R291 B.n239 B.n238 585
R292 B.n237 B.n236 585
R293 B.n234 B.n233 585
R294 B.n232 B.n231 585
R295 B.n230 B.n229 585
R296 B.n228 B.n227 585
R297 B.n226 B.n225 585
R298 B.n224 B.n223 585
R299 B.n222 B.n221 585
R300 B.n220 B.n219 585
R301 B.n218 B.n217 585
R302 B.n216 B.n215 585
R303 B.n214 B.n213 585
R304 B.n212 B.n211 585
R305 B.n210 B.n209 585
R306 B.n208 B.n207 585
R307 B.n206 B.n205 585
R308 B.n204 B.n203 585
R309 B.n202 B.n201 585
R310 B.n200 B.n199 585
R311 B.n198 B.n197 585
R312 B.n196 B.n195 585
R313 B.n194 B.n193 585
R314 B.n192 B.n191 585
R315 B.n190 B.n189 585
R316 B.n188 B.n187 585
R317 B.n186 B.n185 585
R318 B.n184 B.n183 585
R319 B.n144 B.n143 585
R320 B.n966 B.n145 585
R321 B.n970 B.n145 585
R322 B.n965 B.n964 585
R323 B.n964 B.n141 585
R324 B.n963 B.n140 585
R325 B.n976 B.n140 585
R326 B.n962 B.n139 585
R327 B.n977 B.n139 585
R328 B.n961 B.n138 585
R329 B.n978 B.n138 585
R330 B.n960 B.n959 585
R331 B.n959 B.n134 585
R332 B.n958 B.n133 585
R333 B.n984 B.n133 585
R334 B.n957 B.n132 585
R335 B.n985 B.n132 585
R336 B.n956 B.n131 585
R337 B.n986 B.n131 585
R338 B.n955 B.n954 585
R339 B.n954 B.n130 585
R340 B.n953 B.n126 585
R341 B.n992 B.n126 585
R342 B.n952 B.n125 585
R343 B.n993 B.n125 585
R344 B.n951 B.n124 585
R345 B.n994 B.n124 585
R346 B.n950 B.n949 585
R347 B.n949 B.n120 585
R348 B.n948 B.n119 585
R349 B.n1000 B.n119 585
R350 B.n947 B.n118 585
R351 B.n1001 B.n118 585
R352 B.n946 B.n117 585
R353 B.n1002 B.n117 585
R354 B.n945 B.n944 585
R355 B.n944 B.n113 585
R356 B.n943 B.n112 585
R357 B.n1008 B.n112 585
R358 B.n942 B.n111 585
R359 B.n1009 B.n111 585
R360 B.n941 B.n110 585
R361 B.n1010 B.n110 585
R362 B.n940 B.n939 585
R363 B.n939 B.n106 585
R364 B.n938 B.n105 585
R365 B.n1016 B.n105 585
R366 B.n937 B.n104 585
R367 B.n1017 B.n104 585
R368 B.n936 B.n103 585
R369 B.n1018 B.n103 585
R370 B.n935 B.n934 585
R371 B.n934 B.n99 585
R372 B.n933 B.n98 585
R373 B.n1024 B.n98 585
R374 B.n932 B.n97 585
R375 B.n1025 B.n97 585
R376 B.n931 B.n96 585
R377 B.n1026 B.n96 585
R378 B.n930 B.n929 585
R379 B.n929 B.n92 585
R380 B.n928 B.n91 585
R381 B.n1032 B.n91 585
R382 B.n927 B.n90 585
R383 B.n1033 B.n90 585
R384 B.n926 B.n89 585
R385 B.n1034 B.n89 585
R386 B.n925 B.n924 585
R387 B.n924 B.n85 585
R388 B.n923 B.n84 585
R389 B.n1040 B.n84 585
R390 B.n922 B.n83 585
R391 B.n1041 B.n83 585
R392 B.n921 B.n82 585
R393 B.n1042 B.n82 585
R394 B.n920 B.n919 585
R395 B.n919 B.n78 585
R396 B.n918 B.n77 585
R397 B.n1048 B.n77 585
R398 B.n917 B.n76 585
R399 B.n1049 B.n76 585
R400 B.n916 B.n75 585
R401 B.n1050 B.n75 585
R402 B.n915 B.n914 585
R403 B.n914 B.n71 585
R404 B.n913 B.n70 585
R405 B.n1056 B.n70 585
R406 B.n912 B.n69 585
R407 B.n1057 B.n69 585
R408 B.n911 B.n68 585
R409 B.n1058 B.n68 585
R410 B.n910 B.n909 585
R411 B.n909 B.n64 585
R412 B.n908 B.n63 585
R413 B.n1064 B.n63 585
R414 B.n907 B.n62 585
R415 B.n1065 B.n62 585
R416 B.n906 B.n61 585
R417 B.n1066 B.n61 585
R418 B.n905 B.n904 585
R419 B.n904 B.n57 585
R420 B.n903 B.n56 585
R421 B.n1072 B.n56 585
R422 B.n902 B.n55 585
R423 B.n1073 B.n55 585
R424 B.n901 B.n54 585
R425 B.n1074 B.n54 585
R426 B.n900 B.n899 585
R427 B.n899 B.n50 585
R428 B.n898 B.n49 585
R429 B.n1080 B.n49 585
R430 B.n897 B.n48 585
R431 B.n1081 B.n48 585
R432 B.n896 B.n47 585
R433 B.n1082 B.n47 585
R434 B.n895 B.n894 585
R435 B.n894 B.n43 585
R436 B.n893 B.n42 585
R437 B.n1088 B.n42 585
R438 B.n892 B.n41 585
R439 B.n1089 B.n41 585
R440 B.n891 B.n40 585
R441 B.n1090 B.n40 585
R442 B.n890 B.n889 585
R443 B.n889 B.n36 585
R444 B.n888 B.n35 585
R445 B.n1096 B.n35 585
R446 B.n887 B.n34 585
R447 B.n1097 B.n34 585
R448 B.n886 B.n33 585
R449 B.n1098 B.n33 585
R450 B.n885 B.n884 585
R451 B.n884 B.n29 585
R452 B.n883 B.n28 585
R453 B.n1104 B.n28 585
R454 B.n882 B.n27 585
R455 B.n1105 B.n27 585
R456 B.n881 B.n26 585
R457 B.n1106 B.n26 585
R458 B.n880 B.n879 585
R459 B.n879 B.n22 585
R460 B.n878 B.n21 585
R461 B.n1112 B.n21 585
R462 B.n877 B.n20 585
R463 B.n1113 B.n20 585
R464 B.n876 B.n19 585
R465 B.n1114 B.n19 585
R466 B.n875 B.n874 585
R467 B.n874 B.n15 585
R468 B.n873 B.n14 585
R469 B.n1120 B.n14 585
R470 B.n872 B.n13 585
R471 B.n1121 B.n13 585
R472 B.n871 B.n12 585
R473 B.n1122 B.n12 585
R474 B.n870 B.n869 585
R475 B.n869 B.n8 585
R476 B.n868 B.n7 585
R477 B.n1128 B.n7 585
R478 B.n867 B.n6 585
R479 B.n1129 B.n6 585
R480 B.n866 B.n5 585
R481 B.n1130 B.n5 585
R482 B.n865 B.n864 585
R483 B.n864 B.n4 585
R484 B.n863 B.n305 585
R485 B.n863 B.n862 585
R486 B.n853 B.n306 585
R487 B.n307 B.n306 585
R488 B.n855 B.n854 585
R489 B.n856 B.n855 585
R490 B.n852 B.n312 585
R491 B.n312 B.n311 585
R492 B.n851 B.n850 585
R493 B.n850 B.n849 585
R494 B.n314 B.n313 585
R495 B.n315 B.n314 585
R496 B.n842 B.n841 585
R497 B.n843 B.n842 585
R498 B.n840 B.n320 585
R499 B.n320 B.n319 585
R500 B.n839 B.n838 585
R501 B.n838 B.n837 585
R502 B.n322 B.n321 585
R503 B.n323 B.n322 585
R504 B.n830 B.n829 585
R505 B.n831 B.n830 585
R506 B.n828 B.n328 585
R507 B.n328 B.n327 585
R508 B.n827 B.n826 585
R509 B.n826 B.n825 585
R510 B.n330 B.n329 585
R511 B.n331 B.n330 585
R512 B.n818 B.n817 585
R513 B.n819 B.n818 585
R514 B.n816 B.n336 585
R515 B.n336 B.n335 585
R516 B.n815 B.n814 585
R517 B.n814 B.n813 585
R518 B.n338 B.n337 585
R519 B.n339 B.n338 585
R520 B.n806 B.n805 585
R521 B.n807 B.n806 585
R522 B.n804 B.n344 585
R523 B.n344 B.n343 585
R524 B.n803 B.n802 585
R525 B.n802 B.n801 585
R526 B.n346 B.n345 585
R527 B.n347 B.n346 585
R528 B.n794 B.n793 585
R529 B.n795 B.n794 585
R530 B.n792 B.n352 585
R531 B.n352 B.n351 585
R532 B.n791 B.n790 585
R533 B.n790 B.n789 585
R534 B.n354 B.n353 585
R535 B.n355 B.n354 585
R536 B.n782 B.n781 585
R537 B.n783 B.n782 585
R538 B.n780 B.n360 585
R539 B.n360 B.n359 585
R540 B.n779 B.n778 585
R541 B.n778 B.n777 585
R542 B.n362 B.n361 585
R543 B.n363 B.n362 585
R544 B.n770 B.n769 585
R545 B.n771 B.n770 585
R546 B.n768 B.n368 585
R547 B.n368 B.n367 585
R548 B.n767 B.n766 585
R549 B.n766 B.n765 585
R550 B.n370 B.n369 585
R551 B.n371 B.n370 585
R552 B.n758 B.n757 585
R553 B.n759 B.n758 585
R554 B.n756 B.n376 585
R555 B.n376 B.n375 585
R556 B.n755 B.n754 585
R557 B.n754 B.n753 585
R558 B.n378 B.n377 585
R559 B.n379 B.n378 585
R560 B.n746 B.n745 585
R561 B.n747 B.n746 585
R562 B.n744 B.n384 585
R563 B.n384 B.n383 585
R564 B.n743 B.n742 585
R565 B.n742 B.n741 585
R566 B.n386 B.n385 585
R567 B.n387 B.n386 585
R568 B.n734 B.n733 585
R569 B.n735 B.n734 585
R570 B.n732 B.n392 585
R571 B.n392 B.n391 585
R572 B.n731 B.n730 585
R573 B.n730 B.n729 585
R574 B.n394 B.n393 585
R575 B.n395 B.n394 585
R576 B.n722 B.n721 585
R577 B.n723 B.n722 585
R578 B.n720 B.n400 585
R579 B.n400 B.n399 585
R580 B.n719 B.n718 585
R581 B.n718 B.n717 585
R582 B.n402 B.n401 585
R583 B.n403 B.n402 585
R584 B.n710 B.n709 585
R585 B.n711 B.n710 585
R586 B.n708 B.n408 585
R587 B.n408 B.n407 585
R588 B.n707 B.n706 585
R589 B.n706 B.n705 585
R590 B.n410 B.n409 585
R591 B.n411 B.n410 585
R592 B.n698 B.n697 585
R593 B.n699 B.n698 585
R594 B.n696 B.n416 585
R595 B.n416 B.n415 585
R596 B.n695 B.n694 585
R597 B.n694 B.n693 585
R598 B.n418 B.n417 585
R599 B.n419 B.n418 585
R600 B.n686 B.n685 585
R601 B.n687 B.n686 585
R602 B.n684 B.n424 585
R603 B.n424 B.n423 585
R604 B.n683 B.n682 585
R605 B.n682 B.n681 585
R606 B.n426 B.n425 585
R607 B.n427 B.n426 585
R608 B.n674 B.n673 585
R609 B.n675 B.n674 585
R610 B.n672 B.n432 585
R611 B.n432 B.n431 585
R612 B.n671 B.n670 585
R613 B.n670 B.n669 585
R614 B.n434 B.n433 585
R615 B.n435 B.n434 585
R616 B.n662 B.n661 585
R617 B.n663 B.n662 585
R618 B.n660 B.n440 585
R619 B.n440 B.n439 585
R620 B.n659 B.n658 585
R621 B.n658 B.n657 585
R622 B.n442 B.n441 585
R623 B.n650 B.n442 585
R624 B.n649 B.n648 585
R625 B.n651 B.n649 585
R626 B.n647 B.n447 585
R627 B.n447 B.n446 585
R628 B.n646 B.n645 585
R629 B.n645 B.n644 585
R630 B.n449 B.n448 585
R631 B.n450 B.n449 585
R632 B.n637 B.n636 585
R633 B.n638 B.n637 585
R634 B.n635 B.n455 585
R635 B.n455 B.n454 585
R636 B.n634 B.n633 585
R637 B.n633 B.n632 585
R638 B.n457 B.n456 585
R639 B.n458 B.n457 585
R640 B.n625 B.n624 585
R641 B.n626 B.n625 585
R642 B.n461 B.n460 585
R643 B.n498 B.n497 585
R644 B.n499 B.n495 585
R645 B.n495 B.n462 585
R646 B.n501 B.n500 585
R647 B.n503 B.n494 585
R648 B.n506 B.n505 585
R649 B.n507 B.n493 585
R650 B.n509 B.n508 585
R651 B.n511 B.n492 585
R652 B.n514 B.n513 585
R653 B.n515 B.n491 585
R654 B.n517 B.n516 585
R655 B.n519 B.n490 585
R656 B.n522 B.n521 585
R657 B.n523 B.n489 585
R658 B.n525 B.n524 585
R659 B.n527 B.n488 585
R660 B.n530 B.n529 585
R661 B.n531 B.n487 585
R662 B.n533 B.n532 585
R663 B.n535 B.n486 585
R664 B.n538 B.n537 585
R665 B.n539 B.n485 585
R666 B.n541 B.n540 585
R667 B.n543 B.n484 585
R668 B.n546 B.n545 585
R669 B.n547 B.n481 585
R670 B.n550 B.n549 585
R671 B.n552 B.n480 585
R672 B.n555 B.n554 585
R673 B.n556 B.n479 585
R674 B.n558 B.n557 585
R675 B.n560 B.n478 585
R676 B.n563 B.n562 585
R677 B.n564 B.n477 585
R678 B.n569 B.n568 585
R679 B.n571 B.n476 585
R680 B.n574 B.n573 585
R681 B.n575 B.n475 585
R682 B.n577 B.n576 585
R683 B.n579 B.n474 585
R684 B.n582 B.n581 585
R685 B.n583 B.n473 585
R686 B.n585 B.n584 585
R687 B.n587 B.n472 585
R688 B.n590 B.n589 585
R689 B.n591 B.n471 585
R690 B.n593 B.n592 585
R691 B.n595 B.n470 585
R692 B.n598 B.n597 585
R693 B.n599 B.n469 585
R694 B.n601 B.n600 585
R695 B.n603 B.n468 585
R696 B.n606 B.n605 585
R697 B.n607 B.n467 585
R698 B.n609 B.n608 585
R699 B.n611 B.n466 585
R700 B.n614 B.n613 585
R701 B.n615 B.n465 585
R702 B.n617 B.n616 585
R703 B.n619 B.n464 585
R704 B.n622 B.n621 585
R705 B.n623 B.n463 585
R706 B.n628 B.n627 585
R707 B.n627 B.n626 585
R708 B.n629 B.n459 585
R709 B.n459 B.n458 585
R710 B.n631 B.n630 585
R711 B.n632 B.n631 585
R712 B.n453 B.n452 585
R713 B.n454 B.n453 585
R714 B.n640 B.n639 585
R715 B.n639 B.n638 585
R716 B.n641 B.n451 585
R717 B.n451 B.n450 585
R718 B.n643 B.n642 585
R719 B.n644 B.n643 585
R720 B.n445 B.n444 585
R721 B.n446 B.n445 585
R722 B.n653 B.n652 585
R723 B.n652 B.n651 585
R724 B.n654 B.n443 585
R725 B.n650 B.n443 585
R726 B.n656 B.n655 585
R727 B.n657 B.n656 585
R728 B.n438 B.n437 585
R729 B.n439 B.n438 585
R730 B.n665 B.n664 585
R731 B.n664 B.n663 585
R732 B.n666 B.n436 585
R733 B.n436 B.n435 585
R734 B.n668 B.n667 585
R735 B.n669 B.n668 585
R736 B.n430 B.n429 585
R737 B.n431 B.n430 585
R738 B.n677 B.n676 585
R739 B.n676 B.n675 585
R740 B.n678 B.n428 585
R741 B.n428 B.n427 585
R742 B.n680 B.n679 585
R743 B.n681 B.n680 585
R744 B.n422 B.n421 585
R745 B.n423 B.n422 585
R746 B.n689 B.n688 585
R747 B.n688 B.n687 585
R748 B.n690 B.n420 585
R749 B.n420 B.n419 585
R750 B.n692 B.n691 585
R751 B.n693 B.n692 585
R752 B.n414 B.n413 585
R753 B.n415 B.n414 585
R754 B.n701 B.n700 585
R755 B.n700 B.n699 585
R756 B.n702 B.n412 585
R757 B.n412 B.n411 585
R758 B.n704 B.n703 585
R759 B.n705 B.n704 585
R760 B.n406 B.n405 585
R761 B.n407 B.n406 585
R762 B.n713 B.n712 585
R763 B.n712 B.n711 585
R764 B.n714 B.n404 585
R765 B.n404 B.n403 585
R766 B.n716 B.n715 585
R767 B.n717 B.n716 585
R768 B.n398 B.n397 585
R769 B.n399 B.n398 585
R770 B.n725 B.n724 585
R771 B.n724 B.n723 585
R772 B.n726 B.n396 585
R773 B.n396 B.n395 585
R774 B.n728 B.n727 585
R775 B.n729 B.n728 585
R776 B.n390 B.n389 585
R777 B.n391 B.n390 585
R778 B.n737 B.n736 585
R779 B.n736 B.n735 585
R780 B.n738 B.n388 585
R781 B.n388 B.n387 585
R782 B.n740 B.n739 585
R783 B.n741 B.n740 585
R784 B.n382 B.n381 585
R785 B.n383 B.n382 585
R786 B.n749 B.n748 585
R787 B.n748 B.n747 585
R788 B.n750 B.n380 585
R789 B.n380 B.n379 585
R790 B.n752 B.n751 585
R791 B.n753 B.n752 585
R792 B.n374 B.n373 585
R793 B.n375 B.n374 585
R794 B.n761 B.n760 585
R795 B.n760 B.n759 585
R796 B.n762 B.n372 585
R797 B.n372 B.n371 585
R798 B.n764 B.n763 585
R799 B.n765 B.n764 585
R800 B.n366 B.n365 585
R801 B.n367 B.n366 585
R802 B.n773 B.n772 585
R803 B.n772 B.n771 585
R804 B.n774 B.n364 585
R805 B.n364 B.n363 585
R806 B.n776 B.n775 585
R807 B.n777 B.n776 585
R808 B.n358 B.n357 585
R809 B.n359 B.n358 585
R810 B.n785 B.n784 585
R811 B.n784 B.n783 585
R812 B.n786 B.n356 585
R813 B.n356 B.n355 585
R814 B.n788 B.n787 585
R815 B.n789 B.n788 585
R816 B.n350 B.n349 585
R817 B.n351 B.n350 585
R818 B.n797 B.n796 585
R819 B.n796 B.n795 585
R820 B.n798 B.n348 585
R821 B.n348 B.n347 585
R822 B.n800 B.n799 585
R823 B.n801 B.n800 585
R824 B.n342 B.n341 585
R825 B.n343 B.n342 585
R826 B.n809 B.n808 585
R827 B.n808 B.n807 585
R828 B.n810 B.n340 585
R829 B.n340 B.n339 585
R830 B.n812 B.n811 585
R831 B.n813 B.n812 585
R832 B.n334 B.n333 585
R833 B.n335 B.n334 585
R834 B.n821 B.n820 585
R835 B.n820 B.n819 585
R836 B.n822 B.n332 585
R837 B.n332 B.n331 585
R838 B.n824 B.n823 585
R839 B.n825 B.n824 585
R840 B.n326 B.n325 585
R841 B.n327 B.n326 585
R842 B.n833 B.n832 585
R843 B.n832 B.n831 585
R844 B.n834 B.n324 585
R845 B.n324 B.n323 585
R846 B.n836 B.n835 585
R847 B.n837 B.n836 585
R848 B.n318 B.n317 585
R849 B.n319 B.n318 585
R850 B.n845 B.n844 585
R851 B.n844 B.n843 585
R852 B.n846 B.n316 585
R853 B.n316 B.n315 585
R854 B.n848 B.n847 585
R855 B.n849 B.n848 585
R856 B.n310 B.n309 585
R857 B.n311 B.n310 585
R858 B.n858 B.n857 585
R859 B.n857 B.n856 585
R860 B.n859 B.n308 585
R861 B.n308 B.n307 585
R862 B.n861 B.n860 585
R863 B.n862 B.n861 585
R864 B.n2 B.n0 585
R865 B.n4 B.n2 585
R866 B.n3 B.n1 585
R867 B.n1129 B.n3 585
R868 B.n1127 B.n1126 585
R869 B.n1128 B.n1127 585
R870 B.n1125 B.n9 585
R871 B.n9 B.n8 585
R872 B.n1124 B.n1123 585
R873 B.n1123 B.n1122 585
R874 B.n11 B.n10 585
R875 B.n1121 B.n11 585
R876 B.n1119 B.n1118 585
R877 B.n1120 B.n1119 585
R878 B.n1117 B.n16 585
R879 B.n16 B.n15 585
R880 B.n1116 B.n1115 585
R881 B.n1115 B.n1114 585
R882 B.n18 B.n17 585
R883 B.n1113 B.n18 585
R884 B.n1111 B.n1110 585
R885 B.n1112 B.n1111 585
R886 B.n1109 B.n23 585
R887 B.n23 B.n22 585
R888 B.n1108 B.n1107 585
R889 B.n1107 B.n1106 585
R890 B.n25 B.n24 585
R891 B.n1105 B.n25 585
R892 B.n1103 B.n1102 585
R893 B.n1104 B.n1103 585
R894 B.n1101 B.n30 585
R895 B.n30 B.n29 585
R896 B.n1100 B.n1099 585
R897 B.n1099 B.n1098 585
R898 B.n32 B.n31 585
R899 B.n1097 B.n32 585
R900 B.n1095 B.n1094 585
R901 B.n1096 B.n1095 585
R902 B.n1093 B.n37 585
R903 B.n37 B.n36 585
R904 B.n1092 B.n1091 585
R905 B.n1091 B.n1090 585
R906 B.n39 B.n38 585
R907 B.n1089 B.n39 585
R908 B.n1087 B.n1086 585
R909 B.n1088 B.n1087 585
R910 B.n1085 B.n44 585
R911 B.n44 B.n43 585
R912 B.n1084 B.n1083 585
R913 B.n1083 B.n1082 585
R914 B.n46 B.n45 585
R915 B.n1081 B.n46 585
R916 B.n1079 B.n1078 585
R917 B.n1080 B.n1079 585
R918 B.n1077 B.n51 585
R919 B.n51 B.n50 585
R920 B.n1076 B.n1075 585
R921 B.n1075 B.n1074 585
R922 B.n53 B.n52 585
R923 B.n1073 B.n53 585
R924 B.n1071 B.n1070 585
R925 B.n1072 B.n1071 585
R926 B.n1069 B.n58 585
R927 B.n58 B.n57 585
R928 B.n1068 B.n1067 585
R929 B.n1067 B.n1066 585
R930 B.n60 B.n59 585
R931 B.n1065 B.n60 585
R932 B.n1063 B.n1062 585
R933 B.n1064 B.n1063 585
R934 B.n1061 B.n65 585
R935 B.n65 B.n64 585
R936 B.n1060 B.n1059 585
R937 B.n1059 B.n1058 585
R938 B.n67 B.n66 585
R939 B.n1057 B.n67 585
R940 B.n1055 B.n1054 585
R941 B.n1056 B.n1055 585
R942 B.n1053 B.n72 585
R943 B.n72 B.n71 585
R944 B.n1052 B.n1051 585
R945 B.n1051 B.n1050 585
R946 B.n74 B.n73 585
R947 B.n1049 B.n74 585
R948 B.n1047 B.n1046 585
R949 B.n1048 B.n1047 585
R950 B.n1045 B.n79 585
R951 B.n79 B.n78 585
R952 B.n1044 B.n1043 585
R953 B.n1043 B.n1042 585
R954 B.n81 B.n80 585
R955 B.n1041 B.n81 585
R956 B.n1039 B.n1038 585
R957 B.n1040 B.n1039 585
R958 B.n1037 B.n86 585
R959 B.n86 B.n85 585
R960 B.n1036 B.n1035 585
R961 B.n1035 B.n1034 585
R962 B.n88 B.n87 585
R963 B.n1033 B.n88 585
R964 B.n1031 B.n1030 585
R965 B.n1032 B.n1031 585
R966 B.n1029 B.n93 585
R967 B.n93 B.n92 585
R968 B.n1028 B.n1027 585
R969 B.n1027 B.n1026 585
R970 B.n95 B.n94 585
R971 B.n1025 B.n95 585
R972 B.n1023 B.n1022 585
R973 B.n1024 B.n1023 585
R974 B.n1021 B.n100 585
R975 B.n100 B.n99 585
R976 B.n1020 B.n1019 585
R977 B.n1019 B.n1018 585
R978 B.n102 B.n101 585
R979 B.n1017 B.n102 585
R980 B.n1015 B.n1014 585
R981 B.n1016 B.n1015 585
R982 B.n1013 B.n107 585
R983 B.n107 B.n106 585
R984 B.n1012 B.n1011 585
R985 B.n1011 B.n1010 585
R986 B.n109 B.n108 585
R987 B.n1009 B.n109 585
R988 B.n1007 B.n1006 585
R989 B.n1008 B.n1007 585
R990 B.n1005 B.n114 585
R991 B.n114 B.n113 585
R992 B.n1004 B.n1003 585
R993 B.n1003 B.n1002 585
R994 B.n116 B.n115 585
R995 B.n1001 B.n116 585
R996 B.n999 B.n998 585
R997 B.n1000 B.n999 585
R998 B.n997 B.n121 585
R999 B.n121 B.n120 585
R1000 B.n996 B.n995 585
R1001 B.n995 B.n994 585
R1002 B.n123 B.n122 585
R1003 B.n993 B.n123 585
R1004 B.n991 B.n990 585
R1005 B.n992 B.n991 585
R1006 B.n989 B.n127 585
R1007 B.n130 B.n127 585
R1008 B.n988 B.n987 585
R1009 B.n987 B.n986 585
R1010 B.n129 B.n128 585
R1011 B.n985 B.n129 585
R1012 B.n983 B.n982 585
R1013 B.n984 B.n983 585
R1014 B.n981 B.n135 585
R1015 B.n135 B.n134 585
R1016 B.n980 B.n979 585
R1017 B.n979 B.n978 585
R1018 B.n137 B.n136 585
R1019 B.n977 B.n137 585
R1020 B.n975 B.n974 585
R1021 B.n976 B.n975 585
R1022 B.n973 B.n142 585
R1023 B.n142 B.n141 585
R1024 B.n972 B.n971 585
R1025 B.n971 B.n970 585
R1026 B.n1132 B.n1131 585
R1027 B.n1131 B.n1130 585
R1028 B.n627 B.n461 454.062
R1029 B.n971 B.n144 454.062
R1030 B.n625 B.n463 454.062
R1031 B.n968 B.n145 454.062
R1032 B.n969 B.n176 256.663
R1033 B.n969 B.n175 256.663
R1034 B.n969 B.n174 256.663
R1035 B.n969 B.n173 256.663
R1036 B.n969 B.n172 256.663
R1037 B.n969 B.n171 256.663
R1038 B.n969 B.n170 256.663
R1039 B.n969 B.n169 256.663
R1040 B.n969 B.n168 256.663
R1041 B.n969 B.n167 256.663
R1042 B.n969 B.n166 256.663
R1043 B.n969 B.n165 256.663
R1044 B.n969 B.n164 256.663
R1045 B.n969 B.n163 256.663
R1046 B.n969 B.n162 256.663
R1047 B.n969 B.n161 256.663
R1048 B.n969 B.n160 256.663
R1049 B.n969 B.n159 256.663
R1050 B.n969 B.n158 256.663
R1051 B.n969 B.n157 256.663
R1052 B.n969 B.n156 256.663
R1053 B.n969 B.n155 256.663
R1054 B.n969 B.n154 256.663
R1055 B.n969 B.n153 256.663
R1056 B.n969 B.n152 256.663
R1057 B.n969 B.n151 256.663
R1058 B.n969 B.n150 256.663
R1059 B.n969 B.n149 256.663
R1060 B.n969 B.n148 256.663
R1061 B.n969 B.n147 256.663
R1062 B.n969 B.n146 256.663
R1063 B.n496 B.n462 256.663
R1064 B.n502 B.n462 256.663
R1065 B.n504 B.n462 256.663
R1066 B.n510 B.n462 256.663
R1067 B.n512 B.n462 256.663
R1068 B.n518 B.n462 256.663
R1069 B.n520 B.n462 256.663
R1070 B.n526 B.n462 256.663
R1071 B.n528 B.n462 256.663
R1072 B.n534 B.n462 256.663
R1073 B.n536 B.n462 256.663
R1074 B.n542 B.n462 256.663
R1075 B.n544 B.n462 256.663
R1076 B.n551 B.n462 256.663
R1077 B.n553 B.n462 256.663
R1078 B.n559 B.n462 256.663
R1079 B.n561 B.n462 256.663
R1080 B.n570 B.n462 256.663
R1081 B.n572 B.n462 256.663
R1082 B.n578 B.n462 256.663
R1083 B.n580 B.n462 256.663
R1084 B.n586 B.n462 256.663
R1085 B.n588 B.n462 256.663
R1086 B.n594 B.n462 256.663
R1087 B.n596 B.n462 256.663
R1088 B.n602 B.n462 256.663
R1089 B.n604 B.n462 256.663
R1090 B.n610 B.n462 256.663
R1091 B.n612 B.n462 256.663
R1092 B.n618 B.n462 256.663
R1093 B.n620 B.n462 256.663
R1094 B.n565 B.t13 253.501
R1095 B.n482 B.t9 253.501
R1096 B.n181 B.t16 253.501
R1097 B.n178 B.t20 253.501
R1098 B.n627 B.n459 163.367
R1099 B.n631 B.n459 163.367
R1100 B.n631 B.n453 163.367
R1101 B.n639 B.n453 163.367
R1102 B.n639 B.n451 163.367
R1103 B.n643 B.n451 163.367
R1104 B.n643 B.n445 163.367
R1105 B.n652 B.n445 163.367
R1106 B.n652 B.n443 163.367
R1107 B.n656 B.n443 163.367
R1108 B.n656 B.n438 163.367
R1109 B.n664 B.n438 163.367
R1110 B.n664 B.n436 163.367
R1111 B.n668 B.n436 163.367
R1112 B.n668 B.n430 163.367
R1113 B.n676 B.n430 163.367
R1114 B.n676 B.n428 163.367
R1115 B.n680 B.n428 163.367
R1116 B.n680 B.n422 163.367
R1117 B.n688 B.n422 163.367
R1118 B.n688 B.n420 163.367
R1119 B.n692 B.n420 163.367
R1120 B.n692 B.n414 163.367
R1121 B.n700 B.n414 163.367
R1122 B.n700 B.n412 163.367
R1123 B.n704 B.n412 163.367
R1124 B.n704 B.n406 163.367
R1125 B.n712 B.n406 163.367
R1126 B.n712 B.n404 163.367
R1127 B.n716 B.n404 163.367
R1128 B.n716 B.n398 163.367
R1129 B.n724 B.n398 163.367
R1130 B.n724 B.n396 163.367
R1131 B.n728 B.n396 163.367
R1132 B.n728 B.n390 163.367
R1133 B.n736 B.n390 163.367
R1134 B.n736 B.n388 163.367
R1135 B.n740 B.n388 163.367
R1136 B.n740 B.n382 163.367
R1137 B.n748 B.n382 163.367
R1138 B.n748 B.n380 163.367
R1139 B.n752 B.n380 163.367
R1140 B.n752 B.n374 163.367
R1141 B.n760 B.n374 163.367
R1142 B.n760 B.n372 163.367
R1143 B.n764 B.n372 163.367
R1144 B.n764 B.n366 163.367
R1145 B.n772 B.n366 163.367
R1146 B.n772 B.n364 163.367
R1147 B.n776 B.n364 163.367
R1148 B.n776 B.n358 163.367
R1149 B.n784 B.n358 163.367
R1150 B.n784 B.n356 163.367
R1151 B.n788 B.n356 163.367
R1152 B.n788 B.n350 163.367
R1153 B.n796 B.n350 163.367
R1154 B.n796 B.n348 163.367
R1155 B.n800 B.n348 163.367
R1156 B.n800 B.n342 163.367
R1157 B.n808 B.n342 163.367
R1158 B.n808 B.n340 163.367
R1159 B.n812 B.n340 163.367
R1160 B.n812 B.n334 163.367
R1161 B.n820 B.n334 163.367
R1162 B.n820 B.n332 163.367
R1163 B.n824 B.n332 163.367
R1164 B.n824 B.n326 163.367
R1165 B.n832 B.n326 163.367
R1166 B.n832 B.n324 163.367
R1167 B.n836 B.n324 163.367
R1168 B.n836 B.n318 163.367
R1169 B.n844 B.n318 163.367
R1170 B.n844 B.n316 163.367
R1171 B.n848 B.n316 163.367
R1172 B.n848 B.n310 163.367
R1173 B.n857 B.n310 163.367
R1174 B.n857 B.n308 163.367
R1175 B.n861 B.n308 163.367
R1176 B.n861 B.n2 163.367
R1177 B.n1131 B.n2 163.367
R1178 B.n1131 B.n3 163.367
R1179 B.n1127 B.n3 163.367
R1180 B.n1127 B.n9 163.367
R1181 B.n1123 B.n9 163.367
R1182 B.n1123 B.n11 163.367
R1183 B.n1119 B.n11 163.367
R1184 B.n1119 B.n16 163.367
R1185 B.n1115 B.n16 163.367
R1186 B.n1115 B.n18 163.367
R1187 B.n1111 B.n18 163.367
R1188 B.n1111 B.n23 163.367
R1189 B.n1107 B.n23 163.367
R1190 B.n1107 B.n25 163.367
R1191 B.n1103 B.n25 163.367
R1192 B.n1103 B.n30 163.367
R1193 B.n1099 B.n30 163.367
R1194 B.n1099 B.n32 163.367
R1195 B.n1095 B.n32 163.367
R1196 B.n1095 B.n37 163.367
R1197 B.n1091 B.n37 163.367
R1198 B.n1091 B.n39 163.367
R1199 B.n1087 B.n39 163.367
R1200 B.n1087 B.n44 163.367
R1201 B.n1083 B.n44 163.367
R1202 B.n1083 B.n46 163.367
R1203 B.n1079 B.n46 163.367
R1204 B.n1079 B.n51 163.367
R1205 B.n1075 B.n51 163.367
R1206 B.n1075 B.n53 163.367
R1207 B.n1071 B.n53 163.367
R1208 B.n1071 B.n58 163.367
R1209 B.n1067 B.n58 163.367
R1210 B.n1067 B.n60 163.367
R1211 B.n1063 B.n60 163.367
R1212 B.n1063 B.n65 163.367
R1213 B.n1059 B.n65 163.367
R1214 B.n1059 B.n67 163.367
R1215 B.n1055 B.n67 163.367
R1216 B.n1055 B.n72 163.367
R1217 B.n1051 B.n72 163.367
R1218 B.n1051 B.n74 163.367
R1219 B.n1047 B.n74 163.367
R1220 B.n1047 B.n79 163.367
R1221 B.n1043 B.n79 163.367
R1222 B.n1043 B.n81 163.367
R1223 B.n1039 B.n81 163.367
R1224 B.n1039 B.n86 163.367
R1225 B.n1035 B.n86 163.367
R1226 B.n1035 B.n88 163.367
R1227 B.n1031 B.n88 163.367
R1228 B.n1031 B.n93 163.367
R1229 B.n1027 B.n93 163.367
R1230 B.n1027 B.n95 163.367
R1231 B.n1023 B.n95 163.367
R1232 B.n1023 B.n100 163.367
R1233 B.n1019 B.n100 163.367
R1234 B.n1019 B.n102 163.367
R1235 B.n1015 B.n102 163.367
R1236 B.n1015 B.n107 163.367
R1237 B.n1011 B.n107 163.367
R1238 B.n1011 B.n109 163.367
R1239 B.n1007 B.n109 163.367
R1240 B.n1007 B.n114 163.367
R1241 B.n1003 B.n114 163.367
R1242 B.n1003 B.n116 163.367
R1243 B.n999 B.n116 163.367
R1244 B.n999 B.n121 163.367
R1245 B.n995 B.n121 163.367
R1246 B.n995 B.n123 163.367
R1247 B.n991 B.n123 163.367
R1248 B.n991 B.n127 163.367
R1249 B.n987 B.n127 163.367
R1250 B.n987 B.n129 163.367
R1251 B.n983 B.n129 163.367
R1252 B.n983 B.n135 163.367
R1253 B.n979 B.n135 163.367
R1254 B.n979 B.n137 163.367
R1255 B.n975 B.n137 163.367
R1256 B.n975 B.n142 163.367
R1257 B.n971 B.n142 163.367
R1258 B.n497 B.n495 163.367
R1259 B.n501 B.n495 163.367
R1260 B.n505 B.n503 163.367
R1261 B.n509 B.n493 163.367
R1262 B.n513 B.n511 163.367
R1263 B.n517 B.n491 163.367
R1264 B.n521 B.n519 163.367
R1265 B.n525 B.n489 163.367
R1266 B.n529 B.n527 163.367
R1267 B.n533 B.n487 163.367
R1268 B.n537 B.n535 163.367
R1269 B.n541 B.n485 163.367
R1270 B.n545 B.n543 163.367
R1271 B.n550 B.n481 163.367
R1272 B.n554 B.n552 163.367
R1273 B.n558 B.n479 163.367
R1274 B.n562 B.n560 163.367
R1275 B.n569 B.n477 163.367
R1276 B.n573 B.n571 163.367
R1277 B.n577 B.n475 163.367
R1278 B.n581 B.n579 163.367
R1279 B.n585 B.n473 163.367
R1280 B.n589 B.n587 163.367
R1281 B.n593 B.n471 163.367
R1282 B.n597 B.n595 163.367
R1283 B.n601 B.n469 163.367
R1284 B.n605 B.n603 163.367
R1285 B.n609 B.n467 163.367
R1286 B.n613 B.n611 163.367
R1287 B.n617 B.n465 163.367
R1288 B.n621 B.n619 163.367
R1289 B.n625 B.n457 163.367
R1290 B.n633 B.n457 163.367
R1291 B.n633 B.n455 163.367
R1292 B.n637 B.n455 163.367
R1293 B.n637 B.n449 163.367
R1294 B.n645 B.n449 163.367
R1295 B.n645 B.n447 163.367
R1296 B.n649 B.n447 163.367
R1297 B.n649 B.n442 163.367
R1298 B.n658 B.n442 163.367
R1299 B.n658 B.n440 163.367
R1300 B.n662 B.n440 163.367
R1301 B.n662 B.n434 163.367
R1302 B.n670 B.n434 163.367
R1303 B.n670 B.n432 163.367
R1304 B.n674 B.n432 163.367
R1305 B.n674 B.n426 163.367
R1306 B.n682 B.n426 163.367
R1307 B.n682 B.n424 163.367
R1308 B.n686 B.n424 163.367
R1309 B.n686 B.n418 163.367
R1310 B.n694 B.n418 163.367
R1311 B.n694 B.n416 163.367
R1312 B.n698 B.n416 163.367
R1313 B.n698 B.n410 163.367
R1314 B.n706 B.n410 163.367
R1315 B.n706 B.n408 163.367
R1316 B.n710 B.n408 163.367
R1317 B.n710 B.n402 163.367
R1318 B.n718 B.n402 163.367
R1319 B.n718 B.n400 163.367
R1320 B.n722 B.n400 163.367
R1321 B.n722 B.n394 163.367
R1322 B.n730 B.n394 163.367
R1323 B.n730 B.n392 163.367
R1324 B.n734 B.n392 163.367
R1325 B.n734 B.n386 163.367
R1326 B.n742 B.n386 163.367
R1327 B.n742 B.n384 163.367
R1328 B.n746 B.n384 163.367
R1329 B.n746 B.n378 163.367
R1330 B.n754 B.n378 163.367
R1331 B.n754 B.n376 163.367
R1332 B.n758 B.n376 163.367
R1333 B.n758 B.n370 163.367
R1334 B.n766 B.n370 163.367
R1335 B.n766 B.n368 163.367
R1336 B.n770 B.n368 163.367
R1337 B.n770 B.n362 163.367
R1338 B.n778 B.n362 163.367
R1339 B.n778 B.n360 163.367
R1340 B.n782 B.n360 163.367
R1341 B.n782 B.n354 163.367
R1342 B.n790 B.n354 163.367
R1343 B.n790 B.n352 163.367
R1344 B.n794 B.n352 163.367
R1345 B.n794 B.n346 163.367
R1346 B.n802 B.n346 163.367
R1347 B.n802 B.n344 163.367
R1348 B.n806 B.n344 163.367
R1349 B.n806 B.n338 163.367
R1350 B.n814 B.n338 163.367
R1351 B.n814 B.n336 163.367
R1352 B.n818 B.n336 163.367
R1353 B.n818 B.n330 163.367
R1354 B.n826 B.n330 163.367
R1355 B.n826 B.n328 163.367
R1356 B.n830 B.n328 163.367
R1357 B.n830 B.n322 163.367
R1358 B.n838 B.n322 163.367
R1359 B.n838 B.n320 163.367
R1360 B.n842 B.n320 163.367
R1361 B.n842 B.n314 163.367
R1362 B.n850 B.n314 163.367
R1363 B.n850 B.n312 163.367
R1364 B.n855 B.n312 163.367
R1365 B.n855 B.n306 163.367
R1366 B.n863 B.n306 163.367
R1367 B.n864 B.n863 163.367
R1368 B.n864 B.n5 163.367
R1369 B.n6 B.n5 163.367
R1370 B.n7 B.n6 163.367
R1371 B.n869 B.n7 163.367
R1372 B.n869 B.n12 163.367
R1373 B.n13 B.n12 163.367
R1374 B.n14 B.n13 163.367
R1375 B.n874 B.n14 163.367
R1376 B.n874 B.n19 163.367
R1377 B.n20 B.n19 163.367
R1378 B.n21 B.n20 163.367
R1379 B.n879 B.n21 163.367
R1380 B.n879 B.n26 163.367
R1381 B.n27 B.n26 163.367
R1382 B.n28 B.n27 163.367
R1383 B.n884 B.n28 163.367
R1384 B.n884 B.n33 163.367
R1385 B.n34 B.n33 163.367
R1386 B.n35 B.n34 163.367
R1387 B.n889 B.n35 163.367
R1388 B.n889 B.n40 163.367
R1389 B.n41 B.n40 163.367
R1390 B.n42 B.n41 163.367
R1391 B.n894 B.n42 163.367
R1392 B.n894 B.n47 163.367
R1393 B.n48 B.n47 163.367
R1394 B.n49 B.n48 163.367
R1395 B.n899 B.n49 163.367
R1396 B.n899 B.n54 163.367
R1397 B.n55 B.n54 163.367
R1398 B.n56 B.n55 163.367
R1399 B.n904 B.n56 163.367
R1400 B.n904 B.n61 163.367
R1401 B.n62 B.n61 163.367
R1402 B.n63 B.n62 163.367
R1403 B.n909 B.n63 163.367
R1404 B.n909 B.n68 163.367
R1405 B.n69 B.n68 163.367
R1406 B.n70 B.n69 163.367
R1407 B.n914 B.n70 163.367
R1408 B.n914 B.n75 163.367
R1409 B.n76 B.n75 163.367
R1410 B.n77 B.n76 163.367
R1411 B.n919 B.n77 163.367
R1412 B.n919 B.n82 163.367
R1413 B.n83 B.n82 163.367
R1414 B.n84 B.n83 163.367
R1415 B.n924 B.n84 163.367
R1416 B.n924 B.n89 163.367
R1417 B.n90 B.n89 163.367
R1418 B.n91 B.n90 163.367
R1419 B.n929 B.n91 163.367
R1420 B.n929 B.n96 163.367
R1421 B.n97 B.n96 163.367
R1422 B.n98 B.n97 163.367
R1423 B.n934 B.n98 163.367
R1424 B.n934 B.n103 163.367
R1425 B.n104 B.n103 163.367
R1426 B.n105 B.n104 163.367
R1427 B.n939 B.n105 163.367
R1428 B.n939 B.n110 163.367
R1429 B.n111 B.n110 163.367
R1430 B.n112 B.n111 163.367
R1431 B.n944 B.n112 163.367
R1432 B.n944 B.n117 163.367
R1433 B.n118 B.n117 163.367
R1434 B.n119 B.n118 163.367
R1435 B.n949 B.n119 163.367
R1436 B.n949 B.n124 163.367
R1437 B.n125 B.n124 163.367
R1438 B.n126 B.n125 163.367
R1439 B.n954 B.n126 163.367
R1440 B.n954 B.n131 163.367
R1441 B.n132 B.n131 163.367
R1442 B.n133 B.n132 163.367
R1443 B.n959 B.n133 163.367
R1444 B.n959 B.n138 163.367
R1445 B.n139 B.n138 163.367
R1446 B.n140 B.n139 163.367
R1447 B.n964 B.n140 163.367
R1448 B.n964 B.n145 163.367
R1449 B.n185 B.n184 163.367
R1450 B.n189 B.n188 163.367
R1451 B.n193 B.n192 163.367
R1452 B.n197 B.n196 163.367
R1453 B.n201 B.n200 163.367
R1454 B.n205 B.n204 163.367
R1455 B.n209 B.n208 163.367
R1456 B.n213 B.n212 163.367
R1457 B.n217 B.n216 163.367
R1458 B.n221 B.n220 163.367
R1459 B.n225 B.n224 163.367
R1460 B.n229 B.n228 163.367
R1461 B.n233 B.n232 163.367
R1462 B.n238 B.n237 163.367
R1463 B.n242 B.n241 163.367
R1464 B.n246 B.n245 163.367
R1465 B.n250 B.n249 163.367
R1466 B.n254 B.n253 163.367
R1467 B.n258 B.n257 163.367
R1468 B.n262 B.n261 163.367
R1469 B.n266 B.n265 163.367
R1470 B.n270 B.n269 163.367
R1471 B.n274 B.n273 163.367
R1472 B.n278 B.n277 163.367
R1473 B.n282 B.n281 163.367
R1474 B.n286 B.n285 163.367
R1475 B.n290 B.n289 163.367
R1476 B.n294 B.n293 163.367
R1477 B.n298 B.n297 163.367
R1478 B.n302 B.n301 163.367
R1479 B.n968 B.n177 163.367
R1480 B.n565 B.t15 149.119
R1481 B.n178 B.t21 149.119
R1482 B.n482 B.t12 149.112
R1483 B.n181 B.t18 149.112
R1484 B.n626 B.n462 107.871
R1485 B.n970 B.n969 107.871
R1486 B.n566 B.n565 78.9338
R1487 B.n483 B.n482 78.9338
R1488 B.n182 B.n181 78.9338
R1489 B.n179 B.n178 78.9338
R1490 B.n496 B.n461 71.676
R1491 B.n502 B.n501 71.676
R1492 B.n505 B.n504 71.676
R1493 B.n510 B.n509 71.676
R1494 B.n513 B.n512 71.676
R1495 B.n518 B.n517 71.676
R1496 B.n521 B.n520 71.676
R1497 B.n526 B.n525 71.676
R1498 B.n529 B.n528 71.676
R1499 B.n534 B.n533 71.676
R1500 B.n537 B.n536 71.676
R1501 B.n542 B.n541 71.676
R1502 B.n545 B.n544 71.676
R1503 B.n551 B.n550 71.676
R1504 B.n554 B.n553 71.676
R1505 B.n559 B.n558 71.676
R1506 B.n562 B.n561 71.676
R1507 B.n570 B.n569 71.676
R1508 B.n573 B.n572 71.676
R1509 B.n578 B.n577 71.676
R1510 B.n581 B.n580 71.676
R1511 B.n586 B.n585 71.676
R1512 B.n589 B.n588 71.676
R1513 B.n594 B.n593 71.676
R1514 B.n597 B.n596 71.676
R1515 B.n602 B.n601 71.676
R1516 B.n605 B.n604 71.676
R1517 B.n610 B.n609 71.676
R1518 B.n613 B.n612 71.676
R1519 B.n618 B.n617 71.676
R1520 B.n621 B.n620 71.676
R1521 B.n146 B.n144 71.676
R1522 B.n185 B.n147 71.676
R1523 B.n189 B.n148 71.676
R1524 B.n193 B.n149 71.676
R1525 B.n197 B.n150 71.676
R1526 B.n201 B.n151 71.676
R1527 B.n205 B.n152 71.676
R1528 B.n209 B.n153 71.676
R1529 B.n213 B.n154 71.676
R1530 B.n217 B.n155 71.676
R1531 B.n221 B.n156 71.676
R1532 B.n225 B.n157 71.676
R1533 B.n229 B.n158 71.676
R1534 B.n233 B.n159 71.676
R1535 B.n238 B.n160 71.676
R1536 B.n242 B.n161 71.676
R1537 B.n246 B.n162 71.676
R1538 B.n250 B.n163 71.676
R1539 B.n254 B.n164 71.676
R1540 B.n258 B.n165 71.676
R1541 B.n262 B.n166 71.676
R1542 B.n266 B.n167 71.676
R1543 B.n270 B.n168 71.676
R1544 B.n274 B.n169 71.676
R1545 B.n278 B.n170 71.676
R1546 B.n282 B.n171 71.676
R1547 B.n286 B.n172 71.676
R1548 B.n290 B.n173 71.676
R1549 B.n294 B.n174 71.676
R1550 B.n298 B.n175 71.676
R1551 B.n302 B.n176 71.676
R1552 B.n177 B.n176 71.676
R1553 B.n301 B.n175 71.676
R1554 B.n297 B.n174 71.676
R1555 B.n293 B.n173 71.676
R1556 B.n289 B.n172 71.676
R1557 B.n285 B.n171 71.676
R1558 B.n281 B.n170 71.676
R1559 B.n277 B.n169 71.676
R1560 B.n273 B.n168 71.676
R1561 B.n269 B.n167 71.676
R1562 B.n265 B.n166 71.676
R1563 B.n261 B.n165 71.676
R1564 B.n257 B.n164 71.676
R1565 B.n253 B.n163 71.676
R1566 B.n249 B.n162 71.676
R1567 B.n245 B.n161 71.676
R1568 B.n241 B.n160 71.676
R1569 B.n237 B.n159 71.676
R1570 B.n232 B.n158 71.676
R1571 B.n228 B.n157 71.676
R1572 B.n224 B.n156 71.676
R1573 B.n220 B.n155 71.676
R1574 B.n216 B.n154 71.676
R1575 B.n212 B.n153 71.676
R1576 B.n208 B.n152 71.676
R1577 B.n204 B.n151 71.676
R1578 B.n200 B.n150 71.676
R1579 B.n196 B.n149 71.676
R1580 B.n192 B.n148 71.676
R1581 B.n188 B.n147 71.676
R1582 B.n184 B.n146 71.676
R1583 B.n497 B.n496 71.676
R1584 B.n503 B.n502 71.676
R1585 B.n504 B.n493 71.676
R1586 B.n511 B.n510 71.676
R1587 B.n512 B.n491 71.676
R1588 B.n519 B.n518 71.676
R1589 B.n520 B.n489 71.676
R1590 B.n527 B.n526 71.676
R1591 B.n528 B.n487 71.676
R1592 B.n535 B.n534 71.676
R1593 B.n536 B.n485 71.676
R1594 B.n543 B.n542 71.676
R1595 B.n544 B.n481 71.676
R1596 B.n552 B.n551 71.676
R1597 B.n553 B.n479 71.676
R1598 B.n560 B.n559 71.676
R1599 B.n561 B.n477 71.676
R1600 B.n571 B.n570 71.676
R1601 B.n572 B.n475 71.676
R1602 B.n579 B.n578 71.676
R1603 B.n580 B.n473 71.676
R1604 B.n587 B.n586 71.676
R1605 B.n588 B.n471 71.676
R1606 B.n595 B.n594 71.676
R1607 B.n596 B.n469 71.676
R1608 B.n603 B.n602 71.676
R1609 B.n604 B.n467 71.676
R1610 B.n611 B.n610 71.676
R1611 B.n612 B.n465 71.676
R1612 B.n619 B.n618 71.676
R1613 B.n620 B.n463 71.676
R1614 B.n566 B.t14 70.1864
R1615 B.n179 B.t22 70.1864
R1616 B.n483 B.t11 70.1786
R1617 B.n182 B.t19 70.1786
R1618 B.n626 B.n458 61.6404
R1619 B.n632 B.n458 61.6404
R1620 B.n632 B.n454 61.6404
R1621 B.n638 B.n454 61.6404
R1622 B.n638 B.n450 61.6404
R1623 B.n644 B.n450 61.6404
R1624 B.n644 B.n446 61.6404
R1625 B.n651 B.n446 61.6404
R1626 B.n651 B.n650 61.6404
R1627 B.n657 B.n439 61.6404
R1628 B.n663 B.n439 61.6404
R1629 B.n663 B.n435 61.6404
R1630 B.n669 B.n435 61.6404
R1631 B.n669 B.n431 61.6404
R1632 B.n675 B.n431 61.6404
R1633 B.n675 B.n427 61.6404
R1634 B.n681 B.n427 61.6404
R1635 B.n681 B.n423 61.6404
R1636 B.n687 B.n423 61.6404
R1637 B.n687 B.n419 61.6404
R1638 B.n693 B.n419 61.6404
R1639 B.n693 B.n415 61.6404
R1640 B.n699 B.n415 61.6404
R1641 B.n705 B.n411 61.6404
R1642 B.n705 B.n407 61.6404
R1643 B.n711 B.n407 61.6404
R1644 B.n711 B.n403 61.6404
R1645 B.n717 B.n403 61.6404
R1646 B.n717 B.n399 61.6404
R1647 B.n723 B.n399 61.6404
R1648 B.n723 B.n395 61.6404
R1649 B.n729 B.n395 61.6404
R1650 B.n729 B.n391 61.6404
R1651 B.n735 B.n391 61.6404
R1652 B.n741 B.n387 61.6404
R1653 B.n741 B.n383 61.6404
R1654 B.n747 B.n383 61.6404
R1655 B.n747 B.n379 61.6404
R1656 B.n753 B.n379 61.6404
R1657 B.n753 B.n375 61.6404
R1658 B.n759 B.n375 61.6404
R1659 B.n759 B.n371 61.6404
R1660 B.n765 B.n371 61.6404
R1661 B.n765 B.n367 61.6404
R1662 B.n771 B.n367 61.6404
R1663 B.n777 B.n363 61.6404
R1664 B.n777 B.n359 61.6404
R1665 B.n783 B.n359 61.6404
R1666 B.n783 B.n355 61.6404
R1667 B.n789 B.n355 61.6404
R1668 B.n789 B.n351 61.6404
R1669 B.n795 B.n351 61.6404
R1670 B.n795 B.n347 61.6404
R1671 B.n801 B.n347 61.6404
R1672 B.n801 B.n343 61.6404
R1673 B.n807 B.n343 61.6404
R1674 B.n813 B.n339 61.6404
R1675 B.n813 B.n335 61.6404
R1676 B.n819 B.n335 61.6404
R1677 B.n819 B.n331 61.6404
R1678 B.n825 B.n331 61.6404
R1679 B.n825 B.n327 61.6404
R1680 B.n831 B.n327 61.6404
R1681 B.n831 B.n323 61.6404
R1682 B.n837 B.n323 61.6404
R1683 B.n837 B.n319 61.6404
R1684 B.n843 B.n319 61.6404
R1685 B.n849 B.n315 61.6404
R1686 B.n849 B.n311 61.6404
R1687 B.n856 B.n311 61.6404
R1688 B.n856 B.n307 61.6404
R1689 B.n862 B.n307 61.6404
R1690 B.n862 B.n4 61.6404
R1691 B.n1130 B.n4 61.6404
R1692 B.n1130 B.n1129 61.6404
R1693 B.n1129 B.n1128 61.6404
R1694 B.n1128 B.n8 61.6404
R1695 B.n1122 B.n8 61.6404
R1696 B.n1122 B.n1121 61.6404
R1697 B.n1121 B.n1120 61.6404
R1698 B.n1120 B.n15 61.6404
R1699 B.n1114 B.n1113 61.6404
R1700 B.n1113 B.n1112 61.6404
R1701 B.n1112 B.n22 61.6404
R1702 B.n1106 B.n22 61.6404
R1703 B.n1106 B.n1105 61.6404
R1704 B.n1105 B.n1104 61.6404
R1705 B.n1104 B.n29 61.6404
R1706 B.n1098 B.n29 61.6404
R1707 B.n1098 B.n1097 61.6404
R1708 B.n1097 B.n1096 61.6404
R1709 B.n1096 B.n36 61.6404
R1710 B.n1090 B.n1089 61.6404
R1711 B.n1089 B.n1088 61.6404
R1712 B.n1088 B.n43 61.6404
R1713 B.n1082 B.n43 61.6404
R1714 B.n1082 B.n1081 61.6404
R1715 B.n1081 B.n1080 61.6404
R1716 B.n1080 B.n50 61.6404
R1717 B.n1074 B.n50 61.6404
R1718 B.n1074 B.n1073 61.6404
R1719 B.n1073 B.n1072 61.6404
R1720 B.n1072 B.n57 61.6404
R1721 B.n1066 B.n1065 61.6404
R1722 B.n1065 B.n1064 61.6404
R1723 B.n1064 B.n64 61.6404
R1724 B.n1058 B.n64 61.6404
R1725 B.n1058 B.n1057 61.6404
R1726 B.n1057 B.n1056 61.6404
R1727 B.n1056 B.n71 61.6404
R1728 B.n1050 B.n71 61.6404
R1729 B.n1050 B.n1049 61.6404
R1730 B.n1049 B.n1048 61.6404
R1731 B.n1048 B.n78 61.6404
R1732 B.n1042 B.n1041 61.6404
R1733 B.n1041 B.n1040 61.6404
R1734 B.n1040 B.n85 61.6404
R1735 B.n1034 B.n85 61.6404
R1736 B.n1034 B.n1033 61.6404
R1737 B.n1033 B.n1032 61.6404
R1738 B.n1032 B.n92 61.6404
R1739 B.n1026 B.n92 61.6404
R1740 B.n1026 B.n1025 61.6404
R1741 B.n1025 B.n1024 61.6404
R1742 B.n1024 B.n99 61.6404
R1743 B.n1018 B.n1017 61.6404
R1744 B.n1017 B.n1016 61.6404
R1745 B.n1016 B.n106 61.6404
R1746 B.n1010 B.n106 61.6404
R1747 B.n1010 B.n1009 61.6404
R1748 B.n1009 B.n1008 61.6404
R1749 B.n1008 B.n113 61.6404
R1750 B.n1002 B.n113 61.6404
R1751 B.n1002 B.n1001 61.6404
R1752 B.n1001 B.n1000 61.6404
R1753 B.n1000 B.n120 61.6404
R1754 B.n994 B.n120 61.6404
R1755 B.n994 B.n993 61.6404
R1756 B.n993 B.n992 61.6404
R1757 B.n986 B.n130 61.6404
R1758 B.n986 B.n985 61.6404
R1759 B.n985 B.n984 61.6404
R1760 B.n984 B.n134 61.6404
R1761 B.n978 B.n134 61.6404
R1762 B.n978 B.n977 61.6404
R1763 B.n977 B.n976 61.6404
R1764 B.n976 B.n141 61.6404
R1765 B.n970 B.n141 61.6404
R1766 B.n567 B.n566 59.5399
R1767 B.n548 B.n483 59.5399
R1768 B.n235 B.n182 59.5399
R1769 B.n180 B.n179 59.5399
R1770 B.n657 B.t10 39.8851
R1771 B.n992 B.t17 39.8851
R1772 B.t0 B.n315 36.2593
R1773 B.t1 B.n15 36.2593
R1774 B.t2 B.n339 34.4463
R1775 B.t8 B.n36 34.4463
R1776 B.n699 B.t6 32.6334
R1777 B.t7 B.n363 32.6334
R1778 B.t5 B.n57 32.6334
R1779 B.n1018 B.t3 32.6334
R1780 B.n735 B.t4 30.8204
R1781 B.t4 B.n387 30.8204
R1782 B.t23 B.n78 30.8204
R1783 B.n1042 B.t23 30.8204
R1784 B.n967 B.n966 29.5029
R1785 B.n972 B.n143 29.5029
R1786 B.n624 B.n623 29.5029
R1787 B.n628 B.n460 29.5029
R1788 B.t6 B.n411 29.0075
R1789 B.n771 B.t7 29.0075
R1790 B.n1066 B.t5 29.0075
R1791 B.t3 B.n99 29.0075
R1792 B.n807 B.t2 27.1946
R1793 B.n1090 B.t8 27.1946
R1794 B.n843 B.t0 25.3816
R1795 B.n1114 B.t1 25.3816
R1796 B.n650 B.t10 21.7558
R1797 B.n130 B.t17 21.7558
R1798 B B.n1132 18.0485
R1799 B.n183 B.n143 10.6151
R1800 B.n186 B.n183 10.6151
R1801 B.n187 B.n186 10.6151
R1802 B.n190 B.n187 10.6151
R1803 B.n191 B.n190 10.6151
R1804 B.n194 B.n191 10.6151
R1805 B.n195 B.n194 10.6151
R1806 B.n198 B.n195 10.6151
R1807 B.n199 B.n198 10.6151
R1808 B.n202 B.n199 10.6151
R1809 B.n203 B.n202 10.6151
R1810 B.n206 B.n203 10.6151
R1811 B.n207 B.n206 10.6151
R1812 B.n210 B.n207 10.6151
R1813 B.n211 B.n210 10.6151
R1814 B.n214 B.n211 10.6151
R1815 B.n215 B.n214 10.6151
R1816 B.n218 B.n215 10.6151
R1817 B.n219 B.n218 10.6151
R1818 B.n222 B.n219 10.6151
R1819 B.n223 B.n222 10.6151
R1820 B.n226 B.n223 10.6151
R1821 B.n227 B.n226 10.6151
R1822 B.n230 B.n227 10.6151
R1823 B.n231 B.n230 10.6151
R1824 B.n234 B.n231 10.6151
R1825 B.n239 B.n236 10.6151
R1826 B.n240 B.n239 10.6151
R1827 B.n243 B.n240 10.6151
R1828 B.n244 B.n243 10.6151
R1829 B.n247 B.n244 10.6151
R1830 B.n248 B.n247 10.6151
R1831 B.n251 B.n248 10.6151
R1832 B.n252 B.n251 10.6151
R1833 B.n256 B.n255 10.6151
R1834 B.n259 B.n256 10.6151
R1835 B.n260 B.n259 10.6151
R1836 B.n263 B.n260 10.6151
R1837 B.n264 B.n263 10.6151
R1838 B.n267 B.n264 10.6151
R1839 B.n268 B.n267 10.6151
R1840 B.n271 B.n268 10.6151
R1841 B.n272 B.n271 10.6151
R1842 B.n275 B.n272 10.6151
R1843 B.n276 B.n275 10.6151
R1844 B.n279 B.n276 10.6151
R1845 B.n280 B.n279 10.6151
R1846 B.n283 B.n280 10.6151
R1847 B.n284 B.n283 10.6151
R1848 B.n287 B.n284 10.6151
R1849 B.n288 B.n287 10.6151
R1850 B.n291 B.n288 10.6151
R1851 B.n292 B.n291 10.6151
R1852 B.n295 B.n292 10.6151
R1853 B.n296 B.n295 10.6151
R1854 B.n299 B.n296 10.6151
R1855 B.n300 B.n299 10.6151
R1856 B.n303 B.n300 10.6151
R1857 B.n304 B.n303 10.6151
R1858 B.n967 B.n304 10.6151
R1859 B.n624 B.n456 10.6151
R1860 B.n634 B.n456 10.6151
R1861 B.n635 B.n634 10.6151
R1862 B.n636 B.n635 10.6151
R1863 B.n636 B.n448 10.6151
R1864 B.n646 B.n448 10.6151
R1865 B.n647 B.n646 10.6151
R1866 B.n648 B.n647 10.6151
R1867 B.n648 B.n441 10.6151
R1868 B.n659 B.n441 10.6151
R1869 B.n660 B.n659 10.6151
R1870 B.n661 B.n660 10.6151
R1871 B.n661 B.n433 10.6151
R1872 B.n671 B.n433 10.6151
R1873 B.n672 B.n671 10.6151
R1874 B.n673 B.n672 10.6151
R1875 B.n673 B.n425 10.6151
R1876 B.n683 B.n425 10.6151
R1877 B.n684 B.n683 10.6151
R1878 B.n685 B.n684 10.6151
R1879 B.n685 B.n417 10.6151
R1880 B.n695 B.n417 10.6151
R1881 B.n696 B.n695 10.6151
R1882 B.n697 B.n696 10.6151
R1883 B.n697 B.n409 10.6151
R1884 B.n707 B.n409 10.6151
R1885 B.n708 B.n707 10.6151
R1886 B.n709 B.n708 10.6151
R1887 B.n709 B.n401 10.6151
R1888 B.n719 B.n401 10.6151
R1889 B.n720 B.n719 10.6151
R1890 B.n721 B.n720 10.6151
R1891 B.n721 B.n393 10.6151
R1892 B.n731 B.n393 10.6151
R1893 B.n732 B.n731 10.6151
R1894 B.n733 B.n732 10.6151
R1895 B.n733 B.n385 10.6151
R1896 B.n743 B.n385 10.6151
R1897 B.n744 B.n743 10.6151
R1898 B.n745 B.n744 10.6151
R1899 B.n745 B.n377 10.6151
R1900 B.n755 B.n377 10.6151
R1901 B.n756 B.n755 10.6151
R1902 B.n757 B.n756 10.6151
R1903 B.n757 B.n369 10.6151
R1904 B.n767 B.n369 10.6151
R1905 B.n768 B.n767 10.6151
R1906 B.n769 B.n768 10.6151
R1907 B.n769 B.n361 10.6151
R1908 B.n779 B.n361 10.6151
R1909 B.n780 B.n779 10.6151
R1910 B.n781 B.n780 10.6151
R1911 B.n781 B.n353 10.6151
R1912 B.n791 B.n353 10.6151
R1913 B.n792 B.n791 10.6151
R1914 B.n793 B.n792 10.6151
R1915 B.n793 B.n345 10.6151
R1916 B.n803 B.n345 10.6151
R1917 B.n804 B.n803 10.6151
R1918 B.n805 B.n804 10.6151
R1919 B.n805 B.n337 10.6151
R1920 B.n815 B.n337 10.6151
R1921 B.n816 B.n815 10.6151
R1922 B.n817 B.n816 10.6151
R1923 B.n817 B.n329 10.6151
R1924 B.n827 B.n329 10.6151
R1925 B.n828 B.n827 10.6151
R1926 B.n829 B.n828 10.6151
R1927 B.n829 B.n321 10.6151
R1928 B.n839 B.n321 10.6151
R1929 B.n840 B.n839 10.6151
R1930 B.n841 B.n840 10.6151
R1931 B.n841 B.n313 10.6151
R1932 B.n851 B.n313 10.6151
R1933 B.n852 B.n851 10.6151
R1934 B.n854 B.n852 10.6151
R1935 B.n854 B.n853 10.6151
R1936 B.n853 B.n305 10.6151
R1937 B.n865 B.n305 10.6151
R1938 B.n866 B.n865 10.6151
R1939 B.n867 B.n866 10.6151
R1940 B.n868 B.n867 10.6151
R1941 B.n870 B.n868 10.6151
R1942 B.n871 B.n870 10.6151
R1943 B.n872 B.n871 10.6151
R1944 B.n873 B.n872 10.6151
R1945 B.n875 B.n873 10.6151
R1946 B.n876 B.n875 10.6151
R1947 B.n877 B.n876 10.6151
R1948 B.n878 B.n877 10.6151
R1949 B.n880 B.n878 10.6151
R1950 B.n881 B.n880 10.6151
R1951 B.n882 B.n881 10.6151
R1952 B.n883 B.n882 10.6151
R1953 B.n885 B.n883 10.6151
R1954 B.n886 B.n885 10.6151
R1955 B.n887 B.n886 10.6151
R1956 B.n888 B.n887 10.6151
R1957 B.n890 B.n888 10.6151
R1958 B.n891 B.n890 10.6151
R1959 B.n892 B.n891 10.6151
R1960 B.n893 B.n892 10.6151
R1961 B.n895 B.n893 10.6151
R1962 B.n896 B.n895 10.6151
R1963 B.n897 B.n896 10.6151
R1964 B.n898 B.n897 10.6151
R1965 B.n900 B.n898 10.6151
R1966 B.n901 B.n900 10.6151
R1967 B.n902 B.n901 10.6151
R1968 B.n903 B.n902 10.6151
R1969 B.n905 B.n903 10.6151
R1970 B.n906 B.n905 10.6151
R1971 B.n907 B.n906 10.6151
R1972 B.n908 B.n907 10.6151
R1973 B.n910 B.n908 10.6151
R1974 B.n911 B.n910 10.6151
R1975 B.n912 B.n911 10.6151
R1976 B.n913 B.n912 10.6151
R1977 B.n915 B.n913 10.6151
R1978 B.n916 B.n915 10.6151
R1979 B.n917 B.n916 10.6151
R1980 B.n918 B.n917 10.6151
R1981 B.n920 B.n918 10.6151
R1982 B.n921 B.n920 10.6151
R1983 B.n922 B.n921 10.6151
R1984 B.n923 B.n922 10.6151
R1985 B.n925 B.n923 10.6151
R1986 B.n926 B.n925 10.6151
R1987 B.n927 B.n926 10.6151
R1988 B.n928 B.n927 10.6151
R1989 B.n930 B.n928 10.6151
R1990 B.n931 B.n930 10.6151
R1991 B.n932 B.n931 10.6151
R1992 B.n933 B.n932 10.6151
R1993 B.n935 B.n933 10.6151
R1994 B.n936 B.n935 10.6151
R1995 B.n937 B.n936 10.6151
R1996 B.n938 B.n937 10.6151
R1997 B.n940 B.n938 10.6151
R1998 B.n941 B.n940 10.6151
R1999 B.n942 B.n941 10.6151
R2000 B.n943 B.n942 10.6151
R2001 B.n945 B.n943 10.6151
R2002 B.n946 B.n945 10.6151
R2003 B.n947 B.n946 10.6151
R2004 B.n948 B.n947 10.6151
R2005 B.n950 B.n948 10.6151
R2006 B.n951 B.n950 10.6151
R2007 B.n952 B.n951 10.6151
R2008 B.n953 B.n952 10.6151
R2009 B.n955 B.n953 10.6151
R2010 B.n956 B.n955 10.6151
R2011 B.n957 B.n956 10.6151
R2012 B.n958 B.n957 10.6151
R2013 B.n960 B.n958 10.6151
R2014 B.n961 B.n960 10.6151
R2015 B.n962 B.n961 10.6151
R2016 B.n963 B.n962 10.6151
R2017 B.n965 B.n963 10.6151
R2018 B.n966 B.n965 10.6151
R2019 B.n498 B.n460 10.6151
R2020 B.n499 B.n498 10.6151
R2021 B.n500 B.n499 10.6151
R2022 B.n500 B.n494 10.6151
R2023 B.n506 B.n494 10.6151
R2024 B.n507 B.n506 10.6151
R2025 B.n508 B.n507 10.6151
R2026 B.n508 B.n492 10.6151
R2027 B.n514 B.n492 10.6151
R2028 B.n515 B.n514 10.6151
R2029 B.n516 B.n515 10.6151
R2030 B.n516 B.n490 10.6151
R2031 B.n522 B.n490 10.6151
R2032 B.n523 B.n522 10.6151
R2033 B.n524 B.n523 10.6151
R2034 B.n524 B.n488 10.6151
R2035 B.n530 B.n488 10.6151
R2036 B.n531 B.n530 10.6151
R2037 B.n532 B.n531 10.6151
R2038 B.n532 B.n486 10.6151
R2039 B.n538 B.n486 10.6151
R2040 B.n539 B.n538 10.6151
R2041 B.n540 B.n539 10.6151
R2042 B.n540 B.n484 10.6151
R2043 B.n546 B.n484 10.6151
R2044 B.n547 B.n546 10.6151
R2045 B.n549 B.n480 10.6151
R2046 B.n555 B.n480 10.6151
R2047 B.n556 B.n555 10.6151
R2048 B.n557 B.n556 10.6151
R2049 B.n557 B.n478 10.6151
R2050 B.n563 B.n478 10.6151
R2051 B.n564 B.n563 10.6151
R2052 B.n568 B.n564 10.6151
R2053 B.n574 B.n476 10.6151
R2054 B.n575 B.n574 10.6151
R2055 B.n576 B.n575 10.6151
R2056 B.n576 B.n474 10.6151
R2057 B.n582 B.n474 10.6151
R2058 B.n583 B.n582 10.6151
R2059 B.n584 B.n583 10.6151
R2060 B.n584 B.n472 10.6151
R2061 B.n590 B.n472 10.6151
R2062 B.n591 B.n590 10.6151
R2063 B.n592 B.n591 10.6151
R2064 B.n592 B.n470 10.6151
R2065 B.n598 B.n470 10.6151
R2066 B.n599 B.n598 10.6151
R2067 B.n600 B.n599 10.6151
R2068 B.n600 B.n468 10.6151
R2069 B.n606 B.n468 10.6151
R2070 B.n607 B.n606 10.6151
R2071 B.n608 B.n607 10.6151
R2072 B.n608 B.n466 10.6151
R2073 B.n614 B.n466 10.6151
R2074 B.n615 B.n614 10.6151
R2075 B.n616 B.n615 10.6151
R2076 B.n616 B.n464 10.6151
R2077 B.n622 B.n464 10.6151
R2078 B.n623 B.n622 10.6151
R2079 B.n629 B.n628 10.6151
R2080 B.n630 B.n629 10.6151
R2081 B.n630 B.n452 10.6151
R2082 B.n640 B.n452 10.6151
R2083 B.n641 B.n640 10.6151
R2084 B.n642 B.n641 10.6151
R2085 B.n642 B.n444 10.6151
R2086 B.n653 B.n444 10.6151
R2087 B.n654 B.n653 10.6151
R2088 B.n655 B.n654 10.6151
R2089 B.n655 B.n437 10.6151
R2090 B.n665 B.n437 10.6151
R2091 B.n666 B.n665 10.6151
R2092 B.n667 B.n666 10.6151
R2093 B.n667 B.n429 10.6151
R2094 B.n677 B.n429 10.6151
R2095 B.n678 B.n677 10.6151
R2096 B.n679 B.n678 10.6151
R2097 B.n679 B.n421 10.6151
R2098 B.n689 B.n421 10.6151
R2099 B.n690 B.n689 10.6151
R2100 B.n691 B.n690 10.6151
R2101 B.n691 B.n413 10.6151
R2102 B.n701 B.n413 10.6151
R2103 B.n702 B.n701 10.6151
R2104 B.n703 B.n702 10.6151
R2105 B.n703 B.n405 10.6151
R2106 B.n713 B.n405 10.6151
R2107 B.n714 B.n713 10.6151
R2108 B.n715 B.n714 10.6151
R2109 B.n715 B.n397 10.6151
R2110 B.n725 B.n397 10.6151
R2111 B.n726 B.n725 10.6151
R2112 B.n727 B.n726 10.6151
R2113 B.n727 B.n389 10.6151
R2114 B.n737 B.n389 10.6151
R2115 B.n738 B.n737 10.6151
R2116 B.n739 B.n738 10.6151
R2117 B.n739 B.n381 10.6151
R2118 B.n749 B.n381 10.6151
R2119 B.n750 B.n749 10.6151
R2120 B.n751 B.n750 10.6151
R2121 B.n751 B.n373 10.6151
R2122 B.n761 B.n373 10.6151
R2123 B.n762 B.n761 10.6151
R2124 B.n763 B.n762 10.6151
R2125 B.n763 B.n365 10.6151
R2126 B.n773 B.n365 10.6151
R2127 B.n774 B.n773 10.6151
R2128 B.n775 B.n774 10.6151
R2129 B.n775 B.n357 10.6151
R2130 B.n785 B.n357 10.6151
R2131 B.n786 B.n785 10.6151
R2132 B.n787 B.n786 10.6151
R2133 B.n787 B.n349 10.6151
R2134 B.n797 B.n349 10.6151
R2135 B.n798 B.n797 10.6151
R2136 B.n799 B.n798 10.6151
R2137 B.n799 B.n341 10.6151
R2138 B.n809 B.n341 10.6151
R2139 B.n810 B.n809 10.6151
R2140 B.n811 B.n810 10.6151
R2141 B.n811 B.n333 10.6151
R2142 B.n821 B.n333 10.6151
R2143 B.n822 B.n821 10.6151
R2144 B.n823 B.n822 10.6151
R2145 B.n823 B.n325 10.6151
R2146 B.n833 B.n325 10.6151
R2147 B.n834 B.n833 10.6151
R2148 B.n835 B.n834 10.6151
R2149 B.n835 B.n317 10.6151
R2150 B.n845 B.n317 10.6151
R2151 B.n846 B.n845 10.6151
R2152 B.n847 B.n846 10.6151
R2153 B.n847 B.n309 10.6151
R2154 B.n858 B.n309 10.6151
R2155 B.n859 B.n858 10.6151
R2156 B.n860 B.n859 10.6151
R2157 B.n860 B.n0 10.6151
R2158 B.n1126 B.n1 10.6151
R2159 B.n1126 B.n1125 10.6151
R2160 B.n1125 B.n1124 10.6151
R2161 B.n1124 B.n10 10.6151
R2162 B.n1118 B.n10 10.6151
R2163 B.n1118 B.n1117 10.6151
R2164 B.n1117 B.n1116 10.6151
R2165 B.n1116 B.n17 10.6151
R2166 B.n1110 B.n17 10.6151
R2167 B.n1110 B.n1109 10.6151
R2168 B.n1109 B.n1108 10.6151
R2169 B.n1108 B.n24 10.6151
R2170 B.n1102 B.n24 10.6151
R2171 B.n1102 B.n1101 10.6151
R2172 B.n1101 B.n1100 10.6151
R2173 B.n1100 B.n31 10.6151
R2174 B.n1094 B.n31 10.6151
R2175 B.n1094 B.n1093 10.6151
R2176 B.n1093 B.n1092 10.6151
R2177 B.n1092 B.n38 10.6151
R2178 B.n1086 B.n38 10.6151
R2179 B.n1086 B.n1085 10.6151
R2180 B.n1085 B.n1084 10.6151
R2181 B.n1084 B.n45 10.6151
R2182 B.n1078 B.n45 10.6151
R2183 B.n1078 B.n1077 10.6151
R2184 B.n1077 B.n1076 10.6151
R2185 B.n1076 B.n52 10.6151
R2186 B.n1070 B.n52 10.6151
R2187 B.n1070 B.n1069 10.6151
R2188 B.n1069 B.n1068 10.6151
R2189 B.n1068 B.n59 10.6151
R2190 B.n1062 B.n59 10.6151
R2191 B.n1062 B.n1061 10.6151
R2192 B.n1061 B.n1060 10.6151
R2193 B.n1060 B.n66 10.6151
R2194 B.n1054 B.n66 10.6151
R2195 B.n1054 B.n1053 10.6151
R2196 B.n1053 B.n1052 10.6151
R2197 B.n1052 B.n73 10.6151
R2198 B.n1046 B.n73 10.6151
R2199 B.n1046 B.n1045 10.6151
R2200 B.n1045 B.n1044 10.6151
R2201 B.n1044 B.n80 10.6151
R2202 B.n1038 B.n80 10.6151
R2203 B.n1038 B.n1037 10.6151
R2204 B.n1037 B.n1036 10.6151
R2205 B.n1036 B.n87 10.6151
R2206 B.n1030 B.n87 10.6151
R2207 B.n1030 B.n1029 10.6151
R2208 B.n1029 B.n1028 10.6151
R2209 B.n1028 B.n94 10.6151
R2210 B.n1022 B.n94 10.6151
R2211 B.n1022 B.n1021 10.6151
R2212 B.n1021 B.n1020 10.6151
R2213 B.n1020 B.n101 10.6151
R2214 B.n1014 B.n101 10.6151
R2215 B.n1014 B.n1013 10.6151
R2216 B.n1013 B.n1012 10.6151
R2217 B.n1012 B.n108 10.6151
R2218 B.n1006 B.n108 10.6151
R2219 B.n1006 B.n1005 10.6151
R2220 B.n1005 B.n1004 10.6151
R2221 B.n1004 B.n115 10.6151
R2222 B.n998 B.n115 10.6151
R2223 B.n998 B.n997 10.6151
R2224 B.n997 B.n996 10.6151
R2225 B.n996 B.n122 10.6151
R2226 B.n990 B.n122 10.6151
R2227 B.n990 B.n989 10.6151
R2228 B.n989 B.n988 10.6151
R2229 B.n988 B.n128 10.6151
R2230 B.n982 B.n128 10.6151
R2231 B.n982 B.n981 10.6151
R2232 B.n981 B.n980 10.6151
R2233 B.n980 B.n136 10.6151
R2234 B.n974 B.n136 10.6151
R2235 B.n974 B.n973 10.6151
R2236 B.n973 B.n972 10.6151
R2237 B.n236 B.n235 6.5566
R2238 B.n252 B.n180 6.5566
R2239 B.n549 B.n548 6.5566
R2240 B.n568 B.n567 6.5566
R2241 B.n235 B.n234 4.05904
R2242 B.n255 B.n180 4.05904
R2243 B.n548 B.n547 4.05904
R2244 B.n567 B.n476 4.05904
R2245 B.n1132 B.n0 2.81026
R2246 B.n1132 B.n1 2.81026
R2247 VN.n108 VN.n107 161.3
R2248 VN.n106 VN.n56 161.3
R2249 VN.n105 VN.n104 161.3
R2250 VN.n103 VN.n57 161.3
R2251 VN.n102 VN.n101 161.3
R2252 VN.n100 VN.n58 161.3
R2253 VN.n99 VN.n98 161.3
R2254 VN.n97 VN.n59 161.3
R2255 VN.n96 VN.n95 161.3
R2256 VN.n94 VN.n60 161.3
R2257 VN.n93 VN.n92 161.3
R2258 VN.n91 VN.n62 161.3
R2259 VN.n90 VN.n89 161.3
R2260 VN.n88 VN.n63 161.3
R2261 VN.n87 VN.n86 161.3
R2262 VN.n85 VN.n64 161.3
R2263 VN.n84 VN.n83 161.3
R2264 VN.n82 VN.n65 161.3
R2265 VN.n81 VN.n80 161.3
R2266 VN.n79 VN.n66 161.3
R2267 VN.n78 VN.n77 161.3
R2268 VN.n76 VN.n67 161.3
R2269 VN.n75 VN.n74 161.3
R2270 VN.n73 VN.n68 161.3
R2271 VN.n72 VN.n71 161.3
R2272 VN.n53 VN.n52 161.3
R2273 VN.n51 VN.n1 161.3
R2274 VN.n50 VN.n49 161.3
R2275 VN.n48 VN.n2 161.3
R2276 VN.n47 VN.n46 161.3
R2277 VN.n45 VN.n3 161.3
R2278 VN.n44 VN.n43 161.3
R2279 VN.n42 VN.n4 161.3
R2280 VN.n41 VN.n40 161.3
R2281 VN.n38 VN.n5 161.3
R2282 VN.n37 VN.n36 161.3
R2283 VN.n35 VN.n6 161.3
R2284 VN.n34 VN.n33 161.3
R2285 VN.n32 VN.n7 161.3
R2286 VN.n31 VN.n30 161.3
R2287 VN.n29 VN.n8 161.3
R2288 VN.n28 VN.n27 161.3
R2289 VN.n26 VN.n9 161.3
R2290 VN.n25 VN.n24 161.3
R2291 VN.n23 VN.n10 161.3
R2292 VN.n22 VN.n21 161.3
R2293 VN.n20 VN.n11 161.3
R2294 VN.n19 VN.n18 161.3
R2295 VN.n17 VN.n12 161.3
R2296 VN.n16 VN.n15 161.3
R2297 VN.n54 VN.n0 83.3598
R2298 VN.n109 VN.n55 83.3598
R2299 VN.n69 VN.t4 77.093
R2300 VN.n13 VN.t8 77.093
R2301 VN.n14 VN.n13 71.5921
R2302 VN.n70 VN.n69 71.5921
R2303 VN VN.n109 55.6837
R2304 VN.n46 VN.n2 50.7491
R2305 VN.n101 VN.n57 50.7491
R2306 VN.n27 VN.t1 44.2053
R2307 VN.n14 VN.t5 44.2053
R2308 VN.n39 VN.t9 44.2053
R2309 VN.n0 VN.t3 44.2053
R2310 VN.n83 VN.t7 44.2053
R2311 VN.n70 VN.t6 44.2053
R2312 VN.n61 VN.t2 44.2053
R2313 VN.n55 VN.t0 44.2053
R2314 VN.n21 VN.n20 43.9677
R2315 VN.n33 VN.n6 43.9677
R2316 VN.n77 VN.n76 43.9677
R2317 VN.n89 VN.n62 43.9677
R2318 VN.n21 VN.n10 37.1863
R2319 VN.n33 VN.n32 37.1863
R2320 VN.n77 VN.n66 37.1863
R2321 VN.n89 VN.n88 37.1863
R2322 VN.n46 VN.n45 30.405
R2323 VN.n101 VN.n100 30.405
R2324 VN.n15 VN.n12 24.5923
R2325 VN.n19 VN.n12 24.5923
R2326 VN.n20 VN.n19 24.5923
R2327 VN.n25 VN.n10 24.5923
R2328 VN.n26 VN.n25 24.5923
R2329 VN.n27 VN.n26 24.5923
R2330 VN.n27 VN.n8 24.5923
R2331 VN.n31 VN.n8 24.5923
R2332 VN.n32 VN.n31 24.5923
R2333 VN.n37 VN.n6 24.5923
R2334 VN.n38 VN.n37 24.5923
R2335 VN.n40 VN.n38 24.5923
R2336 VN.n44 VN.n4 24.5923
R2337 VN.n45 VN.n44 24.5923
R2338 VN.n50 VN.n2 24.5923
R2339 VN.n51 VN.n50 24.5923
R2340 VN.n52 VN.n51 24.5923
R2341 VN.n76 VN.n75 24.5923
R2342 VN.n75 VN.n68 24.5923
R2343 VN.n71 VN.n68 24.5923
R2344 VN.n88 VN.n87 24.5923
R2345 VN.n87 VN.n64 24.5923
R2346 VN.n83 VN.n64 24.5923
R2347 VN.n83 VN.n82 24.5923
R2348 VN.n82 VN.n81 24.5923
R2349 VN.n81 VN.n66 24.5923
R2350 VN.n100 VN.n99 24.5923
R2351 VN.n99 VN.n59 24.5923
R2352 VN.n95 VN.n94 24.5923
R2353 VN.n94 VN.n93 24.5923
R2354 VN.n93 VN.n62 24.5923
R2355 VN.n107 VN.n106 24.5923
R2356 VN.n106 VN.n105 24.5923
R2357 VN.n105 VN.n57 24.5923
R2358 VN.n39 VN.n4 21.1495
R2359 VN.n61 VN.n59 21.1495
R2360 VN.n52 VN.n0 6.88621
R2361 VN.n107 VN.n55 6.88621
R2362 VN.n15 VN.n14 3.44336
R2363 VN.n40 VN.n39 3.44336
R2364 VN.n71 VN.n70 3.44336
R2365 VN.n95 VN.n61 3.44336
R2366 VN.n72 VN.n69 3.23944
R2367 VN.n16 VN.n13 3.23944
R2368 VN.n109 VN.n108 0.354861
R2369 VN.n54 VN.n53 0.354861
R2370 VN VN.n54 0.267071
R2371 VN.n108 VN.n56 0.189894
R2372 VN.n104 VN.n56 0.189894
R2373 VN.n104 VN.n103 0.189894
R2374 VN.n103 VN.n102 0.189894
R2375 VN.n102 VN.n58 0.189894
R2376 VN.n98 VN.n58 0.189894
R2377 VN.n98 VN.n97 0.189894
R2378 VN.n97 VN.n96 0.189894
R2379 VN.n96 VN.n60 0.189894
R2380 VN.n92 VN.n60 0.189894
R2381 VN.n92 VN.n91 0.189894
R2382 VN.n91 VN.n90 0.189894
R2383 VN.n90 VN.n63 0.189894
R2384 VN.n86 VN.n63 0.189894
R2385 VN.n86 VN.n85 0.189894
R2386 VN.n85 VN.n84 0.189894
R2387 VN.n84 VN.n65 0.189894
R2388 VN.n80 VN.n65 0.189894
R2389 VN.n80 VN.n79 0.189894
R2390 VN.n79 VN.n78 0.189894
R2391 VN.n78 VN.n67 0.189894
R2392 VN.n74 VN.n67 0.189894
R2393 VN.n74 VN.n73 0.189894
R2394 VN.n73 VN.n72 0.189894
R2395 VN.n17 VN.n16 0.189894
R2396 VN.n18 VN.n17 0.189894
R2397 VN.n18 VN.n11 0.189894
R2398 VN.n22 VN.n11 0.189894
R2399 VN.n23 VN.n22 0.189894
R2400 VN.n24 VN.n23 0.189894
R2401 VN.n24 VN.n9 0.189894
R2402 VN.n28 VN.n9 0.189894
R2403 VN.n29 VN.n28 0.189894
R2404 VN.n30 VN.n29 0.189894
R2405 VN.n30 VN.n7 0.189894
R2406 VN.n34 VN.n7 0.189894
R2407 VN.n35 VN.n34 0.189894
R2408 VN.n36 VN.n35 0.189894
R2409 VN.n36 VN.n5 0.189894
R2410 VN.n41 VN.n5 0.189894
R2411 VN.n42 VN.n41 0.189894
R2412 VN.n43 VN.n42 0.189894
R2413 VN.n43 VN.n3 0.189894
R2414 VN.n47 VN.n3 0.189894
R2415 VN.n48 VN.n47 0.189894
R2416 VN.n49 VN.n48 0.189894
R2417 VN.n49 VN.n1 0.189894
R2418 VN.n53 VN.n1 0.189894
R2419 VDD2.n1 VDD2.t1 74.1299
R2420 VDD2.n4 VDD2.t9 70.6214
R2421 VDD2.n3 VDD2.n2 70.3101
R2422 VDD2 VDD2.n7 70.3082
R2423 VDD2.n6 VDD2.n5 67.7351
R2424 VDD2.n1 VDD2.n0 67.734
R2425 VDD2.n4 VDD2.n3 46.295
R2426 VDD2.n6 VDD2.n4 3.50912
R2427 VDD2.n7 VDD2.t3 2.8868
R2428 VDD2.n7 VDD2.t5 2.8868
R2429 VDD2.n5 VDD2.t7 2.8868
R2430 VDD2.n5 VDD2.t2 2.8868
R2431 VDD2.n2 VDD2.t0 2.8868
R2432 VDD2.n2 VDD2.t6 2.8868
R2433 VDD2.n0 VDD2.t4 2.8868
R2434 VDD2.n0 VDD2.t8 2.8868
R2435 VDD2 VDD2.n6 0.935845
R2436 VDD2.n3 VDD2.n1 0.822309
C0 VN VTAIL 8.37265f
C1 VP VTAIL 8.38704f
C2 VN VDD1 0.156125f
C3 VP VDD1 7.2945f
C4 VN VDD2 6.72506f
C5 VP VDD2 0.72869f
C6 VTAIL VDD1 8.96354f
C7 VTAIL VDD2 9.02386f
C8 VDD1 VDD2 2.9155f
C9 VP VN 9.11769f
C10 VDD2 B 7.67567f
C11 VDD1 B 7.61616f
C12 VTAIL B 6.376286f
C13 VN B 22.951448f
C14 VP B 21.512283f
C15 VDD2.t1 B 1.57886f
C16 VDD2.t4 B 0.142993f
C17 VDD2.t8 B 0.142993f
C18 VDD2.n0 B 1.2217f
C19 VDD2.n1 B 1.1225f
C20 VDD2.t0 B 0.142993f
C21 VDD2.t6 B 0.142993f
C22 VDD2.n2 B 1.2486f
C23 VDD2.n3 B 3.34773f
C24 VDD2.t9 B 1.55166f
C25 VDD2.n4 B 3.32609f
C26 VDD2.t7 B 0.142993f
C27 VDD2.t2 B 0.142993f
C28 VDD2.n5 B 1.22171f
C29 VDD2.n6 B 0.583725f
C30 VDD2.t3 B 0.142993f
C31 VDD2.t5 B 0.142993f
C32 VDD2.n7 B 1.24855f
C33 VN.t3 B 1.30367f
C34 VN.n0 B 0.548292f
C35 VN.n1 B 0.019057f
C36 VN.n2 B 0.034621f
C37 VN.n3 B 0.019057f
C38 VN.n4 B 0.032898f
C39 VN.n5 B 0.019057f
C40 VN.n6 B 0.036878f
C41 VN.n7 B 0.019057f
C42 VN.n8 B 0.03534f
C43 VN.n9 B 0.019057f
C44 VN.t1 B 1.30367f
C45 VN.n10 B 0.038176f
C46 VN.n11 B 0.019057f
C47 VN.n12 B 0.03534f
C48 VN.t8 B 1.56833f
C49 VN.n13 B 0.512723f
C50 VN.t5 B 1.30367f
C51 VN.n14 B 0.535616f
C52 VN.n15 B 0.020336f
C53 VN.n16 B 0.241921f
C54 VN.n17 B 0.019057f
C55 VN.n18 B 0.019057f
C56 VN.n19 B 0.03534f
C57 VN.n20 B 0.036878f
C58 VN.n21 B 0.015692f
C59 VN.n22 B 0.019057f
C60 VN.n23 B 0.019057f
C61 VN.n24 B 0.019057f
C62 VN.n25 B 0.03534f
C63 VN.n26 B 0.03534f
C64 VN.n27 B 0.492091f
C65 VN.n28 B 0.019057f
C66 VN.n29 B 0.019057f
C67 VN.n30 B 0.019057f
C68 VN.n31 B 0.03534f
C69 VN.n32 B 0.038176f
C70 VN.n33 B 0.015692f
C71 VN.n34 B 0.019057f
C72 VN.n35 B 0.019057f
C73 VN.n36 B 0.019057f
C74 VN.n37 B 0.03534f
C75 VN.n38 B 0.03534f
C76 VN.t9 B 1.30367f
C77 VN.n39 B 0.474197f
C78 VN.n40 B 0.020336f
C79 VN.n41 B 0.019057f
C80 VN.n42 B 0.019057f
C81 VN.n43 B 0.019057f
C82 VN.n44 B 0.03534f
C83 VN.n45 B 0.037875f
C84 VN.n46 B 0.01825f
C85 VN.n47 B 0.019057f
C86 VN.n48 B 0.019057f
C87 VN.n49 B 0.019057f
C88 VN.n50 B 0.03534f
C89 VN.n51 B 0.03534f
C90 VN.n52 B 0.022779f
C91 VN.n53 B 0.030753f
C92 VN.n54 B 0.055459f
C93 VN.t0 B 1.30367f
C94 VN.n55 B 0.548292f
C95 VN.n56 B 0.019057f
C96 VN.n57 B 0.034621f
C97 VN.n58 B 0.019057f
C98 VN.n59 B 0.032898f
C99 VN.n60 B 0.019057f
C100 VN.t2 B 1.30367f
C101 VN.n61 B 0.474197f
C102 VN.n62 B 0.036878f
C103 VN.n63 B 0.019057f
C104 VN.n64 B 0.03534f
C105 VN.n65 B 0.019057f
C106 VN.t7 B 1.30367f
C107 VN.n66 B 0.038176f
C108 VN.n67 B 0.019057f
C109 VN.n68 B 0.03534f
C110 VN.t4 B 1.56833f
C111 VN.n69 B 0.512723f
C112 VN.t6 B 1.30367f
C113 VN.n70 B 0.535616f
C114 VN.n71 B 0.020336f
C115 VN.n72 B 0.241921f
C116 VN.n73 B 0.019057f
C117 VN.n74 B 0.019057f
C118 VN.n75 B 0.03534f
C119 VN.n76 B 0.036878f
C120 VN.n77 B 0.015692f
C121 VN.n78 B 0.019057f
C122 VN.n79 B 0.019057f
C123 VN.n80 B 0.019057f
C124 VN.n81 B 0.03534f
C125 VN.n82 B 0.03534f
C126 VN.n83 B 0.492091f
C127 VN.n84 B 0.019057f
C128 VN.n85 B 0.019057f
C129 VN.n86 B 0.019057f
C130 VN.n87 B 0.03534f
C131 VN.n88 B 0.038176f
C132 VN.n89 B 0.015692f
C133 VN.n90 B 0.019057f
C134 VN.n91 B 0.019057f
C135 VN.n92 B 0.019057f
C136 VN.n93 B 0.03534f
C137 VN.n94 B 0.03534f
C138 VN.n95 B 0.020336f
C139 VN.n96 B 0.019057f
C140 VN.n97 B 0.019057f
C141 VN.n98 B 0.019057f
C142 VN.n99 B 0.03534f
C143 VN.n100 B 0.037875f
C144 VN.n101 B 0.01825f
C145 VN.n102 B 0.019057f
C146 VN.n103 B 0.019057f
C147 VN.n104 B 0.019057f
C148 VN.n105 B 0.03534f
C149 VN.n106 B 0.03534f
C150 VN.n107 B 0.022779f
C151 VN.n108 B 0.030753f
C152 VN.n109 B 1.27369f
C153 VTAIL.t1 B 0.158927f
C154 VTAIL.t8 B 0.158927f
C155 VTAIL.n0 B 1.28486f
C156 VTAIL.n1 B 0.726292f
C157 VTAIL.t13 B 1.63486f
C158 VTAIL.n2 B 0.8871f
C159 VTAIL.t11 B 0.158927f
C160 VTAIL.t16 B 0.158927f
C161 VTAIL.n3 B 1.28486f
C162 VTAIL.n4 B 0.924997f
C163 VTAIL.t17 B 0.158927f
C164 VTAIL.t14 B 0.158927f
C165 VTAIL.n5 B 1.28486f
C166 VTAIL.n6 B 2.21333f
C167 VTAIL.t6 B 0.158927f
C168 VTAIL.t4 B 0.158927f
C169 VTAIL.n7 B 1.28487f
C170 VTAIL.n8 B 2.21332f
C171 VTAIL.t7 B 0.158927f
C172 VTAIL.t2 B 0.158927f
C173 VTAIL.n9 B 1.28487f
C174 VTAIL.n10 B 0.924987f
C175 VTAIL.t0 B 1.63487f
C176 VTAIL.n11 B 0.887085f
C177 VTAIL.t10 B 0.158927f
C178 VTAIL.t18 B 0.158927f
C179 VTAIL.n12 B 1.28487f
C180 VTAIL.n13 B 0.803647f
C181 VTAIL.t9 B 0.158927f
C182 VTAIL.t12 B 0.158927f
C183 VTAIL.n14 B 1.28487f
C184 VTAIL.n15 B 0.924987f
C185 VTAIL.t15 B 1.63486f
C186 VTAIL.n16 B 1.96533f
C187 VTAIL.t3 B 1.63486f
C188 VTAIL.n17 B 1.96533f
C189 VTAIL.t5 B 0.158927f
C190 VTAIL.t19 B 0.158927f
C191 VTAIL.n18 B 1.28486f
C192 VTAIL.n19 B 0.670915f
C193 VDD1.t7 B 1.62131f
C194 VDD1.t0 B 0.146836f
C195 VDD1.t9 B 0.146836f
C196 VDD1.n0 B 1.25455f
C197 VDD1.n1 B 1.1618f
C198 VDD1.t8 B 1.6213f
C199 VDD1.t4 B 0.146836f
C200 VDD1.t2 B 0.146836f
C201 VDD1.n2 B 1.25454f
C202 VDD1.n3 B 1.15267f
C203 VDD1.t1 B 0.146836f
C204 VDD1.t5 B 0.146836f
C205 VDD1.n4 B 1.28216f
C206 VDD1.n5 B 3.60224f
C207 VDD1.t3 B 0.146836f
C208 VDD1.t6 B 0.146836f
C209 VDD1.n6 B 1.25454f
C210 VDD1.n7 B 3.51398f
C211 VP.t5 B 1.33747f
C212 VP.n0 B 0.562509f
C213 VP.n1 B 0.019552f
C214 VP.n2 B 0.035519f
C215 VP.n3 B 0.019552f
C216 VP.n4 B 0.033751f
C217 VP.n5 B 0.019552f
C218 VP.n6 B 0.037834f
C219 VP.n7 B 0.019552f
C220 VP.n8 B 0.036256f
C221 VP.n9 B 0.019552f
C222 VP.t7 B 1.33747f
C223 VP.n10 B 0.039166f
C224 VP.n11 B 0.019552f
C225 VP.n12 B 0.036256f
C226 VP.n13 B 0.019552f
C227 VP.t4 B 1.33747f
C228 VP.n14 B 0.038857f
C229 VP.n15 B 0.019552f
C230 VP.n16 B 0.036256f
C231 VP.t3 B 1.33747f
C232 VP.n17 B 0.562509f
C233 VP.n18 B 0.019552f
C234 VP.n19 B 0.035519f
C235 VP.n20 B 0.019552f
C236 VP.n21 B 0.033751f
C237 VP.n22 B 0.019552f
C238 VP.n23 B 0.037834f
C239 VP.n24 B 0.019552f
C240 VP.n25 B 0.036256f
C241 VP.n26 B 0.019552f
C242 VP.t9 B 1.33747f
C243 VP.n27 B 0.039166f
C244 VP.n28 B 0.019552f
C245 VP.n29 B 0.036256f
C246 VP.t8 B 1.60899f
C247 VP.n30 B 0.526018f
C248 VP.t0 B 1.33747f
C249 VP.n31 B 0.549504f
C250 VP.n32 B 0.020863f
C251 VP.n33 B 0.248194f
C252 VP.n34 B 0.019552f
C253 VP.n35 B 0.019552f
C254 VP.n36 B 0.036256f
C255 VP.n37 B 0.037834f
C256 VP.n38 B 0.016099f
C257 VP.n39 B 0.019552f
C258 VP.n40 B 0.019552f
C259 VP.n41 B 0.019552f
C260 VP.n42 B 0.036256f
C261 VP.n43 B 0.036256f
C262 VP.n44 B 0.50485f
C263 VP.n45 B 0.019552f
C264 VP.n46 B 0.019552f
C265 VP.n47 B 0.019552f
C266 VP.n48 B 0.036256f
C267 VP.n49 B 0.039166f
C268 VP.n50 B 0.016099f
C269 VP.n51 B 0.019552f
C270 VP.n52 B 0.019552f
C271 VP.n53 B 0.019552f
C272 VP.n54 B 0.036256f
C273 VP.n55 B 0.036256f
C274 VP.t6 B 1.33747f
C275 VP.n56 B 0.486492f
C276 VP.n57 B 0.020863f
C277 VP.n58 B 0.019552f
C278 VP.n59 B 0.019552f
C279 VP.n60 B 0.019552f
C280 VP.n61 B 0.036256f
C281 VP.n62 B 0.038857f
C282 VP.n63 B 0.018723f
C283 VP.n64 B 0.019552f
C284 VP.n65 B 0.019552f
C285 VP.n66 B 0.019552f
C286 VP.n67 B 0.036256f
C287 VP.n68 B 0.036256f
C288 VP.n69 B 0.023369f
C289 VP.n70 B 0.031551f
C290 VP.n71 B 1.299f
C291 VP.n72 B 1.3117f
C292 VP.t1 B 1.33747f
C293 VP.n73 B 0.562509f
C294 VP.n74 B 0.023369f
C295 VP.n75 B 0.031551f
C296 VP.n76 B 0.019552f
C297 VP.n77 B 0.019552f
C298 VP.n78 B 0.036256f
C299 VP.n79 B 0.035519f
C300 VP.n80 B 0.018723f
C301 VP.n81 B 0.019552f
C302 VP.n82 B 0.019552f
C303 VP.n83 B 0.019552f
C304 VP.n84 B 0.036256f
C305 VP.n85 B 0.033751f
C306 VP.n86 B 0.486492f
C307 VP.n87 B 0.020863f
C308 VP.n88 B 0.019552f
C309 VP.n89 B 0.019552f
C310 VP.n90 B 0.019552f
C311 VP.n91 B 0.036256f
C312 VP.n92 B 0.037834f
C313 VP.n93 B 0.016099f
C314 VP.n94 B 0.019552f
C315 VP.n95 B 0.019552f
C316 VP.n96 B 0.019552f
C317 VP.n97 B 0.036256f
C318 VP.n98 B 0.036256f
C319 VP.n99 B 0.50485f
C320 VP.n100 B 0.019552f
C321 VP.n101 B 0.019552f
C322 VP.n102 B 0.019552f
C323 VP.n103 B 0.036256f
C324 VP.n104 B 0.039166f
C325 VP.n105 B 0.016099f
C326 VP.n106 B 0.019552f
C327 VP.n107 B 0.019552f
C328 VP.n108 B 0.019552f
C329 VP.n109 B 0.036256f
C330 VP.n110 B 0.036256f
C331 VP.t2 B 1.33747f
C332 VP.n111 B 0.486492f
C333 VP.n112 B 0.020863f
C334 VP.n113 B 0.019552f
C335 VP.n114 B 0.019552f
C336 VP.n115 B 0.019552f
C337 VP.n116 B 0.036256f
C338 VP.n117 B 0.038857f
C339 VP.n118 B 0.018723f
C340 VP.n119 B 0.019552f
C341 VP.n120 B 0.019552f
C342 VP.n121 B 0.019552f
C343 VP.n122 B 0.036256f
C344 VP.n123 B 0.036256f
C345 VP.n124 B 0.023369f
C346 VP.n125 B 0.031551f
C347 VP.n126 B 0.056897f
.ends

