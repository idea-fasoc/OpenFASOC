* NGSPICE file created from diff_pair_sample_0373.ext - technology: sky130A

.subckt diff_pair_sample_0373 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t3 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X1 VDD2.t2 VN.t1 VTAIL.t18 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X2 VDD1.t9 VP.t0 VTAIL.t6 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=6.0177 ps=31.64 w=15.43 l=2.07
X3 VDD2.t1 VN.t2 VTAIL.t17 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=6.0177 pd=31.64 as=2.54595 ps=15.76 w=15.43 l=2.07
X4 VTAIL.t7 VP.t1 VDD1.t8 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X5 VTAIL.t3 VP.t2 VDD1.t7 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X6 VTAIL.t16 VN.t3 VDD2.t0 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X7 B.t11 B.t9 B.t10 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=6.0177 pd=31.64 as=0 ps=0 w=15.43 l=2.07
X8 VDD1.t6 VP.t3 VTAIL.t9 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X9 VDD2.t9 VN.t4 VTAIL.t15 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=6.0177 ps=31.64 w=15.43 l=2.07
X10 VTAIL.t14 VN.t5 VDD2.t8 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X11 B.t8 B.t6 B.t7 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=6.0177 pd=31.64 as=0 ps=0 w=15.43 l=2.07
X12 VTAIL.t5 VP.t4 VDD1.t5 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X13 VDD1.t4 VP.t5 VTAIL.t8 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=6.0177 ps=31.64 w=15.43 l=2.07
X14 VDD1.t3 VP.t6 VTAIL.t2 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X15 VDD2.t5 VN.t6 VTAIL.t13 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X16 VTAIL.t1 VP.t7 VDD1.t2 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X17 VDD1.t1 VP.t8 VTAIL.t4 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=6.0177 pd=31.64 as=2.54595 ps=15.76 w=15.43 l=2.07
X18 B.t5 B.t3 B.t4 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=6.0177 pd=31.64 as=0 ps=0 w=15.43 l=2.07
X19 VDD2.t4 VN.t7 VTAIL.t12 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=6.0177 ps=31.64 w=15.43 l=2.07
X20 VTAIL.t11 VN.t8 VDD2.t7 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=2.54595 pd=15.76 as=2.54595 ps=15.76 w=15.43 l=2.07
X21 B.t2 B.t0 B.t1 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=6.0177 pd=31.64 as=0 ps=0 w=15.43 l=2.07
X22 VDD2.t6 VN.t9 VTAIL.t10 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=6.0177 pd=31.64 as=2.54595 ps=15.76 w=15.43 l=2.07
X23 VDD1.t0 VP.t9 VTAIL.t0 w_n3850_n4054# sky130_fd_pr__pfet_01v8 ad=6.0177 pd=31.64 as=2.54595 ps=15.76 w=15.43 l=2.07
R0 VN.n8 VN.t9 212.583
R1 VN.n41 VN.t4 212.583
R2 VN.n16 VN.t1 179.644
R3 VN.n7 VN.t0 179.644
R4 VN.n23 VN.t8 179.644
R5 VN.n31 VN.t7 179.644
R6 VN.n49 VN.t6 179.644
R7 VN.n40 VN.t5 179.644
R8 VN.n56 VN.t3 179.644
R9 VN.n64 VN.t2 179.644
R10 VN.n63 VN.n33 161.3
R11 VN.n62 VN.n61 161.3
R12 VN.n60 VN.n34 161.3
R13 VN.n59 VN.n58 161.3
R14 VN.n57 VN.n35 161.3
R15 VN.n55 VN.n54 161.3
R16 VN.n53 VN.n36 161.3
R17 VN.n52 VN.n51 161.3
R18 VN.n50 VN.n37 161.3
R19 VN.n49 VN.n48 161.3
R20 VN.n47 VN.n38 161.3
R21 VN.n46 VN.n45 161.3
R22 VN.n44 VN.n39 161.3
R23 VN.n43 VN.n42 161.3
R24 VN.n30 VN.n0 161.3
R25 VN.n29 VN.n28 161.3
R26 VN.n27 VN.n1 161.3
R27 VN.n26 VN.n25 161.3
R28 VN.n24 VN.n2 161.3
R29 VN.n22 VN.n21 161.3
R30 VN.n20 VN.n3 161.3
R31 VN.n19 VN.n18 161.3
R32 VN.n17 VN.n4 161.3
R33 VN.n16 VN.n15 161.3
R34 VN.n14 VN.n5 161.3
R35 VN.n13 VN.n12 161.3
R36 VN.n11 VN.n6 161.3
R37 VN.n10 VN.n9 161.3
R38 VN.n32 VN.n31 96.0763
R39 VN.n65 VN.n64 96.0763
R40 VN.n12 VN.n11 56.5193
R41 VN.n18 VN.n3 56.5193
R42 VN.n45 VN.n44 56.5193
R43 VN.n51 VN.n36 56.5193
R44 VN VN.n65 53.0739
R45 VN.n8 VN.n7 51.1767
R46 VN.n41 VN.n40 51.1767
R47 VN.n29 VN.n1 50.2061
R48 VN.n62 VN.n34 50.2061
R49 VN.n25 VN.n1 30.7807
R50 VN.n58 VN.n34 30.7807
R51 VN.n11 VN.n10 24.4675
R52 VN.n12 VN.n5 24.4675
R53 VN.n16 VN.n5 24.4675
R54 VN.n17 VN.n16 24.4675
R55 VN.n18 VN.n17 24.4675
R56 VN.n22 VN.n3 24.4675
R57 VN.n25 VN.n24 24.4675
R58 VN.n30 VN.n29 24.4675
R59 VN.n44 VN.n43 24.4675
R60 VN.n51 VN.n50 24.4675
R61 VN.n50 VN.n49 24.4675
R62 VN.n49 VN.n38 24.4675
R63 VN.n45 VN.n38 24.4675
R64 VN.n58 VN.n57 24.4675
R65 VN.n55 VN.n36 24.4675
R66 VN.n63 VN.n62 24.4675
R67 VN.n10 VN.n7 19.5741
R68 VN.n23 VN.n22 19.5741
R69 VN.n43 VN.n40 19.5741
R70 VN.n56 VN.n55 19.5741
R71 VN.n31 VN.n30 14.6807
R72 VN.n64 VN.n63 14.6807
R73 VN.n42 VN.n41 9.46762
R74 VN.n9 VN.n8 9.46762
R75 VN.n24 VN.n23 4.8939
R76 VN.n57 VN.n56 4.8939
R77 VN.n65 VN.n33 0.278367
R78 VN.n32 VN.n0 0.278367
R79 VN.n61 VN.n33 0.189894
R80 VN.n61 VN.n60 0.189894
R81 VN.n60 VN.n59 0.189894
R82 VN.n59 VN.n35 0.189894
R83 VN.n54 VN.n35 0.189894
R84 VN.n54 VN.n53 0.189894
R85 VN.n53 VN.n52 0.189894
R86 VN.n52 VN.n37 0.189894
R87 VN.n48 VN.n37 0.189894
R88 VN.n48 VN.n47 0.189894
R89 VN.n47 VN.n46 0.189894
R90 VN.n46 VN.n39 0.189894
R91 VN.n42 VN.n39 0.189894
R92 VN.n9 VN.n6 0.189894
R93 VN.n13 VN.n6 0.189894
R94 VN.n14 VN.n13 0.189894
R95 VN.n15 VN.n14 0.189894
R96 VN.n15 VN.n4 0.189894
R97 VN.n19 VN.n4 0.189894
R98 VN.n20 VN.n19 0.189894
R99 VN.n21 VN.n20 0.189894
R100 VN.n21 VN.n2 0.189894
R101 VN.n26 VN.n2 0.189894
R102 VN.n27 VN.n26 0.189894
R103 VN.n28 VN.n27 0.189894
R104 VN.n28 VN.n0 0.189894
R105 VN VN.n32 0.153454
R106 VDD2.n169 VDD2.n89 756.745
R107 VDD2.n80 VDD2.n0 756.745
R108 VDD2.n170 VDD2.n169 585
R109 VDD2.n168 VDD2.n167 585
R110 VDD2.n93 VDD2.n92 585
R111 VDD2.n97 VDD2.n95 585
R112 VDD2.n162 VDD2.n161 585
R113 VDD2.n160 VDD2.n159 585
R114 VDD2.n99 VDD2.n98 585
R115 VDD2.n154 VDD2.n153 585
R116 VDD2.n152 VDD2.n151 585
R117 VDD2.n103 VDD2.n102 585
R118 VDD2.n146 VDD2.n145 585
R119 VDD2.n144 VDD2.n143 585
R120 VDD2.n107 VDD2.n106 585
R121 VDD2.n138 VDD2.n137 585
R122 VDD2.n136 VDD2.n135 585
R123 VDD2.n111 VDD2.n110 585
R124 VDD2.n130 VDD2.n129 585
R125 VDD2.n128 VDD2.n127 585
R126 VDD2.n115 VDD2.n114 585
R127 VDD2.n122 VDD2.n121 585
R128 VDD2.n120 VDD2.n119 585
R129 VDD2.n29 VDD2.n28 585
R130 VDD2.n31 VDD2.n30 585
R131 VDD2.n24 VDD2.n23 585
R132 VDD2.n37 VDD2.n36 585
R133 VDD2.n39 VDD2.n38 585
R134 VDD2.n20 VDD2.n19 585
R135 VDD2.n45 VDD2.n44 585
R136 VDD2.n47 VDD2.n46 585
R137 VDD2.n16 VDD2.n15 585
R138 VDD2.n53 VDD2.n52 585
R139 VDD2.n55 VDD2.n54 585
R140 VDD2.n12 VDD2.n11 585
R141 VDD2.n61 VDD2.n60 585
R142 VDD2.n63 VDD2.n62 585
R143 VDD2.n8 VDD2.n7 585
R144 VDD2.n70 VDD2.n69 585
R145 VDD2.n71 VDD2.n6 585
R146 VDD2.n73 VDD2.n72 585
R147 VDD2.n4 VDD2.n3 585
R148 VDD2.n79 VDD2.n78 585
R149 VDD2.n81 VDD2.n80 585
R150 VDD2.n118 VDD2.t1 327.466
R151 VDD2.n27 VDD2.t6 327.466
R152 VDD2.n169 VDD2.n168 171.744
R153 VDD2.n168 VDD2.n92 171.744
R154 VDD2.n97 VDD2.n92 171.744
R155 VDD2.n161 VDD2.n97 171.744
R156 VDD2.n161 VDD2.n160 171.744
R157 VDD2.n160 VDD2.n98 171.744
R158 VDD2.n153 VDD2.n98 171.744
R159 VDD2.n153 VDD2.n152 171.744
R160 VDD2.n152 VDD2.n102 171.744
R161 VDD2.n145 VDD2.n102 171.744
R162 VDD2.n145 VDD2.n144 171.744
R163 VDD2.n144 VDD2.n106 171.744
R164 VDD2.n137 VDD2.n106 171.744
R165 VDD2.n137 VDD2.n136 171.744
R166 VDD2.n136 VDD2.n110 171.744
R167 VDD2.n129 VDD2.n110 171.744
R168 VDD2.n129 VDD2.n128 171.744
R169 VDD2.n128 VDD2.n114 171.744
R170 VDD2.n121 VDD2.n114 171.744
R171 VDD2.n121 VDD2.n120 171.744
R172 VDD2.n30 VDD2.n29 171.744
R173 VDD2.n30 VDD2.n23 171.744
R174 VDD2.n37 VDD2.n23 171.744
R175 VDD2.n38 VDD2.n37 171.744
R176 VDD2.n38 VDD2.n19 171.744
R177 VDD2.n45 VDD2.n19 171.744
R178 VDD2.n46 VDD2.n45 171.744
R179 VDD2.n46 VDD2.n15 171.744
R180 VDD2.n53 VDD2.n15 171.744
R181 VDD2.n54 VDD2.n53 171.744
R182 VDD2.n54 VDD2.n11 171.744
R183 VDD2.n61 VDD2.n11 171.744
R184 VDD2.n62 VDD2.n61 171.744
R185 VDD2.n62 VDD2.n7 171.744
R186 VDD2.n70 VDD2.n7 171.744
R187 VDD2.n71 VDD2.n70 171.744
R188 VDD2.n72 VDD2.n71 171.744
R189 VDD2.n72 VDD2.n3 171.744
R190 VDD2.n79 VDD2.n3 171.744
R191 VDD2.n80 VDD2.n79 171.744
R192 VDD2.n120 VDD2.t1 85.8723
R193 VDD2.n29 VDD2.t6 85.8723
R194 VDD2.n88 VDD2.n87 73.1119
R195 VDD2 VDD2.n177 73.1091
R196 VDD2.n176 VDD2.n175 71.6157
R197 VDD2.n86 VDD2.n85 71.6155
R198 VDD2.n86 VDD2.n84 52.2907
R199 VDD2.n174 VDD2.n173 50.2217
R200 VDD2.n174 VDD2.n88 46.8446
R201 VDD2.n119 VDD2.n118 16.3895
R202 VDD2.n28 VDD2.n27 16.3895
R203 VDD2.n95 VDD2.n93 13.1884
R204 VDD2.n73 VDD2.n4 13.1884
R205 VDD2.n167 VDD2.n166 12.8005
R206 VDD2.n163 VDD2.n162 12.8005
R207 VDD2.n122 VDD2.n117 12.8005
R208 VDD2.n31 VDD2.n26 12.8005
R209 VDD2.n74 VDD2.n6 12.8005
R210 VDD2.n78 VDD2.n77 12.8005
R211 VDD2.n170 VDD2.n91 12.0247
R212 VDD2.n159 VDD2.n96 12.0247
R213 VDD2.n123 VDD2.n115 12.0247
R214 VDD2.n32 VDD2.n24 12.0247
R215 VDD2.n69 VDD2.n68 12.0247
R216 VDD2.n81 VDD2.n2 12.0247
R217 VDD2.n171 VDD2.n89 11.249
R218 VDD2.n158 VDD2.n99 11.249
R219 VDD2.n127 VDD2.n126 11.249
R220 VDD2.n36 VDD2.n35 11.249
R221 VDD2.n67 VDD2.n8 11.249
R222 VDD2.n82 VDD2.n0 11.249
R223 VDD2.n155 VDD2.n154 10.4732
R224 VDD2.n130 VDD2.n113 10.4732
R225 VDD2.n39 VDD2.n22 10.4732
R226 VDD2.n64 VDD2.n63 10.4732
R227 VDD2.n151 VDD2.n101 9.69747
R228 VDD2.n131 VDD2.n111 9.69747
R229 VDD2.n40 VDD2.n20 9.69747
R230 VDD2.n60 VDD2.n10 9.69747
R231 VDD2.n173 VDD2.n172 9.45567
R232 VDD2.n84 VDD2.n83 9.45567
R233 VDD2.n105 VDD2.n104 9.3005
R234 VDD2.n148 VDD2.n147 9.3005
R235 VDD2.n150 VDD2.n149 9.3005
R236 VDD2.n101 VDD2.n100 9.3005
R237 VDD2.n156 VDD2.n155 9.3005
R238 VDD2.n158 VDD2.n157 9.3005
R239 VDD2.n96 VDD2.n94 9.3005
R240 VDD2.n164 VDD2.n163 9.3005
R241 VDD2.n172 VDD2.n171 9.3005
R242 VDD2.n91 VDD2.n90 9.3005
R243 VDD2.n166 VDD2.n165 9.3005
R244 VDD2.n142 VDD2.n141 9.3005
R245 VDD2.n140 VDD2.n139 9.3005
R246 VDD2.n109 VDD2.n108 9.3005
R247 VDD2.n134 VDD2.n133 9.3005
R248 VDD2.n132 VDD2.n131 9.3005
R249 VDD2.n113 VDD2.n112 9.3005
R250 VDD2.n126 VDD2.n125 9.3005
R251 VDD2.n124 VDD2.n123 9.3005
R252 VDD2.n117 VDD2.n116 9.3005
R253 VDD2.n83 VDD2.n82 9.3005
R254 VDD2.n2 VDD2.n1 9.3005
R255 VDD2.n77 VDD2.n76 9.3005
R256 VDD2.n49 VDD2.n48 9.3005
R257 VDD2.n18 VDD2.n17 9.3005
R258 VDD2.n43 VDD2.n42 9.3005
R259 VDD2.n41 VDD2.n40 9.3005
R260 VDD2.n22 VDD2.n21 9.3005
R261 VDD2.n35 VDD2.n34 9.3005
R262 VDD2.n33 VDD2.n32 9.3005
R263 VDD2.n26 VDD2.n25 9.3005
R264 VDD2.n51 VDD2.n50 9.3005
R265 VDD2.n14 VDD2.n13 9.3005
R266 VDD2.n57 VDD2.n56 9.3005
R267 VDD2.n59 VDD2.n58 9.3005
R268 VDD2.n10 VDD2.n9 9.3005
R269 VDD2.n65 VDD2.n64 9.3005
R270 VDD2.n67 VDD2.n66 9.3005
R271 VDD2.n68 VDD2.n5 9.3005
R272 VDD2.n75 VDD2.n74 9.3005
R273 VDD2.n150 VDD2.n103 8.92171
R274 VDD2.n135 VDD2.n134 8.92171
R275 VDD2.n44 VDD2.n43 8.92171
R276 VDD2.n59 VDD2.n12 8.92171
R277 VDD2.n147 VDD2.n146 8.14595
R278 VDD2.n138 VDD2.n109 8.14595
R279 VDD2.n47 VDD2.n18 8.14595
R280 VDD2.n56 VDD2.n55 8.14595
R281 VDD2.n143 VDD2.n105 7.3702
R282 VDD2.n139 VDD2.n107 7.3702
R283 VDD2.n48 VDD2.n16 7.3702
R284 VDD2.n52 VDD2.n14 7.3702
R285 VDD2.n143 VDD2.n142 6.59444
R286 VDD2.n142 VDD2.n107 6.59444
R287 VDD2.n51 VDD2.n16 6.59444
R288 VDD2.n52 VDD2.n51 6.59444
R289 VDD2.n146 VDD2.n105 5.81868
R290 VDD2.n139 VDD2.n138 5.81868
R291 VDD2.n48 VDD2.n47 5.81868
R292 VDD2.n55 VDD2.n14 5.81868
R293 VDD2.n147 VDD2.n103 5.04292
R294 VDD2.n135 VDD2.n109 5.04292
R295 VDD2.n44 VDD2.n18 5.04292
R296 VDD2.n56 VDD2.n12 5.04292
R297 VDD2.n151 VDD2.n150 4.26717
R298 VDD2.n134 VDD2.n111 4.26717
R299 VDD2.n43 VDD2.n20 4.26717
R300 VDD2.n60 VDD2.n59 4.26717
R301 VDD2.n118 VDD2.n116 3.70982
R302 VDD2.n27 VDD2.n25 3.70982
R303 VDD2.n154 VDD2.n101 3.49141
R304 VDD2.n131 VDD2.n130 3.49141
R305 VDD2.n40 VDD2.n39 3.49141
R306 VDD2.n63 VDD2.n10 3.49141
R307 VDD2.n173 VDD2.n89 2.71565
R308 VDD2.n155 VDD2.n99 2.71565
R309 VDD2.n127 VDD2.n113 2.71565
R310 VDD2.n36 VDD2.n22 2.71565
R311 VDD2.n64 VDD2.n8 2.71565
R312 VDD2.n84 VDD2.n0 2.71565
R313 VDD2.n177 VDD2.t8 2.10711
R314 VDD2.n177 VDD2.t9 2.10711
R315 VDD2.n175 VDD2.t0 2.10711
R316 VDD2.n175 VDD2.t5 2.10711
R317 VDD2.n87 VDD2.t7 2.10711
R318 VDD2.n87 VDD2.t4 2.10711
R319 VDD2.n85 VDD2.t3 2.10711
R320 VDD2.n85 VDD2.t2 2.10711
R321 VDD2.n176 VDD2.n174 2.06947
R322 VDD2.n171 VDD2.n170 1.93989
R323 VDD2.n159 VDD2.n158 1.93989
R324 VDD2.n126 VDD2.n115 1.93989
R325 VDD2.n35 VDD2.n24 1.93989
R326 VDD2.n69 VDD2.n67 1.93989
R327 VDD2.n82 VDD2.n81 1.93989
R328 VDD2.n167 VDD2.n91 1.16414
R329 VDD2.n162 VDD2.n96 1.16414
R330 VDD2.n123 VDD2.n122 1.16414
R331 VDD2.n32 VDD2.n31 1.16414
R332 VDD2.n68 VDD2.n6 1.16414
R333 VDD2.n78 VDD2.n2 1.16414
R334 VDD2 VDD2.n176 0.575931
R335 VDD2.n88 VDD2.n86 0.462395
R336 VDD2.n166 VDD2.n93 0.388379
R337 VDD2.n163 VDD2.n95 0.388379
R338 VDD2.n119 VDD2.n117 0.388379
R339 VDD2.n28 VDD2.n26 0.388379
R340 VDD2.n74 VDD2.n73 0.388379
R341 VDD2.n77 VDD2.n4 0.388379
R342 VDD2.n172 VDD2.n90 0.155672
R343 VDD2.n165 VDD2.n90 0.155672
R344 VDD2.n165 VDD2.n164 0.155672
R345 VDD2.n164 VDD2.n94 0.155672
R346 VDD2.n157 VDD2.n94 0.155672
R347 VDD2.n157 VDD2.n156 0.155672
R348 VDD2.n156 VDD2.n100 0.155672
R349 VDD2.n149 VDD2.n100 0.155672
R350 VDD2.n149 VDD2.n148 0.155672
R351 VDD2.n148 VDD2.n104 0.155672
R352 VDD2.n141 VDD2.n104 0.155672
R353 VDD2.n141 VDD2.n140 0.155672
R354 VDD2.n140 VDD2.n108 0.155672
R355 VDD2.n133 VDD2.n108 0.155672
R356 VDD2.n133 VDD2.n132 0.155672
R357 VDD2.n132 VDD2.n112 0.155672
R358 VDD2.n125 VDD2.n112 0.155672
R359 VDD2.n125 VDD2.n124 0.155672
R360 VDD2.n124 VDD2.n116 0.155672
R361 VDD2.n33 VDD2.n25 0.155672
R362 VDD2.n34 VDD2.n33 0.155672
R363 VDD2.n34 VDD2.n21 0.155672
R364 VDD2.n41 VDD2.n21 0.155672
R365 VDD2.n42 VDD2.n41 0.155672
R366 VDD2.n42 VDD2.n17 0.155672
R367 VDD2.n49 VDD2.n17 0.155672
R368 VDD2.n50 VDD2.n49 0.155672
R369 VDD2.n50 VDD2.n13 0.155672
R370 VDD2.n57 VDD2.n13 0.155672
R371 VDD2.n58 VDD2.n57 0.155672
R372 VDD2.n58 VDD2.n9 0.155672
R373 VDD2.n65 VDD2.n9 0.155672
R374 VDD2.n66 VDD2.n65 0.155672
R375 VDD2.n66 VDD2.n5 0.155672
R376 VDD2.n75 VDD2.n5 0.155672
R377 VDD2.n76 VDD2.n75 0.155672
R378 VDD2.n76 VDD2.n1 0.155672
R379 VDD2.n83 VDD2.n1 0.155672
R380 VTAIL.n352 VTAIL.n272 756.745
R381 VTAIL.n82 VTAIL.n2 756.745
R382 VTAIL.n266 VTAIL.n186 756.745
R383 VTAIL.n176 VTAIL.n96 756.745
R384 VTAIL.n301 VTAIL.n300 585
R385 VTAIL.n303 VTAIL.n302 585
R386 VTAIL.n296 VTAIL.n295 585
R387 VTAIL.n309 VTAIL.n308 585
R388 VTAIL.n311 VTAIL.n310 585
R389 VTAIL.n292 VTAIL.n291 585
R390 VTAIL.n317 VTAIL.n316 585
R391 VTAIL.n319 VTAIL.n318 585
R392 VTAIL.n288 VTAIL.n287 585
R393 VTAIL.n325 VTAIL.n324 585
R394 VTAIL.n327 VTAIL.n326 585
R395 VTAIL.n284 VTAIL.n283 585
R396 VTAIL.n333 VTAIL.n332 585
R397 VTAIL.n335 VTAIL.n334 585
R398 VTAIL.n280 VTAIL.n279 585
R399 VTAIL.n342 VTAIL.n341 585
R400 VTAIL.n343 VTAIL.n278 585
R401 VTAIL.n345 VTAIL.n344 585
R402 VTAIL.n276 VTAIL.n275 585
R403 VTAIL.n351 VTAIL.n350 585
R404 VTAIL.n353 VTAIL.n352 585
R405 VTAIL.n31 VTAIL.n30 585
R406 VTAIL.n33 VTAIL.n32 585
R407 VTAIL.n26 VTAIL.n25 585
R408 VTAIL.n39 VTAIL.n38 585
R409 VTAIL.n41 VTAIL.n40 585
R410 VTAIL.n22 VTAIL.n21 585
R411 VTAIL.n47 VTAIL.n46 585
R412 VTAIL.n49 VTAIL.n48 585
R413 VTAIL.n18 VTAIL.n17 585
R414 VTAIL.n55 VTAIL.n54 585
R415 VTAIL.n57 VTAIL.n56 585
R416 VTAIL.n14 VTAIL.n13 585
R417 VTAIL.n63 VTAIL.n62 585
R418 VTAIL.n65 VTAIL.n64 585
R419 VTAIL.n10 VTAIL.n9 585
R420 VTAIL.n72 VTAIL.n71 585
R421 VTAIL.n73 VTAIL.n8 585
R422 VTAIL.n75 VTAIL.n74 585
R423 VTAIL.n6 VTAIL.n5 585
R424 VTAIL.n81 VTAIL.n80 585
R425 VTAIL.n83 VTAIL.n82 585
R426 VTAIL.n267 VTAIL.n266 585
R427 VTAIL.n265 VTAIL.n264 585
R428 VTAIL.n190 VTAIL.n189 585
R429 VTAIL.n194 VTAIL.n192 585
R430 VTAIL.n259 VTAIL.n258 585
R431 VTAIL.n257 VTAIL.n256 585
R432 VTAIL.n196 VTAIL.n195 585
R433 VTAIL.n251 VTAIL.n250 585
R434 VTAIL.n249 VTAIL.n248 585
R435 VTAIL.n200 VTAIL.n199 585
R436 VTAIL.n243 VTAIL.n242 585
R437 VTAIL.n241 VTAIL.n240 585
R438 VTAIL.n204 VTAIL.n203 585
R439 VTAIL.n235 VTAIL.n234 585
R440 VTAIL.n233 VTAIL.n232 585
R441 VTAIL.n208 VTAIL.n207 585
R442 VTAIL.n227 VTAIL.n226 585
R443 VTAIL.n225 VTAIL.n224 585
R444 VTAIL.n212 VTAIL.n211 585
R445 VTAIL.n219 VTAIL.n218 585
R446 VTAIL.n217 VTAIL.n216 585
R447 VTAIL.n177 VTAIL.n176 585
R448 VTAIL.n175 VTAIL.n174 585
R449 VTAIL.n100 VTAIL.n99 585
R450 VTAIL.n104 VTAIL.n102 585
R451 VTAIL.n169 VTAIL.n168 585
R452 VTAIL.n167 VTAIL.n166 585
R453 VTAIL.n106 VTAIL.n105 585
R454 VTAIL.n161 VTAIL.n160 585
R455 VTAIL.n159 VTAIL.n158 585
R456 VTAIL.n110 VTAIL.n109 585
R457 VTAIL.n153 VTAIL.n152 585
R458 VTAIL.n151 VTAIL.n150 585
R459 VTAIL.n114 VTAIL.n113 585
R460 VTAIL.n145 VTAIL.n144 585
R461 VTAIL.n143 VTAIL.n142 585
R462 VTAIL.n118 VTAIL.n117 585
R463 VTAIL.n137 VTAIL.n136 585
R464 VTAIL.n135 VTAIL.n134 585
R465 VTAIL.n122 VTAIL.n121 585
R466 VTAIL.n129 VTAIL.n128 585
R467 VTAIL.n127 VTAIL.n126 585
R468 VTAIL.n299 VTAIL.t12 327.466
R469 VTAIL.n29 VTAIL.t8 327.466
R470 VTAIL.n215 VTAIL.t6 327.466
R471 VTAIL.n125 VTAIL.t15 327.466
R472 VTAIL.n302 VTAIL.n301 171.744
R473 VTAIL.n302 VTAIL.n295 171.744
R474 VTAIL.n309 VTAIL.n295 171.744
R475 VTAIL.n310 VTAIL.n309 171.744
R476 VTAIL.n310 VTAIL.n291 171.744
R477 VTAIL.n317 VTAIL.n291 171.744
R478 VTAIL.n318 VTAIL.n317 171.744
R479 VTAIL.n318 VTAIL.n287 171.744
R480 VTAIL.n325 VTAIL.n287 171.744
R481 VTAIL.n326 VTAIL.n325 171.744
R482 VTAIL.n326 VTAIL.n283 171.744
R483 VTAIL.n333 VTAIL.n283 171.744
R484 VTAIL.n334 VTAIL.n333 171.744
R485 VTAIL.n334 VTAIL.n279 171.744
R486 VTAIL.n342 VTAIL.n279 171.744
R487 VTAIL.n343 VTAIL.n342 171.744
R488 VTAIL.n344 VTAIL.n343 171.744
R489 VTAIL.n344 VTAIL.n275 171.744
R490 VTAIL.n351 VTAIL.n275 171.744
R491 VTAIL.n352 VTAIL.n351 171.744
R492 VTAIL.n32 VTAIL.n31 171.744
R493 VTAIL.n32 VTAIL.n25 171.744
R494 VTAIL.n39 VTAIL.n25 171.744
R495 VTAIL.n40 VTAIL.n39 171.744
R496 VTAIL.n40 VTAIL.n21 171.744
R497 VTAIL.n47 VTAIL.n21 171.744
R498 VTAIL.n48 VTAIL.n47 171.744
R499 VTAIL.n48 VTAIL.n17 171.744
R500 VTAIL.n55 VTAIL.n17 171.744
R501 VTAIL.n56 VTAIL.n55 171.744
R502 VTAIL.n56 VTAIL.n13 171.744
R503 VTAIL.n63 VTAIL.n13 171.744
R504 VTAIL.n64 VTAIL.n63 171.744
R505 VTAIL.n64 VTAIL.n9 171.744
R506 VTAIL.n72 VTAIL.n9 171.744
R507 VTAIL.n73 VTAIL.n72 171.744
R508 VTAIL.n74 VTAIL.n73 171.744
R509 VTAIL.n74 VTAIL.n5 171.744
R510 VTAIL.n81 VTAIL.n5 171.744
R511 VTAIL.n82 VTAIL.n81 171.744
R512 VTAIL.n266 VTAIL.n265 171.744
R513 VTAIL.n265 VTAIL.n189 171.744
R514 VTAIL.n194 VTAIL.n189 171.744
R515 VTAIL.n258 VTAIL.n194 171.744
R516 VTAIL.n258 VTAIL.n257 171.744
R517 VTAIL.n257 VTAIL.n195 171.744
R518 VTAIL.n250 VTAIL.n195 171.744
R519 VTAIL.n250 VTAIL.n249 171.744
R520 VTAIL.n249 VTAIL.n199 171.744
R521 VTAIL.n242 VTAIL.n199 171.744
R522 VTAIL.n242 VTAIL.n241 171.744
R523 VTAIL.n241 VTAIL.n203 171.744
R524 VTAIL.n234 VTAIL.n203 171.744
R525 VTAIL.n234 VTAIL.n233 171.744
R526 VTAIL.n233 VTAIL.n207 171.744
R527 VTAIL.n226 VTAIL.n207 171.744
R528 VTAIL.n226 VTAIL.n225 171.744
R529 VTAIL.n225 VTAIL.n211 171.744
R530 VTAIL.n218 VTAIL.n211 171.744
R531 VTAIL.n218 VTAIL.n217 171.744
R532 VTAIL.n176 VTAIL.n175 171.744
R533 VTAIL.n175 VTAIL.n99 171.744
R534 VTAIL.n104 VTAIL.n99 171.744
R535 VTAIL.n168 VTAIL.n104 171.744
R536 VTAIL.n168 VTAIL.n167 171.744
R537 VTAIL.n167 VTAIL.n105 171.744
R538 VTAIL.n160 VTAIL.n105 171.744
R539 VTAIL.n160 VTAIL.n159 171.744
R540 VTAIL.n159 VTAIL.n109 171.744
R541 VTAIL.n152 VTAIL.n109 171.744
R542 VTAIL.n152 VTAIL.n151 171.744
R543 VTAIL.n151 VTAIL.n113 171.744
R544 VTAIL.n144 VTAIL.n113 171.744
R545 VTAIL.n144 VTAIL.n143 171.744
R546 VTAIL.n143 VTAIL.n117 171.744
R547 VTAIL.n136 VTAIL.n117 171.744
R548 VTAIL.n136 VTAIL.n135 171.744
R549 VTAIL.n135 VTAIL.n121 171.744
R550 VTAIL.n128 VTAIL.n121 171.744
R551 VTAIL.n128 VTAIL.n127 171.744
R552 VTAIL.n301 VTAIL.t12 85.8723
R553 VTAIL.n31 VTAIL.t8 85.8723
R554 VTAIL.n217 VTAIL.t6 85.8723
R555 VTAIL.n127 VTAIL.t15 85.8723
R556 VTAIL.n185 VTAIL.n184 54.9369
R557 VTAIL.n183 VTAIL.n182 54.9369
R558 VTAIL.n95 VTAIL.n94 54.9369
R559 VTAIL.n93 VTAIL.n92 54.9369
R560 VTAIL.n359 VTAIL.n358 54.9367
R561 VTAIL.n1 VTAIL.n0 54.9367
R562 VTAIL.n89 VTAIL.n88 54.9367
R563 VTAIL.n91 VTAIL.n90 54.9367
R564 VTAIL.n357 VTAIL.n356 33.5429
R565 VTAIL.n87 VTAIL.n86 33.5429
R566 VTAIL.n271 VTAIL.n270 33.5429
R567 VTAIL.n181 VTAIL.n180 33.5429
R568 VTAIL.n93 VTAIL.n91 29.8065
R569 VTAIL.n357 VTAIL.n271 27.7376
R570 VTAIL.n300 VTAIL.n299 16.3895
R571 VTAIL.n30 VTAIL.n29 16.3895
R572 VTAIL.n216 VTAIL.n215 16.3895
R573 VTAIL.n126 VTAIL.n125 16.3895
R574 VTAIL.n345 VTAIL.n276 13.1884
R575 VTAIL.n75 VTAIL.n6 13.1884
R576 VTAIL.n192 VTAIL.n190 13.1884
R577 VTAIL.n102 VTAIL.n100 13.1884
R578 VTAIL.n303 VTAIL.n298 12.8005
R579 VTAIL.n346 VTAIL.n278 12.8005
R580 VTAIL.n350 VTAIL.n349 12.8005
R581 VTAIL.n33 VTAIL.n28 12.8005
R582 VTAIL.n76 VTAIL.n8 12.8005
R583 VTAIL.n80 VTAIL.n79 12.8005
R584 VTAIL.n264 VTAIL.n263 12.8005
R585 VTAIL.n260 VTAIL.n259 12.8005
R586 VTAIL.n219 VTAIL.n214 12.8005
R587 VTAIL.n174 VTAIL.n173 12.8005
R588 VTAIL.n170 VTAIL.n169 12.8005
R589 VTAIL.n129 VTAIL.n124 12.8005
R590 VTAIL.n304 VTAIL.n296 12.0247
R591 VTAIL.n341 VTAIL.n340 12.0247
R592 VTAIL.n353 VTAIL.n274 12.0247
R593 VTAIL.n34 VTAIL.n26 12.0247
R594 VTAIL.n71 VTAIL.n70 12.0247
R595 VTAIL.n83 VTAIL.n4 12.0247
R596 VTAIL.n267 VTAIL.n188 12.0247
R597 VTAIL.n256 VTAIL.n193 12.0247
R598 VTAIL.n220 VTAIL.n212 12.0247
R599 VTAIL.n177 VTAIL.n98 12.0247
R600 VTAIL.n166 VTAIL.n103 12.0247
R601 VTAIL.n130 VTAIL.n122 12.0247
R602 VTAIL.n308 VTAIL.n307 11.249
R603 VTAIL.n339 VTAIL.n280 11.249
R604 VTAIL.n354 VTAIL.n272 11.249
R605 VTAIL.n38 VTAIL.n37 11.249
R606 VTAIL.n69 VTAIL.n10 11.249
R607 VTAIL.n84 VTAIL.n2 11.249
R608 VTAIL.n268 VTAIL.n186 11.249
R609 VTAIL.n255 VTAIL.n196 11.249
R610 VTAIL.n224 VTAIL.n223 11.249
R611 VTAIL.n178 VTAIL.n96 11.249
R612 VTAIL.n165 VTAIL.n106 11.249
R613 VTAIL.n134 VTAIL.n133 11.249
R614 VTAIL.n311 VTAIL.n294 10.4732
R615 VTAIL.n336 VTAIL.n335 10.4732
R616 VTAIL.n41 VTAIL.n24 10.4732
R617 VTAIL.n66 VTAIL.n65 10.4732
R618 VTAIL.n252 VTAIL.n251 10.4732
R619 VTAIL.n227 VTAIL.n210 10.4732
R620 VTAIL.n162 VTAIL.n161 10.4732
R621 VTAIL.n137 VTAIL.n120 10.4732
R622 VTAIL.n312 VTAIL.n292 9.69747
R623 VTAIL.n332 VTAIL.n282 9.69747
R624 VTAIL.n42 VTAIL.n22 9.69747
R625 VTAIL.n62 VTAIL.n12 9.69747
R626 VTAIL.n248 VTAIL.n198 9.69747
R627 VTAIL.n228 VTAIL.n208 9.69747
R628 VTAIL.n158 VTAIL.n108 9.69747
R629 VTAIL.n138 VTAIL.n118 9.69747
R630 VTAIL.n356 VTAIL.n355 9.45567
R631 VTAIL.n86 VTAIL.n85 9.45567
R632 VTAIL.n270 VTAIL.n269 9.45567
R633 VTAIL.n180 VTAIL.n179 9.45567
R634 VTAIL.n355 VTAIL.n354 9.3005
R635 VTAIL.n274 VTAIL.n273 9.3005
R636 VTAIL.n349 VTAIL.n348 9.3005
R637 VTAIL.n321 VTAIL.n320 9.3005
R638 VTAIL.n290 VTAIL.n289 9.3005
R639 VTAIL.n315 VTAIL.n314 9.3005
R640 VTAIL.n313 VTAIL.n312 9.3005
R641 VTAIL.n294 VTAIL.n293 9.3005
R642 VTAIL.n307 VTAIL.n306 9.3005
R643 VTAIL.n305 VTAIL.n304 9.3005
R644 VTAIL.n298 VTAIL.n297 9.3005
R645 VTAIL.n323 VTAIL.n322 9.3005
R646 VTAIL.n286 VTAIL.n285 9.3005
R647 VTAIL.n329 VTAIL.n328 9.3005
R648 VTAIL.n331 VTAIL.n330 9.3005
R649 VTAIL.n282 VTAIL.n281 9.3005
R650 VTAIL.n337 VTAIL.n336 9.3005
R651 VTAIL.n339 VTAIL.n338 9.3005
R652 VTAIL.n340 VTAIL.n277 9.3005
R653 VTAIL.n347 VTAIL.n346 9.3005
R654 VTAIL.n85 VTAIL.n84 9.3005
R655 VTAIL.n4 VTAIL.n3 9.3005
R656 VTAIL.n79 VTAIL.n78 9.3005
R657 VTAIL.n51 VTAIL.n50 9.3005
R658 VTAIL.n20 VTAIL.n19 9.3005
R659 VTAIL.n45 VTAIL.n44 9.3005
R660 VTAIL.n43 VTAIL.n42 9.3005
R661 VTAIL.n24 VTAIL.n23 9.3005
R662 VTAIL.n37 VTAIL.n36 9.3005
R663 VTAIL.n35 VTAIL.n34 9.3005
R664 VTAIL.n28 VTAIL.n27 9.3005
R665 VTAIL.n53 VTAIL.n52 9.3005
R666 VTAIL.n16 VTAIL.n15 9.3005
R667 VTAIL.n59 VTAIL.n58 9.3005
R668 VTAIL.n61 VTAIL.n60 9.3005
R669 VTAIL.n12 VTAIL.n11 9.3005
R670 VTAIL.n67 VTAIL.n66 9.3005
R671 VTAIL.n69 VTAIL.n68 9.3005
R672 VTAIL.n70 VTAIL.n7 9.3005
R673 VTAIL.n77 VTAIL.n76 9.3005
R674 VTAIL.n202 VTAIL.n201 9.3005
R675 VTAIL.n245 VTAIL.n244 9.3005
R676 VTAIL.n247 VTAIL.n246 9.3005
R677 VTAIL.n198 VTAIL.n197 9.3005
R678 VTAIL.n253 VTAIL.n252 9.3005
R679 VTAIL.n255 VTAIL.n254 9.3005
R680 VTAIL.n193 VTAIL.n191 9.3005
R681 VTAIL.n261 VTAIL.n260 9.3005
R682 VTAIL.n269 VTAIL.n268 9.3005
R683 VTAIL.n188 VTAIL.n187 9.3005
R684 VTAIL.n263 VTAIL.n262 9.3005
R685 VTAIL.n239 VTAIL.n238 9.3005
R686 VTAIL.n237 VTAIL.n236 9.3005
R687 VTAIL.n206 VTAIL.n205 9.3005
R688 VTAIL.n231 VTAIL.n230 9.3005
R689 VTAIL.n229 VTAIL.n228 9.3005
R690 VTAIL.n210 VTAIL.n209 9.3005
R691 VTAIL.n223 VTAIL.n222 9.3005
R692 VTAIL.n221 VTAIL.n220 9.3005
R693 VTAIL.n214 VTAIL.n213 9.3005
R694 VTAIL.n112 VTAIL.n111 9.3005
R695 VTAIL.n155 VTAIL.n154 9.3005
R696 VTAIL.n157 VTAIL.n156 9.3005
R697 VTAIL.n108 VTAIL.n107 9.3005
R698 VTAIL.n163 VTAIL.n162 9.3005
R699 VTAIL.n165 VTAIL.n164 9.3005
R700 VTAIL.n103 VTAIL.n101 9.3005
R701 VTAIL.n171 VTAIL.n170 9.3005
R702 VTAIL.n179 VTAIL.n178 9.3005
R703 VTAIL.n98 VTAIL.n97 9.3005
R704 VTAIL.n173 VTAIL.n172 9.3005
R705 VTAIL.n149 VTAIL.n148 9.3005
R706 VTAIL.n147 VTAIL.n146 9.3005
R707 VTAIL.n116 VTAIL.n115 9.3005
R708 VTAIL.n141 VTAIL.n140 9.3005
R709 VTAIL.n139 VTAIL.n138 9.3005
R710 VTAIL.n120 VTAIL.n119 9.3005
R711 VTAIL.n133 VTAIL.n132 9.3005
R712 VTAIL.n131 VTAIL.n130 9.3005
R713 VTAIL.n124 VTAIL.n123 9.3005
R714 VTAIL.n316 VTAIL.n315 8.92171
R715 VTAIL.n331 VTAIL.n284 8.92171
R716 VTAIL.n46 VTAIL.n45 8.92171
R717 VTAIL.n61 VTAIL.n14 8.92171
R718 VTAIL.n247 VTAIL.n200 8.92171
R719 VTAIL.n232 VTAIL.n231 8.92171
R720 VTAIL.n157 VTAIL.n110 8.92171
R721 VTAIL.n142 VTAIL.n141 8.92171
R722 VTAIL.n319 VTAIL.n290 8.14595
R723 VTAIL.n328 VTAIL.n327 8.14595
R724 VTAIL.n49 VTAIL.n20 8.14595
R725 VTAIL.n58 VTAIL.n57 8.14595
R726 VTAIL.n244 VTAIL.n243 8.14595
R727 VTAIL.n235 VTAIL.n206 8.14595
R728 VTAIL.n154 VTAIL.n153 8.14595
R729 VTAIL.n145 VTAIL.n116 8.14595
R730 VTAIL.n320 VTAIL.n288 7.3702
R731 VTAIL.n324 VTAIL.n286 7.3702
R732 VTAIL.n50 VTAIL.n18 7.3702
R733 VTAIL.n54 VTAIL.n16 7.3702
R734 VTAIL.n240 VTAIL.n202 7.3702
R735 VTAIL.n236 VTAIL.n204 7.3702
R736 VTAIL.n150 VTAIL.n112 7.3702
R737 VTAIL.n146 VTAIL.n114 7.3702
R738 VTAIL.n323 VTAIL.n288 6.59444
R739 VTAIL.n324 VTAIL.n323 6.59444
R740 VTAIL.n53 VTAIL.n18 6.59444
R741 VTAIL.n54 VTAIL.n53 6.59444
R742 VTAIL.n240 VTAIL.n239 6.59444
R743 VTAIL.n239 VTAIL.n204 6.59444
R744 VTAIL.n150 VTAIL.n149 6.59444
R745 VTAIL.n149 VTAIL.n114 6.59444
R746 VTAIL.n320 VTAIL.n319 5.81868
R747 VTAIL.n327 VTAIL.n286 5.81868
R748 VTAIL.n50 VTAIL.n49 5.81868
R749 VTAIL.n57 VTAIL.n16 5.81868
R750 VTAIL.n243 VTAIL.n202 5.81868
R751 VTAIL.n236 VTAIL.n235 5.81868
R752 VTAIL.n153 VTAIL.n112 5.81868
R753 VTAIL.n146 VTAIL.n145 5.81868
R754 VTAIL.n316 VTAIL.n290 5.04292
R755 VTAIL.n328 VTAIL.n284 5.04292
R756 VTAIL.n46 VTAIL.n20 5.04292
R757 VTAIL.n58 VTAIL.n14 5.04292
R758 VTAIL.n244 VTAIL.n200 5.04292
R759 VTAIL.n232 VTAIL.n206 5.04292
R760 VTAIL.n154 VTAIL.n110 5.04292
R761 VTAIL.n142 VTAIL.n116 5.04292
R762 VTAIL.n315 VTAIL.n292 4.26717
R763 VTAIL.n332 VTAIL.n331 4.26717
R764 VTAIL.n45 VTAIL.n22 4.26717
R765 VTAIL.n62 VTAIL.n61 4.26717
R766 VTAIL.n248 VTAIL.n247 4.26717
R767 VTAIL.n231 VTAIL.n208 4.26717
R768 VTAIL.n158 VTAIL.n157 4.26717
R769 VTAIL.n141 VTAIL.n118 4.26717
R770 VTAIL.n299 VTAIL.n297 3.70982
R771 VTAIL.n29 VTAIL.n27 3.70982
R772 VTAIL.n215 VTAIL.n213 3.70982
R773 VTAIL.n125 VTAIL.n123 3.70982
R774 VTAIL.n312 VTAIL.n311 3.49141
R775 VTAIL.n335 VTAIL.n282 3.49141
R776 VTAIL.n42 VTAIL.n41 3.49141
R777 VTAIL.n65 VTAIL.n12 3.49141
R778 VTAIL.n251 VTAIL.n198 3.49141
R779 VTAIL.n228 VTAIL.n227 3.49141
R780 VTAIL.n161 VTAIL.n108 3.49141
R781 VTAIL.n138 VTAIL.n137 3.49141
R782 VTAIL.n308 VTAIL.n294 2.71565
R783 VTAIL.n336 VTAIL.n280 2.71565
R784 VTAIL.n356 VTAIL.n272 2.71565
R785 VTAIL.n38 VTAIL.n24 2.71565
R786 VTAIL.n66 VTAIL.n10 2.71565
R787 VTAIL.n86 VTAIL.n2 2.71565
R788 VTAIL.n270 VTAIL.n186 2.71565
R789 VTAIL.n252 VTAIL.n196 2.71565
R790 VTAIL.n224 VTAIL.n210 2.71565
R791 VTAIL.n180 VTAIL.n96 2.71565
R792 VTAIL.n162 VTAIL.n106 2.71565
R793 VTAIL.n134 VTAIL.n120 2.71565
R794 VTAIL.n358 VTAIL.t18 2.10711
R795 VTAIL.n358 VTAIL.t11 2.10711
R796 VTAIL.n0 VTAIL.t10 2.10711
R797 VTAIL.n0 VTAIL.t19 2.10711
R798 VTAIL.n88 VTAIL.t9 2.10711
R799 VTAIL.n88 VTAIL.t1 2.10711
R800 VTAIL.n90 VTAIL.t0 2.10711
R801 VTAIL.n90 VTAIL.t7 2.10711
R802 VTAIL.n184 VTAIL.t2 2.10711
R803 VTAIL.n184 VTAIL.t3 2.10711
R804 VTAIL.n182 VTAIL.t4 2.10711
R805 VTAIL.n182 VTAIL.t5 2.10711
R806 VTAIL.n94 VTAIL.t13 2.10711
R807 VTAIL.n94 VTAIL.t14 2.10711
R808 VTAIL.n92 VTAIL.t17 2.10711
R809 VTAIL.n92 VTAIL.t16 2.10711
R810 VTAIL.n95 VTAIL.n93 2.06947
R811 VTAIL.n181 VTAIL.n95 2.06947
R812 VTAIL.n185 VTAIL.n183 2.06947
R813 VTAIL.n271 VTAIL.n185 2.06947
R814 VTAIL.n91 VTAIL.n89 2.06947
R815 VTAIL.n89 VTAIL.n87 2.06947
R816 VTAIL.n359 VTAIL.n357 2.06947
R817 VTAIL.n307 VTAIL.n296 1.93989
R818 VTAIL.n341 VTAIL.n339 1.93989
R819 VTAIL.n354 VTAIL.n353 1.93989
R820 VTAIL.n37 VTAIL.n26 1.93989
R821 VTAIL.n71 VTAIL.n69 1.93989
R822 VTAIL.n84 VTAIL.n83 1.93989
R823 VTAIL.n268 VTAIL.n267 1.93989
R824 VTAIL.n256 VTAIL.n255 1.93989
R825 VTAIL.n223 VTAIL.n212 1.93989
R826 VTAIL.n178 VTAIL.n177 1.93989
R827 VTAIL.n166 VTAIL.n165 1.93989
R828 VTAIL.n133 VTAIL.n122 1.93989
R829 VTAIL VTAIL.n1 1.61041
R830 VTAIL.n183 VTAIL.n181 1.50481
R831 VTAIL.n87 VTAIL.n1 1.50481
R832 VTAIL.n304 VTAIL.n303 1.16414
R833 VTAIL.n340 VTAIL.n278 1.16414
R834 VTAIL.n350 VTAIL.n274 1.16414
R835 VTAIL.n34 VTAIL.n33 1.16414
R836 VTAIL.n70 VTAIL.n8 1.16414
R837 VTAIL.n80 VTAIL.n4 1.16414
R838 VTAIL.n264 VTAIL.n188 1.16414
R839 VTAIL.n259 VTAIL.n193 1.16414
R840 VTAIL.n220 VTAIL.n219 1.16414
R841 VTAIL.n174 VTAIL.n98 1.16414
R842 VTAIL.n169 VTAIL.n103 1.16414
R843 VTAIL.n130 VTAIL.n129 1.16414
R844 VTAIL VTAIL.n359 0.459552
R845 VTAIL.n300 VTAIL.n298 0.388379
R846 VTAIL.n346 VTAIL.n345 0.388379
R847 VTAIL.n349 VTAIL.n276 0.388379
R848 VTAIL.n30 VTAIL.n28 0.388379
R849 VTAIL.n76 VTAIL.n75 0.388379
R850 VTAIL.n79 VTAIL.n6 0.388379
R851 VTAIL.n263 VTAIL.n190 0.388379
R852 VTAIL.n260 VTAIL.n192 0.388379
R853 VTAIL.n216 VTAIL.n214 0.388379
R854 VTAIL.n173 VTAIL.n100 0.388379
R855 VTAIL.n170 VTAIL.n102 0.388379
R856 VTAIL.n126 VTAIL.n124 0.388379
R857 VTAIL.n305 VTAIL.n297 0.155672
R858 VTAIL.n306 VTAIL.n305 0.155672
R859 VTAIL.n306 VTAIL.n293 0.155672
R860 VTAIL.n313 VTAIL.n293 0.155672
R861 VTAIL.n314 VTAIL.n313 0.155672
R862 VTAIL.n314 VTAIL.n289 0.155672
R863 VTAIL.n321 VTAIL.n289 0.155672
R864 VTAIL.n322 VTAIL.n321 0.155672
R865 VTAIL.n322 VTAIL.n285 0.155672
R866 VTAIL.n329 VTAIL.n285 0.155672
R867 VTAIL.n330 VTAIL.n329 0.155672
R868 VTAIL.n330 VTAIL.n281 0.155672
R869 VTAIL.n337 VTAIL.n281 0.155672
R870 VTAIL.n338 VTAIL.n337 0.155672
R871 VTAIL.n338 VTAIL.n277 0.155672
R872 VTAIL.n347 VTAIL.n277 0.155672
R873 VTAIL.n348 VTAIL.n347 0.155672
R874 VTAIL.n348 VTAIL.n273 0.155672
R875 VTAIL.n355 VTAIL.n273 0.155672
R876 VTAIL.n35 VTAIL.n27 0.155672
R877 VTAIL.n36 VTAIL.n35 0.155672
R878 VTAIL.n36 VTAIL.n23 0.155672
R879 VTAIL.n43 VTAIL.n23 0.155672
R880 VTAIL.n44 VTAIL.n43 0.155672
R881 VTAIL.n44 VTAIL.n19 0.155672
R882 VTAIL.n51 VTAIL.n19 0.155672
R883 VTAIL.n52 VTAIL.n51 0.155672
R884 VTAIL.n52 VTAIL.n15 0.155672
R885 VTAIL.n59 VTAIL.n15 0.155672
R886 VTAIL.n60 VTAIL.n59 0.155672
R887 VTAIL.n60 VTAIL.n11 0.155672
R888 VTAIL.n67 VTAIL.n11 0.155672
R889 VTAIL.n68 VTAIL.n67 0.155672
R890 VTAIL.n68 VTAIL.n7 0.155672
R891 VTAIL.n77 VTAIL.n7 0.155672
R892 VTAIL.n78 VTAIL.n77 0.155672
R893 VTAIL.n78 VTAIL.n3 0.155672
R894 VTAIL.n85 VTAIL.n3 0.155672
R895 VTAIL.n269 VTAIL.n187 0.155672
R896 VTAIL.n262 VTAIL.n187 0.155672
R897 VTAIL.n262 VTAIL.n261 0.155672
R898 VTAIL.n261 VTAIL.n191 0.155672
R899 VTAIL.n254 VTAIL.n191 0.155672
R900 VTAIL.n254 VTAIL.n253 0.155672
R901 VTAIL.n253 VTAIL.n197 0.155672
R902 VTAIL.n246 VTAIL.n197 0.155672
R903 VTAIL.n246 VTAIL.n245 0.155672
R904 VTAIL.n245 VTAIL.n201 0.155672
R905 VTAIL.n238 VTAIL.n201 0.155672
R906 VTAIL.n238 VTAIL.n237 0.155672
R907 VTAIL.n237 VTAIL.n205 0.155672
R908 VTAIL.n230 VTAIL.n205 0.155672
R909 VTAIL.n230 VTAIL.n229 0.155672
R910 VTAIL.n229 VTAIL.n209 0.155672
R911 VTAIL.n222 VTAIL.n209 0.155672
R912 VTAIL.n222 VTAIL.n221 0.155672
R913 VTAIL.n221 VTAIL.n213 0.155672
R914 VTAIL.n179 VTAIL.n97 0.155672
R915 VTAIL.n172 VTAIL.n97 0.155672
R916 VTAIL.n172 VTAIL.n171 0.155672
R917 VTAIL.n171 VTAIL.n101 0.155672
R918 VTAIL.n164 VTAIL.n101 0.155672
R919 VTAIL.n164 VTAIL.n163 0.155672
R920 VTAIL.n163 VTAIL.n107 0.155672
R921 VTAIL.n156 VTAIL.n107 0.155672
R922 VTAIL.n156 VTAIL.n155 0.155672
R923 VTAIL.n155 VTAIL.n111 0.155672
R924 VTAIL.n148 VTAIL.n111 0.155672
R925 VTAIL.n148 VTAIL.n147 0.155672
R926 VTAIL.n147 VTAIL.n115 0.155672
R927 VTAIL.n140 VTAIL.n115 0.155672
R928 VTAIL.n140 VTAIL.n139 0.155672
R929 VTAIL.n139 VTAIL.n119 0.155672
R930 VTAIL.n132 VTAIL.n119 0.155672
R931 VTAIL.n132 VTAIL.n131 0.155672
R932 VTAIL.n131 VTAIL.n123 0.155672
R933 VP.n18 VP.t8 212.583
R934 VP.n60 VP.t3 179.644
R935 VP.n44 VP.t9 179.644
R936 VP.n7 VP.t1 179.644
R937 VP.n67 VP.t7 179.644
R938 VP.n75 VP.t5 179.644
R939 VP.n26 VP.t6 179.644
R940 VP.n41 VP.t0 179.644
R941 VP.n33 VP.t2 179.644
R942 VP.n17 VP.t4 179.644
R943 VP.n20 VP.n19 161.3
R944 VP.n21 VP.n16 161.3
R945 VP.n23 VP.n22 161.3
R946 VP.n24 VP.n15 161.3
R947 VP.n26 VP.n25 161.3
R948 VP.n27 VP.n14 161.3
R949 VP.n29 VP.n28 161.3
R950 VP.n30 VP.n13 161.3
R951 VP.n32 VP.n31 161.3
R952 VP.n34 VP.n12 161.3
R953 VP.n36 VP.n35 161.3
R954 VP.n37 VP.n11 161.3
R955 VP.n39 VP.n38 161.3
R956 VP.n40 VP.n10 161.3
R957 VP.n74 VP.n0 161.3
R958 VP.n73 VP.n72 161.3
R959 VP.n71 VP.n1 161.3
R960 VP.n70 VP.n69 161.3
R961 VP.n68 VP.n2 161.3
R962 VP.n66 VP.n65 161.3
R963 VP.n64 VP.n3 161.3
R964 VP.n63 VP.n62 161.3
R965 VP.n61 VP.n4 161.3
R966 VP.n60 VP.n59 161.3
R967 VP.n58 VP.n5 161.3
R968 VP.n57 VP.n56 161.3
R969 VP.n55 VP.n6 161.3
R970 VP.n54 VP.n53 161.3
R971 VP.n52 VP.n51 161.3
R972 VP.n50 VP.n8 161.3
R973 VP.n49 VP.n48 161.3
R974 VP.n47 VP.n9 161.3
R975 VP.n46 VP.n45 161.3
R976 VP.n44 VP.n43 96.0763
R977 VP.n76 VP.n75 96.0763
R978 VP.n42 VP.n41 96.0763
R979 VP.n56 VP.n55 56.5193
R980 VP.n62 VP.n3 56.5193
R981 VP.n28 VP.n13 56.5193
R982 VP.n22 VP.n21 56.5193
R983 VP.n43 VP.n42 52.795
R984 VP.n18 VP.n17 51.1767
R985 VP.n49 VP.n9 50.2061
R986 VP.n73 VP.n1 50.2061
R987 VP.n39 VP.n11 50.2061
R988 VP.n50 VP.n49 30.7807
R989 VP.n69 VP.n1 30.7807
R990 VP.n35 VP.n11 30.7807
R991 VP.n45 VP.n9 24.4675
R992 VP.n51 VP.n50 24.4675
R993 VP.n55 VP.n54 24.4675
R994 VP.n56 VP.n5 24.4675
R995 VP.n60 VP.n5 24.4675
R996 VP.n61 VP.n60 24.4675
R997 VP.n62 VP.n61 24.4675
R998 VP.n66 VP.n3 24.4675
R999 VP.n69 VP.n68 24.4675
R1000 VP.n74 VP.n73 24.4675
R1001 VP.n40 VP.n39 24.4675
R1002 VP.n32 VP.n13 24.4675
R1003 VP.n35 VP.n34 24.4675
R1004 VP.n22 VP.n15 24.4675
R1005 VP.n26 VP.n15 24.4675
R1006 VP.n27 VP.n26 24.4675
R1007 VP.n28 VP.n27 24.4675
R1008 VP.n21 VP.n20 24.4675
R1009 VP.n54 VP.n7 19.5741
R1010 VP.n67 VP.n66 19.5741
R1011 VP.n33 VP.n32 19.5741
R1012 VP.n20 VP.n17 19.5741
R1013 VP.n45 VP.n44 14.6807
R1014 VP.n75 VP.n74 14.6807
R1015 VP.n41 VP.n40 14.6807
R1016 VP.n19 VP.n18 9.46762
R1017 VP.n51 VP.n7 4.8939
R1018 VP.n68 VP.n67 4.8939
R1019 VP.n34 VP.n33 4.8939
R1020 VP.n42 VP.n10 0.278367
R1021 VP.n46 VP.n43 0.278367
R1022 VP.n76 VP.n0 0.278367
R1023 VP.n19 VP.n16 0.189894
R1024 VP.n23 VP.n16 0.189894
R1025 VP.n24 VP.n23 0.189894
R1026 VP.n25 VP.n24 0.189894
R1027 VP.n25 VP.n14 0.189894
R1028 VP.n29 VP.n14 0.189894
R1029 VP.n30 VP.n29 0.189894
R1030 VP.n31 VP.n30 0.189894
R1031 VP.n31 VP.n12 0.189894
R1032 VP.n36 VP.n12 0.189894
R1033 VP.n37 VP.n36 0.189894
R1034 VP.n38 VP.n37 0.189894
R1035 VP.n38 VP.n10 0.189894
R1036 VP.n47 VP.n46 0.189894
R1037 VP.n48 VP.n47 0.189894
R1038 VP.n48 VP.n8 0.189894
R1039 VP.n52 VP.n8 0.189894
R1040 VP.n53 VP.n52 0.189894
R1041 VP.n53 VP.n6 0.189894
R1042 VP.n57 VP.n6 0.189894
R1043 VP.n58 VP.n57 0.189894
R1044 VP.n59 VP.n58 0.189894
R1045 VP.n59 VP.n4 0.189894
R1046 VP.n63 VP.n4 0.189894
R1047 VP.n64 VP.n63 0.189894
R1048 VP.n65 VP.n64 0.189894
R1049 VP.n65 VP.n2 0.189894
R1050 VP.n70 VP.n2 0.189894
R1051 VP.n71 VP.n70 0.189894
R1052 VP.n72 VP.n71 0.189894
R1053 VP.n72 VP.n0 0.189894
R1054 VP VP.n76 0.153454
R1055 VDD1.n80 VDD1.n0 756.745
R1056 VDD1.n167 VDD1.n87 756.745
R1057 VDD1.n81 VDD1.n80 585
R1058 VDD1.n79 VDD1.n78 585
R1059 VDD1.n4 VDD1.n3 585
R1060 VDD1.n8 VDD1.n6 585
R1061 VDD1.n73 VDD1.n72 585
R1062 VDD1.n71 VDD1.n70 585
R1063 VDD1.n10 VDD1.n9 585
R1064 VDD1.n65 VDD1.n64 585
R1065 VDD1.n63 VDD1.n62 585
R1066 VDD1.n14 VDD1.n13 585
R1067 VDD1.n57 VDD1.n56 585
R1068 VDD1.n55 VDD1.n54 585
R1069 VDD1.n18 VDD1.n17 585
R1070 VDD1.n49 VDD1.n48 585
R1071 VDD1.n47 VDD1.n46 585
R1072 VDD1.n22 VDD1.n21 585
R1073 VDD1.n41 VDD1.n40 585
R1074 VDD1.n39 VDD1.n38 585
R1075 VDD1.n26 VDD1.n25 585
R1076 VDD1.n33 VDD1.n32 585
R1077 VDD1.n31 VDD1.n30 585
R1078 VDD1.n116 VDD1.n115 585
R1079 VDD1.n118 VDD1.n117 585
R1080 VDD1.n111 VDD1.n110 585
R1081 VDD1.n124 VDD1.n123 585
R1082 VDD1.n126 VDD1.n125 585
R1083 VDD1.n107 VDD1.n106 585
R1084 VDD1.n132 VDD1.n131 585
R1085 VDD1.n134 VDD1.n133 585
R1086 VDD1.n103 VDD1.n102 585
R1087 VDD1.n140 VDD1.n139 585
R1088 VDD1.n142 VDD1.n141 585
R1089 VDD1.n99 VDD1.n98 585
R1090 VDD1.n148 VDD1.n147 585
R1091 VDD1.n150 VDD1.n149 585
R1092 VDD1.n95 VDD1.n94 585
R1093 VDD1.n157 VDD1.n156 585
R1094 VDD1.n158 VDD1.n93 585
R1095 VDD1.n160 VDD1.n159 585
R1096 VDD1.n91 VDD1.n90 585
R1097 VDD1.n166 VDD1.n165 585
R1098 VDD1.n168 VDD1.n167 585
R1099 VDD1.n29 VDD1.t1 327.466
R1100 VDD1.n114 VDD1.t0 327.466
R1101 VDD1.n80 VDD1.n79 171.744
R1102 VDD1.n79 VDD1.n3 171.744
R1103 VDD1.n8 VDD1.n3 171.744
R1104 VDD1.n72 VDD1.n8 171.744
R1105 VDD1.n72 VDD1.n71 171.744
R1106 VDD1.n71 VDD1.n9 171.744
R1107 VDD1.n64 VDD1.n9 171.744
R1108 VDD1.n64 VDD1.n63 171.744
R1109 VDD1.n63 VDD1.n13 171.744
R1110 VDD1.n56 VDD1.n13 171.744
R1111 VDD1.n56 VDD1.n55 171.744
R1112 VDD1.n55 VDD1.n17 171.744
R1113 VDD1.n48 VDD1.n17 171.744
R1114 VDD1.n48 VDD1.n47 171.744
R1115 VDD1.n47 VDD1.n21 171.744
R1116 VDD1.n40 VDD1.n21 171.744
R1117 VDD1.n40 VDD1.n39 171.744
R1118 VDD1.n39 VDD1.n25 171.744
R1119 VDD1.n32 VDD1.n25 171.744
R1120 VDD1.n32 VDD1.n31 171.744
R1121 VDD1.n117 VDD1.n116 171.744
R1122 VDD1.n117 VDD1.n110 171.744
R1123 VDD1.n124 VDD1.n110 171.744
R1124 VDD1.n125 VDD1.n124 171.744
R1125 VDD1.n125 VDD1.n106 171.744
R1126 VDD1.n132 VDD1.n106 171.744
R1127 VDD1.n133 VDD1.n132 171.744
R1128 VDD1.n133 VDD1.n102 171.744
R1129 VDD1.n140 VDD1.n102 171.744
R1130 VDD1.n141 VDD1.n140 171.744
R1131 VDD1.n141 VDD1.n98 171.744
R1132 VDD1.n148 VDD1.n98 171.744
R1133 VDD1.n149 VDD1.n148 171.744
R1134 VDD1.n149 VDD1.n94 171.744
R1135 VDD1.n157 VDD1.n94 171.744
R1136 VDD1.n158 VDD1.n157 171.744
R1137 VDD1.n159 VDD1.n158 171.744
R1138 VDD1.n159 VDD1.n90 171.744
R1139 VDD1.n166 VDD1.n90 171.744
R1140 VDD1.n167 VDD1.n166 171.744
R1141 VDD1.n31 VDD1.t1 85.8723
R1142 VDD1.n116 VDD1.t0 85.8723
R1143 VDD1.n175 VDD1.n174 73.1119
R1144 VDD1.n86 VDD1.n85 71.6157
R1145 VDD1.n173 VDD1.n172 71.6155
R1146 VDD1.n177 VDD1.n176 71.6155
R1147 VDD1.n86 VDD1.n84 52.2907
R1148 VDD1.n173 VDD1.n171 52.2907
R1149 VDD1.n177 VDD1.n175 48.4621
R1150 VDD1.n30 VDD1.n29 16.3895
R1151 VDD1.n115 VDD1.n114 16.3895
R1152 VDD1.n6 VDD1.n4 13.1884
R1153 VDD1.n160 VDD1.n91 13.1884
R1154 VDD1.n78 VDD1.n77 12.8005
R1155 VDD1.n74 VDD1.n73 12.8005
R1156 VDD1.n33 VDD1.n28 12.8005
R1157 VDD1.n118 VDD1.n113 12.8005
R1158 VDD1.n161 VDD1.n93 12.8005
R1159 VDD1.n165 VDD1.n164 12.8005
R1160 VDD1.n81 VDD1.n2 12.0247
R1161 VDD1.n70 VDD1.n7 12.0247
R1162 VDD1.n34 VDD1.n26 12.0247
R1163 VDD1.n119 VDD1.n111 12.0247
R1164 VDD1.n156 VDD1.n155 12.0247
R1165 VDD1.n168 VDD1.n89 12.0247
R1166 VDD1.n82 VDD1.n0 11.249
R1167 VDD1.n69 VDD1.n10 11.249
R1168 VDD1.n38 VDD1.n37 11.249
R1169 VDD1.n123 VDD1.n122 11.249
R1170 VDD1.n154 VDD1.n95 11.249
R1171 VDD1.n169 VDD1.n87 11.249
R1172 VDD1.n66 VDD1.n65 10.4732
R1173 VDD1.n41 VDD1.n24 10.4732
R1174 VDD1.n126 VDD1.n109 10.4732
R1175 VDD1.n151 VDD1.n150 10.4732
R1176 VDD1.n62 VDD1.n12 9.69747
R1177 VDD1.n42 VDD1.n22 9.69747
R1178 VDD1.n127 VDD1.n107 9.69747
R1179 VDD1.n147 VDD1.n97 9.69747
R1180 VDD1.n84 VDD1.n83 9.45567
R1181 VDD1.n171 VDD1.n170 9.45567
R1182 VDD1.n16 VDD1.n15 9.3005
R1183 VDD1.n59 VDD1.n58 9.3005
R1184 VDD1.n61 VDD1.n60 9.3005
R1185 VDD1.n12 VDD1.n11 9.3005
R1186 VDD1.n67 VDD1.n66 9.3005
R1187 VDD1.n69 VDD1.n68 9.3005
R1188 VDD1.n7 VDD1.n5 9.3005
R1189 VDD1.n75 VDD1.n74 9.3005
R1190 VDD1.n83 VDD1.n82 9.3005
R1191 VDD1.n2 VDD1.n1 9.3005
R1192 VDD1.n77 VDD1.n76 9.3005
R1193 VDD1.n53 VDD1.n52 9.3005
R1194 VDD1.n51 VDD1.n50 9.3005
R1195 VDD1.n20 VDD1.n19 9.3005
R1196 VDD1.n45 VDD1.n44 9.3005
R1197 VDD1.n43 VDD1.n42 9.3005
R1198 VDD1.n24 VDD1.n23 9.3005
R1199 VDD1.n37 VDD1.n36 9.3005
R1200 VDD1.n35 VDD1.n34 9.3005
R1201 VDD1.n28 VDD1.n27 9.3005
R1202 VDD1.n170 VDD1.n169 9.3005
R1203 VDD1.n89 VDD1.n88 9.3005
R1204 VDD1.n164 VDD1.n163 9.3005
R1205 VDD1.n136 VDD1.n135 9.3005
R1206 VDD1.n105 VDD1.n104 9.3005
R1207 VDD1.n130 VDD1.n129 9.3005
R1208 VDD1.n128 VDD1.n127 9.3005
R1209 VDD1.n109 VDD1.n108 9.3005
R1210 VDD1.n122 VDD1.n121 9.3005
R1211 VDD1.n120 VDD1.n119 9.3005
R1212 VDD1.n113 VDD1.n112 9.3005
R1213 VDD1.n138 VDD1.n137 9.3005
R1214 VDD1.n101 VDD1.n100 9.3005
R1215 VDD1.n144 VDD1.n143 9.3005
R1216 VDD1.n146 VDD1.n145 9.3005
R1217 VDD1.n97 VDD1.n96 9.3005
R1218 VDD1.n152 VDD1.n151 9.3005
R1219 VDD1.n154 VDD1.n153 9.3005
R1220 VDD1.n155 VDD1.n92 9.3005
R1221 VDD1.n162 VDD1.n161 9.3005
R1222 VDD1.n61 VDD1.n14 8.92171
R1223 VDD1.n46 VDD1.n45 8.92171
R1224 VDD1.n131 VDD1.n130 8.92171
R1225 VDD1.n146 VDD1.n99 8.92171
R1226 VDD1.n58 VDD1.n57 8.14595
R1227 VDD1.n49 VDD1.n20 8.14595
R1228 VDD1.n134 VDD1.n105 8.14595
R1229 VDD1.n143 VDD1.n142 8.14595
R1230 VDD1.n54 VDD1.n16 7.3702
R1231 VDD1.n50 VDD1.n18 7.3702
R1232 VDD1.n135 VDD1.n103 7.3702
R1233 VDD1.n139 VDD1.n101 7.3702
R1234 VDD1.n54 VDD1.n53 6.59444
R1235 VDD1.n53 VDD1.n18 6.59444
R1236 VDD1.n138 VDD1.n103 6.59444
R1237 VDD1.n139 VDD1.n138 6.59444
R1238 VDD1.n57 VDD1.n16 5.81868
R1239 VDD1.n50 VDD1.n49 5.81868
R1240 VDD1.n135 VDD1.n134 5.81868
R1241 VDD1.n142 VDD1.n101 5.81868
R1242 VDD1.n58 VDD1.n14 5.04292
R1243 VDD1.n46 VDD1.n20 5.04292
R1244 VDD1.n131 VDD1.n105 5.04292
R1245 VDD1.n143 VDD1.n99 5.04292
R1246 VDD1.n62 VDD1.n61 4.26717
R1247 VDD1.n45 VDD1.n22 4.26717
R1248 VDD1.n130 VDD1.n107 4.26717
R1249 VDD1.n147 VDD1.n146 4.26717
R1250 VDD1.n29 VDD1.n27 3.70982
R1251 VDD1.n114 VDD1.n112 3.70982
R1252 VDD1.n65 VDD1.n12 3.49141
R1253 VDD1.n42 VDD1.n41 3.49141
R1254 VDD1.n127 VDD1.n126 3.49141
R1255 VDD1.n150 VDD1.n97 3.49141
R1256 VDD1.n84 VDD1.n0 2.71565
R1257 VDD1.n66 VDD1.n10 2.71565
R1258 VDD1.n38 VDD1.n24 2.71565
R1259 VDD1.n123 VDD1.n109 2.71565
R1260 VDD1.n151 VDD1.n95 2.71565
R1261 VDD1.n171 VDD1.n87 2.71565
R1262 VDD1.n176 VDD1.t7 2.10711
R1263 VDD1.n176 VDD1.t9 2.10711
R1264 VDD1.n85 VDD1.t5 2.10711
R1265 VDD1.n85 VDD1.t3 2.10711
R1266 VDD1.n174 VDD1.t2 2.10711
R1267 VDD1.n174 VDD1.t4 2.10711
R1268 VDD1.n172 VDD1.t8 2.10711
R1269 VDD1.n172 VDD1.t6 2.10711
R1270 VDD1.n82 VDD1.n81 1.93989
R1271 VDD1.n70 VDD1.n69 1.93989
R1272 VDD1.n37 VDD1.n26 1.93989
R1273 VDD1.n122 VDD1.n111 1.93989
R1274 VDD1.n156 VDD1.n154 1.93989
R1275 VDD1.n169 VDD1.n168 1.93989
R1276 VDD1 VDD1.n177 1.49403
R1277 VDD1.n78 VDD1.n2 1.16414
R1278 VDD1.n73 VDD1.n7 1.16414
R1279 VDD1.n34 VDD1.n33 1.16414
R1280 VDD1.n119 VDD1.n118 1.16414
R1281 VDD1.n155 VDD1.n93 1.16414
R1282 VDD1.n165 VDD1.n89 1.16414
R1283 VDD1 VDD1.n86 0.575931
R1284 VDD1.n175 VDD1.n173 0.462395
R1285 VDD1.n77 VDD1.n4 0.388379
R1286 VDD1.n74 VDD1.n6 0.388379
R1287 VDD1.n30 VDD1.n28 0.388379
R1288 VDD1.n115 VDD1.n113 0.388379
R1289 VDD1.n161 VDD1.n160 0.388379
R1290 VDD1.n164 VDD1.n91 0.388379
R1291 VDD1.n83 VDD1.n1 0.155672
R1292 VDD1.n76 VDD1.n1 0.155672
R1293 VDD1.n76 VDD1.n75 0.155672
R1294 VDD1.n75 VDD1.n5 0.155672
R1295 VDD1.n68 VDD1.n5 0.155672
R1296 VDD1.n68 VDD1.n67 0.155672
R1297 VDD1.n67 VDD1.n11 0.155672
R1298 VDD1.n60 VDD1.n11 0.155672
R1299 VDD1.n60 VDD1.n59 0.155672
R1300 VDD1.n59 VDD1.n15 0.155672
R1301 VDD1.n52 VDD1.n15 0.155672
R1302 VDD1.n52 VDD1.n51 0.155672
R1303 VDD1.n51 VDD1.n19 0.155672
R1304 VDD1.n44 VDD1.n19 0.155672
R1305 VDD1.n44 VDD1.n43 0.155672
R1306 VDD1.n43 VDD1.n23 0.155672
R1307 VDD1.n36 VDD1.n23 0.155672
R1308 VDD1.n36 VDD1.n35 0.155672
R1309 VDD1.n35 VDD1.n27 0.155672
R1310 VDD1.n120 VDD1.n112 0.155672
R1311 VDD1.n121 VDD1.n120 0.155672
R1312 VDD1.n121 VDD1.n108 0.155672
R1313 VDD1.n128 VDD1.n108 0.155672
R1314 VDD1.n129 VDD1.n128 0.155672
R1315 VDD1.n129 VDD1.n104 0.155672
R1316 VDD1.n136 VDD1.n104 0.155672
R1317 VDD1.n137 VDD1.n136 0.155672
R1318 VDD1.n137 VDD1.n100 0.155672
R1319 VDD1.n144 VDD1.n100 0.155672
R1320 VDD1.n145 VDD1.n144 0.155672
R1321 VDD1.n145 VDD1.n96 0.155672
R1322 VDD1.n152 VDD1.n96 0.155672
R1323 VDD1.n153 VDD1.n152 0.155672
R1324 VDD1.n153 VDD1.n92 0.155672
R1325 VDD1.n162 VDD1.n92 0.155672
R1326 VDD1.n163 VDD1.n162 0.155672
R1327 VDD1.n163 VDD1.n88 0.155672
R1328 VDD1.n170 VDD1.n88 0.155672
R1329 B.n468 B.n467 585
R1330 B.n466 B.n139 585
R1331 B.n465 B.n464 585
R1332 B.n463 B.n140 585
R1333 B.n462 B.n461 585
R1334 B.n460 B.n141 585
R1335 B.n459 B.n458 585
R1336 B.n457 B.n142 585
R1337 B.n456 B.n455 585
R1338 B.n454 B.n143 585
R1339 B.n453 B.n452 585
R1340 B.n451 B.n144 585
R1341 B.n450 B.n449 585
R1342 B.n448 B.n145 585
R1343 B.n447 B.n446 585
R1344 B.n445 B.n146 585
R1345 B.n444 B.n443 585
R1346 B.n442 B.n147 585
R1347 B.n441 B.n440 585
R1348 B.n439 B.n148 585
R1349 B.n438 B.n437 585
R1350 B.n436 B.n149 585
R1351 B.n435 B.n434 585
R1352 B.n433 B.n150 585
R1353 B.n432 B.n431 585
R1354 B.n430 B.n151 585
R1355 B.n429 B.n428 585
R1356 B.n427 B.n152 585
R1357 B.n426 B.n425 585
R1358 B.n424 B.n153 585
R1359 B.n423 B.n422 585
R1360 B.n421 B.n154 585
R1361 B.n420 B.n419 585
R1362 B.n418 B.n155 585
R1363 B.n417 B.n416 585
R1364 B.n415 B.n156 585
R1365 B.n414 B.n413 585
R1366 B.n412 B.n157 585
R1367 B.n411 B.n410 585
R1368 B.n409 B.n158 585
R1369 B.n408 B.n407 585
R1370 B.n406 B.n159 585
R1371 B.n405 B.n404 585
R1372 B.n403 B.n160 585
R1373 B.n402 B.n401 585
R1374 B.n400 B.n161 585
R1375 B.n399 B.n398 585
R1376 B.n397 B.n162 585
R1377 B.n396 B.n395 585
R1378 B.n394 B.n163 585
R1379 B.n393 B.n392 585
R1380 B.n391 B.n164 585
R1381 B.n390 B.n389 585
R1382 B.n385 B.n165 585
R1383 B.n384 B.n383 585
R1384 B.n382 B.n166 585
R1385 B.n381 B.n380 585
R1386 B.n379 B.n167 585
R1387 B.n378 B.n377 585
R1388 B.n376 B.n168 585
R1389 B.n375 B.n374 585
R1390 B.n372 B.n169 585
R1391 B.n371 B.n370 585
R1392 B.n369 B.n172 585
R1393 B.n368 B.n367 585
R1394 B.n366 B.n173 585
R1395 B.n365 B.n364 585
R1396 B.n363 B.n174 585
R1397 B.n362 B.n361 585
R1398 B.n360 B.n175 585
R1399 B.n359 B.n358 585
R1400 B.n357 B.n176 585
R1401 B.n356 B.n355 585
R1402 B.n354 B.n177 585
R1403 B.n353 B.n352 585
R1404 B.n351 B.n178 585
R1405 B.n350 B.n349 585
R1406 B.n348 B.n179 585
R1407 B.n347 B.n346 585
R1408 B.n345 B.n180 585
R1409 B.n344 B.n343 585
R1410 B.n342 B.n181 585
R1411 B.n341 B.n340 585
R1412 B.n339 B.n182 585
R1413 B.n338 B.n337 585
R1414 B.n336 B.n183 585
R1415 B.n335 B.n334 585
R1416 B.n333 B.n184 585
R1417 B.n332 B.n331 585
R1418 B.n330 B.n185 585
R1419 B.n329 B.n328 585
R1420 B.n327 B.n186 585
R1421 B.n326 B.n325 585
R1422 B.n324 B.n187 585
R1423 B.n323 B.n322 585
R1424 B.n321 B.n188 585
R1425 B.n320 B.n319 585
R1426 B.n318 B.n189 585
R1427 B.n317 B.n316 585
R1428 B.n315 B.n190 585
R1429 B.n314 B.n313 585
R1430 B.n312 B.n191 585
R1431 B.n311 B.n310 585
R1432 B.n309 B.n192 585
R1433 B.n308 B.n307 585
R1434 B.n306 B.n193 585
R1435 B.n305 B.n304 585
R1436 B.n303 B.n194 585
R1437 B.n302 B.n301 585
R1438 B.n300 B.n195 585
R1439 B.n299 B.n298 585
R1440 B.n297 B.n196 585
R1441 B.n296 B.n295 585
R1442 B.n469 B.n138 585
R1443 B.n471 B.n470 585
R1444 B.n472 B.n137 585
R1445 B.n474 B.n473 585
R1446 B.n475 B.n136 585
R1447 B.n477 B.n476 585
R1448 B.n478 B.n135 585
R1449 B.n480 B.n479 585
R1450 B.n481 B.n134 585
R1451 B.n483 B.n482 585
R1452 B.n484 B.n133 585
R1453 B.n486 B.n485 585
R1454 B.n487 B.n132 585
R1455 B.n489 B.n488 585
R1456 B.n490 B.n131 585
R1457 B.n492 B.n491 585
R1458 B.n493 B.n130 585
R1459 B.n495 B.n494 585
R1460 B.n496 B.n129 585
R1461 B.n498 B.n497 585
R1462 B.n499 B.n128 585
R1463 B.n501 B.n500 585
R1464 B.n502 B.n127 585
R1465 B.n504 B.n503 585
R1466 B.n505 B.n126 585
R1467 B.n507 B.n506 585
R1468 B.n508 B.n125 585
R1469 B.n510 B.n509 585
R1470 B.n511 B.n124 585
R1471 B.n513 B.n512 585
R1472 B.n514 B.n123 585
R1473 B.n516 B.n515 585
R1474 B.n517 B.n122 585
R1475 B.n519 B.n518 585
R1476 B.n520 B.n121 585
R1477 B.n522 B.n521 585
R1478 B.n523 B.n120 585
R1479 B.n525 B.n524 585
R1480 B.n526 B.n119 585
R1481 B.n528 B.n527 585
R1482 B.n529 B.n118 585
R1483 B.n531 B.n530 585
R1484 B.n532 B.n117 585
R1485 B.n534 B.n533 585
R1486 B.n535 B.n116 585
R1487 B.n537 B.n536 585
R1488 B.n538 B.n115 585
R1489 B.n540 B.n539 585
R1490 B.n541 B.n114 585
R1491 B.n543 B.n542 585
R1492 B.n544 B.n113 585
R1493 B.n546 B.n545 585
R1494 B.n547 B.n112 585
R1495 B.n549 B.n548 585
R1496 B.n550 B.n111 585
R1497 B.n552 B.n551 585
R1498 B.n553 B.n110 585
R1499 B.n555 B.n554 585
R1500 B.n556 B.n109 585
R1501 B.n558 B.n557 585
R1502 B.n559 B.n108 585
R1503 B.n561 B.n560 585
R1504 B.n562 B.n107 585
R1505 B.n564 B.n563 585
R1506 B.n565 B.n106 585
R1507 B.n567 B.n566 585
R1508 B.n568 B.n105 585
R1509 B.n570 B.n569 585
R1510 B.n571 B.n104 585
R1511 B.n573 B.n572 585
R1512 B.n574 B.n103 585
R1513 B.n576 B.n575 585
R1514 B.n577 B.n102 585
R1515 B.n579 B.n578 585
R1516 B.n580 B.n101 585
R1517 B.n582 B.n581 585
R1518 B.n583 B.n100 585
R1519 B.n585 B.n584 585
R1520 B.n586 B.n99 585
R1521 B.n588 B.n587 585
R1522 B.n589 B.n98 585
R1523 B.n591 B.n590 585
R1524 B.n592 B.n97 585
R1525 B.n594 B.n593 585
R1526 B.n595 B.n96 585
R1527 B.n597 B.n596 585
R1528 B.n598 B.n95 585
R1529 B.n600 B.n599 585
R1530 B.n601 B.n94 585
R1531 B.n603 B.n602 585
R1532 B.n604 B.n93 585
R1533 B.n606 B.n605 585
R1534 B.n607 B.n92 585
R1535 B.n609 B.n608 585
R1536 B.n610 B.n91 585
R1537 B.n612 B.n611 585
R1538 B.n613 B.n90 585
R1539 B.n615 B.n614 585
R1540 B.n616 B.n89 585
R1541 B.n618 B.n617 585
R1542 B.n619 B.n88 585
R1543 B.n621 B.n620 585
R1544 B.n792 B.n27 585
R1545 B.n791 B.n790 585
R1546 B.n789 B.n28 585
R1547 B.n788 B.n787 585
R1548 B.n786 B.n29 585
R1549 B.n785 B.n784 585
R1550 B.n783 B.n30 585
R1551 B.n782 B.n781 585
R1552 B.n780 B.n31 585
R1553 B.n779 B.n778 585
R1554 B.n777 B.n32 585
R1555 B.n776 B.n775 585
R1556 B.n774 B.n33 585
R1557 B.n773 B.n772 585
R1558 B.n771 B.n34 585
R1559 B.n770 B.n769 585
R1560 B.n768 B.n35 585
R1561 B.n767 B.n766 585
R1562 B.n765 B.n36 585
R1563 B.n764 B.n763 585
R1564 B.n762 B.n37 585
R1565 B.n761 B.n760 585
R1566 B.n759 B.n38 585
R1567 B.n758 B.n757 585
R1568 B.n756 B.n39 585
R1569 B.n755 B.n754 585
R1570 B.n753 B.n40 585
R1571 B.n752 B.n751 585
R1572 B.n750 B.n41 585
R1573 B.n749 B.n748 585
R1574 B.n747 B.n42 585
R1575 B.n746 B.n745 585
R1576 B.n744 B.n43 585
R1577 B.n743 B.n742 585
R1578 B.n741 B.n44 585
R1579 B.n740 B.n739 585
R1580 B.n738 B.n45 585
R1581 B.n737 B.n736 585
R1582 B.n735 B.n46 585
R1583 B.n734 B.n733 585
R1584 B.n732 B.n47 585
R1585 B.n731 B.n730 585
R1586 B.n729 B.n48 585
R1587 B.n728 B.n727 585
R1588 B.n726 B.n49 585
R1589 B.n725 B.n724 585
R1590 B.n723 B.n50 585
R1591 B.n722 B.n721 585
R1592 B.n720 B.n51 585
R1593 B.n719 B.n718 585
R1594 B.n717 B.n52 585
R1595 B.n716 B.n715 585
R1596 B.n713 B.n53 585
R1597 B.n712 B.n711 585
R1598 B.n710 B.n56 585
R1599 B.n709 B.n708 585
R1600 B.n707 B.n57 585
R1601 B.n706 B.n705 585
R1602 B.n704 B.n58 585
R1603 B.n703 B.n702 585
R1604 B.n701 B.n59 585
R1605 B.n699 B.n698 585
R1606 B.n697 B.n62 585
R1607 B.n696 B.n695 585
R1608 B.n694 B.n63 585
R1609 B.n693 B.n692 585
R1610 B.n691 B.n64 585
R1611 B.n690 B.n689 585
R1612 B.n688 B.n65 585
R1613 B.n687 B.n686 585
R1614 B.n685 B.n66 585
R1615 B.n684 B.n683 585
R1616 B.n682 B.n67 585
R1617 B.n681 B.n680 585
R1618 B.n679 B.n68 585
R1619 B.n678 B.n677 585
R1620 B.n676 B.n69 585
R1621 B.n675 B.n674 585
R1622 B.n673 B.n70 585
R1623 B.n672 B.n671 585
R1624 B.n670 B.n71 585
R1625 B.n669 B.n668 585
R1626 B.n667 B.n72 585
R1627 B.n666 B.n665 585
R1628 B.n664 B.n73 585
R1629 B.n663 B.n662 585
R1630 B.n661 B.n74 585
R1631 B.n660 B.n659 585
R1632 B.n658 B.n75 585
R1633 B.n657 B.n656 585
R1634 B.n655 B.n76 585
R1635 B.n654 B.n653 585
R1636 B.n652 B.n77 585
R1637 B.n651 B.n650 585
R1638 B.n649 B.n78 585
R1639 B.n648 B.n647 585
R1640 B.n646 B.n79 585
R1641 B.n645 B.n644 585
R1642 B.n643 B.n80 585
R1643 B.n642 B.n641 585
R1644 B.n640 B.n81 585
R1645 B.n639 B.n638 585
R1646 B.n637 B.n82 585
R1647 B.n636 B.n635 585
R1648 B.n634 B.n83 585
R1649 B.n633 B.n632 585
R1650 B.n631 B.n84 585
R1651 B.n630 B.n629 585
R1652 B.n628 B.n85 585
R1653 B.n627 B.n626 585
R1654 B.n625 B.n86 585
R1655 B.n624 B.n623 585
R1656 B.n622 B.n87 585
R1657 B.n794 B.n793 585
R1658 B.n795 B.n26 585
R1659 B.n797 B.n796 585
R1660 B.n798 B.n25 585
R1661 B.n800 B.n799 585
R1662 B.n801 B.n24 585
R1663 B.n803 B.n802 585
R1664 B.n804 B.n23 585
R1665 B.n806 B.n805 585
R1666 B.n807 B.n22 585
R1667 B.n809 B.n808 585
R1668 B.n810 B.n21 585
R1669 B.n812 B.n811 585
R1670 B.n813 B.n20 585
R1671 B.n815 B.n814 585
R1672 B.n816 B.n19 585
R1673 B.n818 B.n817 585
R1674 B.n819 B.n18 585
R1675 B.n821 B.n820 585
R1676 B.n822 B.n17 585
R1677 B.n824 B.n823 585
R1678 B.n825 B.n16 585
R1679 B.n827 B.n826 585
R1680 B.n828 B.n15 585
R1681 B.n830 B.n829 585
R1682 B.n831 B.n14 585
R1683 B.n833 B.n832 585
R1684 B.n834 B.n13 585
R1685 B.n836 B.n835 585
R1686 B.n837 B.n12 585
R1687 B.n839 B.n838 585
R1688 B.n840 B.n11 585
R1689 B.n842 B.n841 585
R1690 B.n843 B.n10 585
R1691 B.n845 B.n844 585
R1692 B.n846 B.n9 585
R1693 B.n848 B.n847 585
R1694 B.n849 B.n8 585
R1695 B.n851 B.n850 585
R1696 B.n852 B.n7 585
R1697 B.n854 B.n853 585
R1698 B.n855 B.n6 585
R1699 B.n857 B.n856 585
R1700 B.n858 B.n5 585
R1701 B.n860 B.n859 585
R1702 B.n861 B.n4 585
R1703 B.n863 B.n862 585
R1704 B.n864 B.n3 585
R1705 B.n866 B.n865 585
R1706 B.n867 B.n0 585
R1707 B.n2 B.n1 585
R1708 B.n222 B.n221 585
R1709 B.n224 B.n223 585
R1710 B.n225 B.n220 585
R1711 B.n227 B.n226 585
R1712 B.n228 B.n219 585
R1713 B.n230 B.n229 585
R1714 B.n231 B.n218 585
R1715 B.n233 B.n232 585
R1716 B.n234 B.n217 585
R1717 B.n236 B.n235 585
R1718 B.n237 B.n216 585
R1719 B.n239 B.n238 585
R1720 B.n240 B.n215 585
R1721 B.n242 B.n241 585
R1722 B.n243 B.n214 585
R1723 B.n245 B.n244 585
R1724 B.n246 B.n213 585
R1725 B.n248 B.n247 585
R1726 B.n249 B.n212 585
R1727 B.n251 B.n250 585
R1728 B.n252 B.n211 585
R1729 B.n254 B.n253 585
R1730 B.n255 B.n210 585
R1731 B.n257 B.n256 585
R1732 B.n258 B.n209 585
R1733 B.n260 B.n259 585
R1734 B.n261 B.n208 585
R1735 B.n263 B.n262 585
R1736 B.n264 B.n207 585
R1737 B.n266 B.n265 585
R1738 B.n267 B.n206 585
R1739 B.n269 B.n268 585
R1740 B.n270 B.n205 585
R1741 B.n272 B.n271 585
R1742 B.n273 B.n204 585
R1743 B.n275 B.n274 585
R1744 B.n276 B.n203 585
R1745 B.n278 B.n277 585
R1746 B.n279 B.n202 585
R1747 B.n281 B.n280 585
R1748 B.n282 B.n201 585
R1749 B.n284 B.n283 585
R1750 B.n285 B.n200 585
R1751 B.n287 B.n286 585
R1752 B.n288 B.n199 585
R1753 B.n290 B.n289 585
R1754 B.n291 B.n198 585
R1755 B.n293 B.n292 585
R1756 B.n294 B.n197 585
R1757 B.n296 B.n197 492.5
R1758 B.n469 B.n468 492.5
R1759 B.n620 B.n87 492.5
R1760 B.n794 B.n27 492.5
R1761 B.n386 B.t7 483.896
R1762 B.n60 B.t2 483.896
R1763 B.n170 B.t10 483.896
R1764 B.n54 B.t5 483.896
R1765 B.n387 B.t8 437.351
R1766 B.n61 B.t1 437.351
R1767 B.n171 B.t11 437.351
R1768 B.n55 B.t4 437.351
R1769 B.n170 B.t9 386.721
R1770 B.n386 B.t6 386.721
R1771 B.n60 B.t0 386.721
R1772 B.n54 B.t3 386.721
R1773 B.n869 B.n868 256.663
R1774 B.n868 B.n867 235.042
R1775 B.n868 B.n2 235.042
R1776 B.n297 B.n296 163.367
R1777 B.n298 B.n297 163.367
R1778 B.n298 B.n195 163.367
R1779 B.n302 B.n195 163.367
R1780 B.n303 B.n302 163.367
R1781 B.n304 B.n303 163.367
R1782 B.n304 B.n193 163.367
R1783 B.n308 B.n193 163.367
R1784 B.n309 B.n308 163.367
R1785 B.n310 B.n309 163.367
R1786 B.n310 B.n191 163.367
R1787 B.n314 B.n191 163.367
R1788 B.n315 B.n314 163.367
R1789 B.n316 B.n315 163.367
R1790 B.n316 B.n189 163.367
R1791 B.n320 B.n189 163.367
R1792 B.n321 B.n320 163.367
R1793 B.n322 B.n321 163.367
R1794 B.n322 B.n187 163.367
R1795 B.n326 B.n187 163.367
R1796 B.n327 B.n326 163.367
R1797 B.n328 B.n327 163.367
R1798 B.n328 B.n185 163.367
R1799 B.n332 B.n185 163.367
R1800 B.n333 B.n332 163.367
R1801 B.n334 B.n333 163.367
R1802 B.n334 B.n183 163.367
R1803 B.n338 B.n183 163.367
R1804 B.n339 B.n338 163.367
R1805 B.n340 B.n339 163.367
R1806 B.n340 B.n181 163.367
R1807 B.n344 B.n181 163.367
R1808 B.n345 B.n344 163.367
R1809 B.n346 B.n345 163.367
R1810 B.n346 B.n179 163.367
R1811 B.n350 B.n179 163.367
R1812 B.n351 B.n350 163.367
R1813 B.n352 B.n351 163.367
R1814 B.n352 B.n177 163.367
R1815 B.n356 B.n177 163.367
R1816 B.n357 B.n356 163.367
R1817 B.n358 B.n357 163.367
R1818 B.n358 B.n175 163.367
R1819 B.n362 B.n175 163.367
R1820 B.n363 B.n362 163.367
R1821 B.n364 B.n363 163.367
R1822 B.n364 B.n173 163.367
R1823 B.n368 B.n173 163.367
R1824 B.n369 B.n368 163.367
R1825 B.n370 B.n369 163.367
R1826 B.n370 B.n169 163.367
R1827 B.n375 B.n169 163.367
R1828 B.n376 B.n375 163.367
R1829 B.n377 B.n376 163.367
R1830 B.n377 B.n167 163.367
R1831 B.n381 B.n167 163.367
R1832 B.n382 B.n381 163.367
R1833 B.n383 B.n382 163.367
R1834 B.n383 B.n165 163.367
R1835 B.n390 B.n165 163.367
R1836 B.n391 B.n390 163.367
R1837 B.n392 B.n391 163.367
R1838 B.n392 B.n163 163.367
R1839 B.n396 B.n163 163.367
R1840 B.n397 B.n396 163.367
R1841 B.n398 B.n397 163.367
R1842 B.n398 B.n161 163.367
R1843 B.n402 B.n161 163.367
R1844 B.n403 B.n402 163.367
R1845 B.n404 B.n403 163.367
R1846 B.n404 B.n159 163.367
R1847 B.n408 B.n159 163.367
R1848 B.n409 B.n408 163.367
R1849 B.n410 B.n409 163.367
R1850 B.n410 B.n157 163.367
R1851 B.n414 B.n157 163.367
R1852 B.n415 B.n414 163.367
R1853 B.n416 B.n415 163.367
R1854 B.n416 B.n155 163.367
R1855 B.n420 B.n155 163.367
R1856 B.n421 B.n420 163.367
R1857 B.n422 B.n421 163.367
R1858 B.n422 B.n153 163.367
R1859 B.n426 B.n153 163.367
R1860 B.n427 B.n426 163.367
R1861 B.n428 B.n427 163.367
R1862 B.n428 B.n151 163.367
R1863 B.n432 B.n151 163.367
R1864 B.n433 B.n432 163.367
R1865 B.n434 B.n433 163.367
R1866 B.n434 B.n149 163.367
R1867 B.n438 B.n149 163.367
R1868 B.n439 B.n438 163.367
R1869 B.n440 B.n439 163.367
R1870 B.n440 B.n147 163.367
R1871 B.n444 B.n147 163.367
R1872 B.n445 B.n444 163.367
R1873 B.n446 B.n445 163.367
R1874 B.n446 B.n145 163.367
R1875 B.n450 B.n145 163.367
R1876 B.n451 B.n450 163.367
R1877 B.n452 B.n451 163.367
R1878 B.n452 B.n143 163.367
R1879 B.n456 B.n143 163.367
R1880 B.n457 B.n456 163.367
R1881 B.n458 B.n457 163.367
R1882 B.n458 B.n141 163.367
R1883 B.n462 B.n141 163.367
R1884 B.n463 B.n462 163.367
R1885 B.n464 B.n463 163.367
R1886 B.n464 B.n139 163.367
R1887 B.n468 B.n139 163.367
R1888 B.n620 B.n619 163.367
R1889 B.n619 B.n618 163.367
R1890 B.n618 B.n89 163.367
R1891 B.n614 B.n89 163.367
R1892 B.n614 B.n613 163.367
R1893 B.n613 B.n612 163.367
R1894 B.n612 B.n91 163.367
R1895 B.n608 B.n91 163.367
R1896 B.n608 B.n607 163.367
R1897 B.n607 B.n606 163.367
R1898 B.n606 B.n93 163.367
R1899 B.n602 B.n93 163.367
R1900 B.n602 B.n601 163.367
R1901 B.n601 B.n600 163.367
R1902 B.n600 B.n95 163.367
R1903 B.n596 B.n95 163.367
R1904 B.n596 B.n595 163.367
R1905 B.n595 B.n594 163.367
R1906 B.n594 B.n97 163.367
R1907 B.n590 B.n97 163.367
R1908 B.n590 B.n589 163.367
R1909 B.n589 B.n588 163.367
R1910 B.n588 B.n99 163.367
R1911 B.n584 B.n99 163.367
R1912 B.n584 B.n583 163.367
R1913 B.n583 B.n582 163.367
R1914 B.n582 B.n101 163.367
R1915 B.n578 B.n101 163.367
R1916 B.n578 B.n577 163.367
R1917 B.n577 B.n576 163.367
R1918 B.n576 B.n103 163.367
R1919 B.n572 B.n103 163.367
R1920 B.n572 B.n571 163.367
R1921 B.n571 B.n570 163.367
R1922 B.n570 B.n105 163.367
R1923 B.n566 B.n105 163.367
R1924 B.n566 B.n565 163.367
R1925 B.n565 B.n564 163.367
R1926 B.n564 B.n107 163.367
R1927 B.n560 B.n107 163.367
R1928 B.n560 B.n559 163.367
R1929 B.n559 B.n558 163.367
R1930 B.n558 B.n109 163.367
R1931 B.n554 B.n109 163.367
R1932 B.n554 B.n553 163.367
R1933 B.n553 B.n552 163.367
R1934 B.n552 B.n111 163.367
R1935 B.n548 B.n111 163.367
R1936 B.n548 B.n547 163.367
R1937 B.n547 B.n546 163.367
R1938 B.n546 B.n113 163.367
R1939 B.n542 B.n113 163.367
R1940 B.n542 B.n541 163.367
R1941 B.n541 B.n540 163.367
R1942 B.n540 B.n115 163.367
R1943 B.n536 B.n115 163.367
R1944 B.n536 B.n535 163.367
R1945 B.n535 B.n534 163.367
R1946 B.n534 B.n117 163.367
R1947 B.n530 B.n117 163.367
R1948 B.n530 B.n529 163.367
R1949 B.n529 B.n528 163.367
R1950 B.n528 B.n119 163.367
R1951 B.n524 B.n119 163.367
R1952 B.n524 B.n523 163.367
R1953 B.n523 B.n522 163.367
R1954 B.n522 B.n121 163.367
R1955 B.n518 B.n121 163.367
R1956 B.n518 B.n517 163.367
R1957 B.n517 B.n516 163.367
R1958 B.n516 B.n123 163.367
R1959 B.n512 B.n123 163.367
R1960 B.n512 B.n511 163.367
R1961 B.n511 B.n510 163.367
R1962 B.n510 B.n125 163.367
R1963 B.n506 B.n125 163.367
R1964 B.n506 B.n505 163.367
R1965 B.n505 B.n504 163.367
R1966 B.n504 B.n127 163.367
R1967 B.n500 B.n127 163.367
R1968 B.n500 B.n499 163.367
R1969 B.n499 B.n498 163.367
R1970 B.n498 B.n129 163.367
R1971 B.n494 B.n129 163.367
R1972 B.n494 B.n493 163.367
R1973 B.n493 B.n492 163.367
R1974 B.n492 B.n131 163.367
R1975 B.n488 B.n131 163.367
R1976 B.n488 B.n487 163.367
R1977 B.n487 B.n486 163.367
R1978 B.n486 B.n133 163.367
R1979 B.n482 B.n133 163.367
R1980 B.n482 B.n481 163.367
R1981 B.n481 B.n480 163.367
R1982 B.n480 B.n135 163.367
R1983 B.n476 B.n135 163.367
R1984 B.n476 B.n475 163.367
R1985 B.n475 B.n474 163.367
R1986 B.n474 B.n137 163.367
R1987 B.n470 B.n137 163.367
R1988 B.n470 B.n469 163.367
R1989 B.n790 B.n27 163.367
R1990 B.n790 B.n789 163.367
R1991 B.n789 B.n788 163.367
R1992 B.n788 B.n29 163.367
R1993 B.n784 B.n29 163.367
R1994 B.n784 B.n783 163.367
R1995 B.n783 B.n782 163.367
R1996 B.n782 B.n31 163.367
R1997 B.n778 B.n31 163.367
R1998 B.n778 B.n777 163.367
R1999 B.n777 B.n776 163.367
R2000 B.n776 B.n33 163.367
R2001 B.n772 B.n33 163.367
R2002 B.n772 B.n771 163.367
R2003 B.n771 B.n770 163.367
R2004 B.n770 B.n35 163.367
R2005 B.n766 B.n35 163.367
R2006 B.n766 B.n765 163.367
R2007 B.n765 B.n764 163.367
R2008 B.n764 B.n37 163.367
R2009 B.n760 B.n37 163.367
R2010 B.n760 B.n759 163.367
R2011 B.n759 B.n758 163.367
R2012 B.n758 B.n39 163.367
R2013 B.n754 B.n39 163.367
R2014 B.n754 B.n753 163.367
R2015 B.n753 B.n752 163.367
R2016 B.n752 B.n41 163.367
R2017 B.n748 B.n41 163.367
R2018 B.n748 B.n747 163.367
R2019 B.n747 B.n746 163.367
R2020 B.n746 B.n43 163.367
R2021 B.n742 B.n43 163.367
R2022 B.n742 B.n741 163.367
R2023 B.n741 B.n740 163.367
R2024 B.n740 B.n45 163.367
R2025 B.n736 B.n45 163.367
R2026 B.n736 B.n735 163.367
R2027 B.n735 B.n734 163.367
R2028 B.n734 B.n47 163.367
R2029 B.n730 B.n47 163.367
R2030 B.n730 B.n729 163.367
R2031 B.n729 B.n728 163.367
R2032 B.n728 B.n49 163.367
R2033 B.n724 B.n49 163.367
R2034 B.n724 B.n723 163.367
R2035 B.n723 B.n722 163.367
R2036 B.n722 B.n51 163.367
R2037 B.n718 B.n51 163.367
R2038 B.n718 B.n717 163.367
R2039 B.n717 B.n716 163.367
R2040 B.n716 B.n53 163.367
R2041 B.n711 B.n53 163.367
R2042 B.n711 B.n710 163.367
R2043 B.n710 B.n709 163.367
R2044 B.n709 B.n57 163.367
R2045 B.n705 B.n57 163.367
R2046 B.n705 B.n704 163.367
R2047 B.n704 B.n703 163.367
R2048 B.n703 B.n59 163.367
R2049 B.n698 B.n59 163.367
R2050 B.n698 B.n697 163.367
R2051 B.n697 B.n696 163.367
R2052 B.n696 B.n63 163.367
R2053 B.n692 B.n63 163.367
R2054 B.n692 B.n691 163.367
R2055 B.n691 B.n690 163.367
R2056 B.n690 B.n65 163.367
R2057 B.n686 B.n65 163.367
R2058 B.n686 B.n685 163.367
R2059 B.n685 B.n684 163.367
R2060 B.n684 B.n67 163.367
R2061 B.n680 B.n67 163.367
R2062 B.n680 B.n679 163.367
R2063 B.n679 B.n678 163.367
R2064 B.n678 B.n69 163.367
R2065 B.n674 B.n69 163.367
R2066 B.n674 B.n673 163.367
R2067 B.n673 B.n672 163.367
R2068 B.n672 B.n71 163.367
R2069 B.n668 B.n71 163.367
R2070 B.n668 B.n667 163.367
R2071 B.n667 B.n666 163.367
R2072 B.n666 B.n73 163.367
R2073 B.n662 B.n73 163.367
R2074 B.n662 B.n661 163.367
R2075 B.n661 B.n660 163.367
R2076 B.n660 B.n75 163.367
R2077 B.n656 B.n75 163.367
R2078 B.n656 B.n655 163.367
R2079 B.n655 B.n654 163.367
R2080 B.n654 B.n77 163.367
R2081 B.n650 B.n77 163.367
R2082 B.n650 B.n649 163.367
R2083 B.n649 B.n648 163.367
R2084 B.n648 B.n79 163.367
R2085 B.n644 B.n79 163.367
R2086 B.n644 B.n643 163.367
R2087 B.n643 B.n642 163.367
R2088 B.n642 B.n81 163.367
R2089 B.n638 B.n81 163.367
R2090 B.n638 B.n637 163.367
R2091 B.n637 B.n636 163.367
R2092 B.n636 B.n83 163.367
R2093 B.n632 B.n83 163.367
R2094 B.n632 B.n631 163.367
R2095 B.n631 B.n630 163.367
R2096 B.n630 B.n85 163.367
R2097 B.n626 B.n85 163.367
R2098 B.n626 B.n625 163.367
R2099 B.n625 B.n624 163.367
R2100 B.n624 B.n87 163.367
R2101 B.n795 B.n794 163.367
R2102 B.n796 B.n795 163.367
R2103 B.n796 B.n25 163.367
R2104 B.n800 B.n25 163.367
R2105 B.n801 B.n800 163.367
R2106 B.n802 B.n801 163.367
R2107 B.n802 B.n23 163.367
R2108 B.n806 B.n23 163.367
R2109 B.n807 B.n806 163.367
R2110 B.n808 B.n807 163.367
R2111 B.n808 B.n21 163.367
R2112 B.n812 B.n21 163.367
R2113 B.n813 B.n812 163.367
R2114 B.n814 B.n813 163.367
R2115 B.n814 B.n19 163.367
R2116 B.n818 B.n19 163.367
R2117 B.n819 B.n818 163.367
R2118 B.n820 B.n819 163.367
R2119 B.n820 B.n17 163.367
R2120 B.n824 B.n17 163.367
R2121 B.n825 B.n824 163.367
R2122 B.n826 B.n825 163.367
R2123 B.n826 B.n15 163.367
R2124 B.n830 B.n15 163.367
R2125 B.n831 B.n830 163.367
R2126 B.n832 B.n831 163.367
R2127 B.n832 B.n13 163.367
R2128 B.n836 B.n13 163.367
R2129 B.n837 B.n836 163.367
R2130 B.n838 B.n837 163.367
R2131 B.n838 B.n11 163.367
R2132 B.n842 B.n11 163.367
R2133 B.n843 B.n842 163.367
R2134 B.n844 B.n843 163.367
R2135 B.n844 B.n9 163.367
R2136 B.n848 B.n9 163.367
R2137 B.n849 B.n848 163.367
R2138 B.n850 B.n849 163.367
R2139 B.n850 B.n7 163.367
R2140 B.n854 B.n7 163.367
R2141 B.n855 B.n854 163.367
R2142 B.n856 B.n855 163.367
R2143 B.n856 B.n5 163.367
R2144 B.n860 B.n5 163.367
R2145 B.n861 B.n860 163.367
R2146 B.n862 B.n861 163.367
R2147 B.n862 B.n3 163.367
R2148 B.n866 B.n3 163.367
R2149 B.n867 B.n866 163.367
R2150 B.n221 B.n2 163.367
R2151 B.n224 B.n221 163.367
R2152 B.n225 B.n224 163.367
R2153 B.n226 B.n225 163.367
R2154 B.n226 B.n219 163.367
R2155 B.n230 B.n219 163.367
R2156 B.n231 B.n230 163.367
R2157 B.n232 B.n231 163.367
R2158 B.n232 B.n217 163.367
R2159 B.n236 B.n217 163.367
R2160 B.n237 B.n236 163.367
R2161 B.n238 B.n237 163.367
R2162 B.n238 B.n215 163.367
R2163 B.n242 B.n215 163.367
R2164 B.n243 B.n242 163.367
R2165 B.n244 B.n243 163.367
R2166 B.n244 B.n213 163.367
R2167 B.n248 B.n213 163.367
R2168 B.n249 B.n248 163.367
R2169 B.n250 B.n249 163.367
R2170 B.n250 B.n211 163.367
R2171 B.n254 B.n211 163.367
R2172 B.n255 B.n254 163.367
R2173 B.n256 B.n255 163.367
R2174 B.n256 B.n209 163.367
R2175 B.n260 B.n209 163.367
R2176 B.n261 B.n260 163.367
R2177 B.n262 B.n261 163.367
R2178 B.n262 B.n207 163.367
R2179 B.n266 B.n207 163.367
R2180 B.n267 B.n266 163.367
R2181 B.n268 B.n267 163.367
R2182 B.n268 B.n205 163.367
R2183 B.n272 B.n205 163.367
R2184 B.n273 B.n272 163.367
R2185 B.n274 B.n273 163.367
R2186 B.n274 B.n203 163.367
R2187 B.n278 B.n203 163.367
R2188 B.n279 B.n278 163.367
R2189 B.n280 B.n279 163.367
R2190 B.n280 B.n201 163.367
R2191 B.n284 B.n201 163.367
R2192 B.n285 B.n284 163.367
R2193 B.n286 B.n285 163.367
R2194 B.n286 B.n199 163.367
R2195 B.n290 B.n199 163.367
R2196 B.n291 B.n290 163.367
R2197 B.n292 B.n291 163.367
R2198 B.n292 B.n197 163.367
R2199 B.n373 B.n171 59.5399
R2200 B.n388 B.n387 59.5399
R2201 B.n700 B.n61 59.5399
R2202 B.n714 B.n55 59.5399
R2203 B.n171 B.n170 46.546
R2204 B.n387 B.n386 46.546
R2205 B.n61 B.n60 46.546
R2206 B.n55 B.n54 46.546
R2207 B.n793 B.n792 32.0005
R2208 B.n622 B.n621 32.0005
R2209 B.n467 B.n138 32.0005
R2210 B.n295 B.n294 32.0005
R2211 B B.n869 18.0485
R2212 B.n793 B.n26 10.6151
R2213 B.n797 B.n26 10.6151
R2214 B.n798 B.n797 10.6151
R2215 B.n799 B.n798 10.6151
R2216 B.n799 B.n24 10.6151
R2217 B.n803 B.n24 10.6151
R2218 B.n804 B.n803 10.6151
R2219 B.n805 B.n804 10.6151
R2220 B.n805 B.n22 10.6151
R2221 B.n809 B.n22 10.6151
R2222 B.n810 B.n809 10.6151
R2223 B.n811 B.n810 10.6151
R2224 B.n811 B.n20 10.6151
R2225 B.n815 B.n20 10.6151
R2226 B.n816 B.n815 10.6151
R2227 B.n817 B.n816 10.6151
R2228 B.n817 B.n18 10.6151
R2229 B.n821 B.n18 10.6151
R2230 B.n822 B.n821 10.6151
R2231 B.n823 B.n822 10.6151
R2232 B.n823 B.n16 10.6151
R2233 B.n827 B.n16 10.6151
R2234 B.n828 B.n827 10.6151
R2235 B.n829 B.n828 10.6151
R2236 B.n829 B.n14 10.6151
R2237 B.n833 B.n14 10.6151
R2238 B.n834 B.n833 10.6151
R2239 B.n835 B.n834 10.6151
R2240 B.n835 B.n12 10.6151
R2241 B.n839 B.n12 10.6151
R2242 B.n840 B.n839 10.6151
R2243 B.n841 B.n840 10.6151
R2244 B.n841 B.n10 10.6151
R2245 B.n845 B.n10 10.6151
R2246 B.n846 B.n845 10.6151
R2247 B.n847 B.n846 10.6151
R2248 B.n847 B.n8 10.6151
R2249 B.n851 B.n8 10.6151
R2250 B.n852 B.n851 10.6151
R2251 B.n853 B.n852 10.6151
R2252 B.n853 B.n6 10.6151
R2253 B.n857 B.n6 10.6151
R2254 B.n858 B.n857 10.6151
R2255 B.n859 B.n858 10.6151
R2256 B.n859 B.n4 10.6151
R2257 B.n863 B.n4 10.6151
R2258 B.n864 B.n863 10.6151
R2259 B.n865 B.n864 10.6151
R2260 B.n865 B.n0 10.6151
R2261 B.n792 B.n791 10.6151
R2262 B.n791 B.n28 10.6151
R2263 B.n787 B.n28 10.6151
R2264 B.n787 B.n786 10.6151
R2265 B.n786 B.n785 10.6151
R2266 B.n785 B.n30 10.6151
R2267 B.n781 B.n30 10.6151
R2268 B.n781 B.n780 10.6151
R2269 B.n780 B.n779 10.6151
R2270 B.n779 B.n32 10.6151
R2271 B.n775 B.n32 10.6151
R2272 B.n775 B.n774 10.6151
R2273 B.n774 B.n773 10.6151
R2274 B.n773 B.n34 10.6151
R2275 B.n769 B.n34 10.6151
R2276 B.n769 B.n768 10.6151
R2277 B.n768 B.n767 10.6151
R2278 B.n767 B.n36 10.6151
R2279 B.n763 B.n36 10.6151
R2280 B.n763 B.n762 10.6151
R2281 B.n762 B.n761 10.6151
R2282 B.n761 B.n38 10.6151
R2283 B.n757 B.n38 10.6151
R2284 B.n757 B.n756 10.6151
R2285 B.n756 B.n755 10.6151
R2286 B.n755 B.n40 10.6151
R2287 B.n751 B.n40 10.6151
R2288 B.n751 B.n750 10.6151
R2289 B.n750 B.n749 10.6151
R2290 B.n749 B.n42 10.6151
R2291 B.n745 B.n42 10.6151
R2292 B.n745 B.n744 10.6151
R2293 B.n744 B.n743 10.6151
R2294 B.n743 B.n44 10.6151
R2295 B.n739 B.n44 10.6151
R2296 B.n739 B.n738 10.6151
R2297 B.n738 B.n737 10.6151
R2298 B.n737 B.n46 10.6151
R2299 B.n733 B.n46 10.6151
R2300 B.n733 B.n732 10.6151
R2301 B.n732 B.n731 10.6151
R2302 B.n731 B.n48 10.6151
R2303 B.n727 B.n48 10.6151
R2304 B.n727 B.n726 10.6151
R2305 B.n726 B.n725 10.6151
R2306 B.n725 B.n50 10.6151
R2307 B.n721 B.n50 10.6151
R2308 B.n721 B.n720 10.6151
R2309 B.n720 B.n719 10.6151
R2310 B.n719 B.n52 10.6151
R2311 B.n715 B.n52 10.6151
R2312 B.n713 B.n712 10.6151
R2313 B.n712 B.n56 10.6151
R2314 B.n708 B.n56 10.6151
R2315 B.n708 B.n707 10.6151
R2316 B.n707 B.n706 10.6151
R2317 B.n706 B.n58 10.6151
R2318 B.n702 B.n58 10.6151
R2319 B.n702 B.n701 10.6151
R2320 B.n699 B.n62 10.6151
R2321 B.n695 B.n62 10.6151
R2322 B.n695 B.n694 10.6151
R2323 B.n694 B.n693 10.6151
R2324 B.n693 B.n64 10.6151
R2325 B.n689 B.n64 10.6151
R2326 B.n689 B.n688 10.6151
R2327 B.n688 B.n687 10.6151
R2328 B.n687 B.n66 10.6151
R2329 B.n683 B.n66 10.6151
R2330 B.n683 B.n682 10.6151
R2331 B.n682 B.n681 10.6151
R2332 B.n681 B.n68 10.6151
R2333 B.n677 B.n68 10.6151
R2334 B.n677 B.n676 10.6151
R2335 B.n676 B.n675 10.6151
R2336 B.n675 B.n70 10.6151
R2337 B.n671 B.n70 10.6151
R2338 B.n671 B.n670 10.6151
R2339 B.n670 B.n669 10.6151
R2340 B.n669 B.n72 10.6151
R2341 B.n665 B.n72 10.6151
R2342 B.n665 B.n664 10.6151
R2343 B.n664 B.n663 10.6151
R2344 B.n663 B.n74 10.6151
R2345 B.n659 B.n74 10.6151
R2346 B.n659 B.n658 10.6151
R2347 B.n658 B.n657 10.6151
R2348 B.n657 B.n76 10.6151
R2349 B.n653 B.n76 10.6151
R2350 B.n653 B.n652 10.6151
R2351 B.n652 B.n651 10.6151
R2352 B.n651 B.n78 10.6151
R2353 B.n647 B.n78 10.6151
R2354 B.n647 B.n646 10.6151
R2355 B.n646 B.n645 10.6151
R2356 B.n645 B.n80 10.6151
R2357 B.n641 B.n80 10.6151
R2358 B.n641 B.n640 10.6151
R2359 B.n640 B.n639 10.6151
R2360 B.n639 B.n82 10.6151
R2361 B.n635 B.n82 10.6151
R2362 B.n635 B.n634 10.6151
R2363 B.n634 B.n633 10.6151
R2364 B.n633 B.n84 10.6151
R2365 B.n629 B.n84 10.6151
R2366 B.n629 B.n628 10.6151
R2367 B.n628 B.n627 10.6151
R2368 B.n627 B.n86 10.6151
R2369 B.n623 B.n86 10.6151
R2370 B.n623 B.n622 10.6151
R2371 B.n621 B.n88 10.6151
R2372 B.n617 B.n88 10.6151
R2373 B.n617 B.n616 10.6151
R2374 B.n616 B.n615 10.6151
R2375 B.n615 B.n90 10.6151
R2376 B.n611 B.n90 10.6151
R2377 B.n611 B.n610 10.6151
R2378 B.n610 B.n609 10.6151
R2379 B.n609 B.n92 10.6151
R2380 B.n605 B.n92 10.6151
R2381 B.n605 B.n604 10.6151
R2382 B.n604 B.n603 10.6151
R2383 B.n603 B.n94 10.6151
R2384 B.n599 B.n94 10.6151
R2385 B.n599 B.n598 10.6151
R2386 B.n598 B.n597 10.6151
R2387 B.n597 B.n96 10.6151
R2388 B.n593 B.n96 10.6151
R2389 B.n593 B.n592 10.6151
R2390 B.n592 B.n591 10.6151
R2391 B.n591 B.n98 10.6151
R2392 B.n587 B.n98 10.6151
R2393 B.n587 B.n586 10.6151
R2394 B.n586 B.n585 10.6151
R2395 B.n585 B.n100 10.6151
R2396 B.n581 B.n100 10.6151
R2397 B.n581 B.n580 10.6151
R2398 B.n580 B.n579 10.6151
R2399 B.n579 B.n102 10.6151
R2400 B.n575 B.n102 10.6151
R2401 B.n575 B.n574 10.6151
R2402 B.n574 B.n573 10.6151
R2403 B.n573 B.n104 10.6151
R2404 B.n569 B.n104 10.6151
R2405 B.n569 B.n568 10.6151
R2406 B.n568 B.n567 10.6151
R2407 B.n567 B.n106 10.6151
R2408 B.n563 B.n106 10.6151
R2409 B.n563 B.n562 10.6151
R2410 B.n562 B.n561 10.6151
R2411 B.n561 B.n108 10.6151
R2412 B.n557 B.n108 10.6151
R2413 B.n557 B.n556 10.6151
R2414 B.n556 B.n555 10.6151
R2415 B.n555 B.n110 10.6151
R2416 B.n551 B.n110 10.6151
R2417 B.n551 B.n550 10.6151
R2418 B.n550 B.n549 10.6151
R2419 B.n549 B.n112 10.6151
R2420 B.n545 B.n112 10.6151
R2421 B.n545 B.n544 10.6151
R2422 B.n544 B.n543 10.6151
R2423 B.n543 B.n114 10.6151
R2424 B.n539 B.n114 10.6151
R2425 B.n539 B.n538 10.6151
R2426 B.n538 B.n537 10.6151
R2427 B.n537 B.n116 10.6151
R2428 B.n533 B.n116 10.6151
R2429 B.n533 B.n532 10.6151
R2430 B.n532 B.n531 10.6151
R2431 B.n531 B.n118 10.6151
R2432 B.n527 B.n118 10.6151
R2433 B.n527 B.n526 10.6151
R2434 B.n526 B.n525 10.6151
R2435 B.n525 B.n120 10.6151
R2436 B.n521 B.n120 10.6151
R2437 B.n521 B.n520 10.6151
R2438 B.n520 B.n519 10.6151
R2439 B.n519 B.n122 10.6151
R2440 B.n515 B.n122 10.6151
R2441 B.n515 B.n514 10.6151
R2442 B.n514 B.n513 10.6151
R2443 B.n513 B.n124 10.6151
R2444 B.n509 B.n124 10.6151
R2445 B.n509 B.n508 10.6151
R2446 B.n508 B.n507 10.6151
R2447 B.n507 B.n126 10.6151
R2448 B.n503 B.n126 10.6151
R2449 B.n503 B.n502 10.6151
R2450 B.n502 B.n501 10.6151
R2451 B.n501 B.n128 10.6151
R2452 B.n497 B.n128 10.6151
R2453 B.n497 B.n496 10.6151
R2454 B.n496 B.n495 10.6151
R2455 B.n495 B.n130 10.6151
R2456 B.n491 B.n130 10.6151
R2457 B.n491 B.n490 10.6151
R2458 B.n490 B.n489 10.6151
R2459 B.n489 B.n132 10.6151
R2460 B.n485 B.n132 10.6151
R2461 B.n485 B.n484 10.6151
R2462 B.n484 B.n483 10.6151
R2463 B.n483 B.n134 10.6151
R2464 B.n479 B.n134 10.6151
R2465 B.n479 B.n478 10.6151
R2466 B.n478 B.n477 10.6151
R2467 B.n477 B.n136 10.6151
R2468 B.n473 B.n136 10.6151
R2469 B.n473 B.n472 10.6151
R2470 B.n472 B.n471 10.6151
R2471 B.n471 B.n138 10.6151
R2472 B.n222 B.n1 10.6151
R2473 B.n223 B.n222 10.6151
R2474 B.n223 B.n220 10.6151
R2475 B.n227 B.n220 10.6151
R2476 B.n228 B.n227 10.6151
R2477 B.n229 B.n228 10.6151
R2478 B.n229 B.n218 10.6151
R2479 B.n233 B.n218 10.6151
R2480 B.n234 B.n233 10.6151
R2481 B.n235 B.n234 10.6151
R2482 B.n235 B.n216 10.6151
R2483 B.n239 B.n216 10.6151
R2484 B.n240 B.n239 10.6151
R2485 B.n241 B.n240 10.6151
R2486 B.n241 B.n214 10.6151
R2487 B.n245 B.n214 10.6151
R2488 B.n246 B.n245 10.6151
R2489 B.n247 B.n246 10.6151
R2490 B.n247 B.n212 10.6151
R2491 B.n251 B.n212 10.6151
R2492 B.n252 B.n251 10.6151
R2493 B.n253 B.n252 10.6151
R2494 B.n253 B.n210 10.6151
R2495 B.n257 B.n210 10.6151
R2496 B.n258 B.n257 10.6151
R2497 B.n259 B.n258 10.6151
R2498 B.n259 B.n208 10.6151
R2499 B.n263 B.n208 10.6151
R2500 B.n264 B.n263 10.6151
R2501 B.n265 B.n264 10.6151
R2502 B.n265 B.n206 10.6151
R2503 B.n269 B.n206 10.6151
R2504 B.n270 B.n269 10.6151
R2505 B.n271 B.n270 10.6151
R2506 B.n271 B.n204 10.6151
R2507 B.n275 B.n204 10.6151
R2508 B.n276 B.n275 10.6151
R2509 B.n277 B.n276 10.6151
R2510 B.n277 B.n202 10.6151
R2511 B.n281 B.n202 10.6151
R2512 B.n282 B.n281 10.6151
R2513 B.n283 B.n282 10.6151
R2514 B.n283 B.n200 10.6151
R2515 B.n287 B.n200 10.6151
R2516 B.n288 B.n287 10.6151
R2517 B.n289 B.n288 10.6151
R2518 B.n289 B.n198 10.6151
R2519 B.n293 B.n198 10.6151
R2520 B.n294 B.n293 10.6151
R2521 B.n295 B.n196 10.6151
R2522 B.n299 B.n196 10.6151
R2523 B.n300 B.n299 10.6151
R2524 B.n301 B.n300 10.6151
R2525 B.n301 B.n194 10.6151
R2526 B.n305 B.n194 10.6151
R2527 B.n306 B.n305 10.6151
R2528 B.n307 B.n306 10.6151
R2529 B.n307 B.n192 10.6151
R2530 B.n311 B.n192 10.6151
R2531 B.n312 B.n311 10.6151
R2532 B.n313 B.n312 10.6151
R2533 B.n313 B.n190 10.6151
R2534 B.n317 B.n190 10.6151
R2535 B.n318 B.n317 10.6151
R2536 B.n319 B.n318 10.6151
R2537 B.n319 B.n188 10.6151
R2538 B.n323 B.n188 10.6151
R2539 B.n324 B.n323 10.6151
R2540 B.n325 B.n324 10.6151
R2541 B.n325 B.n186 10.6151
R2542 B.n329 B.n186 10.6151
R2543 B.n330 B.n329 10.6151
R2544 B.n331 B.n330 10.6151
R2545 B.n331 B.n184 10.6151
R2546 B.n335 B.n184 10.6151
R2547 B.n336 B.n335 10.6151
R2548 B.n337 B.n336 10.6151
R2549 B.n337 B.n182 10.6151
R2550 B.n341 B.n182 10.6151
R2551 B.n342 B.n341 10.6151
R2552 B.n343 B.n342 10.6151
R2553 B.n343 B.n180 10.6151
R2554 B.n347 B.n180 10.6151
R2555 B.n348 B.n347 10.6151
R2556 B.n349 B.n348 10.6151
R2557 B.n349 B.n178 10.6151
R2558 B.n353 B.n178 10.6151
R2559 B.n354 B.n353 10.6151
R2560 B.n355 B.n354 10.6151
R2561 B.n355 B.n176 10.6151
R2562 B.n359 B.n176 10.6151
R2563 B.n360 B.n359 10.6151
R2564 B.n361 B.n360 10.6151
R2565 B.n361 B.n174 10.6151
R2566 B.n365 B.n174 10.6151
R2567 B.n366 B.n365 10.6151
R2568 B.n367 B.n366 10.6151
R2569 B.n367 B.n172 10.6151
R2570 B.n371 B.n172 10.6151
R2571 B.n372 B.n371 10.6151
R2572 B.n374 B.n168 10.6151
R2573 B.n378 B.n168 10.6151
R2574 B.n379 B.n378 10.6151
R2575 B.n380 B.n379 10.6151
R2576 B.n380 B.n166 10.6151
R2577 B.n384 B.n166 10.6151
R2578 B.n385 B.n384 10.6151
R2579 B.n389 B.n385 10.6151
R2580 B.n393 B.n164 10.6151
R2581 B.n394 B.n393 10.6151
R2582 B.n395 B.n394 10.6151
R2583 B.n395 B.n162 10.6151
R2584 B.n399 B.n162 10.6151
R2585 B.n400 B.n399 10.6151
R2586 B.n401 B.n400 10.6151
R2587 B.n401 B.n160 10.6151
R2588 B.n405 B.n160 10.6151
R2589 B.n406 B.n405 10.6151
R2590 B.n407 B.n406 10.6151
R2591 B.n407 B.n158 10.6151
R2592 B.n411 B.n158 10.6151
R2593 B.n412 B.n411 10.6151
R2594 B.n413 B.n412 10.6151
R2595 B.n413 B.n156 10.6151
R2596 B.n417 B.n156 10.6151
R2597 B.n418 B.n417 10.6151
R2598 B.n419 B.n418 10.6151
R2599 B.n419 B.n154 10.6151
R2600 B.n423 B.n154 10.6151
R2601 B.n424 B.n423 10.6151
R2602 B.n425 B.n424 10.6151
R2603 B.n425 B.n152 10.6151
R2604 B.n429 B.n152 10.6151
R2605 B.n430 B.n429 10.6151
R2606 B.n431 B.n430 10.6151
R2607 B.n431 B.n150 10.6151
R2608 B.n435 B.n150 10.6151
R2609 B.n436 B.n435 10.6151
R2610 B.n437 B.n436 10.6151
R2611 B.n437 B.n148 10.6151
R2612 B.n441 B.n148 10.6151
R2613 B.n442 B.n441 10.6151
R2614 B.n443 B.n442 10.6151
R2615 B.n443 B.n146 10.6151
R2616 B.n447 B.n146 10.6151
R2617 B.n448 B.n447 10.6151
R2618 B.n449 B.n448 10.6151
R2619 B.n449 B.n144 10.6151
R2620 B.n453 B.n144 10.6151
R2621 B.n454 B.n453 10.6151
R2622 B.n455 B.n454 10.6151
R2623 B.n455 B.n142 10.6151
R2624 B.n459 B.n142 10.6151
R2625 B.n460 B.n459 10.6151
R2626 B.n461 B.n460 10.6151
R2627 B.n461 B.n140 10.6151
R2628 B.n465 B.n140 10.6151
R2629 B.n466 B.n465 10.6151
R2630 B.n467 B.n466 10.6151
R2631 B.n869 B.n0 8.11757
R2632 B.n869 B.n1 8.11757
R2633 B.n714 B.n713 6.5566
R2634 B.n701 B.n700 6.5566
R2635 B.n374 B.n373 6.5566
R2636 B.n389 B.n388 6.5566
R2637 B.n715 B.n714 4.05904
R2638 B.n700 B.n699 4.05904
R2639 B.n373 B.n372 4.05904
R2640 B.n388 B.n164 4.05904
C0 VN VDD2 12.896099f
C1 VTAIL VDD1 12.196099f
C2 VDD1 B 2.53882f
C3 w_n3850_n4054# VDD2 2.9449f
C4 VP VDD1 13.2556f
C5 VTAIL B 4.23549f
C6 VN VDD1 0.152175f
C7 VP VTAIL 13.186f
C8 VN VTAIL 13.171599f
C9 VP B 2.02603f
C10 VDD1 w_n3850_n4054# 2.8288f
C11 VDD1 VDD2 1.83026f
C12 VN B 1.18882f
C13 VP VN 8.25634f
C14 VTAIL w_n3850_n4054# 3.63226f
C15 VTAIL VDD2 12.241799f
C16 w_n3850_n4054# B 10.6171f
C17 B VDD2 2.6361f
C18 VP w_n3850_n4054# 8.64546f
C19 VP VDD2 0.516345f
C20 VN w_n3850_n4054# 8.14584f
C21 VDD2 VSUBS 2.00076f
C22 VDD1 VSUBS 1.826988f
C23 VTAIL VSUBS 1.293141f
C24 VN VSUBS 6.97048f
C25 VP VSUBS 3.690576f
C26 B VSUBS 4.99833f
C27 w_n3850_n4054# VSUBS 0.191314p
C28 B.n0 VSUBS 0.007781f
C29 B.n1 VSUBS 0.007781f
C30 B.n2 VSUBS 0.011507f
C31 B.n3 VSUBS 0.008818f
C32 B.n4 VSUBS 0.008818f
C33 B.n5 VSUBS 0.008818f
C34 B.n6 VSUBS 0.008818f
C35 B.n7 VSUBS 0.008818f
C36 B.n8 VSUBS 0.008818f
C37 B.n9 VSUBS 0.008818f
C38 B.n10 VSUBS 0.008818f
C39 B.n11 VSUBS 0.008818f
C40 B.n12 VSUBS 0.008818f
C41 B.n13 VSUBS 0.008818f
C42 B.n14 VSUBS 0.008818f
C43 B.n15 VSUBS 0.008818f
C44 B.n16 VSUBS 0.008818f
C45 B.n17 VSUBS 0.008818f
C46 B.n18 VSUBS 0.008818f
C47 B.n19 VSUBS 0.008818f
C48 B.n20 VSUBS 0.008818f
C49 B.n21 VSUBS 0.008818f
C50 B.n22 VSUBS 0.008818f
C51 B.n23 VSUBS 0.008818f
C52 B.n24 VSUBS 0.008818f
C53 B.n25 VSUBS 0.008818f
C54 B.n26 VSUBS 0.008818f
C55 B.n27 VSUBS 0.02084f
C56 B.n28 VSUBS 0.008818f
C57 B.n29 VSUBS 0.008818f
C58 B.n30 VSUBS 0.008818f
C59 B.n31 VSUBS 0.008818f
C60 B.n32 VSUBS 0.008818f
C61 B.n33 VSUBS 0.008818f
C62 B.n34 VSUBS 0.008818f
C63 B.n35 VSUBS 0.008818f
C64 B.n36 VSUBS 0.008818f
C65 B.n37 VSUBS 0.008818f
C66 B.n38 VSUBS 0.008818f
C67 B.n39 VSUBS 0.008818f
C68 B.n40 VSUBS 0.008818f
C69 B.n41 VSUBS 0.008818f
C70 B.n42 VSUBS 0.008818f
C71 B.n43 VSUBS 0.008818f
C72 B.n44 VSUBS 0.008818f
C73 B.n45 VSUBS 0.008818f
C74 B.n46 VSUBS 0.008818f
C75 B.n47 VSUBS 0.008818f
C76 B.n48 VSUBS 0.008818f
C77 B.n49 VSUBS 0.008818f
C78 B.n50 VSUBS 0.008818f
C79 B.n51 VSUBS 0.008818f
C80 B.n52 VSUBS 0.008818f
C81 B.n53 VSUBS 0.008818f
C82 B.t4 VSUBS 0.364886f
C83 B.t5 VSUBS 0.399426f
C84 B.t3 VSUBS 1.77303f
C85 B.n54 VSUBS 0.603933f
C86 B.n55 VSUBS 0.371658f
C87 B.n56 VSUBS 0.008818f
C88 B.n57 VSUBS 0.008818f
C89 B.n58 VSUBS 0.008818f
C90 B.n59 VSUBS 0.008818f
C91 B.t1 VSUBS 0.36489f
C92 B.t2 VSUBS 0.399429f
C93 B.t0 VSUBS 1.77303f
C94 B.n60 VSUBS 0.603929f
C95 B.n61 VSUBS 0.371653f
C96 B.n62 VSUBS 0.008818f
C97 B.n63 VSUBS 0.008818f
C98 B.n64 VSUBS 0.008818f
C99 B.n65 VSUBS 0.008818f
C100 B.n66 VSUBS 0.008818f
C101 B.n67 VSUBS 0.008818f
C102 B.n68 VSUBS 0.008818f
C103 B.n69 VSUBS 0.008818f
C104 B.n70 VSUBS 0.008818f
C105 B.n71 VSUBS 0.008818f
C106 B.n72 VSUBS 0.008818f
C107 B.n73 VSUBS 0.008818f
C108 B.n74 VSUBS 0.008818f
C109 B.n75 VSUBS 0.008818f
C110 B.n76 VSUBS 0.008818f
C111 B.n77 VSUBS 0.008818f
C112 B.n78 VSUBS 0.008818f
C113 B.n79 VSUBS 0.008818f
C114 B.n80 VSUBS 0.008818f
C115 B.n81 VSUBS 0.008818f
C116 B.n82 VSUBS 0.008818f
C117 B.n83 VSUBS 0.008818f
C118 B.n84 VSUBS 0.008818f
C119 B.n85 VSUBS 0.008818f
C120 B.n86 VSUBS 0.008818f
C121 B.n87 VSUBS 0.02084f
C122 B.n88 VSUBS 0.008818f
C123 B.n89 VSUBS 0.008818f
C124 B.n90 VSUBS 0.008818f
C125 B.n91 VSUBS 0.008818f
C126 B.n92 VSUBS 0.008818f
C127 B.n93 VSUBS 0.008818f
C128 B.n94 VSUBS 0.008818f
C129 B.n95 VSUBS 0.008818f
C130 B.n96 VSUBS 0.008818f
C131 B.n97 VSUBS 0.008818f
C132 B.n98 VSUBS 0.008818f
C133 B.n99 VSUBS 0.008818f
C134 B.n100 VSUBS 0.008818f
C135 B.n101 VSUBS 0.008818f
C136 B.n102 VSUBS 0.008818f
C137 B.n103 VSUBS 0.008818f
C138 B.n104 VSUBS 0.008818f
C139 B.n105 VSUBS 0.008818f
C140 B.n106 VSUBS 0.008818f
C141 B.n107 VSUBS 0.008818f
C142 B.n108 VSUBS 0.008818f
C143 B.n109 VSUBS 0.008818f
C144 B.n110 VSUBS 0.008818f
C145 B.n111 VSUBS 0.008818f
C146 B.n112 VSUBS 0.008818f
C147 B.n113 VSUBS 0.008818f
C148 B.n114 VSUBS 0.008818f
C149 B.n115 VSUBS 0.008818f
C150 B.n116 VSUBS 0.008818f
C151 B.n117 VSUBS 0.008818f
C152 B.n118 VSUBS 0.008818f
C153 B.n119 VSUBS 0.008818f
C154 B.n120 VSUBS 0.008818f
C155 B.n121 VSUBS 0.008818f
C156 B.n122 VSUBS 0.008818f
C157 B.n123 VSUBS 0.008818f
C158 B.n124 VSUBS 0.008818f
C159 B.n125 VSUBS 0.008818f
C160 B.n126 VSUBS 0.008818f
C161 B.n127 VSUBS 0.008818f
C162 B.n128 VSUBS 0.008818f
C163 B.n129 VSUBS 0.008818f
C164 B.n130 VSUBS 0.008818f
C165 B.n131 VSUBS 0.008818f
C166 B.n132 VSUBS 0.008818f
C167 B.n133 VSUBS 0.008818f
C168 B.n134 VSUBS 0.008818f
C169 B.n135 VSUBS 0.008818f
C170 B.n136 VSUBS 0.008818f
C171 B.n137 VSUBS 0.008818f
C172 B.n138 VSUBS 0.020943f
C173 B.n139 VSUBS 0.008818f
C174 B.n140 VSUBS 0.008818f
C175 B.n141 VSUBS 0.008818f
C176 B.n142 VSUBS 0.008818f
C177 B.n143 VSUBS 0.008818f
C178 B.n144 VSUBS 0.008818f
C179 B.n145 VSUBS 0.008818f
C180 B.n146 VSUBS 0.008818f
C181 B.n147 VSUBS 0.008818f
C182 B.n148 VSUBS 0.008818f
C183 B.n149 VSUBS 0.008818f
C184 B.n150 VSUBS 0.008818f
C185 B.n151 VSUBS 0.008818f
C186 B.n152 VSUBS 0.008818f
C187 B.n153 VSUBS 0.008818f
C188 B.n154 VSUBS 0.008818f
C189 B.n155 VSUBS 0.008818f
C190 B.n156 VSUBS 0.008818f
C191 B.n157 VSUBS 0.008818f
C192 B.n158 VSUBS 0.008818f
C193 B.n159 VSUBS 0.008818f
C194 B.n160 VSUBS 0.008818f
C195 B.n161 VSUBS 0.008818f
C196 B.n162 VSUBS 0.008818f
C197 B.n163 VSUBS 0.008818f
C198 B.n164 VSUBS 0.006095f
C199 B.n165 VSUBS 0.008818f
C200 B.n166 VSUBS 0.008818f
C201 B.n167 VSUBS 0.008818f
C202 B.n168 VSUBS 0.008818f
C203 B.n169 VSUBS 0.008818f
C204 B.t11 VSUBS 0.364886f
C205 B.t10 VSUBS 0.399426f
C206 B.t9 VSUBS 1.77303f
C207 B.n170 VSUBS 0.603933f
C208 B.n171 VSUBS 0.371658f
C209 B.n172 VSUBS 0.008818f
C210 B.n173 VSUBS 0.008818f
C211 B.n174 VSUBS 0.008818f
C212 B.n175 VSUBS 0.008818f
C213 B.n176 VSUBS 0.008818f
C214 B.n177 VSUBS 0.008818f
C215 B.n178 VSUBS 0.008818f
C216 B.n179 VSUBS 0.008818f
C217 B.n180 VSUBS 0.008818f
C218 B.n181 VSUBS 0.008818f
C219 B.n182 VSUBS 0.008818f
C220 B.n183 VSUBS 0.008818f
C221 B.n184 VSUBS 0.008818f
C222 B.n185 VSUBS 0.008818f
C223 B.n186 VSUBS 0.008818f
C224 B.n187 VSUBS 0.008818f
C225 B.n188 VSUBS 0.008818f
C226 B.n189 VSUBS 0.008818f
C227 B.n190 VSUBS 0.008818f
C228 B.n191 VSUBS 0.008818f
C229 B.n192 VSUBS 0.008818f
C230 B.n193 VSUBS 0.008818f
C231 B.n194 VSUBS 0.008818f
C232 B.n195 VSUBS 0.008818f
C233 B.n196 VSUBS 0.008818f
C234 B.n197 VSUBS 0.01988f
C235 B.n198 VSUBS 0.008818f
C236 B.n199 VSUBS 0.008818f
C237 B.n200 VSUBS 0.008818f
C238 B.n201 VSUBS 0.008818f
C239 B.n202 VSUBS 0.008818f
C240 B.n203 VSUBS 0.008818f
C241 B.n204 VSUBS 0.008818f
C242 B.n205 VSUBS 0.008818f
C243 B.n206 VSUBS 0.008818f
C244 B.n207 VSUBS 0.008818f
C245 B.n208 VSUBS 0.008818f
C246 B.n209 VSUBS 0.008818f
C247 B.n210 VSUBS 0.008818f
C248 B.n211 VSUBS 0.008818f
C249 B.n212 VSUBS 0.008818f
C250 B.n213 VSUBS 0.008818f
C251 B.n214 VSUBS 0.008818f
C252 B.n215 VSUBS 0.008818f
C253 B.n216 VSUBS 0.008818f
C254 B.n217 VSUBS 0.008818f
C255 B.n218 VSUBS 0.008818f
C256 B.n219 VSUBS 0.008818f
C257 B.n220 VSUBS 0.008818f
C258 B.n221 VSUBS 0.008818f
C259 B.n222 VSUBS 0.008818f
C260 B.n223 VSUBS 0.008818f
C261 B.n224 VSUBS 0.008818f
C262 B.n225 VSUBS 0.008818f
C263 B.n226 VSUBS 0.008818f
C264 B.n227 VSUBS 0.008818f
C265 B.n228 VSUBS 0.008818f
C266 B.n229 VSUBS 0.008818f
C267 B.n230 VSUBS 0.008818f
C268 B.n231 VSUBS 0.008818f
C269 B.n232 VSUBS 0.008818f
C270 B.n233 VSUBS 0.008818f
C271 B.n234 VSUBS 0.008818f
C272 B.n235 VSUBS 0.008818f
C273 B.n236 VSUBS 0.008818f
C274 B.n237 VSUBS 0.008818f
C275 B.n238 VSUBS 0.008818f
C276 B.n239 VSUBS 0.008818f
C277 B.n240 VSUBS 0.008818f
C278 B.n241 VSUBS 0.008818f
C279 B.n242 VSUBS 0.008818f
C280 B.n243 VSUBS 0.008818f
C281 B.n244 VSUBS 0.008818f
C282 B.n245 VSUBS 0.008818f
C283 B.n246 VSUBS 0.008818f
C284 B.n247 VSUBS 0.008818f
C285 B.n248 VSUBS 0.008818f
C286 B.n249 VSUBS 0.008818f
C287 B.n250 VSUBS 0.008818f
C288 B.n251 VSUBS 0.008818f
C289 B.n252 VSUBS 0.008818f
C290 B.n253 VSUBS 0.008818f
C291 B.n254 VSUBS 0.008818f
C292 B.n255 VSUBS 0.008818f
C293 B.n256 VSUBS 0.008818f
C294 B.n257 VSUBS 0.008818f
C295 B.n258 VSUBS 0.008818f
C296 B.n259 VSUBS 0.008818f
C297 B.n260 VSUBS 0.008818f
C298 B.n261 VSUBS 0.008818f
C299 B.n262 VSUBS 0.008818f
C300 B.n263 VSUBS 0.008818f
C301 B.n264 VSUBS 0.008818f
C302 B.n265 VSUBS 0.008818f
C303 B.n266 VSUBS 0.008818f
C304 B.n267 VSUBS 0.008818f
C305 B.n268 VSUBS 0.008818f
C306 B.n269 VSUBS 0.008818f
C307 B.n270 VSUBS 0.008818f
C308 B.n271 VSUBS 0.008818f
C309 B.n272 VSUBS 0.008818f
C310 B.n273 VSUBS 0.008818f
C311 B.n274 VSUBS 0.008818f
C312 B.n275 VSUBS 0.008818f
C313 B.n276 VSUBS 0.008818f
C314 B.n277 VSUBS 0.008818f
C315 B.n278 VSUBS 0.008818f
C316 B.n279 VSUBS 0.008818f
C317 B.n280 VSUBS 0.008818f
C318 B.n281 VSUBS 0.008818f
C319 B.n282 VSUBS 0.008818f
C320 B.n283 VSUBS 0.008818f
C321 B.n284 VSUBS 0.008818f
C322 B.n285 VSUBS 0.008818f
C323 B.n286 VSUBS 0.008818f
C324 B.n287 VSUBS 0.008818f
C325 B.n288 VSUBS 0.008818f
C326 B.n289 VSUBS 0.008818f
C327 B.n290 VSUBS 0.008818f
C328 B.n291 VSUBS 0.008818f
C329 B.n292 VSUBS 0.008818f
C330 B.n293 VSUBS 0.008818f
C331 B.n294 VSUBS 0.01988f
C332 B.n295 VSUBS 0.02084f
C333 B.n296 VSUBS 0.02084f
C334 B.n297 VSUBS 0.008818f
C335 B.n298 VSUBS 0.008818f
C336 B.n299 VSUBS 0.008818f
C337 B.n300 VSUBS 0.008818f
C338 B.n301 VSUBS 0.008818f
C339 B.n302 VSUBS 0.008818f
C340 B.n303 VSUBS 0.008818f
C341 B.n304 VSUBS 0.008818f
C342 B.n305 VSUBS 0.008818f
C343 B.n306 VSUBS 0.008818f
C344 B.n307 VSUBS 0.008818f
C345 B.n308 VSUBS 0.008818f
C346 B.n309 VSUBS 0.008818f
C347 B.n310 VSUBS 0.008818f
C348 B.n311 VSUBS 0.008818f
C349 B.n312 VSUBS 0.008818f
C350 B.n313 VSUBS 0.008818f
C351 B.n314 VSUBS 0.008818f
C352 B.n315 VSUBS 0.008818f
C353 B.n316 VSUBS 0.008818f
C354 B.n317 VSUBS 0.008818f
C355 B.n318 VSUBS 0.008818f
C356 B.n319 VSUBS 0.008818f
C357 B.n320 VSUBS 0.008818f
C358 B.n321 VSUBS 0.008818f
C359 B.n322 VSUBS 0.008818f
C360 B.n323 VSUBS 0.008818f
C361 B.n324 VSUBS 0.008818f
C362 B.n325 VSUBS 0.008818f
C363 B.n326 VSUBS 0.008818f
C364 B.n327 VSUBS 0.008818f
C365 B.n328 VSUBS 0.008818f
C366 B.n329 VSUBS 0.008818f
C367 B.n330 VSUBS 0.008818f
C368 B.n331 VSUBS 0.008818f
C369 B.n332 VSUBS 0.008818f
C370 B.n333 VSUBS 0.008818f
C371 B.n334 VSUBS 0.008818f
C372 B.n335 VSUBS 0.008818f
C373 B.n336 VSUBS 0.008818f
C374 B.n337 VSUBS 0.008818f
C375 B.n338 VSUBS 0.008818f
C376 B.n339 VSUBS 0.008818f
C377 B.n340 VSUBS 0.008818f
C378 B.n341 VSUBS 0.008818f
C379 B.n342 VSUBS 0.008818f
C380 B.n343 VSUBS 0.008818f
C381 B.n344 VSUBS 0.008818f
C382 B.n345 VSUBS 0.008818f
C383 B.n346 VSUBS 0.008818f
C384 B.n347 VSUBS 0.008818f
C385 B.n348 VSUBS 0.008818f
C386 B.n349 VSUBS 0.008818f
C387 B.n350 VSUBS 0.008818f
C388 B.n351 VSUBS 0.008818f
C389 B.n352 VSUBS 0.008818f
C390 B.n353 VSUBS 0.008818f
C391 B.n354 VSUBS 0.008818f
C392 B.n355 VSUBS 0.008818f
C393 B.n356 VSUBS 0.008818f
C394 B.n357 VSUBS 0.008818f
C395 B.n358 VSUBS 0.008818f
C396 B.n359 VSUBS 0.008818f
C397 B.n360 VSUBS 0.008818f
C398 B.n361 VSUBS 0.008818f
C399 B.n362 VSUBS 0.008818f
C400 B.n363 VSUBS 0.008818f
C401 B.n364 VSUBS 0.008818f
C402 B.n365 VSUBS 0.008818f
C403 B.n366 VSUBS 0.008818f
C404 B.n367 VSUBS 0.008818f
C405 B.n368 VSUBS 0.008818f
C406 B.n369 VSUBS 0.008818f
C407 B.n370 VSUBS 0.008818f
C408 B.n371 VSUBS 0.008818f
C409 B.n372 VSUBS 0.006095f
C410 B.n373 VSUBS 0.020431f
C411 B.n374 VSUBS 0.007132f
C412 B.n375 VSUBS 0.008818f
C413 B.n376 VSUBS 0.008818f
C414 B.n377 VSUBS 0.008818f
C415 B.n378 VSUBS 0.008818f
C416 B.n379 VSUBS 0.008818f
C417 B.n380 VSUBS 0.008818f
C418 B.n381 VSUBS 0.008818f
C419 B.n382 VSUBS 0.008818f
C420 B.n383 VSUBS 0.008818f
C421 B.n384 VSUBS 0.008818f
C422 B.n385 VSUBS 0.008818f
C423 B.t8 VSUBS 0.36489f
C424 B.t7 VSUBS 0.399429f
C425 B.t6 VSUBS 1.77303f
C426 B.n386 VSUBS 0.603929f
C427 B.n387 VSUBS 0.371653f
C428 B.n388 VSUBS 0.020431f
C429 B.n389 VSUBS 0.007132f
C430 B.n390 VSUBS 0.008818f
C431 B.n391 VSUBS 0.008818f
C432 B.n392 VSUBS 0.008818f
C433 B.n393 VSUBS 0.008818f
C434 B.n394 VSUBS 0.008818f
C435 B.n395 VSUBS 0.008818f
C436 B.n396 VSUBS 0.008818f
C437 B.n397 VSUBS 0.008818f
C438 B.n398 VSUBS 0.008818f
C439 B.n399 VSUBS 0.008818f
C440 B.n400 VSUBS 0.008818f
C441 B.n401 VSUBS 0.008818f
C442 B.n402 VSUBS 0.008818f
C443 B.n403 VSUBS 0.008818f
C444 B.n404 VSUBS 0.008818f
C445 B.n405 VSUBS 0.008818f
C446 B.n406 VSUBS 0.008818f
C447 B.n407 VSUBS 0.008818f
C448 B.n408 VSUBS 0.008818f
C449 B.n409 VSUBS 0.008818f
C450 B.n410 VSUBS 0.008818f
C451 B.n411 VSUBS 0.008818f
C452 B.n412 VSUBS 0.008818f
C453 B.n413 VSUBS 0.008818f
C454 B.n414 VSUBS 0.008818f
C455 B.n415 VSUBS 0.008818f
C456 B.n416 VSUBS 0.008818f
C457 B.n417 VSUBS 0.008818f
C458 B.n418 VSUBS 0.008818f
C459 B.n419 VSUBS 0.008818f
C460 B.n420 VSUBS 0.008818f
C461 B.n421 VSUBS 0.008818f
C462 B.n422 VSUBS 0.008818f
C463 B.n423 VSUBS 0.008818f
C464 B.n424 VSUBS 0.008818f
C465 B.n425 VSUBS 0.008818f
C466 B.n426 VSUBS 0.008818f
C467 B.n427 VSUBS 0.008818f
C468 B.n428 VSUBS 0.008818f
C469 B.n429 VSUBS 0.008818f
C470 B.n430 VSUBS 0.008818f
C471 B.n431 VSUBS 0.008818f
C472 B.n432 VSUBS 0.008818f
C473 B.n433 VSUBS 0.008818f
C474 B.n434 VSUBS 0.008818f
C475 B.n435 VSUBS 0.008818f
C476 B.n436 VSUBS 0.008818f
C477 B.n437 VSUBS 0.008818f
C478 B.n438 VSUBS 0.008818f
C479 B.n439 VSUBS 0.008818f
C480 B.n440 VSUBS 0.008818f
C481 B.n441 VSUBS 0.008818f
C482 B.n442 VSUBS 0.008818f
C483 B.n443 VSUBS 0.008818f
C484 B.n444 VSUBS 0.008818f
C485 B.n445 VSUBS 0.008818f
C486 B.n446 VSUBS 0.008818f
C487 B.n447 VSUBS 0.008818f
C488 B.n448 VSUBS 0.008818f
C489 B.n449 VSUBS 0.008818f
C490 B.n450 VSUBS 0.008818f
C491 B.n451 VSUBS 0.008818f
C492 B.n452 VSUBS 0.008818f
C493 B.n453 VSUBS 0.008818f
C494 B.n454 VSUBS 0.008818f
C495 B.n455 VSUBS 0.008818f
C496 B.n456 VSUBS 0.008818f
C497 B.n457 VSUBS 0.008818f
C498 B.n458 VSUBS 0.008818f
C499 B.n459 VSUBS 0.008818f
C500 B.n460 VSUBS 0.008818f
C501 B.n461 VSUBS 0.008818f
C502 B.n462 VSUBS 0.008818f
C503 B.n463 VSUBS 0.008818f
C504 B.n464 VSUBS 0.008818f
C505 B.n465 VSUBS 0.008818f
C506 B.n466 VSUBS 0.008818f
C507 B.n467 VSUBS 0.019776f
C508 B.n468 VSUBS 0.02084f
C509 B.n469 VSUBS 0.01988f
C510 B.n470 VSUBS 0.008818f
C511 B.n471 VSUBS 0.008818f
C512 B.n472 VSUBS 0.008818f
C513 B.n473 VSUBS 0.008818f
C514 B.n474 VSUBS 0.008818f
C515 B.n475 VSUBS 0.008818f
C516 B.n476 VSUBS 0.008818f
C517 B.n477 VSUBS 0.008818f
C518 B.n478 VSUBS 0.008818f
C519 B.n479 VSUBS 0.008818f
C520 B.n480 VSUBS 0.008818f
C521 B.n481 VSUBS 0.008818f
C522 B.n482 VSUBS 0.008818f
C523 B.n483 VSUBS 0.008818f
C524 B.n484 VSUBS 0.008818f
C525 B.n485 VSUBS 0.008818f
C526 B.n486 VSUBS 0.008818f
C527 B.n487 VSUBS 0.008818f
C528 B.n488 VSUBS 0.008818f
C529 B.n489 VSUBS 0.008818f
C530 B.n490 VSUBS 0.008818f
C531 B.n491 VSUBS 0.008818f
C532 B.n492 VSUBS 0.008818f
C533 B.n493 VSUBS 0.008818f
C534 B.n494 VSUBS 0.008818f
C535 B.n495 VSUBS 0.008818f
C536 B.n496 VSUBS 0.008818f
C537 B.n497 VSUBS 0.008818f
C538 B.n498 VSUBS 0.008818f
C539 B.n499 VSUBS 0.008818f
C540 B.n500 VSUBS 0.008818f
C541 B.n501 VSUBS 0.008818f
C542 B.n502 VSUBS 0.008818f
C543 B.n503 VSUBS 0.008818f
C544 B.n504 VSUBS 0.008818f
C545 B.n505 VSUBS 0.008818f
C546 B.n506 VSUBS 0.008818f
C547 B.n507 VSUBS 0.008818f
C548 B.n508 VSUBS 0.008818f
C549 B.n509 VSUBS 0.008818f
C550 B.n510 VSUBS 0.008818f
C551 B.n511 VSUBS 0.008818f
C552 B.n512 VSUBS 0.008818f
C553 B.n513 VSUBS 0.008818f
C554 B.n514 VSUBS 0.008818f
C555 B.n515 VSUBS 0.008818f
C556 B.n516 VSUBS 0.008818f
C557 B.n517 VSUBS 0.008818f
C558 B.n518 VSUBS 0.008818f
C559 B.n519 VSUBS 0.008818f
C560 B.n520 VSUBS 0.008818f
C561 B.n521 VSUBS 0.008818f
C562 B.n522 VSUBS 0.008818f
C563 B.n523 VSUBS 0.008818f
C564 B.n524 VSUBS 0.008818f
C565 B.n525 VSUBS 0.008818f
C566 B.n526 VSUBS 0.008818f
C567 B.n527 VSUBS 0.008818f
C568 B.n528 VSUBS 0.008818f
C569 B.n529 VSUBS 0.008818f
C570 B.n530 VSUBS 0.008818f
C571 B.n531 VSUBS 0.008818f
C572 B.n532 VSUBS 0.008818f
C573 B.n533 VSUBS 0.008818f
C574 B.n534 VSUBS 0.008818f
C575 B.n535 VSUBS 0.008818f
C576 B.n536 VSUBS 0.008818f
C577 B.n537 VSUBS 0.008818f
C578 B.n538 VSUBS 0.008818f
C579 B.n539 VSUBS 0.008818f
C580 B.n540 VSUBS 0.008818f
C581 B.n541 VSUBS 0.008818f
C582 B.n542 VSUBS 0.008818f
C583 B.n543 VSUBS 0.008818f
C584 B.n544 VSUBS 0.008818f
C585 B.n545 VSUBS 0.008818f
C586 B.n546 VSUBS 0.008818f
C587 B.n547 VSUBS 0.008818f
C588 B.n548 VSUBS 0.008818f
C589 B.n549 VSUBS 0.008818f
C590 B.n550 VSUBS 0.008818f
C591 B.n551 VSUBS 0.008818f
C592 B.n552 VSUBS 0.008818f
C593 B.n553 VSUBS 0.008818f
C594 B.n554 VSUBS 0.008818f
C595 B.n555 VSUBS 0.008818f
C596 B.n556 VSUBS 0.008818f
C597 B.n557 VSUBS 0.008818f
C598 B.n558 VSUBS 0.008818f
C599 B.n559 VSUBS 0.008818f
C600 B.n560 VSUBS 0.008818f
C601 B.n561 VSUBS 0.008818f
C602 B.n562 VSUBS 0.008818f
C603 B.n563 VSUBS 0.008818f
C604 B.n564 VSUBS 0.008818f
C605 B.n565 VSUBS 0.008818f
C606 B.n566 VSUBS 0.008818f
C607 B.n567 VSUBS 0.008818f
C608 B.n568 VSUBS 0.008818f
C609 B.n569 VSUBS 0.008818f
C610 B.n570 VSUBS 0.008818f
C611 B.n571 VSUBS 0.008818f
C612 B.n572 VSUBS 0.008818f
C613 B.n573 VSUBS 0.008818f
C614 B.n574 VSUBS 0.008818f
C615 B.n575 VSUBS 0.008818f
C616 B.n576 VSUBS 0.008818f
C617 B.n577 VSUBS 0.008818f
C618 B.n578 VSUBS 0.008818f
C619 B.n579 VSUBS 0.008818f
C620 B.n580 VSUBS 0.008818f
C621 B.n581 VSUBS 0.008818f
C622 B.n582 VSUBS 0.008818f
C623 B.n583 VSUBS 0.008818f
C624 B.n584 VSUBS 0.008818f
C625 B.n585 VSUBS 0.008818f
C626 B.n586 VSUBS 0.008818f
C627 B.n587 VSUBS 0.008818f
C628 B.n588 VSUBS 0.008818f
C629 B.n589 VSUBS 0.008818f
C630 B.n590 VSUBS 0.008818f
C631 B.n591 VSUBS 0.008818f
C632 B.n592 VSUBS 0.008818f
C633 B.n593 VSUBS 0.008818f
C634 B.n594 VSUBS 0.008818f
C635 B.n595 VSUBS 0.008818f
C636 B.n596 VSUBS 0.008818f
C637 B.n597 VSUBS 0.008818f
C638 B.n598 VSUBS 0.008818f
C639 B.n599 VSUBS 0.008818f
C640 B.n600 VSUBS 0.008818f
C641 B.n601 VSUBS 0.008818f
C642 B.n602 VSUBS 0.008818f
C643 B.n603 VSUBS 0.008818f
C644 B.n604 VSUBS 0.008818f
C645 B.n605 VSUBS 0.008818f
C646 B.n606 VSUBS 0.008818f
C647 B.n607 VSUBS 0.008818f
C648 B.n608 VSUBS 0.008818f
C649 B.n609 VSUBS 0.008818f
C650 B.n610 VSUBS 0.008818f
C651 B.n611 VSUBS 0.008818f
C652 B.n612 VSUBS 0.008818f
C653 B.n613 VSUBS 0.008818f
C654 B.n614 VSUBS 0.008818f
C655 B.n615 VSUBS 0.008818f
C656 B.n616 VSUBS 0.008818f
C657 B.n617 VSUBS 0.008818f
C658 B.n618 VSUBS 0.008818f
C659 B.n619 VSUBS 0.008818f
C660 B.n620 VSUBS 0.01988f
C661 B.n621 VSUBS 0.01988f
C662 B.n622 VSUBS 0.02084f
C663 B.n623 VSUBS 0.008818f
C664 B.n624 VSUBS 0.008818f
C665 B.n625 VSUBS 0.008818f
C666 B.n626 VSUBS 0.008818f
C667 B.n627 VSUBS 0.008818f
C668 B.n628 VSUBS 0.008818f
C669 B.n629 VSUBS 0.008818f
C670 B.n630 VSUBS 0.008818f
C671 B.n631 VSUBS 0.008818f
C672 B.n632 VSUBS 0.008818f
C673 B.n633 VSUBS 0.008818f
C674 B.n634 VSUBS 0.008818f
C675 B.n635 VSUBS 0.008818f
C676 B.n636 VSUBS 0.008818f
C677 B.n637 VSUBS 0.008818f
C678 B.n638 VSUBS 0.008818f
C679 B.n639 VSUBS 0.008818f
C680 B.n640 VSUBS 0.008818f
C681 B.n641 VSUBS 0.008818f
C682 B.n642 VSUBS 0.008818f
C683 B.n643 VSUBS 0.008818f
C684 B.n644 VSUBS 0.008818f
C685 B.n645 VSUBS 0.008818f
C686 B.n646 VSUBS 0.008818f
C687 B.n647 VSUBS 0.008818f
C688 B.n648 VSUBS 0.008818f
C689 B.n649 VSUBS 0.008818f
C690 B.n650 VSUBS 0.008818f
C691 B.n651 VSUBS 0.008818f
C692 B.n652 VSUBS 0.008818f
C693 B.n653 VSUBS 0.008818f
C694 B.n654 VSUBS 0.008818f
C695 B.n655 VSUBS 0.008818f
C696 B.n656 VSUBS 0.008818f
C697 B.n657 VSUBS 0.008818f
C698 B.n658 VSUBS 0.008818f
C699 B.n659 VSUBS 0.008818f
C700 B.n660 VSUBS 0.008818f
C701 B.n661 VSUBS 0.008818f
C702 B.n662 VSUBS 0.008818f
C703 B.n663 VSUBS 0.008818f
C704 B.n664 VSUBS 0.008818f
C705 B.n665 VSUBS 0.008818f
C706 B.n666 VSUBS 0.008818f
C707 B.n667 VSUBS 0.008818f
C708 B.n668 VSUBS 0.008818f
C709 B.n669 VSUBS 0.008818f
C710 B.n670 VSUBS 0.008818f
C711 B.n671 VSUBS 0.008818f
C712 B.n672 VSUBS 0.008818f
C713 B.n673 VSUBS 0.008818f
C714 B.n674 VSUBS 0.008818f
C715 B.n675 VSUBS 0.008818f
C716 B.n676 VSUBS 0.008818f
C717 B.n677 VSUBS 0.008818f
C718 B.n678 VSUBS 0.008818f
C719 B.n679 VSUBS 0.008818f
C720 B.n680 VSUBS 0.008818f
C721 B.n681 VSUBS 0.008818f
C722 B.n682 VSUBS 0.008818f
C723 B.n683 VSUBS 0.008818f
C724 B.n684 VSUBS 0.008818f
C725 B.n685 VSUBS 0.008818f
C726 B.n686 VSUBS 0.008818f
C727 B.n687 VSUBS 0.008818f
C728 B.n688 VSUBS 0.008818f
C729 B.n689 VSUBS 0.008818f
C730 B.n690 VSUBS 0.008818f
C731 B.n691 VSUBS 0.008818f
C732 B.n692 VSUBS 0.008818f
C733 B.n693 VSUBS 0.008818f
C734 B.n694 VSUBS 0.008818f
C735 B.n695 VSUBS 0.008818f
C736 B.n696 VSUBS 0.008818f
C737 B.n697 VSUBS 0.008818f
C738 B.n698 VSUBS 0.008818f
C739 B.n699 VSUBS 0.006095f
C740 B.n700 VSUBS 0.020431f
C741 B.n701 VSUBS 0.007132f
C742 B.n702 VSUBS 0.008818f
C743 B.n703 VSUBS 0.008818f
C744 B.n704 VSUBS 0.008818f
C745 B.n705 VSUBS 0.008818f
C746 B.n706 VSUBS 0.008818f
C747 B.n707 VSUBS 0.008818f
C748 B.n708 VSUBS 0.008818f
C749 B.n709 VSUBS 0.008818f
C750 B.n710 VSUBS 0.008818f
C751 B.n711 VSUBS 0.008818f
C752 B.n712 VSUBS 0.008818f
C753 B.n713 VSUBS 0.007132f
C754 B.n714 VSUBS 0.020431f
C755 B.n715 VSUBS 0.006095f
C756 B.n716 VSUBS 0.008818f
C757 B.n717 VSUBS 0.008818f
C758 B.n718 VSUBS 0.008818f
C759 B.n719 VSUBS 0.008818f
C760 B.n720 VSUBS 0.008818f
C761 B.n721 VSUBS 0.008818f
C762 B.n722 VSUBS 0.008818f
C763 B.n723 VSUBS 0.008818f
C764 B.n724 VSUBS 0.008818f
C765 B.n725 VSUBS 0.008818f
C766 B.n726 VSUBS 0.008818f
C767 B.n727 VSUBS 0.008818f
C768 B.n728 VSUBS 0.008818f
C769 B.n729 VSUBS 0.008818f
C770 B.n730 VSUBS 0.008818f
C771 B.n731 VSUBS 0.008818f
C772 B.n732 VSUBS 0.008818f
C773 B.n733 VSUBS 0.008818f
C774 B.n734 VSUBS 0.008818f
C775 B.n735 VSUBS 0.008818f
C776 B.n736 VSUBS 0.008818f
C777 B.n737 VSUBS 0.008818f
C778 B.n738 VSUBS 0.008818f
C779 B.n739 VSUBS 0.008818f
C780 B.n740 VSUBS 0.008818f
C781 B.n741 VSUBS 0.008818f
C782 B.n742 VSUBS 0.008818f
C783 B.n743 VSUBS 0.008818f
C784 B.n744 VSUBS 0.008818f
C785 B.n745 VSUBS 0.008818f
C786 B.n746 VSUBS 0.008818f
C787 B.n747 VSUBS 0.008818f
C788 B.n748 VSUBS 0.008818f
C789 B.n749 VSUBS 0.008818f
C790 B.n750 VSUBS 0.008818f
C791 B.n751 VSUBS 0.008818f
C792 B.n752 VSUBS 0.008818f
C793 B.n753 VSUBS 0.008818f
C794 B.n754 VSUBS 0.008818f
C795 B.n755 VSUBS 0.008818f
C796 B.n756 VSUBS 0.008818f
C797 B.n757 VSUBS 0.008818f
C798 B.n758 VSUBS 0.008818f
C799 B.n759 VSUBS 0.008818f
C800 B.n760 VSUBS 0.008818f
C801 B.n761 VSUBS 0.008818f
C802 B.n762 VSUBS 0.008818f
C803 B.n763 VSUBS 0.008818f
C804 B.n764 VSUBS 0.008818f
C805 B.n765 VSUBS 0.008818f
C806 B.n766 VSUBS 0.008818f
C807 B.n767 VSUBS 0.008818f
C808 B.n768 VSUBS 0.008818f
C809 B.n769 VSUBS 0.008818f
C810 B.n770 VSUBS 0.008818f
C811 B.n771 VSUBS 0.008818f
C812 B.n772 VSUBS 0.008818f
C813 B.n773 VSUBS 0.008818f
C814 B.n774 VSUBS 0.008818f
C815 B.n775 VSUBS 0.008818f
C816 B.n776 VSUBS 0.008818f
C817 B.n777 VSUBS 0.008818f
C818 B.n778 VSUBS 0.008818f
C819 B.n779 VSUBS 0.008818f
C820 B.n780 VSUBS 0.008818f
C821 B.n781 VSUBS 0.008818f
C822 B.n782 VSUBS 0.008818f
C823 B.n783 VSUBS 0.008818f
C824 B.n784 VSUBS 0.008818f
C825 B.n785 VSUBS 0.008818f
C826 B.n786 VSUBS 0.008818f
C827 B.n787 VSUBS 0.008818f
C828 B.n788 VSUBS 0.008818f
C829 B.n789 VSUBS 0.008818f
C830 B.n790 VSUBS 0.008818f
C831 B.n791 VSUBS 0.008818f
C832 B.n792 VSUBS 0.02084f
C833 B.n793 VSUBS 0.01988f
C834 B.n794 VSUBS 0.01988f
C835 B.n795 VSUBS 0.008818f
C836 B.n796 VSUBS 0.008818f
C837 B.n797 VSUBS 0.008818f
C838 B.n798 VSUBS 0.008818f
C839 B.n799 VSUBS 0.008818f
C840 B.n800 VSUBS 0.008818f
C841 B.n801 VSUBS 0.008818f
C842 B.n802 VSUBS 0.008818f
C843 B.n803 VSUBS 0.008818f
C844 B.n804 VSUBS 0.008818f
C845 B.n805 VSUBS 0.008818f
C846 B.n806 VSUBS 0.008818f
C847 B.n807 VSUBS 0.008818f
C848 B.n808 VSUBS 0.008818f
C849 B.n809 VSUBS 0.008818f
C850 B.n810 VSUBS 0.008818f
C851 B.n811 VSUBS 0.008818f
C852 B.n812 VSUBS 0.008818f
C853 B.n813 VSUBS 0.008818f
C854 B.n814 VSUBS 0.008818f
C855 B.n815 VSUBS 0.008818f
C856 B.n816 VSUBS 0.008818f
C857 B.n817 VSUBS 0.008818f
C858 B.n818 VSUBS 0.008818f
C859 B.n819 VSUBS 0.008818f
C860 B.n820 VSUBS 0.008818f
C861 B.n821 VSUBS 0.008818f
C862 B.n822 VSUBS 0.008818f
C863 B.n823 VSUBS 0.008818f
C864 B.n824 VSUBS 0.008818f
C865 B.n825 VSUBS 0.008818f
C866 B.n826 VSUBS 0.008818f
C867 B.n827 VSUBS 0.008818f
C868 B.n828 VSUBS 0.008818f
C869 B.n829 VSUBS 0.008818f
C870 B.n830 VSUBS 0.008818f
C871 B.n831 VSUBS 0.008818f
C872 B.n832 VSUBS 0.008818f
C873 B.n833 VSUBS 0.008818f
C874 B.n834 VSUBS 0.008818f
C875 B.n835 VSUBS 0.008818f
C876 B.n836 VSUBS 0.008818f
C877 B.n837 VSUBS 0.008818f
C878 B.n838 VSUBS 0.008818f
C879 B.n839 VSUBS 0.008818f
C880 B.n840 VSUBS 0.008818f
C881 B.n841 VSUBS 0.008818f
C882 B.n842 VSUBS 0.008818f
C883 B.n843 VSUBS 0.008818f
C884 B.n844 VSUBS 0.008818f
C885 B.n845 VSUBS 0.008818f
C886 B.n846 VSUBS 0.008818f
C887 B.n847 VSUBS 0.008818f
C888 B.n848 VSUBS 0.008818f
C889 B.n849 VSUBS 0.008818f
C890 B.n850 VSUBS 0.008818f
C891 B.n851 VSUBS 0.008818f
C892 B.n852 VSUBS 0.008818f
C893 B.n853 VSUBS 0.008818f
C894 B.n854 VSUBS 0.008818f
C895 B.n855 VSUBS 0.008818f
C896 B.n856 VSUBS 0.008818f
C897 B.n857 VSUBS 0.008818f
C898 B.n858 VSUBS 0.008818f
C899 B.n859 VSUBS 0.008818f
C900 B.n860 VSUBS 0.008818f
C901 B.n861 VSUBS 0.008818f
C902 B.n862 VSUBS 0.008818f
C903 B.n863 VSUBS 0.008818f
C904 B.n864 VSUBS 0.008818f
C905 B.n865 VSUBS 0.008818f
C906 B.n866 VSUBS 0.008818f
C907 B.n867 VSUBS 0.011507f
C908 B.n868 VSUBS 0.012258f
C909 B.n869 VSUBS 0.024377f
C910 VDD1.n0 VSUBS 0.028449f
C911 VDD1.n1 VSUBS 0.026929f
C912 VDD1.n2 VSUBS 0.014471f
C913 VDD1.n3 VSUBS 0.034203f
C914 VDD1.n4 VSUBS 0.014896f
C915 VDD1.n5 VSUBS 0.026929f
C916 VDD1.n6 VSUBS 0.014896f
C917 VDD1.n7 VSUBS 0.014471f
C918 VDD1.n8 VSUBS 0.034203f
C919 VDD1.n9 VSUBS 0.034203f
C920 VDD1.n10 VSUBS 0.015322f
C921 VDD1.n11 VSUBS 0.026929f
C922 VDD1.n12 VSUBS 0.014471f
C923 VDD1.n13 VSUBS 0.034203f
C924 VDD1.n14 VSUBS 0.015322f
C925 VDD1.n15 VSUBS 0.026929f
C926 VDD1.n16 VSUBS 0.014471f
C927 VDD1.n17 VSUBS 0.034203f
C928 VDD1.n18 VSUBS 0.015322f
C929 VDD1.n19 VSUBS 0.026929f
C930 VDD1.n20 VSUBS 0.014471f
C931 VDD1.n21 VSUBS 0.034203f
C932 VDD1.n22 VSUBS 0.015322f
C933 VDD1.n23 VSUBS 0.026929f
C934 VDD1.n24 VSUBS 0.014471f
C935 VDD1.n25 VSUBS 0.034203f
C936 VDD1.n26 VSUBS 0.015322f
C937 VDD1.n27 VSUBS 1.77205f
C938 VDD1.n28 VSUBS 0.014471f
C939 VDD1.t1 VSUBS 0.073251f
C940 VDD1.n29 VSUBS 0.193243f
C941 VDD1.n30 VSUBS 0.021759f
C942 VDD1.n31 VSUBS 0.025652f
C943 VDD1.n32 VSUBS 0.034203f
C944 VDD1.n33 VSUBS 0.015322f
C945 VDD1.n34 VSUBS 0.014471f
C946 VDD1.n35 VSUBS 0.026929f
C947 VDD1.n36 VSUBS 0.026929f
C948 VDD1.n37 VSUBS 0.014471f
C949 VDD1.n38 VSUBS 0.015322f
C950 VDD1.n39 VSUBS 0.034203f
C951 VDD1.n40 VSUBS 0.034203f
C952 VDD1.n41 VSUBS 0.015322f
C953 VDD1.n42 VSUBS 0.014471f
C954 VDD1.n43 VSUBS 0.026929f
C955 VDD1.n44 VSUBS 0.026929f
C956 VDD1.n45 VSUBS 0.014471f
C957 VDD1.n46 VSUBS 0.015322f
C958 VDD1.n47 VSUBS 0.034203f
C959 VDD1.n48 VSUBS 0.034203f
C960 VDD1.n49 VSUBS 0.015322f
C961 VDD1.n50 VSUBS 0.014471f
C962 VDD1.n51 VSUBS 0.026929f
C963 VDD1.n52 VSUBS 0.026929f
C964 VDD1.n53 VSUBS 0.014471f
C965 VDD1.n54 VSUBS 0.015322f
C966 VDD1.n55 VSUBS 0.034203f
C967 VDD1.n56 VSUBS 0.034203f
C968 VDD1.n57 VSUBS 0.015322f
C969 VDD1.n58 VSUBS 0.014471f
C970 VDD1.n59 VSUBS 0.026929f
C971 VDD1.n60 VSUBS 0.026929f
C972 VDD1.n61 VSUBS 0.014471f
C973 VDD1.n62 VSUBS 0.015322f
C974 VDD1.n63 VSUBS 0.034203f
C975 VDD1.n64 VSUBS 0.034203f
C976 VDD1.n65 VSUBS 0.015322f
C977 VDD1.n66 VSUBS 0.014471f
C978 VDD1.n67 VSUBS 0.026929f
C979 VDD1.n68 VSUBS 0.026929f
C980 VDD1.n69 VSUBS 0.014471f
C981 VDD1.n70 VSUBS 0.015322f
C982 VDD1.n71 VSUBS 0.034203f
C983 VDD1.n72 VSUBS 0.034203f
C984 VDD1.n73 VSUBS 0.015322f
C985 VDD1.n74 VSUBS 0.014471f
C986 VDD1.n75 VSUBS 0.026929f
C987 VDD1.n76 VSUBS 0.026929f
C988 VDD1.n77 VSUBS 0.014471f
C989 VDD1.n78 VSUBS 0.015322f
C990 VDD1.n79 VSUBS 0.034203f
C991 VDD1.n80 VSUBS 0.078919f
C992 VDD1.n81 VSUBS 0.015322f
C993 VDD1.n82 VSUBS 0.014471f
C994 VDD1.n83 VSUBS 0.064821f
C995 VDD1.n84 VSUBS 0.067381f
C996 VDD1.t5 VSUBS 0.328354f
C997 VDD1.t3 VSUBS 0.328354f
C998 VDD1.n85 VSUBS 2.67982f
C999 VDD1.n86 VSUBS 0.966139f
C1000 VDD1.n87 VSUBS 0.028449f
C1001 VDD1.n88 VSUBS 0.026929f
C1002 VDD1.n89 VSUBS 0.014471f
C1003 VDD1.n90 VSUBS 0.034203f
C1004 VDD1.n91 VSUBS 0.014896f
C1005 VDD1.n92 VSUBS 0.026929f
C1006 VDD1.n93 VSUBS 0.015322f
C1007 VDD1.n94 VSUBS 0.034203f
C1008 VDD1.n95 VSUBS 0.015322f
C1009 VDD1.n96 VSUBS 0.026929f
C1010 VDD1.n97 VSUBS 0.014471f
C1011 VDD1.n98 VSUBS 0.034203f
C1012 VDD1.n99 VSUBS 0.015322f
C1013 VDD1.n100 VSUBS 0.026929f
C1014 VDD1.n101 VSUBS 0.014471f
C1015 VDD1.n102 VSUBS 0.034203f
C1016 VDD1.n103 VSUBS 0.015322f
C1017 VDD1.n104 VSUBS 0.026929f
C1018 VDD1.n105 VSUBS 0.014471f
C1019 VDD1.n106 VSUBS 0.034203f
C1020 VDD1.n107 VSUBS 0.015322f
C1021 VDD1.n108 VSUBS 0.026929f
C1022 VDD1.n109 VSUBS 0.014471f
C1023 VDD1.n110 VSUBS 0.034203f
C1024 VDD1.n111 VSUBS 0.015322f
C1025 VDD1.n112 VSUBS 1.77205f
C1026 VDD1.n113 VSUBS 0.014471f
C1027 VDD1.t0 VSUBS 0.073251f
C1028 VDD1.n114 VSUBS 0.193243f
C1029 VDD1.n115 VSUBS 0.021759f
C1030 VDD1.n116 VSUBS 0.025652f
C1031 VDD1.n117 VSUBS 0.034203f
C1032 VDD1.n118 VSUBS 0.015322f
C1033 VDD1.n119 VSUBS 0.014471f
C1034 VDD1.n120 VSUBS 0.026929f
C1035 VDD1.n121 VSUBS 0.026929f
C1036 VDD1.n122 VSUBS 0.014471f
C1037 VDD1.n123 VSUBS 0.015322f
C1038 VDD1.n124 VSUBS 0.034203f
C1039 VDD1.n125 VSUBS 0.034203f
C1040 VDD1.n126 VSUBS 0.015322f
C1041 VDD1.n127 VSUBS 0.014471f
C1042 VDD1.n128 VSUBS 0.026929f
C1043 VDD1.n129 VSUBS 0.026929f
C1044 VDD1.n130 VSUBS 0.014471f
C1045 VDD1.n131 VSUBS 0.015322f
C1046 VDD1.n132 VSUBS 0.034203f
C1047 VDD1.n133 VSUBS 0.034203f
C1048 VDD1.n134 VSUBS 0.015322f
C1049 VDD1.n135 VSUBS 0.014471f
C1050 VDD1.n136 VSUBS 0.026929f
C1051 VDD1.n137 VSUBS 0.026929f
C1052 VDD1.n138 VSUBS 0.014471f
C1053 VDD1.n139 VSUBS 0.015322f
C1054 VDD1.n140 VSUBS 0.034203f
C1055 VDD1.n141 VSUBS 0.034203f
C1056 VDD1.n142 VSUBS 0.015322f
C1057 VDD1.n143 VSUBS 0.014471f
C1058 VDD1.n144 VSUBS 0.026929f
C1059 VDD1.n145 VSUBS 0.026929f
C1060 VDD1.n146 VSUBS 0.014471f
C1061 VDD1.n147 VSUBS 0.015322f
C1062 VDD1.n148 VSUBS 0.034203f
C1063 VDD1.n149 VSUBS 0.034203f
C1064 VDD1.n150 VSUBS 0.015322f
C1065 VDD1.n151 VSUBS 0.014471f
C1066 VDD1.n152 VSUBS 0.026929f
C1067 VDD1.n153 VSUBS 0.026929f
C1068 VDD1.n154 VSUBS 0.014471f
C1069 VDD1.n155 VSUBS 0.014471f
C1070 VDD1.n156 VSUBS 0.015322f
C1071 VDD1.n157 VSUBS 0.034203f
C1072 VDD1.n158 VSUBS 0.034203f
C1073 VDD1.n159 VSUBS 0.034203f
C1074 VDD1.n160 VSUBS 0.014896f
C1075 VDD1.n161 VSUBS 0.014471f
C1076 VDD1.n162 VSUBS 0.026929f
C1077 VDD1.n163 VSUBS 0.026929f
C1078 VDD1.n164 VSUBS 0.014471f
C1079 VDD1.n165 VSUBS 0.015322f
C1080 VDD1.n166 VSUBS 0.034203f
C1081 VDD1.n167 VSUBS 0.078919f
C1082 VDD1.n168 VSUBS 0.015322f
C1083 VDD1.n169 VSUBS 0.014471f
C1084 VDD1.n170 VSUBS 0.064821f
C1085 VDD1.n171 VSUBS 0.067381f
C1086 VDD1.t8 VSUBS 0.328354f
C1087 VDD1.t6 VSUBS 0.328354f
C1088 VDD1.n172 VSUBS 2.67981f
C1089 VDD1.n173 VSUBS 0.957651f
C1090 VDD1.t2 VSUBS 0.328354f
C1091 VDD1.t4 VSUBS 0.328354f
C1092 VDD1.n174 VSUBS 2.69688f
C1093 VDD1.n175 VSUBS 3.46881f
C1094 VDD1.t7 VSUBS 0.328354f
C1095 VDD1.t9 VSUBS 0.328354f
C1096 VDD1.n176 VSUBS 2.67981f
C1097 VDD1.n177 VSUBS 3.75449f
C1098 VP.n0 VSUBS 0.042248f
C1099 VP.t5 VSUBS 2.80641f
C1100 VP.n1 VSUBS 0.030272f
C1101 VP.n2 VSUBS 0.032045f
C1102 VP.t7 VSUBS 2.80641f
C1103 VP.n3 VSUBS 0.051245f
C1104 VP.n4 VSUBS 0.032045f
C1105 VP.t3 VSUBS 2.80641f
C1106 VP.n5 VSUBS 0.059724f
C1107 VP.n6 VSUBS 0.032045f
C1108 VP.t1 VSUBS 2.80641f
C1109 VP.n7 VSUBS 0.98561f
C1110 VP.n8 VSUBS 0.032045f
C1111 VP.n9 VSUBS 0.058814f
C1112 VP.n10 VSUBS 0.042248f
C1113 VP.t0 VSUBS 2.80641f
C1114 VP.n11 VSUBS 0.030272f
C1115 VP.n12 VSUBS 0.032045f
C1116 VP.t2 VSUBS 2.80641f
C1117 VP.n13 VSUBS 0.051245f
C1118 VP.n14 VSUBS 0.032045f
C1119 VP.t6 VSUBS 2.80641f
C1120 VP.n15 VSUBS 0.059724f
C1121 VP.n16 VSUBS 0.032045f
C1122 VP.t4 VSUBS 2.80641f
C1123 VP.n17 VSUBS 1.07392f
C1124 VP.t8 VSUBS 2.98475f
C1125 VP.n18 VSUBS 1.05905f
C1126 VP.n19 VSUBS 0.268746f
C1127 VP.n20 VSUBS 0.053826f
C1128 VP.n21 VSUBS 0.051245f
C1129 VP.n22 VSUBS 0.042315f
C1130 VP.n23 VSUBS 0.032045f
C1131 VP.n24 VSUBS 0.032045f
C1132 VP.n25 VSUBS 0.032045f
C1133 VP.n26 VSUBS 1.01585f
C1134 VP.n27 VSUBS 0.059724f
C1135 VP.n28 VSUBS 0.042315f
C1136 VP.n29 VSUBS 0.032045f
C1137 VP.n30 VSUBS 0.032045f
C1138 VP.n31 VSUBS 0.032045f
C1139 VP.n32 VSUBS 0.053826f
C1140 VP.n33 VSUBS 0.98561f
C1141 VP.n34 VSUBS 0.036135f
C1142 VP.n35 VSUBS 0.064197f
C1143 VP.n36 VSUBS 0.032045f
C1144 VP.n37 VSUBS 0.032045f
C1145 VP.n38 VSUBS 0.032045f
C1146 VP.n39 VSUBS 0.058814f
C1147 VP.n40 VSUBS 0.047929f
C1148 VP.n41 VSUBS 1.07775f
C1149 VP.n42 VSUBS 1.91943f
C1150 VP.n43 VSUBS 1.94125f
C1151 VP.t9 VSUBS 2.80641f
C1152 VP.n44 VSUBS 1.07775f
C1153 VP.n45 VSUBS 0.047929f
C1154 VP.n46 VSUBS 0.042248f
C1155 VP.n47 VSUBS 0.032045f
C1156 VP.n48 VSUBS 0.032045f
C1157 VP.n49 VSUBS 0.030272f
C1158 VP.n50 VSUBS 0.064197f
C1159 VP.n51 VSUBS 0.036135f
C1160 VP.n52 VSUBS 0.032045f
C1161 VP.n53 VSUBS 0.032045f
C1162 VP.n54 VSUBS 0.053826f
C1163 VP.n55 VSUBS 0.051245f
C1164 VP.n56 VSUBS 0.042315f
C1165 VP.n57 VSUBS 0.032045f
C1166 VP.n58 VSUBS 0.032045f
C1167 VP.n59 VSUBS 0.032045f
C1168 VP.n60 VSUBS 1.01585f
C1169 VP.n61 VSUBS 0.059724f
C1170 VP.n62 VSUBS 0.042315f
C1171 VP.n63 VSUBS 0.032045f
C1172 VP.n64 VSUBS 0.032045f
C1173 VP.n65 VSUBS 0.032045f
C1174 VP.n66 VSUBS 0.053826f
C1175 VP.n67 VSUBS 0.98561f
C1176 VP.n68 VSUBS 0.036135f
C1177 VP.n69 VSUBS 0.064197f
C1178 VP.n70 VSUBS 0.032045f
C1179 VP.n71 VSUBS 0.032045f
C1180 VP.n72 VSUBS 0.032045f
C1181 VP.n73 VSUBS 0.058814f
C1182 VP.n74 VSUBS 0.047929f
C1183 VP.n75 VSUBS 1.07775f
C1184 VP.n76 VSUBS 0.043666f
C1185 VTAIL.t10 VSUBS 0.336023f
C1186 VTAIL.t19 VSUBS 0.336023f
C1187 VTAIL.n0 VSUBS 2.58459f
C1188 VTAIL.n1 VSUBS 0.92192f
C1189 VTAIL.n2 VSUBS 0.029114f
C1190 VTAIL.n3 VSUBS 0.027558f
C1191 VTAIL.n4 VSUBS 0.014809f
C1192 VTAIL.n5 VSUBS 0.035002f
C1193 VTAIL.n6 VSUBS 0.015244f
C1194 VTAIL.n7 VSUBS 0.027558f
C1195 VTAIL.n8 VSUBS 0.01568f
C1196 VTAIL.n9 VSUBS 0.035002f
C1197 VTAIL.n10 VSUBS 0.01568f
C1198 VTAIL.n11 VSUBS 0.027558f
C1199 VTAIL.n12 VSUBS 0.014809f
C1200 VTAIL.n13 VSUBS 0.035002f
C1201 VTAIL.n14 VSUBS 0.01568f
C1202 VTAIL.n15 VSUBS 0.027558f
C1203 VTAIL.n16 VSUBS 0.014809f
C1204 VTAIL.n17 VSUBS 0.035002f
C1205 VTAIL.n18 VSUBS 0.01568f
C1206 VTAIL.n19 VSUBS 0.027558f
C1207 VTAIL.n20 VSUBS 0.014809f
C1208 VTAIL.n21 VSUBS 0.035002f
C1209 VTAIL.n22 VSUBS 0.01568f
C1210 VTAIL.n23 VSUBS 0.027558f
C1211 VTAIL.n24 VSUBS 0.014809f
C1212 VTAIL.n25 VSUBS 0.035002f
C1213 VTAIL.n26 VSUBS 0.01568f
C1214 VTAIL.n27 VSUBS 1.81344f
C1215 VTAIL.n28 VSUBS 0.014809f
C1216 VTAIL.t8 VSUBS 0.074962f
C1217 VTAIL.n29 VSUBS 0.197756f
C1218 VTAIL.n30 VSUBS 0.022267f
C1219 VTAIL.n31 VSUBS 0.026252f
C1220 VTAIL.n32 VSUBS 0.035002f
C1221 VTAIL.n33 VSUBS 0.01568f
C1222 VTAIL.n34 VSUBS 0.014809f
C1223 VTAIL.n35 VSUBS 0.027558f
C1224 VTAIL.n36 VSUBS 0.027558f
C1225 VTAIL.n37 VSUBS 0.014809f
C1226 VTAIL.n38 VSUBS 0.01568f
C1227 VTAIL.n39 VSUBS 0.035002f
C1228 VTAIL.n40 VSUBS 0.035002f
C1229 VTAIL.n41 VSUBS 0.01568f
C1230 VTAIL.n42 VSUBS 0.014809f
C1231 VTAIL.n43 VSUBS 0.027558f
C1232 VTAIL.n44 VSUBS 0.027558f
C1233 VTAIL.n45 VSUBS 0.014809f
C1234 VTAIL.n46 VSUBS 0.01568f
C1235 VTAIL.n47 VSUBS 0.035002f
C1236 VTAIL.n48 VSUBS 0.035002f
C1237 VTAIL.n49 VSUBS 0.01568f
C1238 VTAIL.n50 VSUBS 0.014809f
C1239 VTAIL.n51 VSUBS 0.027558f
C1240 VTAIL.n52 VSUBS 0.027558f
C1241 VTAIL.n53 VSUBS 0.014809f
C1242 VTAIL.n54 VSUBS 0.01568f
C1243 VTAIL.n55 VSUBS 0.035002f
C1244 VTAIL.n56 VSUBS 0.035002f
C1245 VTAIL.n57 VSUBS 0.01568f
C1246 VTAIL.n58 VSUBS 0.014809f
C1247 VTAIL.n59 VSUBS 0.027558f
C1248 VTAIL.n60 VSUBS 0.027558f
C1249 VTAIL.n61 VSUBS 0.014809f
C1250 VTAIL.n62 VSUBS 0.01568f
C1251 VTAIL.n63 VSUBS 0.035002f
C1252 VTAIL.n64 VSUBS 0.035002f
C1253 VTAIL.n65 VSUBS 0.01568f
C1254 VTAIL.n66 VSUBS 0.014809f
C1255 VTAIL.n67 VSUBS 0.027558f
C1256 VTAIL.n68 VSUBS 0.027558f
C1257 VTAIL.n69 VSUBS 0.014809f
C1258 VTAIL.n70 VSUBS 0.014809f
C1259 VTAIL.n71 VSUBS 0.01568f
C1260 VTAIL.n72 VSUBS 0.035002f
C1261 VTAIL.n73 VSUBS 0.035002f
C1262 VTAIL.n74 VSUBS 0.035002f
C1263 VTAIL.n75 VSUBS 0.015244f
C1264 VTAIL.n76 VSUBS 0.014809f
C1265 VTAIL.n77 VSUBS 0.027558f
C1266 VTAIL.n78 VSUBS 0.027558f
C1267 VTAIL.n79 VSUBS 0.014809f
C1268 VTAIL.n80 VSUBS 0.01568f
C1269 VTAIL.n81 VSUBS 0.035002f
C1270 VTAIL.n82 VSUBS 0.080762f
C1271 VTAIL.n83 VSUBS 0.01568f
C1272 VTAIL.n84 VSUBS 0.014809f
C1273 VTAIL.n85 VSUBS 0.066335f
C1274 VTAIL.n86 VSUBS 0.040518f
C1275 VTAIL.n87 VSUBS 0.342326f
C1276 VTAIL.t9 VSUBS 0.336023f
C1277 VTAIL.t1 VSUBS 0.336023f
C1278 VTAIL.n88 VSUBS 2.58459f
C1279 VTAIL.n89 VSUBS 1.01282f
C1280 VTAIL.t0 VSUBS 0.336023f
C1281 VTAIL.t7 VSUBS 0.336023f
C1282 VTAIL.n90 VSUBS 2.58459f
C1283 VTAIL.n91 VSUBS 2.75206f
C1284 VTAIL.t17 VSUBS 0.336023f
C1285 VTAIL.t16 VSUBS 0.336023f
C1286 VTAIL.n92 VSUBS 2.58461f
C1287 VTAIL.n93 VSUBS 2.75204f
C1288 VTAIL.t13 VSUBS 0.336023f
C1289 VTAIL.t14 VSUBS 0.336023f
C1290 VTAIL.n94 VSUBS 2.58461f
C1291 VTAIL.n95 VSUBS 1.01281f
C1292 VTAIL.n96 VSUBS 0.029114f
C1293 VTAIL.n97 VSUBS 0.027558f
C1294 VTAIL.n98 VSUBS 0.014809f
C1295 VTAIL.n99 VSUBS 0.035002f
C1296 VTAIL.n100 VSUBS 0.015244f
C1297 VTAIL.n101 VSUBS 0.027558f
C1298 VTAIL.n102 VSUBS 0.015244f
C1299 VTAIL.n103 VSUBS 0.014809f
C1300 VTAIL.n104 VSUBS 0.035002f
C1301 VTAIL.n105 VSUBS 0.035002f
C1302 VTAIL.n106 VSUBS 0.01568f
C1303 VTAIL.n107 VSUBS 0.027558f
C1304 VTAIL.n108 VSUBS 0.014809f
C1305 VTAIL.n109 VSUBS 0.035002f
C1306 VTAIL.n110 VSUBS 0.01568f
C1307 VTAIL.n111 VSUBS 0.027558f
C1308 VTAIL.n112 VSUBS 0.014809f
C1309 VTAIL.n113 VSUBS 0.035002f
C1310 VTAIL.n114 VSUBS 0.01568f
C1311 VTAIL.n115 VSUBS 0.027558f
C1312 VTAIL.n116 VSUBS 0.014809f
C1313 VTAIL.n117 VSUBS 0.035002f
C1314 VTAIL.n118 VSUBS 0.01568f
C1315 VTAIL.n119 VSUBS 0.027558f
C1316 VTAIL.n120 VSUBS 0.014809f
C1317 VTAIL.n121 VSUBS 0.035002f
C1318 VTAIL.n122 VSUBS 0.01568f
C1319 VTAIL.n123 VSUBS 1.81344f
C1320 VTAIL.n124 VSUBS 0.014809f
C1321 VTAIL.t15 VSUBS 0.074962f
C1322 VTAIL.n125 VSUBS 0.197756f
C1323 VTAIL.n126 VSUBS 0.022267f
C1324 VTAIL.n127 VSUBS 0.026252f
C1325 VTAIL.n128 VSUBS 0.035002f
C1326 VTAIL.n129 VSUBS 0.01568f
C1327 VTAIL.n130 VSUBS 0.014809f
C1328 VTAIL.n131 VSUBS 0.027558f
C1329 VTAIL.n132 VSUBS 0.027558f
C1330 VTAIL.n133 VSUBS 0.014809f
C1331 VTAIL.n134 VSUBS 0.01568f
C1332 VTAIL.n135 VSUBS 0.035002f
C1333 VTAIL.n136 VSUBS 0.035002f
C1334 VTAIL.n137 VSUBS 0.01568f
C1335 VTAIL.n138 VSUBS 0.014809f
C1336 VTAIL.n139 VSUBS 0.027558f
C1337 VTAIL.n140 VSUBS 0.027558f
C1338 VTAIL.n141 VSUBS 0.014809f
C1339 VTAIL.n142 VSUBS 0.01568f
C1340 VTAIL.n143 VSUBS 0.035002f
C1341 VTAIL.n144 VSUBS 0.035002f
C1342 VTAIL.n145 VSUBS 0.01568f
C1343 VTAIL.n146 VSUBS 0.014809f
C1344 VTAIL.n147 VSUBS 0.027558f
C1345 VTAIL.n148 VSUBS 0.027558f
C1346 VTAIL.n149 VSUBS 0.014809f
C1347 VTAIL.n150 VSUBS 0.01568f
C1348 VTAIL.n151 VSUBS 0.035002f
C1349 VTAIL.n152 VSUBS 0.035002f
C1350 VTAIL.n153 VSUBS 0.01568f
C1351 VTAIL.n154 VSUBS 0.014809f
C1352 VTAIL.n155 VSUBS 0.027558f
C1353 VTAIL.n156 VSUBS 0.027558f
C1354 VTAIL.n157 VSUBS 0.014809f
C1355 VTAIL.n158 VSUBS 0.01568f
C1356 VTAIL.n159 VSUBS 0.035002f
C1357 VTAIL.n160 VSUBS 0.035002f
C1358 VTAIL.n161 VSUBS 0.01568f
C1359 VTAIL.n162 VSUBS 0.014809f
C1360 VTAIL.n163 VSUBS 0.027558f
C1361 VTAIL.n164 VSUBS 0.027558f
C1362 VTAIL.n165 VSUBS 0.014809f
C1363 VTAIL.n166 VSUBS 0.01568f
C1364 VTAIL.n167 VSUBS 0.035002f
C1365 VTAIL.n168 VSUBS 0.035002f
C1366 VTAIL.n169 VSUBS 0.01568f
C1367 VTAIL.n170 VSUBS 0.014809f
C1368 VTAIL.n171 VSUBS 0.027558f
C1369 VTAIL.n172 VSUBS 0.027558f
C1370 VTAIL.n173 VSUBS 0.014809f
C1371 VTAIL.n174 VSUBS 0.01568f
C1372 VTAIL.n175 VSUBS 0.035002f
C1373 VTAIL.n176 VSUBS 0.080762f
C1374 VTAIL.n177 VSUBS 0.01568f
C1375 VTAIL.n178 VSUBS 0.014809f
C1376 VTAIL.n179 VSUBS 0.066335f
C1377 VTAIL.n180 VSUBS 0.040518f
C1378 VTAIL.n181 VSUBS 0.342326f
C1379 VTAIL.t4 VSUBS 0.336023f
C1380 VTAIL.t5 VSUBS 0.336023f
C1381 VTAIL.n182 VSUBS 2.58461f
C1382 VTAIL.n183 VSUBS 0.962667f
C1383 VTAIL.t2 VSUBS 0.336023f
C1384 VTAIL.t3 VSUBS 0.336023f
C1385 VTAIL.n184 VSUBS 2.58461f
C1386 VTAIL.n185 VSUBS 1.01281f
C1387 VTAIL.n186 VSUBS 0.029114f
C1388 VTAIL.n187 VSUBS 0.027558f
C1389 VTAIL.n188 VSUBS 0.014809f
C1390 VTAIL.n189 VSUBS 0.035002f
C1391 VTAIL.n190 VSUBS 0.015244f
C1392 VTAIL.n191 VSUBS 0.027558f
C1393 VTAIL.n192 VSUBS 0.015244f
C1394 VTAIL.n193 VSUBS 0.014809f
C1395 VTAIL.n194 VSUBS 0.035002f
C1396 VTAIL.n195 VSUBS 0.035002f
C1397 VTAIL.n196 VSUBS 0.01568f
C1398 VTAIL.n197 VSUBS 0.027558f
C1399 VTAIL.n198 VSUBS 0.014809f
C1400 VTAIL.n199 VSUBS 0.035002f
C1401 VTAIL.n200 VSUBS 0.01568f
C1402 VTAIL.n201 VSUBS 0.027558f
C1403 VTAIL.n202 VSUBS 0.014809f
C1404 VTAIL.n203 VSUBS 0.035002f
C1405 VTAIL.n204 VSUBS 0.01568f
C1406 VTAIL.n205 VSUBS 0.027558f
C1407 VTAIL.n206 VSUBS 0.014809f
C1408 VTAIL.n207 VSUBS 0.035002f
C1409 VTAIL.n208 VSUBS 0.01568f
C1410 VTAIL.n209 VSUBS 0.027558f
C1411 VTAIL.n210 VSUBS 0.014809f
C1412 VTAIL.n211 VSUBS 0.035002f
C1413 VTAIL.n212 VSUBS 0.01568f
C1414 VTAIL.n213 VSUBS 1.81344f
C1415 VTAIL.n214 VSUBS 0.014809f
C1416 VTAIL.t6 VSUBS 0.074962f
C1417 VTAIL.n215 VSUBS 0.197756f
C1418 VTAIL.n216 VSUBS 0.022267f
C1419 VTAIL.n217 VSUBS 0.026252f
C1420 VTAIL.n218 VSUBS 0.035002f
C1421 VTAIL.n219 VSUBS 0.01568f
C1422 VTAIL.n220 VSUBS 0.014809f
C1423 VTAIL.n221 VSUBS 0.027558f
C1424 VTAIL.n222 VSUBS 0.027558f
C1425 VTAIL.n223 VSUBS 0.014809f
C1426 VTAIL.n224 VSUBS 0.01568f
C1427 VTAIL.n225 VSUBS 0.035002f
C1428 VTAIL.n226 VSUBS 0.035002f
C1429 VTAIL.n227 VSUBS 0.01568f
C1430 VTAIL.n228 VSUBS 0.014809f
C1431 VTAIL.n229 VSUBS 0.027558f
C1432 VTAIL.n230 VSUBS 0.027558f
C1433 VTAIL.n231 VSUBS 0.014809f
C1434 VTAIL.n232 VSUBS 0.01568f
C1435 VTAIL.n233 VSUBS 0.035002f
C1436 VTAIL.n234 VSUBS 0.035002f
C1437 VTAIL.n235 VSUBS 0.01568f
C1438 VTAIL.n236 VSUBS 0.014809f
C1439 VTAIL.n237 VSUBS 0.027558f
C1440 VTAIL.n238 VSUBS 0.027558f
C1441 VTAIL.n239 VSUBS 0.014809f
C1442 VTAIL.n240 VSUBS 0.01568f
C1443 VTAIL.n241 VSUBS 0.035002f
C1444 VTAIL.n242 VSUBS 0.035002f
C1445 VTAIL.n243 VSUBS 0.01568f
C1446 VTAIL.n244 VSUBS 0.014809f
C1447 VTAIL.n245 VSUBS 0.027558f
C1448 VTAIL.n246 VSUBS 0.027558f
C1449 VTAIL.n247 VSUBS 0.014809f
C1450 VTAIL.n248 VSUBS 0.01568f
C1451 VTAIL.n249 VSUBS 0.035002f
C1452 VTAIL.n250 VSUBS 0.035002f
C1453 VTAIL.n251 VSUBS 0.01568f
C1454 VTAIL.n252 VSUBS 0.014809f
C1455 VTAIL.n253 VSUBS 0.027558f
C1456 VTAIL.n254 VSUBS 0.027558f
C1457 VTAIL.n255 VSUBS 0.014809f
C1458 VTAIL.n256 VSUBS 0.01568f
C1459 VTAIL.n257 VSUBS 0.035002f
C1460 VTAIL.n258 VSUBS 0.035002f
C1461 VTAIL.n259 VSUBS 0.01568f
C1462 VTAIL.n260 VSUBS 0.014809f
C1463 VTAIL.n261 VSUBS 0.027558f
C1464 VTAIL.n262 VSUBS 0.027558f
C1465 VTAIL.n263 VSUBS 0.014809f
C1466 VTAIL.n264 VSUBS 0.01568f
C1467 VTAIL.n265 VSUBS 0.035002f
C1468 VTAIL.n266 VSUBS 0.080762f
C1469 VTAIL.n267 VSUBS 0.01568f
C1470 VTAIL.n268 VSUBS 0.014809f
C1471 VTAIL.n269 VSUBS 0.066335f
C1472 VTAIL.n270 VSUBS 0.040518f
C1473 VTAIL.n271 VSUBS 1.94798f
C1474 VTAIL.n272 VSUBS 0.029114f
C1475 VTAIL.n273 VSUBS 0.027558f
C1476 VTAIL.n274 VSUBS 0.014809f
C1477 VTAIL.n275 VSUBS 0.035002f
C1478 VTAIL.n276 VSUBS 0.015244f
C1479 VTAIL.n277 VSUBS 0.027558f
C1480 VTAIL.n278 VSUBS 0.01568f
C1481 VTAIL.n279 VSUBS 0.035002f
C1482 VTAIL.n280 VSUBS 0.01568f
C1483 VTAIL.n281 VSUBS 0.027558f
C1484 VTAIL.n282 VSUBS 0.014809f
C1485 VTAIL.n283 VSUBS 0.035002f
C1486 VTAIL.n284 VSUBS 0.01568f
C1487 VTAIL.n285 VSUBS 0.027558f
C1488 VTAIL.n286 VSUBS 0.014809f
C1489 VTAIL.n287 VSUBS 0.035002f
C1490 VTAIL.n288 VSUBS 0.01568f
C1491 VTAIL.n289 VSUBS 0.027558f
C1492 VTAIL.n290 VSUBS 0.014809f
C1493 VTAIL.n291 VSUBS 0.035002f
C1494 VTAIL.n292 VSUBS 0.01568f
C1495 VTAIL.n293 VSUBS 0.027558f
C1496 VTAIL.n294 VSUBS 0.014809f
C1497 VTAIL.n295 VSUBS 0.035002f
C1498 VTAIL.n296 VSUBS 0.01568f
C1499 VTAIL.n297 VSUBS 1.81344f
C1500 VTAIL.n298 VSUBS 0.014809f
C1501 VTAIL.t12 VSUBS 0.074962f
C1502 VTAIL.n299 VSUBS 0.197756f
C1503 VTAIL.n300 VSUBS 0.022267f
C1504 VTAIL.n301 VSUBS 0.026252f
C1505 VTAIL.n302 VSUBS 0.035002f
C1506 VTAIL.n303 VSUBS 0.01568f
C1507 VTAIL.n304 VSUBS 0.014809f
C1508 VTAIL.n305 VSUBS 0.027558f
C1509 VTAIL.n306 VSUBS 0.027558f
C1510 VTAIL.n307 VSUBS 0.014809f
C1511 VTAIL.n308 VSUBS 0.01568f
C1512 VTAIL.n309 VSUBS 0.035002f
C1513 VTAIL.n310 VSUBS 0.035002f
C1514 VTAIL.n311 VSUBS 0.01568f
C1515 VTAIL.n312 VSUBS 0.014809f
C1516 VTAIL.n313 VSUBS 0.027558f
C1517 VTAIL.n314 VSUBS 0.027558f
C1518 VTAIL.n315 VSUBS 0.014809f
C1519 VTAIL.n316 VSUBS 0.01568f
C1520 VTAIL.n317 VSUBS 0.035002f
C1521 VTAIL.n318 VSUBS 0.035002f
C1522 VTAIL.n319 VSUBS 0.01568f
C1523 VTAIL.n320 VSUBS 0.014809f
C1524 VTAIL.n321 VSUBS 0.027558f
C1525 VTAIL.n322 VSUBS 0.027558f
C1526 VTAIL.n323 VSUBS 0.014809f
C1527 VTAIL.n324 VSUBS 0.01568f
C1528 VTAIL.n325 VSUBS 0.035002f
C1529 VTAIL.n326 VSUBS 0.035002f
C1530 VTAIL.n327 VSUBS 0.01568f
C1531 VTAIL.n328 VSUBS 0.014809f
C1532 VTAIL.n329 VSUBS 0.027558f
C1533 VTAIL.n330 VSUBS 0.027558f
C1534 VTAIL.n331 VSUBS 0.014809f
C1535 VTAIL.n332 VSUBS 0.01568f
C1536 VTAIL.n333 VSUBS 0.035002f
C1537 VTAIL.n334 VSUBS 0.035002f
C1538 VTAIL.n335 VSUBS 0.01568f
C1539 VTAIL.n336 VSUBS 0.014809f
C1540 VTAIL.n337 VSUBS 0.027558f
C1541 VTAIL.n338 VSUBS 0.027558f
C1542 VTAIL.n339 VSUBS 0.014809f
C1543 VTAIL.n340 VSUBS 0.014809f
C1544 VTAIL.n341 VSUBS 0.01568f
C1545 VTAIL.n342 VSUBS 0.035002f
C1546 VTAIL.n343 VSUBS 0.035002f
C1547 VTAIL.n344 VSUBS 0.035002f
C1548 VTAIL.n345 VSUBS 0.015244f
C1549 VTAIL.n346 VSUBS 0.014809f
C1550 VTAIL.n347 VSUBS 0.027558f
C1551 VTAIL.n348 VSUBS 0.027558f
C1552 VTAIL.n349 VSUBS 0.014809f
C1553 VTAIL.n350 VSUBS 0.01568f
C1554 VTAIL.n351 VSUBS 0.035002f
C1555 VTAIL.n352 VSUBS 0.080762f
C1556 VTAIL.n353 VSUBS 0.01568f
C1557 VTAIL.n354 VSUBS 0.014809f
C1558 VTAIL.n355 VSUBS 0.066335f
C1559 VTAIL.n356 VSUBS 0.040518f
C1560 VTAIL.n357 VSUBS 1.94798f
C1561 VTAIL.t18 VSUBS 0.336023f
C1562 VTAIL.t11 VSUBS 0.336023f
C1563 VTAIL.n358 VSUBS 2.58459f
C1564 VTAIL.n359 VSUBS 0.869866f
C1565 VDD2.n0 VSUBS 0.028356f
C1566 VDD2.n1 VSUBS 0.026841f
C1567 VDD2.n2 VSUBS 0.014423f
C1568 VDD2.n3 VSUBS 0.034091f
C1569 VDD2.n4 VSUBS 0.014847f
C1570 VDD2.n5 VSUBS 0.026841f
C1571 VDD2.n6 VSUBS 0.015272f
C1572 VDD2.n7 VSUBS 0.034091f
C1573 VDD2.n8 VSUBS 0.015272f
C1574 VDD2.n9 VSUBS 0.026841f
C1575 VDD2.n10 VSUBS 0.014423f
C1576 VDD2.n11 VSUBS 0.034091f
C1577 VDD2.n12 VSUBS 0.015272f
C1578 VDD2.n13 VSUBS 0.026841f
C1579 VDD2.n14 VSUBS 0.014423f
C1580 VDD2.n15 VSUBS 0.034091f
C1581 VDD2.n16 VSUBS 0.015272f
C1582 VDD2.n17 VSUBS 0.026841f
C1583 VDD2.n18 VSUBS 0.014423f
C1584 VDD2.n19 VSUBS 0.034091f
C1585 VDD2.n20 VSUBS 0.015272f
C1586 VDD2.n21 VSUBS 0.026841f
C1587 VDD2.n22 VSUBS 0.014423f
C1588 VDD2.n23 VSUBS 0.034091f
C1589 VDD2.n24 VSUBS 0.015272f
C1590 VDD2.n25 VSUBS 1.76625f
C1591 VDD2.n26 VSUBS 0.014423f
C1592 VDD2.t6 VSUBS 0.073011f
C1593 VDD2.n27 VSUBS 0.19261f
C1594 VDD2.n28 VSUBS 0.021687f
C1595 VDD2.n29 VSUBS 0.025568f
C1596 VDD2.n30 VSUBS 0.034091f
C1597 VDD2.n31 VSUBS 0.015272f
C1598 VDD2.n32 VSUBS 0.014423f
C1599 VDD2.n33 VSUBS 0.026841f
C1600 VDD2.n34 VSUBS 0.026841f
C1601 VDD2.n35 VSUBS 0.014423f
C1602 VDD2.n36 VSUBS 0.015272f
C1603 VDD2.n37 VSUBS 0.034091f
C1604 VDD2.n38 VSUBS 0.034091f
C1605 VDD2.n39 VSUBS 0.015272f
C1606 VDD2.n40 VSUBS 0.014423f
C1607 VDD2.n41 VSUBS 0.026841f
C1608 VDD2.n42 VSUBS 0.026841f
C1609 VDD2.n43 VSUBS 0.014423f
C1610 VDD2.n44 VSUBS 0.015272f
C1611 VDD2.n45 VSUBS 0.034091f
C1612 VDD2.n46 VSUBS 0.034091f
C1613 VDD2.n47 VSUBS 0.015272f
C1614 VDD2.n48 VSUBS 0.014423f
C1615 VDD2.n49 VSUBS 0.026841f
C1616 VDD2.n50 VSUBS 0.026841f
C1617 VDD2.n51 VSUBS 0.014423f
C1618 VDD2.n52 VSUBS 0.015272f
C1619 VDD2.n53 VSUBS 0.034091f
C1620 VDD2.n54 VSUBS 0.034091f
C1621 VDD2.n55 VSUBS 0.015272f
C1622 VDD2.n56 VSUBS 0.014423f
C1623 VDD2.n57 VSUBS 0.026841f
C1624 VDD2.n58 VSUBS 0.026841f
C1625 VDD2.n59 VSUBS 0.014423f
C1626 VDD2.n60 VSUBS 0.015272f
C1627 VDD2.n61 VSUBS 0.034091f
C1628 VDD2.n62 VSUBS 0.034091f
C1629 VDD2.n63 VSUBS 0.015272f
C1630 VDD2.n64 VSUBS 0.014423f
C1631 VDD2.n65 VSUBS 0.026841f
C1632 VDD2.n66 VSUBS 0.026841f
C1633 VDD2.n67 VSUBS 0.014423f
C1634 VDD2.n68 VSUBS 0.014423f
C1635 VDD2.n69 VSUBS 0.015272f
C1636 VDD2.n70 VSUBS 0.034091f
C1637 VDD2.n71 VSUBS 0.034091f
C1638 VDD2.n72 VSUBS 0.034091f
C1639 VDD2.n73 VSUBS 0.014847f
C1640 VDD2.n74 VSUBS 0.014423f
C1641 VDD2.n75 VSUBS 0.026841f
C1642 VDD2.n76 VSUBS 0.026841f
C1643 VDD2.n77 VSUBS 0.014423f
C1644 VDD2.n78 VSUBS 0.015272f
C1645 VDD2.n79 VSUBS 0.034091f
C1646 VDD2.n80 VSUBS 0.078661f
C1647 VDD2.n81 VSUBS 0.015272f
C1648 VDD2.n82 VSUBS 0.014423f
C1649 VDD2.n83 VSUBS 0.064608f
C1650 VDD2.n84 VSUBS 0.06716f
C1651 VDD2.t3 VSUBS 0.327279f
C1652 VDD2.t2 VSUBS 0.327279f
C1653 VDD2.n85 VSUBS 2.67104f
C1654 VDD2.n86 VSUBS 0.954515f
C1655 VDD2.t7 VSUBS 0.327279f
C1656 VDD2.t4 VSUBS 0.327279f
C1657 VDD2.n87 VSUBS 2.68804f
C1658 VDD2.n88 VSUBS 3.33618f
C1659 VDD2.n89 VSUBS 0.028356f
C1660 VDD2.n90 VSUBS 0.026841f
C1661 VDD2.n91 VSUBS 0.014423f
C1662 VDD2.n92 VSUBS 0.034091f
C1663 VDD2.n93 VSUBS 0.014847f
C1664 VDD2.n94 VSUBS 0.026841f
C1665 VDD2.n95 VSUBS 0.014847f
C1666 VDD2.n96 VSUBS 0.014423f
C1667 VDD2.n97 VSUBS 0.034091f
C1668 VDD2.n98 VSUBS 0.034091f
C1669 VDD2.n99 VSUBS 0.015272f
C1670 VDD2.n100 VSUBS 0.026841f
C1671 VDD2.n101 VSUBS 0.014423f
C1672 VDD2.n102 VSUBS 0.034091f
C1673 VDD2.n103 VSUBS 0.015272f
C1674 VDD2.n104 VSUBS 0.026841f
C1675 VDD2.n105 VSUBS 0.014423f
C1676 VDD2.n106 VSUBS 0.034091f
C1677 VDD2.n107 VSUBS 0.015272f
C1678 VDD2.n108 VSUBS 0.026841f
C1679 VDD2.n109 VSUBS 0.014423f
C1680 VDD2.n110 VSUBS 0.034091f
C1681 VDD2.n111 VSUBS 0.015272f
C1682 VDD2.n112 VSUBS 0.026841f
C1683 VDD2.n113 VSUBS 0.014423f
C1684 VDD2.n114 VSUBS 0.034091f
C1685 VDD2.n115 VSUBS 0.015272f
C1686 VDD2.n116 VSUBS 1.76625f
C1687 VDD2.n117 VSUBS 0.014423f
C1688 VDD2.t1 VSUBS 0.073011f
C1689 VDD2.n118 VSUBS 0.19261f
C1690 VDD2.n119 VSUBS 0.021687f
C1691 VDD2.n120 VSUBS 0.025568f
C1692 VDD2.n121 VSUBS 0.034091f
C1693 VDD2.n122 VSUBS 0.015272f
C1694 VDD2.n123 VSUBS 0.014423f
C1695 VDD2.n124 VSUBS 0.026841f
C1696 VDD2.n125 VSUBS 0.026841f
C1697 VDD2.n126 VSUBS 0.014423f
C1698 VDD2.n127 VSUBS 0.015272f
C1699 VDD2.n128 VSUBS 0.034091f
C1700 VDD2.n129 VSUBS 0.034091f
C1701 VDD2.n130 VSUBS 0.015272f
C1702 VDD2.n131 VSUBS 0.014423f
C1703 VDD2.n132 VSUBS 0.026841f
C1704 VDD2.n133 VSUBS 0.026841f
C1705 VDD2.n134 VSUBS 0.014423f
C1706 VDD2.n135 VSUBS 0.015272f
C1707 VDD2.n136 VSUBS 0.034091f
C1708 VDD2.n137 VSUBS 0.034091f
C1709 VDD2.n138 VSUBS 0.015272f
C1710 VDD2.n139 VSUBS 0.014423f
C1711 VDD2.n140 VSUBS 0.026841f
C1712 VDD2.n141 VSUBS 0.026841f
C1713 VDD2.n142 VSUBS 0.014423f
C1714 VDD2.n143 VSUBS 0.015272f
C1715 VDD2.n144 VSUBS 0.034091f
C1716 VDD2.n145 VSUBS 0.034091f
C1717 VDD2.n146 VSUBS 0.015272f
C1718 VDD2.n147 VSUBS 0.014423f
C1719 VDD2.n148 VSUBS 0.026841f
C1720 VDD2.n149 VSUBS 0.026841f
C1721 VDD2.n150 VSUBS 0.014423f
C1722 VDD2.n151 VSUBS 0.015272f
C1723 VDD2.n152 VSUBS 0.034091f
C1724 VDD2.n153 VSUBS 0.034091f
C1725 VDD2.n154 VSUBS 0.015272f
C1726 VDD2.n155 VSUBS 0.014423f
C1727 VDD2.n156 VSUBS 0.026841f
C1728 VDD2.n157 VSUBS 0.026841f
C1729 VDD2.n158 VSUBS 0.014423f
C1730 VDD2.n159 VSUBS 0.015272f
C1731 VDD2.n160 VSUBS 0.034091f
C1732 VDD2.n161 VSUBS 0.034091f
C1733 VDD2.n162 VSUBS 0.015272f
C1734 VDD2.n163 VSUBS 0.014423f
C1735 VDD2.n164 VSUBS 0.026841f
C1736 VDD2.n165 VSUBS 0.026841f
C1737 VDD2.n166 VSUBS 0.014423f
C1738 VDD2.n167 VSUBS 0.015272f
C1739 VDD2.n168 VSUBS 0.034091f
C1740 VDD2.n169 VSUBS 0.078661f
C1741 VDD2.n170 VSUBS 0.015272f
C1742 VDD2.n171 VSUBS 0.014423f
C1743 VDD2.n172 VSUBS 0.064608f
C1744 VDD2.n173 VSUBS 0.057977f
C1745 VDD2.n174 VSUBS 3.16613f
C1746 VDD2.t0 VSUBS 0.327279f
C1747 VDD2.t5 VSUBS 0.327279f
C1748 VDD2.n175 VSUBS 2.67105f
C1749 VDD2.n176 VSUBS 0.740065f
C1750 VDD2.t8 VSUBS 0.327279f
C1751 VDD2.t9 VSUBS 0.327279f
C1752 VDD2.n177 VSUBS 2.688f
C1753 VN.n0 VSUBS 0.03951f
C1754 VN.t7 VSUBS 2.62454f
C1755 VN.n1 VSUBS 0.02831f
C1756 VN.n2 VSUBS 0.029968f
C1757 VN.t8 VSUBS 2.62454f
C1758 VN.n3 VSUBS 0.047924f
C1759 VN.n4 VSUBS 0.029968f
C1760 VN.t1 VSUBS 2.62454f
C1761 VN.n5 VSUBS 0.055853f
C1762 VN.n6 VSUBS 0.029968f
C1763 VN.t0 VSUBS 2.62454f
C1764 VN.n7 VSUBS 1.00433f
C1765 VN.t9 VSUBS 2.79132f
C1766 VN.n8 VSUBS 0.990423f
C1767 VN.n9 VSUBS 0.251329f
C1768 VN.n10 VSUBS 0.050338f
C1769 VN.n11 VSUBS 0.047924f
C1770 VN.n12 VSUBS 0.039573f
C1771 VN.n13 VSUBS 0.029968f
C1772 VN.n14 VSUBS 0.029968f
C1773 VN.n15 VSUBS 0.029968f
C1774 VN.n16 VSUBS 0.950016f
C1775 VN.n17 VSUBS 0.055853f
C1776 VN.n18 VSUBS 0.039573f
C1777 VN.n19 VSUBS 0.029968f
C1778 VN.n20 VSUBS 0.029968f
C1779 VN.n21 VSUBS 0.029968f
C1780 VN.n22 VSUBS 0.050338f
C1781 VN.n23 VSUBS 0.921738f
C1782 VN.n24 VSUBS 0.033793f
C1783 VN.n25 VSUBS 0.060037f
C1784 VN.n26 VSUBS 0.029968f
C1785 VN.n27 VSUBS 0.029968f
C1786 VN.n28 VSUBS 0.029968f
C1787 VN.n29 VSUBS 0.055002f
C1788 VN.n30 VSUBS 0.044823f
C1789 VN.n31 VSUBS 1.00791f
C1790 VN.n32 VSUBS 0.040836f
C1791 VN.n33 VSUBS 0.03951f
C1792 VN.t2 VSUBS 2.62454f
C1793 VN.n34 VSUBS 0.02831f
C1794 VN.n35 VSUBS 0.029968f
C1795 VN.t3 VSUBS 2.62454f
C1796 VN.n36 VSUBS 0.047924f
C1797 VN.n37 VSUBS 0.029968f
C1798 VN.t6 VSUBS 2.62454f
C1799 VN.n38 VSUBS 0.055853f
C1800 VN.n39 VSUBS 0.029968f
C1801 VN.t5 VSUBS 2.62454f
C1802 VN.n40 VSUBS 1.00433f
C1803 VN.t4 VSUBS 2.79132f
C1804 VN.n41 VSUBS 0.990423f
C1805 VN.n42 VSUBS 0.251329f
C1806 VN.n43 VSUBS 0.050338f
C1807 VN.n44 VSUBS 0.047924f
C1808 VN.n45 VSUBS 0.039573f
C1809 VN.n46 VSUBS 0.029968f
C1810 VN.n47 VSUBS 0.029968f
C1811 VN.n48 VSUBS 0.029968f
C1812 VN.n49 VSUBS 0.950016f
C1813 VN.n50 VSUBS 0.055853f
C1814 VN.n51 VSUBS 0.039573f
C1815 VN.n52 VSUBS 0.029968f
C1816 VN.n53 VSUBS 0.029968f
C1817 VN.n54 VSUBS 0.029968f
C1818 VN.n55 VSUBS 0.050338f
C1819 VN.n56 VSUBS 0.921738f
C1820 VN.n57 VSUBS 0.033793f
C1821 VN.n58 VSUBS 0.060037f
C1822 VN.n59 VSUBS 0.029968f
C1823 VN.n60 VSUBS 0.029968f
C1824 VN.n61 VSUBS 0.029968f
C1825 VN.n62 VSUBS 0.055002f
C1826 VN.n63 VSUBS 0.044823f
C1827 VN.n64 VSUBS 1.00791f
C1828 VN.n65 VSUBS 1.81101f
.ends

