* NGSPICE file created from diff_pair_sample_1698.ext - technology: sky130A

.subckt diff_pair_sample_1698 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9748 pd=31.42 as=0 ps=0 w=15.32 l=2.64
X1 VTAIL.t7 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=5.9748 pd=31.42 as=2.5278 ps=15.65 w=15.32 l=2.64
X2 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9748 pd=31.42 as=0 ps=0 w=15.32 l=2.64
X3 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9748 pd=31.42 as=0 ps=0 w=15.32 l=2.64
X4 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9748 pd=31.42 as=0 ps=0 w=15.32 l=2.64
X5 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9748 pd=31.42 as=2.5278 ps=15.65 w=15.32 l=2.64
X6 VDD2.t2 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5278 pd=15.65 as=5.9748 ps=31.42 w=15.32 l=2.64
X7 VDD1.t0 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5278 pd=15.65 as=5.9748 ps=31.42 w=15.32 l=2.64
X8 VTAIL.t2 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.9748 pd=31.42 as=2.5278 ps=15.65 w=15.32 l=2.64
X9 VDD2.t0 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5278 pd=15.65 as=5.9748 ps=31.42 w=15.32 l=2.64
X10 VTAIL.t5 VP.t2 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9748 pd=31.42 as=2.5278 ps=15.65 w=15.32 l=2.64
X11 VDD1.t1 VP.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5278 pd=15.65 as=5.9748 ps=31.42 w=15.32 l=2.64
R0 B.n626 B.n625 585
R1 B.n628 B.n126 585
R2 B.n631 B.n630 585
R3 B.n632 B.n125 585
R4 B.n634 B.n633 585
R5 B.n636 B.n124 585
R6 B.n639 B.n638 585
R7 B.n640 B.n123 585
R8 B.n642 B.n641 585
R9 B.n644 B.n122 585
R10 B.n647 B.n646 585
R11 B.n648 B.n121 585
R12 B.n650 B.n649 585
R13 B.n652 B.n120 585
R14 B.n655 B.n654 585
R15 B.n656 B.n119 585
R16 B.n658 B.n657 585
R17 B.n660 B.n118 585
R18 B.n663 B.n662 585
R19 B.n664 B.n117 585
R20 B.n666 B.n665 585
R21 B.n668 B.n116 585
R22 B.n671 B.n670 585
R23 B.n672 B.n115 585
R24 B.n674 B.n673 585
R25 B.n676 B.n114 585
R26 B.n679 B.n678 585
R27 B.n680 B.n113 585
R28 B.n682 B.n681 585
R29 B.n684 B.n112 585
R30 B.n687 B.n686 585
R31 B.n688 B.n111 585
R32 B.n690 B.n689 585
R33 B.n692 B.n110 585
R34 B.n695 B.n694 585
R35 B.n696 B.n109 585
R36 B.n698 B.n697 585
R37 B.n700 B.n108 585
R38 B.n703 B.n702 585
R39 B.n704 B.n107 585
R40 B.n706 B.n705 585
R41 B.n708 B.n106 585
R42 B.n711 B.n710 585
R43 B.n712 B.n105 585
R44 B.n714 B.n713 585
R45 B.n716 B.n104 585
R46 B.n719 B.n718 585
R47 B.n720 B.n103 585
R48 B.n722 B.n721 585
R49 B.n724 B.n102 585
R50 B.n727 B.n726 585
R51 B.n729 B.n99 585
R52 B.n731 B.n730 585
R53 B.n733 B.n98 585
R54 B.n736 B.n735 585
R55 B.n737 B.n97 585
R56 B.n739 B.n738 585
R57 B.n741 B.n96 585
R58 B.n744 B.n743 585
R59 B.n745 B.n92 585
R60 B.n747 B.n746 585
R61 B.n749 B.n91 585
R62 B.n752 B.n751 585
R63 B.n753 B.n90 585
R64 B.n755 B.n754 585
R65 B.n757 B.n89 585
R66 B.n760 B.n759 585
R67 B.n761 B.n88 585
R68 B.n763 B.n762 585
R69 B.n765 B.n87 585
R70 B.n768 B.n767 585
R71 B.n769 B.n86 585
R72 B.n771 B.n770 585
R73 B.n773 B.n85 585
R74 B.n776 B.n775 585
R75 B.n777 B.n84 585
R76 B.n779 B.n778 585
R77 B.n781 B.n83 585
R78 B.n784 B.n783 585
R79 B.n785 B.n82 585
R80 B.n787 B.n786 585
R81 B.n789 B.n81 585
R82 B.n792 B.n791 585
R83 B.n793 B.n80 585
R84 B.n795 B.n794 585
R85 B.n797 B.n79 585
R86 B.n800 B.n799 585
R87 B.n801 B.n78 585
R88 B.n803 B.n802 585
R89 B.n805 B.n77 585
R90 B.n808 B.n807 585
R91 B.n809 B.n76 585
R92 B.n811 B.n810 585
R93 B.n813 B.n75 585
R94 B.n816 B.n815 585
R95 B.n817 B.n74 585
R96 B.n819 B.n818 585
R97 B.n821 B.n73 585
R98 B.n824 B.n823 585
R99 B.n825 B.n72 585
R100 B.n827 B.n826 585
R101 B.n829 B.n71 585
R102 B.n832 B.n831 585
R103 B.n833 B.n70 585
R104 B.n835 B.n834 585
R105 B.n837 B.n69 585
R106 B.n840 B.n839 585
R107 B.n841 B.n68 585
R108 B.n843 B.n842 585
R109 B.n845 B.n67 585
R110 B.n848 B.n847 585
R111 B.n849 B.n66 585
R112 B.n624 B.n64 585
R113 B.n852 B.n64 585
R114 B.n623 B.n63 585
R115 B.n853 B.n63 585
R116 B.n622 B.n62 585
R117 B.n854 B.n62 585
R118 B.n621 B.n620 585
R119 B.n620 B.n58 585
R120 B.n619 B.n57 585
R121 B.n860 B.n57 585
R122 B.n618 B.n56 585
R123 B.n861 B.n56 585
R124 B.n617 B.n55 585
R125 B.n862 B.n55 585
R126 B.n616 B.n615 585
R127 B.n615 B.n54 585
R128 B.n614 B.n50 585
R129 B.n868 B.n50 585
R130 B.n613 B.n49 585
R131 B.n869 B.n49 585
R132 B.n612 B.n48 585
R133 B.n870 B.n48 585
R134 B.n611 B.n610 585
R135 B.n610 B.n44 585
R136 B.n609 B.n43 585
R137 B.n876 B.n43 585
R138 B.n608 B.n42 585
R139 B.n877 B.n42 585
R140 B.n607 B.n41 585
R141 B.n878 B.n41 585
R142 B.n606 B.n605 585
R143 B.n605 B.n37 585
R144 B.n604 B.n36 585
R145 B.n884 B.n36 585
R146 B.n603 B.n35 585
R147 B.n885 B.n35 585
R148 B.n602 B.n34 585
R149 B.n886 B.n34 585
R150 B.n601 B.n600 585
R151 B.n600 B.n33 585
R152 B.n599 B.n29 585
R153 B.n892 B.n29 585
R154 B.n598 B.n28 585
R155 B.n893 B.n28 585
R156 B.n597 B.n27 585
R157 B.n894 B.n27 585
R158 B.n596 B.n595 585
R159 B.n595 B.n23 585
R160 B.n594 B.n22 585
R161 B.n900 B.n22 585
R162 B.n593 B.n21 585
R163 B.n901 B.n21 585
R164 B.n592 B.n20 585
R165 B.n902 B.n20 585
R166 B.n591 B.n590 585
R167 B.n590 B.n16 585
R168 B.n589 B.n15 585
R169 B.n908 B.n15 585
R170 B.n588 B.n14 585
R171 B.n909 B.n14 585
R172 B.n587 B.n13 585
R173 B.n910 B.n13 585
R174 B.n586 B.n585 585
R175 B.n585 B.n12 585
R176 B.n584 B.n583 585
R177 B.n584 B.n8 585
R178 B.n582 B.n7 585
R179 B.n917 B.n7 585
R180 B.n581 B.n6 585
R181 B.n918 B.n6 585
R182 B.n580 B.n5 585
R183 B.n919 B.n5 585
R184 B.n579 B.n578 585
R185 B.n578 B.n4 585
R186 B.n577 B.n127 585
R187 B.n577 B.n576 585
R188 B.n567 B.n128 585
R189 B.n129 B.n128 585
R190 B.n569 B.n568 585
R191 B.n570 B.n569 585
R192 B.n566 B.n134 585
R193 B.n134 B.n133 585
R194 B.n565 B.n564 585
R195 B.n564 B.n563 585
R196 B.n136 B.n135 585
R197 B.n137 B.n136 585
R198 B.n556 B.n555 585
R199 B.n557 B.n556 585
R200 B.n554 B.n142 585
R201 B.n142 B.n141 585
R202 B.n553 B.n552 585
R203 B.n552 B.n551 585
R204 B.n144 B.n143 585
R205 B.n145 B.n144 585
R206 B.n544 B.n543 585
R207 B.n545 B.n544 585
R208 B.n542 B.n150 585
R209 B.n150 B.n149 585
R210 B.n541 B.n540 585
R211 B.n540 B.n539 585
R212 B.n152 B.n151 585
R213 B.n532 B.n152 585
R214 B.n531 B.n530 585
R215 B.n533 B.n531 585
R216 B.n529 B.n157 585
R217 B.n157 B.n156 585
R218 B.n528 B.n527 585
R219 B.n527 B.n526 585
R220 B.n159 B.n158 585
R221 B.n160 B.n159 585
R222 B.n519 B.n518 585
R223 B.n520 B.n519 585
R224 B.n517 B.n165 585
R225 B.n165 B.n164 585
R226 B.n516 B.n515 585
R227 B.n515 B.n514 585
R228 B.n167 B.n166 585
R229 B.n168 B.n167 585
R230 B.n507 B.n506 585
R231 B.n508 B.n507 585
R232 B.n505 B.n173 585
R233 B.n173 B.n172 585
R234 B.n504 B.n503 585
R235 B.n503 B.n502 585
R236 B.n175 B.n174 585
R237 B.n495 B.n175 585
R238 B.n494 B.n493 585
R239 B.n496 B.n494 585
R240 B.n492 B.n180 585
R241 B.n180 B.n179 585
R242 B.n491 B.n490 585
R243 B.n490 B.n489 585
R244 B.n182 B.n181 585
R245 B.n183 B.n182 585
R246 B.n482 B.n481 585
R247 B.n483 B.n482 585
R248 B.n480 B.n188 585
R249 B.n188 B.n187 585
R250 B.n479 B.n478 585
R251 B.n478 B.n477 585
R252 B.n474 B.n192 585
R253 B.n473 B.n472 585
R254 B.n470 B.n193 585
R255 B.n470 B.n191 585
R256 B.n469 B.n468 585
R257 B.n467 B.n466 585
R258 B.n465 B.n195 585
R259 B.n463 B.n462 585
R260 B.n461 B.n196 585
R261 B.n460 B.n459 585
R262 B.n457 B.n197 585
R263 B.n455 B.n454 585
R264 B.n453 B.n198 585
R265 B.n452 B.n451 585
R266 B.n449 B.n199 585
R267 B.n447 B.n446 585
R268 B.n445 B.n200 585
R269 B.n444 B.n443 585
R270 B.n441 B.n201 585
R271 B.n439 B.n438 585
R272 B.n437 B.n202 585
R273 B.n436 B.n435 585
R274 B.n433 B.n203 585
R275 B.n431 B.n430 585
R276 B.n429 B.n204 585
R277 B.n428 B.n427 585
R278 B.n425 B.n205 585
R279 B.n423 B.n422 585
R280 B.n421 B.n206 585
R281 B.n420 B.n419 585
R282 B.n417 B.n207 585
R283 B.n415 B.n414 585
R284 B.n413 B.n208 585
R285 B.n412 B.n411 585
R286 B.n409 B.n209 585
R287 B.n407 B.n406 585
R288 B.n405 B.n210 585
R289 B.n404 B.n403 585
R290 B.n401 B.n211 585
R291 B.n399 B.n398 585
R292 B.n397 B.n212 585
R293 B.n396 B.n395 585
R294 B.n393 B.n213 585
R295 B.n391 B.n390 585
R296 B.n389 B.n214 585
R297 B.n388 B.n387 585
R298 B.n385 B.n215 585
R299 B.n383 B.n382 585
R300 B.n381 B.n216 585
R301 B.n380 B.n379 585
R302 B.n377 B.n217 585
R303 B.n375 B.n374 585
R304 B.n372 B.n218 585
R305 B.n371 B.n370 585
R306 B.n368 B.n221 585
R307 B.n366 B.n365 585
R308 B.n364 B.n222 585
R309 B.n363 B.n362 585
R310 B.n360 B.n223 585
R311 B.n358 B.n357 585
R312 B.n356 B.n224 585
R313 B.n355 B.n354 585
R314 B.n352 B.n351 585
R315 B.n350 B.n349 585
R316 B.n348 B.n229 585
R317 B.n346 B.n345 585
R318 B.n344 B.n230 585
R319 B.n343 B.n342 585
R320 B.n340 B.n231 585
R321 B.n338 B.n337 585
R322 B.n336 B.n232 585
R323 B.n335 B.n334 585
R324 B.n332 B.n233 585
R325 B.n330 B.n329 585
R326 B.n328 B.n234 585
R327 B.n327 B.n326 585
R328 B.n324 B.n235 585
R329 B.n322 B.n321 585
R330 B.n320 B.n236 585
R331 B.n319 B.n318 585
R332 B.n316 B.n237 585
R333 B.n314 B.n313 585
R334 B.n312 B.n238 585
R335 B.n311 B.n310 585
R336 B.n308 B.n239 585
R337 B.n306 B.n305 585
R338 B.n304 B.n240 585
R339 B.n303 B.n302 585
R340 B.n300 B.n241 585
R341 B.n298 B.n297 585
R342 B.n296 B.n242 585
R343 B.n295 B.n294 585
R344 B.n292 B.n243 585
R345 B.n290 B.n289 585
R346 B.n288 B.n244 585
R347 B.n287 B.n286 585
R348 B.n284 B.n245 585
R349 B.n282 B.n281 585
R350 B.n280 B.n246 585
R351 B.n279 B.n278 585
R352 B.n276 B.n247 585
R353 B.n274 B.n273 585
R354 B.n272 B.n248 585
R355 B.n271 B.n270 585
R356 B.n268 B.n249 585
R357 B.n266 B.n265 585
R358 B.n264 B.n250 585
R359 B.n263 B.n262 585
R360 B.n260 B.n251 585
R361 B.n258 B.n257 585
R362 B.n256 B.n252 585
R363 B.n255 B.n254 585
R364 B.n190 B.n189 585
R365 B.n191 B.n190 585
R366 B.n476 B.n475 585
R367 B.n477 B.n476 585
R368 B.n186 B.n185 585
R369 B.n187 B.n186 585
R370 B.n485 B.n484 585
R371 B.n484 B.n483 585
R372 B.n486 B.n184 585
R373 B.n184 B.n183 585
R374 B.n488 B.n487 585
R375 B.n489 B.n488 585
R376 B.n178 B.n177 585
R377 B.n179 B.n178 585
R378 B.n498 B.n497 585
R379 B.n497 B.n496 585
R380 B.n499 B.n176 585
R381 B.n495 B.n176 585
R382 B.n501 B.n500 585
R383 B.n502 B.n501 585
R384 B.n171 B.n170 585
R385 B.n172 B.n171 585
R386 B.n510 B.n509 585
R387 B.n509 B.n508 585
R388 B.n511 B.n169 585
R389 B.n169 B.n168 585
R390 B.n513 B.n512 585
R391 B.n514 B.n513 585
R392 B.n163 B.n162 585
R393 B.n164 B.n163 585
R394 B.n522 B.n521 585
R395 B.n521 B.n520 585
R396 B.n523 B.n161 585
R397 B.n161 B.n160 585
R398 B.n525 B.n524 585
R399 B.n526 B.n525 585
R400 B.n155 B.n154 585
R401 B.n156 B.n155 585
R402 B.n535 B.n534 585
R403 B.n534 B.n533 585
R404 B.n536 B.n153 585
R405 B.n532 B.n153 585
R406 B.n538 B.n537 585
R407 B.n539 B.n538 585
R408 B.n148 B.n147 585
R409 B.n149 B.n148 585
R410 B.n547 B.n546 585
R411 B.n546 B.n545 585
R412 B.n548 B.n146 585
R413 B.n146 B.n145 585
R414 B.n550 B.n549 585
R415 B.n551 B.n550 585
R416 B.n140 B.n139 585
R417 B.n141 B.n140 585
R418 B.n559 B.n558 585
R419 B.n558 B.n557 585
R420 B.n560 B.n138 585
R421 B.n138 B.n137 585
R422 B.n562 B.n561 585
R423 B.n563 B.n562 585
R424 B.n132 B.n131 585
R425 B.n133 B.n132 585
R426 B.n572 B.n571 585
R427 B.n571 B.n570 585
R428 B.n573 B.n130 585
R429 B.n130 B.n129 585
R430 B.n575 B.n574 585
R431 B.n576 B.n575 585
R432 B.n3 B.n0 585
R433 B.n4 B.n3 585
R434 B.n916 B.n1 585
R435 B.n917 B.n916 585
R436 B.n915 B.n914 585
R437 B.n915 B.n8 585
R438 B.n913 B.n9 585
R439 B.n12 B.n9 585
R440 B.n912 B.n911 585
R441 B.n911 B.n910 585
R442 B.n11 B.n10 585
R443 B.n909 B.n11 585
R444 B.n907 B.n906 585
R445 B.n908 B.n907 585
R446 B.n905 B.n17 585
R447 B.n17 B.n16 585
R448 B.n904 B.n903 585
R449 B.n903 B.n902 585
R450 B.n19 B.n18 585
R451 B.n901 B.n19 585
R452 B.n899 B.n898 585
R453 B.n900 B.n899 585
R454 B.n897 B.n24 585
R455 B.n24 B.n23 585
R456 B.n896 B.n895 585
R457 B.n895 B.n894 585
R458 B.n26 B.n25 585
R459 B.n893 B.n26 585
R460 B.n891 B.n890 585
R461 B.n892 B.n891 585
R462 B.n889 B.n30 585
R463 B.n33 B.n30 585
R464 B.n888 B.n887 585
R465 B.n887 B.n886 585
R466 B.n32 B.n31 585
R467 B.n885 B.n32 585
R468 B.n883 B.n882 585
R469 B.n884 B.n883 585
R470 B.n881 B.n38 585
R471 B.n38 B.n37 585
R472 B.n880 B.n879 585
R473 B.n879 B.n878 585
R474 B.n40 B.n39 585
R475 B.n877 B.n40 585
R476 B.n875 B.n874 585
R477 B.n876 B.n875 585
R478 B.n873 B.n45 585
R479 B.n45 B.n44 585
R480 B.n872 B.n871 585
R481 B.n871 B.n870 585
R482 B.n47 B.n46 585
R483 B.n869 B.n47 585
R484 B.n867 B.n866 585
R485 B.n868 B.n867 585
R486 B.n865 B.n51 585
R487 B.n54 B.n51 585
R488 B.n864 B.n863 585
R489 B.n863 B.n862 585
R490 B.n53 B.n52 585
R491 B.n861 B.n53 585
R492 B.n859 B.n858 585
R493 B.n860 B.n859 585
R494 B.n857 B.n59 585
R495 B.n59 B.n58 585
R496 B.n856 B.n855 585
R497 B.n855 B.n854 585
R498 B.n61 B.n60 585
R499 B.n853 B.n61 585
R500 B.n851 B.n850 585
R501 B.n852 B.n851 585
R502 B.n920 B.n919 585
R503 B.n918 B.n2 585
R504 B.n851 B.n66 497.305
R505 B.n626 B.n64 497.305
R506 B.n478 B.n190 497.305
R507 B.n476 B.n192 497.305
R508 B.n100 B.t16 396.618
R509 B.n225 B.t14 396.618
R510 B.n93 B.t10 396.618
R511 B.n219 B.t7 396.618
R512 B.n93 B.t8 347.959
R513 B.n100 B.t15 347.959
R514 B.n225 B.t12 347.959
R515 B.n219 B.t4 347.959
R516 B.n101 B.t17 339.019
R517 B.n226 B.t13 339.019
R518 B.n94 B.t11 339.019
R519 B.n220 B.t6 339.019
R520 B.n627 B.n65 256.663
R521 B.n629 B.n65 256.663
R522 B.n635 B.n65 256.663
R523 B.n637 B.n65 256.663
R524 B.n643 B.n65 256.663
R525 B.n645 B.n65 256.663
R526 B.n651 B.n65 256.663
R527 B.n653 B.n65 256.663
R528 B.n659 B.n65 256.663
R529 B.n661 B.n65 256.663
R530 B.n667 B.n65 256.663
R531 B.n669 B.n65 256.663
R532 B.n675 B.n65 256.663
R533 B.n677 B.n65 256.663
R534 B.n683 B.n65 256.663
R535 B.n685 B.n65 256.663
R536 B.n691 B.n65 256.663
R537 B.n693 B.n65 256.663
R538 B.n699 B.n65 256.663
R539 B.n701 B.n65 256.663
R540 B.n707 B.n65 256.663
R541 B.n709 B.n65 256.663
R542 B.n715 B.n65 256.663
R543 B.n717 B.n65 256.663
R544 B.n723 B.n65 256.663
R545 B.n725 B.n65 256.663
R546 B.n732 B.n65 256.663
R547 B.n734 B.n65 256.663
R548 B.n740 B.n65 256.663
R549 B.n742 B.n65 256.663
R550 B.n748 B.n65 256.663
R551 B.n750 B.n65 256.663
R552 B.n756 B.n65 256.663
R553 B.n758 B.n65 256.663
R554 B.n764 B.n65 256.663
R555 B.n766 B.n65 256.663
R556 B.n772 B.n65 256.663
R557 B.n774 B.n65 256.663
R558 B.n780 B.n65 256.663
R559 B.n782 B.n65 256.663
R560 B.n788 B.n65 256.663
R561 B.n790 B.n65 256.663
R562 B.n796 B.n65 256.663
R563 B.n798 B.n65 256.663
R564 B.n804 B.n65 256.663
R565 B.n806 B.n65 256.663
R566 B.n812 B.n65 256.663
R567 B.n814 B.n65 256.663
R568 B.n820 B.n65 256.663
R569 B.n822 B.n65 256.663
R570 B.n828 B.n65 256.663
R571 B.n830 B.n65 256.663
R572 B.n836 B.n65 256.663
R573 B.n838 B.n65 256.663
R574 B.n844 B.n65 256.663
R575 B.n846 B.n65 256.663
R576 B.n471 B.n191 256.663
R577 B.n194 B.n191 256.663
R578 B.n464 B.n191 256.663
R579 B.n458 B.n191 256.663
R580 B.n456 B.n191 256.663
R581 B.n450 B.n191 256.663
R582 B.n448 B.n191 256.663
R583 B.n442 B.n191 256.663
R584 B.n440 B.n191 256.663
R585 B.n434 B.n191 256.663
R586 B.n432 B.n191 256.663
R587 B.n426 B.n191 256.663
R588 B.n424 B.n191 256.663
R589 B.n418 B.n191 256.663
R590 B.n416 B.n191 256.663
R591 B.n410 B.n191 256.663
R592 B.n408 B.n191 256.663
R593 B.n402 B.n191 256.663
R594 B.n400 B.n191 256.663
R595 B.n394 B.n191 256.663
R596 B.n392 B.n191 256.663
R597 B.n386 B.n191 256.663
R598 B.n384 B.n191 256.663
R599 B.n378 B.n191 256.663
R600 B.n376 B.n191 256.663
R601 B.n369 B.n191 256.663
R602 B.n367 B.n191 256.663
R603 B.n361 B.n191 256.663
R604 B.n359 B.n191 256.663
R605 B.n353 B.n191 256.663
R606 B.n228 B.n191 256.663
R607 B.n347 B.n191 256.663
R608 B.n341 B.n191 256.663
R609 B.n339 B.n191 256.663
R610 B.n333 B.n191 256.663
R611 B.n331 B.n191 256.663
R612 B.n325 B.n191 256.663
R613 B.n323 B.n191 256.663
R614 B.n317 B.n191 256.663
R615 B.n315 B.n191 256.663
R616 B.n309 B.n191 256.663
R617 B.n307 B.n191 256.663
R618 B.n301 B.n191 256.663
R619 B.n299 B.n191 256.663
R620 B.n293 B.n191 256.663
R621 B.n291 B.n191 256.663
R622 B.n285 B.n191 256.663
R623 B.n283 B.n191 256.663
R624 B.n277 B.n191 256.663
R625 B.n275 B.n191 256.663
R626 B.n269 B.n191 256.663
R627 B.n267 B.n191 256.663
R628 B.n261 B.n191 256.663
R629 B.n259 B.n191 256.663
R630 B.n253 B.n191 256.663
R631 B.n922 B.n921 256.663
R632 B.n847 B.n845 163.367
R633 B.n843 B.n68 163.367
R634 B.n839 B.n837 163.367
R635 B.n835 B.n70 163.367
R636 B.n831 B.n829 163.367
R637 B.n827 B.n72 163.367
R638 B.n823 B.n821 163.367
R639 B.n819 B.n74 163.367
R640 B.n815 B.n813 163.367
R641 B.n811 B.n76 163.367
R642 B.n807 B.n805 163.367
R643 B.n803 B.n78 163.367
R644 B.n799 B.n797 163.367
R645 B.n795 B.n80 163.367
R646 B.n791 B.n789 163.367
R647 B.n787 B.n82 163.367
R648 B.n783 B.n781 163.367
R649 B.n779 B.n84 163.367
R650 B.n775 B.n773 163.367
R651 B.n771 B.n86 163.367
R652 B.n767 B.n765 163.367
R653 B.n763 B.n88 163.367
R654 B.n759 B.n757 163.367
R655 B.n755 B.n90 163.367
R656 B.n751 B.n749 163.367
R657 B.n747 B.n92 163.367
R658 B.n743 B.n741 163.367
R659 B.n739 B.n97 163.367
R660 B.n735 B.n733 163.367
R661 B.n731 B.n99 163.367
R662 B.n726 B.n724 163.367
R663 B.n722 B.n103 163.367
R664 B.n718 B.n716 163.367
R665 B.n714 B.n105 163.367
R666 B.n710 B.n708 163.367
R667 B.n706 B.n107 163.367
R668 B.n702 B.n700 163.367
R669 B.n698 B.n109 163.367
R670 B.n694 B.n692 163.367
R671 B.n690 B.n111 163.367
R672 B.n686 B.n684 163.367
R673 B.n682 B.n113 163.367
R674 B.n678 B.n676 163.367
R675 B.n674 B.n115 163.367
R676 B.n670 B.n668 163.367
R677 B.n666 B.n117 163.367
R678 B.n662 B.n660 163.367
R679 B.n658 B.n119 163.367
R680 B.n654 B.n652 163.367
R681 B.n650 B.n121 163.367
R682 B.n646 B.n644 163.367
R683 B.n642 B.n123 163.367
R684 B.n638 B.n636 163.367
R685 B.n634 B.n125 163.367
R686 B.n630 B.n628 163.367
R687 B.n478 B.n188 163.367
R688 B.n482 B.n188 163.367
R689 B.n482 B.n182 163.367
R690 B.n490 B.n182 163.367
R691 B.n490 B.n180 163.367
R692 B.n494 B.n180 163.367
R693 B.n494 B.n175 163.367
R694 B.n503 B.n175 163.367
R695 B.n503 B.n173 163.367
R696 B.n507 B.n173 163.367
R697 B.n507 B.n167 163.367
R698 B.n515 B.n167 163.367
R699 B.n515 B.n165 163.367
R700 B.n519 B.n165 163.367
R701 B.n519 B.n159 163.367
R702 B.n527 B.n159 163.367
R703 B.n527 B.n157 163.367
R704 B.n531 B.n157 163.367
R705 B.n531 B.n152 163.367
R706 B.n540 B.n152 163.367
R707 B.n540 B.n150 163.367
R708 B.n544 B.n150 163.367
R709 B.n544 B.n144 163.367
R710 B.n552 B.n144 163.367
R711 B.n552 B.n142 163.367
R712 B.n556 B.n142 163.367
R713 B.n556 B.n136 163.367
R714 B.n564 B.n136 163.367
R715 B.n564 B.n134 163.367
R716 B.n569 B.n134 163.367
R717 B.n569 B.n128 163.367
R718 B.n577 B.n128 163.367
R719 B.n578 B.n577 163.367
R720 B.n578 B.n5 163.367
R721 B.n6 B.n5 163.367
R722 B.n7 B.n6 163.367
R723 B.n584 B.n7 163.367
R724 B.n585 B.n584 163.367
R725 B.n585 B.n13 163.367
R726 B.n14 B.n13 163.367
R727 B.n15 B.n14 163.367
R728 B.n590 B.n15 163.367
R729 B.n590 B.n20 163.367
R730 B.n21 B.n20 163.367
R731 B.n22 B.n21 163.367
R732 B.n595 B.n22 163.367
R733 B.n595 B.n27 163.367
R734 B.n28 B.n27 163.367
R735 B.n29 B.n28 163.367
R736 B.n600 B.n29 163.367
R737 B.n600 B.n34 163.367
R738 B.n35 B.n34 163.367
R739 B.n36 B.n35 163.367
R740 B.n605 B.n36 163.367
R741 B.n605 B.n41 163.367
R742 B.n42 B.n41 163.367
R743 B.n43 B.n42 163.367
R744 B.n610 B.n43 163.367
R745 B.n610 B.n48 163.367
R746 B.n49 B.n48 163.367
R747 B.n50 B.n49 163.367
R748 B.n615 B.n50 163.367
R749 B.n615 B.n55 163.367
R750 B.n56 B.n55 163.367
R751 B.n57 B.n56 163.367
R752 B.n620 B.n57 163.367
R753 B.n620 B.n62 163.367
R754 B.n63 B.n62 163.367
R755 B.n64 B.n63 163.367
R756 B.n472 B.n470 163.367
R757 B.n470 B.n469 163.367
R758 B.n466 B.n465 163.367
R759 B.n463 B.n196 163.367
R760 B.n459 B.n457 163.367
R761 B.n455 B.n198 163.367
R762 B.n451 B.n449 163.367
R763 B.n447 B.n200 163.367
R764 B.n443 B.n441 163.367
R765 B.n439 B.n202 163.367
R766 B.n435 B.n433 163.367
R767 B.n431 B.n204 163.367
R768 B.n427 B.n425 163.367
R769 B.n423 B.n206 163.367
R770 B.n419 B.n417 163.367
R771 B.n415 B.n208 163.367
R772 B.n411 B.n409 163.367
R773 B.n407 B.n210 163.367
R774 B.n403 B.n401 163.367
R775 B.n399 B.n212 163.367
R776 B.n395 B.n393 163.367
R777 B.n391 B.n214 163.367
R778 B.n387 B.n385 163.367
R779 B.n383 B.n216 163.367
R780 B.n379 B.n377 163.367
R781 B.n375 B.n218 163.367
R782 B.n370 B.n368 163.367
R783 B.n366 B.n222 163.367
R784 B.n362 B.n360 163.367
R785 B.n358 B.n224 163.367
R786 B.n354 B.n352 163.367
R787 B.n349 B.n348 163.367
R788 B.n346 B.n230 163.367
R789 B.n342 B.n340 163.367
R790 B.n338 B.n232 163.367
R791 B.n334 B.n332 163.367
R792 B.n330 B.n234 163.367
R793 B.n326 B.n324 163.367
R794 B.n322 B.n236 163.367
R795 B.n318 B.n316 163.367
R796 B.n314 B.n238 163.367
R797 B.n310 B.n308 163.367
R798 B.n306 B.n240 163.367
R799 B.n302 B.n300 163.367
R800 B.n298 B.n242 163.367
R801 B.n294 B.n292 163.367
R802 B.n290 B.n244 163.367
R803 B.n286 B.n284 163.367
R804 B.n282 B.n246 163.367
R805 B.n278 B.n276 163.367
R806 B.n274 B.n248 163.367
R807 B.n270 B.n268 163.367
R808 B.n266 B.n250 163.367
R809 B.n262 B.n260 163.367
R810 B.n258 B.n252 163.367
R811 B.n254 B.n190 163.367
R812 B.n476 B.n186 163.367
R813 B.n484 B.n186 163.367
R814 B.n484 B.n184 163.367
R815 B.n488 B.n184 163.367
R816 B.n488 B.n178 163.367
R817 B.n497 B.n178 163.367
R818 B.n497 B.n176 163.367
R819 B.n501 B.n176 163.367
R820 B.n501 B.n171 163.367
R821 B.n509 B.n171 163.367
R822 B.n509 B.n169 163.367
R823 B.n513 B.n169 163.367
R824 B.n513 B.n163 163.367
R825 B.n521 B.n163 163.367
R826 B.n521 B.n161 163.367
R827 B.n525 B.n161 163.367
R828 B.n525 B.n155 163.367
R829 B.n534 B.n155 163.367
R830 B.n534 B.n153 163.367
R831 B.n538 B.n153 163.367
R832 B.n538 B.n148 163.367
R833 B.n546 B.n148 163.367
R834 B.n546 B.n146 163.367
R835 B.n550 B.n146 163.367
R836 B.n550 B.n140 163.367
R837 B.n558 B.n140 163.367
R838 B.n558 B.n138 163.367
R839 B.n562 B.n138 163.367
R840 B.n562 B.n132 163.367
R841 B.n571 B.n132 163.367
R842 B.n571 B.n130 163.367
R843 B.n575 B.n130 163.367
R844 B.n575 B.n3 163.367
R845 B.n920 B.n3 163.367
R846 B.n916 B.n2 163.367
R847 B.n916 B.n915 163.367
R848 B.n915 B.n9 163.367
R849 B.n911 B.n9 163.367
R850 B.n911 B.n11 163.367
R851 B.n907 B.n11 163.367
R852 B.n907 B.n17 163.367
R853 B.n903 B.n17 163.367
R854 B.n903 B.n19 163.367
R855 B.n899 B.n19 163.367
R856 B.n899 B.n24 163.367
R857 B.n895 B.n24 163.367
R858 B.n895 B.n26 163.367
R859 B.n891 B.n26 163.367
R860 B.n891 B.n30 163.367
R861 B.n887 B.n30 163.367
R862 B.n887 B.n32 163.367
R863 B.n883 B.n32 163.367
R864 B.n883 B.n38 163.367
R865 B.n879 B.n38 163.367
R866 B.n879 B.n40 163.367
R867 B.n875 B.n40 163.367
R868 B.n875 B.n45 163.367
R869 B.n871 B.n45 163.367
R870 B.n871 B.n47 163.367
R871 B.n867 B.n47 163.367
R872 B.n867 B.n51 163.367
R873 B.n863 B.n51 163.367
R874 B.n863 B.n53 163.367
R875 B.n859 B.n53 163.367
R876 B.n859 B.n59 163.367
R877 B.n855 B.n59 163.367
R878 B.n855 B.n61 163.367
R879 B.n851 B.n61 163.367
R880 B.n846 B.n66 71.676
R881 B.n845 B.n844 71.676
R882 B.n838 B.n68 71.676
R883 B.n837 B.n836 71.676
R884 B.n830 B.n70 71.676
R885 B.n829 B.n828 71.676
R886 B.n822 B.n72 71.676
R887 B.n821 B.n820 71.676
R888 B.n814 B.n74 71.676
R889 B.n813 B.n812 71.676
R890 B.n806 B.n76 71.676
R891 B.n805 B.n804 71.676
R892 B.n798 B.n78 71.676
R893 B.n797 B.n796 71.676
R894 B.n790 B.n80 71.676
R895 B.n789 B.n788 71.676
R896 B.n782 B.n82 71.676
R897 B.n781 B.n780 71.676
R898 B.n774 B.n84 71.676
R899 B.n773 B.n772 71.676
R900 B.n766 B.n86 71.676
R901 B.n765 B.n764 71.676
R902 B.n758 B.n88 71.676
R903 B.n757 B.n756 71.676
R904 B.n750 B.n90 71.676
R905 B.n749 B.n748 71.676
R906 B.n742 B.n92 71.676
R907 B.n741 B.n740 71.676
R908 B.n734 B.n97 71.676
R909 B.n733 B.n732 71.676
R910 B.n725 B.n99 71.676
R911 B.n724 B.n723 71.676
R912 B.n717 B.n103 71.676
R913 B.n716 B.n715 71.676
R914 B.n709 B.n105 71.676
R915 B.n708 B.n707 71.676
R916 B.n701 B.n107 71.676
R917 B.n700 B.n699 71.676
R918 B.n693 B.n109 71.676
R919 B.n692 B.n691 71.676
R920 B.n685 B.n111 71.676
R921 B.n684 B.n683 71.676
R922 B.n677 B.n113 71.676
R923 B.n676 B.n675 71.676
R924 B.n669 B.n115 71.676
R925 B.n668 B.n667 71.676
R926 B.n661 B.n117 71.676
R927 B.n660 B.n659 71.676
R928 B.n653 B.n119 71.676
R929 B.n652 B.n651 71.676
R930 B.n645 B.n121 71.676
R931 B.n644 B.n643 71.676
R932 B.n637 B.n123 71.676
R933 B.n636 B.n635 71.676
R934 B.n629 B.n125 71.676
R935 B.n628 B.n627 71.676
R936 B.n627 B.n626 71.676
R937 B.n630 B.n629 71.676
R938 B.n635 B.n634 71.676
R939 B.n638 B.n637 71.676
R940 B.n643 B.n642 71.676
R941 B.n646 B.n645 71.676
R942 B.n651 B.n650 71.676
R943 B.n654 B.n653 71.676
R944 B.n659 B.n658 71.676
R945 B.n662 B.n661 71.676
R946 B.n667 B.n666 71.676
R947 B.n670 B.n669 71.676
R948 B.n675 B.n674 71.676
R949 B.n678 B.n677 71.676
R950 B.n683 B.n682 71.676
R951 B.n686 B.n685 71.676
R952 B.n691 B.n690 71.676
R953 B.n694 B.n693 71.676
R954 B.n699 B.n698 71.676
R955 B.n702 B.n701 71.676
R956 B.n707 B.n706 71.676
R957 B.n710 B.n709 71.676
R958 B.n715 B.n714 71.676
R959 B.n718 B.n717 71.676
R960 B.n723 B.n722 71.676
R961 B.n726 B.n725 71.676
R962 B.n732 B.n731 71.676
R963 B.n735 B.n734 71.676
R964 B.n740 B.n739 71.676
R965 B.n743 B.n742 71.676
R966 B.n748 B.n747 71.676
R967 B.n751 B.n750 71.676
R968 B.n756 B.n755 71.676
R969 B.n759 B.n758 71.676
R970 B.n764 B.n763 71.676
R971 B.n767 B.n766 71.676
R972 B.n772 B.n771 71.676
R973 B.n775 B.n774 71.676
R974 B.n780 B.n779 71.676
R975 B.n783 B.n782 71.676
R976 B.n788 B.n787 71.676
R977 B.n791 B.n790 71.676
R978 B.n796 B.n795 71.676
R979 B.n799 B.n798 71.676
R980 B.n804 B.n803 71.676
R981 B.n807 B.n806 71.676
R982 B.n812 B.n811 71.676
R983 B.n815 B.n814 71.676
R984 B.n820 B.n819 71.676
R985 B.n823 B.n822 71.676
R986 B.n828 B.n827 71.676
R987 B.n831 B.n830 71.676
R988 B.n836 B.n835 71.676
R989 B.n839 B.n838 71.676
R990 B.n844 B.n843 71.676
R991 B.n847 B.n846 71.676
R992 B.n471 B.n192 71.676
R993 B.n469 B.n194 71.676
R994 B.n465 B.n464 71.676
R995 B.n458 B.n196 71.676
R996 B.n457 B.n456 71.676
R997 B.n450 B.n198 71.676
R998 B.n449 B.n448 71.676
R999 B.n442 B.n200 71.676
R1000 B.n441 B.n440 71.676
R1001 B.n434 B.n202 71.676
R1002 B.n433 B.n432 71.676
R1003 B.n426 B.n204 71.676
R1004 B.n425 B.n424 71.676
R1005 B.n418 B.n206 71.676
R1006 B.n417 B.n416 71.676
R1007 B.n410 B.n208 71.676
R1008 B.n409 B.n408 71.676
R1009 B.n402 B.n210 71.676
R1010 B.n401 B.n400 71.676
R1011 B.n394 B.n212 71.676
R1012 B.n393 B.n392 71.676
R1013 B.n386 B.n214 71.676
R1014 B.n385 B.n384 71.676
R1015 B.n378 B.n216 71.676
R1016 B.n377 B.n376 71.676
R1017 B.n369 B.n218 71.676
R1018 B.n368 B.n367 71.676
R1019 B.n361 B.n222 71.676
R1020 B.n360 B.n359 71.676
R1021 B.n353 B.n224 71.676
R1022 B.n352 B.n228 71.676
R1023 B.n348 B.n347 71.676
R1024 B.n341 B.n230 71.676
R1025 B.n340 B.n339 71.676
R1026 B.n333 B.n232 71.676
R1027 B.n332 B.n331 71.676
R1028 B.n325 B.n234 71.676
R1029 B.n324 B.n323 71.676
R1030 B.n317 B.n236 71.676
R1031 B.n316 B.n315 71.676
R1032 B.n309 B.n238 71.676
R1033 B.n308 B.n307 71.676
R1034 B.n301 B.n240 71.676
R1035 B.n300 B.n299 71.676
R1036 B.n293 B.n242 71.676
R1037 B.n292 B.n291 71.676
R1038 B.n285 B.n244 71.676
R1039 B.n284 B.n283 71.676
R1040 B.n277 B.n246 71.676
R1041 B.n276 B.n275 71.676
R1042 B.n269 B.n248 71.676
R1043 B.n268 B.n267 71.676
R1044 B.n261 B.n250 71.676
R1045 B.n260 B.n259 71.676
R1046 B.n253 B.n252 71.676
R1047 B.n472 B.n471 71.676
R1048 B.n466 B.n194 71.676
R1049 B.n464 B.n463 71.676
R1050 B.n459 B.n458 71.676
R1051 B.n456 B.n455 71.676
R1052 B.n451 B.n450 71.676
R1053 B.n448 B.n447 71.676
R1054 B.n443 B.n442 71.676
R1055 B.n440 B.n439 71.676
R1056 B.n435 B.n434 71.676
R1057 B.n432 B.n431 71.676
R1058 B.n427 B.n426 71.676
R1059 B.n424 B.n423 71.676
R1060 B.n419 B.n418 71.676
R1061 B.n416 B.n415 71.676
R1062 B.n411 B.n410 71.676
R1063 B.n408 B.n407 71.676
R1064 B.n403 B.n402 71.676
R1065 B.n400 B.n399 71.676
R1066 B.n395 B.n394 71.676
R1067 B.n392 B.n391 71.676
R1068 B.n387 B.n386 71.676
R1069 B.n384 B.n383 71.676
R1070 B.n379 B.n378 71.676
R1071 B.n376 B.n375 71.676
R1072 B.n370 B.n369 71.676
R1073 B.n367 B.n366 71.676
R1074 B.n362 B.n361 71.676
R1075 B.n359 B.n358 71.676
R1076 B.n354 B.n353 71.676
R1077 B.n349 B.n228 71.676
R1078 B.n347 B.n346 71.676
R1079 B.n342 B.n341 71.676
R1080 B.n339 B.n338 71.676
R1081 B.n334 B.n333 71.676
R1082 B.n331 B.n330 71.676
R1083 B.n326 B.n325 71.676
R1084 B.n323 B.n322 71.676
R1085 B.n318 B.n317 71.676
R1086 B.n315 B.n314 71.676
R1087 B.n310 B.n309 71.676
R1088 B.n307 B.n306 71.676
R1089 B.n302 B.n301 71.676
R1090 B.n299 B.n298 71.676
R1091 B.n294 B.n293 71.676
R1092 B.n291 B.n290 71.676
R1093 B.n286 B.n285 71.676
R1094 B.n283 B.n282 71.676
R1095 B.n278 B.n277 71.676
R1096 B.n275 B.n274 71.676
R1097 B.n270 B.n269 71.676
R1098 B.n267 B.n266 71.676
R1099 B.n262 B.n261 71.676
R1100 B.n259 B.n258 71.676
R1101 B.n254 B.n253 71.676
R1102 B.n921 B.n920 71.676
R1103 B.n921 B.n2 71.676
R1104 B.n95 B.n94 59.5399
R1105 B.n728 B.n101 59.5399
R1106 B.n227 B.n226 59.5399
R1107 B.n373 B.n220 59.5399
R1108 B.n477 B.n191 59.2867
R1109 B.n852 B.n65 59.2867
R1110 B.n94 B.n93 57.6005
R1111 B.n101 B.n100 57.6005
R1112 B.n226 B.n225 57.6005
R1113 B.n220 B.n219 57.6005
R1114 B.n477 B.n187 36.32
R1115 B.n483 B.n187 36.32
R1116 B.n483 B.n183 36.32
R1117 B.n489 B.n183 36.32
R1118 B.n489 B.n179 36.32
R1119 B.n496 B.n179 36.32
R1120 B.n496 B.n495 36.32
R1121 B.n502 B.n172 36.32
R1122 B.n508 B.n172 36.32
R1123 B.n508 B.n168 36.32
R1124 B.n514 B.n168 36.32
R1125 B.n514 B.n164 36.32
R1126 B.n520 B.n164 36.32
R1127 B.n520 B.n160 36.32
R1128 B.n526 B.n160 36.32
R1129 B.n526 B.n156 36.32
R1130 B.n533 B.n156 36.32
R1131 B.n533 B.n532 36.32
R1132 B.n539 B.n149 36.32
R1133 B.n545 B.n149 36.32
R1134 B.n545 B.n145 36.32
R1135 B.n551 B.n145 36.32
R1136 B.n551 B.n141 36.32
R1137 B.n557 B.n141 36.32
R1138 B.n557 B.n137 36.32
R1139 B.n563 B.n137 36.32
R1140 B.n570 B.n133 36.32
R1141 B.n570 B.n129 36.32
R1142 B.n576 B.n129 36.32
R1143 B.n576 B.n4 36.32
R1144 B.n919 B.n4 36.32
R1145 B.n919 B.n918 36.32
R1146 B.n918 B.n917 36.32
R1147 B.n917 B.n8 36.32
R1148 B.n12 B.n8 36.32
R1149 B.n910 B.n12 36.32
R1150 B.n910 B.n909 36.32
R1151 B.n908 B.n16 36.32
R1152 B.n902 B.n16 36.32
R1153 B.n902 B.n901 36.32
R1154 B.n901 B.n900 36.32
R1155 B.n900 B.n23 36.32
R1156 B.n894 B.n23 36.32
R1157 B.n894 B.n893 36.32
R1158 B.n893 B.n892 36.32
R1159 B.n886 B.n33 36.32
R1160 B.n886 B.n885 36.32
R1161 B.n885 B.n884 36.32
R1162 B.n884 B.n37 36.32
R1163 B.n878 B.n37 36.32
R1164 B.n878 B.n877 36.32
R1165 B.n877 B.n876 36.32
R1166 B.n876 B.n44 36.32
R1167 B.n870 B.n44 36.32
R1168 B.n870 B.n869 36.32
R1169 B.n869 B.n868 36.32
R1170 B.n862 B.n54 36.32
R1171 B.n862 B.n861 36.32
R1172 B.n861 B.n860 36.32
R1173 B.n860 B.n58 36.32
R1174 B.n854 B.n58 36.32
R1175 B.n854 B.n853 36.32
R1176 B.n853 B.n852 36.32
R1177 B.n475 B.n474 32.3127
R1178 B.n479 B.n189 32.3127
R1179 B.n625 B.n624 32.3127
R1180 B.n850 B.n849 32.3127
R1181 B.n495 B.t5 30.9789
R1182 B.n54 B.t9 30.9789
R1183 B.n532 B.t2 28.8425
R1184 B.n33 B.t1 28.8425
R1185 B.n563 B.t3 19.2285
R1186 B.t0 B.n908 19.2285
R1187 B B.n922 18.0485
R1188 B.t3 B.n133 17.092
R1189 B.n909 B.t0 17.092
R1190 B.n475 B.n185 10.6151
R1191 B.n485 B.n185 10.6151
R1192 B.n486 B.n485 10.6151
R1193 B.n487 B.n486 10.6151
R1194 B.n487 B.n177 10.6151
R1195 B.n498 B.n177 10.6151
R1196 B.n499 B.n498 10.6151
R1197 B.n500 B.n499 10.6151
R1198 B.n500 B.n170 10.6151
R1199 B.n510 B.n170 10.6151
R1200 B.n511 B.n510 10.6151
R1201 B.n512 B.n511 10.6151
R1202 B.n512 B.n162 10.6151
R1203 B.n522 B.n162 10.6151
R1204 B.n523 B.n522 10.6151
R1205 B.n524 B.n523 10.6151
R1206 B.n524 B.n154 10.6151
R1207 B.n535 B.n154 10.6151
R1208 B.n536 B.n535 10.6151
R1209 B.n537 B.n536 10.6151
R1210 B.n537 B.n147 10.6151
R1211 B.n547 B.n147 10.6151
R1212 B.n548 B.n547 10.6151
R1213 B.n549 B.n548 10.6151
R1214 B.n549 B.n139 10.6151
R1215 B.n559 B.n139 10.6151
R1216 B.n560 B.n559 10.6151
R1217 B.n561 B.n560 10.6151
R1218 B.n561 B.n131 10.6151
R1219 B.n572 B.n131 10.6151
R1220 B.n573 B.n572 10.6151
R1221 B.n574 B.n573 10.6151
R1222 B.n574 B.n0 10.6151
R1223 B.n474 B.n473 10.6151
R1224 B.n473 B.n193 10.6151
R1225 B.n468 B.n193 10.6151
R1226 B.n468 B.n467 10.6151
R1227 B.n467 B.n195 10.6151
R1228 B.n462 B.n195 10.6151
R1229 B.n462 B.n461 10.6151
R1230 B.n461 B.n460 10.6151
R1231 B.n460 B.n197 10.6151
R1232 B.n454 B.n197 10.6151
R1233 B.n454 B.n453 10.6151
R1234 B.n453 B.n452 10.6151
R1235 B.n452 B.n199 10.6151
R1236 B.n446 B.n199 10.6151
R1237 B.n446 B.n445 10.6151
R1238 B.n445 B.n444 10.6151
R1239 B.n444 B.n201 10.6151
R1240 B.n438 B.n201 10.6151
R1241 B.n438 B.n437 10.6151
R1242 B.n437 B.n436 10.6151
R1243 B.n436 B.n203 10.6151
R1244 B.n430 B.n203 10.6151
R1245 B.n430 B.n429 10.6151
R1246 B.n429 B.n428 10.6151
R1247 B.n428 B.n205 10.6151
R1248 B.n422 B.n205 10.6151
R1249 B.n422 B.n421 10.6151
R1250 B.n421 B.n420 10.6151
R1251 B.n420 B.n207 10.6151
R1252 B.n414 B.n207 10.6151
R1253 B.n414 B.n413 10.6151
R1254 B.n413 B.n412 10.6151
R1255 B.n412 B.n209 10.6151
R1256 B.n406 B.n209 10.6151
R1257 B.n406 B.n405 10.6151
R1258 B.n405 B.n404 10.6151
R1259 B.n404 B.n211 10.6151
R1260 B.n398 B.n211 10.6151
R1261 B.n398 B.n397 10.6151
R1262 B.n397 B.n396 10.6151
R1263 B.n396 B.n213 10.6151
R1264 B.n390 B.n213 10.6151
R1265 B.n390 B.n389 10.6151
R1266 B.n389 B.n388 10.6151
R1267 B.n388 B.n215 10.6151
R1268 B.n382 B.n215 10.6151
R1269 B.n382 B.n381 10.6151
R1270 B.n381 B.n380 10.6151
R1271 B.n380 B.n217 10.6151
R1272 B.n374 B.n217 10.6151
R1273 B.n372 B.n371 10.6151
R1274 B.n371 B.n221 10.6151
R1275 B.n365 B.n221 10.6151
R1276 B.n365 B.n364 10.6151
R1277 B.n364 B.n363 10.6151
R1278 B.n363 B.n223 10.6151
R1279 B.n357 B.n223 10.6151
R1280 B.n357 B.n356 10.6151
R1281 B.n356 B.n355 10.6151
R1282 B.n351 B.n350 10.6151
R1283 B.n350 B.n229 10.6151
R1284 B.n345 B.n229 10.6151
R1285 B.n345 B.n344 10.6151
R1286 B.n344 B.n343 10.6151
R1287 B.n343 B.n231 10.6151
R1288 B.n337 B.n231 10.6151
R1289 B.n337 B.n336 10.6151
R1290 B.n336 B.n335 10.6151
R1291 B.n335 B.n233 10.6151
R1292 B.n329 B.n233 10.6151
R1293 B.n329 B.n328 10.6151
R1294 B.n328 B.n327 10.6151
R1295 B.n327 B.n235 10.6151
R1296 B.n321 B.n235 10.6151
R1297 B.n321 B.n320 10.6151
R1298 B.n320 B.n319 10.6151
R1299 B.n319 B.n237 10.6151
R1300 B.n313 B.n237 10.6151
R1301 B.n313 B.n312 10.6151
R1302 B.n312 B.n311 10.6151
R1303 B.n311 B.n239 10.6151
R1304 B.n305 B.n239 10.6151
R1305 B.n305 B.n304 10.6151
R1306 B.n304 B.n303 10.6151
R1307 B.n303 B.n241 10.6151
R1308 B.n297 B.n241 10.6151
R1309 B.n297 B.n296 10.6151
R1310 B.n296 B.n295 10.6151
R1311 B.n295 B.n243 10.6151
R1312 B.n289 B.n243 10.6151
R1313 B.n289 B.n288 10.6151
R1314 B.n288 B.n287 10.6151
R1315 B.n287 B.n245 10.6151
R1316 B.n281 B.n245 10.6151
R1317 B.n281 B.n280 10.6151
R1318 B.n280 B.n279 10.6151
R1319 B.n279 B.n247 10.6151
R1320 B.n273 B.n247 10.6151
R1321 B.n273 B.n272 10.6151
R1322 B.n272 B.n271 10.6151
R1323 B.n271 B.n249 10.6151
R1324 B.n265 B.n249 10.6151
R1325 B.n265 B.n264 10.6151
R1326 B.n264 B.n263 10.6151
R1327 B.n263 B.n251 10.6151
R1328 B.n257 B.n251 10.6151
R1329 B.n257 B.n256 10.6151
R1330 B.n256 B.n255 10.6151
R1331 B.n255 B.n189 10.6151
R1332 B.n480 B.n479 10.6151
R1333 B.n481 B.n480 10.6151
R1334 B.n481 B.n181 10.6151
R1335 B.n491 B.n181 10.6151
R1336 B.n492 B.n491 10.6151
R1337 B.n493 B.n492 10.6151
R1338 B.n493 B.n174 10.6151
R1339 B.n504 B.n174 10.6151
R1340 B.n505 B.n504 10.6151
R1341 B.n506 B.n505 10.6151
R1342 B.n506 B.n166 10.6151
R1343 B.n516 B.n166 10.6151
R1344 B.n517 B.n516 10.6151
R1345 B.n518 B.n517 10.6151
R1346 B.n518 B.n158 10.6151
R1347 B.n528 B.n158 10.6151
R1348 B.n529 B.n528 10.6151
R1349 B.n530 B.n529 10.6151
R1350 B.n530 B.n151 10.6151
R1351 B.n541 B.n151 10.6151
R1352 B.n542 B.n541 10.6151
R1353 B.n543 B.n542 10.6151
R1354 B.n543 B.n143 10.6151
R1355 B.n553 B.n143 10.6151
R1356 B.n554 B.n553 10.6151
R1357 B.n555 B.n554 10.6151
R1358 B.n555 B.n135 10.6151
R1359 B.n565 B.n135 10.6151
R1360 B.n566 B.n565 10.6151
R1361 B.n568 B.n566 10.6151
R1362 B.n568 B.n567 10.6151
R1363 B.n567 B.n127 10.6151
R1364 B.n579 B.n127 10.6151
R1365 B.n580 B.n579 10.6151
R1366 B.n581 B.n580 10.6151
R1367 B.n582 B.n581 10.6151
R1368 B.n583 B.n582 10.6151
R1369 B.n586 B.n583 10.6151
R1370 B.n587 B.n586 10.6151
R1371 B.n588 B.n587 10.6151
R1372 B.n589 B.n588 10.6151
R1373 B.n591 B.n589 10.6151
R1374 B.n592 B.n591 10.6151
R1375 B.n593 B.n592 10.6151
R1376 B.n594 B.n593 10.6151
R1377 B.n596 B.n594 10.6151
R1378 B.n597 B.n596 10.6151
R1379 B.n598 B.n597 10.6151
R1380 B.n599 B.n598 10.6151
R1381 B.n601 B.n599 10.6151
R1382 B.n602 B.n601 10.6151
R1383 B.n603 B.n602 10.6151
R1384 B.n604 B.n603 10.6151
R1385 B.n606 B.n604 10.6151
R1386 B.n607 B.n606 10.6151
R1387 B.n608 B.n607 10.6151
R1388 B.n609 B.n608 10.6151
R1389 B.n611 B.n609 10.6151
R1390 B.n612 B.n611 10.6151
R1391 B.n613 B.n612 10.6151
R1392 B.n614 B.n613 10.6151
R1393 B.n616 B.n614 10.6151
R1394 B.n617 B.n616 10.6151
R1395 B.n618 B.n617 10.6151
R1396 B.n619 B.n618 10.6151
R1397 B.n621 B.n619 10.6151
R1398 B.n622 B.n621 10.6151
R1399 B.n623 B.n622 10.6151
R1400 B.n624 B.n623 10.6151
R1401 B.n914 B.n1 10.6151
R1402 B.n914 B.n913 10.6151
R1403 B.n913 B.n912 10.6151
R1404 B.n912 B.n10 10.6151
R1405 B.n906 B.n10 10.6151
R1406 B.n906 B.n905 10.6151
R1407 B.n905 B.n904 10.6151
R1408 B.n904 B.n18 10.6151
R1409 B.n898 B.n18 10.6151
R1410 B.n898 B.n897 10.6151
R1411 B.n897 B.n896 10.6151
R1412 B.n896 B.n25 10.6151
R1413 B.n890 B.n25 10.6151
R1414 B.n890 B.n889 10.6151
R1415 B.n889 B.n888 10.6151
R1416 B.n888 B.n31 10.6151
R1417 B.n882 B.n31 10.6151
R1418 B.n882 B.n881 10.6151
R1419 B.n881 B.n880 10.6151
R1420 B.n880 B.n39 10.6151
R1421 B.n874 B.n39 10.6151
R1422 B.n874 B.n873 10.6151
R1423 B.n873 B.n872 10.6151
R1424 B.n872 B.n46 10.6151
R1425 B.n866 B.n46 10.6151
R1426 B.n866 B.n865 10.6151
R1427 B.n865 B.n864 10.6151
R1428 B.n864 B.n52 10.6151
R1429 B.n858 B.n52 10.6151
R1430 B.n858 B.n857 10.6151
R1431 B.n857 B.n856 10.6151
R1432 B.n856 B.n60 10.6151
R1433 B.n850 B.n60 10.6151
R1434 B.n849 B.n848 10.6151
R1435 B.n848 B.n67 10.6151
R1436 B.n842 B.n67 10.6151
R1437 B.n842 B.n841 10.6151
R1438 B.n841 B.n840 10.6151
R1439 B.n840 B.n69 10.6151
R1440 B.n834 B.n69 10.6151
R1441 B.n834 B.n833 10.6151
R1442 B.n833 B.n832 10.6151
R1443 B.n832 B.n71 10.6151
R1444 B.n826 B.n71 10.6151
R1445 B.n826 B.n825 10.6151
R1446 B.n825 B.n824 10.6151
R1447 B.n824 B.n73 10.6151
R1448 B.n818 B.n73 10.6151
R1449 B.n818 B.n817 10.6151
R1450 B.n817 B.n816 10.6151
R1451 B.n816 B.n75 10.6151
R1452 B.n810 B.n75 10.6151
R1453 B.n810 B.n809 10.6151
R1454 B.n809 B.n808 10.6151
R1455 B.n808 B.n77 10.6151
R1456 B.n802 B.n77 10.6151
R1457 B.n802 B.n801 10.6151
R1458 B.n801 B.n800 10.6151
R1459 B.n800 B.n79 10.6151
R1460 B.n794 B.n79 10.6151
R1461 B.n794 B.n793 10.6151
R1462 B.n793 B.n792 10.6151
R1463 B.n792 B.n81 10.6151
R1464 B.n786 B.n81 10.6151
R1465 B.n786 B.n785 10.6151
R1466 B.n785 B.n784 10.6151
R1467 B.n784 B.n83 10.6151
R1468 B.n778 B.n83 10.6151
R1469 B.n778 B.n777 10.6151
R1470 B.n777 B.n776 10.6151
R1471 B.n776 B.n85 10.6151
R1472 B.n770 B.n85 10.6151
R1473 B.n770 B.n769 10.6151
R1474 B.n769 B.n768 10.6151
R1475 B.n768 B.n87 10.6151
R1476 B.n762 B.n87 10.6151
R1477 B.n762 B.n761 10.6151
R1478 B.n761 B.n760 10.6151
R1479 B.n760 B.n89 10.6151
R1480 B.n754 B.n89 10.6151
R1481 B.n754 B.n753 10.6151
R1482 B.n753 B.n752 10.6151
R1483 B.n752 B.n91 10.6151
R1484 B.n746 B.n745 10.6151
R1485 B.n745 B.n744 10.6151
R1486 B.n744 B.n96 10.6151
R1487 B.n738 B.n96 10.6151
R1488 B.n738 B.n737 10.6151
R1489 B.n737 B.n736 10.6151
R1490 B.n736 B.n98 10.6151
R1491 B.n730 B.n98 10.6151
R1492 B.n730 B.n729 10.6151
R1493 B.n727 B.n102 10.6151
R1494 B.n721 B.n102 10.6151
R1495 B.n721 B.n720 10.6151
R1496 B.n720 B.n719 10.6151
R1497 B.n719 B.n104 10.6151
R1498 B.n713 B.n104 10.6151
R1499 B.n713 B.n712 10.6151
R1500 B.n712 B.n711 10.6151
R1501 B.n711 B.n106 10.6151
R1502 B.n705 B.n106 10.6151
R1503 B.n705 B.n704 10.6151
R1504 B.n704 B.n703 10.6151
R1505 B.n703 B.n108 10.6151
R1506 B.n697 B.n108 10.6151
R1507 B.n697 B.n696 10.6151
R1508 B.n696 B.n695 10.6151
R1509 B.n695 B.n110 10.6151
R1510 B.n689 B.n110 10.6151
R1511 B.n689 B.n688 10.6151
R1512 B.n688 B.n687 10.6151
R1513 B.n687 B.n112 10.6151
R1514 B.n681 B.n112 10.6151
R1515 B.n681 B.n680 10.6151
R1516 B.n680 B.n679 10.6151
R1517 B.n679 B.n114 10.6151
R1518 B.n673 B.n114 10.6151
R1519 B.n673 B.n672 10.6151
R1520 B.n672 B.n671 10.6151
R1521 B.n671 B.n116 10.6151
R1522 B.n665 B.n116 10.6151
R1523 B.n665 B.n664 10.6151
R1524 B.n664 B.n663 10.6151
R1525 B.n663 B.n118 10.6151
R1526 B.n657 B.n118 10.6151
R1527 B.n657 B.n656 10.6151
R1528 B.n656 B.n655 10.6151
R1529 B.n655 B.n120 10.6151
R1530 B.n649 B.n120 10.6151
R1531 B.n649 B.n648 10.6151
R1532 B.n648 B.n647 10.6151
R1533 B.n647 B.n122 10.6151
R1534 B.n641 B.n122 10.6151
R1535 B.n641 B.n640 10.6151
R1536 B.n640 B.n639 10.6151
R1537 B.n639 B.n124 10.6151
R1538 B.n633 B.n124 10.6151
R1539 B.n633 B.n632 10.6151
R1540 B.n632 B.n631 10.6151
R1541 B.n631 B.n126 10.6151
R1542 B.n625 B.n126 10.6151
R1543 B.n374 B.n373 9.36635
R1544 B.n351 B.n227 9.36635
R1545 B.n95 B.n91 9.36635
R1546 B.n728 B.n727 9.36635
R1547 B.n922 B.n0 8.11757
R1548 B.n922 B.n1 8.11757
R1549 B.n539 B.t2 7.47804
R1550 B.n892 B.t1 7.47804
R1551 B.n502 B.t5 5.3416
R1552 B.n868 B.t9 5.3416
R1553 B.n373 B.n372 1.24928
R1554 B.n355 B.n227 1.24928
R1555 B.n746 B.n95 1.24928
R1556 B.n729 B.n728 1.24928
R1557 VP.n4 VP.t2 176.411
R1558 VP.n4 VP.t3 175.627
R1559 VP.n14 VP.n0 161.3
R1560 VP.n13 VP.n12 161.3
R1561 VP.n11 VP.n1 161.3
R1562 VP.n10 VP.n9 161.3
R1563 VP.n8 VP.n2 161.3
R1564 VP.n7 VP.n6 161.3
R1565 VP.n3 VP.t0 139.853
R1566 VP.n15 VP.t1 139.853
R1567 VP.n5 VP.n3 99.3501
R1568 VP.n16 VP.n15 99.3501
R1569 VP.n9 VP.n1 56.5617
R1570 VP.n5 VP.n4 53.2378
R1571 VP.n8 VP.n7 24.5923
R1572 VP.n9 VP.n8 24.5923
R1573 VP.n13 VP.n1 24.5923
R1574 VP.n14 VP.n13 24.5923
R1575 VP.n7 VP.n3 11.5587
R1576 VP.n15 VP.n14 11.5587
R1577 VP.n6 VP.n5 0.278335
R1578 VP.n16 VP.n0 0.278335
R1579 VP.n6 VP.n2 0.189894
R1580 VP.n10 VP.n2 0.189894
R1581 VP.n11 VP.n10 0.189894
R1582 VP.n12 VP.n11 0.189894
R1583 VP.n12 VP.n0 0.189894
R1584 VP VP.n16 0.153485
R1585 VDD1 VDD1.n1 105.195
R1586 VDD1 VDD1.n0 60.1248
R1587 VDD1.n0 VDD1.t2 1.29293
R1588 VDD1.n0 VDD1.t1 1.29293
R1589 VDD1.n1 VDD1.t3 1.29293
R1590 VDD1.n1 VDD1.t0 1.29293
R1591 VTAIL.n682 VTAIL.n602 289.615
R1592 VTAIL.n80 VTAIL.n0 289.615
R1593 VTAIL.n166 VTAIL.n86 289.615
R1594 VTAIL.n252 VTAIL.n172 289.615
R1595 VTAIL.n596 VTAIL.n516 289.615
R1596 VTAIL.n510 VTAIL.n430 289.615
R1597 VTAIL.n424 VTAIL.n344 289.615
R1598 VTAIL.n338 VTAIL.n258 289.615
R1599 VTAIL.n631 VTAIL.n630 185
R1600 VTAIL.n633 VTAIL.n632 185
R1601 VTAIL.n626 VTAIL.n625 185
R1602 VTAIL.n639 VTAIL.n638 185
R1603 VTAIL.n641 VTAIL.n640 185
R1604 VTAIL.n622 VTAIL.n621 185
R1605 VTAIL.n647 VTAIL.n646 185
R1606 VTAIL.n649 VTAIL.n648 185
R1607 VTAIL.n618 VTAIL.n617 185
R1608 VTAIL.n655 VTAIL.n654 185
R1609 VTAIL.n657 VTAIL.n656 185
R1610 VTAIL.n614 VTAIL.n613 185
R1611 VTAIL.n663 VTAIL.n662 185
R1612 VTAIL.n665 VTAIL.n664 185
R1613 VTAIL.n610 VTAIL.n609 185
R1614 VTAIL.n672 VTAIL.n671 185
R1615 VTAIL.n673 VTAIL.n608 185
R1616 VTAIL.n675 VTAIL.n674 185
R1617 VTAIL.n606 VTAIL.n605 185
R1618 VTAIL.n681 VTAIL.n680 185
R1619 VTAIL.n683 VTAIL.n682 185
R1620 VTAIL.n29 VTAIL.n28 185
R1621 VTAIL.n31 VTAIL.n30 185
R1622 VTAIL.n24 VTAIL.n23 185
R1623 VTAIL.n37 VTAIL.n36 185
R1624 VTAIL.n39 VTAIL.n38 185
R1625 VTAIL.n20 VTAIL.n19 185
R1626 VTAIL.n45 VTAIL.n44 185
R1627 VTAIL.n47 VTAIL.n46 185
R1628 VTAIL.n16 VTAIL.n15 185
R1629 VTAIL.n53 VTAIL.n52 185
R1630 VTAIL.n55 VTAIL.n54 185
R1631 VTAIL.n12 VTAIL.n11 185
R1632 VTAIL.n61 VTAIL.n60 185
R1633 VTAIL.n63 VTAIL.n62 185
R1634 VTAIL.n8 VTAIL.n7 185
R1635 VTAIL.n70 VTAIL.n69 185
R1636 VTAIL.n71 VTAIL.n6 185
R1637 VTAIL.n73 VTAIL.n72 185
R1638 VTAIL.n4 VTAIL.n3 185
R1639 VTAIL.n79 VTAIL.n78 185
R1640 VTAIL.n81 VTAIL.n80 185
R1641 VTAIL.n115 VTAIL.n114 185
R1642 VTAIL.n117 VTAIL.n116 185
R1643 VTAIL.n110 VTAIL.n109 185
R1644 VTAIL.n123 VTAIL.n122 185
R1645 VTAIL.n125 VTAIL.n124 185
R1646 VTAIL.n106 VTAIL.n105 185
R1647 VTAIL.n131 VTAIL.n130 185
R1648 VTAIL.n133 VTAIL.n132 185
R1649 VTAIL.n102 VTAIL.n101 185
R1650 VTAIL.n139 VTAIL.n138 185
R1651 VTAIL.n141 VTAIL.n140 185
R1652 VTAIL.n98 VTAIL.n97 185
R1653 VTAIL.n147 VTAIL.n146 185
R1654 VTAIL.n149 VTAIL.n148 185
R1655 VTAIL.n94 VTAIL.n93 185
R1656 VTAIL.n156 VTAIL.n155 185
R1657 VTAIL.n157 VTAIL.n92 185
R1658 VTAIL.n159 VTAIL.n158 185
R1659 VTAIL.n90 VTAIL.n89 185
R1660 VTAIL.n165 VTAIL.n164 185
R1661 VTAIL.n167 VTAIL.n166 185
R1662 VTAIL.n201 VTAIL.n200 185
R1663 VTAIL.n203 VTAIL.n202 185
R1664 VTAIL.n196 VTAIL.n195 185
R1665 VTAIL.n209 VTAIL.n208 185
R1666 VTAIL.n211 VTAIL.n210 185
R1667 VTAIL.n192 VTAIL.n191 185
R1668 VTAIL.n217 VTAIL.n216 185
R1669 VTAIL.n219 VTAIL.n218 185
R1670 VTAIL.n188 VTAIL.n187 185
R1671 VTAIL.n225 VTAIL.n224 185
R1672 VTAIL.n227 VTAIL.n226 185
R1673 VTAIL.n184 VTAIL.n183 185
R1674 VTAIL.n233 VTAIL.n232 185
R1675 VTAIL.n235 VTAIL.n234 185
R1676 VTAIL.n180 VTAIL.n179 185
R1677 VTAIL.n242 VTAIL.n241 185
R1678 VTAIL.n243 VTAIL.n178 185
R1679 VTAIL.n245 VTAIL.n244 185
R1680 VTAIL.n176 VTAIL.n175 185
R1681 VTAIL.n251 VTAIL.n250 185
R1682 VTAIL.n253 VTAIL.n252 185
R1683 VTAIL.n597 VTAIL.n596 185
R1684 VTAIL.n595 VTAIL.n594 185
R1685 VTAIL.n520 VTAIL.n519 185
R1686 VTAIL.n524 VTAIL.n522 185
R1687 VTAIL.n589 VTAIL.n588 185
R1688 VTAIL.n587 VTAIL.n586 185
R1689 VTAIL.n526 VTAIL.n525 185
R1690 VTAIL.n581 VTAIL.n580 185
R1691 VTAIL.n579 VTAIL.n578 185
R1692 VTAIL.n530 VTAIL.n529 185
R1693 VTAIL.n573 VTAIL.n572 185
R1694 VTAIL.n571 VTAIL.n570 185
R1695 VTAIL.n534 VTAIL.n533 185
R1696 VTAIL.n565 VTAIL.n564 185
R1697 VTAIL.n563 VTAIL.n562 185
R1698 VTAIL.n538 VTAIL.n537 185
R1699 VTAIL.n557 VTAIL.n556 185
R1700 VTAIL.n555 VTAIL.n554 185
R1701 VTAIL.n542 VTAIL.n541 185
R1702 VTAIL.n549 VTAIL.n548 185
R1703 VTAIL.n547 VTAIL.n546 185
R1704 VTAIL.n511 VTAIL.n510 185
R1705 VTAIL.n509 VTAIL.n508 185
R1706 VTAIL.n434 VTAIL.n433 185
R1707 VTAIL.n438 VTAIL.n436 185
R1708 VTAIL.n503 VTAIL.n502 185
R1709 VTAIL.n501 VTAIL.n500 185
R1710 VTAIL.n440 VTAIL.n439 185
R1711 VTAIL.n495 VTAIL.n494 185
R1712 VTAIL.n493 VTAIL.n492 185
R1713 VTAIL.n444 VTAIL.n443 185
R1714 VTAIL.n487 VTAIL.n486 185
R1715 VTAIL.n485 VTAIL.n484 185
R1716 VTAIL.n448 VTAIL.n447 185
R1717 VTAIL.n479 VTAIL.n478 185
R1718 VTAIL.n477 VTAIL.n476 185
R1719 VTAIL.n452 VTAIL.n451 185
R1720 VTAIL.n471 VTAIL.n470 185
R1721 VTAIL.n469 VTAIL.n468 185
R1722 VTAIL.n456 VTAIL.n455 185
R1723 VTAIL.n463 VTAIL.n462 185
R1724 VTAIL.n461 VTAIL.n460 185
R1725 VTAIL.n425 VTAIL.n424 185
R1726 VTAIL.n423 VTAIL.n422 185
R1727 VTAIL.n348 VTAIL.n347 185
R1728 VTAIL.n352 VTAIL.n350 185
R1729 VTAIL.n417 VTAIL.n416 185
R1730 VTAIL.n415 VTAIL.n414 185
R1731 VTAIL.n354 VTAIL.n353 185
R1732 VTAIL.n409 VTAIL.n408 185
R1733 VTAIL.n407 VTAIL.n406 185
R1734 VTAIL.n358 VTAIL.n357 185
R1735 VTAIL.n401 VTAIL.n400 185
R1736 VTAIL.n399 VTAIL.n398 185
R1737 VTAIL.n362 VTAIL.n361 185
R1738 VTAIL.n393 VTAIL.n392 185
R1739 VTAIL.n391 VTAIL.n390 185
R1740 VTAIL.n366 VTAIL.n365 185
R1741 VTAIL.n385 VTAIL.n384 185
R1742 VTAIL.n383 VTAIL.n382 185
R1743 VTAIL.n370 VTAIL.n369 185
R1744 VTAIL.n377 VTAIL.n376 185
R1745 VTAIL.n375 VTAIL.n374 185
R1746 VTAIL.n339 VTAIL.n338 185
R1747 VTAIL.n337 VTAIL.n336 185
R1748 VTAIL.n262 VTAIL.n261 185
R1749 VTAIL.n266 VTAIL.n264 185
R1750 VTAIL.n331 VTAIL.n330 185
R1751 VTAIL.n329 VTAIL.n328 185
R1752 VTAIL.n268 VTAIL.n267 185
R1753 VTAIL.n323 VTAIL.n322 185
R1754 VTAIL.n321 VTAIL.n320 185
R1755 VTAIL.n272 VTAIL.n271 185
R1756 VTAIL.n315 VTAIL.n314 185
R1757 VTAIL.n313 VTAIL.n312 185
R1758 VTAIL.n276 VTAIL.n275 185
R1759 VTAIL.n307 VTAIL.n306 185
R1760 VTAIL.n305 VTAIL.n304 185
R1761 VTAIL.n280 VTAIL.n279 185
R1762 VTAIL.n299 VTAIL.n298 185
R1763 VTAIL.n297 VTAIL.n296 185
R1764 VTAIL.n284 VTAIL.n283 185
R1765 VTAIL.n291 VTAIL.n290 185
R1766 VTAIL.n289 VTAIL.n288 185
R1767 VTAIL.n629 VTAIL.t1 147.659
R1768 VTAIL.n27 VTAIL.t0 147.659
R1769 VTAIL.n113 VTAIL.t6 147.659
R1770 VTAIL.n199 VTAIL.t7 147.659
R1771 VTAIL.n545 VTAIL.t4 147.659
R1772 VTAIL.n459 VTAIL.t5 147.659
R1773 VTAIL.n373 VTAIL.t3 147.659
R1774 VTAIL.n287 VTAIL.t2 147.659
R1775 VTAIL.n632 VTAIL.n631 104.615
R1776 VTAIL.n632 VTAIL.n625 104.615
R1777 VTAIL.n639 VTAIL.n625 104.615
R1778 VTAIL.n640 VTAIL.n639 104.615
R1779 VTAIL.n640 VTAIL.n621 104.615
R1780 VTAIL.n647 VTAIL.n621 104.615
R1781 VTAIL.n648 VTAIL.n647 104.615
R1782 VTAIL.n648 VTAIL.n617 104.615
R1783 VTAIL.n655 VTAIL.n617 104.615
R1784 VTAIL.n656 VTAIL.n655 104.615
R1785 VTAIL.n656 VTAIL.n613 104.615
R1786 VTAIL.n663 VTAIL.n613 104.615
R1787 VTAIL.n664 VTAIL.n663 104.615
R1788 VTAIL.n664 VTAIL.n609 104.615
R1789 VTAIL.n672 VTAIL.n609 104.615
R1790 VTAIL.n673 VTAIL.n672 104.615
R1791 VTAIL.n674 VTAIL.n673 104.615
R1792 VTAIL.n674 VTAIL.n605 104.615
R1793 VTAIL.n681 VTAIL.n605 104.615
R1794 VTAIL.n682 VTAIL.n681 104.615
R1795 VTAIL.n30 VTAIL.n29 104.615
R1796 VTAIL.n30 VTAIL.n23 104.615
R1797 VTAIL.n37 VTAIL.n23 104.615
R1798 VTAIL.n38 VTAIL.n37 104.615
R1799 VTAIL.n38 VTAIL.n19 104.615
R1800 VTAIL.n45 VTAIL.n19 104.615
R1801 VTAIL.n46 VTAIL.n45 104.615
R1802 VTAIL.n46 VTAIL.n15 104.615
R1803 VTAIL.n53 VTAIL.n15 104.615
R1804 VTAIL.n54 VTAIL.n53 104.615
R1805 VTAIL.n54 VTAIL.n11 104.615
R1806 VTAIL.n61 VTAIL.n11 104.615
R1807 VTAIL.n62 VTAIL.n61 104.615
R1808 VTAIL.n62 VTAIL.n7 104.615
R1809 VTAIL.n70 VTAIL.n7 104.615
R1810 VTAIL.n71 VTAIL.n70 104.615
R1811 VTAIL.n72 VTAIL.n71 104.615
R1812 VTAIL.n72 VTAIL.n3 104.615
R1813 VTAIL.n79 VTAIL.n3 104.615
R1814 VTAIL.n80 VTAIL.n79 104.615
R1815 VTAIL.n116 VTAIL.n115 104.615
R1816 VTAIL.n116 VTAIL.n109 104.615
R1817 VTAIL.n123 VTAIL.n109 104.615
R1818 VTAIL.n124 VTAIL.n123 104.615
R1819 VTAIL.n124 VTAIL.n105 104.615
R1820 VTAIL.n131 VTAIL.n105 104.615
R1821 VTAIL.n132 VTAIL.n131 104.615
R1822 VTAIL.n132 VTAIL.n101 104.615
R1823 VTAIL.n139 VTAIL.n101 104.615
R1824 VTAIL.n140 VTAIL.n139 104.615
R1825 VTAIL.n140 VTAIL.n97 104.615
R1826 VTAIL.n147 VTAIL.n97 104.615
R1827 VTAIL.n148 VTAIL.n147 104.615
R1828 VTAIL.n148 VTAIL.n93 104.615
R1829 VTAIL.n156 VTAIL.n93 104.615
R1830 VTAIL.n157 VTAIL.n156 104.615
R1831 VTAIL.n158 VTAIL.n157 104.615
R1832 VTAIL.n158 VTAIL.n89 104.615
R1833 VTAIL.n165 VTAIL.n89 104.615
R1834 VTAIL.n166 VTAIL.n165 104.615
R1835 VTAIL.n202 VTAIL.n201 104.615
R1836 VTAIL.n202 VTAIL.n195 104.615
R1837 VTAIL.n209 VTAIL.n195 104.615
R1838 VTAIL.n210 VTAIL.n209 104.615
R1839 VTAIL.n210 VTAIL.n191 104.615
R1840 VTAIL.n217 VTAIL.n191 104.615
R1841 VTAIL.n218 VTAIL.n217 104.615
R1842 VTAIL.n218 VTAIL.n187 104.615
R1843 VTAIL.n225 VTAIL.n187 104.615
R1844 VTAIL.n226 VTAIL.n225 104.615
R1845 VTAIL.n226 VTAIL.n183 104.615
R1846 VTAIL.n233 VTAIL.n183 104.615
R1847 VTAIL.n234 VTAIL.n233 104.615
R1848 VTAIL.n234 VTAIL.n179 104.615
R1849 VTAIL.n242 VTAIL.n179 104.615
R1850 VTAIL.n243 VTAIL.n242 104.615
R1851 VTAIL.n244 VTAIL.n243 104.615
R1852 VTAIL.n244 VTAIL.n175 104.615
R1853 VTAIL.n251 VTAIL.n175 104.615
R1854 VTAIL.n252 VTAIL.n251 104.615
R1855 VTAIL.n596 VTAIL.n595 104.615
R1856 VTAIL.n595 VTAIL.n519 104.615
R1857 VTAIL.n524 VTAIL.n519 104.615
R1858 VTAIL.n588 VTAIL.n524 104.615
R1859 VTAIL.n588 VTAIL.n587 104.615
R1860 VTAIL.n587 VTAIL.n525 104.615
R1861 VTAIL.n580 VTAIL.n525 104.615
R1862 VTAIL.n580 VTAIL.n579 104.615
R1863 VTAIL.n579 VTAIL.n529 104.615
R1864 VTAIL.n572 VTAIL.n529 104.615
R1865 VTAIL.n572 VTAIL.n571 104.615
R1866 VTAIL.n571 VTAIL.n533 104.615
R1867 VTAIL.n564 VTAIL.n533 104.615
R1868 VTAIL.n564 VTAIL.n563 104.615
R1869 VTAIL.n563 VTAIL.n537 104.615
R1870 VTAIL.n556 VTAIL.n537 104.615
R1871 VTAIL.n556 VTAIL.n555 104.615
R1872 VTAIL.n555 VTAIL.n541 104.615
R1873 VTAIL.n548 VTAIL.n541 104.615
R1874 VTAIL.n548 VTAIL.n547 104.615
R1875 VTAIL.n510 VTAIL.n509 104.615
R1876 VTAIL.n509 VTAIL.n433 104.615
R1877 VTAIL.n438 VTAIL.n433 104.615
R1878 VTAIL.n502 VTAIL.n438 104.615
R1879 VTAIL.n502 VTAIL.n501 104.615
R1880 VTAIL.n501 VTAIL.n439 104.615
R1881 VTAIL.n494 VTAIL.n439 104.615
R1882 VTAIL.n494 VTAIL.n493 104.615
R1883 VTAIL.n493 VTAIL.n443 104.615
R1884 VTAIL.n486 VTAIL.n443 104.615
R1885 VTAIL.n486 VTAIL.n485 104.615
R1886 VTAIL.n485 VTAIL.n447 104.615
R1887 VTAIL.n478 VTAIL.n447 104.615
R1888 VTAIL.n478 VTAIL.n477 104.615
R1889 VTAIL.n477 VTAIL.n451 104.615
R1890 VTAIL.n470 VTAIL.n451 104.615
R1891 VTAIL.n470 VTAIL.n469 104.615
R1892 VTAIL.n469 VTAIL.n455 104.615
R1893 VTAIL.n462 VTAIL.n455 104.615
R1894 VTAIL.n462 VTAIL.n461 104.615
R1895 VTAIL.n424 VTAIL.n423 104.615
R1896 VTAIL.n423 VTAIL.n347 104.615
R1897 VTAIL.n352 VTAIL.n347 104.615
R1898 VTAIL.n416 VTAIL.n352 104.615
R1899 VTAIL.n416 VTAIL.n415 104.615
R1900 VTAIL.n415 VTAIL.n353 104.615
R1901 VTAIL.n408 VTAIL.n353 104.615
R1902 VTAIL.n408 VTAIL.n407 104.615
R1903 VTAIL.n407 VTAIL.n357 104.615
R1904 VTAIL.n400 VTAIL.n357 104.615
R1905 VTAIL.n400 VTAIL.n399 104.615
R1906 VTAIL.n399 VTAIL.n361 104.615
R1907 VTAIL.n392 VTAIL.n361 104.615
R1908 VTAIL.n392 VTAIL.n391 104.615
R1909 VTAIL.n391 VTAIL.n365 104.615
R1910 VTAIL.n384 VTAIL.n365 104.615
R1911 VTAIL.n384 VTAIL.n383 104.615
R1912 VTAIL.n383 VTAIL.n369 104.615
R1913 VTAIL.n376 VTAIL.n369 104.615
R1914 VTAIL.n376 VTAIL.n375 104.615
R1915 VTAIL.n338 VTAIL.n337 104.615
R1916 VTAIL.n337 VTAIL.n261 104.615
R1917 VTAIL.n266 VTAIL.n261 104.615
R1918 VTAIL.n330 VTAIL.n266 104.615
R1919 VTAIL.n330 VTAIL.n329 104.615
R1920 VTAIL.n329 VTAIL.n267 104.615
R1921 VTAIL.n322 VTAIL.n267 104.615
R1922 VTAIL.n322 VTAIL.n321 104.615
R1923 VTAIL.n321 VTAIL.n271 104.615
R1924 VTAIL.n314 VTAIL.n271 104.615
R1925 VTAIL.n314 VTAIL.n313 104.615
R1926 VTAIL.n313 VTAIL.n275 104.615
R1927 VTAIL.n306 VTAIL.n275 104.615
R1928 VTAIL.n306 VTAIL.n305 104.615
R1929 VTAIL.n305 VTAIL.n279 104.615
R1930 VTAIL.n298 VTAIL.n279 104.615
R1931 VTAIL.n298 VTAIL.n297 104.615
R1932 VTAIL.n297 VTAIL.n283 104.615
R1933 VTAIL.n290 VTAIL.n283 104.615
R1934 VTAIL.n290 VTAIL.n289 104.615
R1935 VTAIL.n631 VTAIL.t1 52.3082
R1936 VTAIL.n29 VTAIL.t0 52.3082
R1937 VTAIL.n115 VTAIL.t6 52.3082
R1938 VTAIL.n201 VTAIL.t7 52.3082
R1939 VTAIL.n547 VTAIL.t4 52.3082
R1940 VTAIL.n461 VTAIL.t5 52.3082
R1941 VTAIL.n375 VTAIL.t3 52.3082
R1942 VTAIL.n289 VTAIL.t2 52.3082
R1943 VTAIL.n687 VTAIL.n686 31.4096
R1944 VTAIL.n85 VTAIL.n84 31.4096
R1945 VTAIL.n171 VTAIL.n170 31.4096
R1946 VTAIL.n257 VTAIL.n256 31.4096
R1947 VTAIL.n601 VTAIL.n600 31.4096
R1948 VTAIL.n515 VTAIL.n514 31.4096
R1949 VTAIL.n429 VTAIL.n428 31.4096
R1950 VTAIL.n343 VTAIL.n342 31.4096
R1951 VTAIL.n687 VTAIL.n601 28.1341
R1952 VTAIL.n343 VTAIL.n257 28.1341
R1953 VTAIL.n630 VTAIL.n629 15.6677
R1954 VTAIL.n28 VTAIL.n27 15.6677
R1955 VTAIL.n114 VTAIL.n113 15.6677
R1956 VTAIL.n200 VTAIL.n199 15.6677
R1957 VTAIL.n546 VTAIL.n545 15.6677
R1958 VTAIL.n460 VTAIL.n459 15.6677
R1959 VTAIL.n374 VTAIL.n373 15.6677
R1960 VTAIL.n288 VTAIL.n287 15.6677
R1961 VTAIL.n675 VTAIL.n606 13.1884
R1962 VTAIL.n73 VTAIL.n4 13.1884
R1963 VTAIL.n159 VTAIL.n90 13.1884
R1964 VTAIL.n245 VTAIL.n176 13.1884
R1965 VTAIL.n522 VTAIL.n520 13.1884
R1966 VTAIL.n436 VTAIL.n434 13.1884
R1967 VTAIL.n350 VTAIL.n348 13.1884
R1968 VTAIL.n264 VTAIL.n262 13.1884
R1969 VTAIL.n633 VTAIL.n628 12.8005
R1970 VTAIL.n676 VTAIL.n608 12.8005
R1971 VTAIL.n680 VTAIL.n679 12.8005
R1972 VTAIL.n31 VTAIL.n26 12.8005
R1973 VTAIL.n74 VTAIL.n6 12.8005
R1974 VTAIL.n78 VTAIL.n77 12.8005
R1975 VTAIL.n117 VTAIL.n112 12.8005
R1976 VTAIL.n160 VTAIL.n92 12.8005
R1977 VTAIL.n164 VTAIL.n163 12.8005
R1978 VTAIL.n203 VTAIL.n198 12.8005
R1979 VTAIL.n246 VTAIL.n178 12.8005
R1980 VTAIL.n250 VTAIL.n249 12.8005
R1981 VTAIL.n594 VTAIL.n593 12.8005
R1982 VTAIL.n590 VTAIL.n589 12.8005
R1983 VTAIL.n549 VTAIL.n544 12.8005
R1984 VTAIL.n508 VTAIL.n507 12.8005
R1985 VTAIL.n504 VTAIL.n503 12.8005
R1986 VTAIL.n463 VTAIL.n458 12.8005
R1987 VTAIL.n422 VTAIL.n421 12.8005
R1988 VTAIL.n418 VTAIL.n417 12.8005
R1989 VTAIL.n377 VTAIL.n372 12.8005
R1990 VTAIL.n336 VTAIL.n335 12.8005
R1991 VTAIL.n332 VTAIL.n331 12.8005
R1992 VTAIL.n291 VTAIL.n286 12.8005
R1993 VTAIL.n634 VTAIL.n626 12.0247
R1994 VTAIL.n671 VTAIL.n670 12.0247
R1995 VTAIL.n683 VTAIL.n604 12.0247
R1996 VTAIL.n32 VTAIL.n24 12.0247
R1997 VTAIL.n69 VTAIL.n68 12.0247
R1998 VTAIL.n81 VTAIL.n2 12.0247
R1999 VTAIL.n118 VTAIL.n110 12.0247
R2000 VTAIL.n155 VTAIL.n154 12.0247
R2001 VTAIL.n167 VTAIL.n88 12.0247
R2002 VTAIL.n204 VTAIL.n196 12.0247
R2003 VTAIL.n241 VTAIL.n240 12.0247
R2004 VTAIL.n253 VTAIL.n174 12.0247
R2005 VTAIL.n597 VTAIL.n518 12.0247
R2006 VTAIL.n586 VTAIL.n523 12.0247
R2007 VTAIL.n550 VTAIL.n542 12.0247
R2008 VTAIL.n511 VTAIL.n432 12.0247
R2009 VTAIL.n500 VTAIL.n437 12.0247
R2010 VTAIL.n464 VTAIL.n456 12.0247
R2011 VTAIL.n425 VTAIL.n346 12.0247
R2012 VTAIL.n414 VTAIL.n351 12.0247
R2013 VTAIL.n378 VTAIL.n370 12.0247
R2014 VTAIL.n339 VTAIL.n260 12.0247
R2015 VTAIL.n328 VTAIL.n265 12.0247
R2016 VTAIL.n292 VTAIL.n284 12.0247
R2017 VTAIL.n638 VTAIL.n637 11.249
R2018 VTAIL.n669 VTAIL.n610 11.249
R2019 VTAIL.n684 VTAIL.n602 11.249
R2020 VTAIL.n36 VTAIL.n35 11.249
R2021 VTAIL.n67 VTAIL.n8 11.249
R2022 VTAIL.n82 VTAIL.n0 11.249
R2023 VTAIL.n122 VTAIL.n121 11.249
R2024 VTAIL.n153 VTAIL.n94 11.249
R2025 VTAIL.n168 VTAIL.n86 11.249
R2026 VTAIL.n208 VTAIL.n207 11.249
R2027 VTAIL.n239 VTAIL.n180 11.249
R2028 VTAIL.n254 VTAIL.n172 11.249
R2029 VTAIL.n598 VTAIL.n516 11.249
R2030 VTAIL.n585 VTAIL.n526 11.249
R2031 VTAIL.n554 VTAIL.n553 11.249
R2032 VTAIL.n512 VTAIL.n430 11.249
R2033 VTAIL.n499 VTAIL.n440 11.249
R2034 VTAIL.n468 VTAIL.n467 11.249
R2035 VTAIL.n426 VTAIL.n344 11.249
R2036 VTAIL.n413 VTAIL.n354 11.249
R2037 VTAIL.n382 VTAIL.n381 11.249
R2038 VTAIL.n340 VTAIL.n258 11.249
R2039 VTAIL.n327 VTAIL.n268 11.249
R2040 VTAIL.n296 VTAIL.n295 11.249
R2041 VTAIL.n641 VTAIL.n624 10.4732
R2042 VTAIL.n666 VTAIL.n665 10.4732
R2043 VTAIL.n39 VTAIL.n22 10.4732
R2044 VTAIL.n64 VTAIL.n63 10.4732
R2045 VTAIL.n125 VTAIL.n108 10.4732
R2046 VTAIL.n150 VTAIL.n149 10.4732
R2047 VTAIL.n211 VTAIL.n194 10.4732
R2048 VTAIL.n236 VTAIL.n235 10.4732
R2049 VTAIL.n582 VTAIL.n581 10.4732
R2050 VTAIL.n557 VTAIL.n540 10.4732
R2051 VTAIL.n496 VTAIL.n495 10.4732
R2052 VTAIL.n471 VTAIL.n454 10.4732
R2053 VTAIL.n410 VTAIL.n409 10.4732
R2054 VTAIL.n385 VTAIL.n368 10.4732
R2055 VTAIL.n324 VTAIL.n323 10.4732
R2056 VTAIL.n299 VTAIL.n282 10.4732
R2057 VTAIL.n642 VTAIL.n622 9.69747
R2058 VTAIL.n662 VTAIL.n612 9.69747
R2059 VTAIL.n40 VTAIL.n20 9.69747
R2060 VTAIL.n60 VTAIL.n10 9.69747
R2061 VTAIL.n126 VTAIL.n106 9.69747
R2062 VTAIL.n146 VTAIL.n96 9.69747
R2063 VTAIL.n212 VTAIL.n192 9.69747
R2064 VTAIL.n232 VTAIL.n182 9.69747
R2065 VTAIL.n578 VTAIL.n528 9.69747
R2066 VTAIL.n558 VTAIL.n538 9.69747
R2067 VTAIL.n492 VTAIL.n442 9.69747
R2068 VTAIL.n472 VTAIL.n452 9.69747
R2069 VTAIL.n406 VTAIL.n356 9.69747
R2070 VTAIL.n386 VTAIL.n366 9.69747
R2071 VTAIL.n320 VTAIL.n270 9.69747
R2072 VTAIL.n300 VTAIL.n280 9.69747
R2073 VTAIL.n686 VTAIL.n685 9.45567
R2074 VTAIL.n84 VTAIL.n83 9.45567
R2075 VTAIL.n170 VTAIL.n169 9.45567
R2076 VTAIL.n256 VTAIL.n255 9.45567
R2077 VTAIL.n600 VTAIL.n599 9.45567
R2078 VTAIL.n514 VTAIL.n513 9.45567
R2079 VTAIL.n428 VTAIL.n427 9.45567
R2080 VTAIL.n342 VTAIL.n341 9.45567
R2081 VTAIL.n685 VTAIL.n684 9.3005
R2082 VTAIL.n604 VTAIL.n603 9.3005
R2083 VTAIL.n679 VTAIL.n678 9.3005
R2084 VTAIL.n651 VTAIL.n650 9.3005
R2085 VTAIL.n620 VTAIL.n619 9.3005
R2086 VTAIL.n645 VTAIL.n644 9.3005
R2087 VTAIL.n643 VTAIL.n642 9.3005
R2088 VTAIL.n624 VTAIL.n623 9.3005
R2089 VTAIL.n637 VTAIL.n636 9.3005
R2090 VTAIL.n635 VTAIL.n634 9.3005
R2091 VTAIL.n628 VTAIL.n627 9.3005
R2092 VTAIL.n653 VTAIL.n652 9.3005
R2093 VTAIL.n616 VTAIL.n615 9.3005
R2094 VTAIL.n659 VTAIL.n658 9.3005
R2095 VTAIL.n661 VTAIL.n660 9.3005
R2096 VTAIL.n612 VTAIL.n611 9.3005
R2097 VTAIL.n667 VTAIL.n666 9.3005
R2098 VTAIL.n669 VTAIL.n668 9.3005
R2099 VTAIL.n670 VTAIL.n607 9.3005
R2100 VTAIL.n677 VTAIL.n676 9.3005
R2101 VTAIL.n83 VTAIL.n82 9.3005
R2102 VTAIL.n2 VTAIL.n1 9.3005
R2103 VTAIL.n77 VTAIL.n76 9.3005
R2104 VTAIL.n49 VTAIL.n48 9.3005
R2105 VTAIL.n18 VTAIL.n17 9.3005
R2106 VTAIL.n43 VTAIL.n42 9.3005
R2107 VTAIL.n41 VTAIL.n40 9.3005
R2108 VTAIL.n22 VTAIL.n21 9.3005
R2109 VTAIL.n35 VTAIL.n34 9.3005
R2110 VTAIL.n33 VTAIL.n32 9.3005
R2111 VTAIL.n26 VTAIL.n25 9.3005
R2112 VTAIL.n51 VTAIL.n50 9.3005
R2113 VTAIL.n14 VTAIL.n13 9.3005
R2114 VTAIL.n57 VTAIL.n56 9.3005
R2115 VTAIL.n59 VTAIL.n58 9.3005
R2116 VTAIL.n10 VTAIL.n9 9.3005
R2117 VTAIL.n65 VTAIL.n64 9.3005
R2118 VTAIL.n67 VTAIL.n66 9.3005
R2119 VTAIL.n68 VTAIL.n5 9.3005
R2120 VTAIL.n75 VTAIL.n74 9.3005
R2121 VTAIL.n169 VTAIL.n168 9.3005
R2122 VTAIL.n88 VTAIL.n87 9.3005
R2123 VTAIL.n163 VTAIL.n162 9.3005
R2124 VTAIL.n135 VTAIL.n134 9.3005
R2125 VTAIL.n104 VTAIL.n103 9.3005
R2126 VTAIL.n129 VTAIL.n128 9.3005
R2127 VTAIL.n127 VTAIL.n126 9.3005
R2128 VTAIL.n108 VTAIL.n107 9.3005
R2129 VTAIL.n121 VTAIL.n120 9.3005
R2130 VTAIL.n119 VTAIL.n118 9.3005
R2131 VTAIL.n112 VTAIL.n111 9.3005
R2132 VTAIL.n137 VTAIL.n136 9.3005
R2133 VTAIL.n100 VTAIL.n99 9.3005
R2134 VTAIL.n143 VTAIL.n142 9.3005
R2135 VTAIL.n145 VTAIL.n144 9.3005
R2136 VTAIL.n96 VTAIL.n95 9.3005
R2137 VTAIL.n151 VTAIL.n150 9.3005
R2138 VTAIL.n153 VTAIL.n152 9.3005
R2139 VTAIL.n154 VTAIL.n91 9.3005
R2140 VTAIL.n161 VTAIL.n160 9.3005
R2141 VTAIL.n255 VTAIL.n254 9.3005
R2142 VTAIL.n174 VTAIL.n173 9.3005
R2143 VTAIL.n249 VTAIL.n248 9.3005
R2144 VTAIL.n221 VTAIL.n220 9.3005
R2145 VTAIL.n190 VTAIL.n189 9.3005
R2146 VTAIL.n215 VTAIL.n214 9.3005
R2147 VTAIL.n213 VTAIL.n212 9.3005
R2148 VTAIL.n194 VTAIL.n193 9.3005
R2149 VTAIL.n207 VTAIL.n206 9.3005
R2150 VTAIL.n205 VTAIL.n204 9.3005
R2151 VTAIL.n198 VTAIL.n197 9.3005
R2152 VTAIL.n223 VTAIL.n222 9.3005
R2153 VTAIL.n186 VTAIL.n185 9.3005
R2154 VTAIL.n229 VTAIL.n228 9.3005
R2155 VTAIL.n231 VTAIL.n230 9.3005
R2156 VTAIL.n182 VTAIL.n181 9.3005
R2157 VTAIL.n237 VTAIL.n236 9.3005
R2158 VTAIL.n239 VTAIL.n238 9.3005
R2159 VTAIL.n240 VTAIL.n177 9.3005
R2160 VTAIL.n247 VTAIL.n246 9.3005
R2161 VTAIL.n532 VTAIL.n531 9.3005
R2162 VTAIL.n575 VTAIL.n574 9.3005
R2163 VTAIL.n577 VTAIL.n576 9.3005
R2164 VTAIL.n528 VTAIL.n527 9.3005
R2165 VTAIL.n583 VTAIL.n582 9.3005
R2166 VTAIL.n585 VTAIL.n584 9.3005
R2167 VTAIL.n523 VTAIL.n521 9.3005
R2168 VTAIL.n591 VTAIL.n590 9.3005
R2169 VTAIL.n599 VTAIL.n598 9.3005
R2170 VTAIL.n518 VTAIL.n517 9.3005
R2171 VTAIL.n593 VTAIL.n592 9.3005
R2172 VTAIL.n569 VTAIL.n568 9.3005
R2173 VTAIL.n567 VTAIL.n566 9.3005
R2174 VTAIL.n536 VTAIL.n535 9.3005
R2175 VTAIL.n561 VTAIL.n560 9.3005
R2176 VTAIL.n559 VTAIL.n558 9.3005
R2177 VTAIL.n540 VTAIL.n539 9.3005
R2178 VTAIL.n553 VTAIL.n552 9.3005
R2179 VTAIL.n551 VTAIL.n550 9.3005
R2180 VTAIL.n544 VTAIL.n543 9.3005
R2181 VTAIL.n446 VTAIL.n445 9.3005
R2182 VTAIL.n489 VTAIL.n488 9.3005
R2183 VTAIL.n491 VTAIL.n490 9.3005
R2184 VTAIL.n442 VTAIL.n441 9.3005
R2185 VTAIL.n497 VTAIL.n496 9.3005
R2186 VTAIL.n499 VTAIL.n498 9.3005
R2187 VTAIL.n437 VTAIL.n435 9.3005
R2188 VTAIL.n505 VTAIL.n504 9.3005
R2189 VTAIL.n513 VTAIL.n512 9.3005
R2190 VTAIL.n432 VTAIL.n431 9.3005
R2191 VTAIL.n507 VTAIL.n506 9.3005
R2192 VTAIL.n483 VTAIL.n482 9.3005
R2193 VTAIL.n481 VTAIL.n480 9.3005
R2194 VTAIL.n450 VTAIL.n449 9.3005
R2195 VTAIL.n475 VTAIL.n474 9.3005
R2196 VTAIL.n473 VTAIL.n472 9.3005
R2197 VTAIL.n454 VTAIL.n453 9.3005
R2198 VTAIL.n467 VTAIL.n466 9.3005
R2199 VTAIL.n465 VTAIL.n464 9.3005
R2200 VTAIL.n458 VTAIL.n457 9.3005
R2201 VTAIL.n360 VTAIL.n359 9.3005
R2202 VTAIL.n403 VTAIL.n402 9.3005
R2203 VTAIL.n405 VTAIL.n404 9.3005
R2204 VTAIL.n356 VTAIL.n355 9.3005
R2205 VTAIL.n411 VTAIL.n410 9.3005
R2206 VTAIL.n413 VTAIL.n412 9.3005
R2207 VTAIL.n351 VTAIL.n349 9.3005
R2208 VTAIL.n419 VTAIL.n418 9.3005
R2209 VTAIL.n427 VTAIL.n426 9.3005
R2210 VTAIL.n346 VTAIL.n345 9.3005
R2211 VTAIL.n421 VTAIL.n420 9.3005
R2212 VTAIL.n397 VTAIL.n396 9.3005
R2213 VTAIL.n395 VTAIL.n394 9.3005
R2214 VTAIL.n364 VTAIL.n363 9.3005
R2215 VTAIL.n389 VTAIL.n388 9.3005
R2216 VTAIL.n387 VTAIL.n386 9.3005
R2217 VTAIL.n368 VTAIL.n367 9.3005
R2218 VTAIL.n381 VTAIL.n380 9.3005
R2219 VTAIL.n379 VTAIL.n378 9.3005
R2220 VTAIL.n372 VTAIL.n371 9.3005
R2221 VTAIL.n274 VTAIL.n273 9.3005
R2222 VTAIL.n317 VTAIL.n316 9.3005
R2223 VTAIL.n319 VTAIL.n318 9.3005
R2224 VTAIL.n270 VTAIL.n269 9.3005
R2225 VTAIL.n325 VTAIL.n324 9.3005
R2226 VTAIL.n327 VTAIL.n326 9.3005
R2227 VTAIL.n265 VTAIL.n263 9.3005
R2228 VTAIL.n333 VTAIL.n332 9.3005
R2229 VTAIL.n341 VTAIL.n340 9.3005
R2230 VTAIL.n260 VTAIL.n259 9.3005
R2231 VTAIL.n335 VTAIL.n334 9.3005
R2232 VTAIL.n311 VTAIL.n310 9.3005
R2233 VTAIL.n309 VTAIL.n308 9.3005
R2234 VTAIL.n278 VTAIL.n277 9.3005
R2235 VTAIL.n303 VTAIL.n302 9.3005
R2236 VTAIL.n301 VTAIL.n300 9.3005
R2237 VTAIL.n282 VTAIL.n281 9.3005
R2238 VTAIL.n295 VTAIL.n294 9.3005
R2239 VTAIL.n293 VTAIL.n292 9.3005
R2240 VTAIL.n286 VTAIL.n285 9.3005
R2241 VTAIL.n646 VTAIL.n645 8.92171
R2242 VTAIL.n661 VTAIL.n614 8.92171
R2243 VTAIL.n44 VTAIL.n43 8.92171
R2244 VTAIL.n59 VTAIL.n12 8.92171
R2245 VTAIL.n130 VTAIL.n129 8.92171
R2246 VTAIL.n145 VTAIL.n98 8.92171
R2247 VTAIL.n216 VTAIL.n215 8.92171
R2248 VTAIL.n231 VTAIL.n184 8.92171
R2249 VTAIL.n577 VTAIL.n530 8.92171
R2250 VTAIL.n562 VTAIL.n561 8.92171
R2251 VTAIL.n491 VTAIL.n444 8.92171
R2252 VTAIL.n476 VTAIL.n475 8.92171
R2253 VTAIL.n405 VTAIL.n358 8.92171
R2254 VTAIL.n390 VTAIL.n389 8.92171
R2255 VTAIL.n319 VTAIL.n272 8.92171
R2256 VTAIL.n304 VTAIL.n303 8.92171
R2257 VTAIL.n649 VTAIL.n620 8.14595
R2258 VTAIL.n658 VTAIL.n657 8.14595
R2259 VTAIL.n47 VTAIL.n18 8.14595
R2260 VTAIL.n56 VTAIL.n55 8.14595
R2261 VTAIL.n133 VTAIL.n104 8.14595
R2262 VTAIL.n142 VTAIL.n141 8.14595
R2263 VTAIL.n219 VTAIL.n190 8.14595
R2264 VTAIL.n228 VTAIL.n227 8.14595
R2265 VTAIL.n574 VTAIL.n573 8.14595
R2266 VTAIL.n565 VTAIL.n536 8.14595
R2267 VTAIL.n488 VTAIL.n487 8.14595
R2268 VTAIL.n479 VTAIL.n450 8.14595
R2269 VTAIL.n402 VTAIL.n401 8.14595
R2270 VTAIL.n393 VTAIL.n364 8.14595
R2271 VTAIL.n316 VTAIL.n315 8.14595
R2272 VTAIL.n307 VTAIL.n278 8.14595
R2273 VTAIL.n650 VTAIL.n618 7.3702
R2274 VTAIL.n654 VTAIL.n616 7.3702
R2275 VTAIL.n48 VTAIL.n16 7.3702
R2276 VTAIL.n52 VTAIL.n14 7.3702
R2277 VTAIL.n134 VTAIL.n102 7.3702
R2278 VTAIL.n138 VTAIL.n100 7.3702
R2279 VTAIL.n220 VTAIL.n188 7.3702
R2280 VTAIL.n224 VTAIL.n186 7.3702
R2281 VTAIL.n570 VTAIL.n532 7.3702
R2282 VTAIL.n566 VTAIL.n534 7.3702
R2283 VTAIL.n484 VTAIL.n446 7.3702
R2284 VTAIL.n480 VTAIL.n448 7.3702
R2285 VTAIL.n398 VTAIL.n360 7.3702
R2286 VTAIL.n394 VTAIL.n362 7.3702
R2287 VTAIL.n312 VTAIL.n274 7.3702
R2288 VTAIL.n308 VTAIL.n276 7.3702
R2289 VTAIL.n653 VTAIL.n618 6.59444
R2290 VTAIL.n654 VTAIL.n653 6.59444
R2291 VTAIL.n51 VTAIL.n16 6.59444
R2292 VTAIL.n52 VTAIL.n51 6.59444
R2293 VTAIL.n137 VTAIL.n102 6.59444
R2294 VTAIL.n138 VTAIL.n137 6.59444
R2295 VTAIL.n223 VTAIL.n188 6.59444
R2296 VTAIL.n224 VTAIL.n223 6.59444
R2297 VTAIL.n570 VTAIL.n569 6.59444
R2298 VTAIL.n569 VTAIL.n534 6.59444
R2299 VTAIL.n484 VTAIL.n483 6.59444
R2300 VTAIL.n483 VTAIL.n448 6.59444
R2301 VTAIL.n398 VTAIL.n397 6.59444
R2302 VTAIL.n397 VTAIL.n362 6.59444
R2303 VTAIL.n312 VTAIL.n311 6.59444
R2304 VTAIL.n311 VTAIL.n276 6.59444
R2305 VTAIL.n650 VTAIL.n649 5.81868
R2306 VTAIL.n657 VTAIL.n616 5.81868
R2307 VTAIL.n48 VTAIL.n47 5.81868
R2308 VTAIL.n55 VTAIL.n14 5.81868
R2309 VTAIL.n134 VTAIL.n133 5.81868
R2310 VTAIL.n141 VTAIL.n100 5.81868
R2311 VTAIL.n220 VTAIL.n219 5.81868
R2312 VTAIL.n227 VTAIL.n186 5.81868
R2313 VTAIL.n573 VTAIL.n532 5.81868
R2314 VTAIL.n566 VTAIL.n565 5.81868
R2315 VTAIL.n487 VTAIL.n446 5.81868
R2316 VTAIL.n480 VTAIL.n479 5.81868
R2317 VTAIL.n401 VTAIL.n360 5.81868
R2318 VTAIL.n394 VTAIL.n393 5.81868
R2319 VTAIL.n315 VTAIL.n274 5.81868
R2320 VTAIL.n308 VTAIL.n307 5.81868
R2321 VTAIL.n646 VTAIL.n620 5.04292
R2322 VTAIL.n658 VTAIL.n614 5.04292
R2323 VTAIL.n44 VTAIL.n18 5.04292
R2324 VTAIL.n56 VTAIL.n12 5.04292
R2325 VTAIL.n130 VTAIL.n104 5.04292
R2326 VTAIL.n142 VTAIL.n98 5.04292
R2327 VTAIL.n216 VTAIL.n190 5.04292
R2328 VTAIL.n228 VTAIL.n184 5.04292
R2329 VTAIL.n574 VTAIL.n530 5.04292
R2330 VTAIL.n562 VTAIL.n536 5.04292
R2331 VTAIL.n488 VTAIL.n444 5.04292
R2332 VTAIL.n476 VTAIL.n450 5.04292
R2333 VTAIL.n402 VTAIL.n358 5.04292
R2334 VTAIL.n390 VTAIL.n364 5.04292
R2335 VTAIL.n316 VTAIL.n272 5.04292
R2336 VTAIL.n304 VTAIL.n278 5.04292
R2337 VTAIL.n629 VTAIL.n627 4.38563
R2338 VTAIL.n27 VTAIL.n25 4.38563
R2339 VTAIL.n113 VTAIL.n111 4.38563
R2340 VTAIL.n199 VTAIL.n197 4.38563
R2341 VTAIL.n545 VTAIL.n543 4.38563
R2342 VTAIL.n459 VTAIL.n457 4.38563
R2343 VTAIL.n373 VTAIL.n371 4.38563
R2344 VTAIL.n287 VTAIL.n285 4.38563
R2345 VTAIL.n645 VTAIL.n622 4.26717
R2346 VTAIL.n662 VTAIL.n661 4.26717
R2347 VTAIL.n43 VTAIL.n20 4.26717
R2348 VTAIL.n60 VTAIL.n59 4.26717
R2349 VTAIL.n129 VTAIL.n106 4.26717
R2350 VTAIL.n146 VTAIL.n145 4.26717
R2351 VTAIL.n215 VTAIL.n192 4.26717
R2352 VTAIL.n232 VTAIL.n231 4.26717
R2353 VTAIL.n578 VTAIL.n577 4.26717
R2354 VTAIL.n561 VTAIL.n538 4.26717
R2355 VTAIL.n492 VTAIL.n491 4.26717
R2356 VTAIL.n475 VTAIL.n452 4.26717
R2357 VTAIL.n406 VTAIL.n405 4.26717
R2358 VTAIL.n389 VTAIL.n366 4.26717
R2359 VTAIL.n320 VTAIL.n319 4.26717
R2360 VTAIL.n303 VTAIL.n280 4.26717
R2361 VTAIL.n642 VTAIL.n641 3.49141
R2362 VTAIL.n665 VTAIL.n612 3.49141
R2363 VTAIL.n40 VTAIL.n39 3.49141
R2364 VTAIL.n63 VTAIL.n10 3.49141
R2365 VTAIL.n126 VTAIL.n125 3.49141
R2366 VTAIL.n149 VTAIL.n96 3.49141
R2367 VTAIL.n212 VTAIL.n211 3.49141
R2368 VTAIL.n235 VTAIL.n182 3.49141
R2369 VTAIL.n581 VTAIL.n528 3.49141
R2370 VTAIL.n558 VTAIL.n557 3.49141
R2371 VTAIL.n495 VTAIL.n442 3.49141
R2372 VTAIL.n472 VTAIL.n471 3.49141
R2373 VTAIL.n409 VTAIL.n356 3.49141
R2374 VTAIL.n386 VTAIL.n385 3.49141
R2375 VTAIL.n323 VTAIL.n270 3.49141
R2376 VTAIL.n300 VTAIL.n299 3.49141
R2377 VTAIL.n638 VTAIL.n624 2.71565
R2378 VTAIL.n666 VTAIL.n610 2.71565
R2379 VTAIL.n686 VTAIL.n602 2.71565
R2380 VTAIL.n36 VTAIL.n22 2.71565
R2381 VTAIL.n64 VTAIL.n8 2.71565
R2382 VTAIL.n84 VTAIL.n0 2.71565
R2383 VTAIL.n122 VTAIL.n108 2.71565
R2384 VTAIL.n150 VTAIL.n94 2.71565
R2385 VTAIL.n170 VTAIL.n86 2.71565
R2386 VTAIL.n208 VTAIL.n194 2.71565
R2387 VTAIL.n236 VTAIL.n180 2.71565
R2388 VTAIL.n256 VTAIL.n172 2.71565
R2389 VTAIL.n600 VTAIL.n516 2.71565
R2390 VTAIL.n582 VTAIL.n526 2.71565
R2391 VTAIL.n554 VTAIL.n540 2.71565
R2392 VTAIL.n514 VTAIL.n430 2.71565
R2393 VTAIL.n496 VTAIL.n440 2.71565
R2394 VTAIL.n468 VTAIL.n454 2.71565
R2395 VTAIL.n428 VTAIL.n344 2.71565
R2396 VTAIL.n410 VTAIL.n354 2.71565
R2397 VTAIL.n382 VTAIL.n368 2.71565
R2398 VTAIL.n342 VTAIL.n258 2.71565
R2399 VTAIL.n324 VTAIL.n268 2.71565
R2400 VTAIL.n296 VTAIL.n282 2.71565
R2401 VTAIL.n429 VTAIL.n343 2.56084
R2402 VTAIL.n601 VTAIL.n515 2.56084
R2403 VTAIL.n257 VTAIL.n171 2.56084
R2404 VTAIL.n637 VTAIL.n626 1.93989
R2405 VTAIL.n671 VTAIL.n669 1.93989
R2406 VTAIL.n684 VTAIL.n683 1.93989
R2407 VTAIL.n35 VTAIL.n24 1.93989
R2408 VTAIL.n69 VTAIL.n67 1.93989
R2409 VTAIL.n82 VTAIL.n81 1.93989
R2410 VTAIL.n121 VTAIL.n110 1.93989
R2411 VTAIL.n155 VTAIL.n153 1.93989
R2412 VTAIL.n168 VTAIL.n167 1.93989
R2413 VTAIL.n207 VTAIL.n196 1.93989
R2414 VTAIL.n241 VTAIL.n239 1.93989
R2415 VTAIL.n254 VTAIL.n253 1.93989
R2416 VTAIL.n598 VTAIL.n597 1.93989
R2417 VTAIL.n586 VTAIL.n585 1.93989
R2418 VTAIL.n553 VTAIL.n542 1.93989
R2419 VTAIL.n512 VTAIL.n511 1.93989
R2420 VTAIL.n500 VTAIL.n499 1.93989
R2421 VTAIL.n467 VTAIL.n456 1.93989
R2422 VTAIL.n426 VTAIL.n425 1.93989
R2423 VTAIL.n414 VTAIL.n413 1.93989
R2424 VTAIL.n381 VTAIL.n370 1.93989
R2425 VTAIL.n340 VTAIL.n339 1.93989
R2426 VTAIL.n328 VTAIL.n327 1.93989
R2427 VTAIL.n295 VTAIL.n284 1.93989
R2428 VTAIL VTAIL.n85 1.33886
R2429 VTAIL VTAIL.n687 1.22248
R2430 VTAIL.n634 VTAIL.n633 1.16414
R2431 VTAIL.n670 VTAIL.n608 1.16414
R2432 VTAIL.n680 VTAIL.n604 1.16414
R2433 VTAIL.n32 VTAIL.n31 1.16414
R2434 VTAIL.n68 VTAIL.n6 1.16414
R2435 VTAIL.n78 VTAIL.n2 1.16414
R2436 VTAIL.n118 VTAIL.n117 1.16414
R2437 VTAIL.n154 VTAIL.n92 1.16414
R2438 VTAIL.n164 VTAIL.n88 1.16414
R2439 VTAIL.n204 VTAIL.n203 1.16414
R2440 VTAIL.n240 VTAIL.n178 1.16414
R2441 VTAIL.n250 VTAIL.n174 1.16414
R2442 VTAIL.n594 VTAIL.n518 1.16414
R2443 VTAIL.n589 VTAIL.n523 1.16414
R2444 VTAIL.n550 VTAIL.n549 1.16414
R2445 VTAIL.n508 VTAIL.n432 1.16414
R2446 VTAIL.n503 VTAIL.n437 1.16414
R2447 VTAIL.n464 VTAIL.n463 1.16414
R2448 VTAIL.n422 VTAIL.n346 1.16414
R2449 VTAIL.n417 VTAIL.n351 1.16414
R2450 VTAIL.n378 VTAIL.n377 1.16414
R2451 VTAIL.n336 VTAIL.n260 1.16414
R2452 VTAIL.n331 VTAIL.n265 1.16414
R2453 VTAIL.n292 VTAIL.n291 1.16414
R2454 VTAIL.n515 VTAIL.n429 0.470328
R2455 VTAIL.n171 VTAIL.n85 0.470328
R2456 VTAIL.n630 VTAIL.n628 0.388379
R2457 VTAIL.n676 VTAIL.n675 0.388379
R2458 VTAIL.n679 VTAIL.n606 0.388379
R2459 VTAIL.n28 VTAIL.n26 0.388379
R2460 VTAIL.n74 VTAIL.n73 0.388379
R2461 VTAIL.n77 VTAIL.n4 0.388379
R2462 VTAIL.n114 VTAIL.n112 0.388379
R2463 VTAIL.n160 VTAIL.n159 0.388379
R2464 VTAIL.n163 VTAIL.n90 0.388379
R2465 VTAIL.n200 VTAIL.n198 0.388379
R2466 VTAIL.n246 VTAIL.n245 0.388379
R2467 VTAIL.n249 VTAIL.n176 0.388379
R2468 VTAIL.n593 VTAIL.n520 0.388379
R2469 VTAIL.n590 VTAIL.n522 0.388379
R2470 VTAIL.n546 VTAIL.n544 0.388379
R2471 VTAIL.n507 VTAIL.n434 0.388379
R2472 VTAIL.n504 VTAIL.n436 0.388379
R2473 VTAIL.n460 VTAIL.n458 0.388379
R2474 VTAIL.n421 VTAIL.n348 0.388379
R2475 VTAIL.n418 VTAIL.n350 0.388379
R2476 VTAIL.n374 VTAIL.n372 0.388379
R2477 VTAIL.n335 VTAIL.n262 0.388379
R2478 VTAIL.n332 VTAIL.n264 0.388379
R2479 VTAIL.n288 VTAIL.n286 0.388379
R2480 VTAIL.n635 VTAIL.n627 0.155672
R2481 VTAIL.n636 VTAIL.n635 0.155672
R2482 VTAIL.n636 VTAIL.n623 0.155672
R2483 VTAIL.n643 VTAIL.n623 0.155672
R2484 VTAIL.n644 VTAIL.n643 0.155672
R2485 VTAIL.n644 VTAIL.n619 0.155672
R2486 VTAIL.n651 VTAIL.n619 0.155672
R2487 VTAIL.n652 VTAIL.n651 0.155672
R2488 VTAIL.n652 VTAIL.n615 0.155672
R2489 VTAIL.n659 VTAIL.n615 0.155672
R2490 VTAIL.n660 VTAIL.n659 0.155672
R2491 VTAIL.n660 VTAIL.n611 0.155672
R2492 VTAIL.n667 VTAIL.n611 0.155672
R2493 VTAIL.n668 VTAIL.n667 0.155672
R2494 VTAIL.n668 VTAIL.n607 0.155672
R2495 VTAIL.n677 VTAIL.n607 0.155672
R2496 VTAIL.n678 VTAIL.n677 0.155672
R2497 VTAIL.n678 VTAIL.n603 0.155672
R2498 VTAIL.n685 VTAIL.n603 0.155672
R2499 VTAIL.n33 VTAIL.n25 0.155672
R2500 VTAIL.n34 VTAIL.n33 0.155672
R2501 VTAIL.n34 VTAIL.n21 0.155672
R2502 VTAIL.n41 VTAIL.n21 0.155672
R2503 VTAIL.n42 VTAIL.n41 0.155672
R2504 VTAIL.n42 VTAIL.n17 0.155672
R2505 VTAIL.n49 VTAIL.n17 0.155672
R2506 VTAIL.n50 VTAIL.n49 0.155672
R2507 VTAIL.n50 VTAIL.n13 0.155672
R2508 VTAIL.n57 VTAIL.n13 0.155672
R2509 VTAIL.n58 VTAIL.n57 0.155672
R2510 VTAIL.n58 VTAIL.n9 0.155672
R2511 VTAIL.n65 VTAIL.n9 0.155672
R2512 VTAIL.n66 VTAIL.n65 0.155672
R2513 VTAIL.n66 VTAIL.n5 0.155672
R2514 VTAIL.n75 VTAIL.n5 0.155672
R2515 VTAIL.n76 VTAIL.n75 0.155672
R2516 VTAIL.n76 VTAIL.n1 0.155672
R2517 VTAIL.n83 VTAIL.n1 0.155672
R2518 VTAIL.n119 VTAIL.n111 0.155672
R2519 VTAIL.n120 VTAIL.n119 0.155672
R2520 VTAIL.n120 VTAIL.n107 0.155672
R2521 VTAIL.n127 VTAIL.n107 0.155672
R2522 VTAIL.n128 VTAIL.n127 0.155672
R2523 VTAIL.n128 VTAIL.n103 0.155672
R2524 VTAIL.n135 VTAIL.n103 0.155672
R2525 VTAIL.n136 VTAIL.n135 0.155672
R2526 VTAIL.n136 VTAIL.n99 0.155672
R2527 VTAIL.n143 VTAIL.n99 0.155672
R2528 VTAIL.n144 VTAIL.n143 0.155672
R2529 VTAIL.n144 VTAIL.n95 0.155672
R2530 VTAIL.n151 VTAIL.n95 0.155672
R2531 VTAIL.n152 VTAIL.n151 0.155672
R2532 VTAIL.n152 VTAIL.n91 0.155672
R2533 VTAIL.n161 VTAIL.n91 0.155672
R2534 VTAIL.n162 VTAIL.n161 0.155672
R2535 VTAIL.n162 VTAIL.n87 0.155672
R2536 VTAIL.n169 VTAIL.n87 0.155672
R2537 VTAIL.n205 VTAIL.n197 0.155672
R2538 VTAIL.n206 VTAIL.n205 0.155672
R2539 VTAIL.n206 VTAIL.n193 0.155672
R2540 VTAIL.n213 VTAIL.n193 0.155672
R2541 VTAIL.n214 VTAIL.n213 0.155672
R2542 VTAIL.n214 VTAIL.n189 0.155672
R2543 VTAIL.n221 VTAIL.n189 0.155672
R2544 VTAIL.n222 VTAIL.n221 0.155672
R2545 VTAIL.n222 VTAIL.n185 0.155672
R2546 VTAIL.n229 VTAIL.n185 0.155672
R2547 VTAIL.n230 VTAIL.n229 0.155672
R2548 VTAIL.n230 VTAIL.n181 0.155672
R2549 VTAIL.n237 VTAIL.n181 0.155672
R2550 VTAIL.n238 VTAIL.n237 0.155672
R2551 VTAIL.n238 VTAIL.n177 0.155672
R2552 VTAIL.n247 VTAIL.n177 0.155672
R2553 VTAIL.n248 VTAIL.n247 0.155672
R2554 VTAIL.n248 VTAIL.n173 0.155672
R2555 VTAIL.n255 VTAIL.n173 0.155672
R2556 VTAIL.n599 VTAIL.n517 0.155672
R2557 VTAIL.n592 VTAIL.n517 0.155672
R2558 VTAIL.n592 VTAIL.n591 0.155672
R2559 VTAIL.n591 VTAIL.n521 0.155672
R2560 VTAIL.n584 VTAIL.n521 0.155672
R2561 VTAIL.n584 VTAIL.n583 0.155672
R2562 VTAIL.n583 VTAIL.n527 0.155672
R2563 VTAIL.n576 VTAIL.n527 0.155672
R2564 VTAIL.n576 VTAIL.n575 0.155672
R2565 VTAIL.n575 VTAIL.n531 0.155672
R2566 VTAIL.n568 VTAIL.n531 0.155672
R2567 VTAIL.n568 VTAIL.n567 0.155672
R2568 VTAIL.n567 VTAIL.n535 0.155672
R2569 VTAIL.n560 VTAIL.n535 0.155672
R2570 VTAIL.n560 VTAIL.n559 0.155672
R2571 VTAIL.n559 VTAIL.n539 0.155672
R2572 VTAIL.n552 VTAIL.n539 0.155672
R2573 VTAIL.n552 VTAIL.n551 0.155672
R2574 VTAIL.n551 VTAIL.n543 0.155672
R2575 VTAIL.n513 VTAIL.n431 0.155672
R2576 VTAIL.n506 VTAIL.n431 0.155672
R2577 VTAIL.n506 VTAIL.n505 0.155672
R2578 VTAIL.n505 VTAIL.n435 0.155672
R2579 VTAIL.n498 VTAIL.n435 0.155672
R2580 VTAIL.n498 VTAIL.n497 0.155672
R2581 VTAIL.n497 VTAIL.n441 0.155672
R2582 VTAIL.n490 VTAIL.n441 0.155672
R2583 VTAIL.n490 VTAIL.n489 0.155672
R2584 VTAIL.n489 VTAIL.n445 0.155672
R2585 VTAIL.n482 VTAIL.n445 0.155672
R2586 VTAIL.n482 VTAIL.n481 0.155672
R2587 VTAIL.n481 VTAIL.n449 0.155672
R2588 VTAIL.n474 VTAIL.n449 0.155672
R2589 VTAIL.n474 VTAIL.n473 0.155672
R2590 VTAIL.n473 VTAIL.n453 0.155672
R2591 VTAIL.n466 VTAIL.n453 0.155672
R2592 VTAIL.n466 VTAIL.n465 0.155672
R2593 VTAIL.n465 VTAIL.n457 0.155672
R2594 VTAIL.n427 VTAIL.n345 0.155672
R2595 VTAIL.n420 VTAIL.n345 0.155672
R2596 VTAIL.n420 VTAIL.n419 0.155672
R2597 VTAIL.n419 VTAIL.n349 0.155672
R2598 VTAIL.n412 VTAIL.n349 0.155672
R2599 VTAIL.n412 VTAIL.n411 0.155672
R2600 VTAIL.n411 VTAIL.n355 0.155672
R2601 VTAIL.n404 VTAIL.n355 0.155672
R2602 VTAIL.n404 VTAIL.n403 0.155672
R2603 VTAIL.n403 VTAIL.n359 0.155672
R2604 VTAIL.n396 VTAIL.n359 0.155672
R2605 VTAIL.n396 VTAIL.n395 0.155672
R2606 VTAIL.n395 VTAIL.n363 0.155672
R2607 VTAIL.n388 VTAIL.n363 0.155672
R2608 VTAIL.n388 VTAIL.n387 0.155672
R2609 VTAIL.n387 VTAIL.n367 0.155672
R2610 VTAIL.n380 VTAIL.n367 0.155672
R2611 VTAIL.n380 VTAIL.n379 0.155672
R2612 VTAIL.n379 VTAIL.n371 0.155672
R2613 VTAIL.n341 VTAIL.n259 0.155672
R2614 VTAIL.n334 VTAIL.n259 0.155672
R2615 VTAIL.n334 VTAIL.n333 0.155672
R2616 VTAIL.n333 VTAIL.n263 0.155672
R2617 VTAIL.n326 VTAIL.n263 0.155672
R2618 VTAIL.n326 VTAIL.n325 0.155672
R2619 VTAIL.n325 VTAIL.n269 0.155672
R2620 VTAIL.n318 VTAIL.n269 0.155672
R2621 VTAIL.n318 VTAIL.n317 0.155672
R2622 VTAIL.n317 VTAIL.n273 0.155672
R2623 VTAIL.n310 VTAIL.n273 0.155672
R2624 VTAIL.n310 VTAIL.n309 0.155672
R2625 VTAIL.n309 VTAIL.n277 0.155672
R2626 VTAIL.n302 VTAIL.n277 0.155672
R2627 VTAIL.n302 VTAIL.n301 0.155672
R2628 VTAIL.n301 VTAIL.n281 0.155672
R2629 VTAIL.n294 VTAIL.n281 0.155672
R2630 VTAIL.n294 VTAIL.n293 0.155672
R2631 VTAIL.n293 VTAIL.n285 0.155672
R2632 VN.n0 VN.t0 176.411
R2633 VN.n1 VN.t1 176.411
R2634 VN.n0 VN.t3 175.627
R2635 VN.n1 VN.t2 175.627
R2636 VN VN.n1 53.5166
R2637 VN VN.n0 4.24007
R2638 VDD2.n2 VDD2.n0 104.669
R2639 VDD2.n2 VDD2.n1 60.0666
R2640 VDD2.n1 VDD2.t1 1.29293
R2641 VDD2.n1 VDD2.t2 1.29293
R2642 VDD2.n0 VDD2.t3 1.29293
R2643 VDD2.n0 VDD2.t0 1.29293
R2644 VDD2 VDD2.n2 0.0586897
C0 VTAIL VDD1 6.19892f
C1 VN VDD2 5.990819f
C2 VDD1 VDD2 1.03068f
C3 VTAIL VDD2 6.25339f
C4 VP VN 6.82755f
C5 VP VDD1 6.23788f
C6 VP VTAIL 5.7746f
C7 VP VDD2 0.39732f
C8 VN VDD1 0.149505f
C9 VN VTAIL 5.7605f
C10 VDD2 B 4.059964f
C11 VDD1 B 8.522449f
C12 VTAIL B 12.095297f
C13 VN B 11.032001f
C14 VP B 9.233464f
C15 VDD2.t3 B 0.323769f
C16 VDD2.t0 B 0.323769f
C17 VDD2.n0 B 3.73524f
C18 VDD2.t1 B 0.323769f
C19 VDD2.t2 B 0.323769f
C20 VDD2.n1 B 2.92828f
C21 VDD2.n2 B 4.11501f
C22 VN.t0 B 2.94017f
C23 VN.t3 B 2.93541f
C24 VN.n0 B 1.86381f
C25 VN.t1 B 2.94017f
C26 VN.t2 B 2.93541f
C27 VN.n1 B 3.29255f
C28 VTAIL.n0 B 0.020083f
C29 VTAIL.n1 B 0.015806f
C30 VTAIL.n2 B 0.008493f
C31 VTAIL.n3 B 0.020075f
C32 VTAIL.n4 B 0.008743f
C33 VTAIL.n5 B 0.015806f
C34 VTAIL.n6 B 0.008993f
C35 VTAIL.n7 B 0.020075f
C36 VTAIL.n8 B 0.008993f
C37 VTAIL.n9 B 0.015806f
C38 VTAIL.n10 B 0.008493f
C39 VTAIL.n11 B 0.020075f
C40 VTAIL.n12 B 0.008993f
C41 VTAIL.n13 B 0.015806f
C42 VTAIL.n14 B 0.008493f
C43 VTAIL.n15 B 0.020075f
C44 VTAIL.n16 B 0.008993f
C45 VTAIL.n17 B 0.015806f
C46 VTAIL.n18 B 0.008493f
C47 VTAIL.n19 B 0.020075f
C48 VTAIL.n20 B 0.008993f
C49 VTAIL.n21 B 0.015806f
C50 VTAIL.n22 B 0.008493f
C51 VTAIL.n23 B 0.020075f
C52 VTAIL.n24 B 0.008993f
C53 VTAIL.n25 B 1.05151f
C54 VTAIL.n26 B 0.008493f
C55 VTAIL.t0 B 0.033118f
C56 VTAIL.n27 B 0.104355f
C57 VTAIL.n28 B 0.011859f
C58 VTAIL.n29 B 0.015056f
C59 VTAIL.n30 B 0.020075f
C60 VTAIL.n31 B 0.008993f
C61 VTAIL.n32 B 0.008493f
C62 VTAIL.n33 B 0.015806f
C63 VTAIL.n34 B 0.015806f
C64 VTAIL.n35 B 0.008493f
C65 VTAIL.n36 B 0.008993f
C66 VTAIL.n37 B 0.020075f
C67 VTAIL.n38 B 0.020075f
C68 VTAIL.n39 B 0.008993f
C69 VTAIL.n40 B 0.008493f
C70 VTAIL.n41 B 0.015806f
C71 VTAIL.n42 B 0.015806f
C72 VTAIL.n43 B 0.008493f
C73 VTAIL.n44 B 0.008993f
C74 VTAIL.n45 B 0.020075f
C75 VTAIL.n46 B 0.020075f
C76 VTAIL.n47 B 0.008993f
C77 VTAIL.n48 B 0.008493f
C78 VTAIL.n49 B 0.015806f
C79 VTAIL.n50 B 0.015806f
C80 VTAIL.n51 B 0.008493f
C81 VTAIL.n52 B 0.008993f
C82 VTAIL.n53 B 0.020075f
C83 VTAIL.n54 B 0.020075f
C84 VTAIL.n55 B 0.008993f
C85 VTAIL.n56 B 0.008493f
C86 VTAIL.n57 B 0.015806f
C87 VTAIL.n58 B 0.015806f
C88 VTAIL.n59 B 0.008493f
C89 VTAIL.n60 B 0.008993f
C90 VTAIL.n61 B 0.020075f
C91 VTAIL.n62 B 0.020075f
C92 VTAIL.n63 B 0.008993f
C93 VTAIL.n64 B 0.008493f
C94 VTAIL.n65 B 0.015806f
C95 VTAIL.n66 B 0.015806f
C96 VTAIL.n67 B 0.008493f
C97 VTAIL.n68 B 0.008493f
C98 VTAIL.n69 B 0.008993f
C99 VTAIL.n70 B 0.020075f
C100 VTAIL.n71 B 0.020075f
C101 VTAIL.n72 B 0.020075f
C102 VTAIL.n73 B 0.008743f
C103 VTAIL.n74 B 0.008493f
C104 VTAIL.n75 B 0.015806f
C105 VTAIL.n76 B 0.015806f
C106 VTAIL.n77 B 0.008493f
C107 VTAIL.n78 B 0.008993f
C108 VTAIL.n79 B 0.020075f
C109 VTAIL.n80 B 0.039687f
C110 VTAIL.n81 B 0.008993f
C111 VTAIL.n82 B 0.008493f
C112 VTAIL.n83 B 0.03567f
C113 VTAIL.n84 B 0.021792f
C114 VTAIL.n85 B 0.105101f
C115 VTAIL.n86 B 0.020083f
C116 VTAIL.n87 B 0.015806f
C117 VTAIL.n88 B 0.008493f
C118 VTAIL.n89 B 0.020075f
C119 VTAIL.n90 B 0.008743f
C120 VTAIL.n91 B 0.015806f
C121 VTAIL.n92 B 0.008993f
C122 VTAIL.n93 B 0.020075f
C123 VTAIL.n94 B 0.008993f
C124 VTAIL.n95 B 0.015806f
C125 VTAIL.n96 B 0.008493f
C126 VTAIL.n97 B 0.020075f
C127 VTAIL.n98 B 0.008993f
C128 VTAIL.n99 B 0.015806f
C129 VTAIL.n100 B 0.008493f
C130 VTAIL.n101 B 0.020075f
C131 VTAIL.n102 B 0.008993f
C132 VTAIL.n103 B 0.015806f
C133 VTAIL.n104 B 0.008493f
C134 VTAIL.n105 B 0.020075f
C135 VTAIL.n106 B 0.008993f
C136 VTAIL.n107 B 0.015806f
C137 VTAIL.n108 B 0.008493f
C138 VTAIL.n109 B 0.020075f
C139 VTAIL.n110 B 0.008993f
C140 VTAIL.n111 B 1.05151f
C141 VTAIL.n112 B 0.008493f
C142 VTAIL.t6 B 0.033118f
C143 VTAIL.n113 B 0.104355f
C144 VTAIL.n114 B 0.011859f
C145 VTAIL.n115 B 0.015056f
C146 VTAIL.n116 B 0.020075f
C147 VTAIL.n117 B 0.008993f
C148 VTAIL.n118 B 0.008493f
C149 VTAIL.n119 B 0.015806f
C150 VTAIL.n120 B 0.015806f
C151 VTAIL.n121 B 0.008493f
C152 VTAIL.n122 B 0.008993f
C153 VTAIL.n123 B 0.020075f
C154 VTAIL.n124 B 0.020075f
C155 VTAIL.n125 B 0.008993f
C156 VTAIL.n126 B 0.008493f
C157 VTAIL.n127 B 0.015806f
C158 VTAIL.n128 B 0.015806f
C159 VTAIL.n129 B 0.008493f
C160 VTAIL.n130 B 0.008993f
C161 VTAIL.n131 B 0.020075f
C162 VTAIL.n132 B 0.020075f
C163 VTAIL.n133 B 0.008993f
C164 VTAIL.n134 B 0.008493f
C165 VTAIL.n135 B 0.015806f
C166 VTAIL.n136 B 0.015806f
C167 VTAIL.n137 B 0.008493f
C168 VTAIL.n138 B 0.008993f
C169 VTAIL.n139 B 0.020075f
C170 VTAIL.n140 B 0.020075f
C171 VTAIL.n141 B 0.008993f
C172 VTAIL.n142 B 0.008493f
C173 VTAIL.n143 B 0.015806f
C174 VTAIL.n144 B 0.015806f
C175 VTAIL.n145 B 0.008493f
C176 VTAIL.n146 B 0.008993f
C177 VTAIL.n147 B 0.020075f
C178 VTAIL.n148 B 0.020075f
C179 VTAIL.n149 B 0.008993f
C180 VTAIL.n150 B 0.008493f
C181 VTAIL.n151 B 0.015806f
C182 VTAIL.n152 B 0.015806f
C183 VTAIL.n153 B 0.008493f
C184 VTAIL.n154 B 0.008493f
C185 VTAIL.n155 B 0.008993f
C186 VTAIL.n156 B 0.020075f
C187 VTAIL.n157 B 0.020075f
C188 VTAIL.n158 B 0.020075f
C189 VTAIL.n159 B 0.008743f
C190 VTAIL.n160 B 0.008493f
C191 VTAIL.n161 B 0.015806f
C192 VTAIL.n162 B 0.015806f
C193 VTAIL.n163 B 0.008493f
C194 VTAIL.n164 B 0.008993f
C195 VTAIL.n165 B 0.020075f
C196 VTAIL.n166 B 0.039687f
C197 VTAIL.n167 B 0.008993f
C198 VTAIL.n168 B 0.008493f
C199 VTAIL.n169 B 0.03567f
C200 VTAIL.n170 B 0.021792f
C201 VTAIL.n171 B 0.167335f
C202 VTAIL.n172 B 0.020083f
C203 VTAIL.n173 B 0.015806f
C204 VTAIL.n174 B 0.008493f
C205 VTAIL.n175 B 0.020075f
C206 VTAIL.n176 B 0.008743f
C207 VTAIL.n177 B 0.015806f
C208 VTAIL.n178 B 0.008993f
C209 VTAIL.n179 B 0.020075f
C210 VTAIL.n180 B 0.008993f
C211 VTAIL.n181 B 0.015806f
C212 VTAIL.n182 B 0.008493f
C213 VTAIL.n183 B 0.020075f
C214 VTAIL.n184 B 0.008993f
C215 VTAIL.n185 B 0.015806f
C216 VTAIL.n186 B 0.008493f
C217 VTAIL.n187 B 0.020075f
C218 VTAIL.n188 B 0.008993f
C219 VTAIL.n189 B 0.015806f
C220 VTAIL.n190 B 0.008493f
C221 VTAIL.n191 B 0.020075f
C222 VTAIL.n192 B 0.008993f
C223 VTAIL.n193 B 0.015806f
C224 VTAIL.n194 B 0.008493f
C225 VTAIL.n195 B 0.020075f
C226 VTAIL.n196 B 0.008993f
C227 VTAIL.n197 B 1.05151f
C228 VTAIL.n198 B 0.008493f
C229 VTAIL.t7 B 0.033118f
C230 VTAIL.n199 B 0.104355f
C231 VTAIL.n200 B 0.011859f
C232 VTAIL.n201 B 0.015056f
C233 VTAIL.n202 B 0.020075f
C234 VTAIL.n203 B 0.008993f
C235 VTAIL.n204 B 0.008493f
C236 VTAIL.n205 B 0.015806f
C237 VTAIL.n206 B 0.015806f
C238 VTAIL.n207 B 0.008493f
C239 VTAIL.n208 B 0.008993f
C240 VTAIL.n209 B 0.020075f
C241 VTAIL.n210 B 0.020075f
C242 VTAIL.n211 B 0.008993f
C243 VTAIL.n212 B 0.008493f
C244 VTAIL.n213 B 0.015806f
C245 VTAIL.n214 B 0.015806f
C246 VTAIL.n215 B 0.008493f
C247 VTAIL.n216 B 0.008993f
C248 VTAIL.n217 B 0.020075f
C249 VTAIL.n218 B 0.020075f
C250 VTAIL.n219 B 0.008993f
C251 VTAIL.n220 B 0.008493f
C252 VTAIL.n221 B 0.015806f
C253 VTAIL.n222 B 0.015806f
C254 VTAIL.n223 B 0.008493f
C255 VTAIL.n224 B 0.008993f
C256 VTAIL.n225 B 0.020075f
C257 VTAIL.n226 B 0.020075f
C258 VTAIL.n227 B 0.008993f
C259 VTAIL.n228 B 0.008493f
C260 VTAIL.n229 B 0.015806f
C261 VTAIL.n230 B 0.015806f
C262 VTAIL.n231 B 0.008493f
C263 VTAIL.n232 B 0.008993f
C264 VTAIL.n233 B 0.020075f
C265 VTAIL.n234 B 0.020075f
C266 VTAIL.n235 B 0.008993f
C267 VTAIL.n236 B 0.008493f
C268 VTAIL.n237 B 0.015806f
C269 VTAIL.n238 B 0.015806f
C270 VTAIL.n239 B 0.008493f
C271 VTAIL.n240 B 0.008493f
C272 VTAIL.n241 B 0.008993f
C273 VTAIL.n242 B 0.020075f
C274 VTAIL.n243 B 0.020075f
C275 VTAIL.n244 B 0.020075f
C276 VTAIL.n245 B 0.008743f
C277 VTAIL.n246 B 0.008493f
C278 VTAIL.n247 B 0.015806f
C279 VTAIL.n248 B 0.015806f
C280 VTAIL.n249 B 0.008493f
C281 VTAIL.n250 B 0.008993f
C282 VTAIL.n251 B 0.020075f
C283 VTAIL.n252 B 0.039687f
C284 VTAIL.n253 B 0.008993f
C285 VTAIL.n254 B 0.008493f
C286 VTAIL.n255 B 0.03567f
C287 VTAIL.n256 B 0.021792f
C288 VTAIL.n257 B 1.16112f
C289 VTAIL.n258 B 0.020083f
C290 VTAIL.n259 B 0.015806f
C291 VTAIL.n260 B 0.008493f
C292 VTAIL.n261 B 0.020075f
C293 VTAIL.n262 B 0.008743f
C294 VTAIL.n263 B 0.015806f
C295 VTAIL.n264 B 0.008743f
C296 VTAIL.n265 B 0.008493f
C297 VTAIL.n266 B 0.020075f
C298 VTAIL.n267 B 0.020075f
C299 VTAIL.n268 B 0.008993f
C300 VTAIL.n269 B 0.015806f
C301 VTAIL.n270 B 0.008493f
C302 VTAIL.n271 B 0.020075f
C303 VTAIL.n272 B 0.008993f
C304 VTAIL.n273 B 0.015806f
C305 VTAIL.n274 B 0.008493f
C306 VTAIL.n275 B 0.020075f
C307 VTAIL.n276 B 0.008993f
C308 VTAIL.n277 B 0.015806f
C309 VTAIL.n278 B 0.008493f
C310 VTAIL.n279 B 0.020075f
C311 VTAIL.n280 B 0.008993f
C312 VTAIL.n281 B 0.015806f
C313 VTAIL.n282 B 0.008493f
C314 VTAIL.n283 B 0.020075f
C315 VTAIL.n284 B 0.008993f
C316 VTAIL.n285 B 1.05151f
C317 VTAIL.n286 B 0.008493f
C318 VTAIL.t2 B 0.033118f
C319 VTAIL.n287 B 0.104355f
C320 VTAIL.n288 B 0.011859f
C321 VTAIL.n289 B 0.015056f
C322 VTAIL.n290 B 0.020075f
C323 VTAIL.n291 B 0.008993f
C324 VTAIL.n292 B 0.008493f
C325 VTAIL.n293 B 0.015806f
C326 VTAIL.n294 B 0.015806f
C327 VTAIL.n295 B 0.008493f
C328 VTAIL.n296 B 0.008993f
C329 VTAIL.n297 B 0.020075f
C330 VTAIL.n298 B 0.020075f
C331 VTAIL.n299 B 0.008993f
C332 VTAIL.n300 B 0.008493f
C333 VTAIL.n301 B 0.015806f
C334 VTAIL.n302 B 0.015806f
C335 VTAIL.n303 B 0.008493f
C336 VTAIL.n304 B 0.008993f
C337 VTAIL.n305 B 0.020075f
C338 VTAIL.n306 B 0.020075f
C339 VTAIL.n307 B 0.008993f
C340 VTAIL.n308 B 0.008493f
C341 VTAIL.n309 B 0.015806f
C342 VTAIL.n310 B 0.015806f
C343 VTAIL.n311 B 0.008493f
C344 VTAIL.n312 B 0.008993f
C345 VTAIL.n313 B 0.020075f
C346 VTAIL.n314 B 0.020075f
C347 VTAIL.n315 B 0.008993f
C348 VTAIL.n316 B 0.008493f
C349 VTAIL.n317 B 0.015806f
C350 VTAIL.n318 B 0.015806f
C351 VTAIL.n319 B 0.008493f
C352 VTAIL.n320 B 0.008993f
C353 VTAIL.n321 B 0.020075f
C354 VTAIL.n322 B 0.020075f
C355 VTAIL.n323 B 0.008993f
C356 VTAIL.n324 B 0.008493f
C357 VTAIL.n325 B 0.015806f
C358 VTAIL.n326 B 0.015806f
C359 VTAIL.n327 B 0.008493f
C360 VTAIL.n328 B 0.008993f
C361 VTAIL.n329 B 0.020075f
C362 VTAIL.n330 B 0.020075f
C363 VTAIL.n331 B 0.008993f
C364 VTAIL.n332 B 0.008493f
C365 VTAIL.n333 B 0.015806f
C366 VTAIL.n334 B 0.015806f
C367 VTAIL.n335 B 0.008493f
C368 VTAIL.n336 B 0.008993f
C369 VTAIL.n337 B 0.020075f
C370 VTAIL.n338 B 0.039687f
C371 VTAIL.n339 B 0.008993f
C372 VTAIL.n340 B 0.008493f
C373 VTAIL.n341 B 0.03567f
C374 VTAIL.n342 B 0.021792f
C375 VTAIL.n343 B 1.16112f
C376 VTAIL.n344 B 0.020083f
C377 VTAIL.n345 B 0.015806f
C378 VTAIL.n346 B 0.008493f
C379 VTAIL.n347 B 0.020075f
C380 VTAIL.n348 B 0.008743f
C381 VTAIL.n349 B 0.015806f
C382 VTAIL.n350 B 0.008743f
C383 VTAIL.n351 B 0.008493f
C384 VTAIL.n352 B 0.020075f
C385 VTAIL.n353 B 0.020075f
C386 VTAIL.n354 B 0.008993f
C387 VTAIL.n355 B 0.015806f
C388 VTAIL.n356 B 0.008493f
C389 VTAIL.n357 B 0.020075f
C390 VTAIL.n358 B 0.008993f
C391 VTAIL.n359 B 0.015806f
C392 VTAIL.n360 B 0.008493f
C393 VTAIL.n361 B 0.020075f
C394 VTAIL.n362 B 0.008993f
C395 VTAIL.n363 B 0.015806f
C396 VTAIL.n364 B 0.008493f
C397 VTAIL.n365 B 0.020075f
C398 VTAIL.n366 B 0.008993f
C399 VTAIL.n367 B 0.015806f
C400 VTAIL.n368 B 0.008493f
C401 VTAIL.n369 B 0.020075f
C402 VTAIL.n370 B 0.008993f
C403 VTAIL.n371 B 1.05151f
C404 VTAIL.n372 B 0.008493f
C405 VTAIL.t3 B 0.033118f
C406 VTAIL.n373 B 0.104355f
C407 VTAIL.n374 B 0.011859f
C408 VTAIL.n375 B 0.015056f
C409 VTAIL.n376 B 0.020075f
C410 VTAIL.n377 B 0.008993f
C411 VTAIL.n378 B 0.008493f
C412 VTAIL.n379 B 0.015806f
C413 VTAIL.n380 B 0.015806f
C414 VTAIL.n381 B 0.008493f
C415 VTAIL.n382 B 0.008993f
C416 VTAIL.n383 B 0.020075f
C417 VTAIL.n384 B 0.020075f
C418 VTAIL.n385 B 0.008993f
C419 VTAIL.n386 B 0.008493f
C420 VTAIL.n387 B 0.015806f
C421 VTAIL.n388 B 0.015806f
C422 VTAIL.n389 B 0.008493f
C423 VTAIL.n390 B 0.008993f
C424 VTAIL.n391 B 0.020075f
C425 VTAIL.n392 B 0.020075f
C426 VTAIL.n393 B 0.008993f
C427 VTAIL.n394 B 0.008493f
C428 VTAIL.n395 B 0.015806f
C429 VTAIL.n396 B 0.015806f
C430 VTAIL.n397 B 0.008493f
C431 VTAIL.n398 B 0.008993f
C432 VTAIL.n399 B 0.020075f
C433 VTAIL.n400 B 0.020075f
C434 VTAIL.n401 B 0.008993f
C435 VTAIL.n402 B 0.008493f
C436 VTAIL.n403 B 0.015806f
C437 VTAIL.n404 B 0.015806f
C438 VTAIL.n405 B 0.008493f
C439 VTAIL.n406 B 0.008993f
C440 VTAIL.n407 B 0.020075f
C441 VTAIL.n408 B 0.020075f
C442 VTAIL.n409 B 0.008993f
C443 VTAIL.n410 B 0.008493f
C444 VTAIL.n411 B 0.015806f
C445 VTAIL.n412 B 0.015806f
C446 VTAIL.n413 B 0.008493f
C447 VTAIL.n414 B 0.008993f
C448 VTAIL.n415 B 0.020075f
C449 VTAIL.n416 B 0.020075f
C450 VTAIL.n417 B 0.008993f
C451 VTAIL.n418 B 0.008493f
C452 VTAIL.n419 B 0.015806f
C453 VTAIL.n420 B 0.015806f
C454 VTAIL.n421 B 0.008493f
C455 VTAIL.n422 B 0.008993f
C456 VTAIL.n423 B 0.020075f
C457 VTAIL.n424 B 0.039687f
C458 VTAIL.n425 B 0.008993f
C459 VTAIL.n426 B 0.008493f
C460 VTAIL.n427 B 0.03567f
C461 VTAIL.n428 B 0.021792f
C462 VTAIL.n429 B 0.167335f
C463 VTAIL.n430 B 0.020083f
C464 VTAIL.n431 B 0.015806f
C465 VTAIL.n432 B 0.008493f
C466 VTAIL.n433 B 0.020075f
C467 VTAIL.n434 B 0.008743f
C468 VTAIL.n435 B 0.015806f
C469 VTAIL.n436 B 0.008743f
C470 VTAIL.n437 B 0.008493f
C471 VTAIL.n438 B 0.020075f
C472 VTAIL.n439 B 0.020075f
C473 VTAIL.n440 B 0.008993f
C474 VTAIL.n441 B 0.015806f
C475 VTAIL.n442 B 0.008493f
C476 VTAIL.n443 B 0.020075f
C477 VTAIL.n444 B 0.008993f
C478 VTAIL.n445 B 0.015806f
C479 VTAIL.n446 B 0.008493f
C480 VTAIL.n447 B 0.020075f
C481 VTAIL.n448 B 0.008993f
C482 VTAIL.n449 B 0.015806f
C483 VTAIL.n450 B 0.008493f
C484 VTAIL.n451 B 0.020075f
C485 VTAIL.n452 B 0.008993f
C486 VTAIL.n453 B 0.015806f
C487 VTAIL.n454 B 0.008493f
C488 VTAIL.n455 B 0.020075f
C489 VTAIL.n456 B 0.008993f
C490 VTAIL.n457 B 1.05151f
C491 VTAIL.n458 B 0.008493f
C492 VTAIL.t5 B 0.033118f
C493 VTAIL.n459 B 0.104355f
C494 VTAIL.n460 B 0.011859f
C495 VTAIL.n461 B 0.015056f
C496 VTAIL.n462 B 0.020075f
C497 VTAIL.n463 B 0.008993f
C498 VTAIL.n464 B 0.008493f
C499 VTAIL.n465 B 0.015806f
C500 VTAIL.n466 B 0.015806f
C501 VTAIL.n467 B 0.008493f
C502 VTAIL.n468 B 0.008993f
C503 VTAIL.n469 B 0.020075f
C504 VTAIL.n470 B 0.020075f
C505 VTAIL.n471 B 0.008993f
C506 VTAIL.n472 B 0.008493f
C507 VTAIL.n473 B 0.015806f
C508 VTAIL.n474 B 0.015806f
C509 VTAIL.n475 B 0.008493f
C510 VTAIL.n476 B 0.008993f
C511 VTAIL.n477 B 0.020075f
C512 VTAIL.n478 B 0.020075f
C513 VTAIL.n479 B 0.008993f
C514 VTAIL.n480 B 0.008493f
C515 VTAIL.n481 B 0.015806f
C516 VTAIL.n482 B 0.015806f
C517 VTAIL.n483 B 0.008493f
C518 VTAIL.n484 B 0.008993f
C519 VTAIL.n485 B 0.020075f
C520 VTAIL.n486 B 0.020075f
C521 VTAIL.n487 B 0.008993f
C522 VTAIL.n488 B 0.008493f
C523 VTAIL.n489 B 0.015806f
C524 VTAIL.n490 B 0.015806f
C525 VTAIL.n491 B 0.008493f
C526 VTAIL.n492 B 0.008993f
C527 VTAIL.n493 B 0.020075f
C528 VTAIL.n494 B 0.020075f
C529 VTAIL.n495 B 0.008993f
C530 VTAIL.n496 B 0.008493f
C531 VTAIL.n497 B 0.015806f
C532 VTAIL.n498 B 0.015806f
C533 VTAIL.n499 B 0.008493f
C534 VTAIL.n500 B 0.008993f
C535 VTAIL.n501 B 0.020075f
C536 VTAIL.n502 B 0.020075f
C537 VTAIL.n503 B 0.008993f
C538 VTAIL.n504 B 0.008493f
C539 VTAIL.n505 B 0.015806f
C540 VTAIL.n506 B 0.015806f
C541 VTAIL.n507 B 0.008493f
C542 VTAIL.n508 B 0.008993f
C543 VTAIL.n509 B 0.020075f
C544 VTAIL.n510 B 0.039687f
C545 VTAIL.n511 B 0.008993f
C546 VTAIL.n512 B 0.008493f
C547 VTAIL.n513 B 0.03567f
C548 VTAIL.n514 B 0.021792f
C549 VTAIL.n515 B 0.167335f
C550 VTAIL.n516 B 0.020083f
C551 VTAIL.n517 B 0.015806f
C552 VTAIL.n518 B 0.008493f
C553 VTAIL.n519 B 0.020075f
C554 VTAIL.n520 B 0.008743f
C555 VTAIL.n521 B 0.015806f
C556 VTAIL.n522 B 0.008743f
C557 VTAIL.n523 B 0.008493f
C558 VTAIL.n524 B 0.020075f
C559 VTAIL.n525 B 0.020075f
C560 VTAIL.n526 B 0.008993f
C561 VTAIL.n527 B 0.015806f
C562 VTAIL.n528 B 0.008493f
C563 VTAIL.n529 B 0.020075f
C564 VTAIL.n530 B 0.008993f
C565 VTAIL.n531 B 0.015806f
C566 VTAIL.n532 B 0.008493f
C567 VTAIL.n533 B 0.020075f
C568 VTAIL.n534 B 0.008993f
C569 VTAIL.n535 B 0.015806f
C570 VTAIL.n536 B 0.008493f
C571 VTAIL.n537 B 0.020075f
C572 VTAIL.n538 B 0.008993f
C573 VTAIL.n539 B 0.015806f
C574 VTAIL.n540 B 0.008493f
C575 VTAIL.n541 B 0.020075f
C576 VTAIL.n542 B 0.008993f
C577 VTAIL.n543 B 1.05151f
C578 VTAIL.n544 B 0.008493f
C579 VTAIL.t4 B 0.033118f
C580 VTAIL.n545 B 0.104355f
C581 VTAIL.n546 B 0.011859f
C582 VTAIL.n547 B 0.015056f
C583 VTAIL.n548 B 0.020075f
C584 VTAIL.n549 B 0.008993f
C585 VTAIL.n550 B 0.008493f
C586 VTAIL.n551 B 0.015806f
C587 VTAIL.n552 B 0.015806f
C588 VTAIL.n553 B 0.008493f
C589 VTAIL.n554 B 0.008993f
C590 VTAIL.n555 B 0.020075f
C591 VTAIL.n556 B 0.020075f
C592 VTAIL.n557 B 0.008993f
C593 VTAIL.n558 B 0.008493f
C594 VTAIL.n559 B 0.015806f
C595 VTAIL.n560 B 0.015806f
C596 VTAIL.n561 B 0.008493f
C597 VTAIL.n562 B 0.008993f
C598 VTAIL.n563 B 0.020075f
C599 VTAIL.n564 B 0.020075f
C600 VTAIL.n565 B 0.008993f
C601 VTAIL.n566 B 0.008493f
C602 VTAIL.n567 B 0.015806f
C603 VTAIL.n568 B 0.015806f
C604 VTAIL.n569 B 0.008493f
C605 VTAIL.n570 B 0.008993f
C606 VTAIL.n571 B 0.020075f
C607 VTAIL.n572 B 0.020075f
C608 VTAIL.n573 B 0.008993f
C609 VTAIL.n574 B 0.008493f
C610 VTAIL.n575 B 0.015806f
C611 VTAIL.n576 B 0.015806f
C612 VTAIL.n577 B 0.008493f
C613 VTAIL.n578 B 0.008993f
C614 VTAIL.n579 B 0.020075f
C615 VTAIL.n580 B 0.020075f
C616 VTAIL.n581 B 0.008993f
C617 VTAIL.n582 B 0.008493f
C618 VTAIL.n583 B 0.015806f
C619 VTAIL.n584 B 0.015806f
C620 VTAIL.n585 B 0.008493f
C621 VTAIL.n586 B 0.008993f
C622 VTAIL.n587 B 0.020075f
C623 VTAIL.n588 B 0.020075f
C624 VTAIL.n589 B 0.008993f
C625 VTAIL.n590 B 0.008493f
C626 VTAIL.n591 B 0.015806f
C627 VTAIL.n592 B 0.015806f
C628 VTAIL.n593 B 0.008493f
C629 VTAIL.n594 B 0.008993f
C630 VTAIL.n595 B 0.020075f
C631 VTAIL.n596 B 0.039687f
C632 VTAIL.n597 B 0.008993f
C633 VTAIL.n598 B 0.008493f
C634 VTAIL.n599 B 0.03567f
C635 VTAIL.n600 B 0.021792f
C636 VTAIL.n601 B 1.16112f
C637 VTAIL.n602 B 0.020083f
C638 VTAIL.n603 B 0.015806f
C639 VTAIL.n604 B 0.008493f
C640 VTAIL.n605 B 0.020075f
C641 VTAIL.n606 B 0.008743f
C642 VTAIL.n607 B 0.015806f
C643 VTAIL.n608 B 0.008993f
C644 VTAIL.n609 B 0.020075f
C645 VTAIL.n610 B 0.008993f
C646 VTAIL.n611 B 0.015806f
C647 VTAIL.n612 B 0.008493f
C648 VTAIL.n613 B 0.020075f
C649 VTAIL.n614 B 0.008993f
C650 VTAIL.n615 B 0.015806f
C651 VTAIL.n616 B 0.008493f
C652 VTAIL.n617 B 0.020075f
C653 VTAIL.n618 B 0.008993f
C654 VTAIL.n619 B 0.015806f
C655 VTAIL.n620 B 0.008493f
C656 VTAIL.n621 B 0.020075f
C657 VTAIL.n622 B 0.008993f
C658 VTAIL.n623 B 0.015806f
C659 VTAIL.n624 B 0.008493f
C660 VTAIL.n625 B 0.020075f
C661 VTAIL.n626 B 0.008993f
C662 VTAIL.n627 B 1.05151f
C663 VTAIL.n628 B 0.008493f
C664 VTAIL.t1 B 0.033118f
C665 VTAIL.n629 B 0.104355f
C666 VTAIL.n630 B 0.011859f
C667 VTAIL.n631 B 0.015056f
C668 VTAIL.n632 B 0.020075f
C669 VTAIL.n633 B 0.008993f
C670 VTAIL.n634 B 0.008493f
C671 VTAIL.n635 B 0.015806f
C672 VTAIL.n636 B 0.015806f
C673 VTAIL.n637 B 0.008493f
C674 VTAIL.n638 B 0.008993f
C675 VTAIL.n639 B 0.020075f
C676 VTAIL.n640 B 0.020075f
C677 VTAIL.n641 B 0.008993f
C678 VTAIL.n642 B 0.008493f
C679 VTAIL.n643 B 0.015806f
C680 VTAIL.n644 B 0.015806f
C681 VTAIL.n645 B 0.008493f
C682 VTAIL.n646 B 0.008993f
C683 VTAIL.n647 B 0.020075f
C684 VTAIL.n648 B 0.020075f
C685 VTAIL.n649 B 0.008993f
C686 VTAIL.n650 B 0.008493f
C687 VTAIL.n651 B 0.015806f
C688 VTAIL.n652 B 0.015806f
C689 VTAIL.n653 B 0.008493f
C690 VTAIL.n654 B 0.008993f
C691 VTAIL.n655 B 0.020075f
C692 VTAIL.n656 B 0.020075f
C693 VTAIL.n657 B 0.008993f
C694 VTAIL.n658 B 0.008493f
C695 VTAIL.n659 B 0.015806f
C696 VTAIL.n660 B 0.015806f
C697 VTAIL.n661 B 0.008493f
C698 VTAIL.n662 B 0.008993f
C699 VTAIL.n663 B 0.020075f
C700 VTAIL.n664 B 0.020075f
C701 VTAIL.n665 B 0.008993f
C702 VTAIL.n666 B 0.008493f
C703 VTAIL.n667 B 0.015806f
C704 VTAIL.n668 B 0.015806f
C705 VTAIL.n669 B 0.008493f
C706 VTAIL.n670 B 0.008493f
C707 VTAIL.n671 B 0.008993f
C708 VTAIL.n672 B 0.020075f
C709 VTAIL.n673 B 0.020075f
C710 VTAIL.n674 B 0.020075f
C711 VTAIL.n675 B 0.008743f
C712 VTAIL.n676 B 0.008493f
C713 VTAIL.n677 B 0.015806f
C714 VTAIL.n678 B 0.015806f
C715 VTAIL.n679 B 0.008493f
C716 VTAIL.n680 B 0.008993f
C717 VTAIL.n681 B 0.020075f
C718 VTAIL.n682 B 0.039687f
C719 VTAIL.n683 B 0.008993f
C720 VTAIL.n684 B 0.008493f
C721 VTAIL.n685 B 0.03567f
C722 VTAIL.n686 B 0.021792f
C723 VTAIL.n687 B 1.09295f
C724 VDD1.t2 B 0.323801f
C725 VDD1.t1 B 0.323801f
C726 VDD1.n0 B 2.92901f
C727 VDD1.t3 B 0.323801f
C728 VDD1.t0 B 0.323801f
C729 VDD1.n1 B 3.7637f
C730 VP.n0 B 0.032638f
C731 VP.t1 B 2.74506f
C732 VP.n1 B 0.035988f
C733 VP.n2 B 0.024757f
C734 VP.t0 B 2.74506f
C735 VP.n3 B 1.04412f
C736 VP.t3 B 2.97246f
C737 VP.t2 B 2.97729f
C738 VP.n4 B 3.32118f
C739 VP.n5 B 1.48114f
C740 VP.n6 B 0.032638f
C741 VP.n7 B 0.033898f
C742 VP.n8 B 0.04591f
C743 VP.n9 B 0.035988f
C744 VP.n10 B 0.024757f
C745 VP.n11 B 0.024757f
C746 VP.n12 B 0.024757f
C747 VP.n13 B 0.04591f
C748 VP.n14 B 0.033898f
C749 VP.n15 B 1.04412f
C750 VP.n16 B 0.039541f
.ends

