* NGSPICE file created from diff_pair_sample_0592.ext - technology: sky130A

.subckt diff_pair_sample_0592 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t4 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=0.93555 pd=6 as=2.2113 ps=12.12 w=5.67 l=1.89
X1 B.t11 B.t9 B.t10 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=2.2113 pd=12.12 as=0 ps=0 w=5.67 l=1.89
X2 VDD1.t4 VP.t1 VTAIL.t3 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=2.2113 pd=12.12 as=0.93555 ps=6 w=5.67 l=1.89
X3 B.t8 B.t6 B.t7 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=2.2113 pd=12.12 as=0 ps=0 w=5.67 l=1.89
X4 VDD2.t5 VN.t0 VTAIL.t2 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=0.93555 pd=6 as=2.2113 ps=12.12 w=5.67 l=1.89
X5 VDD2.t4 VN.t1 VTAIL.t1 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=2.2113 pd=12.12 as=0.93555 ps=6 w=5.67 l=1.89
X6 VDD2.t3 VN.t2 VTAIL.t0 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=0.93555 pd=6 as=2.2113 ps=12.12 w=5.67 l=1.89
X7 VDD1.t3 VP.t2 VTAIL.t6 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=0.93555 pd=6 as=2.2113 ps=12.12 w=5.67 l=1.89
X8 VTAIL.t9 VN.t3 VDD2.t2 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=0.93555 pd=6 as=0.93555 ps=6 w=5.67 l=1.89
X9 VTAIL.t8 VP.t3 VDD1.t2 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=0.93555 pd=6 as=0.93555 ps=6 w=5.67 l=1.89
X10 B.t5 B.t3 B.t4 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=2.2113 pd=12.12 as=0 ps=0 w=5.67 l=1.89
X11 VDD2.t1 VN.t4 VTAIL.t11 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=2.2113 pd=12.12 as=0.93555 ps=6 w=5.67 l=1.89
X12 VTAIL.t7 VP.t4 VDD1.t1 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=0.93555 pd=6 as=0.93555 ps=6 w=5.67 l=1.89
X13 B.t2 B.t0 B.t1 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=2.2113 pd=12.12 as=0 ps=0 w=5.67 l=1.89
X14 VTAIL.t10 VN.t5 VDD2.t0 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=0.93555 pd=6 as=0.93555 ps=6 w=5.67 l=1.89
X15 VDD1.t0 VP.t5 VTAIL.t5 w_n2746_n2102# sky130_fd_pr__pfet_01v8 ad=2.2113 pd=12.12 as=0.93555 ps=6 w=5.67 l=1.89
R0 VP.n9 VP.n8 161.3
R1 VP.n10 VP.n5 161.3
R2 VP.n12 VP.n11 161.3
R3 VP.n13 VP.n4 161.3
R4 VP.n30 VP.n0 161.3
R5 VP.n29 VP.n28 161.3
R6 VP.n27 VP.n1 161.3
R7 VP.n26 VP.n25 161.3
R8 VP.n23 VP.n2 161.3
R9 VP.n22 VP.n21 161.3
R10 VP.n20 VP.n3 161.3
R11 VP.n19 VP.n18 161.3
R12 VP.n6 VP.t1 103.392
R13 VP.n17 VP.n16 87.7575
R14 VP.n32 VP.n31 87.7575
R15 VP.n15 VP.n14 87.7575
R16 VP.n17 VP.t5 72.3005
R17 VP.n24 VP.t3 72.3005
R18 VP.n31 VP.t0 72.3005
R19 VP.n14 VP.t2 72.3005
R20 VP.n7 VP.t4 72.3005
R21 VP.n7 VP.n6 57.8248
R22 VP.n22 VP.n3 54.0911
R23 VP.n29 VP.n1 54.0911
R24 VP.n12 VP.n5 54.0911
R25 VP.n16 VP.n15 41.1435
R26 VP.n18 VP.n3 26.8957
R27 VP.n30 VP.n29 26.8957
R28 VP.n13 VP.n12 26.8957
R29 VP.n23 VP.n22 24.4675
R30 VP.n25 VP.n1 24.4675
R31 VP.n8 VP.n5 24.4675
R32 VP.n18 VP.n17 22.9995
R33 VP.n31 VP.n30 22.9995
R34 VP.n14 VP.n13 22.9995
R35 VP.n9 VP.n6 12.851
R36 VP.n24 VP.n23 12.234
R37 VP.n25 VP.n24 12.234
R38 VP.n8 VP.n7 12.234
R39 VP.n15 VP.n4 0.278367
R40 VP.n19 VP.n16 0.278367
R41 VP.n32 VP.n0 0.278367
R42 VP.n10 VP.n9 0.189894
R43 VP.n11 VP.n10 0.189894
R44 VP.n11 VP.n4 0.189894
R45 VP.n20 VP.n19 0.189894
R46 VP.n21 VP.n20 0.189894
R47 VP.n21 VP.n2 0.189894
R48 VP.n26 VP.n2 0.189894
R49 VP.n27 VP.n26 0.189894
R50 VP.n28 VP.n27 0.189894
R51 VP.n28 VP.n0 0.189894
R52 VP VP.n32 0.153454
R53 VTAIL.n7 VTAIL.t0 84.2763
R54 VTAIL.n11 VTAIL.t2 84.2761
R55 VTAIL.n2 VTAIL.t4 84.2761
R56 VTAIL.n10 VTAIL.t6 84.2761
R57 VTAIL.n9 VTAIL.n8 78.5435
R58 VTAIL.n6 VTAIL.n5 78.5435
R59 VTAIL.n1 VTAIL.n0 78.5433
R60 VTAIL.n4 VTAIL.n3 78.5433
R61 VTAIL.n6 VTAIL.n4 21.0824
R62 VTAIL.n11 VTAIL.n10 19.1686
R63 VTAIL.n0 VTAIL.t1 5.7333
R64 VTAIL.n0 VTAIL.t9 5.7333
R65 VTAIL.n3 VTAIL.t5 5.7333
R66 VTAIL.n3 VTAIL.t8 5.7333
R67 VTAIL.n8 VTAIL.t3 5.7333
R68 VTAIL.n8 VTAIL.t7 5.7333
R69 VTAIL.n5 VTAIL.t11 5.7333
R70 VTAIL.n5 VTAIL.t10 5.7333
R71 VTAIL.n7 VTAIL.n6 1.91429
R72 VTAIL.n10 VTAIL.n9 1.91429
R73 VTAIL.n4 VTAIL.n2 1.91429
R74 VTAIL.n9 VTAIL.n7 1.42722
R75 VTAIL.n2 VTAIL.n1 1.42722
R76 VTAIL VTAIL.n11 1.37766
R77 VTAIL VTAIL.n1 0.537138
R78 VDD1 VDD1.t4 102.448
R79 VDD1.n1 VDD1.t0 102.335
R80 VDD1.n1 VDD1.n0 95.6452
R81 VDD1.n3 VDD1.n2 95.2222
R82 VDD1.n3 VDD1.n1 36.363
R83 VDD1.n2 VDD1.t1 5.7333
R84 VDD1.n2 VDD1.t3 5.7333
R85 VDD1.n0 VDD1.t2 5.7333
R86 VDD1.n0 VDD1.t5 5.7333
R87 VDD1 VDD1.n3 0.420759
R88 B.n375 B.n374 585
R89 B.n376 B.n51 585
R90 B.n378 B.n377 585
R91 B.n379 B.n50 585
R92 B.n381 B.n380 585
R93 B.n382 B.n49 585
R94 B.n384 B.n383 585
R95 B.n385 B.n48 585
R96 B.n387 B.n386 585
R97 B.n388 B.n47 585
R98 B.n390 B.n389 585
R99 B.n391 B.n46 585
R100 B.n393 B.n392 585
R101 B.n394 B.n45 585
R102 B.n396 B.n395 585
R103 B.n397 B.n44 585
R104 B.n399 B.n398 585
R105 B.n400 B.n43 585
R106 B.n402 B.n401 585
R107 B.n403 B.n42 585
R108 B.n405 B.n404 585
R109 B.n406 B.n41 585
R110 B.n408 B.n407 585
R111 B.n410 B.n38 585
R112 B.n412 B.n411 585
R113 B.n413 B.n37 585
R114 B.n415 B.n414 585
R115 B.n416 B.n36 585
R116 B.n418 B.n417 585
R117 B.n419 B.n35 585
R118 B.n421 B.n420 585
R119 B.n422 B.n31 585
R120 B.n424 B.n423 585
R121 B.n425 B.n30 585
R122 B.n427 B.n426 585
R123 B.n428 B.n29 585
R124 B.n430 B.n429 585
R125 B.n431 B.n28 585
R126 B.n433 B.n432 585
R127 B.n434 B.n27 585
R128 B.n436 B.n435 585
R129 B.n437 B.n26 585
R130 B.n439 B.n438 585
R131 B.n440 B.n25 585
R132 B.n442 B.n441 585
R133 B.n443 B.n24 585
R134 B.n445 B.n444 585
R135 B.n446 B.n23 585
R136 B.n448 B.n447 585
R137 B.n449 B.n22 585
R138 B.n451 B.n450 585
R139 B.n452 B.n21 585
R140 B.n454 B.n453 585
R141 B.n455 B.n20 585
R142 B.n457 B.n456 585
R143 B.n458 B.n19 585
R144 B.n373 B.n52 585
R145 B.n372 B.n371 585
R146 B.n370 B.n53 585
R147 B.n369 B.n368 585
R148 B.n367 B.n54 585
R149 B.n366 B.n365 585
R150 B.n364 B.n55 585
R151 B.n363 B.n362 585
R152 B.n361 B.n56 585
R153 B.n360 B.n359 585
R154 B.n358 B.n57 585
R155 B.n357 B.n356 585
R156 B.n355 B.n58 585
R157 B.n354 B.n353 585
R158 B.n352 B.n59 585
R159 B.n351 B.n350 585
R160 B.n349 B.n60 585
R161 B.n348 B.n347 585
R162 B.n346 B.n61 585
R163 B.n345 B.n344 585
R164 B.n343 B.n62 585
R165 B.n342 B.n341 585
R166 B.n340 B.n63 585
R167 B.n339 B.n338 585
R168 B.n337 B.n64 585
R169 B.n336 B.n335 585
R170 B.n334 B.n65 585
R171 B.n333 B.n332 585
R172 B.n331 B.n66 585
R173 B.n330 B.n329 585
R174 B.n328 B.n67 585
R175 B.n327 B.n326 585
R176 B.n325 B.n68 585
R177 B.n324 B.n323 585
R178 B.n322 B.n69 585
R179 B.n321 B.n320 585
R180 B.n319 B.n70 585
R181 B.n318 B.n317 585
R182 B.n316 B.n71 585
R183 B.n315 B.n314 585
R184 B.n313 B.n72 585
R185 B.n312 B.n311 585
R186 B.n310 B.n73 585
R187 B.n309 B.n308 585
R188 B.n307 B.n74 585
R189 B.n306 B.n305 585
R190 B.n304 B.n75 585
R191 B.n303 B.n302 585
R192 B.n301 B.n76 585
R193 B.n300 B.n299 585
R194 B.n298 B.n77 585
R195 B.n297 B.n296 585
R196 B.n295 B.n78 585
R197 B.n294 B.n293 585
R198 B.n292 B.n79 585
R199 B.n291 B.n290 585
R200 B.n289 B.n80 585
R201 B.n288 B.n287 585
R202 B.n286 B.n81 585
R203 B.n285 B.n284 585
R204 B.n283 B.n82 585
R205 B.n282 B.n281 585
R206 B.n280 B.n83 585
R207 B.n279 B.n278 585
R208 B.n277 B.n84 585
R209 B.n276 B.n275 585
R210 B.n274 B.n85 585
R211 B.n273 B.n272 585
R212 B.n271 B.n86 585
R213 B.n186 B.n185 585
R214 B.n187 B.n118 585
R215 B.n189 B.n188 585
R216 B.n190 B.n117 585
R217 B.n192 B.n191 585
R218 B.n193 B.n116 585
R219 B.n195 B.n194 585
R220 B.n196 B.n115 585
R221 B.n198 B.n197 585
R222 B.n199 B.n114 585
R223 B.n201 B.n200 585
R224 B.n202 B.n113 585
R225 B.n204 B.n203 585
R226 B.n205 B.n112 585
R227 B.n207 B.n206 585
R228 B.n208 B.n111 585
R229 B.n210 B.n209 585
R230 B.n211 B.n110 585
R231 B.n213 B.n212 585
R232 B.n214 B.n109 585
R233 B.n216 B.n215 585
R234 B.n217 B.n108 585
R235 B.n219 B.n218 585
R236 B.n221 B.n220 585
R237 B.n222 B.n104 585
R238 B.n224 B.n223 585
R239 B.n225 B.n103 585
R240 B.n227 B.n226 585
R241 B.n228 B.n102 585
R242 B.n230 B.n229 585
R243 B.n231 B.n101 585
R244 B.n233 B.n232 585
R245 B.n234 B.n98 585
R246 B.n237 B.n236 585
R247 B.n238 B.n97 585
R248 B.n240 B.n239 585
R249 B.n241 B.n96 585
R250 B.n243 B.n242 585
R251 B.n244 B.n95 585
R252 B.n246 B.n245 585
R253 B.n247 B.n94 585
R254 B.n249 B.n248 585
R255 B.n250 B.n93 585
R256 B.n252 B.n251 585
R257 B.n253 B.n92 585
R258 B.n255 B.n254 585
R259 B.n256 B.n91 585
R260 B.n258 B.n257 585
R261 B.n259 B.n90 585
R262 B.n261 B.n260 585
R263 B.n262 B.n89 585
R264 B.n264 B.n263 585
R265 B.n265 B.n88 585
R266 B.n267 B.n266 585
R267 B.n268 B.n87 585
R268 B.n270 B.n269 585
R269 B.n184 B.n119 585
R270 B.n183 B.n182 585
R271 B.n181 B.n120 585
R272 B.n180 B.n179 585
R273 B.n178 B.n121 585
R274 B.n177 B.n176 585
R275 B.n175 B.n122 585
R276 B.n174 B.n173 585
R277 B.n172 B.n123 585
R278 B.n171 B.n170 585
R279 B.n169 B.n124 585
R280 B.n168 B.n167 585
R281 B.n166 B.n125 585
R282 B.n165 B.n164 585
R283 B.n163 B.n126 585
R284 B.n162 B.n161 585
R285 B.n160 B.n127 585
R286 B.n159 B.n158 585
R287 B.n157 B.n128 585
R288 B.n156 B.n155 585
R289 B.n154 B.n129 585
R290 B.n153 B.n152 585
R291 B.n151 B.n130 585
R292 B.n150 B.n149 585
R293 B.n148 B.n131 585
R294 B.n147 B.n146 585
R295 B.n145 B.n132 585
R296 B.n144 B.n143 585
R297 B.n142 B.n133 585
R298 B.n141 B.n140 585
R299 B.n139 B.n134 585
R300 B.n138 B.n137 585
R301 B.n136 B.n135 585
R302 B.n2 B.n0 585
R303 B.n509 B.n1 585
R304 B.n508 B.n507 585
R305 B.n506 B.n3 585
R306 B.n505 B.n504 585
R307 B.n503 B.n4 585
R308 B.n502 B.n501 585
R309 B.n500 B.n5 585
R310 B.n499 B.n498 585
R311 B.n497 B.n6 585
R312 B.n496 B.n495 585
R313 B.n494 B.n7 585
R314 B.n493 B.n492 585
R315 B.n491 B.n8 585
R316 B.n490 B.n489 585
R317 B.n488 B.n9 585
R318 B.n487 B.n486 585
R319 B.n485 B.n10 585
R320 B.n484 B.n483 585
R321 B.n482 B.n11 585
R322 B.n481 B.n480 585
R323 B.n479 B.n12 585
R324 B.n478 B.n477 585
R325 B.n476 B.n13 585
R326 B.n475 B.n474 585
R327 B.n473 B.n14 585
R328 B.n472 B.n471 585
R329 B.n470 B.n15 585
R330 B.n469 B.n468 585
R331 B.n467 B.n16 585
R332 B.n466 B.n465 585
R333 B.n464 B.n17 585
R334 B.n463 B.n462 585
R335 B.n461 B.n18 585
R336 B.n460 B.n459 585
R337 B.n511 B.n510 585
R338 B.n185 B.n184 502.111
R339 B.n460 B.n19 502.111
R340 B.n269 B.n86 502.111
R341 B.n375 B.n52 502.111
R342 B.n99 B.t6 278.947
R343 B.n105 B.t0 278.947
R344 B.n32 B.t9 278.947
R345 B.n39 B.t3 278.947
R346 B.n184 B.n183 163.367
R347 B.n183 B.n120 163.367
R348 B.n179 B.n120 163.367
R349 B.n179 B.n178 163.367
R350 B.n178 B.n177 163.367
R351 B.n177 B.n122 163.367
R352 B.n173 B.n122 163.367
R353 B.n173 B.n172 163.367
R354 B.n172 B.n171 163.367
R355 B.n171 B.n124 163.367
R356 B.n167 B.n124 163.367
R357 B.n167 B.n166 163.367
R358 B.n166 B.n165 163.367
R359 B.n165 B.n126 163.367
R360 B.n161 B.n126 163.367
R361 B.n161 B.n160 163.367
R362 B.n160 B.n159 163.367
R363 B.n159 B.n128 163.367
R364 B.n155 B.n128 163.367
R365 B.n155 B.n154 163.367
R366 B.n154 B.n153 163.367
R367 B.n153 B.n130 163.367
R368 B.n149 B.n130 163.367
R369 B.n149 B.n148 163.367
R370 B.n148 B.n147 163.367
R371 B.n147 B.n132 163.367
R372 B.n143 B.n132 163.367
R373 B.n143 B.n142 163.367
R374 B.n142 B.n141 163.367
R375 B.n141 B.n134 163.367
R376 B.n137 B.n134 163.367
R377 B.n137 B.n136 163.367
R378 B.n136 B.n2 163.367
R379 B.n510 B.n2 163.367
R380 B.n510 B.n509 163.367
R381 B.n509 B.n508 163.367
R382 B.n508 B.n3 163.367
R383 B.n504 B.n3 163.367
R384 B.n504 B.n503 163.367
R385 B.n503 B.n502 163.367
R386 B.n502 B.n5 163.367
R387 B.n498 B.n5 163.367
R388 B.n498 B.n497 163.367
R389 B.n497 B.n496 163.367
R390 B.n496 B.n7 163.367
R391 B.n492 B.n7 163.367
R392 B.n492 B.n491 163.367
R393 B.n491 B.n490 163.367
R394 B.n490 B.n9 163.367
R395 B.n486 B.n9 163.367
R396 B.n486 B.n485 163.367
R397 B.n485 B.n484 163.367
R398 B.n484 B.n11 163.367
R399 B.n480 B.n11 163.367
R400 B.n480 B.n479 163.367
R401 B.n479 B.n478 163.367
R402 B.n478 B.n13 163.367
R403 B.n474 B.n13 163.367
R404 B.n474 B.n473 163.367
R405 B.n473 B.n472 163.367
R406 B.n472 B.n15 163.367
R407 B.n468 B.n15 163.367
R408 B.n468 B.n467 163.367
R409 B.n467 B.n466 163.367
R410 B.n466 B.n17 163.367
R411 B.n462 B.n17 163.367
R412 B.n462 B.n461 163.367
R413 B.n461 B.n460 163.367
R414 B.n185 B.n118 163.367
R415 B.n189 B.n118 163.367
R416 B.n190 B.n189 163.367
R417 B.n191 B.n190 163.367
R418 B.n191 B.n116 163.367
R419 B.n195 B.n116 163.367
R420 B.n196 B.n195 163.367
R421 B.n197 B.n196 163.367
R422 B.n197 B.n114 163.367
R423 B.n201 B.n114 163.367
R424 B.n202 B.n201 163.367
R425 B.n203 B.n202 163.367
R426 B.n203 B.n112 163.367
R427 B.n207 B.n112 163.367
R428 B.n208 B.n207 163.367
R429 B.n209 B.n208 163.367
R430 B.n209 B.n110 163.367
R431 B.n213 B.n110 163.367
R432 B.n214 B.n213 163.367
R433 B.n215 B.n214 163.367
R434 B.n215 B.n108 163.367
R435 B.n219 B.n108 163.367
R436 B.n220 B.n219 163.367
R437 B.n220 B.n104 163.367
R438 B.n224 B.n104 163.367
R439 B.n225 B.n224 163.367
R440 B.n226 B.n225 163.367
R441 B.n226 B.n102 163.367
R442 B.n230 B.n102 163.367
R443 B.n231 B.n230 163.367
R444 B.n232 B.n231 163.367
R445 B.n232 B.n98 163.367
R446 B.n237 B.n98 163.367
R447 B.n238 B.n237 163.367
R448 B.n239 B.n238 163.367
R449 B.n239 B.n96 163.367
R450 B.n243 B.n96 163.367
R451 B.n244 B.n243 163.367
R452 B.n245 B.n244 163.367
R453 B.n245 B.n94 163.367
R454 B.n249 B.n94 163.367
R455 B.n250 B.n249 163.367
R456 B.n251 B.n250 163.367
R457 B.n251 B.n92 163.367
R458 B.n255 B.n92 163.367
R459 B.n256 B.n255 163.367
R460 B.n257 B.n256 163.367
R461 B.n257 B.n90 163.367
R462 B.n261 B.n90 163.367
R463 B.n262 B.n261 163.367
R464 B.n263 B.n262 163.367
R465 B.n263 B.n88 163.367
R466 B.n267 B.n88 163.367
R467 B.n268 B.n267 163.367
R468 B.n269 B.n268 163.367
R469 B.n273 B.n86 163.367
R470 B.n274 B.n273 163.367
R471 B.n275 B.n274 163.367
R472 B.n275 B.n84 163.367
R473 B.n279 B.n84 163.367
R474 B.n280 B.n279 163.367
R475 B.n281 B.n280 163.367
R476 B.n281 B.n82 163.367
R477 B.n285 B.n82 163.367
R478 B.n286 B.n285 163.367
R479 B.n287 B.n286 163.367
R480 B.n287 B.n80 163.367
R481 B.n291 B.n80 163.367
R482 B.n292 B.n291 163.367
R483 B.n293 B.n292 163.367
R484 B.n293 B.n78 163.367
R485 B.n297 B.n78 163.367
R486 B.n298 B.n297 163.367
R487 B.n299 B.n298 163.367
R488 B.n299 B.n76 163.367
R489 B.n303 B.n76 163.367
R490 B.n304 B.n303 163.367
R491 B.n305 B.n304 163.367
R492 B.n305 B.n74 163.367
R493 B.n309 B.n74 163.367
R494 B.n310 B.n309 163.367
R495 B.n311 B.n310 163.367
R496 B.n311 B.n72 163.367
R497 B.n315 B.n72 163.367
R498 B.n316 B.n315 163.367
R499 B.n317 B.n316 163.367
R500 B.n317 B.n70 163.367
R501 B.n321 B.n70 163.367
R502 B.n322 B.n321 163.367
R503 B.n323 B.n322 163.367
R504 B.n323 B.n68 163.367
R505 B.n327 B.n68 163.367
R506 B.n328 B.n327 163.367
R507 B.n329 B.n328 163.367
R508 B.n329 B.n66 163.367
R509 B.n333 B.n66 163.367
R510 B.n334 B.n333 163.367
R511 B.n335 B.n334 163.367
R512 B.n335 B.n64 163.367
R513 B.n339 B.n64 163.367
R514 B.n340 B.n339 163.367
R515 B.n341 B.n340 163.367
R516 B.n341 B.n62 163.367
R517 B.n345 B.n62 163.367
R518 B.n346 B.n345 163.367
R519 B.n347 B.n346 163.367
R520 B.n347 B.n60 163.367
R521 B.n351 B.n60 163.367
R522 B.n352 B.n351 163.367
R523 B.n353 B.n352 163.367
R524 B.n353 B.n58 163.367
R525 B.n357 B.n58 163.367
R526 B.n358 B.n357 163.367
R527 B.n359 B.n358 163.367
R528 B.n359 B.n56 163.367
R529 B.n363 B.n56 163.367
R530 B.n364 B.n363 163.367
R531 B.n365 B.n364 163.367
R532 B.n365 B.n54 163.367
R533 B.n369 B.n54 163.367
R534 B.n370 B.n369 163.367
R535 B.n371 B.n370 163.367
R536 B.n371 B.n52 163.367
R537 B.n456 B.n19 163.367
R538 B.n456 B.n455 163.367
R539 B.n455 B.n454 163.367
R540 B.n454 B.n21 163.367
R541 B.n450 B.n21 163.367
R542 B.n450 B.n449 163.367
R543 B.n449 B.n448 163.367
R544 B.n448 B.n23 163.367
R545 B.n444 B.n23 163.367
R546 B.n444 B.n443 163.367
R547 B.n443 B.n442 163.367
R548 B.n442 B.n25 163.367
R549 B.n438 B.n25 163.367
R550 B.n438 B.n437 163.367
R551 B.n437 B.n436 163.367
R552 B.n436 B.n27 163.367
R553 B.n432 B.n27 163.367
R554 B.n432 B.n431 163.367
R555 B.n431 B.n430 163.367
R556 B.n430 B.n29 163.367
R557 B.n426 B.n29 163.367
R558 B.n426 B.n425 163.367
R559 B.n425 B.n424 163.367
R560 B.n424 B.n31 163.367
R561 B.n420 B.n31 163.367
R562 B.n420 B.n419 163.367
R563 B.n419 B.n418 163.367
R564 B.n418 B.n36 163.367
R565 B.n414 B.n36 163.367
R566 B.n414 B.n413 163.367
R567 B.n413 B.n412 163.367
R568 B.n412 B.n38 163.367
R569 B.n407 B.n38 163.367
R570 B.n407 B.n406 163.367
R571 B.n406 B.n405 163.367
R572 B.n405 B.n42 163.367
R573 B.n401 B.n42 163.367
R574 B.n401 B.n400 163.367
R575 B.n400 B.n399 163.367
R576 B.n399 B.n44 163.367
R577 B.n395 B.n44 163.367
R578 B.n395 B.n394 163.367
R579 B.n394 B.n393 163.367
R580 B.n393 B.n46 163.367
R581 B.n389 B.n46 163.367
R582 B.n389 B.n388 163.367
R583 B.n388 B.n387 163.367
R584 B.n387 B.n48 163.367
R585 B.n383 B.n48 163.367
R586 B.n383 B.n382 163.367
R587 B.n382 B.n381 163.367
R588 B.n381 B.n50 163.367
R589 B.n377 B.n50 163.367
R590 B.n377 B.n376 163.367
R591 B.n376 B.n375 163.367
R592 B.n99 B.t8 159.607
R593 B.n39 B.t4 159.607
R594 B.n105 B.t2 159.601
R595 B.n32 B.t10 159.601
R596 B.n100 B.t7 116.552
R597 B.n40 B.t5 116.552
R598 B.n106 B.t1 116.547
R599 B.n33 B.t11 116.547
R600 B.n235 B.n100 59.5399
R601 B.n107 B.n106 59.5399
R602 B.n34 B.n33 59.5399
R603 B.n409 B.n40 59.5399
R604 B.n100 B.n99 43.055
R605 B.n106 B.n105 43.055
R606 B.n33 B.n32 43.055
R607 B.n40 B.n39 43.055
R608 B.n459 B.n458 32.6249
R609 B.n374 B.n373 32.6249
R610 B.n271 B.n270 32.6249
R611 B.n186 B.n119 32.6249
R612 B B.n511 18.0485
R613 B.n458 B.n457 10.6151
R614 B.n457 B.n20 10.6151
R615 B.n453 B.n20 10.6151
R616 B.n453 B.n452 10.6151
R617 B.n452 B.n451 10.6151
R618 B.n451 B.n22 10.6151
R619 B.n447 B.n22 10.6151
R620 B.n447 B.n446 10.6151
R621 B.n446 B.n445 10.6151
R622 B.n445 B.n24 10.6151
R623 B.n441 B.n24 10.6151
R624 B.n441 B.n440 10.6151
R625 B.n440 B.n439 10.6151
R626 B.n439 B.n26 10.6151
R627 B.n435 B.n26 10.6151
R628 B.n435 B.n434 10.6151
R629 B.n434 B.n433 10.6151
R630 B.n433 B.n28 10.6151
R631 B.n429 B.n28 10.6151
R632 B.n429 B.n428 10.6151
R633 B.n428 B.n427 10.6151
R634 B.n427 B.n30 10.6151
R635 B.n423 B.n422 10.6151
R636 B.n422 B.n421 10.6151
R637 B.n421 B.n35 10.6151
R638 B.n417 B.n35 10.6151
R639 B.n417 B.n416 10.6151
R640 B.n416 B.n415 10.6151
R641 B.n415 B.n37 10.6151
R642 B.n411 B.n37 10.6151
R643 B.n411 B.n410 10.6151
R644 B.n408 B.n41 10.6151
R645 B.n404 B.n41 10.6151
R646 B.n404 B.n403 10.6151
R647 B.n403 B.n402 10.6151
R648 B.n402 B.n43 10.6151
R649 B.n398 B.n43 10.6151
R650 B.n398 B.n397 10.6151
R651 B.n397 B.n396 10.6151
R652 B.n396 B.n45 10.6151
R653 B.n392 B.n45 10.6151
R654 B.n392 B.n391 10.6151
R655 B.n391 B.n390 10.6151
R656 B.n390 B.n47 10.6151
R657 B.n386 B.n47 10.6151
R658 B.n386 B.n385 10.6151
R659 B.n385 B.n384 10.6151
R660 B.n384 B.n49 10.6151
R661 B.n380 B.n49 10.6151
R662 B.n380 B.n379 10.6151
R663 B.n379 B.n378 10.6151
R664 B.n378 B.n51 10.6151
R665 B.n374 B.n51 10.6151
R666 B.n272 B.n271 10.6151
R667 B.n272 B.n85 10.6151
R668 B.n276 B.n85 10.6151
R669 B.n277 B.n276 10.6151
R670 B.n278 B.n277 10.6151
R671 B.n278 B.n83 10.6151
R672 B.n282 B.n83 10.6151
R673 B.n283 B.n282 10.6151
R674 B.n284 B.n283 10.6151
R675 B.n284 B.n81 10.6151
R676 B.n288 B.n81 10.6151
R677 B.n289 B.n288 10.6151
R678 B.n290 B.n289 10.6151
R679 B.n290 B.n79 10.6151
R680 B.n294 B.n79 10.6151
R681 B.n295 B.n294 10.6151
R682 B.n296 B.n295 10.6151
R683 B.n296 B.n77 10.6151
R684 B.n300 B.n77 10.6151
R685 B.n301 B.n300 10.6151
R686 B.n302 B.n301 10.6151
R687 B.n302 B.n75 10.6151
R688 B.n306 B.n75 10.6151
R689 B.n307 B.n306 10.6151
R690 B.n308 B.n307 10.6151
R691 B.n308 B.n73 10.6151
R692 B.n312 B.n73 10.6151
R693 B.n313 B.n312 10.6151
R694 B.n314 B.n313 10.6151
R695 B.n314 B.n71 10.6151
R696 B.n318 B.n71 10.6151
R697 B.n319 B.n318 10.6151
R698 B.n320 B.n319 10.6151
R699 B.n320 B.n69 10.6151
R700 B.n324 B.n69 10.6151
R701 B.n325 B.n324 10.6151
R702 B.n326 B.n325 10.6151
R703 B.n326 B.n67 10.6151
R704 B.n330 B.n67 10.6151
R705 B.n331 B.n330 10.6151
R706 B.n332 B.n331 10.6151
R707 B.n332 B.n65 10.6151
R708 B.n336 B.n65 10.6151
R709 B.n337 B.n336 10.6151
R710 B.n338 B.n337 10.6151
R711 B.n338 B.n63 10.6151
R712 B.n342 B.n63 10.6151
R713 B.n343 B.n342 10.6151
R714 B.n344 B.n343 10.6151
R715 B.n344 B.n61 10.6151
R716 B.n348 B.n61 10.6151
R717 B.n349 B.n348 10.6151
R718 B.n350 B.n349 10.6151
R719 B.n350 B.n59 10.6151
R720 B.n354 B.n59 10.6151
R721 B.n355 B.n354 10.6151
R722 B.n356 B.n355 10.6151
R723 B.n356 B.n57 10.6151
R724 B.n360 B.n57 10.6151
R725 B.n361 B.n360 10.6151
R726 B.n362 B.n361 10.6151
R727 B.n362 B.n55 10.6151
R728 B.n366 B.n55 10.6151
R729 B.n367 B.n366 10.6151
R730 B.n368 B.n367 10.6151
R731 B.n368 B.n53 10.6151
R732 B.n372 B.n53 10.6151
R733 B.n373 B.n372 10.6151
R734 B.n187 B.n186 10.6151
R735 B.n188 B.n187 10.6151
R736 B.n188 B.n117 10.6151
R737 B.n192 B.n117 10.6151
R738 B.n193 B.n192 10.6151
R739 B.n194 B.n193 10.6151
R740 B.n194 B.n115 10.6151
R741 B.n198 B.n115 10.6151
R742 B.n199 B.n198 10.6151
R743 B.n200 B.n199 10.6151
R744 B.n200 B.n113 10.6151
R745 B.n204 B.n113 10.6151
R746 B.n205 B.n204 10.6151
R747 B.n206 B.n205 10.6151
R748 B.n206 B.n111 10.6151
R749 B.n210 B.n111 10.6151
R750 B.n211 B.n210 10.6151
R751 B.n212 B.n211 10.6151
R752 B.n212 B.n109 10.6151
R753 B.n216 B.n109 10.6151
R754 B.n217 B.n216 10.6151
R755 B.n218 B.n217 10.6151
R756 B.n222 B.n221 10.6151
R757 B.n223 B.n222 10.6151
R758 B.n223 B.n103 10.6151
R759 B.n227 B.n103 10.6151
R760 B.n228 B.n227 10.6151
R761 B.n229 B.n228 10.6151
R762 B.n229 B.n101 10.6151
R763 B.n233 B.n101 10.6151
R764 B.n234 B.n233 10.6151
R765 B.n236 B.n97 10.6151
R766 B.n240 B.n97 10.6151
R767 B.n241 B.n240 10.6151
R768 B.n242 B.n241 10.6151
R769 B.n242 B.n95 10.6151
R770 B.n246 B.n95 10.6151
R771 B.n247 B.n246 10.6151
R772 B.n248 B.n247 10.6151
R773 B.n248 B.n93 10.6151
R774 B.n252 B.n93 10.6151
R775 B.n253 B.n252 10.6151
R776 B.n254 B.n253 10.6151
R777 B.n254 B.n91 10.6151
R778 B.n258 B.n91 10.6151
R779 B.n259 B.n258 10.6151
R780 B.n260 B.n259 10.6151
R781 B.n260 B.n89 10.6151
R782 B.n264 B.n89 10.6151
R783 B.n265 B.n264 10.6151
R784 B.n266 B.n265 10.6151
R785 B.n266 B.n87 10.6151
R786 B.n270 B.n87 10.6151
R787 B.n182 B.n119 10.6151
R788 B.n182 B.n181 10.6151
R789 B.n181 B.n180 10.6151
R790 B.n180 B.n121 10.6151
R791 B.n176 B.n121 10.6151
R792 B.n176 B.n175 10.6151
R793 B.n175 B.n174 10.6151
R794 B.n174 B.n123 10.6151
R795 B.n170 B.n123 10.6151
R796 B.n170 B.n169 10.6151
R797 B.n169 B.n168 10.6151
R798 B.n168 B.n125 10.6151
R799 B.n164 B.n125 10.6151
R800 B.n164 B.n163 10.6151
R801 B.n163 B.n162 10.6151
R802 B.n162 B.n127 10.6151
R803 B.n158 B.n127 10.6151
R804 B.n158 B.n157 10.6151
R805 B.n157 B.n156 10.6151
R806 B.n156 B.n129 10.6151
R807 B.n152 B.n129 10.6151
R808 B.n152 B.n151 10.6151
R809 B.n151 B.n150 10.6151
R810 B.n150 B.n131 10.6151
R811 B.n146 B.n131 10.6151
R812 B.n146 B.n145 10.6151
R813 B.n145 B.n144 10.6151
R814 B.n144 B.n133 10.6151
R815 B.n140 B.n133 10.6151
R816 B.n140 B.n139 10.6151
R817 B.n139 B.n138 10.6151
R818 B.n138 B.n135 10.6151
R819 B.n135 B.n0 10.6151
R820 B.n507 B.n1 10.6151
R821 B.n507 B.n506 10.6151
R822 B.n506 B.n505 10.6151
R823 B.n505 B.n4 10.6151
R824 B.n501 B.n4 10.6151
R825 B.n501 B.n500 10.6151
R826 B.n500 B.n499 10.6151
R827 B.n499 B.n6 10.6151
R828 B.n495 B.n6 10.6151
R829 B.n495 B.n494 10.6151
R830 B.n494 B.n493 10.6151
R831 B.n493 B.n8 10.6151
R832 B.n489 B.n8 10.6151
R833 B.n489 B.n488 10.6151
R834 B.n488 B.n487 10.6151
R835 B.n487 B.n10 10.6151
R836 B.n483 B.n10 10.6151
R837 B.n483 B.n482 10.6151
R838 B.n482 B.n481 10.6151
R839 B.n481 B.n12 10.6151
R840 B.n477 B.n12 10.6151
R841 B.n477 B.n476 10.6151
R842 B.n476 B.n475 10.6151
R843 B.n475 B.n14 10.6151
R844 B.n471 B.n14 10.6151
R845 B.n471 B.n470 10.6151
R846 B.n470 B.n469 10.6151
R847 B.n469 B.n16 10.6151
R848 B.n465 B.n16 10.6151
R849 B.n465 B.n464 10.6151
R850 B.n464 B.n463 10.6151
R851 B.n463 B.n18 10.6151
R852 B.n459 B.n18 10.6151
R853 B.n34 B.n30 9.36635
R854 B.n409 B.n408 9.36635
R855 B.n218 B.n107 9.36635
R856 B.n236 B.n235 9.36635
R857 B.n511 B.n0 2.81026
R858 B.n511 B.n1 2.81026
R859 B.n423 B.n34 1.24928
R860 B.n410 B.n409 1.24928
R861 B.n221 B.n107 1.24928
R862 B.n235 B.n234 1.24928
R863 VN.n21 VN.n12 161.3
R864 VN.n20 VN.n19 161.3
R865 VN.n18 VN.n13 161.3
R866 VN.n17 VN.n16 161.3
R867 VN.n9 VN.n0 161.3
R868 VN.n8 VN.n7 161.3
R869 VN.n6 VN.n1 161.3
R870 VN.n5 VN.n4 161.3
R871 VN.n2 VN.t1 103.392
R872 VN.n14 VN.t2 103.392
R873 VN.n11 VN.n10 87.7575
R874 VN.n23 VN.n22 87.7575
R875 VN.n3 VN.t3 72.3005
R876 VN.n10 VN.t0 72.3005
R877 VN.n15 VN.t5 72.3005
R878 VN.n22 VN.t4 72.3005
R879 VN.n3 VN.n2 57.8248
R880 VN.n15 VN.n14 57.8248
R881 VN.n8 VN.n1 54.0911
R882 VN.n20 VN.n13 54.0911
R883 VN VN.n23 41.4224
R884 VN.n9 VN.n8 26.8957
R885 VN.n21 VN.n20 26.8957
R886 VN.n4 VN.n1 24.4675
R887 VN.n16 VN.n13 24.4675
R888 VN.n10 VN.n9 22.9995
R889 VN.n22 VN.n21 22.9995
R890 VN.n17 VN.n14 12.851
R891 VN.n5 VN.n2 12.851
R892 VN.n4 VN.n3 12.234
R893 VN.n16 VN.n15 12.234
R894 VN.n23 VN.n12 0.278367
R895 VN.n11 VN.n0 0.278367
R896 VN.n19 VN.n12 0.189894
R897 VN.n19 VN.n18 0.189894
R898 VN.n18 VN.n17 0.189894
R899 VN.n6 VN.n5 0.189894
R900 VN.n7 VN.n6 0.189894
R901 VN.n7 VN.n0 0.189894
R902 VN VN.n11 0.153454
R903 VDD2.n1 VDD2.t4 102.335
R904 VDD2.n2 VDD2.t1 100.956
R905 VDD2.n1 VDD2.n0 95.6452
R906 VDD2 VDD2.n3 95.6424
R907 VDD2.n2 VDD2.n1 34.8231
R908 VDD2.n3 VDD2.t0 5.7333
R909 VDD2.n3 VDD2.t3 5.7333
R910 VDD2.n0 VDD2.t2 5.7333
R911 VDD2.n0 VDD2.t5 5.7333
R912 VDD2 VDD2.n2 1.49403
C0 B VP 1.52398f
C1 VDD1 B 1.41324f
C2 VN w_n2746_n2102# 4.91648f
C3 VDD1 VP 3.40365f
C4 VTAIL VDD2 5.1955f
C5 VTAIL w_n2746_n2102# 2.01091f
C6 VN B 0.938115f
C7 w_n2746_n2102# VDD2 1.73397f
C8 VN VP 5.06583f
C9 VDD1 VN 0.149787f
C10 VTAIL B 2.03384f
C11 VTAIL VP 3.54651f
C12 VDD1 VTAIL 5.14842f
C13 B VDD2 1.47044f
C14 VP VDD2 0.397571f
C15 VDD1 VDD2 1.15407f
C16 B w_n2746_n2102# 6.93012f
C17 VP w_n2746_n2102# 5.26952f
C18 VDD1 w_n2746_n2102# 1.67164f
C19 VTAIL VN 3.53229f
C20 VN VDD2 3.15794f
C21 VDD2 VSUBS 1.256635f
C22 VDD1 VSUBS 1.651167f
C23 VTAIL VSUBS 0.595332f
C24 VN VSUBS 4.89268f
C25 VP VSUBS 2.042605f
C26 B VSUBS 3.286648f
C27 w_n2746_n2102# VSUBS 72.1319f
C28 VDD2.t4 VSUBS 0.875535f
C29 VDD2.t2 VSUBS 0.098905f
C30 VDD2.t5 VSUBS 0.098905f
C31 VDD2.n0 VSUBS 0.647657f
C32 VDD2.n1 VSUBS 2.28943f
C33 VDD2.t1 VSUBS 0.868718f
C34 VDD2.n2 VSUBS 2.01475f
C35 VDD2.t0 VSUBS 0.098905f
C36 VDD2.t3 VSUBS 0.098905f
C37 VDD2.n3 VSUBS 0.647635f
C38 VN.n0 VSUBS 0.058345f
C39 VN.t0 VSUBS 1.25092f
C40 VN.n1 VSUBS 0.077569f
C41 VN.t1 VSUBS 1.46028f
C42 VN.n2 VSUBS 0.589258f
C43 VN.t3 VSUBS 1.25092f
C44 VN.n3 VSUBS 0.585653f
C45 VN.n4 VSUBS 0.062119f
C46 VN.n5 VSUBS 0.326914f
C47 VN.n6 VSUBS 0.044255f
C48 VN.n7 VSUBS 0.044255f
C49 VN.n8 VSUBS 0.048332f
C50 VN.n9 VSUBS 0.083343f
C51 VN.n10 VSUBS 0.620565f
C52 VN.n11 VSUBS 0.048773f
C53 VN.n12 VSUBS 0.058345f
C54 VN.t4 VSUBS 1.25092f
C55 VN.n13 VSUBS 0.077569f
C56 VN.t2 VSUBS 1.46028f
C57 VN.n14 VSUBS 0.589258f
C58 VN.t5 VSUBS 1.25092f
C59 VN.n15 VSUBS 0.585653f
C60 VN.n16 VSUBS 0.062119f
C61 VN.n17 VSUBS 0.326914f
C62 VN.n18 VSUBS 0.044255f
C63 VN.n19 VSUBS 0.044255f
C64 VN.n20 VSUBS 0.048332f
C65 VN.n21 VSUBS 0.083343f
C66 VN.n22 VSUBS 0.620565f
C67 VN.n23 VSUBS 1.82142f
C68 B.n0 VSUBS 0.00507f
C69 B.n1 VSUBS 0.00507f
C70 B.n2 VSUBS 0.008018f
C71 B.n3 VSUBS 0.008018f
C72 B.n4 VSUBS 0.008018f
C73 B.n5 VSUBS 0.008018f
C74 B.n6 VSUBS 0.008018f
C75 B.n7 VSUBS 0.008018f
C76 B.n8 VSUBS 0.008018f
C77 B.n9 VSUBS 0.008018f
C78 B.n10 VSUBS 0.008018f
C79 B.n11 VSUBS 0.008018f
C80 B.n12 VSUBS 0.008018f
C81 B.n13 VSUBS 0.008018f
C82 B.n14 VSUBS 0.008018f
C83 B.n15 VSUBS 0.008018f
C84 B.n16 VSUBS 0.008018f
C85 B.n17 VSUBS 0.008018f
C86 B.n18 VSUBS 0.008018f
C87 B.n19 VSUBS 0.019547f
C88 B.n20 VSUBS 0.008018f
C89 B.n21 VSUBS 0.008018f
C90 B.n22 VSUBS 0.008018f
C91 B.n23 VSUBS 0.008018f
C92 B.n24 VSUBS 0.008018f
C93 B.n25 VSUBS 0.008018f
C94 B.n26 VSUBS 0.008018f
C95 B.n27 VSUBS 0.008018f
C96 B.n28 VSUBS 0.008018f
C97 B.n29 VSUBS 0.008018f
C98 B.n30 VSUBS 0.007547f
C99 B.n31 VSUBS 0.008018f
C100 B.t11 VSUBS 0.186995f
C101 B.t10 VSUBS 0.204863f
C102 B.t9 VSUBS 0.572482f
C103 B.n32 VSUBS 0.119619f
C104 B.n33 VSUBS 0.077672f
C105 B.n34 VSUBS 0.018577f
C106 B.n35 VSUBS 0.008018f
C107 B.n36 VSUBS 0.008018f
C108 B.n37 VSUBS 0.008018f
C109 B.n38 VSUBS 0.008018f
C110 B.t5 VSUBS 0.186995f
C111 B.t4 VSUBS 0.204862f
C112 B.t3 VSUBS 0.572482f
C113 B.n39 VSUBS 0.11962f
C114 B.n40 VSUBS 0.077672f
C115 B.n41 VSUBS 0.008018f
C116 B.n42 VSUBS 0.008018f
C117 B.n43 VSUBS 0.008018f
C118 B.n44 VSUBS 0.008018f
C119 B.n45 VSUBS 0.008018f
C120 B.n46 VSUBS 0.008018f
C121 B.n47 VSUBS 0.008018f
C122 B.n48 VSUBS 0.008018f
C123 B.n49 VSUBS 0.008018f
C124 B.n50 VSUBS 0.008018f
C125 B.n51 VSUBS 0.008018f
C126 B.n52 VSUBS 0.017951f
C127 B.n53 VSUBS 0.008018f
C128 B.n54 VSUBS 0.008018f
C129 B.n55 VSUBS 0.008018f
C130 B.n56 VSUBS 0.008018f
C131 B.n57 VSUBS 0.008018f
C132 B.n58 VSUBS 0.008018f
C133 B.n59 VSUBS 0.008018f
C134 B.n60 VSUBS 0.008018f
C135 B.n61 VSUBS 0.008018f
C136 B.n62 VSUBS 0.008018f
C137 B.n63 VSUBS 0.008018f
C138 B.n64 VSUBS 0.008018f
C139 B.n65 VSUBS 0.008018f
C140 B.n66 VSUBS 0.008018f
C141 B.n67 VSUBS 0.008018f
C142 B.n68 VSUBS 0.008018f
C143 B.n69 VSUBS 0.008018f
C144 B.n70 VSUBS 0.008018f
C145 B.n71 VSUBS 0.008018f
C146 B.n72 VSUBS 0.008018f
C147 B.n73 VSUBS 0.008018f
C148 B.n74 VSUBS 0.008018f
C149 B.n75 VSUBS 0.008018f
C150 B.n76 VSUBS 0.008018f
C151 B.n77 VSUBS 0.008018f
C152 B.n78 VSUBS 0.008018f
C153 B.n79 VSUBS 0.008018f
C154 B.n80 VSUBS 0.008018f
C155 B.n81 VSUBS 0.008018f
C156 B.n82 VSUBS 0.008018f
C157 B.n83 VSUBS 0.008018f
C158 B.n84 VSUBS 0.008018f
C159 B.n85 VSUBS 0.008018f
C160 B.n86 VSUBS 0.017951f
C161 B.n87 VSUBS 0.008018f
C162 B.n88 VSUBS 0.008018f
C163 B.n89 VSUBS 0.008018f
C164 B.n90 VSUBS 0.008018f
C165 B.n91 VSUBS 0.008018f
C166 B.n92 VSUBS 0.008018f
C167 B.n93 VSUBS 0.008018f
C168 B.n94 VSUBS 0.008018f
C169 B.n95 VSUBS 0.008018f
C170 B.n96 VSUBS 0.008018f
C171 B.n97 VSUBS 0.008018f
C172 B.n98 VSUBS 0.008018f
C173 B.t7 VSUBS 0.186995f
C174 B.t8 VSUBS 0.204862f
C175 B.t6 VSUBS 0.572482f
C176 B.n99 VSUBS 0.11962f
C177 B.n100 VSUBS 0.077672f
C178 B.n101 VSUBS 0.008018f
C179 B.n102 VSUBS 0.008018f
C180 B.n103 VSUBS 0.008018f
C181 B.n104 VSUBS 0.008018f
C182 B.t1 VSUBS 0.186995f
C183 B.t2 VSUBS 0.204863f
C184 B.t0 VSUBS 0.572482f
C185 B.n105 VSUBS 0.119619f
C186 B.n106 VSUBS 0.077672f
C187 B.n107 VSUBS 0.018577f
C188 B.n108 VSUBS 0.008018f
C189 B.n109 VSUBS 0.008018f
C190 B.n110 VSUBS 0.008018f
C191 B.n111 VSUBS 0.008018f
C192 B.n112 VSUBS 0.008018f
C193 B.n113 VSUBS 0.008018f
C194 B.n114 VSUBS 0.008018f
C195 B.n115 VSUBS 0.008018f
C196 B.n116 VSUBS 0.008018f
C197 B.n117 VSUBS 0.008018f
C198 B.n118 VSUBS 0.008018f
C199 B.n119 VSUBS 0.017951f
C200 B.n120 VSUBS 0.008018f
C201 B.n121 VSUBS 0.008018f
C202 B.n122 VSUBS 0.008018f
C203 B.n123 VSUBS 0.008018f
C204 B.n124 VSUBS 0.008018f
C205 B.n125 VSUBS 0.008018f
C206 B.n126 VSUBS 0.008018f
C207 B.n127 VSUBS 0.008018f
C208 B.n128 VSUBS 0.008018f
C209 B.n129 VSUBS 0.008018f
C210 B.n130 VSUBS 0.008018f
C211 B.n131 VSUBS 0.008018f
C212 B.n132 VSUBS 0.008018f
C213 B.n133 VSUBS 0.008018f
C214 B.n134 VSUBS 0.008018f
C215 B.n135 VSUBS 0.008018f
C216 B.n136 VSUBS 0.008018f
C217 B.n137 VSUBS 0.008018f
C218 B.n138 VSUBS 0.008018f
C219 B.n139 VSUBS 0.008018f
C220 B.n140 VSUBS 0.008018f
C221 B.n141 VSUBS 0.008018f
C222 B.n142 VSUBS 0.008018f
C223 B.n143 VSUBS 0.008018f
C224 B.n144 VSUBS 0.008018f
C225 B.n145 VSUBS 0.008018f
C226 B.n146 VSUBS 0.008018f
C227 B.n147 VSUBS 0.008018f
C228 B.n148 VSUBS 0.008018f
C229 B.n149 VSUBS 0.008018f
C230 B.n150 VSUBS 0.008018f
C231 B.n151 VSUBS 0.008018f
C232 B.n152 VSUBS 0.008018f
C233 B.n153 VSUBS 0.008018f
C234 B.n154 VSUBS 0.008018f
C235 B.n155 VSUBS 0.008018f
C236 B.n156 VSUBS 0.008018f
C237 B.n157 VSUBS 0.008018f
C238 B.n158 VSUBS 0.008018f
C239 B.n159 VSUBS 0.008018f
C240 B.n160 VSUBS 0.008018f
C241 B.n161 VSUBS 0.008018f
C242 B.n162 VSUBS 0.008018f
C243 B.n163 VSUBS 0.008018f
C244 B.n164 VSUBS 0.008018f
C245 B.n165 VSUBS 0.008018f
C246 B.n166 VSUBS 0.008018f
C247 B.n167 VSUBS 0.008018f
C248 B.n168 VSUBS 0.008018f
C249 B.n169 VSUBS 0.008018f
C250 B.n170 VSUBS 0.008018f
C251 B.n171 VSUBS 0.008018f
C252 B.n172 VSUBS 0.008018f
C253 B.n173 VSUBS 0.008018f
C254 B.n174 VSUBS 0.008018f
C255 B.n175 VSUBS 0.008018f
C256 B.n176 VSUBS 0.008018f
C257 B.n177 VSUBS 0.008018f
C258 B.n178 VSUBS 0.008018f
C259 B.n179 VSUBS 0.008018f
C260 B.n180 VSUBS 0.008018f
C261 B.n181 VSUBS 0.008018f
C262 B.n182 VSUBS 0.008018f
C263 B.n183 VSUBS 0.008018f
C264 B.n184 VSUBS 0.017951f
C265 B.n185 VSUBS 0.019547f
C266 B.n186 VSUBS 0.019547f
C267 B.n187 VSUBS 0.008018f
C268 B.n188 VSUBS 0.008018f
C269 B.n189 VSUBS 0.008018f
C270 B.n190 VSUBS 0.008018f
C271 B.n191 VSUBS 0.008018f
C272 B.n192 VSUBS 0.008018f
C273 B.n193 VSUBS 0.008018f
C274 B.n194 VSUBS 0.008018f
C275 B.n195 VSUBS 0.008018f
C276 B.n196 VSUBS 0.008018f
C277 B.n197 VSUBS 0.008018f
C278 B.n198 VSUBS 0.008018f
C279 B.n199 VSUBS 0.008018f
C280 B.n200 VSUBS 0.008018f
C281 B.n201 VSUBS 0.008018f
C282 B.n202 VSUBS 0.008018f
C283 B.n203 VSUBS 0.008018f
C284 B.n204 VSUBS 0.008018f
C285 B.n205 VSUBS 0.008018f
C286 B.n206 VSUBS 0.008018f
C287 B.n207 VSUBS 0.008018f
C288 B.n208 VSUBS 0.008018f
C289 B.n209 VSUBS 0.008018f
C290 B.n210 VSUBS 0.008018f
C291 B.n211 VSUBS 0.008018f
C292 B.n212 VSUBS 0.008018f
C293 B.n213 VSUBS 0.008018f
C294 B.n214 VSUBS 0.008018f
C295 B.n215 VSUBS 0.008018f
C296 B.n216 VSUBS 0.008018f
C297 B.n217 VSUBS 0.008018f
C298 B.n218 VSUBS 0.007547f
C299 B.n219 VSUBS 0.008018f
C300 B.n220 VSUBS 0.008018f
C301 B.n221 VSUBS 0.004481f
C302 B.n222 VSUBS 0.008018f
C303 B.n223 VSUBS 0.008018f
C304 B.n224 VSUBS 0.008018f
C305 B.n225 VSUBS 0.008018f
C306 B.n226 VSUBS 0.008018f
C307 B.n227 VSUBS 0.008018f
C308 B.n228 VSUBS 0.008018f
C309 B.n229 VSUBS 0.008018f
C310 B.n230 VSUBS 0.008018f
C311 B.n231 VSUBS 0.008018f
C312 B.n232 VSUBS 0.008018f
C313 B.n233 VSUBS 0.008018f
C314 B.n234 VSUBS 0.004481f
C315 B.n235 VSUBS 0.018577f
C316 B.n236 VSUBS 0.007547f
C317 B.n237 VSUBS 0.008018f
C318 B.n238 VSUBS 0.008018f
C319 B.n239 VSUBS 0.008018f
C320 B.n240 VSUBS 0.008018f
C321 B.n241 VSUBS 0.008018f
C322 B.n242 VSUBS 0.008018f
C323 B.n243 VSUBS 0.008018f
C324 B.n244 VSUBS 0.008018f
C325 B.n245 VSUBS 0.008018f
C326 B.n246 VSUBS 0.008018f
C327 B.n247 VSUBS 0.008018f
C328 B.n248 VSUBS 0.008018f
C329 B.n249 VSUBS 0.008018f
C330 B.n250 VSUBS 0.008018f
C331 B.n251 VSUBS 0.008018f
C332 B.n252 VSUBS 0.008018f
C333 B.n253 VSUBS 0.008018f
C334 B.n254 VSUBS 0.008018f
C335 B.n255 VSUBS 0.008018f
C336 B.n256 VSUBS 0.008018f
C337 B.n257 VSUBS 0.008018f
C338 B.n258 VSUBS 0.008018f
C339 B.n259 VSUBS 0.008018f
C340 B.n260 VSUBS 0.008018f
C341 B.n261 VSUBS 0.008018f
C342 B.n262 VSUBS 0.008018f
C343 B.n263 VSUBS 0.008018f
C344 B.n264 VSUBS 0.008018f
C345 B.n265 VSUBS 0.008018f
C346 B.n266 VSUBS 0.008018f
C347 B.n267 VSUBS 0.008018f
C348 B.n268 VSUBS 0.008018f
C349 B.n269 VSUBS 0.019547f
C350 B.n270 VSUBS 0.019547f
C351 B.n271 VSUBS 0.017951f
C352 B.n272 VSUBS 0.008018f
C353 B.n273 VSUBS 0.008018f
C354 B.n274 VSUBS 0.008018f
C355 B.n275 VSUBS 0.008018f
C356 B.n276 VSUBS 0.008018f
C357 B.n277 VSUBS 0.008018f
C358 B.n278 VSUBS 0.008018f
C359 B.n279 VSUBS 0.008018f
C360 B.n280 VSUBS 0.008018f
C361 B.n281 VSUBS 0.008018f
C362 B.n282 VSUBS 0.008018f
C363 B.n283 VSUBS 0.008018f
C364 B.n284 VSUBS 0.008018f
C365 B.n285 VSUBS 0.008018f
C366 B.n286 VSUBS 0.008018f
C367 B.n287 VSUBS 0.008018f
C368 B.n288 VSUBS 0.008018f
C369 B.n289 VSUBS 0.008018f
C370 B.n290 VSUBS 0.008018f
C371 B.n291 VSUBS 0.008018f
C372 B.n292 VSUBS 0.008018f
C373 B.n293 VSUBS 0.008018f
C374 B.n294 VSUBS 0.008018f
C375 B.n295 VSUBS 0.008018f
C376 B.n296 VSUBS 0.008018f
C377 B.n297 VSUBS 0.008018f
C378 B.n298 VSUBS 0.008018f
C379 B.n299 VSUBS 0.008018f
C380 B.n300 VSUBS 0.008018f
C381 B.n301 VSUBS 0.008018f
C382 B.n302 VSUBS 0.008018f
C383 B.n303 VSUBS 0.008018f
C384 B.n304 VSUBS 0.008018f
C385 B.n305 VSUBS 0.008018f
C386 B.n306 VSUBS 0.008018f
C387 B.n307 VSUBS 0.008018f
C388 B.n308 VSUBS 0.008018f
C389 B.n309 VSUBS 0.008018f
C390 B.n310 VSUBS 0.008018f
C391 B.n311 VSUBS 0.008018f
C392 B.n312 VSUBS 0.008018f
C393 B.n313 VSUBS 0.008018f
C394 B.n314 VSUBS 0.008018f
C395 B.n315 VSUBS 0.008018f
C396 B.n316 VSUBS 0.008018f
C397 B.n317 VSUBS 0.008018f
C398 B.n318 VSUBS 0.008018f
C399 B.n319 VSUBS 0.008018f
C400 B.n320 VSUBS 0.008018f
C401 B.n321 VSUBS 0.008018f
C402 B.n322 VSUBS 0.008018f
C403 B.n323 VSUBS 0.008018f
C404 B.n324 VSUBS 0.008018f
C405 B.n325 VSUBS 0.008018f
C406 B.n326 VSUBS 0.008018f
C407 B.n327 VSUBS 0.008018f
C408 B.n328 VSUBS 0.008018f
C409 B.n329 VSUBS 0.008018f
C410 B.n330 VSUBS 0.008018f
C411 B.n331 VSUBS 0.008018f
C412 B.n332 VSUBS 0.008018f
C413 B.n333 VSUBS 0.008018f
C414 B.n334 VSUBS 0.008018f
C415 B.n335 VSUBS 0.008018f
C416 B.n336 VSUBS 0.008018f
C417 B.n337 VSUBS 0.008018f
C418 B.n338 VSUBS 0.008018f
C419 B.n339 VSUBS 0.008018f
C420 B.n340 VSUBS 0.008018f
C421 B.n341 VSUBS 0.008018f
C422 B.n342 VSUBS 0.008018f
C423 B.n343 VSUBS 0.008018f
C424 B.n344 VSUBS 0.008018f
C425 B.n345 VSUBS 0.008018f
C426 B.n346 VSUBS 0.008018f
C427 B.n347 VSUBS 0.008018f
C428 B.n348 VSUBS 0.008018f
C429 B.n349 VSUBS 0.008018f
C430 B.n350 VSUBS 0.008018f
C431 B.n351 VSUBS 0.008018f
C432 B.n352 VSUBS 0.008018f
C433 B.n353 VSUBS 0.008018f
C434 B.n354 VSUBS 0.008018f
C435 B.n355 VSUBS 0.008018f
C436 B.n356 VSUBS 0.008018f
C437 B.n357 VSUBS 0.008018f
C438 B.n358 VSUBS 0.008018f
C439 B.n359 VSUBS 0.008018f
C440 B.n360 VSUBS 0.008018f
C441 B.n361 VSUBS 0.008018f
C442 B.n362 VSUBS 0.008018f
C443 B.n363 VSUBS 0.008018f
C444 B.n364 VSUBS 0.008018f
C445 B.n365 VSUBS 0.008018f
C446 B.n366 VSUBS 0.008018f
C447 B.n367 VSUBS 0.008018f
C448 B.n368 VSUBS 0.008018f
C449 B.n369 VSUBS 0.008018f
C450 B.n370 VSUBS 0.008018f
C451 B.n371 VSUBS 0.008018f
C452 B.n372 VSUBS 0.008018f
C453 B.n373 VSUBS 0.018899f
C454 B.n374 VSUBS 0.018598f
C455 B.n375 VSUBS 0.019547f
C456 B.n376 VSUBS 0.008018f
C457 B.n377 VSUBS 0.008018f
C458 B.n378 VSUBS 0.008018f
C459 B.n379 VSUBS 0.008018f
C460 B.n380 VSUBS 0.008018f
C461 B.n381 VSUBS 0.008018f
C462 B.n382 VSUBS 0.008018f
C463 B.n383 VSUBS 0.008018f
C464 B.n384 VSUBS 0.008018f
C465 B.n385 VSUBS 0.008018f
C466 B.n386 VSUBS 0.008018f
C467 B.n387 VSUBS 0.008018f
C468 B.n388 VSUBS 0.008018f
C469 B.n389 VSUBS 0.008018f
C470 B.n390 VSUBS 0.008018f
C471 B.n391 VSUBS 0.008018f
C472 B.n392 VSUBS 0.008018f
C473 B.n393 VSUBS 0.008018f
C474 B.n394 VSUBS 0.008018f
C475 B.n395 VSUBS 0.008018f
C476 B.n396 VSUBS 0.008018f
C477 B.n397 VSUBS 0.008018f
C478 B.n398 VSUBS 0.008018f
C479 B.n399 VSUBS 0.008018f
C480 B.n400 VSUBS 0.008018f
C481 B.n401 VSUBS 0.008018f
C482 B.n402 VSUBS 0.008018f
C483 B.n403 VSUBS 0.008018f
C484 B.n404 VSUBS 0.008018f
C485 B.n405 VSUBS 0.008018f
C486 B.n406 VSUBS 0.008018f
C487 B.n407 VSUBS 0.008018f
C488 B.n408 VSUBS 0.007547f
C489 B.n409 VSUBS 0.018577f
C490 B.n410 VSUBS 0.004481f
C491 B.n411 VSUBS 0.008018f
C492 B.n412 VSUBS 0.008018f
C493 B.n413 VSUBS 0.008018f
C494 B.n414 VSUBS 0.008018f
C495 B.n415 VSUBS 0.008018f
C496 B.n416 VSUBS 0.008018f
C497 B.n417 VSUBS 0.008018f
C498 B.n418 VSUBS 0.008018f
C499 B.n419 VSUBS 0.008018f
C500 B.n420 VSUBS 0.008018f
C501 B.n421 VSUBS 0.008018f
C502 B.n422 VSUBS 0.008018f
C503 B.n423 VSUBS 0.004481f
C504 B.n424 VSUBS 0.008018f
C505 B.n425 VSUBS 0.008018f
C506 B.n426 VSUBS 0.008018f
C507 B.n427 VSUBS 0.008018f
C508 B.n428 VSUBS 0.008018f
C509 B.n429 VSUBS 0.008018f
C510 B.n430 VSUBS 0.008018f
C511 B.n431 VSUBS 0.008018f
C512 B.n432 VSUBS 0.008018f
C513 B.n433 VSUBS 0.008018f
C514 B.n434 VSUBS 0.008018f
C515 B.n435 VSUBS 0.008018f
C516 B.n436 VSUBS 0.008018f
C517 B.n437 VSUBS 0.008018f
C518 B.n438 VSUBS 0.008018f
C519 B.n439 VSUBS 0.008018f
C520 B.n440 VSUBS 0.008018f
C521 B.n441 VSUBS 0.008018f
C522 B.n442 VSUBS 0.008018f
C523 B.n443 VSUBS 0.008018f
C524 B.n444 VSUBS 0.008018f
C525 B.n445 VSUBS 0.008018f
C526 B.n446 VSUBS 0.008018f
C527 B.n447 VSUBS 0.008018f
C528 B.n448 VSUBS 0.008018f
C529 B.n449 VSUBS 0.008018f
C530 B.n450 VSUBS 0.008018f
C531 B.n451 VSUBS 0.008018f
C532 B.n452 VSUBS 0.008018f
C533 B.n453 VSUBS 0.008018f
C534 B.n454 VSUBS 0.008018f
C535 B.n455 VSUBS 0.008018f
C536 B.n456 VSUBS 0.008018f
C537 B.n457 VSUBS 0.008018f
C538 B.n458 VSUBS 0.019547f
C539 B.n459 VSUBS 0.017951f
C540 B.n460 VSUBS 0.017951f
C541 B.n461 VSUBS 0.008018f
C542 B.n462 VSUBS 0.008018f
C543 B.n463 VSUBS 0.008018f
C544 B.n464 VSUBS 0.008018f
C545 B.n465 VSUBS 0.008018f
C546 B.n466 VSUBS 0.008018f
C547 B.n467 VSUBS 0.008018f
C548 B.n468 VSUBS 0.008018f
C549 B.n469 VSUBS 0.008018f
C550 B.n470 VSUBS 0.008018f
C551 B.n471 VSUBS 0.008018f
C552 B.n472 VSUBS 0.008018f
C553 B.n473 VSUBS 0.008018f
C554 B.n474 VSUBS 0.008018f
C555 B.n475 VSUBS 0.008018f
C556 B.n476 VSUBS 0.008018f
C557 B.n477 VSUBS 0.008018f
C558 B.n478 VSUBS 0.008018f
C559 B.n479 VSUBS 0.008018f
C560 B.n480 VSUBS 0.008018f
C561 B.n481 VSUBS 0.008018f
C562 B.n482 VSUBS 0.008018f
C563 B.n483 VSUBS 0.008018f
C564 B.n484 VSUBS 0.008018f
C565 B.n485 VSUBS 0.008018f
C566 B.n486 VSUBS 0.008018f
C567 B.n487 VSUBS 0.008018f
C568 B.n488 VSUBS 0.008018f
C569 B.n489 VSUBS 0.008018f
C570 B.n490 VSUBS 0.008018f
C571 B.n491 VSUBS 0.008018f
C572 B.n492 VSUBS 0.008018f
C573 B.n493 VSUBS 0.008018f
C574 B.n494 VSUBS 0.008018f
C575 B.n495 VSUBS 0.008018f
C576 B.n496 VSUBS 0.008018f
C577 B.n497 VSUBS 0.008018f
C578 B.n498 VSUBS 0.008018f
C579 B.n499 VSUBS 0.008018f
C580 B.n500 VSUBS 0.008018f
C581 B.n501 VSUBS 0.008018f
C582 B.n502 VSUBS 0.008018f
C583 B.n503 VSUBS 0.008018f
C584 B.n504 VSUBS 0.008018f
C585 B.n505 VSUBS 0.008018f
C586 B.n506 VSUBS 0.008018f
C587 B.n507 VSUBS 0.008018f
C588 B.n508 VSUBS 0.008018f
C589 B.n509 VSUBS 0.008018f
C590 B.n510 VSUBS 0.008018f
C591 B.n511 VSUBS 0.018156f
C592 VDD1.t4 VSUBS 0.878111f
C593 VDD1.t0 VSUBS 0.877441f
C594 VDD1.t2 VSUBS 0.09912f
C595 VDD1.t5 VSUBS 0.09912f
C596 VDD1.n0 VSUBS 0.649068f
C597 VDD1.n1 VSUBS 2.38374f
C598 VDD1.t1 VSUBS 0.09912f
C599 VDD1.t3 VSUBS 0.09912f
C600 VDD1.n2 VSUBS 0.646725f
C601 VDD1.n3 VSUBS 2.02499f
C602 VTAIL.t1 VSUBS 0.145188f
C603 VTAIL.t9 VSUBS 0.145188f
C604 VTAIL.n0 VSUBS 0.838901f
C605 VTAIL.n1 VSUBS 0.785992f
C606 VTAIL.t4 VSUBS 1.16074f
C607 VTAIL.n2 VSUBS 1.00391f
C608 VTAIL.t5 VSUBS 0.145188f
C609 VTAIL.t8 VSUBS 0.145188f
C610 VTAIL.n3 VSUBS 0.838901f
C611 VTAIL.n4 VSUBS 2.13098f
C612 VTAIL.t11 VSUBS 0.145188f
C613 VTAIL.t10 VSUBS 0.145188f
C614 VTAIL.n5 VSUBS 0.838905f
C615 VTAIL.n6 VSUBS 2.13098f
C616 VTAIL.t0 VSUBS 1.16075f
C617 VTAIL.n7 VSUBS 1.0039f
C618 VTAIL.t3 VSUBS 0.145188f
C619 VTAIL.t7 VSUBS 0.145188f
C620 VTAIL.n8 VSUBS 0.838905f
C621 VTAIL.n9 VSUBS 0.929778f
C622 VTAIL.t6 VSUBS 1.16074f
C623 VTAIL.n10 VSUBS 2.00529f
C624 VTAIL.t2 VSUBS 1.16074f
C625 VTAIL.n11 VSUBS 1.94926f
C626 VP.n0 VSUBS 0.060667f
C627 VP.t0 VSUBS 1.30071f
C628 VP.n1 VSUBS 0.080657f
C629 VP.n2 VSUBS 0.046016f
C630 VP.t3 VSUBS 1.30071f
C631 VP.n3 VSUBS 0.050255f
C632 VP.n4 VSUBS 0.060667f
C633 VP.t2 VSUBS 1.30071f
C634 VP.n5 VSUBS 0.080657f
C635 VP.t1 VSUBS 1.5184f
C636 VP.n6 VSUBS 0.612711f
C637 VP.t4 VSUBS 1.30071f
C638 VP.n7 VSUBS 0.608963f
C639 VP.n8 VSUBS 0.064591f
C640 VP.n9 VSUBS 0.339926f
C641 VP.n10 VSUBS 0.046016f
C642 VP.n11 VSUBS 0.046016f
C643 VP.n12 VSUBS 0.050255f
C644 VP.n13 VSUBS 0.08666f
C645 VP.n14 VSUBS 0.645265f
C646 VP.n15 VSUBS 1.86835f
C647 VP.n16 VSUBS 1.90855f
C648 VP.t5 VSUBS 1.30071f
C649 VP.n17 VSUBS 0.645265f
C650 VP.n18 VSUBS 0.08666f
C651 VP.n19 VSUBS 0.060667f
C652 VP.n20 VSUBS 0.046016f
C653 VP.n21 VSUBS 0.046016f
C654 VP.n22 VSUBS 0.080657f
C655 VP.n23 VSUBS 0.064591f
C656 VP.n24 VSUBS 0.502993f
C657 VP.n25 VSUBS 0.064591f
C658 VP.n26 VSUBS 0.046016f
C659 VP.n27 VSUBS 0.046016f
C660 VP.n28 VSUBS 0.046016f
C661 VP.n29 VSUBS 0.050255f
C662 VP.n30 VSUBS 0.08666f
C663 VP.n31 VSUBS 0.645265f
C664 VP.n32 VSUBS 0.050714f
.ends

