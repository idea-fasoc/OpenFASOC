* NGSPICE file created from diff_pair_sample_0177.ext - technology: sky130A

.subckt diff_pair_sample_0177 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t9 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8347 pd=17.51 as=6.7002 ps=35.14 w=17.18 l=0.55
X1 VTAIL.t5 VP.t1 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8347 pd=17.51 as=2.8347 ps=17.51 w=17.18 l=0.55
X2 VDD2.t5 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8347 pd=17.51 as=6.7002 ps=35.14 w=17.18 l=0.55
X3 VDD1.t3 VP.t2 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=2.8347 pd=17.51 as=6.7002 ps=35.14 w=17.18 l=0.55
X4 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7002 pd=35.14 as=0 ps=0 w=17.18 l=0.55
X5 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=6.7002 pd=35.14 as=0 ps=0 w=17.18 l=0.55
X6 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.7002 pd=35.14 as=0 ps=0 w=17.18 l=0.55
X7 VDD2.t4 VN.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.8347 pd=17.51 as=6.7002 ps=35.14 w=17.18 l=0.55
X8 VTAIL.t11 VN.t2 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8347 pd=17.51 as=2.8347 ps=17.51 w=17.18 l=0.55
X9 VTAIL.t6 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8347 pd=17.51 as=2.8347 ps=17.51 w=17.18 l=0.55
X10 VDD2.t2 VN.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=6.7002 pd=35.14 as=2.8347 ps=17.51 w=17.18 l=0.55
X11 VTAIL.t1 VN.t4 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.8347 pd=17.51 as=2.8347 ps=17.51 w=17.18 l=0.55
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.7002 pd=35.14 as=0 ps=0 w=17.18 l=0.55
X13 VDD1.t1 VP.t4 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=6.7002 pd=35.14 as=2.8347 ps=17.51 w=17.18 l=0.55
X14 VDD1.t0 VP.t5 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=6.7002 pd=35.14 as=2.8347 ps=17.51 w=17.18 l=0.55
X15 VDD2.t0 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=6.7002 pd=35.14 as=2.8347 ps=17.51 w=17.18 l=0.55
R0 VP.n1 VP.t5 851.042
R1 VP.n6 VP.t4 824.221
R2 VP.n7 VP.t3 824.221
R3 VP.n8 VP.t0 824.221
R4 VP.n3 VP.t2 824.221
R5 VP.n2 VP.t1 824.221
R6 VP.n9 VP.n8 161.3
R7 VP.n4 VP.n3 161.3
R8 VP.n6 VP.n5 161.3
R9 VP.n7 VP.n0 80.6037
R10 VP.n7 VP.n6 48.2005
R11 VP.n8 VP.n7 48.2005
R12 VP.n3 VP.n2 48.2005
R13 VP.n4 VP.n1 45.1367
R14 VP.n5 VP.n4 44.5763
R15 VP.n2 VP.n1 13.3799
R16 VP.n5 VP.n0 0.285035
R17 VP.n9 VP.n0 0.285035
R18 VP VP.n9 0.0516364
R19 VTAIL.n7 VTAIL.t4 45.5636
R20 VTAIL.n11 VTAIL.t3 45.5635
R21 VTAIL.n2 VTAIL.t9 45.5635
R22 VTAIL.n10 VTAIL.t10 45.5635
R23 VTAIL.n9 VTAIL.n8 44.4112
R24 VTAIL.n6 VTAIL.n5 44.4112
R25 VTAIL.n1 VTAIL.n0 44.4109
R26 VTAIL.n4 VTAIL.n3 44.4109
R27 VTAIL.n6 VTAIL.n4 28.6945
R28 VTAIL.n11 VTAIL.n10 27.9358
R29 VTAIL.n0 VTAIL.t0 1.153
R30 VTAIL.n0 VTAIL.t11 1.153
R31 VTAIL.n3 VTAIL.t8 1.153
R32 VTAIL.n3 VTAIL.t6 1.153
R33 VTAIL.n8 VTAIL.t7 1.153
R34 VTAIL.n8 VTAIL.t5 1.153
R35 VTAIL.n5 VTAIL.t2 1.153
R36 VTAIL.n5 VTAIL.t1 1.153
R37 VTAIL.n9 VTAIL.n7 0.849638
R38 VTAIL.n2 VTAIL.n1 0.849638
R39 VTAIL.n7 VTAIL.n6 0.759121
R40 VTAIL.n10 VTAIL.n9 0.759121
R41 VTAIL.n4 VTAIL.n2 0.759121
R42 VTAIL VTAIL.n11 0.511276
R43 VTAIL VTAIL.n1 0.248345
R44 VDD1 VDD1.t0 62.8695
R45 VDD1.n1 VDD1.t1 62.7559
R46 VDD1.n1 VDD1.n0 61.224
R47 VDD1.n3 VDD1.n2 61.0898
R48 VDD1.n3 VDD1.n1 41.9535
R49 VDD1.n2 VDD1.t4 1.153
R50 VDD1.n2 VDD1.t3 1.153
R51 VDD1.n0 VDD1.t2 1.153
R52 VDD1.n0 VDD1.t5 1.153
R53 VDD1 VDD1.n3 0.131966
R54 B.n67 B.t6 958.11
R55 B.n73 B.t17 958.11
R56 B.n176 B.t10 958.11
R57 B.n168 B.t14 958.11
R58 B.n531 B.n104 585
R59 B.n104 B.n37 585
R60 B.n533 B.n532 585
R61 B.n535 B.n103 585
R62 B.n538 B.n537 585
R63 B.n539 B.n102 585
R64 B.n541 B.n540 585
R65 B.n543 B.n101 585
R66 B.n546 B.n545 585
R67 B.n547 B.n100 585
R68 B.n549 B.n548 585
R69 B.n551 B.n99 585
R70 B.n554 B.n553 585
R71 B.n555 B.n98 585
R72 B.n557 B.n556 585
R73 B.n559 B.n97 585
R74 B.n562 B.n561 585
R75 B.n563 B.n96 585
R76 B.n565 B.n564 585
R77 B.n567 B.n95 585
R78 B.n570 B.n569 585
R79 B.n571 B.n94 585
R80 B.n573 B.n572 585
R81 B.n575 B.n93 585
R82 B.n578 B.n577 585
R83 B.n579 B.n92 585
R84 B.n581 B.n580 585
R85 B.n583 B.n91 585
R86 B.n586 B.n585 585
R87 B.n587 B.n90 585
R88 B.n589 B.n588 585
R89 B.n591 B.n89 585
R90 B.n594 B.n593 585
R91 B.n595 B.n88 585
R92 B.n597 B.n596 585
R93 B.n599 B.n87 585
R94 B.n602 B.n601 585
R95 B.n603 B.n86 585
R96 B.n605 B.n604 585
R97 B.n607 B.n85 585
R98 B.n610 B.n609 585
R99 B.n611 B.n84 585
R100 B.n613 B.n612 585
R101 B.n615 B.n83 585
R102 B.n618 B.n617 585
R103 B.n619 B.n82 585
R104 B.n621 B.n620 585
R105 B.n623 B.n81 585
R106 B.n626 B.n625 585
R107 B.n627 B.n80 585
R108 B.n629 B.n628 585
R109 B.n631 B.n79 585
R110 B.n634 B.n633 585
R111 B.n635 B.n78 585
R112 B.n637 B.n636 585
R113 B.n639 B.n77 585
R114 B.n641 B.n640 585
R115 B.n643 B.n642 585
R116 B.n646 B.n645 585
R117 B.n647 B.n72 585
R118 B.n649 B.n648 585
R119 B.n651 B.n71 585
R120 B.n654 B.n653 585
R121 B.n655 B.n70 585
R122 B.n657 B.n656 585
R123 B.n659 B.n69 585
R124 B.n662 B.n661 585
R125 B.n664 B.n66 585
R126 B.n666 B.n665 585
R127 B.n668 B.n65 585
R128 B.n671 B.n670 585
R129 B.n672 B.n64 585
R130 B.n674 B.n673 585
R131 B.n676 B.n63 585
R132 B.n679 B.n678 585
R133 B.n680 B.n62 585
R134 B.n682 B.n681 585
R135 B.n684 B.n61 585
R136 B.n687 B.n686 585
R137 B.n688 B.n60 585
R138 B.n690 B.n689 585
R139 B.n692 B.n59 585
R140 B.n695 B.n694 585
R141 B.n696 B.n58 585
R142 B.n698 B.n697 585
R143 B.n700 B.n57 585
R144 B.n703 B.n702 585
R145 B.n704 B.n56 585
R146 B.n706 B.n705 585
R147 B.n708 B.n55 585
R148 B.n711 B.n710 585
R149 B.n712 B.n54 585
R150 B.n714 B.n713 585
R151 B.n716 B.n53 585
R152 B.n719 B.n718 585
R153 B.n720 B.n52 585
R154 B.n722 B.n721 585
R155 B.n724 B.n51 585
R156 B.n727 B.n726 585
R157 B.n728 B.n50 585
R158 B.n730 B.n729 585
R159 B.n732 B.n49 585
R160 B.n735 B.n734 585
R161 B.n736 B.n48 585
R162 B.n738 B.n737 585
R163 B.n740 B.n47 585
R164 B.n743 B.n742 585
R165 B.n744 B.n46 585
R166 B.n746 B.n745 585
R167 B.n748 B.n45 585
R168 B.n751 B.n750 585
R169 B.n752 B.n44 585
R170 B.n754 B.n753 585
R171 B.n756 B.n43 585
R172 B.n759 B.n758 585
R173 B.n760 B.n42 585
R174 B.n762 B.n761 585
R175 B.n764 B.n41 585
R176 B.n767 B.n766 585
R177 B.n768 B.n40 585
R178 B.n770 B.n769 585
R179 B.n772 B.n39 585
R180 B.n775 B.n774 585
R181 B.n776 B.n38 585
R182 B.n530 B.n36 585
R183 B.n779 B.n36 585
R184 B.n529 B.n35 585
R185 B.n780 B.n35 585
R186 B.n528 B.n34 585
R187 B.n781 B.n34 585
R188 B.n527 B.n526 585
R189 B.n526 B.n30 585
R190 B.n525 B.n29 585
R191 B.n787 B.n29 585
R192 B.n524 B.n28 585
R193 B.n788 B.n28 585
R194 B.n523 B.n27 585
R195 B.n789 B.n27 585
R196 B.n522 B.n521 585
R197 B.n521 B.n23 585
R198 B.n520 B.n22 585
R199 B.n795 B.n22 585
R200 B.n519 B.n21 585
R201 B.n796 B.n21 585
R202 B.n518 B.n20 585
R203 B.n797 B.n20 585
R204 B.n517 B.n516 585
R205 B.n516 B.n16 585
R206 B.n515 B.n15 585
R207 B.n803 B.n15 585
R208 B.n514 B.n14 585
R209 B.n804 B.n14 585
R210 B.n513 B.n13 585
R211 B.n805 B.n13 585
R212 B.n512 B.n511 585
R213 B.n511 B.n12 585
R214 B.n510 B.n509 585
R215 B.n510 B.n8 585
R216 B.n508 B.n7 585
R217 B.n812 B.n7 585
R218 B.n507 B.n6 585
R219 B.n813 B.n6 585
R220 B.n506 B.n5 585
R221 B.n814 B.n5 585
R222 B.n505 B.n504 585
R223 B.n504 B.n4 585
R224 B.n503 B.n105 585
R225 B.n503 B.n502 585
R226 B.n492 B.n106 585
R227 B.n495 B.n106 585
R228 B.n494 B.n493 585
R229 B.n496 B.n494 585
R230 B.n491 B.n110 585
R231 B.n114 B.n110 585
R232 B.n490 B.n489 585
R233 B.n489 B.n488 585
R234 B.n112 B.n111 585
R235 B.n113 B.n112 585
R236 B.n481 B.n480 585
R237 B.n482 B.n481 585
R238 B.n479 B.n119 585
R239 B.n119 B.n118 585
R240 B.n478 B.n477 585
R241 B.n477 B.n476 585
R242 B.n121 B.n120 585
R243 B.n122 B.n121 585
R244 B.n469 B.n468 585
R245 B.n470 B.n469 585
R246 B.n467 B.n127 585
R247 B.n127 B.n126 585
R248 B.n466 B.n465 585
R249 B.n465 B.n464 585
R250 B.n129 B.n128 585
R251 B.n130 B.n129 585
R252 B.n457 B.n456 585
R253 B.n458 B.n457 585
R254 B.n455 B.n135 585
R255 B.n135 B.n134 585
R256 B.n454 B.n453 585
R257 B.n453 B.n452 585
R258 B.n449 B.n139 585
R259 B.n448 B.n447 585
R260 B.n445 B.n140 585
R261 B.n445 B.n138 585
R262 B.n444 B.n443 585
R263 B.n442 B.n441 585
R264 B.n440 B.n142 585
R265 B.n438 B.n437 585
R266 B.n436 B.n143 585
R267 B.n435 B.n434 585
R268 B.n432 B.n144 585
R269 B.n430 B.n429 585
R270 B.n428 B.n145 585
R271 B.n427 B.n426 585
R272 B.n424 B.n146 585
R273 B.n422 B.n421 585
R274 B.n420 B.n147 585
R275 B.n419 B.n418 585
R276 B.n416 B.n148 585
R277 B.n414 B.n413 585
R278 B.n412 B.n149 585
R279 B.n411 B.n410 585
R280 B.n408 B.n150 585
R281 B.n406 B.n405 585
R282 B.n404 B.n151 585
R283 B.n403 B.n402 585
R284 B.n400 B.n152 585
R285 B.n398 B.n397 585
R286 B.n396 B.n153 585
R287 B.n395 B.n394 585
R288 B.n392 B.n154 585
R289 B.n390 B.n389 585
R290 B.n388 B.n155 585
R291 B.n387 B.n386 585
R292 B.n384 B.n156 585
R293 B.n382 B.n381 585
R294 B.n380 B.n157 585
R295 B.n379 B.n378 585
R296 B.n376 B.n158 585
R297 B.n374 B.n373 585
R298 B.n372 B.n159 585
R299 B.n371 B.n370 585
R300 B.n368 B.n160 585
R301 B.n366 B.n365 585
R302 B.n364 B.n161 585
R303 B.n363 B.n362 585
R304 B.n360 B.n162 585
R305 B.n358 B.n357 585
R306 B.n356 B.n163 585
R307 B.n355 B.n354 585
R308 B.n352 B.n164 585
R309 B.n350 B.n349 585
R310 B.n348 B.n165 585
R311 B.n347 B.n346 585
R312 B.n344 B.n166 585
R313 B.n342 B.n341 585
R314 B.n340 B.n167 585
R315 B.n339 B.n338 585
R316 B.n336 B.n335 585
R317 B.n334 B.n333 585
R318 B.n332 B.n172 585
R319 B.n330 B.n329 585
R320 B.n328 B.n173 585
R321 B.n327 B.n326 585
R322 B.n324 B.n174 585
R323 B.n322 B.n321 585
R324 B.n320 B.n175 585
R325 B.n318 B.n317 585
R326 B.n315 B.n178 585
R327 B.n313 B.n312 585
R328 B.n311 B.n179 585
R329 B.n310 B.n309 585
R330 B.n307 B.n180 585
R331 B.n305 B.n304 585
R332 B.n303 B.n181 585
R333 B.n302 B.n301 585
R334 B.n299 B.n182 585
R335 B.n297 B.n296 585
R336 B.n295 B.n183 585
R337 B.n294 B.n293 585
R338 B.n291 B.n184 585
R339 B.n289 B.n288 585
R340 B.n287 B.n185 585
R341 B.n286 B.n285 585
R342 B.n283 B.n186 585
R343 B.n281 B.n280 585
R344 B.n279 B.n187 585
R345 B.n278 B.n277 585
R346 B.n275 B.n188 585
R347 B.n273 B.n272 585
R348 B.n271 B.n189 585
R349 B.n270 B.n269 585
R350 B.n267 B.n190 585
R351 B.n265 B.n264 585
R352 B.n263 B.n191 585
R353 B.n262 B.n261 585
R354 B.n259 B.n192 585
R355 B.n257 B.n256 585
R356 B.n255 B.n193 585
R357 B.n254 B.n253 585
R358 B.n251 B.n194 585
R359 B.n249 B.n248 585
R360 B.n247 B.n195 585
R361 B.n246 B.n245 585
R362 B.n243 B.n196 585
R363 B.n241 B.n240 585
R364 B.n239 B.n197 585
R365 B.n238 B.n237 585
R366 B.n235 B.n198 585
R367 B.n233 B.n232 585
R368 B.n231 B.n199 585
R369 B.n230 B.n229 585
R370 B.n227 B.n200 585
R371 B.n225 B.n224 585
R372 B.n223 B.n201 585
R373 B.n222 B.n221 585
R374 B.n219 B.n202 585
R375 B.n217 B.n216 585
R376 B.n215 B.n203 585
R377 B.n214 B.n213 585
R378 B.n211 B.n204 585
R379 B.n209 B.n208 585
R380 B.n207 B.n206 585
R381 B.n137 B.n136 585
R382 B.n451 B.n450 585
R383 B.n452 B.n451 585
R384 B.n133 B.n132 585
R385 B.n134 B.n133 585
R386 B.n460 B.n459 585
R387 B.n459 B.n458 585
R388 B.n461 B.n131 585
R389 B.n131 B.n130 585
R390 B.n463 B.n462 585
R391 B.n464 B.n463 585
R392 B.n125 B.n124 585
R393 B.n126 B.n125 585
R394 B.n472 B.n471 585
R395 B.n471 B.n470 585
R396 B.n473 B.n123 585
R397 B.n123 B.n122 585
R398 B.n475 B.n474 585
R399 B.n476 B.n475 585
R400 B.n117 B.n116 585
R401 B.n118 B.n117 585
R402 B.n484 B.n483 585
R403 B.n483 B.n482 585
R404 B.n485 B.n115 585
R405 B.n115 B.n113 585
R406 B.n487 B.n486 585
R407 B.n488 B.n487 585
R408 B.n109 B.n108 585
R409 B.n114 B.n109 585
R410 B.n498 B.n497 585
R411 B.n497 B.n496 585
R412 B.n499 B.n107 585
R413 B.n495 B.n107 585
R414 B.n501 B.n500 585
R415 B.n502 B.n501 585
R416 B.n3 B.n0 585
R417 B.n4 B.n3 585
R418 B.n811 B.n1 585
R419 B.n812 B.n811 585
R420 B.n810 B.n809 585
R421 B.n810 B.n8 585
R422 B.n808 B.n9 585
R423 B.n12 B.n9 585
R424 B.n807 B.n806 585
R425 B.n806 B.n805 585
R426 B.n11 B.n10 585
R427 B.n804 B.n11 585
R428 B.n802 B.n801 585
R429 B.n803 B.n802 585
R430 B.n800 B.n17 585
R431 B.n17 B.n16 585
R432 B.n799 B.n798 585
R433 B.n798 B.n797 585
R434 B.n19 B.n18 585
R435 B.n796 B.n19 585
R436 B.n794 B.n793 585
R437 B.n795 B.n794 585
R438 B.n792 B.n24 585
R439 B.n24 B.n23 585
R440 B.n791 B.n790 585
R441 B.n790 B.n789 585
R442 B.n26 B.n25 585
R443 B.n788 B.n26 585
R444 B.n786 B.n785 585
R445 B.n787 B.n786 585
R446 B.n784 B.n31 585
R447 B.n31 B.n30 585
R448 B.n783 B.n782 585
R449 B.n782 B.n781 585
R450 B.n33 B.n32 585
R451 B.n780 B.n33 585
R452 B.n778 B.n777 585
R453 B.n779 B.n778 585
R454 B.n815 B.n814 585
R455 B.n813 B.n2 585
R456 B.n778 B.n38 516.524
R457 B.n104 B.n36 516.524
R458 B.n453 B.n137 516.524
R459 B.n451 B.n139 516.524
R460 B.n534 B.n37 256.663
R461 B.n536 B.n37 256.663
R462 B.n542 B.n37 256.663
R463 B.n544 B.n37 256.663
R464 B.n550 B.n37 256.663
R465 B.n552 B.n37 256.663
R466 B.n558 B.n37 256.663
R467 B.n560 B.n37 256.663
R468 B.n566 B.n37 256.663
R469 B.n568 B.n37 256.663
R470 B.n574 B.n37 256.663
R471 B.n576 B.n37 256.663
R472 B.n582 B.n37 256.663
R473 B.n584 B.n37 256.663
R474 B.n590 B.n37 256.663
R475 B.n592 B.n37 256.663
R476 B.n598 B.n37 256.663
R477 B.n600 B.n37 256.663
R478 B.n606 B.n37 256.663
R479 B.n608 B.n37 256.663
R480 B.n614 B.n37 256.663
R481 B.n616 B.n37 256.663
R482 B.n622 B.n37 256.663
R483 B.n624 B.n37 256.663
R484 B.n630 B.n37 256.663
R485 B.n632 B.n37 256.663
R486 B.n638 B.n37 256.663
R487 B.n76 B.n37 256.663
R488 B.n644 B.n37 256.663
R489 B.n650 B.n37 256.663
R490 B.n652 B.n37 256.663
R491 B.n658 B.n37 256.663
R492 B.n660 B.n37 256.663
R493 B.n667 B.n37 256.663
R494 B.n669 B.n37 256.663
R495 B.n675 B.n37 256.663
R496 B.n677 B.n37 256.663
R497 B.n683 B.n37 256.663
R498 B.n685 B.n37 256.663
R499 B.n691 B.n37 256.663
R500 B.n693 B.n37 256.663
R501 B.n699 B.n37 256.663
R502 B.n701 B.n37 256.663
R503 B.n707 B.n37 256.663
R504 B.n709 B.n37 256.663
R505 B.n715 B.n37 256.663
R506 B.n717 B.n37 256.663
R507 B.n723 B.n37 256.663
R508 B.n725 B.n37 256.663
R509 B.n731 B.n37 256.663
R510 B.n733 B.n37 256.663
R511 B.n739 B.n37 256.663
R512 B.n741 B.n37 256.663
R513 B.n747 B.n37 256.663
R514 B.n749 B.n37 256.663
R515 B.n755 B.n37 256.663
R516 B.n757 B.n37 256.663
R517 B.n763 B.n37 256.663
R518 B.n765 B.n37 256.663
R519 B.n771 B.n37 256.663
R520 B.n773 B.n37 256.663
R521 B.n446 B.n138 256.663
R522 B.n141 B.n138 256.663
R523 B.n439 B.n138 256.663
R524 B.n433 B.n138 256.663
R525 B.n431 B.n138 256.663
R526 B.n425 B.n138 256.663
R527 B.n423 B.n138 256.663
R528 B.n417 B.n138 256.663
R529 B.n415 B.n138 256.663
R530 B.n409 B.n138 256.663
R531 B.n407 B.n138 256.663
R532 B.n401 B.n138 256.663
R533 B.n399 B.n138 256.663
R534 B.n393 B.n138 256.663
R535 B.n391 B.n138 256.663
R536 B.n385 B.n138 256.663
R537 B.n383 B.n138 256.663
R538 B.n377 B.n138 256.663
R539 B.n375 B.n138 256.663
R540 B.n369 B.n138 256.663
R541 B.n367 B.n138 256.663
R542 B.n361 B.n138 256.663
R543 B.n359 B.n138 256.663
R544 B.n353 B.n138 256.663
R545 B.n351 B.n138 256.663
R546 B.n345 B.n138 256.663
R547 B.n343 B.n138 256.663
R548 B.n337 B.n138 256.663
R549 B.n171 B.n138 256.663
R550 B.n331 B.n138 256.663
R551 B.n325 B.n138 256.663
R552 B.n323 B.n138 256.663
R553 B.n316 B.n138 256.663
R554 B.n314 B.n138 256.663
R555 B.n308 B.n138 256.663
R556 B.n306 B.n138 256.663
R557 B.n300 B.n138 256.663
R558 B.n298 B.n138 256.663
R559 B.n292 B.n138 256.663
R560 B.n290 B.n138 256.663
R561 B.n284 B.n138 256.663
R562 B.n282 B.n138 256.663
R563 B.n276 B.n138 256.663
R564 B.n274 B.n138 256.663
R565 B.n268 B.n138 256.663
R566 B.n266 B.n138 256.663
R567 B.n260 B.n138 256.663
R568 B.n258 B.n138 256.663
R569 B.n252 B.n138 256.663
R570 B.n250 B.n138 256.663
R571 B.n244 B.n138 256.663
R572 B.n242 B.n138 256.663
R573 B.n236 B.n138 256.663
R574 B.n234 B.n138 256.663
R575 B.n228 B.n138 256.663
R576 B.n226 B.n138 256.663
R577 B.n220 B.n138 256.663
R578 B.n218 B.n138 256.663
R579 B.n212 B.n138 256.663
R580 B.n210 B.n138 256.663
R581 B.n205 B.n138 256.663
R582 B.n817 B.n816 256.663
R583 B.n774 B.n772 163.367
R584 B.n770 B.n40 163.367
R585 B.n766 B.n764 163.367
R586 B.n762 B.n42 163.367
R587 B.n758 B.n756 163.367
R588 B.n754 B.n44 163.367
R589 B.n750 B.n748 163.367
R590 B.n746 B.n46 163.367
R591 B.n742 B.n740 163.367
R592 B.n738 B.n48 163.367
R593 B.n734 B.n732 163.367
R594 B.n730 B.n50 163.367
R595 B.n726 B.n724 163.367
R596 B.n722 B.n52 163.367
R597 B.n718 B.n716 163.367
R598 B.n714 B.n54 163.367
R599 B.n710 B.n708 163.367
R600 B.n706 B.n56 163.367
R601 B.n702 B.n700 163.367
R602 B.n698 B.n58 163.367
R603 B.n694 B.n692 163.367
R604 B.n690 B.n60 163.367
R605 B.n686 B.n684 163.367
R606 B.n682 B.n62 163.367
R607 B.n678 B.n676 163.367
R608 B.n674 B.n64 163.367
R609 B.n670 B.n668 163.367
R610 B.n666 B.n66 163.367
R611 B.n661 B.n659 163.367
R612 B.n657 B.n70 163.367
R613 B.n653 B.n651 163.367
R614 B.n649 B.n72 163.367
R615 B.n645 B.n643 163.367
R616 B.n640 B.n639 163.367
R617 B.n637 B.n78 163.367
R618 B.n633 B.n631 163.367
R619 B.n629 B.n80 163.367
R620 B.n625 B.n623 163.367
R621 B.n621 B.n82 163.367
R622 B.n617 B.n615 163.367
R623 B.n613 B.n84 163.367
R624 B.n609 B.n607 163.367
R625 B.n605 B.n86 163.367
R626 B.n601 B.n599 163.367
R627 B.n597 B.n88 163.367
R628 B.n593 B.n591 163.367
R629 B.n589 B.n90 163.367
R630 B.n585 B.n583 163.367
R631 B.n581 B.n92 163.367
R632 B.n577 B.n575 163.367
R633 B.n573 B.n94 163.367
R634 B.n569 B.n567 163.367
R635 B.n565 B.n96 163.367
R636 B.n561 B.n559 163.367
R637 B.n557 B.n98 163.367
R638 B.n553 B.n551 163.367
R639 B.n549 B.n100 163.367
R640 B.n545 B.n543 163.367
R641 B.n541 B.n102 163.367
R642 B.n537 B.n535 163.367
R643 B.n533 B.n104 163.367
R644 B.n453 B.n135 163.367
R645 B.n457 B.n135 163.367
R646 B.n457 B.n129 163.367
R647 B.n465 B.n129 163.367
R648 B.n465 B.n127 163.367
R649 B.n469 B.n127 163.367
R650 B.n469 B.n121 163.367
R651 B.n477 B.n121 163.367
R652 B.n477 B.n119 163.367
R653 B.n481 B.n119 163.367
R654 B.n481 B.n112 163.367
R655 B.n489 B.n112 163.367
R656 B.n489 B.n110 163.367
R657 B.n494 B.n110 163.367
R658 B.n494 B.n106 163.367
R659 B.n503 B.n106 163.367
R660 B.n504 B.n503 163.367
R661 B.n504 B.n5 163.367
R662 B.n6 B.n5 163.367
R663 B.n7 B.n6 163.367
R664 B.n510 B.n7 163.367
R665 B.n511 B.n510 163.367
R666 B.n511 B.n13 163.367
R667 B.n14 B.n13 163.367
R668 B.n15 B.n14 163.367
R669 B.n516 B.n15 163.367
R670 B.n516 B.n20 163.367
R671 B.n21 B.n20 163.367
R672 B.n22 B.n21 163.367
R673 B.n521 B.n22 163.367
R674 B.n521 B.n27 163.367
R675 B.n28 B.n27 163.367
R676 B.n29 B.n28 163.367
R677 B.n526 B.n29 163.367
R678 B.n526 B.n34 163.367
R679 B.n35 B.n34 163.367
R680 B.n36 B.n35 163.367
R681 B.n447 B.n445 163.367
R682 B.n445 B.n444 163.367
R683 B.n441 B.n440 163.367
R684 B.n438 B.n143 163.367
R685 B.n434 B.n432 163.367
R686 B.n430 B.n145 163.367
R687 B.n426 B.n424 163.367
R688 B.n422 B.n147 163.367
R689 B.n418 B.n416 163.367
R690 B.n414 B.n149 163.367
R691 B.n410 B.n408 163.367
R692 B.n406 B.n151 163.367
R693 B.n402 B.n400 163.367
R694 B.n398 B.n153 163.367
R695 B.n394 B.n392 163.367
R696 B.n390 B.n155 163.367
R697 B.n386 B.n384 163.367
R698 B.n382 B.n157 163.367
R699 B.n378 B.n376 163.367
R700 B.n374 B.n159 163.367
R701 B.n370 B.n368 163.367
R702 B.n366 B.n161 163.367
R703 B.n362 B.n360 163.367
R704 B.n358 B.n163 163.367
R705 B.n354 B.n352 163.367
R706 B.n350 B.n165 163.367
R707 B.n346 B.n344 163.367
R708 B.n342 B.n167 163.367
R709 B.n338 B.n336 163.367
R710 B.n333 B.n332 163.367
R711 B.n330 B.n173 163.367
R712 B.n326 B.n324 163.367
R713 B.n322 B.n175 163.367
R714 B.n317 B.n315 163.367
R715 B.n313 B.n179 163.367
R716 B.n309 B.n307 163.367
R717 B.n305 B.n181 163.367
R718 B.n301 B.n299 163.367
R719 B.n297 B.n183 163.367
R720 B.n293 B.n291 163.367
R721 B.n289 B.n185 163.367
R722 B.n285 B.n283 163.367
R723 B.n281 B.n187 163.367
R724 B.n277 B.n275 163.367
R725 B.n273 B.n189 163.367
R726 B.n269 B.n267 163.367
R727 B.n265 B.n191 163.367
R728 B.n261 B.n259 163.367
R729 B.n257 B.n193 163.367
R730 B.n253 B.n251 163.367
R731 B.n249 B.n195 163.367
R732 B.n245 B.n243 163.367
R733 B.n241 B.n197 163.367
R734 B.n237 B.n235 163.367
R735 B.n233 B.n199 163.367
R736 B.n229 B.n227 163.367
R737 B.n225 B.n201 163.367
R738 B.n221 B.n219 163.367
R739 B.n217 B.n203 163.367
R740 B.n213 B.n211 163.367
R741 B.n209 B.n206 163.367
R742 B.n451 B.n133 163.367
R743 B.n459 B.n133 163.367
R744 B.n459 B.n131 163.367
R745 B.n463 B.n131 163.367
R746 B.n463 B.n125 163.367
R747 B.n471 B.n125 163.367
R748 B.n471 B.n123 163.367
R749 B.n475 B.n123 163.367
R750 B.n475 B.n117 163.367
R751 B.n483 B.n117 163.367
R752 B.n483 B.n115 163.367
R753 B.n487 B.n115 163.367
R754 B.n487 B.n109 163.367
R755 B.n497 B.n109 163.367
R756 B.n497 B.n107 163.367
R757 B.n501 B.n107 163.367
R758 B.n501 B.n3 163.367
R759 B.n815 B.n3 163.367
R760 B.n811 B.n2 163.367
R761 B.n811 B.n810 163.367
R762 B.n810 B.n9 163.367
R763 B.n806 B.n9 163.367
R764 B.n806 B.n11 163.367
R765 B.n802 B.n11 163.367
R766 B.n802 B.n17 163.367
R767 B.n798 B.n17 163.367
R768 B.n798 B.n19 163.367
R769 B.n794 B.n19 163.367
R770 B.n794 B.n24 163.367
R771 B.n790 B.n24 163.367
R772 B.n790 B.n26 163.367
R773 B.n786 B.n26 163.367
R774 B.n786 B.n31 163.367
R775 B.n782 B.n31 163.367
R776 B.n782 B.n33 163.367
R777 B.n778 B.n33 163.367
R778 B.n73 B.t18 87.8575
R779 B.n176 B.t13 87.8575
R780 B.n67 B.t8 87.8347
R781 B.n168 B.t16 87.8347
R782 B.n773 B.n38 71.676
R783 B.n772 B.n771 71.676
R784 B.n765 B.n40 71.676
R785 B.n764 B.n763 71.676
R786 B.n757 B.n42 71.676
R787 B.n756 B.n755 71.676
R788 B.n749 B.n44 71.676
R789 B.n748 B.n747 71.676
R790 B.n741 B.n46 71.676
R791 B.n740 B.n739 71.676
R792 B.n733 B.n48 71.676
R793 B.n732 B.n731 71.676
R794 B.n725 B.n50 71.676
R795 B.n724 B.n723 71.676
R796 B.n717 B.n52 71.676
R797 B.n716 B.n715 71.676
R798 B.n709 B.n54 71.676
R799 B.n708 B.n707 71.676
R800 B.n701 B.n56 71.676
R801 B.n700 B.n699 71.676
R802 B.n693 B.n58 71.676
R803 B.n692 B.n691 71.676
R804 B.n685 B.n60 71.676
R805 B.n684 B.n683 71.676
R806 B.n677 B.n62 71.676
R807 B.n676 B.n675 71.676
R808 B.n669 B.n64 71.676
R809 B.n668 B.n667 71.676
R810 B.n660 B.n66 71.676
R811 B.n659 B.n658 71.676
R812 B.n652 B.n70 71.676
R813 B.n651 B.n650 71.676
R814 B.n644 B.n72 71.676
R815 B.n643 B.n76 71.676
R816 B.n639 B.n638 71.676
R817 B.n632 B.n78 71.676
R818 B.n631 B.n630 71.676
R819 B.n624 B.n80 71.676
R820 B.n623 B.n622 71.676
R821 B.n616 B.n82 71.676
R822 B.n615 B.n614 71.676
R823 B.n608 B.n84 71.676
R824 B.n607 B.n606 71.676
R825 B.n600 B.n86 71.676
R826 B.n599 B.n598 71.676
R827 B.n592 B.n88 71.676
R828 B.n591 B.n590 71.676
R829 B.n584 B.n90 71.676
R830 B.n583 B.n582 71.676
R831 B.n576 B.n92 71.676
R832 B.n575 B.n574 71.676
R833 B.n568 B.n94 71.676
R834 B.n567 B.n566 71.676
R835 B.n560 B.n96 71.676
R836 B.n559 B.n558 71.676
R837 B.n552 B.n98 71.676
R838 B.n551 B.n550 71.676
R839 B.n544 B.n100 71.676
R840 B.n543 B.n542 71.676
R841 B.n536 B.n102 71.676
R842 B.n535 B.n534 71.676
R843 B.n534 B.n533 71.676
R844 B.n537 B.n536 71.676
R845 B.n542 B.n541 71.676
R846 B.n545 B.n544 71.676
R847 B.n550 B.n549 71.676
R848 B.n553 B.n552 71.676
R849 B.n558 B.n557 71.676
R850 B.n561 B.n560 71.676
R851 B.n566 B.n565 71.676
R852 B.n569 B.n568 71.676
R853 B.n574 B.n573 71.676
R854 B.n577 B.n576 71.676
R855 B.n582 B.n581 71.676
R856 B.n585 B.n584 71.676
R857 B.n590 B.n589 71.676
R858 B.n593 B.n592 71.676
R859 B.n598 B.n597 71.676
R860 B.n601 B.n600 71.676
R861 B.n606 B.n605 71.676
R862 B.n609 B.n608 71.676
R863 B.n614 B.n613 71.676
R864 B.n617 B.n616 71.676
R865 B.n622 B.n621 71.676
R866 B.n625 B.n624 71.676
R867 B.n630 B.n629 71.676
R868 B.n633 B.n632 71.676
R869 B.n638 B.n637 71.676
R870 B.n640 B.n76 71.676
R871 B.n645 B.n644 71.676
R872 B.n650 B.n649 71.676
R873 B.n653 B.n652 71.676
R874 B.n658 B.n657 71.676
R875 B.n661 B.n660 71.676
R876 B.n667 B.n666 71.676
R877 B.n670 B.n669 71.676
R878 B.n675 B.n674 71.676
R879 B.n678 B.n677 71.676
R880 B.n683 B.n682 71.676
R881 B.n686 B.n685 71.676
R882 B.n691 B.n690 71.676
R883 B.n694 B.n693 71.676
R884 B.n699 B.n698 71.676
R885 B.n702 B.n701 71.676
R886 B.n707 B.n706 71.676
R887 B.n710 B.n709 71.676
R888 B.n715 B.n714 71.676
R889 B.n718 B.n717 71.676
R890 B.n723 B.n722 71.676
R891 B.n726 B.n725 71.676
R892 B.n731 B.n730 71.676
R893 B.n734 B.n733 71.676
R894 B.n739 B.n738 71.676
R895 B.n742 B.n741 71.676
R896 B.n747 B.n746 71.676
R897 B.n750 B.n749 71.676
R898 B.n755 B.n754 71.676
R899 B.n758 B.n757 71.676
R900 B.n763 B.n762 71.676
R901 B.n766 B.n765 71.676
R902 B.n771 B.n770 71.676
R903 B.n774 B.n773 71.676
R904 B.n446 B.n139 71.676
R905 B.n444 B.n141 71.676
R906 B.n440 B.n439 71.676
R907 B.n433 B.n143 71.676
R908 B.n432 B.n431 71.676
R909 B.n425 B.n145 71.676
R910 B.n424 B.n423 71.676
R911 B.n417 B.n147 71.676
R912 B.n416 B.n415 71.676
R913 B.n409 B.n149 71.676
R914 B.n408 B.n407 71.676
R915 B.n401 B.n151 71.676
R916 B.n400 B.n399 71.676
R917 B.n393 B.n153 71.676
R918 B.n392 B.n391 71.676
R919 B.n385 B.n155 71.676
R920 B.n384 B.n383 71.676
R921 B.n377 B.n157 71.676
R922 B.n376 B.n375 71.676
R923 B.n369 B.n159 71.676
R924 B.n368 B.n367 71.676
R925 B.n361 B.n161 71.676
R926 B.n360 B.n359 71.676
R927 B.n353 B.n163 71.676
R928 B.n352 B.n351 71.676
R929 B.n345 B.n165 71.676
R930 B.n344 B.n343 71.676
R931 B.n337 B.n167 71.676
R932 B.n336 B.n171 71.676
R933 B.n332 B.n331 71.676
R934 B.n325 B.n173 71.676
R935 B.n324 B.n323 71.676
R936 B.n316 B.n175 71.676
R937 B.n315 B.n314 71.676
R938 B.n308 B.n179 71.676
R939 B.n307 B.n306 71.676
R940 B.n300 B.n181 71.676
R941 B.n299 B.n298 71.676
R942 B.n292 B.n183 71.676
R943 B.n291 B.n290 71.676
R944 B.n284 B.n185 71.676
R945 B.n283 B.n282 71.676
R946 B.n276 B.n187 71.676
R947 B.n275 B.n274 71.676
R948 B.n268 B.n189 71.676
R949 B.n267 B.n266 71.676
R950 B.n260 B.n191 71.676
R951 B.n259 B.n258 71.676
R952 B.n252 B.n193 71.676
R953 B.n251 B.n250 71.676
R954 B.n244 B.n195 71.676
R955 B.n243 B.n242 71.676
R956 B.n236 B.n197 71.676
R957 B.n235 B.n234 71.676
R958 B.n228 B.n199 71.676
R959 B.n227 B.n226 71.676
R960 B.n220 B.n201 71.676
R961 B.n219 B.n218 71.676
R962 B.n212 B.n203 71.676
R963 B.n211 B.n210 71.676
R964 B.n206 B.n205 71.676
R965 B.n447 B.n446 71.676
R966 B.n441 B.n141 71.676
R967 B.n439 B.n438 71.676
R968 B.n434 B.n433 71.676
R969 B.n431 B.n430 71.676
R970 B.n426 B.n425 71.676
R971 B.n423 B.n422 71.676
R972 B.n418 B.n417 71.676
R973 B.n415 B.n414 71.676
R974 B.n410 B.n409 71.676
R975 B.n407 B.n406 71.676
R976 B.n402 B.n401 71.676
R977 B.n399 B.n398 71.676
R978 B.n394 B.n393 71.676
R979 B.n391 B.n390 71.676
R980 B.n386 B.n385 71.676
R981 B.n383 B.n382 71.676
R982 B.n378 B.n377 71.676
R983 B.n375 B.n374 71.676
R984 B.n370 B.n369 71.676
R985 B.n367 B.n366 71.676
R986 B.n362 B.n361 71.676
R987 B.n359 B.n358 71.676
R988 B.n354 B.n353 71.676
R989 B.n351 B.n350 71.676
R990 B.n346 B.n345 71.676
R991 B.n343 B.n342 71.676
R992 B.n338 B.n337 71.676
R993 B.n333 B.n171 71.676
R994 B.n331 B.n330 71.676
R995 B.n326 B.n325 71.676
R996 B.n323 B.n322 71.676
R997 B.n317 B.n316 71.676
R998 B.n314 B.n313 71.676
R999 B.n309 B.n308 71.676
R1000 B.n306 B.n305 71.676
R1001 B.n301 B.n300 71.676
R1002 B.n298 B.n297 71.676
R1003 B.n293 B.n292 71.676
R1004 B.n290 B.n289 71.676
R1005 B.n285 B.n284 71.676
R1006 B.n282 B.n281 71.676
R1007 B.n277 B.n276 71.676
R1008 B.n274 B.n273 71.676
R1009 B.n269 B.n268 71.676
R1010 B.n266 B.n265 71.676
R1011 B.n261 B.n260 71.676
R1012 B.n258 B.n257 71.676
R1013 B.n253 B.n252 71.676
R1014 B.n250 B.n249 71.676
R1015 B.n245 B.n244 71.676
R1016 B.n242 B.n241 71.676
R1017 B.n237 B.n236 71.676
R1018 B.n234 B.n233 71.676
R1019 B.n229 B.n228 71.676
R1020 B.n226 B.n225 71.676
R1021 B.n221 B.n220 71.676
R1022 B.n218 B.n217 71.676
R1023 B.n213 B.n212 71.676
R1024 B.n210 B.n209 71.676
R1025 B.n205 B.n137 71.676
R1026 B.n816 B.n815 71.676
R1027 B.n816 B.n2 71.676
R1028 B.n74 B.t19 70.7908
R1029 B.n177 B.t12 70.7908
R1030 B.n68 B.t9 70.7681
R1031 B.n169 B.t15 70.7681
R1032 B.n663 B.n68 59.5399
R1033 B.n75 B.n74 59.5399
R1034 B.n319 B.n177 59.5399
R1035 B.n170 B.n169 59.5399
R1036 B.n452 B.n138 59.2746
R1037 B.n779 B.n37 59.2746
R1038 B.n450 B.n449 33.5615
R1039 B.n454 B.n136 33.5615
R1040 B.n531 B.n530 33.5615
R1041 B.n777 B.n776 33.5615
R1042 B.n452 B.n134 33.3116
R1043 B.n458 B.n134 33.3116
R1044 B.n458 B.n130 33.3116
R1045 B.n464 B.n130 33.3116
R1046 B.n470 B.n126 33.3116
R1047 B.n470 B.n122 33.3116
R1048 B.n476 B.n122 33.3116
R1049 B.n476 B.n118 33.3116
R1050 B.n482 B.n118 33.3116
R1051 B.n488 B.n113 33.3116
R1052 B.n488 B.n114 33.3116
R1053 B.n496 B.n495 33.3116
R1054 B.n502 B.n4 33.3116
R1055 B.n814 B.n4 33.3116
R1056 B.n814 B.n813 33.3116
R1057 B.n813 B.n812 33.3116
R1058 B.n812 B.n8 33.3116
R1059 B.n805 B.n12 33.3116
R1060 B.n804 B.n803 33.3116
R1061 B.n803 B.n16 33.3116
R1062 B.n797 B.n796 33.3116
R1063 B.n796 B.n795 33.3116
R1064 B.n795 B.n23 33.3116
R1065 B.n789 B.n23 33.3116
R1066 B.n789 B.n788 33.3116
R1067 B.n787 B.n30 33.3116
R1068 B.n781 B.n30 33.3116
R1069 B.n781 B.n780 33.3116
R1070 B.n780 B.n779 33.3116
R1071 B.n496 B.t1 32.8217
R1072 B.n805 B.t5 32.8217
R1073 B.n464 B.t11 21.0649
R1074 B.t7 B.n787 21.0649
R1075 B.n495 B.t4 20.0851
R1076 B.n12 B.t0 20.0851
R1077 B.t2 B.n113 19.1054
R1078 B.t3 B.n16 19.1054
R1079 B B.n817 18.0485
R1080 B.n68 B.n67 17.0672
R1081 B.n74 B.n73 17.0672
R1082 B.n177 B.n176 17.0672
R1083 B.n169 B.n168 17.0672
R1084 B.n482 B.t2 14.2067
R1085 B.n797 B.t3 14.2067
R1086 B.n502 B.t4 13.227
R1087 B.t0 B.n8 13.227
R1088 B.t11 B.n126 12.2472
R1089 B.n788 B.t7 12.2472
R1090 B.n450 B.n132 10.6151
R1091 B.n460 B.n132 10.6151
R1092 B.n461 B.n460 10.6151
R1093 B.n462 B.n461 10.6151
R1094 B.n462 B.n124 10.6151
R1095 B.n472 B.n124 10.6151
R1096 B.n473 B.n472 10.6151
R1097 B.n474 B.n473 10.6151
R1098 B.n474 B.n116 10.6151
R1099 B.n484 B.n116 10.6151
R1100 B.n485 B.n484 10.6151
R1101 B.n486 B.n485 10.6151
R1102 B.n486 B.n108 10.6151
R1103 B.n498 B.n108 10.6151
R1104 B.n499 B.n498 10.6151
R1105 B.n500 B.n499 10.6151
R1106 B.n500 B.n0 10.6151
R1107 B.n449 B.n448 10.6151
R1108 B.n448 B.n140 10.6151
R1109 B.n443 B.n140 10.6151
R1110 B.n443 B.n442 10.6151
R1111 B.n442 B.n142 10.6151
R1112 B.n437 B.n142 10.6151
R1113 B.n437 B.n436 10.6151
R1114 B.n436 B.n435 10.6151
R1115 B.n435 B.n144 10.6151
R1116 B.n429 B.n144 10.6151
R1117 B.n429 B.n428 10.6151
R1118 B.n428 B.n427 10.6151
R1119 B.n427 B.n146 10.6151
R1120 B.n421 B.n146 10.6151
R1121 B.n421 B.n420 10.6151
R1122 B.n420 B.n419 10.6151
R1123 B.n419 B.n148 10.6151
R1124 B.n413 B.n148 10.6151
R1125 B.n413 B.n412 10.6151
R1126 B.n412 B.n411 10.6151
R1127 B.n411 B.n150 10.6151
R1128 B.n405 B.n150 10.6151
R1129 B.n405 B.n404 10.6151
R1130 B.n404 B.n403 10.6151
R1131 B.n403 B.n152 10.6151
R1132 B.n397 B.n152 10.6151
R1133 B.n397 B.n396 10.6151
R1134 B.n396 B.n395 10.6151
R1135 B.n395 B.n154 10.6151
R1136 B.n389 B.n154 10.6151
R1137 B.n389 B.n388 10.6151
R1138 B.n388 B.n387 10.6151
R1139 B.n387 B.n156 10.6151
R1140 B.n381 B.n156 10.6151
R1141 B.n381 B.n380 10.6151
R1142 B.n380 B.n379 10.6151
R1143 B.n379 B.n158 10.6151
R1144 B.n373 B.n158 10.6151
R1145 B.n373 B.n372 10.6151
R1146 B.n372 B.n371 10.6151
R1147 B.n371 B.n160 10.6151
R1148 B.n365 B.n160 10.6151
R1149 B.n365 B.n364 10.6151
R1150 B.n364 B.n363 10.6151
R1151 B.n363 B.n162 10.6151
R1152 B.n357 B.n162 10.6151
R1153 B.n357 B.n356 10.6151
R1154 B.n356 B.n355 10.6151
R1155 B.n355 B.n164 10.6151
R1156 B.n349 B.n164 10.6151
R1157 B.n349 B.n348 10.6151
R1158 B.n348 B.n347 10.6151
R1159 B.n347 B.n166 10.6151
R1160 B.n341 B.n166 10.6151
R1161 B.n341 B.n340 10.6151
R1162 B.n340 B.n339 10.6151
R1163 B.n335 B.n334 10.6151
R1164 B.n334 B.n172 10.6151
R1165 B.n329 B.n172 10.6151
R1166 B.n329 B.n328 10.6151
R1167 B.n328 B.n327 10.6151
R1168 B.n327 B.n174 10.6151
R1169 B.n321 B.n174 10.6151
R1170 B.n321 B.n320 10.6151
R1171 B.n318 B.n178 10.6151
R1172 B.n312 B.n178 10.6151
R1173 B.n312 B.n311 10.6151
R1174 B.n311 B.n310 10.6151
R1175 B.n310 B.n180 10.6151
R1176 B.n304 B.n180 10.6151
R1177 B.n304 B.n303 10.6151
R1178 B.n303 B.n302 10.6151
R1179 B.n302 B.n182 10.6151
R1180 B.n296 B.n182 10.6151
R1181 B.n296 B.n295 10.6151
R1182 B.n295 B.n294 10.6151
R1183 B.n294 B.n184 10.6151
R1184 B.n288 B.n184 10.6151
R1185 B.n288 B.n287 10.6151
R1186 B.n287 B.n286 10.6151
R1187 B.n286 B.n186 10.6151
R1188 B.n280 B.n186 10.6151
R1189 B.n280 B.n279 10.6151
R1190 B.n279 B.n278 10.6151
R1191 B.n278 B.n188 10.6151
R1192 B.n272 B.n188 10.6151
R1193 B.n272 B.n271 10.6151
R1194 B.n271 B.n270 10.6151
R1195 B.n270 B.n190 10.6151
R1196 B.n264 B.n190 10.6151
R1197 B.n264 B.n263 10.6151
R1198 B.n263 B.n262 10.6151
R1199 B.n262 B.n192 10.6151
R1200 B.n256 B.n192 10.6151
R1201 B.n256 B.n255 10.6151
R1202 B.n255 B.n254 10.6151
R1203 B.n254 B.n194 10.6151
R1204 B.n248 B.n194 10.6151
R1205 B.n248 B.n247 10.6151
R1206 B.n247 B.n246 10.6151
R1207 B.n246 B.n196 10.6151
R1208 B.n240 B.n196 10.6151
R1209 B.n240 B.n239 10.6151
R1210 B.n239 B.n238 10.6151
R1211 B.n238 B.n198 10.6151
R1212 B.n232 B.n198 10.6151
R1213 B.n232 B.n231 10.6151
R1214 B.n231 B.n230 10.6151
R1215 B.n230 B.n200 10.6151
R1216 B.n224 B.n200 10.6151
R1217 B.n224 B.n223 10.6151
R1218 B.n223 B.n222 10.6151
R1219 B.n222 B.n202 10.6151
R1220 B.n216 B.n202 10.6151
R1221 B.n216 B.n215 10.6151
R1222 B.n215 B.n214 10.6151
R1223 B.n214 B.n204 10.6151
R1224 B.n208 B.n204 10.6151
R1225 B.n208 B.n207 10.6151
R1226 B.n207 B.n136 10.6151
R1227 B.n455 B.n454 10.6151
R1228 B.n456 B.n455 10.6151
R1229 B.n456 B.n128 10.6151
R1230 B.n466 B.n128 10.6151
R1231 B.n467 B.n466 10.6151
R1232 B.n468 B.n467 10.6151
R1233 B.n468 B.n120 10.6151
R1234 B.n478 B.n120 10.6151
R1235 B.n479 B.n478 10.6151
R1236 B.n480 B.n479 10.6151
R1237 B.n480 B.n111 10.6151
R1238 B.n490 B.n111 10.6151
R1239 B.n491 B.n490 10.6151
R1240 B.n493 B.n491 10.6151
R1241 B.n493 B.n492 10.6151
R1242 B.n492 B.n105 10.6151
R1243 B.n505 B.n105 10.6151
R1244 B.n506 B.n505 10.6151
R1245 B.n507 B.n506 10.6151
R1246 B.n508 B.n507 10.6151
R1247 B.n509 B.n508 10.6151
R1248 B.n512 B.n509 10.6151
R1249 B.n513 B.n512 10.6151
R1250 B.n514 B.n513 10.6151
R1251 B.n515 B.n514 10.6151
R1252 B.n517 B.n515 10.6151
R1253 B.n518 B.n517 10.6151
R1254 B.n519 B.n518 10.6151
R1255 B.n520 B.n519 10.6151
R1256 B.n522 B.n520 10.6151
R1257 B.n523 B.n522 10.6151
R1258 B.n524 B.n523 10.6151
R1259 B.n525 B.n524 10.6151
R1260 B.n527 B.n525 10.6151
R1261 B.n528 B.n527 10.6151
R1262 B.n529 B.n528 10.6151
R1263 B.n530 B.n529 10.6151
R1264 B.n809 B.n1 10.6151
R1265 B.n809 B.n808 10.6151
R1266 B.n808 B.n807 10.6151
R1267 B.n807 B.n10 10.6151
R1268 B.n801 B.n10 10.6151
R1269 B.n801 B.n800 10.6151
R1270 B.n800 B.n799 10.6151
R1271 B.n799 B.n18 10.6151
R1272 B.n793 B.n18 10.6151
R1273 B.n793 B.n792 10.6151
R1274 B.n792 B.n791 10.6151
R1275 B.n791 B.n25 10.6151
R1276 B.n785 B.n25 10.6151
R1277 B.n785 B.n784 10.6151
R1278 B.n784 B.n783 10.6151
R1279 B.n783 B.n32 10.6151
R1280 B.n777 B.n32 10.6151
R1281 B.n776 B.n775 10.6151
R1282 B.n775 B.n39 10.6151
R1283 B.n769 B.n39 10.6151
R1284 B.n769 B.n768 10.6151
R1285 B.n768 B.n767 10.6151
R1286 B.n767 B.n41 10.6151
R1287 B.n761 B.n41 10.6151
R1288 B.n761 B.n760 10.6151
R1289 B.n760 B.n759 10.6151
R1290 B.n759 B.n43 10.6151
R1291 B.n753 B.n43 10.6151
R1292 B.n753 B.n752 10.6151
R1293 B.n752 B.n751 10.6151
R1294 B.n751 B.n45 10.6151
R1295 B.n745 B.n45 10.6151
R1296 B.n745 B.n744 10.6151
R1297 B.n744 B.n743 10.6151
R1298 B.n743 B.n47 10.6151
R1299 B.n737 B.n47 10.6151
R1300 B.n737 B.n736 10.6151
R1301 B.n736 B.n735 10.6151
R1302 B.n735 B.n49 10.6151
R1303 B.n729 B.n49 10.6151
R1304 B.n729 B.n728 10.6151
R1305 B.n728 B.n727 10.6151
R1306 B.n727 B.n51 10.6151
R1307 B.n721 B.n51 10.6151
R1308 B.n721 B.n720 10.6151
R1309 B.n720 B.n719 10.6151
R1310 B.n719 B.n53 10.6151
R1311 B.n713 B.n53 10.6151
R1312 B.n713 B.n712 10.6151
R1313 B.n712 B.n711 10.6151
R1314 B.n711 B.n55 10.6151
R1315 B.n705 B.n55 10.6151
R1316 B.n705 B.n704 10.6151
R1317 B.n704 B.n703 10.6151
R1318 B.n703 B.n57 10.6151
R1319 B.n697 B.n57 10.6151
R1320 B.n697 B.n696 10.6151
R1321 B.n696 B.n695 10.6151
R1322 B.n695 B.n59 10.6151
R1323 B.n689 B.n59 10.6151
R1324 B.n689 B.n688 10.6151
R1325 B.n688 B.n687 10.6151
R1326 B.n687 B.n61 10.6151
R1327 B.n681 B.n61 10.6151
R1328 B.n681 B.n680 10.6151
R1329 B.n680 B.n679 10.6151
R1330 B.n679 B.n63 10.6151
R1331 B.n673 B.n63 10.6151
R1332 B.n673 B.n672 10.6151
R1333 B.n672 B.n671 10.6151
R1334 B.n671 B.n65 10.6151
R1335 B.n665 B.n65 10.6151
R1336 B.n665 B.n664 10.6151
R1337 B.n662 B.n69 10.6151
R1338 B.n656 B.n69 10.6151
R1339 B.n656 B.n655 10.6151
R1340 B.n655 B.n654 10.6151
R1341 B.n654 B.n71 10.6151
R1342 B.n648 B.n71 10.6151
R1343 B.n648 B.n647 10.6151
R1344 B.n647 B.n646 10.6151
R1345 B.n642 B.n641 10.6151
R1346 B.n641 B.n77 10.6151
R1347 B.n636 B.n77 10.6151
R1348 B.n636 B.n635 10.6151
R1349 B.n635 B.n634 10.6151
R1350 B.n634 B.n79 10.6151
R1351 B.n628 B.n79 10.6151
R1352 B.n628 B.n627 10.6151
R1353 B.n627 B.n626 10.6151
R1354 B.n626 B.n81 10.6151
R1355 B.n620 B.n81 10.6151
R1356 B.n620 B.n619 10.6151
R1357 B.n619 B.n618 10.6151
R1358 B.n618 B.n83 10.6151
R1359 B.n612 B.n83 10.6151
R1360 B.n612 B.n611 10.6151
R1361 B.n611 B.n610 10.6151
R1362 B.n610 B.n85 10.6151
R1363 B.n604 B.n85 10.6151
R1364 B.n604 B.n603 10.6151
R1365 B.n603 B.n602 10.6151
R1366 B.n602 B.n87 10.6151
R1367 B.n596 B.n87 10.6151
R1368 B.n596 B.n595 10.6151
R1369 B.n595 B.n594 10.6151
R1370 B.n594 B.n89 10.6151
R1371 B.n588 B.n89 10.6151
R1372 B.n588 B.n587 10.6151
R1373 B.n587 B.n586 10.6151
R1374 B.n586 B.n91 10.6151
R1375 B.n580 B.n91 10.6151
R1376 B.n580 B.n579 10.6151
R1377 B.n579 B.n578 10.6151
R1378 B.n578 B.n93 10.6151
R1379 B.n572 B.n93 10.6151
R1380 B.n572 B.n571 10.6151
R1381 B.n571 B.n570 10.6151
R1382 B.n570 B.n95 10.6151
R1383 B.n564 B.n95 10.6151
R1384 B.n564 B.n563 10.6151
R1385 B.n563 B.n562 10.6151
R1386 B.n562 B.n97 10.6151
R1387 B.n556 B.n97 10.6151
R1388 B.n556 B.n555 10.6151
R1389 B.n555 B.n554 10.6151
R1390 B.n554 B.n99 10.6151
R1391 B.n548 B.n99 10.6151
R1392 B.n548 B.n547 10.6151
R1393 B.n547 B.n546 10.6151
R1394 B.n546 B.n101 10.6151
R1395 B.n540 B.n101 10.6151
R1396 B.n540 B.n539 10.6151
R1397 B.n539 B.n538 10.6151
R1398 B.n538 B.n103 10.6151
R1399 B.n532 B.n103 10.6151
R1400 B.n532 B.n531 10.6151
R1401 B.n817 B.n0 8.11757
R1402 B.n817 B.n1 8.11757
R1403 B.n335 B.n170 6.5566
R1404 B.n320 B.n319 6.5566
R1405 B.n663 B.n662 6.5566
R1406 B.n646 B.n75 6.5566
R1407 B.n339 B.n170 4.05904
R1408 B.n319 B.n318 4.05904
R1409 B.n664 B.n663 4.05904
R1410 B.n642 B.n75 4.05904
R1411 B.n114 B.t1 0.490369
R1412 B.t5 B.n804 0.490369
R1413 VN.n0 VN.t5 851.042
R1414 VN.n4 VN.t1 851.042
R1415 VN.n1 VN.t2 824.221
R1416 VN.n2 VN.t0 824.221
R1417 VN.n5 VN.t4 824.221
R1418 VN.n6 VN.t3 824.221
R1419 VN.n3 VN.n2 161.3
R1420 VN.n7 VN.n6 161.3
R1421 VN.n2 VN.n1 48.2005
R1422 VN.n6 VN.n5 48.2005
R1423 VN.n7 VN.n4 45.1367
R1424 VN.n3 VN.n0 45.1367
R1425 VN VN.n7 44.9569
R1426 VN.n5 VN.n4 13.3799
R1427 VN.n1 VN.n0 13.3799
R1428 VN VN.n3 0.0516364
R1429 VDD2.n1 VDD2.t0 62.7559
R1430 VDD2.n2 VDD2.t2 62.2424
R1431 VDD2.n1 VDD2.n0 61.224
R1432 VDD2 VDD2.n3 61.2212
R1433 VDD2.n2 VDD2.n1 40.9912
R1434 VDD2.n3 VDD2.t1 1.153
R1435 VDD2.n3 VDD2.t4 1.153
R1436 VDD2.n0 VDD2.t3 1.153
R1437 VDD2.n0 VDD2.t5 1.153
R1438 VDD2 VDD2.n2 0.627655
C0 VDD1 VTAIL 14.8446f
C1 VN VP 5.89198f
C2 VDD2 VP 0.286212f
C3 VDD2 VN 5.34276f
C4 VTAIL VP 4.78861f
C5 VTAIL VN 4.77372f
C6 VDD2 VTAIL 14.8739f
C7 VDD1 VP 5.47399f
C8 VDD1 VN 0.148325f
C9 VDD1 VDD2 0.659222f
C10 VDD2 B 5.309386f
C11 VDD1 B 5.540463f
C12 VTAIL B 8.123399f
C13 VN B 8.0432f
C14 VP B 5.660073f
C15 VDD2.t0 B 3.84151f
C16 VDD2.t3 B 0.330356f
C17 VDD2.t5 B 0.330356f
C18 VDD2.n0 B 3.00476f
C19 VDD2.n1 B 2.27934f
C20 VDD2.t2 B 3.83892f
C21 VDD2.n2 B 2.56967f
C22 VDD2.t1 B 0.330356f
C23 VDD2.t4 B 0.330356f
C24 VDD2.n3 B 3.00473f
C25 VN.t5 B 1.34688f
C26 VN.n0 B 0.492966f
C27 VN.t2 B 1.33087f
C28 VN.n1 B 0.519219f
C29 VN.t0 B 1.33087f
C30 VN.n2 B 0.507952f
C31 VN.n3 B 0.195896f
C32 VN.t1 B 1.34688f
C33 VN.n4 B 0.492966f
C34 VN.t4 B 1.33087f
C35 VN.n5 B 0.519219f
C36 VN.t3 B 1.33087f
C37 VN.n6 B 0.507952f
C38 VN.n7 B 2.44874f
C39 VDD1.t0 B 3.84409f
C40 VDD1.t1 B 3.84343f
C41 VDD1.t2 B 0.33052f
C42 VDD1.t5 B 0.33052f
C43 VDD1.n0 B 3.00626f
C44 VDD1.n1 B 2.35335f
C45 VDD1.t4 B 0.33052f
C46 VDD1.t3 B 0.33052f
C47 VDD1.n2 B 3.00562f
C48 VDD1.n3 B 2.54242f
C49 VTAIL.t0 B 0.335557f
C50 VTAIL.t11 B 0.335557f
C51 VTAIL.n0 B 2.97646f
C52 VTAIL.n1 B 0.333081f
C53 VTAIL.t9 B 3.80166f
C54 VTAIL.n2 B 0.46372f
C55 VTAIL.t8 B 0.335557f
C56 VTAIL.t6 B 0.335557f
C57 VTAIL.n3 B 2.97646f
C58 VTAIL.n4 B 1.94225f
C59 VTAIL.t2 B 0.335557f
C60 VTAIL.t1 B 0.335557f
C61 VTAIL.n5 B 2.97647f
C62 VTAIL.n6 B 1.94225f
C63 VTAIL.t4 B 3.80168f
C64 VTAIL.n7 B 0.463697f
C65 VTAIL.t7 B 0.335557f
C66 VTAIL.t5 B 0.335557f
C67 VTAIL.n8 B 2.97647f
C68 VTAIL.n9 B 0.373757f
C69 VTAIL.t10 B 3.80166f
C70 VTAIL.n10 B 1.97179f
C71 VTAIL.t3 B 3.80166f
C72 VTAIL.n11 B 1.95205f
C73 VP.n0 B 0.067218f
C74 VP.t5 B 1.3697f
C75 VP.n1 B 0.501315f
C76 VP.t2 B 1.35341f
C77 VP.t1 B 1.35341f
C78 VP.n2 B 0.528013f
C79 VP.n3 B 0.516555f
C80 VP.n4 B 2.45718f
C81 VP.n5 B 2.35481f
C82 VP.t4 B 1.35341f
C83 VP.n6 B 0.516555f
C84 VP.t3 B 1.35341f
C85 VP.n7 B 0.528013f
C86 VP.t0 B 1.35341f
C87 VP.n8 B 0.516555f
C88 VP.n9 B 0.056013f
.ends

