* NGSPICE file created from diff_pair_sample_0533.ext - technology: sky130A

.subckt diff_pair_sample_0533 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1306_n1636# sky130_fd_pr__pfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=0.51
X1 VDD1.t1 VP.t0 VTAIL.t2 w_n1306_n1636# sky130_fd_pr__pfet_01v8 ad=1.2948 pd=7.42 as=1.2948 ps=7.42 w=3.32 l=0.51
X2 B.t8 B.t6 B.t7 w_n1306_n1636# sky130_fd_pr__pfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=0.51
X3 B.t5 B.t3 B.t4 w_n1306_n1636# sky130_fd_pr__pfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=0.51
X4 B.t2 B.t0 B.t1 w_n1306_n1636# sky130_fd_pr__pfet_01v8 ad=1.2948 pd=7.42 as=0 ps=0 w=3.32 l=0.51
X5 VDD2.t1 VN.t0 VTAIL.t0 w_n1306_n1636# sky130_fd_pr__pfet_01v8 ad=1.2948 pd=7.42 as=1.2948 ps=7.42 w=3.32 l=0.51
X6 VDD1.t0 VP.t1 VTAIL.t3 w_n1306_n1636# sky130_fd_pr__pfet_01v8 ad=1.2948 pd=7.42 as=1.2948 ps=7.42 w=3.32 l=0.51
X7 VDD2.t0 VN.t1 VTAIL.t1 w_n1306_n1636# sky130_fd_pr__pfet_01v8 ad=1.2948 pd=7.42 as=1.2948 ps=7.42 w=3.32 l=0.51
R0 B.n203 B.n34 585
R1 B.n205 B.n204 585
R2 B.n206 B.n33 585
R3 B.n208 B.n207 585
R4 B.n209 B.n32 585
R5 B.n211 B.n210 585
R6 B.n212 B.n31 585
R7 B.n214 B.n213 585
R8 B.n215 B.n30 585
R9 B.n217 B.n216 585
R10 B.n218 B.n29 585
R11 B.n220 B.n219 585
R12 B.n221 B.n28 585
R13 B.n223 B.n222 585
R14 B.n224 B.n27 585
R15 B.n226 B.n225 585
R16 B.n228 B.n24 585
R17 B.n230 B.n229 585
R18 B.n231 B.n23 585
R19 B.n233 B.n232 585
R20 B.n234 B.n22 585
R21 B.n236 B.n235 585
R22 B.n237 B.n21 585
R23 B.n239 B.n238 585
R24 B.n240 B.n17 585
R25 B.n242 B.n241 585
R26 B.n243 B.n16 585
R27 B.n245 B.n244 585
R28 B.n246 B.n15 585
R29 B.n248 B.n247 585
R30 B.n249 B.n14 585
R31 B.n251 B.n250 585
R32 B.n252 B.n13 585
R33 B.n254 B.n253 585
R34 B.n255 B.n12 585
R35 B.n257 B.n256 585
R36 B.n258 B.n11 585
R37 B.n260 B.n259 585
R38 B.n261 B.n10 585
R39 B.n263 B.n262 585
R40 B.n264 B.n9 585
R41 B.n266 B.n265 585
R42 B.n202 B.n201 585
R43 B.n200 B.n35 585
R44 B.n199 B.n198 585
R45 B.n197 B.n36 585
R46 B.n196 B.n195 585
R47 B.n194 B.n37 585
R48 B.n193 B.n192 585
R49 B.n191 B.n38 585
R50 B.n190 B.n189 585
R51 B.n188 B.n39 585
R52 B.n187 B.n186 585
R53 B.n185 B.n40 585
R54 B.n184 B.n183 585
R55 B.n182 B.n41 585
R56 B.n181 B.n180 585
R57 B.n179 B.n42 585
R58 B.n178 B.n177 585
R59 B.n176 B.n43 585
R60 B.n175 B.n174 585
R61 B.n173 B.n44 585
R62 B.n172 B.n171 585
R63 B.n170 B.n45 585
R64 B.n169 B.n168 585
R65 B.n167 B.n46 585
R66 B.n166 B.n165 585
R67 B.n164 B.n47 585
R68 B.n163 B.n162 585
R69 B.n98 B.n73 585
R70 B.n100 B.n99 585
R71 B.n101 B.n72 585
R72 B.n103 B.n102 585
R73 B.n104 B.n71 585
R74 B.n106 B.n105 585
R75 B.n107 B.n70 585
R76 B.n109 B.n108 585
R77 B.n110 B.n69 585
R78 B.n112 B.n111 585
R79 B.n113 B.n68 585
R80 B.n115 B.n114 585
R81 B.n116 B.n67 585
R82 B.n118 B.n117 585
R83 B.n119 B.n66 585
R84 B.n121 B.n120 585
R85 B.n123 B.n122 585
R86 B.n124 B.n62 585
R87 B.n126 B.n125 585
R88 B.n127 B.n61 585
R89 B.n129 B.n128 585
R90 B.n130 B.n60 585
R91 B.n132 B.n131 585
R92 B.n133 B.n59 585
R93 B.n135 B.n134 585
R94 B.n136 B.n56 585
R95 B.n139 B.n138 585
R96 B.n140 B.n55 585
R97 B.n142 B.n141 585
R98 B.n143 B.n54 585
R99 B.n145 B.n144 585
R100 B.n146 B.n53 585
R101 B.n148 B.n147 585
R102 B.n149 B.n52 585
R103 B.n151 B.n150 585
R104 B.n152 B.n51 585
R105 B.n154 B.n153 585
R106 B.n155 B.n50 585
R107 B.n157 B.n156 585
R108 B.n158 B.n49 585
R109 B.n160 B.n159 585
R110 B.n161 B.n48 585
R111 B.n97 B.n96 585
R112 B.n95 B.n74 585
R113 B.n94 B.n93 585
R114 B.n92 B.n75 585
R115 B.n91 B.n90 585
R116 B.n89 B.n76 585
R117 B.n88 B.n87 585
R118 B.n86 B.n77 585
R119 B.n85 B.n84 585
R120 B.n83 B.n78 585
R121 B.n82 B.n81 585
R122 B.n80 B.n79 585
R123 B.n2 B.n0 585
R124 B.n285 B.n1 585
R125 B.n284 B.n283 585
R126 B.n282 B.n3 585
R127 B.n281 B.n280 585
R128 B.n279 B.n4 585
R129 B.n278 B.n277 585
R130 B.n276 B.n5 585
R131 B.n275 B.n274 585
R132 B.n273 B.n6 585
R133 B.n272 B.n271 585
R134 B.n270 B.n7 585
R135 B.n269 B.n268 585
R136 B.n267 B.n8 585
R137 B.n287 B.n286 585
R138 B.n98 B.n97 497.305
R139 B.n267 B.n266 497.305
R140 B.n163 B.n48 497.305
R141 B.n201 B.n34 497.305
R142 B.n57 B.t0 363.058
R143 B.n63 B.t3 363.058
R144 B.n18 B.t6 363.058
R145 B.n25 B.t9 363.058
R146 B.n57 B.t2 244.179
R147 B.n25 B.t10 244.179
R148 B.n63 B.t5 244.179
R149 B.n18 B.t7 244.179
R150 B.n58 B.t1 227.888
R151 B.n26 B.t11 227.888
R152 B.n64 B.t4 227.887
R153 B.n19 B.t8 227.887
R154 B.n97 B.n74 163.367
R155 B.n93 B.n74 163.367
R156 B.n93 B.n92 163.367
R157 B.n92 B.n91 163.367
R158 B.n91 B.n76 163.367
R159 B.n87 B.n76 163.367
R160 B.n87 B.n86 163.367
R161 B.n86 B.n85 163.367
R162 B.n85 B.n78 163.367
R163 B.n81 B.n78 163.367
R164 B.n81 B.n80 163.367
R165 B.n80 B.n2 163.367
R166 B.n286 B.n2 163.367
R167 B.n286 B.n285 163.367
R168 B.n285 B.n284 163.367
R169 B.n284 B.n3 163.367
R170 B.n280 B.n3 163.367
R171 B.n280 B.n279 163.367
R172 B.n279 B.n278 163.367
R173 B.n278 B.n5 163.367
R174 B.n274 B.n5 163.367
R175 B.n274 B.n273 163.367
R176 B.n273 B.n272 163.367
R177 B.n272 B.n7 163.367
R178 B.n268 B.n7 163.367
R179 B.n268 B.n267 163.367
R180 B.n99 B.n98 163.367
R181 B.n99 B.n72 163.367
R182 B.n103 B.n72 163.367
R183 B.n104 B.n103 163.367
R184 B.n105 B.n104 163.367
R185 B.n105 B.n70 163.367
R186 B.n109 B.n70 163.367
R187 B.n110 B.n109 163.367
R188 B.n111 B.n110 163.367
R189 B.n111 B.n68 163.367
R190 B.n115 B.n68 163.367
R191 B.n116 B.n115 163.367
R192 B.n117 B.n116 163.367
R193 B.n117 B.n66 163.367
R194 B.n121 B.n66 163.367
R195 B.n122 B.n121 163.367
R196 B.n122 B.n62 163.367
R197 B.n126 B.n62 163.367
R198 B.n127 B.n126 163.367
R199 B.n128 B.n127 163.367
R200 B.n128 B.n60 163.367
R201 B.n132 B.n60 163.367
R202 B.n133 B.n132 163.367
R203 B.n134 B.n133 163.367
R204 B.n134 B.n56 163.367
R205 B.n139 B.n56 163.367
R206 B.n140 B.n139 163.367
R207 B.n141 B.n140 163.367
R208 B.n141 B.n54 163.367
R209 B.n145 B.n54 163.367
R210 B.n146 B.n145 163.367
R211 B.n147 B.n146 163.367
R212 B.n147 B.n52 163.367
R213 B.n151 B.n52 163.367
R214 B.n152 B.n151 163.367
R215 B.n153 B.n152 163.367
R216 B.n153 B.n50 163.367
R217 B.n157 B.n50 163.367
R218 B.n158 B.n157 163.367
R219 B.n159 B.n158 163.367
R220 B.n159 B.n48 163.367
R221 B.n164 B.n163 163.367
R222 B.n165 B.n164 163.367
R223 B.n165 B.n46 163.367
R224 B.n169 B.n46 163.367
R225 B.n170 B.n169 163.367
R226 B.n171 B.n170 163.367
R227 B.n171 B.n44 163.367
R228 B.n175 B.n44 163.367
R229 B.n176 B.n175 163.367
R230 B.n177 B.n176 163.367
R231 B.n177 B.n42 163.367
R232 B.n181 B.n42 163.367
R233 B.n182 B.n181 163.367
R234 B.n183 B.n182 163.367
R235 B.n183 B.n40 163.367
R236 B.n187 B.n40 163.367
R237 B.n188 B.n187 163.367
R238 B.n189 B.n188 163.367
R239 B.n189 B.n38 163.367
R240 B.n193 B.n38 163.367
R241 B.n194 B.n193 163.367
R242 B.n195 B.n194 163.367
R243 B.n195 B.n36 163.367
R244 B.n199 B.n36 163.367
R245 B.n200 B.n199 163.367
R246 B.n201 B.n200 163.367
R247 B.n266 B.n9 163.367
R248 B.n262 B.n9 163.367
R249 B.n262 B.n261 163.367
R250 B.n261 B.n260 163.367
R251 B.n260 B.n11 163.367
R252 B.n256 B.n11 163.367
R253 B.n256 B.n255 163.367
R254 B.n255 B.n254 163.367
R255 B.n254 B.n13 163.367
R256 B.n250 B.n13 163.367
R257 B.n250 B.n249 163.367
R258 B.n249 B.n248 163.367
R259 B.n248 B.n15 163.367
R260 B.n244 B.n15 163.367
R261 B.n244 B.n243 163.367
R262 B.n243 B.n242 163.367
R263 B.n242 B.n17 163.367
R264 B.n238 B.n17 163.367
R265 B.n238 B.n237 163.367
R266 B.n237 B.n236 163.367
R267 B.n236 B.n22 163.367
R268 B.n232 B.n22 163.367
R269 B.n232 B.n231 163.367
R270 B.n231 B.n230 163.367
R271 B.n230 B.n24 163.367
R272 B.n225 B.n24 163.367
R273 B.n225 B.n224 163.367
R274 B.n224 B.n223 163.367
R275 B.n223 B.n28 163.367
R276 B.n219 B.n28 163.367
R277 B.n219 B.n218 163.367
R278 B.n218 B.n217 163.367
R279 B.n217 B.n30 163.367
R280 B.n213 B.n30 163.367
R281 B.n213 B.n212 163.367
R282 B.n212 B.n211 163.367
R283 B.n211 B.n32 163.367
R284 B.n207 B.n32 163.367
R285 B.n207 B.n206 163.367
R286 B.n206 B.n205 163.367
R287 B.n205 B.n34 163.367
R288 B.n137 B.n58 59.5399
R289 B.n65 B.n64 59.5399
R290 B.n20 B.n19 59.5399
R291 B.n227 B.n26 59.5399
R292 B.n265 B.n8 32.3127
R293 B.n203 B.n202 32.3127
R294 B.n162 B.n161 32.3127
R295 B.n96 B.n73 32.3127
R296 B B.n287 18.0485
R297 B.n58 B.n57 16.2914
R298 B.n64 B.n63 16.2914
R299 B.n19 B.n18 16.2914
R300 B.n26 B.n25 16.2914
R301 B.n265 B.n264 10.6151
R302 B.n264 B.n263 10.6151
R303 B.n263 B.n10 10.6151
R304 B.n259 B.n10 10.6151
R305 B.n259 B.n258 10.6151
R306 B.n258 B.n257 10.6151
R307 B.n257 B.n12 10.6151
R308 B.n253 B.n12 10.6151
R309 B.n253 B.n252 10.6151
R310 B.n252 B.n251 10.6151
R311 B.n251 B.n14 10.6151
R312 B.n247 B.n14 10.6151
R313 B.n247 B.n246 10.6151
R314 B.n246 B.n245 10.6151
R315 B.n245 B.n16 10.6151
R316 B.n241 B.n240 10.6151
R317 B.n240 B.n239 10.6151
R318 B.n239 B.n21 10.6151
R319 B.n235 B.n21 10.6151
R320 B.n235 B.n234 10.6151
R321 B.n234 B.n233 10.6151
R322 B.n233 B.n23 10.6151
R323 B.n229 B.n23 10.6151
R324 B.n229 B.n228 10.6151
R325 B.n226 B.n27 10.6151
R326 B.n222 B.n27 10.6151
R327 B.n222 B.n221 10.6151
R328 B.n221 B.n220 10.6151
R329 B.n220 B.n29 10.6151
R330 B.n216 B.n29 10.6151
R331 B.n216 B.n215 10.6151
R332 B.n215 B.n214 10.6151
R333 B.n214 B.n31 10.6151
R334 B.n210 B.n31 10.6151
R335 B.n210 B.n209 10.6151
R336 B.n209 B.n208 10.6151
R337 B.n208 B.n33 10.6151
R338 B.n204 B.n33 10.6151
R339 B.n204 B.n203 10.6151
R340 B.n162 B.n47 10.6151
R341 B.n166 B.n47 10.6151
R342 B.n167 B.n166 10.6151
R343 B.n168 B.n167 10.6151
R344 B.n168 B.n45 10.6151
R345 B.n172 B.n45 10.6151
R346 B.n173 B.n172 10.6151
R347 B.n174 B.n173 10.6151
R348 B.n174 B.n43 10.6151
R349 B.n178 B.n43 10.6151
R350 B.n179 B.n178 10.6151
R351 B.n180 B.n179 10.6151
R352 B.n180 B.n41 10.6151
R353 B.n184 B.n41 10.6151
R354 B.n185 B.n184 10.6151
R355 B.n186 B.n185 10.6151
R356 B.n186 B.n39 10.6151
R357 B.n190 B.n39 10.6151
R358 B.n191 B.n190 10.6151
R359 B.n192 B.n191 10.6151
R360 B.n192 B.n37 10.6151
R361 B.n196 B.n37 10.6151
R362 B.n197 B.n196 10.6151
R363 B.n198 B.n197 10.6151
R364 B.n198 B.n35 10.6151
R365 B.n202 B.n35 10.6151
R366 B.n100 B.n73 10.6151
R367 B.n101 B.n100 10.6151
R368 B.n102 B.n101 10.6151
R369 B.n102 B.n71 10.6151
R370 B.n106 B.n71 10.6151
R371 B.n107 B.n106 10.6151
R372 B.n108 B.n107 10.6151
R373 B.n108 B.n69 10.6151
R374 B.n112 B.n69 10.6151
R375 B.n113 B.n112 10.6151
R376 B.n114 B.n113 10.6151
R377 B.n114 B.n67 10.6151
R378 B.n118 B.n67 10.6151
R379 B.n119 B.n118 10.6151
R380 B.n120 B.n119 10.6151
R381 B.n124 B.n123 10.6151
R382 B.n125 B.n124 10.6151
R383 B.n125 B.n61 10.6151
R384 B.n129 B.n61 10.6151
R385 B.n130 B.n129 10.6151
R386 B.n131 B.n130 10.6151
R387 B.n131 B.n59 10.6151
R388 B.n135 B.n59 10.6151
R389 B.n136 B.n135 10.6151
R390 B.n138 B.n55 10.6151
R391 B.n142 B.n55 10.6151
R392 B.n143 B.n142 10.6151
R393 B.n144 B.n143 10.6151
R394 B.n144 B.n53 10.6151
R395 B.n148 B.n53 10.6151
R396 B.n149 B.n148 10.6151
R397 B.n150 B.n149 10.6151
R398 B.n150 B.n51 10.6151
R399 B.n154 B.n51 10.6151
R400 B.n155 B.n154 10.6151
R401 B.n156 B.n155 10.6151
R402 B.n156 B.n49 10.6151
R403 B.n160 B.n49 10.6151
R404 B.n161 B.n160 10.6151
R405 B.n96 B.n95 10.6151
R406 B.n95 B.n94 10.6151
R407 B.n94 B.n75 10.6151
R408 B.n90 B.n75 10.6151
R409 B.n90 B.n89 10.6151
R410 B.n89 B.n88 10.6151
R411 B.n88 B.n77 10.6151
R412 B.n84 B.n77 10.6151
R413 B.n84 B.n83 10.6151
R414 B.n83 B.n82 10.6151
R415 B.n82 B.n79 10.6151
R416 B.n79 B.n0 10.6151
R417 B.n283 B.n1 10.6151
R418 B.n283 B.n282 10.6151
R419 B.n282 B.n281 10.6151
R420 B.n281 B.n4 10.6151
R421 B.n277 B.n4 10.6151
R422 B.n277 B.n276 10.6151
R423 B.n276 B.n275 10.6151
R424 B.n275 B.n6 10.6151
R425 B.n271 B.n6 10.6151
R426 B.n271 B.n270 10.6151
R427 B.n270 B.n269 10.6151
R428 B.n269 B.n8 10.6151
R429 B.n20 B.n16 8.74196
R430 B.n227 B.n226 8.74196
R431 B.n120 B.n65 8.74196
R432 B.n138 B.n137 8.74196
R433 B.n287 B.n0 2.81026
R434 B.n287 B.n1 2.81026
R435 B.n241 B.n20 1.87367
R436 B.n228 B.n227 1.87367
R437 B.n123 B.n65 1.87367
R438 B.n137 B.n136 1.87367
R439 VP.n0 VP.t1 427.765
R440 VP.n0 VP.t0 395.212
R441 VP VP.n0 0.0516364
R442 VTAIL.n58 VTAIL.n48 756.745
R443 VTAIL.n10 VTAIL.n0 756.745
R444 VTAIL.n42 VTAIL.n32 756.745
R445 VTAIL.n26 VTAIL.n16 756.745
R446 VTAIL.n52 VTAIL.n51 585
R447 VTAIL.n57 VTAIL.n56 585
R448 VTAIL.n59 VTAIL.n58 585
R449 VTAIL.n4 VTAIL.n3 585
R450 VTAIL.n9 VTAIL.n8 585
R451 VTAIL.n11 VTAIL.n10 585
R452 VTAIL.n43 VTAIL.n42 585
R453 VTAIL.n41 VTAIL.n40 585
R454 VTAIL.n36 VTAIL.n35 585
R455 VTAIL.n27 VTAIL.n26 585
R456 VTAIL.n25 VTAIL.n24 585
R457 VTAIL.n20 VTAIL.n19 585
R458 VTAIL.n53 VTAIL.t0 336.901
R459 VTAIL.n5 VTAIL.t2 336.901
R460 VTAIL.n37 VTAIL.t3 336.901
R461 VTAIL.n21 VTAIL.t1 336.901
R462 VTAIL.n57 VTAIL.n51 171.744
R463 VTAIL.n58 VTAIL.n57 171.744
R464 VTAIL.n9 VTAIL.n3 171.744
R465 VTAIL.n10 VTAIL.n9 171.744
R466 VTAIL.n42 VTAIL.n41 171.744
R467 VTAIL.n41 VTAIL.n35 171.744
R468 VTAIL.n26 VTAIL.n25 171.744
R469 VTAIL.n25 VTAIL.n19 171.744
R470 VTAIL.t0 VTAIL.n51 85.8723
R471 VTAIL.t2 VTAIL.n3 85.8723
R472 VTAIL.t3 VTAIL.n35 85.8723
R473 VTAIL.t1 VTAIL.n19 85.8723
R474 VTAIL.n63 VTAIL.n62 36.0641
R475 VTAIL.n15 VTAIL.n14 36.0641
R476 VTAIL.n47 VTAIL.n46 36.0641
R477 VTAIL.n31 VTAIL.n30 36.0641
R478 VTAIL.n31 VTAIL.n15 16.6945
R479 VTAIL.n53 VTAIL.n52 16.193
R480 VTAIL.n5 VTAIL.n4 16.193
R481 VTAIL.n37 VTAIL.n36 16.193
R482 VTAIL.n21 VTAIL.n20 16.193
R483 VTAIL.n63 VTAIL.n47 15.9703
R484 VTAIL.n56 VTAIL.n55 12.8005
R485 VTAIL.n8 VTAIL.n7 12.8005
R486 VTAIL.n40 VTAIL.n39 12.8005
R487 VTAIL.n24 VTAIL.n23 12.8005
R488 VTAIL.n59 VTAIL.n50 12.0247
R489 VTAIL.n11 VTAIL.n2 12.0247
R490 VTAIL.n43 VTAIL.n34 12.0247
R491 VTAIL.n27 VTAIL.n18 12.0247
R492 VTAIL.n60 VTAIL.n48 11.249
R493 VTAIL.n12 VTAIL.n0 11.249
R494 VTAIL.n44 VTAIL.n32 11.249
R495 VTAIL.n28 VTAIL.n16 11.249
R496 VTAIL.n62 VTAIL.n61 9.45567
R497 VTAIL.n14 VTAIL.n13 9.45567
R498 VTAIL.n46 VTAIL.n45 9.45567
R499 VTAIL.n30 VTAIL.n29 9.45567
R500 VTAIL.n61 VTAIL.n60 9.3005
R501 VTAIL.n50 VTAIL.n49 9.3005
R502 VTAIL.n55 VTAIL.n54 9.3005
R503 VTAIL.n13 VTAIL.n12 9.3005
R504 VTAIL.n2 VTAIL.n1 9.3005
R505 VTAIL.n7 VTAIL.n6 9.3005
R506 VTAIL.n45 VTAIL.n44 9.3005
R507 VTAIL.n34 VTAIL.n33 9.3005
R508 VTAIL.n39 VTAIL.n38 9.3005
R509 VTAIL.n29 VTAIL.n28 9.3005
R510 VTAIL.n18 VTAIL.n17 9.3005
R511 VTAIL.n23 VTAIL.n22 9.3005
R512 VTAIL.n38 VTAIL.n37 3.91276
R513 VTAIL.n22 VTAIL.n21 3.91276
R514 VTAIL.n54 VTAIL.n53 3.91276
R515 VTAIL.n6 VTAIL.n5 3.91276
R516 VTAIL.n62 VTAIL.n48 2.71565
R517 VTAIL.n14 VTAIL.n0 2.71565
R518 VTAIL.n46 VTAIL.n32 2.71565
R519 VTAIL.n30 VTAIL.n16 2.71565
R520 VTAIL.n60 VTAIL.n59 1.93989
R521 VTAIL.n12 VTAIL.n11 1.93989
R522 VTAIL.n44 VTAIL.n43 1.93989
R523 VTAIL.n28 VTAIL.n27 1.93989
R524 VTAIL.n56 VTAIL.n50 1.16414
R525 VTAIL.n8 VTAIL.n2 1.16414
R526 VTAIL.n40 VTAIL.n34 1.16414
R527 VTAIL.n24 VTAIL.n18 1.16414
R528 VTAIL.n47 VTAIL.n31 0.832397
R529 VTAIL VTAIL.n15 0.709552
R530 VTAIL.n55 VTAIL.n52 0.388379
R531 VTAIL.n7 VTAIL.n4 0.388379
R532 VTAIL.n39 VTAIL.n36 0.388379
R533 VTAIL.n23 VTAIL.n20 0.388379
R534 VTAIL.n54 VTAIL.n49 0.155672
R535 VTAIL.n61 VTAIL.n49 0.155672
R536 VTAIL.n6 VTAIL.n1 0.155672
R537 VTAIL.n13 VTAIL.n1 0.155672
R538 VTAIL.n45 VTAIL.n33 0.155672
R539 VTAIL.n38 VTAIL.n33 0.155672
R540 VTAIL.n29 VTAIL.n17 0.155672
R541 VTAIL.n22 VTAIL.n17 0.155672
R542 VTAIL VTAIL.n63 0.123345
R543 VDD1.n10 VDD1.n0 756.745
R544 VDD1.n25 VDD1.n15 756.745
R545 VDD1.n11 VDD1.n10 585
R546 VDD1.n9 VDD1.n8 585
R547 VDD1.n4 VDD1.n3 585
R548 VDD1.n19 VDD1.n18 585
R549 VDD1.n24 VDD1.n23 585
R550 VDD1.n26 VDD1.n25 585
R551 VDD1.n5 VDD1.t0 336.901
R552 VDD1.n20 VDD1.t1 336.901
R553 VDD1.n10 VDD1.n9 171.744
R554 VDD1.n9 VDD1.n3 171.744
R555 VDD1.n24 VDD1.n18 171.744
R556 VDD1.n25 VDD1.n24 171.744
R557 VDD1.t0 VDD1.n3 85.8723
R558 VDD1.t1 VDD1.n18 85.8723
R559 VDD1 VDD1.n29 81.4358
R560 VDD1 VDD1.n14 52.9821
R561 VDD1.n5 VDD1.n4 16.193
R562 VDD1.n20 VDD1.n19 16.193
R563 VDD1.n8 VDD1.n7 12.8005
R564 VDD1.n23 VDD1.n22 12.8005
R565 VDD1.n11 VDD1.n2 12.0247
R566 VDD1.n26 VDD1.n17 12.0247
R567 VDD1.n12 VDD1.n0 11.249
R568 VDD1.n27 VDD1.n15 11.249
R569 VDD1.n14 VDD1.n13 9.45567
R570 VDD1.n29 VDD1.n28 9.45567
R571 VDD1.n13 VDD1.n12 9.3005
R572 VDD1.n2 VDD1.n1 9.3005
R573 VDD1.n7 VDD1.n6 9.3005
R574 VDD1.n28 VDD1.n27 9.3005
R575 VDD1.n17 VDD1.n16 9.3005
R576 VDD1.n22 VDD1.n21 9.3005
R577 VDD1.n6 VDD1.n5 3.91276
R578 VDD1.n21 VDD1.n20 3.91276
R579 VDD1.n14 VDD1.n0 2.71565
R580 VDD1.n29 VDD1.n15 2.71565
R581 VDD1.n12 VDD1.n11 1.93989
R582 VDD1.n27 VDD1.n26 1.93989
R583 VDD1.n8 VDD1.n2 1.16414
R584 VDD1.n23 VDD1.n17 1.16414
R585 VDD1.n7 VDD1.n4 0.388379
R586 VDD1.n22 VDD1.n19 0.388379
R587 VDD1.n13 VDD1.n1 0.155672
R588 VDD1.n6 VDD1.n1 0.155672
R589 VDD1.n21 VDD1.n16 0.155672
R590 VDD1.n28 VDD1.n16 0.155672
R591 VN VN.t1 428.147
R592 VN VN.t0 395.264
R593 VDD2.n25 VDD2.n15 756.745
R594 VDD2.n10 VDD2.n0 756.745
R595 VDD2.n26 VDD2.n25 585
R596 VDD2.n24 VDD2.n23 585
R597 VDD2.n19 VDD2.n18 585
R598 VDD2.n4 VDD2.n3 585
R599 VDD2.n9 VDD2.n8 585
R600 VDD2.n11 VDD2.n10 585
R601 VDD2.n20 VDD2.t0 336.901
R602 VDD2.n5 VDD2.t1 336.901
R603 VDD2.n25 VDD2.n24 171.744
R604 VDD2.n24 VDD2.n18 171.744
R605 VDD2.n9 VDD2.n3 171.744
R606 VDD2.n10 VDD2.n9 171.744
R607 VDD2.t0 VDD2.n18 85.8723
R608 VDD2.t1 VDD2.n3 85.8723
R609 VDD2.n30 VDD2.n14 80.73
R610 VDD2.n30 VDD2.n29 52.7429
R611 VDD2.n20 VDD2.n19 16.193
R612 VDD2.n5 VDD2.n4 16.193
R613 VDD2.n23 VDD2.n22 12.8005
R614 VDD2.n8 VDD2.n7 12.8005
R615 VDD2.n26 VDD2.n17 12.0247
R616 VDD2.n11 VDD2.n2 12.0247
R617 VDD2.n27 VDD2.n15 11.249
R618 VDD2.n12 VDD2.n0 11.249
R619 VDD2.n29 VDD2.n28 9.45567
R620 VDD2.n14 VDD2.n13 9.45567
R621 VDD2.n28 VDD2.n27 9.3005
R622 VDD2.n17 VDD2.n16 9.3005
R623 VDD2.n22 VDD2.n21 9.3005
R624 VDD2.n13 VDD2.n12 9.3005
R625 VDD2.n2 VDD2.n1 9.3005
R626 VDD2.n7 VDD2.n6 9.3005
R627 VDD2.n21 VDD2.n20 3.91276
R628 VDD2.n6 VDD2.n5 3.91276
R629 VDD2.n29 VDD2.n15 2.71565
R630 VDD2.n14 VDD2.n0 2.71565
R631 VDD2.n27 VDD2.n26 1.93989
R632 VDD2.n12 VDD2.n11 1.93989
R633 VDD2.n23 VDD2.n17 1.16414
R634 VDD2.n8 VDD2.n2 1.16414
R635 VDD2.n22 VDD2.n19 0.388379
R636 VDD2.n7 VDD2.n4 0.388379
R637 VDD2 VDD2.n30 0.239724
R638 VDD2.n28 VDD2.n16 0.155672
R639 VDD2.n21 VDD2.n16 0.155672
R640 VDD2.n6 VDD2.n1 0.155672
R641 VDD2.n13 VDD2.n1 0.155672
C0 VDD2 VTAIL 2.56199f
C1 VDD2 VP 0.251207f
C2 VDD1 VN 0.153606f
C3 w_n1306_n1636# VDD1 0.902215f
C4 VTAIL B 1.07063f
C5 VP B 0.845937f
C6 w_n1306_n1636# VN 1.45022f
C7 VTAIL VP 0.587334f
C8 VDD2 VDD1 0.441854f
C9 VDD2 VN 0.657788f
C10 w_n1306_n1636# VDD2 0.904507f
C11 VDD1 B 0.757422f
C12 VDD1 VTAIL 2.52482f
C13 VDD1 VP 0.753563f
C14 B VN 0.588573f
C15 VTAIL VN 0.573071f
C16 w_n1306_n1636# B 4.11056f
C17 VP VN 2.87246f
C18 w_n1306_n1636# VTAIL 1.45856f
C19 w_n1306_n1636# VP 1.61024f
C20 VDD2 B 0.770723f
C21 VDD2 VSUBS 0.426512f
C22 VDD1 VSUBS 1.743173f
C23 VTAIL VSUBS 0.145284f
C24 VN VSUBS 3.47403f
C25 VP VSUBS 0.660221f
C26 B VSUBS 1.552664f
C27 w_n1306_n1636# VSUBS 27.002901f
C28 VDD2.n0 VSUBS 0.019574f
C29 VDD2.n1 VSUBS 0.017609f
C30 VDD2.n2 VSUBS 0.009462f
C31 VDD2.n3 VSUBS 0.016774f
C32 VDD2.n4 VSUBS 0.013808f
C33 VDD2.t1 VSUBS 0.050796f
C34 VDD2.n5 VSUBS 0.065558f
C35 VDD2.n6 VSUBS 0.185572f
C36 VDD2.n7 VSUBS 0.009462f
C37 VDD2.n8 VSUBS 0.010019f
C38 VDD2.n9 VSUBS 0.022366f
C39 VDD2.n10 VSUBS 0.054911f
C40 VDD2.n11 VSUBS 0.010019f
C41 VDD2.n12 VSUBS 0.009462f
C42 VDD2.n13 VSUBS 0.045514f
C43 VDD2.n14 VSUBS 0.235145f
C44 VDD2.n15 VSUBS 0.019574f
C45 VDD2.n16 VSUBS 0.017609f
C46 VDD2.n17 VSUBS 0.009462f
C47 VDD2.n18 VSUBS 0.016774f
C48 VDD2.n19 VSUBS 0.013808f
C49 VDD2.t0 VSUBS 0.050796f
C50 VDD2.n20 VSUBS 0.065558f
C51 VDD2.n21 VSUBS 0.185572f
C52 VDD2.n22 VSUBS 0.009462f
C53 VDD2.n23 VSUBS 0.010019f
C54 VDD2.n24 VSUBS 0.022366f
C55 VDD2.n25 VSUBS 0.054911f
C56 VDD2.n26 VSUBS 0.010019f
C57 VDD2.n27 VSUBS 0.009462f
C58 VDD2.n28 VSUBS 0.045514f
C59 VDD2.n29 VSUBS 0.039914f
C60 VDD2.n30 VSUBS 1.20852f
C61 VN.t0 VSUBS 0.256234f
C62 VN.t1 VSUBS 0.346142f
C63 VDD1.n0 VSUBS 0.018362f
C64 VDD1.n1 VSUBS 0.016519f
C65 VDD1.n2 VSUBS 0.008876f
C66 VDD1.n3 VSUBS 0.015735f
C67 VDD1.n4 VSUBS 0.012953f
C68 VDD1.t0 VSUBS 0.047651f
C69 VDD1.n5 VSUBS 0.061498f
C70 VDD1.n6 VSUBS 0.17408f
C71 VDD1.n7 VSUBS 0.008876f
C72 VDD1.n8 VSUBS 0.009399f
C73 VDD1.n9 VSUBS 0.020981f
C74 VDD1.n10 VSUBS 0.051511f
C75 VDD1.n11 VSUBS 0.009399f
C76 VDD1.n12 VSUBS 0.008876f
C77 VDD1.n13 VSUBS 0.042695f
C78 VDD1.n14 VSUBS 0.037655f
C79 VDD1.n15 VSUBS 0.018362f
C80 VDD1.n16 VSUBS 0.016519f
C81 VDD1.n17 VSUBS 0.008876f
C82 VDD1.n18 VSUBS 0.015735f
C83 VDD1.n19 VSUBS 0.012953f
C84 VDD1.t1 VSUBS 0.047651f
C85 VDD1.n20 VSUBS 0.061498f
C86 VDD1.n21 VSUBS 0.17408f
C87 VDD1.n22 VSUBS 0.008876f
C88 VDD1.n23 VSUBS 0.009399f
C89 VDD1.n24 VSUBS 0.020981f
C90 VDD1.n25 VSUBS 0.051511f
C91 VDD1.n26 VSUBS 0.009399f
C92 VDD1.n27 VSUBS 0.008876f
C93 VDD1.n28 VSUBS 0.042695f
C94 VDD1.n29 VSUBS 0.237348f
C95 VTAIL.n0 VSUBS 0.022732f
C96 VTAIL.n1 VSUBS 0.02045f
C97 VTAIL.n2 VSUBS 0.010989f
C98 VTAIL.n3 VSUBS 0.019481f
C99 VTAIL.n4 VSUBS 0.016036f
C100 VTAIL.t2 VSUBS 0.058992f
C101 VTAIL.n5 VSUBS 0.076135f
C102 VTAIL.n6 VSUBS 0.215513f
C103 VTAIL.n7 VSUBS 0.010989f
C104 VTAIL.n8 VSUBS 0.011636f
C105 VTAIL.n9 VSUBS 0.025974f
C106 VTAIL.n10 VSUBS 0.063771f
C107 VTAIL.n11 VSUBS 0.011636f
C108 VTAIL.n12 VSUBS 0.010989f
C109 VTAIL.n13 VSUBS 0.052857f
C110 VTAIL.n14 VSUBS 0.032272f
C111 VTAIL.n15 VSUBS 0.630312f
C112 VTAIL.n16 VSUBS 0.022732f
C113 VTAIL.n17 VSUBS 0.02045f
C114 VTAIL.n18 VSUBS 0.010989f
C115 VTAIL.n19 VSUBS 0.019481f
C116 VTAIL.n20 VSUBS 0.016036f
C117 VTAIL.t1 VSUBS 0.058992f
C118 VTAIL.n21 VSUBS 0.076135f
C119 VTAIL.n22 VSUBS 0.215513f
C120 VTAIL.n23 VSUBS 0.010989f
C121 VTAIL.n24 VSUBS 0.011636f
C122 VTAIL.n25 VSUBS 0.025974f
C123 VTAIL.n26 VSUBS 0.063771f
C124 VTAIL.n27 VSUBS 0.011636f
C125 VTAIL.n28 VSUBS 0.010989f
C126 VTAIL.n29 VSUBS 0.052857f
C127 VTAIL.n30 VSUBS 0.032272f
C128 VTAIL.n31 VSUBS 0.638407f
C129 VTAIL.n32 VSUBS 0.022732f
C130 VTAIL.n33 VSUBS 0.02045f
C131 VTAIL.n34 VSUBS 0.010989f
C132 VTAIL.n35 VSUBS 0.019481f
C133 VTAIL.n36 VSUBS 0.016036f
C134 VTAIL.t3 VSUBS 0.058992f
C135 VTAIL.n37 VSUBS 0.076135f
C136 VTAIL.n38 VSUBS 0.215513f
C137 VTAIL.n39 VSUBS 0.010989f
C138 VTAIL.n40 VSUBS 0.011636f
C139 VTAIL.n41 VSUBS 0.025974f
C140 VTAIL.n42 VSUBS 0.063771f
C141 VTAIL.n43 VSUBS 0.011636f
C142 VTAIL.n44 VSUBS 0.010989f
C143 VTAIL.n45 VSUBS 0.052857f
C144 VTAIL.n46 VSUBS 0.032272f
C145 VTAIL.n47 VSUBS 0.59069f
C146 VTAIL.n48 VSUBS 0.022732f
C147 VTAIL.n49 VSUBS 0.02045f
C148 VTAIL.n50 VSUBS 0.010989f
C149 VTAIL.n51 VSUBS 0.019481f
C150 VTAIL.n52 VSUBS 0.016036f
C151 VTAIL.t0 VSUBS 0.058992f
C152 VTAIL.n53 VSUBS 0.076135f
C153 VTAIL.n54 VSUBS 0.215513f
C154 VTAIL.n55 VSUBS 0.010989f
C155 VTAIL.n56 VSUBS 0.011636f
C156 VTAIL.n57 VSUBS 0.025974f
C157 VTAIL.n58 VSUBS 0.063771f
C158 VTAIL.n59 VSUBS 0.011636f
C159 VTAIL.n60 VSUBS 0.010989f
C160 VTAIL.n61 VSUBS 0.052857f
C161 VTAIL.n62 VSUBS 0.032272f
C162 VTAIL.n63 VSUBS 0.543967f
C163 VP.t1 VSUBS 0.350137f
C164 VP.t0 VSUBS 0.261506f
C165 VP.n0 VSUBS 2.27852f
C166 B.n0 VSUBS 0.005018f
C167 B.n1 VSUBS 0.005018f
C168 B.n2 VSUBS 0.007936f
C169 B.n3 VSUBS 0.007936f
C170 B.n4 VSUBS 0.007936f
C171 B.n5 VSUBS 0.007936f
C172 B.n6 VSUBS 0.007936f
C173 B.n7 VSUBS 0.007936f
C174 B.n8 VSUBS 0.017896f
C175 B.n9 VSUBS 0.007936f
C176 B.n10 VSUBS 0.007936f
C177 B.n11 VSUBS 0.007936f
C178 B.n12 VSUBS 0.007936f
C179 B.n13 VSUBS 0.007936f
C180 B.n14 VSUBS 0.007936f
C181 B.n15 VSUBS 0.007936f
C182 B.n16 VSUBS 0.007236f
C183 B.n17 VSUBS 0.007936f
C184 B.t8 VSUBS 0.055731f
C185 B.t7 VSUBS 0.061875f
C186 B.t6 VSUBS 0.085303f
C187 B.n18 VSUBS 0.111125f
C188 B.n19 VSUBS 0.10341f
C189 B.n20 VSUBS 0.018386f
C190 B.n21 VSUBS 0.007936f
C191 B.n22 VSUBS 0.007936f
C192 B.n23 VSUBS 0.007936f
C193 B.n24 VSUBS 0.007936f
C194 B.t11 VSUBS 0.055731f
C195 B.t10 VSUBS 0.061875f
C196 B.t9 VSUBS 0.085303f
C197 B.n25 VSUBS 0.111124f
C198 B.n26 VSUBS 0.103409f
C199 B.n27 VSUBS 0.007936f
C200 B.n28 VSUBS 0.007936f
C201 B.n29 VSUBS 0.007936f
C202 B.n30 VSUBS 0.007936f
C203 B.n31 VSUBS 0.007936f
C204 B.n32 VSUBS 0.007936f
C205 B.n33 VSUBS 0.007936f
C206 B.n34 VSUBS 0.018982f
C207 B.n35 VSUBS 0.007936f
C208 B.n36 VSUBS 0.007936f
C209 B.n37 VSUBS 0.007936f
C210 B.n38 VSUBS 0.007936f
C211 B.n39 VSUBS 0.007936f
C212 B.n40 VSUBS 0.007936f
C213 B.n41 VSUBS 0.007936f
C214 B.n42 VSUBS 0.007936f
C215 B.n43 VSUBS 0.007936f
C216 B.n44 VSUBS 0.007936f
C217 B.n45 VSUBS 0.007936f
C218 B.n46 VSUBS 0.007936f
C219 B.n47 VSUBS 0.007936f
C220 B.n48 VSUBS 0.018982f
C221 B.n49 VSUBS 0.007936f
C222 B.n50 VSUBS 0.007936f
C223 B.n51 VSUBS 0.007936f
C224 B.n52 VSUBS 0.007936f
C225 B.n53 VSUBS 0.007936f
C226 B.n54 VSUBS 0.007936f
C227 B.n55 VSUBS 0.007936f
C228 B.n56 VSUBS 0.007936f
C229 B.t1 VSUBS 0.055731f
C230 B.t2 VSUBS 0.061875f
C231 B.t0 VSUBS 0.085303f
C232 B.n57 VSUBS 0.111124f
C233 B.n58 VSUBS 0.103409f
C234 B.n59 VSUBS 0.007936f
C235 B.n60 VSUBS 0.007936f
C236 B.n61 VSUBS 0.007936f
C237 B.n62 VSUBS 0.007936f
C238 B.t4 VSUBS 0.055731f
C239 B.t5 VSUBS 0.061875f
C240 B.t3 VSUBS 0.085303f
C241 B.n63 VSUBS 0.111125f
C242 B.n64 VSUBS 0.10341f
C243 B.n65 VSUBS 0.018386f
C244 B.n66 VSUBS 0.007936f
C245 B.n67 VSUBS 0.007936f
C246 B.n68 VSUBS 0.007936f
C247 B.n69 VSUBS 0.007936f
C248 B.n70 VSUBS 0.007936f
C249 B.n71 VSUBS 0.007936f
C250 B.n72 VSUBS 0.007936f
C251 B.n73 VSUBS 0.018982f
C252 B.n74 VSUBS 0.007936f
C253 B.n75 VSUBS 0.007936f
C254 B.n76 VSUBS 0.007936f
C255 B.n77 VSUBS 0.007936f
C256 B.n78 VSUBS 0.007936f
C257 B.n79 VSUBS 0.007936f
C258 B.n80 VSUBS 0.007936f
C259 B.n81 VSUBS 0.007936f
C260 B.n82 VSUBS 0.007936f
C261 B.n83 VSUBS 0.007936f
C262 B.n84 VSUBS 0.007936f
C263 B.n85 VSUBS 0.007936f
C264 B.n86 VSUBS 0.007936f
C265 B.n87 VSUBS 0.007936f
C266 B.n88 VSUBS 0.007936f
C267 B.n89 VSUBS 0.007936f
C268 B.n90 VSUBS 0.007936f
C269 B.n91 VSUBS 0.007936f
C270 B.n92 VSUBS 0.007936f
C271 B.n93 VSUBS 0.007936f
C272 B.n94 VSUBS 0.007936f
C273 B.n95 VSUBS 0.007936f
C274 B.n96 VSUBS 0.017896f
C275 B.n97 VSUBS 0.017896f
C276 B.n98 VSUBS 0.018982f
C277 B.n99 VSUBS 0.007936f
C278 B.n100 VSUBS 0.007936f
C279 B.n101 VSUBS 0.007936f
C280 B.n102 VSUBS 0.007936f
C281 B.n103 VSUBS 0.007936f
C282 B.n104 VSUBS 0.007936f
C283 B.n105 VSUBS 0.007936f
C284 B.n106 VSUBS 0.007936f
C285 B.n107 VSUBS 0.007936f
C286 B.n108 VSUBS 0.007936f
C287 B.n109 VSUBS 0.007936f
C288 B.n110 VSUBS 0.007936f
C289 B.n111 VSUBS 0.007936f
C290 B.n112 VSUBS 0.007936f
C291 B.n113 VSUBS 0.007936f
C292 B.n114 VSUBS 0.007936f
C293 B.n115 VSUBS 0.007936f
C294 B.n116 VSUBS 0.007936f
C295 B.n117 VSUBS 0.007936f
C296 B.n118 VSUBS 0.007936f
C297 B.n119 VSUBS 0.007936f
C298 B.n120 VSUBS 0.007236f
C299 B.n121 VSUBS 0.007936f
C300 B.n122 VSUBS 0.007936f
C301 B.n123 VSUBS 0.004668f
C302 B.n124 VSUBS 0.007936f
C303 B.n125 VSUBS 0.007936f
C304 B.n126 VSUBS 0.007936f
C305 B.n127 VSUBS 0.007936f
C306 B.n128 VSUBS 0.007936f
C307 B.n129 VSUBS 0.007936f
C308 B.n130 VSUBS 0.007936f
C309 B.n131 VSUBS 0.007936f
C310 B.n132 VSUBS 0.007936f
C311 B.n133 VSUBS 0.007936f
C312 B.n134 VSUBS 0.007936f
C313 B.n135 VSUBS 0.007936f
C314 B.n136 VSUBS 0.004668f
C315 B.n137 VSUBS 0.018386f
C316 B.n138 VSUBS 0.007236f
C317 B.n139 VSUBS 0.007936f
C318 B.n140 VSUBS 0.007936f
C319 B.n141 VSUBS 0.007936f
C320 B.n142 VSUBS 0.007936f
C321 B.n143 VSUBS 0.007936f
C322 B.n144 VSUBS 0.007936f
C323 B.n145 VSUBS 0.007936f
C324 B.n146 VSUBS 0.007936f
C325 B.n147 VSUBS 0.007936f
C326 B.n148 VSUBS 0.007936f
C327 B.n149 VSUBS 0.007936f
C328 B.n150 VSUBS 0.007936f
C329 B.n151 VSUBS 0.007936f
C330 B.n152 VSUBS 0.007936f
C331 B.n153 VSUBS 0.007936f
C332 B.n154 VSUBS 0.007936f
C333 B.n155 VSUBS 0.007936f
C334 B.n156 VSUBS 0.007936f
C335 B.n157 VSUBS 0.007936f
C336 B.n158 VSUBS 0.007936f
C337 B.n159 VSUBS 0.007936f
C338 B.n160 VSUBS 0.007936f
C339 B.n161 VSUBS 0.018982f
C340 B.n162 VSUBS 0.017896f
C341 B.n163 VSUBS 0.017896f
C342 B.n164 VSUBS 0.007936f
C343 B.n165 VSUBS 0.007936f
C344 B.n166 VSUBS 0.007936f
C345 B.n167 VSUBS 0.007936f
C346 B.n168 VSUBS 0.007936f
C347 B.n169 VSUBS 0.007936f
C348 B.n170 VSUBS 0.007936f
C349 B.n171 VSUBS 0.007936f
C350 B.n172 VSUBS 0.007936f
C351 B.n173 VSUBS 0.007936f
C352 B.n174 VSUBS 0.007936f
C353 B.n175 VSUBS 0.007936f
C354 B.n176 VSUBS 0.007936f
C355 B.n177 VSUBS 0.007936f
C356 B.n178 VSUBS 0.007936f
C357 B.n179 VSUBS 0.007936f
C358 B.n180 VSUBS 0.007936f
C359 B.n181 VSUBS 0.007936f
C360 B.n182 VSUBS 0.007936f
C361 B.n183 VSUBS 0.007936f
C362 B.n184 VSUBS 0.007936f
C363 B.n185 VSUBS 0.007936f
C364 B.n186 VSUBS 0.007936f
C365 B.n187 VSUBS 0.007936f
C366 B.n188 VSUBS 0.007936f
C367 B.n189 VSUBS 0.007936f
C368 B.n190 VSUBS 0.007936f
C369 B.n191 VSUBS 0.007936f
C370 B.n192 VSUBS 0.007936f
C371 B.n193 VSUBS 0.007936f
C372 B.n194 VSUBS 0.007936f
C373 B.n195 VSUBS 0.007936f
C374 B.n196 VSUBS 0.007936f
C375 B.n197 VSUBS 0.007936f
C376 B.n198 VSUBS 0.007936f
C377 B.n199 VSUBS 0.007936f
C378 B.n200 VSUBS 0.007936f
C379 B.n201 VSUBS 0.017896f
C380 B.n202 VSUBS 0.018843f
C381 B.n203 VSUBS 0.018034f
C382 B.n204 VSUBS 0.007936f
C383 B.n205 VSUBS 0.007936f
C384 B.n206 VSUBS 0.007936f
C385 B.n207 VSUBS 0.007936f
C386 B.n208 VSUBS 0.007936f
C387 B.n209 VSUBS 0.007936f
C388 B.n210 VSUBS 0.007936f
C389 B.n211 VSUBS 0.007936f
C390 B.n212 VSUBS 0.007936f
C391 B.n213 VSUBS 0.007936f
C392 B.n214 VSUBS 0.007936f
C393 B.n215 VSUBS 0.007936f
C394 B.n216 VSUBS 0.007936f
C395 B.n217 VSUBS 0.007936f
C396 B.n218 VSUBS 0.007936f
C397 B.n219 VSUBS 0.007936f
C398 B.n220 VSUBS 0.007936f
C399 B.n221 VSUBS 0.007936f
C400 B.n222 VSUBS 0.007936f
C401 B.n223 VSUBS 0.007936f
C402 B.n224 VSUBS 0.007936f
C403 B.n225 VSUBS 0.007936f
C404 B.n226 VSUBS 0.007236f
C405 B.n227 VSUBS 0.018386f
C406 B.n228 VSUBS 0.004668f
C407 B.n229 VSUBS 0.007936f
C408 B.n230 VSUBS 0.007936f
C409 B.n231 VSUBS 0.007936f
C410 B.n232 VSUBS 0.007936f
C411 B.n233 VSUBS 0.007936f
C412 B.n234 VSUBS 0.007936f
C413 B.n235 VSUBS 0.007936f
C414 B.n236 VSUBS 0.007936f
C415 B.n237 VSUBS 0.007936f
C416 B.n238 VSUBS 0.007936f
C417 B.n239 VSUBS 0.007936f
C418 B.n240 VSUBS 0.007936f
C419 B.n241 VSUBS 0.004668f
C420 B.n242 VSUBS 0.007936f
C421 B.n243 VSUBS 0.007936f
C422 B.n244 VSUBS 0.007936f
C423 B.n245 VSUBS 0.007936f
C424 B.n246 VSUBS 0.007936f
C425 B.n247 VSUBS 0.007936f
C426 B.n248 VSUBS 0.007936f
C427 B.n249 VSUBS 0.007936f
C428 B.n250 VSUBS 0.007936f
C429 B.n251 VSUBS 0.007936f
C430 B.n252 VSUBS 0.007936f
C431 B.n253 VSUBS 0.007936f
C432 B.n254 VSUBS 0.007936f
C433 B.n255 VSUBS 0.007936f
C434 B.n256 VSUBS 0.007936f
C435 B.n257 VSUBS 0.007936f
C436 B.n258 VSUBS 0.007936f
C437 B.n259 VSUBS 0.007936f
C438 B.n260 VSUBS 0.007936f
C439 B.n261 VSUBS 0.007936f
C440 B.n262 VSUBS 0.007936f
C441 B.n263 VSUBS 0.007936f
C442 B.n264 VSUBS 0.007936f
C443 B.n265 VSUBS 0.018982f
C444 B.n266 VSUBS 0.018982f
C445 B.n267 VSUBS 0.017896f
C446 B.n268 VSUBS 0.007936f
C447 B.n269 VSUBS 0.007936f
C448 B.n270 VSUBS 0.007936f
C449 B.n271 VSUBS 0.007936f
C450 B.n272 VSUBS 0.007936f
C451 B.n273 VSUBS 0.007936f
C452 B.n274 VSUBS 0.007936f
C453 B.n275 VSUBS 0.007936f
C454 B.n276 VSUBS 0.007936f
C455 B.n277 VSUBS 0.007936f
C456 B.n278 VSUBS 0.007936f
C457 B.n279 VSUBS 0.007936f
C458 B.n280 VSUBS 0.007936f
C459 B.n281 VSUBS 0.007936f
C460 B.n282 VSUBS 0.007936f
C461 B.n283 VSUBS 0.007936f
C462 B.n284 VSUBS 0.007936f
C463 B.n285 VSUBS 0.007936f
C464 B.n286 VSUBS 0.007936f
C465 B.n287 VSUBS 0.017969f
.ends

