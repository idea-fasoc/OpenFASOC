* NGSPICE file created from diff_pair_sample_0846.ext - technology: sky130A

.subckt diff_pair_sample_0846 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t13 VN.t0 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5382 pd=3.54 as=0.2277 ps=1.71 w=1.38 l=1.65
X1 VTAIL.t12 VN.t1 VDD2.t4 B.t21 sky130_fd_pr__nfet_01v8 ad=0.5382 pd=3.54 as=0.2277 ps=1.71 w=1.38 l=1.65
X2 VDD1.t7 VP.t0 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.5382 ps=3.54 w=1.38 l=1.65
X3 VTAIL.t4 VP.t1 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=1.65
X4 VDD1.t5 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=1.65
X5 VTAIL.t2 VP.t3 VDD1.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5382 pd=3.54 as=0.2277 ps=1.71 w=1.38 l=1.65
X6 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=0.5382 pd=3.54 as=0 ps=0 w=1.38 l=1.65
X7 VDD1.t3 VP.t4 VTAIL.t14 B.t20 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.5382 ps=3.54 w=1.38 l=1.65
X8 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=0.5382 pd=3.54 as=0 ps=0 w=1.38 l=1.65
X9 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5382 pd=3.54 as=0 ps=0 w=1.38 l=1.65
X10 VDD2.t5 VN.t2 VTAIL.t11 B.t20 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.5382 ps=3.54 w=1.38 l=1.65
X11 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.5382 pd=3.54 as=0 ps=0 w=1.38 l=1.65
X12 VDD2.t2 VN.t3 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.5382 ps=3.54 w=1.38 l=1.65
X13 VTAIL.t9 VN.t4 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=1.65
X14 VDD2.t7 VN.t5 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=1.65
X15 VTAIL.t15 VP.t5 VDD1.t2 B.t21 sky130_fd_pr__nfet_01v8 ad=0.5382 pd=3.54 as=0.2277 ps=1.71 w=1.38 l=1.65
X16 VDD2.t0 VN.t6 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=1.65
X17 VTAIL.t6 VN.t7 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=1.65
X18 VTAIL.t1 VP.t6 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=1.65
X19 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.2277 pd=1.71 as=0.2277 ps=1.71 w=1.38 l=1.65
R0 VN.n20 VN.n19 175.071
R1 VN.n41 VN.n40 175.071
R2 VN.n39 VN.n21 161.3
R3 VN.n38 VN.n37 161.3
R4 VN.n36 VN.n22 161.3
R5 VN.n35 VN.n34 161.3
R6 VN.n32 VN.n23 161.3
R7 VN.n31 VN.n30 161.3
R8 VN.n29 VN.n24 161.3
R9 VN.n28 VN.n27 161.3
R10 VN.n18 VN.n0 161.3
R11 VN.n17 VN.n16 161.3
R12 VN.n15 VN.n1 161.3
R13 VN.n14 VN.n13 161.3
R14 VN.n11 VN.n2 161.3
R15 VN.n10 VN.n9 161.3
R16 VN.n8 VN.n3 161.3
R17 VN.n7 VN.n6 161.3
R18 VN.n10 VN.n3 56.5617
R19 VN.n31 VN.n24 56.5617
R20 VN.n17 VN.n1 56.5617
R21 VN.n38 VN.n22 56.5617
R22 VN.n5 VN.n4 54.8557
R23 VN.n26 VN.n25 54.8557
R24 VN.n4 VN.t1 54.3696
R25 VN.n25 VN.t2 54.3696
R26 VN VN.n41 38.76
R27 VN.n6 VN.n3 24.5923
R28 VN.n11 VN.n10 24.5923
R29 VN.n13 VN.n1 24.5923
R30 VN.n18 VN.n17 24.5923
R31 VN.n27 VN.n24 24.5923
R32 VN.n34 VN.n22 24.5923
R33 VN.n32 VN.n31 24.5923
R34 VN.n39 VN.n38 24.5923
R35 VN.n5 VN.t5 20.1569
R36 VN.n12 VN.t7 20.1569
R37 VN.n19 VN.t3 20.1569
R38 VN.n26 VN.t4 20.1569
R39 VN.n33 VN.t6 20.1569
R40 VN.n40 VN.t0 20.1569
R41 VN.n28 VN.n25 17.6839
R42 VN.n7 VN.n4 17.6839
R43 VN.n13 VN.n12 12.7883
R44 VN.n34 VN.n33 12.7883
R45 VN.n6 VN.n5 11.8046
R46 VN.n12 VN.n11 11.8046
R47 VN.n27 VN.n26 11.8046
R48 VN.n33 VN.n32 11.8046
R49 VN.n19 VN.n18 10.8209
R50 VN.n40 VN.n39 10.8209
R51 VN.n41 VN.n21 0.189894
R52 VN.n37 VN.n21 0.189894
R53 VN.n37 VN.n36 0.189894
R54 VN.n36 VN.n35 0.189894
R55 VN.n35 VN.n23 0.189894
R56 VN.n30 VN.n23 0.189894
R57 VN.n30 VN.n29 0.189894
R58 VN.n29 VN.n28 0.189894
R59 VN.n8 VN.n7 0.189894
R60 VN.n9 VN.n8 0.189894
R61 VN.n9 VN.n2 0.189894
R62 VN.n14 VN.n2 0.189894
R63 VN.n15 VN.n14 0.189894
R64 VN.n16 VN.n15 0.189894
R65 VN.n16 VN.n0 0.189894
R66 VN.n20 VN.n0 0.189894
R67 VN VN.n20 0.0516364
R68 VDD2.n2 VDD2.n1 116.034
R69 VDD2.n2 VDD2.n0 116.034
R70 VDD2 VDD2.n5 116.032
R71 VDD2.n4 VDD2.n3 115.237
R72 VDD2.n4 VDD2.n2 32.586
R73 VDD2.n5 VDD2.t3 14.3483
R74 VDD2.n5 VDD2.t5 14.3483
R75 VDD2.n3 VDD2.t1 14.3483
R76 VDD2.n3 VDD2.t0 14.3483
R77 VDD2.n1 VDD2.t6 14.3483
R78 VDD2.n1 VDD2.t2 14.3483
R79 VDD2.n0 VDD2.t4 14.3483
R80 VDD2.n0 VDD2.t7 14.3483
R81 VDD2 VDD2.n4 0.912138
R82 VTAIL.n11 VTAIL.t15 112.906
R83 VTAIL.n10 VTAIL.t11 112.906
R84 VTAIL.n7 VTAIL.t13 112.906
R85 VTAIL.n15 VTAIL.t10 112.906
R86 VTAIL.n2 VTAIL.t12 112.906
R87 VTAIL.n3 VTAIL.t14 112.906
R88 VTAIL.n6 VTAIL.t2 112.906
R89 VTAIL.n14 VTAIL.t5 112.906
R90 VTAIL.n13 VTAIL.n12 98.5581
R91 VTAIL.n9 VTAIL.n8 98.5581
R92 VTAIL.n1 VTAIL.n0 98.558
R93 VTAIL.n5 VTAIL.n4 98.558
R94 VTAIL.n15 VTAIL.n14 15.2634
R95 VTAIL.n7 VTAIL.n6 15.2634
R96 VTAIL.n0 VTAIL.t8 14.3483
R97 VTAIL.n0 VTAIL.t6 14.3483
R98 VTAIL.n4 VTAIL.t3 14.3483
R99 VTAIL.n4 VTAIL.t4 14.3483
R100 VTAIL.n12 VTAIL.t0 14.3483
R101 VTAIL.n12 VTAIL.t1 14.3483
R102 VTAIL.n8 VTAIL.t7 14.3483
R103 VTAIL.n8 VTAIL.t9 14.3483
R104 VTAIL.n9 VTAIL.n7 1.7074
R105 VTAIL.n10 VTAIL.n9 1.7074
R106 VTAIL.n13 VTAIL.n11 1.7074
R107 VTAIL.n14 VTAIL.n13 1.7074
R108 VTAIL.n6 VTAIL.n5 1.7074
R109 VTAIL.n5 VTAIL.n3 1.7074
R110 VTAIL.n2 VTAIL.n1 1.7074
R111 VTAIL VTAIL.n15 1.64921
R112 VTAIL.n11 VTAIL.n10 0.470328
R113 VTAIL.n3 VTAIL.n2 0.470328
R114 VTAIL VTAIL.n1 0.0586897
R115 B.n459 B.n458 585
R116 B.n147 B.n84 585
R117 B.n146 B.n145 585
R118 B.n144 B.n143 585
R119 B.n142 B.n141 585
R120 B.n140 B.n139 585
R121 B.n138 B.n137 585
R122 B.n136 B.n135 585
R123 B.n134 B.n133 585
R124 B.n132 B.n131 585
R125 B.n130 B.n129 585
R126 B.n128 B.n127 585
R127 B.n126 B.n125 585
R128 B.n124 B.n123 585
R129 B.n122 B.n121 585
R130 B.n120 B.n119 585
R131 B.n118 B.n117 585
R132 B.n116 B.n115 585
R133 B.n114 B.n113 585
R134 B.n112 B.n111 585
R135 B.n110 B.n109 585
R136 B.n108 B.n107 585
R137 B.n106 B.n105 585
R138 B.n104 B.n103 585
R139 B.n102 B.n101 585
R140 B.n100 B.n99 585
R141 B.n98 B.n97 585
R142 B.n96 B.n95 585
R143 B.n94 B.n93 585
R144 B.n92 B.n91 585
R145 B.n457 B.n69 585
R146 B.n462 B.n69 585
R147 B.n456 B.n68 585
R148 B.n463 B.n68 585
R149 B.n455 B.n454 585
R150 B.n454 B.n64 585
R151 B.n453 B.n63 585
R152 B.n469 B.n63 585
R153 B.n452 B.n62 585
R154 B.n470 B.n62 585
R155 B.n451 B.n61 585
R156 B.n471 B.n61 585
R157 B.n450 B.n449 585
R158 B.n449 B.n57 585
R159 B.n448 B.n56 585
R160 B.n477 B.n56 585
R161 B.n447 B.n55 585
R162 B.n478 B.n55 585
R163 B.n446 B.n54 585
R164 B.n479 B.n54 585
R165 B.n445 B.n444 585
R166 B.n444 B.n50 585
R167 B.n443 B.n49 585
R168 B.n485 B.n49 585
R169 B.n442 B.n48 585
R170 B.n486 B.n48 585
R171 B.n441 B.n47 585
R172 B.n487 B.n47 585
R173 B.n440 B.n439 585
R174 B.n439 B.n43 585
R175 B.n438 B.n42 585
R176 B.n493 B.n42 585
R177 B.n437 B.n41 585
R178 B.n494 B.n41 585
R179 B.n436 B.n40 585
R180 B.n495 B.n40 585
R181 B.n435 B.n434 585
R182 B.n434 B.n36 585
R183 B.n433 B.n35 585
R184 B.n501 B.n35 585
R185 B.n432 B.n34 585
R186 B.n502 B.n34 585
R187 B.n431 B.n33 585
R188 B.n503 B.n33 585
R189 B.n430 B.n429 585
R190 B.n429 B.n29 585
R191 B.n428 B.n28 585
R192 B.n509 B.n28 585
R193 B.n427 B.n27 585
R194 B.n510 B.n27 585
R195 B.n426 B.n26 585
R196 B.n511 B.n26 585
R197 B.n425 B.n424 585
R198 B.n424 B.n25 585
R199 B.n423 B.n21 585
R200 B.n517 B.n21 585
R201 B.n422 B.n20 585
R202 B.n518 B.n20 585
R203 B.n421 B.n19 585
R204 B.n519 B.n19 585
R205 B.n420 B.n419 585
R206 B.n419 B.n15 585
R207 B.n418 B.n14 585
R208 B.n525 B.n14 585
R209 B.n417 B.n13 585
R210 B.n526 B.n13 585
R211 B.n416 B.n12 585
R212 B.n527 B.n12 585
R213 B.n415 B.n414 585
R214 B.n414 B.n8 585
R215 B.n413 B.n7 585
R216 B.n533 B.n7 585
R217 B.n412 B.n6 585
R218 B.n534 B.n6 585
R219 B.n411 B.n5 585
R220 B.n535 B.n5 585
R221 B.n410 B.n409 585
R222 B.n409 B.n4 585
R223 B.n408 B.n148 585
R224 B.n408 B.n407 585
R225 B.n398 B.n149 585
R226 B.n150 B.n149 585
R227 B.n400 B.n399 585
R228 B.n401 B.n400 585
R229 B.n397 B.n154 585
R230 B.n158 B.n154 585
R231 B.n396 B.n395 585
R232 B.n395 B.n394 585
R233 B.n156 B.n155 585
R234 B.n157 B.n156 585
R235 B.n387 B.n386 585
R236 B.n388 B.n387 585
R237 B.n385 B.n163 585
R238 B.n163 B.n162 585
R239 B.n384 B.n383 585
R240 B.n383 B.n382 585
R241 B.n165 B.n164 585
R242 B.n375 B.n165 585
R243 B.n374 B.n373 585
R244 B.n376 B.n374 585
R245 B.n372 B.n170 585
R246 B.n170 B.n169 585
R247 B.n371 B.n370 585
R248 B.n370 B.n369 585
R249 B.n172 B.n171 585
R250 B.n173 B.n172 585
R251 B.n362 B.n361 585
R252 B.n363 B.n362 585
R253 B.n360 B.n177 585
R254 B.n181 B.n177 585
R255 B.n359 B.n358 585
R256 B.n358 B.n357 585
R257 B.n179 B.n178 585
R258 B.n180 B.n179 585
R259 B.n350 B.n349 585
R260 B.n351 B.n350 585
R261 B.n348 B.n186 585
R262 B.n186 B.n185 585
R263 B.n347 B.n346 585
R264 B.n346 B.n345 585
R265 B.n188 B.n187 585
R266 B.n189 B.n188 585
R267 B.n338 B.n337 585
R268 B.n339 B.n338 585
R269 B.n336 B.n194 585
R270 B.n194 B.n193 585
R271 B.n335 B.n334 585
R272 B.n334 B.n333 585
R273 B.n196 B.n195 585
R274 B.n197 B.n196 585
R275 B.n326 B.n325 585
R276 B.n327 B.n326 585
R277 B.n324 B.n202 585
R278 B.n202 B.n201 585
R279 B.n323 B.n322 585
R280 B.n322 B.n321 585
R281 B.n204 B.n203 585
R282 B.n205 B.n204 585
R283 B.n314 B.n313 585
R284 B.n315 B.n314 585
R285 B.n312 B.n210 585
R286 B.n210 B.n209 585
R287 B.n311 B.n310 585
R288 B.n310 B.n309 585
R289 B.n212 B.n211 585
R290 B.n213 B.n212 585
R291 B.n302 B.n301 585
R292 B.n303 B.n302 585
R293 B.n300 B.n218 585
R294 B.n218 B.n217 585
R295 B.n295 B.n294 585
R296 B.n293 B.n235 585
R297 B.n292 B.n234 585
R298 B.n297 B.n234 585
R299 B.n291 B.n290 585
R300 B.n289 B.n288 585
R301 B.n287 B.n286 585
R302 B.n285 B.n284 585
R303 B.n283 B.n282 585
R304 B.n281 B.n280 585
R305 B.n279 B.n278 585
R306 B.n276 B.n275 585
R307 B.n274 B.n273 585
R308 B.n272 B.n271 585
R309 B.n270 B.n269 585
R310 B.n268 B.n267 585
R311 B.n266 B.n265 585
R312 B.n264 B.n263 585
R313 B.n262 B.n261 585
R314 B.n260 B.n259 585
R315 B.n258 B.n257 585
R316 B.n255 B.n254 585
R317 B.n253 B.n252 585
R318 B.n251 B.n250 585
R319 B.n249 B.n248 585
R320 B.n247 B.n246 585
R321 B.n245 B.n244 585
R322 B.n243 B.n242 585
R323 B.n241 B.n240 585
R324 B.n220 B.n219 585
R325 B.n299 B.n298 585
R326 B.n298 B.n297 585
R327 B.n216 B.n215 585
R328 B.n217 B.n216 585
R329 B.n305 B.n304 585
R330 B.n304 B.n303 585
R331 B.n306 B.n214 585
R332 B.n214 B.n213 585
R333 B.n308 B.n307 585
R334 B.n309 B.n308 585
R335 B.n208 B.n207 585
R336 B.n209 B.n208 585
R337 B.n317 B.n316 585
R338 B.n316 B.n315 585
R339 B.n318 B.n206 585
R340 B.n206 B.n205 585
R341 B.n320 B.n319 585
R342 B.n321 B.n320 585
R343 B.n200 B.n199 585
R344 B.n201 B.n200 585
R345 B.n329 B.n328 585
R346 B.n328 B.n327 585
R347 B.n330 B.n198 585
R348 B.n198 B.n197 585
R349 B.n332 B.n331 585
R350 B.n333 B.n332 585
R351 B.n192 B.n191 585
R352 B.n193 B.n192 585
R353 B.n341 B.n340 585
R354 B.n340 B.n339 585
R355 B.n342 B.n190 585
R356 B.n190 B.n189 585
R357 B.n344 B.n343 585
R358 B.n345 B.n344 585
R359 B.n184 B.n183 585
R360 B.n185 B.n184 585
R361 B.n353 B.n352 585
R362 B.n352 B.n351 585
R363 B.n354 B.n182 585
R364 B.n182 B.n180 585
R365 B.n356 B.n355 585
R366 B.n357 B.n356 585
R367 B.n176 B.n175 585
R368 B.n181 B.n176 585
R369 B.n365 B.n364 585
R370 B.n364 B.n363 585
R371 B.n366 B.n174 585
R372 B.n174 B.n173 585
R373 B.n368 B.n367 585
R374 B.n369 B.n368 585
R375 B.n168 B.n167 585
R376 B.n169 B.n168 585
R377 B.n378 B.n377 585
R378 B.n377 B.n376 585
R379 B.n379 B.n166 585
R380 B.n375 B.n166 585
R381 B.n381 B.n380 585
R382 B.n382 B.n381 585
R383 B.n161 B.n160 585
R384 B.n162 B.n161 585
R385 B.n390 B.n389 585
R386 B.n389 B.n388 585
R387 B.n391 B.n159 585
R388 B.n159 B.n157 585
R389 B.n393 B.n392 585
R390 B.n394 B.n393 585
R391 B.n153 B.n152 585
R392 B.n158 B.n153 585
R393 B.n403 B.n402 585
R394 B.n402 B.n401 585
R395 B.n404 B.n151 585
R396 B.n151 B.n150 585
R397 B.n406 B.n405 585
R398 B.n407 B.n406 585
R399 B.n2 B.n0 585
R400 B.n4 B.n2 585
R401 B.n3 B.n1 585
R402 B.n534 B.n3 585
R403 B.n532 B.n531 585
R404 B.n533 B.n532 585
R405 B.n530 B.n9 585
R406 B.n9 B.n8 585
R407 B.n529 B.n528 585
R408 B.n528 B.n527 585
R409 B.n11 B.n10 585
R410 B.n526 B.n11 585
R411 B.n524 B.n523 585
R412 B.n525 B.n524 585
R413 B.n522 B.n16 585
R414 B.n16 B.n15 585
R415 B.n521 B.n520 585
R416 B.n520 B.n519 585
R417 B.n18 B.n17 585
R418 B.n518 B.n18 585
R419 B.n516 B.n515 585
R420 B.n517 B.n516 585
R421 B.n514 B.n22 585
R422 B.n25 B.n22 585
R423 B.n513 B.n512 585
R424 B.n512 B.n511 585
R425 B.n24 B.n23 585
R426 B.n510 B.n24 585
R427 B.n508 B.n507 585
R428 B.n509 B.n508 585
R429 B.n506 B.n30 585
R430 B.n30 B.n29 585
R431 B.n505 B.n504 585
R432 B.n504 B.n503 585
R433 B.n32 B.n31 585
R434 B.n502 B.n32 585
R435 B.n500 B.n499 585
R436 B.n501 B.n500 585
R437 B.n498 B.n37 585
R438 B.n37 B.n36 585
R439 B.n497 B.n496 585
R440 B.n496 B.n495 585
R441 B.n39 B.n38 585
R442 B.n494 B.n39 585
R443 B.n492 B.n491 585
R444 B.n493 B.n492 585
R445 B.n490 B.n44 585
R446 B.n44 B.n43 585
R447 B.n489 B.n488 585
R448 B.n488 B.n487 585
R449 B.n46 B.n45 585
R450 B.n486 B.n46 585
R451 B.n484 B.n483 585
R452 B.n485 B.n484 585
R453 B.n482 B.n51 585
R454 B.n51 B.n50 585
R455 B.n481 B.n480 585
R456 B.n480 B.n479 585
R457 B.n53 B.n52 585
R458 B.n478 B.n53 585
R459 B.n476 B.n475 585
R460 B.n477 B.n476 585
R461 B.n474 B.n58 585
R462 B.n58 B.n57 585
R463 B.n473 B.n472 585
R464 B.n472 B.n471 585
R465 B.n60 B.n59 585
R466 B.n470 B.n60 585
R467 B.n468 B.n467 585
R468 B.n469 B.n468 585
R469 B.n466 B.n65 585
R470 B.n65 B.n64 585
R471 B.n465 B.n464 585
R472 B.n464 B.n463 585
R473 B.n67 B.n66 585
R474 B.n462 B.n67 585
R475 B.n537 B.n536 585
R476 B.n536 B.n535 585
R477 B.n295 B.n216 564.573
R478 B.n91 B.n67 564.573
R479 B.n298 B.n218 564.573
R480 B.n459 B.n69 564.573
R481 B.n461 B.n460 256.663
R482 B.n461 B.n83 256.663
R483 B.n461 B.n82 256.663
R484 B.n461 B.n81 256.663
R485 B.n461 B.n80 256.663
R486 B.n461 B.n79 256.663
R487 B.n461 B.n78 256.663
R488 B.n461 B.n77 256.663
R489 B.n461 B.n76 256.663
R490 B.n461 B.n75 256.663
R491 B.n461 B.n74 256.663
R492 B.n461 B.n73 256.663
R493 B.n461 B.n72 256.663
R494 B.n461 B.n71 256.663
R495 B.n461 B.n70 256.663
R496 B.n297 B.n296 256.663
R497 B.n297 B.n221 256.663
R498 B.n297 B.n222 256.663
R499 B.n297 B.n223 256.663
R500 B.n297 B.n224 256.663
R501 B.n297 B.n225 256.663
R502 B.n297 B.n226 256.663
R503 B.n297 B.n227 256.663
R504 B.n297 B.n228 256.663
R505 B.n297 B.n229 256.663
R506 B.n297 B.n230 256.663
R507 B.n297 B.n231 256.663
R508 B.n297 B.n232 256.663
R509 B.n297 B.n233 256.663
R510 B.n297 B.n217 229.752
R511 B.n462 B.n461 229.752
R512 B.n238 B.t10 226.114
R513 B.n236 B.t6 226.114
R514 B.n88 B.t17 226.114
R515 B.n85 B.t13 226.114
R516 B.n304 B.n216 163.367
R517 B.n304 B.n214 163.367
R518 B.n308 B.n214 163.367
R519 B.n308 B.n208 163.367
R520 B.n316 B.n208 163.367
R521 B.n316 B.n206 163.367
R522 B.n320 B.n206 163.367
R523 B.n320 B.n200 163.367
R524 B.n328 B.n200 163.367
R525 B.n328 B.n198 163.367
R526 B.n332 B.n198 163.367
R527 B.n332 B.n192 163.367
R528 B.n340 B.n192 163.367
R529 B.n340 B.n190 163.367
R530 B.n344 B.n190 163.367
R531 B.n344 B.n184 163.367
R532 B.n352 B.n184 163.367
R533 B.n352 B.n182 163.367
R534 B.n356 B.n182 163.367
R535 B.n356 B.n176 163.367
R536 B.n364 B.n176 163.367
R537 B.n364 B.n174 163.367
R538 B.n368 B.n174 163.367
R539 B.n368 B.n168 163.367
R540 B.n377 B.n168 163.367
R541 B.n377 B.n166 163.367
R542 B.n381 B.n166 163.367
R543 B.n381 B.n161 163.367
R544 B.n389 B.n161 163.367
R545 B.n389 B.n159 163.367
R546 B.n393 B.n159 163.367
R547 B.n393 B.n153 163.367
R548 B.n402 B.n153 163.367
R549 B.n402 B.n151 163.367
R550 B.n406 B.n151 163.367
R551 B.n406 B.n2 163.367
R552 B.n536 B.n2 163.367
R553 B.n536 B.n3 163.367
R554 B.n532 B.n3 163.367
R555 B.n532 B.n9 163.367
R556 B.n528 B.n9 163.367
R557 B.n528 B.n11 163.367
R558 B.n524 B.n11 163.367
R559 B.n524 B.n16 163.367
R560 B.n520 B.n16 163.367
R561 B.n520 B.n18 163.367
R562 B.n516 B.n18 163.367
R563 B.n516 B.n22 163.367
R564 B.n512 B.n22 163.367
R565 B.n512 B.n24 163.367
R566 B.n508 B.n24 163.367
R567 B.n508 B.n30 163.367
R568 B.n504 B.n30 163.367
R569 B.n504 B.n32 163.367
R570 B.n500 B.n32 163.367
R571 B.n500 B.n37 163.367
R572 B.n496 B.n37 163.367
R573 B.n496 B.n39 163.367
R574 B.n492 B.n39 163.367
R575 B.n492 B.n44 163.367
R576 B.n488 B.n44 163.367
R577 B.n488 B.n46 163.367
R578 B.n484 B.n46 163.367
R579 B.n484 B.n51 163.367
R580 B.n480 B.n51 163.367
R581 B.n480 B.n53 163.367
R582 B.n476 B.n53 163.367
R583 B.n476 B.n58 163.367
R584 B.n472 B.n58 163.367
R585 B.n472 B.n60 163.367
R586 B.n468 B.n60 163.367
R587 B.n468 B.n65 163.367
R588 B.n464 B.n65 163.367
R589 B.n464 B.n67 163.367
R590 B.n235 B.n234 163.367
R591 B.n290 B.n234 163.367
R592 B.n288 B.n287 163.367
R593 B.n284 B.n283 163.367
R594 B.n280 B.n279 163.367
R595 B.n275 B.n274 163.367
R596 B.n271 B.n270 163.367
R597 B.n267 B.n266 163.367
R598 B.n263 B.n262 163.367
R599 B.n259 B.n258 163.367
R600 B.n254 B.n253 163.367
R601 B.n250 B.n249 163.367
R602 B.n246 B.n245 163.367
R603 B.n242 B.n241 163.367
R604 B.n298 B.n220 163.367
R605 B.n302 B.n218 163.367
R606 B.n302 B.n212 163.367
R607 B.n310 B.n212 163.367
R608 B.n310 B.n210 163.367
R609 B.n314 B.n210 163.367
R610 B.n314 B.n204 163.367
R611 B.n322 B.n204 163.367
R612 B.n322 B.n202 163.367
R613 B.n326 B.n202 163.367
R614 B.n326 B.n196 163.367
R615 B.n334 B.n196 163.367
R616 B.n334 B.n194 163.367
R617 B.n338 B.n194 163.367
R618 B.n338 B.n188 163.367
R619 B.n346 B.n188 163.367
R620 B.n346 B.n186 163.367
R621 B.n350 B.n186 163.367
R622 B.n350 B.n179 163.367
R623 B.n358 B.n179 163.367
R624 B.n358 B.n177 163.367
R625 B.n362 B.n177 163.367
R626 B.n362 B.n172 163.367
R627 B.n370 B.n172 163.367
R628 B.n370 B.n170 163.367
R629 B.n374 B.n170 163.367
R630 B.n374 B.n165 163.367
R631 B.n383 B.n165 163.367
R632 B.n383 B.n163 163.367
R633 B.n387 B.n163 163.367
R634 B.n387 B.n156 163.367
R635 B.n395 B.n156 163.367
R636 B.n395 B.n154 163.367
R637 B.n400 B.n154 163.367
R638 B.n400 B.n149 163.367
R639 B.n408 B.n149 163.367
R640 B.n409 B.n408 163.367
R641 B.n409 B.n5 163.367
R642 B.n6 B.n5 163.367
R643 B.n7 B.n6 163.367
R644 B.n414 B.n7 163.367
R645 B.n414 B.n12 163.367
R646 B.n13 B.n12 163.367
R647 B.n14 B.n13 163.367
R648 B.n419 B.n14 163.367
R649 B.n419 B.n19 163.367
R650 B.n20 B.n19 163.367
R651 B.n21 B.n20 163.367
R652 B.n424 B.n21 163.367
R653 B.n424 B.n26 163.367
R654 B.n27 B.n26 163.367
R655 B.n28 B.n27 163.367
R656 B.n429 B.n28 163.367
R657 B.n429 B.n33 163.367
R658 B.n34 B.n33 163.367
R659 B.n35 B.n34 163.367
R660 B.n434 B.n35 163.367
R661 B.n434 B.n40 163.367
R662 B.n41 B.n40 163.367
R663 B.n42 B.n41 163.367
R664 B.n439 B.n42 163.367
R665 B.n439 B.n47 163.367
R666 B.n48 B.n47 163.367
R667 B.n49 B.n48 163.367
R668 B.n444 B.n49 163.367
R669 B.n444 B.n54 163.367
R670 B.n55 B.n54 163.367
R671 B.n56 B.n55 163.367
R672 B.n449 B.n56 163.367
R673 B.n449 B.n61 163.367
R674 B.n62 B.n61 163.367
R675 B.n63 B.n62 163.367
R676 B.n454 B.n63 163.367
R677 B.n454 B.n68 163.367
R678 B.n69 B.n68 163.367
R679 B.n95 B.n94 163.367
R680 B.n99 B.n98 163.367
R681 B.n103 B.n102 163.367
R682 B.n107 B.n106 163.367
R683 B.n111 B.n110 163.367
R684 B.n115 B.n114 163.367
R685 B.n119 B.n118 163.367
R686 B.n123 B.n122 163.367
R687 B.n127 B.n126 163.367
R688 B.n131 B.n130 163.367
R689 B.n135 B.n134 163.367
R690 B.n139 B.n138 163.367
R691 B.n143 B.n142 163.367
R692 B.n145 B.n84 163.367
R693 B.n238 B.t12 144.56
R694 B.n85 B.t15 144.56
R695 B.n236 B.t9 144.56
R696 B.n88 B.t18 144.56
R697 B.n303 B.n217 112.397
R698 B.n303 B.n213 112.397
R699 B.n309 B.n213 112.397
R700 B.n309 B.n209 112.397
R701 B.n315 B.n209 112.397
R702 B.n321 B.n205 112.397
R703 B.n321 B.n201 112.397
R704 B.n327 B.n201 112.397
R705 B.n327 B.n197 112.397
R706 B.n333 B.n197 112.397
R707 B.n333 B.n193 112.397
R708 B.n339 B.n193 112.397
R709 B.n339 B.n189 112.397
R710 B.n345 B.n189 112.397
R711 B.n351 B.n185 112.397
R712 B.n351 B.n180 112.397
R713 B.n357 B.n180 112.397
R714 B.n357 B.n181 112.397
R715 B.n363 B.n173 112.397
R716 B.n369 B.n173 112.397
R717 B.n369 B.n169 112.397
R718 B.n376 B.n169 112.397
R719 B.n376 B.n375 112.397
R720 B.n382 B.n162 112.397
R721 B.n388 B.n162 112.397
R722 B.n388 B.n157 112.397
R723 B.n394 B.n157 112.397
R724 B.n394 B.n158 112.397
R725 B.n401 B.n150 112.397
R726 B.n407 B.n150 112.397
R727 B.n407 B.n4 112.397
R728 B.n535 B.n4 112.397
R729 B.n535 B.n534 112.397
R730 B.n534 B.n533 112.397
R731 B.n533 B.n8 112.397
R732 B.n527 B.n8 112.397
R733 B.n526 B.n525 112.397
R734 B.n525 B.n15 112.397
R735 B.n519 B.n15 112.397
R736 B.n519 B.n518 112.397
R737 B.n518 B.n517 112.397
R738 B.n511 B.n25 112.397
R739 B.n511 B.n510 112.397
R740 B.n510 B.n509 112.397
R741 B.n509 B.n29 112.397
R742 B.n503 B.n29 112.397
R743 B.n502 B.n501 112.397
R744 B.n501 B.n36 112.397
R745 B.n495 B.n36 112.397
R746 B.n495 B.n494 112.397
R747 B.n493 B.n43 112.397
R748 B.n487 B.n43 112.397
R749 B.n487 B.n486 112.397
R750 B.n486 B.n485 112.397
R751 B.n485 B.n50 112.397
R752 B.n479 B.n50 112.397
R753 B.n479 B.n478 112.397
R754 B.n478 B.n477 112.397
R755 B.n477 B.n57 112.397
R756 B.n471 B.n470 112.397
R757 B.n470 B.n469 112.397
R758 B.n469 B.n64 112.397
R759 B.n463 B.n64 112.397
R760 B.n463 B.n462 112.397
R761 B.n315 B.t7 110.745
R762 B.t2 B.n185 110.745
R763 B.n494 B.t5 110.745
R764 B.n471 B.t14 110.745
R765 B.n239 B.t11 106.159
R766 B.n86 B.t16 106.159
R767 B.n237 B.t8 106.159
R768 B.n89 B.t19 106.159
R769 B.n181 B.t3 94.2154
R770 B.t1 B.n502 94.2154
R771 B.n375 B.t4 74.3807
R772 B.n25 B.t0 74.3807
R773 B.n296 B.n295 71.676
R774 B.n290 B.n221 71.676
R775 B.n287 B.n222 71.676
R776 B.n283 B.n223 71.676
R777 B.n279 B.n224 71.676
R778 B.n274 B.n225 71.676
R779 B.n270 B.n226 71.676
R780 B.n266 B.n227 71.676
R781 B.n262 B.n228 71.676
R782 B.n258 B.n229 71.676
R783 B.n253 B.n230 71.676
R784 B.n249 B.n231 71.676
R785 B.n245 B.n232 71.676
R786 B.n241 B.n233 71.676
R787 B.n91 B.n70 71.676
R788 B.n95 B.n71 71.676
R789 B.n99 B.n72 71.676
R790 B.n103 B.n73 71.676
R791 B.n107 B.n74 71.676
R792 B.n111 B.n75 71.676
R793 B.n115 B.n76 71.676
R794 B.n119 B.n77 71.676
R795 B.n123 B.n78 71.676
R796 B.n127 B.n79 71.676
R797 B.n131 B.n80 71.676
R798 B.n135 B.n81 71.676
R799 B.n139 B.n82 71.676
R800 B.n143 B.n83 71.676
R801 B.n460 B.n84 71.676
R802 B.n460 B.n459 71.676
R803 B.n145 B.n83 71.676
R804 B.n142 B.n82 71.676
R805 B.n138 B.n81 71.676
R806 B.n134 B.n80 71.676
R807 B.n130 B.n79 71.676
R808 B.n126 B.n78 71.676
R809 B.n122 B.n77 71.676
R810 B.n118 B.n76 71.676
R811 B.n114 B.n75 71.676
R812 B.n110 B.n74 71.676
R813 B.n106 B.n73 71.676
R814 B.n102 B.n72 71.676
R815 B.n98 B.n71 71.676
R816 B.n94 B.n70 71.676
R817 B.n296 B.n235 71.676
R818 B.n288 B.n221 71.676
R819 B.n284 B.n222 71.676
R820 B.n280 B.n223 71.676
R821 B.n275 B.n224 71.676
R822 B.n271 B.n225 71.676
R823 B.n267 B.n226 71.676
R824 B.n263 B.n227 71.676
R825 B.n259 B.n228 71.676
R826 B.n254 B.n229 71.676
R827 B.n250 B.n230 71.676
R828 B.n246 B.n231 71.676
R829 B.n242 B.n232 71.676
R830 B.n233 B.n220 71.676
R831 B.n256 B.n239 59.5399
R832 B.n277 B.n237 59.5399
R833 B.n90 B.n89 59.5399
R834 B.n87 B.n86 59.5399
R835 B.n401 B.t20 57.8517
R836 B.n527 B.t21 57.8517
R837 B.n158 B.t20 54.546
R838 B.t21 B.n526 54.546
R839 B.n239 B.n238 38.4005
R840 B.n237 B.n236 38.4005
R841 B.n89 B.n88 38.4005
R842 B.n86 B.n85 38.4005
R843 B.n382 B.t4 38.017
R844 B.n517 B.t0 38.017
R845 B.n92 B.n66 36.6834
R846 B.n458 B.n457 36.6834
R847 B.n300 B.n299 36.6834
R848 B.n294 B.n215 36.6834
R849 B.n363 B.t3 18.1823
R850 B.n503 B.t1 18.1823
R851 B B.n537 18.0485
R852 B.n93 B.n92 10.6151
R853 B.n96 B.n93 10.6151
R854 B.n97 B.n96 10.6151
R855 B.n100 B.n97 10.6151
R856 B.n101 B.n100 10.6151
R857 B.n104 B.n101 10.6151
R858 B.n105 B.n104 10.6151
R859 B.n108 B.n105 10.6151
R860 B.n109 B.n108 10.6151
R861 B.n113 B.n112 10.6151
R862 B.n116 B.n113 10.6151
R863 B.n117 B.n116 10.6151
R864 B.n120 B.n117 10.6151
R865 B.n121 B.n120 10.6151
R866 B.n124 B.n121 10.6151
R867 B.n125 B.n124 10.6151
R868 B.n128 B.n125 10.6151
R869 B.n129 B.n128 10.6151
R870 B.n133 B.n132 10.6151
R871 B.n136 B.n133 10.6151
R872 B.n137 B.n136 10.6151
R873 B.n140 B.n137 10.6151
R874 B.n141 B.n140 10.6151
R875 B.n144 B.n141 10.6151
R876 B.n146 B.n144 10.6151
R877 B.n147 B.n146 10.6151
R878 B.n458 B.n147 10.6151
R879 B.n301 B.n300 10.6151
R880 B.n301 B.n211 10.6151
R881 B.n311 B.n211 10.6151
R882 B.n312 B.n311 10.6151
R883 B.n313 B.n312 10.6151
R884 B.n313 B.n203 10.6151
R885 B.n323 B.n203 10.6151
R886 B.n324 B.n323 10.6151
R887 B.n325 B.n324 10.6151
R888 B.n325 B.n195 10.6151
R889 B.n335 B.n195 10.6151
R890 B.n336 B.n335 10.6151
R891 B.n337 B.n336 10.6151
R892 B.n337 B.n187 10.6151
R893 B.n347 B.n187 10.6151
R894 B.n348 B.n347 10.6151
R895 B.n349 B.n348 10.6151
R896 B.n349 B.n178 10.6151
R897 B.n359 B.n178 10.6151
R898 B.n360 B.n359 10.6151
R899 B.n361 B.n360 10.6151
R900 B.n361 B.n171 10.6151
R901 B.n371 B.n171 10.6151
R902 B.n372 B.n371 10.6151
R903 B.n373 B.n372 10.6151
R904 B.n373 B.n164 10.6151
R905 B.n384 B.n164 10.6151
R906 B.n385 B.n384 10.6151
R907 B.n386 B.n385 10.6151
R908 B.n386 B.n155 10.6151
R909 B.n396 B.n155 10.6151
R910 B.n397 B.n396 10.6151
R911 B.n399 B.n397 10.6151
R912 B.n399 B.n398 10.6151
R913 B.n398 B.n148 10.6151
R914 B.n410 B.n148 10.6151
R915 B.n411 B.n410 10.6151
R916 B.n412 B.n411 10.6151
R917 B.n413 B.n412 10.6151
R918 B.n415 B.n413 10.6151
R919 B.n416 B.n415 10.6151
R920 B.n417 B.n416 10.6151
R921 B.n418 B.n417 10.6151
R922 B.n420 B.n418 10.6151
R923 B.n421 B.n420 10.6151
R924 B.n422 B.n421 10.6151
R925 B.n423 B.n422 10.6151
R926 B.n425 B.n423 10.6151
R927 B.n426 B.n425 10.6151
R928 B.n427 B.n426 10.6151
R929 B.n428 B.n427 10.6151
R930 B.n430 B.n428 10.6151
R931 B.n431 B.n430 10.6151
R932 B.n432 B.n431 10.6151
R933 B.n433 B.n432 10.6151
R934 B.n435 B.n433 10.6151
R935 B.n436 B.n435 10.6151
R936 B.n437 B.n436 10.6151
R937 B.n438 B.n437 10.6151
R938 B.n440 B.n438 10.6151
R939 B.n441 B.n440 10.6151
R940 B.n442 B.n441 10.6151
R941 B.n443 B.n442 10.6151
R942 B.n445 B.n443 10.6151
R943 B.n446 B.n445 10.6151
R944 B.n447 B.n446 10.6151
R945 B.n448 B.n447 10.6151
R946 B.n450 B.n448 10.6151
R947 B.n451 B.n450 10.6151
R948 B.n452 B.n451 10.6151
R949 B.n453 B.n452 10.6151
R950 B.n455 B.n453 10.6151
R951 B.n456 B.n455 10.6151
R952 B.n457 B.n456 10.6151
R953 B.n294 B.n293 10.6151
R954 B.n293 B.n292 10.6151
R955 B.n292 B.n291 10.6151
R956 B.n291 B.n289 10.6151
R957 B.n289 B.n286 10.6151
R958 B.n286 B.n285 10.6151
R959 B.n285 B.n282 10.6151
R960 B.n282 B.n281 10.6151
R961 B.n281 B.n278 10.6151
R962 B.n276 B.n273 10.6151
R963 B.n273 B.n272 10.6151
R964 B.n272 B.n269 10.6151
R965 B.n269 B.n268 10.6151
R966 B.n268 B.n265 10.6151
R967 B.n265 B.n264 10.6151
R968 B.n264 B.n261 10.6151
R969 B.n261 B.n260 10.6151
R970 B.n260 B.n257 10.6151
R971 B.n255 B.n252 10.6151
R972 B.n252 B.n251 10.6151
R973 B.n251 B.n248 10.6151
R974 B.n248 B.n247 10.6151
R975 B.n247 B.n244 10.6151
R976 B.n244 B.n243 10.6151
R977 B.n243 B.n240 10.6151
R978 B.n240 B.n219 10.6151
R979 B.n299 B.n219 10.6151
R980 B.n305 B.n215 10.6151
R981 B.n306 B.n305 10.6151
R982 B.n307 B.n306 10.6151
R983 B.n307 B.n207 10.6151
R984 B.n317 B.n207 10.6151
R985 B.n318 B.n317 10.6151
R986 B.n319 B.n318 10.6151
R987 B.n319 B.n199 10.6151
R988 B.n329 B.n199 10.6151
R989 B.n330 B.n329 10.6151
R990 B.n331 B.n330 10.6151
R991 B.n331 B.n191 10.6151
R992 B.n341 B.n191 10.6151
R993 B.n342 B.n341 10.6151
R994 B.n343 B.n342 10.6151
R995 B.n343 B.n183 10.6151
R996 B.n353 B.n183 10.6151
R997 B.n354 B.n353 10.6151
R998 B.n355 B.n354 10.6151
R999 B.n355 B.n175 10.6151
R1000 B.n365 B.n175 10.6151
R1001 B.n366 B.n365 10.6151
R1002 B.n367 B.n366 10.6151
R1003 B.n367 B.n167 10.6151
R1004 B.n378 B.n167 10.6151
R1005 B.n379 B.n378 10.6151
R1006 B.n380 B.n379 10.6151
R1007 B.n380 B.n160 10.6151
R1008 B.n390 B.n160 10.6151
R1009 B.n391 B.n390 10.6151
R1010 B.n392 B.n391 10.6151
R1011 B.n392 B.n152 10.6151
R1012 B.n403 B.n152 10.6151
R1013 B.n404 B.n403 10.6151
R1014 B.n405 B.n404 10.6151
R1015 B.n405 B.n0 10.6151
R1016 B.n531 B.n1 10.6151
R1017 B.n531 B.n530 10.6151
R1018 B.n530 B.n529 10.6151
R1019 B.n529 B.n10 10.6151
R1020 B.n523 B.n10 10.6151
R1021 B.n523 B.n522 10.6151
R1022 B.n522 B.n521 10.6151
R1023 B.n521 B.n17 10.6151
R1024 B.n515 B.n17 10.6151
R1025 B.n515 B.n514 10.6151
R1026 B.n514 B.n513 10.6151
R1027 B.n513 B.n23 10.6151
R1028 B.n507 B.n23 10.6151
R1029 B.n507 B.n506 10.6151
R1030 B.n506 B.n505 10.6151
R1031 B.n505 B.n31 10.6151
R1032 B.n499 B.n31 10.6151
R1033 B.n499 B.n498 10.6151
R1034 B.n498 B.n497 10.6151
R1035 B.n497 B.n38 10.6151
R1036 B.n491 B.n38 10.6151
R1037 B.n491 B.n490 10.6151
R1038 B.n490 B.n489 10.6151
R1039 B.n489 B.n45 10.6151
R1040 B.n483 B.n45 10.6151
R1041 B.n483 B.n482 10.6151
R1042 B.n482 B.n481 10.6151
R1043 B.n481 B.n52 10.6151
R1044 B.n475 B.n52 10.6151
R1045 B.n475 B.n474 10.6151
R1046 B.n474 B.n473 10.6151
R1047 B.n473 B.n59 10.6151
R1048 B.n467 B.n59 10.6151
R1049 B.n467 B.n466 10.6151
R1050 B.n466 B.n465 10.6151
R1051 B.n465 B.n66 10.6151
R1052 B.n109 B.n90 9.36635
R1053 B.n132 B.n87 9.36635
R1054 B.n278 B.n277 9.36635
R1055 B.n256 B.n255 9.36635
R1056 B.n537 B.n0 2.81026
R1057 B.n537 B.n1 2.81026
R1058 B.t7 B.n205 1.65339
R1059 B.n345 B.t2 1.65339
R1060 B.t5 B.n493 1.65339
R1061 B.t14 B.n57 1.65339
R1062 B.n112 B.n90 1.24928
R1063 B.n129 B.n87 1.24928
R1064 B.n277 B.n276 1.24928
R1065 B.n257 B.n256 1.24928
R1066 VP.n28 VP.n27 175.071
R1067 VP.n50 VP.n49 175.071
R1068 VP.n26 VP.n25 175.071
R1069 VP.n13 VP.n12 161.3
R1070 VP.n14 VP.n9 161.3
R1071 VP.n16 VP.n15 161.3
R1072 VP.n17 VP.n8 161.3
R1073 VP.n20 VP.n19 161.3
R1074 VP.n21 VP.n7 161.3
R1075 VP.n23 VP.n22 161.3
R1076 VP.n24 VP.n6 161.3
R1077 VP.n48 VP.n0 161.3
R1078 VP.n47 VP.n46 161.3
R1079 VP.n45 VP.n1 161.3
R1080 VP.n44 VP.n43 161.3
R1081 VP.n41 VP.n2 161.3
R1082 VP.n40 VP.n39 161.3
R1083 VP.n38 VP.n3 161.3
R1084 VP.n37 VP.n36 161.3
R1085 VP.n34 VP.n4 161.3
R1086 VP.n33 VP.n32 161.3
R1087 VP.n31 VP.n5 161.3
R1088 VP.n30 VP.n29 161.3
R1089 VP.n40 VP.n3 56.5617
R1090 VP.n16 VP.n9 56.5617
R1091 VP.n33 VP.n5 56.5617
R1092 VP.n47 VP.n1 56.5617
R1093 VP.n23 VP.n7 56.5617
R1094 VP.n11 VP.n10 54.8557
R1095 VP.n10 VP.t5 54.3696
R1096 VP.n27 VP.n26 38.3793
R1097 VP.n29 VP.n5 24.5923
R1098 VP.n34 VP.n33 24.5923
R1099 VP.n36 VP.n3 24.5923
R1100 VP.n41 VP.n40 24.5923
R1101 VP.n43 VP.n1 24.5923
R1102 VP.n48 VP.n47 24.5923
R1103 VP.n24 VP.n23 24.5923
R1104 VP.n17 VP.n16 24.5923
R1105 VP.n19 VP.n7 24.5923
R1106 VP.n12 VP.n9 24.5923
R1107 VP.n28 VP.t3 20.1569
R1108 VP.n35 VP.t2 20.1569
R1109 VP.n42 VP.t1 20.1569
R1110 VP.n49 VP.t4 20.1569
R1111 VP.n25 VP.t0 20.1569
R1112 VP.n18 VP.t6 20.1569
R1113 VP.n11 VP.t7 20.1569
R1114 VP.n13 VP.n10 17.6839
R1115 VP.n35 VP.n34 12.7883
R1116 VP.n43 VP.n42 12.7883
R1117 VP.n19 VP.n18 12.7883
R1118 VP.n36 VP.n35 11.8046
R1119 VP.n42 VP.n41 11.8046
R1120 VP.n18 VP.n17 11.8046
R1121 VP.n12 VP.n11 11.8046
R1122 VP.n29 VP.n28 10.8209
R1123 VP.n49 VP.n48 10.8209
R1124 VP.n25 VP.n24 10.8209
R1125 VP.n14 VP.n13 0.189894
R1126 VP.n15 VP.n14 0.189894
R1127 VP.n15 VP.n8 0.189894
R1128 VP.n20 VP.n8 0.189894
R1129 VP.n21 VP.n20 0.189894
R1130 VP.n22 VP.n21 0.189894
R1131 VP.n22 VP.n6 0.189894
R1132 VP.n26 VP.n6 0.189894
R1133 VP.n30 VP.n27 0.189894
R1134 VP.n31 VP.n30 0.189894
R1135 VP.n32 VP.n31 0.189894
R1136 VP.n32 VP.n4 0.189894
R1137 VP.n37 VP.n4 0.189894
R1138 VP.n38 VP.n37 0.189894
R1139 VP.n39 VP.n38 0.189894
R1140 VP.n39 VP.n2 0.189894
R1141 VP.n44 VP.n2 0.189894
R1142 VP.n45 VP.n44 0.189894
R1143 VP.n46 VP.n45 0.189894
R1144 VP.n46 VP.n0 0.189894
R1145 VP.n50 VP.n0 0.189894
R1146 VP VP.n50 0.0516364
R1147 VDD1 VDD1.n0 116.148
R1148 VDD1.n3 VDD1.n2 116.034
R1149 VDD1.n3 VDD1.n1 116.034
R1150 VDD1.n5 VDD1.n4 115.237
R1151 VDD1.n5 VDD1.n3 33.169
R1152 VDD1.n4 VDD1.t1 14.3483
R1153 VDD1.n4 VDD1.t7 14.3483
R1154 VDD1.n0 VDD1.t2 14.3483
R1155 VDD1.n0 VDD1.t0 14.3483
R1156 VDD1.n2 VDD1.t6 14.3483
R1157 VDD1.n2 VDD1.t3 14.3483
R1158 VDD1.n1 VDD1.t4 14.3483
R1159 VDD1.n1 VDD1.t5 14.3483
R1160 VDD1 VDD1.n5 0.795759
C0 VDD2 VP 0.42684f
C1 VTAIL VN 2.03813f
C2 VP VTAIL 2.05224f
C3 VDD2 VTAIL 3.71754f
C4 VN VDD1 0.156983f
C5 VP VDD1 1.54011f
C6 VDD2 VDD1 1.28375f
C7 VTAIL VDD1 3.66949f
C8 VP VN 4.53487f
C9 VDD2 VN 1.27269f
C10 VDD2 B 3.425892f
C11 VDD1 B 3.748519f
C12 VTAIL B 3.186319f
C13 VN B 10.679581f
C14 VP B 9.393478f
C15 VDD1.t2 B 0.019338f
C16 VDD1.t0 B 0.019338f
C17 VDD1.n0 B 0.115551f
C18 VDD1.t4 B 0.019338f
C19 VDD1.t5 B 0.019338f
C20 VDD1.n1 B 0.115246f
C21 VDD1.t6 B 0.019338f
C22 VDD1.t3 B 0.019338f
C23 VDD1.n2 B 0.115246f
C24 VDD1.n3 B 1.46416f
C25 VDD1.t1 B 0.019338f
C26 VDD1.t7 B 0.019338f
C27 VDD1.n4 B 0.113412f
C28 VDD1.n5 B 1.2538f
C29 VP.n0 B 0.032113f
C30 VP.t4 B 0.155425f
C31 VP.n1 B 0.044905f
C32 VP.n2 B 0.032113f
C33 VP.t1 B 0.155425f
C34 VP.n3 B 0.046682f
C35 VP.n4 B 0.032113f
C36 VP.t2 B 0.155425f
C37 VP.n5 B 0.048459f
C38 VP.n6 B 0.032113f
C39 VP.t0 B 0.155425f
C40 VP.n7 B 0.044905f
C41 VP.n8 B 0.032113f
C42 VP.t6 B 0.155425f
C43 VP.n9 B 0.046682f
C44 VP.t5 B 0.301822f
C45 VP.n10 B 0.14872f
C46 VP.t7 B 0.155425f
C47 VP.n11 B 0.160681f
C48 VP.n12 B 0.044264f
C49 VP.n13 B 0.207175f
C50 VP.n14 B 0.032113f
C51 VP.n15 B 0.032113f
C52 VP.n16 B 0.046682f
C53 VP.n17 B 0.044264f
C54 VP.n18 B 0.097707f
C55 VP.n19 B 0.04544f
C56 VP.n20 B 0.032113f
C57 VP.n21 B 0.032113f
C58 VP.n22 B 0.032113f
C59 VP.n23 B 0.048459f
C60 VP.n24 B 0.043088f
C61 VP.n25 B 0.172618f
C62 VP.n26 B 1.14134f
C63 VP.n27 B 1.17151f
C64 VP.t3 B 0.155425f
C65 VP.n28 B 0.172618f
C66 VP.n29 B 0.043088f
C67 VP.n30 B 0.032113f
C68 VP.n31 B 0.032113f
C69 VP.n32 B 0.032113f
C70 VP.n33 B 0.044905f
C71 VP.n34 B 0.04544f
C72 VP.n35 B 0.097707f
C73 VP.n36 B 0.044264f
C74 VP.n37 B 0.032113f
C75 VP.n38 B 0.032113f
C76 VP.n39 B 0.032113f
C77 VP.n40 B 0.046682f
C78 VP.n41 B 0.044264f
C79 VP.n42 B 0.097707f
C80 VP.n43 B 0.04544f
C81 VP.n44 B 0.032113f
C82 VP.n45 B 0.032113f
C83 VP.n46 B 0.032113f
C84 VP.n47 B 0.048459f
C85 VP.n48 B 0.043088f
C86 VP.n49 B 0.172618f
C87 VP.n50 B 0.031282f
C88 VTAIL.t8 B 0.03513f
C89 VTAIL.t6 B 0.03513f
C90 VTAIL.n0 B 0.17149f
C91 VTAIL.n1 B 0.384186f
C92 VTAIL.t12 B 0.237796f
C93 VTAIL.n2 B 0.456419f
C94 VTAIL.t14 B 0.237796f
C95 VTAIL.n3 B 0.456419f
C96 VTAIL.t3 B 0.03513f
C97 VTAIL.t4 B 0.03513f
C98 VTAIL.n4 B 0.17149f
C99 VTAIL.n5 B 0.555325f
C100 VTAIL.t2 B 0.237796f
C101 VTAIL.n6 B 1.14591f
C102 VTAIL.t13 B 0.237797f
C103 VTAIL.n7 B 1.14591f
C104 VTAIL.t7 B 0.03513f
C105 VTAIL.t9 B 0.03513f
C106 VTAIL.n8 B 0.17149f
C107 VTAIL.n9 B 0.555325f
C108 VTAIL.t11 B 0.237797f
C109 VTAIL.n10 B 0.456418f
C110 VTAIL.t15 B 0.237797f
C111 VTAIL.n11 B 0.456418f
C112 VTAIL.t0 B 0.03513f
C113 VTAIL.t1 B 0.03513f
C114 VTAIL.n12 B 0.17149f
C115 VTAIL.n13 B 0.555325f
C116 VTAIL.t5 B 0.237796f
C117 VTAIL.n14 B 1.14591f
C118 VTAIL.t10 B 0.237796f
C119 VTAIL.n15 B 1.13987f
C120 VDD2.t4 B 0.019687f
C121 VDD2.t7 B 0.019687f
C122 VDD2.n0 B 0.117322f
C123 VDD2.t6 B 0.019687f
C124 VDD2.t2 B 0.019687f
C125 VDD2.n1 B 0.117322f
C126 VDD2.n2 B 1.45237f
C127 VDD2.t1 B 0.019687f
C128 VDD2.t0 B 0.019687f
C129 VDD2.n3 B 0.115456f
C130 VDD2.n4 B 1.25466f
C131 VDD2.t3 B 0.019687f
C132 VDD2.t5 B 0.019687f
C133 VDD2.n5 B 0.117311f
C134 VN.n0 B 0.031412f
C135 VN.t3 B 0.15203f
C136 VN.n1 B 0.043924f
C137 VN.n2 B 0.031412f
C138 VN.t7 B 0.15203f
C139 VN.n3 B 0.045662f
C140 VN.t1 B 0.295229f
C141 VN.n4 B 0.145472f
C142 VN.t5 B 0.15203f
C143 VN.n5 B 0.157171f
C144 VN.n6 B 0.043297f
C145 VN.n7 B 0.20265f
C146 VN.n8 B 0.031412f
C147 VN.n9 B 0.031412f
C148 VN.n10 B 0.045662f
C149 VN.n11 B 0.043297f
C150 VN.n12 B 0.095573f
C151 VN.n13 B 0.044447f
C152 VN.n14 B 0.031412f
C153 VN.n15 B 0.031412f
C154 VN.n16 B 0.031412f
C155 VN.n17 B 0.0474f
C156 VN.n18 B 0.042147f
C157 VN.n19 B 0.168847f
C158 VN.n20 B 0.030599f
C159 VN.n21 B 0.031412f
C160 VN.t0 B 0.15203f
C161 VN.n22 B 0.043924f
C162 VN.n23 B 0.031412f
C163 VN.t6 B 0.15203f
C164 VN.n24 B 0.045662f
C165 VN.t2 B 0.295229f
C166 VN.n25 B 0.145472f
C167 VN.t4 B 0.15203f
C168 VN.n26 B 0.157171f
C169 VN.n27 B 0.043297f
C170 VN.n28 B 0.20265f
C171 VN.n29 B 0.031412f
C172 VN.n30 B 0.031412f
C173 VN.n31 B 0.045662f
C174 VN.n32 B 0.043297f
C175 VN.n33 B 0.095573f
C176 VN.n34 B 0.044447f
C177 VN.n35 B 0.031412f
C178 VN.n36 B 0.031412f
C179 VN.n37 B 0.031412f
C180 VN.n38 B 0.0474f
C181 VN.n39 B 0.042147f
C182 VN.n40 B 0.168847f
C183 VN.n41 B 1.13716f
.ends

