* NGSPICE file created from diff_pair_sample_0531.ext - technology: sky130A

.subckt diff_pair_sample_0531 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t4 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.1782 pd=1.41 as=0.4212 ps=2.94 w=1.08 l=3.3
X1 VDD1.t3 VP.t0 VTAIL.t2 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.1782 pd=1.41 as=0.4212 ps=2.94 w=1.08 l=3.3
X2 B.t11 B.t9 B.t10 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.4212 pd=2.94 as=0 ps=0 w=1.08 l=3.3
X3 B.t8 B.t6 B.t7 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.4212 pd=2.94 as=0 ps=0 w=1.08 l=3.3
X4 VTAIL.t1 VP.t1 VDD1.t2 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.4212 pd=2.94 as=0.1782 ps=1.41 w=1.08 l=3.3
X5 VTAIL.t3 VP.t2 VDD1.t1 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.4212 pd=2.94 as=0.1782 ps=1.41 w=1.08 l=3.3
X6 B.t5 B.t3 B.t4 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.4212 pd=2.94 as=0 ps=0 w=1.08 l=3.3
X7 VDD2.t2 VN.t1 VTAIL.t6 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.1782 pd=1.41 as=0.4212 ps=2.94 w=1.08 l=3.3
X8 VDD1.t0 VP.t3 VTAIL.t0 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.1782 pd=1.41 as=0.4212 ps=2.94 w=1.08 l=3.3
X9 VTAIL.t5 VN.t2 VDD2.t1 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.4212 pd=2.94 as=0.1782 ps=1.41 w=1.08 l=3.3
X10 B.t2 B.t0 B.t1 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.4212 pd=2.94 as=0 ps=0 w=1.08 l=3.3
X11 VTAIL.t7 VN.t3 VDD2.t0 w_n3148_n1184# sky130_fd_pr__pfet_01v8 ad=0.4212 pd=2.94 as=0.1782 ps=1.41 w=1.08 l=3.3
R0 VN.n1 VN.t1 42.9001
R1 VN.n0 VN.t2 42.9001
R2 VN VN.n1 42.8981
R3 VN.n0 VN.t0 41.78
R4 VN.n1 VN.t3 41.78
R5 VN VN.n0 2.4776
R6 VTAIL.n7 VTAIL.t4 372.135
R7 VTAIL.n0 VTAIL.t5 372.135
R8 VTAIL.n1 VTAIL.t2 372.135
R9 VTAIL.n2 VTAIL.t3 372.135
R10 VTAIL.n6 VTAIL.t0 372.135
R11 VTAIL.n5 VTAIL.t1 372.135
R12 VTAIL.n4 VTAIL.t6 372.135
R13 VTAIL.n3 VTAIL.t7 372.135
R14 VTAIL.n7 VTAIL.n6 16.4272
R15 VTAIL.n3 VTAIL.n2 16.4272
R16 VTAIL.n4 VTAIL.n3 3.12981
R17 VTAIL.n6 VTAIL.n5 3.12981
R18 VTAIL.n2 VTAIL.n1 3.12981
R19 VTAIL VTAIL.n0 1.62334
R20 VTAIL VTAIL.n7 1.50697
R21 VTAIL.n5 VTAIL.n4 0.470328
R22 VTAIL.n1 VTAIL.n0 0.470328
R23 VDD2.n2 VDD2.n0 379.909
R24 VDD2.n2 VDD2.n1 345.875
R25 VDD2.n1 VDD2.t0 30.0977
R26 VDD2.n1 VDD2.t2 30.0977
R27 VDD2.n0 VDD2.t1 30.0977
R28 VDD2.n0 VDD2.t3 30.0977
R29 VDD2 VDD2.n2 0.0586897
R30 VP.n17 VP.n16 161.3
R31 VP.n15 VP.n1 161.3
R32 VP.n14 VP.n13 161.3
R33 VP.n12 VP.n2 161.3
R34 VP.n11 VP.n10 161.3
R35 VP.n9 VP.n3 161.3
R36 VP.n8 VP.n7 161.3
R37 VP.n6 VP.n4 74.7527
R38 VP.n18 VP.n0 74.7527
R39 VP.n5 VP.t1 42.8999
R40 VP.n6 VP.n5 42.7328
R41 VP.n5 VP.t3 41.78
R42 VP.n10 VP.n2 40.577
R43 VP.n14 VP.n2 40.577
R44 VP.n9 VP.n8 24.5923
R45 VP.n10 VP.n9 24.5923
R46 VP.n15 VP.n14 24.5923
R47 VP.n16 VP.n15 24.5923
R48 VP.n8 VP.n4 15.4934
R49 VP.n16 VP.n0 15.4934
R50 VP.n4 VP.t2 7.88777
R51 VP.n0 VP.t0 7.88777
R52 VP.n7 VP.n6 0.354861
R53 VP.n18 VP.n17 0.354861
R54 VP VP.n18 0.267071
R55 VP.n7 VP.n3 0.189894
R56 VP.n11 VP.n3 0.189894
R57 VP.n12 VP.n11 0.189894
R58 VP.n13 VP.n12 0.189894
R59 VP.n13 VP.n1 0.189894
R60 VP.n17 VP.n1 0.189894
R61 VDD1 VDD1.n1 380.435
R62 VDD1 VDD1.n0 345.935
R63 VDD1.n0 VDD1.t2 30.0977
R64 VDD1.n0 VDD1.t0 30.0977
R65 VDD1.n1 VDD1.t1 30.0977
R66 VDD1.n1 VDD1.t3 30.0977
R67 B.n345 B.n40 585
R68 B.n347 B.n346 585
R69 B.n348 B.n39 585
R70 B.n350 B.n349 585
R71 B.n351 B.n38 585
R72 B.n353 B.n352 585
R73 B.n354 B.n37 585
R74 B.n356 B.n355 585
R75 B.n357 B.n36 585
R76 B.n359 B.n358 585
R77 B.n361 B.n33 585
R78 B.n363 B.n362 585
R79 B.n364 B.n32 585
R80 B.n366 B.n365 585
R81 B.n367 B.n31 585
R82 B.n369 B.n368 585
R83 B.n370 B.n30 585
R84 B.n372 B.n371 585
R85 B.n373 B.n27 585
R86 B.n376 B.n375 585
R87 B.n377 B.n26 585
R88 B.n379 B.n378 585
R89 B.n380 B.n25 585
R90 B.n382 B.n381 585
R91 B.n383 B.n24 585
R92 B.n385 B.n384 585
R93 B.n386 B.n23 585
R94 B.n388 B.n387 585
R95 B.n389 B.n22 585
R96 B.n344 B.n343 585
R97 B.n342 B.n41 585
R98 B.n341 B.n340 585
R99 B.n339 B.n42 585
R100 B.n338 B.n337 585
R101 B.n336 B.n43 585
R102 B.n335 B.n334 585
R103 B.n333 B.n44 585
R104 B.n332 B.n331 585
R105 B.n330 B.n45 585
R106 B.n329 B.n328 585
R107 B.n327 B.n46 585
R108 B.n326 B.n325 585
R109 B.n324 B.n47 585
R110 B.n323 B.n322 585
R111 B.n321 B.n48 585
R112 B.n320 B.n319 585
R113 B.n318 B.n49 585
R114 B.n317 B.n316 585
R115 B.n315 B.n50 585
R116 B.n314 B.n313 585
R117 B.n312 B.n51 585
R118 B.n311 B.n310 585
R119 B.n309 B.n52 585
R120 B.n308 B.n307 585
R121 B.n306 B.n53 585
R122 B.n305 B.n304 585
R123 B.n303 B.n54 585
R124 B.n302 B.n301 585
R125 B.n300 B.n55 585
R126 B.n299 B.n298 585
R127 B.n297 B.n56 585
R128 B.n296 B.n295 585
R129 B.n294 B.n57 585
R130 B.n293 B.n292 585
R131 B.n291 B.n58 585
R132 B.n290 B.n289 585
R133 B.n288 B.n59 585
R134 B.n287 B.n286 585
R135 B.n285 B.n60 585
R136 B.n284 B.n283 585
R137 B.n282 B.n61 585
R138 B.n281 B.n280 585
R139 B.n279 B.n62 585
R140 B.n278 B.n277 585
R141 B.n276 B.n63 585
R142 B.n275 B.n274 585
R143 B.n273 B.n64 585
R144 B.n272 B.n271 585
R145 B.n270 B.n65 585
R146 B.n269 B.n268 585
R147 B.n267 B.n66 585
R148 B.n266 B.n265 585
R149 B.n264 B.n67 585
R150 B.n263 B.n262 585
R151 B.n261 B.n68 585
R152 B.n260 B.n259 585
R153 B.n258 B.n69 585
R154 B.n257 B.n256 585
R155 B.n255 B.n70 585
R156 B.n254 B.n253 585
R157 B.n252 B.n71 585
R158 B.n251 B.n250 585
R159 B.n249 B.n72 585
R160 B.n248 B.n247 585
R161 B.n246 B.n73 585
R162 B.n245 B.n244 585
R163 B.n243 B.n74 585
R164 B.n242 B.n241 585
R165 B.n240 B.n75 585
R166 B.n239 B.n238 585
R167 B.n237 B.n76 585
R168 B.n236 B.n235 585
R169 B.n234 B.n77 585
R170 B.n233 B.n232 585
R171 B.n231 B.n78 585
R172 B.n230 B.n229 585
R173 B.n228 B.n79 585
R174 B.n227 B.n226 585
R175 B.n225 B.n80 585
R176 B.n224 B.n223 585
R177 B.n179 B.n178 585
R178 B.n180 B.n99 585
R179 B.n182 B.n181 585
R180 B.n183 B.n98 585
R181 B.n185 B.n184 585
R182 B.n186 B.n97 585
R183 B.n188 B.n187 585
R184 B.n189 B.n96 585
R185 B.n191 B.n190 585
R186 B.n192 B.n93 585
R187 B.n195 B.n194 585
R188 B.n196 B.n92 585
R189 B.n198 B.n197 585
R190 B.n199 B.n91 585
R191 B.n201 B.n200 585
R192 B.n202 B.n90 585
R193 B.n204 B.n203 585
R194 B.n205 B.n89 585
R195 B.n207 B.n206 585
R196 B.n209 B.n208 585
R197 B.n210 B.n85 585
R198 B.n212 B.n211 585
R199 B.n213 B.n84 585
R200 B.n215 B.n214 585
R201 B.n216 B.n83 585
R202 B.n218 B.n217 585
R203 B.n219 B.n82 585
R204 B.n221 B.n220 585
R205 B.n222 B.n81 585
R206 B.n177 B.n100 585
R207 B.n176 B.n175 585
R208 B.n174 B.n101 585
R209 B.n173 B.n172 585
R210 B.n171 B.n102 585
R211 B.n170 B.n169 585
R212 B.n168 B.n103 585
R213 B.n167 B.n166 585
R214 B.n165 B.n104 585
R215 B.n164 B.n163 585
R216 B.n162 B.n105 585
R217 B.n161 B.n160 585
R218 B.n159 B.n106 585
R219 B.n158 B.n157 585
R220 B.n156 B.n107 585
R221 B.n155 B.n154 585
R222 B.n153 B.n108 585
R223 B.n152 B.n151 585
R224 B.n150 B.n109 585
R225 B.n149 B.n148 585
R226 B.n147 B.n110 585
R227 B.n146 B.n145 585
R228 B.n144 B.n111 585
R229 B.n143 B.n142 585
R230 B.n141 B.n112 585
R231 B.n140 B.n139 585
R232 B.n138 B.n113 585
R233 B.n137 B.n136 585
R234 B.n135 B.n114 585
R235 B.n134 B.n133 585
R236 B.n132 B.n115 585
R237 B.n131 B.n130 585
R238 B.n129 B.n116 585
R239 B.n128 B.n127 585
R240 B.n126 B.n117 585
R241 B.n125 B.n124 585
R242 B.n123 B.n118 585
R243 B.n122 B.n121 585
R244 B.n120 B.n119 585
R245 B.n2 B.n0 585
R246 B.n449 B.n1 585
R247 B.n448 B.n447 585
R248 B.n446 B.n3 585
R249 B.n445 B.n444 585
R250 B.n443 B.n4 585
R251 B.n442 B.n441 585
R252 B.n440 B.n5 585
R253 B.n439 B.n438 585
R254 B.n437 B.n6 585
R255 B.n436 B.n435 585
R256 B.n434 B.n7 585
R257 B.n433 B.n432 585
R258 B.n431 B.n8 585
R259 B.n430 B.n429 585
R260 B.n428 B.n9 585
R261 B.n427 B.n426 585
R262 B.n425 B.n10 585
R263 B.n424 B.n423 585
R264 B.n422 B.n11 585
R265 B.n421 B.n420 585
R266 B.n419 B.n12 585
R267 B.n418 B.n417 585
R268 B.n416 B.n13 585
R269 B.n415 B.n414 585
R270 B.n413 B.n14 585
R271 B.n412 B.n411 585
R272 B.n410 B.n15 585
R273 B.n409 B.n408 585
R274 B.n407 B.n16 585
R275 B.n406 B.n405 585
R276 B.n404 B.n17 585
R277 B.n403 B.n402 585
R278 B.n401 B.n18 585
R279 B.n400 B.n399 585
R280 B.n398 B.n19 585
R281 B.n397 B.n396 585
R282 B.n395 B.n20 585
R283 B.n394 B.n393 585
R284 B.n392 B.n21 585
R285 B.n391 B.n390 585
R286 B.n451 B.n450 585
R287 B.n178 B.n177 487.695
R288 B.n390 B.n389 487.695
R289 B.n224 B.n81 487.695
R290 B.n345 B.n344 487.695
R291 B.n86 B.t2 433.151
R292 B.n94 B.t11 433.151
R293 B.n28 B.t4 433.151
R294 B.n34 B.t7 433.151
R295 B.n87 B.t1 362.75
R296 B.n95 B.t10 362.75
R297 B.n29 B.t5 362.75
R298 B.n35 B.t8 362.75
R299 B.n86 B.t0 209.588
R300 B.n94 B.t9 209.588
R301 B.n28 B.t3 209.588
R302 B.n34 B.t6 209.588
R303 B.n177 B.n176 163.367
R304 B.n176 B.n101 163.367
R305 B.n172 B.n101 163.367
R306 B.n172 B.n171 163.367
R307 B.n171 B.n170 163.367
R308 B.n170 B.n103 163.367
R309 B.n166 B.n103 163.367
R310 B.n166 B.n165 163.367
R311 B.n165 B.n164 163.367
R312 B.n164 B.n105 163.367
R313 B.n160 B.n105 163.367
R314 B.n160 B.n159 163.367
R315 B.n159 B.n158 163.367
R316 B.n158 B.n107 163.367
R317 B.n154 B.n107 163.367
R318 B.n154 B.n153 163.367
R319 B.n153 B.n152 163.367
R320 B.n152 B.n109 163.367
R321 B.n148 B.n109 163.367
R322 B.n148 B.n147 163.367
R323 B.n147 B.n146 163.367
R324 B.n146 B.n111 163.367
R325 B.n142 B.n111 163.367
R326 B.n142 B.n141 163.367
R327 B.n141 B.n140 163.367
R328 B.n140 B.n113 163.367
R329 B.n136 B.n113 163.367
R330 B.n136 B.n135 163.367
R331 B.n135 B.n134 163.367
R332 B.n134 B.n115 163.367
R333 B.n130 B.n115 163.367
R334 B.n130 B.n129 163.367
R335 B.n129 B.n128 163.367
R336 B.n128 B.n117 163.367
R337 B.n124 B.n117 163.367
R338 B.n124 B.n123 163.367
R339 B.n123 B.n122 163.367
R340 B.n122 B.n119 163.367
R341 B.n119 B.n2 163.367
R342 B.n450 B.n2 163.367
R343 B.n450 B.n449 163.367
R344 B.n449 B.n448 163.367
R345 B.n448 B.n3 163.367
R346 B.n444 B.n3 163.367
R347 B.n444 B.n443 163.367
R348 B.n443 B.n442 163.367
R349 B.n442 B.n5 163.367
R350 B.n438 B.n5 163.367
R351 B.n438 B.n437 163.367
R352 B.n437 B.n436 163.367
R353 B.n436 B.n7 163.367
R354 B.n432 B.n7 163.367
R355 B.n432 B.n431 163.367
R356 B.n431 B.n430 163.367
R357 B.n430 B.n9 163.367
R358 B.n426 B.n9 163.367
R359 B.n426 B.n425 163.367
R360 B.n425 B.n424 163.367
R361 B.n424 B.n11 163.367
R362 B.n420 B.n11 163.367
R363 B.n420 B.n419 163.367
R364 B.n419 B.n418 163.367
R365 B.n418 B.n13 163.367
R366 B.n414 B.n13 163.367
R367 B.n414 B.n413 163.367
R368 B.n413 B.n412 163.367
R369 B.n412 B.n15 163.367
R370 B.n408 B.n15 163.367
R371 B.n408 B.n407 163.367
R372 B.n407 B.n406 163.367
R373 B.n406 B.n17 163.367
R374 B.n402 B.n17 163.367
R375 B.n402 B.n401 163.367
R376 B.n401 B.n400 163.367
R377 B.n400 B.n19 163.367
R378 B.n396 B.n19 163.367
R379 B.n396 B.n395 163.367
R380 B.n395 B.n394 163.367
R381 B.n394 B.n21 163.367
R382 B.n390 B.n21 163.367
R383 B.n178 B.n99 163.367
R384 B.n182 B.n99 163.367
R385 B.n183 B.n182 163.367
R386 B.n184 B.n183 163.367
R387 B.n184 B.n97 163.367
R388 B.n188 B.n97 163.367
R389 B.n189 B.n188 163.367
R390 B.n190 B.n189 163.367
R391 B.n190 B.n93 163.367
R392 B.n195 B.n93 163.367
R393 B.n196 B.n195 163.367
R394 B.n197 B.n196 163.367
R395 B.n197 B.n91 163.367
R396 B.n201 B.n91 163.367
R397 B.n202 B.n201 163.367
R398 B.n203 B.n202 163.367
R399 B.n203 B.n89 163.367
R400 B.n207 B.n89 163.367
R401 B.n208 B.n207 163.367
R402 B.n208 B.n85 163.367
R403 B.n212 B.n85 163.367
R404 B.n213 B.n212 163.367
R405 B.n214 B.n213 163.367
R406 B.n214 B.n83 163.367
R407 B.n218 B.n83 163.367
R408 B.n219 B.n218 163.367
R409 B.n220 B.n219 163.367
R410 B.n220 B.n81 163.367
R411 B.n225 B.n224 163.367
R412 B.n226 B.n225 163.367
R413 B.n226 B.n79 163.367
R414 B.n230 B.n79 163.367
R415 B.n231 B.n230 163.367
R416 B.n232 B.n231 163.367
R417 B.n232 B.n77 163.367
R418 B.n236 B.n77 163.367
R419 B.n237 B.n236 163.367
R420 B.n238 B.n237 163.367
R421 B.n238 B.n75 163.367
R422 B.n242 B.n75 163.367
R423 B.n243 B.n242 163.367
R424 B.n244 B.n243 163.367
R425 B.n244 B.n73 163.367
R426 B.n248 B.n73 163.367
R427 B.n249 B.n248 163.367
R428 B.n250 B.n249 163.367
R429 B.n250 B.n71 163.367
R430 B.n254 B.n71 163.367
R431 B.n255 B.n254 163.367
R432 B.n256 B.n255 163.367
R433 B.n256 B.n69 163.367
R434 B.n260 B.n69 163.367
R435 B.n261 B.n260 163.367
R436 B.n262 B.n261 163.367
R437 B.n262 B.n67 163.367
R438 B.n266 B.n67 163.367
R439 B.n267 B.n266 163.367
R440 B.n268 B.n267 163.367
R441 B.n268 B.n65 163.367
R442 B.n272 B.n65 163.367
R443 B.n273 B.n272 163.367
R444 B.n274 B.n273 163.367
R445 B.n274 B.n63 163.367
R446 B.n278 B.n63 163.367
R447 B.n279 B.n278 163.367
R448 B.n280 B.n279 163.367
R449 B.n280 B.n61 163.367
R450 B.n284 B.n61 163.367
R451 B.n285 B.n284 163.367
R452 B.n286 B.n285 163.367
R453 B.n286 B.n59 163.367
R454 B.n290 B.n59 163.367
R455 B.n291 B.n290 163.367
R456 B.n292 B.n291 163.367
R457 B.n292 B.n57 163.367
R458 B.n296 B.n57 163.367
R459 B.n297 B.n296 163.367
R460 B.n298 B.n297 163.367
R461 B.n298 B.n55 163.367
R462 B.n302 B.n55 163.367
R463 B.n303 B.n302 163.367
R464 B.n304 B.n303 163.367
R465 B.n304 B.n53 163.367
R466 B.n308 B.n53 163.367
R467 B.n309 B.n308 163.367
R468 B.n310 B.n309 163.367
R469 B.n310 B.n51 163.367
R470 B.n314 B.n51 163.367
R471 B.n315 B.n314 163.367
R472 B.n316 B.n315 163.367
R473 B.n316 B.n49 163.367
R474 B.n320 B.n49 163.367
R475 B.n321 B.n320 163.367
R476 B.n322 B.n321 163.367
R477 B.n322 B.n47 163.367
R478 B.n326 B.n47 163.367
R479 B.n327 B.n326 163.367
R480 B.n328 B.n327 163.367
R481 B.n328 B.n45 163.367
R482 B.n332 B.n45 163.367
R483 B.n333 B.n332 163.367
R484 B.n334 B.n333 163.367
R485 B.n334 B.n43 163.367
R486 B.n338 B.n43 163.367
R487 B.n339 B.n338 163.367
R488 B.n340 B.n339 163.367
R489 B.n340 B.n41 163.367
R490 B.n344 B.n41 163.367
R491 B.n389 B.n388 163.367
R492 B.n388 B.n23 163.367
R493 B.n384 B.n23 163.367
R494 B.n384 B.n383 163.367
R495 B.n383 B.n382 163.367
R496 B.n382 B.n25 163.367
R497 B.n378 B.n25 163.367
R498 B.n378 B.n377 163.367
R499 B.n377 B.n376 163.367
R500 B.n376 B.n27 163.367
R501 B.n371 B.n27 163.367
R502 B.n371 B.n370 163.367
R503 B.n370 B.n369 163.367
R504 B.n369 B.n31 163.367
R505 B.n365 B.n31 163.367
R506 B.n365 B.n364 163.367
R507 B.n364 B.n363 163.367
R508 B.n363 B.n33 163.367
R509 B.n358 B.n33 163.367
R510 B.n358 B.n357 163.367
R511 B.n357 B.n356 163.367
R512 B.n356 B.n37 163.367
R513 B.n352 B.n37 163.367
R514 B.n352 B.n351 163.367
R515 B.n351 B.n350 163.367
R516 B.n350 B.n39 163.367
R517 B.n346 B.n39 163.367
R518 B.n346 B.n345 163.367
R519 B.n87 B.n86 70.4005
R520 B.n95 B.n94 70.4005
R521 B.n29 B.n28 70.4005
R522 B.n35 B.n34 70.4005
R523 B.n88 B.n87 59.5399
R524 B.n193 B.n95 59.5399
R525 B.n374 B.n29 59.5399
R526 B.n360 B.n35 59.5399
R527 B.n391 B.n22 31.6883
R528 B.n343 B.n40 31.6883
R529 B.n223 B.n222 31.6883
R530 B.n179 B.n100 31.6883
R531 B B.n451 18.0485
R532 B.n387 B.n22 10.6151
R533 B.n387 B.n386 10.6151
R534 B.n386 B.n385 10.6151
R535 B.n385 B.n24 10.6151
R536 B.n381 B.n24 10.6151
R537 B.n381 B.n380 10.6151
R538 B.n380 B.n379 10.6151
R539 B.n379 B.n26 10.6151
R540 B.n375 B.n26 10.6151
R541 B.n373 B.n372 10.6151
R542 B.n372 B.n30 10.6151
R543 B.n368 B.n30 10.6151
R544 B.n368 B.n367 10.6151
R545 B.n367 B.n366 10.6151
R546 B.n366 B.n32 10.6151
R547 B.n362 B.n32 10.6151
R548 B.n362 B.n361 10.6151
R549 B.n359 B.n36 10.6151
R550 B.n355 B.n36 10.6151
R551 B.n355 B.n354 10.6151
R552 B.n354 B.n353 10.6151
R553 B.n353 B.n38 10.6151
R554 B.n349 B.n38 10.6151
R555 B.n349 B.n348 10.6151
R556 B.n348 B.n347 10.6151
R557 B.n347 B.n40 10.6151
R558 B.n223 B.n80 10.6151
R559 B.n227 B.n80 10.6151
R560 B.n228 B.n227 10.6151
R561 B.n229 B.n228 10.6151
R562 B.n229 B.n78 10.6151
R563 B.n233 B.n78 10.6151
R564 B.n234 B.n233 10.6151
R565 B.n235 B.n234 10.6151
R566 B.n235 B.n76 10.6151
R567 B.n239 B.n76 10.6151
R568 B.n240 B.n239 10.6151
R569 B.n241 B.n240 10.6151
R570 B.n241 B.n74 10.6151
R571 B.n245 B.n74 10.6151
R572 B.n246 B.n245 10.6151
R573 B.n247 B.n246 10.6151
R574 B.n247 B.n72 10.6151
R575 B.n251 B.n72 10.6151
R576 B.n252 B.n251 10.6151
R577 B.n253 B.n252 10.6151
R578 B.n253 B.n70 10.6151
R579 B.n257 B.n70 10.6151
R580 B.n258 B.n257 10.6151
R581 B.n259 B.n258 10.6151
R582 B.n259 B.n68 10.6151
R583 B.n263 B.n68 10.6151
R584 B.n264 B.n263 10.6151
R585 B.n265 B.n264 10.6151
R586 B.n265 B.n66 10.6151
R587 B.n269 B.n66 10.6151
R588 B.n270 B.n269 10.6151
R589 B.n271 B.n270 10.6151
R590 B.n271 B.n64 10.6151
R591 B.n275 B.n64 10.6151
R592 B.n276 B.n275 10.6151
R593 B.n277 B.n276 10.6151
R594 B.n277 B.n62 10.6151
R595 B.n281 B.n62 10.6151
R596 B.n282 B.n281 10.6151
R597 B.n283 B.n282 10.6151
R598 B.n283 B.n60 10.6151
R599 B.n287 B.n60 10.6151
R600 B.n288 B.n287 10.6151
R601 B.n289 B.n288 10.6151
R602 B.n289 B.n58 10.6151
R603 B.n293 B.n58 10.6151
R604 B.n294 B.n293 10.6151
R605 B.n295 B.n294 10.6151
R606 B.n295 B.n56 10.6151
R607 B.n299 B.n56 10.6151
R608 B.n300 B.n299 10.6151
R609 B.n301 B.n300 10.6151
R610 B.n301 B.n54 10.6151
R611 B.n305 B.n54 10.6151
R612 B.n306 B.n305 10.6151
R613 B.n307 B.n306 10.6151
R614 B.n307 B.n52 10.6151
R615 B.n311 B.n52 10.6151
R616 B.n312 B.n311 10.6151
R617 B.n313 B.n312 10.6151
R618 B.n313 B.n50 10.6151
R619 B.n317 B.n50 10.6151
R620 B.n318 B.n317 10.6151
R621 B.n319 B.n318 10.6151
R622 B.n319 B.n48 10.6151
R623 B.n323 B.n48 10.6151
R624 B.n324 B.n323 10.6151
R625 B.n325 B.n324 10.6151
R626 B.n325 B.n46 10.6151
R627 B.n329 B.n46 10.6151
R628 B.n330 B.n329 10.6151
R629 B.n331 B.n330 10.6151
R630 B.n331 B.n44 10.6151
R631 B.n335 B.n44 10.6151
R632 B.n336 B.n335 10.6151
R633 B.n337 B.n336 10.6151
R634 B.n337 B.n42 10.6151
R635 B.n341 B.n42 10.6151
R636 B.n342 B.n341 10.6151
R637 B.n343 B.n342 10.6151
R638 B.n180 B.n179 10.6151
R639 B.n181 B.n180 10.6151
R640 B.n181 B.n98 10.6151
R641 B.n185 B.n98 10.6151
R642 B.n186 B.n185 10.6151
R643 B.n187 B.n186 10.6151
R644 B.n187 B.n96 10.6151
R645 B.n191 B.n96 10.6151
R646 B.n192 B.n191 10.6151
R647 B.n194 B.n92 10.6151
R648 B.n198 B.n92 10.6151
R649 B.n199 B.n198 10.6151
R650 B.n200 B.n199 10.6151
R651 B.n200 B.n90 10.6151
R652 B.n204 B.n90 10.6151
R653 B.n205 B.n204 10.6151
R654 B.n206 B.n205 10.6151
R655 B.n210 B.n209 10.6151
R656 B.n211 B.n210 10.6151
R657 B.n211 B.n84 10.6151
R658 B.n215 B.n84 10.6151
R659 B.n216 B.n215 10.6151
R660 B.n217 B.n216 10.6151
R661 B.n217 B.n82 10.6151
R662 B.n221 B.n82 10.6151
R663 B.n222 B.n221 10.6151
R664 B.n175 B.n100 10.6151
R665 B.n175 B.n174 10.6151
R666 B.n174 B.n173 10.6151
R667 B.n173 B.n102 10.6151
R668 B.n169 B.n102 10.6151
R669 B.n169 B.n168 10.6151
R670 B.n168 B.n167 10.6151
R671 B.n167 B.n104 10.6151
R672 B.n163 B.n104 10.6151
R673 B.n163 B.n162 10.6151
R674 B.n162 B.n161 10.6151
R675 B.n161 B.n106 10.6151
R676 B.n157 B.n106 10.6151
R677 B.n157 B.n156 10.6151
R678 B.n156 B.n155 10.6151
R679 B.n155 B.n108 10.6151
R680 B.n151 B.n108 10.6151
R681 B.n151 B.n150 10.6151
R682 B.n150 B.n149 10.6151
R683 B.n149 B.n110 10.6151
R684 B.n145 B.n110 10.6151
R685 B.n145 B.n144 10.6151
R686 B.n144 B.n143 10.6151
R687 B.n143 B.n112 10.6151
R688 B.n139 B.n112 10.6151
R689 B.n139 B.n138 10.6151
R690 B.n138 B.n137 10.6151
R691 B.n137 B.n114 10.6151
R692 B.n133 B.n114 10.6151
R693 B.n133 B.n132 10.6151
R694 B.n132 B.n131 10.6151
R695 B.n131 B.n116 10.6151
R696 B.n127 B.n116 10.6151
R697 B.n127 B.n126 10.6151
R698 B.n126 B.n125 10.6151
R699 B.n125 B.n118 10.6151
R700 B.n121 B.n118 10.6151
R701 B.n121 B.n120 10.6151
R702 B.n120 B.n0 10.6151
R703 B.n447 B.n1 10.6151
R704 B.n447 B.n446 10.6151
R705 B.n446 B.n445 10.6151
R706 B.n445 B.n4 10.6151
R707 B.n441 B.n4 10.6151
R708 B.n441 B.n440 10.6151
R709 B.n440 B.n439 10.6151
R710 B.n439 B.n6 10.6151
R711 B.n435 B.n6 10.6151
R712 B.n435 B.n434 10.6151
R713 B.n434 B.n433 10.6151
R714 B.n433 B.n8 10.6151
R715 B.n429 B.n8 10.6151
R716 B.n429 B.n428 10.6151
R717 B.n428 B.n427 10.6151
R718 B.n427 B.n10 10.6151
R719 B.n423 B.n10 10.6151
R720 B.n423 B.n422 10.6151
R721 B.n422 B.n421 10.6151
R722 B.n421 B.n12 10.6151
R723 B.n417 B.n12 10.6151
R724 B.n417 B.n416 10.6151
R725 B.n416 B.n415 10.6151
R726 B.n415 B.n14 10.6151
R727 B.n411 B.n14 10.6151
R728 B.n411 B.n410 10.6151
R729 B.n410 B.n409 10.6151
R730 B.n409 B.n16 10.6151
R731 B.n405 B.n16 10.6151
R732 B.n405 B.n404 10.6151
R733 B.n404 B.n403 10.6151
R734 B.n403 B.n18 10.6151
R735 B.n399 B.n18 10.6151
R736 B.n399 B.n398 10.6151
R737 B.n398 B.n397 10.6151
R738 B.n397 B.n20 10.6151
R739 B.n393 B.n20 10.6151
R740 B.n393 B.n392 10.6151
R741 B.n392 B.n391 10.6151
R742 B.n374 B.n373 6.5566
R743 B.n361 B.n360 6.5566
R744 B.n194 B.n193 6.5566
R745 B.n206 B.n88 6.5566
R746 B.n375 B.n374 4.05904
R747 B.n360 B.n359 4.05904
R748 B.n193 B.n192 4.05904
R749 B.n209 B.n88 4.05904
R750 B.n451 B.n0 2.81026
R751 B.n451 B.n1 2.81026
C0 VTAIL w_n3148_n1184# 1.51677f
C1 VDD2 VP 0.447395f
C2 VDD1 VP 1.04347f
C3 VTAIL VP 1.62302f
C4 VN B 1.05186f
C5 VDD2 VN 0.755415f
C6 VDD2 B 1.15542f
C7 VDD1 VN 0.15671f
C8 VDD1 B 1.09095f
C9 w_n3148_n1184# VP 5.64095f
C10 VTAIL VN 1.60891f
C11 VTAIL B 1.33634f
C12 VDD1 VDD2 1.19017f
C13 VTAIL VDD2 3.25319f
C14 VDD1 VTAIL 3.19429f
C15 w_n3148_n1184# VN 5.24197f
C16 w_n3148_n1184# B 7.13268f
C17 VN VP 4.67776f
C18 VP B 1.72842f
C19 VDD2 w_n3148_n1184# 1.35184f
C20 VDD1 w_n3148_n1184# 1.2813f
C21 VDD2 VSUBS 0.780964f
C22 VDD1 VSUBS 3.867977f
C23 VTAIL VSUBS 0.448917f
C24 VN VSUBS 6.05609f
C25 VP VSUBS 2.090166f
C26 B VSUBS 3.728904f
C27 w_n3148_n1184# VSUBS 48.0133f
C28 B.n0 VSUBS 0.006724f
C29 B.n1 VSUBS 0.006724f
C30 B.n2 VSUBS 0.010633f
C31 B.n3 VSUBS 0.010633f
C32 B.n4 VSUBS 0.010633f
C33 B.n5 VSUBS 0.010633f
C34 B.n6 VSUBS 0.010633f
C35 B.n7 VSUBS 0.010633f
C36 B.n8 VSUBS 0.010633f
C37 B.n9 VSUBS 0.010633f
C38 B.n10 VSUBS 0.010633f
C39 B.n11 VSUBS 0.010633f
C40 B.n12 VSUBS 0.010633f
C41 B.n13 VSUBS 0.010633f
C42 B.n14 VSUBS 0.010633f
C43 B.n15 VSUBS 0.010633f
C44 B.n16 VSUBS 0.010633f
C45 B.n17 VSUBS 0.010633f
C46 B.n18 VSUBS 0.010633f
C47 B.n19 VSUBS 0.010633f
C48 B.n20 VSUBS 0.010633f
C49 B.n21 VSUBS 0.010633f
C50 B.n22 VSUBS 0.025389f
C51 B.n23 VSUBS 0.010633f
C52 B.n24 VSUBS 0.010633f
C53 B.n25 VSUBS 0.010633f
C54 B.n26 VSUBS 0.010633f
C55 B.n27 VSUBS 0.010633f
C56 B.t5 VSUBS 0.030871f
C57 B.t4 VSUBS 0.040904f
C58 B.t3 VSUBS 0.27277f
C59 B.n28 VSUBS 0.104778f
C60 B.n29 VSUBS 0.076899f
C61 B.n30 VSUBS 0.010633f
C62 B.n31 VSUBS 0.010633f
C63 B.n32 VSUBS 0.010633f
C64 B.n33 VSUBS 0.010633f
C65 B.t8 VSUBS 0.030871f
C66 B.t7 VSUBS 0.040904f
C67 B.t6 VSUBS 0.27277f
C68 B.n34 VSUBS 0.104778f
C69 B.n35 VSUBS 0.076899f
C70 B.n36 VSUBS 0.010633f
C71 B.n37 VSUBS 0.010633f
C72 B.n38 VSUBS 0.010633f
C73 B.n39 VSUBS 0.010633f
C74 B.n40 VSUBS 0.024094f
C75 B.n41 VSUBS 0.010633f
C76 B.n42 VSUBS 0.010633f
C77 B.n43 VSUBS 0.010633f
C78 B.n44 VSUBS 0.010633f
C79 B.n45 VSUBS 0.010633f
C80 B.n46 VSUBS 0.010633f
C81 B.n47 VSUBS 0.010633f
C82 B.n48 VSUBS 0.010633f
C83 B.n49 VSUBS 0.010633f
C84 B.n50 VSUBS 0.010633f
C85 B.n51 VSUBS 0.010633f
C86 B.n52 VSUBS 0.010633f
C87 B.n53 VSUBS 0.010633f
C88 B.n54 VSUBS 0.010633f
C89 B.n55 VSUBS 0.010633f
C90 B.n56 VSUBS 0.010633f
C91 B.n57 VSUBS 0.010633f
C92 B.n58 VSUBS 0.010633f
C93 B.n59 VSUBS 0.010633f
C94 B.n60 VSUBS 0.010633f
C95 B.n61 VSUBS 0.010633f
C96 B.n62 VSUBS 0.010633f
C97 B.n63 VSUBS 0.010633f
C98 B.n64 VSUBS 0.010633f
C99 B.n65 VSUBS 0.010633f
C100 B.n66 VSUBS 0.010633f
C101 B.n67 VSUBS 0.010633f
C102 B.n68 VSUBS 0.010633f
C103 B.n69 VSUBS 0.010633f
C104 B.n70 VSUBS 0.010633f
C105 B.n71 VSUBS 0.010633f
C106 B.n72 VSUBS 0.010633f
C107 B.n73 VSUBS 0.010633f
C108 B.n74 VSUBS 0.010633f
C109 B.n75 VSUBS 0.010633f
C110 B.n76 VSUBS 0.010633f
C111 B.n77 VSUBS 0.010633f
C112 B.n78 VSUBS 0.010633f
C113 B.n79 VSUBS 0.010633f
C114 B.n80 VSUBS 0.010633f
C115 B.n81 VSUBS 0.025389f
C116 B.n82 VSUBS 0.010633f
C117 B.n83 VSUBS 0.010633f
C118 B.n84 VSUBS 0.010633f
C119 B.n85 VSUBS 0.010633f
C120 B.t1 VSUBS 0.030871f
C121 B.t2 VSUBS 0.040904f
C122 B.t0 VSUBS 0.27277f
C123 B.n86 VSUBS 0.104778f
C124 B.n87 VSUBS 0.076899f
C125 B.n88 VSUBS 0.024636f
C126 B.n89 VSUBS 0.010633f
C127 B.n90 VSUBS 0.010633f
C128 B.n91 VSUBS 0.010633f
C129 B.n92 VSUBS 0.010633f
C130 B.n93 VSUBS 0.010633f
C131 B.t10 VSUBS 0.030871f
C132 B.t11 VSUBS 0.040904f
C133 B.t9 VSUBS 0.27277f
C134 B.n94 VSUBS 0.104778f
C135 B.n95 VSUBS 0.076899f
C136 B.n96 VSUBS 0.010633f
C137 B.n97 VSUBS 0.010633f
C138 B.n98 VSUBS 0.010633f
C139 B.n99 VSUBS 0.010633f
C140 B.n100 VSUBS 0.023399f
C141 B.n101 VSUBS 0.010633f
C142 B.n102 VSUBS 0.010633f
C143 B.n103 VSUBS 0.010633f
C144 B.n104 VSUBS 0.010633f
C145 B.n105 VSUBS 0.010633f
C146 B.n106 VSUBS 0.010633f
C147 B.n107 VSUBS 0.010633f
C148 B.n108 VSUBS 0.010633f
C149 B.n109 VSUBS 0.010633f
C150 B.n110 VSUBS 0.010633f
C151 B.n111 VSUBS 0.010633f
C152 B.n112 VSUBS 0.010633f
C153 B.n113 VSUBS 0.010633f
C154 B.n114 VSUBS 0.010633f
C155 B.n115 VSUBS 0.010633f
C156 B.n116 VSUBS 0.010633f
C157 B.n117 VSUBS 0.010633f
C158 B.n118 VSUBS 0.010633f
C159 B.n119 VSUBS 0.010633f
C160 B.n120 VSUBS 0.010633f
C161 B.n121 VSUBS 0.010633f
C162 B.n122 VSUBS 0.010633f
C163 B.n123 VSUBS 0.010633f
C164 B.n124 VSUBS 0.010633f
C165 B.n125 VSUBS 0.010633f
C166 B.n126 VSUBS 0.010633f
C167 B.n127 VSUBS 0.010633f
C168 B.n128 VSUBS 0.010633f
C169 B.n129 VSUBS 0.010633f
C170 B.n130 VSUBS 0.010633f
C171 B.n131 VSUBS 0.010633f
C172 B.n132 VSUBS 0.010633f
C173 B.n133 VSUBS 0.010633f
C174 B.n134 VSUBS 0.010633f
C175 B.n135 VSUBS 0.010633f
C176 B.n136 VSUBS 0.010633f
C177 B.n137 VSUBS 0.010633f
C178 B.n138 VSUBS 0.010633f
C179 B.n139 VSUBS 0.010633f
C180 B.n140 VSUBS 0.010633f
C181 B.n141 VSUBS 0.010633f
C182 B.n142 VSUBS 0.010633f
C183 B.n143 VSUBS 0.010633f
C184 B.n144 VSUBS 0.010633f
C185 B.n145 VSUBS 0.010633f
C186 B.n146 VSUBS 0.010633f
C187 B.n147 VSUBS 0.010633f
C188 B.n148 VSUBS 0.010633f
C189 B.n149 VSUBS 0.010633f
C190 B.n150 VSUBS 0.010633f
C191 B.n151 VSUBS 0.010633f
C192 B.n152 VSUBS 0.010633f
C193 B.n153 VSUBS 0.010633f
C194 B.n154 VSUBS 0.010633f
C195 B.n155 VSUBS 0.010633f
C196 B.n156 VSUBS 0.010633f
C197 B.n157 VSUBS 0.010633f
C198 B.n158 VSUBS 0.010633f
C199 B.n159 VSUBS 0.010633f
C200 B.n160 VSUBS 0.010633f
C201 B.n161 VSUBS 0.010633f
C202 B.n162 VSUBS 0.010633f
C203 B.n163 VSUBS 0.010633f
C204 B.n164 VSUBS 0.010633f
C205 B.n165 VSUBS 0.010633f
C206 B.n166 VSUBS 0.010633f
C207 B.n167 VSUBS 0.010633f
C208 B.n168 VSUBS 0.010633f
C209 B.n169 VSUBS 0.010633f
C210 B.n170 VSUBS 0.010633f
C211 B.n171 VSUBS 0.010633f
C212 B.n172 VSUBS 0.010633f
C213 B.n173 VSUBS 0.010633f
C214 B.n174 VSUBS 0.010633f
C215 B.n175 VSUBS 0.010633f
C216 B.n176 VSUBS 0.010633f
C217 B.n177 VSUBS 0.023399f
C218 B.n178 VSUBS 0.025389f
C219 B.n179 VSUBS 0.025389f
C220 B.n180 VSUBS 0.010633f
C221 B.n181 VSUBS 0.010633f
C222 B.n182 VSUBS 0.010633f
C223 B.n183 VSUBS 0.010633f
C224 B.n184 VSUBS 0.010633f
C225 B.n185 VSUBS 0.010633f
C226 B.n186 VSUBS 0.010633f
C227 B.n187 VSUBS 0.010633f
C228 B.n188 VSUBS 0.010633f
C229 B.n189 VSUBS 0.010633f
C230 B.n190 VSUBS 0.010633f
C231 B.n191 VSUBS 0.010633f
C232 B.n192 VSUBS 0.007349f
C233 B.n193 VSUBS 0.024636f
C234 B.n194 VSUBS 0.0086f
C235 B.n195 VSUBS 0.010633f
C236 B.n196 VSUBS 0.010633f
C237 B.n197 VSUBS 0.010633f
C238 B.n198 VSUBS 0.010633f
C239 B.n199 VSUBS 0.010633f
C240 B.n200 VSUBS 0.010633f
C241 B.n201 VSUBS 0.010633f
C242 B.n202 VSUBS 0.010633f
C243 B.n203 VSUBS 0.010633f
C244 B.n204 VSUBS 0.010633f
C245 B.n205 VSUBS 0.010633f
C246 B.n206 VSUBS 0.0086f
C247 B.n207 VSUBS 0.010633f
C248 B.n208 VSUBS 0.010633f
C249 B.n209 VSUBS 0.007349f
C250 B.n210 VSUBS 0.010633f
C251 B.n211 VSUBS 0.010633f
C252 B.n212 VSUBS 0.010633f
C253 B.n213 VSUBS 0.010633f
C254 B.n214 VSUBS 0.010633f
C255 B.n215 VSUBS 0.010633f
C256 B.n216 VSUBS 0.010633f
C257 B.n217 VSUBS 0.010633f
C258 B.n218 VSUBS 0.010633f
C259 B.n219 VSUBS 0.010633f
C260 B.n220 VSUBS 0.010633f
C261 B.n221 VSUBS 0.010633f
C262 B.n222 VSUBS 0.025389f
C263 B.n223 VSUBS 0.023399f
C264 B.n224 VSUBS 0.023399f
C265 B.n225 VSUBS 0.010633f
C266 B.n226 VSUBS 0.010633f
C267 B.n227 VSUBS 0.010633f
C268 B.n228 VSUBS 0.010633f
C269 B.n229 VSUBS 0.010633f
C270 B.n230 VSUBS 0.010633f
C271 B.n231 VSUBS 0.010633f
C272 B.n232 VSUBS 0.010633f
C273 B.n233 VSUBS 0.010633f
C274 B.n234 VSUBS 0.010633f
C275 B.n235 VSUBS 0.010633f
C276 B.n236 VSUBS 0.010633f
C277 B.n237 VSUBS 0.010633f
C278 B.n238 VSUBS 0.010633f
C279 B.n239 VSUBS 0.010633f
C280 B.n240 VSUBS 0.010633f
C281 B.n241 VSUBS 0.010633f
C282 B.n242 VSUBS 0.010633f
C283 B.n243 VSUBS 0.010633f
C284 B.n244 VSUBS 0.010633f
C285 B.n245 VSUBS 0.010633f
C286 B.n246 VSUBS 0.010633f
C287 B.n247 VSUBS 0.010633f
C288 B.n248 VSUBS 0.010633f
C289 B.n249 VSUBS 0.010633f
C290 B.n250 VSUBS 0.010633f
C291 B.n251 VSUBS 0.010633f
C292 B.n252 VSUBS 0.010633f
C293 B.n253 VSUBS 0.010633f
C294 B.n254 VSUBS 0.010633f
C295 B.n255 VSUBS 0.010633f
C296 B.n256 VSUBS 0.010633f
C297 B.n257 VSUBS 0.010633f
C298 B.n258 VSUBS 0.010633f
C299 B.n259 VSUBS 0.010633f
C300 B.n260 VSUBS 0.010633f
C301 B.n261 VSUBS 0.010633f
C302 B.n262 VSUBS 0.010633f
C303 B.n263 VSUBS 0.010633f
C304 B.n264 VSUBS 0.010633f
C305 B.n265 VSUBS 0.010633f
C306 B.n266 VSUBS 0.010633f
C307 B.n267 VSUBS 0.010633f
C308 B.n268 VSUBS 0.010633f
C309 B.n269 VSUBS 0.010633f
C310 B.n270 VSUBS 0.010633f
C311 B.n271 VSUBS 0.010633f
C312 B.n272 VSUBS 0.010633f
C313 B.n273 VSUBS 0.010633f
C314 B.n274 VSUBS 0.010633f
C315 B.n275 VSUBS 0.010633f
C316 B.n276 VSUBS 0.010633f
C317 B.n277 VSUBS 0.010633f
C318 B.n278 VSUBS 0.010633f
C319 B.n279 VSUBS 0.010633f
C320 B.n280 VSUBS 0.010633f
C321 B.n281 VSUBS 0.010633f
C322 B.n282 VSUBS 0.010633f
C323 B.n283 VSUBS 0.010633f
C324 B.n284 VSUBS 0.010633f
C325 B.n285 VSUBS 0.010633f
C326 B.n286 VSUBS 0.010633f
C327 B.n287 VSUBS 0.010633f
C328 B.n288 VSUBS 0.010633f
C329 B.n289 VSUBS 0.010633f
C330 B.n290 VSUBS 0.010633f
C331 B.n291 VSUBS 0.010633f
C332 B.n292 VSUBS 0.010633f
C333 B.n293 VSUBS 0.010633f
C334 B.n294 VSUBS 0.010633f
C335 B.n295 VSUBS 0.010633f
C336 B.n296 VSUBS 0.010633f
C337 B.n297 VSUBS 0.010633f
C338 B.n298 VSUBS 0.010633f
C339 B.n299 VSUBS 0.010633f
C340 B.n300 VSUBS 0.010633f
C341 B.n301 VSUBS 0.010633f
C342 B.n302 VSUBS 0.010633f
C343 B.n303 VSUBS 0.010633f
C344 B.n304 VSUBS 0.010633f
C345 B.n305 VSUBS 0.010633f
C346 B.n306 VSUBS 0.010633f
C347 B.n307 VSUBS 0.010633f
C348 B.n308 VSUBS 0.010633f
C349 B.n309 VSUBS 0.010633f
C350 B.n310 VSUBS 0.010633f
C351 B.n311 VSUBS 0.010633f
C352 B.n312 VSUBS 0.010633f
C353 B.n313 VSUBS 0.010633f
C354 B.n314 VSUBS 0.010633f
C355 B.n315 VSUBS 0.010633f
C356 B.n316 VSUBS 0.010633f
C357 B.n317 VSUBS 0.010633f
C358 B.n318 VSUBS 0.010633f
C359 B.n319 VSUBS 0.010633f
C360 B.n320 VSUBS 0.010633f
C361 B.n321 VSUBS 0.010633f
C362 B.n322 VSUBS 0.010633f
C363 B.n323 VSUBS 0.010633f
C364 B.n324 VSUBS 0.010633f
C365 B.n325 VSUBS 0.010633f
C366 B.n326 VSUBS 0.010633f
C367 B.n327 VSUBS 0.010633f
C368 B.n328 VSUBS 0.010633f
C369 B.n329 VSUBS 0.010633f
C370 B.n330 VSUBS 0.010633f
C371 B.n331 VSUBS 0.010633f
C372 B.n332 VSUBS 0.010633f
C373 B.n333 VSUBS 0.010633f
C374 B.n334 VSUBS 0.010633f
C375 B.n335 VSUBS 0.010633f
C376 B.n336 VSUBS 0.010633f
C377 B.n337 VSUBS 0.010633f
C378 B.n338 VSUBS 0.010633f
C379 B.n339 VSUBS 0.010633f
C380 B.n340 VSUBS 0.010633f
C381 B.n341 VSUBS 0.010633f
C382 B.n342 VSUBS 0.010633f
C383 B.n343 VSUBS 0.024694f
C384 B.n344 VSUBS 0.023399f
C385 B.n345 VSUBS 0.025389f
C386 B.n346 VSUBS 0.010633f
C387 B.n347 VSUBS 0.010633f
C388 B.n348 VSUBS 0.010633f
C389 B.n349 VSUBS 0.010633f
C390 B.n350 VSUBS 0.010633f
C391 B.n351 VSUBS 0.010633f
C392 B.n352 VSUBS 0.010633f
C393 B.n353 VSUBS 0.010633f
C394 B.n354 VSUBS 0.010633f
C395 B.n355 VSUBS 0.010633f
C396 B.n356 VSUBS 0.010633f
C397 B.n357 VSUBS 0.010633f
C398 B.n358 VSUBS 0.010633f
C399 B.n359 VSUBS 0.007349f
C400 B.n360 VSUBS 0.024636f
C401 B.n361 VSUBS 0.0086f
C402 B.n362 VSUBS 0.010633f
C403 B.n363 VSUBS 0.010633f
C404 B.n364 VSUBS 0.010633f
C405 B.n365 VSUBS 0.010633f
C406 B.n366 VSUBS 0.010633f
C407 B.n367 VSUBS 0.010633f
C408 B.n368 VSUBS 0.010633f
C409 B.n369 VSUBS 0.010633f
C410 B.n370 VSUBS 0.010633f
C411 B.n371 VSUBS 0.010633f
C412 B.n372 VSUBS 0.010633f
C413 B.n373 VSUBS 0.0086f
C414 B.n374 VSUBS 0.024636f
C415 B.n375 VSUBS 0.007349f
C416 B.n376 VSUBS 0.010633f
C417 B.n377 VSUBS 0.010633f
C418 B.n378 VSUBS 0.010633f
C419 B.n379 VSUBS 0.010633f
C420 B.n380 VSUBS 0.010633f
C421 B.n381 VSUBS 0.010633f
C422 B.n382 VSUBS 0.010633f
C423 B.n383 VSUBS 0.010633f
C424 B.n384 VSUBS 0.010633f
C425 B.n385 VSUBS 0.010633f
C426 B.n386 VSUBS 0.010633f
C427 B.n387 VSUBS 0.010633f
C428 B.n388 VSUBS 0.010633f
C429 B.n389 VSUBS 0.025389f
C430 B.n390 VSUBS 0.023399f
C431 B.n391 VSUBS 0.023399f
C432 B.n392 VSUBS 0.010633f
C433 B.n393 VSUBS 0.010633f
C434 B.n394 VSUBS 0.010633f
C435 B.n395 VSUBS 0.010633f
C436 B.n396 VSUBS 0.010633f
C437 B.n397 VSUBS 0.010633f
C438 B.n398 VSUBS 0.010633f
C439 B.n399 VSUBS 0.010633f
C440 B.n400 VSUBS 0.010633f
C441 B.n401 VSUBS 0.010633f
C442 B.n402 VSUBS 0.010633f
C443 B.n403 VSUBS 0.010633f
C444 B.n404 VSUBS 0.010633f
C445 B.n405 VSUBS 0.010633f
C446 B.n406 VSUBS 0.010633f
C447 B.n407 VSUBS 0.010633f
C448 B.n408 VSUBS 0.010633f
C449 B.n409 VSUBS 0.010633f
C450 B.n410 VSUBS 0.010633f
C451 B.n411 VSUBS 0.010633f
C452 B.n412 VSUBS 0.010633f
C453 B.n413 VSUBS 0.010633f
C454 B.n414 VSUBS 0.010633f
C455 B.n415 VSUBS 0.010633f
C456 B.n416 VSUBS 0.010633f
C457 B.n417 VSUBS 0.010633f
C458 B.n418 VSUBS 0.010633f
C459 B.n419 VSUBS 0.010633f
C460 B.n420 VSUBS 0.010633f
C461 B.n421 VSUBS 0.010633f
C462 B.n422 VSUBS 0.010633f
C463 B.n423 VSUBS 0.010633f
C464 B.n424 VSUBS 0.010633f
C465 B.n425 VSUBS 0.010633f
C466 B.n426 VSUBS 0.010633f
C467 B.n427 VSUBS 0.010633f
C468 B.n428 VSUBS 0.010633f
C469 B.n429 VSUBS 0.010633f
C470 B.n430 VSUBS 0.010633f
C471 B.n431 VSUBS 0.010633f
C472 B.n432 VSUBS 0.010633f
C473 B.n433 VSUBS 0.010633f
C474 B.n434 VSUBS 0.010633f
C475 B.n435 VSUBS 0.010633f
C476 B.n436 VSUBS 0.010633f
C477 B.n437 VSUBS 0.010633f
C478 B.n438 VSUBS 0.010633f
C479 B.n439 VSUBS 0.010633f
C480 B.n440 VSUBS 0.010633f
C481 B.n441 VSUBS 0.010633f
C482 B.n442 VSUBS 0.010633f
C483 B.n443 VSUBS 0.010633f
C484 B.n444 VSUBS 0.010633f
C485 B.n445 VSUBS 0.010633f
C486 B.n446 VSUBS 0.010633f
C487 B.n447 VSUBS 0.010633f
C488 B.n448 VSUBS 0.010633f
C489 B.n449 VSUBS 0.010633f
C490 B.n450 VSUBS 0.010633f
C491 B.n451 VSUBS 0.024077f
C492 VDD1.t2 VSUBS 0.020303f
C493 VDD1.t0 VSUBS 0.020303f
C494 VDD1.n0 VSUBS 0.067423f
C495 VDD1.t1 VSUBS 0.020303f
C496 VDD1.t3 VSUBS 0.020303f
C497 VDD1.n1 VSUBS 0.151762f
C498 VP.t0 VSUBS 0.369619f
C499 VP.n0 VSUBS 0.438993f
C500 VP.n1 VSUBS 0.053527f
C501 VP.n2 VSUBS 0.043232f
C502 VP.n3 VSUBS 0.053527f
C503 VP.t2 VSUBS 0.369619f
C504 VP.n4 VSUBS 0.438993f
C505 VP.t1 VSUBS 0.883515f
C506 VP.t3 VSUBS 0.865026f
C507 VP.n5 VSUBS 3.233f
C508 VP.n6 VSUBS 2.40598f
C509 VP.n7 VSUBS 0.086378f
C510 VP.n8 VSUBS 0.08113f
C511 VP.n9 VSUBS 0.099261f
C512 VP.n10 VSUBS 0.105824f
C513 VP.n11 VSUBS 0.053527f
C514 VP.n12 VSUBS 0.053527f
C515 VP.n13 VSUBS 0.053527f
C516 VP.n14 VSUBS 0.105824f
C517 VP.n15 VSUBS 0.099261f
C518 VP.n16 VSUBS 0.08113f
C519 VP.n17 VSUBS 0.086378f
C520 VP.n18 VSUBS 0.127797f
C521 VDD2.t1 VSUBS 0.021529f
C522 VDD2.t3 VSUBS 0.021529f
C523 VDD2.n0 VSUBS 0.15513f
C524 VDD2.t0 VSUBS 0.021529f
C525 VDD2.t2 VSUBS 0.021529f
C526 VDD2.n1 VSUBS 0.071415f
C527 VDD2.n2 VSUBS 2.72755f
C528 VTAIL.t5 VSUBS 0.097437f
C529 VTAIL.n0 VSUBS 0.319545f
C530 VTAIL.t2 VSUBS 0.097437f
C531 VTAIL.n1 VSUBS 0.42969f
C532 VTAIL.t3 VSUBS 0.097437f
C533 VTAIL.n2 VSUBS 1.00044f
C534 VTAIL.t7 VSUBS 0.097437f
C535 VTAIL.n3 VSUBS 1.00044f
C536 VTAIL.t6 VSUBS 0.097437f
C537 VTAIL.n4 VSUBS 0.42969f
C538 VTAIL.t1 VSUBS 0.097437f
C539 VTAIL.n5 VSUBS 0.42969f
C540 VTAIL.t0 VSUBS 0.097437f
C541 VTAIL.n6 VSUBS 1.00044f
C542 VTAIL.t4 VSUBS 0.097437f
C543 VTAIL.n7 VSUBS 0.881783f
C544 VN.t0 VSUBS 0.825403f
C545 VN.t2 VSUBS 0.843047f
C546 VN.n0 VSUBS 0.627751f
C547 VN.t3 VSUBS 0.825403f
C548 VN.t1 VSUBS 0.843047f
C549 VN.n1 VSUBS 3.10685f
.ends

