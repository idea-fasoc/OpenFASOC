* NGSPICE file created from diff_pair_sample_1680.ext - technology: sky130A

.subckt diff_pair_sample_1680 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5958 pd=19.22 as=1.5213 ps=9.55 w=9.22 l=1.14
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=3.5958 pd=19.22 as=0 ps=0 w=9.22 l=1.14
X2 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.5958 pd=19.22 as=0 ps=0 w=9.22 l=1.14
X3 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.5958 pd=19.22 as=0 ps=0 w=9.22 l=1.14
X4 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.5958 pd=19.22 as=0 ps=0 w=9.22 l=1.14
X5 VDD2.t1 VN.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5213 pd=9.55 as=3.5958 ps=19.22 w=9.22 l=1.14
X6 VDD2.t3 VN.t2 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5213 pd=9.55 as=3.5958 ps=19.22 w=9.22 l=1.14
X7 VTAIL.t2 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=3.5958 pd=19.22 as=1.5213 ps=9.55 w=9.22 l=1.14
X8 VTAIL.t4 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.5958 pd=19.22 as=1.5213 ps=9.55 w=9.22 l=1.14
X9 VTAIL.t0 VP.t1 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5958 pd=19.22 as=1.5213 ps=9.55 w=9.22 l=1.14
X10 VDD1.t1 VP.t2 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5213 pd=9.55 as=3.5958 ps=19.22 w=9.22 l=1.14
X11 VDD1.t0 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5213 pd=9.55 as=3.5958 ps=19.22 w=9.22 l=1.14
R0 VN.n0 VN.t0 248.404
R1 VN.n1 VN.t1 248.404
R2 VN.n1 VN.t3 248.315
R3 VN.n0 VN.t2 248.315
R4 VN VN.n1 71.372
R5 VN VN.n0 31.2622
R6 VDD2.n2 VDD2.n0 98.0788
R7 VDD2.n2 VDD2.n1 62.614
R8 VDD2.n1 VDD2.t2 2.14801
R9 VDD2.n1 VDD2.t1 2.14801
R10 VDD2.n0 VDD2.t0 2.14801
R11 VDD2.n0 VDD2.t3 2.14801
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n394 VTAIL.n350 289.615
R14 VTAIL.n44 VTAIL.n0 289.615
R15 VTAIL.n94 VTAIL.n50 289.615
R16 VTAIL.n144 VTAIL.n100 289.615
R17 VTAIL.n344 VTAIL.n300 289.615
R18 VTAIL.n294 VTAIL.n250 289.615
R19 VTAIL.n244 VTAIL.n200 289.615
R20 VTAIL.n194 VTAIL.n150 289.615
R21 VTAIL.n367 VTAIL.n366 185
R22 VTAIL.n369 VTAIL.n368 185
R23 VTAIL.n362 VTAIL.n361 185
R24 VTAIL.n375 VTAIL.n374 185
R25 VTAIL.n377 VTAIL.n376 185
R26 VTAIL.n358 VTAIL.n357 185
R27 VTAIL.n384 VTAIL.n383 185
R28 VTAIL.n385 VTAIL.n356 185
R29 VTAIL.n387 VTAIL.n386 185
R30 VTAIL.n354 VTAIL.n353 185
R31 VTAIL.n393 VTAIL.n392 185
R32 VTAIL.n395 VTAIL.n394 185
R33 VTAIL.n17 VTAIL.n16 185
R34 VTAIL.n19 VTAIL.n18 185
R35 VTAIL.n12 VTAIL.n11 185
R36 VTAIL.n25 VTAIL.n24 185
R37 VTAIL.n27 VTAIL.n26 185
R38 VTAIL.n8 VTAIL.n7 185
R39 VTAIL.n34 VTAIL.n33 185
R40 VTAIL.n35 VTAIL.n6 185
R41 VTAIL.n37 VTAIL.n36 185
R42 VTAIL.n4 VTAIL.n3 185
R43 VTAIL.n43 VTAIL.n42 185
R44 VTAIL.n45 VTAIL.n44 185
R45 VTAIL.n67 VTAIL.n66 185
R46 VTAIL.n69 VTAIL.n68 185
R47 VTAIL.n62 VTAIL.n61 185
R48 VTAIL.n75 VTAIL.n74 185
R49 VTAIL.n77 VTAIL.n76 185
R50 VTAIL.n58 VTAIL.n57 185
R51 VTAIL.n84 VTAIL.n83 185
R52 VTAIL.n85 VTAIL.n56 185
R53 VTAIL.n87 VTAIL.n86 185
R54 VTAIL.n54 VTAIL.n53 185
R55 VTAIL.n93 VTAIL.n92 185
R56 VTAIL.n95 VTAIL.n94 185
R57 VTAIL.n117 VTAIL.n116 185
R58 VTAIL.n119 VTAIL.n118 185
R59 VTAIL.n112 VTAIL.n111 185
R60 VTAIL.n125 VTAIL.n124 185
R61 VTAIL.n127 VTAIL.n126 185
R62 VTAIL.n108 VTAIL.n107 185
R63 VTAIL.n134 VTAIL.n133 185
R64 VTAIL.n135 VTAIL.n106 185
R65 VTAIL.n137 VTAIL.n136 185
R66 VTAIL.n104 VTAIL.n103 185
R67 VTAIL.n143 VTAIL.n142 185
R68 VTAIL.n145 VTAIL.n144 185
R69 VTAIL.n345 VTAIL.n344 185
R70 VTAIL.n343 VTAIL.n342 185
R71 VTAIL.n304 VTAIL.n303 185
R72 VTAIL.n308 VTAIL.n306 185
R73 VTAIL.n337 VTAIL.n336 185
R74 VTAIL.n335 VTAIL.n334 185
R75 VTAIL.n310 VTAIL.n309 185
R76 VTAIL.n329 VTAIL.n328 185
R77 VTAIL.n327 VTAIL.n326 185
R78 VTAIL.n314 VTAIL.n313 185
R79 VTAIL.n321 VTAIL.n320 185
R80 VTAIL.n319 VTAIL.n318 185
R81 VTAIL.n295 VTAIL.n294 185
R82 VTAIL.n293 VTAIL.n292 185
R83 VTAIL.n254 VTAIL.n253 185
R84 VTAIL.n258 VTAIL.n256 185
R85 VTAIL.n287 VTAIL.n286 185
R86 VTAIL.n285 VTAIL.n284 185
R87 VTAIL.n260 VTAIL.n259 185
R88 VTAIL.n279 VTAIL.n278 185
R89 VTAIL.n277 VTAIL.n276 185
R90 VTAIL.n264 VTAIL.n263 185
R91 VTAIL.n271 VTAIL.n270 185
R92 VTAIL.n269 VTAIL.n268 185
R93 VTAIL.n245 VTAIL.n244 185
R94 VTAIL.n243 VTAIL.n242 185
R95 VTAIL.n204 VTAIL.n203 185
R96 VTAIL.n208 VTAIL.n206 185
R97 VTAIL.n237 VTAIL.n236 185
R98 VTAIL.n235 VTAIL.n234 185
R99 VTAIL.n210 VTAIL.n209 185
R100 VTAIL.n229 VTAIL.n228 185
R101 VTAIL.n227 VTAIL.n226 185
R102 VTAIL.n214 VTAIL.n213 185
R103 VTAIL.n221 VTAIL.n220 185
R104 VTAIL.n219 VTAIL.n218 185
R105 VTAIL.n195 VTAIL.n194 185
R106 VTAIL.n193 VTAIL.n192 185
R107 VTAIL.n154 VTAIL.n153 185
R108 VTAIL.n158 VTAIL.n156 185
R109 VTAIL.n187 VTAIL.n186 185
R110 VTAIL.n185 VTAIL.n184 185
R111 VTAIL.n160 VTAIL.n159 185
R112 VTAIL.n179 VTAIL.n178 185
R113 VTAIL.n177 VTAIL.n176 185
R114 VTAIL.n164 VTAIL.n163 185
R115 VTAIL.n171 VTAIL.n170 185
R116 VTAIL.n169 VTAIL.n168 185
R117 VTAIL.n365 VTAIL.t5 149.524
R118 VTAIL.n15 VTAIL.t7 149.524
R119 VTAIL.n65 VTAIL.t1 149.524
R120 VTAIL.n115 VTAIL.t2 149.524
R121 VTAIL.n317 VTAIL.t3 149.524
R122 VTAIL.n267 VTAIL.t0 149.524
R123 VTAIL.n217 VTAIL.t6 149.524
R124 VTAIL.n167 VTAIL.t4 149.524
R125 VTAIL.n368 VTAIL.n367 104.615
R126 VTAIL.n368 VTAIL.n361 104.615
R127 VTAIL.n375 VTAIL.n361 104.615
R128 VTAIL.n376 VTAIL.n375 104.615
R129 VTAIL.n376 VTAIL.n357 104.615
R130 VTAIL.n384 VTAIL.n357 104.615
R131 VTAIL.n385 VTAIL.n384 104.615
R132 VTAIL.n386 VTAIL.n385 104.615
R133 VTAIL.n386 VTAIL.n353 104.615
R134 VTAIL.n393 VTAIL.n353 104.615
R135 VTAIL.n394 VTAIL.n393 104.615
R136 VTAIL.n18 VTAIL.n17 104.615
R137 VTAIL.n18 VTAIL.n11 104.615
R138 VTAIL.n25 VTAIL.n11 104.615
R139 VTAIL.n26 VTAIL.n25 104.615
R140 VTAIL.n26 VTAIL.n7 104.615
R141 VTAIL.n34 VTAIL.n7 104.615
R142 VTAIL.n35 VTAIL.n34 104.615
R143 VTAIL.n36 VTAIL.n35 104.615
R144 VTAIL.n36 VTAIL.n3 104.615
R145 VTAIL.n43 VTAIL.n3 104.615
R146 VTAIL.n44 VTAIL.n43 104.615
R147 VTAIL.n68 VTAIL.n67 104.615
R148 VTAIL.n68 VTAIL.n61 104.615
R149 VTAIL.n75 VTAIL.n61 104.615
R150 VTAIL.n76 VTAIL.n75 104.615
R151 VTAIL.n76 VTAIL.n57 104.615
R152 VTAIL.n84 VTAIL.n57 104.615
R153 VTAIL.n85 VTAIL.n84 104.615
R154 VTAIL.n86 VTAIL.n85 104.615
R155 VTAIL.n86 VTAIL.n53 104.615
R156 VTAIL.n93 VTAIL.n53 104.615
R157 VTAIL.n94 VTAIL.n93 104.615
R158 VTAIL.n118 VTAIL.n117 104.615
R159 VTAIL.n118 VTAIL.n111 104.615
R160 VTAIL.n125 VTAIL.n111 104.615
R161 VTAIL.n126 VTAIL.n125 104.615
R162 VTAIL.n126 VTAIL.n107 104.615
R163 VTAIL.n134 VTAIL.n107 104.615
R164 VTAIL.n135 VTAIL.n134 104.615
R165 VTAIL.n136 VTAIL.n135 104.615
R166 VTAIL.n136 VTAIL.n103 104.615
R167 VTAIL.n143 VTAIL.n103 104.615
R168 VTAIL.n144 VTAIL.n143 104.615
R169 VTAIL.n344 VTAIL.n343 104.615
R170 VTAIL.n343 VTAIL.n303 104.615
R171 VTAIL.n308 VTAIL.n303 104.615
R172 VTAIL.n336 VTAIL.n308 104.615
R173 VTAIL.n336 VTAIL.n335 104.615
R174 VTAIL.n335 VTAIL.n309 104.615
R175 VTAIL.n328 VTAIL.n309 104.615
R176 VTAIL.n328 VTAIL.n327 104.615
R177 VTAIL.n327 VTAIL.n313 104.615
R178 VTAIL.n320 VTAIL.n313 104.615
R179 VTAIL.n320 VTAIL.n319 104.615
R180 VTAIL.n294 VTAIL.n293 104.615
R181 VTAIL.n293 VTAIL.n253 104.615
R182 VTAIL.n258 VTAIL.n253 104.615
R183 VTAIL.n286 VTAIL.n258 104.615
R184 VTAIL.n286 VTAIL.n285 104.615
R185 VTAIL.n285 VTAIL.n259 104.615
R186 VTAIL.n278 VTAIL.n259 104.615
R187 VTAIL.n278 VTAIL.n277 104.615
R188 VTAIL.n277 VTAIL.n263 104.615
R189 VTAIL.n270 VTAIL.n263 104.615
R190 VTAIL.n270 VTAIL.n269 104.615
R191 VTAIL.n244 VTAIL.n243 104.615
R192 VTAIL.n243 VTAIL.n203 104.615
R193 VTAIL.n208 VTAIL.n203 104.615
R194 VTAIL.n236 VTAIL.n208 104.615
R195 VTAIL.n236 VTAIL.n235 104.615
R196 VTAIL.n235 VTAIL.n209 104.615
R197 VTAIL.n228 VTAIL.n209 104.615
R198 VTAIL.n228 VTAIL.n227 104.615
R199 VTAIL.n227 VTAIL.n213 104.615
R200 VTAIL.n220 VTAIL.n213 104.615
R201 VTAIL.n220 VTAIL.n219 104.615
R202 VTAIL.n194 VTAIL.n193 104.615
R203 VTAIL.n193 VTAIL.n153 104.615
R204 VTAIL.n158 VTAIL.n153 104.615
R205 VTAIL.n186 VTAIL.n158 104.615
R206 VTAIL.n186 VTAIL.n185 104.615
R207 VTAIL.n185 VTAIL.n159 104.615
R208 VTAIL.n178 VTAIL.n159 104.615
R209 VTAIL.n178 VTAIL.n177 104.615
R210 VTAIL.n177 VTAIL.n163 104.615
R211 VTAIL.n170 VTAIL.n163 104.615
R212 VTAIL.n170 VTAIL.n169 104.615
R213 VTAIL.n367 VTAIL.t5 52.3082
R214 VTAIL.n17 VTAIL.t7 52.3082
R215 VTAIL.n67 VTAIL.t1 52.3082
R216 VTAIL.n117 VTAIL.t2 52.3082
R217 VTAIL.n319 VTAIL.t3 52.3082
R218 VTAIL.n269 VTAIL.t0 52.3082
R219 VTAIL.n219 VTAIL.t6 52.3082
R220 VTAIL.n169 VTAIL.t4 52.3082
R221 VTAIL.n399 VTAIL.n398 31.7975
R222 VTAIL.n49 VTAIL.n48 31.7975
R223 VTAIL.n99 VTAIL.n98 31.7975
R224 VTAIL.n149 VTAIL.n148 31.7975
R225 VTAIL.n349 VTAIL.n348 31.7975
R226 VTAIL.n299 VTAIL.n298 31.7975
R227 VTAIL.n249 VTAIL.n248 31.7975
R228 VTAIL.n199 VTAIL.n198 31.7975
R229 VTAIL.n399 VTAIL.n349 21.5824
R230 VTAIL.n199 VTAIL.n149 21.5824
R231 VTAIL.n387 VTAIL.n354 13.1884
R232 VTAIL.n37 VTAIL.n4 13.1884
R233 VTAIL.n87 VTAIL.n54 13.1884
R234 VTAIL.n137 VTAIL.n104 13.1884
R235 VTAIL.n306 VTAIL.n304 13.1884
R236 VTAIL.n256 VTAIL.n254 13.1884
R237 VTAIL.n206 VTAIL.n204 13.1884
R238 VTAIL.n156 VTAIL.n154 13.1884
R239 VTAIL.n388 VTAIL.n356 12.8005
R240 VTAIL.n392 VTAIL.n391 12.8005
R241 VTAIL.n38 VTAIL.n6 12.8005
R242 VTAIL.n42 VTAIL.n41 12.8005
R243 VTAIL.n88 VTAIL.n56 12.8005
R244 VTAIL.n92 VTAIL.n91 12.8005
R245 VTAIL.n138 VTAIL.n106 12.8005
R246 VTAIL.n142 VTAIL.n141 12.8005
R247 VTAIL.n342 VTAIL.n341 12.8005
R248 VTAIL.n338 VTAIL.n337 12.8005
R249 VTAIL.n292 VTAIL.n291 12.8005
R250 VTAIL.n288 VTAIL.n287 12.8005
R251 VTAIL.n242 VTAIL.n241 12.8005
R252 VTAIL.n238 VTAIL.n237 12.8005
R253 VTAIL.n192 VTAIL.n191 12.8005
R254 VTAIL.n188 VTAIL.n187 12.8005
R255 VTAIL.n383 VTAIL.n382 12.0247
R256 VTAIL.n395 VTAIL.n352 12.0247
R257 VTAIL.n33 VTAIL.n32 12.0247
R258 VTAIL.n45 VTAIL.n2 12.0247
R259 VTAIL.n83 VTAIL.n82 12.0247
R260 VTAIL.n95 VTAIL.n52 12.0247
R261 VTAIL.n133 VTAIL.n132 12.0247
R262 VTAIL.n145 VTAIL.n102 12.0247
R263 VTAIL.n345 VTAIL.n302 12.0247
R264 VTAIL.n334 VTAIL.n307 12.0247
R265 VTAIL.n295 VTAIL.n252 12.0247
R266 VTAIL.n284 VTAIL.n257 12.0247
R267 VTAIL.n245 VTAIL.n202 12.0247
R268 VTAIL.n234 VTAIL.n207 12.0247
R269 VTAIL.n195 VTAIL.n152 12.0247
R270 VTAIL.n184 VTAIL.n157 12.0247
R271 VTAIL.n381 VTAIL.n358 11.249
R272 VTAIL.n396 VTAIL.n350 11.249
R273 VTAIL.n31 VTAIL.n8 11.249
R274 VTAIL.n46 VTAIL.n0 11.249
R275 VTAIL.n81 VTAIL.n58 11.249
R276 VTAIL.n96 VTAIL.n50 11.249
R277 VTAIL.n131 VTAIL.n108 11.249
R278 VTAIL.n146 VTAIL.n100 11.249
R279 VTAIL.n346 VTAIL.n300 11.249
R280 VTAIL.n333 VTAIL.n310 11.249
R281 VTAIL.n296 VTAIL.n250 11.249
R282 VTAIL.n283 VTAIL.n260 11.249
R283 VTAIL.n246 VTAIL.n200 11.249
R284 VTAIL.n233 VTAIL.n210 11.249
R285 VTAIL.n196 VTAIL.n150 11.249
R286 VTAIL.n183 VTAIL.n160 11.249
R287 VTAIL.n378 VTAIL.n377 10.4732
R288 VTAIL.n28 VTAIL.n27 10.4732
R289 VTAIL.n78 VTAIL.n77 10.4732
R290 VTAIL.n128 VTAIL.n127 10.4732
R291 VTAIL.n330 VTAIL.n329 10.4732
R292 VTAIL.n280 VTAIL.n279 10.4732
R293 VTAIL.n230 VTAIL.n229 10.4732
R294 VTAIL.n180 VTAIL.n179 10.4732
R295 VTAIL.n366 VTAIL.n365 10.2747
R296 VTAIL.n16 VTAIL.n15 10.2747
R297 VTAIL.n66 VTAIL.n65 10.2747
R298 VTAIL.n116 VTAIL.n115 10.2747
R299 VTAIL.n318 VTAIL.n317 10.2747
R300 VTAIL.n268 VTAIL.n267 10.2747
R301 VTAIL.n218 VTAIL.n217 10.2747
R302 VTAIL.n168 VTAIL.n167 10.2747
R303 VTAIL.n374 VTAIL.n360 9.69747
R304 VTAIL.n24 VTAIL.n10 9.69747
R305 VTAIL.n74 VTAIL.n60 9.69747
R306 VTAIL.n124 VTAIL.n110 9.69747
R307 VTAIL.n326 VTAIL.n312 9.69747
R308 VTAIL.n276 VTAIL.n262 9.69747
R309 VTAIL.n226 VTAIL.n212 9.69747
R310 VTAIL.n176 VTAIL.n162 9.69747
R311 VTAIL.n398 VTAIL.n397 9.45567
R312 VTAIL.n48 VTAIL.n47 9.45567
R313 VTAIL.n98 VTAIL.n97 9.45567
R314 VTAIL.n148 VTAIL.n147 9.45567
R315 VTAIL.n348 VTAIL.n347 9.45567
R316 VTAIL.n298 VTAIL.n297 9.45567
R317 VTAIL.n248 VTAIL.n247 9.45567
R318 VTAIL.n198 VTAIL.n197 9.45567
R319 VTAIL.n397 VTAIL.n396 9.3005
R320 VTAIL.n352 VTAIL.n351 9.3005
R321 VTAIL.n391 VTAIL.n390 9.3005
R322 VTAIL.n364 VTAIL.n363 9.3005
R323 VTAIL.n371 VTAIL.n370 9.3005
R324 VTAIL.n373 VTAIL.n372 9.3005
R325 VTAIL.n360 VTAIL.n359 9.3005
R326 VTAIL.n379 VTAIL.n378 9.3005
R327 VTAIL.n381 VTAIL.n380 9.3005
R328 VTAIL.n382 VTAIL.n355 9.3005
R329 VTAIL.n389 VTAIL.n388 9.3005
R330 VTAIL.n47 VTAIL.n46 9.3005
R331 VTAIL.n2 VTAIL.n1 9.3005
R332 VTAIL.n41 VTAIL.n40 9.3005
R333 VTAIL.n14 VTAIL.n13 9.3005
R334 VTAIL.n21 VTAIL.n20 9.3005
R335 VTAIL.n23 VTAIL.n22 9.3005
R336 VTAIL.n10 VTAIL.n9 9.3005
R337 VTAIL.n29 VTAIL.n28 9.3005
R338 VTAIL.n31 VTAIL.n30 9.3005
R339 VTAIL.n32 VTAIL.n5 9.3005
R340 VTAIL.n39 VTAIL.n38 9.3005
R341 VTAIL.n97 VTAIL.n96 9.3005
R342 VTAIL.n52 VTAIL.n51 9.3005
R343 VTAIL.n91 VTAIL.n90 9.3005
R344 VTAIL.n64 VTAIL.n63 9.3005
R345 VTAIL.n71 VTAIL.n70 9.3005
R346 VTAIL.n73 VTAIL.n72 9.3005
R347 VTAIL.n60 VTAIL.n59 9.3005
R348 VTAIL.n79 VTAIL.n78 9.3005
R349 VTAIL.n81 VTAIL.n80 9.3005
R350 VTAIL.n82 VTAIL.n55 9.3005
R351 VTAIL.n89 VTAIL.n88 9.3005
R352 VTAIL.n147 VTAIL.n146 9.3005
R353 VTAIL.n102 VTAIL.n101 9.3005
R354 VTAIL.n141 VTAIL.n140 9.3005
R355 VTAIL.n114 VTAIL.n113 9.3005
R356 VTAIL.n121 VTAIL.n120 9.3005
R357 VTAIL.n123 VTAIL.n122 9.3005
R358 VTAIL.n110 VTAIL.n109 9.3005
R359 VTAIL.n129 VTAIL.n128 9.3005
R360 VTAIL.n131 VTAIL.n130 9.3005
R361 VTAIL.n132 VTAIL.n105 9.3005
R362 VTAIL.n139 VTAIL.n138 9.3005
R363 VTAIL.n316 VTAIL.n315 9.3005
R364 VTAIL.n323 VTAIL.n322 9.3005
R365 VTAIL.n325 VTAIL.n324 9.3005
R366 VTAIL.n312 VTAIL.n311 9.3005
R367 VTAIL.n331 VTAIL.n330 9.3005
R368 VTAIL.n333 VTAIL.n332 9.3005
R369 VTAIL.n307 VTAIL.n305 9.3005
R370 VTAIL.n339 VTAIL.n338 9.3005
R371 VTAIL.n347 VTAIL.n346 9.3005
R372 VTAIL.n302 VTAIL.n301 9.3005
R373 VTAIL.n341 VTAIL.n340 9.3005
R374 VTAIL.n266 VTAIL.n265 9.3005
R375 VTAIL.n273 VTAIL.n272 9.3005
R376 VTAIL.n275 VTAIL.n274 9.3005
R377 VTAIL.n262 VTAIL.n261 9.3005
R378 VTAIL.n281 VTAIL.n280 9.3005
R379 VTAIL.n283 VTAIL.n282 9.3005
R380 VTAIL.n257 VTAIL.n255 9.3005
R381 VTAIL.n289 VTAIL.n288 9.3005
R382 VTAIL.n297 VTAIL.n296 9.3005
R383 VTAIL.n252 VTAIL.n251 9.3005
R384 VTAIL.n291 VTAIL.n290 9.3005
R385 VTAIL.n216 VTAIL.n215 9.3005
R386 VTAIL.n223 VTAIL.n222 9.3005
R387 VTAIL.n225 VTAIL.n224 9.3005
R388 VTAIL.n212 VTAIL.n211 9.3005
R389 VTAIL.n231 VTAIL.n230 9.3005
R390 VTAIL.n233 VTAIL.n232 9.3005
R391 VTAIL.n207 VTAIL.n205 9.3005
R392 VTAIL.n239 VTAIL.n238 9.3005
R393 VTAIL.n247 VTAIL.n246 9.3005
R394 VTAIL.n202 VTAIL.n201 9.3005
R395 VTAIL.n241 VTAIL.n240 9.3005
R396 VTAIL.n166 VTAIL.n165 9.3005
R397 VTAIL.n173 VTAIL.n172 9.3005
R398 VTAIL.n175 VTAIL.n174 9.3005
R399 VTAIL.n162 VTAIL.n161 9.3005
R400 VTAIL.n181 VTAIL.n180 9.3005
R401 VTAIL.n183 VTAIL.n182 9.3005
R402 VTAIL.n157 VTAIL.n155 9.3005
R403 VTAIL.n189 VTAIL.n188 9.3005
R404 VTAIL.n197 VTAIL.n196 9.3005
R405 VTAIL.n152 VTAIL.n151 9.3005
R406 VTAIL.n191 VTAIL.n190 9.3005
R407 VTAIL.n373 VTAIL.n362 8.92171
R408 VTAIL.n23 VTAIL.n12 8.92171
R409 VTAIL.n73 VTAIL.n62 8.92171
R410 VTAIL.n123 VTAIL.n112 8.92171
R411 VTAIL.n325 VTAIL.n314 8.92171
R412 VTAIL.n275 VTAIL.n264 8.92171
R413 VTAIL.n225 VTAIL.n214 8.92171
R414 VTAIL.n175 VTAIL.n164 8.92171
R415 VTAIL.n370 VTAIL.n369 8.14595
R416 VTAIL.n20 VTAIL.n19 8.14595
R417 VTAIL.n70 VTAIL.n69 8.14595
R418 VTAIL.n120 VTAIL.n119 8.14595
R419 VTAIL.n322 VTAIL.n321 8.14595
R420 VTAIL.n272 VTAIL.n271 8.14595
R421 VTAIL.n222 VTAIL.n221 8.14595
R422 VTAIL.n172 VTAIL.n171 8.14595
R423 VTAIL.n366 VTAIL.n364 7.3702
R424 VTAIL.n16 VTAIL.n14 7.3702
R425 VTAIL.n66 VTAIL.n64 7.3702
R426 VTAIL.n116 VTAIL.n114 7.3702
R427 VTAIL.n318 VTAIL.n316 7.3702
R428 VTAIL.n268 VTAIL.n266 7.3702
R429 VTAIL.n218 VTAIL.n216 7.3702
R430 VTAIL.n168 VTAIL.n166 7.3702
R431 VTAIL.n369 VTAIL.n364 5.81868
R432 VTAIL.n19 VTAIL.n14 5.81868
R433 VTAIL.n69 VTAIL.n64 5.81868
R434 VTAIL.n119 VTAIL.n114 5.81868
R435 VTAIL.n321 VTAIL.n316 5.81868
R436 VTAIL.n271 VTAIL.n266 5.81868
R437 VTAIL.n221 VTAIL.n216 5.81868
R438 VTAIL.n171 VTAIL.n166 5.81868
R439 VTAIL.n370 VTAIL.n362 5.04292
R440 VTAIL.n20 VTAIL.n12 5.04292
R441 VTAIL.n70 VTAIL.n62 5.04292
R442 VTAIL.n120 VTAIL.n112 5.04292
R443 VTAIL.n322 VTAIL.n314 5.04292
R444 VTAIL.n272 VTAIL.n264 5.04292
R445 VTAIL.n222 VTAIL.n214 5.04292
R446 VTAIL.n172 VTAIL.n164 5.04292
R447 VTAIL.n374 VTAIL.n373 4.26717
R448 VTAIL.n24 VTAIL.n23 4.26717
R449 VTAIL.n74 VTAIL.n73 4.26717
R450 VTAIL.n124 VTAIL.n123 4.26717
R451 VTAIL.n326 VTAIL.n325 4.26717
R452 VTAIL.n276 VTAIL.n275 4.26717
R453 VTAIL.n226 VTAIL.n225 4.26717
R454 VTAIL.n176 VTAIL.n175 4.26717
R455 VTAIL.n377 VTAIL.n360 3.49141
R456 VTAIL.n27 VTAIL.n10 3.49141
R457 VTAIL.n77 VTAIL.n60 3.49141
R458 VTAIL.n127 VTAIL.n110 3.49141
R459 VTAIL.n329 VTAIL.n312 3.49141
R460 VTAIL.n279 VTAIL.n262 3.49141
R461 VTAIL.n229 VTAIL.n212 3.49141
R462 VTAIL.n179 VTAIL.n162 3.49141
R463 VTAIL.n365 VTAIL.n363 2.84303
R464 VTAIL.n15 VTAIL.n13 2.84303
R465 VTAIL.n65 VTAIL.n63 2.84303
R466 VTAIL.n115 VTAIL.n113 2.84303
R467 VTAIL.n317 VTAIL.n315 2.84303
R468 VTAIL.n267 VTAIL.n265 2.84303
R469 VTAIL.n217 VTAIL.n215 2.84303
R470 VTAIL.n167 VTAIL.n165 2.84303
R471 VTAIL.n378 VTAIL.n358 2.71565
R472 VTAIL.n398 VTAIL.n350 2.71565
R473 VTAIL.n28 VTAIL.n8 2.71565
R474 VTAIL.n48 VTAIL.n0 2.71565
R475 VTAIL.n78 VTAIL.n58 2.71565
R476 VTAIL.n98 VTAIL.n50 2.71565
R477 VTAIL.n128 VTAIL.n108 2.71565
R478 VTAIL.n148 VTAIL.n100 2.71565
R479 VTAIL.n348 VTAIL.n300 2.71565
R480 VTAIL.n330 VTAIL.n310 2.71565
R481 VTAIL.n298 VTAIL.n250 2.71565
R482 VTAIL.n280 VTAIL.n260 2.71565
R483 VTAIL.n248 VTAIL.n200 2.71565
R484 VTAIL.n230 VTAIL.n210 2.71565
R485 VTAIL.n198 VTAIL.n150 2.71565
R486 VTAIL.n180 VTAIL.n160 2.71565
R487 VTAIL.n383 VTAIL.n381 1.93989
R488 VTAIL.n396 VTAIL.n395 1.93989
R489 VTAIL.n33 VTAIL.n31 1.93989
R490 VTAIL.n46 VTAIL.n45 1.93989
R491 VTAIL.n83 VTAIL.n81 1.93989
R492 VTAIL.n96 VTAIL.n95 1.93989
R493 VTAIL.n133 VTAIL.n131 1.93989
R494 VTAIL.n146 VTAIL.n145 1.93989
R495 VTAIL.n346 VTAIL.n345 1.93989
R496 VTAIL.n334 VTAIL.n333 1.93989
R497 VTAIL.n296 VTAIL.n295 1.93989
R498 VTAIL.n284 VTAIL.n283 1.93989
R499 VTAIL.n246 VTAIL.n245 1.93989
R500 VTAIL.n234 VTAIL.n233 1.93989
R501 VTAIL.n196 VTAIL.n195 1.93989
R502 VTAIL.n184 VTAIL.n183 1.93989
R503 VTAIL.n249 VTAIL.n199 1.26774
R504 VTAIL.n349 VTAIL.n299 1.26774
R505 VTAIL.n149 VTAIL.n99 1.26774
R506 VTAIL.n382 VTAIL.n356 1.16414
R507 VTAIL.n392 VTAIL.n352 1.16414
R508 VTAIL.n32 VTAIL.n6 1.16414
R509 VTAIL.n42 VTAIL.n2 1.16414
R510 VTAIL.n82 VTAIL.n56 1.16414
R511 VTAIL.n92 VTAIL.n52 1.16414
R512 VTAIL.n132 VTAIL.n106 1.16414
R513 VTAIL.n142 VTAIL.n102 1.16414
R514 VTAIL.n342 VTAIL.n302 1.16414
R515 VTAIL.n337 VTAIL.n307 1.16414
R516 VTAIL.n292 VTAIL.n252 1.16414
R517 VTAIL.n287 VTAIL.n257 1.16414
R518 VTAIL.n242 VTAIL.n202 1.16414
R519 VTAIL.n237 VTAIL.n207 1.16414
R520 VTAIL.n192 VTAIL.n152 1.16414
R521 VTAIL.n187 VTAIL.n157 1.16414
R522 VTAIL VTAIL.n49 0.69231
R523 VTAIL VTAIL.n399 0.575931
R524 VTAIL.n299 VTAIL.n249 0.470328
R525 VTAIL.n99 VTAIL.n49 0.470328
R526 VTAIL.n388 VTAIL.n387 0.388379
R527 VTAIL.n391 VTAIL.n354 0.388379
R528 VTAIL.n38 VTAIL.n37 0.388379
R529 VTAIL.n41 VTAIL.n4 0.388379
R530 VTAIL.n88 VTAIL.n87 0.388379
R531 VTAIL.n91 VTAIL.n54 0.388379
R532 VTAIL.n138 VTAIL.n137 0.388379
R533 VTAIL.n141 VTAIL.n104 0.388379
R534 VTAIL.n341 VTAIL.n304 0.388379
R535 VTAIL.n338 VTAIL.n306 0.388379
R536 VTAIL.n291 VTAIL.n254 0.388379
R537 VTAIL.n288 VTAIL.n256 0.388379
R538 VTAIL.n241 VTAIL.n204 0.388379
R539 VTAIL.n238 VTAIL.n206 0.388379
R540 VTAIL.n191 VTAIL.n154 0.388379
R541 VTAIL.n188 VTAIL.n156 0.388379
R542 VTAIL.n371 VTAIL.n363 0.155672
R543 VTAIL.n372 VTAIL.n371 0.155672
R544 VTAIL.n372 VTAIL.n359 0.155672
R545 VTAIL.n379 VTAIL.n359 0.155672
R546 VTAIL.n380 VTAIL.n379 0.155672
R547 VTAIL.n380 VTAIL.n355 0.155672
R548 VTAIL.n389 VTAIL.n355 0.155672
R549 VTAIL.n390 VTAIL.n389 0.155672
R550 VTAIL.n390 VTAIL.n351 0.155672
R551 VTAIL.n397 VTAIL.n351 0.155672
R552 VTAIL.n21 VTAIL.n13 0.155672
R553 VTAIL.n22 VTAIL.n21 0.155672
R554 VTAIL.n22 VTAIL.n9 0.155672
R555 VTAIL.n29 VTAIL.n9 0.155672
R556 VTAIL.n30 VTAIL.n29 0.155672
R557 VTAIL.n30 VTAIL.n5 0.155672
R558 VTAIL.n39 VTAIL.n5 0.155672
R559 VTAIL.n40 VTAIL.n39 0.155672
R560 VTAIL.n40 VTAIL.n1 0.155672
R561 VTAIL.n47 VTAIL.n1 0.155672
R562 VTAIL.n71 VTAIL.n63 0.155672
R563 VTAIL.n72 VTAIL.n71 0.155672
R564 VTAIL.n72 VTAIL.n59 0.155672
R565 VTAIL.n79 VTAIL.n59 0.155672
R566 VTAIL.n80 VTAIL.n79 0.155672
R567 VTAIL.n80 VTAIL.n55 0.155672
R568 VTAIL.n89 VTAIL.n55 0.155672
R569 VTAIL.n90 VTAIL.n89 0.155672
R570 VTAIL.n90 VTAIL.n51 0.155672
R571 VTAIL.n97 VTAIL.n51 0.155672
R572 VTAIL.n121 VTAIL.n113 0.155672
R573 VTAIL.n122 VTAIL.n121 0.155672
R574 VTAIL.n122 VTAIL.n109 0.155672
R575 VTAIL.n129 VTAIL.n109 0.155672
R576 VTAIL.n130 VTAIL.n129 0.155672
R577 VTAIL.n130 VTAIL.n105 0.155672
R578 VTAIL.n139 VTAIL.n105 0.155672
R579 VTAIL.n140 VTAIL.n139 0.155672
R580 VTAIL.n140 VTAIL.n101 0.155672
R581 VTAIL.n147 VTAIL.n101 0.155672
R582 VTAIL.n347 VTAIL.n301 0.155672
R583 VTAIL.n340 VTAIL.n301 0.155672
R584 VTAIL.n340 VTAIL.n339 0.155672
R585 VTAIL.n339 VTAIL.n305 0.155672
R586 VTAIL.n332 VTAIL.n305 0.155672
R587 VTAIL.n332 VTAIL.n331 0.155672
R588 VTAIL.n331 VTAIL.n311 0.155672
R589 VTAIL.n324 VTAIL.n311 0.155672
R590 VTAIL.n324 VTAIL.n323 0.155672
R591 VTAIL.n323 VTAIL.n315 0.155672
R592 VTAIL.n297 VTAIL.n251 0.155672
R593 VTAIL.n290 VTAIL.n251 0.155672
R594 VTAIL.n290 VTAIL.n289 0.155672
R595 VTAIL.n289 VTAIL.n255 0.155672
R596 VTAIL.n282 VTAIL.n255 0.155672
R597 VTAIL.n282 VTAIL.n281 0.155672
R598 VTAIL.n281 VTAIL.n261 0.155672
R599 VTAIL.n274 VTAIL.n261 0.155672
R600 VTAIL.n274 VTAIL.n273 0.155672
R601 VTAIL.n273 VTAIL.n265 0.155672
R602 VTAIL.n247 VTAIL.n201 0.155672
R603 VTAIL.n240 VTAIL.n201 0.155672
R604 VTAIL.n240 VTAIL.n239 0.155672
R605 VTAIL.n239 VTAIL.n205 0.155672
R606 VTAIL.n232 VTAIL.n205 0.155672
R607 VTAIL.n232 VTAIL.n231 0.155672
R608 VTAIL.n231 VTAIL.n211 0.155672
R609 VTAIL.n224 VTAIL.n211 0.155672
R610 VTAIL.n224 VTAIL.n223 0.155672
R611 VTAIL.n223 VTAIL.n215 0.155672
R612 VTAIL.n197 VTAIL.n151 0.155672
R613 VTAIL.n190 VTAIL.n151 0.155672
R614 VTAIL.n190 VTAIL.n189 0.155672
R615 VTAIL.n189 VTAIL.n155 0.155672
R616 VTAIL.n182 VTAIL.n155 0.155672
R617 VTAIL.n182 VTAIL.n181 0.155672
R618 VTAIL.n181 VTAIL.n161 0.155672
R619 VTAIL.n174 VTAIL.n161 0.155672
R620 VTAIL.n174 VTAIL.n173 0.155672
R621 VTAIL.n173 VTAIL.n165 0.155672
R622 B.n561 B.n560 585
R623 B.n234 B.n79 585
R624 B.n233 B.n232 585
R625 B.n231 B.n230 585
R626 B.n229 B.n228 585
R627 B.n227 B.n226 585
R628 B.n225 B.n224 585
R629 B.n223 B.n222 585
R630 B.n221 B.n220 585
R631 B.n219 B.n218 585
R632 B.n217 B.n216 585
R633 B.n215 B.n214 585
R634 B.n213 B.n212 585
R635 B.n211 B.n210 585
R636 B.n209 B.n208 585
R637 B.n207 B.n206 585
R638 B.n205 B.n204 585
R639 B.n203 B.n202 585
R640 B.n201 B.n200 585
R641 B.n199 B.n198 585
R642 B.n197 B.n196 585
R643 B.n195 B.n194 585
R644 B.n193 B.n192 585
R645 B.n191 B.n190 585
R646 B.n189 B.n188 585
R647 B.n187 B.n186 585
R648 B.n185 B.n184 585
R649 B.n183 B.n182 585
R650 B.n181 B.n180 585
R651 B.n179 B.n178 585
R652 B.n177 B.n176 585
R653 B.n175 B.n174 585
R654 B.n173 B.n172 585
R655 B.n170 B.n169 585
R656 B.n168 B.n167 585
R657 B.n166 B.n165 585
R658 B.n164 B.n163 585
R659 B.n162 B.n161 585
R660 B.n160 B.n159 585
R661 B.n158 B.n157 585
R662 B.n156 B.n155 585
R663 B.n154 B.n153 585
R664 B.n152 B.n151 585
R665 B.n149 B.n148 585
R666 B.n147 B.n146 585
R667 B.n145 B.n144 585
R668 B.n143 B.n142 585
R669 B.n141 B.n140 585
R670 B.n139 B.n138 585
R671 B.n137 B.n136 585
R672 B.n135 B.n134 585
R673 B.n133 B.n132 585
R674 B.n131 B.n130 585
R675 B.n129 B.n128 585
R676 B.n127 B.n126 585
R677 B.n125 B.n124 585
R678 B.n123 B.n122 585
R679 B.n121 B.n120 585
R680 B.n119 B.n118 585
R681 B.n117 B.n116 585
R682 B.n115 B.n114 585
R683 B.n113 B.n112 585
R684 B.n111 B.n110 585
R685 B.n109 B.n108 585
R686 B.n107 B.n106 585
R687 B.n105 B.n104 585
R688 B.n103 B.n102 585
R689 B.n101 B.n100 585
R690 B.n99 B.n98 585
R691 B.n97 B.n96 585
R692 B.n95 B.n94 585
R693 B.n93 B.n92 585
R694 B.n91 B.n90 585
R695 B.n89 B.n88 585
R696 B.n87 B.n86 585
R697 B.n85 B.n84 585
R698 B.n559 B.n41 585
R699 B.n564 B.n41 585
R700 B.n558 B.n40 585
R701 B.n565 B.n40 585
R702 B.n557 B.n556 585
R703 B.n556 B.n36 585
R704 B.n555 B.n35 585
R705 B.n571 B.n35 585
R706 B.n554 B.n34 585
R707 B.n572 B.n34 585
R708 B.n553 B.n33 585
R709 B.n573 B.n33 585
R710 B.n552 B.n551 585
R711 B.n551 B.n29 585
R712 B.n550 B.n28 585
R713 B.n579 B.n28 585
R714 B.n549 B.n27 585
R715 B.n580 B.n27 585
R716 B.n548 B.n26 585
R717 B.n581 B.n26 585
R718 B.n547 B.n546 585
R719 B.n546 B.n22 585
R720 B.n545 B.n21 585
R721 B.n587 B.n21 585
R722 B.n544 B.n20 585
R723 B.n588 B.n20 585
R724 B.n543 B.n19 585
R725 B.n589 B.n19 585
R726 B.n542 B.n541 585
R727 B.n541 B.n15 585
R728 B.n540 B.n14 585
R729 B.n595 B.n14 585
R730 B.n539 B.n13 585
R731 B.n596 B.n13 585
R732 B.n538 B.n12 585
R733 B.n597 B.n12 585
R734 B.n537 B.n536 585
R735 B.n536 B.n8 585
R736 B.n535 B.n7 585
R737 B.n603 B.n7 585
R738 B.n534 B.n6 585
R739 B.n604 B.n6 585
R740 B.n533 B.n5 585
R741 B.n605 B.n5 585
R742 B.n532 B.n531 585
R743 B.n531 B.n4 585
R744 B.n530 B.n235 585
R745 B.n530 B.n529 585
R746 B.n520 B.n236 585
R747 B.n237 B.n236 585
R748 B.n522 B.n521 585
R749 B.n523 B.n522 585
R750 B.n519 B.n242 585
R751 B.n242 B.n241 585
R752 B.n518 B.n517 585
R753 B.n517 B.n516 585
R754 B.n244 B.n243 585
R755 B.n245 B.n244 585
R756 B.n509 B.n508 585
R757 B.n510 B.n509 585
R758 B.n507 B.n249 585
R759 B.n253 B.n249 585
R760 B.n506 B.n505 585
R761 B.n505 B.n504 585
R762 B.n251 B.n250 585
R763 B.n252 B.n251 585
R764 B.n497 B.n496 585
R765 B.n498 B.n497 585
R766 B.n495 B.n258 585
R767 B.n258 B.n257 585
R768 B.n494 B.n493 585
R769 B.n493 B.n492 585
R770 B.n260 B.n259 585
R771 B.n261 B.n260 585
R772 B.n485 B.n484 585
R773 B.n486 B.n485 585
R774 B.n483 B.n266 585
R775 B.n266 B.n265 585
R776 B.n482 B.n481 585
R777 B.n481 B.n480 585
R778 B.n268 B.n267 585
R779 B.n269 B.n268 585
R780 B.n473 B.n472 585
R781 B.n474 B.n473 585
R782 B.n471 B.n274 585
R783 B.n274 B.n273 585
R784 B.n466 B.n465 585
R785 B.n464 B.n314 585
R786 B.n463 B.n313 585
R787 B.n468 B.n313 585
R788 B.n462 B.n461 585
R789 B.n460 B.n459 585
R790 B.n458 B.n457 585
R791 B.n456 B.n455 585
R792 B.n454 B.n453 585
R793 B.n452 B.n451 585
R794 B.n450 B.n449 585
R795 B.n448 B.n447 585
R796 B.n446 B.n445 585
R797 B.n444 B.n443 585
R798 B.n442 B.n441 585
R799 B.n440 B.n439 585
R800 B.n438 B.n437 585
R801 B.n436 B.n435 585
R802 B.n434 B.n433 585
R803 B.n432 B.n431 585
R804 B.n430 B.n429 585
R805 B.n428 B.n427 585
R806 B.n426 B.n425 585
R807 B.n424 B.n423 585
R808 B.n422 B.n421 585
R809 B.n420 B.n419 585
R810 B.n418 B.n417 585
R811 B.n416 B.n415 585
R812 B.n414 B.n413 585
R813 B.n412 B.n411 585
R814 B.n410 B.n409 585
R815 B.n408 B.n407 585
R816 B.n406 B.n405 585
R817 B.n404 B.n403 585
R818 B.n402 B.n401 585
R819 B.n400 B.n399 585
R820 B.n398 B.n397 585
R821 B.n396 B.n395 585
R822 B.n394 B.n393 585
R823 B.n392 B.n391 585
R824 B.n390 B.n389 585
R825 B.n388 B.n387 585
R826 B.n386 B.n385 585
R827 B.n384 B.n383 585
R828 B.n382 B.n381 585
R829 B.n380 B.n379 585
R830 B.n378 B.n377 585
R831 B.n376 B.n375 585
R832 B.n374 B.n373 585
R833 B.n372 B.n371 585
R834 B.n370 B.n369 585
R835 B.n368 B.n367 585
R836 B.n366 B.n365 585
R837 B.n364 B.n363 585
R838 B.n362 B.n361 585
R839 B.n360 B.n359 585
R840 B.n358 B.n357 585
R841 B.n356 B.n355 585
R842 B.n354 B.n353 585
R843 B.n352 B.n351 585
R844 B.n350 B.n349 585
R845 B.n348 B.n347 585
R846 B.n346 B.n345 585
R847 B.n344 B.n343 585
R848 B.n342 B.n341 585
R849 B.n340 B.n339 585
R850 B.n338 B.n337 585
R851 B.n336 B.n335 585
R852 B.n334 B.n333 585
R853 B.n332 B.n331 585
R854 B.n330 B.n329 585
R855 B.n328 B.n327 585
R856 B.n326 B.n325 585
R857 B.n324 B.n323 585
R858 B.n322 B.n321 585
R859 B.n276 B.n275 585
R860 B.n470 B.n469 585
R861 B.n469 B.n468 585
R862 B.n272 B.n271 585
R863 B.n273 B.n272 585
R864 B.n476 B.n475 585
R865 B.n475 B.n474 585
R866 B.n477 B.n270 585
R867 B.n270 B.n269 585
R868 B.n479 B.n478 585
R869 B.n480 B.n479 585
R870 B.n264 B.n263 585
R871 B.n265 B.n264 585
R872 B.n488 B.n487 585
R873 B.n487 B.n486 585
R874 B.n489 B.n262 585
R875 B.n262 B.n261 585
R876 B.n491 B.n490 585
R877 B.n492 B.n491 585
R878 B.n256 B.n255 585
R879 B.n257 B.n256 585
R880 B.n500 B.n499 585
R881 B.n499 B.n498 585
R882 B.n501 B.n254 585
R883 B.n254 B.n252 585
R884 B.n503 B.n502 585
R885 B.n504 B.n503 585
R886 B.n248 B.n247 585
R887 B.n253 B.n248 585
R888 B.n512 B.n511 585
R889 B.n511 B.n510 585
R890 B.n513 B.n246 585
R891 B.n246 B.n245 585
R892 B.n515 B.n514 585
R893 B.n516 B.n515 585
R894 B.n240 B.n239 585
R895 B.n241 B.n240 585
R896 B.n525 B.n524 585
R897 B.n524 B.n523 585
R898 B.n526 B.n238 585
R899 B.n238 B.n237 585
R900 B.n528 B.n527 585
R901 B.n529 B.n528 585
R902 B.n2 B.n0 585
R903 B.n4 B.n2 585
R904 B.n3 B.n1 585
R905 B.n604 B.n3 585
R906 B.n602 B.n601 585
R907 B.n603 B.n602 585
R908 B.n600 B.n9 585
R909 B.n9 B.n8 585
R910 B.n599 B.n598 585
R911 B.n598 B.n597 585
R912 B.n11 B.n10 585
R913 B.n596 B.n11 585
R914 B.n594 B.n593 585
R915 B.n595 B.n594 585
R916 B.n592 B.n16 585
R917 B.n16 B.n15 585
R918 B.n591 B.n590 585
R919 B.n590 B.n589 585
R920 B.n18 B.n17 585
R921 B.n588 B.n18 585
R922 B.n586 B.n585 585
R923 B.n587 B.n586 585
R924 B.n584 B.n23 585
R925 B.n23 B.n22 585
R926 B.n583 B.n582 585
R927 B.n582 B.n581 585
R928 B.n25 B.n24 585
R929 B.n580 B.n25 585
R930 B.n578 B.n577 585
R931 B.n579 B.n578 585
R932 B.n576 B.n30 585
R933 B.n30 B.n29 585
R934 B.n575 B.n574 585
R935 B.n574 B.n573 585
R936 B.n32 B.n31 585
R937 B.n572 B.n32 585
R938 B.n570 B.n569 585
R939 B.n571 B.n570 585
R940 B.n568 B.n37 585
R941 B.n37 B.n36 585
R942 B.n567 B.n566 585
R943 B.n566 B.n565 585
R944 B.n39 B.n38 585
R945 B.n564 B.n39 585
R946 B.n607 B.n606 585
R947 B.n606 B.n605 585
R948 B.n466 B.n272 550.159
R949 B.n84 B.n39 550.159
R950 B.n469 B.n274 550.159
R951 B.n561 B.n41 550.159
R952 B.n318 B.t4 398.705
R953 B.n315 B.t15 398.705
R954 B.n82 B.t8 398.705
R955 B.n80 B.t12 398.705
R956 B.n318 B.t7 262.505
R957 B.n80 B.t13 262.505
R958 B.n315 B.t17 262.505
R959 B.n82 B.t10 262.505
R960 B.n563 B.n562 256.663
R961 B.n563 B.n78 256.663
R962 B.n563 B.n77 256.663
R963 B.n563 B.n76 256.663
R964 B.n563 B.n75 256.663
R965 B.n563 B.n74 256.663
R966 B.n563 B.n73 256.663
R967 B.n563 B.n72 256.663
R968 B.n563 B.n71 256.663
R969 B.n563 B.n70 256.663
R970 B.n563 B.n69 256.663
R971 B.n563 B.n68 256.663
R972 B.n563 B.n67 256.663
R973 B.n563 B.n66 256.663
R974 B.n563 B.n65 256.663
R975 B.n563 B.n64 256.663
R976 B.n563 B.n63 256.663
R977 B.n563 B.n62 256.663
R978 B.n563 B.n61 256.663
R979 B.n563 B.n60 256.663
R980 B.n563 B.n59 256.663
R981 B.n563 B.n58 256.663
R982 B.n563 B.n57 256.663
R983 B.n563 B.n56 256.663
R984 B.n563 B.n55 256.663
R985 B.n563 B.n54 256.663
R986 B.n563 B.n53 256.663
R987 B.n563 B.n52 256.663
R988 B.n563 B.n51 256.663
R989 B.n563 B.n50 256.663
R990 B.n563 B.n49 256.663
R991 B.n563 B.n48 256.663
R992 B.n563 B.n47 256.663
R993 B.n563 B.n46 256.663
R994 B.n563 B.n45 256.663
R995 B.n563 B.n44 256.663
R996 B.n563 B.n43 256.663
R997 B.n563 B.n42 256.663
R998 B.n468 B.n467 256.663
R999 B.n468 B.n277 256.663
R1000 B.n468 B.n278 256.663
R1001 B.n468 B.n279 256.663
R1002 B.n468 B.n280 256.663
R1003 B.n468 B.n281 256.663
R1004 B.n468 B.n282 256.663
R1005 B.n468 B.n283 256.663
R1006 B.n468 B.n284 256.663
R1007 B.n468 B.n285 256.663
R1008 B.n468 B.n286 256.663
R1009 B.n468 B.n287 256.663
R1010 B.n468 B.n288 256.663
R1011 B.n468 B.n289 256.663
R1012 B.n468 B.n290 256.663
R1013 B.n468 B.n291 256.663
R1014 B.n468 B.n292 256.663
R1015 B.n468 B.n293 256.663
R1016 B.n468 B.n294 256.663
R1017 B.n468 B.n295 256.663
R1018 B.n468 B.n296 256.663
R1019 B.n468 B.n297 256.663
R1020 B.n468 B.n298 256.663
R1021 B.n468 B.n299 256.663
R1022 B.n468 B.n300 256.663
R1023 B.n468 B.n301 256.663
R1024 B.n468 B.n302 256.663
R1025 B.n468 B.n303 256.663
R1026 B.n468 B.n304 256.663
R1027 B.n468 B.n305 256.663
R1028 B.n468 B.n306 256.663
R1029 B.n468 B.n307 256.663
R1030 B.n468 B.n308 256.663
R1031 B.n468 B.n309 256.663
R1032 B.n468 B.n310 256.663
R1033 B.n468 B.n311 256.663
R1034 B.n468 B.n312 256.663
R1035 B.n319 B.t6 233.996
R1036 B.n81 B.t14 233.996
R1037 B.n316 B.t16 233.995
R1038 B.n83 B.t11 233.995
R1039 B.n475 B.n272 163.367
R1040 B.n475 B.n270 163.367
R1041 B.n479 B.n270 163.367
R1042 B.n479 B.n264 163.367
R1043 B.n487 B.n264 163.367
R1044 B.n487 B.n262 163.367
R1045 B.n491 B.n262 163.367
R1046 B.n491 B.n256 163.367
R1047 B.n499 B.n256 163.367
R1048 B.n499 B.n254 163.367
R1049 B.n503 B.n254 163.367
R1050 B.n503 B.n248 163.367
R1051 B.n511 B.n248 163.367
R1052 B.n511 B.n246 163.367
R1053 B.n515 B.n246 163.367
R1054 B.n515 B.n240 163.367
R1055 B.n524 B.n240 163.367
R1056 B.n524 B.n238 163.367
R1057 B.n528 B.n238 163.367
R1058 B.n528 B.n2 163.367
R1059 B.n606 B.n2 163.367
R1060 B.n606 B.n3 163.367
R1061 B.n602 B.n3 163.367
R1062 B.n602 B.n9 163.367
R1063 B.n598 B.n9 163.367
R1064 B.n598 B.n11 163.367
R1065 B.n594 B.n11 163.367
R1066 B.n594 B.n16 163.367
R1067 B.n590 B.n16 163.367
R1068 B.n590 B.n18 163.367
R1069 B.n586 B.n18 163.367
R1070 B.n586 B.n23 163.367
R1071 B.n582 B.n23 163.367
R1072 B.n582 B.n25 163.367
R1073 B.n578 B.n25 163.367
R1074 B.n578 B.n30 163.367
R1075 B.n574 B.n30 163.367
R1076 B.n574 B.n32 163.367
R1077 B.n570 B.n32 163.367
R1078 B.n570 B.n37 163.367
R1079 B.n566 B.n37 163.367
R1080 B.n566 B.n39 163.367
R1081 B.n314 B.n313 163.367
R1082 B.n461 B.n313 163.367
R1083 B.n459 B.n458 163.367
R1084 B.n455 B.n454 163.367
R1085 B.n451 B.n450 163.367
R1086 B.n447 B.n446 163.367
R1087 B.n443 B.n442 163.367
R1088 B.n439 B.n438 163.367
R1089 B.n435 B.n434 163.367
R1090 B.n431 B.n430 163.367
R1091 B.n427 B.n426 163.367
R1092 B.n423 B.n422 163.367
R1093 B.n419 B.n418 163.367
R1094 B.n415 B.n414 163.367
R1095 B.n411 B.n410 163.367
R1096 B.n407 B.n406 163.367
R1097 B.n403 B.n402 163.367
R1098 B.n399 B.n398 163.367
R1099 B.n395 B.n394 163.367
R1100 B.n391 B.n390 163.367
R1101 B.n387 B.n386 163.367
R1102 B.n383 B.n382 163.367
R1103 B.n379 B.n378 163.367
R1104 B.n375 B.n374 163.367
R1105 B.n371 B.n370 163.367
R1106 B.n367 B.n366 163.367
R1107 B.n363 B.n362 163.367
R1108 B.n359 B.n358 163.367
R1109 B.n355 B.n354 163.367
R1110 B.n351 B.n350 163.367
R1111 B.n347 B.n346 163.367
R1112 B.n343 B.n342 163.367
R1113 B.n339 B.n338 163.367
R1114 B.n335 B.n334 163.367
R1115 B.n331 B.n330 163.367
R1116 B.n327 B.n326 163.367
R1117 B.n323 B.n322 163.367
R1118 B.n469 B.n276 163.367
R1119 B.n473 B.n274 163.367
R1120 B.n473 B.n268 163.367
R1121 B.n481 B.n268 163.367
R1122 B.n481 B.n266 163.367
R1123 B.n485 B.n266 163.367
R1124 B.n485 B.n260 163.367
R1125 B.n493 B.n260 163.367
R1126 B.n493 B.n258 163.367
R1127 B.n497 B.n258 163.367
R1128 B.n497 B.n251 163.367
R1129 B.n505 B.n251 163.367
R1130 B.n505 B.n249 163.367
R1131 B.n509 B.n249 163.367
R1132 B.n509 B.n244 163.367
R1133 B.n517 B.n244 163.367
R1134 B.n517 B.n242 163.367
R1135 B.n522 B.n242 163.367
R1136 B.n522 B.n236 163.367
R1137 B.n530 B.n236 163.367
R1138 B.n531 B.n530 163.367
R1139 B.n531 B.n5 163.367
R1140 B.n6 B.n5 163.367
R1141 B.n7 B.n6 163.367
R1142 B.n536 B.n7 163.367
R1143 B.n536 B.n12 163.367
R1144 B.n13 B.n12 163.367
R1145 B.n14 B.n13 163.367
R1146 B.n541 B.n14 163.367
R1147 B.n541 B.n19 163.367
R1148 B.n20 B.n19 163.367
R1149 B.n21 B.n20 163.367
R1150 B.n546 B.n21 163.367
R1151 B.n546 B.n26 163.367
R1152 B.n27 B.n26 163.367
R1153 B.n28 B.n27 163.367
R1154 B.n551 B.n28 163.367
R1155 B.n551 B.n33 163.367
R1156 B.n34 B.n33 163.367
R1157 B.n35 B.n34 163.367
R1158 B.n556 B.n35 163.367
R1159 B.n556 B.n40 163.367
R1160 B.n41 B.n40 163.367
R1161 B.n88 B.n87 163.367
R1162 B.n92 B.n91 163.367
R1163 B.n96 B.n95 163.367
R1164 B.n100 B.n99 163.367
R1165 B.n104 B.n103 163.367
R1166 B.n108 B.n107 163.367
R1167 B.n112 B.n111 163.367
R1168 B.n116 B.n115 163.367
R1169 B.n120 B.n119 163.367
R1170 B.n124 B.n123 163.367
R1171 B.n128 B.n127 163.367
R1172 B.n132 B.n131 163.367
R1173 B.n136 B.n135 163.367
R1174 B.n140 B.n139 163.367
R1175 B.n144 B.n143 163.367
R1176 B.n148 B.n147 163.367
R1177 B.n153 B.n152 163.367
R1178 B.n157 B.n156 163.367
R1179 B.n161 B.n160 163.367
R1180 B.n165 B.n164 163.367
R1181 B.n169 B.n168 163.367
R1182 B.n174 B.n173 163.367
R1183 B.n178 B.n177 163.367
R1184 B.n182 B.n181 163.367
R1185 B.n186 B.n185 163.367
R1186 B.n190 B.n189 163.367
R1187 B.n194 B.n193 163.367
R1188 B.n198 B.n197 163.367
R1189 B.n202 B.n201 163.367
R1190 B.n206 B.n205 163.367
R1191 B.n210 B.n209 163.367
R1192 B.n214 B.n213 163.367
R1193 B.n218 B.n217 163.367
R1194 B.n222 B.n221 163.367
R1195 B.n226 B.n225 163.367
R1196 B.n230 B.n229 163.367
R1197 B.n232 B.n79 163.367
R1198 B.n468 B.n273 97.8963
R1199 B.n564 B.n563 97.8963
R1200 B.n467 B.n466 71.676
R1201 B.n461 B.n277 71.676
R1202 B.n458 B.n278 71.676
R1203 B.n454 B.n279 71.676
R1204 B.n450 B.n280 71.676
R1205 B.n446 B.n281 71.676
R1206 B.n442 B.n282 71.676
R1207 B.n438 B.n283 71.676
R1208 B.n434 B.n284 71.676
R1209 B.n430 B.n285 71.676
R1210 B.n426 B.n286 71.676
R1211 B.n422 B.n287 71.676
R1212 B.n418 B.n288 71.676
R1213 B.n414 B.n289 71.676
R1214 B.n410 B.n290 71.676
R1215 B.n406 B.n291 71.676
R1216 B.n402 B.n292 71.676
R1217 B.n398 B.n293 71.676
R1218 B.n394 B.n294 71.676
R1219 B.n390 B.n295 71.676
R1220 B.n386 B.n296 71.676
R1221 B.n382 B.n297 71.676
R1222 B.n378 B.n298 71.676
R1223 B.n374 B.n299 71.676
R1224 B.n370 B.n300 71.676
R1225 B.n366 B.n301 71.676
R1226 B.n362 B.n302 71.676
R1227 B.n358 B.n303 71.676
R1228 B.n354 B.n304 71.676
R1229 B.n350 B.n305 71.676
R1230 B.n346 B.n306 71.676
R1231 B.n342 B.n307 71.676
R1232 B.n338 B.n308 71.676
R1233 B.n334 B.n309 71.676
R1234 B.n330 B.n310 71.676
R1235 B.n326 B.n311 71.676
R1236 B.n322 B.n312 71.676
R1237 B.n84 B.n42 71.676
R1238 B.n88 B.n43 71.676
R1239 B.n92 B.n44 71.676
R1240 B.n96 B.n45 71.676
R1241 B.n100 B.n46 71.676
R1242 B.n104 B.n47 71.676
R1243 B.n108 B.n48 71.676
R1244 B.n112 B.n49 71.676
R1245 B.n116 B.n50 71.676
R1246 B.n120 B.n51 71.676
R1247 B.n124 B.n52 71.676
R1248 B.n128 B.n53 71.676
R1249 B.n132 B.n54 71.676
R1250 B.n136 B.n55 71.676
R1251 B.n140 B.n56 71.676
R1252 B.n144 B.n57 71.676
R1253 B.n148 B.n58 71.676
R1254 B.n153 B.n59 71.676
R1255 B.n157 B.n60 71.676
R1256 B.n161 B.n61 71.676
R1257 B.n165 B.n62 71.676
R1258 B.n169 B.n63 71.676
R1259 B.n174 B.n64 71.676
R1260 B.n178 B.n65 71.676
R1261 B.n182 B.n66 71.676
R1262 B.n186 B.n67 71.676
R1263 B.n190 B.n68 71.676
R1264 B.n194 B.n69 71.676
R1265 B.n198 B.n70 71.676
R1266 B.n202 B.n71 71.676
R1267 B.n206 B.n72 71.676
R1268 B.n210 B.n73 71.676
R1269 B.n214 B.n74 71.676
R1270 B.n218 B.n75 71.676
R1271 B.n222 B.n76 71.676
R1272 B.n226 B.n77 71.676
R1273 B.n230 B.n78 71.676
R1274 B.n562 B.n79 71.676
R1275 B.n562 B.n561 71.676
R1276 B.n232 B.n78 71.676
R1277 B.n229 B.n77 71.676
R1278 B.n225 B.n76 71.676
R1279 B.n221 B.n75 71.676
R1280 B.n217 B.n74 71.676
R1281 B.n213 B.n73 71.676
R1282 B.n209 B.n72 71.676
R1283 B.n205 B.n71 71.676
R1284 B.n201 B.n70 71.676
R1285 B.n197 B.n69 71.676
R1286 B.n193 B.n68 71.676
R1287 B.n189 B.n67 71.676
R1288 B.n185 B.n66 71.676
R1289 B.n181 B.n65 71.676
R1290 B.n177 B.n64 71.676
R1291 B.n173 B.n63 71.676
R1292 B.n168 B.n62 71.676
R1293 B.n164 B.n61 71.676
R1294 B.n160 B.n60 71.676
R1295 B.n156 B.n59 71.676
R1296 B.n152 B.n58 71.676
R1297 B.n147 B.n57 71.676
R1298 B.n143 B.n56 71.676
R1299 B.n139 B.n55 71.676
R1300 B.n135 B.n54 71.676
R1301 B.n131 B.n53 71.676
R1302 B.n127 B.n52 71.676
R1303 B.n123 B.n51 71.676
R1304 B.n119 B.n50 71.676
R1305 B.n115 B.n49 71.676
R1306 B.n111 B.n48 71.676
R1307 B.n107 B.n47 71.676
R1308 B.n103 B.n46 71.676
R1309 B.n99 B.n45 71.676
R1310 B.n95 B.n44 71.676
R1311 B.n91 B.n43 71.676
R1312 B.n87 B.n42 71.676
R1313 B.n467 B.n314 71.676
R1314 B.n459 B.n277 71.676
R1315 B.n455 B.n278 71.676
R1316 B.n451 B.n279 71.676
R1317 B.n447 B.n280 71.676
R1318 B.n443 B.n281 71.676
R1319 B.n439 B.n282 71.676
R1320 B.n435 B.n283 71.676
R1321 B.n431 B.n284 71.676
R1322 B.n427 B.n285 71.676
R1323 B.n423 B.n286 71.676
R1324 B.n419 B.n287 71.676
R1325 B.n415 B.n288 71.676
R1326 B.n411 B.n289 71.676
R1327 B.n407 B.n290 71.676
R1328 B.n403 B.n291 71.676
R1329 B.n399 B.n292 71.676
R1330 B.n395 B.n293 71.676
R1331 B.n391 B.n294 71.676
R1332 B.n387 B.n295 71.676
R1333 B.n383 B.n296 71.676
R1334 B.n379 B.n297 71.676
R1335 B.n375 B.n298 71.676
R1336 B.n371 B.n299 71.676
R1337 B.n367 B.n300 71.676
R1338 B.n363 B.n301 71.676
R1339 B.n359 B.n302 71.676
R1340 B.n355 B.n303 71.676
R1341 B.n351 B.n304 71.676
R1342 B.n347 B.n305 71.676
R1343 B.n343 B.n306 71.676
R1344 B.n339 B.n307 71.676
R1345 B.n335 B.n308 71.676
R1346 B.n331 B.n309 71.676
R1347 B.n327 B.n310 71.676
R1348 B.n323 B.n311 71.676
R1349 B.n312 B.n276 71.676
R1350 B.n320 B.n319 59.5399
R1351 B.n317 B.n316 59.5399
R1352 B.n150 B.n83 59.5399
R1353 B.n171 B.n81 59.5399
R1354 B.n474 B.n273 51.6045
R1355 B.n474 B.n269 51.6045
R1356 B.n480 B.n269 51.6045
R1357 B.n480 B.n265 51.6045
R1358 B.n486 B.n265 51.6045
R1359 B.n492 B.n261 51.6045
R1360 B.n492 B.n257 51.6045
R1361 B.n498 B.n257 51.6045
R1362 B.n498 B.n252 51.6045
R1363 B.n504 B.n252 51.6045
R1364 B.n504 B.n253 51.6045
R1365 B.n510 B.n245 51.6045
R1366 B.n516 B.n245 51.6045
R1367 B.n516 B.n241 51.6045
R1368 B.n523 B.n241 51.6045
R1369 B.n529 B.n237 51.6045
R1370 B.n529 B.n4 51.6045
R1371 B.n605 B.n4 51.6045
R1372 B.n605 B.n604 51.6045
R1373 B.n604 B.n603 51.6045
R1374 B.n603 B.n8 51.6045
R1375 B.n597 B.n596 51.6045
R1376 B.n596 B.n595 51.6045
R1377 B.n595 B.n15 51.6045
R1378 B.n589 B.n15 51.6045
R1379 B.n588 B.n587 51.6045
R1380 B.n587 B.n22 51.6045
R1381 B.n581 B.n22 51.6045
R1382 B.n581 B.n580 51.6045
R1383 B.n580 B.n579 51.6045
R1384 B.n579 B.n29 51.6045
R1385 B.n573 B.n572 51.6045
R1386 B.n572 B.n571 51.6045
R1387 B.n571 B.n36 51.6045
R1388 B.n565 B.n36 51.6045
R1389 B.n565 B.n564 51.6045
R1390 B.n253 B.t2 47.0512
R1391 B.t3 B.n588 47.0512
R1392 B.t1 B.n237 39.4624
R1393 B.t0 B.n8 39.4624
R1394 B.n85 B.n38 35.7468
R1395 B.n471 B.n470 35.7468
R1396 B.n465 B.n271 35.7468
R1397 B.n560 B.n559 35.7468
R1398 B.t5 B.n261 31.8736
R1399 B.t9 B.n29 31.8736
R1400 B.n319 B.n318 28.5096
R1401 B.n316 B.n315 28.5096
R1402 B.n83 B.n82 28.5096
R1403 B.n81 B.n80 28.5096
R1404 B.n486 B.t5 19.7314
R1405 B.n573 B.t9 19.7314
R1406 B B.n607 18.0485
R1407 B.n523 B.t1 12.1426
R1408 B.n597 B.t0 12.1426
R1409 B.n86 B.n85 10.6151
R1410 B.n89 B.n86 10.6151
R1411 B.n90 B.n89 10.6151
R1412 B.n93 B.n90 10.6151
R1413 B.n94 B.n93 10.6151
R1414 B.n97 B.n94 10.6151
R1415 B.n98 B.n97 10.6151
R1416 B.n101 B.n98 10.6151
R1417 B.n102 B.n101 10.6151
R1418 B.n105 B.n102 10.6151
R1419 B.n106 B.n105 10.6151
R1420 B.n109 B.n106 10.6151
R1421 B.n110 B.n109 10.6151
R1422 B.n113 B.n110 10.6151
R1423 B.n114 B.n113 10.6151
R1424 B.n117 B.n114 10.6151
R1425 B.n118 B.n117 10.6151
R1426 B.n121 B.n118 10.6151
R1427 B.n122 B.n121 10.6151
R1428 B.n125 B.n122 10.6151
R1429 B.n126 B.n125 10.6151
R1430 B.n129 B.n126 10.6151
R1431 B.n130 B.n129 10.6151
R1432 B.n133 B.n130 10.6151
R1433 B.n134 B.n133 10.6151
R1434 B.n137 B.n134 10.6151
R1435 B.n138 B.n137 10.6151
R1436 B.n141 B.n138 10.6151
R1437 B.n142 B.n141 10.6151
R1438 B.n145 B.n142 10.6151
R1439 B.n146 B.n145 10.6151
R1440 B.n149 B.n146 10.6151
R1441 B.n154 B.n151 10.6151
R1442 B.n155 B.n154 10.6151
R1443 B.n158 B.n155 10.6151
R1444 B.n159 B.n158 10.6151
R1445 B.n162 B.n159 10.6151
R1446 B.n163 B.n162 10.6151
R1447 B.n166 B.n163 10.6151
R1448 B.n167 B.n166 10.6151
R1449 B.n170 B.n167 10.6151
R1450 B.n175 B.n172 10.6151
R1451 B.n176 B.n175 10.6151
R1452 B.n179 B.n176 10.6151
R1453 B.n180 B.n179 10.6151
R1454 B.n183 B.n180 10.6151
R1455 B.n184 B.n183 10.6151
R1456 B.n187 B.n184 10.6151
R1457 B.n188 B.n187 10.6151
R1458 B.n191 B.n188 10.6151
R1459 B.n192 B.n191 10.6151
R1460 B.n195 B.n192 10.6151
R1461 B.n196 B.n195 10.6151
R1462 B.n199 B.n196 10.6151
R1463 B.n200 B.n199 10.6151
R1464 B.n203 B.n200 10.6151
R1465 B.n204 B.n203 10.6151
R1466 B.n207 B.n204 10.6151
R1467 B.n208 B.n207 10.6151
R1468 B.n211 B.n208 10.6151
R1469 B.n212 B.n211 10.6151
R1470 B.n215 B.n212 10.6151
R1471 B.n216 B.n215 10.6151
R1472 B.n219 B.n216 10.6151
R1473 B.n220 B.n219 10.6151
R1474 B.n223 B.n220 10.6151
R1475 B.n224 B.n223 10.6151
R1476 B.n227 B.n224 10.6151
R1477 B.n228 B.n227 10.6151
R1478 B.n231 B.n228 10.6151
R1479 B.n233 B.n231 10.6151
R1480 B.n234 B.n233 10.6151
R1481 B.n560 B.n234 10.6151
R1482 B.n472 B.n471 10.6151
R1483 B.n472 B.n267 10.6151
R1484 B.n482 B.n267 10.6151
R1485 B.n483 B.n482 10.6151
R1486 B.n484 B.n483 10.6151
R1487 B.n484 B.n259 10.6151
R1488 B.n494 B.n259 10.6151
R1489 B.n495 B.n494 10.6151
R1490 B.n496 B.n495 10.6151
R1491 B.n496 B.n250 10.6151
R1492 B.n506 B.n250 10.6151
R1493 B.n507 B.n506 10.6151
R1494 B.n508 B.n507 10.6151
R1495 B.n508 B.n243 10.6151
R1496 B.n518 B.n243 10.6151
R1497 B.n519 B.n518 10.6151
R1498 B.n521 B.n519 10.6151
R1499 B.n521 B.n520 10.6151
R1500 B.n520 B.n235 10.6151
R1501 B.n532 B.n235 10.6151
R1502 B.n533 B.n532 10.6151
R1503 B.n534 B.n533 10.6151
R1504 B.n535 B.n534 10.6151
R1505 B.n537 B.n535 10.6151
R1506 B.n538 B.n537 10.6151
R1507 B.n539 B.n538 10.6151
R1508 B.n540 B.n539 10.6151
R1509 B.n542 B.n540 10.6151
R1510 B.n543 B.n542 10.6151
R1511 B.n544 B.n543 10.6151
R1512 B.n545 B.n544 10.6151
R1513 B.n547 B.n545 10.6151
R1514 B.n548 B.n547 10.6151
R1515 B.n549 B.n548 10.6151
R1516 B.n550 B.n549 10.6151
R1517 B.n552 B.n550 10.6151
R1518 B.n553 B.n552 10.6151
R1519 B.n554 B.n553 10.6151
R1520 B.n555 B.n554 10.6151
R1521 B.n557 B.n555 10.6151
R1522 B.n558 B.n557 10.6151
R1523 B.n559 B.n558 10.6151
R1524 B.n465 B.n464 10.6151
R1525 B.n464 B.n463 10.6151
R1526 B.n463 B.n462 10.6151
R1527 B.n462 B.n460 10.6151
R1528 B.n460 B.n457 10.6151
R1529 B.n457 B.n456 10.6151
R1530 B.n456 B.n453 10.6151
R1531 B.n453 B.n452 10.6151
R1532 B.n452 B.n449 10.6151
R1533 B.n449 B.n448 10.6151
R1534 B.n448 B.n445 10.6151
R1535 B.n445 B.n444 10.6151
R1536 B.n444 B.n441 10.6151
R1537 B.n441 B.n440 10.6151
R1538 B.n440 B.n437 10.6151
R1539 B.n437 B.n436 10.6151
R1540 B.n436 B.n433 10.6151
R1541 B.n433 B.n432 10.6151
R1542 B.n432 B.n429 10.6151
R1543 B.n429 B.n428 10.6151
R1544 B.n428 B.n425 10.6151
R1545 B.n425 B.n424 10.6151
R1546 B.n424 B.n421 10.6151
R1547 B.n421 B.n420 10.6151
R1548 B.n420 B.n417 10.6151
R1549 B.n417 B.n416 10.6151
R1550 B.n416 B.n413 10.6151
R1551 B.n413 B.n412 10.6151
R1552 B.n412 B.n409 10.6151
R1553 B.n409 B.n408 10.6151
R1554 B.n408 B.n405 10.6151
R1555 B.n405 B.n404 10.6151
R1556 B.n401 B.n400 10.6151
R1557 B.n400 B.n397 10.6151
R1558 B.n397 B.n396 10.6151
R1559 B.n396 B.n393 10.6151
R1560 B.n393 B.n392 10.6151
R1561 B.n392 B.n389 10.6151
R1562 B.n389 B.n388 10.6151
R1563 B.n388 B.n385 10.6151
R1564 B.n385 B.n384 10.6151
R1565 B.n381 B.n380 10.6151
R1566 B.n380 B.n377 10.6151
R1567 B.n377 B.n376 10.6151
R1568 B.n376 B.n373 10.6151
R1569 B.n373 B.n372 10.6151
R1570 B.n372 B.n369 10.6151
R1571 B.n369 B.n368 10.6151
R1572 B.n368 B.n365 10.6151
R1573 B.n365 B.n364 10.6151
R1574 B.n364 B.n361 10.6151
R1575 B.n361 B.n360 10.6151
R1576 B.n360 B.n357 10.6151
R1577 B.n357 B.n356 10.6151
R1578 B.n356 B.n353 10.6151
R1579 B.n353 B.n352 10.6151
R1580 B.n352 B.n349 10.6151
R1581 B.n349 B.n348 10.6151
R1582 B.n348 B.n345 10.6151
R1583 B.n345 B.n344 10.6151
R1584 B.n344 B.n341 10.6151
R1585 B.n341 B.n340 10.6151
R1586 B.n340 B.n337 10.6151
R1587 B.n337 B.n336 10.6151
R1588 B.n336 B.n333 10.6151
R1589 B.n333 B.n332 10.6151
R1590 B.n332 B.n329 10.6151
R1591 B.n329 B.n328 10.6151
R1592 B.n328 B.n325 10.6151
R1593 B.n325 B.n324 10.6151
R1594 B.n324 B.n321 10.6151
R1595 B.n321 B.n275 10.6151
R1596 B.n470 B.n275 10.6151
R1597 B.n476 B.n271 10.6151
R1598 B.n477 B.n476 10.6151
R1599 B.n478 B.n477 10.6151
R1600 B.n478 B.n263 10.6151
R1601 B.n488 B.n263 10.6151
R1602 B.n489 B.n488 10.6151
R1603 B.n490 B.n489 10.6151
R1604 B.n490 B.n255 10.6151
R1605 B.n500 B.n255 10.6151
R1606 B.n501 B.n500 10.6151
R1607 B.n502 B.n501 10.6151
R1608 B.n502 B.n247 10.6151
R1609 B.n512 B.n247 10.6151
R1610 B.n513 B.n512 10.6151
R1611 B.n514 B.n513 10.6151
R1612 B.n514 B.n239 10.6151
R1613 B.n525 B.n239 10.6151
R1614 B.n526 B.n525 10.6151
R1615 B.n527 B.n526 10.6151
R1616 B.n527 B.n0 10.6151
R1617 B.n601 B.n1 10.6151
R1618 B.n601 B.n600 10.6151
R1619 B.n600 B.n599 10.6151
R1620 B.n599 B.n10 10.6151
R1621 B.n593 B.n10 10.6151
R1622 B.n593 B.n592 10.6151
R1623 B.n592 B.n591 10.6151
R1624 B.n591 B.n17 10.6151
R1625 B.n585 B.n17 10.6151
R1626 B.n585 B.n584 10.6151
R1627 B.n584 B.n583 10.6151
R1628 B.n583 B.n24 10.6151
R1629 B.n577 B.n24 10.6151
R1630 B.n577 B.n576 10.6151
R1631 B.n576 B.n575 10.6151
R1632 B.n575 B.n31 10.6151
R1633 B.n569 B.n31 10.6151
R1634 B.n569 B.n568 10.6151
R1635 B.n568 B.n567 10.6151
R1636 B.n567 B.n38 10.6151
R1637 B.n150 B.n149 9.36635
R1638 B.n172 B.n171 9.36635
R1639 B.n404 B.n317 9.36635
R1640 B.n381 B.n320 9.36635
R1641 B.n510 B.t2 4.55379
R1642 B.n589 B.t3 4.55379
R1643 B.n607 B.n0 2.81026
R1644 B.n607 B.n1 2.81026
R1645 B.n151 B.n150 1.24928
R1646 B.n171 B.n170 1.24928
R1647 B.n401 B.n317 1.24928
R1648 B.n384 B.n320 1.24928
R1649 VP.n0 VP.t1 248.404
R1650 VP.n0 VP.t2 248.315
R1651 VP.n2 VP.t0 229.797
R1652 VP.n3 VP.t3 229.797
R1653 VP.n4 VP.n3 80.6037
R1654 VP.n2 VP.n1 80.6037
R1655 VP.n1 VP.n0 71.0865
R1656 VP.n3 VP.n2 48.2005
R1657 VP.n4 VP.n1 0.380177
R1658 VP VP.n4 0.146778
R1659 VDD1 VDD1.n1 98.6036
R1660 VDD1 VDD1.n0 62.6722
R1661 VDD1.n0 VDD1.t2 2.14801
R1662 VDD1.n0 VDD1.t1 2.14801
R1663 VDD1.n1 VDD1.t3 2.14801
R1664 VDD1.n1 VDD1.t0 2.14801
C0 VDD2 VTAIL 4.93228f
C1 VTAIL VP 2.82923f
C2 VDD1 VN 0.14746f
C3 VDD2 VP 0.301183f
C4 VDD1 VTAIL 4.88786f
C5 VDD2 VDD1 0.672052f
C6 VDD1 VP 3.1662f
C7 VTAIL VN 2.81512f
C8 VDD2 VN 3.01284f
C9 VN VP 4.62299f
C10 VDD2 B 2.733505f
C11 VDD1 B 6.11981f
C12 VTAIL B 7.526012f
C13 VN B 8.199349f
C14 VP B 5.652375f
C15 VDD1.t2 B 0.198123f
C16 VDD1.t1 B 0.198123f
C17 VDD1.n0 B 1.73414f
C18 VDD1.t3 B 0.198123f
C19 VDD1.t0 B 0.198123f
C20 VDD1.n1 B 2.26875f
C21 VP.t2 B 1.29896f
C22 VP.t1 B 1.29916f
C23 VP.n0 B 1.93299f
C24 VP.n1 B 2.40258f
C25 VP.t0 B 1.25991f
C26 VP.n2 B 0.523595f
C27 VP.t3 B 1.25991f
C28 VP.n3 B 0.523595f
C29 VP.n4 B 0.053112f
C30 VTAIL.n0 B 0.021153f
C31 VTAIL.n1 B 0.016472f
C32 VTAIL.n2 B 0.008852f
C33 VTAIL.n3 B 0.020922f
C34 VTAIL.n4 B 0.009112f
C35 VTAIL.n5 B 0.016472f
C36 VTAIL.n6 B 0.009372f
C37 VTAIL.n7 B 0.020922f
C38 VTAIL.n8 B 0.009372f
C39 VTAIL.n9 B 0.016472f
C40 VTAIL.n10 B 0.008852f
C41 VTAIL.n11 B 0.020922f
C42 VTAIL.n12 B 0.009372f
C43 VTAIL.n13 B 0.627317f
C44 VTAIL.n14 B 0.008852f
C45 VTAIL.t7 B 0.035091f
C46 VTAIL.n15 B 0.101187f
C47 VTAIL.n16 B 0.01479f
C48 VTAIL.n17 B 0.015691f
C49 VTAIL.n18 B 0.020922f
C50 VTAIL.n19 B 0.009372f
C51 VTAIL.n20 B 0.008852f
C52 VTAIL.n21 B 0.016472f
C53 VTAIL.n22 B 0.016472f
C54 VTAIL.n23 B 0.008852f
C55 VTAIL.n24 B 0.009372f
C56 VTAIL.n25 B 0.020922f
C57 VTAIL.n26 B 0.020922f
C58 VTAIL.n27 B 0.009372f
C59 VTAIL.n28 B 0.008852f
C60 VTAIL.n29 B 0.016472f
C61 VTAIL.n30 B 0.016472f
C62 VTAIL.n31 B 0.008852f
C63 VTAIL.n32 B 0.008852f
C64 VTAIL.n33 B 0.009372f
C65 VTAIL.n34 B 0.020922f
C66 VTAIL.n35 B 0.020922f
C67 VTAIL.n36 B 0.020922f
C68 VTAIL.n37 B 0.009112f
C69 VTAIL.n38 B 0.008852f
C70 VTAIL.n39 B 0.016472f
C71 VTAIL.n40 B 0.016472f
C72 VTAIL.n41 B 0.008852f
C73 VTAIL.n42 B 0.009372f
C74 VTAIL.n43 B 0.020922f
C75 VTAIL.n44 B 0.041755f
C76 VTAIL.n45 B 0.009372f
C77 VTAIL.n46 B 0.008852f
C78 VTAIL.n47 B 0.037625f
C79 VTAIL.n48 B 0.022986f
C80 VTAIL.n49 B 0.075472f
C81 VTAIL.n50 B 0.021153f
C82 VTAIL.n51 B 0.016472f
C83 VTAIL.n52 B 0.008852f
C84 VTAIL.n53 B 0.020922f
C85 VTAIL.n54 B 0.009112f
C86 VTAIL.n55 B 0.016472f
C87 VTAIL.n56 B 0.009372f
C88 VTAIL.n57 B 0.020922f
C89 VTAIL.n58 B 0.009372f
C90 VTAIL.n59 B 0.016472f
C91 VTAIL.n60 B 0.008852f
C92 VTAIL.n61 B 0.020922f
C93 VTAIL.n62 B 0.009372f
C94 VTAIL.n63 B 0.627317f
C95 VTAIL.n64 B 0.008852f
C96 VTAIL.t1 B 0.035091f
C97 VTAIL.n65 B 0.101187f
C98 VTAIL.n66 B 0.01479f
C99 VTAIL.n67 B 0.015691f
C100 VTAIL.n68 B 0.020922f
C101 VTAIL.n69 B 0.009372f
C102 VTAIL.n70 B 0.008852f
C103 VTAIL.n71 B 0.016472f
C104 VTAIL.n72 B 0.016472f
C105 VTAIL.n73 B 0.008852f
C106 VTAIL.n74 B 0.009372f
C107 VTAIL.n75 B 0.020922f
C108 VTAIL.n76 B 0.020922f
C109 VTAIL.n77 B 0.009372f
C110 VTAIL.n78 B 0.008852f
C111 VTAIL.n79 B 0.016472f
C112 VTAIL.n80 B 0.016472f
C113 VTAIL.n81 B 0.008852f
C114 VTAIL.n82 B 0.008852f
C115 VTAIL.n83 B 0.009372f
C116 VTAIL.n84 B 0.020922f
C117 VTAIL.n85 B 0.020922f
C118 VTAIL.n86 B 0.020922f
C119 VTAIL.n87 B 0.009112f
C120 VTAIL.n88 B 0.008852f
C121 VTAIL.n89 B 0.016472f
C122 VTAIL.n90 B 0.016472f
C123 VTAIL.n91 B 0.008852f
C124 VTAIL.n92 B 0.009372f
C125 VTAIL.n93 B 0.020922f
C126 VTAIL.n94 B 0.041755f
C127 VTAIL.n95 B 0.009372f
C128 VTAIL.n96 B 0.008852f
C129 VTAIL.n97 B 0.037625f
C130 VTAIL.n98 B 0.022986f
C131 VTAIL.n99 B 0.106014f
C132 VTAIL.n100 B 0.021153f
C133 VTAIL.n101 B 0.016472f
C134 VTAIL.n102 B 0.008852f
C135 VTAIL.n103 B 0.020922f
C136 VTAIL.n104 B 0.009112f
C137 VTAIL.n105 B 0.016472f
C138 VTAIL.n106 B 0.009372f
C139 VTAIL.n107 B 0.020922f
C140 VTAIL.n108 B 0.009372f
C141 VTAIL.n109 B 0.016472f
C142 VTAIL.n110 B 0.008852f
C143 VTAIL.n111 B 0.020922f
C144 VTAIL.n112 B 0.009372f
C145 VTAIL.n113 B 0.627317f
C146 VTAIL.n114 B 0.008852f
C147 VTAIL.t2 B 0.035091f
C148 VTAIL.n115 B 0.101187f
C149 VTAIL.n116 B 0.01479f
C150 VTAIL.n117 B 0.015691f
C151 VTAIL.n118 B 0.020922f
C152 VTAIL.n119 B 0.009372f
C153 VTAIL.n120 B 0.008852f
C154 VTAIL.n121 B 0.016472f
C155 VTAIL.n122 B 0.016472f
C156 VTAIL.n123 B 0.008852f
C157 VTAIL.n124 B 0.009372f
C158 VTAIL.n125 B 0.020922f
C159 VTAIL.n126 B 0.020922f
C160 VTAIL.n127 B 0.009372f
C161 VTAIL.n128 B 0.008852f
C162 VTAIL.n129 B 0.016472f
C163 VTAIL.n130 B 0.016472f
C164 VTAIL.n131 B 0.008852f
C165 VTAIL.n132 B 0.008852f
C166 VTAIL.n133 B 0.009372f
C167 VTAIL.n134 B 0.020922f
C168 VTAIL.n135 B 0.020922f
C169 VTAIL.n136 B 0.020922f
C170 VTAIL.n137 B 0.009112f
C171 VTAIL.n138 B 0.008852f
C172 VTAIL.n139 B 0.016472f
C173 VTAIL.n140 B 0.016472f
C174 VTAIL.n141 B 0.008852f
C175 VTAIL.n142 B 0.009372f
C176 VTAIL.n143 B 0.020922f
C177 VTAIL.n144 B 0.041755f
C178 VTAIL.n145 B 0.009372f
C179 VTAIL.n146 B 0.008852f
C180 VTAIL.n147 B 0.037625f
C181 VTAIL.n148 B 0.022986f
C182 VTAIL.n149 B 0.793974f
C183 VTAIL.n150 B 0.021153f
C184 VTAIL.n151 B 0.016472f
C185 VTAIL.n152 B 0.008852f
C186 VTAIL.n153 B 0.020922f
C187 VTAIL.n154 B 0.009112f
C188 VTAIL.n155 B 0.016472f
C189 VTAIL.n156 B 0.009112f
C190 VTAIL.n157 B 0.008852f
C191 VTAIL.n158 B 0.020922f
C192 VTAIL.n159 B 0.020922f
C193 VTAIL.n160 B 0.009372f
C194 VTAIL.n161 B 0.016472f
C195 VTAIL.n162 B 0.008852f
C196 VTAIL.n163 B 0.020922f
C197 VTAIL.n164 B 0.009372f
C198 VTAIL.n165 B 0.627317f
C199 VTAIL.n166 B 0.008852f
C200 VTAIL.t4 B 0.035091f
C201 VTAIL.n167 B 0.101187f
C202 VTAIL.n168 B 0.01479f
C203 VTAIL.n169 B 0.015691f
C204 VTAIL.n170 B 0.020922f
C205 VTAIL.n171 B 0.009372f
C206 VTAIL.n172 B 0.008852f
C207 VTAIL.n173 B 0.016472f
C208 VTAIL.n174 B 0.016472f
C209 VTAIL.n175 B 0.008852f
C210 VTAIL.n176 B 0.009372f
C211 VTAIL.n177 B 0.020922f
C212 VTAIL.n178 B 0.020922f
C213 VTAIL.n179 B 0.009372f
C214 VTAIL.n180 B 0.008852f
C215 VTAIL.n181 B 0.016472f
C216 VTAIL.n182 B 0.016472f
C217 VTAIL.n183 B 0.008852f
C218 VTAIL.n184 B 0.009372f
C219 VTAIL.n185 B 0.020922f
C220 VTAIL.n186 B 0.020922f
C221 VTAIL.n187 B 0.009372f
C222 VTAIL.n188 B 0.008852f
C223 VTAIL.n189 B 0.016472f
C224 VTAIL.n190 B 0.016472f
C225 VTAIL.n191 B 0.008852f
C226 VTAIL.n192 B 0.009372f
C227 VTAIL.n193 B 0.020922f
C228 VTAIL.n194 B 0.041755f
C229 VTAIL.n195 B 0.009372f
C230 VTAIL.n196 B 0.008852f
C231 VTAIL.n197 B 0.037625f
C232 VTAIL.n198 B 0.022986f
C233 VTAIL.n199 B 0.793974f
C234 VTAIL.n200 B 0.021153f
C235 VTAIL.n201 B 0.016472f
C236 VTAIL.n202 B 0.008852f
C237 VTAIL.n203 B 0.020922f
C238 VTAIL.n204 B 0.009112f
C239 VTAIL.n205 B 0.016472f
C240 VTAIL.n206 B 0.009112f
C241 VTAIL.n207 B 0.008852f
C242 VTAIL.n208 B 0.020922f
C243 VTAIL.n209 B 0.020922f
C244 VTAIL.n210 B 0.009372f
C245 VTAIL.n211 B 0.016472f
C246 VTAIL.n212 B 0.008852f
C247 VTAIL.n213 B 0.020922f
C248 VTAIL.n214 B 0.009372f
C249 VTAIL.n215 B 0.627317f
C250 VTAIL.n216 B 0.008852f
C251 VTAIL.t6 B 0.035091f
C252 VTAIL.n217 B 0.101187f
C253 VTAIL.n218 B 0.01479f
C254 VTAIL.n219 B 0.015691f
C255 VTAIL.n220 B 0.020922f
C256 VTAIL.n221 B 0.009372f
C257 VTAIL.n222 B 0.008852f
C258 VTAIL.n223 B 0.016472f
C259 VTAIL.n224 B 0.016472f
C260 VTAIL.n225 B 0.008852f
C261 VTAIL.n226 B 0.009372f
C262 VTAIL.n227 B 0.020922f
C263 VTAIL.n228 B 0.020922f
C264 VTAIL.n229 B 0.009372f
C265 VTAIL.n230 B 0.008852f
C266 VTAIL.n231 B 0.016472f
C267 VTAIL.n232 B 0.016472f
C268 VTAIL.n233 B 0.008852f
C269 VTAIL.n234 B 0.009372f
C270 VTAIL.n235 B 0.020922f
C271 VTAIL.n236 B 0.020922f
C272 VTAIL.n237 B 0.009372f
C273 VTAIL.n238 B 0.008852f
C274 VTAIL.n239 B 0.016472f
C275 VTAIL.n240 B 0.016472f
C276 VTAIL.n241 B 0.008852f
C277 VTAIL.n242 B 0.009372f
C278 VTAIL.n243 B 0.020922f
C279 VTAIL.n244 B 0.041755f
C280 VTAIL.n245 B 0.009372f
C281 VTAIL.n246 B 0.008852f
C282 VTAIL.n247 B 0.037625f
C283 VTAIL.n248 B 0.022986f
C284 VTAIL.n249 B 0.106014f
C285 VTAIL.n250 B 0.021153f
C286 VTAIL.n251 B 0.016472f
C287 VTAIL.n252 B 0.008852f
C288 VTAIL.n253 B 0.020922f
C289 VTAIL.n254 B 0.009112f
C290 VTAIL.n255 B 0.016472f
C291 VTAIL.n256 B 0.009112f
C292 VTAIL.n257 B 0.008852f
C293 VTAIL.n258 B 0.020922f
C294 VTAIL.n259 B 0.020922f
C295 VTAIL.n260 B 0.009372f
C296 VTAIL.n261 B 0.016472f
C297 VTAIL.n262 B 0.008852f
C298 VTAIL.n263 B 0.020922f
C299 VTAIL.n264 B 0.009372f
C300 VTAIL.n265 B 0.627317f
C301 VTAIL.n266 B 0.008852f
C302 VTAIL.t0 B 0.035091f
C303 VTAIL.n267 B 0.101187f
C304 VTAIL.n268 B 0.01479f
C305 VTAIL.n269 B 0.015691f
C306 VTAIL.n270 B 0.020922f
C307 VTAIL.n271 B 0.009372f
C308 VTAIL.n272 B 0.008852f
C309 VTAIL.n273 B 0.016472f
C310 VTAIL.n274 B 0.016472f
C311 VTAIL.n275 B 0.008852f
C312 VTAIL.n276 B 0.009372f
C313 VTAIL.n277 B 0.020922f
C314 VTAIL.n278 B 0.020922f
C315 VTAIL.n279 B 0.009372f
C316 VTAIL.n280 B 0.008852f
C317 VTAIL.n281 B 0.016472f
C318 VTAIL.n282 B 0.016472f
C319 VTAIL.n283 B 0.008852f
C320 VTAIL.n284 B 0.009372f
C321 VTAIL.n285 B 0.020922f
C322 VTAIL.n286 B 0.020922f
C323 VTAIL.n287 B 0.009372f
C324 VTAIL.n288 B 0.008852f
C325 VTAIL.n289 B 0.016472f
C326 VTAIL.n290 B 0.016472f
C327 VTAIL.n291 B 0.008852f
C328 VTAIL.n292 B 0.009372f
C329 VTAIL.n293 B 0.020922f
C330 VTAIL.n294 B 0.041755f
C331 VTAIL.n295 B 0.009372f
C332 VTAIL.n296 B 0.008852f
C333 VTAIL.n297 B 0.037625f
C334 VTAIL.n298 B 0.022986f
C335 VTAIL.n299 B 0.106014f
C336 VTAIL.n300 B 0.021153f
C337 VTAIL.n301 B 0.016472f
C338 VTAIL.n302 B 0.008852f
C339 VTAIL.n303 B 0.020922f
C340 VTAIL.n304 B 0.009112f
C341 VTAIL.n305 B 0.016472f
C342 VTAIL.n306 B 0.009112f
C343 VTAIL.n307 B 0.008852f
C344 VTAIL.n308 B 0.020922f
C345 VTAIL.n309 B 0.020922f
C346 VTAIL.n310 B 0.009372f
C347 VTAIL.n311 B 0.016472f
C348 VTAIL.n312 B 0.008852f
C349 VTAIL.n313 B 0.020922f
C350 VTAIL.n314 B 0.009372f
C351 VTAIL.n315 B 0.627317f
C352 VTAIL.n316 B 0.008852f
C353 VTAIL.t3 B 0.035091f
C354 VTAIL.n317 B 0.101187f
C355 VTAIL.n318 B 0.01479f
C356 VTAIL.n319 B 0.015691f
C357 VTAIL.n320 B 0.020922f
C358 VTAIL.n321 B 0.009372f
C359 VTAIL.n322 B 0.008852f
C360 VTAIL.n323 B 0.016472f
C361 VTAIL.n324 B 0.016472f
C362 VTAIL.n325 B 0.008852f
C363 VTAIL.n326 B 0.009372f
C364 VTAIL.n327 B 0.020922f
C365 VTAIL.n328 B 0.020922f
C366 VTAIL.n329 B 0.009372f
C367 VTAIL.n330 B 0.008852f
C368 VTAIL.n331 B 0.016472f
C369 VTAIL.n332 B 0.016472f
C370 VTAIL.n333 B 0.008852f
C371 VTAIL.n334 B 0.009372f
C372 VTAIL.n335 B 0.020922f
C373 VTAIL.n336 B 0.020922f
C374 VTAIL.n337 B 0.009372f
C375 VTAIL.n338 B 0.008852f
C376 VTAIL.n339 B 0.016472f
C377 VTAIL.n340 B 0.016472f
C378 VTAIL.n341 B 0.008852f
C379 VTAIL.n342 B 0.009372f
C380 VTAIL.n343 B 0.020922f
C381 VTAIL.n344 B 0.041755f
C382 VTAIL.n345 B 0.009372f
C383 VTAIL.n346 B 0.008852f
C384 VTAIL.n347 B 0.037625f
C385 VTAIL.n348 B 0.022986f
C386 VTAIL.n349 B 0.793974f
C387 VTAIL.n350 B 0.021153f
C388 VTAIL.n351 B 0.016472f
C389 VTAIL.n352 B 0.008852f
C390 VTAIL.n353 B 0.020922f
C391 VTAIL.n354 B 0.009112f
C392 VTAIL.n355 B 0.016472f
C393 VTAIL.n356 B 0.009372f
C394 VTAIL.n357 B 0.020922f
C395 VTAIL.n358 B 0.009372f
C396 VTAIL.n359 B 0.016472f
C397 VTAIL.n360 B 0.008852f
C398 VTAIL.n361 B 0.020922f
C399 VTAIL.n362 B 0.009372f
C400 VTAIL.n363 B 0.627317f
C401 VTAIL.n364 B 0.008852f
C402 VTAIL.t5 B 0.035091f
C403 VTAIL.n365 B 0.101187f
C404 VTAIL.n366 B 0.01479f
C405 VTAIL.n367 B 0.015691f
C406 VTAIL.n368 B 0.020922f
C407 VTAIL.n369 B 0.009372f
C408 VTAIL.n370 B 0.008852f
C409 VTAIL.n371 B 0.016472f
C410 VTAIL.n372 B 0.016472f
C411 VTAIL.n373 B 0.008852f
C412 VTAIL.n374 B 0.009372f
C413 VTAIL.n375 B 0.020922f
C414 VTAIL.n376 B 0.020922f
C415 VTAIL.n377 B 0.009372f
C416 VTAIL.n378 B 0.008852f
C417 VTAIL.n379 B 0.016472f
C418 VTAIL.n380 B 0.016472f
C419 VTAIL.n381 B 0.008852f
C420 VTAIL.n382 B 0.008852f
C421 VTAIL.n383 B 0.009372f
C422 VTAIL.n384 B 0.020922f
C423 VTAIL.n385 B 0.020922f
C424 VTAIL.n386 B 0.020922f
C425 VTAIL.n387 B 0.009112f
C426 VTAIL.n388 B 0.008852f
C427 VTAIL.n389 B 0.016472f
C428 VTAIL.n390 B 0.016472f
C429 VTAIL.n391 B 0.008852f
C430 VTAIL.n392 B 0.009372f
C431 VTAIL.n393 B 0.020922f
C432 VTAIL.n394 B 0.041755f
C433 VTAIL.n395 B 0.009372f
C434 VTAIL.n396 B 0.008852f
C435 VTAIL.n397 B 0.037625f
C436 VTAIL.n398 B 0.022986f
C437 VTAIL.n399 B 0.757255f
C438 VDD2.t0 B 0.195657f
C439 VDD2.t3 B 0.195657f
C440 VDD2.n0 B 2.21588f
C441 VDD2.t2 B 0.195657f
C442 VDD2.t1 B 0.195657f
C443 VDD2.n1 B 1.71224f
C444 VDD2.n2 B 3.07382f
C445 VN.t0 B 1.26763f
C446 VN.t2 B 1.26743f
C447 VN.n0 B 0.946512f
C448 VN.t1 B 1.26763f
C449 VN.t3 B 1.26743f
C450 VN.n1 B 1.90201f
.ends

