* NGSPICE file created from diff_pair_sample_0210.ext - technology: sky130A

.subckt diff_pair_sample_0210 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.21945 pd=1.66 as=0.5187 ps=3.44 w=1.33 l=3.12
X1 VTAIL.t5 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5187 pd=3.44 as=0.21945 ps=1.66 w=1.33 l=3.12
X2 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5187 pd=3.44 as=0 ps=0 w=1.33 l=3.12
X3 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5187 pd=3.44 as=0 ps=0 w=1.33 l=3.12
X4 VDD2.t3 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.21945 pd=1.66 as=0.5187 ps=3.44 w=1.33 l=3.12
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5187 pd=3.44 as=0 ps=0 w=1.33 l=3.12
X6 VDD2.t2 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.21945 pd=1.66 as=0.5187 ps=3.44 w=1.33 l=3.12
X7 VTAIL.t1 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.5187 pd=3.44 as=0.21945 ps=1.66 w=1.33 l=3.12
X8 VDD1.t1 VP.t2 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.21945 pd=1.66 as=0.5187 ps=3.44 w=1.33 l=3.12
X9 VTAIL.t2 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5187 pd=3.44 as=0.21945 ps=1.66 w=1.33 l=3.12
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=0.5187 pd=3.44 as=0 ps=0 w=1.33 l=3.12
X11 VTAIL.t7 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.5187 pd=3.44 as=0.21945 ps=1.66 w=1.33 l=3.12
R0 VP.n15 VP.n14 161.3
R1 VP.n13 VP.n1 161.3
R2 VP.n12 VP.n11 161.3
R3 VP.n10 VP.n2 161.3
R4 VP.n9 VP.n8 161.3
R5 VP.n7 VP.n3 161.3
R6 VP.n6 VP.n5 66.8237
R7 VP.n16 VP.n0 66.8237
R8 VP.n12 VP.n2 56.5193
R9 VP.n4 VP.t3 44.7874
R10 VP.n4 VP.t0 43.7682
R11 VP.n5 VP.n4 42.7479
R12 VP.n8 VP.n7 24.4675
R13 VP.n8 VP.n2 24.4675
R14 VP.n13 VP.n12 24.4675
R15 VP.n14 VP.n13 24.4675
R16 VP.n7 VP.n6 23.2442
R17 VP.n14 VP.n0 23.2442
R18 VP.n6 VP.t1 10.2739
R19 VP.n0 VP.t2 10.2739
R20 VP.n5 VP.n3 0.354971
R21 VP.n16 VP.n15 0.354971
R22 VP VP.n16 0.26696
R23 VP.n9 VP.n3 0.189894
R24 VP.n10 VP.n9 0.189894
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n1 0.189894
R27 VP.n15 VP.n1 0.189894
R28 VTAIL.n7 VTAIL.t3 156.877
R29 VTAIL.n0 VTAIL.t2 156.877
R30 VTAIL.n1 VTAIL.t6 156.877
R31 VTAIL.n2 VTAIL.t5 156.877
R32 VTAIL.n6 VTAIL.t4 156.877
R33 VTAIL.n5 VTAIL.t7 156.877
R34 VTAIL.n4 VTAIL.t0 156.877
R35 VTAIL.n3 VTAIL.t1 156.877
R36 VTAIL.n7 VTAIL.n6 16.4876
R37 VTAIL.n3 VTAIL.n2 16.4876
R38 VTAIL.n4 VTAIL.n3 2.97464
R39 VTAIL.n6 VTAIL.n5 2.97464
R40 VTAIL.n2 VTAIL.n1 2.97464
R41 VTAIL VTAIL.n0 1.54576
R42 VTAIL VTAIL.n7 1.42938
R43 VTAIL.n5 VTAIL.n4 0.470328
R44 VTAIL.n1 VTAIL.n0 0.470328
R45 VDD1 VDD1.n1 181.708
R46 VDD1 VDD1.n0 147.457
R47 VDD1.n0 VDD1.t0 14.8877
R48 VDD1.n0 VDD1.t3 14.8877
R49 VDD1.n1 VDD1.t2 14.8877
R50 VDD1.n1 VDD1.t1 14.8877
R51 B.n414 B.n413 585
R52 B.n415 B.n93 585
R53 B.n417 B.n416 585
R54 B.n419 B.n92 585
R55 B.n422 B.n421 585
R56 B.n423 B.n91 585
R57 B.n425 B.n424 585
R58 B.n427 B.n90 585
R59 B.n429 B.n428 585
R60 B.n431 B.n430 585
R61 B.n434 B.n433 585
R62 B.n435 B.n85 585
R63 B.n437 B.n436 585
R64 B.n439 B.n84 585
R65 B.n442 B.n441 585
R66 B.n443 B.n83 585
R67 B.n445 B.n444 585
R68 B.n447 B.n82 585
R69 B.n449 B.n448 585
R70 B.n451 B.n450 585
R71 B.n454 B.n453 585
R72 B.n455 B.n77 585
R73 B.n457 B.n456 585
R74 B.n459 B.n76 585
R75 B.n462 B.n461 585
R76 B.n463 B.n75 585
R77 B.n465 B.n464 585
R78 B.n467 B.n74 585
R79 B.n470 B.n469 585
R80 B.n471 B.n73 585
R81 B.n411 B.n71 585
R82 B.n474 B.n71 585
R83 B.n410 B.n70 585
R84 B.n475 B.n70 585
R85 B.n409 B.n69 585
R86 B.n476 B.n69 585
R87 B.n408 B.n407 585
R88 B.n407 B.n65 585
R89 B.n406 B.n64 585
R90 B.n482 B.n64 585
R91 B.n405 B.n63 585
R92 B.n483 B.n63 585
R93 B.n404 B.n62 585
R94 B.n484 B.n62 585
R95 B.n403 B.n402 585
R96 B.n402 B.n58 585
R97 B.n401 B.n57 585
R98 B.n490 B.n57 585
R99 B.n400 B.n56 585
R100 B.n491 B.n56 585
R101 B.n399 B.n55 585
R102 B.n492 B.n55 585
R103 B.n398 B.n397 585
R104 B.n397 B.n51 585
R105 B.n396 B.n50 585
R106 B.n498 B.n50 585
R107 B.n395 B.n49 585
R108 B.n499 B.n49 585
R109 B.n394 B.n48 585
R110 B.n500 B.n48 585
R111 B.n393 B.n392 585
R112 B.n392 B.n44 585
R113 B.n391 B.n43 585
R114 B.n506 B.n43 585
R115 B.n390 B.n42 585
R116 B.n507 B.n42 585
R117 B.n389 B.n41 585
R118 B.n508 B.n41 585
R119 B.n388 B.n387 585
R120 B.n387 B.n37 585
R121 B.n386 B.n36 585
R122 B.n514 B.n36 585
R123 B.n385 B.n35 585
R124 B.n515 B.n35 585
R125 B.n384 B.n34 585
R126 B.n516 B.n34 585
R127 B.n383 B.n382 585
R128 B.n382 B.n30 585
R129 B.n381 B.n29 585
R130 B.n522 B.n29 585
R131 B.n380 B.n28 585
R132 B.n523 B.n28 585
R133 B.n379 B.n27 585
R134 B.n524 B.n27 585
R135 B.n378 B.n377 585
R136 B.n377 B.n23 585
R137 B.n376 B.n22 585
R138 B.n530 B.n22 585
R139 B.n375 B.n21 585
R140 B.n531 B.n21 585
R141 B.n374 B.n20 585
R142 B.n532 B.n20 585
R143 B.n373 B.n372 585
R144 B.n372 B.n19 585
R145 B.n371 B.n15 585
R146 B.n538 B.n15 585
R147 B.n370 B.n14 585
R148 B.n539 B.n14 585
R149 B.n369 B.n13 585
R150 B.n540 B.n13 585
R151 B.n368 B.n367 585
R152 B.n367 B.n12 585
R153 B.n366 B.n365 585
R154 B.n366 B.n8 585
R155 B.n364 B.n7 585
R156 B.n547 B.n7 585
R157 B.n363 B.n6 585
R158 B.n548 B.n6 585
R159 B.n362 B.n5 585
R160 B.n549 B.n5 585
R161 B.n361 B.n360 585
R162 B.n360 B.n4 585
R163 B.n359 B.n94 585
R164 B.n359 B.n358 585
R165 B.n349 B.n95 585
R166 B.n96 B.n95 585
R167 B.n351 B.n350 585
R168 B.n352 B.n351 585
R169 B.n348 B.n101 585
R170 B.n101 B.n100 585
R171 B.n347 B.n346 585
R172 B.n346 B.n345 585
R173 B.n103 B.n102 585
R174 B.n338 B.n103 585
R175 B.n337 B.n336 585
R176 B.n339 B.n337 585
R177 B.n335 B.n108 585
R178 B.n108 B.n107 585
R179 B.n334 B.n333 585
R180 B.n333 B.n332 585
R181 B.n110 B.n109 585
R182 B.n111 B.n110 585
R183 B.n325 B.n324 585
R184 B.n326 B.n325 585
R185 B.n323 B.n116 585
R186 B.n116 B.n115 585
R187 B.n322 B.n321 585
R188 B.n321 B.n320 585
R189 B.n118 B.n117 585
R190 B.n119 B.n118 585
R191 B.n313 B.n312 585
R192 B.n314 B.n313 585
R193 B.n311 B.n123 585
R194 B.n127 B.n123 585
R195 B.n310 B.n309 585
R196 B.n309 B.n308 585
R197 B.n125 B.n124 585
R198 B.n126 B.n125 585
R199 B.n301 B.n300 585
R200 B.n302 B.n301 585
R201 B.n299 B.n132 585
R202 B.n132 B.n131 585
R203 B.n298 B.n297 585
R204 B.n297 B.n296 585
R205 B.n134 B.n133 585
R206 B.n135 B.n134 585
R207 B.n289 B.n288 585
R208 B.n290 B.n289 585
R209 B.n287 B.n140 585
R210 B.n140 B.n139 585
R211 B.n286 B.n285 585
R212 B.n285 B.n284 585
R213 B.n142 B.n141 585
R214 B.n143 B.n142 585
R215 B.n277 B.n276 585
R216 B.n278 B.n277 585
R217 B.n275 B.n148 585
R218 B.n148 B.n147 585
R219 B.n274 B.n273 585
R220 B.n273 B.n272 585
R221 B.n150 B.n149 585
R222 B.n151 B.n150 585
R223 B.n265 B.n264 585
R224 B.n266 B.n265 585
R225 B.n263 B.n156 585
R226 B.n156 B.n155 585
R227 B.n262 B.n261 585
R228 B.n261 B.n260 585
R229 B.n158 B.n157 585
R230 B.n159 B.n158 585
R231 B.n253 B.n252 585
R232 B.n254 B.n253 585
R233 B.n251 B.n164 585
R234 B.n164 B.n163 585
R235 B.n250 B.n249 585
R236 B.n249 B.n248 585
R237 B.n245 B.n168 585
R238 B.n244 B.n243 585
R239 B.n241 B.n169 585
R240 B.n241 B.n167 585
R241 B.n240 B.n239 585
R242 B.n238 B.n237 585
R243 B.n236 B.n171 585
R244 B.n234 B.n233 585
R245 B.n232 B.n172 585
R246 B.n231 B.n230 585
R247 B.n228 B.n173 585
R248 B.n226 B.n225 585
R249 B.n224 B.n174 585
R250 B.n223 B.n222 585
R251 B.n220 B.n178 585
R252 B.n218 B.n217 585
R253 B.n216 B.n179 585
R254 B.n215 B.n214 585
R255 B.n212 B.n180 585
R256 B.n210 B.n209 585
R257 B.n208 B.n181 585
R258 B.n206 B.n205 585
R259 B.n203 B.n184 585
R260 B.n201 B.n200 585
R261 B.n199 B.n185 585
R262 B.n198 B.n197 585
R263 B.n195 B.n186 585
R264 B.n193 B.n192 585
R265 B.n191 B.n187 585
R266 B.n190 B.n189 585
R267 B.n166 B.n165 585
R268 B.n167 B.n166 585
R269 B.n247 B.n246 585
R270 B.n248 B.n247 585
R271 B.n162 B.n161 585
R272 B.n163 B.n162 585
R273 B.n256 B.n255 585
R274 B.n255 B.n254 585
R275 B.n257 B.n160 585
R276 B.n160 B.n159 585
R277 B.n259 B.n258 585
R278 B.n260 B.n259 585
R279 B.n154 B.n153 585
R280 B.n155 B.n154 585
R281 B.n268 B.n267 585
R282 B.n267 B.n266 585
R283 B.n269 B.n152 585
R284 B.n152 B.n151 585
R285 B.n271 B.n270 585
R286 B.n272 B.n271 585
R287 B.n146 B.n145 585
R288 B.n147 B.n146 585
R289 B.n280 B.n279 585
R290 B.n279 B.n278 585
R291 B.n281 B.n144 585
R292 B.n144 B.n143 585
R293 B.n283 B.n282 585
R294 B.n284 B.n283 585
R295 B.n138 B.n137 585
R296 B.n139 B.n138 585
R297 B.n292 B.n291 585
R298 B.n291 B.n290 585
R299 B.n293 B.n136 585
R300 B.n136 B.n135 585
R301 B.n295 B.n294 585
R302 B.n296 B.n295 585
R303 B.n130 B.n129 585
R304 B.n131 B.n130 585
R305 B.n304 B.n303 585
R306 B.n303 B.n302 585
R307 B.n305 B.n128 585
R308 B.n128 B.n126 585
R309 B.n307 B.n306 585
R310 B.n308 B.n307 585
R311 B.n122 B.n121 585
R312 B.n127 B.n122 585
R313 B.n316 B.n315 585
R314 B.n315 B.n314 585
R315 B.n317 B.n120 585
R316 B.n120 B.n119 585
R317 B.n319 B.n318 585
R318 B.n320 B.n319 585
R319 B.n114 B.n113 585
R320 B.n115 B.n114 585
R321 B.n328 B.n327 585
R322 B.n327 B.n326 585
R323 B.n329 B.n112 585
R324 B.n112 B.n111 585
R325 B.n331 B.n330 585
R326 B.n332 B.n331 585
R327 B.n106 B.n105 585
R328 B.n107 B.n106 585
R329 B.n341 B.n340 585
R330 B.n340 B.n339 585
R331 B.n342 B.n104 585
R332 B.n338 B.n104 585
R333 B.n344 B.n343 585
R334 B.n345 B.n344 585
R335 B.n99 B.n98 585
R336 B.n100 B.n99 585
R337 B.n354 B.n353 585
R338 B.n353 B.n352 585
R339 B.n355 B.n97 585
R340 B.n97 B.n96 585
R341 B.n357 B.n356 585
R342 B.n358 B.n357 585
R343 B.n3 B.n0 585
R344 B.n4 B.n3 585
R345 B.n546 B.n1 585
R346 B.n547 B.n546 585
R347 B.n545 B.n544 585
R348 B.n545 B.n8 585
R349 B.n543 B.n9 585
R350 B.n12 B.n9 585
R351 B.n542 B.n541 585
R352 B.n541 B.n540 585
R353 B.n11 B.n10 585
R354 B.n539 B.n11 585
R355 B.n537 B.n536 585
R356 B.n538 B.n537 585
R357 B.n535 B.n16 585
R358 B.n19 B.n16 585
R359 B.n534 B.n533 585
R360 B.n533 B.n532 585
R361 B.n18 B.n17 585
R362 B.n531 B.n18 585
R363 B.n529 B.n528 585
R364 B.n530 B.n529 585
R365 B.n527 B.n24 585
R366 B.n24 B.n23 585
R367 B.n526 B.n525 585
R368 B.n525 B.n524 585
R369 B.n26 B.n25 585
R370 B.n523 B.n26 585
R371 B.n521 B.n520 585
R372 B.n522 B.n521 585
R373 B.n519 B.n31 585
R374 B.n31 B.n30 585
R375 B.n518 B.n517 585
R376 B.n517 B.n516 585
R377 B.n33 B.n32 585
R378 B.n515 B.n33 585
R379 B.n513 B.n512 585
R380 B.n514 B.n513 585
R381 B.n511 B.n38 585
R382 B.n38 B.n37 585
R383 B.n510 B.n509 585
R384 B.n509 B.n508 585
R385 B.n40 B.n39 585
R386 B.n507 B.n40 585
R387 B.n505 B.n504 585
R388 B.n506 B.n505 585
R389 B.n503 B.n45 585
R390 B.n45 B.n44 585
R391 B.n502 B.n501 585
R392 B.n501 B.n500 585
R393 B.n47 B.n46 585
R394 B.n499 B.n47 585
R395 B.n497 B.n496 585
R396 B.n498 B.n497 585
R397 B.n495 B.n52 585
R398 B.n52 B.n51 585
R399 B.n494 B.n493 585
R400 B.n493 B.n492 585
R401 B.n54 B.n53 585
R402 B.n491 B.n54 585
R403 B.n489 B.n488 585
R404 B.n490 B.n489 585
R405 B.n487 B.n59 585
R406 B.n59 B.n58 585
R407 B.n486 B.n485 585
R408 B.n485 B.n484 585
R409 B.n61 B.n60 585
R410 B.n483 B.n61 585
R411 B.n481 B.n480 585
R412 B.n482 B.n481 585
R413 B.n479 B.n66 585
R414 B.n66 B.n65 585
R415 B.n478 B.n477 585
R416 B.n477 B.n476 585
R417 B.n68 B.n67 585
R418 B.n475 B.n68 585
R419 B.n473 B.n472 585
R420 B.n474 B.n473 585
R421 B.n550 B.n549 585
R422 B.n548 B.n2 585
R423 B.n473 B.n73 511.721
R424 B.n413 B.n71 511.721
R425 B.n249 B.n166 511.721
R426 B.n247 B.n168 511.721
R427 B.n412 B.n72 256.663
R428 B.n418 B.n72 256.663
R429 B.n420 B.n72 256.663
R430 B.n426 B.n72 256.663
R431 B.n89 B.n72 256.663
R432 B.n432 B.n72 256.663
R433 B.n438 B.n72 256.663
R434 B.n440 B.n72 256.663
R435 B.n446 B.n72 256.663
R436 B.n81 B.n72 256.663
R437 B.n452 B.n72 256.663
R438 B.n458 B.n72 256.663
R439 B.n460 B.n72 256.663
R440 B.n466 B.n72 256.663
R441 B.n468 B.n72 256.663
R442 B.n242 B.n167 256.663
R443 B.n170 B.n167 256.663
R444 B.n235 B.n167 256.663
R445 B.n229 B.n167 256.663
R446 B.n227 B.n167 256.663
R447 B.n221 B.n167 256.663
R448 B.n219 B.n167 256.663
R449 B.n213 B.n167 256.663
R450 B.n211 B.n167 256.663
R451 B.n204 B.n167 256.663
R452 B.n202 B.n167 256.663
R453 B.n196 B.n167 256.663
R454 B.n194 B.n167 256.663
R455 B.n188 B.n167 256.663
R456 B.n552 B.n551 256.663
R457 B.n78 B.t13 217.669
R458 B.n86 B.t6 217.669
R459 B.n182 B.t17 217.669
R460 B.n175 B.t11 217.669
R461 B.n248 B.n167 211.506
R462 B.n474 B.n72 211.506
R463 B.n78 B.t12 209.32
R464 B.n86 B.t4 209.32
R465 B.n182 B.t15 209.32
R466 B.n175 B.t8 209.32
R467 B.n469 B.n467 163.367
R468 B.n465 B.n75 163.367
R469 B.n461 B.n459 163.367
R470 B.n457 B.n77 163.367
R471 B.n453 B.n451 163.367
R472 B.n448 B.n447 163.367
R473 B.n445 B.n83 163.367
R474 B.n441 B.n439 163.367
R475 B.n437 B.n85 163.367
R476 B.n433 B.n431 163.367
R477 B.n428 B.n427 163.367
R478 B.n425 B.n91 163.367
R479 B.n421 B.n419 163.367
R480 B.n417 B.n93 163.367
R481 B.n249 B.n164 163.367
R482 B.n253 B.n164 163.367
R483 B.n253 B.n158 163.367
R484 B.n261 B.n158 163.367
R485 B.n261 B.n156 163.367
R486 B.n265 B.n156 163.367
R487 B.n265 B.n150 163.367
R488 B.n273 B.n150 163.367
R489 B.n273 B.n148 163.367
R490 B.n277 B.n148 163.367
R491 B.n277 B.n142 163.367
R492 B.n285 B.n142 163.367
R493 B.n285 B.n140 163.367
R494 B.n289 B.n140 163.367
R495 B.n289 B.n134 163.367
R496 B.n297 B.n134 163.367
R497 B.n297 B.n132 163.367
R498 B.n301 B.n132 163.367
R499 B.n301 B.n125 163.367
R500 B.n309 B.n125 163.367
R501 B.n309 B.n123 163.367
R502 B.n313 B.n123 163.367
R503 B.n313 B.n118 163.367
R504 B.n321 B.n118 163.367
R505 B.n321 B.n116 163.367
R506 B.n325 B.n116 163.367
R507 B.n325 B.n110 163.367
R508 B.n333 B.n110 163.367
R509 B.n333 B.n108 163.367
R510 B.n337 B.n108 163.367
R511 B.n337 B.n103 163.367
R512 B.n346 B.n103 163.367
R513 B.n346 B.n101 163.367
R514 B.n351 B.n101 163.367
R515 B.n351 B.n95 163.367
R516 B.n359 B.n95 163.367
R517 B.n360 B.n359 163.367
R518 B.n360 B.n5 163.367
R519 B.n6 B.n5 163.367
R520 B.n7 B.n6 163.367
R521 B.n366 B.n7 163.367
R522 B.n367 B.n366 163.367
R523 B.n367 B.n13 163.367
R524 B.n14 B.n13 163.367
R525 B.n15 B.n14 163.367
R526 B.n372 B.n15 163.367
R527 B.n372 B.n20 163.367
R528 B.n21 B.n20 163.367
R529 B.n22 B.n21 163.367
R530 B.n377 B.n22 163.367
R531 B.n377 B.n27 163.367
R532 B.n28 B.n27 163.367
R533 B.n29 B.n28 163.367
R534 B.n382 B.n29 163.367
R535 B.n382 B.n34 163.367
R536 B.n35 B.n34 163.367
R537 B.n36 B.n35 163.367
R538 B.n387 B.n36 163.367
R539 B.n387 B.n41 163.367
R540 B.n42 B.n41 163.367
R541 B.n43 B.n42 163.367
R542 B.n392 B.n43 163.367
R543 B.n392 B.n48 163.367
R544 B.n49 B.n48 163.367
R545 B.n50 B.n49 163.367
R546 B.n397 B.n50 163.367
R547 B.n397 B.n55 163.367
R548 B.n56 B.n55 163.367
R549 B.n57 B.n56 163.367
R550 B.n402 B.n57 163.367
R551 B.n402 B.n62 163.367
R552 B.n63 B.n62 163.367
R553 B.n64 B.n63 163.367
R554 B.n407 B.n64 163.367
R555 B.n407 B.n69 163.367
R556 B.n70 B.n69 163.367
R557 B.n71 B.n70 163.367
R558 B.n243 B.n241 163.367
R559 B.n241 B.n240 163.367
R560 B.n237 B.n236 163.367
R561 B.n234 B.n172 163.367
R562 B.n230 B.n228 163.367
R563 B.n226 B.n174 163.367
R564 B.n222 B.n220 163.367
R565 B.n218 B.n179 163.367
R566 B.n214 B.n212 163.367
R567 B.n210 B.n181 163.367
R568 B.n205 B.n203 163.367
R569 B.n201 B.n185 163.367
R570 B.n197 B.n195 163.367
R571 B.n193 B.n187 163.367
R572 B.n189 B.n166 163.367
R573 B.n247 B.n162 163.367
R574 B.n255 B.n162 163.367
R575 B.n255 B.n160 163.367
R576 B.n259 B.n160 163.367
R577 B.n259 B.n154 163.367
R578 B.n267 B.n154 163.367
R579 B.n267 B.n152 163.367
R580 B.n271 B.n152 163.367
R581 B.n271 B.n146 163.367
R582 B.n279 B.n146 163.367
R583 B.n279 B.n144 163.367
R584 B.n283 B.n144 163.367
R585 B.n283 B.n138 163.367
R586 B.n291 B.n138 163.367
R587 B.n291 B.n136 163.367
R588 B.n295 B.n136 163.367
R589 B.n295 B.n130 163.367
R590 B.n303 B.n130 163.367
R591 B.n303 B.n128 163.367
R592 B.n307 B.n128 163.367
R593 B.n307 B.n122 163.367
R594 B.n315 B.n122 163.367
R595 B.n315 B.n120 163.367
R596 B.n319 B.n120 163.367
R597 B.n319 B.n114 163.367
R598 B.n327 B.n114 163.367
R599 B.n327 B.n112 163.367
R600 B.n331 B.n112 163.367
R601 B.n331 B.n106 163.367
R602 B.n340 B.n106 163.367
R603 B.n340 B.n104 163.367
R604 B.n344 B.n104 163.367
R605 B.n344 B.n99 163.367
R606 B.n353 B.n99 163.367
R607 B.n353 B.n97 163.367
R608 B.n357 B.n97 163.367
R609 B.n357 B.n3 163.367
R610 B.n550 B.n3 163.367
R611 B.n546 B.n2 163.367
R612 B.n546 B.n545 163.367
R613 B.n545 B.n9 163.367
R614 B.n541 B.n9 163.367
R615 B.n541 B.n11 163.367
R616 B.n537 B.n11 163.367
R617 B.n537 B.n16 163.367
R618 B.n533 B.n16 163.367
R619 B.n533 B.n18 163.367
R620 B.n529 B.n18 163.367
R621 B.n529 B.n24 163.367
R622 B.n525 B.n24 163.367
R623 B.n525 B.n26 163.367
R624 B.n521 B.n26 163.367
R625 B.n521 B.n31 163.367
R626 B.n517 B.n31 163.367
R627 B.n517 B.n33 163.367
R628 B.n513 B.n33 163.367
R629 B.n513 B.n38 163.367
R630 B.n509 B.n38 163.367
R631 B.n509 B.n40 163.367
R632 B.n505 B.n40 163.367
R633 B.n505 B.n45 163.367
R634 B.n501 B.n45 163.367
R635 B.n501 B.n47 163.367
R636 B.n497 B.n47 163.367
R637 B.n497 B.n52 163.367
R638 B.n493 B.n52 163.367
R639 B.n493 B.n54 163.367
R640 B.n489 B.n54 163.367
R641 B.n489 B.n59 163.367
R642 B.n485 B.n59 163.367
R643 B.n485 B.n61 163.367
R644 B.n481 B.n61 163.367
R645 B.n481 B.n66 163.367
R646 B.n477 B.n66 163.367
R647 B.n477 B.n68 163.367
R648 B.n473 B.n68 163.367
R649 B.n79 B.t14 150.761
R650 B.n87 B.t7 150.761
R651 B.n183 B.t16 150.761
R652 B.n176 B.t10 150.761
R653 B.n248 B.n163 113.249
R654 B.n254 B.n163 113.249
R655 B.n254 B.n159 113.249
R656 B.n260 B.n159 113.249
R657 B.n260 B.n155 113.249
R658 B.n266 B.n155 113.249
R659 B.n266 B.n151 113.249
R660 B.n272 B.n151 113.249
R661 B.n278 B.n147 113.249
R662 B.n278 B.n143 113.249
R663 B.n284 B.n143 113.249
R664 B.n284 B.n139 113.249
R665 B.n290 B.n139 113.249
R666 B.n290 B.n135 113.249
R667 B.n296 B.n135 113.249
R668 B.n296 B.n131 113.249
R669 B.n302 B.n131 113.249
R670 B.n302 B.n126 113.249
R671 B.n308 B.n126 113.249
R672 B.n308 B.n127 113.249
R673 B.n314 B.n119 113.249
R674 B.n320 B.n119 113.249
R675 B.n320 B.n115 113.249
R676 B.n326 B.n115 113.249
R677 B.n326 B.n111 113.249
R678 B.n332 B.n111 113.249
R679 B.n332 B.n107 113.249
R680 B.n339 B.n107 113.249
R681 B.n339 B.n338 113.249
R682 B.n345 B.n100 113.249
R683 B.n352 B.n100 113.249
R684 B.n352 B.n96 113.249
R685 B.n358 B.n96 113.249
R686 B.n358 B.n4 113.249
R687 B.n549 B.n4 113.249
R688 B.n549 B.n548 113.249
R689 B.n548 B.n547 113.249
R690 B.n547 B.n8 113.249
R691 B.n12 B.n8 113.249
R692 B.n540 B.n12 113.249
R693 B.n540 B.n539 113.249
R694 B.n539 B.n538 113.249
R695 B.n532 B.n19 113.249
R696 B.n532 B.n531 113.249
R697 B.n531 B.n530 113.249
R698 B.n530 B.n23 113.249
R699 B.n524 B.n23 113.249
R700 B.n524 B.n523 113.249
R701 B.n523 B.n522 113.249
R702 B.n522 B.n30 113.249
R703 B.n516 B.n30 113.249
R704 B.n515 B.n514 113.249
R705 B.n514 B.n37 113.249
R706 B.n508 B.n37 113.249
R707 B.n508 B.n507 113.249
R708 B.n507 B.n506 113.249
R709 B.n506 B.n44 113.249
R710 B.n500 B.n44 113.249
R711 B.n500 B.n499 113.249
R712 B.n499 B.n498 113.249
R713 B.n498 B.n51 113.249
R714 B.n492 B.n51 113.249
R715 B.n492 B.n491 113.249
R716 B.n490 B.n58 113.249
R717 B.n484 B.n58 113.249
R718 B.n484 B.n483 113.249
R719 B.n483 B.n482 113.249
R720 B.n482 B.n65 113.249
R721 B.n476 B.n65 113.249
R722 B.n476 B.n475 113.249
R723 B.n475 B.n474 113.249
R724 B.n338 B.t0 93.2632
R725 B.n19 B.t2 93.2632
R726 B.t9 B.n147 76.6091
R727 B.n127 B.t1 76.6091
R728 B.t3 B.n515 76.6091
R729 B.n491 B.t5 76.6091
R730 B.n468 B.n73 71.676
R731 B.n467 B.n466 71.676
R732 B.n460 B.n75 71.676
R733 B.n459 B.n458 71.676
R734 B.n452 B.n77 71.676
R735 B.n451 B.n81 71.676
R736 B.n447 B.n446 71.676
R737 B.n440 B.n83 71.676
R738 B.n439 B.n438 71.676
R739 B.n432 B.n85 71.676
R740 B.n431 B.n89 71.676
R741 B.n427 B.n426 71.676
R742 B.n420 B.n91 71.676
R743 B.n419 B.n418 71.676
R744 B.n412 B.n93 71.676
R745 B.n413 B.n412 71.676
R746 B.n418 B.n417 71.676
R747 B.n421 B.n420 71.676
R748 B.n426 B.n425 71.676
R749 B.n428 B.n89 71.676
R750 B.n433 B.n432 71.676
R751 B.n438 B.n437 71.676
R752 B.n441 B.n440 71.676
R753 B.n446 B.n445 71.676
R754 B.n448 B.n81 71.676
R755 B.n453 B.n452 71.676
R756 B.n458 B.n457 71.676
R757 B.n461 B.n460 71.676
R758 B.n466 B.n465 71.676
R759 B.n469 B.n468 71.676
R760 B.n242 B.n168 71.676
R761 B.n240 B.n170 71.676
R762 B.n236 B.n235 71.676
R763 B.n229 B.n172 71.676
R764 B.n228 B.n227 71.676
R765 B.n221 B.n174 71.676
R766 B.n220 B.n219 71.676
R767 B.n213 B.n179 71.676
R768 B.n212 B.n211 71.676
R769 B.n204 B.n181 71.676
R770 B.n203 B.n202 71.676
R771 B.n196 B.n185 71.676
R772 B.n195 B.n194 71.676
R773 B.n188 B.n187 71.676
R774 B.n243 B.n242 71.676
R775 B.n237 B.n170 71.676
R776 B.n235 B.n234 71.676
R777 B.n230 B.n229 71.676
R778 B.n227 B.n226 71.676
R779 B.n222 B.n221 71.676
R780 B.n219 B.n218 71.676
R781 B.n214 B.n213 71.676
R782 B.n211 B.n210 71.676
R783 B.n205 B.n204 71.676
R784 B.n202 B.n201 71.676
R785 B.n197 B.n196 71.676
R786 B.n194 B.n193 71.676
R787 B.n189 B.n188 71.676
R788 B.n551 B.n550 71.676
R789 B.n551 B.n2 71.676
R790 B.n79 B.n78 66.9096
R791 B.n87 B.n86 66.9096
R792 B.n183 B.n182 66.9096
R793 B.n176 B.n175 66.9096
R794 B.n80 B.n79 59.5399
R795 B.n88 B.n87 59.5399
R796 B.n207 B.n183 59.5399
R797 B.n177 B.n176 59.5399
R798 B.n272 B.t9 36.6394
R799 B.n314 B.t1 36.6394
R800 B.n516 B.t3 36.6394
R801 B.t5 B.n490 36.6394
R802 B.n246 B.n245 33.2493
R803 B.n250 B.n165 33.2493
R804 B.n414 B.n411 33.2493
R805 B.n472 B.n471 33.2493
R806 B.n345 B.t0 19.9854
R807 B.n538 B.t2 19.9854
R808 B B.n552 18.0485
R809 B.n246 B.n161 10.6151
R810 B.n256 B.n161 10.6151
R811 B.n257 B.n256 10.6151
R812 B.n258 B.n257 10.6151
R813 B.n258 B.n153 10.6151
R814 B.n268 B.n153 10.6151
R815 B.n269 B.n268 10.6151
R816 B.n270 B.n269 10.6151
R817 B.n270 B.n145 10.6151
R818 B.n280 B.n145 10.6151
R819 B.n281 B.n280 10.6151
R820 B.n282 B.n281 10.6151
R821 B.n282 B.n137 10.6151
R822 B.n292 B.n137 10.6151
R823 B.n293 B.n292 10.6151
R824 B.n294 B.n293 10.6151
R825 B.n294 B.n129 10.6151
R826 B.n304 B.n129 10.6151
R827 B.n305 B.n304 10.6151
R828 B.n306 B.n305 10.6151
R829 B.n306 B.n121 10.6151
R830 B.n316 B.n121 10.6151
R831 B.n317 B.n316 10.6151
R832 B.n318 B.n317 10.6151
R833 B.n318 B.n113 10.6151
R834 B.n328 B.n113 10.6151
R835 B.n329 B.n328 10.6151
R836 B.n330 B.n329 10.6151
R837 B.n330 B.n105 10.6151
R838 B.n341 B.n105 10.6151
R839 B.n342 B.n341 10.6151
R840 B.n343 B.n342 10.6151
R841 B.n343 B.n98 10.6151
R842 B.n354 B.n98 10.6151
R843 B.n355 B.n354 10.6151
R844 B.n356 B.n355 10.6151
R845 B.n356 B.n0 10.6151
R846 B.n245 B.n244 10.6151
R847 B.n244 B.n169 10.6151
R848 B.n239 B.n169 10.6151
R849 B.n239 B.n238 10.6151
R850 B.n238 B.n171 10.6151
R851 B.n233 B.n171 10.6151
R852 B.n233 B.n232 10.6151
R853 B.n232 B.n231 10.6151
R854 B.n231 B.n173 10.6151
R855 B.n225 B.n224 10.6151
R856 B.n224 B.n223 10.6151
R857 B.n223 B.n178 10.6151
R858 B.n217 B.n178 10.6151
R859 B.n217 B.n216 10.6151
R860 B.n216 B.n215 10.6151
R861 B.n215 B.n180 10.6151
R862 B.n209 B.n180 10.6151
R863 B.n209 B.n208 10.6151
R864 B.n206 B.n184 10.6151
R865 B.n200 B.n184 10.6151
R866 B.n200 B.n199 10.6151
R867 B.n199 B.n198 10.6151
R868 B.n198 B.n186 10.6151
R869 B.n192 B.n186 10.6151
R870 B.n192 B.n191 10.6151
R871 B.n191 B.n190 10.6151
R872 B.n190 B.n165 10.6151
R873 B.n251 B.n250 10.6151
R874 B.n252 B.n251 10.6151
R875 B.n252 B.n157 10.6151
R876 B.n262 B.n157 10.6151
R877 B.n263 B.n262 10.6151
R878 B.n264 B.n263 10.6151
R879 B.n264 B.n149 10.6151
R880 B.n274 B.n149 10.6151
R881 B.n275 B.n274 10.6151
R882 B.n276 B.n275 10.6151
R883 B.n276 B.n141 10.6151
R884 B.n286 B.n141 10.6151
R885 B.n287 B.n286 10.6151
R886 B.n288 B.n287 10.6151
R887 B.n288 B.n133 10.6151
R888 B.n298 B.n133 10.6151
R889 B.n299 B.n298 10.6151
R890 B.n300 B.n299 10.6151
R891 B.n300 B.n124 10.6151
R892 B.n310 B.n124 10.6151
R893 B.n311 B.n310 10.6151
R894 B.n312 B.n311 10.6151
R895 B.n312 B.n117 10.6151
R896 B.n322 B.n117 10.6151
R897 B.n323 B.n322 10.6151
R898 B.n324 B.n323 10.6151
R899 B.n324 B.n109 10.6151
R900 B.n334 B.n109 10.6151
R901 B.n335 B.n334 10.6151
R902 B.n336 B.n335 10.6151
R903 B.n336 B.n102 10.6151
R904 B.n347 B.n102 10.6151
R905 B.n348 B.n347 10.6151
R906 B.n350 B.n348 10.6151
R907 B.n350 B.n349 10.6151
R908 B.n349 B.n94 10.6151
R909 B.n361 B.n94 10.6151
R910 B.n362 B.n361 10.6151
R911 B.n363 B.n362 10.6151
R912 B.n364 B.n363 10.6151
R913 B.n365 B.n364 10.6151
R914 B.n368 B.n365 10.6151
R915 B.n369 B.n368 10.6151
R916 B.n370 B.n369 10.6151
R917 B.n371 B.n370 10.6151
R918 B.n373 B.n371 10.6151
R919 B.n374 B.n373 10.6151
R920 B.n375 B.n374 10.6151
R921 B.n376 B.n375 10.6151
R922 B.n378 B.n376 10.6151
R923 B.n379 B.n378 10.6151
R924 B.n380 B.n379 10.6151
R925 B.n381 B.n380 10.6151
R926 B.n383 B.n381 10.6151
R927 B.n384 B.n383 10.6151
R928 B.n385 B.n384 10.6151
R929 B.n386 B.n385 10.6151
R930 B.n388 B.n386 10.6151
R931 B.n389 B.n388 10.6151
R932 B.n390 B.n389 10.6151
R933 B.n391 B.n390 10.6151
R934 B.n393 B.n391 10.6151
R935 B.n394 B.n393 10.6151
R936 B.n395 B.n394 10.6151
R937 B.n396 B.n395 10.6151
R938 B.n398 B.n396 10.6151
R939 B.n399 B.n398 10.6151
R940 B.n400 B.n399 10.6151
R941 B.n401 B.n400 10.6151
R942 B.n403 B.n401 10.6151
R943 B.n404 B.n403 10.6151
R944 B.n405 B.n404 10.6151
R945 B.n406 B.n405 10.6151
R946 B.n408 B.n406 10.6151
R947 B.n409 B.n408 10.6151
R948 B.n410 B.n409 10.6151
R949 B.n411 B.n410 10.6151
R950 B.n544 B.n1 10.6151
R951 B.n544 B.n543 10.6151
R952 B.n543 B.n542 10.6151
R953 B.n542 B.n10 10.6151
R954 B.n536 B.n10 10.6151
R955 B.n536 B.n535 10.6151
R956 B.n535 B.n534 10.6151
R957 B.n534 B.n17 10.6151
R958 B.n528 B.n17 10.6151
R959 B.n528 B.n527 10.6151
R960 B.n527 B.n526 10.6151
R961 B.n526 B.n25 10.6151
R962 B.n520 B.n25 10.6151
R963 B.n520 B.n519 10.6151
R964 B.n519 B.n518 10.6151
R965 B.n518 B.n32 10.6151
R966 B.n512 B.n32 10.6151
R967 B.n512 B.n511 10.6151
R968 B.n511 B.n510 10.6151
R969 B.n510 B.n39 10.6151
R970 B.n504 B.n39 10.6151
R971 B.n504 B.n503 10.6151
R972 B.n503 B.n502 10.6151
R973 B.n502 B.n46 10.6151
R974 B.n496 B.n46 10.6151
R975 B.n496 B.n495 10.6151
R976 B.n495 B.n494 10.6151
R977 B.n494 B.n53 10.6151
R978 B.n488 B.n53 10.6151
R979 B.n488 B.n487 10.6151
R980 B.n487 B.n486 10.6151
R981 B.n486 B.n60 10.6151
R982 B.n480 B.n60 10.6151
R983 B.n480 B.n479 10.6151
R984 B.n479 B.n478 10.6151
R985 B.n478 B.n67 10.6151
R986 B.n472 B.n67 10.6151
R987 B.n471 B.n470 10.6151
R988 B.n470 B.n74 10.6151
R989 B.n464 B.n74 10.6151
R990 B.n464 B.n463 10.6151
R991 B.n463 B.n462 10.6151
R992 B.n462 B.n76 10.6151
R993 B.n456 B.n76 10.6151
R994 B.n456 B.n455 10.6151
R995 B.n455 B.n454 10.6151
R996 B.n450 B.n449 10.6151
R997 B.n449 B.n82 10.6151
R998 B.n444 B.n82 10.6151
R999 B.n444 B.n443 10.6151
R1000 B.n443 B.n442 10.6151
R1001 B.n442 B.n84 10.6151
R1002 B.n436 B.n84 10.6151
R1003 B.n436 B.n435 10.6151
R1004 B.n435 B.n434 10.6151
R1005 B.n430 B.n429 10.6151
R1006 B.n429 B.n90 10.6151
R1007 B.n424 B.n90 10.6151
R1008 B.n424 B.n423 10.6151
R1009 B.n423 B.n422 10.6151
R1010 B.n422 B.n92 10.6151
R1011 B.n416 B.n92 10.6151
R1012 B.n416 B.n415 10.6151
R1013 B.n415 B.n414 10.6151
R1014 B.n177 B.n173 9.36635
R1015 B.n207 B.n206 9.36635
R1016 B.n454 B.n80 9.36635
R1017 B.n430 B.n88 9.36635
R1018 B.n552 B.n0 8.11757
R1019 B.n552 B.n1 8.11757
R1020 B.n225 B.n177 1.24928
R1021 B.n208 B.n207 1.24928
R1022 B.n450 B.n80 1.24928
R1023 B.n434 B.n88 1.24928
R1024 VN.n0 VN.t3 44.7876
R1025 VN.n1 VN.t1 44.7876
R1026 VN.n0 VN.t0 43.7682
R1027 VN.n1 VN.t2 43.7682
R1028 VN VN.n1 42.9133
R1029 VN VN.n0 2.79586
R1030 VDD2.n2 VDD2.n0 181.183
R1031 VDD2.n2 VDD2.n1 147.399
R1032 VDD2.n1 VDD2.t1 14.8877
R1033 VDD2.n1 VDD2.t2 14.8877
R1034 VDD2.n0 VDD2.t0 14.8877
R1035 VDD2.n0 VDD2.t3 14.8877
R1036 VDD2 VDD2.n2 0.0586897
C0 VDD1 VTAIL 3.15f
C1 VTAIL VN 1.60841f
C2 VP VTAIL 1.62251f
C3 VDD2 VTAIL 3.2077f
C4 VDD1 VN 0.15615f
C5 VP VDD1 1.11285f
C6 VDD2 VDD1 1.15471f
C7 VP VN 4.59607f
C8 VDD2 VN 0.83602f
C9 VP VDD2 0.435352f
C10 VDD2 B 3.190249f
C11 VDD1 B 5.86355f
C12 VTAIL B 3.40333f
C13 VN B 10.429111f
C14 VP B 9.049264f
C15 VDD2.t0 B 0.025051f
C16 VDD2.t3 B 0.025051f
C17 VDD2.n0 B 0.288679f
C18 VDD2.t1 B 0.025051f
C19 VDD2.t2 B 0.025051f
C20 VDD2.n1 B 0.125641f
C21 VDD2.n2 B 2.45193f
C22 VN.t0 B 0.415856f
C23 VN.t3 B 0.42264f
C24 VN.n0 B 0.28508f
C25 VN.t1 B 0.42264f
C26 VN.t2 B 0.415856f
C27 VN.n1 B 1.37514f
C28 VDD1.t0 B 0.023618f
C29 VDD1.t3 B 0.023618f
C30 VDD1.n0 B 0.118611f
C31 VDD1.t2 B 0.023618f
C32 VDD1.t1 B 0.023618f
C33 VDD1.n1 B 0.282673f
C34 VTAIL.t2 B 0.127711f
C35 VTAIL.n0 B 0.300052f
C36 VTAIL.t6 B 0.127711f
C37 VTAIL.n1 B 0.395913f
C38 VTAIL.t5 B 0.127711f
C39 VTAIL.n2 B 0.923665f
C40 VTAIL.t1 B 0.127711f
C41 VTAIL.n3 B 0.923665f
C42 VTAIL.t0 B 0.127711f
C43 VTAIL.n4 B 0.395913f
C44 VTAIL.t7 B 0.127711f
C45 VTAIL.n5 B 0.395913f
C46 VTAIL.t4 B 0.127711f
C47 VTAIL.n6 B 0.923665f
C48 VTAIL.t3 B 0.127711f
C49 VTAIL.n7 B 0.819996f
C50 VP.t2 B 0.203916f
C51 VP.n0 B 0.213581f
C52 VP.n1 B 0.023399f
C53 VP.n2 B 0.034159f
C54 VP.n3 B 0.037766f
C55 VP.t1 B 0.203916f
C56 VP.t3 B 0.425661f
C57 VP.t0 B 0.418829f
C58 VP.n4 B 1.37495f
C59 VP.n5 B 1.0382f
C60 VP.n6 B 0.213581f
C61 VP.n7 B 0.042533f
C62 VP.n8 B 0.043611f
C63 VP.n9 B 0.023399f
C64 VP.n10 B 0.023399f
C65 VP.n11 B 0.023399f
C66 VP.n12 B 0.034159f
C67 VP.n13 B 0.043611f
C68 VP.n14 B 0.042533f
C69 VP.n15 B 0.037766f
C70 VP.n16 B 0.045765f
.ends

