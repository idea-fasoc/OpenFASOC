* NGSPICE file created from diff_pair_sample_0707.ext - technology: sky130A

.subckt diff_pair_sample_0707 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=2.31825 pd=14.38 as=5.4795 ps=28.88 w=14.05 l=3.49
X1 VDD2.t3 VN.t0 VTAIL.t0 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=2.31825 pd=14.38 as=5.4795 ps=28.88 w=14.05 l=3.49
X2 VDD2.t2 VN.t1 VTAIL.t2 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=2.31825 pd=14.38 as=5.4795 ps=28.88 w=14.05 l=3.49
X3 VTAIL.t1 VN.t2 VDD2.t1 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=5.4795 pd=28.88 as=2.31825 ps=14.38 w=14.05 l=3.49
X4 B.t11 B.t9 B.t10 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=5.4795 pd=28.88 as=0 ps=0 w=14.05 l=3.49
X5 B.t8 B.t6 B.t7 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=5.4795 pd=28.88 as=0 ps=0 w=14.05 l=3.49
X6 B.t5 B.t3 B.t4 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=5.4795 pd=28.88 as=0 ps=0 w=14.05 l=3.49
X7 B.t2 B.t0 B.t1 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=5.4795 pd=28.88 as=0 ps=0 w=14.05 l=3.49
X8 VTAIL.t3 VN.t3 VDD2.t0 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=5.4795 pd=28.88 as=2.31825 ps=14.38 w=14.05 l=3.49
X9 VTAIL.t7 VP.t1 VDD1.t2 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=5.4795 pd=28.88 as=2.31825 ps=14.38 w=14.05 l=3.49
X10 VDD1.t1 VP.t2 VTAIL.t6 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=2.31825 pd=14.38 as=5.4795 ps=28.88 w=14.05 l=3.49
X11 VTAIL.t4 VP.t3 VDD1.t0 w_n3262_n3778# sky130_fd_pr__pfet_01v8 ad=5.4795 pd=28.88 as=2.31825 ps=14.38 w=14.05 l=3.49
R0 VP.n19 VP.n18 161.3
R1 VP.n17 VP.n1 161.3
R2 VP.n16 VP.n15 161.3
R3 VP.n14 VP.n2 161.3
R4 VP.n13 VP.n12 161.3
R5 VP.n11 VP.n3 161.3
R6 VP.n10 VP.n9 161.3
R7 VP.n8 VP.n4 161.3
R8 VP.n5 VP.t1 131.412
R9 VP.n5 VP.t0 130.196
R10 VP.n6 VP.t3 97.022
R11 VP.n0 VP.t2 97.022
R12 VP.n7 VP.n6 82.238
R13 VP.n20 VP.n0 82.238
R14 VP.n12 VP.n2 56.5193
R15 VP.n7 VP.n5 52.8224
R16 VP.n10 VP.n4 24.4675
R17 VP.n11 VP.n10 24.4675
R18 VP.n12 VP.n11 24.4675
R19 VP.n16 VP.n2 24.4675
R20 VP.n17 VP.n16 24.4675
R21 VP.n18 VP.n17 24.4675
R22 VP.n6 VP.n4 7.82994
R23 VP.n18 VP.n0 7.82994
R24 VP.n8 VP.n7 0.354971
R25 VP.n20 VP.n19 0.354971
R26 VP VP.n20 0.26696
R27 VP.n9 VP.n8 0.189894
R28 VP.n9 VP.n3 0.189894
R29 VP.n13 VP.n3 0.189894
R30 VP.n14 VP.n13 0.189894
R31 VP.n15 VP.n14 0.189894
R32 VP.n15 VP.n1 0.189894
R33 VP.n19 VP.n1 0.189894
R34 VTAIL.n618 VTAIL.n546 756.745
R35 VTAIL.n72 VTAIL.n0 756.745
R36 VTAIL.n150 VTAIL.n78 756.745
R37 VTAIL.n228 VTAIL.n156 756.745
R38 VTAIL.n540 VTAIL.n468 756.745
R39 VTAIL.n462 VTAIL.n390 756.745
R40 VTAIL.n384 VTAIL.n312 756.745
R41 VTAIL.n306 VTAIL.n234 756.745
R42 VTAIL.n570 VTAIL.n569 585
R43 VTAIL.n575 VTAIL.n574 585
R44 VTAIL.n577 VTAIL.n576 585
R45 VTAIL.n566 VTAIL.n565 585
R46 VTAIL.n583 VTAIL.n582 585
R47 VTAIL.n585 VTAIL.n584 585
R48 VTAIL.n562 VTAIL.n561 585
R49 VTAIL.n591 VTAIL.n590 585
R50 VTAIL.n593 VTAIL.n592 585
R51 VTAIL.n558 VTAIL.n557 585
R52 VTAIL.n599 VTAIL.n598 585
R53 VTAIL.n601 VTAIL.n600 585
R54 VTAIL.n554 VTAIL.n553 585
R55 VTAIL.n607 VTAIL.n606 585
R56 VTAIL.n609 VTAIL.n608 585
R57 VTAIL.n550 VTAIL.n549 585
R58 VTAIL.n616 VTAIL.n615 585
R59 VTAIL.n617 VTAIL.n548 585
R60 VTAIL.n619 VTAIL.n618 585
R61 VTAIL.n24 VTAIL.n23 585
R62 VTAIL.n29 VTAIL.n28 585
R63 VTAIL.n31 VTAIL.n30 585
R64 VTAIL.n20 VTAIL.n19 585
R65 VTAIL.n37 VTAIL.n36 585
R66 VTAIL.n39 VTAIL.n38 585
R67 VTAIL.n16 VTAIL.n15 585
R68 VTAIL.n45 VTAIL.n44 585
R69 VTAIL.n47 VTAIL.n46 585
R70 VTAIL.n12 VTAIL.n11 585
R71 VTAIL.n53 VTAIL.n52 585
R72 VTAIL.n55 VTAIL.n54 585
R73 VTAIL.n8 VTAIL.n7 585
R74 VTAIL.n61 VTAIL.n60 585
R75 VTAIL.n63 VTAIL.n62 585
R76 VTAIL.n4 VTAIL.n3 585
R77 VTAIL.n70 VTAIL.n69 585
R78 VTAIL.n71 VTAIL.n2 585
R79 VTAIL.n73 VTAIL.n72 585
R80 VTAIL.n102 VTAIL.n101 585
R81 VTAIL.n107 VTAIL.n106 585
R82 VTAIL.n109 VTAIL.n108 585
R83 VTAIL.n98 VTAIL.n97 585
R84 VTAIL.n115 VTAIL.n114 585
R85 VTAIL.n117 VTAIL.n116 585
R86 VTAIL.n94 VTAIL.n93 585
R87 VTAIL.n123 VTAIL.n122 585
R88 VTAIL.n125 VTAIL.n124 585
R89 VTAIL.n90 VTAIL.n89 585
R90 VTAIL.n131 VTAIL.n130 585
R91 VTAIL.n133 VTAIL.n132 585
R92 VTAIL.n86 VTAIL.n85 585
R93 VTAIL.n139 VTAIL.n138 585
R94 VTAIL.n141 VTAIL.n140 585
R95 VTAIL.n82 VTAIL.n81 585
R96 VTAIL.n148 VTAIL.n147 585
R97 VTAIL.n149 VTAIL.n80 585
R98 VTAIL.n151 VTAIL.n150 585
R99 VTAIL.n180 VTAIL.n179 585
R100 VTAIL.n185 VTAIL.n184 585
R101 VTAIL.n187 VTAIL.n186 585
R102 VTAIL.n176 VTAIL.n175 585
R103 VTAIL.n193 VTAIL.n192 585
R104 VTAIL.n195 VTAIL.n194 585
R105 VTAIL.n172 VTAIL.n171 585
R106 VTAIL.n201 VTAIL.n200 585
R107 VTAIL.n203 VTAIL.n202 585
R108 VTAIL.n168 VTAIL.n167 585
R109 VTAIL.n209 VTAIL.n208 585
R110 VTAIL.n211 VTAIL.n210 585
R111 VTAIL.n164 VTAIL.n163 585
R112 VTAIL.n217 VTAIL.n216 585
R113 VTAIL.n219 VTAIL.n218 585
R114 VTAIL.n160 VTAIL.n159 585
R115 VTAIL.n226 VTAIL.n225 585
R116 VTAIL.n227 VTAIL.n158 585
R117 VTAIL.n229 VTAIL.n228 585
R118 VTAIL.n541 VTAIL.n540 585
R119 VTAIL.n539 VTAIL.n470 585
R120 VTAIL.n538 VTAIL.n537 585
R121 VTAIL.n473 VTAIL.n471 585
R122 VTAIL.n532 VTAIL.n531 585
R123 VTAIL.n530 VTAIL.n529 585
R124 VTAIL.n477 VTAIL.n476 585
R125 VTAIL.n524 VTAIL.n523 585
R126 VTAIL.n522 VTAIL.n521 585
R127 VTAIL.n481 VTAIL.n480 585
R128 VTAIL.n516 VTAIL.n515 585
R129 VTAIL.n514 VTAIL.n513 585
R130 VTAIL.n485 VTAIL.n484 585
R131 VTAIL.n508 VTAIL.n507 585
R132 VTAIL.n506 VTAIL.n505 585
R133 VTAIL.n489 VTAIL.n488 585
R134 VTAIL.n500 VTAIL.n499 585
R135 VTAIL.n498 VTAIL.n497 585
R136 VTAIL.n493 VTAIL.n492 585
R137 VTAIL.n463 VTAIL.n462 585
R138 VTAIL.n461 VTAIL.n392 585
R139 VTAIL.n460 VTAIL.n459 585
R140 VTAIL.n395 VTAIL.n393 585
R141 VTAIL.n454 VTAIL.n453 585
R142 VTAIL.n452 VTAIL.n451 585
R143 VTAIL.n399 VTAIL.n398 585
R144 VTAIL.n446 VTAIL.n445 585
R145 VTAIL.n444 VTAIL.n443 585
R146 VTAIL.n403 VTAIL.n402 585
R147 VTAIL.n438 VTAIL.n437 585
R148 VTAIL.n436 VTAIL.n435 585
R149 VTAIL.n407 VTAIL.n406 585
R150 VTAIL.n430 VTAIL.n429 585
R151 VTAIL.n428 VTAIL.n427 585
R152 VTAIL.n411 VTAIL.n410 585
R153 VTAIL.n422 VTAIL.n421 585
R154 VTAIL.n420 VTAIL.n419 585
R155 VTAIL.n415 VTAIL.n414 585
R156 VTAIL.n385 VTAIL.n384 585
R157 VTAIL.n383 VTAIL.n314 585
R158 VTAIL.n382 VTAIL.n381 585
R159 VTAIL.n317 VTAIL.n315 585
R160 VTAIL.n376 VTAIL.n375 585
R161 VTAIL.n374 VTAIL.n373 585
R162 VTAIL.n321 VTAIL.n320 585
R163 VTAIL.n368 VTAIL.n367 585
R164 VTAIL.n366 VTAIL.n365 585
R165 VTAIL.n325 VTAIL.n324 585
R166 VTAIL.n360 VTAIL.n359 585
R167 VTAIL.n358 VTAIL.n357 585
R168 VTAIL.n329 VTAIL.n328 585
R169 VTAIL.n352 VTAIL.n351 585
R170 VTAIL.n350 VTAIL.n349 585
R171 VTAIL.n333 VTAIL.n332 585
R172 VTAIL.n344 VTAIL.n343 585
R173 VTAIL.n342 VTAIL.n341 585
R174 VTAIL.n337 VTAIL.n336 585
R175 VTAIL.n307 VTAIL.n306 585
R176 VTAIL.n305 VTAIL.n236 585
R177 VTAIL.n304 VTAIL.n303 585
R178 VTAIL.n239 VTAIL.n237 585
R179 VTAIL.n298 VTAIL.n297 585
R180 VTAIL.n296 VTAIL.n295 585
R181 VTAIL.n243 VTAIL.n242 585
R182 VTAIL.n290 VTAIL.n289 585
R183 VTAIL.n288 VTAIL.n287 585
R184 VTAIL.n247 VTAIL.n246 585
R185 VTAIL.n282 VTAIL.n281 585
R186 VTAIL.n280 VTAIL.n279 585
R187 VTAIL.n251 VTAIL.n250 585
R188 VTAIL.n274 VTAIL.n273 585
R189 VTAIL.n272 VTAIL.n271 585
R190 VTAIL.n255 VTAIL.n254 585
R191 VTAIL.n266 VTAIL.n265 585
R192 VTAIL.n264 VTAIL.n263 585
R193 VTAIL.n259 VTAIL.n258 585
R194 VTAIL.n571 VTAIL.t0 327.466
R195 VTAIL.n25 VTAIL.t1 327.466
R196 VTAIL.n103 VTAIL.t6 327.466
R197 VTAIL.n181 VTAIL.t4 327.466
R198 VTAIL.n494 VTAIL.t5 327.466
R199 VTAIL.n416 VTAIL.t7 327.466
R200 VTAIL.n338 VTAIL.t2 327.466
R201 VTAIL.n260 VTAIL.t3 327.466
R202 VTAIL.n575 VTAIL.n569 171.744
R203 VTAIL.n576 VTAIL.n575 171.744
R204 VTAIL.n576 VTAIL.n565 171.744
R205 VTAIL.n583 VTAIL.n565 171.744
R206 VTAIL.n584 VTAIL.n583 171.744
R207 VTAIL.n584 VTAIL.n561 171.744
R208 VTAIL.n591 VTAIL.n561 171.744
R209 VTAIL.n592 VTAIL.n591 171.744
R210 VTAIL.n592 VTAIL.n557 171.744
R211 VTAIL.n599 VTAIL.n557 171.744
R212 VTAIL.n600 VTAIL.n599 171.744
R213 VTAIL.n600 VTAIL.n553 171.744
R214 VTAIL.n607 VTAIL.n553 171.744
R215 VTAIL.n608 VTAIL.n607 171.744
R216 VTAIL.n608 VTAIL.n549 171.744
R217 VTAIL.n616 VTAIL.n549 171.744
R218 VTAIL.n617 VTAIL.n616 171.744
R219 VTAIL.n618 VTAIL.n617 171.744
R220 VTAIL.n29 VTAIL.n23 171.744
R221 VTAIL.n30 VTAIL.n29 171.744
R222 VTAIL.n30 VTAIL.n19 171.744
R223 VTAIL.n37 VTAIL.n19 171.744
R224 VTAIL.n38 VTAIL.n37 171.744
R225 VTAIL.n38 VTAIL.n15 171.744
R226 VTAIL.n45 VTAIL.n15 171.744
R227 VTAIL.n46 VTAIL.n45 171.744
R228 VTAIL.n46 VTAIL.n11 171.744
R229 VTAIL.n53 VTAIL.n11 171.744
R230 VTAIL.n54 VTAIL.n53 171.744
R231 VTAIL.n54 VTAIL.n7 171.744
R232 VTAIL.n61 VTAIL.n7 171.744
R233 VTAIL.n62 VTAIL.n61 171.744
R234 VTAIL.n62 VTAIL.n3 171.744
R235 VTAIL.n70 VTAIL.n3 171.744
R236 VTAIL.n71 VTAIL.n70 171.744
R237 VTAIL.n72 VTAIL.n71 171.744
R238 VTAIL.n107 VTAIL.n101 171.744
R239 VTAIL.n108 VTAIL.n107 171.744
R240 VTAIL.n108 VTAIL.n97 171.744
R241 VTAIL.n115 VTAIL.n97 171.744
R242 VTAIL.n116 VTAIL.n115 171.744
R243 VTAIL.n116 VTAIL.n93 171.744
R244 VTAIL.n123 VTAIL.n93 171.744
R245 VTAIL.n124 VTAIL.n123 171.744
R246 VTAIL.n124 VTAIL.n89 171.744
R247 VTAIL.n131 VTAIL.n89 171.744
R248 VTAIL.n132 VTAIL.n131 171.744
R249 VTAIL.n132 VTAIL.n85 171.744
R250 VTAIL.n139 VTAIL.n85 171.744
R251 VTAIL.n140 VTAIL.n139 171.744
R252 VTAIL.n140 VTAIL.n81 171.744
R253 VTAIL.n148 VTAIL.n81 171.744
R254 VTAIL.n149 VTAIL.n148 171.744
R255 VTAIL.n150 VTAIL.n149 171.744
R256 VTAIL.n185 VTAIL.n179 171.744
R257 VTAIL.n186 VTAIL.n185 171.744
R258 VTAIL.n186 VTAIL.n175 171.744
R259 VTAIL.n193 VTAIL.n175 171.744
R260 VTAIL.n194 VTAIL.n193 171.744
R261 VTAIL.n194 VTAIL.n171 171.744
R262 VTAIL.n201 VTAIL.n171 171.744
R263 VTAIL.n202 VTAIL.n201 171.744
R264 VTAIL.n202 VTAIL.n167 171.744
R265 VTAIL.n209 VTAIL.n167 171.744
R266 VTAIL.n210 VTAIL.n209 171.744
R267 VTAIL.n210 VTAIL.n163 171.744
R268 VTAIL.n217 VTAIL.n163 171.744
R269 VTAIL.n218 VTAIL.n217 171.744
R270 VTAIL.n218 VTAIL.n159 171.744
R271 VTAIL.n226 VTAIL.n159 171.744
R272 VTAIL.n227 VTAIL.n226 171.744
R273 VTAIL.n228 VTAIL.n227 171.744
R274 VTAIL.n540 VTAIL.n539 171.744
R275 VTAIL.n539 VTAIL.n538 171.744
R276 VTAIL.n538 VTAIL.n471 171.744
R277 VTAIL.n531 VTAIL.n471 171.744
R278 VTAIL.n531 VTAIL.n530 171.744
R279 VTAIL.n530 VTAIL.n476 171.744
R280 VTAIL.n523 VTAIL.n476 171.744
R281 VTAIL.n523 VTAIL.n522 171.744
R282 VTAIL.n522 VTAIL.n480 171.744
R283 VTAIL.n515 VTAIL.n480 171.744
R284 VTAIL.n515 VTAIL.n514 171.744
R285 VTAIL.n514 VTAIL.n484 171.744
R286 VTAIL.n507 VTAIL.n484 171.744
R287 VTAIL.n507 VTAIL.n506 171.744
R288 VTAIL.n506 VTAIL.n488 171.744
R289 VTAIL.n499 VTAIL.n488 171.744
R290 VTAIL.n499 VTAIL.n498 171.744
R291 VTAIL.n498 VTAIL.n492 171.744
R292 VTAIL.n462 VTAIL.n461 171.744
R293 VTAIL.n461 VTAIL.n460 171.744
R294 VTAIL.n460 VTAIL.n393 171.744
R295 VTAIL.n453 VTAIL.n393 171.744
R296 VTAIL.n453 VTAIL.n452 171.744
R297 VTAIL.n452 VTAIL.n398 171.744
R298 VTAIL.n445 VTAIL.n398 171.744
R299 VTAIL.n445 VTAIL.n444 171.744
R300 VTAIL.n444 VTAIL.n402 171.744
R301 VTAIL.n437 VTAIL.n402 171.744
R302 VTAIL.n437 VTAIL.n436 171.744
R303 VTAIL.n436 VTAIL.n406 171.744
R304 VTAIL.n429 VTAIL.n406 171.744
R305 VTAIL.n429 VTAIL.n428 171.744
R306 VTAIL.n428 VTAIL.n410 171.744
R307 VTAIL.n421 VTAIL.n410 171.744
R308 VTAIL.n421 VTAIL.n420 171.744
R309 VTAIL.n420 VTAIL.n414 171.744
R310 VTAIL.n384 VTAIL.n383 171.744
R311 VTAIL.n383 VTAIL.n382 171.744
R312 VTAIL.n382 VTAIL.n315 171.744
R313 VTAIL.n375 VTAIL.n315 171.744
R314 VTAIL.n375 VTAIL.n374 171.744
R315 VTAIL.n374 VTAIL.n320 171.744
R316 VTAIL.n367 VTAIL.n320 171.744
R317 VTAIL.n367 VTAIL.n366 171.744
R318 VTAIL.n366 VTAIL.n324 171.744
R319 VTAIL.n359 VTAIL.n324 171.744
R320 VTAIL.n359 VTAIL.n358 171.744
R321 VTAIL.n358 VTAIL.n328 171.744
R322 VTAIL.n351 VTAIL.n328 171.744
R323 VTAIL.n351 VTAIL.n350 171.744
R324 VTAIL.n350 VTAIL.n332 171.744
R325 VTAIL.n343 VTAIL.n332 171.744
R326 VTAIL.n343 VTAIL.n342 171.744
R327 VTAIL.n342 VTAIL.n336 171.744
R328 VTAIL.n306 VTAIL.n305 171.744
R329 VTAIL.n305 VTAIL.n304 171.744
R330 VTAIL.n304 VTAIL.n237 171.744
R331 VTAIL.n297 VTAIL.n237 171.744
R332 VTAIL.n297 VTAIL.n296 171.744
R333 VTAIL.n296 VTAIL.n242 171.744
R334 VTAIL.n289 VTAIL.n242 171.744
R335 VTAIL.n289 VTAIL.n288 171.744
R336 VTAIL.n288 VTAIL.n246 171.744
R337 VTAIL.n281 VTAIL.n246 171.744
R338 VTAIL.n281 VTAIL.n280 171.744
R339 VTAIL.n280 VTAIL.n250 171.744
R340 VTAIL.n273 VTAIL.n250 171.744
R341 VTAIL.n273 VTAIL.n272 171.744
R342 VTAIL.n272 VTAIL.n254 171.744
R343 VTAIL.n265 VTAIL.n254 171.744
R344 VTAIL.n265 VTAIL.n264 171.744
R345 VTAIL.n264 VTAIL.n258 171.744
R346 VTAIL.t0 VTAIL.n569 85.8723
R347 VTAIL.t1 VTAIL.n23 85.8723
R348 VTAIL.t6 VTAIL.n101 85.8723
R349 VTAIL.t4 VTAIL.n179 85.8723
R350 VTAIL.t5 VTAIL.n492 85.8723
R351 VTAIL.t7 VTAIL.n414 85.8723
R352 VTAIL.t2 VTAIL.n336 85.8723
R353 VTAIL.t3 VTAIL.n258 85.8723
R354 VTAIL.n623 VTAIL.n622 34.7066
R355 VTAIL.n77 VTAIL.n76 34.7066
R356 VTAIL.n155 VTAIL.n154 34.7066
R357 VTAIL.n233 VTAIL.n232 34.7066
R358 VTAIL.n545 VTAIL.n544 34.7066
R359 VTAIL.n467 VTAIL.n466 34.7066
R360 VTAIL.n389 VTAIL.n388 34.7066
R361 VTAIL.n311 VTAIL.n310 34.7066
R362 VTAIL.n623 VTAIL.n545 27.7721
R363 VTAIL.n311 VTAIL.n233 27.7721
R364 VTAIL.n571 VTAIL.n570 16.3895
R365 VTAIL.n25 VTAIL.n24 16.3895
R366 VTAIL.n103 VTAIL.n102 16.3895
R367 VTAIL.n181 VTAIL.n180 16.3895
R368 VTAIL.n494 VTAIL.n493 16.3895
R369 VTAIL.n416 VTAIL.n415 16.3895
R370 VTAIL.n338 VTAIL.n337 16.3895
R371 VTAIL.n260 VTAIL.n259 16.3895
R372 VTAIL.n619 VTAIL.n548 13.1884
R373 VTAIL.n73 VTAIL.n2 13.1884
R374 VTAIL.n151 VTAIL.n80 13.1884
R375 VTAIL.n229 VTAIL.n158 13.1884
R376 VTAIL.n541 VTAIL.n470 13.1884
R377 VTAIL.n463 VTAIL.n392 13.1884
R378 VTAIL.n385 VTAIL.n314 13.1884
R379 VTAIL.n307 VTAIL.n236 13.1884
R380 VTAIL.n574 VTAIL.n573 12.8005
R381 VTAIL.n615 VTAIL.n614 12.8005
R382 VTAIL.n620 VTAIL.n546 12.8005
R383 VTAIL.n28 VTAIL.n27 12.8005
R384 VTAIL.n69 VTAIL.n68 12.8005
R385 VTAIL.n74 VTAIL.n0 12.8005
R386 VTAIL.n106 VTAIL.n105 12.8005
R387 VTAIL.n147 VTAIL.n146 12.8005
R388 VTAIL.n152 VTAIL.n78 12.8005
R389 VTAIL.n184 VTAIL.n183 12.8005
R390 VTAIL.n225 VTAIL.n224 12.8005
R391 VTAIL.n230 VTAIL.n156 12.8005
R392 VTAIL.n542 VTAIL.n468 12.8005
R393 VTAIL.n537 VTAIL.n472 12.8005
R394 VTAIL.n497 VTAIL.n496 12.8005
R395 VTAIL.n464 VTAIL.n390 12.8005
R396 VTAIL.n459 VTAIL.n394 12.8005
R397 VTAIL.n419 VTAIL.n418 12.8005
R398 VTAIL.n386 VTAIL.n312 12.8005
R399 VTAIL.n381 VTAIL.n316 12.8005
R400 VTAIL.n341 VTAIL.n340 12.8005
R401 VTAIL.n308 VTAIL.n234 12.8005
R402 VTAIL.n303 VTAIL.n238 12.8005
R403 VTAIL.n263 VTAIL.n262 12.8005
R404 VTAIL.n577 VTAIL.n568 12.0247
R405 VTAIL.n613 VTAIL.n550 12.0247
R406 VTAIL.n31 VTAIL.n22 12.0247
R407 VTAIL.n67 VTAIL.n4 12.0247
R408 VTAIL.n109 VTAIL.n100 12.0247
R409 VTAIL.n145 VTAIL.n82 12.0247
R410 VTAIL.n187 VTAIL.n178 12.0247
R411 VTAIL.n223 VTAIL.n160 12.0247
R412 VTAIL.n536 VTAIL.n473 12.0247
R413 VTAIL.n500 VTAIL.n491 12.0247
R414 VTAIL.n458 VTAIL.n395 12.0247
R415 VTAIL.n422 VTAIL.n413 12.0247
R416 VTAIL.n380 VTAIL.n317 12.0247
R417 VTAIL.n344 VTAIL.n335 12.0247
R418 VTAIL.n302 VTAIL.n239 12.0247
R419 VTAIL.n266 VTAIL.n257 12.0247
R420 VTAIL.n578 VTAIL.n566 11.249
R421 VTAIL.n610 VTAIL.n609 11.249
R422 VTAIL.n32 VTAIL.n20 11.249
R423 VTAIL.n64 VTAIL.n63 11.249
R424 VTAIL.n110 VTAIL.n98 11.249
R425 VTAIL.n142 VTAIL.n141 11.249
R426 VTAIL.n188 VTAIL.n176 11.249
R427 VTAIL.n220 VTAIL.n219 11.249
R428 VTAIL.n533 VTAIL.n532 11.249
R429 VTAIL.n501 VTAIL.n489 11.249
R430 VTAIL.n455 VTAIL.n454 11.249
R431 VTAIL.n423 VTAIL.n411 11.249
R432 VTAIL.n377 VTAIL.n376 11.249
R433 VTAIL.n345 VTAIL.n333 11.249
R434 VTAIL.n299 VTAIL.n298 11.249
R435 VTAIL.n267 VTAIL.n255 11.249
R436 VTAIL.n582 VTAIL.n581 10.4732
R437 VTAIL.n606 VTAIL.n552 10.4732
R438 VTAIL.n36 VTAIL.n35 10.4732
R439 VTAIL.n60 VTAIL.n6 10.4732
R440 VTAIL.n114 VTAIL.n113 10.4732
R441 VTAIL.n138 VTAIL.n84 10.4732
R442 VTAIL.n192 VTAIL.n191 10.4732
R443 VTAIL.n216 VTAIL.n162 10.4732
R444 VTAIL.n529 VTAIL.n475 10.4732
R445 VTAIL.n505 VTAIL.n504 10.4732
R446 VTAIL.n451 VTAIL.n397 10.4732
R447 VTAIL.n427 VTAIL.n426 10.4732
R448 VTAIL.n373 VTAIL.n319 10.4732
R449 VTAIL.n349 VTAIL.n348 10.4732
R450 VTAIL.n295 VTAIL.n241 10.4732
R451 VTAIL.n271 VTAIL.n270 10.4732
R452 VTAIL.n585 VTAIL.n564 9.69747
R453 VTAIL.n605 VTAIL.n554 9.69747
R454 VTAIL.n39 VTAIL.n18 9.69747
R455 VTAIL.n59 VTAIL.n8 9.69747
R456 VTAIL.n117 VTAIL.n96 9.69747
R457 VTAIL.n137 VTAIL.n86 9.69747
R458 VTAIL.n195 VTAIL.n174 9.69747
R459 VTAIL.n215 VTAIL.n164 9.69747
R460 VTAIL.n528 VTAIL.n477 9.69747
R461 VTAIL.n508 VTAIL.n487 9.69747
R462 VTAIL.n450 VTAIL.n399 9.69747
R463 VTAIL.n430 VTAIL.n409 9.69747
R464 VTAIL.n372 VTAIL.n321 9.69747
R465 VTAIL.n352 VTAIL.n331 9.69747
R466 VTAIL.n294 VTAIL.n243 9.69747
R467 VTAIL.n274 VTAIL.n253 9.69747
R468 VTAIL.n622 VTAIL.n621 9.45567
R469 VTAIL.n76 VTAIL.n75 9.45567
R470 VTAIL.n154 VTAIL.n153 9.45567
R471 VTAIL.n232 VTAIL.n231 9.45567
R472 VTAIL.n544 VTAIL.n543 9.45567
R473 VTAIL.n466 VTAIL.n465 9.45567
R474 VTAIL.n388 VTAIL.n387 9.45567
R475 VTAIL.n310 VTAIL.n309 9.45567
R476 VTAIL.n621 VTAIL.n620 9.3005
R477 VTAIL.n560 VTAIL.n559 9.3005
R478 VTAIL.n589 VTAIL.n588 9.3005
R479 VTAIL.n587 VTAIL.n586 9.3005
R480 VTAIL.n564 VTAIL.n563 9.3005
R481 VTAIL.n581 VTAIL.n580 9.3005
R482 VTAIL.n579 VTAIL.n578 9.3005
R483 VTAIL.n568 VTAIL.n567 9.3005
R484 VTAIL.n573 VTAIL.n572 9.3005
R485 VTAIL.n595 VTAIL.n594 9.3005
R486 VTAIL.n597 VTAIL.n596 9.3005
R487 VTAIL.n556 VTAIL.n555 9.3005
R488 VTAIL.n603 VTAIL.n602 9.3005
R489 VTAIL.n605 VTAIL.n604 9.3005
R490 VTAIL.n552 VTAIL.n551 9.3005
R491 VTAIL.n611 VTAIL.n610 9.3005
R492 VTAIL.n613 VTAIL.n612 9.3005
R493 VTAIL.n614 VTAIL.n547 9.3005
R494 VTAIL.n75 VTAIL.n74 9.3005
R495 VTAIL.n14 VTAIL.n13 9.3005
R496 VTAIL.n43 VTAIL.n42 9.3005
R497 VTAIL.n41 VTAIL.n40 9.3005
R498 VTAIL.n18 VTAIL.n17 9.3005
R499 VTAIL.n35 VTAIL.n34 9.3005
R500 VTAIL.n33 VTAIL.n32 9.3005
R501 VTAIL.n22 VTAIL.n21 9.3005
R502 VTAIL.n27 VTAIL.n26 9.3005
R503 VTAIL.n49 VTAIL.n48 9.3005
R504 VTAIL.n51 VTAIL.n50 9.3005
R505 VTAIL.n10 VTAIL.n9 9.3005
R506 VTAIL.n57 VTAIL.n56 9.3005
R507 VTAIL.n59 VTAIL.n58 9.3005
R508 VTAIL.n6 VTAIL.n5 9.3005
R509 VTAIL.n65 VTAIL.n64 9.3005
R510 VTAIL.n67 VTAIL.n66 9.3005
R511 VTAIL.n68 VTAIL.n1 9.3005
R512 VTAIL.n153 VTAIL.n152 9.3005
R513 VTAIL.n92 VTAIL.n91 9.3005
R514 VTAIL.n121 VTAIL.n120 9.3005
R515 VTAIL.n119 VTAIL.n118 9.3005
R516 VTAIL.n96 VTAIL.n95 9.3005
R517 VTAIL.n113 VTAIL.n112 9.3005
R518 VTAIL.n111 VTAIL.n110 9.3005
R519 VTAIL.n100 VTAIL.n99 9.3005
R520 VTAIL.n105 VTAIL.n104 9.3005
R521 VTAIL.n127 VTAIL.n126 9.3005
R522 VTAIL.n129 VTAIL.n128 9.3005
R523 VTAIL.n88 VTAIL.n87 9.3005
R524 VTAIL.n135 VTAIL.n134 9.3005
R525 VTAIL.n137 VTAIL.n136 9.3005
R526 VTAIL.n84 VTAIL.n83 9.3005
R527 VTAIL.n143 VTAIL.n142 9.3005
R528 VTAIL.n145 VTAIL.n144 9.3005
R529 VTAIL.n146 VTAIL.n79 9.3005
R530 VTAIL.n231 VTAIL.n230 9.3005
R531 VTAIL.n170 VTAIL.n169 9.3005
R532 VTAIL.n199 VTAIL.n198 9.3005
R533 VTAIL.n197 VTAIL.n196 9.3005
R534 VTAIL.n174 VTAIL.n173 9.3005
R535 VTAIL.n191 VTAIL.n190 9.3005
R536 VTAIL.n189 VTAIL.n188 9.3005
R537 VTAIL.n178 VTAIL.n177 9.3005
R538 VTAIL.n183 VTAIL.n182 9.3005
R539 VTAIL.n205 VTAIL.n204 9.3005
R540 VTAIL.n207 VTAIL.n206 9.3005
R541 VTAIL.n166 VTAIL.n165 9.3005
R542 VTAIL.n213 VTAIL.n212 9.3005
R543 VTAIL.n215 VTAIL.n214 9.3005
R544 VTAIL.n162 VTAIL.n161 9.3005
R545 VTAIL.n221 VTAIL.n220 9.3005
R546 VTAIL.n223 VTAIL.n222 9.3005
R547 VTAIL.n224 VTAIL.n157 9.3005
R548 VTAIL.n520 VTAIL.n519 9.3005
R549 VTAIL.n479 VTAIL.n478 9.3005
R550 VTAIL.n526 VTAIL.n525 9.3005
R551 VTAIL.n528 VTAIL.n527 9.3005
R552 VTAIL.n475 VTAIL.n474 9.3005
R553 VTAIL.n534 VTAIL.n533 9.3005
R554 VTAIL.n536 VTAIL.n535 9.3005
R555 VTAIL.n472 VTAIL.n469 9.3005
R556 VTAIL.n543 VTAIL.n542 9.3005
R557 VTAIL.n518 VTAIL.n517 9.3005
R558 VTAIL.n483 VTAIL.n482 9.3005
R559 VTAIL.n512 VTAIL.n511 9.3005
R560 VTAIL.n510 VTAIL.n509 9.3005
R561 VTAIL.n487 VTAIL.n486 9.3005
R562 VTAIL.n504 VTAIL.n503 9.3005
R563 VTAIL.n502 VTAIL.n501 9.3005
R564 VTAIL.n491 VTAIL.n490 9.3005
R565 VTAIL.n496 VTAIL.n495 9.3005
R566 VTAIL.n442 VTAIL.n441 9.3005
R567 VTAIL.n401 VTAIL.n400 9.3005
R568 VTAIL.n448 VTAIL.n447 9.3005
R569 VTAIL.n450 VTAIL.n449 9.3005
R570 VTAIL.n397 VTAIL.n396 9.3005
R571 VTAIL.n456 VTAIL.n455 9.3005
R572 VTAIL.n458 VTAIL.n457 9.3005
R573 VTAIL.n394 VTAIL.n391 9.3005
R574 VTAIL.n465 VTAIL.n464 9.3005
R575 VTAIL.n440 VTAIL.n439 9.3005
R576 VTAIL.n405 VTAIL.n404 9.3005
R577 VTAIL.n434 VTAIL.n433 9.3005
R578 VTAIL.n432 VTAIL.n431 9.3005
R579 VTAIL.n409 VTAIL.n408 9.3005
R580 VTAIL.n426 VTAIL.n425 9.3005
R581 VTAIL.n424 VTAIL.n423 9.3005
R582 VTAIL.n413 VTAIL.n412 9.3005
R583 VTAIL.n418 VTAIL.n417 9.3005
R584 VTAIL.n364 VTAIL.n363 9.3005
R585 VTAIL.n323 VTAIL.n322 9.3005
R586 VTAIL.n370 VTAIL.n369 9.3005
R587 VTAIL.n372 VTAIL.n371 9.3005
R588 VTAIL.n319 VTAIL.n318 9.3005
R589 VTAIL.n378 VTAIL.n377 9.3005
R590 VTAIL.n380 VTAIL.n379 9.3005
R591 VTAIL.n316 VTAIL.n313 9.3005
R592 VTAIL.n387 VTAIL.n386 9.3005
R593 VTAIL.n362 VTAIL.n361 9.3005
R594 VTAIL.n327 VTAIL.n326 9.3005
R595 VTAIL.n356 VTAIL.n355 9.3005
R596 VTAIL.n354 VTAIL.n353 9.3005
R597 VTAIL.n331 VTAIL.n330 9.3005
R598 VTAIL.n348 VTAIL.n347 9.3005
R599 VTAIL.n346 VTAIL.n345 9.3005
R600 VTAIL.n335 VTAIL.n334 9.3005
R601 VTAIL.n340 VTAIL.n339 9.3005
R602 VTAIL.n286 VTAIL.n285 9.3005
R603 VTAIL.n245 VTAIL.n244 9.3005
R604 VTAIL.n292 VTAIL.n291 9.3005
R605 VTAIL.n294 VTAIL.n293 9.3005
R606 VTAIL.n241 VTAIL.n240 9.3005
R607 VTAIL.n300 VTAIL.n299 9.3005
R608 VTAIL.n302 VTAIL.n301 9.3005
R609 VTAIL.n238 VTAIL.n235 9.3005
R610 VTAIL.n309 VTAIL.n308 9.3005
R611 VTAIL.n284 VTAIL.n283 9.3005
R612 VTAIL.n249 VTAIL.n248 9.3005
R613 VTAIL.n278 VTAIL.n277 9.3005
R614 VTAIL.n276 VTAIL.n275 9.3005
R615 VTAIL.n253 VTAIL.n252 9.3005
R616 VTAIL.n270 VTAIL.n269 9.3005
R617 VTAIL.n268 VTAIL.n267 9.3005
R618 VTAIL.n257 VTAIL.n256 9.3005
R619 VTAIL.n262 VTAIL.n261 9.3005
R620 VTAIL.n586 VTAIL.n562 8.92171
R621 VTAIL.n602 VTAIL.n601 8.92171
R622 VTAIL.n40 VTAIL.n16 8.92171
R623 VTAIL.n56 VTAIL.n55 8.92171
R624 VTAIL.n118 VTAIL.n94 8.92171
R625 VTAIL.n134 VTAIL.n133 8.92171
R626 VTAIL.n196 VTAIL.n172 8.92171
R627 VTAIL.n212 VTAIL.n211 8.92171
R628 VTAIL.n525 VTAIL.n524 8.92171
R629 VTAIL.n509 VTAIL.n485 8.92171
R630 VTAIL.n447 VTAIL.n446 8.92171
R631 VTAIL.n431 VTAIL.n407 8.92171
R632 VTAIL.n369 VTAIL.n368 8.92171
R633 VTAIL.n353 VTAIL.n329 8.92171
R634 VTAIL.n291 VTAIL.n290 8.92171
R635 VTAIL.n275 VTAIL.n251 8.92171
R636 VTAIL.n590 VTAIL.n589 8.14595
R637 VTAIL.n598 VTAIL.n556 8.14595
R638 VTAIL.n44 VTAIL.n43 8.14595
R639 VTAIL.n52 VTAIL.n10 8.14595
R640 VTAIL.n122 VTAIL.n121 8.14595
R641 VTAIL.n130 VTAIL.n88 8.14595
R642 VTAIL.n200 VTAIL.n199 8.14595
R643 VTAIL.n208 VTAIL.n166 8.14595
R644 VTAIL.n521 VTAIL.n479 8.14595
R645 VTAIL.n513 VTAIL.n512 8.14595
R646 VTAIL.n443 VTAIL.n401 8.14595
R647 VTAIL.n435 VTAIL.n434 8.14595
R648 VTAIL.n365 VTAIL.n323 8.14595
R649 VTAIL.n357 VTAIL.n356 8.14595
R650 VTAIL.n287 VTAIL.n245 8.14595
R651 VTAIL.n279 VTAIL.n278 8.14595
R652 VTAIL.n593 VTAIL.n560 7.3702
R653 VTAIL.n597 VTAIL.n558 7.3702
R654 VTAIL.n47 VTAIL.n14 7.3702
R655 VTAIL.n51 VTAIL.n12 7.3702
R656 VTAIL.n125 VTAIL.n92 7.3702
R657 VTAIL.n129 VTAIL.n90 7.3702
R658 VTAIL.n203 VTAIL.n170 7.3702
R659 VTAIL.n207 VTAIL.n168 7.3702
R660 VTAIL.n520 VTAIL.n481 7.3702
R661 VTAIL.n516 VTAIL.n483 7.3702
R662 VTAIL.n442 VTAIL.n403 7.3702
R663 VTAIL.n438 VTAIL.n405 7.3702
R664 VTAIL.n364 VTAIL.n325 7.3702
R665 VTAIL.n360 VTAIL.n327 7.3702
R666 VTAIL.n286 VTAIL.n247 7.3702
R667 VTAIL.n282 VTAIL.n249 7.3702
R668 VTAIL.n594 VTAIL.n593 6.59444
R669 VTAIL.n594 VTAIL.n558 6.59444
R670 VTAIL.n48 VTAIL.n47 6.59444
R671 VTAIL.n48 VTAIL.n12 6.59444
R672 VTAIL.n126 VTAIL.n125 6.59444
R673 VTAIL.n126 VTAIL.n90 6.59444
R674 VTAIL.n204 VTAIL.n203 6.59444
R675 VTAIL.n204 VTAIL.n168 6.59444
R676 VTAIL.n517 VTAIL.n481 6.59444
R677 VTAIL.n517 VTAIL.n516 6.59444
R678 VTAIL.n439 VTAIL.n403 6.59444
R679 VTAIL.n439 VTAIL.n438 6.59444
R680 VTAIL.n361 VTAIL.n325 6.59444
R681 VTAIL.n361 VTAIL.n360 6.59444
R682 VTAIL.n283 VTAIL.n247 6.59444
R683 VTAIL.n283 VTAIL.n282 6.59444
R684 VTAIL.n590 VTAIL.n560 5.81868
R685 VTAIL.n598 VTAIL.n597 5.81868
R686 VTAIL.n44 VTAIL.n14 5.81868
R687 VTAIL.n52 VTAIL.n51 5.81868
R688 VTAIL.n122 VTAIL.n92 5.81868
R689 VTAIL.n130 VTAIL.n129 5.81868
R690 VTAIL.n200 VTAIL.n170 5.81868
R691 VTAIL.n208 VTAIL.n207 5.81868
R692 VTAIL.n521 VTAIL.n520 5.81868
R693 VTAIL.n513 VTAIL.n483 5.81868
R694 VTAIL.n443 VTAIL.n442 5.81868
R695 VTAIL.n435 VTAIL.n405 5.81868
R696 VTAIL.n365 VTAIL.n364 5.81868
R697 VTAIL.n357 VTAIL.n327 5.81868
R698 VTAIL.n287 VTAIL.n286 5.81868
R699 VTAIL.n279 VTAIL.n249 5.81868
R700 VTAIL.n589 VTAIL.n562 5.04292
R701 VTAIL.n601 VTAIL.n556 5.04292
R702 VTAIL.n43 VTAIL.n16 5.04292
R703 VTAIL.n55 VTAIL.n10 5.04292
R704 VTAIL.n121 VTAIL.n94 5.04292
R705 VTAIL.n133 VTAIL.n88 5.04292
R706 VTAIL.n199 VTAIL.n172 5.04292
R707 VTAIL.n211 VTAIL.n166 5.04292
R708 VTAIL.n524 VTAIL.n479 5.04292
R709 VTAIL.n512 VTAIL.n485 5.04292
R710 VTAIL.n446 VTAIL.n401 5.04292
R711 VTAIL.n434 VTAIL.n407 5.04292
R712 VTAIL.n368 VTAIL.n323 5.04292
R713 VTAIL.n356 VTAIL.n329 5.04292
R714 VTAIL.n290 VTAIL.n245 5.04292
R715 VTAIL.n278 VTAIL.n251 5.04292
R716 VTAIL.n586 VTAIL.n585 4.26717
R717 VTAIL.n602 VTAIL.n554 4.26717
R718 VTAIL.n40 VTAIL.n39 4.26717
R719 VTAIL.n56 VTAIL.n8 4.26717
R720 VTAIL.n118 VTAIL.n117 4.26717
R721 VTAIL.n134 VTAIL.n86 4.26717
R722 VTAIL.n196 VTAIL.n195 4.26717
R723 VTAIL.n212 VTAIL.n164 4.26717
R724 VTAIL.n525 VTAIL.n477 4.26717
R725 VTAIL.n509 VTAIL.n508 4.26717
R726 VTAIL.n447 VTAIL.n399 4.26717
R727 VTAIL.n431 VTAIL.n430 4.26717
R728 VTAIL.n369 VTAIL.n321 4.26717
R729 VTAIL.n353 VTAIL.n352 4.26717
R730 VTAIL.n291 VTAIL.n243 4.26717
R731 VTAIL.n275 VTAIL.n274 4.26717
R732 VTAIL.n572 VTAIL.n571 3.70982
R733 VTAIL.n26 VTAIL.n25 3.70982
R734 VTAIL.n104 VTAIL.n103 3.70982
R735 VTAIL.n182 VTAIL.n181 3.70982
R736 VTAIL.n495 VTAIL.n494 3.70982
R737 VTAIL.n417 VTAIL.n416 3.70982
R738 VTAIL.n339 VTAIL.n338 3.70982
R739 VTAIL.n261 VTAIL.n260 3.70982
R740 VTAIL.n582 VTAIL.n564 3.49141
R741 VTAIL.n606 VTAIL.n605 3.49141
R742 VTAIL.n36 VTAIL.n18 3.49141
R743 VTAIL.n60 VTAIL.n59 3.49141
R744 VTAIL.n114 VTAIL.n96 3.49141
R745 VTAIL.n138 VTAIL.n137 3.49141
R746 VTAIL.n192 VTAIL.n174 3.49141
R747 VTAIL.n216 VTAIL.n215 3.49141
R748 VTAIL.n529 VTAIL.n528 3.49141
R749 VTAIL.n505 VTAIL.n487 3.49141
R750 VTAIL.n451 VTAIL.n450 3.49141
R751 VTAIL.n427 VTAIL.n409 3.49141
R752 VTAIL.n373 VTAIL.n372 3.49141
R753 VTAIL.n349 VTAIL.n331 3.49141
R754 VTAIL.n295 VTAIL.n294 3.49141
R755 VTAIL.n271 VTAIL.n253 3.49141
R756 VTAIL.n389 VTAIL.n311 3.2936
R757 VTAIL.n545 VTAIL.n467 3.2936
R758 VTAIL.n233 VTAIL.n155 3.2936
R759 VTAIL.n581 VTAIL.n566 2.71565
R760 VTAIL.n609 VTAIL.n552 2.71565
R761 VTAIL.n35 VTAIL.n20 2.71565
R762 VTAIL.n63 VTAIL.n6 2.71565
R763 VTAIL.n113 VTAIL.n98 2.71565
R764 VTAIL.n141 VTAIL.n84 2.71565
R765 VTAIL.n191 VTAIL.n176 2.71565
R766 VTAIL.n219 VTAIL.n162 2.71565
R767 VTAIL.n532 VTAIL.n475 2.71565
R768 VTAIL.n504 VTAIL.n489 2.71565
R769 VTAIL.n454 VTAIL.n397 2.71565
R770 VTAIL.n426 VTAIL.n411 2.71565
R771 VTAIL.n376 VTAIL.n319 2.71565
R772 VTAIL.n348 VTAIL.n333 2.71565
R773 VTAIL.n298 VTAIL.n241 2.71565
R774 VTAIL.n270 VTAIL.n255 2.71565
R775 VTAIL.n578 VTAIL.n577 1.93989
R776 VTAIL.n610 VTAIL.n550 1.93989
R777 VTAIL.n32 VTAIL.n31 1.93989
R778 VTAIL.n64 VTAIL.n4 1.93989
R779 VTAIL.n110 VTAIL.n109 1.93989
R780 VTAIL.n142 VTAIL.n82 1.93989
R781 VTAIL.n188 VTAIL.n187 1.93989
R782 VTAIL.n220 VTAIL.n160 1.93989
R783 VTAIL.n533 VTAIL.n473 1.93989
R784 VTAIL.n501 VTAIL.n500 1.93989
R785 VTAIL.n455 VTAIL.n395 1.93989
R786 VTAIL.n423 VTAIL.n422 1.93989
R787 VTAIL.n377 VTAIL.n317 1.93989
R788 VTAIL.n345 VTAIL.n344 1.93989
R789 VTAIL.n299 VTAIL.n239 1.93989
R790 VTAIL.n267 VTAIL.n266 1.93989
R791 VTAIL VTAIL.n77 1.70524
R792 VTAIL VTAIL.n623 1.58886
R793 VTAIL.n574 VTAIL.n568 1.16414
R794 VTAIL.n615 VTAIL.n613 1.16414
R795 VTAIL.n622 VTAIL.n546 1.16414
R796 VTAIL.n28 VTAIL.n22 1.16414
R797 VTAIL.n69 VTAIL.n67 1.16414
R798 VTAIL.n76 VTAIL.n0 1.16414
R799 VTAIL.n106 VTAIL.n100 1.16414
R800 VTAIL.n147 VTAIL.n145 1.16414
R801 VTAIL.n154 VTAIL.n78 1.16414
R802 VTAIL.n184 VTAIL.n178 1.16414
R803 VTAIL.n225 VTAIL.n223 1.16414
R804 VTAIL.n232 VTAIL.n156 1.16414
R805 VTAIL.n544 VTAIL.n468 1.16414
R806 VTAIL.n537 VTAIL.n536 1.16414
R807 VTAIL.n497 VTAIL.n491 1.16414
R808 VTAIL.n466 VTAIL.n390 1.16414
R809 VTAIL.n459 VTAIL.n458 1.16414
R810 VTAIL.n419 VTAIL.n413 1.16414
R811 VTAIL.n388 VTAIL.n312 1.16414
R812 VTAIL.n381 VTAIL.n380 1.16414
R813 VTAIL.n341 VTAIL.n335 1.16414
R814 VTAIL.n310 VTAIL.n234 1.16414
R815 VTAIL.n303 VTAIL.n302 1.16414
R816 VTAIL.n263 VTAIL.n257 1.16414
R817 VTAIL.n467 VTAIL.n389 0.470328
R818 VTAIL.n155 VTAIL.n77 0.470328
R819 VTAIL.n573 VTAIL.n570 0.388379
R820 VTAIL.n614 VTAIL.n548 0.388379
R821 VTAIL.n620 VTAIL.n619 0.388379
R822 VTAIL.n27 VTAIL.n24 0.388379
R823 VTAIL.n68 VTAIL.n2 0.388379
R824 VTAIL.n74 VTAIL.n73 0.388379
R825 VTAIL.n105 VTAIL.n102 0.388379
R826 VTAIL.n146 VTAIL.n80 0.388379
R827 VTAIL.n152 VTAIL.n151 0.388379
R828 VTAIL.n183 VTAIL.n180 0.388379
R829 VTAIL.n224 VTAIL.n158 0.388379
R830 VTAIL.n230 VTAIL.n229 0.388379
R831 VTAIL.n542 VTAIL.n541 0.388379
R832 VTAIL.n472 VTAIL.n470 0.388379
R833 VTAIL.n496 VTAIL.n493 0.388379
R834 VTAIL.n464 VTAIL.n463 0.388379
R835 VTAIL.n394 VTAIL.n392 0.388379
R836 VTAIL.n418 VTAIL.n415 0.388379
R837 VTAIL.n386 VTAIL.n385 0.388379
R838 VTAIL.n316 VTAIL.n314 0.388379
R839 VTAIL.n340 VTAIL.n337 0.388379
R840 VTAIL.n308 VTAIL.n307 0.388379
R841 VTAIL.n238 VTAIL.n236 0.388379
R842 VTAIL.n262 VTAIL.n259 0.388379
R843 VTAIL.n572 VTAIL.n567 0.155672
R844 VTAIL.n579 VTAIL.n567 0.155672
R845 VTAIL.n580 VTAIL.n579 0.155672
R846 VTAIL.n580 VTAIL.n563 0.155672
R847 VTAIL.n587 VTAIL.n563 0.155672
R848 VTAIL.n588 VTAIL.n587 0.155672
R849 VTAIL.n588 VTAIL.n559 0.155672
R850 VTAIL.n595 VTAIL.n559 0.155672
R851 VTAIL.n596 VTAIL.n595 0.155672
R852 VTAIL.n596 VTAIL.n555 0.155672
R853 VTAIL.n603 VTAIL.n555 0.155672
R854 VTAIL.n604 VTAIL.n603 0.155672
R855 VTAIL.n604 VTAIL.n551 0.155672
R856 VTAIL.n611 VTAIL.n551 0.155672
R857 VTAIL.n612 VTAIL.n611 0.155672
R858 VTAIL.n612 VTAIL.n547 0.155672
R859 VTAIL.n621 VTAIL.n547 0.155672
R860 VTAIL.n26 VTAIL.n21 0.155672
R861 VTAIL.n33 VTAIL.n21 0.155672
R862 VTAIL.n34 VTAIL.n33 0.155672
R863 VTAIL.n34 VTAIL.n17 0.155672
R864 VTAIL.n41 VTAIL.n17 0.155672
R865 VTAIL.n42 VTAIL.n41 0.155672
R866 VTAIL.n42 VTAIL.n13 0.155672
R867 VTAIL.n49 VTAIL.n13 0.155672
R868 VTAIL.n50 VTAIL.n49 0.155672
R869 VTAIL.n50 VTAIL.n9 0.155672
R870 VTAIL.n57 VTAIL.n9 0.155672
R871 VTAIL.n58 VTAIL.n57 0.155672
R872 VTAIL.n58 VTAIL.n5 0.155672
R873 VTAIL.n65 VTAIL.n5 0.155672
R874 VTAIL.n66 VTAIL.n65 0.155672
R875 VTAIL.n66 VTAIL.n1 0.155672
R876 VTAIL.n75 VTAIL.n1 0.155672
R877 VTAIL.n104 VTAIL.n99 0.155672
R878 VTAIL.n111 VTAIL.n99 0.155672
R879 VTAIL.n112 VTAIL.n111 0.155672
R880 VTAIL.n112 VTAIL.n95 0.155672
R881 VTAIL.n119 VTAIL.n95 0.155672
R882 VTAIL.n120 VTAIL.n119 0.155672
R883 VTAIL.n120 VTAIL.n91 0.155672
R884 VTAIL.n127 VTAIL.n91 0.155672
R885 VTAIL.n128 VTAIL.n127 0.155672
R886 VTAIL.n128 VTAIL.n87 0.155672
R887 VTAIL.n135 VTAIL.n87 0.155672
R888 VTAIL.n136 VTAIL.n135 0.155672
R889 VTAIL.n136 VTAIL.n83 0.155672
R890 VTAIL.n143 VTAIL.n83 0.155672
R891 VTAIL.n144 VTAIL.n143 0.155672
R892 VTAIL.n144 VTAIL.n79 0.155672
R893 VTAIL.n153 VTAIL.n79 0.155672
R894 VTAIL.n182 VTAIL.n177 0.155672
R895 VTAIL.n189 VTAIL.n177 0.155672
R896 VTAIL.n190 VTAIL.n189 0.155672
R897 VTAIL.n190 VTAIL.n173 0.155672
R898 VTAIL.n197 VTAIL.n173 0.155672
R899 VTAIL.n198 VTAIL.n197 0.155672
R900 VTAIL.n198 VTAIL.n169 0.155672
R901 VTAIL.n205 VTAIL.n169 0.155672
R902 VTAIL.n206 VTAIL.n205 0.155672
R903 VTAIL.n206 VTAIL.n165 0.155672
R904 VTAIL.n213 VTAIL.n165 0.155672
R905 VTAIL.n214 VTAIL.n213 0.155672
R906 VTAIL.n214 VTAIL.n161 0.155672
R907 VTAIL.n221 VTAIL.n161 0.155672
R908 VTAIL.n222 VTAIL.n221 0.155672
R909 VTAIL.n222 VTAIL.n157 0.155672
R910 VTAIL.n231 VTAIL.n157 0.155672
R911 VTAIL.n543 VTAIL.n469 0.155672
R912 VTAIL.n535 VTAIL.n469 0.155672
R913 VTAIL.n535 VTAIL.n534 0.155672
R914 VTAIL.n534 VTAIL.n474 0.155672
R915 VTAIL.n527 VTAIL.n474 0.155672
R916 VTAIL.n527 VTAIL.n526 0.155672
R917 VTAIL.n526 VTAIL.n478 0.155672
R918 VTAIL.n519 VTAIL.n478 0.155672
R919 VTAIL.n519 VTAIL.n518 0.155672
R920 VTAIL.n518 VTAIL.n482 0.155672
R921 VTAIL.n511 VTAIL.n482 0.155672
R922 VTAIL.n511 VTAIL.n510 0.155672
R923 VTAIL.n510 VTAIL.n486 0.155672
R924 VTAIL.n503 VTAIL.n486 0.155672
R925 VTAIL.n503 VTAIL.n502 0.155672
R926 VTAIL.n502 VTAIL.n490 0.155672
R927 VTAIL.n495 VTAIL.n490 0.155672
R928 VTAIL.n465 VTAIL.n391 0.155672
R929 VTAIL.n457 VTAIL.n391 0.155672
R930 VTAIL.n457 VTAIL.n456 0.155672
R931 VTAIL.n456 VTAIL.n396 0.155672
R932 VTAIL.n449 VTAIL.n396 0.155672
R933 VTAIL.n449 VTAIL.n448 0.155672
R934 VTAIL.n448 VTAIL.n400 0.155672
R935 VTAIL.n441 VTAIL.n400 0.155672
R936 VTAIL.n441 VTAIL.n440 0.155672
R937 VTAIL.n440 VTAIL.n404 0.155672
R938 VTAIL.n433 VTAIL.n404 0.155672
R939 VTAIL.n433 VTAIL.n432 0.155672
R940 VTAIL.n432 VTAIL.n408 0.155672
R941 VTAIL.n425 VTAIL.n408 0.155672
R942 VTAIL.n425 VTAIL.n424 0.155672
R943 VTAIL.n424 VTAIL.n412 0.155672
R944 VTAIL.n417 VTAIL.n412 0.155672
R945 VTAIL.n387 VTAIL.n313 0.155672
R946 VTAIL.n379 VTAIL.n313 0.155672
R947 VTAIL.n379 VTAIL.n378 0.155672
R948 VTAIL.n378 VTAIL.n318 0.155672
R949 VTAIL.n371 VTAIL.n318 0.155672
R950 VTAIL.n371 VTAIL.n370 0.155672
R951 VTAIL.n370 VTAIL.n322 0.155672
R952 VTAIL.n363 VTAIL.n322 0.155672
R953 VTAIL.n363 VTAIL.n362 0.155672
R954 VTAIL.n362 VTAIL.n326 0.155672
R955 VTAIL.n355 VTAIL.n326 0.155672
R956 VTAIL.n355 VTAIL.n354 0.155672
R957 VTAIL.n354 VTAIL.n330 0.155672
R958 VTAIL.n347 VTAIL.n330 0.155672
R959 VTAIL.n347 VTAIL.n346 0.155672
R960 VTAIL.n346 VTAIL.n334 0.155672
R961 VTAIL.n339 VTAIL.n334 0.155672
R962 VTAIL.n309 VTAIL.n235 0.155672
R963 VTAIL.n301 VTAIL.n235 0.155672
R964 VTAIL.n301 VTAIL.n300 0.155672
R965 VTAIL.n300 VTAIL.n240 0.155672
R966 VTAIL.n293 VTAIL.n240 0.155672
R967 VTAIL.n293 VTAIL.n292 0.155672
R968 VTAIL.n292 VTAIL.n244 0.155672
R969 VTAIL.n285 VTAIL.n244 0.155672
R970 VTAIL.n285 VTAIL.n284 0.155672
R971 VTAIL.n284 VTAIL.n248 0.155672
R972 VTAIL.n277 VTAIL.n248 0.155672
R973 VTAIL.n277 VTAIL.n276 0.155672
R974 VTAIL.n276 VTAIL.n252 0.155672
R975 VTAIL.n269 VTAIL.n252 0.155672
R976 VTAIL.n269 VTAIL.n268 0.155672
R977 VTAIL.n268 VTAIL.n256 0.155672
R978 VTAIL.n261 VTAIL.n256 0.155672
R979 VDD1 VDD1.n1 120.087
R980 VDD1 VDD1.n0 73.9135
R981 VDD1.n0 VDD1.t2 2.31402
R982 VDD1.n0 VDD1.t3 2.31402
R983 VDD1.n1 VDD1.t0 2.31402
R984 VDD1.n1 VDD1.t1 2.31402
R985 VN.n1 VN.t1 131.413
R986 VN.n0 VN.t2 131.413
R987 VN.n0 VN.t0 130.196
R988 VN.n1 VN.t3 130.196
R989 VN VN.n1 52.9877
R990 VN VN.n0 2.21123
R991 VDD2.n2 VDD2.n0 119.561
R992 VDD2.n2 VDD2.n1 73.8553
R993 VDD2.n1 VDD2.t0 2.31402
R994 VDD2.n1 VDD2.t2 2.31402
R995 VDD2.n0 VDD2.t1 2.31402
R996 VDD2.n0 VDD2.t3 2.31402
R997 VDD2 VDD2.n2 0.0586897
R998 B.n548 B.n79 585
R999 B.n550 B.n549 585
R1000 B.n551 B.n78 585
R1001 B.n553 B.n552 585
R1002 B.n554 B.n77 585
R1003 B.n556 B.n555 585
R1004 B.n557 B.n76 585
R1005 B.n559 B.n558 585
R1006 B.n560 B.n75 585
R1007 B.n562 B.n561 585
R1008 B.n563 B.n74 585
R1009 B.n565 B.n564 585
R1010 B.n566 B.n73 585
R1011 B.n568 B.n567 585
R1012 B.n569 B.n72 585
R1013 B.n571 B.n570 585
R1014 B.n572 B.n71 585
R1015 B.n574 B.n573 585
R1016 B.n575 B.n70 585
R1017 B.n577 B.n576 585
R1018 B.n578 B.n69 585
R1019 B.n580 B.n579 585
R1020 B.n581 B.n68 585
R1021 B.n583 B.n582 585
R1022 B.n584 B.n67 585
R1023 B.n586 B.n585 585
R1024 B.n587 B.n66 585
R1025 B.n589 B.n588 585
R1026 B.n590 B.n65 585
R1027 B.n592 B.n591 585
R1028 B.n593 B.n64 585
R1029 B.n595 B.n594 585
R1030 B.n596 B.n63 585
R1031 B.n598 B.n597 585
R1032 B.n599 B.n62 585
R1033 B.n601 B.n600 585
R1034 B.n602 B.n61 585
R1035 B.n604 B.n603 585
R1036 B.n605 B.n60 585
R1037 B.n607 B.n606 585
R1038 B.n608 B.n59 585
R1039 B.n610 B.n609 585
R1040 B.n611 B.n58 585
R1041 B.n613 B.n612 585
R1042 B.n614 B.n57 585
R1043 B.n616 B.n615 585
R1044 B.n617 B.n56 585
R1045 B.n619 B.n618 585
R1046 B.n621 B.n53 585
R1047 B.n623 B.n622 585
R1048 B.n624 B.n52 585
R1049 B.n626 B.n625 585
R1050 B.n627 B.n51 585
R1051 B.n629 B.n628 585
R1052 B.n630 B.n50 585
R1053 B.n632 B.n631 585
R1054 B.n633 B.n47 585
R1055 B.n636 B.n635 585
R1056 B.n637 B.n46 585
R1057 B.n639 B.n638 585
R1058 B.n640 B.n45 585
R1059 B.n642 B.n641 585
R1060 B.n643 B.n44 585
R1061 B.n645 B.n644 585
R1062 B.n646 B.n43 585
R1063 B.n648 B.n647 585
R1064 B.n649 B.n42 585
R1065 B.n651 B.n650 585
R1066 B.n652 B.n41 585
R1067 B.n654 B.n653 585
R1068 B.n655 B.n40 585
R1069 B.n657 B.n656 585
R1070 B.n658 B.n39 585
R1071 B.n660 B.n659 585
R1072 B.n661 B.n38 585
R1073 B.n663 B.n662 585
R1074 B.n664 B.n37 585
R1075 B.n666 B.n665 585
R1076 B.n667 B.n36 585
R1077 B.n669 B.n668 585
R1078 B.n670 B.n35 585
R1079 B.n672 B.n671 585
R1080 B.n673 B.n34 585
R1081 B.n675 B.n674 585
R1082 B.n676 B.n33 585
R1083 B.n678 B.n677 585
R1084 B.n679 B.n32 585
R1085 B.n681 B.n680 585
R1086 B.n682 B.n31 585
R1087 B.n684 B.n683 585
R1088 B.n685 B.n30 585
R1089 B.n687 B.n686 585
R1090 B.n688 B.n29 585
R1091 B.n690 B.n689 585
R1092 B.n691 B.n28 585
R1093 B.n693 B.n692 585
R1094 B.n694 B.n27 585
R1095 B.n696 B.n695 585
R1096 B.n697 B.n26 585
R1097 B.n699 B.n698 585
R1098 B.n700 B.n25 585
R1099 B.n702 B.n701 585
R1100 B.n703 B.n24 585
R1101 B.n705 B.n704 585
R1102 B.n706 B.n23 585
R1103 B.n547 B.n546 585
R1104 B.n545 B.n80 585
R1105 B.n544 B.n543 585
R1106 B.n542 B.n81 585
R1107 B.n541 B.n540 585
R1108 B.n539 B.n82 585
R1109 B.n538 B.n537 585
R1110 B.n536 B.n83 585
R1111 B.n535 B.n534 585
R1112 B.n533 B.n84 585
R1113 B.n532 B.n531 585
R1114 B.n530 B.n85 585
R1115 B.n529 B.n528 585
R1116 B.n527 B.n86 585
R1117 B.n526 B.n525 585
R1118 B.n524 B.n87 585
R1119 B.n523 B.n522 585
R1120 B.n521 B.n88 585
R1121 B.n520 B.n519 585
R1122 B.n518 B.n89 585
R1123 B.n517 B.n516 585
R1124 B.n515 B.n90 585
R1125 B.n514 B.n513 585
R1126 B.n512 B.n91 585
R1127 B.n511 B.n510 585
R1128 B.n509 B.n92 585
R1129 B.n508 B.n507 585
R1130 B.n506 B.n93 585
R1131 B.n505 B.n504 585
R1132 B.n503 B.n94 585
R1133 B.n502 B.n501 585
R1134 B.n500 B.n95 585
R1135 B.n499 B.n498 585
R1136 B.n497 B.n96 585
R1137 B.n496 B.n495 585
R1138 B.n494 B.n97 585
R1139 B.n493 B.n492 585
R1140 B.n491 B.n98 585
R1141 B.n490 B.n489 585
R1142 B.n488 B.n99 585
R1143 B.n487 B.n486 585
R1144 B.n485 B.n100 585
R1145 B.n484 B.n483 585
R1146 B.n482 B.n101 585
R1147 B.n481 B.n480 585
R1148 B.n479 B.n102 585
R1149 B.n478 B.n477 585
R1150 B.n476 B.n103 585
R1151 B.n475 B.n474 585
R1152 B.n473 B.n104 585
R1153 B.n472 B.n471 585
R1154 B.n470 B.n105 585
R1155 B.n469 B.n468 585
R1156 B.n467 B.n106 585
R1157 B.n466 B.n465 585
R1158 B.n464 B.n107 585
R1159 B.n463 B.n462 585
R1160 B.n461 B.n108 585
R1161 B.n460 B.n459 585
R1162 B.n458 B.n109 585
R1163 B.n457 B.n456 585
R1164 B.n455 B.n110 585
R1165 B.n454 B.n453 585
R1166 B.n452 B.n111 585
R1167 B.n451 B.n450 585
R1168 B.n449 B.n112 585
R1169 B.n448 B.n447 585
R1170 B.n446 B.n113 585
R1171 B.n445 B.n444 585
R1172 B.n443 B.n114 585
R1173 B.n442 B.n441 585
R1174 B.n440 B.n115 585
R1175 B.n439 B.n438 585
R1176 B.n437 B.n116 585
R1177 B.n436 B.n435 585
R1178 B.n434 B.n117 585
R1179 B.n433 B.n432 585
R1180 B.n431 B.n118 585
R1181 B.n430 B.n429 585
R1182 B.n428 B.n119 585
R1183 B.n427 B.n426 585
R1184 B.n425 B.n120 585
R1185 B.n424 B.n423 585
R1186 B.n422 B.n121 585
R1187 B.n421 B.n420 585
R1188 B.n262 B.n261 585
R1189 B.n263 B.n178 585
R1190 B.n265 B.n264 585
R1191 B.n266 B.n177 585
R1192 B.n268 B.n267 585
R1193 B.n269 B.n176 585
R1194 B.n271 B.n270 585
R1195 B.n272 B.n175 585
R1196 B.n274 B.n273 585
R1197 B.n275 B.n174 585
R1198 B.n277 B.n276 585
R1199 B.n278 B.n173 585
R1200 B.n280 B.n279 585
R1201 B.n281 B.n172 585
R1202 B.n283 B.n282 585
R1203 B.n284 B.n171 585
R1204 B.n286 B.n285 585
R1205 B.n287 B.n170 585
R1206 B.n289 B.n288 585
R1207 B.n290 B.n169 585
R1208 B.n292 B.n291 585
R1209 B.n293 B.n168 585
R1210 B.n295 B.n294 585
R1211 B.n296 B.n167 585
R1212 B.n298 B.n297 585
R1213 B.n299 B.n166 585
R1214 B.n301 B.n300 585
R1215 B.n302 B.n165 585
R1216 B.n304 B.n303 585
R1217 B.n305 B.n164 585
R1218 B.n307 B.n306 585
R1219 B.n308 B.n163 585
R1220 B.n310 B.n309 585
R1221 B.n311 B.n162 585
R1222 B.n313 B.n312 585
R1223 B.n314 B.n161 585
R1224 B.n316 B.n315 585
R1225 B.n317 B.n160 585
R1226 B.n319 B.n318 585
R1227 B.n320 B.n159 585
R1228 B.n322 B.n321 585
R1229 B.n323 B.n158 585
R1230 B.n325 B.n324 585
R1231 B.n326 B.n157 585
R1232 B.n328 B.n327 585
R1233 B.n329 B.n156 585
R1234 B.n331 B.n330 585
R1235 B.n332 B.n153 585
R1236 B.n335 B.n334 585
R1237 B.n336 B.n152 585
R1238 B.n338 B.n337 585
R1239 B.n339 B.n151 585
R1240 B.n341 B.n340 585
R1241 B.n342 B.n150 585
R1242 B.n344 B.n343 585
R1243 B.n345 B.n149 585
R1244 B.n347 B.n346 585
R1245 B.n349 B.n348 585
R1246 B.n350 B.n145 585
R1247 B.n352 B.n351 585
R1248 B.n353 B.n144 585
R1249 B.n355 B.n354 585
R1250 B.n356 B.n143 585
R1251 B.n358 B.n357 585
R1252 B.n359 B.n142 585
R1253 B.n361 B.n360 585
R1254 B.n362 B.n141 585
R1255 B.n364 B.n363 585
R1256 B.n365 B.n140 585
R1257 B.n367 B.n366 585
R1258 B.n368 B.n139 585
R1259 B.n370 B.n369 585
R1260 B.n371 B.n138 585
R1261 B.n373 B.n372 585
R1262 B.n374 B.n137 585
R1263 B.n376 B.n375 585
R1264 B.n377 B.n136 585
R1265 B.n379 B.n378 585
R1266 B.n380 B.n135 585
R1267 B.n382 B.n381 585
R1268 B.n383 B.n134 585
R1269 B.n385 B.n384 585
R1270 B.n386 B.n133 585
R1271 B.n388 B.n387 585
R1272 B.n389 B.n132 585
R1273 B.n391 B.n390 585
R1274 B.n392 B.n131 585
R1275 B.n394 B.n393 585
R1276 B.n395 B.n130 585
R1277 B.n397 B.n396 585
R1278 B.n398 B.n129 585
R1279 B.n400 B.n399 585
R1280 B.n401 B.n128 585
R1281 B.n403 B.n402 585
R1282 B.n404 B.n127 585
R1283 B.n406 B.n405 585
R1284 B.n407 B.n126 585
R1285 B.n409 B.n408 585
R1286 B.n410 B.n125 585
R1287 B.n412 B.n411 585
R1288 B.n413 B.n124 585
R1289 B.n415 B.n414 585
R1290 B.n416 B.n123 585
R1291 B.n418 B.n417 585
R1292 B.n419 B.n122 585
R1293 B.n260 B.n179 585
R1294 B.n259 B.n258 585
R1295 B.n257 B.n180 585
R1296 B.n256 B.n255 585
R1297 B.n254 B.n181 585
R1298 B.n253 B.n252 585
R1299 B.n251 B.n182 585
R1300 B.n250 B.n249 585
R1301 B.n248 B.n183 585
R1302 B.n247 B.n246 585
R1303 B.n245 B.n184 585
R1304 B.n244 B.n243 585
R1305 B.n242 B.n185 585
R1306 B.n241 B.n240 585
R1307 B.n239 B.n186 585
R1308 B.n238 B.n237 585
R1309 B.n236 B.n187 585
R1310 B.n235 B.n234 585
R1311 B.n233 B.n188 585
R1312 B.n232 B.n231 585
R1313 B.n230 B.n189 585
R1314 B.n229 B.n228 585
R1315 B.n227 B.n190 585
R1316 B.n226 B.n225 585
R1317 B.n224 B.n191 585
R1318 B.n223 B.n222 585
R1319 B.n221 B.n192 585
R1320 B.n220 B.n219 585
R1321 B.n218 B.n193 585
R1322 B.n217 B.n216 585
R1323 B.n215 B.n194 585
R1324 B.n214 B.n213 585
R1325 B.n212 B.n195 585
R1326 B.n211 B.n210 585
R1327 B.n209 B.n196 585
R1328 B.n208 B.n207 585
R1329 B.n206 B.n197 585
R1330 B.n205 B.n204 585
R1331 B.n203 B.n198 585
R1332 B.n202 B.n201 585
R1333 B.n200 B.n199 585
R1334 B.n2 B.n0 585
R1335 B.n769 B.n1 585
R1336 B.n768 B.n767 585
R1337 B.n766 B.n3 585
R1338 B.n765 B.n764 585
R1339 B.n763 B.n4 585
R1340 B.n762 B.n761 585
R1341 B.n760 B.n5 585
R1342 B.n759 B.n758 585
R1343 B.n757 B.n6 585
R1344 B.n756 B.n755 585
R1345 B.n754 B.n7 585
R1346 B.n753 B.n752 585
R1347 B.n751 B.n8 585
R1348 B.n750 B.n749 585
R1349 B.n748 B.n9 585
R1350 B.n747 B.n746 585
R1351 B.n745 B.n10 585
R1352 B.n744 B.n743 585
R1353 B.n742 B.n11 585
R1354 B.n741 B.n740 585
R1355 B.n739 B.n12 585
R1356 B.n738 B.n737 585
R1357 B.n736 B.n13 585
R1358 B.n735 B.n734 585
R1359 B.n733 B.n14 585
R1360 B.n732 B.n731 585
R1361 B.n730 B.n15 585
R1362 B.n729 B.n728 585
R1363 B.n727 B.n16 585
R1364 B.n726 B.n725 585
R1365 B.n724 B.n17 585
R1366 B.n723 B.n722 585
R1367 B.n721 B.n18 585
R1368 B.n720 B.n719 585
R1369 B.n718 B.n19 585
R1370 B.n717 B.n716 585
R1371 B.n715 B.n20 585
R1372 B.n714 B.n713 585
R1373 B.n712 B.n21 585
R1374 B.n711 B.n710 585
R1375 B.n709 B.n22 585
R1376 B.n708 B.n707 585
R1377 B.n771 B.n770 585
R1378 B.n146 B.t11 486.55
R1379 B.n54 B.t1 486.55
R1380 B.n154 B.t8 486.55
R1381 B.n48 B.t4 486.55
R1382 B.n262 B.n179 458.866
R1383 B.n708 B.n23 458.866
R1384 B.n420 B.n419 458.866
R1385 B.n546 B.n79 458.866
R1386 B.n147 B.t10 412.466
R1387 B.n55 B.t2 412.466
R1388 B.n155 B.t7 412.466
R1389 B.n49 B.t5 412.466
R1390 B.n146 B.t9 306.106
R1391 B.n154 B.t6 306.106
R1392 B.n48 B.t3 306.106
R1393 B.n54 B.t0 306.106
R1394 B.n258 B.n179 163.367
R1395 B.n258 B.n257 163.367
R1396 B.n257 B.n256 163.367
R1397 B.n256 B.n181 163.367
R1398 B.n252 B.n181 163.367
R1399 B.n252 B.n251 163.367
R1400 B.n251 B.n250 163.367
R1401 B.n250 B.n183 163.367
R1402 B.n246 B.n183 163.367
R1403 B.n246 B.n245 163.367
R1404 B.n245 B.n244 163.367
R1405 B.n244 B.n185 163.367
R1406 B.n240 B.n185 163.367
R1407 B.n240 B.n239 163.367
R1408 B.n239 B.n238 163.367
R1409 B.n238 B.n187 163.367
R1410 B.n234 B.n187 163.367
R1411 B.n234 B.n233 163.367
R1412 B.n233 B.n232 163.367
R1413 B.n232 B.n189 163.367
R1414 B.n228 B.n189 163.367
R1415 B.n228 B.n227 163.367
R1416 B.n227 B.n226 163.367
R1417 B.n226 B.n191 163.367
R1418 B.n222 B.n191 163.367
R1419 B.n222 B.n221 163.367
R1420 B.n221 B.n220 163.367
R1421 B.n220 B.n193 163.367
R1422 B.n216 B.n193 163.367
R1423 B.n216 B.n215 163.367
R1424 B.n215 B.n214 163.367
R1425 B.n214 B.n195 163.367
R1426 B.n210 B.n195 163.367
R1427 B.n210 B.n209 163.367
R1428 B.n209 B.n208 163.367
R1429 B.n208 B.n197 163.367
R1430 B.n204 B.n197 163.367
R1431 B.n204 B.n203 163.367
R1432 B.n203 B.n202 163.367
R1433 B.n202 B.n199 163.367
R1434 B.n199 B.n2 163.367
R1435 B.n770 B.n2 163.367
R1436 B.n770 B.n769 163.367
R1437 B.n769 B.n768 163.367
R1438 B.n768 B.n3 163.367
R1439 B.n764 B.n3 163.367
R1440 B.n764 B.n763 163.367
R1441 B.n763 B.n762 163.367
R1442 B.n762 B.n5 163.367
R1443 B.n758 B.n5 163.367
R1444 B.n758 B.n757 163.367
R1445 B.n757 B.n756 163.367
R1446 B.n756 B.n7 163.367
R1447 B.n752 B.n7 163.367
R1448 B.n752 B.n751 163.367
R1449 B.n751 B.n750 163.367
R1450 B.n750 B.n9 163.367
R1451 B.n746 B.n9 163.367
R1452 B.n746 B.n745 163.367
R1453 B.n745 B.n744 163.367
R1454 B.n744 B.n11 163.367
R1455 B.n740 B.n11 163.367
R1456 B.n740 B.n739 163.367
R1457 B.n739 B.n738 163.367
R1458 B.n738 B.n13 163.367
R1459 B.n734 B.n13 163.367
R1460 B.n734 B.n733 163.367
R1461 B.n733 B.n732 163.367
R1462 B.n732 B.n15 163.367
R1463 B.n728 B.n15 163.367
R1464 B.n728 B.n727 163.367
R1465 B.n727 B.n726 163.367
R1466 B.n726 B.n17 163.367
R1467 B.n722 B.n17 163.367
R1468 B.n722 B.n721 163.367
R1469 B.n721 B.n720 163.367
R1470 B.n720 B.n19 163.367
R1471 B.n716 B.n19 163.367
R1472 B.n716 B.n715 163.367
R1473 B.n715 B.n714 163.367
R1474 B.n714 B.n21 163.367
R1475 B.n710 B.n21 163.367
R1476 B.n710 B.n709 163.367
R1477 B.n709 B.n708 163.367
R1478 B.n263 B.n262 163.367
R1479 B.n264 B.n263 163.367
R1480 B.n264 B.n177 163.367
R1481 B.n268 B.n177 163.367
R1482 B.n269 B.n268 163.367
R1483 B.n270 B.n269 163.367
R1484 B.n270 B.n175 163.367
R1485 B.n274 B.n175 163.367
R1486 B.n275 B.n274 163.367
R1487 B.n276 B.n275 163.367
R1488 B.n276 B.n173 163.367
R1489 B.n280 B.n173 163.367
R1490 B.n281 B.n280 163.367
R1491 B.n282 B.n281 163.367
R1492 B.n282 B.n171 163.367
R1493 B.n286 B.n171 163.367
R1494 B.n287 B.n286 163.367
R1495 B.n288 B.n287 163.367
R1496 B.n288 B.n169 163.367
R1497 B.n292 B.n169 163.367
R1498 B.n293 B.n292 163.367
R1499 B.n294 B.n293 163.367
R1500 B.n294 B.n167 163.367
R1501 B.n298 B.n167 163.367
R1502 B.n299 B.n298 163.367
R1503 B.n300 B.n299 163.367
R1504 B.n300 B.n165 163.367
R1505 B.n304 B.n165 163.367
R1506 B.n305 B.n304 163.367
R1507 B.n306 B.n305 163.367
R1508 B.n306 B.n163 163.367
R1509 B.n310 B.n163 163.367
R1510 B.n311 B.n310 163.367
R1511 B.n312 B.n311 163.367
R1512 B.n312 B.n161 163.367
R1513 B.n316 B.n161 163.367
R1514 B.n317 B.n316 163.367
R1515 B.n318 B.n317 163.367
R1516 B.n318 B.n159 163.367
R1517 B.n322 B.n159 163.367
R1518 B.n323 B.n322 163.367
R1519 B.n324 B.n323 163.367
R1520 B.n324 B.n157 163.367
R1521 B.n328 B.n157 163.367
R1522 B.n329 B.n328 163.367
R1523 B.n330 B.n329 163.367
R1524 B.n330 B.n153 163.367
R1525 B.n335 B.n153 163.367
R1526 B.n336 B.n335 163.367
R1527 B.n337 B.n336 163.367
R1528 B.n337 B.n151 163.367
R1529 B.n341 B.n151 163.367
R1530 B.n342 B.n341 163.367
R1531 B.n343 B.n342 163.367
R1532 B.n343 B.n149 163.367
R1533 B.n347 B.n149 163.367
R1534 B.n348 B.n347 163.367
R1535 B.n348 B.n145 163.367
R1536 B.n352 B.n145 163.367
R1537 B.n353 B.n352 163.367
R1538 B.n354 B.n353 163.367
R1539 B.n354 B.n143 163.367
R1540 B.n358 B.n143 163.367
R1541 B.n359 B.n358 163.367
R1542 B.n360 B.n359 163.367
R1543 B.n360 B.n141 163.367
R1544 B.n364 B.n141 163.367
R1545 B.n365 B.n364 163.367
R1546 B.n366 B.n365 163.367
R1547 B.n366 B.n139 163.367
R1548 B.n370 B.n139 163.367
R1549 B.n371 B.n370 163.367
R1550 B.n372 B.n371 163.367
R1551 B.n372 B.n137 163.367
R1552 B.n376 B.n137 163.367
R1553 B.n377 B.n376 163.367
R1554 B.n378 B.n377 163.367
R1555 B.n378 B.n135 163.367
R1556 B.n382 B.n135 163.367
R1557 B.n383 B.n382 163.367
R1558 B.n384 B.n383 163.367
R1559 B.n384 B.n133 163.367
R1560 B.n388 B.n133 163.367
R1561 B.n389 B.n388 163.367
R1562 B.n390 B.n389 163.367
R1563 B.n390 B.n131 163.367
R1564 B.n394 B.n131 163.367
R1565 B.n395 B.n394 163.367
R1566 B.n396 B.n395 163.367
R1567 B.n396 B.n129 163.367
R1568 B.n400 B.n129 163.367
R1569 B.n401 B.n400 163.367
R1570 B.n402 B.n401 163.367
R1571 B.n402 B.n127 163.367
R1572 B.n406 B.n127 163.367
R1573 B.n407 B.n406 163.367
R1574 B.n408 B.n407 163.367
R1575 B.n408 B.n125 163.367
R1576 B.n412 B.n125 163.367
R1577 B.n413 B.n412 163.367
R1578 B.n414 B.n413 163.367
R1579 B.n414 B.n123 163.367
R1580 B.n418 B.n123 163.367
R1581 B.n419 B.n418 163.367
R1582 B.n420 B.n121 163.367
R1583 B.n424 B.n121 163.367
R1584 B.n425 B.n424 163.367
R1585 B.n426 B.n425 163.367
R1586 B.n426 B.n119 163.367
R1587 B.n430 B.n119 163.367
R1588 B.n431 B.n430 163.367
R1589 B.n432 B.n431 163.367
R1590 B.n432 B.n117 163.367
R1591 B.n436 B.n117 163.367
R1592 B.n437 B.n436 163.367
R1593 B.n438 B.n437 163.367
R1594 B.n438 B.n115 163.367
R1595 B.n442 B.n115 163.367
R1596 B.n443 B.n442 163.367
R1597 B.n444 B.n443 163.367
R1598 B.n444 B.n113 163.367
R1599 B.n448 B.n113 163.367
R1600 B.n449 B.n448 163.367
R1601 B.n450 B.n449 163.367
R1602 B.n450 B.n111 163.367
R1603 B.n454 B.n111 163.367
R1604 B.n455 B.n454 163.367
R1605 B.n456 B.n455 163.367
R1606 B.n456 B.n109 163.367
R1607 B.n460 B.n109 163.367
R1608 B.n461 B.n460 163.367
R1609 B.n462 B.n461 163.367
R1610 B.n462 B.n107 163.367
R1611 B.n466 B.n107 163.367
R1612 B.n467 B.n466 163.367
R1613 B.n468 B.n467 163.367
R1614 B.n468 B.n105 163.367
R1615 B.n472 B.n105 163.367
R1616 B.n473 B.n472 163.367
R1617 B.n474 B.n473 163.367
R1618 B.n474 B.n103 163.367
R1619 B.n478 B.n103 163.367
R1620 B.n479 B.n478 163.367
R1621 B.n480 B.n479 163.367
R1622 B.n480 B.n101 163.367
R1623 B.n484 B.n101 163.367
R1624 B.n485 B.n484 163.367
R1625 B.n486 B.n485 163.367
R1626 B.n486 B.n99 163.367
R1627 B.n490 B.n99 163.367
R1628 B.n491 B.n490 163.367
R1629 B.n492 B.n491 163.367
R1630 B.n492 B.n97 163.367
R1631 B.n496 B.n97 163.367
R1632 B.n497 B.n496 163.367
R1633 B.n498 B.n497 163.367
R1634 B.n498 B.n95 163.367
R1635 B.n502 B.n95 163.367
R1636 B.n503 B.n502 163.367
R1637 B.n504 B.n503 163.367
R1638 B.n504 B.n93 163.367
R1639 B.n508 B.n93 163.367
R1640 B.n509 B.n508 163.367
R1641 B.n510 B.n509 163.367
R1642 B.n510 B.n91 163.367
R1643 B.n514 B.n91 163.367
R1644 B.n515 B.n514 163.367
R1645 B.n516 B.n515 163.367
R1646 B.n516 B.n89 163.367
R1647 B.n520 B.n89 163.367
R1648 B.n521 B.n520 163.367
R1649 B.n522 B.n521 163.367
R1650 B.n522 B.n87 163.367
R1651 B.n526 B.n87 163.367
R1652 B.n527 B.n526 163.367
R1653 B.n528 B.n527 163.367
R1654 B.n528 B.n85 163.367
R1655 B.n532 B.n85 163.367
R1656 B.n533 B.n532 163.367
R1657 B.n534 B.n533 163.367
R1658 B.n534 B.n83 163.367
R1659 B.n538 B.n83 163.367
R1660 B.n539 B.n538 163.367
R1661 B.n540 B.n539 163.367
R1662 B.n540 B.n81 163.367
R1663 B.n544 B.n81 163.367
R1664 B.n545 B.n544 163.367
R1665 B.n546 B.n545 163.367
R1666 B.n704 B.n23 163.367
R1667 B.n704 B.n703 163.367
R1668 B.n703 B.n702 163.367
R1669 B.n702 B.n25 163.367
R1670 B.n698 B.n25 163.367
R1671 B.n698 B.n697 163.367
R1672 B.n697 B.n696 163.367
R1673 B.n696 B.n27 163.367
R1674 B.n692 B.n27 163.367
R1675 B.n692 B.n691 163.367
R1676 B.n691 B.n690 163.367
R1677 B.n690 B.n29 163.367
R1678 B.n686 B.n29 163.367
R1679 B.n686 B.n685 163.367
R1680 B.n685 B.n684 163.367
R1681 B.n684 B.n31 163.367
R1682 B.n680 B.n31 163.367
R1683 B.n680 B.n679 163.367
R1684 B.n679 B.n678 163.367
R1685 B.n678 B.n33 163.367
R1686 B.n674 B.n33 163.367
R1687 B.n674 B.n673 163.367
R1688 B.n673 B.n672 163.367
R1689 B.n672 B.n35 163.367
R1690 B.n668 B.n35 163.367
R1691 B.n668 B.n667 163.367
R1692 B.n667 B.n666 163.367
R1693 B.n666 B.n37 163.367
R1694 B.n662 B.n37 163.367
R1695 B.n662 B.n661 163.367
R1696 B.n661 B.n660 163.367
R1697 B.n660 B.n39 163.367
R1698 B.n656 B.n39 163.367
R1699 B.n656 B.n655 163.367
R1700 B.n655 B.n654 163.367
R1701 B.n654 B.n41 163.367
R1702 B.n650 B.n41 163.367
R1703 B.n650 B.n649 163.367
R1704 B.n649 B.n648 163.367
R1705 B.n648 B.n43 163.367
R1706 B.n644 B.n43 163.367
R1707 B.n644 B.n643 163.367
R1708 B.n643 B.n642 163.367
R1709 B.n642 B.n45 163.367
R1710 B.n638 B.n45 163.367
R1711 B.n638 B.n637 163.367
R1712 B.n637 B.n636 163.367
R1713 B.n636 B.n47 163.367
R1714 B.n631 B.n47 163.367
R1715 B.n631 B.n630 163.367
R1716 B.n630 B.n629 163.367
R1717 B.n629 B.n51 163.367
R1718 B.n625 B.n51 163.367
R1719 B.n625 B.n624 163.367
R1720 B.n624 B.n623 163.367
R1721 B.n623 B.n53 163.367
R1722 B.n618 B.n53 163.367
R1723 B.n618 B.n617 163.367
R1724 B.n617 B.n616 163.367
R1725 B.n616 B.n57 163.367
R1726 B.n612 B.n57 163.367
R1727 B.n612 B.n611 163.367
R1728 B.n611 B.n610 163.367
R1729 B.n610 B.n59 163.367
R1730 B.n606 B.n59 163.367
R1731 B.n606 B.n605 163.367
R1732 B.n605 B.n604 163.367
R1733 B.n604 B.n61 163.367
R1734 B.n600 B.n61 163.367
R1735 B.n600 B.n599 163.367
R1736 B.n599 B.n598 163.367
R1737 B.n598 B.n63 163.367
R1738 B.n594 B.n63 163.367
R1739 B.n594 B.n593 163.367
R1740 B.n593 B.n592 163.367
R1741 B.n592 B.n65 163.367
R1742 B.n588 B.n65 163.367
R1743 B.n588 B.n587 163.367
R1744 B.n587 B.n586 163.367
R1745 B.n586 B.n67 163.367
R1746 B.n582 B.n67 163.367
R1747 B.n582 B.n581 163.367
R1748 B.n581 B.n580 163.367
R1749 B.n580 B.n69 163.367
R1750 B.n576 B.n69 163.367
R1751 B.n576 B.n575 163.367
R1752 B.n575 B.n574 163.367
R1753 B.n574 B.n71 163.367
R1754 B.n570 B.n71 163.367
R1755 B.n570 B.n569 163.367
R1756 B.n569 B.n568 163.367
R1757 B.n568 B.n73 163.367
R1758 B.n564 B.n73 163.367
R1759 B.n564 B.n563 163.367
R1760 B.n563 B.n562 163.367
R1761 B.n562 B.n75 163.367
R1762 B.n558 B.n75 163.367
R1763 B.n558 B.n557 163.367
R1764 B.n557 B.n556 163.367
R1765 B.n556 B.n77 163.367
R1766 B.n552 B.n77 163.367
R1767 B.n552 B.n551 163.367
R1768 B.n551 B.n550 163.367
R1769 B.n550 B.n79 163.367
R1770 B.n147 B.n146 74.0854
R1771 B.n155 B.n154 74.0854
R1772 B.n49 B.n48 74.0854
R1773 B.n55 B.n54 74.0854
R1774 B.n148 B.n147 59.5399
R1775 B.n333 B.n155 59.5399
R1776 B.n634 B.n49 59.5399
R1777 B.n620 B.n55 59.5399
R1778 B.n707 B.n706 29.8151
R1779 B.n421 B.n122 29.8151
R1780 B.n261 B.n260 29.8151
R1781 B.n548 B.n547 29.8151
R1782 B B.n771 18.0485
R1783 B.n706 B.n705 10.6151
R1784 B.n705 B.n24 10.6151
R1785 B.n701 B.n24 10.6151
R1786 B.n701 B.n700 10.6151
R1787 B.n700 B.n699 10.6151
R1788 B.n699 B.n26 10.6151
R1789 B.n695 B.n26 10.6151
R1790 B.n695 B.n694 10.6151
R1791 B.n694 B.n693 10.6151
R1792 B.n693 B.n28 10.6151
R1793 B.n689 B.n28 10.6151
R1794 B.n689 B.n688 10.6151
R1795 B.n688 B.n687 10.6151
R1796 B.n687 B.n30 10.6151
R1797 B.n683 B.n30 10.6151
R1798 B.n683 B.n682 10.6151
R1799 B.n682 B.n681 10.6151
R1800 B.n681 B.n32 10.6151
R1801 B.n677 B.n32 10.6151
R1802 B.n677 B.n676 10.6151
R1803 B.n676 B.n675 10.6151
R1804 B.n675 B.n34 10.6151
R1805 B.n671 B.n34 10.6151
R1806 B.n671 B.n670 10.6151
R1807 B.n670 B.n669 10.6151
R1808 B.n669 B.n36 10.6151
R1809 B.n665 B.n36 10.6151
R1810 B.n665 B.n664 10.6151
R1811 B.n664 B.n663 10.6151
R1812 B.n663 B.n38 10.6151
R1813 B.n659 B.n38 10.6151
R1814 B.n659 B.n658 10.6151
R1815 B.n658 B.n657 10.6151
R1816 B.n657 B.n40 10.6151
R1817 B.n653 B.n40 10.6151
R1818 B.n653 B.n652 10.6151
R1819 B.n652 B.n651 10.6151
R1820 B.n651 B.n42 10.6151
R1821 B.n647 B.n42 10.6151
R1822 B.n647 B.n646 10.6151
R1823 B.n646 B.n645 10.6151
R1824 B.n645 B.n44 10.6151
R1825 B.n641 B.n44 10.6151
R1826 B.n641 B.n640 10.6151
R1827 B.n640 B.n639 10.6151
R1828 B.n639 B.n46 10.6151
R1829 B.n635 B.n46 10.6151
R1830 B.n633 B.n632 10.6151
R1831 B.n632 B.n50 10.6151
R1832 B.n628 B.n50 10.6151
R1833 B.n628 B.n627 10.6151
R1834 B.n627 B.n626 10.6151
R1835 B.n626 B.n52 10.6151
R1836 B.n622 B.n52 10.6151
R1837 B.n622 B.n621 10.6151
R1838 B.n619 B.n56 10.6151
R1839 B.n615 B.n56 10.6151
R1840 B.n615 B.n614 10.6151
R1841 B.n614 B.n613 10.6151
R1842 B.n613 B.n58 10.6151
R1843 B.n609 B.n58 10.6151
R1844 B.n609 B.n608 10.6151
R1845 B.n608 B.n607 10.6151
R1846 B.n607 B.n60 10.6151
R1847 B.n603 B.n60 10.6151
R1848 B.n603 B.n602 10.6151
R1849 B.n602 B.n601 10.6151
R1850 B.n601 B.n62 10.6151
R1851 B.n597 B.n62 10.6151
R1852 B.n597 B.n596 10.6151
R1853 B.n596 B.n595 10.6151
R1854 B.n595 B.n64 10.6151
R1855 B.n591 B.n64 10.6151
R1856 B.n591 B.n590 10.6151
R1857 B.n590 B.n589 10.6151
R1858 B.n589 B.n66 10.6151
R1859 B.n585 B.n66 10.6151
R1860 B.n585 B.n584 10.6151
R1861 B.n584 B.n583 10.6151
R1862 B.n583 B.n68 10.6151
R1863 B.n579 B.n68 10.6151
R1864 B.n579 B.n578 10.6151
R1865 B.n578 B.n577 10.6151
R1866 B.n577 B.n70 10.6151
R1867 B.n573 B.n70 10.6151
R1868 B.n573 B.n572 10.6151
R1869 B.n572 B.n571 10.6151
R1870 B.n571 B.n72 10.6151
R1871 B.n567 B.n72 10.6151
R1872 B.n567 B.n566 10.6151
R1873 B.n566 B.n565 10.6151
R1874 B.n565 B.n74 10.6151
R1875 B.n561 B.n74 10.6151
R1876 B.n561 B.n560 10.6151
R1877 B.n560 B.n559 10.6151
R1878 B.n559 B.n76 10.6151
R1879 B.n555 B.n76 10.6151
R1880 B.n555 B.n554 10.6151
R1881 B.n554 B.n553 10.6151
R1882 B.n553 B.n78 10.6151
R1883 B.n549 B.n78 10.6151
R1884 B.n549 B.n548 10.6151
R1885 B.n422 B.n421 10.6151
R1886 B.n423 B.n422 10.6151
R1887 B.n423 B.n120 10.6151
R1888 B.n427 B.n120 10.6151
R1889 B.n428 B.n427 10.6151
R1890 B.n429 B.n428 10.6151
R1891 B.n429 B.n118 10.6151
R1892 B.n433 B.n118 10.6151
R1893 B.n434 B.n433 10.6151
R1894 B.n435 B.n434 10.6151
R1895 B.n435 B.n116 10.6151
R1896 B.n439 B.n116 10.6151
R1897 B.n440 B.n439 10.6151
R1898 B.n441 B.n440 10.6151
R1899 B.n441 B.n114 10.6151
R1900 B.n445 B.n114 10.6151
R1901 B.n446 B.n445 10.6151
R1902 B.n447 B.n446 10.6151
R1903 B.n447 B.n112 10.6151
R1904 B.n451 B.n112 10.6151
R1905 B.n452 B.n451 10.6151
R1906 B.n453 B.n452 10.6151
R1907 B.n453 B.n110 10.6151
R1908 B.n457 B.n110 10.6151
R1909 B.n458 B.n457 10.6151
R1910 B.n459 B.n458 10.6151
R1911 B.n459 B.n108 10.6151
R1912 B.n463 B.n108 10.6151
R1913 B.n464 B.n463 10.6151
R1914 B.n465 B.n464 10.6151
R1915 B.n465 B.n106 10.6151
R1916 B.n469 B.n106 10.6151
R1917 B.n470 B.n469 10.6151
R1918 B.n471 B.n470 10.6151
R1919 B.n471 B.n104 10.6151
R1920 B.n475 B.n104 10.6151
R1921 B.n476 B.n475 10.6151
R1922 B.n477 B.n476 10.6151
R1923 B.n477 B.n102 10.6151
R1924 B.n481 B.n102 10.6151
R1925 B.n482 B.n481 10.6151
R1926 B.n483 B.n482 10.6151
R1927 B.n483 B.n100 10.6151
R1928 B.n487 B.n100 10.6151
R1929 B.n488 B.n487 10.6151
R1930 B.n489 B.n488 10.6151
R1931 B.n489 B.n98 10.6151
R1932 B.n493 B.n98 10.6151
R1933 B.n494 B.n493 10.6151
R1934 B.n495 B.n494 10.6151
R1935 B.n495 B.n96 10.6151
R1936 B.n499 B.n96 10.6151
R1937 B.n500 B.n499 10.6151
R1938 B.n501 B.n500 10.6151
R1939 B.n501 B.n94 10.6151
R1940 B.n505 B.n94 10.6151
R1941 B.n506 B.n505 10.6151
R1942 B.n507 B.n506 10.6151
R1943 B.n507 B.n92 10.6151
R1944 B.n511 B.n92 10.6151
R1945 B.n512 B.n511 10.6151
R1946 B.n513 B.n512 10.6151
R1947 B.n513 B.n90 10.6151
R1948 B.n517 B.n90 10.6151
R1949 B.n518 B.n517 10.6151
R1950 B.n519 B.n518 10.6151
R1951 B.n519 B.n88 10.6151
R1952 B.n523 B.n88 10.6151
R1953 B.n524 B.n523 10.6151
R1954 B.n525 B.n524 10.6151
R1955 B.n525 B.n86 10.6151
R1956 B.n529 B.n86 10.6151
R1957 B.n530 B.n529 10.6151
R1958 B.n531 B.n530 10.6151
R1959 B.n531 B.n84 10.6151
R1960 B.n535 B.n84 10.6151
R1961 B.n536 B.n535 10.6151
R1962 B.n537 B.n536 10.6151
R1963 B.n537 B.n82 10.6151
R1964 B.n541 B.n82 10.6151
R1965 B.n542 B.n541 10.6151
R1966 B.n543 B.n542 10.6151
R1967 B.n543 B.n80 10.6151
R1968 B.n547 B.n80 10.6151
R1969 B.n261 B.n178 10.6151
R1970 B.n265 B.n178 10.6151
R1971 B.n266 B.n265 10.6151
R1972 B.n267 B.n266 10.6151
R1973 B.n267 B.n176 10.6151
R1974 B.n271 B.n176 10.6151
R1975 B.n272 B.n271 10.6151
R1976 B.n273 B.n272 10.6151
R1977 B.n273 B.n174 10.6151
R1978 B.n277 B.n174 10.6151
R1979 B.n278 B.n277 10.6151
R1980 B.n279 B.n278 10.6151
R1981 B.n279 B.n172 10.6151
R1982 B.n283 B.n172 10.6151
R1983 B.n284 B.n283 10.6151
R1984 B.n285 B.n284 10.6151
R1985 B.n285 B.n170 10.6151
R1986 B.n289 B.n170 10.6151
R1987 B.n290 B.n289 10.6151
R1988 B.n291 B.n290 10.6151
R1989 B.n291 B.n168 10.6151
R1990 B.n295 B.n168 10.6151
R1991 B.n296 B.n295 10.6151
R1992 B.n297 B.n296 10.6151
R1993 B.n297 B.n166 10.6151
R1994 B.n301 B.n166 10.6151
R1995 B.n302 B.n301 10.6151
R1996 B.n303 B.n302 10.6151
R1997 B.n303 B.n164 10.6151
R1998 B.n307 B.n164 10.6151
R1999 B.n308 B.n307 10.6151
R2000 B.n309 B.n308 10.6151
R2001 B.n309 B.n162 10.6151
R2002 B.n313 B.n162 10.6151
R2003 B.n314 B.n313 10.6151
R2004 B.n315 B.n314 10.6151
R2005 B.n315 B.n160 10.6151
R2006 B.n319 B.n160 10.6151
R2007 B.n320 B.n319 10.6151
R2008 B.n321 B.n320 10.6151
R2009 B.n321 B.n158 10.6151
R2010 B.n325 B.n158 10.6151
R2011 B.n326 B.n325 10.6151
R2012 B.n327 B.n326 10.6151
R2013 B.n327 B.n156 10.6151
R2014 B.n331 B.n156 10.6151
R2015 B.n332 B.n331 10.6151
R2016 B.n334 B.n152 10.6151
R2017 B.n338 B.n152 10.6151
R2018 B.n339 B.n338 10.6151
R2019 B.n340 B.n339 10.6151
R2020 B.n340 B.n150 10.6151
R2021 B.n344 B.n150 10.6151
R2022 B.n345 B.n344 10.6151
R2023 B.n346 B.n345 10.6151
R2024 B.n350 B.n349 10.6151
R2025 B.n351 B.n350 10.6151
R2026 B.n351 B.n144 10.6151
R2027 B.n355 B.n144 10.6151
R2028 B.n356 B.n355 10.6151
R2029 B.n357 B.n356 10.6151
R2030 B.n357 B.n142 10.6151
R2031 B.n361 B.n142 10.6151
R2032 B.n362 B.n361 10.6151
R2033 B.n363 B.n362 10.6151
R2034 B.n363 B.n140 10.6151
R2035 B.n367 B.n140 10.6151
R2036 B.n368 B.n367 10.6151
R2037 B.n369 B.n368 10.6151
R2038 B.n369 B.n138 10.6151
R2039 B.n373 B.n138 10.6151
R2040 B.n374 B.n373 10.6151
R2041 B.n375 B.n374 10.6151
R2042 B.n375 B.n136 10.6151
R2043 B.n379 B.n136 10.6151
R2044 B.n380 B.n379 10.6151
R2045 B.n381 B.n380 10.6151
R2046 B.n381 B.n134 10.6151
R2047 B.n385 B.n134 10.6151
R2048 B.n386 B.n385 10.6151
R2049 B.n387 B.n386 10.6151
R2050 B.n387 B.n132 10.6151
R2051 B.n391 B.n132 10.6151
R2052 B.n392 B.n391 10.6151
R2053 B.n393 B.n392 10.6151
R2054 B.n393 B.n130 10.6151
R2055 B.n397 B.n130 10.6151
R2056 B.n398 B.n397 10.6151
R2057 B.n399 B.n398 10.6151
R2058 B.n399 B.n128 10.6151
R2059 B.n403 B.n128 10.6151
R2060 B.n404 B.n403 10.6151
R2061 B.n405 B.n404 10.6151
R2062 B.n405 B.n126 10.6151
R2063 B.n409 B.n126 10.6151
R2064 B.n410 B.n409 10.6151
R2065 B.n411 B.n410 10.6151
R2066 B.n411 B.n124 10.6151
R2067 B.n415 B.n124 10.6151
R2068 B.n416 B.n415 10.6151
R2069 B.n417 B.n416 10.6151
R2070 B.n417 B.n122 10.6151
R2071 B.n260 B.n259 10.6151
R2072 B.n259 B.n180 10.6151
R2073 B.n255 B.n180 10.6151
R2074 B.n255 B.n254 10.6151
R2075 B.n254 B.n253 10.6151
R2076 B.n253 B.n182 10.6151
R2077 B.n249 B.n182 10.6151
R2078 B.n249 B.n248 10.6151
R2079 B.n248 B.n247 10.6151
R2080 B.n247 B.n184 10.6151
R2081 B.n243 B.n184 10.6151
R2082 B.n243 B.n242 10.6151
R2083 B.n242 B.n241 10.6151
R2084 B.n241 B.n186 10.6151
R2085 B.n237 B.n186 10.6151
R2086 B.n237 B.n236 10.6151
R2087 B.n236 B.n235 10.6151
R2088 B.n235 B.n188 10.6151
R2089 B.n231 B.n188 10.6151
R2090 B.n231 B.n230 10.6151
R2091 B.n230 B.n229 10.6151
R2092 B.n229 B.n190 10.6151
R2093 B.n225 B.n190 10.6151
R2094 B.n225 B.n224 10.6151
R2095 B.n224 B.n223 10.6151
R2096 B.n223 B.n192 10.6151
R2097 B.n219 B.n192 10.6151
R2098 B.n219 B.n218 10.6151
R2099 B.n218 B.n217 10.6151
R2100 B.n217 B.n194 10.6151
R2101 B.n213 B.n194 10.6151
R2102 B.n213 B.n212 10.6151
R2103 B.n212 B.n211 10.6151
R2104 B.n211 B.n196 10.6151
R2105 B.n207 B.n196 10.6151
R2106 B.n207 B.n206 10.6151
R2107 B.n206 B.n205 10.6151
R2108 B.n205 B.n198 10.6151
R2109 B.n201 B.n198 10.6151
R2110 B.n201 B.n200 10.6151
R2111 B.n200 B.n0 10.6151
R2112 B.n767 B.n1 10.6151
R2113 B.n767 B.n766 10.6151
R2114 B.n766 B.n765 10.6151
R2115 B.n765 B.n4 10.6151
R2116 B.n761 B.n4 10.6151
R2117 B.n761 B.n760 10.6151
R2118 B.n760 B.n759 10.6151
R2119 B.n759 B.n6 10.6151
R2120 B.n755 B.n6 10.6151
R2121 B.n755 B.n754 10.6151
R2122 B.n754 B.n753 10.6151
R2123 B.n753 B.n8 10.6151
R2124 B.n749 B.n8 10.6151
R2125 B.n749 B.n748 10.6151
R2126 B.n748 B.n747 10.6151
R2127 B.n747 B.n10 10.6151
R2128 B.n743 B.n10 10.6151
R2129 B.n743 B.n742 10.6151
R2130 B.n742 B.n741 10.6151
R2131 B.n741 B.n12 10.6151
R2132 B.n737 B.n12 10.6151
R2133 B.n737 B.n736 10.6151
R2134 B.n736 B.n735 10.6151
R2135 B.n735 B.n14 10.6151
R2136 B.n731 B.n14 10.6151
R2137 B.n731 B.n730 10.6151
R2138 B.n730 B.n729 10.6151
R2139 B.n729 B.n16 10.6151
R2140 B.n725 B.n16 10.6151
R2141 B.n725 B.n724 10.6151
R2142 B.n724 B.n723 10.6151
R2143 B.n723 B.n18 10.6151
R2144 B.n719 B.n18 10.6151
R2145 B.n719 B.n718 10.6151
R2146 B.n718 B.n717 10.6151
R2147 B.n717 B.n20 10.6151
R2148 B.n713 B.n20 10.6151
R2149 B.n713 B.n712 10.6151
R2150 B.n712 B.n711 10.6151
R2151 B.n711 B.n22 10.6151
R2152 B.n707 B.n22 10.6151
R2153 B.n634 B.n633 6.5566
R2154 B.n621 B.n620 6.5566
R2155 B.n334 B.n333 6.5566
R2156 B.n346 B.n148 6.5566
R2157 B.n635 B.n634 4.05904
R2158 B.n620 B.n619 4.05904
R2159 B.n333 B.n332 4.05904
R2160 B.n349 B.n148 4.05904
R2161 B.n771 B.n0 2.81026
R2162 B.n771 B.n1 2.81026
C0 VDD1 VTAIL 6.07591f
C1 VN w_n3262_n3778# 5.73061f
C2 VDD2 VDD1 1.23897f
C3 VDD2 VTAIL 6.13609f
C4 B w_n3262_n3778# 10.914701f
C5 VP w_n3262_n3778# 6.1522f
C6 B VN 1.30169f
C7 VN VP 7.21436f
C8 B VP 2.00545f
C9 VDD1 w_n3262_n3778# 1.67768f
C10 VN VDD1 0.149954f
C11 w_n3262_n3778# VTAIL 4.45491f
C12 VN VTAIL 5.71686f
C13 VDD2 w_n3262_n3778# 1.75343f
C14 VDD2 VN 5.76742f
C15 B VDD1 1.47448f
C16 VDD1 VP 6.06759f
C17 B VTAIL 6.01531f
C18 VP VTAIL 5.73097f
C19 B VDD2 1.54137f
C20 VDD2 VP 0.451088f
C21 VDD2 VSUBS 1.1431f
C22 VDD1 VSUBS 6.522f
C23 VTAIL VSUBS 1.416573f
C24 VN VSUBS 5.99847f
C25 VP VSUBS 2.832158f
C26 B VSUBS 5.215698f
C27 w_n3262_n3778# VSUBS 0.151292p
C28 B.n0 VSUBS 0.004225f
C29 B.n1 VSUBS 0.004225f
C30 B.n2 VSUBS 0.006681f
C31 B.n3 VSUBS 0.006681f
C32 B.n4 VSUBS 0.006681f
C33 B.n5 VSUBS 0.006681f
C34 B.n6 VSUBS 0.006681f
C35 B.n7 VSUBS 0.006681f
C36 B.n8 VSUBS 0.006681f
C37 B.n9 VSUBS 0.006681f
C38 B.n10 VSUBS 0.006681f
C39 B.n11 VSUBS 0.006681f
C40 B.n12 VSUBS 0.006681f
C41 B.n13 VSUBS 0.006681f
C42 B.n14 VSUBS 0.006681f
C43 B.n15 VSUBS 0.006681f
C44 B.n16 VSUBS 0.006681f
C45 B.n17 VSUBS 0.006681f
C46 B.n18 VSUBS 0.006681f
C47 B.n19 VSUBS 0.006681f
C48 B.n20 VSUBS 0.006681f
C49 B.n21 VSUBS 0.006681f
C50 B.n22 VSUBS 0.006681f
C51 B.n23 VSUBS 0.015065f
C52 B.n24 VSUBS 0.006681f
C53 B.n25 VSUBS 0.006681f
C54 B.n26 VSUBS 0.006681f
C55 B.n27 VSUBS 0.006681f
C56 B.n28 VSUBS 0.006681f
C57 B.n29 VSUBS 0.006681f
C58 B.n30 VSUBS 0.006681f
C59 B.n31 VSUBS 0.006681f
C60 B.n32 VSUBS 0.006681f
C61 B.n33 VSUBS 0.006681f
C62 B.n34 VSUBS 0.006681f
C63 B.n35 VSUBS 0.006681f
C64 B.n36 VSUBS 0.006681f
C65 B.n37 VSUBS 0.006681f
C66 B.n38 VSUBS 0.006681f
C67 B.n39 VSUBS 0.006681f
C68 B.n40 VSUBS 0.006681f
C69 B.n41 VSUBS 0.006681f
C70 B.n42 VSUBS 0.006681f
C71 B.n43 VSUBS 0.006681f
C72 B.n44 VSUBS 0.006681f
C73 B.n45 VSUBS 0.006681f
C74 B.n46 VSUBS 0.006681f
C75 B.n47 VSUBS 0.006681f
C76 B.t5 VSUBS 0.245721f
C77 B.t4 VSUBS 0.285432f
C78 B.t3 VSUBS 2.15274f
C79 B.n48 VSUBS 0.45396f
C80 B.n49 VSUBS 0.270329f
C81 B.n50 VSUBS 0.006681f
C82 B.n51 VSUBS 0.006681f
C83 B.n52 VSUBS 0.006681f
C84 B.n53 VSUBS 0.006681f
C85 B.t2 VSUBS 0.245724f
C86 B.t1 VSUBS 0.285435f
C87 B.t0 VSUBS 2.15274f
C88 B.n54 VSUBS 0.453957f
C89 B.n55 VSUBS 0.270326f
C90 B.n56 VSUBS 0.006681f
C91 B.n57 VSUBS 0.006681f
C92 B.n58 VSUBS 0.006681f
C93 B.n59 VSUBS 0.006681f
C94 B.n60 VSUBS 0.006681f
C95 B.n61 VSUBS 0.006681f
C96 B.n62 VSUBS 0.006681f
C97 B.n63 VSUBS 0.006681f
C98 B.n64 VSUBS 0.006681f
C99 B.n65 VSUBS 0.006681f
C100 B.n66 VSUBS 0.006681f
C101 B.n67 VSUBS 0.006681f
C102 B.n68 VSUBS 0.006681f
C103 B.n69 VSUBS 0.006681f
C104 B.n70 VSUBS 0.006681f
C105 B.n71 VSUBS 0.006681f
C106 B.n72 VSUBS 0.006681f
C107 B.n73 VSUBS 0.006681f
C108 B.n74 VSUBS 0.006681f
C109 B.n75 VSUBS 0.006681f
C110 B.n76 VSUBS 0.006681f
C111 B.n77 VSUBS 0.006681f
C112 B.n78 VSUBS 0.006681f
C113 B.n79 VSUBS 0.015065f
C114 B.n80 VSUBS 0.006681f
C115 B.n81 VSUBS 0.006681f
C116 B.n82 VSUBS 0.006681f
C117 B.n83 VSUBS 0.006681f
C118 B.n84 VSUBS 0.006681f
C119 B.n85 VSUBS 0.006681f
C120 B.n86 VSUBS 0.006681f
C121 B.n87 VSUBS 0.006681f
C122 B.n88 VSUBS 0.006681f
C123 B.n89 VSUBS 0.006681f
C124 B.n90 VSUBS 0.006681f
C125 B.n91 VSUBS 0.006681f
C126 B.n92 VSUBS 0.006681f
C127 B.n93 VSUBS 0.006681f
C128 B.n94 VSUBS 0.006681f
C129 B.n95 VSUBS 0.006681f
C130 B.n96 VSUBS 0.006681f
C131 B.n97 VSUBS 0.006681f
C132 B.n98 VSUBS 0.006681f
C133 B.n99 VSUBS 0.006681f
C134 B.n100 VSUBS 0.006681f
C135 B.n101 VSUBS 0.006681f
C136 B.n102 VSUBS 0.006681f
C137 B.n103 VSUBS 0.006681f
C138 B.n104 VSUBS 0.006681f
C139 B.n105 VSUBS 0.006681f
C140 B.n106 VSUBS 0.006681f
C141 B.n107 VSUBS 0.006681f
C142 B.n108 VSUBS 0.006681f
C143 B.n109 VSUBS 0.006681f
C144 B.n110 VSUBS 0.006681f
C145 B.n111 VSUBS 0.006681f
C146 B.n112 VSUBS 0.006681f
C147 B.n113 VSUBS 0.006681f
C148 B.n114 VSUBS 0.006681f
C149 B.n115 VSUBS 0.006681f
C150 B.n116 VSUBS 0.006681f
C151 B.n117 VSUBS 0.006681f
C152 B.n118 VSUBS 0.006681f
C153 B.n119 VSUBS 0.006681f
C154 B.n120 VSUBS 0.006681f
C155 B.n121 VSUBS 0.006681f
C156 B.n122 VSUBS 0.015065f
C157 B.n123 VSUBS 0.006681f
C158 B.n124 VSUBS 0.006681f
C159 B.n125 VSUBS 0.006681f
C160 B.n126 VSUBS 0.006681f
C161 B.n127 VSUBS 0.006681f
C162 B.n128 VSUBS 0.006681f
C163 B.n129 VSUBS 0.006681f
C164 B.n130 VSUBS 0.006681f
C165 B.n131 VSUBS 0.006681f
C166 B.n132 VSUBS 0.006681f
C167 B.n133 VSUBS 0.006681f
C168 B.n134 VSUBS 0.006681f
C169 B.n135 VSUBS 0.006681f
C170 B.n136 VSUBS 0.006681f
C171 B.n137 VSUBS 0.006681f
C172 B.n138 VSUBS 0.006681f
C173 B.n139 VSUBS 0.006681f
C174 B.n140 VSUBS 0.006681f
C175 B.n141 VSUBS 0.006681f
C176 B.n142 VSUBS 0.006681f
C177 B.n143 VSUBS 0.006681f
C178 B.n144 VSUBS 0.006681f
C179 B.n145 VSUBS 0.006681f
C180 B.t10 VSUBS 0.245724f
C181 B.t11 VSUBS 0.285435f
C182 B.t9 VSUBS 2.15274f
C183 B.n146 VSUBS 0.453957f
C184 B.n147 VSUBS 0.270326f
C185 B.n148 VSUBS 0.01548f
C186 B.n149 VSUBS 0.006681f
C187 B.n150 VSUBS 0.006681f
C188 B.n151 VSUBS 0.006681f
C189 B.n152 VSUBS 0.006681f
C190 B.n153 VSUBS 0.006681f
C191 B.t7 VSUBS 0.245721f
C192 B.t8 VSUBS 0.285432f
C193 B.t6 VSUBS 2.15274f
C194 B.n154 VSUBS 0.45396f
C195 B.n155 VSUBS 0.270329f
C196 B.n156 VSUBS 0.006681f
C197 B.n157 VSUBS 0.006681f
C198 B.n158 VSUBS 0.006681f
C199 B.n159 VSUBS 0.006681f
C200 B.n160 VSUBS 0.006681f
C201 B.n161 VSUBS 0.006681f
C202 B.n162 VSUBS 0.006681f
C203 B.n163 VSUBS 0.006681f
C204 B.n164 VSUBS 0.006681f
C205 B.n165 VSUBS 0.006681f
C206 B.n166 VSUBS 0.006681f
C207 B.n167 VSUBS 0.006681f
C208 B.n168 VSUBS 0.006681f
C209 B.n169 VSUBS 0.006681f
C210 B.n170 VSUBS 0.006681f
C211 B.n171 VSUBS 0.006681f
C212 B.n172 VSUBS 0.006681f
C213 B.n173 VSUBS 0.006681f
C214 B.n174 VSUBS 0.006681f
C215 B.n175 VSUBS 0.006681f
C216 B.n176 VSUBS 0.006681f
C217 B.n177 VSUBS 0.006681f
C218 B.n178 VSUBS 0.006681f
C219 B.n179 VSUBS 0.014411f
C220 B.n180 VSUBS 0.006681f
C221 B.n181 VSUBS 0.006681f
C222 B.n182 VSUBS 0.006681f
C223 B.n183 VSUBS 0.006681f
C224 B.n184 VSUBS 0.006681f
C225 B.n185 VSUBS 0.006681f
C226 B.n186 VSUBS 0.006681f
C227 B.n187 VSUBS 0.006681f
C228 B.n188 VSUBS 0.006681f
C229 B.n189 VSUBS 0.006681f
C230 B.n190 VSUBS 0.006681f
C231 B.n191 VSUBS 0.006681f
C232 B.n192 VSUBS 0.006681f
C233 B.n193 VSUBS 0.006681f
C234 B.n194 VSUBS 0.006681f
C235 B.n195 VSUBS 0.006681f
C236 B.n196 VSUBS 0.006681f
C237 B.n197 VSUBS 0.006681f
C238 B.n198 VSUBS 0.006681f
C239 B.n199 VSUBS 0.006681f
C240 B.n200 VSUBS 0.006681f
C241 B.n201 VSUBS 0.006681f
C242 B.n202 VSUBS 0.006681f
C243 B.n203 VSUBS 0.006681f
C244 B.n204 VSUBS 0.006681f
C245 B.n205 VSUBS 0.006681f
C246 B.n206 VSUBS 0.006681f
C247 B.n207 VSUBS 0.006681f
C248 B.n208 VSUBS 0.006681f
C249 B.n209 VSUBS 0.006681f
C250 B.n210 VSUBS 0.006681f
C251 B.n211 VSUBS 0.006681f
C252 B.n212 VSUBS 0.006681f
C253 B.n213 VSUBS 0.006681f
C254 B.n214 VSUBS 0.006681f
C255 B.n215 VSUBS 0.006681f
C256 B.n216 VSUBS 0.006681f
C257 B.n217 VSUBS 0.006681f
C258 B.n218 VSUBS 0.006681f
C259 B.n219 VSUBS 0.006681f
C260 B.n220 VSUBS 0.006681f
C261 B.n221 VSUBS 0.006681f
C262 B.n222 VSUBS 0.006681f
C263 B.n223 VSUBS 0.006681f
C264 B.n224 VSUBS 0.006681f
C265 B.n225 VSUBS 0.006681f
C266 B.n226 VSUBS 0.006681f
C267 B.n227 VSUBS 0.006681f
C268 B.n228 VSUBS 0.006681f
C269 B.n229 VSUBS 0.006681f
C270 B.n230 VSUBS 0.006681f
C271 B.n231 VSUBS 0.006681f
C272 B.n232 VSUBS 0.006681f
C273 B.n233 VSUBS 0.006681f
C274 B.n234 VSUBS 0.006681f
C275 B.n235 VSUBS 0.006681f
C276 B.n236 VSUBS 0.006681f
C277 B.n237 VSUBS 0.006681f
C278 B.n238 VSUBS 0.006681f
C279 B.n239 VSUBS 0.006681f
C280 B.n240 VSUBS 0.006681f
C281 B.n241 VSUBS 0.006681f
C282 B.n242 VSUBS 0.006681f
C283 B.n243 VSUBS 0.006681f
C284 B.n244 VSUBS 0.006681f
C285 B.n245 VSUBS 0.006681f
C286 B.n246 VSUBS 0.006681f
C287 B.n247 VSUBS 0.006681f
C288 B.n248 VSUBS 0.006681f
C289 B.n249 VSUBS 0.006681f
C290 B.n250 VSUBS 0.006681f
C291 B.n251 VSUBS 0.006681f
C292 B.n252 VSUBS 0.006681f
C293 B.n253 VSUBS 0.006681f
C294 B.n254 VSUBS 0.006681f
C295 B.n255 VSUBS 0.006681f
C296 B.n256 VSUBS 0.006681f
C297 B.n257 VSUBS 0.006681f
C298 B.n258 VSUBS 0.006681f
C299 B.n259 VSUBS 0.006681f
C300 B.n260 VSUBS 0.014411f
C301 B.n261 VSUBS 0.015065f
C302 B.n262 VSUBS 0.015065f
C303 B.n263 VSUBS 0.006681f
C304 B.n264 VSUBS 0.006681f
C305 B.n265 VSUBS 0.006681f
C306 B.n266 VSUBS 0.006681f
C307 B.n267 VSUBS 0.006681f
C308 B.n268 VSUBS 0.006681f
C309 B.n269 VSUBS 0.006681f
C310 B.n270 VSUBS 0.006681f
C311 B.n271 VSUBS 0.006681f
C312 B.n272 VSUBS 0.006681f
C313 B.n273 VSUBS 0.006681f
C314 B.n274 VSUBS 0.006681f
C315 B.n275 VSUBS 0.006681f
C316 B.n276 VSUBS 0.006681f
C317 B.n277 VSUBS 0.006681f
C318 B.n278 VSUBS 0.006681f
C319 B.n279 VSUBS 0.006681f
C320 B.n280 VSUBS 0.006681f
C321 B.n281 VSUBS 0.006681f
C322 B.n282 VSUBS 0.006681f
C323 B.n283 VSUBS 0.006681f
C324 B.n284 VSUBS 0.006681f
C325 B.n285 VSUBS 0.006681f
C326 B.n286 VSUBS 0.006681f
C327 B.n287 VSUBS 0.006681f
C328 B.n288 VSUBS 0.006681f
C329 B.n289 VSUBS 0.006681f
C330 B.n290 VSUBS 0.006681f
C331 B.n291 VSUBS 0.006681f
C332 B.n292 VSUBS 0.006681f
C333 B.n293 VSUBS 0.006681f
C334 B.n294 VSUBS 0.006681f
C335 B.n295 VSUBS 0.006681f
C336 B.n296 VSUBS 0.006681f
C337 B.n297 VSUBS 0.006681f
C338 B.n298 VSUBS 0.006681f
C339 B.n299 VSUBS 0.006681f
C340 B.n300 VSUBS 0.006681f
C341 B.n301 VSUBS 0.006681f
C342 B.n302 VSUBS 0.006681f
C343 B.n303 VSUBS 0.006681f
C344 B.n304 VSUBS 0.006681f
C345 B.n305 VSUBS 0.006681f
C346 B.n306 VSUBS 0.006681f
C347 B.n307 VSUBS 0.006681f
C348 B.n308 VSUBS 0.006681f
C349 B.n309 VSUBS 0.006681f
C350 B.n310 VSUBS 0.006681f
C351 B.n311 VSUBS 0.006681f
C352 B.n312 VSUBS 0.006681f
C353 B.n313 VSUBS 0.006681f
C354 B.n314 VSUBS 0.006681f
C355 B.n315 VSUBS 0.006681f
C356 B.n316 VSUBS 0.006681f
C357 B.n317 VSUBS 0.006681f
C358 B.n318 VSUBS 0.006681f
C359 B.n319 VSUBS 0.006681f
C360 B.n320 VSUBS 0.006681f
C361 B.n321 VSUBS 0.006681f
C362 B.n322 VSUBS 0.006681f
C363 B.n323 VSUBS 0.006681f
C364 B.n324 VSUBS 0.006681f
C365 B.n325 VSUBS 0.006681f
C366 B.n326 VSUBS 0.006681f
C367 B.n327 VSUBS 0.006681f
C368 B.n328 VSUBS 0.006681f
C369 B.n329 VSUBS 0.006681f
C370 B.n330 VSUBS 0.006681f
C371 B.n331 VSUBS 0.006681f
C372 B.n332 VSUBS 0.004618f
C373 B.n333 VSUBS 0.01548f
C374 B.n334 VSUBS 0.005404f
C375 B.n335 VSUBS 0.006681f
C376 B.n336 VSUBS 0.006681f
C377 B.n337 VSUBS 0.006681f
C378 B.n338 VSUBS 0.006681f
C379 B.n339 VSUBS 0.006681f
C380 B.n340 VSUBS 0.006681f
C381 B.n341 VSUBS 0.006681f
C382 B.n342 VSUBS 0.006681f
C383 B.n343 VSUBS 0.006681f
C384 B.n344 VSUBS 0.006681f
C385 B.n345 VSUBS 0.006681f
C386 B.n346 VSUBS 0.005404f
C387 B.n347 VSUBS 0.006681f
C388 B.n348 VSUBS 0.006681f
C389 B.n349 VSUBS 0.004618f
C390 B.n350 VSUBS 0.006681f
C391 B.n351 VSUBS 0.006681f
C392 B.n352 VSUBS 0.006681f
C393 B.n353 VSUBS 0.006681f
C394 B.n354 VSUBS 0.006681f
C395 B.n355 VSUBS 0.006681f
C396 B.n356 VSUBS 0.006681f
C397 B.n357 VSUBS 0.006681f
C398 B.n358 VSUBS 0.006681f
C399 B.n359 VSUBS 0.006681f
C400 B.n360 VSUBS 0.006681f
C401 B.n361 VSUBS 0.006681f
C402 B.n362 VSUBS 0.006681f
C403 B.n363 VSUBS 0.006681f
C404 B.n364 VSUBS 0.006681f
C405 B.n365 VSUBS 0.006681f
C406 B.n366 VSUBS 0.006681f
C407 B.n367 VSUBS 0.006681f
C408 B.n368 VSUBS 0.006681f
C409 B.n369 VSUBS 0.006681f
C410 B.n370 VSUBS 0.006681f
C411 B.n371 VSUBS 0.006681f
C412 B.n372 VSUBS 0.006681f
C413 B.n373 VSUBS 0.006681f
C414 B.n374 VSUBS 0.006681f
C415 B.n375 VSUBS 0.006681f
C416 B.n376 VSUBS 0.006681f
C417 B.n377 VSUBS 0.006681f
C418 B.n378 VSUBS 0.006681f
C419 B.n379 VSUBS 0.006681f
C420 B.n380 VSUBS 0.006681f
C421 B.n381 VSUBS 0.006681f
C422 B.n382 VSUBS 0.006681f
C423 B.n383 VSUBS 0.006681f
C424 B.n384 VSUBS 0.006681f
C425 B.n385 VSUBS 0.006681f
C426 B.n386 VSUBS 0.006681f
C427 B.n387 VSUBS 0.006681f
C428 B.n388 VSUBS 0.006681f
C429 B.n389 VSUBS 0.006681f
C430 B.n390 VSUBS 0.006681f
C431 B.n391 VSUBS 0.006681f
C432 B.n392 VSUBS 0.006681f
C433 B.n393 VSUBS 0.006681f
C434 B.n394 VSUBS 0.006681f
C435 B.n395 VSUBS 0.006681f
C436 B.n396 VSUBS 0.006681f
C437 B.n397 VSUBS 0.006681f
C438 B.n398 VSUBS 0.006681f
C439 B.n399 VSUBS 0.006681f
C440 B.n400 VSUBS 0.006681f
C441 B.n401 VSUBS 0.006681f
C442 B.n402 VSUBS 0.006681f
C443 B.n403 VSUBS 0.006681f
C444 B.n404 VSUBS 0.006681f
C445 B.n405 VSUBS 0.006681f
C446 B.n406 VSUBS 0.006681f
C447 B.n407 VSUBS 0.006681f
C448 B.n408 VSUBS 0.006681f
C449 B.n409 VSUBS 0.006681f
C450 B.n410 VSUBS 0.006681f
C451 B.n411 VSUBS 0.006681f
C452 B.n412 VSUBS 0.006681f
C453 B.n413 VSUBS 0.006681f
C454 B.n414 VSUBS 0.006681f
C455 B.n415 VSUBS 0.006681f
C456 B.n416 VSUBS 0.006681f
C457 B.n417 VSUBS 0.006681f
C458 B.n418 VSUBS 0.006681f
C459 B.n419 VSUBS 0.015065f
C460 B.n420 VSUBS 0.014411f
C461 B.n421 VSUBS 0.014411f
C462 B.n422 VSUBS 0.006681f
C463 B.n423 VSUBS 0.006681f
C464 B.n424 VSUBS 0.006681f
C465 B.n425 VSUBS 0.006681f
C466 B.n426 VSUBS 0.006681f
C467 B.n427 VSUBS 0.006681f
C468 B.n428 VSUBS 0.006681f
C469 B.n429 VSUBS 0.006681f
C470 B.n430 VSUBS 0.006681f
C471 B.n431 VSUBS 0.006681f
C472 B.n432 VSUBS 0.006681f
C473 B.n433 VSUBS 0.006681f
C474 B.n434 VSUBS 0.006681f
C475 B.n435 VSUBS 0.006681f
C476 B.n436 VSUBS 0.006681f
C477 B.n437 VSUBS 0.006681f
C478 B.n438 VSUBS 0.006681f
C479 B.n439 VSUBS 0.006681f
C480 B.n440 VSUBS 0.006681f
C481 B.n441 VSUBS 0.006681f
C482 B.n442 VSUBS 0.006681f
C483 B.n443 VSUBS 0.006681f
C484 B.n444 VSUBS 0.006681f
C485 B.n445 VSUBS 0.006681f
C486 B.n446 VSUBS 0.006681f
C487 B.n447 VSUBS 0.006681f
C488 B.n448 VSUBS 0.006681f
C489 B.n449 VSUBS 0.006681f
C490 B.n450 VSUBS 0.006681f
C491 B.n451 VSUBS 0.006681f
C492 B.n452 VSUBS 0.006681f
C493 B.n453 VSUBS 0.006681f
C494 B.n454 VSUBS 0.006681f
C495 B.n455 VSUBS 0.006681f
C496 B.n456 VSUBS 0.006681f
C497 B.n457 VSUBS 0.006681f
C498 B.n458 VSUBS 0.006681f
C499 B.n459 VSUBS 0.006681f
C500 B.n460 VSUBS 0.006681f
C501 B.n461 VSUBS 0.006681f
C502 B.n462 VSUBS 0.006681f
C503 B.n463 VSUBS 0.006681f
C504 B.n464 VSUBS 0.006681f
C505 B.n465 VSUBS 0.006681f
C506 B.n466 VSUBS 0.006681f
C507 B.n467 VSUBS 0.006681f
C508 B.n468 VSUBS 0.006681f
C509 B.n469 VSUBS 0.006681f
C510 B.n470 VSUBS 0.006681f
C511 B.n471 VSUBS 0.006681f
C512 B.n472 VSUBS 0.006681f
C513 B.n473 VSUBS 0.006681f
C514 B.n474 VSUBS 0.006681f
C515 B.n475 VSUBS 0.006681f
C516 B.n476 VSUBS 0.006681f
C517 B.n477 VSUBS 0.006681f
C518 B.n478 VSUBS 0.006681f
C519 B.n479 VSUBS 0.006681f
C520 B.n480 VSUBS 0.006681f
C521 B.n481 VSUBS 0.006681f
C522 B.n482 VSUBS 0.006681f
C523 B.n483 VSUBS 0.006681f
C524 B.n484 VSUBS 0.006681f
C525 B.n485 VSUBS 0.006681f
C526 B.n486 VSUBS 0.006681f
C527 B.n487 VSUBS 0.006681f
C528 B.n488 VSUBS 0.006681f
C529 B.n489 VSUBS 0.006681f
C530 B.n490 VSUBS 0.006681f
C531 B.n491 VSUBS 0.006681f
C532 B.n492 VSUBS 0.006681f
C533 B.n493 VSUBS 0.006681f
C534 B.n494 VSUBS 0.006681f
C535 B.n495 VSUBS 0.006681f
C536 B.n496 VSUBS 0.006681f
C537 B.n497 VSUBS 0.006681f
C538 B.n498 VSUBS 0.006681f
C539 B.n499 VSUBS 0.006681f
C540 B.n500 VSUBS 0.006681f
C541 B.n501 VSUBS 0.006681f
C542 B.n502 VSUBS 0.006681f
C543 B.n503 VSUBS 0.006681f
C544 B.n504 VSUBS 0.006681f
C545 B.n505 VSUBS 0.006681f
C546 B.n506 VSUBS 0.006681f
C547 B.n507 VSUBS 0.006681f
C548 B.n508 VSUBS 0.006681f
C549 B.n509 VSUBS 0.006681f
C550 B.n510 VSUBS 0.006681f
C551 B.n511 VSUBS 0.006681f
C552 B.n512 VSUBS 0.006681f
C553 B.n513 VSUBS 0.006681f
C554 B.n514 VSUBS 0.006681f
C555 B.n515 VSUBS 0.006681f
C556 B.n516 VSUBS 0.006681f
C557 B.n517 VSUBS 0.006681f
C558 B.n518 VSUBS 0.006681f
C559 B.n519 VSUBS 0.006681f
C560 B.n520 VSUBS 0.006681f
C561 B.n521 VSUBS 0.006681f
C562 B.n522 VSUBS 0.006681f
C563 B.n523 VSUBS 0.006681f
C564 B.n524 VSUBS 0.006681f
C565 B.n525 VSUBS 0.006681f
C566 B.n526 VSUBS 0.006681f
C567 B.n527 VSUBS 0.006681f
C568 B.n528 VSUBS 0.006681f
C569 B.n529 VSUBS 0.006681f
C570 B.n530 VSUBS 0.006681f
C571 B.n531 VSUBS 0.006681f
C572 B.n532 VSUBS 0.006681f
C573 B.n533 VSUBS 0.006681f
C574 B.n534 VSUBS 0.006681f
C575 B.n535 VSUBS 0.006681f
C576 B.n536 VSUBS 0.006681f
C577 B.n537 VSUBS 0.006681f
C578 B.n538 VSUBS 0.006681f
C579 B.n539 VSUBS 0.006681f
C580 B.n540 VSUBS 0.006681f
C581 B.n541 VSUBS 0.006681f
C582 B.n542 VSUBS 0.006681f
C583 B.n543 VSUBS 0.006681f
C584 B.n544 VSUBS 0.006681f
C585 B.n545 VSUBS 0.006681f
C586 B.n546 VSUBS 0.014411f
C587 B.n547 VSUBS 0.015276f
C588 B.n548 VSUBS 0.0142f
C589 B.n549 VSUBS 0.006681f
C590 B.n550 VSUBS 0.006681f
C591 B.n551 VSUBS 0.006681f
C592 B.n552 VSUBS 0.006681f
C593 B.n553 VSUBS 0.006681f
C594 B.n554 VSUBS 0.006681f
C595 B.n555 VSUBS 0.006681f
C596 B.n556 VSUBS 0.006681f
C597 B.n557 VSUBS 0.006681f
C598 B.n558 VSUBS 0.006681f
C599 B.n559 VSUBS 0.006681f
C600 B.n560 VSUBS 0.006681f
C601 B.n561 VSUBS 0.006681f
C602 B.n562 VSUBS 0.006681f
C603 B.n563 VSUBS 0.006681f
C604 B.n564 VSUBS 0.006681f
C605 B.n565 VSUBS 0.006681f
C606 B.n566 VSUBS 0.006681f
C607 B.n567 VSUBS 0.006681f
C608 B.n568 VSUBS 0.006681f
C609 B.n569 VSUBS 0.006681f
C610 B.n570 VSUBS 0.006681f
C611 B.n571 VSUBS 0.006681f
C612 B.n572 VSUBS 0.006681f
C613 B.n573 VSUBS 0.006681f
C614 B.n574 VSUBS 0.006681f
C615 B.n575 VSUBS 0.006681f
C616 B.n576 VSUBS 0.006681f
C617 B.n577 VSUBS 0.006681f
C618 B.n578 VSUBS 0.006681f
C619 B.n579 VSUBS 0.006681f
C620 B.n580 VSUBS 0.006681f
C621 B.n581 VSUBS 0.006681f
C622 B.n582 VSUBS 0.006681f
C623 B.n583 VSUBS 0.006681f
C624 B.n584 VSUBS 0.006681f
C625 B.n585 VSUBS 0.006681f
C626 B.n586 VSUBS 0.006681f
C627 B.n587 VSUBS 0.006681f
C628 B.n588 VSUBS 0.006681f
C629 B.n589 VSUBS 0.006681f
C630 B.n590 VSUBS 0.006681f
C631 B.n591 VSUBS 0.006681f
C632 B.n592 VSUBS 0.006681f
C633 B.n593 VSUBS 0.006681f
C634 B.n594 VSUBS 0.006681f
C635 B.n595 VSUBS 0.006681f
C636 B.n596 VSUBS 0.006681f
C637 B.n597 VSUBS 0.006681f
C638 B.n598 VSUBS 0.006681f
C639 B.n599 VSUBS 0.006681f
C640 B.n600 VSUBS 0.006681f
C641 B.n601 VSUBS 0.006681f
C642 B.n602 VSUBS 0.006681f
C643 B.n603 VSUBS 0.006681f
C644 B.n604 VSUBS 0.006681f
C645 B.n605 VSUBS 0.006681f
C646 B.n606 VSUBS 0.006681f
C647 B.n607 VSUBS 0.006681f
C648 B.n608 VSUBS 0.006681f
C649 B.n609 VSUBS 0.006681f
C650 B.n610 VSUBS 0.006681f
C651 B.n611 VSUBS 0.006681f
C652 B.n612 VSUBS 0.006681f
C653 B.n613 VSUBS 0.006681f
C654 B.n614 VSUBS 0.006681f
C655 B.n615 VSUBS 0.006681f
C656 B.n616 VSUBS 0.006681f
C657 B.n617 VSUBS 0.006681f
C658 B.n618 VSUBS 0.006681f
C659 B.n619 VSUBS 0.004618f
C660 B.n620 VSUBS 0.01548f
C661 B.n621 VSUBS 0.005404f
C662 B.n622 VSUBS 0.006681f
C663 B.n623 VSUBS 0.006681f
C664 B.n624 VSUBS 0.006681f
C665 B.n625 VSUBS 0.006681f
C666 B.n626 VSUBS 0.006681f
C667 B.n627 VSUBS 0.006681f
C668 B.n628 VSUBS 0.006681f
C669 B.n629 VSUBS 0.006681f
C670 B.n630 VSUBS 0.006681f
C671 B.n631 VSUBS 0.006681f
C672 B.n632 VSUBS 0.006681f
C673 B.n633 VSUBS 0.005404f
C674 B.n634 VSUBS 0.01548f
C675 B.n635 VSUBS 0.004618f
C676 B.n636 VSUBS 0.006681f
C677 B.n637 VSUBS 0.006681f
C678 B.n638 VSUBS 0.006681f
C679 B.n639 VSUBS 0.006681f
C680 B.n640 VSUBS 0.006681f
C681 B.n641 VSUBS 0.006681f
C682 B.n642 VSUBS 0.006681f
C683 B.n643 VSUBS 0.006681f
C684 B.n644 VSUBS 0.006681f
C685 B.n645 VSUBS 0.006681f
C686 B.n646 VSUBS 0.006681f
C687 B.n647 VSUBS 0.006681f
C688 B.n648 VSUBS 0.006681f
C689 B.n649 VSUBS 0.006681f
C690 B.n650 VSUBS 0.006681f
C691 B.n651 VSUBS 0.006681f
C692 B.n652 VSUBS 0.006681f
C693 B.n653 VSUBS 0.006681f
C694 B.n654 VSUBS 0.006681f
C695 B.n655 VSUBS 0.006681f
C696 B.n656 VSUBS 0.006681f
C697 B.n657 VSUBS 0.006681f
C698 B.n658 VSUBS 0.006681f
C699 B.n659 VSUBS 0.006681f
C700 B.n660 VSUBS 0.006681f
C701 B.n661 VSUBS 0.006681f
C702 B.n662 VSUBS 0.006681f
C703 B.n663 VSUBS 0.006681f
C704 B.n664 VSUBS 0.006681f
C705 B.n665 VSUBS 0.006681f
C706 B.n666 VSUBS 0.006681f
C707 B.n667 VSUBS 0.006681f
C708 B.n668 VSUBS 0.006681f
C709 B.n669 VSUBS 0.006681f
C710 B.n670 VSUBS 0.006681f
C711 B.n671 VSUBS 0.006681f
C712 B.n672 VSUBS 0.006681f
C713 B.n673 VSUBS 0.006681f
C714 B.n674 VSUBS 0.006681f
C715 B.n675 VSUBS 0.006681f
C716 B.n676 VSUBS 0.006681f
C717 B.n677 VSUBS 0.006681f
C718 B.n678 VSUBS 0.006681f
C719 B.n679 VSUBS 0.006681f
C720 B.n680 VSUBS 0.006681f
C721 B.n681 VSUBS 0.006681f
C722 B.n682 VSUBS 0.006681f
C723 B.n683 VSUBS 0.006681f
C724 B.n684 VSUBS 0.006681f
C725 B.n685 VSUBS 0.006681f
C726 B.n686 VSUBS 0.006681f
C727 B.n687 VSUBS 0.006681f
C728 B.n688 VSUBS 0.006681f
C729 B.n689 VSUBS 0.006681f
C730 B.n690 VSUBS 0.006681f
C731 B.n691 VSUBS 0.006681f
C732 B.n692 VSUBS 0.006681f
C733 B.n693 VSUBS 0.006681f
C734 B.n694 VSUBS 0.006681f
C735 B.n695 VSUBS 0.006681f
C736 B.n696 VSUBS 0.006681f
C737 B.n697 VSUBS 0.006681f
C738 B.n698 VSUBS 0.006681f
C739 B.n699 VSUBS 0.006681f
C740 B.n700 VSUBS 0.006681f
C741 B.n701 VSUBS 0.006681f
C742 B.n702 VSUBS 0.006681f
C743 B.n703 VSUBS 0.006681f
C744 B.n704 VSUBS 0.006681f
C745 B.n705 VSUBS 0.006681f
C746 B.n706 VSUBS 0.015065f
C747 B.n707 VSUBS 0.014411f
C748 B.n708 VSUBS 0.014411f
C749 B.n709 VSUBS 0.006681f
C750 B.n710 VSUBS 0.006681f
C751 B.n711 VSUBS 0.006681f
C752 B.n712 VSUBS 0.006681f
C753 B.n713 VSUBS 0.006681f
C754 B.n714 VSUBS 0.006681f
C755 B.n715 VSUBS 0.006681f
C756 B.n716 VSUBS 0.006681f
C757 B.n717 VSUBS 0.006681f
C758 B.n718 VSUBS 0.006681f
C759 B.n719 VSUBS 0.006681f
C760 B.n720 VSUBS 0.006681f
C761 B.n721 VSUBS 0.006681f
C762 B.n722 VSUBS 0.006681f
C763 B.n723 VSUBS 0.006681f
C764 B.n724 VSUBS 0.006681f
C765 B.n725 VSUBS 0.006681f
C766 B.n726 VSUBS 0.006681f
C767 B.n727 VSUBS 0.006681f
C768 B.n728 VSUBS 0.006681f
C769 B.n729 VSUBS 0.006681f
C770 B.n730 VSUBS 0.006681f
C771 B.n731 VSUBS 0.006681f
C772 B.n732 VSUBS 0.006681f
C773 B.n733 VSUBS 0.006681f
C774 B.n734 VSUBS 0.006681f
C775 B.n735 VSUBS 0.006681f
C776 B.n736 VSUBS 0.006681f
C777 B.n737 VSUBS 0.006681f
C778 B.n738 VSUBS 0.006681f
C779 B.n739 VSUBS 0.006681f
C780 B.n740 VSUBS 0.006681f
C781 B.n741 VSUBS 0.006681f
C782 B.n742 VSUBS 0.006681f
C783 B.n743 VSUBS 0.006681f
C784 B.n744 VSUBS 0.006681f
C785 B.n745 VSUBS 0.006681f
C786 B.n746 VSUBS 0.006681f
C787 B.n747 VSUBS 0.006681f
C788 B.n748 VSUBS 0.006681f
C789 B.n749 VSUBS 0.006681f
C790 B.n750 VSUBS 0.006681f
C791 B.n751 VSUBS 0.006681f
C792 B.n752 VSUBS 0.006681f
C793 B.n753 VSUBS 0.006681f
C794 B.n754 VSUBS 0.006681f
C795 B.n755 VSUBS 0.006681f
C796 B.n756 VSUBS 0.006681f
C797 B.n757 VSUBS 0.006681f
C798 B.n758 VSUBS 0.006681f
C799 B.n759 VSUBS 0.006681f
C800 B.n760 VSUBS 0.006681f
C801 B.n761 VSUBS 0.006681f
C802 B.n762 VSUBS 0.006681f
C803 B.n763 VSUBS 0.006681f
C804 B.n764 VSUBS 0.006681f
C805 B.n765 VSUBS 0.006681f
C806 B.n766 VSUBS 0.006681f
C807 B.n767 VSUBS 0.006681f
C808 B.n768 VSUBS 0.006681f
C809 B.n769 VSUBS 0.006681f
C810 B.n770 VSUBS 0.006681f
C811 B.n771 VSUBS 0.015129f
C812 VDD2.t1 VSUBS 0.29922f
C813 VDD2.t3 VSUBS 0.29922f
C814 VDD2.n0 VSUBS 3.24021f
C815 VDD2.t0 VSUBS 0.29922f
C816 VDD2.t2 VSUBS 0.29922f
C817 VDD2.n1 VSUBS 2.4151f
C818 VDD2.n2 VSUBS 4.75603f
C819 VN.t0 VSUBS 3.96039f
C820 VN.t2 VSUBS 3.97338f
C821 VN.n0 VSUBS 2.40934f
C822 VN.t1 VSUBS 3.97338f
C823 VN.t3 VSUBS 3.96039f
C824 VN.n1 VSUBS 4.17968f
C825 VDD1.t2 VSUBS 0.304219f
C826 VDD1.t3 VSUBS 0.304219f
C827 VDD1.n0 VSUBS 2.45609f
C828 VDD1.t0 VSUBS 0.304219f
C829 VDD1.t1 VSUBS 0.304219f
C830 VDD1.n1 VSUBS 3.32101f
C831 VTAIL.n0 VSUBS 0.024804f
C832 VTAIL.n1 VSUBS 0.023669f
C833 VTAIL.n2 VSUBS 0.013093f
C834 VTAIL.n3 VSUBS 0.030062f
C835 VTAIL.n4 VSUBS 0.013467f
C836 VTAIL.n5 VSUBS 0.023669f
C837 VTAIL.n6 VSUBS 0.012719f
C838 VTAIL.n7 VSUBS 0.030062f
C839 VTAIL.n8 VSUBS 0.013467f
C840 VTAIL.n9 VSUBS 0.023669f
C841 VTAIL.n10 VSUBS 0.012719f
C842 VTAIL.n11 VSUBS 0.030062f
C843 VTAIL.n12 VSUBS 0.013467f
C844 VTAIL.n13 VSUBS 0.023669f
C845 VTAIL.n14 VSUBS 0.012719f
C846 VTAIL.n15 VSUBS 0.030062f
C847 VTAIL.n16 VSUBS 0.013467f
C848 VTAIL.n17 VSUBS 0.023669f
C849 VTAIL.n18 VSUBS 0.012719f
C850 VTAIL.n19 VSUBS 0.030062f
C851 VTAIL.n20 VSUBS 0.013467f
C852 VTAIL.n21 VSUBS 0.023669f
C853 VTAIL.n22 VSUBS 0.012719f
C854 VTAIL.n23 VSUBS 0.022547f
C855 VTAIL.n24 VSUBS 0.019124f
C856 VTAIL.t1 VSUBS 0.064302f
C857 VTAIL.n25 VSUBS 0.160213f
C858 VTAIL.n26 VSUBS 1.40922f
C859 VTAIL.n27 VSUBS 0.012719f
C860 VTAIL.n28 VSUBS 0.013467f
C861 VTAIL.n29 VSUBS 0.030062f
C862 VTAIL.n30 VSUBS 0.030062f
C863 VTAIL.n31 VSUBS 0.013467f
C864 VTAIL.n32 VSUBS 0.012719f
C865 VTAIL.n33 VSUBS 0.023669f
C866 VTAIL.n34 VSUBS 0.023669f
C867 VTAIL.n35 VSUBS 0.012719f
C868 VTAIL.n36 VSUBS 0.013467f
C869 VTAIL.n37 VSUBS 0.030062f
C870 VTAIL.n38 VSUBS 0.030062f
C871 VTAIL.n39 VSUBS 0.013467f
C872 VTAIL.n40 VSUBS 0.012719f
C873 VTAIL.n41 VSUBS 0.023669f
C874 VTAIL.n42 VSUBS 0.023669f
C875 VTAIL.n43 VSUBS 0.012719f
C876 VTAIL.n44 VSUBS 0.013467f
C877 VTAIL.n45 VSUBS 0.030062f
C878 VTAIL.n46 VSUBS 0.030062f
C879 VTAIL.n47 VSUBS 0.013467f
C880 VTAIL.n48 VSUBS 0.012719f
C881 VTAIL.n49 VSUBS 0.023669f
C882 VTAIL.n50 VSUBS 0.023669f
C883 VTAIL.n51 VSUBS 0.012719f
C884 VTAIL.n52 VSUBS 0.013467f
C885 VTAIL.n53 VSUBS 0.030062f
C886 VTAIL.n54 VSUBS 0.030062f
C887 VTAIL.n55 VSUBS 0.013467f
C888 VTAIL.n56 VSUBS 0.012719f
C889 VTAIL.n57 VSUBS 0.023669f
C890 VTAIL.n58 VSUBS 0.023669f
C891 VTAIL.n59 VSUBS 0.012719f
C892 VTAIL.n60 VSUBS 0.013467f
C893 VTAIL.n61 VSUBS 0.030062f
C894 VTAIL.n62 VSUBS 0.030062f
C895 VTAIL.n63 VSUBS 0.013467f
C896 VTAIL.n64 VSUBS 0.012719f
C897 VTAIL.n65 VSUBS 0.023669f
C898 VTAIL.n66 VSUBS 0.023669f
C899 VTAIL.n67 VSUBS 0.012719f
C900 VTAIL.n68 VSUBS 0.012719f
C901 VTAIL.n69 VSUBS 0.013467f
C902 VTAIL.n70 VSUBS 0.030062f
C903 VTAIL.n71 VSUBS 0.030062f
C904 VTAIL.n72 VSUBS 0.068681f
C905 VTAIL.n73 VSUBS 0.013093f
C906 VTAIL.n74 VSUBS 0.012719f
C907 VTAIL.n75 VSUBS 0.058913f
C908 VTAIL.n76 VSUBS 0.034482f
C909 VTAIL.n77 VSUBS 0.188438f
C910 VTAIL.n78 VSUBS 0.024804f
C911 VTAIL.n79 VSUBS 0.023669f
C912 VTAIL.n80 VSUBS 0.013093f
C913 VTAIL.n81 VSUBS 0.030062f
C914 VTAIL.n82 VSUBS 0.013467f
C915 VTAIL.n83 VSUBS 0.023669f
C916 VTAIL.n84 VSUBS 0.012719f
C917 VTAIL.n85 VSUBS 0.030062f
C918 VTAIL.n86 VSUBS 0.013467f
C919 VTAIL.n87 VSUBS 0.023669f
C920 VTAIL.n88 VSUBS 0.012719f
C921 VTAIL.n89 VSUBS 0.030062f
C922 VTAIL.n90 VSUBS 0.013467f
C923 VTAIL.n91 VSUBS 0.023669f
C924 VTAIL.n92 VSUBS 0.012719f
C925 VTAIL.n93 VSUBS 0.030062f
C926 VTAIL.n94 VSUBS 0.013467f
C927 VTAIL.n95 VSUBS 0.023669f
C928 VTAIL.n96 VSUBS 0.012719f
C929 VTAIL.n97 VSUBS 0.030062f
C930 VTAIL.n98 VSUBS 0.013467f
C931 VTAIL.n99 VSUBS 0.023669f
C932 VTAIL.n100 VSUBS 0.012719f
C933 VTAIL.n101 VSUBS 0.022547f
C934 VTAIL.n102 VSUBS 0.019124f
C935 VTAIL.t6 VSUBS 0.064302f
C936 VTAIL.n103 VSUBS 0.160213f
C937 VTAIL.n104 VSUBS 1.40922f
C938 VTAIL.n105 VSUBS 0.012719f
C939 VTAIL.n106 VSUBS 0.013467f
C940 VTAIL.n107 VSUBS 0.030062f
C941 VTAIL.n108 VSUBS 0.030062f
C942 VTAIL.n109 VSUBS 0.013467f
C943 VTAIL.n110 VSUBS 0.012719f
C944 VTAIL.n111 VSUBS 0.023669f
C945 VTAIL.n112 VSUBS 0.023669f
C946 VTAIL.n113 VSUBS 0.012719f
C947 VTAIL.n114 VSUBS 0.013467f
C948 VTAIL.n115 VSUBS 0.030062f
C949 VTAIL.n116 VSUBS 0.030062f
C950 VTAIL.n117 VSUBS 0.013467f
C951 VTAIL.n118 VSUBS 0.012719f
C952 VTAIL.n119 VSUBS 0.023669f
C953 VTAIL.n120 VSUBS 0.023669f
C954 VTAIL.n121 VSUBS 0.012719f
C955 VTAIL.n122 VSUBS 0.013467f
C956 VTAIL.n123 VSUBS 0.030062f
C957 VTAIL.n124 VSUBS 0.030062f
C958 VTAIL.n125 VSUBS 0.013467f
C959 VTAIL.n126 VSUBS 0.012719f
C960 VTAIL.n127 VSUBS 0.023669f
C961 VTAIL.n128 VSUBS 0.023669f
C962 VTAIL.n129 VSUBS 0.012719f
C963 VTAIL.n130 VSUBS 0.013467f
C964 VTAIL.n131 VSUBS 0.030062f
C965 VTAIL.n132 VSUBS 0.030062f
C966 VTAIL.n133 VSUBS 0.013467f
C967 VTAIL.n134 VSUBS 0.012719f
C968 VTAIL.n135 VSUBS 0.023669f
C969 VTAIL.n136 VSUBS 0.023669f
C970 VTAIL.n137 VSUBS 0.012719f
C971 VTAIL.n138 VSUBS 0.013467f
C972 VTAIL.n139 VSUBS 0.030062f
C973 VTAIL.n140 VSUBS 0.030062f
C974 VTAIL.n141 VSUBS 0.013467f
C975 VTAIL.n142 VSUBS 0.012719f
C976 VTAIL.n143 VSUBS 0.023669f
C977 VTAIL.n144 VSUBS 0.023669f
C978 VTAIL.n145 VSUBS 0.012719f
C979 VTAIL.n146 VSUBS 0.012719f
C980 VTAIL.n147 VSUBS 0.013467f
C981 VTAIL.n148 VSUBS 0.030062f
C982 VTAIL.n149 VSUBS 0.030062f
C983 VTAIL.n150 VSUBS 0.068681f
C984 VTAIL.n151 VSUBS 0.013093f
C985 VTAIL.n152 VSUBS 0.012719f
C986 VTAIL.n153 VSUBS 0.058913f
C987 VTAIL.n154 VSUBS 0.034482f
C988 VTAIL.n155 VSUBS 0.309576f
C989 VTAIL.n156 VSUBS 0.024804f
C990 VTAIL.n157 VSUBS 0.023669f
C991 VTAIL.n158 VSUBS 0.013093f
C992 VTAIL.n159 VSUBS 0.030062f
C993 VTAIL.n160 VSUBS 0.013467f
C994 VTAIL.n161 VSUBS 0.023669f
C995 VTAIL.n162 VSUBS 0.012719f
C996 VTAIL.n163 VSUBS 0.030062f
C997 VTAIL.n164 VSUBS 0.013467f
C998 VTAIL.n165 VSUBS 0.023669f
C999 VTAIL.n166 VSUBS 0.012719f
C1000 VTAIL.n167 VSUBS 0.030062f
C1001 VTAIL.n168 VSUBS 0.013467f
C1002 VTAIL.n169 VSUBS 0.023669f
C1003 VTAIL.n170 VSUBS 0.012719f
C1004 VTAIL.n171 VSUBS 0.030062f
C1005 VTAIL.n172 VSUBS 0.013467f
C1006 VTAIL.n173 VSUBS 0.023669f
C1007 VTAIL.n174 VSUBS 0.012719f
C1008 VTAIL.n175 VSUBS 0.030062f
C1009 VTAIL.n176 VSUBS 0.013467f
C1010 VTAIL.n177 VSUBS 0.023669f
C1011 VTAIL.n178 VSUBS 0.012719f
C1012 VTAIL.n179 VSUBS 0.022547f
C1013 VTAIL.n180 VSUBS 0.019124f
C1014 VTAIL.t4 VSUBS 0.064302f
C1015 VTAIL.n181 VSUBS 0.160213f
C1016 VTAIL.n182 VSUBS 1.40922f
C1017 VTAIL.n183 VSUBS 0.012719f
C1018 VTAIL.n184 VSUBS 0.013467f
C1019 VTAIL.n185 VSUBS 0.030062f
C1020 VTAIL.n186 VSUBS 0.030062f
C1021 VTAIL.n187 VSUBS 0.013467f
C1022 VTAIL.n188 VSUBS 0.012719f
C1023 VTAIL.n189 VSUBS 0.023669f
C1024 VTAIL.n190 VSUBS 0.023669f
C1025 VTAIL.n191 VSUBS 0.012719f
C1026 VTAIL.n192 VSUBS 0.013467f
C1027 VTAIL.n193 VSUBS 0.030062f
C1028 VTAIL.n194 VSUBS 0.030062f
C1029 VTAIL.n195 VSUBS 0.013467f
C1030 VTAIL.n196 VSUBS 0.012719f
C1031 VTAIL.n197 VSUBS 0.023669f
C1032 VTAIL.n198 VSUBS 0.023669f
C1033 VTAIL.n199 VSUBS 0.012719f
C1034 VTAIL.n200 VSUBS 0.013467f
C1035 VTAIL.n201 VSUBS 0.030062f
C1036 VTAIL.n202 VSUBS 0.030062f
C1037 VTAIL.n203 VSUBS 0.013467f
C1038 VTAIL.n204 VSUBS 0.012719f
C1039 VTAIL.n205 VSUBS 0.023669f
C1040 VTAIL.n206 VSUBS 0.023669f
C1041 VTAIL.n207 VSUBS 0.012719f
C1042 VTAIL.n208 VSUBS 0.013467f
C1043 VTAIL.n209 VSUBS 0.030062f
C1044 VTAIL.n210 VSUBS 0.030062f
C1045 VTAIL.n211 VSUBS 0.013467f
C1046 VTAIL.n212 VSUBS 0.012719f
C1047 VTAIL.n213 VSUBS 0.023669f
C1048 VTAIL.n214 VSUBS 0.023669f
C1049 VTAIL.n215 VSUBS 0.012719f
C1050 VTAIL.n216 VSUBS 0.013467f
C1051 VTAIL.n217 VSUBS 0.030062f
C1052 VTAIL.n218 VSUBS 0.030062f
C1053 VTAIL.n219 VSUBS 0.013467f
C1054 VTAIL.n220 VSUBS 0.012719f
C1055 VTAIL.n221 VSUBS 0.023669f
C1056 VTAIL.n222 VSUBS 0.023669f
C1057 VTAIL.n223 VSUBS 0.012719f
C1058 VTAIL.n224 VSUBS 0.012719f
C1059 VTAIL.n225 VSUBS 0.013467f
C1060 VTAIL.n226 VSUBS 0.030062f
C1061 VTAIL.n227 VSUBS 0.030062f
C1062 VTAIL.n228 VSUBS 0.068681f
C1063 VTAIL.n229 VSUBS 0.013093f
C1064 VTAIL.n230 VSUBS 0.012719f
C1065 VTAIL.n231 VSUBS 0.058913f
C1066 VTAIL.n232 VSUBS 0.034482f
C1067 VTAIL.n233 VSUBS 1.77015f
C1068 VTAIL.n234 VSUBS 0.024804f
C1069 VTAIL.n235 VSUBS 0.023669f
C1070 VTAIL.n236 VSUBS 0.013093f
C1071 VTAIL.n237 VSUBS 0.030062f
C1072 VTAIL.n238 VSUBS 0.012719f
C1073 VTAIL.n239 VSUBS 0.013467f
C1074 VTAIL.n240 VSUBS 0.023669f
C1075 VTAIL.n241 VSUBS 0.012719f
C1076 VTAIL.n242 VSUBS 0.030062f
C1077 VTAIL.n243 VSUBS 0.013467f
C1078 VTAIL.n244 VSUBS 0.023669f
C1079 VTAIL.n245 VSUBS 0.012719f
C1080 VTAIL.n246 VSUBS 0.030062f
C1081 VTAIL.n247 VSUBS 0.013467f
C1082 VTAIL.n248 VSUBS 0.023669f
C1083 VTAIL.n249 VSUBS 0.012719f
C1084 VTAIL.n250 VSUBS 0.030062f
C1085 VTAIL.n251 VSUBS 0.013467f
C1086 VTAIL.n252 VSUBS 0.023669f
C1087 VTAIL.n253 VSUBS 0.012719f
C1088 VTAIL.n254 VSUBS 0.030062f
C1089 VTAIL.n255 VSUBS 0.013467f
C1090 VTAIL.n256 VSUBS 0.023669f
C1091 VTAIL.n257 VSUBS 0.012719f
C1092 VTAIL.n258 VSUBS 0.022547f
C1093 VTAIL.n259 VSUBS 0.019124f
C1094 VTAIL.t3 VSUBS 0.064302f
C1095 VTAIL.n260 VSUBS 0.160213f
C1096 VTAIL.n261 VSUBS 1.40922f
C1097 VTAIL.n262 VSUBS 0.012719f
C1098 VTAIL.n263 VSUBS 0.013467f
C1099 VTAIL.n264 VSUBS 0.030062f
C1100 VTAIL.n265 VSUBS 0.030062f
C1101 VTAIL.n266 VSUBS 0.013467f
C1102 VTAIL.n267 VSUBS 0.012719f
C1103 VTAIL.n268 VSUBS 0.023669f
C1104 VTAIL.n269 VSUBS 0.023669f
C1105 VTAIL.n270 VSUBS 0.012719f
C1106 VTAIL.n271 VSUBS 0.013467f
C1107 VTAIL.n272 VSUBS 0.030062f
C1108 VTAIL.n273 VSUBS 0.030062f
C1109 VTAIL.n274 VSUBS 0.013467f
C1110 VTAIL.n275 VSUBS 0.012719f
C1111 VTAIL.n276 VSUBS 0.023669f
C1112 VTAIL.n277 VSUBS 0.023669f
C1113 VTAIL.n278 VSUBS 0.012719f
C1114 VTAIL.n279 VSUBS 0.013467f
C1115 VTAIL.n280 VSUBS 0.030062f
C1116 VTAIL.n281 VSUBS 0.030062f
C1117 VTAIL.n282 VSUBS 0.013467f
C1118 VTAIL.n283 VSUBS 0.012719f
C1119 VTAIL.n284 VSUBS 0.023669f
C1120 VTAIL.n285 VSUBS 0.023669f
C1121 VTAIL.n286 VSUBS 0.012719f
C1122 VTAIL.n287 VSUBS 0.013467f
C1123 VTAIL.n288 VSUBS 0.030062f
C1124 VTAIL.n289 VSUBS 0.030062f
C1125 VTAIL.n290 VSUBS 0.013467f
C1126 VTAIL.n291 VSUBS 0.012719f
C1127 VTAIL.n292 VSUBS 0.023669f
C1128 VTAIL.n293 VSUBS 0.023669f
C1129 VTAIL.n294 VSUBS 0.012719f
C1130 VTAIL.n295 VSUBS 0.013467f
C1131 VTAIL.n296 VSUBS 0.030062f
C1132 VTAIL.n297 VSUBS 0.030062f
C1133 VTAIL.n298 VSUBS 0.013467f
C1134 VTAIL.n299 VSUBS 0.012719f
C1135 VTAIL.n300 VSUBS 0.023669f
C1136 VTAIL.n301 VSUBS 0.023669f
C1137 VTAIL.n302 VSUBS 0.012719f
C1138 VTAIL.n303 VSUBS 0.013467f
C1139 VTAIL.n304 VSUBS 0.030062f
C1140 VTAIL.n305 VSUBS 0.030062f
C1141 VTAIL.n306 VSUBS 0.068681f
C1142 VTAIL.n307 VSUBS 0.013093f
C1143 VTAIL.n308 VSUBS 0.012719f
C1144 VTAIL.n309 VSUBS 0.058913f
C1145 VTAIL.n310 VSUBS 0.034482f
C1146 VTAIL.n311 VSUBS 1.77015f
C1147 VTAIL.n312 VSUBS 0.024804f
C1148 VTAIL.n313 VSUBS 0.023669f
C1149 VTAIL.n314 VSUBS 0.013093f
C1150 VTAIL.n315 VSUBS 0.030062f
C1151 VTAIL.n316 VSUBS 0.012719f
C1152 VTAIL.n317 VSUBS 0.013467f
C1153 VTAIL.n318 VSUBS 0.023669f
C1154 VTAIL.n319 VSUBS 0.012719f
C1155 VTAIL.n320 VSUBS 0.030062f
C1156 VTAIL.n321 VSUBS 0.013467f
C1157 VTAIL.n322 VSUBS 0.023669f
C1158 VTAIL.n323 VSUBS 0.012719f
C1159 VTAIL.n324 VSUBS 0.030062f
C1160 VTAIL.n325 VSUBS 0.013467f
C1161 VTAIL.n326 VSUBS 0.023669f
C1162 VTAIL.n327 VSUBS 0.012719f
C1163 VTAIL.n328 VSUBS 0.030062f
C1164 VTAIL.n329 VSUBS 0.013467f
C1165 VTAIL.n330 VSUBS 0.023669f
C1166 VTAIL.n331 VSUBS 0.012719f
C1167 VTAIL.n332 VSUBS 0.030062f
C1168 VTAIL.n333 VSUBS 0.013467f
C1169 VTAIL.n334 VSUBS 0.023669f
C1170 VTAIL.n335 VSUBS 0.012719f
C1171 VTAIL.n336 VSUBS 0.022547f
C1172 VTAIL.n337 VSUBS 0.019124f
C1173 VTAIL.t2 VSUBS 0.064302f
C1174 VTAIL.n338 VSUBS 0.160213f
C1175 VTAIL.n339 VSUBS 1.40922f
C1176 VTAIL.n340 VSUBS 0.012719f
C1177 VTAIL.n341 VSUBS 0.013467f
C1178 VTAIL.n342 VSUBS 0.030062f
C1179 VTAIL.n343 VSUBS 0.030062f
C1180 VTAIL.n344 VSUBS 0.013467f
C1181 VTAIL.n345 VSUBS 0.012719f
C1182 VTAIL.n346 VSUBS 0.023669f
C1183 VTAIL.n347 VSUBS 0.023669f
C1184 VTAIL.n348 VSUBS 0.012719f
C1185 VTAIL.n349 VSUBS 0.013467f
C1186 VTAIL.n350 VSUBS 0.030062f
C1187 VTAIL.n351 VSUBS 0.030062f
C1188 VTAIL.n352 VSUBS 0.013467f
C1189 VTAIL.n353 VSUBS 0.012719f
C1190 VTAIL.n354 VSUBS 0.023669f
C1191 VTAIL.n355 VSUBS 0.023669f
C1192 VTAIL.n356 VSUBS 0.012719f
C1193 VTAIL.n357 VSUBS 0.013467f
C1194 VTAIL.n358 VSUBS 0.030062f
C1195 VTAIL.n359 VSUBS 0.030062f
C1196 VTAIL.n360 VSUBS 0.013467f
C1197 VTAIL.n361 VSUBS 0.012719f
C1198 VTAIL.n362 VSUBS 0.023669f
C1199 VTAIL.n363 VSUBS 0.023669f
C1200 VTAIL.n364 VSUBS 0.012719f
C1201 VTAIL.n365 VSUBS 0.013467f
C1202 VTAIL.n366 VSUBS 0.030062f
C1203 VTAIL.n367 VSUBS 0.030062f
C1204 VTAIL.n368 VSUBS 0.013467f
C1205 VTAIL.n369 VSUBS 0.012719f
C1206 VTAIL.n370 VSUBS 0.023669f
C1207 VTAIL.n371 VSUBS 0.023669f
C1208 VTAIL.n372 VSUBS 0.012719f
C1209 VTAIL.n373 VSUBS 0.013467f
C1210 VTAIL.n374 VSUBS 0.030062f
C1211 VTAIL.n375 VSUBS 0.030062f
C1212 VTAIL.n376 VSUBS 0.013467f
C1213 VTAIL.n377 VSUBS 0.012719f
C1214 VTAIL.n378 VSUBS 0.023669f
C1215 VTAIL.n379 VSUBS 0.023669f
C1216 VTAIL.n380 VSUBS 0.012719f
C1217 VTAIL.n381 VSUBS 0.013467f
C1218 VTAIL.n382 VSUBS 0.030062f
C1219 VTAIL.n383 VSUBS 0.030062f
C1220 VTAIL.n384 VSUBS 0.068681f
C1221 VTAIL.n385 VSUBS 0.013093f
C1222 VTAIL.n386 VSUBS 0.012719f
C1223 VTAIL.n387 VSUBS 0.058913f
C1224 VTAIL.n388 VSUBS 0.034482f
C1225 VTAIL.n389 VSUBS 0.309576f
C1226 VTAIL.n390 VSUBS 0.024804f
C1227 VTAIL.n391 VSUBS 0.023669f
C1228 VTAIL.n392 VSUBS 0.013093f
C1229 VTAIL.n393 VSUBS 0.030062f
C1230 VTAIL.n394 VSUBS 0.012719f
C1231 VTAIL.n395 VSUBS 0.013467f
C1232 VTAIL.n396 VSUBS 0.023669f
C1233 VTAIL.n397 VSUBS 0.012719f
C1234 VTAIL.n398 VSUBS 0.030062f
C1235 VTAIL.n399 VSUBS 0.013467f
C1236 VTAIL.n400 VSUBS 0.023669f
C1237 VTAIL.n401 VSUBS 0.012719f
C1238 VTAIL.n402 VSUBS 0.030062f
C1239 VTAIL.n403 VSUBS 0.013467f
C1240 VTAIL.n404 VSUBS 0.023669f
C1241 VTAIL.n405 VSUBS 0.012719f
C1242 VTAIL.n406 VSUBS 0.030062f
C1243 VTAIL.n407 VSUBS 0.013467f
C1244 VTAIL.n408 VSUBS 0.023669f
C1245 VTAIL.n409 VSUBS 0.012719f
C1246 VTAIL.n410 VSUBS 0.030062f
C1247 VTAIL.n411 VSUBS 0.013467f
C1248 VTAIL.n412 VSUBS 0.023669f
C1249 VTAIL.n413 VSUBS 0.012719f
C1250 VTAIL.n414 VSUBS 0.022547f
C1251 VTAIL.n415 VSUBS 0.019124f
C1252 VTAIL.t7 VSUBS 0.064302f
C1253 VTAIL.n416 VSUBS 0.160213f
C1254 VTAIL.n417 VSUBS 1.40922f
C1255 VTAIL.n418 VSUBS 0.012719f
C1256 VTAIL.n419 VSUBS 0.013467f
C1257 VTAIL.n420 VSUBS 0.030062f
C1258 VTAIL.n421 VSUBS 0.030062f
C1259 VTAIL.n422 VSUBS 0.013467f
C1260 VTAIL.n423 VSUBS 0.012719f
C1261 VTAIL.n424 VSUBS 0.023669f
C1262 VTAIL.n425 VSUBS 0.023669f
C1263 VTAIL.n426 VSUBS 0.012719f
C1264 VTAIL.n427 VSUBS 0.013467f
C1265 VTAIL.n428 VSUBS 0.030062f
C1266 VTAIL.n429 VSUBS 0.030062f
C1267 VTAIL.n430 VSUBS 0.013467f
C1268 VTAIL.n431 VSUBS 0.012719f
C1269 VTAIL.n432 VSUBS 0.023669f
C1270 VTAIL.n433 VSUBS 0.023669f
C1271 VTAIL.n434 VSUBS 0.012719f
C1272 VTAIL.n435 VSUBS 0.013467f
C1273 VTAIL.n436 VSUBS 0.030062f
C1274 VTAIL.n437 VSUBS 0.030062f
C1275 VTAIL.n438 VSUBS 0.013467f
C1276 VTAIL.n439 VSUBS 0.012719f
C1277 VTAIL.n440 VSUBS 0.023669f
C1278 VTAIL.n441 VSUBS 0.023669f
C1279 VTAIL.n442 VSUBS 0.012719f
C1280 VTAIL.n443 VSUBS 0.013467f
C1281 VTAIL.n444 VSUBS 0.030062f
C1282 VTAIL.n445 VSUBS 0.030062f
C1283 VTAIL.n446 VSUBS 0.013467f
C1284 VTAIL.n447 VSUBS 0.012719f
C1285 VTAIL.n448 VSUBS 0.023669f
C1286 VTAIL.n449 VSUBS 0.023669f
C1287 VTAIL.n450 VSUBS 0.012719f
C1288 VTAIL.n451 VSUBS 0.013467f
C1289 VTAIL.n452 VSUBS 0.030062f
C1290 VTAIL.n453 VSUBS 0.030062f
C1291 VTAIL.n454 VSUBS 0.013467f
C1292 VTAIL.n455 VSUBS 0.012719f
C1293 VTAIL.n456 VSUBS 0.023669f
C1294 VTAIL.n457 VSUBS 0.023669f
C1295 VTAIL.n458 VSUBS 0.012719f
C1296 VTAIL.n459 VSUBS 0.013467f
C1297 VTAIL.n460 VSUBS 0.030062f
C1298 VTAIL.n461 VSUBS 0.030062f
C1299 VTAIL.n462 VSUBS 0.068681f
C1300 VTAIL.n463 VSUBS 0.013093f
C1301 VTAIL.n464 VSUBS 0.012719f
C1302 VTAIL.n465 VSUBS 0.058913f
C1303 VTAIL.n466 VSUBS 0.034482f
C1304 VTAIL.n467 VSUBS 0.309576f
C1305 VTAIL.n468 VSUBS 0.024804f
C1306 VTAIL.n469 VSUBS 0.023669f
C1307 VTAIL.n470 VSUBS 0.013093f
C1308 VTAIL.n471 VSUBS 0.030062f
C1309 VTAIL.n472 VSUBS 0.012719f
C1310 VTAIL.n473 VSUBS 0.013467f
C1311 VTAIL.n474 VSUBS 0.023669f
C1312 VTAIL.n475 VSUBS 0.012719f
C1313 VTAIL.n476 VSUBS 0.030062f
C1314 VTAIL.n477 VSUBS 0.013467f
C1315 VTAIL.n478 VSUBS 0.023669f
C1316 VTAIL.n479 VSUBS 0.012719f
C1317 VTAIL.n480 VSUBS 0.030062f
C1318 VTAIL.n481 VSUBS 0.013467f
C1319 VTAIL.n482 VSUBS 0.023669f
C1320 VTAIL.n483 VSUBS 0.012719f
C1321 VTAIL.n484 VSUBS 0.030062f
C1322 VTAIL.n485 VSUBS 0.013467f
C1323 VTAIL.n486 VSUBS 0.023669f
C1324 VTAIL.n487 VSUBS 0.012719f
C1325 VTAIL.n488 VSUBS 0.030062f
C1326 VTAIL.n489 VSUBS 0.013467f
C1327 VTAIL.n490 VSUBS 0.023669f
C1328 VTAIL.n491 VSUBS 0.012719f
C1329 VTAIL.n492 VSUBS 0.022547f
C1330 VTAIL.n493 VSUBS 0.019124f
C1331 VTAIL.t5 VSUBS 0.064302f
C1332 VTAIL.n494 VSUBS 0.160213f
C1333 VTAIL.n495 VSUBS 1.40922f
C1334 VTAIL.n496 VSUBS 0.012719f
C1335 VTAIL.n497 VSUBS 0.013467f
C1336 VTAIL.n498 VSUBS 0.030062f
C1337 VTAIL.n499 VSUBS 0.030062f
C1338 VTAIL.n500 VSUBS 0.013467f
C1339 VTAIL.n501 VSUBS 0.012719f
C1340 VTAIL.n502 VSUBS 0.023669f
C1341 VTAIL.n503 VSUBS 0.023669f
C1342 VTAIL.n504 VSUBS 0.012719f
C1343 VTAIL.n505 VSUBS 0.013467f
C1344 VTAIL.n506 VSUBS 0.030062f
C1345 VTAIL.n507 VSUBS 0.030062f
C1346 VTAIL.n508 VSUBS 0.013467f
C1347 VTAIL.n509 VSUBS 0.012719f
C1348 VTAIL.n510 VSUBS 0.023669f
C1349 VTAIL.n511 VSUBS 0.023669f
C1350 VTAIL.n512 VSUBS 0.012719f
C1351 VTAIL.n513 VSUBS 0.013467f
C1352 VTAIL.n514 VSUBS 0.030062f
C1353 VTAIL.n515 VSUBS 0.030062f
C1354 VTAIL.n516 VSUBS 0.013467f
C1355 VTAIL.n517 VSUBS 0.012719f
C1356 VTAIL.n518 VSUBS 0.023669f
C1357 VTAIL.n519 VSUBS 0.023669f
C1358 VTAIL.n520 VSUBS 0.012719f
C1359 VTAIL.n521 VSUBS 0.013467f
C1360 VTAIL.n522 VSUBS 0.030062f
C1361 VTAIL.n523 VSUBS 0.030062f
C1362 VTAIL.n524 VSUBS 0.013467f
C1363 VTAIL.n525 VSUBS 0.012719f
C1364 VTAIL.n526 VSUBS 0.023669f
C1365 VTAIL.n527 VSUBS 0.023669f
C1366 VTAIL.n528 VSUBS 0.012719f
C1367 VTAIL.n529 VSUBS 0.013467f
C1368 VTAIL.n530 VSUBS 0.030062f
C1369 VTAIL.n531 VSUBS 0.030062f
C1370 VTAIL.n532 VSUBS 0.013467f
C1371 VTAIL.n533 VSUBS 0.012719f
C1372 VTAIL.n534 VSUBS 0.023669f
C1373 VTAIL.n535 VSUBS 0.023669f
C1374 VTAIL.n536 VSUBS 0.012719f
C1375 VTAIL.n537 VSUBS 0.013467f
C1376 VTAIL.n538 VSUBS 0.030062f
C1377 VTAIL.n539 VSUBS 0.030062f
C1378 VTAIL.n540 VSUBS 0.068681f
C1379 VTAIL.n541 VSUBS 0.013093f
C1380 VTAIL.n542 VSUBS 0.012719f
C1381 VTAIL.n543 VSUBS 0.058913f
C1382 VTAIL.n544 VSUBS 0.034482f
C1383 VTAIL.n545 VSUBS 1.77015f
C1384 VTAIL.n546 VSUBS 0.024804f
C1385 VTAIL.n547 VSUBS 0.023669f
C1386 VTAIL.n548 VSUBS 0.013093f
C1387 VTAIL.n549 VSUBS 0.030062f
C1388 VTAIL.n550 VSUBS 0.013467f
C1389 VTAIL.n551 VSUBS 0.023669f
C1390 VTAIL.n552 VSUBS 0.012719f
C1391 VTAIL.n553 VSUBS 0.030062f
C1392 VTAIL.n554 VSUBS 0.013467f
C1393 VTAIL.n555 VSUBS 0.023669f
C1394 VTAIL.n556 VSUBS 0.012719f
C1395 VTAIL.n557 VSUBS 0.030062f
C1396 VTAIL.n558 VSUBS 0.013467f
C1397 VTAIL.n559 VSUBS 0.023669f
C1398 VTAIL.n560 VSUBS 0.012719f
C1399 VTAIL.n561 VSUBS 0.030062f
C1400 VTAIL.n562 VSUBS 0.013467f
C1401 VTAIL.n563 VSUBS 0.023669f
C1402 VTAIL.n564 VSUBS 0.012719f
C1403 VTAIL.n565 VSUBS 0.030062f
C1404 VTAIL.n566 VSUBS 0.013467f
C1405 VTAIL.n567 VSUBS 0.023669f
C1406 VTAIL.n568 VSUBS 0.012719f
C1407 VTAIL.n569 VSUBS 0.022547f
C1408 VTAIL.n570 VSUBS 0.019124f
C1409 VTAIL.t0 VSUBS 0.064302f
C1410 VTAIL.n571 VSUBS 0.160213f
C1411 VTAIL.n572 VSUBS 1.40922f
C1412 VTAIL.n573 VSUBS 0.012719f
C1413 VTAIL.n574 VSUBS 0.013467f
C1414 VTAIL.n575 VSUBS 0.030062f
C1415 VTAIL.n576 VSUBS 0.030062f
C1416 VTAIL.n577 VSUBS 0.013467f
C1417 VTAIL.n578 VSUBS 0.012719f
C1418 VTAIL.n579 VSUBS 0.023669f
C1419 VTAIL.n580 VSUBS 0.023669f
C1420 VTAIL.n581 VSUBS 0.012719f
C1421 VTAIL.n582 VSUBS 0.013467f
C1422 VTAIL.n583 VSUBS 0.030062f
C1423 VTAIL.n584 VSUBS 0.030062f
C1424 VTAIL.n585 VSUBS 0.013467f
C1425 VTAIL.n586 VSUBS 0.012719f
C1426 VTAIL.n587 VSUBS 0.023669f
C1427 VTAIL.n588 VSUBS 0.023669f
C1428 VTAIL.n589 VSUBS 0.012719f
C1429 VTAIL.n590 VSUBS 0.013467f
C1430 VTAIL.n591 VSUBS 0.030062f
C1431 VTAIL.n592 VSUBS 0.030062f
C1432 VTAIL.n593 VSUBS 0.013467f
C1433 VTAIL.n594 VSUBS 0.012719f
C1434 VTAIL.n595 VSUBS 0.023669f
C1435 VTAIL.n596 VSUBS 0.023669f
C1436 VTAIL.n597 VSUBS 0.012719f
C1437 VTAIL.n598 VSUBS 0.013467f
C1438 VTAIL.n599 VSUBS 0.030062f
C1439 VTAIL.n600 VSUBS 0.030062f
C1440 VTAIL.n601 VSUBS 0.013467f
C1441 VTAIL.n602 VSUBS 0.012719f
C1442 VTAIL.n603 VSUBS 0.023669f
C1443 VTAIL.n604 VSUBS 0.023669f
C1444 VTAIL.n605 VSUBS 0.012719f
C1445 VTAIL.n606 VSUBS 0.013467f
C1446 VTAIL.n607 VSUBS 0.030062f
C1447 VTAIL.n608 VSUBS 0.030062f
C1448 VTAIL.n609 VSUBS 0.013467f
C1449 VTAIL.n610 VSUBS 0.012719f
C1450 VTAIL.n611 VSUBS 0.023669f
C1451 VTAIL.n612 VSUBS 0.023669f
C1452 VTAIL.n613 VSUBS 0.012719f
C1453 VTAIL.n614 VSUBS 0.012719f
C1454 VTAIL.n615 VSUBS 0.013467f
C1455 VTAIL.n616 VSUBS 0.030062f
C1456 VTAIL.n617 VSUBS 0.030062f
C1457 VTAIL.n618 VSUBS 0.068681f
C1458 VTAIL.n619 VSUBS 0.013093f
C1459 VTAIL.n620 VSUBS 0.012719f
C1460 VTAIL.n621 VSUBS 0.058913f
C1461 VTAIL.n622 VSUBS 0.034482f
C1462 VTAIL.n623 VSUBS 1.64014f
C1463 VP.t2 VSUBS 4.01f
C1464 VP.n0 VSUBS 1.50795f
C1465 VP.n1 VSUBS 0.02989f
C1466 VP.n2 VSUBS 0.043634f
C1467 VP.n3 VSUBS 0.02989f
C1468 VP.n4 VSUBS 0.037006f
C1469 VP.t1 VSUBS 4.43618f
C1470 VP.t0 VSUBS 4.42168f
C1471 VP.n5 VSUBS 4.65456f
C1472 VP.t3 VSUBS 4.01f
C1473 VP.n6 VSUBS 1.50795f
C1474 VP.n7 VSUBS 1.85063f
C1475 VP.n8 VSUBS 0.048242f
C1476 VP.n9 VSUBS 0.02989f
C1477 VP.n10 VSUBS 0.055708f
C1478 VP.n11 VSUBS 0.055708f
C1479 VP.n12 VSUBS 0.043634f
C1480 VP.n13 VSUBS 0.02989f
C1481 VP.n14 VSUBS 0.02989f
C1482 VP.n15 VSUBS 0.02989f
C1483 VP.n16 VSUBS 0.055708f
C1484 VP.n17 VSUBS 0.055708f
C1485 VP.n18 VSUBS 0.037006f
C1486 VP.n19 VSUBS 0.048242f
C1487 VP.n20 VSUBS 0.082338f
.ends

