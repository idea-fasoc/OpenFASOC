* NGSPICE file created from diff_pair_sample_1505.ext - technology: sky130A

.subckt diff_pair_sample_1505 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=6.5442 pd=34.34 as=0 ps=0 w=16.78 l=1.92
X1 B.t8 B.t6 B.t7 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=6.5442 pd=34.34 as=0 ps=0 w=16.78 l=1.92
X2 VTAIL.t11 VN.t0 VDD2.t1 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=2.7687 pd=17.11 as=2.7687 ps=17.11 w=16.78 l=1.92
X3 B.t5 B.t3 B.t4 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=6.5442 pd=34.34 as=0 ps=0 w=16.78 l=1.92
X4 VDD1.t5 VP.t0 VTAIL.t5 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=6.5442 pd=34.34 as=2.7687 ps=17.11 w=16.78 l=1.92
X5 B.t2 B.t0 B.t1 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=6.5442 pd=34.34 as=0 ps=0 w=16.78 l=1.92
X6 VDD2.t3 VN.t1 VTAIL.t10 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=2.7687 pd=17.11 as=6.5442 ps=34.34 w=16.78 l=1.92
X7 VDD1.t4 VP.t1 VTAIL.t4 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=6.5442 pd=34.34 as=2.7687 ps=17.11 w=16.78 l=1.92
X8 VDD1.t3 VP.t2 VTAIL.t3 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=2.7687 pd=17.11 as=6.5442 ps=34.34 w=16.78 l=1.92
X9 VDD1.t2 VP.t3 VTAIL.t1 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=2.7687 pd=17.11 as=6.5442 ps=34.34 w=16.78 l=1.92
X10 VDD2.t0 VN.t2 VTAIL.t9 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=6.5442 pd=34.34 as=2.7687 ps=17.11 w=16.78 l=1.92
X11 VDD2.t5 VN.t3 VTAIL.t8 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=6.5442 pd=34.34 as=2.7687 ps=17.11 w=16.78 l=1.92
X12 VTAIL.t2 VP.t4 VDD1.t1 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=2.7687 pd=17.11 as=2.7687 ps=17.11 w=16.78 l=1.92
X13 VDD2.t2 VN.t4 VTAIL.t7 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=2.7687 pd=17.11 as=6.5442 ps=34.34 w=16.78 l=1.92
X14 VTAIL.t0 VP.t5 VDD1.t0 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=2.7687 pd=17.11 as=2.7687 ps=17.11 w=16.78 l=1.92
X15 VTAIL.t6 VN.t5 VDD2.t4 w_n2770_n4324# sky130_fd_pr__pfet_01v8 ad=2.7687 pd=17.11 as=2.7687 ps=17.11 w=16.78 l=1.92
R0 B.n432 B.n431 585
R1 B.n430 B.n119 585
R2 B.n429 B.n428 585
R3 B.n427 B.n120 585
R4 B.n426 B.n425 585
R5 B.n424 B.n121 585
R6 B.n423 B.n422 585
R7 B.n421 B.n122 585
R8 B.n420 B.n419 585
R9 B.n418 B.n123 585
R10 B.n417 B.n416 585
R11 B.n415 B.n124 585
R12 B.n414 B.n413 585
R13 B.n412 B.n125 585
R14 B.n411 B.n410 585
R15 B.n409 B.n126 585
R16 B.n408 B.n407 585
R17 B.n406 B.n127 585
R18 B.n405 B.n404 585
R19 B.n403 B.n128 585
R20 B.n402 B.n401 585
R21 B.n400 B.n129 585
R22 B.n399 B.n398 585
R23 B.n397 B.n130 585
R24 B.n396 B.n395 585
R25 B.n394 B.n131 585
R26 B.n393 B.n392 585
R27 B.n391 B.n132 585
R28 B.n390 B.n389 585
R29 B.n388 B.n133 585
R30 B.n387 B.n386 585
R31 B.n385 B.n134 585
R32 B.n384 B.n383 585
R33 B.n382 B.n135 585
R34 B.n381 B.n380 585
R35 B.n379 B.n136 585
R36 B.n378 B.n377 585
R37 B.n376 B.n137 585
R38 B.n375 B.n374 585
R39 B.n373 B.n138 585
R40 B.n372 B.n371 585
R41 B.n370 B.n139 585
R42 B.n369 B.n368 585
R43 B.n367 B.n140 585
R44 B.n366 B.n365 585
R45 B.n364 B.n141 585
R46 B.n363 B.n362 585
R47 B.n361 B.n142 585
R48 B.n360 B.n359 585
R49 B.n358 B.n143 585
R50 B.n357 B.n356 585
R51 B.n355 B.n144 585
R52 B.n354 B.n353 585
R53 B.n352 B.n145 585
R54 B.n351 B.n350 585
R55 B.n349 B.n146 585
R56 B.n348 B.n347 585
R57 B.n343 B.n147 585
R58 B.n342 B.n341 585
R59 B.n340 B.n148 585
R60 B.n339 B.n338 585
R61 B.n337 B.n149 585
R62 B.n336 B.n335 585
R63 B.n334 B.n150 585
R64 B.n333 B.n332 585
R65 B.n330 B.n151 585
R66 B.n329 B.n328 585
R67 B.n327 B.n154 585
R68 B.n326 B.n325 585
R69 B.n324 B.n155 585
R70 B.n323 B.n322 585
R71 B.n321 B.n156 585
R72 B.n320 B.n319 585
R73 B.n318 B.n157 585
R74 B.n317 B.n316 585
R75 B.n315 B.n158 585
R76 B.n314 B.n313 585
R77 B.n312 B.n159 585
R78 B.n311 B.n310 585
R79 B.n309 B.n160 585
R80 B.n308 B.n307 585
R81 B.n306 B.n161 585
R82 B.n305 B.n304 585
R83 B.n303 B.n162 585
R84 B.n302 B.n301 585
R85 B.n300 B.n163 585
R86 B.n299 B.n298 585
R87 B.n297 B.n164 585
R88 B.n296 B.n295 585
R89 B.n294 B.n165 585
R90 B.n293 B.n292 585
R91 B.n291 B.n166 585
R92 B.n290 B.n289 585
R93 B.n288 B.n167 585
R94 B.n287 B.n286 585
R95 B.n285 B.n168 585
R96 B.n284 B.n283 585
R97 B.n282 B.n169 585
R98 B.n281 B.n280 585
R99 B.n279 B.n170 585
R100 B.n278 B.n277 585
R101 B.n276 B.n171 585
R102 B.n275 B.n274 585
R103 B.n273 B.n172 585
R104 B.n272 B.n271 585
R105 B.n270 B.n173 585
R106 B.n269 B.n268 585
R107 B.n267 B.n174 585
R108 B.n266 B.n265 585
R109 B.n264 B.n175 585
R110 B.n263 B.n262 585
R111 B.n261 B.n176 585
R112 B.n260 B.n259 585
R113 B.n258 B.n177 585
R114 B.n257 B.n256 585
R115 B.n255 B.n178 585
R116 B.n254 B.n253 585
R117 B.n252 B.n179 585
R118 B.n251 B.n250 585
R119 B.n249 B.n180 585
R120 B.n248 B.n247 585
R121 B.n433 B.n118 585
R122 B.n435 B.n434 585
R123 B.n436 B.n117 585
R124 B.n438 B.n437 585
R125 B.n439 B.n116 585
R126 B.n441 B.n440 585
R127 B.n442 B.n115 585
R128 B.n444 B.n443 585
R129 B.n445 B.n114 585
R130 B.n447 B.n446 585
R131 B.n448 B.n113 585
R132 B.n450 B.n449 585
R133 B.n451 B.n112 585
R134 B.n453 B.n452 585
R135 B.n454 B.n111 585
R136 B.n456 B.n455 585
R137 B.n457 B.n110 585
R138 B.n459 B.n458 585
R139 B.n460 B.n109 585
R140 B.n462 B.n461 585
R141 B.n463 B.n108 585
R142 B.n465 B.n464 585
R143 B.n466 B.n107 585
R144 B.n468 B.n467 585
R145 B.n469 B.n106 585
R146 B.n471 B.n470 585
R147 B.n472 B.n105 585
R148 B.n474 B.n473 585
R149 B.n475 B.n104 585
R150 B.n477 B.n476 585
R151 B.n478 B.n103 585
R152 B.n480 B.n479 585
R153 B.n481 B.n102 585
R154 B.n483 B.n482 585
R155 B.n484 B.n101 585
R156 B.n486 B.n485 585
R157 B.n487 B.n100 585
R158 B.n489 B.n488 585
R159 B.n490 B.n99 585
R160 B.n492 B.n491 585
R161 B.n493 B.n98 585
R162 B.n495 B.n494 585
R163 B.n496 B.n97 585
R164 B.n498 B.n497 585
R165 B.n499 B.n96 585
R166 B.n501 B.n500 585
R167 B.n502 B.n95 585
R168 B.n504 B.n503 585
R169 B.n505 B.n94 585
R170 B.n507 B.n506 585
R171 B.n508 B.n93 585
R172 B.n510 B.n509 585
R173 B.n511 B.n92 585
R174 B.n513 B.n512 585
R175 B.n514 B.n91 585
R176 B.n516 B.n515 585
R177 B.n517 B.n90 585
R178 B.n519 B.n518 585
R179 B.n520 B.n89 585
R180 B.n522 B.n521 585
R181 B.n523 B.n88 585
R182 B.n525 B.n524 585
R183 B.n526 B.n87 585
R184 B.n528 B.n527 585
R185 B.n529 B.n86 585
R186 B.n531 B.n530 585
R187 B.n532 B.n85 585
R188 B.n534 B.n533 585
R189 B.n535 B.n84 585
R190 B.n537 B.n536 585
R191 B.n720 B.n19 585
R192 B.n719 B.n718 585
R193 B.n717 B.n20 585
R194 B.n716 B.n715 585
R195 B.n714 B.n21 585
R196 B.n713 B.n712 585
R197 B.n711 B.n22 585
R198 B.n710 B.n709 585
R199 B.n708 B.n23 585
R200 B.n707 B.n706 585
R201 B.n705 B.n24 585
R202 B.n704 B.n703 585
R203 B.n702 B.n25 585
R204 B.n701 B.n700 585
R205 B.n699 B.n26 585
R206 B.n698 B.n697 585
R207 B.n696 B.n27 585
R208 B.n695 B.n694 585
R209 B.n693 B.n28 585
R210 B.n692 B.n691 585
R211 B.n690 B.n29 585
R212 B.n689 B.n688 585
R213 B.n687 B.n30 585
R214 B.n686 B.n685 585
R215 B.n684 B.n31 585
R216 B.n683 B.n682 585
R217 B.n681 B.n32 585
R218 B.n680 B.n679 585
R219 B.n678 B.n33 585
R220 B.n677 B.n676 585
R221 B.n675 B.n34 585
R222 B.n674 B.n673 585
R223 B.n672 B.n35 585
R224 B.n671 B.n670 585
R225 B.n669 B.n36 585
R226 B.n668 B.n667 585
R227 B.n666 B.n37 585
R228 B.n665 B.n664 585
R229 B.n663 B.n38 585
R230 B.n662 B.n661 585
R231 B.n660 B.n39 585
R232 B.n659 B.n658 585
R233 B.n657 B.n40 585
R234 B.n656 B.n655 585
R235 B.n654 B.n41 585
R236 B.n653 B.n652 585
R237 B.n651 B.n42 585
R238 B.n650 B.n649 585
R239 B.n648 B.n43 585
R240 B.n647 B.n646 585
R241 B.n645 B.n44 585
R242 B.n644 B.n643 585
R243 B.n642 B.n45 585
R244 B.n641 B.n640 585
R245 B.n639 B.n46 585
R246 B.n638 B.n637 585
R247 B.n635 B.n47 585
R248 B.n634 B.n633 585
R249 B.n632 B.n50 585
R250 B.n631 B.n630 585
R251 B.n629 B.n51 585
R252 B.n628 B.n627 585
R253 B.n626 B.n52 585
R254 B.n625 B.n624 585
R255 B.n623 B.n53 585
R256 B.n621 B.n620 585
R257 B.n619 B.n56 585
R258 B.n618 B.n617 585
R259 B.n616 B.n57 585
R260 B.n615 B.n614 585
R261 B.n613 B.n58 585
R262 B.n612 B.n611 585
R263 B.n610 B.n59 585
R264 B.n609 B.n608 585
R265 B.n607 B.n60 585
R266 B.n606 B.n605 585
R267 B.n604 B.n61 585
R268 B.n603 B.n602 585
R269 B.n601 B.n62 585
R270 B.n600 B.n599 585
R271 B.n598 B.n63 585
R272 B.n597 B.n596 585
R273 B.n595 B.n64 585
R274 B.n594 B.n593 585
R275 B.n592 B.n65 585
R276 B.n591 B.n590 585
R277 B.n589 B.n66 585
R278 B.n588 B.n587 585
R279 B.n586 B.n67 585
R280 B.n585 B.n584 585
R281 B.n583 B.n68 585
R282 B.n582 B.n581 585
R283 B.n580 B.n69 585
R284 B.n579 B.n578 585
R285 B.n577 B.n70 585
R286 B.n576 B.n575 585
R287 B.n574 B.n71 585
R288 B.n573 B.n572 585
R289 B.n571 B.n72 585
R290 B.n570 B.n569 585
R291 B.n568 B.n73 585
R292 B.n567 B.n566 585
R293 B.n565 B.n74 585
R294 B.n564 B.n563 585
R295 B.n562 B.n75 585
R296 B.n561 B.n560 585
R297 B.n559 B.n76 585
R298 B.n558 B.n557 585
R299 B.n556 B.n77 585
R300 B.n555 B.n554 585
R301 B.n553 B.n78 585
R302 B.n552 B.n551 585
R303 B.n550 B.n79 585
R304 B.n549 B.n548 585
R305 B.n547 B.n80 585
R306 B.n546 B.n545 585
R307 B.n544 B.n81 585
R308 B.n543 B.n542 585
R309 B.n541 B.n82 585
R310 B.n540 B.n539 585
R311 B.n538 B.n83 585
R312 B.n722 B.n721 585
R313 B.n723 B.n18 585
R314 B.n725 B.n724 585
R315 B.n726 B.n17 585
R316 B.n728 B.n727 585
R317 B.n729 B.n16 585
R318 B.n731 B.n730 585
R319 B.n732 B.n15 585
R320 B.n734 B.n733 585
R321 B.n735 B.n14 585
R322 B.n737 B.n736 585
R323 B.n738 B.n13 585
R324 B.n740 B.n739 585
R325 B.n741 B.n12 585
R326 B.n743 B.n742 585
R327 B.n744 B.n11 585
R328 B.n746 B.n745 585
R329 B.n747 B.n10 585
R330 B.n749 B.n748 585
R331 B.n750 B.n9 585
R332 B.n752 B.n751 585
R333 B.n753 B.n8 585
R334 B.n755 B.n754 585
R335 B.n756 B.n7 585
R336 B.n758 B.n757 585
R337 B.n759 B.n6 585
R338 B.n761 B.n760 585
R339 B.n762 B.n5 585
R340 B.n764 B.n763 585
R341 B.n765 B.n4 585
R342 B.n767 B.n766 585
R343 B.n768 B.n3 585
R344 B.n770 B.n769 585
R345 B.n771 B.n0 585
R346 B.n2 B.n1 585
R347 B.n198 B.n197 585
R348 B.n200 B.n199 585
R349 B.n201 B.n196 585
R350 B.n203 B.n202 585
R351 B.n204 B.n195 585
R352 B.n206 B.n205 585
R353 B.n207 B.n194 585
R354 B.n209 B.n208 585
R355 B.n210 B.n193 585
R356 B.n212 B.n211 585
R357 B.n213 B.n192 585
R358 B.n215 B.n214 585
R359 B.n216 B.n191 585
R360 B.n218 B.n217 585
R361 B.n219 B.n190 585
R362 B.n221 B.n220 585
R363 B.n222 B.n189 585
R364 B.n224 B.n223 585
R365 B.n225 B.n188 585
R366 B.n227 B.n226 585
R367 B.n228 B.n187 585
R368 B.n230 B.n229 585
R369 B.n231 B.n186 585
R370 B.n233 B.n232 585
R371 B.n234 B.n185 585
R372 B.n236 B.n235 585
R373 B.n237 B.n184 585
R374 B.n239 B.n238 585
R375 B.n240 B.n183 585
R376 B.n242 B.n241 585
R377 B.n243 B.n182 585
R378 B.n245 B.n244 585
R379 B.n246 B.n181 585
R380 B.n248 B.n181 506.916
R381 B.n433 B.n432 506.916
R382 B.n536 B.n83 506.916
R383 B.n722 B.n19 506.916
R384 B.n344 B.t10 505.289
R385 B.n54 B.t5 505.289
R386 B.n152 B.t1 505.289
R387 B.n48 B.t8 505.289
R388 B.n345 B.t11 461.652
R389 B.n55 B.t4 461.652
R390 B.n153 B.t2 461.652
R391 B.n49 B.t7 461.652
R392 B.n152 B.t0 417.348
R393 B.n344 B.t9 417.348
R394 B.n54 B.t3 417.348
R395 B.n48 B.t6 417.348
R396 B.n773 B.n772 256.663
R397 B.n772 B.n771 235.042
R398 B.n772 B.n2 235.042
R399 B.n249 B.n248 163.367
R400 B.n250 B.n249 163.367
R401 B.n250 B.n179 163.367
R402 B.n254 B.n179 163.367
R403 B.n255 B.n254 163.367
R404 B.n256 B.n255 163.367
R405 B.n256 B.n177 163.367
R406 B.n260 B.n177 163.367
R407 B.n261 B.n260 163.367
R408 B.n262 B.n261 163.367
R409 B.n262 B.n175 163.367
R410 B.n266 B.n175 163.367
R411 B.n267 B.n266 163.367
R412 B.n268 B.n267 163.367
R413 B.n268 B.n173 163.367
R414 B.n272 B.n173 163.367
R415 B.n273 B.n272 163.367
R416 B.n274 B.n273 163.367
R417 B.n274 B.n171 163.367
R418 B.n278 B.n171 163.367
R419 B.n279 B.n278 163.367
R420 B.n280 B.n279 163.367
R421 B.n280 B.n169 163.367
R422 B.n284 B.n169 163.367
R423 B.n285 B.n284 163.367
R424 B.n286 B.n285 163.367
R425 B.n286 B.n167 163.367
R426 B.n290 B.n167 163.367
R427 B.n291 B.n290 163.367
R428 B.n292 B.n291 163.367
R429 B.n292 B.n165 163.367
R430 B.n296 B.n165 163.367
R431 B.n297 B.n296 163.367
R432 B.n298 B.n297 163.367
R433 B.n298 B.n163 163.367
R434 B.n302 B.n163 163.367
R435 B.n303 B.n302 163.367
R436 B.n304 B.n303 163.367
R437 B.n304 B.n161 163.367
R438 B.n308 B.n161 163.367
R439 B.n309 B.n308 163.367
R440 B.n310 B.n309 163.367
R441 B.n310 B.n159 163.367
R442 B.n314 B.n159 163.367
R443 B.n315 B.n314 163.367
R444 B.n316 B.n315 163.367
R445 B.n316 B.n157 163.367
R446 B.n320 B.n157 163.367
R447 B.n321 B.n320 163.367
R448 B.n322 B.n321 163.367
R449 B.n322 B.n155 163.367
R450 B.n326 B.n155 163.367
R451 B.n327 B.n326 163.367
R452 B.n328 B.n327 163.367
R453 B.n328 B.n151 163.367
R454 B.n333 B.n151 163.367
R455 B.n334 B.n333 163.367
R456 B.n335 B.n334 163.367
R457 B.n335 B.n149 163.367
R458 B.n339 B.n149 163.367
R459 B.n340 B.n339 163.367
R460 B.n341 B.n340 163.367
R461 B.n341 B.n147 163.367
R462 B.n348 B.n147 163.367
R463 B.n349 B.n348 163.367
R464 B.n350 B.n349 163.367
R465 B.n350 B.n145 163.367
R466 B.n354 B.n145 163.367
R467 B.n355 B.n354 163.367
R468 B.n356 B.n355 163.367
R469 B.n356 B.n143 163.367
R470 B.n360 B.n143 163.367
R471 B.n361 B.n360 163.367
R472 B.n362 B.n361 163.367
R473 B.n362 B.n141 163.367
R474 B.n366 B.n141 163.367
R475 B.n367 B.n366 163.367
R476 B.n368 B.n367 163.367
R477 B.n368 B.n139 163.367
R478 B.n372 B.n139 163.367
R479 B.n373 B.n372 163.367
R480 B.n374 B.n373 163.367
R481 B.n374 B.n137 163.367
R482 B.n378 B.n137 163.367
R483 B.n379 B.n378 163.367
R484 B.n380 B.n379 163.367
R485 B.n380 B.n135 163.367
R486 B.n384 B.n135 163.367
R487 B.n385 B.n384 163.367
R488 B.n386 B.n385 163.367
R489 B.n386 B.n133 163.367
R490 B.n390 B.n133 163.367
R491 B.n391 B.n390 163.367
R492 B.n392 B.n391 163.367
R493 B.n392 B.n131 163.367
R494 B.n396 B.n131 163.367
R495 B.n397 B.n396 163.367
R496 B.n398 B.n397 163.367
R497 B.n398 B.n129 163.367
R498 B.n402 B.n129 163.367
R499 B.n403 B.n402 163.367
R500 B.n404 B.n403 163.367
R501 B.n404 B.n127 163.367
R502 B.n408 B.n127 163.367
R503 B.n409 B.n408 163.367
R504 B.n410 B.n409 163.367
R505 B.n410 B.n125 163.367
R506 B.n414 B.n125 163.367
R507 B.n415 B.n414 163.367
R508 B.n416 B.n415 163.367
R509 B.n416 B.n123 163.367
R510 B.n420 B.n123 163.367
R511 B.n421 B.n420 163.367
R512 B.n422 B.n421 163.367
R513 B.n422 B.n121 163.367
R514 B.n426 B.n121 163.367
R515 B.n427 B.n426 163.367
R516 B.n428 B.n427 163.367
R517 B.n428 B.n119 163.367
R518 B.n432 B.n119 163.367
R519 B.n536 B.n535 163.367
R520 B.n535 B.n534 163.367
R521 B.n534 B.n85 163.367
R522 B.n530 B.n85 163.367
R523 B.n530 B.n529 163.367
R524 B.n529 B.n528 163.367
R525 B.n528 B.n87 163.367
R526 B.n524 B.n87 163.367
R527 B.n524 B.n523 163.367
R528 B.n523 B.n522 163.367
R529 B.n522 B.n89 163.367
R530 B.n518 B.n89 163.367
R531 B.n518 B.n517 163.367
R532 B.n517 B.n516 163.367
R533 B.n516 B.n91 163.367
R534 B.n512 B.n91 163.367
R535 B.n512 B.n511 163.367
R536 B.n511 B.n510 163.367
R537 B.n510 B.n93 163.367
R538 B.n506 B.n93 163.367
R539 B.n506 B.n505 163.367
R540 B.n505 B.n504 163.367
R541 B.n504 B.n95 163.367
R542 B.n500 B.n95 163.367
R543 B.n500 B.n499 163.367
R544 B.n499 B.n498 163.367
R545 B.n498 B.n97 163.367
R546 B.n494 B.n97 163.367
R547 B.n494 B.n493 163.367
R548 B.n493 B.n492 163.367
R549 B.n492 B.n99 163.367
R550 B.n488 B.n99 163.367
R551 B.n488 B.n487 163.367
R552 B.n487 B.n486 163.367
R553 B.n486 B.n101 163.367
R554 B.n482 B.n101 163.367
R555 B.n482 B.n481 163.367
R556 B.n481 B.n480 163.367
R557 B.n480 B.n103 163.367
R558 B.n476 B.n103 163.367
R559 B.n476 B.n475 163.367
R560 B.n475 B.n474 163.367
R561 B.n474 B.n105 163.367
R562 B.n470 B.n105 163.367
R563 B.n470 B.n469 163.367
R564 B.n469 B.n468 163.367
R565 B.n468 B.n107 163.367
R566 B.n464 B.n107 163.367
R567 B.n464 B.n463 163.367
R568 B.n463 B.n462 163.367
R569 B.n462 B.n109 163.367
R570 B.n458 B.n109 163.367
R571 B.n458 B.n457 163.367
R572 B.n457 B.n456 163.367
R573 B.n456 B.n111 163.367
R574 B.n452 B.n111 163.367
R575 B.n452 B.n451 163.367
R576 B.n451 B.n450 163.367
R577 B.n450 B.n113 163.367
R578 B.n446 B.n113 163.367
R579 B.n446 B.n445 163.367
R580 B.n445 B.n444 163.367
R581 B.n444 B.n115 163.367
R582 B.n440 B.n115 163.367
R583 B.n440 B.n439 163.367
R584 B.n439 B.n438 163.367
R585 B.n438 B.n117 163.367
R586 B.n434 B.n117 163.367
R587 B.n434 B.n433 163.367
R588 B.n718 B.n19 163.367
R589 B.n718 B.n717 163.367
R590 B.n717 B.n716 163.367
R591 B.n716 B.n21 163.367
R592 B.n712 B.n21 163.367
R593 B.n712 B.n711 163.367
R594 B.n711 B.n710 163.367
R595 B.n710 B.n23 163.367
R596 B.n706 B.n23 163.367
R597 B.n706 B.n705 163.367
R598 B.n705 B.n704 163.367
R599 B.n704 B.n25 163.367
R600 B.n700 B.n25 163.367
R601 B.n700 B.n699 163.367
R602 B.n699 B.n698 163.367
R603 B.n698 B.n27 163.367
R604 B.n694 B.n27 163.367
R605 B.n694 B.n693 163.367
R606 B.n693 B.n692 163.367
R607 B.n692 B.n29 163.367
R608 B.n688 B.n29 163.367
R609 B.n688 B.n687 163.367
R610 B.n687 B.n686 163.367
R611 B.n686 B.n31 163.367
R612 B.n682 B.n31 163.367
R613 B.n682 B.n681 163.367
R614 B.n681 B.n680 163.367
R615 B.n680 B.n33 163.367
R616 B.n676 B.n33 163.367
R617 B.n676 B.n675 163.367
R618 B.n675 B.n674 163.367
R619 B.n674 B.n35 163.367
R620 B.n670 B.n35 163.367
R621 B.n670 B.n669 163.367
R622 B.n669 B.n668 163.367
R623 B.n668 B.n37 163.367
R624 B.n664 B.n37 163.367
R625 B.n664 B.n663 163.367
R626 B.n663 B.n662 163.367
R627 B.n662 B.n39 163.367
R628 B.n658 B.n39 163.367
R629 B.n658 B.n657 163.367
R630 B.n657 B.n656 163.367
R631 B.n656 B.n41 163.367
R632 B.n652 B.n41 163.367
R633 B.n652 B.n651 163.367
R634 B.n651 B.n650 163.367
R635 B.n650 B.n43 163.367
R636 B.n646 B.n43 163.367
R637 B.n646 B.n645 163.367
R638 B.n645 B.n644 163.367
R639 B.n644 B.n45 163.367
R640 B.n640 B.n45 163.367
R641 B.n640 B.n639 163.367
R642 B.n639 B.n638 163.367
R643 B.n638 B.n47 163.367
R644 B.n633 B.n47 163.367
R645 B.n633 B.n632 163.367
R646 B.n632 B.n631 163.367
R647 B.n631 B.n51 163.367
R648 B.n627 B.n51 163.367
R649 B.n627 B.n626 163.367
R650 B.n626 B.n625 163.367
R651 B.n625 B.n53 163.367
R652 B.n620 B.n53 163.367
R653 B.n620 B.n619 163.367
R654 B.n619 B.n618 163.367
R655 B.n618 B.n57 163.367
R656 B.n614 B.n57 163.367
R657 B.n614 B.n613 163.367
R658 B.n613 B.n612 163.367
R659 B.n612 B.n59 163.367
R660 B.n608 B.n59 163.367
R661 B.n608 B.n607 163.367
R662 B.n607 B.n606 163.367
R663 B.n606 B.n61 163.367
R664 B.n602 B.n61 163.367
R665 B.n602 B.n601 163.367
R666 B.n601 B.n600 163.367
R667 B.n600 B.n63 163.367
R668 B.n596 B.n63 163.367
R669 B.n596 B.n595 163.367
R670 B.n595 B.n594 163.367
R671 B.n594 B.n65 163.367
R672 B.n590 B.n65 163.367
R673 B.n590 B.n589 163.367
R674 B.n589 B.n588 163.367
R675 B.n588 B.n67 163.367
R676 B.n584 B.n67 163.367
R677 B.n584 B.n583 163.367
R678 B.n583 B.n582 163.367
R679 B.n582 B.n69 163.367
R680 B.n578 B.n69 163.367
R681 B.n578 B.n577 163.367
R682 B.n577 B.n576 163.367
R683 B.n576 B.n71 163.367
R684 B.n572 B.n71 163.367
R685 B.n572 B.n571 163.367
R686 B.n571 B.n570 163.367
R687 B.n570 B.n73 163.367
R688 B.n566 B.n73 163.367
R689 B.n566 B.n565 163.367
R690 B.n565 B.n564 163.367
R691 B.n564 B.n75 163.367
R692 B.n560 B.n75 163.367
R693 B.n560 B.n559 163.367
R694 B.n559 B.n558 163.367
R695 B.n558 B.n77 163.367
R696 B.n554 B.n77 163.367
R697 B.n554 B.n553 163.367
R698 B.n553 B.n552 163.367
R699 B.n552 B.n79 163.367
R700 B.n548 B.n79 163.367
R701 B.n548 B.n547 163.367
R702 B.n547 B.n546 163.367
R703 B.n546 B.n81 163.367
R704 B.n542 B.n81 163.367
R705 B.n542 B.n541 163.367
R706 B.n541 B.n540 163.367
R707 B.n540 B.n83 163.367
R708 B.n723 B.n722 163.367
R709 B.n724 B.n723 163.367
R710 B.n724 B.n17 163.367
R711 B.n728 B.n17 163.367
R712 B.n729 B.n728 163.367
R713 B.n730 B.n729 163.367
R714 B.n730 B.n15 163.367
R715 B.n734 B.n15 163.367
R716 B.n735 B.n734 163.367
R717 B.n736 B.n735 163.367
R718 B.n736 B.n13 163.367
R719 B.n740 B.n13 163.367
R720 B.n741 B.n740 163.367
R721 B.n742 B.n741 163.367
R722 B.n742 B.n11 163.367
R723 B.n746 B.n11 163.367
R724 B.n747 B.n746 163.367
R725 B.n748 B.n747 163.367
R726 B.n748 B.n9 163.367
R727 B.n752 B.n9 163.367
R728 B.n753 B.n752 163.367
R729 B.n754 B.n753 163.367
R730 B.n754 B.n7 163.367
R731 B.n758 B.n7 163.367
R732 B.n759 B.n758 163.367
R733 B.n760 B.n759 163.367
R734 B.n760 B.n5 163.367
R735 B.n764 B.n5 163.367
R736 B.n765 B.n764 163.367
R737 B.n766 B.n765 163.367
R738 B.n766 B.n3 163.367
R739 B.n770 B.n3 163.367
R740 B.n771 B.n770 163.367
R741 B.n197 B.n2 163.367
R742 B.n200 B.n197 163.367
R743 B.n201 B.n200 163.367
R744 B.n202 B.n201 163.367
R745 B.n202 B.n195 163.367
R746 B.n206 B.n195 163.367
R747 B.n207 B.n206 163.367
R748 B.n208 B.n207 163.367
R749 B.n208 B.n193 163.367
R750 B.n212 B.n193 163.367
R751 B.n213 B.n212 163.367
R752 B.n214 B.n213 163.367
R753 B.n214 B.n191 163.367
R754 B.n218 B.n191 163.367
R755 B.n219 B.n218 163.367
R756 B.n220 B.n219 163.367
R757 B.n220 B.n189 163.367
R758 B.n224 B.n189 163.367
R759 B.n225 B.n224 163.367
R760 B.n226 B.n225 163.367
R761 B.n226 B.n187 163.367
R762 B.n230 B.n187 163.367
R763 B.n231 B.n230 163.367
R764 B.n232 B.n231 163.367
R765 B.n232 B.n185 163.367
R766 B.n236 B.n185 163.367
R767 B.n237 B.n236 163.367
R768 B.n238 B.n237 163.367
R769 B.n238 B.n183 163.367
R770 B.n242 B.n183 163.367
R771 B.n243 B.n242 163.367
R772 B.n244 B.n243 163.367
R773 B.n244 B.n181 163.367
R774 B.n331 B.n153 59.5399
R775 B.n346 B.n345 59.5399
R776 B.n622 B.n55 59.5399
R777 B.n636 B.n49 59.5399
R778 B.n153 B.n152 43.6369
R779 B.n345 B.n344 43.6369
R780 B.n55 B.n54 43.6369
R781 B.n49 B.n48 43.6369
R782 B.n721 B.n720 32.9371
R783 B.n538 B.n537 32.9371
R784 B.n431 B.n118 32.9371
R785 B.n247 B.n246 32.9371
R786 B B.n773 18.0485
R787 B.n721 B.n18 10.6151
R788 B.n725 B.n18 10.6151
R789 B.n726 B.n725 10.6151
R790 B.n727 B.n726 10.6151
R791 B.n727 B.n16 10.6151
R792 B.n731 B.n16 10.6151
R793 B.n732 B.n731 10.6151
R794 B.n733 B.n732 10.6151
R795 B.n733 B.n14 10.6151
R796 B.n737 B.n14 10.6151
R797 B.n738 B.n737 10.6151
R798 B.n739 B.n738 10.6151
R799 B.n739 B.n12 10.6151
R800 B.n743 B.n12 10.6151
R801 B.n744 B.n743 10.6151
R802 B.n745 B.n744 10.6151
R803 B.n745 B.n10 10.6151
R804 B.n749 B.n10 10.6151
R805 B.n750 B.n749 10.6151
R806 B.n751 B.n750 10.6151
R807 B.n751 B.n8 10.6151
R808 B.n755 B.n8 10.6151
R809 B.n756 B.n755 10.6151
R810 B.n757 B.n756 10.6151
R811 B.n757 B.n6 10.6151
R812 B.n761 B.n6 10.6151
R813 B.n762 B.n761 10.6151
R814 B.n763 B.n762 10.6151
R815 B.n763 B.n4 10.6151
R816 B.n767 B.n4 10.6151
R817 B.n768 B.n767 10.6151
R818 B.n769 B.n768 10.6151
R819 B.n769 B.n0 10.6151
R820 B.n720 B.n719 10.6151
R821 B.n719 B.n20 10.6151
R822 B.n715 B.n20 10.6151
R823 B.n715 B.n714 10.6151
R824 B.n714 B.n713 10.6151
R825 B.n713 B.n22 10.6151
R826 B.n709 B.n22 10.6151
R827 B.n709 B.n708 10.6151
R828 B.n708 B.n707 10.6151
R829 B.n707 B.n24 10.6151
R830 B.n703 B.n24 10.6151
R831 B.n703 B.n702 10.6151
R832 B.n702 B.n701 10.6151
R833 B.n701 B.n26 10.6151
R834 B.n697 B.n26 10.6151
R835 B.n697 B.n696 10.6151
R836 B.n696 B.n695 10.6151
R837 B.n695 B.n28 10.6151
R838 B.n691 B.n28 10.6151
R839 B.n691 B.n690 10.6151
R840 B.n690 B.n689 10.6151
R841 B.n689 B.n30 10.6151
R842 B.n685 B.n30 10.6151
R843 B.n685 B.n684 10.6151
R844 B.n684 B.n683 10.6151
R845 B.n683 B.n32 10.6151
R846 B.n679 B.n32 10.6151
R847 B.n679 B.n678 10.6151
R848 B.n678 B.n677 10.6151
R849 B.n677 B.n34 10.6151
R850 B.n673 B.n34 10.6151
R851 B.n673 B.n672 10.6151
R852 B.n672 B.n671 10.6151
R853 B.n671 B.n36 10.6151
R854 B.n667 B.n36 10.6151
R855 B.n667 B.n666 10.6151
R856 B.n666 B.n665 10.6151
R857 B.n665 B.n38 10.6151
R858 B.n661 B.n38 10.6151
R859 B.n661 B.n660 10.6151
R860 B.n660 B.n659 10.6151
R861 B.n659 B.n40 10.6151
R862 B.n655 B.n40 10.6151
R863 B.n655 B.n654 10.6151
R864 B.n654 B.n653 10.6151
R865 B.n653 B.n42 10.6151
R866 B.n649 B.n42 10.6151
R867 B.n649 B.n648 10.6151
R868 B.n648 B.n647 10.6151
R869 B.n647 B.n44 10.6151
R870 B.n643 B.n44 10.6151
R871 B.n643 B.n642 10.6151
R872 B.n642 B.n641 10.6151
R873 B.n641 B.n46 10.6151
R874 B.n637 B.n46 10.6151
R875 B.n635 B.n634 10.6151
R876 B.n634 B.n50 10.6151
R877 B.n630 B.n50 10.6151
R878 B.n630 B.n629 10.6151
R879 B.n629 B.n628 10.6151
R880 B.n628 B.n52 10.6151
R881 B.n624 B.n52 10.6151
R882 B.n624 B.n623 10.6151
R883 B.n621 B.n56 10.6151
R884 B.n617 B.n56 10.6151
R885 B.n617 B.n616 10.6151
R886 B.n616 B.n615 10.6151
R887 B.n615 B.n58 10.6151
R888 B.n611 B.n58 10.6151
R889 B.n611 B.n610 10.6151
R890 B.n610 B.n609 10.6151
R891 B.n609 B.n60 10.6151
R892 B.n605 B.n60 10.6151
R893 B.n605 B.n604 10.6151
R894 B.n604 B.n603 10.6151
R895 B.n603 B.n62 10.6151
R896 B.n599 B.n62 10.6151
R897 B.n599 B.n598 10.6151
R898 B.n598 B.n597 10.6151
R899 B.n597 B.n64 10.6151
R900 B.n593 B.n64 10.6151
R901 B.n593 B.n592 10.6151
R902 B.n592 B.n591 10.6151
R903 B.n591 B.n66 10.6151
R904 B.n587 B.n66 10.6151
R905 B.n587 B.n586 10.6151
R906 B.n586 B.n585 10.6151
R907 B.n585 B.n68 10.6151
R908 B.n581 B.n68 10.6151
R909 B.n581 B.n580 10.6151
R910 B.n580 B.n579 10.6151
R911 B.n579 B.n70 10.6151
R912 B.n575 B.n70 10.6151
R913 B.n575 B.n574 10.6151
R914 B.n574 B.n573 10.6151
R915 B.n573 B.n72 10.6151
R916 B.n569 B.n72 10.6151
R917 B.n569 B.n568 10.6151
R918 B.n568 B.n567 10.6151
R919 B.n567 B.n74 10.6151
R920 B.n563 B.n74 10.6151
R921 B.n563 B.n562 10.6151
R922 B.n562 B.n561 10.6151
R923 B.n561 B.n76 10.6151
R924 B.n557 B.n76 10.6151
R925 B.n557 B.n556 10.6151
R926 B.n556 B.n555 10.6151
R927 B.n555 B.n78 10.6151
R928 B.n551 B.n78 10.6151
R929 B.n551 B.n550 10.6151
R930 B.n550 B.n549 10.6151
R931 B.n549 B.n80 10.6151
R932 B.n545 B.n80 10.6151
R933 B.n545 B.n544 10.6151
R934 B.n544 B.n543 10.6151
R935 B.n543 B.n82 10.6151
R936 B.n539 B.n82 10.6151
R937 B.n539 B.n538 10.6151
R938 B.n537 B.n84 10.6151
R939 B.n533 B.n84 10.6151
R940 B.n533 B.n532 10.6151
R941 B.n532 B.n531 10.6151
R942 B.n531 B.n86 10.6151
R943 B.n527 B.n86 10.6151
R944 B.n527 B.n526 10.6151
R945 B.n526 B.n525 10.6151
R946 B.n525 B.n88 10.6151
R947 B.n521 B.n88 10.6151
R948 B.n521 B.n520 10.6151
R949 B.n520 B.n519 10.6151
R950 B.n519 B.n90 10.6151
R951 B.n515 B.n90 10.6151
R952 B.n515 B.n514 10.6151
R953 B.n514 B.n513 10.6151
R954 B.n513 B.n92 10.6151
R955 B.n509 B.n92 10.6151
R956 B.n509 B.n508 10.6151
R957 B.n508 B.n507 10.6151
R958 B.n507 B.n94 10.6151
R959 B.n503 B.n94 10.6151
R960 B.n503 B.n502 10.6151
R961 B.n502 B.n501 10.6151
R962 B.n501 B.n96 10.6151
R963 B.n497 B.n96 10.6151
R964 B.n497 B.n496 10.6151
R965 B.n496 B.n495 10.6151
R966 B.n495 B.n98 10.6151
R967 B.n491 B.n98 10.6151
R968 B.n491 B.n490 10.6151
R969 B.n490 B.n489 10.6151
R970 B.n489 B.n100 10.6151
R971 B.n485 B.n100 10.6151
R972 B.n485 B.n484 10.6151
R973 B.n484 B.n483 10.6151
R974 B.n483 B.n102 10.6151
R975 B.n479 B.n102 10.6151
R976 B.n479 B.n478 10.6151
R977 B.n478 B.n477 10.6151
R978 B.n477 B.n104 10.6151
R979 B.n473 B.n104 10.6151
R980 B.n473 B.n472 10.6151
R981 B.n472 B.n471 10.6151
R982 B.n471 B.n106 10.6151
R983 B.n467 B.n106 10.6151
R984 B.n467 B.n466 10.6151
R985 B.n466 B.n465 10.6151
R986 B.n465 B.n108 10.6151
R987 B.n461 B.n108 10.6151
R988 B.n461 B.n460 10.6151
R989 B.n460 B.n459 10.6151
R990 B.n459 B.n110 10.6151
R991 B.n455 B.n110 10.6151
R992 B.n455 B.n454 10.6151
R993 B.n454 B.n453 10.6151
R994 B.n453 B.n112 10.6151
R995 B.n449 B.n112 10.6151
R996 B.n449 B.n448 10.6151
R997 B.n448 B.n447 10.6151
R998 B.n447 B.n114 10.6151
R999 B.n443 B.n114 10.6151
R1000 B.n443 B.n442 10.6151
R1001 B.n442 B.n441 10.6151
R1002 B.n441 B.n116 10.6151
R1003 B.n437 B.n116 10.6151
R1004 B.n437 B.n436 10.6151
R1005 B.n436 B.n435 10.6151
R1006 B.n435 B.n118 10.6151
R1007 B.n198 B.n1 10.6151
R1008 B.n199 B.n198 10.6151
R1009 B.n199 B.n196 10.6151
R1010 B.n203 B.n196 10.6151
R1011 B.n204 B.n203 10.6151
R1012 B.n205 B.n204 10.6151
R1013 B.n205 B.n194 10.6151
R1014 B.n209 B.n194 10.6151
R1015 B.n210 B.n209 10.6151
R1016 B.n211 B.n210 10.6151
R1017 B.n211 B.n192 10.6151
R1018 B.n215 B.n192 10.6151
R1019 B.n216 B.n215 10.6151
R1020 B.n217 B.n216 10.6151
R1021 B.n217 B.n190 10.6151
R1022 B.n221 B.n190 10.6151
R1023 B.n222 B.n221 10.6151
R1024 B.n223 B.n222 10.6151
R1025 B.n223 B.n188 10.6151
R1026 B.n227 B.n188 10.6151
R1027 B.n228 B.n227 10.6151
R1028 B.n229 B.n228 10.6151
R1029 B.n229 B.n186 10.6151
R1030 B.n233 B.n186 10.6151
R1031 B.n234 B.n233 10.6151
R1032 B.n235 B.n234 10.6151
R1033 B.n235 B.n184 10.6151
R1034 B.n239 B.n184 10.6151
R1035 B.n240 B.n239 10.6151
R1036 B.n241 B.n240 10.6151
R1037 B.n241 B.n182 10.6151
R1038 B.n245 B.n182 10.6151
R1039 B.n246 B.n245 10.6151
R1040 B.n247 B.n180 10.6151
R1041 B.n251 B.n180 10.6151
R1042 B.n252 B.n251 10.6151
R1043 B.n253 B.n252 10.6151
R1044 B.n253 B.n178 10.6151
R1045 B.n257 B.n178 10.6151
R1046 B.n258 B.n257 10.6151
R1047 B.n259 B.n258 10.6151
R1048 B.n259 B.n176 10.6151
R1049 B.n263 B.n176 10.6151
R1050 B.n264 B.n263 10.6151
R1051 B.n265 B.n264 10.6151
R1052 B.n265 B.n174 10.6151
R1053 B.n269 B.n174 10.6151
R1054 B.n270 B.n269 10.6151
R1055 B.n271 B.n270 10.6151
R1056 B.n271 B.n172 10.6151
R1057 B.n275 B.n172 10.6151
R1058 B.n276 B.n275 10.6151
R1059 B.n277 B.n276 10.6151
R1060 B.n277 B.n170 10.6151
R1061 B.n281 B.n170 10.6151
R1062 B.n282 B.n281 10.6151
R1063 B.n283 B.n282 10.6151
R1064 B.n283 B.n168 10.6151
R1065 B.n287 B.n168 10.6151
R1066 B.n288 B.n287 10.6151
R1067 B.n289 B.n288 10.6151
R1068 B.n289 B.n166 10.6151
R1069 B.n293 B.n166 10.6151
R1070 B.n294 B.n293 10.6151
R1071 B.n295 B.n294 10.6151
R1072 B.n295 B.n164 10.6151
R1073 B.n299 B.n164 10.6151
R1074 B.n300 B.n299 10.6151
R1075 B.n301 B.n300 10.6151
R1076 B.n301 B.n162 10.6151
R1077 B.n305 B.n162 10.6151
R1078 B.n306 B.n305 10.6151
R1079 B.n307 B.n306 10.6151
R1080 B.n307 B.n160 10.6151
R1081 B.n311 B.n160 10.6151
R1082 B.n312 B.n311 10.6151
R1083 B.n313 B.n312 10.6151
R1084 B.n313 B.n158 10.6151
R1085 B.n317 B.n158 10.6151
R1086 B.n318 B.n317 10.6151
R1087 B.n319 B.n318 10.6151
R1088 B.n319 B.n156 10.6151
R1089 B.n323 B.n156 10.6151
R1090 B.n324 B.n323 10.6151
R1091 B.n325 B.n324 10.6151
R1092 B.n325 B.n154 10.6151
R1093 B.n329 B.n154 10.6151
R1094 B.n330 B.n329 10.6151
R1095 B.n332 B.n150 10.6151
R1096 B.n336 B.n150 10.6151
R1097 B.n337 B.n336 10.6151
R1098 B.n338 B.n337 10.6151
R1099 B.n338 B.n148 10.6151
R1100 B.n342 B.n148 10.6151
R1101 B.n343 B.n342 10.6151
R1102 B.n347 B.n343 10.6151
R1103 B.n351 B.n146 10.6151
R1104 B.n352 B.n351 10.6151
R1105 B.n353 B.n352 10.6151
R1106 B.n353 B.n144 10.6151
R1107 B.n357 B.n144 10.6151
R1108 B.n358 B.n357 10.6151
R1109 B.n359 B.n358 10.6151
R1110 B.n359 B.n142 10.6151
R1111 B.n363 B.n142 10.6151
R1112 B.n364 B.n363 10.6151
R1113 B.n365 B.n364 10.6151
R1114 B.n365 B.n140 10.6151
R1115 B.n369 B.n140 10.6151
R1116 B.n370 B.n369 10.6151
R1117 B.n371 B.n370 10.6151
R1118 B.n371 B.n138 10.6151
R1119 B.n375 B.n138 10.6151
R1120 B.n376 B.n375 10.6151
R1121 B.n377 B.n376 10.6151
R1122 B.n377 B.n136 10.6151
R1123 B.n381 B.n136 10.6151
R1124 B.n382 B.n381 10.6151
R1125 B.n383 B.n382 10.6151
R1126 B.n383 B.n134 10.6151
R1127 B.n387 B.n134 10.6151
R1128 B.n388 B.n387 10.6151
R1129 B.n389 B.n388 10.6151
R1130 B.n389 B.n132 10.6151
R1131 B.n393 B.n132 10.6151
R1132 B.n394 B.n393 10.6151
R1133 B.n395 B.n394 10.6151
R1134 B.n395 B.n130 10.6151
R1135 B.n399 B.n130 10.6151
R1136 B.n400 B.n399 10.6151
R1137 B.n401 B.n400 10.6151
R1138 B.n401 B.n128 10.6151
R1139 B.n405 B.n128 10.6151
R1140 B.n406 B.n405 10.6151
R1141 B.n407 B.n406 10.6151
R1142 B.n407 B.n126 10.6151
R1143 B.n411 B.n126 10.6151
R1144 B.n412 B.n411 10.6151
R1145 B.n413 B.n412 10.6151
R1146 B.n413 B.n124 10.6151
R1147 B.n417 B.n124 10.6151
R1148 B.n418 B.n417 10.6151
R1149 B.n419 B.n418 10.6151
R1150 B.n419 B.n122 10.6151
R1151 B.n423 B.n122 10.6151
R1152 B.n424 B.n423 10.6151
R1153 B.n425 B.n424 10.6151
R1154 B.n425 B.n120 10.6151
R1155 B.n429 B.n120 10.6151
R1156 B.n430 B.n429 10.6151
R1157 B.n431 B.n430 10.6151
R1158 B.n773 B.n0 8.11757
R1159 B.n773 B.n1 8.11757
R1160 B.n636 B.n635 6.5566
R1161 B.n623 B.n622 6.5566
R1162 B.n332 B.n331 6.5566
R1163 B.n347 B.n346 6.5566
R1164 B.n637 B.n636 4.05904
R1165 B.n622 B.n621 4.05904
R1166 B.n331 B.n330 4.05904
R1167 B.n346 B.n146 4.05904
R1168 VN.n2 VN.t2 241.974
R1169 VN.n14 VN.t1 241.974
R1170 VN.n10 VN.t4 210.625
R1171 VN.n3 VN.t0 210.625
R1172 VN.n22 VN.t3 210.625
R1173 VN.n15 VN.t5 210.625
R1174 VN.n21 VN.n12 161.3
R1175 VN.n20 VN.n19 161.3
R1176 VN.n18 VN.n13 161.3
R1177 VN.n17 VN.n16 161.3
R1178 VN.n9 VN.n0 161.3
R1179 VN.n8 VN.n7 161.3
R1180 VN.n6 VN.n1 161.3
R1181 VN.n5 VN.n4 161.3
R1182 VN.n11 VN.n10 86.2628
R1183 VN.n23 VN.n22 86.2628
R1184 VN.n3 VN.n2 57.7705
R1185 VN.n15 VN.n14 57.7705
R1186 VN.n8 VN.n1 52.5823
R1187 VN.n20 VN.n13 52.5823
R1188 VN VN.n23 49.9868
R1189 VN.n9 VN.n8 28.2389
R1190 VN.n21 VN.n20 28.2389
R1191 VN.n4 VN.n1 24.3439
R1192 VN.n10 VN.n9 24.3439
R1193 VN.n16 VN.n13 24.3439
R1194 VN.n22 VN.n21 24.3439
R1195 VN.n17 VN.n14 12.6525
R1196 VN.n5 VN.n2 12.6525
R1197 VN.n4 VN.n3 12.1722
R1198 VN.n16 VN.n15 12.1722
R1199 VN.n23 VN.n12 0.278398
R1200 VN.n11 VN.n0 0.278398
R1201 VN.n19 VN.n12 0.189894
R1202 VN.n19 VN.n18 0.189894
R1203 VN.n18 VN.n17 0.189894
R1204 VN.n6 VN.n5 0.189894
R1205 VN.n7 VN.n6 0.189894
R1206 VN.n7 VN.n0 0.189894
R1207 VN VN.n11 0.153422
R1208 VDD2.n183 VDD2.n95 756.745
R1209 VDD2.n88 VDD2.n0 756.745
R1210 VDD2.n184 VDD2.n183 585
R1211 VDD2.n182 VDD2.n181 585
R1212 VDD2.n99 VDD2.n98 585
R1213 VDD2.n176 VDD2.n175 585
R1214 VDD2.n174 VDD2.n173 585
R1215 VDD2.n172 VDD2.n102 585
R1216 VDD2.n106 VDD2.n103 585
R1217 VDD2.n167 VDD2.n166 585
R1218 VDD2.n165 VDD2.n164 585
R1219 VDD2.n108 VDD2.n107 585
R1220 VDD2.n159 VDD2.n158 585
R1221 VDD2.n157 VDD2.n156 585
R1222 VDD2.n112 VDD2.n111 585
R1223 VDD2.n151 VDD2.n150 585
R1224 VDD2.n149 VDD2.n148 585
R1225 VDD2.n116 VDD2.n115 585
R1226 VDD2.n143 VDD2.n142 585
R1227 VDD2.n141 VDD2.n140 585
R1228 VDD2.n120 VDD2.n119 585
R1229 VDD2.n135 VDD2.n134 585
R1230 VDD2.n133 VDD2.n132 585
R1231 VDD2.n124 VDD2.n123 585
R1232 VDD2.n127 VDD2.n126 585
R1233 VDD2.n31 VDD2.n30 585
R1234 VDD2.n28 VDD2.n27 585
R1235 VDD2.n37 VDD2.n36 585
R1236 VDD2.n39 VDD2.n38 585
R1237 VDD2.n24 VDD2.n23 585
R1238 VDD2.n45 VDD2.n44 585
R1239 VDD2.n47 VDD2.n46 585
R1240 VDD2.n20 VDD2.n19 585
R1241 VDD2.n53 VDD2.n52 585
R1242 VDD2.n55 VDD2.n54 585
R1243 VDD2.n16 VDD2.n15 585
R1244 VDD2.n61 VDD2.n60 585
R1245 VDD2.n63 VDD2.n62 585
R1246 VDD2.n12 VDD2.n11 585
R1247 VDD2.n69 VDD2.n68 585
R1248 VDD2.n72 VDD2.n71 585
R1249 VDD2.n70 VDD2.n8 585
R1250 VDD2.n77 VDD2.n7 585
R1251 VDD2.n79 VDD2.n78 585
R1252 VDD2.n81 VDD2.n80 585
R1253 VDD2.n4 VDD2.n3 585
R1254 VDD2.n87 VDD2.n86 585
R1255 VDD2.n89 VDD2.n88 585
R1256 VDD2.t5 VDD2.n125 327.466
R1257 VDD2.t0 VDD2.n29 327.466
R1258 VDD2.n183 VDD2.n182 171.744
R1259 VDD2.n182 VDD2.n98 171.744
R1260 VDD2.n175 VDD2.n98 171.744
R1261 VDD2.n175 VDD2.n174 171.744
R1262 VDD2.n174 VDD2.n102 171.744
R1263 VDD2.n106 VDD2.n102 171.744
R1264 VDD2.n166 VDD2.n106 171.744
R1265 VDD2.n166 VDD2.n165 171.744
R1266 VDD2.n165 VDD2.n107 171.744
R1267 VDD2.n158 VDD2.n107 171.744
R1268 VDD2.n158 VDD2.n157 171.744
R1269 VDD2.n157 VDD2.n111 171.744
R1270 VDD2.n150 VDD2.n111 171.744
R1271 VDD2.n150 VDD2.n149 171.744
R1272 VDD2.n149 VDD2.n115 171.744
R1273 VDD2.n142 VDD2.n115 171.744
R1274 VDD2.n142 VDD2.n141 171.744
R1275 VDD2.n141 VDD2.n119 171.744
R1276 VDD2.n134 VDD2.n119 171.744
R1277 VDD2.n134 VDD2.n133 171.744
R1278 VDD2.n133 VDD2.n123 171.744
R1279 VDD2.n126 VDD2.n123 171.744
R1280 VDD2.n30 VDD2.n27 171.744
R1281 VDD2.n37 VDD2.n27 171.744
R1282 VDD2.n38 VDD2.n37 171.744
R1283 VDD2.n38 VDD2.n23 171.744
R1284 VDD2.n45 VDD2.n23 171.744
R1285 VDD2.n46 VDD2.n45 171.744
R1286 VDD2.n46 VDD2.n19 171.744
R1287 VDD2.n53 VDD2.n19 171.744
R1288 VDD2.n54 VDD2.n53 171.744
R1289 VDD2.n54 VDD2.n15 171.744
R1290 VDD2.n61 VDD2.n15 171.744
R1291 VDD2.n62 VDD2.n61 171.744
R1292 VDD2.n62 VDD2.n11 171.744
R1293 VDD2.n69 VDD2.n11 171.744
R1294 VDD2.n71 VDD2.n69 171.744
R1295 VDD2.n71 VDD2.n70 171.744
R1296 VDD2.n70 VDD2.n7 171.744
R1297 VDD2.n79 VDD2.n7 171.744
R1298 VDD2.n80 VDD2.n79 171.744
R1299 VDD2.n80 VDD2.n3 171.744
R1300 VDD2.n87 VDD2.n3 171.744
R1301 VDD2.n88 VDD2.n87 171.744
R1302 VDD2.n126 VDD2.t5 85.8723
R1303 VDD2.n30 VDD2.t0 85.8723
R1304 VDD2.n94 VDD2.n93 69.4335
R1305 VDD2 VDD2.n189 69.4307
R1306 VDD2.n94 VDD2.n92 49.8757
R1307 VDD2.n188 VDD2.n187 48.4763
R1308 VDD2.n188 VDD2.n94 44.4847
R1309 VDD2.n127 VDD2.n125 16.3895
R1310 VDD2.n31 VDD2.n29 16.3895
R1311 VDD2.n173 VDD2.n172 13.1884
R1312 VDD2.n78 VDD2.n77 13.1884
R1313 VDD2.n176 VDD2.n101 12.8005
R1314 VDD2.n171 VDD2.n103 12.8005
R1315 VDD2.n128 VDD2.n124 12.8005
R1316 VDD2.n32 VDD2.n28 12.8005
R1317 VDD2.n76 VDD2.n8 12.8005
R1318 VDD2.n81 VDD2.n6 12.8005
R1319 VDD2.n177 VDD2.n99 12.0247
R1320 VDD2.n168 VDD2.n167 12.0247
R1321 VDD2.n132 VDD2.n131 12.0247
R1322 VDD2.n36 VDD2.n35 12.0247
R1323 VDD2.n73 VDD2.n72 12.0247
R1324 VDD2.n82 VDD2.n4 12.0247
R1325 VDD2.n181 VDD2.n180 11.249
R1326 VDD2.n164 VDD2.n105 11.249
R1327 VDD2.n135 VDD2.n122 11.249
R1328 VDD2.n39 VDD2.n26 11.249
R1329 VDD2.n68 VDD2.n10 11.249
R1330 VDD2.n86 VDD2.n85 11.249
R1331 VDD2.n184 VDD2.n97 10.4732
R1332 VDD2.n163 VDD2.n108 10.4732
R1333 VDD2.n136 VDD2.n120 10.4732
R1334 VDD2.n40 VDD2.n24 10.4732
R1335 VDD2.n67 VDD2.n12 10.4732
R1336 VDD2.n89 VDD2.n2 10.4732
R1337 VDD2.n185 VDD2.n95 9.69747
R1338 VDD2.n160 VDD2.n159 9.69747
R1339 VDD2.n140 VDD2.n139 9.69747
R1340 VDD2.n44 VDD2.n43 9.69747
R1341 VDD2.n64 VDD2.n63 9.69747
R1342 VDD2.n90 VDD2.n0 9.69747
R1343 VDD2.n187 VDD2.n186 9.45567
R1344 VDD2.n92 VDD2.n91 9.45567
R1345 VDD2.n153 VDD2.n152 9.3005
R1346 VDD2.n155 VDD2.n154 9.3005
R1347 VDD2.n110 VDD2.n109 9.3005
R1348 VDD2.n161 VDD2.n160 9.3005
R1349 VDD2.n163 VDD2.n162 9.3005
R1350 VDD2.n105 VDD2.n104 9.3005
R1351 VDD2.n169 VDD2.n168 9.3005
R1352 VDD2.n171 VDD2.n170 9.3005
R1353 VDD2.n186 VDD2.n185 9.3005
R1354 VDD2.n97 VDD2.n96 9.3005
R1355 VDD2.n180 VDD2.n179 9.3005
R1356 VDD2.n178 VDD2.n177 9.3005
R1357 VDD2.n101 VDD2.n100 9.3005
R1358 VDD2.n114 VDD2.n113 9.3005
R1359 VDD2.n147 VDD2.n146 9.3005
R1360 VDD2.n145 VDD2.n144 9.3005
R1361 VDD2.n118 VDD2.n117 9.3005
R1362 VDD2.n139 VDD2.n138 9.3005
R1363 VDD2.n137 VDD2.n136 9.3005
R1364 VDD2.n122 VDD2.n121 9.3005
R1365 VDD2.n131 VDD2.n130 9.3005
R1366 VDD2.n129 VDD2.n128 9.3005
R1367 VDD2.n91 VDD2.n90 9.3005
R1368 VDD2.n2 VDD2.n1 9.3005
R1369 VDD2.n85 VDD2.n84 9.3005
R1370 VDD2.n83 VDD2.n82 9.3005
R1371 VDD2.n6 VDD2.n5 9.3005
R1372 VDD2.n51 VDD2.n50 9.3005
R1373 VDD2.n49 VDD2.n48 9.3005
R1374 VDD2.n22 VDD2.n21 9.3005
R1375 VDD2.n43 VDD2.n42 9.3005
R1376 VDD2.n41 VDD2.n40 9.3005
R1377 VDD2.n26 VDD2.n25 9.3005
R1378 VDD2.n35 VDD2.n34 9.3005
R1379 VDD2.n33 VDD2.n32 9.3005
R1380 VDD2.n18 VDD2.n17 9.3005
R1381 VDD2.n57 VDD2.n56 9.3005
R1382 VDD2.n59 VDD2.n58 9.3005
R1383 VDD2.n14 VDD2.n13 9.3005
R1384 VDD2.n65 VDD2.n64 9.3005
R1385 VDD2.n67 VDD2.n66 9.3005
R1386 VDD2.n10 VDD2.n9 9.3005
R1387 VDD2.n74 VDD2.n73 9.3005
R1388 VDD2.n76 VDD2.n75 9.3005
R1389 VDD2.n156 VDD2.n110 8.92171
R1390 VDD2.n143 VDD2.n118 8.92171
R1391 VDD2.n47 VDD2.n22 8.92171
R1392 VDD2.n60 VDD2.n14 8.92171
R1393 VDD2.n155 VDD2.n112 8.14595
R1394 VDD2.n144 VDD2.n116 8.14595
R1395 VDD2.n48 VDD2.n20 8.14595
R1396 VDD2.n59 VDD2.n16 8.14595
R1397 VDD2.n152 VDD2.n151 7.3702
R1398 VDD2.n148 VDD2.n147 7.3702
R1399 VDD2.n52 VDD2.n51 7.3702
R1400 VDD2.n56 VDD2.n55 7.3702
R1401 VDD2.n151 VDD2.n114 6.59444
R1402 VDD2.n148 VDD2.n114 6.59444
R1403 VDD2.n52 VDD2.n18 6.59444
R1404 VDD2.n55 VDD2.n18 6.59444
R1405 VDD2.n152 VDD2.n112 5.81868
R1406 VDD2.n147 VDD2.n116 5.81868
R1407 VDD2.n51 VDD2.n20 5.81868
R1408 VDD2.n56 VDD2.n16 5.81868
R1409 VDD2.n156 VDD2.n155 5.04292
R1410 VDD2.n144 VDD2.n143 5.04292
R1411 VDD2.n48 VDD2.n47 5.04292
R1412 VDD2.n60 VDD2.n59 5.04292
R1413 VDD2.n187 VDD2.n95 4.26717
R1414 VDD2.n159 VDD2.n110 4.26717
R1415 VDD2.n140 VDD2.n118 4.26717
R1416 VDD2.n44 VDD2.n22 4.26717
R1417 VDD2.n63 VDD2.n14 4.26717
R1418 VDD2.n92 VDD2.n0 4.26717
R1419 VDD2.n129 VDD2.n125 3.70982
R1420 VDD2.n33 VDD2.n29 3.70982
R1421 VDD2.n185 VDD2.n184 3.49141
R1422 VDD2.n160 VDD2.n108 3.49141
R1423 VDD2.n139 VDD2.n120 3.49141
R1424 VDD2.n43 VDD2.n24 3.49141
R1425 VDD2.n64 VDD2.n12 3.49141
R1426 VDD2.n90 VDD2.n89 3.49141
R1427 VDD2.n181 VDD2.n97 2.71565
R1428 VDD2.n164 VDD2.n163 2.71565
R1429 VDD2.n136 VDD2.n135 2.71565
R1430 VDD2.n40 VDD2.n39 2.71565
R1431 VDD2.n68 VDD2.n67 2.71565
R1432 VDD2.n86 VDD2.n2 2.71565
R1433 VDD2.n180 VDD2.n99 1.93989
R1434 VDD2.n167 VDD2.n105 1.93989
R1435 VDD2.n132 VDD2.n122 1.93989
R1436 VDD2.n36 VDD2.n26 1.93989
R1437 VDD2.n72 VDD2.n10 1.93989
R1438 VDD2.n85 VDD2.n4 1.93989
R1439 VDD2.n189 VDD2.t4 1.93763
R1440 VDD2.n189 VDD2.t3 1.93763
R1441 VDD2.n93 VDD2.t1 1.93763
R1442 VDD2.n93 VDD2.t2 1.93763
R1443 VDD2 VDD2.n188 1.51343
R1444 VDD2.n177 VDD2.n176 1.16414
R1445 VDD2.n168 VDD2.n103 1.16414
R1446 VDD2.n131 VDD2.n124 1.16414
R1447 VDD2.n35 VDD2.n28 1.16414
R1448 VDD2.n73 VDD2.n8 1.16414
R1449 VDD2.n82 VDD2.n81 1.16414
R1450 VDD2.n173 VDD2.n101 0.388379
R1451 VDD2.n172 VDD2.n171 0.388379
R1452 VDD2.n128 VDD2.n127 0.388379
R1453 VDD2.n32 VDD2.n31 0.388379
R1454 VDD2.n77 VDD2.n76 0.388379
R1455 VDD2.n78 VDD2.n6 0.388379
R1456 VDD2.n186 VDD2.n96 0.155672
R1457 VDD2.n179 VDD2.n96 0.155672
R1458 VDD2.n179 VDD2.n178 0.155672
R1459 VDD2.n178 VDD2.n100 0.155672
R1460 VDD2.n170 VDD2.n100 0.155672
R1461 VDD2.n170 VDD2.n169 0.155672
R1462 VDD2.n169 VDD2.n104 0.155672
R1463 VDD2.n162 VDD2.n104 0.155672
R1464 VDD2.n162 VDD2.n161 0.155672
R1465 VDD2.n161 VDD2.n109 0.155672
R1466 VDD2.n154 VDD2.n109 0.155672
R1467 VDD2.n154 VDD2.n153 0.155672
R1468 VDD2.n153 VDD2.n113 0.155672
R1469 VDD2.n146 VDD2.n113 0.155672
R1470 VDD2.n146 VDD2.n145 0.155672
R1471 VDD2.n145 VDD2.n117 0.155672
R1472 VDD2.n138 VDD2.n117 0.155672
R1473 VDD2.n138 VDD2.n137 0.155672
R1474 VDD2.n137 VDD2.n121 0.155672
R1475 VDD2.n130 VDD2.n121 0.155672
R1476 VDD2.n130 VDD2.n129 0.155672
R1477 VDD2.n34 VDD2.n33 0.155672
R1478 VDD2.n34 VDD2.n25 0.155672
R1479 VDD2.n41 VDD2.n25 0.155672
R1480 VDD2.n42 VDD2.n41 0.155672
R1481 VDD2.n42 VDD2.n21 0.155672
R1482 VDD2.n49 VDD2.n21 0.155672
R1483 VDD2.n50 VDD2.n49 0.155672
R1484 VDD2.n50 VDD2.n17 0.155672
R1485 VDD2.n57 VDD2.n17 0.155672
R1486 VDD2.n58 VDD2.n57 0.155672
R1487 VDD2.n58 VDD2.n13 0.155672
R1488 VDD2.n65 VDD2.n13 0.155672
R1489 VDD2.n66 VDD2.n65 0.155672
R1490 VDD2.n66 VDD2.n9 0.155672
R1491 VDD2.n74 VDD2.n9 0.155672
R1492 VDD2.n75 VDD2.n74 0.155672
R1493 VDD2.n75 VDD2.n5 0.155672
R1494 VDD2.n83 VDD2.n5 0.155672
R1495 VDD2.n84 VDD2.n83 0.155672
R1496 VDD2.n84 VDD2.n1 0.155672
R1497 VDD2.n91 VDD2.n1 0.155672
R1498 VTAIL.n378 VTAIL.n290 756.745
R1499 VTAIL.n90 VTAIL.n2 756.745
R1500 VTAIL.n284 VTAIL.n196 756.745
R1501 VTAIL.n188 VTAIL.n100 756.745
R1502 VTAIL.n321 VTAIL.n320 585
R1503 VTAIL.n318 VTAIL.n317 585
R1504 VTAIL.n327 VTAIL.n326 585
R1505 VTAIL.n329 VTAIL.n328 585
R1506 VTAIL.n314 VTAIL.n313 585
R1507 VTAIL.n335 VTAIL.n334 585
R1508 VTAIL.n337 VTAIL.n336 585
R1509 VTAIL.n310 VTAIL.n309 585
R1510 VTAIL.n343 VTAIL.n342 585
R1511 VTAIL.n345 VTAIL.n344 585
R1512 VTAIL.n306 VTAIL.n305 585
R1513 VTAIL.n351 VTAIL.n350 585
R1514 VTAIL.n353 VTAIL.n352 585
R1515 VTAIL.n302 VTAIL.n301 585
R1516 VTAIL.n359 VTAIL.n358 585
R1517 VTAIL.n362 VTAIL.n361 585
R1518 VTAIL.n360 VTAIL.n298 585
R1519 VTAIL.n367 VTAIL.n297 585
R1520 VTAIL.n369 VTAIL.n368 585
R1521 VTAIL.n371 VTAIL.n370 585
R1522 VTAIL.n294 VTAIL.n293 585
R1523 VTAIL.n377 VTAIL.n376 585
R1524 VTAIL.n379 VTAIL.n378 585
R1525 VTAIL.n33 VTAIL.n32 585
R1526 VTAIL.n30 VTAIL.n29 585
R1527 VTAIL.n39 VTAIL.n38 585
R1528 VTAIL.n41 VTAIL.n40 585
R1529 VTAIL.n26 VTAIL.n25 585
R1530 VTAIL.n47 VTAIL.n46 585
R1531 VTAIL.n49 VTAIL.n48 585
R1532 VTAIL.n22 VTAIL.n21 585
R1533 VTAIL.n55 VTAIL.n54 585
R1534 VTAIL.n57 VTAIL.n56 585
R1535 VTAIL.n18 VTAIL.n17 585
R1536 VTAIL.n63 VTAIL.n62 585
R1537 VTAIL.n65 VTAIL.n64 585
R1538 VTAIL.n14 VTAIL.n13 585
R1539 VTAIL.n71 VTAIL.n70 585
R1540 VTAIL.n74 VTAIL.n73 585
R1541 VTAIL.n72 VTAIL.n10 585
R1542 VTAIL.n79 VTAIL.n9 585
R1543 VTAIL.n81 VTAIL.n80 585
R1544 VTAIL.n83 VTAIL.n82 585
R1545 VTAIL.n6 VTAIL.n5 585
R1546 VTAIL.n89 VTAIL.n88 585
R1547 VTAIL.n91 VTAIL.n90 585
R1548 VTAIL.n285 VTAIL.n284 585
R1549 VTAIL.n283 VTAIL.n282 585
R1550 VTAIL.n200 VTAIL.n199 585
R1551 VTAIL.n277 VTAIL.n276 585
R1552 VTAIL.n275 VTAIL.n274 585
R1553 VTAIL.n273 VTAIL.n203 585
R1554 VTAIL.n207 VTAIL.n204 585
R1555 VTAIL.n268 VTAIL.n267 585
R1556 VTAIL.n266 VTAIL.n265 585
R1557 VTAIL.n209 VTAIL.n208 585
R1558 VTAIL.n260 VTAIL.n259 585
R1559 VTAIL.n258 VTAIL.n257 585
R1560 VTAIL.n213 VTAIL.n212 585
R1561 VTAIL.n252 VTAIL.n251 585
R1562 VTAIL.n250 VTAIL.n249 585
R1563 VTAIL.n217 VTAIL.n216 585
R1564 VTAIL.n244 VTAIL.n243 585
R1565 VTAIL.n242 VTAIL.n241 585
R1566 VTAIL.n221 VTAIL.n220 585
R1567 VTAIL.n236 VTAIL.n235 585
R1568 VTAIL.n234 VTAIL.n233 585
R1569 VTAIL.n225 VTAIL.n224 585
R1570 VTAIL.n228 VTAIL.n227 585
R1571 VTAIL.n189 VTAIL.n188 585
R1572 VTAIL.n187 VTAIL.n186 585
R1573 VTAIL.n104 VTAIL.n103 585
R1574 VTAIL.n181 VTAIL.n180 585
R1575 VTAIL.n179 VTAIL.n178 585
R1576 VTAIL.n177 VTAIL.n107 585
R1577 VTAIL.n111 VTAIL.n108 585
R1578 VTAIL.n172 VTAIL.n171 585
R1579 VTAIL.n170 VTAIL.n169 585
R1580 VTAIL.n113 VTAIL.n112 585
R1581 VTAIL.n164 VTAIL.n163 585
R1582 VTAIL.n162 VTAIL.n161 585
R1583 VTAIL.n117 VTAIL.n116 585
R1584 VTAIL.n156 VTAIL.n155 585
R1585 VTAIL.n154 VTAIL.n153 585
R1586 VTAIL.n121 VTAIL.n120 585
R1587 VTAIL.n148 VTAIL.n147 585
R1588 VTAIL.n146 VTAIL.n145 585
R1589 VTAIL.n125 VTAIL.n124 585
R1590 VTAIL.n140 VTAIL.n139 585
R1591 VTAIL.n138 VTAIL.n137 585
R1592 VTAIL.n129 VTAIL.n128 585
R1593 VTAIL.n132 VTAIL.n131 585
R1594 VTAIL.t1 VTAIL.n226 327.466
R1595 VTAIL.t10 VTAIL.n130 327.466
R1596 VTAIL.t7 VTAIL.n319 327.466
R1597 VTAIL.t3 VTAIL.n31 327.466
R1598 VTAIL.n320 VTAIL.n317 171.744
R1599 VTAIL.n327 VTAIL.n317 171.744
R1600 VTAIL.n328 VTAIL.n327 171.744
R1601 VTAIL.n328 VTAIL.n313 171.744
R1602 VTAIL.n335 VTAIL.n313 171.744
R1603 VTAIL.n336 VTAIL.n335 171.744
R1604 VTAIL.n336 VTAIL.n309 171.744
R1605 VTAIL.n343 VTAIL.n309 171.744
R1606 VTAIL.n344 VTAIL.n343 171.744
R1607 VTAIL.n344 VTAIL.n305 171.744
R1608 VTAIL.n351 VTAIL.n305 171.744
R1609 VTAIL.n352 VTAIL.n351 171.744
R1610 VTAIL.n352 VTAIL.n301 171.744
R1611 VTAIL.n359 VTAIL.n301 171.744
R1612 VTAIL.n361 VTAIL.n359 171.744
R1613 VTAIL.n361 VTAIL.n360 171.744
R1614 VTAIL.n360 VTAIL.n297 171.744
R1615 VTAIL.n369 VTAIL.n297 171.744
R1616 VTAIL.n370 VTAIL.n369 171.744
R1617 VTAIL.n370 VTAIL.n293 171.744
R1618 VTAIL.n377 VTAIL.n293 171.744
R1619 VTAIL.n378 VTAIL.n377 171.744
R1620 VTAIL.n32 VTAIL.n29 171.744
R1621 VTAIL.n39 VTAIL.n29 171.744
R1622 VTAIL.n40 VTAIL.n39 171.744
R1623 VTAIL.n40 VTAIL.n25 171.744
R1624 VTAIL.n47 VTAIL.n25 171.744
R1625 VTAIL.n48 VTAIL.n47 171.744
R1626 VTAIL.n48 VTAIL.n21 171.744
R1627 VTAIL.n55 VTAIL.n21 171.744
R1628 VTAIL.n56 VTAIL.n55 171.744
R1629 VTAIL.n56 VTAIL.n17 171.744
R1630 VTAIL.n63 VTAIL.n17 171.744
R1631 VTAIL.n64 VTAIL.n63 171.744
R1632 VTAIL.n64 VTAIL.n13 171.744
R1633 VTAIL.n71 VTAIL.n13 171.744
R1634 VTAIL.n73 VTAIL.n71 171.744
R1635 VTAIL.n73 VTAIL.n72 171.744
R1636 VTAIL.n72 VTAIL.n9 171.744
R1637 VTAIL.n81 VTAIL.n9 171.744
R1638 VTAIL.n82 VTAIL.n81 171.744
R1639 VTAIL.n82 VTAIL.n5 171.744
R1640 VTAIL.n89 VTAIL.n5 171.744
R1641 VTAIL.n90 VTAIL.n89 171.744
R1642 VTAIL.n284 VTAIL.n283 171.744
R1643 VTAIL.n283 VTAIL.n199 171.744
R1644 VTAIL.n276 VTAIL.n199 171.744
R1645 VTAIL.n276 VTAIL.n275 171.744
R1646 VTAIL.n275 VTAIL.n203 171.744
R1647 VTAIL.n207 VTAIL.n203 171.744
R1648 VTAIL.n267 VTAIL.n207 171.744
R1649 VTAIL.n267 VTAIL.n266 171.744
R1650 VTAIL.n266 VTAIL.n208 171.744
R1651 VTAIL.n259 VTAIL.n208 171.744
R1652 VTAIL.n259 VTAIL.n258 171.744
R1653 VTAIL.n258 VTAIL.n212 171.744
R1654 VTAIL.n251 VTAIL.n212 171.744
R1655 VTAIL.n251 VTAIL.n250 171.744
R1656 VTAIL.n250 VTAIL.n216 171.744
R1657 VTAIL.n243 VTAIL.n216 171.744
R1658 VTAIL.n243 VTAIL.n242 171.744
R1659 VTAIL.n242 VTAIL.n220 171.744
R1660 VTAIL.n235 VTAIL.n220 171.744
R1661 VTAIL.n235 VTAIL.n234 171.744
R1662 VTAIL.n234 VTAIL.n224 171.744
R1663 VTAIL.n227 VTAIL.n224 171.744
R1664 VTAIL.n188 VTAIL.n187 171.744
R1665 VTAIL.n187 VTAIL.n103 171.744
R1666 VTAIL.n180 VTAIL.n103 171.744
R1667 VTAIL.n180 VTAIL.n179 171.744
R1668 VTAIL.n179 VTAIL.n107 171.744
R1669 VTAIL.n111 VTAIL.n107 171.744
R1670 VTAIL.n171 VTAIL.n111 171.744
R1671 VTAIL.n171 VTAIL.n170 171.744
R1672 VTAIL.n170 VTAIL.n112 171.744
R1673 VTAIL.n163 VTAIL.n112 171.744
R1674 VTAIL.n163 VTAIL.n162 171.744
R1675 VTAIL.n162 VTAIL.n116 171.744
R1676 VTAIL.n155 VTAIL.n116 171.744
R1677 VTAIL.n155 VTAIL.n154 171.744
R1678 VTAIL.n154 VTAIL.n120 171.744
R1679 VTAIL.n147 VTAIL.n120 171.744
R1680 VTAIL.n147 VTAIL.n146 171.744
R1681 VTAIL.n146 VTAIL.n124 171.744
R1682 VTAIL.n139 VTAIL.n124 171.744
R1683 VTAIL.n139 VTAIL.n138 171.744
R1684 VTAIL.n138 VTAIL.n128 171.744
R1685 VTAIL.n131 VTAIL.n128 171.744
R1686 VTAIL.n320 VTAIL.t7 85.8723
R1687 VTAIL.n32 VTAIL.t3 85.8723
R1688 VTAIL.n227 VTAIL.t1 85.8723
R1689 VTAIL.n131 VTAIL.t10 85.8723
R1690 VTAIL.n195 VTAIL.n194 52.3254
R1691 VTAIL.n99 VTAIL.n98 52.3254
R1692 VTAIL.n1 VTAIL.n0 52.3252
R1693 VTAIL.n97 VTAIL.n96 52.3252
R1694 VTAIL.n383 VTAIL.n382 31.7975
R1695 VTAIL.n95 VTAIL.n94 31.7975
R1696 VTAIL.n289 VTAIL.n288 31.7975
R1697 VTAIL.n193 VTAIL.n192 31.7975
R1698 VTAIL.n99 VTAIL.n97 30.7117
R1699 VTAIL.n383 VTAIL.n289 28.7721
R1700 VTAIL.n321 VTAIL.n319 16.3895
R1701 VTAIL.n33 VTAIL.n31 16.3895
R1702 VTAIL.n228 VTAIL.n226 16.3895
R1703 VTAIL.n132 VTAIL.n130 16.3895
R1704 VTAIL.n368 VTAIL.n367 13.1884
R1705 VTAIL.n80 VTAIL.n79 13.1884
R1706 VTAIL.n274 VTAIL.n273 13.1884
R1707 VTAIL.n178 VTAIL.n177 13.1884
R1708 VTAIL.n322 VTAIL.n318 12.8005
R1709 VTAIL.n366 VTAIL.n298 12.8005
R1710 VTAIL.n371 VTAIL.n296 12.8005
R1711 VTAIL.n34 VTAIL.n30 12.8005
R1712 VTAIL.n78 VTAIL.n10 12.8005
R1713 VTAIL.n83 VTAIL.n8 12.8005
R1714 VTAIL.n277 VTAIL.n202 12.8005
R1715 VTAIL.n272 VTAIL.n204 12.8005
R1716 VTAIL.n229 VTAIL.n225 12.8005
R1717 VTAIL.n181 VTAIL.n106 12.8005
R1718 VTAIL.n176 VTAIL.n108 12.8005
R1719 VTAIL.n133 VTAIL.n129 12.8005
R1720 VTAIL.n326 VTAIL.n325 12.0247
R1721 VTAIL.n363 VTAIL.n362 12.0247
R1722 VTAIL.n372 VTAIL.n294 12.0247
R1723 VTAIL.n38 VTAIL.n37 12.0247
R1724 VTAIL.n75 VTAIL.n74 12.0247
R1725 VTAIL.n84 VTAIL.n6 12.0247
R1726 VTAIL.n278 VTAIL.n200 12.0247
R1727 VTAIL.n269 VTAIL.n268 12.0247
R1728 VTAIL.n233 VTAIL.n232 12.0247
R1729 VTAIL.n182 VTAIL.n104 12.0247
R1730 VTAIL.n173 VTAIL.n172 12.0247
R1731 VTAIL.n137 VTAIL.n136 12.0247
R1732 VTAIL.n329 VTAIL.n316 11.249
R1733 VTAIL.n358 VTAIL.n300 11.249
R1734 VTAIL.n376 VTAIL.n375 11.249
R1735 VTAIL.n41 VTAIL.n28 11.249
R1736 VTAIL.n70 VTAIL.n12 11.249
R1737 VTAIL.n88 VTAIL.n87 11.249
R1738 VTAIL.n282 VTAIL.n281 11.249
R1739 VTAIL.n265 VTAIL.n206 11.249
R1740 VTAIL.n236 VTAIL.n223 11.249
R1741 VTAIL.n186 VTAIL.n185 11.249
R1742 VTAIL.n169 VTAIL.n110 11.249
R1743 VTAIL.n140 VTAIL.n127 11.249
R1744 VTAIL.n330 VTAIL.n314 10.4732
R1745 VTAIL.n357 VTAIL.n302 10.4732
R1746 VTAIL.n379 VTAIL.n292 10.4732
R1747 VTAIL.n42 VTAIL.n26 10.4732
R1748 VTAIL.n69 VTAIL.n14 10.4732
R1749 VTAIL.n91 VTAIL.n4 10.4732
R1750 VTAIL.n285 VTAIL.n198 10.4732
R1751 VTAIL.n264 VTAIL.n209 10.4732
R1752 VTAIL.n237 VTAIL.n221 10.4732
R1753 VTAIL.n189 VTAIL.n102 10.4732
R1754 VTAIL.n168 VTAIL.n113 10.4732
R1755 VTAIL.n141 VTAIL.n125 10.4732
R1756 VTAIL.n334 VTAIL.n333 9.69747
R1757 VTAIL.n354 VTAIL.n353 9.69747
R1758 VTAIL.n380 VTAIL.n290 9.69747
R1759 VTAIL.n46 VTAIL.n45 9.69747
R1760 VTAIL.n66 VTAIL.n65 9.69747
R1761 VTAIL.n92 VTAIL.n2 9.69747
R1762 VTAIL.n286 VTAIL.n196 9.69747
R1763 VTAIL.n261 VTAIL.n260 9.69747
R1764 VTAIL.n241 VTAIL.n240 9.69747
R1765 VTAIL.n190 VTAIL.n100 9.69747
R1766 VTAIL.n165 VTAIL.n164 9.69747
R1767 VTAIL.n145 VTAIL.n144 9.69747
R1768 VTAIL.n382 VTAIL.n381 9.45567
R1769 VTAIL.n94 VTAIL.n93 9.45567
R1770 VTAIL.n288 VTAIL.n287 9.45567
R1771 VTAIL.n192 VTAIL.n191 9.45567
R1772 VTAIL.n381 VTAIL.n380 9.3005
R1773 VTAIL.n292 VTAIL.n291 9.3005
R1774 VTAIL.n375 VTAIL.n374 9.3005
R1775 VTAIL.n373 VTAIL.n372 9.3005
R1776 VTAIL.n296 VTAIL.n295 9.3005
R1777 VTAIL.n341 VTAIL.n340 9.3005
R1778 VTAIL.n339 VTAIL.n338 9.3005
R1779 VTAIL.n312 VTAIL.n311 9.3005
R1780 VTAIL.n333 VTAIL.n332 9.3005
R1781 VTAIL.n331 VTAIL.n330 9.3005
R1782 VTAIL.n316 VTAIL.n315 9.3005
R1783 VTAIL.n325 VTAIL.n324 9.3005
R1784 VTAIL.n323 VTAIL.n322 9.3005
R1785 VTAIL.n308 VTAIL.n307 9.3005
R1786 VTAIL.n347 VTAIL.n346 9.3005
R1787 VTAIL.n349 VTAIL.n348 9.3005
R1788 VTAIL.n304 VTAIL.n303 9.3005
R1789 VTAIL.n355 VTAIL.n354 9.3005
R1790 VTAIL.n357 VTAIL.n356 9.3005
R1791 VTAIL.n300 VTAIL.n299 9.3005
R1792 VTAIL.n364 VTAIL.n363 9.3005
R1793 VTAIL.n366 VTAIL.n365 9.3005
R1794 VTAIL.n93 VTAIL.n92 9.3005
R1795 VTAIL.n4 VTAIL.n3 9.3005
R1796 VTAIL.n87 VTAIL.n86 9.3005
R1797 VTAIL.n85 VTAIL.n84 9.3005
R1798 VTAIL.n8 VTAIL.n7 9.3005
R1799 VTAIL.n53 VTAIL.n52 9.3005
R1800 VTAIL.n51 VTAIL.n50 9.3005
R1801 VTAIL.n24 VTAIL.n23 9.3005
R1802 VTAIL.n45 VTAIL.n44 9.3005
R1803 VTAIL.n43 VTAIL.n42 9.3005
R1804 VTAIL.n28 VTAIL.n27 9.3005
R1805 VTAIL.n37 VTAIL.n36 9.3005
R1806 VTAIL.n35 VTAIL.n34 9.3005
R1807 VTAIL.n20 VTAIL.n19 9.3005
R1808 VTAIL.n59 VTAIL.n58 9.3005
R1809 VTAIL.n61 VTAIL.n60 9.3005
R1810 VTAIL.n16 VTAIL.n15 9.3005
R1811 VTAIL.n67 VTAIL.n66 9.3005
R1812 VTAIL.n69 VTAIL.n68 9.3005
R1813 VTAIL.n12 VTAIL.n11 9.3005
R1814 VTAIL.n76 VTAIL.n75 9.3005
R1815 VTAIL.n78 VTAIL.n77 9.3005
R1816 VTAIL.n254 VTAIL.n253 9.3005
R1817 VTAIL.n256 VTAIL.n255 9.3005
R1818 VTAIL.n211 VTAIL.n210 9.3005
R1819 VTAIL.n262 VTAIL.n261 9.3005
R1820 VTAIL.n264 VTAIL.n263 9.3005
R1821 VTAIL.n206 VTAIL.n205 9.3005
R1822 VTAIL.n270 VTAIL.n269 9.3005
R1823 VTAIL.n272 VTAIL.n271 9.3005
R1824 VTAIL.n287 VTAIL.n286 9.3005
R1825 VTAIL.n198 VTAIL.n197 9.3005
R1826 VTAIL.n281 VTAIL.n280 9.3005
R1827 VTAIL.n279 VTAIL.n278 9.3005
R1828 VTAIL.n202 VTAIL.n201 9.3005
R1829 VTAIL.n215 VTAIL.n214 9.3005
R1830 VTAIL.n248 VTAIL.n247 9.3005
R1831 VTAIL.n246 VTAIL.n245 9.3005
R1832 VTAIL.n219 VTAIL.n218 9.3005
R1833 VTAIL.n240 VTAIL.n239 9.3005
R1834 VTAIL.n238 VTAIL.n237 9.3005
R1835 VTAIL.n223 VTAIL.n222 9.3005
R1836 VTAIL.n232 VTAIL.n231 9.3005
R1837 VTAIL.n230 VTAIL.n229 9.3005
R1838 VTAIL.n158 VTAIL.n157 9.3005
R1839 VTAIL.n160 VTAIL.n159 9.3005
R1840 VTAIL.n115 VTAIL.n114 9.3005
R1841 VTAIL.n166 VTAIL.n165 9.3005
R1842 VTAIL.n168 VTAIL.n167 9.3005
R1843 VTAIL.n110 VTAIL.n109 9.3005
R1844 VTAIL.n174 VTAIL.n173 9.3005
R1845 VTAIL.n176 VTAIL.n175 9.3005
R1846 VTAIL.n191 VTAIL.n190 9.3005
R1847 VTAIL.n102 VTAIL.n101 9.3005
R1848 VTAIL.n185 VTAIL.n184 9.3005
R1849 VTAIL.n183 VTAIL.n182 9.3005
R1850 VTAIL.n106 VTAIL.n105 9.3005
R1851 VTAIL.n119 VTAIL.n118 9.3005
R1852 VTAIL.n152 VTAIL.n151 9.3005
R1853 VTAIL.n150 VTAIL.n149 9.3005
R1854 VTAIL.n123 VTAIL.n122 9.3005
R1855 VTAIL.n144 VTAIL.n143 9.3005
R1856 VTAIL.n142 VTAIL.n141 9.3005
R1857 VTAIL.n127 VTAIL.n126 9.3005
R1858 VTAIL.n136 VTAIL.n135 9.3005
R1859 VTAIL.n134 VTAIL.n133 9.3005
R1860 VTAIL.n337 VTAIL.n312 8.92171
R1861 VTAIL.n350 VTAIL.n304 8.92171
R1862 VTAIL.n49 VTAIL.n24 8.92171
R1863 VTAIL.n62 VTAIL.n16 8.92171
R1864 VTAIL.n257 VTAIL.n211 8.92171
R1865 VTAIL.n244 VTAIL.n219 8.92171
R1866 VTAIL.n161 VTAIL.n115 8.92171
R1867 VTAIL.n148 VTAIL.n123 8.92171
R1868 VTAIL.n338 VTAIL.n310 8.14595
R1869 VTAIL.n349 VTAIL.n306 8.14595
R1870 VTAIL.n50 VTAIL.n22 8.14595
R1871 VTAIL.n61 VTAIL.n18 8.14595
R1872 VTAIL.n256 VTAIL.n213 8.14595
R1873 VTAIL.n245 VTAIL.n217 8.14595
R1874 VTAIL.n160 VTAIL.n117 8.14595
R1875 VTAIL.n149 VTAIL.n121 8.14595
R1876 VTAIL.n342 VTAIL.n341 7.3702
R1877 VTAIL.n346 VTAIL.n345 7.3702
R1878 VTAIL.n54 VTAIL.n53 7.3702
R1879 VTAIL.n58 VTAIL.n57 7.3702
R1880 VTAIL.n253 VTAIL.n252 7.3702
R1881 VTAIL.n249 VTAIL.n248 7.3702
R1882 VTAIL.n157 VTAIL.n156 7.3702
R1883 VTAIL.n153 VTAIL.n152 7.3702
R1884 VTAIL.n342 VTAIL.n308 6.59444
R1885 VTAIL.n345 VTAIL.n308 6.59444
R1886 VTAIL.n54 VTAIL.n20 6.59444
R1887 VTAIL.n57 VTAIL.n20 6.59444
R1888 VTAIL.n252 VTAIL.n215 6.59444
R1889 VTAIL.n249 VTAIL.n215 6.59444
R1890 VTAIL.n156 VTAIL.n119 6.59444
R1891 VTAIL.n153 VTAIL.n119 6.59444
R1892 VTAIL.n341 VTAIL.n310 5.81868
R1893 VTAIL.n346 VTAIL.n306 5.81868
R1894 VTAIL.n53 VTAIL.n22 5.81868
R1895 VTAIL.n58 VTAIL.n18 5.81868
R1896 VTAIL.n253 VTAIL.n213 5.81868
R1897 VTAIL.n248 VTAIL.n217 5.81868
R1898 VTAIL.n157 VTAIL.n117 5.81868
R1899 VTAIL.n152 VTAIL.n121 5.81868
R1900 VTAIL.n338 VTAIL.n337 5.04292
R1901 VTAIL.n350 VTAIL.n349 5.04292
R1902 VTAIL.n50 VTAIL.n49 5.04292
R1903 VTAIL.n62 VTAIL.n61 5.04292
R1904 VTAIL.n257 VTAIL.n256 5.04292
R1905 VTAIL.n245 VTAIL.n244 5.04292
R1906 VTAIL.n161 VTAIL.n160 5.04292
R1907 VTAIL.n149 VTAIL.n148 5.04292
R1908 VTAIL.n334 VTAIL.n312 4.26717
R1909 VTAIL.n353 VTAIL.n304 4.26717
R1910 VTAIL.n382 VTAIL.n290 4.26717
R1911 VTAIL.n46 VTAIL.n24 4.26717
R1912 VTAIL.n65 VTAIL.n16 4.26717
R1913 VTAIL.n94 VTAIL.n2 4.26717
R1914 VTAIL.n288 VTAIL.n196 4.26717
R1915 VTAIL.n260 VTAIL.n211 4.26717
R1916 VTAIL.n241 VTAIL.n219 4.26717
R1917 VTAIL.n192 VTAIL.n100 4.26717
R1918 VTAIL.n164 VTAIL.n115 4.26717
R1919 VTAIL.n145 VTAIL.n123 4.26717
R1920 VTAIL.n323 VTAIL.n319 3.70982
R1921 VTAIL.n35 VTAIL.n31 3.70982
R1922 VTAIL.n230 VTAIL.n226 3.70982
R1923 VTAIL.n134 VTAIL.n130 3.70982
R1924 VTAIL.n333 VTAIL.n314 3.49141
R1925 VTAIL.n354 VTAIL.n302 3.49141
R1926 VTAIL.n380 VTAIL.n379 3.49141
R1927 VTAIL.n45 VTAIL.n26 3.49141
R1928 VTAIL.n66 VTAIL.n14 3.49141
R1929 VTAIL.n92 VTAIL.n91 3.49141
R1930 VTAIL.n286 VTAIL.n285 3.49141
R1931 VTAIL.n261 VTAIL.n209 3.49141
R1932 VTAIL.n240 VTAIL.n221 3.49141
R1933 VTAIL.n190 VTAIL.n189 3.49141
R1934 VTAIL.n165 VTAIL.n113 3.49141
R1935 VTAIL.n144 VTAIL.n125 3.49141
R1936 VTAIL.n330 VTAIL.n329 2.71565
R1937 VTAIL.n358 VTAIL.n357 2.71565
R1938 VTAIL.n376 VTAIL.n292 2.71565
R1939 VTAIL.n42 VTAIL.n41 2.71565
R1940 VTAIL.n70 VTAIL.n69 2.71565
R1941 VTAIL.n88 VTAIL.n4 2.71565
R1942 VTAIL.n282 VTAIL.n198 2.71565
R1943 VTAIL.n265 VTAIL.n264 2.71565
R1944 VTAIL.n237 VTAIL.n236 2.71565
R1945 VTAIL.n186 VTAIL.n102 2.71565
R1946 VTAIL.n169 VTAIL.n168 2.71565
R1947 VTAIL.n141 VTAIL.n140 2.71565
R1948 VTAIL.n193 VTAIL.n99 1.94016
R1949 VTAIL.n289 VTAIL.n195 1.94016
R1950 VTAIL.n97 VTAIL.n95 1.94016
R1951 VTAIL.n326 VTAIL.n316 1.93989
R1952 VTAIL.n362 VTAIL.n300 1.93989
R1953 VTAIL.n375 VTAIL.n294 1.93989
R1954 VTAIL.n38 VTAIL.n28 1.93989
R1955 VTAIL.n74 VTAIL.n12 1.93989
R1956 VTAIL.n87 VTAIL.n6 1.93989
R1957 VTAIL.n281 VTAIL.n200 1.93989
R1958 VTAIL.n268 VTAIL.n206 1.93989
R1959 VTAIL.n233 VTAIL.n223 1.93989
R1960 VTAIL.n185 VTAIL.n104 1.93989
R1961 VTAIL.n172 VTAIL.n110 1.93989
R1962 VTAIL.n137 VTAIL.n127 1.93989
R1963 VTAIL.n0 VTAIL.t9 1.93763
R1964 VTAIL.n0 VTAIL.t11 1.93763
R1965 VTAIL.n96 VTAIL.t4 1.93763
R1966 VTAIL.n96 VTAIL.t0 1.93763
R1967 VTAIL.n194 VTAIL.t5 1.93763
R1968 VTAIL.n194 VTAIL.t2 1.93763
R1969 VTAIL.n98 VTAIL.t8 1.93763
R1970 VTAIL.n98 VTAIL.t6 1.93763
R1971 VTAIL.n195 VTAIL.n193 1.44016
R1972 VTAIL.n95 VTAIL.n1 1.44016
R1973 VTAIL VTAIL.n383 1.39705
R1974 VTAIL.n325 VTAIL.n318 1.16414
R1975 VTAIL.n363 VTAIL.n298 1.16414
R1976 VTAIL.n372 VTAIL.n371 1.16414
R1977 VTAIL.n37 VTAIL.n30 1.16414
R1978 VTAIL.n75 VTAIL.n10 1.16414
R1979 VTAIL.n84 VTAIL.n83 1.16414
R1980 VTAIL.n278 VTAIL.n277 1.16414
R1981 VTAIL.n269 VTAIL.n204 1.16414
R1982 VTAIL.n232 VTAIL.n225 1.16414
R1983 VTAIL.n182 VTAIL.n181 1.16414
R1984 VTAIL.n173 VTAIL.n108 1.16414
R1985 VTAIL.n136 VTAIL.n129 1.16414
R1986 VTAIL VTAIL.n1 0.543603
R1987 VTAIL.n322 VTAIL.n321 0.388379
R1988 VTAIL.n367 VTAIL.n366 0.388379
R1989 VTAIL.n368 VTAIL.n296 0.388379
R1990 VTAIL.n34 VTAIL.n33 0.388379
R1991 VTAIL.n79 VTAIL.n78 0.388379
R1992 VTAIL.n80 VTAIL.n8 0.388379
R1993 VTAIL.n274 VTAIL.n202 0.388379
R1994 VTAIL.n273 VTAIL.n272 0.388379
R1995 VTAIL.n229 VTAIL.n228 0.388379
R1996 VTAIL.n178 VTAIL.n106 0.388379
R1997 VTAIL.n177 VTAIL.n176 0.388379
R1998 VTAIL.n133 VTAIL.n132 0.388379
R1999 VTAIL.n324 VTAIL.n323 0.155672
R2000 VTAIL.n324 VTAIL.n315 0.155672
R2001 VTAIL.n331 VTAIL.n315 0.155672
R2002 VTAIL.n332 VTAIL.n331 0.155672
R2003 VTAIL.n332 VTAIL.n311 0.155672
R2004 VTAIL.n339 VTAIL.n311 0.155672
R2005 VTAIL.n340 VTAIL.n339 0.155672
R2006 VTAIL.n340 VTAIL.n307 0.155672
R2007 VTAIL.n347 VTAIL.n307 0.155672
R2008 VTAIL.n348 VTAIL.n347 0.155672
R2009 VTAIL.n348 VTAIL.n303 0.155672
R2010 VTAIL.n355 VTAIL.n303 0.155672
R2011 VTAIL.n356 VTAIL.n355 0.155672
R2012 VTAIL.n356 VTAIL.n299 0.155672
R2013 VTAIL.n364 VTAIL.n299 0.155672
R2014 VTAIL.n365 VTAIL.n364 0.155672
R2015 VTAIL.n365 VTAIL.n295 0.155672
R2016 VTAIL.n373 VTAIL.n295 0.155672
R2017 VTAIL.n374 VTAIL.n373 0.155672
R2018 VTAIL.n374 VTAIL.n291 0.155672
R2019 VTAIL.n381 VTAIL.n291 0.155672
R2020 VTAIL.n36 VTAIL.n35 0.155672
R2021 VTAIL.n36 VTAIL.n27 0.155672
R2022 VTAIL.n43 VTAIL.n27 0.155672
R2023 VTAIL.n44 VTAIL.n43 0.155672
R2024 VTAIL.n44 VTAIL.n23 0.155672
R2025 VTAIL.n51 VTAIL.n23 0.155672
R2026 VTAIL.n52 VTAIL.n51 0.155672
R2027 VTAIL.n52 VTAIL.n19 0.155672
R2028 VTAIL.n59 VTAIL.n19 0.155672
R2029 VTAIL.n60 VTAIL.n59 0.155672
R2030 VTAIL.n60 VTAIL.n15 0.155672
R2031 VTAIL.n67 VTAIL.n15 0.155672
R2032 VTAIL.n68 VTAIL.n67 0.155672
R2033 VTAIL.n68 VTAIL.n11 0.155672
R2034 VTAIL.n76 VTAIL.n11 0.155672
R2035 VTAIL.n77 VTAIL.n76 0.155672
R2036 VTAIL.n77 VTAIL.n7 0.155672
R2037 VTAIL.n85 VTAIL.n7 0.155672
R2038 VTAIL.n86 VTAIL.n85 0.155672
R2039 VTAIL.n86 VTAIL.n3 0.155672
R2040 VTAIL.n93 VTAIL.n3 0.155672
R2041 VTAIL.n287 VTAIL.n197 0.155672
R2042 VTAIL.n280 VTAIL.n197 0.155672
R2043 VTAIL.n280 VTAIL.n279 0.155672
R2044 VTAIL.n279 VTAIL.n201 0.155672
R2045 VTAIL.n271 VTAIL.n201 0.155672
R2046 VTAIL.n271 VTAIL.n270 0.155672
R2047 VTAIL.n270 VTAIL.n205 0.155672
R2048 VTAIL.n263 VTAIL.n205 0.155672
R2049 VTAIL.n263 VTAIL.n262 0.155672
R2050 VTAIL.n262 VTAIL.n210 0.155672
R2051 VTAIL.n255 VTAIL.n210 0.155672
R2052 VTAIL.n255 VTAIL.n254 0.155672
R2053 VTAIL.n254 VTAIL.n214 0.155672
R2054 VTAIL.n247 VTAIL.n214 0.155672
R2055 VTAIL.n247 VTAIL.n246 0.155672
R2056 VTAIL.n246 VTAIL.n218 0.155672
R2057 VTAIL.n239 VTAIL.n218 0.155672
R2058 VTAIL.n239 VTAIL.n238 0.155672
R2059 VTAIL.n238 VTAIL.n222 0.155672
R2060 VTAIL.n231 VTAIL.n222 0.155672
R2061 VTAIL.n231 VTAIL.n230 0.155672
R2062 VTAIL.n191 VTAIL.n101 0.155672
R2063 VTAIL.n184 VTAIL.n101 0.155672
R2064 VTAIL.n184 VTAIL.n183 0.155672
R2065 VTAIL.n183 VTAIL.n105 0.155672
R2066 VTAIL.n175 VTAIL.n105 0.155672
R2067 VTAIL.n175 VTAIL.n174 0.155672
R2068 VTAIL.n174 VTAIL.n109 0.155672
R2069 VTAIL.n167 VTAIL.n109 0.155672
R2070 VTAIL.n167 VTAIL.n166 0.155672
R2071 VTAIL.n166 VTAIL.n114 0.155672
R2072 VTAIL.n159 VTAIL.n114 0.155672
R2073 VTAIL.n159 VTAIL.n158 0.155672
R2074 VTAIL.n158 VTAIL.n118 0.155672
R2075 VTAIL.n151 VTAIL.n118 0.155672
R2076 VTAIL.n151 VTAIL.n150 0.155672
R2077 VTAIL.n150 VTAIL.n122 0.155672
R2078 VTAIL.n143 VTAIL.n122 0.155672
R2079 VTAIL.n143 VTAIL.n142 0.155672
R2080 VTAIL.n142 VTAIL.n126 0.155672
R2081 VTAIL.n135 VTAIL.n126 0.155672
R2082 VTAIL.n135 VTAIL.n134 0.155672
R2083 VP.n6 VP.t0 241.974
R2084 VP.n31 VP.t2 210.625
R2085 VP.n17 VP.t1 210.625
R2086 VP.n24 VP.t5 210.625
R2087 VP.n14 VP.t3 210.625
R2088 VP.n7 VP.t4 210.625
R2089 VP.n9 VP.n8 161.3
R2090 VP.n10 VP.n5 161.3
R2091 VP.n12 VP.n11 161.3
R2092 VP.n13 VP.n4 161.3
R2093 VP.n30 VP.n0 161.3
R2094 VP.n29 VP.n28 161.3
R2095 VP.n27 VP.n1 161.3
R2096 VP.n26 VP.n25 161.3
R2097 VP.n23 VP.n2 161.3
R2098 VP.n22 VP.n21 161.3
R2099 VP.n20 VP.n3 161.3
R2100 VP.n19 VP.n18 161.3
R2101 VP.n17 VP.n16 86.2628
R2102 VP.n32 VP.n31 86.2628
R2103 VP.n15 VP.n14 86.2628
R2104 VP.n7 VP.n6 57.7705
R2105 VP.n22 VP.n3 52.5823
R2106 VP.n29 VP.n1 52.5823
R2107 VP.n12 VP.n5 52.5823
R2108 VP.n16 VP.n15 49.7079
R2109 VP.n18 VP.n3 28.2389
R2110 VP.n30 VP.n29 28.2389
R2111 VP.n13 VP.n12 28.2389
R2112 VP.n18 VP.n17 24.3439
R2113 VP.n23 VP.n22 24.3439
R2114 VP.n25 VP.n1 24.3439
R2115 VP.n31 VP.n30 24.3439
R2116 VP.n14 VP.n13 24.3439
R2117 VP.n8 VP.n5 24.3439
R2118 VP.n9 VP.n6 12.6525
R2119 VP.n24 VP.n23 12.1722
R2120 VP.n25 VP.n24 12.1722
R2121 VP.n8 VP.n7 12.1722
R2122 VP.n15 VP.n4 0.278398
R2123 VP.n19 VP.n16 0.278398
R2124 VP.n32 VP.n0 0.278398
R2125 VP.n10 VP.n9 0.189894
R2126 VP.n11 VP.n10 0.189894
R2127 VP.n11 VP.n4 0.189894
R2128 VP.n20 VP.n19 0.189894
R2129 VP.n21 VP.n20 0.189894
R2130 VP.n21 VP.n2 0.189894
R2131 VP.n26 VP.n2 0.189894
R2132 VP.n27 VP.n26 0.189894
R2133 VP.n28 VP.n27 0.189894
R2134 VP.n28 VP.n0 0.189894
R2135 VP VP.n32 0.153422
R2136 VDD1.n88 VDD1.n0 756.745
R2137 VDD1.n181 VDD1.n93 756.745
R2138 VDD1.n89 VDD1.n88 585
R2139 VDD1.n87 VDD1.n86 585
R2140 VDD1.n4 VDD1.n3 585
R2141 VDD1.n81 VDD1.n80 585
R2142 VDD1.n79 VDD1.n78 585
R2143 VDD1.n77 VDD1.n7 585
R2144 VDD1.n11 VDD1.n8 585
R2145 VDD1.n72 VDD1.n71 585
R2146 VDD1.n70 VDD1.n69 585
R2147 VDD1.n13 VDD1.n12 585
R2148 VDD1.n64 VDD1.n63 585
R2149 VDD1.n62 VDD1.n61 585
R2150 VDD1.n17 VDD1.n16 585
R2151 VDD1.n56 VDD1.n55 585
R2152 VDD1.n54 VDD1.n53 585
R2153 VDD1.n21 VDD1.n20 585
R2154 VDD1.n48 VDD1.n47 585
R2155 VDD1.n46 VDD1.n45 585
R2156 VDD1.n25 VDD1.n24 585
R2157 VDD1.n40 VDD1.n39 585
R2158 VDD1.n38 VDD1.n37 585
R2159 VDD1.n29 VDD1.n28 585
R2160 VDD1.n32 VDD1.n31 585
R2161 VDD1.n124 VDD1.n123 585
R2162 VDD1.n121 VDD1.n120 585
R2163 VDD1.n130 VDD1.n129 585
R2164 VDD1.n132 VDD1.n131 585
R2165 VDD1.n117 VDD1.n116 585
R2166 VDD1.n138 VDD1.n137 585
R2167 VDD1.n140 VDD1.n139 585
R2168 VDD1.n113 VDD1.n112 585
R2169 VDD1.n146 VDD1.n145 585
R2170 VDD1.n148 VDD1.n147 585
R2171 VDD1.n109 VDD1.n108 585
R2172 VDD1.n154 VDD1.n153 585
R2173 VDD1.n156 VDD1.n155 585
R2174 VDD1.n105 VDD1.n104 585
R2175 VDD1.n162 VDD1.n161 585
R2176 VDD1.n165 VDD1.n164 585
R2177 VDD1.n163 VDD1.n101 585
R2178 VDD1.n170 VDD1.n100 585
R2179 VDD1.n172 VDD1.n171 585
R2180 VDD1.n174 VDD1.n173 585
R2181 VDD1.n97 VDD1.n96 585
R2182 VDD1.n180 VDD1.n179 585
R2183 VDD1.n182 VDD1.n181 585
R2184 VDD1.t5 VDD1.n30 327.466
R2185 VDD1.t4 VDD1.n122 327.466
R2186 VDD1.n88 VDD1.n87 171.744
R2187 VDD1.n87 VDD1.n3 171.744
R2188 VDD1.n80 VDD1.n3 171.744
R2189 VDD1.n80 VDD1.n79 171.744
R2190 VDD1.n79 VDD1.n7 171.744
R2191 VDD1.n11 VDD1.n7 171.744
R2192 VDD1.n71 VDD1.n11 171.744
R2193 VDD1.n71 VDD1.n70 171.744
R2194 VDD1.n70 VDD1.n12 171.744
R2195 VDD1.n63 VDD1.n12 171.744
R2196 VDD1.n63 VDD1.n62 171.744
R2197 VDD1.n62 VDD1.n16 171.744
R2198 VDD1.n55 VDD1.n16 171.744
R2199 VDD1.n55 VDD1.n54 171.744
R2200 VDD1.n54 VDD1.n20 171.744
R2201 VDD1.n47 VDD1.n20 171.744
R2202 VDD1.n47 VDD1.n46 171.744
R2203 VDD1.n46 VDD1.n24 171.744
R2204 VDD1.n39 VDD1.n24 171.744
R2205 VDD1.n39 VDD1.n38 171.744
R2206 VDD1.n38 VDD1.n28 171.744
R2207 VDD1.n31 VDD1.n28 171.744
R2208 VDD1.n123 VDD1.n120 171.744
R2209 VDD1.n130 VDD1.n120 171.744
R2210 VDD1.n131 VDD1.n130 171.744
R2211 VDD1.n131 VDD1.n116 171.744
R2212 VDD1.n138 VDD1.n116 171.744
R2213 VDD1.n139 VDD1.n138 171.744
R2214 VDD1.n139 VDD1.n112 171.744
R2215 VDD1.n146 VDD1.n112 171.744
R2216 VDD1.n147 VDD1.n146 171.744
R2217 VDD1.n147 VDD1.n108 171.744
R2218 VDD1.n154 VDD1.n108 171.744
R2219 VDD1.n155 VDD1.n154 171.744
R2220 VDD1.n155 VDD1.n104 171.744
R2221 VDD1.n162 VDD1.n104 171.744
R2222 VDD1.n164 VDD1.n162 171.744
R2223 VDD1.n164 VDD1.n163 171.744
R2224 VDD1.n163 VDD1.n100 171.744
R2225 VDD1.n172 VDD1.n100 171.744
R2226 VDD1.n173 VDD1.n172 171.744
R2227 VDD1.n173 VDD1.n96 171.744
R2228 VDD1.n180 VDD1.n96 171.744
R2229 VDD1.n181 VDD1.n180 171.744
R2230 VDD1.n31 VDD1.t5 85.8723
R2231 VDD1.n123 VDD1.t4 85.8723
R2232 VDD1.n187 VDD1.n186 69.4335
R2233 VDD1.n189 VDD1.n188 69.004
R2234 VDD1 VDD1.n92 49.9892
R2235 VDD1.n187 VDD1.n185 49.8757
R2236 VDD1.n189 VDD1.n187 46.0375
R2237 VDD1.n32 VDD1.n30 16.3895
R2238 VDD1.n124 VDD1.n122 16.3895
R2239 VDD1.n78 VDD1.n77 13.1884
R2240 VDD1.n171 VDD1.n170 13.1884
R2241 VDD1.n81 VDD1.n6 12.8005
R2242 VDD1.n76 VDD1.n8 12.8005
R2243 VDD1.n33 VDD1.n29 12.8005
R2244 VDD1.n125 VDD1.n121 12.8005
R2245 VDD1.n169 VDD1.n101 12.8005
R2246 VDD1.n174 VDD1.n99 12.8005
R2247 VDD1.n82 VDD1.n4 12.0247
R2248 VDD1.n73 VDD1.n72 12.0247
R2249 VDD1.n37 VDD1.n36 12.0247
R2250 VDD1.n129 VDD1.n128 12.0247
R2251 VDD1.n166 VDD1.n165 12.0247
R2252 VDD1.n175 VDD1.n97 12.0247
R2253 VDD1.n86 VDD1.n85 11.249
R2254 VDD1.n69 VDD1.n10 11.249
R2255 VDD1.n40 VDD1.n27 11.249
R2256 VDD1.n132 VDD1.n119 11.249
R2257 VDD1.n161 VDD1.n103 11.249
R2258 VDD1.n179 VDD1.n178 11.249
R2259 VDD1.n89 VDD1.n2 10.4732
R2260 VDD1.n68 VDD1.n13 10.4732
R2261 VDD1.n41 VDD1.n25 10.4732
R2262 VDD1.n133 VDD1.n117 10.4732
R2263 VDD1.n160 VDD1.n105 10.4732
R2264 VDD1.n182 VDD1.n95 10.4732
R2265 VDD1.n90 VDD1.n0 9.69747
R2266 VDD1.n65 VDD1.n64 9.69747
R2267 VDD1.n45 VDD1.n44 9.69747
R2268 VDD1.n137 VDD1.n136 9.69747
R2269 VDD1.n157 VDD1.n156 9.69747
R2270 VDD1.n183 VDD1.n93 9.69747
R2271 VDD1.n92 VDD1.n91 9.45567
R2272 VDD1.n185 VDD1.n184 9.45567
R2273 VDD1.n58 VDD1.n57 9.3005
R2274 VDD1.n60 VDD1.n59 9.3005
R2275 VDD1.n15 VDD1.n14 9.3005
R2276 VDD1.n66 VDD1.n65 9.3005
R2277 VDD1.n68 VDD1.n67 9.3005
R2278 VDD1.n10 VDD1.n9 9.3005
R2279 VDD1.n74 VDD1.n73 9.3005
R2280 VDD1.n76 VDD1.n75 9.3005
R2281 VDD1.n91 VDD1.n90 9.3005
R2282 VDD1.n2 VDD1.n1 9.3005
R2283 VDD1.n85 VDD1.n84 9.3005
R2284 VDD1.n83 VDD1.n82 9.3005
R2285 VDD1.n6 VDD1.n5 9.3005
R2286 VDD1.n19 VDD1.n18 9.3005
R2287 VDD1.n52 VDD1.n51 9.3005
R2288 VDD1.n50 VDD1.n49 9.3005
R2289 VDD1.n23 VDD1.n22 9.3005
R2290 VDD1.n44 VDD1.n43 9.3005
R2291 VDD1.n42 VDD1.n41 9.3005
R2292 VDD1.n27 VDD1.n26 9.3005
R2293 VDD1.n36 VDD1.n35 9.3005
R2294 VDD1.n34 VDD1.n33 9.3005
R2295 VDD1.n184 VDD1.n183 9.3005
R2296 VDD1.n95 VDD1.n94 9.3005
R2297 VDD1.n178 VDD1.n177 9.3005
R2298 VDD1.n176 VDD1.n175 9.3005
R2299 VDD1.n99 VDD1.n98 9.3005
R2300 VDD1.n144 VDD1.n143 9.3005
R2301 VDD1.n142 VDD1.n141 9.3005
R2302 VDD1.n115 VDD1.n114 9.3005
R2303 VDD1.n136 VDD1.n135 9.3005
R2304 VDD1.n134 VDD1.n133 9.3005
R2305 VDD1.n119 VDD1.n118 9.3005
R2306 VDD1.n128 VDD1.n127 9.3005
R2307 VDD1.n126 VDD1.n125 9.3005
R2308 VDD1.n111 VDD1.n110 9.3005
R2309 VDD1.n150 VDD1.n149 9.3005
R2310 VDD1.n152 VDD1.n151 9.3005
R2311 VDD1.n107 VDD1.n106 9.3005
R2312 VDD1.n158 VDD1.n157 9.3005
R2313 VDD1.n160 VDD1.n159 9.3005
R2314 VDD1.n103 VDD1.n102 9.3005
R2315 VDD1.n167 VDD1.n166 9.3005
R2316 VDD1.n169 VDD1.n168 9.3005
R2317 VDD1.n61 VDD1.n15 8.92171
R2318 VDD1.n48 VDD1.n23 8.92171
R2319 VDD1.n140 VDD1.n115 8.92171
R2320 VDD1.n153 VDD1.n107 8.92171
R2321 VDD1.n60 VDD1.n17 8.14595
R2322 VDD1.n49 VDD1.n21 8.14595
R2323 VDD1.n141 VDD1.n113 8.14595
R2324 VDD1.n152 VDD1.n109 8.14595
R2325 VDD1.n57 VDD1.n56 7.3702
R2326 VDD1.n53 VDD1.n52 7.3702
R2327 VDD1.n145 VDD1.n144 7.3702
R2328 VDD1.n149 VDD1.n148 7.3702
R2329 VDD1.n56 VDD1.n19 6.59444
R2330 VDD1.n53 VDD1.n19 6.59444
R2331 VDD1.n145 VDD1.n111 6.59444
R2332 VDD1.n148 VDD1.n111 6.59444
R2333 VDD1.n57 VDD1.n17 5.81868
R2334 VDD1.n52 VDD1.n21 5.81868
R2335 VDD1.n144 VDD1.n113 5.81868
R2336 VDD1.n149 VDD1.n109 5.81868
R2337 VDD1.n61 VDD1.n60 5.04292
R2338 VDD1.n49 VDD1.n48 5.04292
R2339 VDD1.n141 VDD1.n140 5.04292
R2340 VDD1.n153 VDD1.n152 5.04292
R2341 VDD1.n92 VDD1.n0 4.26717
R2342 VDD1.n64 VDD1.n15 4.26717
R2343 VDD1.n45 VDD1.n23 4.26717
R2344 VDD1.n137 VDD1.n115 4.26717
R2345 VDD1.n156 VDD1.n107 4.26717
R2346 VDD1.n185 VDD1.n93 4.26717
R2347 VDD1.n34 VDD1.n30 3.70982
R2348 VDD1.n126 VDD1.n122 3.70982
R2349 VDD1.n90 VDD1.n89 3.49141
R2350 VDD1.n65 VDD1.n13 3.49141
R2351 VDD1.n44 VDD1.n25 3.49141
R2352 VDD1.n136 VDD1.n117 3.49141
R2353 VDD1.n157 VDD1.n105 3.49141
R2354 VDD1.n183 VDD1.n182 3.49141
R2355 VDD1.n86 VDD1.n2 2.71565
R2356 VDD1.n69 VDD1.n68 2.71565
R2357 VDD1.n41 VDD1.n40 2.71565
R2358 VDD1.n133 VDD1.n132 2.71565
R2359 VDD1.n161 VDD1.n160 2.71565
R2360 VDD1.n179 VDD1.n95 2.71565
R2361 VDD1.n85 VDD1.n4 1.93989
R2362 VDD1.n72 VDD1.n10 1.93989
R2363 VDD1.n37 VDD1.n27 1.93989
R2364 VDD1.n129 VDD1.n119 1.93989
R2365 VDD1.n165 VDD1.n103 1.93989
R2366 VDD1.n178 VDD1.n97 1.93989
R2367 VDD1.n188 VDD1.t1 1.93763
R2368 VDD1.n188 VDD1.t2 1.93763
R2369 VDD1.n186 VDD1.t0 1.93763
R2370 VDD1.n186 VDD1.t3 1.93763
R2371 VDD1.n82 VDD1.n81 1.16414
R2372 VDD1.n73 VDD1.n8 1.16414
R2373 VDD1.n36 VDD1.n29 1.16414
R2374 VDD1.n128 VDD1.n121 1.16414
R2375 VDD1.n166 VDD1.n101 1.16414
R2376 VDD1.n175 VDD1.n174 1.16414
R2377 VDD1 VDD1.n189 0.427224
R2378 VDD1.n78 VDD1.n6 0.388379
R2379 VDD1.n77 VDD1.n76 0.388379
R2380 VDD1.n33 VDD1.n32 0.388379
R2381 VDD1.n125 VDD1.n124 0.388379
R2382 VDD1.n170 VDD1.n169 0.388379
R2383 VDD1.n171 VDD1.n99 0.388379
R2384 VDD1.n91 VDD1.n1 0.155672
R2385 VDD1.n84 VDD1.n1 0.155672
R2386 VDD1.n84 VDD1.n83 0.155672
R2387 VDD1.n83 VDD1.n5 0.155672
R2388 VDD1.n75 VDD1.n5 0.155672
R2389 VDD1.n75 VDD1.n74 0.155672
R2390 VDD1.n74 VDD1.n9 0.155672
R2391 VDD1.n67 VDD1.n9 0.155672
R2392 VDD1.n67 VDD1.n66 0.155672
R2393 VDD1.n66 VDD1.n14 0.155672
R2394 VDD1.n59 VDD1.n14 0.155672
R2395 VDD1.n59 VDD1.n58 0.155672
R2396 VDD1.n58 VDD1.n18 0.155672
R2397 VDD1.n51 VDD1.n18 0.155672
R2398 VDD1.n51 VDD1.n50 0.155672
R2399 VDD1.n50 VDD1.n22 0.155672
R2400 VDD1.n43 VDD1.n22 0.155672
R2401 VDD1.n43 VDD1.n42 0.155672
R2402 VDD1.n42 VDD1.n26 0.155672
R2403 VDD1.n35 VDD1.n26 0.155672
R2404 VDD1.n35 VDD1.n34 0.155672
R2405 VDD1.n127 VDD1.n126 0.155672
R2406 VDD1.n127 VDD1.n118 0.155672
R2407 VDD1.n134 VDD1.n118 0.155672
R2408 VDD1.n135 VDD1.n134 0.155672
R2409 VDD1.n135 VDD1.n114 0.155672
R2410 VDD1.n142 VDD1.n114 0.155672
R2411 VDD1.n143 VDD1.n142 0.155672
R2412 VDD1.n143 VDD1.n110 0.155672
R2413 VDD1.n150 VDD1.n110 0.155672
R2414 VDD1.n151 VDD1.n150 0.155672
R2415 VDD1.n151 VDD1.n106 0.155672
R2416 VDD1.n158 VDD1.n106 0.155672
R2417 VDD1.n159 VDD1.n158 0.155672
R2418 VDD1.n159 VDD1.n102 0.155672
R2419 VDD1.n167 VDD1.n102 0.155672
R2420 VDD1.n168 VDD1.n167 0.155672
R2421 VDD1.n168 VDD1.n98 0.155672
R2422 VDD1.n176 VDD1.n98 0.155672
R2423 VDD1.n177 VDD1.n176 0.155672
R2424 VDD1.n177 VDD1.n94 0.155672
R2425 VDD1.n184 VDD1.n94 0.155672
C0 VN VDD1 0.149469f
C1 B VDD1 2.28177f
C2 VN VDD2 8.65248f
C3 VP w_n2770_n4324# 5.53348f
C4 B VDD2 2.33955f
C5 VTAIL VDD1 9.711361f
C6 w_n2770_n4324# VN 5.17725f
C7 VP VN 7.155129f
C8 VTAIL VDD2 9.755269f
C9 B w_n2770_n4324# 10.0767f
C10 B VP 1.66776f
C11 w_n2770_n4324# VTAIL 3.61309f
C12 VP VTAIL 8.46898f
C13 B VN 1.07642f
C14 VN VTAIL 8.454531f
C15 VDD1 VDD2 1.16699f
C16 B VTAIL 4.4081f
C17 w_n2770_n4324# VDD1 2.4632f
C18 VP VDD1 8.89938f
C19 w_n2770_n4324# VDD2 2.52661f
C20 VP VDD2 0.400849f
C21 VDD2 VSUBS 1.858854f
C22 VDD1 VSUBS 1.708927f
C23 VTAIL VSUBS 1.240682f
C24 VN VSUBS 5.47763f
C25 VP VSUBS 2.59377f
C26 B VSUBS 4.369325f
C27 w_n2770_n4324# VSUBS 0.146622p
C28 VDD1.n0 VSUBS 0.028493f
C29 VDD1.n1 VSUBS 0.027079f
C30 VDD1.n2 VSUBS 0.014551f
C31 VDD1.n3 VSUBS 0.034393f
C32 VDD1.n4 VSUBS 0.015407f
C33 VDD1.n5 VSUBS 0.027079f
C34 VDD1.n6 VSUBS 0.014551f
C35 VDD1.n7 VSUBS 0.034393f
C36 VDD1.n8 VSUBS 0.015407f
C37 VDD1.n9 VSUBS 0.027079f
C38 VDD1.n10 VSUBS 0.014551f
C39 VDD1.n11 VSUBS 0.034393f
C40 VDD1.n12 VSUBS 0.034393f
C41 VDD1.n13 VSUBS 0.015407f
C42 VDD1.n14 VSUBS 0.027079f
C43 VDD1.n15 VSUBS 0.014551f
C44 VDD1.n16 VSUBS 0.034393f
C45 VDD1.n17 VSUBS 0.015407f
C46 VDD1.n18 VSUBS 0.027079f
C47 VDD1.n19 VSUBS 0.014551f
C48 VDD1.n20 VSUBS 0.034393f
C49 VDD1.n21 VSUBS 0.015407f
C50 VDD1.n22 VSUBS 0.027079f
C51 VDD1.n23 VSUBS 0.014551f
C52 VDD1.n24 VSUBS 0.034393f
C53 VDD1.n25 VSUBS 0.015407f
C54 VDD1.n26 VSUBS 0.027079f
C55 VDD1.n27 VSUBS 0.014551f
C56 VDD1.n28 VSUBS 0.034393f
C57 VDD1.n29 VSUBS 0.015407f
C58 VDD1.n30 VSUBS 0.205097f
C59 VDD1.t5 VSUBS 0.073748f
C60 VDD1.n31 VSUBS 0.025795f
C61 VDD1.n32 VSUBS 0.021879f
C62 VDD1.n33 VSUBS 0.014551f
C63 VDD1.n34 VSUBS 1.94783f
C64 VDD1.n35 VSUBS 0.027079f
C65 VDD1.n36 VSUBS 0.014551f
C66 VDD1.n37 VSUBS 0.015407f
C67 VDD1.n38 VSUBS 0.034393f
C68 VDD1.n39 VSUBS 0.034393f
C69 VDD1.n40 VSUBS 0.015407f
C70 VDD1.n41 VSUBS 0.014551f
C71 VDD1.n42 VSUBS 0.027079f
C72 VDD1.n43 VSUBS 0.027079f
C73 VDD1.n44 VSUBS 0.014551f
C74 VDD1.n45 VSUBS 0.015407f
C75 VDD1.n46 VSUBS 0.034393f
C76 VDD1.n47 VSUBS 0.034393f
C77 VDD1.n48 VSUBS 0.015407f
C78 VDD1.n49 VSUBS 0.014551f
C79 VDD1.n50 VSUBS 0.027079f
C80 VDD1.n51 VSUBS 0.027079f
C81 VDD1.n52 VSUBS 0.014551f
C82 VDD1.n53 VSUBS 0.015407f
C83 VDD1.n54 VSUBS 0.034393f
C84 VDD1.n55 VSUBS 0.034393f
C85 VDD1.n56 VSUBS 0.015407f
C86 VDD1.n57 VSUBS 0.014551f
C87 VDD1.n58 VSUBS 0.027079f
C88 VDD1.n59 VSUBS 0.027079f
C89 VDD1.n60 VSUBS 0.014551f
C90 VDD1.n61 VSUBS 0.015407f
C91 VDD1.n62 VSUBS 0.034393f
C92 VDD1.n63 VSUBS 0.034393f
C93 VDD1.n64 VSUBS 0.015407f
C94 VDD1.n65 VSUBS 0.014551f
C95 VDD1.n66 VSUBS 0.027079f
C96 VDD1.n67 VSUBS 0.027079f
C97 VDD1.n68 VSUBS 0.014551f
C98 VDD1.n69 VSUBS 0.015407f
C99 VDD1.n70 VSUBS 0.034393f
C100 VDD1.n71 VSUBS 0.034393f
C101 VDD1.n72 VSUBS 0.015407f
C102 VDD1.n73 VSUBS 0.014551f
C103 VDD1.n74 VSUBS 0.027079f
C104 VDD1.n75 VSUBS 0.027079f
C105 VDD1.n76 VSUBS 0.014551f
C106 VDD1.n77 VSUBS 0.014979f
C107 VDD1.n78 VSUBS 0.014979f
C108 VDD1.n79 VSUBS 0.034393f
C109 VDD1.n80 VSUBS 0.034393f
C110 VDD1.n81 VSUBS 0.015407f
C111 VDD1.n82 VSUBS 0.014551f
C112 VDD1.n83 VSUBS 0.027079f
C113 VDD1.n84 VSUBS 0.027079f
C114 VDD1.n85 VSUBS 0.014551f
C115 VDD1.n86 VSUBS 0.015407f
C116 VDD1.n87 VSUBS 0.034393f
C117 VDD1.n88 VSUBS 0.078966f
C118 VDD1.n89 VSUBS 0.015407f
C119 VDD1.n90 VSUBS 0.014551f
C120 VDD1.n91 VSUBS 0.061851f
C121 VDD1.n92 VSUBS 0.063761f
C122 VDD1.n93 VSUBS 0.028493f
C123 VDD1.n94 VSUBS 0.027079f
C124 VDD1.n95 VSUBS 0.014551f
C125 VDD1.n96 VSUBS 0.034393f
C126 VDD1.n97 VSUBS 0.015407f
C127 VDD1.n98 VSUBS 0.027079f
C128 VDD1.n99 VSUBS 0.014551f
C129 VDD1.n100 VSUBS 0.034393f
C130 VDD1.n101 VSUBS 0.015407f
C131 VDD1.n102 VSUBS 0.027079f
C132 VDD1.n103 VSUBS 0.014551f
C133 VDD1.n104 VSUBS 0.034393f
C134 VDD1.n105 VSUBS 0.015407f
C135 VDD1.n106 VSUBS 0.027079f
C136 VDD1.n107 VSUBS 0.014551f
C137 VDD1.n108 VSUBS 0.034393f
C138 VDD1.n109 VSUBS 0.015407f
C139 VDD1.n110 VSUBS 0.027079f
C140 VDD1.n111 VSUBS 0.014551f
C141 VDD1.n112 VSUBS 0.034393f
C142 VDD1.n113 VSUBS 0.015407f
C143 VDD1.n114 VSUBS 0.027079f
C144 VDD1.n115 VSUBS 0.014551f
C145 VDD1.n116 VSUBS 0.034393f
C146 VDD1.n117 VSUBS 0.015407f
C147 VDD1.n118 VSUBS 0.027079f
C148 VDD1.n119 VSUBS 0.014551f
C149 VDD1.n120 VSUBS 0.034393f
C150 VDD1.n121 VSUBS 0.015407f
C151 VDD1.n122 VSUBS 0.205097f
C152 VDD1.t4 VSUBS 0.073748f
C153 VDD1.n123 VSUBS 0.025795f
C154 VDD1.n124 VSUBS 0.021879f
C155 VDD1.n125 VSUBS 0.014551f
C156 VDD1.n126 VSUBS 1.94783f
C157 VDD1.n127 VSUBS 0.027079f
C158 VDD1.n128 VSUBS 0.014551f
C159 VDD1.n129 VSUBS 0.015407f
C160 VDD1.n130 VSUBS 0.034393f
C161 VDD1.n131 VSUBS 0.034393f
C162 VDD1.n132 VSUBS 0.015407f
C163 VDD1.n133 VSUBS 0.014551f
C164 VDD1.n134 VSUBS 0.027079f
C165 VDD1.n135 VSUBS 0.027079f
C166 VDD1.n136 VSUBS 0.014551f
C167 VDD1.n137 VSUBS 0.015407f
C168 VDD1.n138 VSUBS 0.034393f
C169 VDD1.n139 VSUBS 0.034393f
C170 VDD1.n140 VSUBS 0.015407f
C171 VDD1.n141 VSUBS 0.014551f
C172 VDD1.n142 VSUBS 0.027079f
C173 VDD1.n143 VSUBS 0.027079f
C174 VDD1.n144 VSUBS 0.014551f
C175 VDD1.n145 VSUBS 0.015407f
C176 VDD1.n146 VSUBS 0.034393f
C177 VDD1.n147 VSUBS 0.034393f
C178 VDD1.n148 VSUBS 0.015407f
C179 VDD1.n149 VSUBS 0.014551f
C180 VDD1.n150 VSUBS 0.027079f
C181 VDD1.n151 VSUBS 0.027079f
C182 VDD1.n152 VSUBS 0.014551f
C183 VDD1.n153 VSUBS 0.015407f
C184 VDD1.n154 VSUBS 0.034393f
C185 VDD1.n155 VSUBS 0.034393f
C186 VDD1.n156 VSUBS 0.015407f
C187 VDD1.n157 VSUBS 0.014551f
C188 VDD1.n158 VSUBS 0.027079f
C189 VDD1.n159 VSUBS 0.027079f
C190 VDD1.n160 VSUBS 0.014551f
C191 VDD1.n161 VSUBS 0.015407f
C192 VDD1.n162 VSUBS 0.034393f
C193 VDD1.n163 VSUBS 0.034393f
C194 VDD1.n164 VSUBS 0.034393f
C195 VDD1.n165 VSUBS 0.015407f
C196 VDD1.n166 VSUBS 0.014551f
C197 VDD1.n167 VSUBS 0.027079f
C198 VDD1.n168 VSUBS 0.027079f
C199 VDD1.n169 VSUBS 0.014551f
C200 VDD1.n170 VSUBS 0.014979f
C201 VDD1.n171 VSUBS 0.014979f
C202 VDD1.n172 VSUBS 0.034393f
C203 VDD1.n173 VSUBS 0.034393f
C204 VDD1.n174 VSUBS 0.015407f
C205 VDD1.n175 VSUBS 0.014551f
C206 VDD1.n176 VSUBS 0.027079f
C207 VDD1.n177 VSUBS 0.027079f
C208 VDD1.n178 VSUBS 0.014551f
C209 VDD1.n179 VSUBS 0.015407f
C210 VDD1.n180 VSUBS 0.034393f
C211 VDD1.n181 VSUBS 0.078966f
C212 VDD1.n182 VSUBS 0.015407f
C213 VDD1.n183 VSUBS 0.014551f
C214 VDD1.n184 VSUBS 0.061851f
C215 VDD1.n185 VSUBS 0.06309f
C216 VDD1.t0 VSUBS 0.359063f
C217 VDD1.t3 VSUBS 0.359063f
C218 VDD1.n186 VSUBS 2.959f
C219 VDD1.n187 VSUBS 3.32785f
C220 VDD1.t1 VSUBS 0.359063f
C221 VDD1.t2 VSUBS 0.359063f
C222 VDD1.n188 VSUBS 2.95436f
C223 VDD1.n189 VSUBS 3.51687f
C224 VP.n0 VSUBS 0.044757f
C225 VP.t2 VSUBS 3.00403f
C226 VP.n1 VSUBS 0.060886f
C227 VP.n2 VSUBS 0.033946f
C228 VP.t5 VSUBS 3.00403f
C229 VP.n3 VSUBS 0.035017f
C230 VP.n4 VSUBS 0.044757f
C231 VP.t3 VSUBS 3.00403f
C232 VP.n5 VSUBS 0.060886f
C233 VP.t0 VSUBS 3.16226f
C234 VP.n6 VSUBS 1.1433f
C235 VP.t4 VSUBS 3.00403f
C236 VP.n7 VSUBS 1.13263f
C237 VP.n8 VSUBS 0.047887f
C238 VP.n9 VSUBS 0.251463f
C239 VP.n10 VSUBS 0.033946f
C240 VP.n11 VSUBS 0.033946f
C241 VP.n12 VSUBS 0.035017f
C242 VP.n13 VSUBS 0.067221f
C243 VP.n14 VSUBS 1.16338f
C244 VP.n15 VSUBS 1.85302f
C245 VP.n16 VSUBS 1.8775f
C246 VP.t1 VSUBS 3.00403f
C247 VP.n17 VSUBS 1.16338f
C248 VP.n18 VSUBS 0.067221f
C249 VP.n19 VSUBS 0.044757f
C250 VP.n20 VSUBS 0.033946f
C251 VP.n21 VSUBS 0.033946f
C252 VP.n22 VSUBS 0.060886f
C253 VP.n23 VSUBS 0.047887f
C254 VP.n24 VSUBS 1.05303f
C255 VP.n25 VSUBS 0.047887f
C256 VP.n26 VSUBS 0.033946f
C257 VP.n27 VSUBS 0.033946f
C258 VP.n28 VSUBS 0.033946f
C259 VP.n29 VSUBS 0.035017f
C260 VP.n30 VSUBS 0.067221f
C261 VP.n31 VSUBS 1.16338f
C262 VP.n32 VSUBS 0.035876f
C263 VTAIL.t9 VSUBS 0.365048f
C264 VTAIL.t11 VSUBS 0.365048f
C265 VTAIL.n0 VSUBS 2.83317f
C266 VTAIL.n1 VSUBS 0.848836f
C267 VTAIL.n2 VSUBS 0.028967f
C268 VTAIL.n3 VSUBS 0.02753f
C269 VTAIL.n4 VSUBS 0.014793f
C270 VTAIL.n5 VSUBS 0.034966f
C271 VTAIL.n6 VSUBS 0.015664f
C272 VTAIL.n7 VSUBS 0.02753f
C273 VTAIL.n8 VSUBS 0.014793f
C274 VTAIL.n9 VSUBS 0.034966f
C275 VTAIL.n10 VSUBS 0.015664f
C276 VTAIL.n11 VSUBS 0.02753f
C277 VTAIL.n12 VSUBS 0.014793f
C278 VTAIL.n13 VSUBS 0.034966f
C279 VTAIL.n14 VSUBS 0.015664f
C280 VTAIL.n15 VSUBS 0.02753f
C281 VTAIL.n16 VSUBS 0.014793f
C282 VTAIL.n17 VSUBS 0.034966f
C283 VTAIL.n18 VSUBS 0.015664f
C284 VTAIL.n19 VSUBS 0.02753f
C285 VTAIL.n20 VSUBS 0.014793f
C286 VTAIL.n21 VSUBS 0.034966f
C287 VTAIL.n22 VSUBS 0.015664f
C288 VTAIL.n23 VSUBS 0.02753f
C289 VTAIL.n24 VSUBS 0.014793f
C290 VTAIL.n25 VSUBS 0.034966f
C291 VTAIL.n26 VSUBS 0.015664f
C292 VTAIL.n27 VSUBS 0.02753f
C293 VTAIL.n28 VSUBS 0.014793f
C294 VTAIL.n29 VSUBS 0.034966f
C295 VTAIL.n30 VSUBS 0.015664f
C296 VTAIL.n31 VSUBS 0.208515f
C297 VTAIL.t3 VSUBS 0.074977f
C298 VTAIL.n32 VSUBS 0.026225f
C299 VTAIL.n33 VSUBS 0.022244f
C300 VTAIL.n34 VSUBS 0.014793f
C301 VTAIL.n35 VSUBS 1.9803f
C302 VTAIL.n36 VSUBS 0.02753f
C303 VTAIL.n37 VSUBS 0.014793f
C304 VTAIL.n38 VSUBS 0.015664f
C305 VTAIL.n39 VSUBS 0.034966f
C306 VTAIL.n40 VSUBS 0.034966f
C307 VTAIL.n41 VSUBS 0.015664f
C308 VTAIL.n42 VSUBS 0.014793f
C309 VTAIL.n43 VSUBS 0.02753f
C310 VTAIL.n44 VSUBS 0.02753f
C311 VTAIL.n45 VSUBS 0.014793f
C312 VTAIL.n46 VSUBS 0.015664f
C313 VTAIL.n47 VSUBS 0.034966f
C314 VTAIL.n48 VSUBS 0.034966f
C315 VTAIL.n49 VSUBS 0.015664f
C316 VTAIL.n50 VSUBS 0.014793f
C317 VTAIL.n51 VSUBS 0.02753f
C318 VTAIL.n52 VSUBS 0.02753f
C319 VTAIL.n53 VSUBS 0.014793f
C320 VTAIL.n54 VSUBS 0.015664f
C321 VTAIL.n55 VSUBS 0.034966f
C322 VTAIL.n56 VSUBS 0.034966f
C323 VTAIL.n57 VSUBS 0.015664f
C324 VTAIL.n58 VSUBS 0.014793f
C325 VTAIL.n59 VSUBS 0.02753f
C326 VTAIL.n60 VSUBS 0.02753f
C327 VTAIL.n61 VSUBS 0.014793f
C328 VTAIL.n62 VSUBS 0.015664f
C329 VTAIL.n63 VSUBS 0.034966f
C330 VTAIL.n64 VSUBS 0.034966f
C331 VTAIL.n65 VSUBS 0.015664f
C332 VTAIL.n66 VSUBS 0.014793f
C333 VTAIL.n67 VSUBS 0.02753f
C334 VTAIL.n68 VSUBS 0.02753f
C335 VTAIL.n69 VSUBS 0.014793f
C336 VTAIL.n70 VSUBS 0.015664f
C337 VTAIL.n71 VSUBS 0.034966f
C338 VTAIL.n72 VSUBS 0.034966f
C339 VTAIL.n73 VSUBS 0.034966f
C340 VTAIL.n74 VSUBS 0.015664f
C341 VTAIL.n75 VSUBS 0.014793f
C342 VTAIL.n76 VSUBS 0.02753f
C343 VTAIL.n77 VSUBS 0.02753f
C344 VTAIL.n78 VSUBS 0.014793f
C345 VTAIL.n79 VSUBS 0.015229f
C346 VTAIL.n80 VSUBS 0.015229f
C347 VTAIL.n81 VSUBS 0.034966f
C348 VTAIL.n82 VSUBS 0.034966f
C349 VTAIL.n83 VSUBS 0.015664f
C350 VTAIL.n84 VSUBS 0.014793f
C351 VTAIL.n85 VSUBS 0.02753f
C352 VTAIL.n86 VSUBS 0.02753f
C353 VTAIL.n87 VSUBS 0.014793f
C354 VTAIL.n88 VSUBS 0.015664f
C355 VTAIL.n89 VSUBS 0.034966f
C356 VTAIL.n90 VSUBS 0.080282f
C357 VTAIL.n91 VSUBS 0.015664f
C358 VTAIL.n92 VSUBS 0.014793f
C359 VTAIL.n93 VSUBS 0.062882f
C360 VTAIL.n94 VSUBS 0.040156f
C361 VTAIL.n95 VSUBS 0.322858f
C362 VTAIL.t4 VSUBS 0.365048f
C363 VTAIL.t0 VSUBS 0.365048f
C364 VTAIL.n96 VSUBS 2.83317f
C365 VTAIL.n97 VSUBS 2.8463f
C366 VTAIL.t8 VSUBS 0.365048f
C367 VTAIL.t6 VSUBS 0.365048f
C368 VTAIL.n98 VSUBS 2.83319f
C369 VTAIL.n99 VSUBS 2.84628f
C370 VTAIL.n100 VSUBS 0.028967f
C371 VTAIL.n101 VSUBS 0.02753f
C372 VTAIL.n102 VSUBS 0.014793f
C373 VTAIL.n103 VSUBS 0.034966f
C374 VTAIL.n104 VSUBS 0.015664f
C375 VTAIL.n105 VSUBS 0.02753f
C376 VTAIL.n106 VSUBS 0.014793f
C377 VTAIL.n107 VSUBS 0.034966f
C378 VTAIL.n108 VSUBS 0.015664f
C379 VTAIL.n109 VSUBS 0.02753f
C380 VTAIL.n110 VSUBS 0.014793f
C381 VTAIL.n111 VSUBS 0.034966f
C382 VTAIL.n112 VSUBS 0.034966f
C383 VTAIL.n113 VSUBS 0.015664f
C384 VTAIL.n114 VSUBS 0.02753f
C385 VTAIL.n115 VSUBS 0.014793f
C386 VTAIL.n116 VSUBS 0.034966f
C387 VTAIL.n117 VSUBS 0.015664f
C388 VTAIL.n118 VSUBS 0.02753f
C389 VTAIL.n119 VSUBS 0.014793f
C390 VTAIL.n120 VSUBS 0.034966f
C391 VTAIL.n121 VSUBS 0.015664f
C392 VTAIL.n122 VSUBS 0.02753f
C393 VTAIL.n123 VSUBS 0.014793f
C394 VTAIL.n124 VSUBS 0.034966f
C395 VTAIL.n125 VSUBS 0.015664f
C396 VTAIL.n126 VSUBS 0.02753f
C397 VTAIL.n127 VSUBS 0.014793f
C398 VTAIL.n128 VSUBS 0.034966f
C399 VTAIL.n129 VSUBS 0.015664f
C400 VTAIL.n130 VSUBS 0.208515f
C401 VTAIL.t10 VSUBS 0.074977f
C402 VTAIL.n131 VSUBS 0.026225f
C403 VTAIL.n132 VSUBS 0.022244f
C404 VTAIL.n133 VSUBS 0.014793f
C405 VTAIL.n134 VSUBS 1.9803f
C406 VTAIL.n135 VSUBS 0.02753f
C407 VTAIL.n136 VSUBS 0.014793f
C408 VTAIL.n137 VSUBS 0.015664f
C409 VTAIL.n138 VSUBS 0.034966f
C410 VTAIL.n139 VSUBS 0.034966f
C411 VTAIL.n140 VSUBS 0.015664f
C412 VTAIL.n141 VSUBS 0.014793f
C413 VTAIL.n142 VSUBS 0.02753f
C414 VTAIL.n143 VSUBS 0.02753f
C415 VTAIL.n144 VSUBS 0.014793f
C416 VTAIL.n145 VSUBS 0.015664f
C417 VTAIL.n146 VSUBS 0.034966f
C418 VTAIL.n147 VSUBS 0.034966f
C419 VTAIL.n148 VSUBS 0.015664f
C420 VTAIL.n149 VSUBS 0.014793f
C421 VTAIL.n150 VSUBS 0.02753f
C422 VTAIL.n151 VSUBS 0.02753f
C423 VTAIL.n152 VSUBS 0.014793f
C424 VTAIL.n153 VSUBS 0.015664f
C425 VTAIL.n154 VSUBS 0.034966f
C426 VTAIL.n155 VSUBS 0.034966f
C427 VTAIL.n156 VSUBS 0.015664f
C428 VTAIL.n157 VSUBS 0.014793f
C429 VTAIL.n158 VSUBS 0.02753f
C430 VTAIL.n159 VSUBS 0.02753f
C431 VTAIL.n160 VSUBS 0.014793f
C432 VTAIL.n161 VSUBS 0.015664f
C433 VTAIL.n162 VSUBS 0.034966f
C434 VTAIL.n163 VSUBS 0.034966f
C435 VTAIL.n164 VSUBS 0.015664f
C436 VTAIL.n165 VSUBS 0.014793f
C437 VTAIL.n166 VSUBS 0.02753f
C438 VTAIL.n167 VSUBS 0.02753f
C439 VTAIL.n168 VSUBS 0.014793f
C440 VTAIL.n169 VSUBS 0.015664f
C441 VTAIL.n170 VSUBS 0.034966f
C442 VTAIL.n171 VSUBS 0.034966f
C443 VTAIL.n172 VSUBS 0.015664f
C444 VTAIL.n173 VSUBS 0.014793f
C445 VTAIL.n174 VSUBS 0.02753f
C446 VTAIL.n175 VSUBS 0.02753f
C447 VTAIL.n176 VSUBS 0.014793f
C448 VTAIL.n177 VSUBS 0.015229f
C449 VTAIL.n178 VSUBS 0.015229f
C450 VTAIL.n179 VSUBS 0.034966f
C451 VTAIL.n180 VSUBS 0.034966f
C452 VTAIL.n181 VSUBS 0.015664f
C453 VTAIL.n182 VSUBS 0.014793f
C454 VTAIL.n183 VSUBS 0.02753f
C455 VTAIL.n184 VSUBS 0.02753f
C456 VTAIL.n185 VSUBS 0.014793f
C457 VTAIL.n186 VSUBS 0.015664f
C458 VTAIL.n187 VSUBS 0.034966f
C459 VTAIL.n188 VSUBS 0.080282f
C460 VTAIL.n189 VSUBS 0.015664f
C461 VTAIL.n190 VSUBS 0.014793f
C462 VTAIL.n191 VSUBS 0.062882f
C463 VTAIL.n192 VSUBS 0.040156f
C464 VTAIL.n193 VSUBS 0.322858f
C465 VTAIL.t5 VSUBS 0.365048f
C466 VTAIL.t2 VSUBS 0.365048f
C467 VTAIL.n194 VSUBS 2.83319f
C468 VTAIL.n195 VSUBS 0.972703f
C469 VTAIL.n196 VSUBS 0.028967f
C470 VTAIL.n197 VSUBS 0.02753f
C471 VTAIL.n198 VSUBS 0.014793f
C472 VTAIL.n199 VSUBS 0.034966f
C473 VTAIL.n200 VSUBS 0.015664f
C474 VTAIL.n201 VSUBS 0.02753f
C475 VTAIL.n202 VSUBS 0.014793f
C476 VTAIL.n203 VSUBS 0.034966f
C477 VTAIL.n204 VSUBS 0.015664f
C478 VTAIL.n205 VSUBS 0.02753f
C479 VTAIL.n206 VSUBS 0.014793f
C480 VTAIL.n207 VSUBS 0.034966f
C481 VTAIL.n208 VSUBS 0.034966f
C482 VTAIL.n209 VSUBS 0.015664f
C483 VTAIL.n210 VSUBS 0.02753f
C484 VTAIL.n211 VSUBS 0.014793f
C485 VTAIL.n212 VSUBS 0.034966f
C486 VTAIL.n213 VSUBS 0.015664f
C487 VTAIL.n214 VSUBS 0.02753f
C488 VTAIL.n215 VSUBS 0.014793f
C489 VTAIL.n216 VSUBS 0.034966f
C490 VTAIL.n217 VSUBS 0.015664f
C491 VTAIL.n218 VSUBS 0.02753f
C492 VTAIL.n219 VSUBS 0.014793f
C493 VTAIL.n220 VSUBS 0.034966f
C494 VTAIL.n221 VSUBS 0.015664f
C495 VTAIL.n222 VSUBS 0.02753f
C496 VTAIL.n223 VSUBS 0.014793f
C497 VTAIL.n224 VSUBS 0.034966f
C498 VTAIL.n225 VSUBS 0.015664f
C499 VTAIL.n226 VSUBS 0.208515f
C500 VTAIL.t1 VSUBS 0.074977f
C501 VTAIL.n227 VSUBS 0.026225f
C502 VTAIL.n228 VSUBS 0.022244f
C503 VTAIL.n229 VSUBS 0.014793f
C504 VTAIL.n230 VSUBS 1.9803f
C505 VTAIL.n231 VSUBS 0.02753f
C506 VTAIL.n232 VSUBS 0.014793f
C507 VTAIL.n233 VSUBS 0.015664f
C508 VTAIL.n234 VSUBS 0.034966f
C509 VTAIL.n235 VSUBS 0.034966f
C510 VTAIL.n236 VSUBS 0.015664f
C511 VTAIL.n237 VSUBS 0.014793f
C512 VTAIL.n238 VSUBS 0.02753f
C513 VTAIL.n239 VSUBS 0.02753f
C514 VTAIL.n240 VSUBS 0.014793f
C515 VTAIL.n241 VSUBS 0.015664f
C516 VTAIL.n242 VSUBS 0.034966f
C517 VTAIL.n243 VSUBS 0.034966f
C518 VTAIL.n244 VSUBS 0.015664f
C519 VTAIL.n245 VSUBS 0.014793f
C520 VTAIL.n246 VSUBS 0.02753f
C521 VTAIL.n247 VSUBS 0.02753f
C522 VTAIL.n248 VSUBS 0.014793f
C523 VTAIL.n249 VSUBS 0.015664f
C524 VTAIL.n250 VSUBS 0.034966f
C525 VTAIL.n251 VSUBS 0.034966f
C526 VTAIL.n252 VSUBS 0.015664f
C527 VTAIL.n253 VSUBS 0.014793f
C528 VTAIL.n254 VSUBS 0.02753f
C529 VTAIL.n255 VSUBS 0.02753f
C530 VTAIL.n256 VSUBS 0.014793f
C531 VTAIL.n257 VSUBS 0.015664f
C532 VTAIL.n258 VSUBS 0.034966f
C533 VTAIL.n259 VSUBS 0.034966f
C534 VTAIL.n260 VSUBS 0.015664f
C535 VTAIL.n261 VSUBS 0.014793f
C536 VTAIL.n262 VSUBS 0.02753f
C537 VTAIL.n263 VSUBS 0.02753f
C538 VTAIL.n264 VSUBS 0.014793f
C539 VTAIL.n265 VSUBS 0.015664f
C540 VTAIL.n266 VSUBS 0.034966f
C541 VTAIL.n267 VSUBS 0.034966f
C542 VTAIL.n268 VSUBS 0.015664f
C543 VTAIL.n269 VSUBS 0.014793f
C544 VTAIL.n270 VSUBS 0.02753f
C545 VTAIL.n271 VSUBS 0.02753f
C546 VTAIL.n272 VSUBS 0.014793f
C547 VTAIL.n273 VSUBS 0.015229f
C548 VTAIL.n274 VSUBS 0.015229f
C549 VTAIL.n275 VSUBS 0.034966f
C550 VTAIL.n276 VSUBS 0.034966f
C551 VTAIL.n277 VSUBS 0.015664f
C552 VTAIL.n278 VSUBS 0.014793f
C553 VTAIL.n279 VSUBS 0.02753f
C554 VTAIL.n280 VSUBS 0.02753f
C555 VTAIL.n281 VSUBS 0.014793f
C556 VTAIL.n282 VSUBS 0.015664f
C557 VTAIL.n283 VSUBS 0.034966f
C558 VTAIL.n284 VSUBS 0.080282f
C559 VTAIL.n285 VSUBS 0.015664f
C560 VTAIL.n286 VSUBS 0.014793f
C561 VTAIL.n287 VSUBS 0.062882f
C562 VTAIL.n288 VSUBS 0.040156f
C563 VTAIL.n289 VSUBS 2.02437f
C564 VTAIL.n290 VSUBS 0.028967f
C565 VTAIL.n291 VSUBS 0.02753f
C566 VTAIL.n292 VSUBS 0.014793f
C567 VTAIL.n293 VSUBS 0.034966f
C568 VTAIL.n294 VSUBS 0.015664f
C569 VTAIL.n295 VSUBS 0.02753f
C570 VTAIL.n296 VSUBS 0.014793f
C571 VTAIL.n297 VSUBS 0.034966f
C572 VTAIL.n298 VSUBS 0.015664f
C573 VTAIL.n299 VSUBS 0.02753f
C574 VTAIL.n300 VSUBS 0.014793f
C575 VTAIL.n301 VSUBS 0.034966f
C576 VTAIL.n302 VSUBS 0.015664f
C577 VTAIL.n303 VSUBS 0.02753f
C578 VTAIL.n304 VSUBS 0.014793f
C579 VTAIL.n305 VSUBS 0.034966f
C580 VTAIL.n306 VSUBS 0.015664f
C581 VTAIL.n307 VSUBS 0.02753f
C582 VTAIL.n308 VSUBS 0.014793f
C583 VTAIL.n309 VSUBS 0.034966f
C584 VTAIL.n310 VSUBS 0.015664f
C585 VTAIL.n311 VSUBS 0.02753f
C586 VTAIL.n312 VSUBS 0.014793f
C587 VTAIL.n313 VSUBS 0.034966f
C588 VTAIL.n314 VSUBS 0.015664f
C589 VTAIL.n315 VSUBS 0.02753f
C590 VTAIL.n316 VSUBS 0.014793f
C591 VTAIL.n317 VSUBS 0.034966f
C592 VTAIL.n318 VSUBS 0.015664f
C593 VTAIL.n319 VSUBS 0.208515f
C594 VTAIL.t7 VSUBS 0.074977f
C595 VTAIL.n320 VSUBS 0.026225f
C596 VTAIL.n321 VSUBS 0.022244f
C597 VTAIL.n322 VSUBS 0.014793f
C598 VTAIL.n323 VSUBS 1.9803f
C599 VTAIL.n324 VSUBS 0.02753f
C600 VTAIL.n325 VSUBS 0.014793f
C601 VTAIL.n326 VSUBS 0.015664f
C602 VTAIL.n327 VSUBS 0.034966f
C603 VTAIL.n328 VSUBS 0.034966f
C604 VTAIL.n329 VSUBS 0.015664f
C605 VTAIL.n330 VSUBS 0.014793f
C606 VTAIL.n331 VSUBS 0.02753f
C607 VTAIL.n332 VSUBS 0.02753f
C608 VTAIL.n333 VSUBS 0.014793f
C609 VTAIL.n334 VSUBS 0.015664f
C610 VTAIL.n335 VSUBS 0.034966f
C611 VTAIL.n336 VSUBS 0.034966f
C612 VTAIL.n337 VSUBS 0.015664f
C613 VTAIL.n338 VSUBS 0.014793f
C614 VTAIL.n339 VSUBS 0.02753f
C615 VTAIL.n340 VSUBS 0.02753f
C616 VTAIL.n341 VSUBS 0.014793f
C617 VTAIL.n342 VSUBS 0.015664f
C618 VTAIL.n343 VSUBS 0.034966f
C619 VTAIL.n344 VSUBS 0.034966f
C620 VTAIL.n345 VSUBS 0.015664f
C621 VTAIL.n346 VSUBS 0.014793f
C622 VTAIL.n347 VSUBS 0.02753f
C623 VTAIL.n348 VSUBS 0.02753f
C624 VTAIL.n349 VSUBS 0.014793f
C625 VTAIL.n350 VSUBS 0.015664f
C626 VTAIL.n351 VSUBS 0.034966f
C627 VTAIL.n352 VSUBS 0.034966f
C628 VTAIL.n353 VSUBS 0.015664f
C629 VTAIL.n354 VSUBS 0.014793f
C630 VTAIL.n355 VSUBS 0.02753f
C631 VTAIL.n356 VSUBS 0.02753f
C632 VTAIL.n357 VSUBS 0.014793f
C633 VTAIL.n358 VSUBS 0.015664f
C634 VTAIL.n359 VSUBS 0.034966f
C635 VTAIL.n360 VSUBS 0.034966f
C636 VTAIL.n361 VSUBS 0.034966f
C637 VTAIL.n362 VSUBS 0.015664f
C638 VTAIL.n363 VSUBS 0.014793f
C639 VTAIL.n364 VSUBS 0.02753f
C640 VTAIL.n365 VSUBS 0.02753f
C641 VTAIL.n366 VSUBS 0.014793f
C642 VTAIL.n367 VSUBS 0.015229f
C643 VTAIL.n368 VSUBS 0.015229f
C644 VTAIL.n369 VSUBS 0.034966f
C645 VTAIL.n370 VSUBS 0.034966f
C646 VTAIL.n371 VSUBS 0.015664f
C647 VTAIL.n372 VSUBS 0.014793f
C648 VTAIL.n373 VSUBS 0.02753f
C649 VTAIL.n374 VSUBS 0.02753f
C650 VTAIL.n375 VSUBS 0.014793f
C651 VTAIL.n376 VSUBS 0.015664f
C652 VTAIL.n377 VSUBS 0.034966f
C653 VTAIL.n378 VSUBS 0.080282f
C654 VTAIL.n379 VSUBS 0.015664f
C655 VTAIL.n380 VSUBS 0.014793f
C656 VTAIL.n381 VSUBS 0.062882f
C657 VTAIL.n382 VSUBS 0.040156f
C658 VTAIL.n383 VSUBS 1.97619f
C659 VDD2.n0 VSUBS 0.028493f
C660 VDD2.n1 VSUBS 0.027079f
C661 VDD2.n2 VSUBS 0.014551f
C662 VDD2.n3 VSUBS 0.034393f
C663 VDD2.n4 VSUBS 0.015407f
C664 VDD2.n5 VSUBS 0.027079f
C665 VDD2.n6 VSUBS 0.014551f
C666 VDD2.n7 VSUBS 0.034393f
C667 VDD2.n8 VSUBS 0.015407f
C668 VDD2.n9 VSUBS 0.027079f
C669 VDD2.n10 VSUBS 0.014551f
C670 VDD2.n11 VSUBS 0.034393f
C671 VDD2.n12 VSUBS 0.015407f
C672 VDD2.n13 VSUBS 0.027079f
C673 VDD2.n14 VSUBS 0.014551f
C674 VDD2.n15 VSUBS 0.034393f
C675 VDD2.n16 VSUBS 0.015407f
C676 VDD2.n17 VSUBS 0.027079f
C677 VDD2.n18 VSUBS 0.014551f
C678 VDD2.n19 VSUBS 0.034393f
C679 VDD2.n20 VSUBS 0.015407f
C680 VDD2.n21 VSUBS 0.027079f
C681 VDD2.n22 VSUBS 0.014551f
C682 VDD2.n23 VSUBS 0.034393f
C683 VDD2.n24 VSUBS 0.015407f
C684 VDD2.n25 VSUBS 0.027079f
C685 VDD2.n26 VSUBS 0.014551f
C686 VDD2.n27 VSUBS 0.034393f
C687 VDD2.n28 VSUBS 0.015407f
C688 VDD2.n29 VSUBS 0.205097f
C689 VDD2.t0 VSUBS 0.073748f
C690 VDD2.n30 VSUBS 0.025795f
C691 VDD2.n31 VSUBS 0.021879f
C692 VDD2.n32 VSUBS 0.014551f
C693 VDD2.n33 VSUBS 1.94784f
C694 VDD2.n34 VSUBS 0.027079f
C695 VDD2.n35 VSUBS 0.014551f
C696 VDD2.n36 VSUBS 0.015407f
C697 VDD2.n37 VSUBS 0.034393f
C698 VDD2.n38 VSUBS 0.034393f
C699 VDD2.n39 VSUBS 0.015407f
C700 VDD2.n40 VSUBS 0.014551f
C701 VDD2.n41 VSUBS 0.027079f
C702 VDD2.n42 VSUBS 0.027079f
C703 VDD2.n43 VSUBS 0.014551f
C704 VDD2.n44 VSUBS 0.015407f
C705 VDD2.n45 VSUBS 0.034393f
C706 VDD2.n46 VSUBS 0.034393f
C707 VDD2.n47 VSUBS 0.015407f
C708 VDD2.n48 VSUBS 0.014551f
C709 VDD2.n49 VSUBS 0.027079f
C710 VDD2.n50 VSUBS 0.027079f
C711 VDD2.n51 VSUBS 0.014551f
C712 VDD2.n52 VSUBS 0.015407f
C713 VDD2.n53 VSUBS 0.034393f
C714 VDD2.n54 VSUBS 0.034393f
C715 VDD2.n55 VSUBS 0.015407f
C716 VDD2.n56 VSUBS 0.014551f
C717 VDD2.n57 VSUBS 0.027079f
C718 VDD2.n58 VSUBS 0.027079f
C719 VDD2.n59 VSUBS 0.014551f
C720 VDD2.n60 VSUBS 0.015407f
C721 VDD2.n61 VSUBS 0.034393f
C722 VDD2.n62 VSUBS 0.034393f
C723 VDD2.n63 VSUBS 0.015407f
C724 VDD2.n64 VSUBS 0.014551f
C725 VDD2.n65 VSUBS 0.027079f
C726 VDD2.n66 VSUBS 0.027079f
C727 VDD2.n67 VSUBS 0.014551f
C728 VDD2.n68 VSUBS 0.015407f
C729 VDD2.n69 VSUBS 0.034393f
C730 VDD2.n70 VSUBS 0.034393f
C731 VDD2.n71 VSUBS 0.034393f
C732 VDD2.n72 VSUBS 0.015407f
C733 VDD2.n73 VSUBS 0.014551f
C734 VDD2.n74 VSUBS 0.027079f
C735 VDD2.n75 VSUBS 0.027079f
C736 VDD2.n76 VSUBS 0.014551f
C737 VDD2.n77 VSUBS 0.014979f
C738 VDD2.n78 VSUBS 0.014979f
C739 VDD2.n79 VSUBS 0.034393f
C740 VDD2.n80 VSUBS 0.034393f
C741 VDD2.n81 VSUBS 0.015407f
C742 VDD2.n82 VSUBS 0.014551f
C743 VDD2.n83 VSUBS 0.027079f
C744 VDD2.n84 VSUBS 0.027079f
C745 VDD2.n85 VSUBS 0.014551f
C746 VDD2.n86 VSUBS 0.015407f
C747 VDD2.n87 VSUBS 0.034393f
C748 VDD2.n88 VSUBS 0.078966f
C749 VDD2.n89 VSUBS 0.015407f
C750 VDD2.n90 VSUBS 0.014551f
C751 VDD2.n91 VSUBS 0.061851f
C752 VDD2.n92 VSUBS 0.06309f
C753 VDD2.t1 VSUBS 0.359064f
C754 VDD2.t2 VSUBS 0.359064f
C755 VDD2.n93 VSUBS 2.95901f
C756 VDD2.n94 VSUBS 3.20938f
C757 VDD2.n95 VSUBS 0.028493f
C758 VDD2.n96 VSUBS 0.027079f
C759 VDD2.n97 VSUBS 0.014551f
C760 VDD2.n98 VSUBS 0.034393f
C761 VDD2.n99 VSUBS 0.015407f
C762 VDD2.n100 VSUBS 0.027079f
C763 VDD2.n101 VSUBS 0.014551f
C764 VDD2.n102 VSUBS 0.034393f
C765 VDD2.n103 VSUBS 0.015407f
C766 VDD2.n104 VSUBS 0.027079f
C767 VDD2.n105 VSUBS 0.014551f
C768 VDD2.n106 VSUBS 0.034393f
C769 VDD2.n107 VSUBS 0.034393f
C770 VDD2.n108 VSUBS 0.015407f
C771 VDD2.n109 VSUBS 0.027079f
C772 VDD2.n110 VSUBS 0.014551f
C773 VDD2.n111 VSUBS 0.034393f
C774 VDD2.n112 VSUBS 0.015407f
C775 VDD2.n113 VSUBS 0.027079f
C776 VDD2.n114 VSUBS 0.014551f
C777 VDD2.n115 VSUBS 0.034393f
C778 VDD2.n116 VSUBS 0.015407f
C779 VDD2.n117 VSUBS 0.027079f
C780 VDD2.n118 VSUBS 0.014551f
C781 VDD2.n119 VSUBS 0.034393f
C782 VDD2.n120 VSUBS 0.015407f
C783 VDD2.n121 VSUBS 0.027079f
C784 VDD2.n122 VSUBS 0.014551f
C785 VDD2.n123 VSUBS 0.034393f
C786 VDD2.n124 VSUBS 0.015407f
C787 VDD2.n125 VSUBS 0.205097f
C788 VDD2.t5 VSUBS 0.073748f
C789 VDD2.n126 VSUBS 0.025795f
C790 VDD2.n127 VSUBS 0.021879f
C791 VDD2.n128 VSUBS 0.014551f
C792 VDD2.n129 VSUBS 1.94784f
C793 VDD2.n130 VSUBS 0.027079f
C794 VDD2.n131 VSUBS 0.014551f
C795 VDD2.n132 VSUBS 0.015407f
C796 VDD2.n133 VSUBS 0.034393f
C797 VDD2.n134 VSUBS 0.034393f
C798 VDD2.n135 VSUBS 0.015407f
C799 VDD2.n136 VSUBS 0.014551f
C800 VDD2.n137 VSUBS 0.027079f
C801 VDD2.n138 VSUBS 0.027079f
C802 VDD2.n139 VSUBS 0.014551f
C803 VDD2.n140 VSUBS 0.015407f
C804 VDD2.n141 VSUBS 0.034393f
C805 VDD2.n142 VSUBS 0.034393f
C806 VDD2.n143 VSUBS 0.015407f
C807 VDD2.n144 VSUBS 0.014551f
C808 VDD2.n145 VSUBS 0.027079f
C809 VDD2.n146 VSUBS 0.027079f
C810 VDD2.n147 VSUBS 0.014551f
C811 VDD2.n148 VSUBS 0.015407f
C812 VDD2.n149 VSUBS 0.034393f
C813 VDD2.n150 VSUBS 0.034393f
C814 VDD2.n151 VSUBS 0.015407f
C815 VDD2.n152 VSUBS 0.014551f
C816 VDD2.n153 VSUBS 0.027079f
C817 VDD2.n154 VSUBS 0.027079f
C818 VDD2.n155 VSUBS 0.014551f
C819 VDD2.n156 VSUBS 0.015407f
C820 VDD2.n157 VSUBS 0.034393f
C821 VDD2.n158 VSUBS 0.034393f
C822 VDD2.n159 VSUBS 0.015407f
C823 VDD2.n160 VSUBS 0.014551f
C824 VDD2.n161 VSUBS 0.027079f
C825 VDD2.n162 VSUBS 0.027079f
C826 VDD2.n163 VSUBS 0.014551f
C827 VDD2.n164 VSUBS 0.015407f
C828 VDD2.n165 VSUBS 0.034393f
C829 VDD2.n166 VSUBS 0.034393f
C830 VDD2.n167 VSUBS 0.015407f
C831 VDD2.n168 VSUBS 0.014551f
C832 VDD2.n169 VSUBS 0.027079f
C833 VDD2.n170 VSUBS 0.027079f
C834 VDD2.n171 VSUBS 0.014551f
C835 VDD2.n172 VSUBS 0.014979f
C836 VDD2.n173 VSUBS 0.014979f
C837 VDD2.n174 VSUBS 0.034393f
C838 VDD2.n175 VSUBS 0.034393f
C839 VDD2.n176 VSUBS 0.015407f
C840 VDD2.n177 VSUBS 0.014551f
C841 VDD2.n178 VSUBS 0.027079f
C842 VDD2.n179 VSUBS 0.027079f
C843 VDD2.n180 VSUBS 0.014551f
C844 VDD2.n181 VSUBS 0.015407f
C845 VDD2.n182 VSUBS 0.034393f
C846 VDD2.n183 VSUBS 0.078966f
C847 VDD2.n184 VSUBS 0.015407f
C848 VDD2.n185 VSUBS 0.014551f
C849 VDD2.n186 VSUBS 0.061851f
C850 VDD2.n187 VSUBS 0.058201f
C851 VDD2.n188 VSUBS 2.9706f
C852 VDD2.t4 VSUBS 0.359064f
C853 VDD2.t3 VSUBS 0.359064f
C854 VDD2.n189 VSUBS 2.95897f
C855 VN.n0 VSUBS 0.043943f
C856 VN.t4 VSUBS 2.94945f
C857 VN.n1 VSUBS 0.05978f
C858 VN.t2 VSUBS 3.10481f
C859 VN.n2 VSUBS 1.12253f
C860 VN.t0 VSUBS 2.94945f
C861 VN.n3 VSUBS 1.11205f
C862 VN.n4 VSUBS 0.047017f
C863 VN.n5 VSUBS 0.246895f
C864 VN.n6 VSUBS 0.033329f
C865 VN.n7 VSUBS 0.033329f
C866 VN.n8 VSUBS 0.034381f
C867 VN.n9 VSUBS 0.065999f
C868 VN.n10 VSUBS 1.14224f
C869 VN.n11 VSUBS 0.035224f
C870 VN.n12 VSUBS 0.043943f
C871 VN.t3 VSUBS 2.94945f
C872 VN.n13 VSUBS 0.05978f
C873 VN.t1 VSUBS 3.10481f
C874 VN.n14 VSUBS 1.12253f
C875 VN.t5 VSUBS 2.94945f
C876 VN.n15 VSUBS 1.11205f
C877 VN.n16 VSUBS 0.047017f
C878 VN.n17 VSUBS 0.246895f
C879 VN.n18 VSUBS 0.033329f
C880 VN.n19 VSUBS 0.033329f
C881 VN.n20 VSUBS 0.034381f
C882 VN.n21 VSUBS 0.065999f
C883 VN.n22 VSUBS 1.14224f
C884 VN.n23 VSUBS 1.83728f
C885 B.n0 VSUBS 0.006877f
C886 B.n1 VSUBS 0.006877f
C887 B.n2 VSUBS 0.010171f
C888 B.n3 VSUBS 0.007794f
C889 B.n4 VSUBS 0.007794f
C890 B.n5 VSUBS 0.007794f
C891 B.n6 VSUBS 0.007794f
C892 B.n7 VSUBS 0.007794f
C893 B.n8 VSUBS 0.007794f
C894 B.n9 VSUBS 0.007794f
C895 B.n10 VSUBS 0.007794f
C896 B.n11 VSUBS 0.007794f
C897 B.n12 VSUBS 0.007794f
C898 B.n13 VSUBS 0.007794f
C899 B.n14 VSUBS 0.007794f
C900 B.n15 VSUBS 0.007794f
C901 B.n16 VSUBS 0.007794f
C902 B.n17 VSUBS 0.007794f
C903 B.n18 VSUBS 0.007794f
C904 B.n19 VSUBS 0.018863f
C905 B.n20 VSUBS 0.007794f
C906 B.n21 VSUBS 0.007794f
C907 B.n22 VSUBS 0.007794f
C908 B.n23 VSUBS 0.007794f
C909 B.n24 VSUBS 0.007794f
C910 B.n25 VSUBS 0.007794f
C911 B.n26 VSUBS 0.007794f
C912 B.n27 VSUBS 0.007794f
C913 B.n28 VSUBS 0.007794f
C914 B.n29 VSUBS 0.007794f
C915 B.n30 VSUBS 0.007794f
C916 B.n31 VSUBS 0.007794f
C917 B.n32 VSUBS 0.007794f
C918 B.n33 VSUBS 0.007794f
C919 B.n34 VSUBS 0.007794f
C920 B.n35 VSUBS 0.007794f
C921 B.n36 VSUBS 0.007794f
C922 B.n37 VSUBS 0.007794f
C923 B.n38 VSUBS 0.007794f
C924 B.n39 VSUBS 0.007794f
C925 B.n40 VSUBS 0.007794f
C926 B.n41 VSUBS 0.007794f
C927 B.n42 VSUBS 0.007794f
C928 B.n43 VSUBS 0.007794f
C929 B.n44 VSUBS 0.007794f
C930 B.n45 VSUBS 0.007794f
C931 B.n46 VSUBS 0.007794f
C932 B.n47 VSUBS 0.007794f
C933 B.t7 VSUBS 0.358158f
C934 B.t8 VSUBS 0.387123f
C935 B.t6 VSUBS 1.56255f
C936 B.n48 VSUBS 0.572113f
C937 B.n49 VSUBS 0.346514f
C938 B.n50 VSUBS 0.007794f
C939 B.n51 VSUBS 0.007794f
C940 B.n52 VSUBS 0.007794f
C941 B.n53 VSUBS 0.007794f
C942 B.t4 VSUBS 0.358162f
C943 B.t5 VSUBS 0.387126f
C944 B.t3 VSUBS 1.56255f
C945 B.n54 VSUBS 0.57211f
C946 B.n55 VSUBS 0.34651f
C947 B.n56 VSUBS 0.007794f
C948 B.n57 VSUBS 0.007794f
C949 B.n58 VSUBS 0.007794f
C950 B.n59 VSUBS 0.007794f
C951 B.n60 VSUBS 0.007794f
C952 B.n61 VSUBS 0.007794f
C953 B.n62 VSUBS 0.007794f
C954 B.n63 VSUBS 0.007794f
C955 B.n64 VSUBS 0.007794f
C956 B.n65 VSUBS 0.007794f
C957 B.n66 VSUBS 0.007794f
C958 B.n67 VSUBS 0.007794f
C959 B.n68 VSUBS 0.007794f
C960 B.n69 VSUBS 0.007794f
C961 B.n70 VSUBS 0.007794f
C962 B.n71 VSUBS 0.007794f
C963 B.n72 VSUBS 0.007794f
C964 B.n73 VSUBS 0.007794f
C965 B.n74 VSUBS 0.007794f
C966 B.n75 VSUBS 0.007794f
C967 B.n76 VSUBS 0.007794f
C968 B.n77 VSUBS 0.007794f
C969 B.n78 VSUBS 0.007794f
C970 B.n79 VSUBS 0.007794f
C971 B.n80 VSUBS 0.007794f
C972 B.n81 VSUBS 0.007794f
C973 B.n82 VSUBS 0.007794f
C974 B.n83 VSUBS 0.018863f
C975 B.n84 VSUBS 0.007794f
C976 B.n85 VSUBS 0.007794f
C977 B.n86 VSUBS 0.007794f
C978 B.n87 VSUBS 0.007794f
C979 B.n88 VSUBS 0.007794f
C980 B.n89 VSUBS 0.007794f
C981 B.n90 VSUBS 0.007794f
C982 B.n91 VSUBS 0.007794f
C983 B.n92 VSUBS 0.007794f
C984 B.n93 VSUBS 0.007794f
C985 B.n94 VSUBS 0.007794f
C986 B.n95 VSUBS 0.007794f
C987 B.n96 VSUBS 0.007794f
C988 B.n97 VSUBS 0.007794f
C989 B.n98 VSUBS 0.007794f
C990 B.n99 VSUBS 0.007794f
C991 B.n100 VSUBS 0.007794f
C992 B.n101 VSUBS 0.007794f
C993 B.n102 VSUBS 0.007794f
C994 B.n103 VSUBS 0.007794f
C995 B.n104 VSUBS 0.007794f
C996 B.n105 VSUBS 0.007794f
C997 B.n106 VSUBS 0.007794f
C998 B.n107 VSUBS 0.007794f
C999 B.n108 VSUBS 0.007794f
C1000 B.n109 VSUBS 0.007794f
C1001 B.n110 VSUBS 0.007794f
C1002 B.n111 VSUBS 0.007794f
C1003 B.n112 VSUBS 0.007794f
C1004 B.n113 VSUBS 0.007794f
C1005 B.n114 VSUBS 0.007794f
C1006 B.n115 VSUBS 0.007794f
C1007 B.n116 VSUBS 0.007794f
C1008 B.n117 VSUBS 0.007794f
C1009 B.n118 VSUBS 0.018729f
C1010 B.n119 VSUBS 0.007794f
C1011 B.n120 VSUBS 0.007794f
C1012 B.n121 VSUBS 0.007794f
C1013 B.n122 VSUBS 0.007794f
C1014 B.n123 VSUBS 0.007794f
C1015 B.n124 VSUBS 0.007794f
C1016 B.n125 VSUBS 0.007794f
C1017 B.n126 VSUBS 0.007794f
C1018 B.n127 VSUBS 0.007794f
C1019 B.n128 VSUBS 0.007794f
C1020 B.n129 VSUBS 0.007794f
C1021 B.n130 VSUBS 0.007794f
C1022 B.n131 VSUBS 0.007794f
C1023 B.n132 VSUBS 0.007794f
C1024 B.n133 VSUBS 0.007794f
C1025 B.n134 VSUBS 0.007794f
C1026 B.n135 VSUBS 0.007794f
C1027 B.n136 VSUBS 0.007794f
C1028 B.n137 VSUBS 0.007794f
C1029 B.n138 VSUBS 0.007794f
C1030 B.n139 VSUBS 0.007794f
C1031 B.n140 VSUBS 0.007794f
C1032 B.n141 VSUBS 0.007794f
C1033 B.n142 VSUBS 0.007794f
C1034 B.n143 VSUBS 0.007794f
C1035 B.n144 VSUBS 0.007794f
C1036 B.n145 VSUBS 0.007794f
C1037 B.n146 VSUBS 0.005387f
C1038 B.n147 VSUBS 0.007794f
C1039 B.n148 VSUBS 0.007794f
C1040 B.n149 VSUBS 0.007794f
C1041 B.n150 VSUBS 0.007794f
C1042 B.n151 VSUBS 0.007794f
C1043 B.t2 VSUBS 0.358158f
C1044 B.t1 VSUBS 0.387123f
C1045 B.t0 VSUBS 1.56255f
C1046 B.n152 VSUBS 0.572113f
C1047 B.n153 VSUBS 0.346514f
C1048 B.n154 VSUBS 0.007794f
C1049 B.n155 VSUBS 0.007794f
C1050 B.n156 VSUBS 0.007794f
C1051 B.n157 VSUBS 0.007794f
C1052 B.n158 VSUBS 0.007794f
C1053 B.n159 VSUBS 0.007794f
C1054 B.n160 VSUBS 0.007794f
C1055 B.n161 VSUBS 0.007794f
C1056 B.n162 VSUBS 0.007794f
C1057 B.n163 VSUBS 0.007794f
C1058 B.n164 VSUBS 0.007794f
C1059 B.n165 VSUBS 0.007794f
C1060 B.n166 VSUBS 0.007794f
C1061 B.n167 VSUBS 0.007794f
C1062 B.n168 VSUBS 0.007794f
C1063 B.n169 VSUBS 0.007794f
C1064 B.n170 VSUBS 0.007794f
C1065 B.n171 VSUBS 0.007794f
C1066 B.n172 VSUBS 0.007794f
C1067 B.n173 VSUBS 0.007794f
C1068 B.n174 VSUBS 0.007794f
C1069 B.n175 VSUBS 0.007794f
C1070 B.n176 VSUBS 0.007794f
C1071 B.n177 VSUBS 0.007794f
C1072 B.n178 VSUBS 0.007794f
C1073 B.n179 VSUBS 0.007794f
C1074 B.n180 VSUBS 0.007794f
C1075 B.n181 VSUBS 0.017816f
C1076 B.n182 VSUBS 0.007794f
C1077 B.n183 VSUBS 0.007794f
C1078 B.n184 VSUBS 0.007794f
C1079 B.n185 VSUBS 0.007794f
C1080 B.n186 VSUBS 0.007794f
C1081 B.n187 VSUBS 0.007794f
C1082 B.n188 VSUBS 0.007794f
C1083 B.n189 VSUBS 0.007794f
C1084 B.n190 VSUBS 0.007794f
C1085 B.n191 VSUBS 0.007794f
C1086 B.n192 VSUBS 0.007794f
C1087 B.n193 VSUBS 0.007794f
C1088 B.n194 VSUBS 0.007794f
C1089 B.n195 VSUBS 0.007794f
C1090 B.n196 VSUBS 0.007794f
C1091 B.n197 VSUBS 0.007794f
C1092 B.n198 VSUBS 0.007794f
C1093 B.n199 VSUBS 0.007794f
C1094 B.n200 VSUBS 0.007794f
C1095 B.n201 VSUBS 0.007794f
C1096 B.n202 VSUBS 0.007794f
C1097 B.n203 VSUBS 0.007794f
C1098 B.n204 VSUBS 0.007794f
C1099 B.n205 VSUBS 0.007794f
C1100 B.n206 VSUBS 0.007794f
C1101 B.n207 VSUBS 0.007794f
C1102 B.n208 VSUBS 0.007794f
C1103 B.n209 VSUBS 0.007794f
C1104 B.n210 VSUBS 0.007794f
C1105 B.n211 VSUBS 0.007794f
C1106 B.n212 VSUBS 0.007794f
C1107 B.n213 VSUBS 0.007794f
C1108 B.n214 VSUBS 0.007794f
C1109 B.n215 VSUBS 0.007794f
C1110 B.n216 VSUBS 0.007794f
C1111 B.n217 VSUBS 0.007794f
C1112 B.n218 VSUBS 0.007794f
C1113 B.n219 VSUBS 0.007794f
C1114 B.n220 VSUBS 0.007794f
C1115 B.n221 VSUBS 0.007794f
C1116 B.n222 VSUBS 0.007794f
C1117 B.n223 VSUBS 0.007794f
C1118 B.n224 VSUBS 0.007794f
C1119 B.n225 VSUBS 0.007794f
C1120 B.n226 VSUBS 0.007794f
C1121 B.n227 VSUBS 0.007794f
C1122 B.n228 VSUBS 0.007794f
C1123 B.n229 VSUBS 0.007794f
C1124 B.n230 VSUBS 0.007794f
C1125 B.n231 VSUBS 0.007794f
C1126 B.n232 VSUBS 0.007794f
C1127 B.n233 VSUBS 0.007794f
C1128 B.n234 VSUBS 0.007794f
C1129 B.n235 VSUBS 0.007794f
C1130 B.n236 VSUBS 0.007794f
C1131 B.n237 VSUBS 0.007794f
C1132 B.n238 VSUBS 0.007794f
C1133 B.n239 VSUBS 0.007794f
C1134 B.n240 VSUBS 0.007794f
C1135 B.n241 VSUBS 0.007794f
C1136 B.n242 VSUBS 0.007794f
C1137 B.n243 VSUBS 0.007794f
C1138 B.n244 VSUBS 0.007794f
C1139 B.n245 VSUBS 0.007794f
C1140 B.n246 VSUBS 0.017816f
C1141 B.n247 VSUBS 0.018863f
C1142 B.n248 VSUBS 0.018863f
C1143 B.n249 VSUBS 0.007794f
C1144 B.n250 VSUBS 0.007794f
C1145 B.n251 VSUBS 0.007794f
C1146 B.n252 VSUBS 0.007794f
C1147 B.n253 VSUBS 0.007794f
C1148 B.n254 VSUBS 0.007794f
C1149 B.n255 VSUBS 0.007794f
C1150 B.n256 VSUBS 0.007794f
C1151 B.n257 VSUBS 0.007794f
C1152 B.n258 VSUBS 0.007794f
C1153 B.n259 VSUBS 0.007794f
C1154 B.n260 VSUBS 0.007794f
C1155 B.n261 VSUBS 0.007794f
C1156 B.n262 VSUBS 0.007794f
C1157 B.n263 VSUBS 0.007794f
C1158 B.n264 VSUBS 0.007794f
C1159 B.n265 VSUBS 0.007794f
C1160 B.n266 VSUBS 0.007794f
C1161 B.n267 VSUBS 0.007794f
C1162 B.n268 VSUBS 0.007794f
C1163 B.n269 VSUBS 0.007794f
C1164 B.n270 VSUBS 0.007794f
C1165 B.n271 VSUBS 0.007794f
C1166 B.n272 VSUBS 0.007794f
C1167 B.n273 VSUBS 0.007794f
C1168 B.n274 VSUBS 0.007794f
C1169 B.n275 VSUBS 0.007794f
C1170 B.n276 VSUBS 0.007794f
C1171 B.n277 VSUBS 0.007794f
C1172 B.n278 VSUBS 0.007794f
C1173 B.n279 VSUBS 0.007794f
C1174 B.n280 VSUBS 0.007794f
C1175 B.n281 VSUBS 0.007794f
C1176 B.n282 VSUBS 0.007794f
C1177 B.n283 VSUBS 0.007794f
C1178 B.n284 VSUBS 0.007794f
C1179 B.n285 VSUBS 0.007794f
C1180 B.n286 VSUBS 0.007794f
C1181 B.n287 VSUBS 0.007794f
C1182 B.n288 VSUBS 0.007794f
C1183 B.n289 VSUBS 0.007794f
C1184 B.n290 VSUBS 0.007794f
C1185 B.n291 VSUBS 0.007794f
C1186 B.n292 VSUBS 0.007794f
C1187 B.n293 VSUBS 0.007794f
C1188 B.n294 VSUBS 0.007794f
C1189 B.n295 VSUBS 0.007794f
C1190 B.n296 VSUBS 0.007794f
C1191 B.n297 VSUBS 0.007794f
C1192 B.n298 VSUBS 0.007794f
C1193 B.n299 VSUBS 0.007794f
C1194 B.n300 VSUBS 0.007794f
C1195 B.n301 VSUBS 0.007794f
C1196 B.n302 VSUBS 0.007794f
C1197 B.n303 VSUBS 0.007794f
C1198 B.n304 VSUBS 0.007794f
C1199 B.n305 VSUBS 0.007794f
C1200 B.n306 VSUBS 0.007794f
C1201 B.n307 VSUBS 0.007794f
C1202 B.n308 VSUBS 0.007794f
C1203 B.n309 VSUBS 0.007794f
C1204 B.n310 VSUBS 0.007794f
C1205 B.n311 VSUBS 0.007794f
C1206 B.n312 VSUBS 0.007794f
C1207 B.n313 VSUBS 0.007794f
C1208 B.n314 VSUBS 0.007794f
C1209 B.n315 VSUBS 0.007794f
C1210 B.n316 VSUBS 0.007794f
C1211 B.n317 VSUBS 0.007794f
C1212 B.n318 VSUBS 0.007794f
C1213 B.n319 VSUBS 0.007794f
C1214 B.n320 VSUBS 0.007794f
C1215 B.n321 VSUBS 0.007794f
C1216 B.n322 VSUBS 0.007794f
C1217 B.n323 VSUBS 0.007794f
C1218 B.n324 VSUBS 0.007794f
C1219 B.n325 VSUBS 0.007794f
C1220 B.n326 VSUBS 0.007794f
C1221 B.n327 VSUBS 0.007794f
C1222 B.n328 VSUBS 0.007794f
C1223 B.n329 VSUBS 0.007794f
C1224 B.n330 VSUBS 0.005387f
C1225 B.n331 VSUBS 0.018059f
C1226 B.n332 VSUBS 0.006304f
C1227 B.n333 VSUBS 0.007794f
C1228 B.n334 VSUBS 0.007794f
C1229 B.n335 VSUBS 0.007794f
C1230 B.n336 VSUBS 0.007794f
C1231 B.n337 VSUBS 0.007794f
C1232 B.n338 VSUBS 0.007794f
C1233 B.n339 VSUBS 0.007794f
C1234 B.n340 VSUBS 0.007794f
C1235 B.n341 VSUBS 0.007794f
C1236 B.n342 VSUBS 0.007794f
C1237 B.n343 VSUBS 0.007794f
C1238 B.t11 VSUBS 0.358162f
C1239 B.t10 VSUBS 0.387126f
C1240 B.t9 VSUBS 1.56255f
C1241 B.n344 VSUBS 0.57211f
C1242 B.n345 VSUBS 0.34651f
C1243 B.n346 VSUBS 0.018059f
C1244 B.n347 VSUBS 0.006304f
C1245 B.n348 VSUBS 0.007794f
C1246 B.n349 VSUBS 0.007794f
C1247 B.n350 VSUBS 0.007794f
C1248 B.n351 VSUBS 0.007794f
C1249 B.n352 VSUBS 0.007794f
C1250 B.n353 VSUBS 0.007794f
C1251 B.n354 VSUBS 0.007794f
C1252 B.n355 VSUBS 0.007794f
C1253 B.n356 VSUBS 0.007794f
C1254 B.n357 VSUBS 0.007794f
C1255 B.n358 VSUBS 0.007794f
C1256 B.n359 VSUBS 0.007794f
C1257 B.n360 VSUBS 0.007794f
C1258 B.n361 VSUBS 0.007794f
C1259 B.n362 VSUBS 0.007794f
C1260 B.n363 VSUBS 0.007794f
C1261 B.n364 VSUBS 0.007794f
C1262 B.n365 VSUBS 0.007794f
C1263 B.n366 VSUBS 0.007794f
C1264 B.n367 VSUBS 0.007794f
C1265 B.n368 VSUBS 0.007794f
C1266 B.n369 VSUBS 0.007794f
C1267 B.n370 VSUBS 0.007794f
C1268 B.n371 VSUBS 0.007794f
C1269 B.n372 VSUBS 0.007794f
C1270 B.n373 VSUBS 0.007794f
C1271 B.n374 VSUBS 0.007794f
C1272 B.n375 VSUBS 0.007794f
C1273 B.n376 VSUBS 0.007794f
C1274 B.n377 VSUBS 0.007794f
C1275 B.n378 VSUBS 0.007794f
C1276 B.n379 VSUBS 0.007794f
C1277 B.n380 VSUBS 0.007794f
C1278 B.n381 VSUBS 0.007794f
C1279 B.n382 VSUBS 0.007794f
C1280 B.n383 VSUBS 0.007794f
C1281 B.n384 VSUBS 0.007794f
C1282 B.n385 VSUBS 0.007794f
C1283 B.n386 VSUBS 0.007794f
C1284 B.n387 VSUBS 0.007794f
C1285 B.n388 VSUBS 0.007794f
C1286 B.n389 VSUBS 0.007794f
C1287 B.n390 VSUBS 0.007794f
C1288 B.n391 VSUBS 0.007794f
C1289 B.n392 VSUBS 0.007794f
C1290 B.n393 VSUBS 0.007794f
C1291 B.n394 VSUBS 0.007794f
C1292 B.n395 VSUBS 0.007794f
C1293 B.n396 VSUBS 0.007794f
C1294 B.n397 VSUBS 0.007794f
C1295 B.n398 VSUBS 0.007794f
C1296 B.n399 VSUBS 0.007794f
C1297 B.n400 VSUBS 0.007794f
C1298 B.n401 VSUBS 0.007794f
C1299 B.n402 VSUBS 0.007794f
C1300 B.n403 VSUBS 0.007794f
C1301 B.n404 VSUBS 0.007794f
C1302 B.n405 VSUBS 0.007794f
C1303 B.n406 VSUBS 0.007794f
C1304 B.n407 VSUBS 0.007794f
C1305 B.n408 VSUBS 0.007794f
C1306 B.n409 VSUBS 0.007794f
C1307 B.n410 VSUBS 0.007794f
C1308 B.n411 VSUBS 0.007794f
C1309 B.n412 VSUBS 0.007794f
C1310 B.n413 VSUBS 0.007794f
C1311 B.n414 VSUBS 0.007794f
C1312 B.n415 VSUBS 0.007794f
C1313 B.n416 VSUBS 0.007794f
C1314 B.n417 VSUBS 0.007794f
C1315 B.n418 VSUBS 0.007794f
C1316 B.n419 VSUBS 0.007794f
C1317 B.n420 VSUBS 0.007794f
C1318 B.n421 VSUBS 0.007794f
C1319 B.n422 VSUBS 0.007794f
C1320 B.n423 VSUBS 0.007794f
C1321 B.n424 VSUBS 0.007794f
C1322 B.n425 VSUBS 0.007794f
C1323 B.n426 VSUBS 0.007794f
C1324 B.n427 VSUBS 0.007794f
C1325 B.n428 VSUBS 0.007794f
C1326 B.n429 VSUBS 0.007794f
C1327 B.n430 VSUBS 0.007794f
C1328 B.n431 VSUBS 0.01795f
C1329 B.n432 VSUBS 0.018863f
C1330 B.n433 VSUBS 0.017816f
C1331 B.n434 VSUBS 0.007794f
C1332 B.n435 VSUBS 0.007794f
C1333 B.n436 VSUBS 0.007794f
C1334 B.n437 VSUBS 0.007794f
C1335 B.n438 VSUBS 0.007794f
C1336 B.n439 VSUBS 0.007794f
C1337 B.n440 VSUBS 0.007794f
C1338 B.n441 VSUBS 0.007794f
C1339 B.n442 VSUBS 0.007794f
C1340 B.n443 VSUBS 0.007794f
C1341 B.n444 VSUBS 0.007794f
C1342 B.n445 VSUBS 0.007794f
C1343 B.n446 VSUBS 0.007794f
C1344 B.n447 VSUBS 0.007794f
C1345 B.n448 VSUBS 0.007794f
C1346 B.n449 VSUBS 0.007794f
C1347 B.n450 VSUBS 0.007794f
C1348 B.n451 VSUBS 0.007794f
C1349 B.n452 VSUBS 0.007794f
C1350 B.n453 VSUBS 0.007794f
C1351 B.n454 VSUBS 0.007794f
C1352 B.n455 VSUBS 0.007794f
C1353 B.n456 VSUBS 0.007794f
C1354 B.n457 VSUBS 0.007794f
C1355 B.n458 VSUBS 0.007794f
C1356 B.n459 VSUBS 0.007794f
C1357 B.n460 VSUBS 0.007794f
C1358 B.n461 VSUBS 0.007794f
C1359 B.n462 VSUBS 0.007794f
C1360 B.n463 VSUBS 0.007794f
C1361 B.n464 VSUBS 0.007794f
C1362 B.n465 VSUBS 0.007794f
C1363 B.n466 VSUBS 0.007794f
C1364 B.n467 VSUBS 0.007794f
C1365 B.n468 VSUBS 0.007794f
C1366 B.n469 VSUBS 0.007794f
C1367 B.n470 VSUBS 0.007794f
C1368 B.n471 VSUBS 0.007794f
C1369 B.n472 VSUBS 0.007794f
C1370 B.n473 VSUBS 0.007794f
C1371 B.n474 VSUBS 0.007794f
C1372 B.n475 VSUBS 0.007794f
C1373 B.n476 VSUBS 0.007794f
C1374 B.n477 VSUBS 0.007794f
C1375 B.n478 VSUBS 0.007794f
C1376 B.n479 VSUBS 0.007794f
C1377 B.n480 VSUBS 0.007794f
C1378 B.n481 VSUBS 0.007794f
C1379 B.n482 VSUBS 0.007794f
C1380 B.n483 VSUBS 0.007794f
C1381 B.n484 VSUBS 0.007794f
C1382 B.n485 VSUBS 0.007794f
C1383 B.n486 VSUBS 0.007794f
C1384 B.n487 VSUBS 0.007794f
C1385 B.n488 VSUBS 0.007794f
C1386 B.n489 VSUBS 0.007794f
C1387 B.n490 VSUBS 0.007794f
C1388 B.n491 VSUBS 0.007794f
C1389 B.n492 VSUBS 0.007794f
C1390 B.n493 VSUBS 0.007794f
C1391 B.n494 VSUBS 0.007794f
C1392 B.n495 VSUBS 0.007794f
C1393 B.n496 VSUBS 0.007794f
C1394 B.n497 VSUBS 0.007794f
C1395 B.n498 VSUBS 0.007794f
C1396 B.n499 VSUBS 0.007794f
C1397 B.n500 VSUBS 0.007794f
C1398 B.n501 VSUBS 0.007794f
C1399 B.n502 VSUBS 0.007794f
C1400 B.n503 VSUBS 0.007794f
C1401 B.n504 VSUBS 0.007794f
C1402 B.n505 VSUBS 0.007794f
C1403 B.n506 VSUBS 0.007794f
C1404 B.n507 VSUBS 0.007794f
C1405 B.n508 VSUBS 0.007794f
C1406 B.n509 VSUBS 0.007794f
C1407 B.n510 VSUBS 0.007794f
C1408 B.n511 VSUBS 0.007794f
C1409 B.n512 VSUBS 0.007794f
C1410 B.n513 VSUBS 0.007794f
C1411 B.n514 VSUBS 0.007794f
C1412 B.n515 VSUBS 0.007794f
C1413 B.n516 VSUBS 0.007794f
C1414 B.n517 VSUBS 0.007794f
C1415 B.n518 VSUBS 0.007794f
C1416 B.n519 VSUBS 0.007794f
C1417 B.n520 VSUBS 0.007794f
C1418 B.n521 VSUBS 0.007794f
C1419 B.n522 VSUBS 0.007794f
C1420 B.n523 VSUBS 0.007794f
C1421 B.n524 VSUBS 0.007794f
C1422 B.n525 VSUBS 0.007794f
C1423 B.n526 VSUBS 0.007794f
C1424 B.n527 VSUBS 0.007794f
C1425 B.n528 VSUBS 0.007794f
C1426 B.n529 VSUBS 0.007794f
C1427 B.n530 VSUBS 0.007794f
C1428 B.n531 VSUBS 0.007794f
C1429 B.n532 VSUBS 0.007794f
C1430 B.n533 VSUBS 0.007794f
C1431 B.n534 VSUBS 0.007794f
C1432 B.n535 VSUBS 0.007794f
C1433 B.n536 VSUBS 0.017816f
C1434 B.n537 VSUBS 0.017816f
C1435 B.n538 VSUBS 0.018863f
C1436 B.n539 VSUBS 0.007794f
C1437 B.n540 VSUBS 0.007794f
C1438 B.n541 VSUBS 0.007794f
C1439 B.n542 VSUBS 0.007794f
C1440 B.n543 VSUBS 0.007794f
C1441 B.n544 VSUBS 0.007794f
C1442 B.n545 VSUBS 0.007794f
C1443 B.n546 VSUBS 0.007794f
C1444 B.n547 VSUBS 0.007794f
C1445 B.n548 VSUBS 0.007794f
C1446 B.n549 VSUBS 0.007794f
C1447 B.n550 VSUBS 0.007794f
C1448 B.n551 VSUBS 0.007794f
C1449 B.n552 VSUBS 0.007794f
C1450 B.n553 VSUBS 0.007794f
C1451 B.n554 VSUBS 0.007794f
C1452 B.n555 VSUBS 0.007794f
C1453 B.n556 VSUBS 0.007794f
C1454 B.n557 VSUBS 0.007794f
C1455 B.n558 VSUBS 0.007794f
C1456 B.n559 VSUBS 0.007794f
C1457 B.n560 VSUBS 0.007794f
C1458 B.n561 VSUBS 0.007794f
C1459 B.n562 VSUBS 0.007794f
C1460 B.n563 VSUBS 0.007794f
C1461 B.n564 VSUBS 0.007794f
C1462 B.n565 VSUBS 0.007794f
C1463 B.n566 VSUBS 0.007794f
C1464 B.n567 VSUBS 0.007794f
C1465 B.n568 VSUBS 0.007794f
C1466 B.n569 VSUBS 0.007794f
C1467 B.n570 VSUBS 0.007794f
C1468 B.n571 VSUBS 0.007794f
C1469 B.n572 VSUBS 0.007794f
C1470 B.n573 VSUBS 0.007794f
C1471 B.n574 VSUBS 0.007794f
C1472 B.n575 VSUBS 0.007794f
C1473 B.n576 VSUBS 0.007794f
C1474 B.n577 VSUBS 0.007794f
C1475 B.n578 VSUBS 0.007794f
C1476 B.n579 VSUBS 0.007794f
C1477 B.n580 VSUBS 0.007794f
C1478 B.n581 VSUBS 0.007794f
C1479 B.n582 VSUBS 0.007794f
C1480 B.n583 VSUBS 0.007794f
C1481 B.n584 VSUBS 0.007794f
C1482 B.n585 VSUBS 0.007794f
C1483 B.n586 VSUBS 0.007794f
C1484 B.n587 VSUBS 0.007794f
C1485 B.n588 VSUBS 0.007794f
C1486 B.n589 VSUBS 0.007794f
C1487 B.n590 VSUBS 0.007794f
C1488 B.n591 VSUBS 0.007794f
C1489 B.n592 VSUBS 0.007794f
C1490 B.n593 VSUBS 0.007794f
C1491 B.n594 VSUBS 0.007794f
C1492 B.n595 VSUBS 0.007794f
C1493 B.n596 VSUBS 0.007794f
C1494 B.n597 VSUBS 0.007794f
C1495 B.n598 VSUBS 0.007794f
C1496 B.n599 VSUBS 0.007794f
C1497 B.n600 VSUBS 0.007794f
C1498 B.n601 VSUBS 0.007794f
C1499 B.n602 VSUBS 0.007794f
C1500 B.n603 VSUBS 0.007794f
C1501 B.n604 VSUBS 0.007794f
C1502 B.n605 VSUBS 0.007794f
C1503 B.n606 VSUBS 0.007794f
C1504 B.n607 VSUBS 0.007794f
C1505 B.n608 VSUBS 0.007794f
C1506 B.n609 VSUBS 0.007794f
C1507 B.n610 VSUBS 0.007794f
C1508 B.n611 VSUBS 0.007794f
C1509 B.n612 VSUBS 0.007794f
C1510 B.n613 VSUBS 0.007794f
C1511 B.n614 VSUBS 0.007794f
C1512 B.n615 VSUBS 0.007794f
C1513 B.n616 VSUBS 0.007794f
C1514 B.n617 VSUBS 0.007794f
C1515 B.n618 VSUBS 0.007794f
C1516 B.n619 VSUBS 0.007794f
C1517 B.n620 VSUBS 0.007794f
C1518 B.n621 VSUBS 0.005387f
C1519 B.n622 VSUBS 0.018059f
C1520 B.n623 VSUBS 0.006304f
C1521 B.n624 VSUBS 0.007794f
C1522 B.n625 VSUBS 0.007794f
C1523 B.n626 VSUBS 0.007794f
C1524 B.n627 VSUBS 0.007794f
C1525 B.n628 VSUBS 0.007794f
C1526 B.n629 VSUBS 0.007794f
C1527 B.n630 VSUBS 0.007794f
C1528 B.n631 VSUBS 0.007794f
C1529 B.n632 VSUBS 0.007794f
C1530 B.n633 VSUBS 0.007794f
C1531 B.n634 VSUBS 0.007794f
C1532 B.n635 VSUBS 0.006304f
C1533 B.n636 VSUBS 0.018059f
C1534 B.n637 VSUBS 0.005387f
C1535 B.n638 VSUBS 0.007794f
C1536 B.n639 VSUBS 0.007794f
C1537 B.n640 VSUBS 0.007794f
C1538 B.n641 VSUBS 0.007794f
C1539 B.n642 VSUBS 0.007794f
C1540 B.n643 VSUBS 0.007794f
C1541 B.n644 VSUBS 0.007794f
C1542 B.n645 VSUBS 0.007794f
C1543 B.n646 VSUBS 0.007794f
C1544 B.n647 VSUBS 0.007794f
C1545 B.n648 VSUBS 0.007794f
C1546 B.n649 VSUBS 0.007794f
C1547 B.n650 VSUBS 0.007794f
C1548 B.n651 VSUBS 0.007794f
C1549 B.n652 VSUBS 0.007794f
C1550 B.n653 VSUBS 0.007794f
C1551 B.n654 VSUBS 0.007794f
C1552 B.n655 VSUBS 0.007794f
C1553 B.n656 VSUBS 0.007794f
C1554 B.n657 VSUBS 0.007794f
C1555 B.n658 VSUBS 0.007794f
C1556 B.n659 VSUBS 0.007794f
C1557 B.n660 VSUBS 0.007794f
C1558 B.n661 VSUBS 0.007794f
C1559 B.n662 VSUBS 0.007794f
C1560 B.n663 VSUBS 0.007794f
C1561 B.n664 VSUBS 0.007794f
C1562 B.n665 VSUBS 0.007794f
C1563 B.n666 VSUBS 0.007794f
C1564 B.n667 VSUBS 0.007794f
C1565 B.n668 VSUBS 0.007794f
C1566 B.n669 VSUBS 0.007794f
C1567 B.n670 VSUBS 0.007794f
C1568 B.n671 VSUBS 0.007794f
C1569 B.n672 VSUBS 0.007794f
C1570 B.n673 VSUBS 0.007794f
C1571 B.n674 VSUBS 0.007794f
C1572 B.n675 VSUBS 0.007794f
C1573 B.n676 VSUBS 0.007794f
C1574 B.n677 VSUBS 0.007794f
C1575 B.n678 VSUBS 0.007794f
C1576 B.n679 VSUBS 0.007794f
C1577 B.n680 VSUBS 0.007794f
C1578 B.n681 VSUBS 0.007794f
C1579 B.n682 VSUBS 0.007794f
C1580 B.n683 VSUBS 0.007794f
C1581 B.n684 VSUBS 0.007794f
C1582 B.n685 VSUBS 0.007794f
C1583 B.n686 VSUBS 0.007794f
C1584 B.n687 VSUBS 0.007794f
C1585 B.n688 VSUBS 0.007794f
C1586 B.n689 VSUBS 0.007794f
C1587 B.n690 VSUBS 0.007794f
C1588 B.n691 VSUBS 0.007794f
C1589 B.n692 VSUBS 0.007794f
C1590 B.n693 VSUBS 0.007794f
C1591 B.n694 VSUBS 0.007794f
C1592 B.n695 VSUBS 0.007794f
C1593 B.n696 VSUBS 0.007794f
C1594 B.n697 VSUBS 0.007794f
C1595 B.n698 VSUBS 0.007794f
C1596 B.n699 VSUBS 0.007794f
C1597 B.n700 VSUBS 0.007794f
C1598 B.n701 VSUBS 0.007794f
C1599 B.n702 VSUBS 0.007794f
C1600 B.n703 VSUBS 0.007794f
C1601 B.n704 VSUBS 0.007794f
C1602 B.n705 VSUBS 0.007794f
C1603 B.n706 VSUBS 0.007794f
C1604 B.n707 VSUBS 0.007794f
C1605 B.n708 VSUBS 0.007794f
C1606 B.n709 VSUBS 0.007794f
C1607 B.n710 VSUBS 0.007794f
C1608 B.n711 VSUBS 0.007794f
C1609 B.n712 VSUBS 0.007794f
C1610 B.n713 VSUBS 0.007794f
C1611 B.n714 VSUBS 0.007794f
C1612 B.n715 VSUBS 0.007794f
C1613 B.n716 VSUBS 0.007794f
C1614 B.n717 VSUBS 0.007794f
C1615 B.n718 VSUBS 0.007794f
C1616 B.n719 VSUBS 0.007794f
C1617 B.n720 VSUBS 0.018863f
C1618 B.n721 VSUBS 0.017816f
C1619 B.n722 VSUBS 0.017816f
C1620 B.n723 VSUBS 0.007794f
C1621 B.n724 VSUBS 0.007794f
C1622 B.n725 VSUBS 0.007794f
C1623 B.n726 VSUBS 0.007794f
C1624 B.n727 VSUBS 0.007794f
C1625 B.n728 VSUBS 0.007794f
C1626 B.n729 VSUBS 0.007794f
C1627 B.n730 VSUBS 0.007794f
C1628 B.n731 VSUBS 0.007794f
C1629 B.n732 VSUBS 0.007794f
C1630 B.n733 VSUBS 0.007794f
C1631 B.n734 VSUBS 0.007794f
C1632 B.n735 VSUBS 0.007794f
C1633 B.n736 VSUBS 0.007794f
C1634 B.n737 VSUBS 0.007794f
C1635 B.n738 VSUBS 0.007794f
C1636 B.n739 VSUBS 0.007794f
C1637 B.n740 VSUBS 0.007794f
C1638 B.n741 VSUBS 0.007794f
C1639 B.n742 VSUBS 0.007794f
C1640 B.n743 VSUBS 0.007794f
C1641 B.n744 VSUBS 0.007794f
C1642 B.n745 VSUBS 0.007794f
C1643 B.n746 VSUBS 0.007794f
C1644 B.n747 VSUBS 0.007794f
C1645 B.n748 VSUBS 0.007794f
C1646 B.n749 VSUBS 0.007794f
C1647 B.n750 VSUBS 0.007794f
C1648 B.n751 VSUBS 0.007794f
C1649 B.n752 VSUBS 0.007794f
C1650 B.n753 VSUBS 0.007794f
C1651 B.n754 VSUBS 0.007794f
C1652 B.n755 VSUBS 0.007794f
C1653 B.n756 VSUBS 0.007794f
C1654 B.n757 VSUBS 0.007794f
C1655 B.n758 VSUBS 0.007794f
C1656 B.n759 VSUBS 0.007794f
C1657 B.n760 VSUBS 0.007794f
C1658 B.n761 VSUBS 0.007794f
C1659 B.n762 VSUBS 0.007794f
C1660 B.n763 VSUBS 0.007794f
C1661 B.n764 VSUBS 0.007794f
C1662 B.n765 VSUBS 0.007794f
C1663 B.n766 VSUBS 0.007794f
C1664 B.n767 VSUBS 0.007794f
C1665 B.n768 VSUBS 0.007794f
C1666 B.n769 VSUBS 0.007794f
C1667 B.n770 VSUBS 0.007794f
C1668 B.n771 VSUBS 0.010171f
C1669 B.n772 VSUBS 0.010835f
C1670 B.n773 VSUBS 0.021546f
.ends

