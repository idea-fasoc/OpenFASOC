* NGSPICE file created from diff_pair_sample_0161.ext - technology: sky130A

.subckt diff_pair_sample_0161 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t10 VP.t0 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4784 pd=9.29 as=1.4784 ps=9.29 w=8.96 l=0.25
X1 VTAIL.t11 VN.t0 VDD2.t5 B.t19 sky130_fd_pr__nfet_01v8 ad=1.4784 pd=9.29 as=1.4784 ps=9.29 w=8.96 l=0.25
X2 VDD1.t3 VP.t1 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4944 pd=18.7 as=1.4784 ps=9.29 w=8.96 l=0.25
X3 VDD1.t0 VP.t2 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4944 pd=18.7 as=1.4784 ps=9.29 w=8.96 l=0.25
X4 B.t18 B.t16 B.t17 B.t6 sky130_fd_pr__nfet_01v8 ad=3.4944 pd=18.7 as=0 ps=0 w=8.96 l=0.25
X5 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=3.4944 pd=18.7 as=0 ps=0 w=8.96 l=0.25
X6 VDD1.t4 VP.t3 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4784 pd=9.29 as=3.4944 ps=18.7 w=8.96 l=0.25
X7 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=3.4944 pd=18.7 as=0 ps=0 w=8.96 l=0.25
X8 VTAIL.t6 VP.t4 VDD1.t1 B.t19 sky130_fd_pr__nfet_01v8 ad=1.4784 pd=9.29 as=1.4784 ps=9.29 w=8.96 l=0.25
X9 VDD2.t4 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.4944 pd=18.7 as=1.4784 ps=9.29 w=8.96 l=0.25
X10 VDD2.t3 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4784 pd=9.29 as=3.4944 ps=18.7 w=8.96 l=0.25
X11 VDD2.t2 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4784 pd=9.29 as=3.4944 ps=18.7 w=8.96 l=0.25
X12 VDD1.t2 VP.t5 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.4784 pd=9.29 as=3.4944 ps=18.7 w=8.96 l=0.25
X13 VDD2.t1 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.4944 pd=18.7 as=1.4784 ps=9.29 w=8.96 l=0.25
X14 B.t8 B.t5 B.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=3.4944 pd=18.7 as=0 ps=0 w=8.96 l=0.25
X15 VTAIL.t1 VN.t5 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4784 pd=9.29 as=1.4784 ps=9.29 w=8.96 l=0.25
R0 VP.n7 VP.t5 1039.19
R1 VP.n5 VP.t1 1039.19
R2 VP.n0 VP.t2 1039.19
R3 VP.n2 VP.t3 1039.19
R4 VP.n6 VP.t4 990.992
R5 VP.n1 VP.t0 990.992
R6 VP.n3 VP.n0 161.489
R7 VP.n8 VP.n7 161.3
R8 VP.n3 VP.n2 161.3
R9 VP.n5 VP.n4 161.3
R10 VP.n4 VP.n3 37.2505
R11 VP.n6 VP.n5 36.5157
R12 VP.n7 VP.n6 36.5157
R13 VP.n1 VP.n0 36.5157
R14 VP.n2 VP.n1 36.5157
R15 VP.n8 VP.n4 0.189894
R16 VP VP.n8 0.0516364
R17 VDD1 VDD1.t0 67.4048
R18 VDD1.n1 VDD1.t3 67.2911
R19 VDD1.n1 VDD1.n0 64.8312
R20 VDD1.n3 VDD1.n2 64.7617
R21 VDD1.n3 VDD1.n1 33.8974
R22 VDD1.n2 VDD1.t5 2.21032
R23 VDD1.n2 VDD1.t4 2.21032
R24 VDD1.n0 VDD1.t1 2.21032
R25 VDD1.n0 VDD1.t2 2.21032
R26 VDD1 VDD1.n3 0.0673103
R27 VTAIL.n7 VTAIL.t4 50.2929
R28 VTAIL.n11 VTAIL.t2 50.2926
R29 VTAIL.n2 VTAIL.t5 50.2926
R30 VTAIL.n10 VTAIL.t7 50.2926
R31 VTAIL.n9 VTAIL.n8 48.083
R32 VTAIL.n6 VTAIL.n5 48.083
R33 VTAIL.n1 VTAIL.n0 48.0828
R34 VTAIL.n4 VTAIL.n3 48.0828
R35 VTAIL.n6 VTAIL.n4 21.091
R36 VTAIL.n11 VTAIL.n10 20.591
R37 VTAIL.n0 VTAIL.t3 2.21032
R38 VTAIL.n0 VTAIL.t1 2.21032
R39 VTAIL.n3 VTAIL.t9 2.21032
R40 VTAIL.n3 VTAIL.t6 2.21032
R41 VTAIL.n8 VTAIL.t8 2.21032
R42 VTAIL.n8 VTAIL.t10 2.21032
R43 VTAIL.n5 VTAIL.t0 2.21032
R44 VTAIL.n5 VTAIL.t11 2.21032
R45 VTAIL.n9 VTAIL.n7 0.720328
R46 VTAIL.n2 VTAIL.n1 0.720328
R47 VTAIL.n7 VTAIL.n6 0.5005
R48 VTAIL.n10 VTAIL.n9 0.5005
R49 VTAIL.n4 VTAIL.n2 0.5005
R50 VTAIL VTAIL.n11 0.31731
R51 VTAIL VTAIL.n1 0.18369
R52 B.n288 B.t16 1088.04
R53 B.n285 B.t5 1088.04
R54 B.n74 B.t9 1088.04
R55 B.n71 B.t13 1088.04
R56 B.n506 B.n505 585
R57 B.n507 B.n506 585
R58 B.n219 B.n69 585
R59 B.n218 B.n217 585
R60 B.n216 B.n215 585
R61 B.n214 B.n213 585
R62 B.n212 B.n211 585
R63 B.n210 B.n209 585
R64 B.n208 B.n207 585
R65 B.n206 B.n205 585
R66 B.n204 B.n203 585
R67 B.n202 B.n201 585
R68 B.n200 B.n199 585
R69 B.n198 B.n197 585
R70 B.n196 B.n195 585
R71 B.n194 B.n193 585
R72 B.n192 B.n191 585
R73 B.n190 B.n189 585
R74 B.n188 B.n187 585
R75 B.n186 B.n185 585
R76 B.n184 B.n183 585
R77 B.n182 B.n181 585
R78 B.n180 B.n179 585
R79 B.n178 B.n177 585
R80 B.n176 B.n175 585
R81 B.n174 B.n173 585
R82 B.n172 B.n171 585
R83 B.n170 B.n169 585
R84 B.n168 B.n167 585
R85 B.n166 B.n165 585
R86 B.n164 B.n163 585
R87 B.n162 B.n161 585
R88 B.n160 B.n159 585
R89 B.n158 B.n157 585
R90 B.n156 B.n155 585
R91 B.n154 B.n153 585
R92 B.n152 B.n151 585
R93 B.n150 B.n149 585
R94 B.n148 B.n147 585
R95 B.n146 B.n145 585
R96 B.n144 B.n143 585
R97 B.n142 B.n141 585
R98 B.n140 B.n139 585
R99 B.n137 B.n136 585
R100 B.n135 B.n134 585
R101 B.n133 B.n132 585
R102 B.n131 B.n130 585
R103 B.n129 B.n128 585
R104 B.n127 B.n126 585
R105 B.n125 B.n124 585
R106 B.n123 B.n122 585
R107 B.n121 B.n120 585
R108 B.n119 B.n118 585
R109 B.n117 B.n116 585
R110 B.n115 B.n114 585
R111 B.n113 B.n112 585
R112 B.n111 B.n110 585
R113 B.n109 B.n108 585
R114 B.n107 B.n106 585
R115 B.n105 B.n104 585
R116 B.n103 B.n102 585
R117 B.n101 B.n100 585
R118 B.n99 B.n98 585
R119 B.n97 B.n96 585
R120 B.n95 B.n94 585
R121 B.n93 B.n92 585
R122 B.n91 B.n90 585
R123 B.n89 B.n88 585
R124 B.n87 B.n86 585
R125 B.n85 B.n84 585
R126 B.n83 B.n82 585
R127 B.n81 B.n80 585
R128 B.n79 B.n78 585
R129 B.n77 B.n76 585
R130 B.n32 B.n31 585
R131 B.n510 B.n509 585
R132 B.n504 B.n70 585
R133 B.n70 B.n29 585
R134 B.n503 B.n28 585
R135 B.n514 B.n28 585
R136 B.n502 B.n27 585
R137 B.n515 B.n27 585
R138 B.n501 B.n26 585
R139 B.n516 B.n26 585
R140 B.n500 B.n499 585
R141 B.n499 B.n25 585
R142 B.n498 B.n21 585
R143 B.n522 B.n21 585
R144 B.n497 B.n20 585
R145 B.n523 B.n20 585
R146 B.n496 B.n19 585
R147 B.n524 B.n19 585
R148 B.n495 B.n494 585
R149 B.n494 B.n15 585
R150 B.n493 B.n14 585
R151 B.n530 B.n14 585
R152 B.n492 B.n13 585
R153 B.n531 B.n13 585
R154 B.n491 B.n12 585
R155 B.n532 B.n12 585
R156 B.n490 B.n489 585
R157 B.n489 B.n11 585
R158 B.n488 B.n7 585
R159 B.n538 B.n7 585
R160 B.n487 B.n6 585
R161 B.n539 B.n6 585
R162 B.n486 B.n5 585
R163 B.n540 B.n5 585
R164 B.n485 B.n484 585
R165 B.n484 B.n4 585
R166 B.n483 B.n220 585
R167 B.n483 B.n482 585
R168 B.n472 B.n221 585
R169 B.n475 B.n221 585
R170 B.n474 B.n473 585
R171 B.n476 B.n474 585
R172 B.n471 B.n225 585
R173 B.n229 B.n225 585
R174 B.n470 B.n469 585
R175 B.n469 B.n468 585
R176 B.n227 B.n226 585
R177 B.n228 B.n227 585
R178 B.n461 B.n460 585
R179 B.n462 B.n461 585
R180 B.n459 B.n234 585
R181 B.n234 B.n233 585
R182 B.n458 B.n457 585
R183 B.n457 B.n456 585
R184 B.n236 B.n235 585
R185 B.n449 B.n236 585
R186 B.n448 B.n447 585
R187 B.n450 B.n448 585
R188 B.n446 B.n241 585
R189 B.n241 B.n240 585
R190 B.n445 B.n444 585
R191 B.n444 B.n443 585
R192 B.n243 B.n242 585
R193 B.n244 B.n243 585
R194 B.n439 B.n438 585
R195 B.n247 B.n246 585
R196 B.n435 B.n434 585
R197 B.n436 B.n435 585
R198 B.n433 B.n284 585
R199 B.n432 B.n431 585
R200 B.n430 B.n429 585
R201 B.n428 B.n427 585
R202 B.n426 B.n425 585
R203 B.n424 B.n423 585
R204 B.n422 B.n421 585
R205 B.n420 B.n419 585
R206 B.n418 B.n417 585
R207 B.n416 B.n415 585
R208 B.n414 B.n413 585
R209 B.n412 B.n411 585
R210 B.n410 B.n409 585
R211 B.n408 B.n407 585
R212 B.n406 B.n405 585
R213 B.n404 B.n403 585
R214 B.n402 B.n401 585
R215 B.n400 B.n399 585
R216 B.n398 B.n397 585
R217 B.n396 B.n395 585
R218 B.n394 B.n393 585
R219 B.n392 B.n391 585
R220 B.n390 B.n389 585
R221 B.n388 B.n387 585
R222 B.n386 B.n385 585
R223 B.n384 B.n383 585
R224 B.n382 B.n381 585
R225 B.n380 B.n379 585
R226 B.n378 B.n377 585
R227 B.n376 B.n375 585
R228 B.n374 B.n373 585
R229 B.n372 B.n371 585
R230 B.n370 B.n369 585
R231 B.n368 B.n367 585
R232 B.n366 B.n365 585
R233 B.n364 B.n363 585
R234 B.n362 B.n361 585
R235 B.n360 B.n359 585
R236 B.n358 B.n357 585
R237 B.n355 B.n354 585
R238 B.n353 B.n352 585
R239 B.n351 B.n350 585
R240 B.n349 B.n348 585
R241 B.n347 B.n346 585
R242 B.n345 B.n344 585
R243 B.n343 B.n342 585
R244 B.n341 B.n340 585
R245 B.n339 B.n338 585
R246 B.n337 B.n336 585
R247 B.n335 B.n334 585
R248 B.n333 B.n332 585
R249 B.n331 B.n330 585
R250 B.n329 B.n328 585
R251 B.n327 B.n326 585
R252 B.n325 B.n324 585
R253 B.n323 B.n322 585
R254 B.n321 B.n320 585
R255 B.n319 B.n318 585
R256 B.n317 B.n316 585
R257 B.n315 B.n314 585
R258 B.n313 B.n312 585
R259 B.n311 B.n310 585
R260 B.n309 B.n308 585
R261 B.n307 B.n306 585
R262 B.n305 B.n304 585
R263 B.n303 B.n302 585
R264 B.n301 B.n300 585
R265 B.n299 B.n298 585
R266 B.n297 B.n296 585
R267 B.n295 B.n294 585
R268 B.n293 B.n292 585
R269 B.n291 B.n290 585
R270 B.n440 B.n245 585
R271 B.n245 B.n244 585
R272 B.n442 B.n441 585
R273 B.n443 B.n442 585
R274 B.n239 B.n238 585
R275 B.n240 B.n239 585
R276 B.n452 B.n451 585
R277 B.n451 B.n450 585
R278 B.n453 B.n237 585
R279 B.n449 B.n237 585
R280 B.n455 B.n454 585
R281 B.n456 B.n455 585
R282 B.n232 B.n231 585
R283 B.n233 B.n232 585
R284 B.n464 B.n463 585
R285 B.n463 B.n462 585
R286 B.n465 B.n230 585
R287 B.n230 B.n228 585
R288 B.n467 B.n466 585
R289 B.n468 B.n467 585
R290 B.n224 B.n223 585
R291 B.n229 B.n224 585
R292 B.n478 B.n477 585
R293 B.n477 B.n476 585
R294 B.n479 B.n222 585
R295 B.n475 B.n222 585
R296 B.n481 B.n480 585
R297 B.n482 B.n481 585
R298 B.n2 B.n0 585
R299 B.n4 B.n2 585
R300 B.n3 B.n1 585
R301 B.n539 B.n3 585
R302 B.n537 B.n536 585
R303 B.n538 B.n537 585
R304 B.n535 B.n8 585
R305 B.n11 B.n8 585
R306 B.n534 B.n533 585
R307 B.n533 B.n532 585
R308 B.n10 B.n9 585
R309 B.n531 B.n10 585
R310 B.n529 B.n528 585
R311 B.n530 B.n529 585
R312 B.n527 B.n16 585
R313 B.n16 B.n15 585
R314 B.n526 B.n525 585
R315 B.n525 B.n524 585
R316 B.n18 B.n17 585
R317 B.n523 B.n18 585
R318 B.n521 B.n520 585
R319 B.n522 B.n521 585
R320 B.n519 B.n22 585
R321 B.n25 B.n22 585
R322 B.n518 B.n517 585
R323 B.n517 B.n516 585
R324 B.n24 B.n23 585
R325 B.n515 B.n24 585
R326 B.n513 B.n512 585
R327 B.n514 B.n513 585
R328 B.n511 B.n30 585
R329 B.n30 B.n29 585
R330 B.n542 B.n541 585
R331 B.n541 B.n540 585
R332 B.n438 B.n245 482.89
R333 B.n509 B.n30 482.89
R334 B.n290 B.n243 482.89
R335 B.n506 B.n70 482.89
R336 B.n507 B.n68 256.663
R337 B.n507 B.n67 256.663
R338 B.n507 B.n66 256.663
R339 B.n507 B.n65 256.663
R340 B.n507 B.n64 256.663
R341 B.n507 B.n63 256.663
R342 B.n507 B.n62 256.663
R343 B.n507 B.n61 256.663
R344 B.n507 B.n60 256.663
R345 B.n507 B.n59 256.663
R346 B.n507 B.n58 256.663
R347 B.n507 B.n57 256.663
R348 B.n507 B.n56 256.663
R349 B.n507 B.n55 256.663
R350 B.n507 B.n54 256.663
R351 B.n507 B.n53 256.663
R352 B.n507 B.n52 256.663
R353 B.n507 B.n51 256.663
R354 B.n507 B.n50 256.663
R355 B.n507 B.n49 256.663
R356 B.n507 B.n48 256.663
R357 B.n507 B.n47 256.663
R358 B.n507 B.n46 256.663
R359 B.n507 B.n45 256.663
R360 B.n507 B.n44 256.663
R361 B.n507 B.n43 256.663
R362 B.n507 B.n42 256.663
R363 B.n507 B.n41 256.663
R364 B.n507 B.n40 256.663
R365 B.n507 B.n39 256.663
R366 B.n507 B.n38 256.663
R367 B.n507 B.n37 256.663
R368 B.n507 B.n36 256.663
R369 B.n507 B.n35 256.663
R370 B.n507 B.n34 256.663
R371 B.n507 B.n33 256.663
R372 B.n508 B.n507 256.663
R373 B.n437 B.n436 256.663
R374 B.n436 B.n248 256.663
R375 B.n436 B.n249 256.663
R376 B.n436 B.n250 256.663
R377 B.n436 B.n251 256.663
R378 B.n436 B.n252 256.663
R379 B.n436 B.n253 256.663
R380 B.n436 B.n254 256.663
R381 B.n436 B.n255 256.663
R382 B.n436 B.n256 256.663
R383 B.n436 B.n257 256.663
R384 B.n436 B.n258 256.663
R385 B.n436 B.n259 256.663
R386 B.n436 B.n260 256.663
R387 B.n436 B.n261 256.663
R388 B.n436 B.n262 256.663
R389 B.n436 B.n263 256.663
R390 B.n436 B.n264 256.663
R391 B.n436 B.n265 256.663
R392 B.n436 B.n266 256.663
R393 B.n436 B.n267 256.663
R394 B.n436 B.n268 256.663
R395 B.n436 B.n269 256.663
R396 B.n436 B.n270 256.663
R397 B.n436 B.n271 256.663
R398 B.n436 B.n272 256.663
R399 B.n436 B.n273 256.663
R400 B.n436 B.n274 256.663
R401 B.n436 B.n275 256.663
R402 B.n436 B.n276 256.663
R403 B.n436 B.n277 256.663
R404 B.n436 B.n278 256.663
R405 B.n436 B.n279 256.663
R406 B.n436 B.n280 256.663
R407 B.n436 B.n281 256.663
R408 B.n436 B.n282 256.663
R409 B.n436 B.n283 256.663
R410 B.n442 B.n245 163.367
R411 B.n442 B.n239 163.367
R412 B.n451 B.n239 163.367
R413 B.n451 B.n237 163.367
R414 B.n455 B.n237 163.367
R415 B.n455 B.n232 163.367
R416 B.n463 B.n232 163.367
R417 B.n463 B.n230 163.367
R418 B.n467 B.n230 163.367
R419 B.n467 B.n224 163.367
R420 B.n477 B.n224 163.367
R421 B.n477 B.n222 163.367
R422 B.n481 B.n222 163.367
R423 B.n481 B.n2 163.367
R424 B.n541 B.n2 163.367
R425 B.n541 B.n3 163.367
R426 B.n537 B.n3 163.367
R427 B.n537 B.n8 163.367
R428 B.n533 B.n8 163.367
R429 B.n533 B.n10 163.367
R430 B.n529 B.n10 163.367
R431 B.n529 B.n16 163.367
R432 B.n525 B.n16 163.367
R433 B.n525 B.n18 163.367
R434 B.n521 B.n18 163.367
R435 B.n521 B.n22 163.367
R436 B.n517 B.n22 163.367
R437 B.n517 B.n24 163.367
R438 B.n513 B.n24 163.367
R439 B.n513 B.n30 163.367
R440 B.n435 B.n247 163.367
R441 B.n435 B.n284 163.367
R442 B.n431 B.n430 163.367
R443 B.n427 B.n426 163.367
R444 B.n423 B.n422 163.367
R445 B.n419 B.n418 163.367
R446 B.n415 B.n414 163.367
R447 B.n411 B.n410 163.367
R448 B.n407 B.n406 163.367
R449 B.n403 B.n402 163.367
R450 B.n399 B.n398 163.367
R451 B.n395 B.n394 163.367
R452 B.n391 B.n390 163.367
R453 B.n387 B.n386 163.367
R454 B.n383 B.n382 163.367
R455 B.n379 B.n378 163.367
R456 B.n375 B.n374 163.367
R457 B.n371 B.n370 163.367
R458 B.n367 B.n366 163.367
R459 B.n363 B.n362 163.367
R460 B.n359 B.n358 163.367
R461 B.n354 B.n353 163.367
R462 B.n350 B.n349 163.367
R463 B.n346 B.n345 163.367
R464 B.n342 B.n341 163.367
R465 B.n338 B.n337 163.367
R466 B.n334 B.n333 163.367
R467 B.n330 B.n329 163.367
R468 B.n326 B.n325 163.367
R469 B.n322 B.n321 163.367
R470 B.n318 B.n317 163.367
R471 B.n314 B.n313 163.367
R472 B.n310 B.n309 163.367
R473 B.n306 B.n305 163.367
R474 B.n302 B.n301 163.367
R475 B.n298 B.n297 163.367
R476 B.n294 B.n293 163.367
R477 B.n444 B.n243 163.367
R478 B.n444 B.n241 163.367
R479 B.n448 B.n241 163.367
R480 B.n448 B.n236 163.367
R481 B.n457 B.n236 163.367
R482 B.n457 B.n234 163.367
R483 B.n461 B.n234 163.367
R484 B.n461 B.n227 163.367
R485 B.n469 B.n227 163.367
R486 B.n469 B.n225 163.367
R487 B.n474 B.n225 163.367
R488 B.n474 B.n221 163.367
R489 B.n483 B.n221 163.367
R490 B.n484 B.n483 163.367
R491 B.n484 B.n5 163.367
R492 B.n6 B.n5 163.367
R493 B.n7 B.n6 163.367
R494 B.n489 B.n7 163.367
R495 B.n489 B.n12 163.367
R496 B.n13 B.n12 163.367
R497 B.n14 B.n13 163.367
R498 B.n494 B.n14 163.367
R499 B.n494 B.n19 163.367
R500 B.n20 B.n19 163.367
R501 B.n21 B.n20 163.367
R502 B.n499 B.n21 163.367
R503 B.n499 B.n26 163.367
R504 B.n27 B.n26 163.367
R505 B.n28 B.n27 163.367
R506 B.n70 B.n28 163.367
R507 B.n76 B.n32 163.367
R508 B.n80 B.n79 163.367
R509 B.n84 B.n83 163.367
R510 B.n88 B.n87 163.367
R511 B.n92 B.n91 163.367
R512 B.n96 B.n95 163.367
R513 B.n100 B.n99 163.367
R514 B.n104 B.n103 163.367
R515 B.n108 B.n107 163.367
R516 B.n112 B.n111 163.367
R517 B.n116 B.n115 163.367
R518 B.n120 B.n119 163.367
R519 B.n124 B.n123 163.367
R520 B.n128 B.n127 163.367
R521 B.n132 B.n131 163.367
R522 B.n136 B.n135 163.367
R523 B.n141 B.n140 163.367
R524 B.n145 B.n144 163.367
R525 B.n149 B.n148 163.367
R526 B.n153 B.n152 163.367
R527 B.n157 B.n156 163.367
R528 B.n161 B.n160 163.367
R529 B.n165 B.n164 163.367
R530 B.n169 B.n168 163.367
R531 B.n173 B.n172 163.367
R532 B.n177 B.n176 163.367
R533 B.n181 B.n180 163.367
R534 B.n185 B.n184 163.367
R535 B.n189 B.n188 163.367
R536 B.n193 B.n192 163.367
R537 B.n197 B.n196 163.367
R538 B.n201 B.n200 163.367
R539 B.n205 B.n204 163.367
R540 B.n209 B.n208 163.367
R541 B.n213 B.n212 163.367
R542 B.n217 B.n216 163.367
R543 B.n506 B.n69 163.367
R544 B.n436 B.n244 91.9569
R545 B.n507 B.n29 91.9569
R546 B.n288 B.t18 81.9211
R547 B.n71 B.t14 81.9211
R548 B.n285 B.t8 81.9104
R549 B.n74 B.t11 81.9104
R550 B.n438 B.n437 71.676
R551 B.n284 B.n248 71.676
R552 B.n430 B.n249 71.676
R553 B.n426 B.n250 71.676
R554 B.n422 B.n251 71.676
R555 B.n418 B.n252 71.676
R556 B.n414 B.n253 71.676
R557 B.n410 B.n254 71.676
R558 B.n406 B.n255 71.676
R559 B.n402 B.n256 71.676
R560 B.n398 B.n257 71.676
R561 B.n394 B.n258 71.676
R562 B.n390 B.n259 71.676
R563 B.n386 B.n260 71.676
R564 B.n382 B.n261 71.676
R565 B.n378 B.n262 71.676
R566 B.n374 B.n263 71.676
R567 B.n370 B.n264 71.676
R568 B.n366 B.n265 71.676
R569 B.n362 B.n266 71.676
R570 B.n358 B.n267 71.676
R571 B.n353 B.n268 71.676
R572 B.n349 B.n269 71.676
R573 B.n345 B.n270 71.676
R574 B.n341 B.n271 71.676
R575 B.n337 B.n272 71.676
R576 B.n333 B.n273 71.676
R577 B.n329 B.n274 71.676
R578 B.n325 B.n275 71.676
R579 B.n321 B.n276 71.676
R580 B.n317 B.n277 71.676
R581 B.n313 B.n278 71.676
R582 B.n309 B.n279 71.676
R583 B.n305 B.n280 71.676
R584 B.n301 B.n281 71.676
R585 B.n297 B.n282 71.676
R586 B.n293 B.n283 71.676
R587 B.n509 B.n508 71.676
R588 B.n76 B.n33 71.676
R589 B.n80 B.n34 71.676
R590 B.n84 B.n35 71.676
R591 B.n88 B.n36 71.676
R592 B.n92 B.n37 71.676
R593 B.n96 B.n38 71.676
R594 B.n100 B.n39 71.676
R595 B.n104 B.n40 71.676
R596 B.n108 B.n41 71.676
R597 B.n112 B.n42 71.676
R598 B.n116 B.n43 71.676
R599 B.n120 B.n44 71.676
R600 B.n124 B.n45 71.676
R601 B.n128 B.n46 71.676
R602 B.n132 B.n47 71.676
R603 B.n136 B.n48 71.676
R604 B.n141 B.n49 71.676
R605 B.n145 B.n50 71.676
R606 B.n149 B.n51 71.676
R607 B.n153 B.n52 71.676
R608 B.n157 B.n53 71.676
R609 B.n161 B.n54 71.676
R610 B.n165 B.n55 71.676
R611 B.n169 B.n56 71.676
R612 B.n173 B.n57 71.676
R613 B.n177 B.n58 71.676
R614 B.n181 B.n59 71.676
R615 B.n185 B.n60 71.676
R616 B.n189 B.n61 71.676
R617 B.n193 B.n62 71.676
R618 B.n197 B.n63 71.676
R619 B.n201 B.n64 71.676
R620 B.n205 B.n65 71.676
R621 B.n209 B.n66 71.676
R622 B.n213 B.n67 71.676
R623 B.n217 B.n68 71.676
R624 B.n69 B.n68 71.676
R625 B.n216 B.n67 71.676
R626 B.n212 B.n66 71.676
R627 B.n208 B.n65 71.676
R628 B.n204 B.n64 71.676
R629 B.n200 B.n63 71.676
R630 B.n196 B.n62 71.676
R631 B.n192 B.n61 71.676
R632 B.n188 B.n60 71.676
R633 B.n184 B.n59 71.676
R634 B.n180 B.n58 71.676
R635 B.n176 B.n57 71.676
R636 B.n172 B.n56 71.676
R637 B.n168 B.n55 71.676
R638 B.n164 B.n54 71.676
R639 B.n160 B.n53 71.676
R640 B.n156 B.n52 71.676
R641 B.n152 B.n51 71.676
R642 B.n148 B.n50 71.676
R643 B.n144 B.n49 71.676
R644 B.n140 B.n48 71.676
R645 B.n135 B.n47 71.676
R646 B.n131 B.n46 71.676
R647 B.n127 B.n45 71.676
R648 B.n123 B.n44 71.676
R649 B.n119 B.n43 71.676
R650 B.n115 B.n42 71.676
R651 B.n111 B.n41 71.676
R652 B.n107 B.n40 71.676
R653 B.n103 B.n39 71.676
R654 B.n99 B.n38 71.676
R655 B.n95 B.n37 71.676
R656 B.n91 B.n36 71.676
R657 B.n87 B.n35 71.676
R658 B.n83 B.n34 71.676
R659 B.n79 B.n33 71.676
R660 B.n508 B.n32 71.676
R661 B.n437 B.n247 71.676
R662 B.n431 B.n248 71.676
R663 B.n427 B.n249 71.676
R664 B.n423 B.n250 71.676
R665 B.n419 B.n251 71.676
R666 B.n415 B.n252 71.676
R667 B.n411 B.n253 71.676
R668 B.n407 B.n254 71.676
R669 B.n403 B.n255 71.676
R670 B.n399 B.n256 71.676
R671 B.n395 B.n257 71.676
R672 B.n391 B.n258 71.676
R673 B.n387 B.n259 71.676
R674 B.n383 B.n260 71.676
R675 B.n379 B.n261 71.676
R676 B.n375 B.n262 71.676
R677 B.n371 B.n263 71.676
R678 B.n367 B.n264 71.676
R679 B.n363 B.n265 71.676
R680 B.n359 B.n266 71.676
R681 B.n354 B.n267 71.676
R682 B.n350 B.n268 71.676
R683 B.n346 B.n269 71.676
R684 B.n342 B.n270 71.676
R685 B.n338 B.n271 71.676
R686 B.n334 B.n272 71.676
R687 B.n330 B.n273 71.676
R688 B.n326 B.n274 71.676
R689 B.n322 B.n275 71.676
R690 B.n318 B.n276 71.676
R691 B.n314 B.n277 71.676
R692 B.n310 B.n278 71.676
R693 B.n306 B.n279 71.676
R694 B.n302 B.n280 71.676
R695 B.n298 B.n281 71.676
R696 B.n294 B.n282 71.676
R697 B.n290 B.n283 71.676
R698 B.n289 B.t17 70.6727
R699 B.n72 B.t15 70.6727
R700 B.n286 B.t7 70.6619
R701 B.n75 B.t12 70.6619
R702 B.n356 B.n289 59.5399
R703 B.n287 B.n286 59.5399
R704 B.n138 B.n75 59.5399
R705 B.n73 B.n72 59.5399
R706 B.n443 B.n244 52.547
R707 B.n443 B.n240 52.547
R708 B.n450 B.n240 52.547
R709 B.n450 B.n449 52.547
R710 B.n456 B.n233 52.547
R711 B.n462 B.n233 52.547
R712 B.n462 B.n228 52.547
R713 B.n468 B.n228 52.547
R714 B.n476 B.n475 52.547
R715 B.n482 B.n4 52.547
R716 B.n540 B.n4 52.547
R717 B.n540 B.n539 52.547
R718 B.n539 B.n538 52.547
R719 B.n532 B.n11 52.547
R720 B.n530 B.n15 52.547
R721 B.n524 B.n15 52.547
R722 B.n524 B.n523 52.547
R723 B.n523 B.n522 52.547
R724 B.n516 B.n25 52.547
R725 B.n516 B.n515 52.547
R726 B.n515 B.n514 52.547
R727 B.n514 B.n29 52.547
R728 B.t0 B.n229 45.5924
R729 B.n531 B.t2 45.5924
R730 B.n229 B.t19 44.0469
R731 B.t1 B.n531 44.0469
R732 B.n456 B.t6 40.9559
R733 B.n522 B.t10 40.9559
R734 B.n511 B.n510 31.3761
R735 B.n505 B.n504 31.3761
R736 B.n291 B.n242 31.3761
R737 B.n440 B.n439 31.3761
R738 B.n475 B.t4 28.592
R739 B.n11 B.t3 28.592
R740 B.n482 B.t4 23.9555
R741 B.n538 B.t3 23.9555
R742 B B.n542 18.0485
R743 B.n449 B.t6 11.5916
R744 B.n25 B.t10 11.5916
R745 B.n289 B.n288 11.249
R746 B.n286 B.n285 11.249
R747 B.n75 B.n74 11.249
R748 B.n72 B.n71 11.249
R749 B.n510 B.n31 10.6151
R750 B.n77 B.n31 10.6151
R751 B.n78 B.n77 10.6151
R752 B.n81 B.n78 10.6151
R753 B.n82 B.n81 10.6151
R754 B.n85 B.n82 10.6151
R755 B.n86 B.n85 10.6151
R756 B.n89 B.n86 10.6151
R757 B.n90 B.n89 10.6151
R758 B.n93 B.n90 10.6151
R759 B.n94 B.n93 10.6151
R760 B.n97 B.n94 10.6151
R761 B.n98 B.n97 10.6151
R762 B.n101 B.n98 10.6151
R763 B.n102 B.n101 10.6151
R764 B.n105 B.n102 10.6151
R765 B.n106 B.n105 10.6151
R766 B.n109 B.n106 10.6151
R767 B.n110 B.n109 10.6151
R768 B.n113 B.n110 10.6151
R769 B.n114 B.n113 10.6151
R770 B.n117 B.n114 10.6151
R771 B.n118 B.n117 10.6151
R772 B.n121 B.n118 10.6151
R773 B.n122 B.n121 10.6151
R774 B.n125 B.n122 10.6151
R775 B.n126 B.n125 10.6151
R776 B.n129 B.n126 10.6151
R777 B.n130 B.n129 10.6151
R778 B.n133 B.n130 10.6151
R779 B.n134 B.n133 10.6151
R780 B.n137 B.n134 10.6151
R781 B.n142 B.n139 10.6151
R782 B.n143 B.n142 10.6151
R783 B.n146 B.n143 10.6151
R784 B.n147 B.n146 10.6151
R785 B.n150 B.n147 10.6151
R786 B.n151 B.n150 10.6151
R787 B.n154 B.n151 10.6151
R788 B.n155 B.n154 10.6151
R789 B.n159 B.n158 10.6151
R790 B.n162 B.n159 10.6151
R791 B.n163 B.n162 10.6151
R792 B.n166 B.n163 10.6151
R793 B.n167 B.n166 10.6151
R794 B.n170 B.n167 10.6151
R795 B.n171 B.n170 10.6151
R796 B.n174 B.n171 10.6151
R797 B.n175 B.n174 10.6151
R798 B.n178 B.n175 10.6151
R799 B.n179 B.n178 10.6151
R800 B.n182 B.n179 10.6151
R801 B.n183 B.n182 10.6151
R802 B.n186 B.n183 10.6151
R803 B.n187 B.n186 10.6151
R804 B.n190 B.n187 10.6151
R805 B.n191 B.n190 10.6151
R806 B.n194 B.n191 10.6151
R807 B.n195 B.n194 10.6151
R808 B.n198 B.n195 10.6151
R809 B.n199 B.n198 10.6151
R810 B.n202 B.n199 10.6151
R811 B.n203 B.n202 10.6151
R812 B.n206 B.n203 10.6151
R813 B.n207 B.n206 10.6151
R814 B.n210 B.n207 10.6151
R815 B.n211 B.n210 10.6151
R816 B.n214 B.n211 10.6151
R817 B.n215 B.n214 10.6151
R818 B.n218 B.n215 10.6151
R819 B.n219 B.n218 10.6151
R820 B.n505 B.n219 10.6151
R821 B.n445 B.n242 10.6151
R822 B.n446 B.n445 10.6151
R823 B.n447 B.n446 10.6151
R824 B.n447 B.n235 10.6151
R825 B.n458 B.n235 10.6151
R826 B.n459 B.n458 10.6151
R827 B.n460 B.n459 10.6151
R828 B.n460 B.n226 10.6151
R829 B.n470 B.n226 10.6151
R830 B.n471 B.n470 10.6151
R831 B.n473 B.n471 10.6151
R832 B.n473 B.n472 10.6151
R833 B.n472 B.n220 10.6151
R834 B.n485 B.n220 10.6151
R835 B.n486 B.n485 10.6151
R836 B.n487 B.n486 10.6151
R837 B.n488 B.n487 10.6151
R838 B.n490 B.n488 10.6151
R839 B.n491 B.n490 10.6151
R840 B.n492 B.n491 10.6151
R841 B.n493 B.n492 10.6151
R842 B.n495 B.n493 10.6151
R843 B.n496 B.n495 10.6151
R844 B.n497 B.n496 10.6151
R845 B.n498 B.n497 10.6151
R846 B.n500 B.n498 10.6151
R847 B.n501 B.n500 10.6151
R848 B.n502 B.n501 10.6151
R849 B.n503 B.n502 10.6151
R850 B.n504 B.n503 10.6151
R851 B.n439 B.n246 10.6151
R852 B.n434 B.n246 10.6151
R853 B.n434 B.n433 10.6151
R854 B.n433 B.n432 10.6151
R855 B.n432 B.n429 10.6151
R856 B.n429 B.n428 10.6151
R857 B.n428 B.n425 10.6151
R858 B.n425 B.n424 10.6151
R859 B.n424 B.n421 10.6151
R860 B.n421 B.n420 10.6151
R861 B.n420 B.n417 10.6151
R862 B.n417 B.n416 10.6151
R863 B.n416 B.n413 10.6151
R864 B.n413 B.n412 10.6151
R865 B.n412 B.n409 10.6151
R866 B.n409 B.n408 10.6151
R867 B.n408 B.n405 10.6151
R868 B.n405 B.n404 10.6151
R869 B.n404 B.n401 10.6151
R870 B.n401 B.n400 10.6151
R871 B.n400 B.n397 10.6151
R872 B.n397 B.n396 10.6151
R873 B.n396 B.n393 10.6151
R874 B.n393 B.n392 10.6151
R875 B.n392 B.n389 10.6151
R876 B.n389 B.n388 10.6151
R877 B.n388 B.n385 10.6151
R878 B.n385 B.n384 10.6151
R879 B.n384 B.n381 10.6151
R880 B.n381 B.n380 10.6151
R881 B.n380 B.n377 10.6151
R882 B.n377 B.n376 10.6151
R883 B.n373 B.n372 10.6151
R884 B.n372 B.n369 10.6151
R885 B.n369 B.n368 10.6151
R886 B.n368 B.n365 10.6151
R887 B.n365 B.n364 10.6151
R888 B.n364 B.n361 10.6151
R889 B.n361 B.n360 10.6151
R890 B.n360 B.n357 10.6151
R891 B.n355 B.n352 10.6151
R892 B.n352 B.n351 10.6151
R893 B.n351 B.n348 10.6151
R894 B.n348 B.n347 10.6151
R895 B.n347 B.n344 10.6151
R896 B.n344 B.n343 10.6151
R897 B.n343 B.n340 10.6151
R898 B.n340 B.n339 10.6151
R899 B.n339 B.n336 10.6151
R900 B.n336 B.n335 10.6151
R901 B.n335 B.n332 10.6151
R902 B.n332 B.n331 10.6151
R903 B.n331 B.n328 10.6151
R904 B.n328 B.n327 10.6151
R905 B.n327 B.n324 10.6151
R906 B.n324 B.n323 10.6151
R907 B.n323 B.n320 10.6151
R908 B.n320 B.n319 10.6151
R909 B.n319 B.n316 10.6151
R910 B.n316 B.n315 10.6151
R911 B.n315 B.n312 10.6151
R912 B.n312 B.n311 10.6151
R913 B.n311 B.n308 10.6151
R914 B.n308 B.n307 10.6151
R915 B.n307 B.n304 10.6151
R916 B.n304 B.n303 10.6151
R917 B.n303 B.n300 10.6151
R918 B.n300 B.n299 10.6151
R919 B.n299 B.n296 10.6151
R920 B.n296 B.n295 10.6151
R921 B.n295 B.n292 10.6151
R922 B.n292 B.n291 10.6151
R923 B.n441 B.n440 10.6151
R924 B.n441 B.n238 10.6151
R925 B.n452 B.n238 10.6151
R926 B.n453 B.n452 10.6151
R927 B.n454 B.n453 10.6151
R928 B.n454 B.n231 10.6151
R929 B.n464 B.n231 10.6151
R930 B.n465 B.n464 10.6151
R931 B.n466 B.n465 10.6151
R932 B.n466 B.n223 10.6151
R933 B.n478 B.n223 10.6151
R934 B.n479 B.n478 10.6151
R935 B.n480 B.n479 10.6151
R936 B.n480 B.n0 10.6151
R937 B.n536 B.n1 10.6151
R938 B.n536 B.n535 10.6151
R939 B.n535 B.n534 10.6151
R940 B.n534 B.n9 10.6151
R941 B.n528 B.n9 10.6151
R942 B.n528 B.n527 10.6151
R943 B.n527 B.n526 10.6151
R944 B.n526 B.n17 10.6151
R945 B.n520 B.n17 10.6151
R946 B.n520 B.n519 10.6151
R947 B.n519 B.n518 10.6151
R948 B.n518 B.n23 10.6151
R949 B.n512 B.n23 10.6151
R950 B.n512 B.n511 10.6151
R951 B.n476 B.t19 8.50068
R952 B.n532 B.t1 8.50068
R953 B.n468 B.t0 6.95519
R954 B.t2 B.n530 6.95519
R955 B.n139 B.n138 6.5566
R956 B.n155 B.n73 6.5566
R957 B.n373 B.n287 6.5566
R958 B.n357 B.n356 6.5566
R959 B.n138 B.n137 4.05904
R960 B.n158 B.n73 4.05904
R961 B.n376 B.n287 4.05904
R962 B.n356 B.n355 4.05904
R963 B.n542 B.n0 2.81026
R964 B.n542 B.n1 2.81026
R965 VN.n2 VN.t2 1039.19
R966 VN.n0 VN.t4 1039.19
R967 VN.n6 VN.t1 1039.19
R968 VN.n4 VN.t3 1039.19
R969 VN.n1 VN.t5 990.992
R970 VN.n5 VN.t0 990.992
R971 VN.n7 VN.n4 161.489
R972 VN.n3 VN.n0 161.489
R973 VN.n3 VN.n2 161.3
R974 VN.n7 VN.n6 161.3
R975 VN VN.n7 37.6312
R976 VN.n1 VN.n0 36.5157
R977 VN.n2 VN.n1 36.5157
R978 VN.n6 VN.n5 36.5157
R979 VN.n5 VN.n4 36.5157
R980 VN VN.n3 0.0516364
R981 VDD2.n1 VDD2.t1 67.2911
R982 VDD2.n2 VDD2.t4 66.9717
R983 VDD2.n1 VDD2.n0 64.8312
R984 VDD2 VDD2.n3 64.8285
R985 VDD2.n2 VDD2.n1 33.0644
R986 VDD2.n3 VDD2.t5 2.21032
R987 VDD2.n3 VDD2.t2 2.21032
R988 VDD2.n0 VDD2.t0 2.21032
R989 VDD2.n0 VDD2.t3 2.21032
R990 VDD2 VDD2.n2 0.43369
C0 VP VN 4.0813f
C1 VP VDD1 2.00797f
C2 VN VDD1 0.147016f
C3 VP VDD2 0.258672f
C4 VN VDD2 1.90021f
C5 VP VTAIL 1.55638f
C6 VDD2 VDD1 0.55141f
C7 VTAIL VN 1.54177f
C8 VTAIL VDD1 11.5685f
C9 VTAIL VDD2 11.5997f
C10 VDD2 B 3.571883f
C11 VDD1 B 3.823967f
C12 VTAIL B 4.896699f
C13 VN B 5.37417f
C14 VP B 4.195393f
C15 VDD2.t1 B 1.96429f
C16 VDD2.t0 B 0.176478f
C17 VDD2.t3 B 0.176478f
C18 VDD2.n0 B 1.54281f
C19 VDD2.n1 B 1.68614f
C20 VDD2.t4 B 1.96288f
C21 VDD2.n2 B 1.89961f
C22 VDD2.t5 B 0.176478f
C23 VDD2.t2 B 0.176478f
C24 VDD2.n3 B 1.54279f
C25 VN.t4 B 0.207651f
C26 VN.n0 B 0.096547f
C27 VN.t5 B 0.203552f
C28 VN.n1 B 0.086809f
C29 VN.t2 B 0.207651f
C30 VN.n2 B 0.0965f
C31 VN.n3 B 0.06493f
C32 VN.t3 B 0.207651f
C33 VN.n4 B 0.096547f
C34 VN.t1 B 0.207651f
C35 VN.t0 B 0.203552f
C36 VN.n5 B 0.086809f
C37 VN.n6 B 0.0965f
C38 VN.n7 B 1.13455f
C39 VTAIL.t3 B 0.189233f
C40 VTAIL.t1 B 0.189233f
C41 VTAIL.n0 B 1.58135f
C42 VTAIL.n1 B 0.328673f
C43 VTAIL.t5 B 2.0136f
C44 VTAIL.n2 B 0.439802f
C45 VTAIL.t9 B 0.189233f
C46 VTAIL.t6 B 0.189233f
C47 VTAIL.n3 B 1.58135f
C48 VTAIL.n4 B 1.40831f
C49 VTAIL.t0 B 0.189233f
C50 VTAIL.t11 B 0.189233f
C51 VTAIL.n5 B 1.58136f
C52 VTAIL.n6 B 1.4083f
C53 VTAIL.t4 B 2.0136f
C54 VTAIL.n7 B 0.439797f
C55 VTAIL.t8 B 0.189233f
C56 VTAIL.t10 B 0.189233f
C57 VTAIL.n8 B 1.58136f
C58 VTAIL.n9 B 0.355951f
C59 VTAIL.t7 B 2.0136f
C60 VTAIL.n10 B 1.4491f
C61 VTAIL.t2 B 2.0136f
C62 VTAIL.n11 B 1.43332f
C63 VDD1.t0 B 2.28547f
C64 VDD1.t3 B 2.28483f
C65 VDD1.t1 B 0.205276f
C66 VDD1.t2 B 0.205276f
C67 VDD1.n0 B 1.79457f
C68 VDD1.n1 B 2.03812f
C69 VDD1.t5 B 0.205276f
C70 VDD1.t4 B 0.205276f
C71 VDD1.n2 B 1.79424f
C72 VDD1.n3 B 2.18144f
C73 VP.t2 B 0.312377f
C74 VP.n0 B 0.145239f
C75 VP.t0 B 0.306209f
C76 VP.n1 B 0.130589f
C77 VP.t3 B 0.312377f
C78 VP.n2 B 0.145168f
C79 VP.n3 B 1.67485f
C80 VP.n4 B 1.66091f
C81 VP.t4 B 0.306209f
C82 VP.t1 B 0.312377f
C83 VP.n5 B 0.145168f
C84 VP.n6 B 0.130589f
C85 VP.t5 B 0.312377f
C86 VP.n7 B 0.145168f
C87 VP.n8 B 0.037357f
.ends

