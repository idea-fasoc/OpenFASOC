* NGSPICE file created from diff_pair_sample_1781.ext - technology: sky130A

.subckt diff_pair_sample_1781 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=5.0739 pd=26.8 as=0 ps=0 w=13.01 l=3.65
X1 VDD1.t9 VP.t0 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
X2 VTAIL.t0 VN.t0 VDD2.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
X3 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=5.0739 pd=26.8 as=0 ps=0 w=13.01 l=3.65
X4 VTAIL.t13 VP.t1 VDD1.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
X5 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.0739 pd=26.8 as=0 ps=0 w=13.01 l=3.65
X6 VDD1.t7 VP.t2 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=5.0739 ps=26.8 w=13.01 l=3.65
X7 VTAIL.t11 VP.t3 VDD1.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
X8 VTAIL.t15 VN.t1 VDD2.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
X9 VDD2.t7 VN.t2 VTAIL.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
X10 VTAIL.t4 VN.t3 VDD2.t6 B.t7 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
X11 VTAIL.t19 VN.t4 VDD2.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
X12 VDD1.t5 VP.t4 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=5.0739 pd=26.8 as=2.14665 ps=13.34 w=13.01 l=3.65
X13 VDD2.t4 VN.t5 VTAIL.t18 B.t4 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=5.0739 ps=26.8 w=13.01 l=3.65
X14 VTAIL.t14 VP.t5 VDD1.t4 B.t8 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
X15 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.0739 pd=26.8 as=0 ps=0 w=13.01 l=3.65
X16 VTAIL.t10 VP.t6 VDD1.t3 B.t9 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
X17 VDD2.t3 VN.t6 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.0739 pd=26.8 as=2.14665 ps=13.34 w=13.01 l=3.65
X18 VDD2.t2 VN.t7 VTAIL.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=5.0739 ps=26.8 w=13.01 l=3.65
X19 VDD2.t1 VN.t8 VTAIL.t16 B.t3 sky130_fd_pr__nfet_01v8 ad=5.0739 pd=26.8 as=2.14665 ps=13.34 w=13.01 l=3.65
X20 VDD1.t2 VP.t7 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=5.0739 pd=26.8 as=2.14665 ps=13.34 w=13.01 l=3.65
X21 VDD2.t0 VN.t9 VTAIL.t17 B.t0 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
X22 VDD1.t1 VP.t8 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=5.0739 ps=26.8 w=13.01 l=3.65
X23 VDD1.t0 VP.t9 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.14665 pd=13.34 as=2.14665 ps=13.34 w=13.01 l=3.65
R0 B.n939 B.n197 585
R1 B.n197 B.n142 585
R2 B.n941 B.n940 585
R3 B.n943 B.n196 585
R4 B.n946 B.n945 585
R5 B.n947 B.n195 585
R6 B.n949 B.n948 585
R7 B.n951 B.n194 585
R8 B.n954 B.n953 585
R9 B.n955 B.n193 585
R10 B.n957 B.n956 585
R11 B.n959 B.n192 585
R12 B.n962 B.n961 585
R13 B.n963 B.n191 585
R14 B.n965 B.n964 585
R15 B.n967 B.n190 585
R16 B.n970 B.n969 585
R17 B.n971 B.n189 585
R18 B.n973 B.n972 585
R19 B.n975 B.n188 585
R20 B.n978 B.n977 585
R21 B.n979 B.n187 585
R22 B.n981 B.n980 585
R23 B.n983 B.n186 585
R24 B.n986 B.n985 585
R25 B.n987 B.n185 585
R26 B.n989 B.n988 585
R27 B.n991 B.n184 585
R28 B.n994 B.n993 585
R29 B.n995 B.n183 585
R30 B.n997 B.n996 585
R31 B.n999 B.n182 585
R32 B.n1002 B.n1001 585
R33 B.n1003 B.n181 585
R34 B.n1005 B.n1004 585
R35 B.n1007 B.n180 585
R36 B.n1010 B.n1009 585
R37 B.n1011 B.n179 585
R38 B.n1013 B.n1012 585
R39 B.n1015 B.n178 585
R40 B.n1018 B.n1017 585
R41 B.n1019 B.n177 585
R42 B.n1021 B.n1020 585
R43 B.n1023 B.n176 585
R44 B.n1025 B.n1024 585
R45 B.n1027 B.n1026 585
R46 B.n1030 B.n1029 585
R47 B.n1031 B.n171 585
R48 B.n1033 B.n1032 585
R49 B.n1035 B.n170 585
R50 B.n1038 B.n1037 585
R51 B.n1039 B.n169 585
R52 B.n1041 B.n1040 585
R53 B.n1043 B.n168 585
R54 B.n1046 B.n1045 585
R55 B.n1048 B.n165 585
R56 B.n1050 B.n1049 585
R57 B.n1052 B.n164 585
R58 B.n1055 B.n1054 585
R59 B.n1056 B.n163 585
R60 B.n1058 B.n1057 585
R61 B.n1060 B.n162 585
R62 B.n1063 B.n1062 585
R63 B.n1064 B.n161 585
R64 B.n1066 B.n1065 585
R65 B.n1068 B.n160 585
R66 B.n1071 B.n1070 585
R67 B.n1072 B.n159 585
R68 B.n1074 B.n1073 585
R69 B.n1076 B.n158 585
R70 B.n1079 B.n1078 585
R71 B.n1080 B.n157 585
R72 B.n1082 B.n1081 585
R73 B.n1084 B.n156 585
R74 B.n1087 B.n1086 585
R75 B.n1088 B.n155 585
R76 B.n1090 B.n1089 585
R77 B.n1092 B.n154 585
R78 B.n1095 B.n1094 585
R79 B.n1096 B.n153 585
R80 B.n1098 B.n1097 585
R81 B.n1100 B.n152 585
R82 B.n1103 B.n1102 585
R83 B.n1104 B.n151 585
R84 B.n1106 B.n1105 585
R85 B.n1108 B.n150 585
R86 B.n1111 B.n1110 585
R87 B.n1112 B.n149 585
R88 B.n1114 B.n1113 585
R89 B.n1116 B.n148 585
R90 B.n1119 B.n1118 585
R91 B.n1120 B.n147 585
R92 B.n1122 B.n1121 585
R93 B.n1124 B.n146 585
R94 B.n1127 B.n1126 585
R95 B.n1128 B.n145 585
R96 B.n1130 B.n1129 585
R97 B.n1132 B.n144 585
R98 B.n1135 B.n1134 585
R99 B.n1136 B.n143 585
R100 B.n938 B.n141 585
R101 B.n1139 B.n141 585
R102 B.n937 B.n140 585
R103 B.n1140 B.n140 585
R104 B.n936 B.n139 585
R105 B.n1141 B.n139 585
R106 B.n935 B.n934 585
R107 B.n934 B.n135 585
R108 B.n933 B.n134 585
R109 B.n1147 B.n134 585
R110 B.n932 B.n133 585
R111 B.n1148 B.n133 585
R112 B.n931 B.n132 585
R113 B.n1149 B.n132 585
R114 B.n930 B.n929 585
R115 B.n929 B.n128 585
R116 B.n928 B.n127 585
R117 B.n1155 B.n127 585
R118 B.n927 B.n126 585
R119 B.n1156 B.n126 585
R120 B.n926 B.n125 585
R121 B.n1157 B.n125 585
R122 B.n925 B.n924 585
R123 B.n924 B.n121 585
R124 B.n923 B.n120 585
R125 B.n1163 B.n120 585
R126 B.n922 B.n119 585
R127 B.n1164 B.n119 585
R128 B.n921 B.n118 585
R129 B.n1165 B.n118 585
R130 B.n920 B.n919 585
R131 B.n919 B.n114 585
R132 B.n918 B.n113 585
R133 B.n1171 B.n113 585
R134 B.n917 B.n112 585
R135 B.n1172 B.n112 585
R136 B.n916 B.n111 585
R137 B.n1173 B.n111 585
R138 B.n915 B.n914 585
R139 B.n914 B.n107 585
R140 B.n913 B.n106 585
R141 B.n1179 B.n106 585
R142 B.n912 B.n105 585
R143 B.n1180 B.n105 585
R144 B.n911 B.n104 585
R145 B.n1181 B.n104 585
R146 B.n910 B.n909 585
R147 B.n909 B.n100 585
R148 B.n908 B.n99 585
R149 B.n1187 B.n99 585
R150 B.n907 B.n98 585
R151 B.n1188 B.n98 585
R152 B.n906 B.n97 585
R153 B.n1189 B.n97 585
R154 B.n905 B.n904 585
R155 B.n904 B.n93 585
R156 B.n903 B.n92 585
R157 B.n1195 B.n92 585
R158 B.n902 B.n91 585
R159 B.n1196 B.n91 585
R160 B.n901 B.n90 585
R161 B.n1197 B.n90 585
R162 B.n900 B.n899 585
R163 B.n899 B.n86 585
R164 B.n898 B.n85 585
R165 B.n1203 B.n85 585
R166 B.n897 B.n84 585
R167 B.n1204 B.n84 585
R168 B.n896 B.n83 585
R169 B.n1205 B.n83 585
R170 B.n895 B.n894 585
R171 B.n894 B.n82 585
R172 B.n893 B.n78 585
R173 B.n1211 B.n78 585
R174 B.n892 B.n77 585
R175 B.n1212 B.n77 585
R176 B.n891 B.n76 585
R177 B.n1213 B.n76 585
R178 B.n890 B.n889 585
R179 B.n889 B.n72 585
R180 B.n888 B.n71 585
R181 B.n1219 B.n71 585
R182 B.n887 B.n70 585
R183 B.n1220 B.n70 585
R184 B.n886 B.n69 585
R185 B.n1221 B.n69 585
R186 B.n885 B.n884 585
R187 B.n884 B.n65 585
R188 B.n883 B.n64 585
R189 B.n1227 B.n64 585
R190 B.n882 B.n63 585
R191 B.n1228 B.n63 585
R192 B.n881 B.n62 585
R193 B.n1229 B.n62 585
R194 B.n880 B.n879 585
R195 B.n879 B.n61 585
R196 B.n878 B.n57 585
R197 B.n1235 B.n57 585
R198 B.n877 B.n56 585
R199 B.n1236 B.n56 585
R200 B.n876 B.n55 585
R201 B.n1237 B.n55 585
R202 B.n875 B.n874 585
R203 B.n874 B.n51 585
R204 B.n873 B.n50 585
R205 B.n1243 B.n50 585
R206 B.n872 B.n49 585
R207 B.n1244 B.n49 585
R208 B.n871 B.n48 585
R209 B.n1245 B.n48 585
R210 B.n870 B.n869 585
R211 B.n869 B.n44 585
R212 B.n868 B.n43 585
R213 B.n1251 B.n43 585
R214 B.n867 B.n42 585
R215 B.n1252 B.n42 585
R216 B.n866 B.n41 585
R217 B.n1253 B.n41 585
R218 B.n865 B.n864 585
R219 B.n864 B.n40 585
R220 B.n863 B.n36 585
R221 B.n1259 B.n36 585
R222 B.n862 B.n35 585
R223 B.n1260 B.n35 585
R224 B.n861 B.n34 585
R225 B.n1261 B.n34 585
R226 B.n860 B.n859 585
R227 B.n859 B.n30 585
R228 B.n858 B.n29 585
R229 B.n1267 B.n29 585
R230 B.n857 B.n28 585
R231 B.n1268 B.n28 585
R232 B.n856 B.n27 585
R233 B.n1269 B.n27 585
R234 B.n855 B.n854 585
R235 B.n854 B.n23 585
R236 B.n853 B.n22 585
R237 B.n1275 B.n22 585
R238 B.n852 B.n21 585
R239 B.n1276 B.n21 585
R240 B.n851 B.n20 585
R241 B.n1277 B.n20 585
R242 B.n850 B.n849 585
R243 B.n849 B.n19 585
R244 B.n848 B.n15 585
R245 B.n1283 B.n15 585
R246 B.n847 B.n14 585
R247 B.n1284 B.n14 585
R248 B.n846 B.n13 585
R249 B.n1285 B.n13 585
R250 B.n845 B.n844 585
R251 B.n844 B.n12 585
R252 B.n843 B.n842 585
R253 B.n843 B.n8 585
R254 B.n841 B.n7 585
R255 B.n1292 B.n7 585
R256 B.n840 B.n6 585
R257 B.n1293 B.n6 585
R258 B.n839 B.n5 585
R259 B.n1294 B.n5 585
R260 B.n838 B.n837 585
R261 B.n837 B.n4 585
R262 B.n836 B.n198 585
R263 B.n836 B.n835 585
R264 B.n826 B.n199 585
R265 B.n200 B.n199 585
R266 B.n828 B.n827 585
R267 B.n829 B.n828 585
R268 B.n825 B.n205 585
R269 B.n205 B.n204 585
R270 B.n824 B.n823 585
R271 B.n823 B.n822 585
R272 B.n207 B.n206 585
R273 B.n815 B.n207 585
R274 B.n814 B.n813 585
R275 B.n816 B.n814 585
R276 B.n812 B.n212 585
R277 B.n212 B.n211 585
R278 B.n811 B.n810 585
R279 B.n810 B.n809 585
R280 B.n214 B.n213 585
R281 B.n215 B.n214 585
R282 B.n802 B.n801 585
R283 B.n803 B.n802 585
R284 B.n800 B.n220 585
R285 B.n220 B.n219 585
R286 B.n799 B.n798 585
R287 B.n798 B.n797 585
R288 B.n222 B.n221 585
R289 B.n223 B.n222 585
R290 B.n790 B.n789 585
R291 B.n791 B.n790 585
R292 B.n788 B.n228 585
R293 B.n228 B.n227 585
R294 B.n787 B.n786 585
R295 B.n786 B.n785 585
R296 B.n230 B.n229 585
R297 B.n778 B.n230 585
R298 B.n777 B.n776 585
R299 B.n779 B.n777 585
R300 B.n775 B.n235 585
R301 B.n235 B.n234 585
R302 B.n774 B.n773 585
R303 B.n773 B.n772 585
R304 B.n237 B.n236 585
R305 B.n238 B.n237 585
R306 B.n765 B.n764 585
R307 B.n766 B.n765 585
R308 B.n763 B.n243 585
R309 B.n243 B.n242 585
R310 B.n762 B.n761 585
R311 B.n761 B.n760 585
R312 B.n245 B.n244 585
R313 B.n246 B.n245 585
R314 B.n753 B.n752 585
R315 B.n754 B.n753 585
R316 B.n751 B.n251 585
R317 B.n251 B.n250 585
R318 B.n750 B.n749 585
R319 B.n749 B.n748 585
R320 B.n253 B.n252 585
R321 B.n741 B.n253 585
R322 B.n740 B.n739 585
R323 B.n742 B.n740 585
R324 B.n738 B.n258 585
R325 B.n258 B.n257 585
R326 B.n737 B.n736 585
R327 B.n736 B.n735 585
R328 B.n260 B.n259 585
R329 B.n261 B.n260 585
R330 B.n728 B.n727 585
R331 B.n729 B.n728 585
R332 B.n726 B.n266 585
R333 B.n266 B.n265 585
R334 B.n725 B.n724 585
R335 B.n724 B.n723 585
R336 B.n268 B.n267 585
R337 B.n269 B.n268 585
R338 B.n716 B.n715 585
R339 B.n717 B.n716 585
R340 B.n714 B.n274 585
R341 B.n274 B.n273 585
R342 B.n713 B.n712 585
R343 B.n712 B.n711 585
R344 B.n276 B.n275 585
R345 B.n704 B.n276 585
R346 B.n703 B.n702 585
R347 B.n705 B.n703 585
R348 B.n701 B.n281 585
R349 B.n281 B.n280 585
R350 B.n700 B.n699 585
R351 B.n699 B.n698 585
R352 B.n283 B.n282 585
R353 B.n284 B.n283 585
R354 B.n691 B.n690 585
R355 B.n692 B.n691 585
R356 B.n689 B.n289 585
R357 B.n289 B.n288 585
R358 B.n688 B.n687 585
R359 B.n687 B.n686 585
R360 B.n291 B.n290 585
R361 B.n292 B.n291 585
R362 B.n679 B.n678 585
R363 B.n680 B.n679 585
R364 B.n677 B.n297 585
R365 B.n297 B.n296 585
R366 B.n676 B.n675 585
R367 B.n675 B.n674 585
R368 B.n299 B.n298 585
R369 B.n300 B.n299 585
R370 B.n667 B.n666 585
R371 B.n668 B.n667 585
R372 B.n665 B.n305 585
R373 B.n305 B.n304 585
R374 B.n664 B.n663 585
R375 B.n663 B.n662 585
R376 B.n307 B.n306 585
R377 B.n308 B.n307 585
R378 B.n655 B.n654 585
R379 B.n656 B.n655 585
R380 B.n653 B.n313 585
R381 B.n313 B.n312 585
R382 B.n652 B.n651 585
R383 B.n651 B.n650 585
R384 B.n315 B.n314 585
R385 B.n316 B.n315 585
R386 B.n643 B.n642 585
R387 B.n644 B.n643 585
R388 B.n641 B.n321 585
R389 B.n321 B.n320 585
R390 B.n640 B.n639 585
R391 B.n639 B.n638 585
R392 B.n323 B.n322 585
R393 B.n324 B.n323 585
R394 B.n631 B.n630 585
R395 B.n632 B.n631 585
R396 B.n629 B.n328 585
R397 B.n332 B.n328 585
R398 B.n628 B.n627 585
R399 B.n627 B.n626 585
R400 B.n330 B.n329 585
R401 B.n331 B.n330 585
R402 B.n619 B.n618 585
R403 B.n620 B.n619 585
R404 B.n617 B.n337 585
R405 B.n337 B.n336 585
R406 B.n616 B.n615 585
R407 B.n615 B.n614 585
R408 B.n339 B.n338 585
R409 B.n340 B.n339 585
R410 B.n607 B.n606 585
R411 B.n608 B.n607 585
R412 B.n605 B.n345 585
R413 B.n345 B.n344 585
R414 B.n604 B.n603 585
R415 B.n603 B.n602 585
R416 B.n599 B.n349 585
R417 B.n598 B.n597 585
R418 B.n595 B.n350 585
R419 B.n595 B.n348 585
R420 B.n594 B.n593 585
R421 B.n592 B.n591 585
R422 B.n590 B.n352 585
R423 B.n588 B.n587 585
R424 B.n586 B.n353 585
R425 B.n585 B.n584 585
R426 B.n582 B.n354 585
R427 B.n580 B.n579 585
R428 B.n578 B.n355 585
R429 B.n577 B.n576 585
R430 B.n574 B.n356 585
R431 B.n572 B.n571 585
R432 B.n570 B.n357 585
R433 B.n569 B.n568 585
R434 B.n566 B.n358 585
R435 B.n564 B.n563 585
R436 B.n562 B.n359 585
R437 B.n561 B.n560 585
R438 B.n558 B.n360 585
R439 B.n556 B.n555 585
R440 B.n554 B.n361 585
R441 B.n553 B.n552 585
R442 B.n550 B.n362 585
R443 B.n548 B.n547 585
R444 B.n546 B.n363 585
R445 B.n545 B.n544 585
R446 B.n542 B.n364 585
R447 B.n540 B.n539 585
R448 B.n538 B.n365 585
R449 B.n537 B.n536 585
R450 B.n534 B.n366 585
R451 B.n532 B.n531 585
R452 B.n530 B.n367 585
R453 B.n529 B.n528 585
R454 B.n526 B.n368 585
R455 B.n524 B.n523 585
R456 B.n522 B.n369 585
R457 B.n521 B.n520 585
R458 B.n518 B.n370 585
R459 B.n516 B.n515 585
R460 B.n514 B.n371 585
R461 B.n513 B.n512 585
R462 B.n510 B.n509 585
R463 B.n508 B.n507 585
R464 B.n506 B.n376 585
R465 B.n504 B.n503 585
R466 B.n502 B.n377 585
R467 B.n501 B.n500 585
R468 B.n498 B.n378 585
R469 B.n496 B.n495 585
R470 B.n494 B.n379 585
R471 B.n492 B.n491 585
R472 B.n489 B.n382 585
R473 B.n487 B.n486 585
R474 B.n485 B.n383 585
R475 B.n484 B.n483 585
R476 B.n481 B.n384 585
R477 B.n479 B.n478 585
R478 B.n477 B.n385 585
R479 B.n476 B.n475 585
R480 B.n473 B.n386 585
R481 B.n471 B.n470 585
R482 B.n469 B.n387 585
R483 B.n468 B.n467 585
R484 B.n465 B.n388 585
R485 B.n463 B.n462 585
R486 B.n461 B.n389 585
R487 B.n460 B.n459 585
R488 B.n457 B.n390 585
R489 B.n455 B.n454 585
R490 B.n453 B.n391 585
R491 B.n452 B.n451 585
R492 B.n449 B.n392 585
R493 B.n447 B.n446 585
R494 B.n445 B.n393 585
R495 B.n444 B.n443 585
R496 B.n441 B.n394 585
R497 B.n439 B.n438 585
R498 B.n437 B.n395 585
R499 B.n436 B.n435 585
R500 B.n433 B.n396 585
R501 B.n431 B.n430 585
R502 B.n429 B.n397 585
R503 B.n428 B.n427 585
R504 B.n425 B.n398 585
R505 B.n423 B.n422 585
R506 B.n421 B.n399 585
R507 B.n420 B.n419 585
R508 B.n417 B.n400 585
R509 B.n415 B.n414 585
R510 B.n413 B.n401 585
R511 B.n412 B.n411 585
R512 B.n409 B.n402 585
R513 B.n407 B.n406 585
R514 B.n405 B.n404 585
R515 B.n347 B.n346 585
R516 B.n601 B.n600 585
R517 B.n602 B.n601 585
R518 B.n343 B.n342 585
R519 B.n344 B.n343 585
R520 B.n610 B.n609 585
R521 B.n609 B.n608 585
R522 B.n611 B.n341 585
R523 B.n341 B.n340 585
R524 B.n613 B.n612 585
R525 B.n614 B.n613 585
R526 B.n335 B.n334 585
R527 B.n336 B.n335 585
R528 B.n622 B.n621 585
R529 B.n621 B.n620 585
R530 B.n623 B.n333 585
R531 B.n333 B.n331 585
R532 B.n625 B.n624 585
R533 B.n626 B.n625 585
R534 B.n327 B.n326 585
R535 B.n332 B.n327 585
R536 B.n634 B.n633 585
R537 B.n633 B.n632 585
R538 B.n635 B.n325 585
R539 B.n325 B.n324 585
R540 B.n637 B.n636 585
R541 B.n638 B.n637 585
R542 B.n319 B.n318 585
R543 B.n320 B.n319 585
R544 B.n646 B.n645 585
R545 B.n645 B.n644 585
R546 B.n647 B.n317 585
R547 B.n317 B.n316 585
R548 B.n649 B.n648 585
R549 B.n650 B.n649 585
R550 B.n311 B.n310 585
R551 B.n312 B.n311 585
R552 B.n658 B.n657 585
R553 B.n657 B.n656 585
R554 B.n659 B.n309 585
R555 B.n309 B.n308 585
R556 B.n661 B.n660 585
R557 B.n662 B.n661 585
R558 B.n303 B.n302 585
R559 B.n304 B.n303 585
R560 B.n670 B.n669 585
R561 B.n669 B.n668 585
R562 B.n671 B.n301 585
R563 B.n301 B.n300 585
R564 B.n673 B.n672 585
R565 B.n674 B.n673 585
R566 B.n295 B.n294 585
R567 B.n296 B.n295 585
R568 B.n682 B.n681 585
R569 B.n681 B.n680 585
R570 B.n683 B.n293 585
R571 B.n293 B.n292 585
R572 B.n685 B.n684 585
R573 B.n686 B.n685 585
R574 B.n287 B.n286 585
R575 B.n288 B.n287 585
R576 B.n694 B.n693 585
R577 B.n693 B.n692 585
R578 B.n695 B.n285 585
R579 B.n285 B.n284 585
R580 B.n697 B.n696 585
R581 B.n698 B.n697 585
R582 B.n279 B.n278 585
R583 B.n280 B.n279 585
R584 B.n707 B.n706 585
R585 B.n706 B.n705 585
R586 B.n708 B.n277 585
R587 B.n704 B.n277 585
R588 B.n710 B.n709 585
R589 B.n711 B.n710 585
R590 B.n272 B.n271 585
R591 B.n273 B.n272 585
R592 B.n719 B.n718 585
R593 B.n718 B.n717 585
R594 B.n720 B.n270 585
R595 B.n270 B.n269 585
R596 B.n722 B.n721 585
R597 B.n723 B.n722 585
R598 B.n264 B.n263 585
R599 B.n265 B.n264 585
R600 B.n731 B.n730 585
R601 B.n730 B.n729 585
R602 B.n732 B.n262 585
R603 B.n262 B.n261 585
R604 B.n734 B.n733 585
R605 B.n735 B.n734 585
R606 B.n256 B.n255 585
R607 B.n257 B.n256 585
R608 B.n744 B.n743 585
R609 B.n743 B.n742 585
R610 B.n745 B.n254 585
R611 B.n741 B.n254 585
R612 B.n747 B.n746 585
R613 B.n748 B.n747 585
R614 B.n249 B.n248 585
R615 B.n250 B.n249 585
R616 B.n756 B.n755 585
R617 B.n755 B.n754 585
R618 B.n757 B.n247 585
R619 B.n247 B.n246 585
R620 B.n759 B.n758 585
R621 B.n760 B.n759 585
R622 B.n241 B.n240 585
R623 B.n242 B.n241 585
R624 B.n768 B.n767 585
R625 B.n767 B.n766 585
R626 B.n769 B.n239 585
R627 B.n239 B.n238 585
R628 B.n771 B.n770 585
R629 B.n772 B.n771 585
R630 B.n233 B.n232 585
R631 B.n234 B.n233 585
R632 B.n781 B.n780 585
R633 B.n780 B.n779 585
R634 B.n782 B.n231 585
R635 B.n778 B.n231 585
R636 B.n784 B.n783 585
R637 B.n785 B.n784 585
R638 B.n226 B.n225 585
R639 B.n227 B.n226 585
R640 B.n793 B.n792 585
R641 B.n792 B.n791 585
R642 B.n794 B.n224 585
R643 B.n224 B.n223 585
R644 B.n796 B.n795 585
R645 B.n797 B.n796 585
R646 B.n218 B.n217 585
R647 B.n219 B.n218 585
R648 B.n805 B.n804 585
R649 B.n804 B.n803 585
R650 B.n806 B.n216 585
R651 B.n216 B.n215 585
R652 B.n808 B.n807 585
R653 B.n809 B.n808 585
R654 B.n210 B.n209 585
R655 B.n211 B.n210 585
R656 B.n818 B.n817 585
R657 B.n817 B.n816 585
R658 B.n819 B.n208 585
R659 B.n815 B.n208 585
R660 B.n821 B.n820 585
R661 B.n822 B.n821 585
R662 B.n203 B.n202 585
R663 B.n204 B.n203 585
R664 B.n831 B.n830 585
R665 B.n830 B.n829 585
R666 B.n832 B.n201 585
R667 B.n201 B.n200 585
R668 B.n834 B.n833 585
R669 B.n835 B.n834 585
R670 B.n3 B.n0 585
R671 B.n4 B.n3 585
R672 B.n1291 B.n1 585
R673 B.n1292 B.n1291 585
R674 B.n1290 B.n1289 585
R675 B.n1290 B.n8 585
R676 B.n1288 B.n9 585
R677 B.n12 B.n9 585
R678 B.n1287 B.n1286 585
R679 B.n1286 B.n1285 585
R680 B.n11 B.n10 585
R681 B.n1284 B.n11 585
R682 B.n1282 B.n1281 585
R683 B.n1283 B.n1282 585
R684 B.n1280 B.n16 585
R685 B.n19 B.n16 585
R686 B.n1279 B.n1278 585
R687 B.n1278 B.n1277 585
R688 B.n18 B.n17 585
R689 B.n1276 B.n18 585
R690 B.n1274 B.n1273 585
R691 B.n1275 B.n1274 585
R692 B.n1272 B.n24 585
R693 B.n24 B.n23 585
R694 B.n1271 B.n1270 585
R695 B.n1270 B.n1269 585
R696 B.n26 B.n25 585
R697 B.n1268 B.n26 585
R698 B.n1266 B.n1265 585
R699 B.n1267 B.n1266 585
R700 B.n1264 B.n31 585
R701 B.n31 B.n30 585
R702 B.n1263 B.n1262 585
R703 B.n1262 B.n1261 585
R704 B.n33 B.n32 585
R705 B.n1260 B.n33 585
R706 B.n1258 B.n1257 585
R707 B.n1259 B.n1258 585
R708 B.n1256 B.n37 585
R709 B.n40 B.n37 585
R710 B.n1255 B.n1254 585
R711 B.n1254 B.n1253 585
R712 B.n39 B.n38 585
R713 B.n1252 B.n39 585
R714 B.n1250 B.n1249 585
R715 B.n1251 B.n1250 585
R716 B.n1248 B.n45 585
R717 B.n45 B.n44 585
R718 B.n1247 B.n1246 585
R719 B.n1246 B.n1245 585
R720 B.n47 B.n46 585
R721 B.n1244 B.n47 585
R722 B.n1242 B.n1241 585
R723 B.n1243 B.n1242 585
R724 B.n1240 B.n52 585
R725 B.n52 B.n51 585
R726 B.n1239 B.n1238 585
R727 B.n1238 B.n1237 585
R728 B.n54 B.n53 585
R729 B.n1236 B.n54 585
R730 B.n1234 B.n1233 585
R731 B.n1235 B.n1234 585
R732 B.n1232 B.n58 585
R733 B.n61 B.n58 585
R734 B.n1231 B.n1230 585
R735 B.n1230 B.n1229 585
R736 B.n60 B.n59 585
R737 B.n1228 B.n60 585
R738 B.n1226 B.n1225 585
R739 B.n1227 B.n1226 585
R740 B.n1224 B.n66 585
R741 B.n66 B.n65 585
R742 B.n1223 B.n1222 585
R743 B.n1222 B.n1221 585
R744 B.n68 B.n67 585
R745 B.n1220 B.n68 585
R746 B.n1218 B.n1217 585
R747 B.n1219 B.n1218 585
R748 B.n1216 B.n73 585
R749 B.n73 B.n72 585
R750 B.n1215 B.n1214 585
R751 B.n1214 B.n1213 585
R752 B.n75 B.n74 585
R753 B.n1212 B.n75 585
R754 B.n1210 B.n1209 585
R755 B.n1211 B.n1210 585
R756 B.n1208 B.n79 585
R757 B.n82 B.n79 585
R758 B.n1207 B.n1206 585
R759 B.n1206 B.n1205 585
R760 B.n81 B.n80 585
R761 B.n1204 B.n81 585
R762 B.n1202 B.n1201 585
R763 B.n1203 B.n1202 585
R764 B.n1200 B.n87 585
R765 B.n87 B.n86 585
R766 B.n1199 B.n1198 585
R767 B.n1198 B.n1197 585
R768 B.n89 B.n88 585
R769 B.n1196 B.n89 585
R770 B.n1194 B.n1193 585
R771 B.n1195 B.n1194 585
R772 B.n1192 B.n94 585
R773 B.n94 B.n93 585
R774 B.n1191 B.n1190 585
R775 B.n1190 B.n1189 585
R776 B.n96 B.n95 585
R777 B.n1188 B.n96 585
R778 B.n1186 B.n1185 585
R779 B.n1187 B.n1186 585
R780 B.n1184 B.n101 585
R781 B.n101 B.n100 585
R782 B.n1183 B.n1182 585
R783 B.n1182 B.n1181 585
R784 B.n103 B.n102 585
R785 B.n1180 B.n103 585
R786 B.n1178 B.n1177 585
R787 B.n1179 B.n1178 585
R788 B.n1176 B.n108 585
R789 B.n108 B.n107 585
R790 B.n1175 B.n1174 585
R791 B.n1174 B.n1173 585
R792 B.n110 B.n109 585
R793 B.n1172 B.n110 585
R794 B.n1170 B.n1169 585
R795 B.n1171 B.n1170 585
R796 B.n1168 B.n115 585
R797 B.n115 B.n114 585
R798 B.n1167 B.n1166 585
R799 B.n1166 B.n1165 585
R800 B.n117 B.n116 585
R801 B.n1164 B.n117 585
R802 B.n1162 B.n1161 585
R803 B.n1163 B.n1162 585
R804 B.n1160 B.n122 585
R805 B.n122 B.n121 585
R806 B.n1159 B.n1158 585
R807 B.n1158 B.n1157 585
R808 B.n124 B.n123 585
R809 B.n1156 B.n124 585
R810 B.n1154 B.n1153 585
R811 B.n1155 B.n1154 585
R812 B.n1152 B.n129 585
R813 B.n129 B.n128 585
R814 B.n1151 B.n1150 585
R815 B.n1150 B.n1149 585
R816 B.n131 B.n130 585
R817 B.n1148 B.n131 585
R818 B.n1146 B.n1145 585
R819 B.n1147 B.n1146 585
R820 B.n1144 B.n136 585
R821 B.n136 B.n135 585
R822 B.n1143 B.n1142 585
R823 B.n1142 B.n1141 585
R824 B.n138 B.n137 585
R825 B.n1140 B.n138 585
R826 B.n1138 B.n1137 585
R827 B.n1139 B.n1138 585
R828 B.n1295 B.n1294 585
R829 B.n1293 B.n2 585
R830 B.n1138 B.n143 454.062
R831 B.n197 B.n141 454.062
R832 B.n603 B.n347 454.062
R833 B.n601 B.n349 454.062
R834 B.n166 B.t10 295.125
R835 B.n172 B.t14 295.125
R836 B.n380 B.t17 295.125
R837 B.n372 B.t21 295.125
R838 B.n942 B.n142 256.663
R839 B.n944 B.n142 256.663
R840 B.n950 B.n142 256.663
R841 B.n952 B.n142 256.663
R842 B.n958 B.n142 256.663
R843 B.n960 B.n142 256.663
R844 B.n966 B.n142 256.663
R845 B.n968 B.n142 256.663
R846 B.n974 B.n142 256.663
R847 B.n976 B.n142 256.663
R848 B.n982 B.n142 256.663
R849 B.n984 B.n142 256.663
R850 B.n990 B.n142 256.663
R851 B.n992 B.n142 256.663
R852 B.n998 B.n142 256.663
R853 B.n1000 B.n142 256.663
R854 B.n1006 B.n142 256.663
R855 B.n1008 B.n142 256.663
R856 B.n1014 B.n142 256.663
R857 B.n1016 B.n142 256.663
R858 B.n1022 B.n142 256.663
R859 B.n175 B.n142 256.663
R860 B.n1028 B.n142 256.663
R861 B.n1034 B.n142 256.663
R862 B.n1036 B.n142 256.663
R863 B.n1042 B.n142 256.663
R864 B.n1044 B.n142 256.663
R865 B.n1051 B.n142 256.663
R866 B.n1053 B.n142 256.663
R867 B.n1059 B.n142 256.663
R868 B.n1061 B.n142 256.663
R869 B.n1067 B.n142 256.663
R870 B.n1069 B.n142 256.663
R871 B.n1075 B.n142 256.663
R872 B.n1077 B.n142 256.663
R873 B.n1083 B.n142 256.663
R874 B.n1085 B.n142 256.663
R875 B.n1091 B.n142 256.663
R876 B.n1093 B.n142 256.663
R877 B.n1099 B.n142 256.663
R878 B.n1101 B.n142 256.663
R879 B.n1107 B.n142 256.663
R880 B.n1109 B.n142 256.663
R881 B.n1115 B.n142 256.663
R882 B.n1117 B.n142 256.663
R883 B.n1123 B.n142 256.663
R884 B.n1125 B.n142 256.663
R885 B.n1131 B.n142 256.663
R886 B.n1133 B.n142 256.663
R887 B.n596 B.n348 256.663
R888 B.n351 B.n348 256.663
R889 B.n589 B.n348 256.663
R890 B.n583 B.n348 256.663
R891 B.n581 B.n348 256.663
R892 B.n575 B.n348 256.663
R893 B.n573 B.n348 256.663
R894 B.n567 B.n348 256.663
R895 B.n565 B.n348 256.663
R896 B.n559 B.n348 256.663
R897 B.n557 B.n348 256.663
R898 B.n551 B.n348 256.663
R899 B.n549 B.n348 256.663
R900 B.n543 B.n348 256.663
R901 B.n541 B.n348 256.663
R902 B.n535 B.n348 256.663
R903 B.n533 B.n348 256.663
R904 B.n527 B.n348 256.663
R905 B.n525 B.n348 256.663
R906 B.n519 B.n348 256.663
R907 B.n517 B.n348 256.663
R908 B.n511 B.n348 256.663
R909 B.n375 B.n348 256.663
R910 B.n505 B.n348 256.663
R911 B.n499 B.n348 256.663
R912 B.n497 B.n348 256.663
R913 B.n490 B.n348 256.663
R914 B.n488 B.n348 256.663
R915 B.n482 B.n348 256.663
R916 B.n480 B.n348 256.663
R917 B.n474 B.n348 256.663
R918 B.n472 B.n348 256.663
R919 B.n466 B.n348 256.663
R920 B.n464 B.n348 256.663
R921 B.n458 B.n348 256.663
R922 B.n456 B.n348 256.663
R923 B.n450 B.n348 256.663
R924 B.n448 B.n348 256.663
R925 B.n442 B.n348 256.663
R926 B.n440 B.n348 256.663
R927 B.n434 B.n348 256.663
R928 B.n432 B.n348 256.663
R929 B.n426 B.n348 256.663
R930 B.n424 B.n348 256.663
R931 B.n418 B.n348 256.663
R932 B.n416 B.n348 256.663
R933 B.n410 B.n348 256.663
R934 B.n408 B.n348 256.663
R935 B.n403 B.n348 256.663
R936 B.n1297 B.n1296 256.663
R937 B.n1134 B.n1132 163.367
R938 B.n1130 B.n145 163.367
R939 B.n1126 B.n1124 163.367
R940 B.n1122 B.n147 163.367
R941 B.n1118 B.n1116 163.367
R942 B.n1114 B.n149 163.367
R943 B.n1110 B.n1108 163.367
R944 B.n1106 B.n151 163.367
R945 B.n1102 B.n1100 163.367
R946 B.n1098 B.n153 163.367
R947 B.n1094 B.n1092 163.367
R948 B.n1090 B.n155 163.367
R949 B.n1086 B.n1084 163.367
R950 B.n1082 B.n157 163.367
R951 B.n1078 B.n1076 163.367
R952 B.n1074 B.n159 163.367
R953 B.n1070 B.n1068 163.367
R954 B.n1066 B.n161 163.367
R955 B.n1062 B.n1060 163.367
R956 B.n1058 B.n163 163.367
R957 B.n1054 B.n1052 163.367
R958 B.n1050 B.n165 163.367
R959 B.n1045 B.n1043 163.367
R960 B.n1041 B.n169 163.367
R961 B.n1037 B.n1035 163.367
R962 B.n1033 B.n171 163.367
R963 B.n1029 B.n1027 163.367
R964 B.n1024 B.n1023 163.367
R965 B.n1021 B.n177 163.367
R966 B.n1017 B.n1015 163.367
R967 B.n1013 B.n179 163.367
R968 B.n1009 B.n1007 163.367
R969 B.n1005 B.n181 163.367
R970 B.n1001 B.n999 163.367
R971 B.n997 B.n183 163.367
R972 B.n993 B.n991 163.367
R973 B.n989 B.n185 163.367
R974 B.n985 B.n983 163.367
R975 B.n981 B.n187 163.367
R976 B.n977 B.n975 163.367
R977 B.n973 B.n189 163.367
R978 B.n969 B.n967 163.367
R979 B.n965 B.n191 163.367
R980 B.n961 B.n959 163.367
R981 B.n957 B.n193 163.367
R982 B.n953 B.n951 163.367
R983 B.n949 B.n195 163.367
R984 B.n945 B.n943 163.367
R985 B.n941 B.n197 163.367
R986 B.n603 B.n345 163.367
R987 B.n607 B.n345 163.367
R988 B.n607 B.n339 163.367
R989 B.n615 B.n339 163.367
R990 B.n615 B.n337 163.367
R991 B.n619 B.n337 163.367
R992 B.n619 B.n330 163.367
R993 B.n627 B.n330 163.367
R994 B.n627 B.n328 163.367
R995 B.n631 B.n328 163.367
R996 B.n631 B.n323 163.367
R997 B.n639 B.n323 163.367
R998 B.n639 B.n321 163.367
R999 B.n643 B.n321 163.367
R1000 B.n643 B.n315 163.367
R1001 B.n651 B.n315 163.367
R1002 B.n651 B.n313 163.367
R1003 B.n655 B.n313 163.367
R1004 B.n655 B.n307 163.367
R1005 B.n663 B.n307 163.367
R1006 B.n663 B.n305 163.367
R1007 B.n667 B.n305 163.367
R1008 B.n667 B.n299 163.367
R1009 B.n675 B.n299 163.367
R1010 B.n675 B.n297 163.367
R1011 B.n679 B.n297 163.367
R1012 B.n679 B.n291 163.367
R1013 B.n687 B.n291 163.367
R1014 B.n687 B.n289 163.367
R1015 B.n691 B.n289 163.367
R1016 B.n691 B.n283 163.367
R1017 B.n699 B.n283 163.367
R1018 B.n699 B.n281 163.367
R1019 B.n703 B.n281 163.367
R1020 B.n703 B.n276 163.367
R1021 B.n712 B.n276 163.367
R1022 B.n712 B.n274 163.367
R1023 B.n716 B.n274 163.367
R1024 B.n716 B.n268 163.367
R1025 B.n724 B.n268 163.367
R1026 B.n724 B.n266 163.367
R1027 B.n728 B.n266 163.367
R1028 B.n728 B.n260 163.367
R1029 B.n736 B.n260 163.367
R1030 B.n736 B.n258 163.367
R1031 B.n740 B.n258 163.367
R1032 B.n740 B.n253 163.367
R1033 B.n749 B.n253 163.367
R1034 B.n749 B.n251 163.367
R1035 B.n753 B.n251 163.367
R1036 B.n753 B.n245 163.367
R1037 B.n761 B.n245 163.367
R1038 B.n761 B.n243 163.367
R1039 B.n765 B.n243 163.367
R1040 B.n765 B.n237 163.367
R1041 B.n773 B.n237 163.367
R1042 B.n773 B.n235 163.367
R1043 B.n777 B.n235 163.367
R1044 B.n777 B.n230 163.367
R1045 B.n786 B.n230 163.367
R1046 B.n786 B.n228 163.367
R1047 B.n790 B.n228 163.367
R1048 B.n790 B.n222 163.367
R1049 B.n798 B.n222 163.367
R1050 B.n798 B.n220 163.367
R1051 B.n802 B.n220 163.367
R1052 B.n802 B.n214 163.367
R1053 B.n810 B.n214 163.367
R1054 B.n810 B.n212 163.367
R1055 B.n814 B.n212 163.367
R1056 B.n814 B.n207 163.367
R1057 B.n823 B.n207 163.367
R1058 B.n823 B.n205 163.367
R1059 B.n828 B.n205 163.367
R1060 B.n828 B.n199 163.367
R1061 B.n836 B.n199 163.367
R1062 B.n837 B.n836 163.367
R1063 B.n837 B.n5 163.367
R1064 B.n6 B.n5 163.367
R1065 B.n7 B.n6 163.367
R1066 B.n843 B.n7 163.367
R1067 B.n844 B.n843 163.367
R1068 B.n844 B.n13 163.367
R1069 B.n14 B.n13 163.367
R1070 B.n15 B.n14 163.367
R1071 B.n849 B.n15 163.367
R1072 B.n849 B.n20 163.367
R1073 B.n21 B.n20 163.367
R1074 B.n22 B.n21 163.367
R1075 B.n854 B.n22 163.367
R1076 B.n854 B.n27 163.367
R1077 B.n28 B.n27 163.367
R1078 B.n29 B.n28 163.367
R1079 B.n859 B.n29 163.367
R1080 B.n859 B.n34 163.367
R1081 B.n35 B.n34 163.367
R1082 B.n36 B.n35 163.367
R1083 B.n864 B.n36 163.367
R1084 B.n864 B.n41 163.367
R1085 B.n42 B.n41 163.367
R1086 B.n43 B.n42 163.367
R1087 B.n869 B.n43 163.367
R1088 B.n869 B.n48 163.367
R1089 B.n49 B.n48 163.367
R1090 B.n50 B.n49 163.367
R1091 B.n874 B.n50 163.367
R1092 B.n874 B.n55 163.367
R1093 B.n56 B.n55 163.367
R1094 B.n57 B.n56 163.367
R1095 B.n879 B.n57 163.367
R1096 B.n879 B.n62 163.367
R1097 B.n63 B.n62 163.367
R1098 B.n64 B.n63 163.367
R1099 B.n884 B.n64 163.367
R1100 B.n884 B.n69 163.367
R1101 B.n70 B.n69 163.367
R1102 B.n71 B.n70 163.367
R1103 B.n889 B.n71 163.367
R1104 B.n889 B.n76 163.367
R1105 B.n77 B.n76 163.367
R1106 B.n78 B.n77 163.367
R1107 B.n894 B.n78 163.367
R1108 B.n894 B.n83 163.367
R1109 B.n84 B.n83 163.367
R1110 B.n85 B.n84 163.367
R1111 B.n899 B.n85 163.367
R1112 B.n899 B.n90 163.367
R1113 B.n91 B.n90 163.367
R1114 B.n92 B.n91 163.367
R1115 B.n904 B.n92 163.367
R1116 B.n904 B.n97 163.367
R1117 B.n98 B.n97 163.367
R1118 B.n99 B.n98 163.367
R1119 B.n909 B.n99 163.367
R1120 B.n909 B.n104 163.367
R1121 B.n105 B.n104 163.367
R1122 B.n106 B.n105 163.367
R1123 B.n914 B.n106 163.367
R1124 B.n914 B.n111 163.367
R1125 B.n112 B.n111 163.367
R1126 B.n113 B.n112 163.367
R1127 B.n919 B.n113 163.367
R1128 B.n919 B.n118 163.367
R1129 B.n119 B.n118 163.367
R1130 B.n120 B.n119 163.367
R1131 B.n924 B.n120 163.367
R1132 B.n924 B.n125 163.367
R1133 B.n126 B.n125 163.367
R1134 B.n127 B.n126 163.367
R1135 B.n929 B.n127 163.367
R1136 B.n929 B.n132 163.367
R1137 B.n133 B.n132 163.367
R1138 B.n134 B.n133 163.367
R1139 B.n934 B.n134 163.367
R1140 B.n934 B.n139 163.367
R1141 B.n140 B.n139 163.367
R1142 B.n141 B.n140 163.367
R1143 B.n597 B.n595 163.367
R1144 B.n595 B.n594 163.367
R1145 B.n591 B.n590 163.367
R1146 B.n588 B.n353 163.367
R1147 B.n584 B.n582 163.367
R1148 B.n580 B.n355 163.367
R1149 B.n576 B.n574 163.367
R1150 B.n572 B.n357 163.367
R1151 B.n568 B.n566 163.367
R1152 B.n564 B.n359 163.367
R1153 B.n560 B.n558 163.367
R1154 B.n556 B.n361 163.367
R1155 B.n552 B.n550 163.367
R1156 B.n548 B.n363 163.367
R1157 B.n544 B.n542 163.367
R1158 B.n540 B.n365 163.367
R1159 B.n536 B.n534 163.367
R1160 B.n532 B.n367 163.367
R1161 B.n528 B.n526 163.367
R1162 B.n524 B.n369 163.367
R1163 B.n520 B.n518 163.367
R1164 B.n516 B.n371 163.367
R1165 B.n512 B.n510 163.367
R1166 B.n507 B.n506 163.367
R1167 B.n504 B.n377 163.367
R1168 B.n500 B.n498 163.367
R1169 B.n496 B.n379 163.367
R1170 B.n491 B.n489 163.367
R1171 B.n487 B.n383 163.367
R1172 B.n483 B.n481 163.367
R1173 B.n479 B.n385 163.367
R1174 B.n475 B.n473 163.367
R1175 B.n471 B.n387 163.367
R1176 B.n467 B.n465 163.367
R1177 B.n463 B.n389 163.367
R1178 B.n459 B.n457 163.367
R1179 B.n455 B.n391 163.367
R1180 B.n451 B.n449 163.367
R1181 B.n447 B.n393 163.367
R1182 B.n443 B.n441 163.367
R1183 B.n439 B.n395 163.367
R1184 B.n435 B.n433 163.367
R1185 B.n431 B.n397 163.367
R1186 B.n427 B.n425 163.367
R1187 B.n423 B.n399 163.367
R1188 B.n419 B.n417 163.367
R1189 B.n415 B.n401 163.367
R1190 B.n411 B.n409 163.367
R1191 B.n407 B.n404 163.367
R1192 B.n601 B.n343 163.367
R1193 B.n609 B.n343 163.367
R1194 B.n609 B.n341 163.367
R1195 B.n613 B.n341 163.367
R1196 B.n613 B.n335 163.367
R1197 B.n621 B.n335 163.367
R1198 B.n621 B.n333 163.367
R1199 B.n625 B.n333 163.367
R1200 B.n625 B.n327 163.367
R1201 B.n633 B.n327 163.367
R1202 B.n633 B.n325 163.367
R1203 B.n637 B.n325 163.367
R1204 B.n637 B.n319 163.367
R1205 B.n645 B.n319 163.367
R1206 B.n645 B.n317 163.367
R1207 B.n649 B.n317 163.367
R1208 B.n649 B.n311 163.367
R1209 B.n657 B.n311 163.367
R1210 B.n657 B.n309 163.367
R1211 B.n661 B.n309 163.367
R1212 B.n661 B.n303 163.367
R1213 B.n669 B.n303 163.367
R1214 B.n669 B.n301 163.367
R1215 B.n673 B.n301 163.367
R1216 B.n673 B.n295 163.367
R1217 B.n681 B.n295 163.367
R1218 B.n681 B.n293 163.367
R1219 B.n685 B.n293 163.367
R1220 B.n685 B.n287 163.367
R1221 B.n693 B.n287 163.367
R1222 B.n693 B.n285 163.367
R1223 B.n697 B.n285 163.367
R1224 B.n697 B.n279 163.367
R1225 B.n706 B.n279 163.367
R1226 B.n706 B.n277 163.367
R1227 B.n710 B.n277 163.367
R1228 B.n710 B.n272 163.367
R1229 B.n718 B.n272 163.367
R1230 B.n718 B.n270 163.367
R1231 B.n722 B.n270 163.367
R1232 B.n722 B.n264 163.367
R1233 B.n730 B.n264 163.367
R1234 B.n730 B.n262 163.367
R1235 B.n734 B.n262 163.367
R1236 B.n734 B.n256 163.367
R1237 B.n743 B.n256 163.367
R1238 B.n743 B.n254 163.367
R1239 B.n747 B.n254 163.367
R1240 B.n747 B.n249 163.367
R1241 B.n755 B.n249 163.367
R1242 B.n755 B.n247 163.367
R1243 B.n759 B.n247 163.367
R1244 B.n759 B.n241 163.367
R1245 B.n767 B.n241 163.367
R1246 B.n767 B.n239 163.367
R1247 B.n771 B.n239 163.367
R1248 B.n771 B.n233 163.367
R1249 B.n780 B.n233 163.367
R1250 B.n780 B.n231 163.367
R1251 B.n784 B.n231 163.367
R1252 B.n784 B.n226 163.367
R1253 B.n792 B.n226 163.367
R1254 B.n792 B.n224 163.367
R1255 B.n796 B.n224 163.367
R1256 B.n796 B.n218 163.367
R1257 B.n804 B.n218 163.367
R1258 B.n804 B.n216 163.367
R1259 B.n808 B.n216 163.367
R1260 B.n808 B.n210 163.367
R1261 B.n817 B.n210 163.367
R1262 B.n817 B.n208 163.367
R1263 B.n821 B.n208 163.367
R1264 B.n821 B.n203 163.367
R1265 B.n830 B.n203 163.367
R1266 B.n830 B.n201 163.367
R1267 B.n834 B.n201 163.367
R1268 B.n834 B.n3 163.367
R1269 B.n1295 B.n3 163.367
R1270 B.n1291 B.n2 163.367
R1271 B.n1291 B.n1290 163.367
R1272 B.n1290 B.n9 163.367
R1273 B.n1286 B.n9 163.367
R1274 B.n1286 B.n11 163.367
R1275 B.n1282 B.n11 163.367
R1276 B.n1282 B.n16 163.367
R1277 B.n1278 B.n16 163.367
R1278 B.n1278 B.n18 163.367
R1279 B.n1274 B.n18 163.367
R1280 B.n1274 B.n24 163.367
R1281 B.n1270 B.n24 163.367
R1282 B.n1270 B.n26 163.367
R1283 B.n1266 B.n26 163.367
R1284 B.n1266 B.n31 163.367
R1285 B.n1262 B.n31 163.367
R1286 B.n1262 B.n33 163.367
R1287 B.n1258 B.n33 163.367
R1288 B.n1258 B.n37 163.367
R1289 B.n1254 B.n37 163.367
R1290 B.n1254 B.n39 163.367
R1291 B.n1250 B.n39 163.367
R1292 B.n1250 B.n45 163.367
R1293 B.n1246 B.n45 163.367
R1294 B.n1246 B.n47 163.367
R1295 B.n1242 B.n47 163.367
R1296 B.n1242 B.n52 163.367
R1297 B.n1238 B.n52 163.367
R1298 B.n1238 B.n54 163.367
R1299 B.n1234 B.n54 163.367
R1300 B.n1234 B.n58 163.367
R1301 B.n1230 B.n58 163.367
R1302 B.n1230 B.n60 163.367
R1303 B.n1226 B.n60 163.367
R1304 B.n1226 B.n66 163.367
R1305 B.n1222 B.n66 163.367
R1306 B.n1222 B.n68 163.367
R1307 B.n1218 B.n68 163.367
R1308 B.n1218 B.n73 163.367
R1309 B.n1214 B.n73 163.367
R1310 B.n1214 B.n75 163.367
R1311 B.n1210 B.n75 163.367
R1312 B.n1210 B.n79 163.367
R1313 B.n1206 B.n79 163.367
R1314 B.n1206 B.n81 163.367
R1315 B.n1202 B.n81 163.367
R1316 B.n1202 B.n87 163.367
R1317 B.n1198 B.n87 163.367
R1318 B.n1198 B.n89 163.367
R1319 B.n1194 B.n89 163.367
R1320 B.n1194 B.n94 163.367
R1321 B.n1190 B.n94 163.367
R1322 B.n1190 B.n96 163.367
R1323 B.n1186 B.n96 163.367
R1324 B.n1186 B.n101 163.367
R1325 B.n1182 B.n101 163.367
R1326 B.n1182 B.n103 163.367
R1327 B.n1178 B.n103 163.367
R1328 B.n1178 B.n108 163.367
R1329 B.n1174 B.n108 163.367
R1330 B.n1174 B.n110 163.367
R1331 B.n1170 B.n110 163.367
R1332 B.n1170 B.n115 163.367
R1333 B.n1166 B.n115 163.367
R1334 B.n1166 B.n117 163.367
R1335 B.n1162 B.n117 163.367
R1336 B.n1162 B.n122 163.367
R1337 B.n1158 B.n122 163.367
R1338 B.n1158 B.n124 163.367
R1339 B.n1154 B.n124 163.367
R1340 B.n1154 B.n129 163.367
R1341 B.n1150 B.n129 163.367
R1342 B.n1150 B.n131 163.367
R1343 B.n1146 B.n131 163.367
R1344 B.n1146 B.n136 163.367
R1345 B.n1142 B.n136 163.367
R1346 B.n1142 B.n138 163.367
R1347 B.n1138 B.n138 163.367
R1348 B.n172 B.t15 146.596
R1349 B.n380 B.t20 146.596
R1350 B.n166 B.t12 146.579
R1351 B.n372 B.t23 146.579
R1352 B.n167 B.n166 77.1884
R1353 B.n173 B.n172 77.1884
R1354 B.n381 B.n380 77.1884
R1355 B.n373 B.n372 77.1884
R1356 B.n1133 B.n143 71.676
R1357 B.n1132 B.n1131 71.676
R1358 B.n1125 B.n145 71.676
R1359 B.n1124 B.n1123 71.676
R1360 B.n1117 B.n147 71.676
R1361 B.n1116 B.n1115 71.676
R1362 B.n1109 B.n149 71.676
R1363 B.n1108 B.n1107 71.676
R1364 B.n1101 B.n151 71.676
R1365 B.n1100 B.n1099 71.676
R1366 B.n1093 B.n153 71.676
R1367 B.n1092 B.n1091 71.676
R1368 B.n1085 B.n155 71.676
R1369 B.n1084 B.n1083 71.676
R1370 B.n1077 B.n157 71.676
R1371 B.n1076 B.n1075 71.676
R1372 B.n1069 B.n159 71.676
R1373 B.n1068 B.n1067 71.676
R1374 B.n1061 B.n161 71.676
R1375 B.n1060 B.n1059 71.676
R1376 B.n1053 B.n163 71.676
R1377 B.n1052 B.n1051 71.676
R1378 B.n1044 B.n165 71.676
R1379 B.n1043 B.n1042 71.676
R1380 B.n1036 B.n169 71.676
R1381 B.n1035 B.n1034 71.676
R1382 B.n1028 B.n171 71.676
R1383 B.n1027 B.n175 71.676
R1384 B.n1023 B.n1022 71.676
R1385 B.n1016 B.n177 71.676
R1386 B.n1015 B.n1014 71.676
R1387 B.n1008 B.n179 71.676
R1388 B.n1007 B.n1006 71.676
R1389 B.n1000 B.n181 71.676
R1390 B.n999 B.n998 71.676
R1391 B.n992 B.n183 71.676
R1392 B.n991 B.n990 71.676
R1393 B.n984 B.n185 71.676
R1394 B.n983 B.n982 71.676
R1395 B.n976 B.n187 71.676
R1396 B.n975 B.n974 71.676
R1397 B.n968 B.n189 71.676
R1398 B.n967 B.n966 71.676
R1399 B.n960 B.n191 71.676
R1400 B.n959 B.n958 71.676
R1401 B.n952 B.n193 71.676
R1402 B.n951 B.n950 71.676
R1403 B.n944 B.n195 71.676
R1404 B.n943 B.n942 71.676
R1405 B.n942 B.n941 71.676
R1406 B.n945 B.n944 71.676
R1407 B.n950 B.n949 71.676
R1408 B.n953 B.n952 71.676
R1409 B.n958 B.n957 71.676
R1410 B.n961 B.n960 71.676
R1411 B.n966 B.n965 71.676
R1412 B.n969 B.n968 71.676
R1413 B.n974 B.n973 71.676
R1414 B.n977 B.n976 71.676
R1415 B.n982 B.n981 71.676
R1416 B.n985 B.n984 71.676
R1417 B.n990 B.n989 71.676
R1418 B.n993 B.n992 71.676
R1419 B.n998 B.n997 71.676
R1420 B.n1001 B.n1000 71.676
R1421 B.n1006 B.n1005 71.676
R1422 B.n1009 B.n1008 71.676
R1423 B.n1014 B.n1013 71.676
R1424 B.n1017 B.n1016 71.676
R1425 B.n1022 B.n1021 71.676
R1426 B.n1024 B.n175 71.676
R1427 B.n1029 B.n1028 71.676
R1428 B.n1034 B.n1033 71.676
R1429 B.n1037 B.n1036 71.676
R1430 B.n1042 B.n1041 71.676
R1431 B.n1045 B.n1044 71.676
R1432 B.n1051 B.n1050 71.676
R1433 B.n1054 B.n1053 71.676
R1434 B.n1059 B.n1058 71.676
R1435 B.n1062 B.n1061 71.676
R1436 B.n1067 B.n1066 71.676
R1437 B.n1070 B.n1069 71.676
R1438 B.n1075 B.n1074 71.676
R1439 B.n1078 B.n1077 71.676
R1440 B.n1083 B.n1082 71.676
R1441 B.n1086 B.n1085 71.676
R1442 B.n1091 B.n1090 71.676
R1443 B.n1094 B.n1093 71.676
R1444 B.n1099 B.n1098 71.676
R1445 B.n1102 B.n1101 71.676
R1446 B.n1107 B.n1106 71.676
R1447 B.n1110 B.n1109 71.676
R1448 B.n1115 B.n1114 71.676
R1449 B.n1118 B.n1117 71.676
R1450 B.n1123 B.n1122 71.676
R1451 B.n1126 B.n1125 71.676
R1452 B.n1131 B.n1130 71.676
R1453 B.n1134 B.n1133 71.676
R1454 B.n596 B.n349 71.676
R1455 B.n594 B.n351 71.676
R1456 B.n590 B.n589 71.676
R1457 B.n583 B.n353 71.676
R1458 B.n582 B.n581 71.676
R1459 B.n575 B.n355 71.676
R1460 B.n574 B.n573 71.676
R1461 B.n567 B.n357 71.676
R1462 B.n566 B.n565 71.676
R1463 B.n559 B.n359 71.676
R1464 B.n558 B.n557 71.676
R1465 B.n551 B.n361 71.676
R1466 B.n550 B.n549 71.676
R1467 B.n543 B.n363 71.676
R1468 B.n542 B.n541 71.676
R1469 B.n535 B.n365 71.676
R1470 B.n534 B.n533 71.676
R1471 B.n527 B.n367 71.676
R1472 B.n526 B.n525 71.676
R1473 B.n519 B.n369 71.676
R1474 B.n518 B.n517 71.676
R1475 B.n511 B.n371 71.676
R1476 B.n510 B.n375 71.676
R1477 B.n506 B.n505 71.676
R1478 B.n499 B.n377 71.676
R1479 B.n498 B.n497 71.676
R1480 B.n490 B.n379 71.676
R1481 B.n489 B.n488 71.676
R1482 B.n482 B.n383 71.676
R1483 B.n481 B.n480 71.676
R1484 B.n474 B.n385 71.676
R1485 B.n473 B.n472 71.676
R1486 B.n466 B.n387 71.676
R1487 B.n465 B.n464 71.676
R1488 B.n458 B.n389 71.676
R1489 B.n457 B.n456 71.676
R1490 B.n450 B.n391 71.676
R1491 B.n449 B.n448 71.676
R1492 B.n442 B.n393 71.676
R1493 B.n441 B.n440 71.676
R1494 B.n434 B.n395 71.676
R1495 B.n433 B.n432 71.676
R1496 B.n426 B.n397 71.676
R1497 B.n425 B.n424 71.676
R1498 B.n418 B.n399 71.676
R1499 B.n417 B.n416 71.676
R1500 B.n410 B.n401 71.676
R1501 B.n409 B.n408 71.676
R1502 B.n404 B.n403 71.676
R1503 B.n597 B.n596 71.676
R1504 B.n591 B.n351 71.676
R1505 B.n589 B.n588 71.676
R1506 B.n584 B.n583 71.676
R1507 B.n581 B.n580 71.676
R1508 B.n576 B.n575 71.676
R1509 B.n573 B.n572 71.676
R1510 B.n568 B.n567 71.676
R1511 B.n565 B.n564 71.676
R1512 B.n560 B.n559 71.676
R1513 B.n557 B.n556 71.676
R1514 B.n552 B.n551 71.676
R1515 B.n549 B.n548 71.676
R1516 B.n544 B.n543 71.676
R1517 B.n541 B.n540 71.676
R1518 B.n536 B.n535 71.676
R1519 B.n533 B.n532 71.676
R1520 B.n528 B.n527 71.676
R1521 B.n525 B.n524 71.676
R1522 B.n520 B.n519 71.676
R1523 B.n517 B.n516 71.676
R1524 B.n512 B.n511 71.676
R1525 B.n507 B.n375 71.676
R1526 B.n505 B.n504 71.676
R1527 B.n500 B.n499 71.676
R1528 B.n497 B.n496 71.676
R1529 B.n491 B.n490 71.676
R1530 B.n488 B.n487 71.676
R1531 B.n483 B.n482 71.676
R1532 B.n480 B.n479 71.676
R1533 B.n475 B.n474 71.676
R1534 B.n472 B.n471 71.676
R1535 B.n467 B.n466 71.676
R1536 B.n464 B.n463 71.676
R1537 B.n459 B.n458 71.676
R1538 B.n456 B.n455 71.676
R1539 B.n451 B.n450 71.676
R1540 B.n448 B.n447 71.676
R1541 B.n443 B.n442 71.676
R1542 B.n440 B.n439 71.676
R1543 B.n435 B.n434 71.676
R1544 B.n432 B.n431 71.676
R1545 B.n427 B.n426 71.676
R1546 B.n424 B.n423 71.676
R1547 B.n419 B.n418 71.676
R1548 B.n416 B.n415 71.676
R1549 B.n411 B.n410 71.676
R1550 B.n408 B.n407 71.676
R1551 B.n403 B.n347 71.676
R1552 B.n1296 B.n1295 71.676
R1553 B.n1296 B.n2 71.676
R1554 B.n173 B.t16 69.4087
R1555 B.n381 B.t19 69.4087
R1556 B.n167 B.t13 69.392
R1557 B.n373 B.t22 69.392
R1558 B.n602 B.n348 67.9797
R1559 B.n1139 B.n142 67.9797
R1560 B.n1047 B.n167 59.5399
R1561 B.n174 B.n173 59.5399
R1562 B.n493 B.n381 59.5399
R1563 B.n374 B.n373 59.5399
R1564 B.n602 B.n344 40.9083
R1565 B.n608 B.n344 40.9083
R1566 B.n608 B.n340 40.9083
R1567 B.n614 B.n340 40.9083
R1568 B.n614 B.n336 40.9083
R1569 B.n620 B.n336 40.9083
R1570 B.n620 B.n331 40.9083
R1571 B.n626 B.n331 40.9083
R1572 B.n626 B.n332 40.9083
R1573 B.n632 B.n324 40.9083
R1574 B.n638 B.n324 40.9083
R1575 B.n638 B.n320 40.9083
R1576 B.n644 B.n320 40.9083
R1577 B.n644 B.n316 40.9083
R1578 B.n650 B.n316 40.9083
R1579 B.n650 B.n312 40.9083
R1580 B.n656 B.n312 40.9083
R1581 B.n656 B.n308 40.9083
R1582 B.n662 B.n308 40.9083
R1583 B.n662 B.n304 40.9083
R1584 B.n668 B.n304 40.9083
R1585 B.n668 B.n300 40.9083
R1586 B.n674 B.n300 40.9083
R1587 B.n680 B.n296 40.9083
R1588 B.n680 B.n292 40.9083
R1589 B.n686 B.n292 40.9083
R1590 B.n686 B.n288 40.9083
R1591 B.n692 B.n288 40.9083
R1592 B.n692 B.n284 40.9083
R1593 B.n698 B.n284 40.9083
R1594 B.n698 B.n280 40.9083
R1595 B.n705 B.n280 40.9083
R1596 B.n705 B.n704 40.9083
R1597 B.n711 B.n273 40.9083
R1598 B.n717 B.n273 40.9083
R1599 B.n717 B.n269 40.9083
R1600 B.n723 B.n269 40.9083
R1601 B.n723 B.n265 40.9083
R1602 B.n729 B.n265 40.9083
R1603 B.n729 B.n261 40.9083
R1604 B.n735 B.n261 40.9083
R1605 B.n735 B.n257 40.9083
R1606 B.n742 B.n257 40.9083
R1607 B.n742 B.n741 40.9083
R1608 B.n748 B.n250 40.9083
R1609 B.n754 B.n250 40.9083
R1610 B.n754 B.n246 40.9083
R1611 B.n760 B.n246 40.9083
R1612 B.n760 B.n242 40.9083
R1613 B.n766 B.n242 40.9083
R1614 B.n766 B.n238 40.9083
R1615 B.n772 B.n238 40.9083
R1616 B.n772 B.n234 40.9083
R1617 B.n779 B.n234 40.9083
R1618 B.n779 B.n778 40.9083
R1619 B.n785 B.n227 40.9083
R1620 B.n791 B.n227 40.9083
R1621 B.n791 B.n223 40.9083
R1622 B.n797 B.n223 40.9083
R1623 B.n797 B.n219 40.9083
R1624 B.n803 B.n219 40.9083
R1625 B.n803 B.n215 40.9083
R1626 B.n809 B.n215 40.9083
R1627 B.n809 B.n211 40.9083
R1628 B.n816 B.n211 40.9083
R1629 B.n816 B.n815 40.9083
R1630 B.n822 B.n204 40.9083
R1631 B.n829 B.n204 40.9083
R1632 B.n829 B.n200 40.9083
R1633 B.n835 B.n200 40.9083
R1634 B.n835 B.n4 40.9083
R1635 B.n1294 B.n4 40.9083
R1636 B.n1294 B.n1293 40.9083
R1637 B.n1293 B.n1292 40.9083
R1638 B.n1292 B.n8 40.9083
R1639 B.n12 B.n8 40.9083
R1640 B.n1285 B.n12 40.9083
R1641 B.n1285 B.n1284 40.9083
R1642 B.n1284 B.n1283 40.9083
R1643 B.n1277 B.n19 40.9083
R1644 B.n1277 B.n1276 40.9083
R1645 B.n1276 B.n1275 40.9083
R1646 B.n1275 B.n23 40.9083
R1647 B.n1269 B.n23 40.9083
R1648 B.n1269 B.n1268 40.9083
R1649 B.n1268 B.n1267 40.9083
R1650 B.n1267 B.n30 40.9083
R1651 B.n1261 B.n30 40.9083
R1652 B.n1261 B.n1260 40.9083
R1653 B.n1260 B.n1259 40.9083
R1654 B.n1253 B.n40 40.9083
R1655 B.n1253 B.n1252 40.9083
R1656 B.n1252 B.n1251 40.9083
R1657 B.n1251 B.n44 40.9083
R1658 B.n1245 B.n44 40.9083
R1659 B.n1245 B.n1244 40.9083
R1660 B.n1244 B.n1243 40.9083
R1661 B.n1243 B.n51 40.9083
R1662 B.n1237 B.n51 40.9083
R1663 B.n1237 B.n1236 40.9083
R1664 B.n1236 B.n1235 40.9083
R1665 B.n1229 B.n61 40.9083
R1666 B.n1229 B.n1228 40.9083
R1667 B.n1228 B.n1227 40.9083
R1668 B.n1227 B.n65 40.9083
R1669 B.n1221 B.n65 40.9083
R1670 B.n1221 B.n1220 40.9083
R1671 B.n1220 B.n1219 40.9083
R1672 B.n1219 B.n72 40.9083
R1673 B.n1213 B.n72 40.9083
R1674 B.n1213 B.n1212 40.9083
R1675 B.n1212 B.n1211 40.9083
R1676 B.n1205 B.n82 40.9083
R1677 B.n1205 B.n1204 40.9083
R1678 B.n1204 B.n1203 40.9083
R1679 B.n1203 B.n86 40.9083
R1680 B.n1197 B.n86 40.9083
R1681 B.n1197 B.n1196 40.9083
R1682 B.n1196 B.n1195 40.9083
R1683 B.n1195 B.n93 40.9083
R1684 B.n1189 B.n93 40.9083
R1685 B.n1189 B.n1188 40.9083
R1686 B.n1187 B.n100 40.9083
R1687 B.n1181 B.n100 40.9083
R1688 B.n1181 B.n1180 40.9083
R1689 B.n1180 B.n1179 40.9083
R1690 B.n1179 B.n107 40.9083
R1691 B.n1173 B.n107 40.9083
R1692 B.n1173 B.n1172 40.9083
R1693 B.n1172 B.n1171 40.9083
R1694 B.n1171 B.n114 40.9083
R1695 B.n1165 B.n114 40.9083
R1696 B.n1165 B.n1164 40.9083
R1697 B.n1164 B.n1163 40.9083
R1698 B.n1163 B.n121 40.9083
R1699 B.n1157 B.n121 40.9083
R1700 B.n1156 B.n1155 40.9083
R1701 B.n1155 B.n128 40.9083
R1702 B.n1149 B.n128 40.9083
R1703 B.n1149 B.n1148 40.9083
R1704 B.n1148 B.n1147 40.9083
R1705 B.n1147 B.n135 40.9083
R1706 B.n1141 B.n135 40.9083
R1707 B.n1141 B.n1140 40.9083
R1708 B.n1140 B.n1139 40.9083
R1709 B.n822 B.t4 39.1036
R1710 B.n1283 B.t3 39.1036
R1711 B.n704 B.t2 37.9004
R1712 B.n82 B.t9 37.9004
R1713 B.t1 B.n296 31.8846
R1714 B.n1188 B.t6 31.8846
R1715 B.n600 B.n599 29.5029
R1716 B.n604 B.n346 29.5029
R1717 B.n939 B.n938 29.5029
R1718 B.n1137 B.n1136 29.5029
R1719 B.n632 B.t18 28.275
R1720 B.n1157 B.t11 28.275
R1721 B.n785 B.t8 27.0719
R1722 B.n1259 B.t7 27.0719
R1723 B.n741 B.t5 25.8687
R1724 B.n61 B.t0 25.8687
R1725 B B.n1297 18.0485
R1726 B.n748 B.t5 15.0401
R1727 B.n1235 B.t0 15.0401
R1728 B.n778 B.t8 13.837
R1729 B.n40 B.t7 13.837
R1730 B.n332 B.t18 12.6338
R1731 B.t11 B.n1156 12.6338
R1732 B.n600 B.n342 10.6151
R1733 B.n610 B.n342 10.6151
R1734 B.n611 B.n610 10.6151
R1735 B.n612 B.n611 10.6151
R1736 B.n612 B.n334 10.6151
R1737 B.n622 B.n334 10.6151
R1738 B.n623 B.n622 10.6151
R1739 B.n624 B.n623 10.6151
R1740 B.n624 B.n326 10.6151
R1741 B.n634 B.n326 10.6151
R1742 B.n635 B.n634 10.6151
R1743 B.n636 B.n635 10.6151
R1744 B.n636 B.n318 10.6151
R1745 B.n646 B.n318 10.6151
R1746 B.n647 B.n646 10.6151
R1747 B.n648 B.n647 10.6151
R1748 B.n648 B.n310 10.6151
R1749 B.n658 B.n310 10.6151
R1750 B.n659 B.n658 10.6151
R1751 B.n660 B.n659 10.6151
R1752 B.n660 B.n302 10.6151
R1753 B.n670 B.n302 10.6151
R1754 B.n671 B.n670 10.6151
R1755 B.n672 B.n671 10.6151
R1756 B.n672 B.n294 10.6151
R1757 B.n682 B.n294 10.6151
R1758 B.n683 B.n682 10.6151
R1759 B.n684 B.n683 10.6151
R1760 B.n684 B.n286 10.6151
R1761 B.n694 B.n286 10.6151
R1762 B.n695 B.n694 10.6151
R1763 B.n696 B.n695 10.6151
R1764 B.n696 B.n278 10.6151
R1765 B.n707 B.n278 10.6151
R1766 B.n708 B.n707 10.6151
R1767 B.n709 B.n708 10.6151
R1768 B.n709 B.n271 10.6151
R1769 B.n719 B.n271 10.6151
R1770 B.n720 B.n719 10.6151
R1771 B.n721 B.n720 10.6151
R1772 B.n721 B.n263 10.6151
R1773 B.n731 B.n263 10.6151
R1774 B.n732 B.n731 10.6151
R1775 B.n733 B.n732 10.6151
R1776 B.n733 B.n255 10.6151
R1777 B.n744 B.n255 10.6151
R1778 B.n745 B.n744 10.6151
R1779 B.n746 B.n745 10.6151
R1780 B.n746 B.n248 10.6151
R1781 B.n756 B.n248 10.6151
R1782 B.n757 B.n756 10.6151
R1783 B.n758 B.n757 10.6151
R1784 B.n758 B.n240 10.6151
R1785 B.n768 B.n240 10.6151
R1786 B.n769 B.n768 10.6151
R1787 B.n770 B.n769 10.6151
R1788 B.n770 B.n232 10.6151
R1789 B.n781 B.n232 10.6151
R1790 B.n782 B.n781 10.6151
R1791 B.n783 B.n782 10.6151
R1792 B.n783 B.n225 10.6151
R1793 B.n793 B.n225 10.6151
R1794 B.n794 B.n793 10.6151
R1795 B.n795 B.n794 10.6151
R1796 B.n795 B.n217 10.6151
R1797 B.n805 B.n217 10.6151
R1798 B.n806 B.n805 10.6151
R1799 B.n807 B.n806 10.6151
R1800 B.n807 B.n209 10.6151
R1801 B.n818 B.n209 10.6151
R1802 B.n819 B.n818 10.6151
R1803 B.n820 B.n819 10.6151
R1804 B.n820 B.n202 10.6151
R1805 B.n831 B.n202 10.6151
R1806 B.n832 B.n831 10.6151
R1807 B.n833 B.n832 10.6151
R1808 B.n833 B.n0 10.6151
R1809 B.n599 B.n598 10.6151
R1810 B.n598 B.n350 10.6151
R1811 B.n593 B.n350 10.6151
R1812 B.n593 B.n592 10.6151
R1813 B.n592 B.n352 10.6151
R1814 B.n587 B.n352 10.6151
R1815 B.n587 B.n586 10.6151
R1816 B.n586 B.n585 10.6151
R1817 B.n585 B.n354 10.6151
R1818 B.n579 B.n354 10.6151
R1819 B.n579 B.n578 10.6151
R1820 B.n578 B.n577 10.6151
R1821 B.n577 B.n356 10.6151
R1822 B.n571 B.n356 10.6151
R1823 B.n571 B.n570 10.6151
R1824 B.n570 B.n569 10.6151
R1825 B.n569 B.n358 10.6151
R1826 B.n563 B.n358 10.6151
R1827 B.n563 B.n562 10.6151
R1828 B.n562 B.n561 10.6151
R1829 B.n561 B.n360 10.6151
R1830 B.n555 B.n360 10.6151
R1831 B.n555 B.n554 10.6151
R1832 B.n554 B.n553 10.6151
R1833 B.n553 B.n362 10.6151
R1834 B.n547 B.n362 10.6151
R1835 B.n547 B.n546 10.6151
R1836 B.n546 B.n545 10.6151
R1837 B.n545 B.n364 10.6151
R1838 B.n539 B.n364 10.6151
R1839 B.n539 B.n538 10.6151
R1840 B.n538 B.n537 10.6151
R1841 B.n537 B.n366 10.6151
R1842 B.n531 B.n366 10.6151
R1843 B.n531 B.n530 10.6151
R1844 B.n530 B.n529 10.6151
R1845 B.n529 B.n368 10.6151
R1846 B.n523 B.n368 10.6151
R1847 B.n523 B.n522 10.6151
R1848 B.n522 B.n521 10.6151
R1849 B.n521 B.n370 10.6151
R1850 B.n515 B.n370 10.6151
R1851 B.n515 B.n514 10.6151
R1852 B.n514 B.n513 10.6151
R1853 B.n509 B.n508 10.6151
R1854 B.n508 B.n376 10.6151
R1855 B.n503 B.n376 10.6151
R1856 B.n503 B.n502 10.6151
R1857 B.n502 B.n501 10.6151
R1858 B.n501 B.n378 10.6151
R1859 B.n495 B.n378 10.6151
R1860 B.n495 B.n494 10.6151
R1861 B.n492 B.n382 10.6151
R1862 B.n486 B.n382 10.6151
R1863 B.n486 B.n485 10.6151
R1864 B.n485 B.n484 10.6151
R1865 B.n484 B.n384 10.6151
R1866 B.n478 B.n384 10.6151
R1867 B.n478 B.n477 10.6151
R1868 B.n477 B.n476 10.6151
R1869 B.n476 B.n386 10.6151
R1870 B.n470 B.n386 10.6151
R1871 B.n470 B.n469 10.6151
R1872 B.n469 B.n468 10.6151
R1873 B.n468 B.n388 10.6151
R1874 B.n462 B.n388 10.6151
R1875 B.n462 B.n461 10.6151
R1876 B.n461 B.n460 10.6151
R1877 B.n460 B.n390 10.6151
R1878 B.n454 B.n390 10.6151
R1879 B.n454 B.n453 10.6151
R1880 B.n453 B.n452 10.6151
R1881 B.n452 B.n392 10.6151
R1882 B.n446 B.n392 10.6151
R1883 B.n446 B.n445 10.6151
R1884 B.n445 B.n444 10.6151
R1885 B.n444 B.n394 10.6151
R1886 B.n438 B.n394 10.6151
R1887 B.n438 B.n437 10.6151
R1888 B.n437 B.n436 10.6151
R1889 B.n436 B.n396 10.6151
R1890 B.n430 B.n396 10.6151
R1891 B.n430 B.n429 10.6151
R1892 B.n429 B.n428 10.6151
R1893 B.n428 B.n398 10.6151
R1894 B.n422 B.n398 10.6151
R1895 B.n422 B.n421 10.6151
R1896 B.n421 B.n420 10.6151
R1897 B.n420 B.n400 10.6151
R1898 B.n414 B.n400 10.6151
R1899 B.n414 B.n413 10.6151
R1900 B.n413 B.n412 10.6151
R1901 B.n412 B.n402 10.6151
R1902 B.n406 B.n402 10.6151
R1903 B.n406 B.n405 10.6151
R1904 B.n405 B.n346 10.6151
R1905 B.n605 B.n604 10.6151
R1906 B.n606 B.n605 10.6151
R1907 B.n606 B.n338 10.6151
R1908 B.n616 B.n338 10.6151
R1909 B.n617 B.n616 10.6151
R1910 B.n618 B.n617 10.6151
R1911 B.n618 B.n329 10.6151
R1912 B.n628 B.n329 10.6151
R1913 B.n629 B.n628 10.6151
R1914 B.n630 B.n629 10.6151
R1915 B.n630 B.n322 10.6151
R1916 B.n640 B.n322 10.6151
R1917 B.n641 B.n640 10.6151
R1918 B.n642 B.n641 10.6151
R1919 B.n642 B.n314 10.6151
R1920 B.n652 B.n314 10.6151
R1921 B.n653 B.n652 10.6151
R1922 B.n654 B.n653 10.6151
R1923 B.n654 B.n306 10.6151
R1924 B.n664 B.n306 10.6151
R1925 B.n665 B.n664 10.6151
R1926 B.n666 B.n665 10.6151
R1927 B.n666 B.n298 10.6151
R1928 B.n676 B.n298 10.6151
R1929 B.n677 B.n676 10.6151
R1930 B.n678 B.n677 10.6151
R1931 B.n678 B.n290 10.6151
R1932 B.n688 B.n290 10.6151
R1933 B.n689 B.n688 10.6151
R1934 B.n690 B.n689 10.6151
R1935 B.n690 B.n282 10.6151
R1936 B.n700 B.n282 10.6151
R1937 B.n701 B.n700 10.6151
R1938 B.n702 B.n701 10.6151
R1939 B.n702 B.n275 10.6151
R1940 B.n713 B.n275 10.6151
R1941 B.n714 B.n713 10.6151
R1942 B.n715 B.n714 10.6151
R1943 B.n715 B.n267 10.6151
R1944 B.n725 B.n267 10.6151
R1945 B.n726 B.n725 10.6151
R1946 B.n727 B.n726 10.6151
R1947 B.n727 B.n259 10.6151
R1948 B.n737 B.n259 10.6151
R1949 B.n738 B.n737 10.6151
R1950 B.n739 B.n738 10.6151
R1951 B.n739 B.n252 10.6151
R1952 B.n750 B.n252 10.6151
R1953 B.n751 B.n750 10.6151
R1954 B.n752 B.n751 10.6151
R1955 B.n752 B.n244 10.6151
R1956 B.n762 B.n244 10.6151
R1957 B.n763 B.n762 10.6151
R1958 B.n764 B.n763 10.6151
R1959 B.n764 B.n236 10.6151
R1960 B.n774 B.n236 10.6151
R1961 B.n775 B.n774 10.6151
R1962 B.n776 B.n775 10.6151
R1963 B.n776 B.n229 10.6151
R1964 B.n787 B.n229 10.6151
R1965 B.n788 B.n787 10.6151
R1966 B.n789 B.n788 10.6151
R1967 B.n789 B.n221 10.6151
R1968 B.n799 B.n221 10.6151
R1969 B.n800 B.n799 10.6151
R1970 B.n801 B.n800 10.6151
R1971 B.n801 B.n213 10.6151
R1972 B.n811 B.n213 10.6151
R1973 B.n812 B.n811 10.6151
R1974 B.n813 B.n812 10.6151
R1975 B.n813 B.n206 10.6151
R1976 B.n824 B.n206 10.6151
R1977 B.n825 B.n824 10.6151
R1978 B.n827 B.n825 10.6151
R1979 B.n827 B.n826 10.6151
R1980 B.n826 B.n198 10.6151
R1981 B.n838 B.n198 10.6151
R1982 B.n839 B.n838 10.6151
R1983 B.n840 B.n839 10.6151
R1984 B.n841 B.n840 10.6151
R1985 B.n842 B.n841 10.6151
R1986 B.n845 B.n842 10.6151
R1987 B.n846 B.n845 10.6151
R1988 B.n847 B.n846 10.6151
R1989 B.n848 B.n847 10.6151
R1990 B.n850 B.n848 10.6151
R1991 B.n851 B.n850 10.6151
R1992 B.n852 B.n851 10.6151
R1993 B.n853 B.n852 10.6151
R1994 B.n855 B.n853 10.6151
R1995 B.n856 B.n855 10.6151
R1996 B.n857 B.n856 10.6151
R1997 B.n858 B.n857 10.6151
R1998 B.n860 B.n858 10.6151
R1999 B.n861 B.n860 10.6151
R2000 B.n862 B.n861 10.6151
R2001 B.n863 B.n862 10.6151
R2002 B.n865 B.n863 10.6151
R2003 B.n866 B.n865 10.6151
R2004 B.n867 B.n866 10.6151
R2005 B.n868 B.n867 10.6151
R2006 B.n870 B.n868 10.6151
R2007 B.n871 B.n870 10.6151
R2008 B.n872 B.n871 10.6151
R2009 B.n873 B.n872 10.6151
R2010 B.n875 B.n873 10.6151
R2011 B.n876 B.n875 10.6151
R2012 B.n877 B.n876 10.6151
R2013 B.n878 B.n877 10.6151
R2014 B.n880 B.n878 10.6151
R2015 B.n881 B.n880 10.6151
R2016 B.n882 B.n881 10.6151
R2017 B.n883 B.n882 10.6151
R2018 B.n885 B.n883 10.6151
R2019 B.n886 B.n885 10.6151
R2020 B.n887 B.n886 10.6151
R2021 B.n888 B.n887 10.6151
R2022 B.n890 B.n888 10.6151
R2023 B.n891 B.n890 10.6151
R2024 B.n892 B.n891 10.6151
R2025 B.n893 B.n892 10.6151
R2026 B.n895 B.n893 10.6151
R2027 B.n896 B.n895 10.6151
R2028 B.n897 B.n896 10.6151
R2029 B.n898 B.n897 10.6151
R2030 B.n900 B.n898 10.6151
R2031 B.n901 B.n900 10.6151
R2032 B.n902 B.n901 10.6151
R2033 B.n903 B.n902 10.6151
R2034 B.n905 B.n903 10.6151
R2035 B.n906 B.n905 10.6151
R2036 B.n907 B.n906 10.6151
R2037 B.n908 B.n907 10.6151
R2038 B.n910 B.n908 10.6151
R2039 B.n911 B.n910 10.6151
R2040 B.n912 B.n911 10.6151
R2041 B.n913 B.n912 10.6151
R2042 B.n915 B.n913 10.6151
R2043 B.n916 B.n915 10.6151
R2044 B.n917 B.n916 10.6151
R2045 B.n918 B.n917 10.6151
R2046 B.n920 B.n918 10.6151
R2047 B.n921 B.n920 10.6151
R2048 B.n922 B.n921 10.6151
R2049 B.n923 B.n922 10.6151
R2050 B.n925 B.n923 10.6151
R2051 B.n926 B.n925 10.6151
R2052 B.n927 B.n926 10.6151
R2053 B.n928 B.n927 10.6151
R2054 B.n930 B.n928 10.6151
R2055 B.n931 B.n930 10.6151
R2056 B.n932 B.n931 10.6151
R2057 B.n933 B.n932 10.6151
R2058 B.n935 B.n933 10.6151
R2059 B.n936 B.n935 10.6151
R2060 B.n937 B.n936 10.6151
R2061 B.n938 B.n937 10.6151
R2062 B.n1289 B.n1 10.6151
R2063 B.n1289 B.n1288 10.6151
R2064 B.n1288 B.n1287 10.6151
R2065 B.n1287 B.n10 10.6151
R2066 B.n1281 B.n10 10.6151
R2067 B.n1281 B.n1280 10.6151
R2068 B.n1280 B.n1279 10.6151
R2069 B.n1279 B.n17 10.6151
R2070 B.n1273 B.n17 10.6151
R2071 B.n1273 B.n1272 10.6151
R2072 B.n1272 B.n1271 10.6151
R2073 B.n1271 B.n25 10.6151
R2074 B.n1265 B.n25 10.6151
R2075 B.n1265 B.n1264 10.6151
R2076 B.n1264 B.n1263 10.6151
R2077 B.n1263 B.n32 10.6151
R2078 B.n1257 B.n32 10.6151
R2079 B.n1257 B.n1256 10.6151
R2080 B.n1256 B.n1255 10.6151
R2081 B.n1255 B.n38 10.6151
R2082 B.n1249 B.n38 10.6151
R2083 B.n1249 B.n1248 10.6151
R2084 B.n1248 B.n1247 10.6151
R2085 B.n1247 B.n46 10.6151
R2086 B.n1241 B.n46 10.6151
R2087 B.n1241 B.n1240 10.6151
R2088 B.n1240 B.n1239 10.6151
R2089 B.n1239 B.n53 10.6151
R2090 B.n1233 B.n53 10.6151
R2091 B.n1233 B.n1232 10.6151
R2092 B.n1232 B.n1231 10.6151
R2093 B.n1231 B.n59 10.6151
R2094 B.n1225 B.n59 10.6151
R2095 B.n1225 B.n1224 10.6151
R2096 B.n1224 B.n1223 10.6151
R2097 B.n1223 B.n67 10.6151
R2098 B.n1217 B.n67 10.6151
R2099 B.n1217 B.n1216 10.6151
R2100 B.n1216 B.n1215 10.6151
R2101 B.n1215 B.n74 10.6151
R2102 B.n1209 B.n74 10.6151
R2103 B.n1209 B.n1208 10.6151
R2104 B.n1208 B.n1207 10.6151
R2105 B.n1207 B.n80 10.6151
R2106 B.n1201 B.n80 10.6151
R2107 B.n1201 B.n1200 10.6151
R2108 B.n1200 B.n1199 10.6151
R2109 B.n1199 B.n88 10.6151
R2110 B.n1193 B.n88 10.6151
R2111 B.n1193 B.n1192 10.6151
R2112 B.n1192 B.n1191 10.6151
R2113 B.n1191 B.n95 10.6151
R2114 B.n1185 B.n95 10.6151
R2115 B.n1185 B.n1184 10.6151
R2116 B.n1184 B.n1183 10.6151
R2117 B.n1183 B.n102 10.6151
R2118 B.n1177 B.n102 10.6151
R2119 B.n1177 B.n1176 10.6151
R2120 B.n1176 B.n1175 10.6151
R2121 B.n1175 B.n109 10.6151
R2122 B.n1169 B.n109 10.6151
R2123 B.n1169 B.n1168 10.6151
R2124 B.n1168 B.n1167 10.6151
R2125 B.n1167 B.n116 10.6151
R2126 B.n1161 B.n116 10.6151
R2127 B.n1161 B.n1160 10.6151
R2128 B.n1160 B.n1159 10.6151
R2129 B.n1159 B.n123 10.6151
R2130 B.n1153 B.n123 10.6151
R2131 B.n1153 B.n1152 10.6151
R2132 B.n1152 B.n1151 10.6151
R2133 B.n1151 B.n130 10.6151
R2134 B.n1145 B.n130 10.6151
R2135 B.n1145 B.n1144 10.6151
R2136 B.n1144 B.n1143 10.6151
R2137 B.n1143 B.n137 10.6151
R2138 B.n1137 B.n137 10.6151
R2139 B.n1136 B.n1135 10.6151
R2140 B.n1135 B.n144 10.6151
R2141 B.n1129 B.n144 10.6151
R2142 B.n1129 B.n1128 10.6151
R2143 B.n1128 B.n1127 10.6151
R2144 B.n1127 B.n146 10.6151
R2145 B.n1121 B.n146 10.6151
R2146 B.n1121 B.n1120 10.6151
R2147 B.n1120 B.n1119 10.6151
R2148 B.n1119 B.n148 10.6151
R2149 B.n1113 B.n148 10.6151
R2150 B.n1113 B.n1112 10.6151
R2151 B.n1112 B.n1111 10.6151
R2152 B.n1111 B.n150 10.6151
R2153 B.n1105 B.n150 10.6151
R2154 B.n1105 B.n1104 10.6151
R2155 B.n1104 B.n1103 10.6151
R2156 B.n1103 B.n152 10.6151
R2157 B.n1097 B.n152 10.6151
R2158 B.n1097 B.n1096 10.6151
R2159 B.n1096 B.n1095 10.6151
R2160 B.n1095 B.n154 10.6151
R2161 B.n1089 B.n154 10.6151
R2162 B.n1089 B.n1088 10.6151
R2163 B.n1088 B.n1087 10.6151
R2164 B.n1087 B.n156 10.6151
R2165 B.n1081 B.n156 10.6151
R2166 B.n1081 B.n1080 10.6151
R2167 B.n1080 B.n1079 10.6151
R2168 B.n1079 B.n158 10.6151
R2169 B.n1073 B.n158 10.6151
R2170 B.n1073 B.n1072 10.6151
R2171 B.n1072 B.n1071 10.6151
R2172 B.n1071 B.n160 10.6151
R2173 B.n1065 B.n160 10.6151
R2174 B.n1065 B.n1064 10.6151
R2175 B.n1064 B.n1063 10.6151
R2176 B.n1063 B.n162 10.6151
R2177 B.n1057 B.n162 10.6151
R2178 B.n1057 B.n1056 10.6151
R2179 B.n1056 B.n1055 10.6151
R2180 B.n1055 B.n164 10.6151
R2181 B.n1049 B.n164 10.6151
R2182 B.n1049 B.n1048 10.6151
R2183 B.n1046 B.n168 10.6151
R2184 B.n1040 B.n168 10.6151
R2185 B.n1040 B.n1039 10.6151
R2186 B.n1039 B.n1038 10.6151
R2187 B.n1038 B.n170 10.6151
R2188 B.n1032 B.n170 10.6151
R2189 B.n1032 B.n1031 10.6151
R2190 B.n1031 B.n1030 10.6151
R2191 B.n1026 B.n1025 10.6151
R2192 B.n1025 B.n176 10.6151
R2193 B.n1020 B.n176 10.6151
R2194 B.n1020 B.n1019 10.6151
R2195 B.n1019 B.n1018 10.6151
R2196 B.n1018 B.n178 10.6151
R2197 B.n1012 B.n178 10.6151
R2198 B.n1012 B.n1011 10.6151
R2199 B.n1011 B.n1010 10.6151
R2200 B.n1010 B.n180 10.6151
R2201 B.n1004 B.n180 10.6151
R2202 B.n1004 B.n1003 10.6151
R2203 B.n1003 B.n1002 10.6151
R2204 B.n1002 B.n182 10.6151
R2205 B.n996 B.n182 10.6151
R2206 B.n996 B.n995 10.6151
R2207 B.n995 B.n994 10.6151
R2208 B.n994 B.n184 10.6151
R2209 B.n988 B.n184 10.6151
R2210 B.n988 B.n987 10.6151
R2211 B.n987 B.n986 10.6151
R2212 B.n986 B.n186 10.6151
R2213 B.n980 B.n186 10.6151
R2214 B.n980 B.n979 10.6151
R2215 B.n979 B.n978 10.6151
R2216 B.n978 B.n188 10.6151
R2217 B.n972 B.n188 10.6151
R2218 B.n972 B.n971 10.6151
R2219 B.n971 B.n970 10.6151
R2220 B.n970 B.n190 10.6151
R2221 B.n964 B.n190 10.6151
R2222 B.n964 B.n963 10.6151
R2223 B.n963 B.n962 10.6151
R2224 B.n962 B.n192 10.6151
R2225 B.n956 B.n192 10.6151
R2226 B.n956 B.n955 10.6151
R2227 B.n955 B.n954 10.6151
R2228 B.n954 B.n194 10.6151
R2229 B.n948 B.n194 10.6151
R2230 B.n948 B.n947 10.6151
R2231 B.n947 B.n946 10.6151
R2232 B.n946 B.n196 10.6151
R2233 B.n940 B.n196 10.6151
R2234 B.n940 B.n939 10.6151
R2235 B.n674 B.t1 9.02429
R2236 B.t6 B.n1187 9.02429
R2237 B.n1297 B.n0 8.11757
R2238 B.n1297 B.n1 8.11757
R2239 B.n509 B.n374 6.5566
R2240 B.n494 B.n493 6.5566
R2241 B.n1047 B.n1046 6.5566
R2242 B.n1030 B.n174 6.5566
R2243 B.n513 B.n374 4.05904
R2244 B.n493 B.n492 4.05904
R2245 B.n1048 B.n1047 4.05904
R2246 B.n1026 B.n174 4.05904
R2247 B.n711 B.t2 3.00843
R2248 B.n1211 B.t9 3.00843
R2249 B.n815 B.t4 1.80526
R2250 B.n19 B.t3 1.80526
R2251 VP.n32 VP.n29 161.3
R2252 VP.n34 VP.n33 161.3
R2253 VP.n35 VP.n28 161.3
R2254 VP.n37 VP.n36 161.3
R2255 VP.n38 VP.n27 161.3
R2256 VP.n40 VP.n39 161.3
R2257 VP.n41 VP.n26 161.3
R2258 VP.n44 VP.n43 161.3
R2259 VP.n45 VP.n25 161.3
R2260 VP.n47 VP.n46 161.3
R2261 VP.n48 VP.n24 161.3
R2262 VP.n50 VP.n49 161.3
R2263 VP.n51 VP.n23 161.3
R2264 VP.n53 VP.n52 161.3
R2265 VP.n54 VP.n22 161.3
R2266 VP.n57 VP.n56 161.3
R2267 VP.n58 VP.n21 161.3
R2268 VP.n60 VP.n59 161.3
R2269 VP.n61 VP.n20 161.3
R2270 VP.n63 VP.n62 161.3
R2271 VP.n64 VP.n19 161.3
R2272 VP.n66 VP.n65 161.3
R2273 VP.n67 VP.n18 161.3
R2274 VP.n69 VP.n68 161.3
R2275 VP.n123 VP.n122 161.3
R2276 VP.n121 VP.n1 161.3
R2277 VP.n120 VP.n119 161.3
R2278 VP.n118 VP.n2 161.3
R2279 VP.n117 VP.n116 161.3
R2280 VP.n115 VP.n3 161.3
R2281 VP.n114 VP.n113 161.3
R2282 VP.n112 VP.n4 161.3
R2283 VP.n111 VP.n110 161.3
R2284 VP.n108 VP.n5 161.3
R2285 VP.n107 VP.n106 161.3
R2286 VP.n105 VP.n6 161.3
R2287 VP.n104 VP.n103 161.3
R2288 VP.n102 VP.n7 161.3
R2289 VP.n101 VP.n100 161.3
R2290 VP.n99 VP.n8 161.3
R2291 VP.n98 VP.n97 161.3
R2292 VP.n95 VP.n9 161.3
R2293 VP.n94 VP.n93 161.3
R2294 VP.n92 VP.n10 161.3
R2295 VP.n91 VP.n90 161.3
R2296 VP.n89 VP.n11 161.3
R2297 VP.n88 VP.n87 161.3
R2298 VP.n86 VP.n12 161.3
R2299 VP.n85 VP.n84 161.3
R2300 VP.n82 VP.n13 161.3
R2301 VP.n81 VP.n80 161.3
R2302 VP.n79 VP.n14 161.3
R2303 VP.n78 VP.n77 161.3
R2304 VP.n76 VP.n15 161.3
R2305 VP.n75 VP.n74 161.3
R2306 VP.n73 VP.n16 161.3
R2307 VP.n31 VP.t4 119.34
R2308 VP.n71 VP.t7 85.9021
R2309 VP.n83 VP.t1 85.9021
R2310 VP.n96 VP.t9 85.9021
R2311 VP.n109 VP.t5 85.9021
R2312 VP.n0 VP.t8 85.9021
R2313 VP.n17 VP.t2 85.9021
R2314 VP.n55 VP.t6 85.9021
R2315 VP.n42 VP.t0 85.9021
R2316 VP.n30 VP.t3 85.9021
R2317 VP.n72 VP.n71 79.7913
R2318 VP.n124 VP.n0 79.7913
R2319 VP.n70 VP.n17 79.7913
R2320 VP.n31 VP.n30 63.3588
R2321 VP.n72 VP.n70 59.719
R2322 VP.n77 VP.n14 56.5193
R2323 VP.n90 VP.n10 56.5193
R2324 VP.n103 VP.n6 56.5193
R2325 VP.n116 VP.n2 56.5193
R2326 VP.n62 VP.n19 56.5193
R2327 VP.n49 VP.n23 56.5193
R2328 VP.n36 VP.n27 56.5193
R2329 VP.n75 VP.n16 24.4675
R2330 VP.n76 VP.n75 24.4675
R2331 VP.n77 VP.n76 24.4675
R2332 VP.n81 VP.n14 24.4675
R2333 VP.n82 VP.n81 24.4675
R2334 VP.n84 VP.n82 24.4675
R2335 VP.n88 VP.n12 24.4675
R2336 VP.n89 VP.n88 24.4675
R2337 VP.n90 VP.n89 24.4675
R2338 VP.n94 VP.n10 24.4675
R2339 VP.n95 VP.n94 24.4675
R2340 VP.n97 VP.n95 24.4675
R2341 VP.n101 VP.n8 24.4675
R2342 VP.n102 VP.n101 24.4675
R2343 VP.n103 VP.n102 24.4675
R2344 VP.n107 VP.n6 24.4675
R2345 VP.n108 VP.n107 24.4675
R2346 VP.n110 VP.n108 24.4675
R2347 VP.n114 VP.n4 24.4675
R2348 VP.n115 VP.n114 24.4675
R2349 VP.n116 VP.n115 24.4675
R2350 VP.n120 VP.n2 24.4675
R2351 VP.n121 VP.n120 24.4675
R2352 VP.n122 VP.n121 24.4675
R2353 VP.n66 VP.n19 24.4675
R2354 VP.n67 VP.n66 24.4675
R2355 VP.n68 VP.n67 24.4675
R2356 VP.n53 VP.n23 24.4675
R2357 VP.n54 VP.n53 24.4675
R2358 VP.n56 VP.n54 24.4675
R2359 VP.n60 VP.n21 24.4675
R2360 VP.n61 VP.n60 24.4675
R2361 VP.n62 VP.n61 24.4675
R2362 VP.n40 VP.n27 24.4675
R2363 VP.n41 VP.n40 24.4675
R2364 VP.n43 VP.n41 24.4675
R2365 VP.n47 VP.n25 24.4675
R2366 VP.n48 VP.n47 24.4675
R2367 VP.n49 VP.n48 24.4675
R2368 VP.n34 VP.n29 24.4675
R2369 VP.n35 VP.n34 24.4675
R2370 VP.n36 VP.n35 24.4675
R2371 VP.n84 VP.n83 13.2127
R2372 VP.n109 VP.n4 13.2127
R2373 VP.n55 VP.n21 13.2127
R2374 VP.n97 VP.n96 12.234
R2375 VP.n96 VP.n8 12.234
R2376 VP.n43 VP.n42 12.234
R2377 VP.n42 VP.n25 12.234
R2378 VP.n83 VP.n12 11.2553
R2379 VP.n110 VP.n109 11.2553
R2380 VP.n56 VP.n55 11.2553
R2381 VP.n30 VP.n29 11.2553
R2382 VP.n71 VP.n16 10.2766
R2383 VP.n122 VP.n0 10.2766
R2384 VP.n68 VP.n17 10.2766
R2385 VP.n32 VP.n31 3.148
R2386 VP.n70 VP.n69 0.354971
R2387 VP.n73 VP.n72 0.354971
R2388 VP.n124 VP.n123 0.354971
R2389 VP VP.n124 0.26696
R2390 VP.n33 VP.n32 0.189894
R2391 VP.n33 VP.n28 0.189894
R2392 VP.n37 VP.n28 0.189894
R2393 VP.n38 VP.n37 0.189894
R2394 VP.n39 VP.n38 0.189894
R2395 VP.n39 VP.n26 0.189894
R2396 VP.n44 VP.n26 0.189894
R2397 VP.n45 VP.n44 0.189894
R2398 VP.n46 VP.n45 0.189894
R2399 VP.n46 VP.n24 0.189894
R2400 VP.n50 VP.n24 0.189894
R2401 VP.n51 VP.n50 0.189894
R2402 VP.n52 VP.n51 0.189894
R2403 VP.n52 VP.n22 0.189894
R2404 VP.n57 VP.n22 0.189894
R2405 VP.n58 VP.n57 0.189894
R2406 VP.n59 VP.n58 0.189894
R2407 VP.n59 VP.n20 0.189894
R2408 VP.n63 VP.n20 0.189894
R2409 VP.n64 VP.n63 0.189894
R2410 VP.n65 VP.n64 0.189894
R2411 VP.n65 VP.n18 0.189894
R2412 VP.n69 VP.n18 0.189894
R2413 VP.n74 VP.n73 0.189894
R2414 VP.n74 VP.n15 0.189894
R2415 VP.n78 VP.n15 0.189894
R2416 VP.n79 VP.n78 0.189894
R2417 VP.n80 VP.n79 0.189894
R2418 VP.n80 VP.n13 0.189894
R2419 VP.n85 VP.n13 0.189894
R2420 VP.n86 VP.n85 0.189894
R2421 VP.n87 VP.n86 0.189894
R2422 VP.n87 VP.n11 0.189894
R2423 VP.n91 VP.n11 0.189894
R2424 VP.n92 VP.n91 0.189894
R2425 VP.n93 VP.n92 0.189894
R2426 VP.n93 VP.n9 0.189894
R2427 VP.n98 VP.n9 0.189894
R2428 VP.n99 VP.n98 0.189894
R2429 VP.n100 VP.n99 0.189894
R2430 VP.n100 VP.n7 0.189894
R2431 VP.n104 VP.n7 0.189894
R2432 VP.n105 VP.n104 0.189894
R2433 VP.n106 VP.n105 0.189894
R2434 VP.n106 VP.n5 0.189894
R2435 VP.n111 VP.n5 0.189894
R2436 VP.n112 VP.n111 0.189894
R2437 VP.n113 VP.n112 0.189894
R2438 VP.n113 VP.n3 0.189894
R2439 VP.n117 VP.n3 0.189894
R2440 VP.n118 VP.n117 0.189894
R2441 VP.n119 VP.n118 0.189894
R2442 VP.n119 VP.n1 0.189894
R2443 VP.n123 VP.n1 0.189894
R2444 VTAIL.n11 VTAIL.t18 49.317
R2445 VTAIL.n17 VTAIL.t2 49.3159
R2446 VTAIL.n2 VTAIL.t5 49.3159
R2447 VTAIL.n16 VTAIL.t12 49.3159
R2448 VTAIL.n15 VTAIL.n14 47.7951
R2449 VTAIL.n13 VTAIL.n12 47.7951
R2450 VTAIL.n10 VTAIL.n9 47.7951
R2451 VTAIL.n8 VTAIL.n7 47.7951
R2452 VTAIL.n19 VTAIL.n18 47.794
R2453 VTAIL.n1 VTAIL.n0 47.794
R2454 VTAIL.n4 VTAIL.n3 47.794
R2455 VTAIL.n6 VTAIL.n5 47.794
R2456 VTAIL.n8 VTAIL.n6 30.4445
R2457 VTAIL.n17 VTAIL.n16 27.0134
R2458 VTAIL.n10 VTAIL.n8 3.43153
R2459 VTAIL.n11 VTAIL.n10 3.43153
R2460 VTAIL.n15 VTAIL.n13 3.43153
R2461 VTAIL.n16 VTAIL.n15 3.43153
R2462 VTAIL.n6 VTAIL.n4 3.43153
R2463 VTAIL.n4 VTAIL.n2 3.43153
R2464 VTAIL.n19 VTAIL.n17 3.43153
R2465 VTAIL VTAIL.n1 2.63197
R2466 VTAIL.n13 VTAIL.n11 2.18584
R2467 VTAIL.n2 VTAIL.n1 2.18584
R2468 VTAIL.n18 VTAIL.t17 1.52241
R2469 VTAIL.n18 VTAIL.t15 1.52241
R2470 VTAIL.n0 VTAIL.t16 1.52241
R2471 VTAIL.n0 VTAIL.t4 1.52241
R2472 VTAIL.n3 VTAIL.t8 1.52241
R2473 VTAIL.n3 VTAIL.t14 1.52241
R2474 VTAIL.n5 VTAIL.t9 1.52241
R2475 VTAIL.n5 VTAIL.t13 1.52241
R2476 VTAIL.n14 VTAIL.t7 1.52241
R2477 VTAIL.n14 VTAIL.t10 1.52241
R2478 VTAIL.n12 VTAIL.t6 1.52241
R2479 VTAIL.n12 VTAIL.t11 1.52241
R2480 VTAIL.n9 VTAIL.t1 1.52241
R2481 VTAIL.n9 VTAIL.t19 1.52241
R2482 VTAIL.n7 VTAIL.t3 1.52241
R2483 VTAIL.n7 VTAIL.t0 1.52241
R2484 VTAIL VTAIL.n19 0.800069
R2485 VDD1.n1 VDD1.t5 69.4268
R2486 VDD1.n3 VDD1.t2 69.4257
R2487 VDD1.n5 VDD1.n4 66.9907
R2488 VDD1.n1 VDD1.n0 64.4739
R2489 VDD1.n7 VDD1.n6 64.4728
R2490 VDD1.n3 VDD1.n2 64.4728
R2491 VDD1.n7 VDD1.n5 53.5268
R2492 VDD1 VDD1.n7 2.51559
R2493 VDD1.n6 VDD1.t3 1.52241
R2494 VDD1.n6 VDD1.t7 1.52241
R2495 VDD1.n0 VDD1.t6 1.52241
R2496 VDD1.n0 VDD1.t9 1.52241
R2497 VDD1.n4 VDD1.t4 1.52241
R2498 VDD1.n4 VDD1.t1 1.52241
R2499 VDD1.n2 VDD1.t8 1.52241
R2500 VDD1.n2 VDD1.t0 1.52241
R2501 VDD1 VDD1.n1 0.916448
R2502 VDD1.n5 VDD1.n3 0.802913
R2503 VN.n106 VN.n105 161.3
R2504 VN.n104 VN.n55 161.3
R2505 VN.n103 VN.n102 161.3
R2506 VN.n101 VN.n56 161.3
R2507 VN.n100 VN.n99 161.3
R2508 VN.n98 VN.n57 161.3
R2509 VN.n97 VN.n96 161.3
R2510 VN.n95 VN.n58 161.3
R2511 VN.n94 VN.n93 161.3
R2512 VN.n92 VN.n59 161.3
R2513 VN.n91 VN.n90 161.3
R2514 VN.n89 VN.n61 161.3
R2515 VN.n88 VN.n87 161.3
R2516 VN.n86 VN.n62 161.3
R2517 VN.n85 VN.n84 161.3
R2518 VN.n83 VN.n63 161.3
R2519 VN.n82 VN.n81 161.3
R2520 VN.n80 VN.n64 161.3
R2521 VN.n79 VN.n78 161.3
R2522 VN.n77 VN.n66 161.3
R2523 VN.n76 VN.n75 161.3
R2524 VN.n74 VN.n67 161.3
R2525 VN.n73 VN.n72 161.3
R2526 VN.n71 VN.n68 161.3
R2527 VN.n52 VN.n51 161.3
R2528 VN.n50 VN.n1 161.3
R2529 VN.n49 VN.n48 161.3
R2530 VN.n47 VN.n2 161.3
R2531 VN.n46 VN.n45 161.3
R2532 VN.n44 VN.n3 161.3
R2533 VN.n43 VN.n42 161.3
R2534 VN.n41 VN.n4 161.3
R2535 VN.n40 VN.n39 161.3
R2536 VN.n37 VN.n5 161.3
R2537 VN.n36 VN.n35 161.3
R2538 VN.n34 VN.n6 161.3
R2539 VN.n33 VN.n32 161.3
R2540 VN.n31 VN.n7 161.3
R2541 VN.n30 VN.n29 161.3
R2542 VN.n28 VN.n8 161.3
R2543 VN.n27 VN.n26 161.3
R2544 VN.n24 VN.n9 161.3
R2545 VN.n23 VN.n22 161.3
R2546 VN.n21 VN.n10 161.3
R2547 VN.n20 VN.n19 161.3
R2548 VN.n18 VN.n11 161.3
R2549 VN.n17 VN.n16 161.3
R2550 VN.n15 VN.n12 161.3
R2551 VN.n70 VN.t5 119.34
R2552 VN.n14 VN.t8 119.34
R2553 VN.n13 VN.t3 85.9021
R2554 VN.n25 VN.t9 85.9021
R2555 VN.n38 VN.t1 85.9021
R2556 VN.n0 VN.t7 85.9021
R2557 VN.n69 VN.t4 85.9021
R2558 VN.n65 VN.t2 85.9021
R2559 VN.n60 VN.t0 85.9021
R2560 VN.n54 VN.t6 85.9021
R2561 VN.n53 VN.n0 79.7913
R2562 VN.n107 VN.n54 79.7913
R2563 VN.n14 VN.n13 63.3588
R2564 VN.n70 VN.n69 63.3588
R2565 VN VN.n107 59.8844
R2566 VN.n19 VN.n10 56.5193
R2567 VN.n32 VN.n6 56.5193
R2568 VN.n45 VN.n2 56.5193
R2569 VN.n75 VN.n66 56.5193
R2570 VN.n87 VN.n61 56.5193
R2571 VN.n99 VN.n56 56.5193
R2572 VN.n17 VN.n12 24.4675
R2573 VN.n18 VN.n17 24.4675
R2574 VN.n19 VN.n18 24.4675
R2575 VN.n23 VN.n10 24.4675
R2576 VN.n24 VN.n23 24.4675
R2577 VN.n26 VN.n24 24.4675
R2578 VN.n30 VN.n8 24.4675
R2579 VN.n31 VN.n30 24.4675
R2580 VN.n32 VN.n31 24.4675
R2581 VN.n36 VN.n6 24.4675
R2582 VN.n37 VN.n36 24.4675
R2583 VN.n39 VN.n37 24.4675
R2584 VN.n43 VN.n4 24.4675
R2585 VN.n44 VN.n43 24.4675
R2586 VN.n45 VN.n44 24.4675
R2587 VN.n49 VN.n2 24.4675
R2588 VN.n50 VN.n49 24.4675
R2589 VN.n51 VN.n50 24.4675
R2590 VN.n75 VN.n74 24.4675
R2591 VN.n74 VN.n73 24.4675
R2592 VN.n73 VN.n68 24.4675
R2593 VN.n87 VN.n86 24.4675
R2594 VN.n86 VN.n85 24.4675
R2595 VN.n85 VN.n63 24.4675
R2596 VN.n81 VN.n80 24.4675
R2597 VN.n80 VN.n79 24.4675
R2598 VN.n79 VN.n66 24.4675
R2599 VN.n99 VN.n98 24.4675
R2600 VN.n98 VN.n97 24.4675
R2601 VN.n97 VN.n58 24.4675
R2602 VN.n93 VN.n92 24.4675
R2603 VN.n92 VN.n91 24.4675
R2604 VN.n91 VN.n61 24.4675
R2605 VN.n105 VN.n104 24.4675
R2606 VN.n104 VN.n103 24.4675
R2607 VN.n103 VN.n56 24.4675
R2608 VN.n38 VN.n4 13.2127
R2609 VN.n60 VN.n58 13.2127
R2610 VN.n26 VN.n25 12.234
R2611 VN.n25 VN.n8 12.234
R2612 VN.n65 VN.n63 12.234
R2613 VN.n81 VN.n65 12.234
R2614 VN.n13 VN.n12 11.2553
R2615 VN.n39 VN.n38 11.2553
R2616 VN.n69 VN.n68 11.2553
R2617 VN.n93 VN.n60 11.2553
R2618 VN.n51 VN.n0 10.2766
R2619 VN.n105 VN.n54 10.2766
R2620 VN.n71 VN.n70 3.14801
R2621 VN.n15 VN.n14 3.14801
R2622 VN.n107 VN.n106 0.354971
R2623 VN.n53 VN.n52 0.354971
R2624 VN VN.n53 0.26696
R2625 VN.n106 VN.n55 0.189894
R2626 VN.n102 VN.n55 0.189894
R2627 VN.n102 VN.n101 0.189894
R2628 VN.n101 VN.n100 0.189894
R2629 VN.n100 VN.n57 0.189894
R2630 VN.n96 VN.n57 0.189894
R2631 VN.n96 VN.n95 0.189894
R2632 VN.n95 VN.n94 0.189894
R2633 VN.n94 VN.n59 0.189894
R2634 VN.n90 VN.n59 0.189894
R2635 VN.n90 VN.n89 0.189894
R2636 VN.n89 VN.n88 0.189894
R2637 VN.n88 VN.n62 0.189894
R2638 VN.n84 VN.n62 0.189894
R2639 VN.n84 VN.n83 0.189894
R2640 VN.n83 VN.n82 0.189894
R2641 VN.n82 VN.n64 0.189894
R2642 VN.n78 VN.n64 0.189894
R2643 VN.n78 VN.n77 0.189894
R2644 VN.n77 VN.n76 0.189894
R2645 VN.n76 VN.n67 0.189894
R2646 VN.n72 VN.n67 0.189894
R2647 VN.n72 VN.n71 0.189894
R2648 VN.n16 VN.n15 0.189894
R2649 VN.n16 VN.n11 0.189894
R2650 VN.n20 VN.n11 0.189894
R2651 VN.n21 VN.n20 0.189894
R2652 VN.n22 VN.n21 0.189894
R2653 VN.n22 VN.n9 0.189894
R2654 VN.n27 VN.n9 0.189894
R2655 VN.n28 VN.n27 0.189894
R2656 VN.n29 VN.n28 0.189894
R2657 VN.n29 VN.n7 0.189894
R2658 VN.n33 VN.n7 0.189894
R2659 VN.n34 VN.n33 0.189894
R2660 VN.n35 VN.n34 0.189894
R2661 VN.n35 VN.n5 0.189894
R2662 VN.n40 VN.n5 0.189894
R2663 VN.n41 VN.n40 0.189894
R2664 VN.n42 VN.n41 0.189894
R2665 VN.n42 VN.n3 0.189894
R2666 VN.n46 VN.n3 0.189894
R2667 VN.n47 VN.n46 0.189894
R2668 VN.n48 VN.n47 0.189894
R2669 VN.n48 VN.n1 0.189894
R2670 VN.n52 VN.n1 0.189894
R2671 VDD2.n1 VDD2.t1 69.4257
R2672 VDD2.n3 VDD2.n2 66.9907
R2673 VDD2 VDD2.n7 66.9879
R2674 VDD2.n4 VDD2.t3 65.9958
R2675 VDD2.n6 VDD2.n5 64.4739
R2676 VDD2.n1 VDD2.n0 64.4728
R2677 VDD2.n4 VDD2.n3 51.2282
R2678 VDD2.n6 VDD2.n4 3.43153
R2679 VDD2.n7 VDD2.t5 1.52241
R2680 VDD2.n7 VDD2.t4 1.52241
R2681 VDD2.n5 VDD2.t9 1.52241
R2682 VDD2.n5 VDD2.t7 1.52241
R2683 VDD2.n2 VDD2.t8 1.52241
R2684 VDD2.n2 VDD2.t2 1.52241
R2685 VDD2.n0 VDD2.t6 1.52241
R2686 VDD2.n0 VDD2.t0 1.52241
R2687 VDD2 VDD2.n6 0.916448
R2688 VDD2.n3 VDD2.n1 0.802913
C0 VDD1 VDD2 2.85979f
C1 VN VP 10.131901f
C2 VTAIL VP 13.2672f
C3 VN VDD2 12.2085f
C4 VTAIL VDD2 11.3603f
C5 VN VDD1 0.155938f
C6 VTAIL VDD1 11.3016f
C7 VDD2 VP 0.717592f
C8 VN VTAIL 13.252701f
C9 VDD1 VP 12.7663f
C10 VDD2 B 8.604037f
C11 VDD1 B 8.584431f
C12 VTAIL B 9.415988f
C13 VN B 23.22063f
C14 VP B 21.799414f
C15 VDD2.t1 B 2.92721f
C16 VDD2.t6 B 0.2529f
C17 VDD2.t0 B 0.2529f
C18 VDD2.n0 B 2.27329f
C19 VDD2.n1 B 1.04532f
C20 VDD2.t8 B 0.2529f
C21 VDD2.t2 B 0.2529f
C22 VDD2.n2 B 2.29875f
C23 VDD2.n3 B 3.45248f
C24 VDD2.t3 B 2.90053f
C25 VDD2.n4 B 3.54355f
C26 VDD2.t9 B 0.2529f
C27 VDD2.t7 B 0.2529f
C28 VDD2.n5 B 2.2733f
C29 VDD2.n6 B 0.540237f
C30 VDD2.t5 B 0.2529f
C31 VDD2.t4 B 0.2529f
C32 VDD2.n7 B 2.2987f
C33 VN.t7 B 2.20296f
C34 VN.n0 B 0.837698f
C35 VN.n1 B 0.016989f
C36 VN.n2 B 0.026221f
C37 VN.n3 B 0.016989f
C38 VN.n4 B 0.024472f
C39 VN.n5 B 0.016989f
C40 VN.n6 B 0.025274f
C41 VN.n7 B 0.016989f
C42 VN.n8 B 0.023847f
C43 VN.n9 B 0.016989f
C44 VN.n10 B 0.024327f
C45 VN.n11 B 0.016989f
C46 VN.n12 B 0.023222f
C47 VN.t3 B 2.20296f
C48 VN.n13 B 0.828016f
C49 VN.t8 B 2.45513f
C50 VN.n14 B 0.784874f
C51 VN.n15 B 0.212877f
C52 VN.n16 B 0.016989f
C53 VN.n17 B 0.031663f
C54 VN.n18 B 0.031663f
C55 VN.n19 B 0.025274f
C56 VN.n20 B 0.016989f
C57 VN.n21 B 0.016989f
C58 VN.n22 B 0.016989f
C59 VN.n23 B 0.031663f
C60 VN.n24 B 0.031663f
C61 VN.t9 B 2.20296f
C62 VN.n25 B 0.769262f
C63 VN.n26 B 0.023847f
C64 VN.n27 B 0.016989f
C65 VN.n28 B 0.016989f
C66 VN.n29 B 0.016989f
C67 VN.n30 B 0.031663f
C68 VN.n31 B 0.031663f
C69 VN.n32 B 0.024327f
C70 VN.n33 B 0.016989f
C71 VN.n34 B 0.016989f
C72 VN.n35 B 0.016989f
C73 VN.n36 B 0.031663f
C74 VN.n37 B 0.031663f
C75 VN.t1 B 2.20296f
C76 VN.n38 B 0.769262f
C77 VN.n39 B 0.023222f
C78 VN.n40 B 0.016989f
C79 VN.n41 B 0.016989f
C80 VN.n42 B 0.016989f
C81 VN.n43 B 0.031663f
C82 VN.n44 B 0.031663f
C83 VN.n45 B 0.023381f
C84 VN.n46 B 0.016989f
C85 VN.n47 B 0.016989f
C86 VN.n48 B 0.016989f
C87 VN.n49 B 0.031663f
C88 VN.n50 B 0.031663f
C89 VN.n51 B 0.022596f
C90 VN.n52 B 0.02742f
C91 VN.n53 B 0.04666f
C92 VN.t6 B 2.20296f
C93 VN.n54 B 0.837698f
C94 VN.n55 B 0.016989f
C95 VN.n56 B 0.026221f
C96 VN.n57 B 0.016989f
C97 VN.n58 B 0.024472f
C98 VN.n59 B 0.016989f
C99 VN.t0 B 2.20296f
C100 VN.n60 B 0.769262f
C101 VN.n61 B 0.025274f
C102 VN.n62 B 0.016989f
C103 VN.n63 B 0.023847f
C104 VN.n64 B 0.016989f
C105 VN.t2 B 2.20296f
C106 VN.n65 B 0.769262f
C107 VN.n66 B 0.024327f
C108 VN.n67 B 0.016989f
C109 VN.n68 B 0.023222f
C110 VN.t5 B 2.45513f
C111 VN.t4 B 2.20296f
C112 VN.n69 B 0.828016f
C113 VN.n70 B 0.784874f
C114 VN.n71 B 0.212877f
C115 VN.n72 B 0.016989f
C116 VN.n73 B 0.031663f
C117 VN.n74 B 0.031663f
C118 VN.n75 B 0.025274f
C119 VN.n76 B 0.016989f
C120 VN.n77 B 0.016989f
C121 VN.n78 B 0.016989f
C122 VN.n79 B 0.031663f
C123 VN.n80 B 0.031663f
C124 VN.n81 B 0.023847f
C125 VN.n82 B 0.016989f
C126 VN.n83 B 0.016989f
C127 VN.n84 B 0.016989f
C128 VN.n85 B 0.031663f
C129 VN.n86 B 0.031663f
C130 VN.n87 B 0.024327f
C131 VN.n88 B 0.016989f
C132 VN.n89 B 0.016989f
C133 VN.n90 B 0.016989f
C134 VN.n91 B 0.031663f
C135 VN.n92 B 0.031663f
C136 VN.n93 B 0.023222f
C137 VN.n94 B 0.016989f
C138 VN.n95 B 0.016989f
C139 VN.n96 B 0.016989f
C140 VN.n97 B 0.031663f
C141 VN.n98 B 0.031663f
C142 VN.n99 B 0.023381f
C143 VN.n100 B 0.016989f
C144 VN.n101 B 0.016989f
C145 VN.n102 B 0.016989f
C146 VN.n103 B 0.031663f
C147 VN.n104 B 0.031663f
C148 VN.n105 B 0.022596f
C149 VN.n106 B 0.02742f
C150 VN.n107 B 1.24939f
C151 VDD1.t5 B 2.97226f
C152 VDD1.t6 B 0.256791f
C153 VDD1.t9 B 0.256791f
C154 VDD1.n0 B 2.30827f
C155 VDD1.n1 B 1.0698f
C156 VDD1.t2 B 2.97225f
C157 VDD1.t8 B 0.256791f
C158 VDD1.t0 B 0.256791f
C159 VDD1.n2 B 2.30827f
C160 VDD1.n3 B 1.0614f
C161 VDD1.t4 B 0.256791f
C162 VDD1.t1 B 0.256791f
C163 VDD1.n4 B 2.33412f
C164 VDD1.n5 B 3.66021f
C165 VDD1.t3 B 0.256791f
C166 VDD1.t7 B 0.256791f
C167 VDD1.n6 B 2.30827f
C168 VDD1.n7 B 3.67469f
C169 VTAIL.t16 B 0.261931f
C170 VTAIL.t4 B 0.261931f
C171 VTAIL.n0 B 2.28543f
C172 VTAIL.n1 B 0.632512f
C173 VTAIL.t5 B 2.91529f
C174 VTAIL.n2 B 0.782646f
C175 VTAIL.t8 B 0.261931f
C176 VTAIL.t14 B 0.261931f
C177 VTAIL.n3 B 2.28543f
C178 VTAIL.n4 B 0.800415f
C179 VTAIL.t9 B 0.261931f
C180 VTAIL.t13 B 0.261931f
C181 VTAIL.n5 B 2.28543f
C182 VTAIL.n6 B 2.34889f
C183 VTAIL.t3 B 0.261931f
C184 VTAIL.t0 B 0.261931f
C185 VTAIL.n7 B 2.28544f
C186 VTAIL.n8 B 2.34888f
C187 VTAIL.t1 B 0.261931f
C188 VTAIL.t19 B 0.261931f
C189 VTAIL.n9 B 2.28544f
C190 VTAIL.n10 B 0.800404f
C191 VTAIL.t18 B 2.91531f
C192 VTAIL.n11 B 0.782629f
C193 VTAIL.t6 B 0.261931f
C194 VTAIL.t11 B 0.261931f
C195 VTAIL.n12 B 2.28544f
C196 VTAIL.n13 B 0.698141f
C197 VTAIL.t7 B 0.261931f
C198 VTAIL.t10 B 0.261931f
C199 VTAIL.n14 B 2.28544f
C200 VTAIL.n15 B 0.800404f
C201 VTAIL.t12 B 2.91529f
C202 VTAIL.n16 B 2.15172f
C203 VTAIL.t2 B 2.91529f
C204 VTAIL.n17 B 2.15172f
C205 VTAIL.t17 B 0.261931f
C206 VTAIL.t15 B 0.261931f
C207 VTAIL.n18 B 2.28543f
C208 VTAIL.n19 B 0.584388f
C209 VP.t8 B 2.24159f
C210 VP.n0 B 0.852389f
C211 VP.n1 B 0.017287f
C212 VP.n2 B 0.026681f
C213 VP.n3 B 0.017287f
C214 VP.n4 B 0.024902f
C215 VP.n5 B 0.017287f
C216 VP.n6 B 0.025718f
C217 VP.n7 B 0.017287f
C218 VP.n8 B 0.024265f
C219 VP.n9 B 0.017287f
C220 VP.n10 B 0.024754f
C221 VP.n11 B 0.017287f
C222 VP.n12 B 0.023629f
C223 VP.n13 B 0.017287f
C224 VP.n14 B 0.023791f
C225 VP.n15 B 0.017287f
C226 VP.n16 B 0.022993f
C227 VP.t2 B 2.24159f
C228 VP.n17 B 0.852389f
C229 VP.n18 B 0.017287f
C230 VP.n19 B 0.026681f
C231 VP.n20 B 0.017287f
C232 VP.n21 B 0.024902f
C233 VP.n22 B 0.017287f
C234 VP.n23 B 0.025718f
C235 VP.n24 B 0.017287f
C236 VP.n25 B 0.024265f
C237 VP.n26 B 0.017287f
C238 VP.n27 B 0.024754f
C239 VP.n28 B 0.017287f
C240 VP.n29 B 0.023629f
C241 VP.t4 B 2.49818f
C242 VP.t3 B 2.24159f
C243 VP.n30 B 0.842536f
C244 VP.n31 B 0.798638f
C245 VP.n32 B 0.216611f
C246 VP.n33 B 0.017287f
C247 VP.n34 B 0.032219f
C248 VP.n35 B 0.032219f
C249 VP.n36 B 0.025718f
C250 VP.n37 B 0.017287f
C251 VP.n38 B 0.017287f
C252 VP.n39 B 0.017287f
C253 VP.n40 B 0.032219f
C254 VP.n41 B 0.032219f
C255 VP.t0 B 2.24159f
C256 VP.n42 B 0.782752f
C257 VP.n43 B 0.024265f
C258 VP.n44 B 0.017287f
C259 VP.n45 B 0.017287f
C260 VP.n46 B 0.017287f
C261 VP.n47 B 0.032219f
C262 VP.n48 B 0.032219f
C263 VP.n49 B 0.024754f
C264 VP.n50 B 0.017287f
C265 VP.n51 B 0.017287f
C266 VP.n52 B 0.017287f
C267 VP.n53 B 0.032219f
C268 VP.n54 B 0.032219f
C269 VP.t6 B 2.24159f
C270 VP.n55 B 0.782752f
C271 VP.n56 B 0.023629f
C272 VP.n57 B 0.017287f
C273 VP.n58 B 0.017287f
C274 VP.n59 B 0.017287f
C275 VP.n60 B 0.032219f
C276 VP.n61 B 0.032219f
C277 VP.n62 B 0.023791f
C278 VP.n63 B 0.017287f
C279 VP.n64 B 0.017287f
C280 VP.n65 B 0.017287f
C281 VP.n66 B 0.032219f
C282 VP.n67 B 0.032219f
C283 VP.n68 B 0.022993f
C284 VP.n69 B 0.027901f
C285 VP.n70 B 1.26463f
C286 VP.t7 B 2.24159f
C287 VP.n71 B 0.852389f
C288 VP.n72 B 1.27504f
C289 VP.n73 B 0.027901f
C290 VP.n74 B 0.017287f
C291 VP.n75 B 0.032219f
C292 VP.n76 B 0.032219f
C293 VP.n77 B 0.026681f
C294 VP.n78 B 0.017287f
C295 VP.n79 B 0.017287f
C296 VP.n80 B 0.017287f
C297 VP.n81 B 0.032219f
C298 VP.n82 B 0.032219f
C299 VP.t1 B 2.24159f
C300 VP.n83 B 0.782752f
C301 VP.n84 B 0.024902f
C302 VP.n85 B 0.017287f
C303 VP.n86 B 0.017287f
C304 VP.n87 B 0.017287f
C305 VP.n88 B 0.032219f
C306 VP.n89 B 0.032219f
C307 VP.n90 B 0.025718f
C308 VP.n91 B 0.017287f
C309 VP.n92 B 0.017287f
C310 VP.n93 B 0.017287f
C311 VP.n94 B 0.032219f
C312 VP.n95 B 0.032219f
C313 VP.t9 B 2.24159f
C314 VP.n96 B 0.782752f
C315 VP.n97 B 0.024265f
C316 VP.n98 B 0.017287f
C317 VP.n99 B 0.017287f
C318 VP.n100 B 0.017287f
C319 VP.n101 B 0.032219f
C320 VP.n102 B 0.032219f
C321 VP.n103 B 0.024754f
C322 VP.n104 B 0.017287f
C323 VP.n105 B 0.017287f
C324 VP.n106 B 0.017287f
C325 VP.n107 B 0.032219f
C326 VP.n108 B 0.032219f
C327 VP.t5 B 2.24159f
C328 VP.n109 B 0.782752f
C329 VP.n110 B 0.023629f
C330 VP.n111 B 0.017287f
C331 VP.n112 B 0.017287f
C332 VP.n113 B 0.017287f
C333 VP.n114 B 0.032219f
C334 VP.n115 B 0.032219f
C335 VP.n116 B 0.023791f
C336 VP.n117 B 0.017287f
C337 VP.n118 B 0.017287f
C338 VP.n119 B 0.017287f
C339 VP.n120 B 0.032219f
C340 VP.n121 B 0.032219f
C341 VP.n122 B 0.022993f
C342 VP.n123 B 0.027901f
C343 VP.n124 B 0.047478f
.ends

