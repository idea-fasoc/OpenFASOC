* NGSPICE file created from diff_pair_sample_1569.ext - technology: sky130A

.subckt diff_pair_sample_1569 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t19 VN.t0 VDD2.t1 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X1 B.t23 B.t21 B.t22 B.t11 sky130_fd_pr__nfet_01v8 ad=7.0122 pd=36.74 as=0 ps=0 w=17.98 l=1.42
X2 VDD2.t0 VN.t1 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=7.0122 pd=36.74 as=2.9667 ps=18.31 w=17.98 l=1.42
X3 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=7.0122 pd=36.74 as=0 ps=0 w=17.98 l=1.42
X4 VDD1.t9 VP.t0 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X5 VTAIL.t8 VP.t1 VDD1.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X6 VDD1.t7 VP.t2 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=7.0122 pd=36.74 as=2.9667 ps=18.31 w=17.98 l=1.42
X7 VTAIL.t17 VN.t2 VDD2.t7 B.t8 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X8 VTAIL.t16 VN.t3 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X9 VTAIL.t6 VP.t3 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X10 VDD2.t3 VN.t4 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=7.0122 pd=36.74 as=2.9667 ps=18.31 w=17.98 l=1.42
X11 VDD2.t2 VN.t5 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X12 VDD2.t9 VN.t6 VTAIL.t13 B.t7 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X13 VTAIL.t2 VP.t4 VDD1.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X14 VDD1.t4 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=7.0122 ps=36.74 w=17.98 l=1.42
X15 VDD2.t8 VN.t7 VTAIL.t12 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=7.0122 ps=36.74 w=17.98 l=1.42
X16 VDD1.t3 VP.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X17 VTAIL.t3 VP.t7 VDD1.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X18 VTAIL.t11 VN.t8 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=2.9667 ps=18.31 w=17.98 l=1.42
X19 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=7.0122 pd=36.74 as=0 ps=0 w=17.98 l=1.42
X20 VDD1.t1 VP.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=7.0122 pd=36.74 as=2.9667 ps=18.31 w=17.98 l=1.42
X21 VDD2.t4 VN.t9 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=7.0122 ps=36.74 w=17.98 l=1.42
X22 VDD1.t0 VP.t9 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9667 pd=18.31 as=7.0122 ps=36.74 w=17.98 l=1.42
X23 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.0122 pd=36.74 as=0 ps=0 w=17.98 l=1.42
R0 VN.n6 VN.t1 340.659
R1 VN.n32 VN.t7 340.659
R2 VN.n17 VN.t0 305.154
R3 VN.n5 VN.t8 305.154
R4 VN.n10 VN.t5 305.154
R5 VN.n23 VN.t9 305.154
R6 VN.n42 VN.t3 305.154
R7 VN.n31 VN.t2 305.154
R8 VN.n30 VN.t6 305.154
R9 VN.n48 VN.t4 305.154
R10 VN.n24 VN.n23 173.596
R11 VN.n49 VN.n48 173.596
R12 VN.n47 VN.n25 161.3
R13 VN.n46 VN.n45 161.3
R14 VN.n44 VN.n26 161.3
R15 VN.n43 VN.n42 161.3
R16 VN.n41 VN.n27 161.3
R17 VN.n40 VN.n39 161.3
R18 VN.n38 VN.n28 161.3
R19 VN.n37 VN.n36 161.3
R20 VN.n35 VN.n29 161.3
R21 VN.n34 VN.n33 161.3
R22 VN.n22 VN.n0 161.3
R23 VN.n21 VN.n20 161.3
R24 VN.n19 VN.n1 161.3
R25 VN.n18 VN.n17 161.3
R26 VN.n16 VN.n2 161.3
R27 VN.n15 VN.n14 161.3
R28 VN.n13 VN.n3 161.3
R29 VN.n12 VN.n11 161.3
R30 VN.n9 VN.n4 161.3
R31 VN.n8 VN.n7 161.3
R32 VN.n9 VN.n8 52.6866
R33 VN.n16 VN.n15 52.6866
R34 VN.n21 VN.n1 52.6866
R35 VN.n35 VN.n34 52.6866
R36 VN.n41 VN.n40 52.6866
R37 VN.n46 VN.n26 52.6866
R38 VN VN.n49 51.5516
R39 VN.n6 VN.n5 41.915
R40 VN.n32 VN.n31 41.915
R41 VN.n11 VN.n9 28.4674
R42 VN.n15 VN.n3 28.4674
R43 VN.n22 VN.n21 28.4674
R44 VN.n36 VN.n35 28.4674
R45 VN.n40 VN.n28 28.4674
R46 VN.n47 VN.n46 28.4674
R47 VN.n8 VN.n5 24.5923
R48 VN.n17 VN.n16 24.5923
R49 VN.n17 VN.n1 24.5923
R50 VN.n34 VN.n31 24.5923
R51 VN.n42 VN.n26 24.5923
R52 VN.n42 VN.n41 24.5923
R53 VN.n33 VN.n32 17.507
R54 VN.n7 VN.n6 17.507
R55 VN.n11 VN.n10 12.2964
R56 VN.n10 VN.n3 12.2964
R57 VN.n23 VN.n22 12.2964
R58 VN.n30 VN.n28 12.2964
R59 VN.n36 VN.n30 12.2964
R60 VN.n48 VN.n47 12.2964
R61 VN.n49 VN.n25 0.189894
R62 VN.n45 VN.n25 0.189894
R63 VN.n45 VN.n44 0.189894
R64 VN.n44 VN.n43 0.189894
R65 VN.n43 VN.n27 0.189894
R66 VN.n39 VN.n27 0.189894
R67 VN.n39 VN.n38 0.189894
R68 VN.n38 VN.n37 0.189894
R69 VN.n37 VN.n29 0.189894
R70 VN.n33 VN.n29 0.189894
R71 VN.n7 VN.n4 0.189894
R72 VN.n12 VN.n4 0.189894
R73 VN.n13 VN.n12 0.189894
R74 VN.n14 VN.n13 0.189894
R75 VN.n14 VN.n2 0.189894
R76 VN.n18 VN.n2 0.189894
R77 VN.n19 VN.n18 0.189894
R78 VN.n20 VN.n19 0.189894
R79 VN.n20 VN.n0 0.189894
R80 VN.n24 VN.n0 0.189894
R81 VN VN.n24 0.0516364
R82 VDD2.n1 VDD2.t0 65.213
R83 VDD2.n4 VDD2.t3 63.7046
R84 VDD2.n3 VDD2.n2 63.6793
R85 VDD2 VDD2.n7 63.6765
R86 VDD2.n6 VDD2.n5 62.6034
R87 VDD2.n1 VDD2.n0 62.6032
R88 VDD2.n4 VDD2.n3 46.3812
R89 VDD2.n6 VDD2.n4 1.50912
R90 VDD2.n7 VDD2.t7 1.10172
R91 VDD2.n7 VDD2.t8 1.10172
R92 VDD2.n5 VDD2.t6 1.10172
R93 VDD2.n5 VDD2.t9 1.10172
R94 VDD2.n2 VDD2.t1 1.10172
R95 VDD2.n2 VDD2.t4 1.10172
R96 VDD2.n0 VDD2.t5 1.10172
R97 VDD2.n0 VDD2.t2 1.10172
R98 VDD2 VDD2.n6 0.435845
R99 VDD2.n3 VDD2.n1 0.322309
R100 VTAIL.n11 VTAIL.t12 47.0258
R101 VTAIL.n17 VTAIL.t10 47.0256
R102 VTAIL.n2 VTAIL.t1 47.0256
R103 VTAIL.n16 VTAIL.t4 47.0256
R104 VTAIL.n15 VTAIL.n14 45.9246
R105 VTAIL.n13 VTAIL.n12 45.9246
R106 VTAIL.n10 VTAIL.n9 45.9246
R107 VTAIL.n8 VTAIL.n7 45.9246
R108 VTAIL.n19 VTAIL.n18 45.9244
R109 VTAIL.n1 VTAIL.n0 45.9244
R110 VTAIL.n4 VTAIL.n3 45.9244
R111 VTAIL.n6 VTAIL.n5 45.9244
R112 VTAIL.n8 VTAIL.n6 30.8841
R113 VTAIL.n17 VTAIL.n16 29.3755
R114 VTAIL.n10 VTAIL.n8 1.50912
R115 VTAIL.n11 VTAIL.n10 1.50912
R116 VTAIL.n15 VTAIL.n13 1.50912
R117 VTAIL.n16 VTAIL.n15 1.50912
R118 VTAIL.n6 VTAIL.n4 1.50912
R119 VTAIL.n4 VTAIL.n2 1.50912
R120 VTAIL.n19 VTAIL.n17 1.50912
R121 VTAIL.n13 VTAIL.n11 1.22464
R122 VTAIL.n2 VTAIL.n1 1.22464
R123 VTAIL VTAIL.n1 1.19016
R124 VTAIL.n18 VTAIL.t14 1.10172
R125 VTAIL.n18 VTAIL.t19 1.10172
R126 VTAIL.n0 VTAIL.t18 1.10172
R127 VTAIL.n0 VTAIL.t11 1.10172
R128 VTAIL.n3 VTAIL.t7 1.10172
R129 VTAIL.n3 VTAIL.t8 1.10172
R130 VTAIL.n5 VTAIL.t9 1.10172
R131 VTAIL.n5 VTAIL.t2 1.10172
R132 VTAIL.n14 VTAIL.t0 1.10172
R133 VTAIL.n14 VTAIL.t6 1.10172
R134 VTAIL.n12 VTAIL.t5 1.10172
R135 VTAIL.n12 VTAIL.t3 1.10172
R136 VTAIL.n9 VTAIL.t13 1.10172
R137 VTAIL.n9 VTAIL.t17 1.10172
R138 VTAIL.n7 VTAIL.t15 1.10172
R139 VTAIL.n7 VTAIL.t16 1.10172
R140 VTAIL VTAIL.n19 0.319466
R141 B.n962 B.n961 585
R142 B.n393 B.n137 585
R143 B.n392 B.n391 585
R144 B.n390 B.n389 585
R145 B.n388 B.n387 585
R146 B.n386 B.n385 585
R147 B.n384 B.n383 585
R148 B.n382 B.n381 585
R149 B.n380 B.n379 585
R150 B.n378 B.n377 585
R151 B.n376 B.n375 585
R152 B.n374 B.n373 585
R153 B.n372 B.n371 585
R154 B.n370 B.n369 585
R155 B.n368 B.n367 585
R156 B.n366 B.n365 585
R157 B.n364 B.n363 585
R158 B.n362 B.n361 585
R159 B.n360 B.n359 585
R160 B.n358 B.n357 585
R161 B.n356 B.n355 585
R162 B.n354 B.n353 585
R163 B.n352 B.n351 585
R164 B.n350 B.n349 585
R165 B.n348 B.n347 585
R166 B.n346 B.n345 585
R167 B.n344 B.n343 585
R168 B.n342 B.n341 585
R169 B.n340 B.n339 585
R170 B.n338 B.n337 585
R171 B.n336 B.n335 585
R172 B.n334 B.n333 585
R173 B.n332 B.n331 585
R174 B.n330 B.n329 585
R175 B.n328 B.n327 585
R176 B.n326 B.n325 585
R177 B.n324 B.n323 585
R178 B.n322 B.n321 585
R179 B.n320 B.n319 585
R180 B.n318 B.n317 585
R181 B.n316 B.n315 585
R182 B.n314 B.n313 585
R183 B.n312 B.n311 585
R184 B.n310 B.n309 585
R185 B.n308 B.n307 585
R186 B.n306 B.n305 585
R187 B.n304 B.n303 585
R188 B.n302 B.n301 585
R189 B.n300 B.n299 585
R190 B.n298 B.n297 585
R191 B.n296 B.n295 585
R192 B.n294 B.n293 585
R193 B.n292 B.n291 585
R194 B.n290 B.n289 585
R195 B.n288 B.n287 585
R196 B.n286 B.n285 585
R197 B.n284 B.n283 585
R198 B.n282 B.n281 585
R199 B.n280 B.n279 585
R200 B.n277 B.n276 585
R201 B.n275 B.n274 585
R202 B.n273 B.n272 585
R203 B.n271 B.n270 585
R204 B.n269 B.n268 585
R205 B.n267 B.n266 585
R206 B.n265 B.n264 585
R207 B.n263 B.n262 585
R208 B.n261 B.n260 585
R209 B.n259 B.n258 585
R210 B.n256 B.n255 585
R211 B.n254 B.n253 585
R212 B.n252 B.n251 585
R213 B.n250 B.n249 585
R214 B.n248 B.n247 585
R215 B.n246 B.n245 585
R216 B.n244 B.n243 585
R217 B.n242 B.n241 585
R218 B.n240 B.n239 585
R219 B.n238 B.n237 585
R220 B.n236 B.n235 585
R221 B.n234 B.n233 585
R222 B.n232 B.n231 585
R223 B.n230 B.n229 585
R224 B.n228 B.n227 585
R225 B.n226 B.n225 585
R226 B.n224 B.n223 585
R227 B.n222 B.n221 585
R228 B.n220 B.n219 585
R229 B.n218 B.n217 585
R230 B.n216 B.n215 585
R231 B.n214 B.n213 585
R232 B.n212 B.n211 585
R233 B.n210 B.n209 585
R234 B.n208 B.n207 585
R235 B.n206 B.n205 585
R236 B.n204 B.n203 585
R237 B.n202 B.n201 585
R238 B.n200 B.n199 585
R239 B.n198 B.n197 585
R240 B.n196 B.n195 585
R241 B.n194 B.n193 585
R242 B.n192 B.n191 585
R243 B.n190 B.n189 585
R244 B.n188 B.n187 585
R245 B.n186 B.n185 585
R246 B.n184 B.n183 585
R247 B.n182 B.n181 585
R248 B.n180 B.n179 585
R249 B.n178 B.n177 585
R250 B.n176 B.n175 585
R251 B.n174 B.n173 585
R252 B.n172 B.n171 585
R253 B.n170 B.n169 585
R254 B.n168 B.n167 585
R255 B.n166 B.n165 585
R256 B.n164 B.n163 585
R257 B.n162 B.n161 585
R258 B.n160 B.n159 585
R259 B.n158 B.n157 585
R260 B.n156 B.n155 585
R261 B.n154 B.n153 585
R262 B.n152 B.n151 585
R263 B.n150 B.n149 585
R264 B.n148 B.n147 585
R265 B.n146 B.n145 585
R266 B.n144 B.n143 585
R267 B.n74 B.n73 585
R268 B.n967 B.n966 585
R269 B.n960 B.n138 585
R270 B.n138 B.n71 585
R271 B.n959 B.n70 585
R272 B.n971 B.n70 585
R273 B.n958 B.n69 585
R274 B.n972 B.n69 585
R275 B.n957 B.n68 585
R276 B.n973 B.n68 585
R277 B.n956 B.n955 585
R278 B.n955 B.n64 585
R279 B.n954 B.n63 585
R280 B.n979 B.n63 585
R281 B.n953 B.n62 585
R282 B.n980 B.n62 585
R283 B.n952 B.n61 585
R284 B.n981 B.n61 585
R285 B.n951 B.n950 585
R286 B.n950 B.n57 585
R287 B.n949 B.n56 585
R288 B.n987 B.n56 585
R289 B.n948 B.n55 585
R290 B.n988 B.n55 585
R291 B.n947 B.n54 585
R292 B.n989 B.n54 585
R293 B.n946 B.n945 585
R294 B.n945 B.n50 585
R295 B.n944 B.n49 585
R296 B.n995 B.n49 585
R297 B.n943 B.n48 585
R298 B.n996 B.n48 585
R299 B.n942 B.n47 585
R300 B.n997 B.n47 585
R301 B.n941 B.n940 585
R302 B.n940 B.n43 585
R303 B.n939 B.n42 585
R304 B.n1003 B.n42 585
R305 B.n938 B.n41 585
R306 B.n1004 B.n41 585
R307 B.n937 B.n40 585
R308 B.n1005 B.n40 585
R309 B.n936 B.n935 585
R310 B.n935 B.n36 585
R311 B.n934 B.n35 585
R312 B.n1011 B.n35 585
R313 B.n933 B.n34 585
R314 B.n1012 B.n34 585
R315 B.n932 B.n33 585
R316 B.n1013 B.n33 585
R317 B.n931 B.n930 585
R318 B.n930 B.n32 585
R319 B.n929 B.n28 585
R320 B.n1019 B.n28 585
R321 B.n928 B.n27 585
R322 B.n1020 B.n27 585
R323 B.n927 B.n26 585
R324 B.n1021 B.n26 585
R325 B.n926 B.n925 585
R326 B.n925 B.n22 585
R327 B.n924 B.n21 585
R328 B.n1027 B.n21 585
R329 B.n923 B.n20 585
R330 B.n1028 B.n20 585
R331 B.n922 B.n19 585
R332 B.n1029 B.n19 585
R333 B.n921 B.n920 585
R334 B.n920 B.n15 585
R335 B.n919 B.n14 585
R336 B.n1035 B.n14 585
R337 B.n918 B.n13 585
R338 B.n1036 B.n13 585
R339 B.n917 B.n12 585
R340 B.n1037 B.n12 585
R341 B.n916 B.n915 585
R342 B.n915 B.n8 585
R343 B.n914 B.n7 585
R344 B.n1043 B.n7 585
R345 B.n913 B.n6 585
R346 B.n1044 B.n6 585
R347 B.n912 B.n5 585
R348 B.n1045 B.n5 585
R349 B.n911 B.n910 585
R350 B.n910 B.n4 585
R351 B.n909 B.n394 585
R352 B.n909 B.n908 585
R353 B.n899 B.n395 585
R354 B.n396 B.n395 585
R355 B.n901 B.n900 585
R356 B.n902 B.n901 585
R357 B.n898 B.n400 585
R358 B.n404 B.n400 585
R359 B.n897 B.n896 585
R360 B.n896 B.n895 585
R361 B.n402 B.n401 585
R362 B.n403 B.n402 585
R363 B.n888 B.n887 585
R364 B.n889 B.n888 585
R365 B.n886 B.n409 585
R366 B.n409 B.n408 585
R367 B.n885 B.n884 585
R368 B.n884 B.n883 585
R369 B.n411 B.n410 585
R370 B.n412 B.n411 585
R371 B.n876 B.n875 585
R372 B.n877 B.n876 585
R373 B.n874 B.n417 585
R374 B.n417 B.n416 585
R375 B.n873 B.n872 585
R376 B.n872 B.n871 585
R377 B.n419 B.n418 585
R378 B.n864 B.n419 585
R379 B.n863 B.n862 585
R380 B.n865 B.n863 585
R381 B.n861 B.n424 585
R382 B.n424 B.n423 585
R383 B.n860 B.n859 585
R384 B.n859 B.n858 585
R385 B.n426 B.n425 585
R386 B.n427 B.n426 585
R387 B.n851 B.n850 585
R388 B.n852 B.n851 585
R389 B.n849 B.n432 585
R390 B.n432 B.n431 585
R391 B.n848 B.n847 585
R392 B.n847 B.n846 585
R393 B.n434 B.n433 585
R394 B.n435 B.n434 585
R395 B.n839 B.n838 585
R396 B.n840 B.n839 585
R397 B.n837 B.n439 585
R398 B.n443 B.n439 585
R399 B.n836 B.n835 585
R400 B.n835 B.n834 585
R401 B.n441 B.n440 585
R402 B.n442 B.n441 585
R403 B.n827 B.n826 585
R404 B.n828 B.n827 585
R405 B.n825 B.n448 585
R406 B.n448 B.n447 585
R407 B.n824 B.n823 585
R408 B.n823 B.n822 585
R409 B.n450 B.n449 585
R410 B.n451 B.n450 585
R411 B.n815 B.n814 585
R412 B.n816 B.n815 585
R413 B.n813 B.n456 585
R414 B.n456 B.n455 585
R415 B.n812 B.n811 585
R416 B.n811 B.n810 585
R417 B.n458 B.n457 585
R418 B.n459 B.n458 585
R419 B.n803 B.n802 585
R420 B.n804 B.n803 585
R421 B.n801 B.n464 585
R422 B.n464 B.n463 585
R423 B.n800 B.n799 585
R424 B.n799 B.n798 585
R425 B.n466 B.n465 585
R426 B.n467 B.n466 585
R427 B.n794 B.n793 585
R428 B.n470 B.n469 585
R429 B.n790 B.n789 585
R430 B.n791 B.n790 585
R431 B.n788 B.n534 585
R432 B.n787 B.n786 585
R433 B.n785 B.n784 585
R434 B.n783 B.n782 585
R435 B.n781 B.n780 585
R436 B.n779 B.n778 585
R437 B.n777 B.n776 585
R438 B.n775 B.n774 585
R439 B.n773 B.n772 585
R440 B.n771 B.n770 585
R441 B.n769 B.n768 585
R442 B.n767 B.n766 585
R443 B.n765 B.n764 585
R444 B.n763 B.n762 585
R445 B.n761 B.n760 585
R446 B.n759 B.n758 585
R447 B.n757 B.n756 585
R448 B.n755 B.n754 585
R449 B.n753 B.n752 585
R450 B.n751 B.n750 585
R451 B.n749 B.n748 585
R452 B.n747 B.n746 585
R453 B.n745 B.n744 585
R454 B.n743 B.n742 585
R455 B.n741 B.n740 585
R456 B.n739 B.n738 585
R457 B.n737 B.n736 585
R458 B.n735 B.n734 585
R459 B.n733 B.n732 585
R460 B.n731 B.n730 585
R461 B.n729 B.n728 585
R462 B.n727 B.n726 585
R463 B.n725 B.n724 585
R464 B.n723 B.n722 585
R465 B.n721 B.n720 585
R466 B.n719 B.n718 585
R467 B.n717 B.n716 585
R468 B.n715 B.n714 585
R469 B.n713 B.n712 585
R470 B.n711 B.n710 585
R471 B.n709 B.n708 585
R472 B.n707 B.n706 585
R473 B.n705 B.n704 585
R474 B.n703 B.n702 585
R475 B.n701 B.n700 585
R476 B.n699 B.n698 585
R477 B.n697 B.n696 585
R478 B.n695 B.n694 585
R479 B.n693 B.n692 585
R480 B.n691 B.n690 585
R481 B.n689 B.n688 585
R482 B.n687 B.n686 585
R483 B.n685 B.n684 585
R484 B.n683 B.n682 585
R485 B.n681 B.n680 585
R486 B.n679 B.n678 585
R487 B.n677 B.n676 585
R488 B.n675 B.n674 585
R489 B.n673 B.n672 585
R490 B.n671 B.n670 585
R491 B.n669 B.n668 585
R492 B.n667 B.n666 585
R493 B.n665 B.n664 585
R494 B.n663 B.n662 585
R495 B.n661 B.n660 585
R496 B.n659 B.n658 585
R497 B.n657 B.n656 585
R498 B.n655 B.n654 585
R499 B.n653 B.n652 585
R500 B.n651 B.n650 585
R501 B.n649 B.n648 585
R502 B.n647 B.n646 585
R503 B.n645 B.n644 585
R504 B.n643 B.n642 585
R505 B.n641 B.n640 585
R506 B.n639 B.n638 585
R507 B.n637 B.n636 585
R508 B.n635 B.n634 585
R509 B.n633 B.n632 585
R510 B.n631 B.n630 585
R511 B.n629 B.n628 585
R512 B.n627 B.n626 585
R513 B.n625 B.n624 585
R514 B.n623 B.n622 585
R515 B.n621 B.n620 585
R516 B.n619 B.n618 585
R517 B.n617 B.n616 585
R518 B.n615 B.n614 585
R519 B.n613 B.n612 585
R520 B.n611 B.n610 585
R521 B.n609 B.n608 585
R522 B.n607 B.n606 585
R523 B.n605 B.n604 585
R524 B.n603 B.n602 585
R525 B.n601 B.n600 585
R526 B.n599 B.n598 585
R527 B.n597 B.n596 585
R528 B.n595 B.n594 585
R529 B.n593 B.n592 585
R530 B.n591 B.n590 585
R531 B.n589 B.n588 585
R532 B.n587 B.n586 585
R533 B.n585 B.n584 585
R534 B.n583 B.n582 585
R535 B.n581 B.n580 585
R536 B.n579 B.n578 585
R537 B.n577 B.n576 585
R538 B.n575 B.n574 585
R539 B.n573 B.n572 585
R540 B.n571 B.n570 585
R541 B.n569 B.n568 585
R542 B.n567 B.n566 585
R543 B.n565 B.n564 585
R544 B.n563 B.n562 585
R545 B.n561 B.n560 585
R546 B.n559 B.n558 585
R547 B.n557 B.n556 585
R548 B.n555 B.n554 585
R549 B.n553 B.n552 585
R550 B.n551 B.n550 585
R551 B.n549 B.n548 585
R552 B.n547 B.n546 585
R553 B.n545 B.n544 585
R554 B.n543 B.n542 585
R555 B.n541 B.n533 585
R556 B.n791 B.n533 585
R557 B.n795 B.n468 585
R558 B.n468 B.n467 585
R559 B.n797 B.n796 585
R560 B.n798 B.n797 585
R561 B.n462 B.n461 585
R562 B.n463 B.n462 585
R563 B.n806 B.n805 585
R564 B.n805 B.n804 585
R565 B.n807 B.n460 585
R566 B.n460 B.n459 585
R567 B.n809 B.n808 585
R568 B.n810 B.n809 585
R569 B.n454 B.n453 585
R570 B.n455 B.n454 585
R571 B.n818 B.n817 585
R572 B.n817 B.n816 585
R573 B.n819 B.n452 585
R574 B.n452 B.n451 585
R575 B.n821 B.n820 585
R576 B.n822 B.n821 585
R577 B.n446 B.n445 585
R578 B.n447 B.n446 585
R579 B.n830 B.n829 585
R580 B.n829 B.n828 585
R581 B.n831 B.n444 585
R582 B.n444 B.n442 585
R583 B.n833 B.n832 585
R584 B.n834 B.n833 585
R585 B.n438 B.n437 585
R586 B.n443 B.n438 585
R587 B.n842 B.n841 585
R588 B.n841 B.n840 585
R589 B.n843 B.n436 585
R590 B.n436 B.n435 585
R591 B.n845 B.n844 585
R592 B.n846 B.n845 585
R593 B.n430 B.n429 585
R594 B.n431 B.n430 585
R595 B.n854 B.n853 585
R596 B.n853 B.n852 585
R597 B.n855 B.n428 585
R598 B.n428 B.n427 585
R599 B.n857 B.n856 585
R600 B.n858 B.n857 585
R601 B.n422 B.n421 585
R602 B.n423 B.n422 585
R603 B.n867 B.n866 585
R604 B.n866 B.n865 585
R605 B.n868 B.n420 585
R606 B.n864 B.n420 585
R607 B.n870 B.n869 585
R608 B.n871 B.n870 585
R609 B.n415 B.n414 585
R610 B.n416 B.n415 585
R611 B.n879 B.n878 585
R612 B.n878 B.n877 585
R613 B.n880 B.n413 585
R614 B.n413 B.n412 585
R615 B.n882 B.n881 585
R616 B.n883 B.n882 585
R617 B.n407 B.n406 585
R618 B.n408 B.n407 585
R619 B.n891 B.n890 585
R620 B.n890 B.n889 585
R621 B.n892 B.n405 585
R622 B.n405 B.n403 585
R623 B.n894 B.n893 585
R624 B.n895 B.n894 585
R625 B.n399 B.n398 585
R626 B.n404 B.n399 585
R627 B.n904 B.n903 585
R628 B.n903 B.n902 585
R629 B.n905 B.n397 585
R630 B.n397 B.n396 585
R631 B.n907 B.n906 585
R632 B.n908 B.n907 585
R633 B.n2 B.n0 585
R634 B.n4 B.n2 585
R635 B.n3 B.n1 585
R636 B.n1044 B.n3 585
R637 B.n1042 B.n1041 585
R638 B.n1043 B.n1042 585
R639 B.n1040 B.n9 585
R640 B.n9 B.n8 585
R641 B.n1039 B.n1038 585
R642 B.n1038 B.n1037 585
R643 B.n11 B.n10 585
R644 B.n1036 B.n11 585
R645 B.n1034 B.n1033 585
R646 B.n1035 B.n1034 585
R647 B.n1032 B.n16 585
R648 B.n16 B.n15 585
R649 B.n1031 B.n1030 585
R650 B.n1030 B.n1029 585
R651 B.n18 B.n17 585
R652 B.n1028 B.n18 585
R653 B.n1026 B.n1025 585
R654 B.n1027 B.n1026 585
R655 B.n1024 B.n23 585
R656 B.n23 B.n22 585
R657 B.n1023 B.n1022 585
R658 B.n1022 B.n1021 585
R659 B.n25 B.n24 585
R660 B.n1020 B.n25 585
R661 B.n1018 B.n1017 585
R662 B.n1019 B.n1018 585
R663 B.n1016 B.n29 585
R664 B.n32 B.n29 585
R665 B.n1015 B.n1014 585
R666 B.n1014 B.n1013 585
R667 B.n31 B.n30 585
R668 B.n1012 B.n31 585
R669 B.n1010 B.n1009 585
R670 B.n1011 B.n1010 585
R671 B.n1008 B.n37 585
R672 B.n37 B.n36 585
R673 B.n1007 B.n1006 585
R674 B.n1006 B.n1005 585
R675 B.n39 B.n38 585
R676 B.n1004 B.n39 585
R677 B.n1002 B.n1001 585
R678 B.n1003 B.n1002 585
R679 B.n1000 B.n44 585
R680 B.n44 B.n43 585
R681 B.n999 B.n998 585
R682 B.n998 B.n997 585
R683 B.n46 B.n45 585
R684 B.n996 B.n46 585
R685 B.n994 B.n993 585
R686 B.n995 B.n994 585
R687 B.n992 B.n51 585
R688 B.n51 B.n50 585
R689 B.n991 B.n990 585
R690 B.n990 B.n989 585
R691 B.n53 B.n52 585
R692 B.n988 B.n53 585
R693 B.n986 B.n985 585
R694 B.n987 B.n986 585
R695 B.n984 B.n58 585
R696 B.n58 B.n57 585
R697 B.n983 B.n982 585
R698 B.n982 B.n981 585
R699 B.n60 B.n59 585
R700 B.n980 B.n60 585
R701 B.n978 B.n977 585
R702 B.n979 B.n978 585
R703 B.n976 B.n65 585
R704 B.n65 B.n64 585
R705 B.n975 B.n974 585
R706 B.n974 B.n973 585
R707 B.n67 B.n66 585
R708 B.n972 B.n67 585
R709 B.n970 B.n969 585
R710 B.n971 B.n970 585
R711 B.n968 B.n72 585
R712 B.n72 B.n71 585
R713 B.n1047 B.n1046 585
R714 B.n1046 B.n1045 585
R715 B.n538 B.t21 510.283
R716 B.n535 B.t10 510.283
R717 B.n141 B.t14 510.283
R718 B.n139 B.t18 510.283
R719 B.n793 B.n468 497.305
R720 B.n966 B.n72 497.305
R721 B.n533 B.n466 497.305
R722 B.n962 B.n138 497.305
R723 B.n964 B.n963 256.663
R724 B.n964 B.n136 256.663
R725 B.n964 B.n135 256.663
R726 B.n964 B.n134 256.663
R727 B.n964 B.n133 256.663
R728 B.n964 B.n132 256.663
R729 B.n964 B.n131 256.663
R730 B.n964 B.n130 256.663
R731 B.n964 B.n129 256.663
R732 B.n964 B.n128 256.663
R733 B.n964 B.n127 256.663
R734 B.n964 B.n126 256.663
R735 B.n964 B.n125 256.663
R736 B.n964 B.n124 256.663
R737 B.n964 B.n123 256.663
R738 B.n964 B.n122 256.663
R739 B.n964 B.n121 256.663
R740 B.n964 B.n120 256.663
R741 B.n964 B.n119 256.663
R742 B.n964 B.n118 256.663
R743 B.n964 B.n117 256.663
R744 B.n964 B.n116 256.663
R745 B.n964 B.n115 256.663
R746 B.n964 B.n114 256.663
R747 B.n964 B.n113 256.663
R748 B.n964 B.n112 256.663
R749 B.n964 B.n111 256.663
R750 B.n964 B.n110 256.663
R751 B.n964 B.n109 256.663
R752 B.n964 B.n108 256.663
R753 B.n964 B.n107 256.663
R754 B.n964 B.n106 256.663
R755 B.n964 B.n105 256.663
R756 B.n964 B.n104 256.663
R757 B.n964 B.n103 256.663
R758 B.n964 B.n102 256.663
R759 B.n964 B.n101 256.663
R760 B.n964 B.n100 256.663
R761 B.n964 B.n99 256.663
R762 B.n964 B.n98 256.663
R763 B.n964 B.n97 256.663
R764 B.n964 B.n96 256.663
R765 B.n964 B.n95 256.663
R766 B.n964 B.n94 256.663
R767 B.n964 B.n93 256.663
R768 B.n964 B.n92 256.663
R769 B.n964 B.n91 256.663
R770 B.n964 B.n90 256.663
R771 B.n964 B.n89 256.663
R772 B.n964 B.n88 256.663
R773 B.n964 B.n87 256.663
R774 B.n964 B.n86 256.663
R775 B.n964 B.n85 256.663
R776 B.n964 B.n84 256.663
R777 B.n964 B.n83 256.663
R778 B.n964 B.n82 256.663
R779 B.n964 B.n81 256.663
R780 B.n964 B.n80 256.663
R781 B.n964 B.n79 256.663
R782 B.n964 B.n78 256.663
R783 B.n964 B.n77 256.663
R784 B.n964 B.n76 256.663
R785 B.n964 B.n75 256.663
R786 B.n965 B.n964 256.663
R787 B.n792 B.n791 256.663
R788 B.n791 B.n471 256.663
R789 B.n791 B.n472 256.663
R790 B.n791 B.n473 256.663
R791 B.n791 B.n474 256.663
R792 B.n791 B.n475 256.663
R793 B.n791 B.n476 256.663
R794 B.n791 B.n477 256.663
R795 B.n791 B.n478 256.663
R796 B.n791 B.n479 256.663
R797 B.n791 B.n480 256.663
R798 B.n791 B.n481 256.663
R799 B.n791 B.n482 256.663
R800 B.n791 B.n483 256.663
R801 B.n791 B.n484 256.663
R802 B.n791 B.n485 256.663
R803 B.n791 B.n486 256.663
R804 B.n791 B.n487 256.663
R805 B.n791 B.n488 256.663
R806 B.n791 B.n489 256.663
R807 B.n791 B.n490 256.663
R808 B.n791 B.n491 256.663
R809 B.n791 B.n492 256.663
R810 B.n791 B.n493 256.663
R811 B.n791 B.n494 256.663
R812 B.n791 B.n495 256.663
R813 B.n791 B.n496 256.663
R814 B.n791 B.n497 256.663
R815 B.n791 B.n498 256.663
R816 B.n791 B.n499 256.663
R817 B.n791 B.n500 256.663
R818 B.n791 B.n501 256.663
R819 B.n791 B.n502 256.663
R820 B.n791 B.n503 256.663
R821 B.n791 B.n504 256.663
R822 B.n791 B.n505 256.663
R823 B.n791 B.n506 256.663
R824 B.n791 B.n507 256.663
R825 B.n791 B.n508 256.663
R826 B.n791 B.n509 256.663
R827 B.n791 B.n510 256.663
R828 B.n791 B.n511 256.663
R829 B.n791 B.n512 256.663
R830 B.n791 B.n513 256.663
R831 B.n791 B.n514 256.663
R832 B.n791 B.n515 256.663
R833 B.n791 B.n516 256.663
R834 B.n791 B.n517 256.663
R835 B.n791 B.n518 256.663
R836 B.n791 B.n519 256.663
R837 B.n791 B.n520 256.663
R838 B.n791 B.n521 256.663
R839 B.n791 B.n522 256.663
R840 B.n791 B.n523 256.663
R841 B.n791 B.n524 256.663
R842 B.n791 B.n525 256.663
R843 B.n791 B.n526 256.663
R844 B.n791 B.n527 256.663
R845 B.n791 B.n528 256.663
R846 B.n791 B.n529 256.663
R847 B.n791 B.n530 256.663
R848 B.n791 B.n531 256.663
R849 B.n791 B.n532 256.663
R850 B.n797 B.n468 163.367
R851 B.n797 B.n462 163.367
R852 B.n805 B.n462 163.367
R853 B.n805 B.n460 163.367
R854 B.n809 B.n460 163.367
R855 B.n809 B.n454 163.367
R856 B.n817 B.n454 163.367
R857 B.n817 B.n452 163.367
R858 B.n821 B.n452 163.367
R859 B.n821 B.n446 163.367
R860 B.n829 B.n446 163.367
R861 B.n829 B.n444 163.367
R862 B.n833 B.n444 163.367
R863 B.n833 B.n438 163.367
R864 B.n841 B.n438 163.367
R865 B.n841 B.n436 163.367
R866 B.n845 B.n436 163.367
R867 B.n845 B.n430 163.367
R868 B.n853 B.n430 163.367
R869 B.n853 B.n428 163.367
R870 B.n857 B.n428 163.367
R871 B.n857 B.n422 163.367
R872 B.n866 B.n422 163.367
R873 B.n866 B.n420 163.367
R874 B.n870 B.n420 163.367
R875 B.n870 B.n415 163.367
R876 B.n878 B.n415 163.367
R877 B.n878 B.n413 163.367
R878 B.n882 B.n413 163.367
R879 B.n882 B.n407 163.367
R880 B.n890 B.n407 163.367
R881 B.n890 B.n405 163.367
R882 B.n894 B.n405 163.367
R883 B.n894 B.n399 163.367
R884 B.n903 B.n399 163.367
R885 B.n903 B.n397 163.367
R886 B.n907 B.n397 163.367
R887 B.n907 B.n2 163.367
R888 B.n1046 B.n2 163.367
R889 B.n1046 B.n3 163.367
R890 B.n1042 B.n3 163.367
R891 B.n1042 B.n9 163.367
R892 B.n1038 B.n9 163.367
R893 B.n1038 B.n11 163.367
R894 B.n1034 B.n11 163.367
R895 B.n1034 B.n16 163.367
R896 B.n1030 B.n16 163.367
R897 B.n1030 B.n18 163.367
R898 B.n1026 B.n18 163.367
R899 B.n1026 B.n23 163.367
R900 B.n1022 B.n23 163.367
R901 B.n1022 B.n25 163.367
R902 B.n1018 B.n25 163.367
R903 B.n1018 B.n29 163.367
R904 B.n1014 B.n29 163.367
R905 B.n1014 B.n31 163.367
R906 B.n1010 B.n31 163.367
R907 B.n1010 B.n37 163.367
R908 B.n1006 B.n37 163.367
R909 B.n1006 B.n39 163.367
R910 B.n1002 B.n39 163.367
R911 B.n1002 B.n44 163.367
R912 B.n998 B.n44 163.367
R913 B.n998 B.n46 163.367
R914 B.n994 B.n46 163.367
R915 B.n994 B.n51 163.367
R916 B.n990 B.n51 163.367
R917 B.n990 B.n53 163.367
R918 B.n986 B.n53 163.367
R919 B.n986 B.n58 163.367
R920 B.n982 B.n58 163.367
R921 B.n982 B.n60 163.367
R922 B.n978 B.n60 163.367
R923 B.n978 B.n65 163.367
R924 B.n974 B.n65 163.367
R925 B.n974 B.n67 163.367
R926 B.n970 B.n67 163.367
R927 B.n970 B.n72 163.367
R928 B.n790 B.n470 163.367
R929 B.n790 B.n534 163.367
R930 B.n786 B.n785 163.367
R931 B.n782 B.n781 163.367
R932 B.n778 B.n777 163.367
R933 B.n774 B.n773 163.367
R934 B.n770 B.n769 163.367
R935 B.n766 B.n765 163.367
R936 B.n762 B.n761 163.367
R937 B.n758 B.n757 163.367
R938 B.n754 B.n753 163.367
R939 B.n750 B.n749 163.367
R940 B.n746 B.n745 163.367
R941 B.n742 B.n741 163.367
R942 B.n738 B.n737 163.367
R943 B.n734 B.n733 163.367
R944 B.n730 B.n729 163.367
R945 B.n726 B.n725 163.367
R946 B.n722 B.n721 163.367
R947 B.n718 B.n717 163.367
R948 B.n714 B.n713 163.367
R949 B.n710 B.n709 163.367
R950 B.n706 B.n705 163.367
R951 B.n702 B.n701 163.367
R952 B.n698 B.n697 163.367
R953 B.n694 B.n693 163.367
R954 B.n690 B.n689 163.367
R955 B.n686 B.n685 163.367
R956 B.n682 B.n681 163.367
R957 B.n678 B.n677 163.367
R958 B.n674 B.n673 163.367
R959 B.n670 B.n669 163.367
R960 B.n666 B.n665 163.367
R961 B.n662 B.n661 163.367
R962 B.n658 B.n657 163.367
R963 B.n654 B.n653 163.367
R964 B.n650 B.n649 163.367
R965 B.n646 B.n645 163.367
R966 B.n642 B.n641 163.367
R967 B.n638 B.n637 163.367
R968 B.n634 B.n633 163.367
R969 B.n630 B.n629 163.367
R970 B.n626 B.n625 163.367
R971 B.n622 B.n621 163.367
R972 B.n618 B.n617 163.367
R973 B.n614 B.n613 163.367
R974 B.n610 B.n609 163.367
R975 B.n606 B.n605 163.367
R976 B.n602 B.n601 163.367
R977 B.n598 B.n597 163.367
R978 B.n594 B.n593 163.367
R979 B.n590 B.n589 163.367
R980 B.n586 B.n585 163.367
R981 B.n582 B.n581 163.367
R982 B.n578 B.n577 163.367
R983 B.n574 B.n573 163.367
R984 B.n570 B.n569 163.367
R985 B.n566 B.n565 163.367
R986 B.n562 B.n561 163.367
R987 B.n558 B.n557 163.367
R988 B.n554 B.n553 163.367
R989 B.n550 B.n549 163.367
R990 B.n546 B.n545 163.367
R991 B.n542 B.n533 163.367
R992 B.n799 B.n466 163.367
R993 B.n799 B.n464 163.367
R994 B.n803 B.n464 163.367
R995 B.n803 B.n458 163.367
R996 B.n811 B.n458 163.367
R997 B.n811 B.n456 163.367
R998 B.n815 B.n456 163.367
R999 B.n815 B.n450 163.367
R1000 B.n823 B.n450 163.367
R1001 B.n823 B.n448 163.367
R1002 B.n827 B.n448 163.367
R1003 B.n827 B.n441 163.367
R1004 B.n835 B.n441 163.367
R1005 B.n835 B.n439 163.367
R1006 B.n839 B.n439 163.367
R1007 B.n839 B.n434 163.367
R1008 B.n847 B.n434 163.367
R1009 B.n847 B.n432 163.367
R1010 B.n851 B.n432 163.367
R1011 B.n851 B.n426 163.367
R1012 B.n859 B.n426 163.367
R1013 B.n859 B.n424 163.367
R1014 B.n863 B.n424 163.367
R1015 B.n863 B.n419 163.367
R1016 B.n872 B.n419 163.367
R1017 B.n872 B.n417 163.367
R1018 B.n876 B.n417 163.367
R1019 B.n876 B.n411 163.367
R1020 B.n884 B.n411 163.367
R1021 B.n884 B.n409 163.367
R1022 B.n888 B.n409 163.367
R1023 B.n888 B.n402 163.367
R1024 B.n896 B.n402 163.367
R1025 B.n896 B.n400 163.367
R1026 B.n901 B.n400 163.367
R1027 B.n901 B.n395 163.367
R1028 B.n909 B.n395 163.367
R1029 B.n910 B.n909 163.367
R1030 B.n910 B.n5 163.367
R1031 B.n6 B.n5 163.367
R1032 B.n7 B.n6 163.367
R1033 B.n915 B.n7 163.367
R1034 B.n915 B.n12 163.367
R1035 B.n13 B.n12 163.367
R1036 B.n14 B.n13 163.367
R1037 B.n920 B.n14 163.367
R1038 B.n920 B.n19 163.367
R1039 B.n20 B.n19 163.367
R1040 B.n21 B.n20 163.367
R1041 B.n925 B.n21 163.367
R1042 B.n925 B.n26 163.367
R1043 B.n27 B.n26 163.367
R1044 B.n28 B.n27 163.367
R1045 B.n930 B.n28 163.367
R1046 B.n930 B.n33 163.367
R1047 B.n34 B.n33 163.367
R1048 B.n35 B.n34 163.367
R1049 B.n935 B.n35 163.367
R1050 B.n935 B.n40 163.367
R1051 B.n41 B.n40 163.367
R1052 B.n42 B.n41 163.367
R1053 B.n940 B.n42 163.367
R1054 B.n940 B.n47 163.367
R1055 B.n48 B.n47 163.367
R1056 B.n49 B.n48 163.367
R1057 B.n945 B.n49 163.367
R1058 B.n945 B.n54 163.367
R1059 B.n55 B.n54 163.367
R1060 B.n56 B.n55 163.367
R1061 B.n950 B.n56 163.367
R1062 B.n950 B.n61 163.367
R1063 B.n62 B.n61 163.367
R1064 B.n63 B.n62 163.367
R1065 B.n955 B.n63 163.367
R1066 B.n955 B.n68 163.367
R1067 B.n69 B.n68 163.367
R1068 B.n70 B.n69 163.367
R1069 B.n138 B.n70 163.367
R1070 B.n143 B.n74 163.367
R1071 B.n147 B.n146 163.367
R1072 B.n151 B.n150 163.367
R1073 B.n155 B.n154 163.367
R1074 B.n159 B.n158 163.367
R1075 B.n163 B.n162 163.367
R1076 B.n167 B.n166 163.367
R1077 B.n171 B.n170 163.367
R1078 B.n175 B.n174 163.367
R1079 B.n179 B.n178 163.367
R1080 B.n183 B.n182 163.367
R1081 B.n187 B.n186 163.367
R1082 B.n191 B.n190 163.367
R1083 B.n195 B.n194 163.367
R1084 B.n199 B.n198 163.367
R1085 B.n203 B.n202 163.367
R1086 B.n207 B.n206 163.367
R1087 B.n211 B.n210 163.367
R1088 B.n215 B.n214 163.367
R1089 B.n219 B.n218 163.367
R1090 B.n223 B.n222 163.367
R1091 B.n227 B.n226 163.367
R1092 B.n231 B.n230 163.367
R1093 B.n235 B.n234 163.367
R1094 B.n239 B.n238 163.367
R1095 B.n243 B.n242 163.367
R1096 B.n247 B.n246 163.367
R1097 B.n251 B.n250 163.367
R1098 B.n255 B.n254 163.367
R1099 B.n260 B.n259 163.367
R1100 B.n264 B.n263 163.367
R1101 B.n268 B.n267 163.367
R1102 B.n272 B.n271 163.367
R1103 B.n276 B.n275 163.367
R1104 B.n281 B.n280 163.367
R1105 B.n285 B.n284 163.367
R1106 B.n289 B.n288 163.367
R1107 B.n293 B.n292 163.367
R1108 B.n297 B.n296 163.367
R1109 B.n301 B.n300 163.367
R1110 B.n305 B.n304 163.367
R1111 B.n309 B.n308 163.367
R1112 B.n313 B.n312 163.367
R1113 B.n317 B.n316 163.367
R1114 B.n321 B.n320 163.367
R1115 B.n325 B.n324 163.367
R1116 B.n329 B.n328 163.367
R1117 B.n333 B.n332 163.367
R1118 B.n337 B.n336 163.367
R1119 B.n341 B.n340 163.367
R1120 B.n345 B.n344 163.367
R1121 B.n349 B.n348 163.367
R1122 B.n353 B.n352 163.367
R1123 B.n357 B.n356 163.367
R1124 B.n361 B.n360 163.367
R1125 B.n365 B.n364 163.367
R1126 B.n369 B.n368 163.367
R1127 B.n373 B.n372 163.367
R1128 B.n377 B.n376 163.367
R1129 B.n381 B.n380 163.367
R1130 B.n385 B.n384 163.367
R1131 B.n389 B.n388 163.367
R1132 B.n391 B.n137 163.367
R1133 B.n538 B.t23 107.007
R1134 B.n139 B.t19 107.007
R1135 B.n535 B.t13 106.984
R1136 B.n141 B.t16 106.984
R1137 B.n539 B.t22 73.0678
R1138 B.n140 B.t20 73.0678
R1139 B.n536 B.t12 73.0441
R1140 B.n142 B.t17 73.0441
R1141 B.n793 B.n792 71.676
R1142 B.n534 B.n471 71.676
R1143 B.n785 B.n472 71.676
R1144 B.n781 B.n473 71.676
R1145 B.n777 B.n474 71.676
R1146 B.n773 B.n475 71.676
R1147 B.n769 B.n476 71.676
R1148 B.n765 B.n477 71.676
R1149 B.n761 B.n478 71.676
R1150 B.n757 B.n479 71.676
R1151 B.n753 B.n480 71.676
R1152 B.n749 B.n481 71.676
R1153 B.n745 B.n482 71.676
R1154 B.n741 B.n483 71.676
R1155 B.n737 B.n484 71.676
R1156 B.n733 B.n485 71.676
R1157 B.n729 B.n486 71.676
R1158 B.n725 B.n487 71.676
R1159 B.n721 B.n488 71.676
R1160 B.n717 B.n489 71.676
R1161 B.n713 B.n490 71.676
R1162 B.n709 B.n491 71.676
R1163 B.n705 B.n492 71.676
R1164 B.n701 B.n493 71.676
R1165 B.n697 B.n494 71.676
R1166 B.n693 B.n495 71.676
R1167 B.n689 B.n496 71.676
R1168 B.n685 B.n497 71.676
R1169 B.n681 B.n498 71.676
R1170 B.n677 B.n499 71.676
R1171 B.n673 B.n500 71.676
R1172 B.n669 B.n501 71.676
R1173 B.n665 B.n502 71.676
R1174 B.n661 B.n503 71.676
R1175 B.n657 B.n504 71.676
R1176 B.n653 B.n505 71.676
R1177 B.n649 B.n506 71.676
R1178 B.n645 B.n507 71.676
R1179 B.n641 B.n508 71.676
R1180 B.n637 B.n509 71.676
R1181 B.n633 B.n510 71.676
R1182 B.n629 B.n511 71.676
R1183 B.n625 B.n512 71.676
R1184 B.n621 B.n513 71.676
R1185 B.n617 B.n514 71.676
R1186 B.n613 B.n515 71.676
R1187 B.n609 B.n516 71.676
R1188 B.n605 B.n517 71.676
R1189 B.n601 B.n518 71.676
R1190 B.n597 B.n519 71.676
R1191 B.n593 B.n520 71.676
R1192 B.n589 B.n521 71.676
R1193 B.n585 B.n522 71.676
R1194 B.n581 B.n523 71.676
R1195 B.n577 B.n524 71.676
R1196 B.n573 B.n525 71.676
R1197 B.n569 B.n526 71.676
R1198 B.n565 B.n527 71.676
R1199 B.n561 B.n528 71.676
R1200 B.n557 B.n529 71.676
R1201 B.n553 B.n530 71.676
R1202 B.n549 B.n531 71.676
R1203 B.n545 B.n532 71.676
R1204 B.n966 B.n965 71.676
R1205 B.n143 B.n75 71.676
R1206 B.n147 B.n76 71.676
R1207 B.n151 B.n77 71.676
R1208 B.n155 B.n78 71.676
R1209 B.n159 B.n79 71.676
R1210 B.n163 B.n80 71.676
R1211 B.n167 B.n81 71.676
R1212 B.n171 B.n82 71.676
R1213 B.n175 B.n83 71.676
R1214 B.n179 B.n84 71.676
R1215 B.n183 B.n85 71.676
R1216 B.n187 B.n86 71.676
R1217 B.n191 B.n87 71.676
R1218 B.n195 B.n88 71.676
R1219 B.n199 B.n89 71.676
R1220 B.n203 B.n90 71.676
R1221 B.n207 B.n91 71.676
R1222 B.n211 B.n92 71.676
R1223 B.n215 B.n93 71.676
R1224 B.n219 B.n94 71.676
R1225 B.n223 B.n95 71.676
R1226 B.n227 B.n96 71.676
R1227 B.n231 B.n97 71.676
R1228 B.n235 B.n98 71.676
R1229 B.n239 B.n99 71.676
R1230 B.n243 B.n100 71.676
R1231 B.n247 B.n101 71.676
R1232 B.n251 B.n102 71.676
R1233 B.n255 B.n103 71.676
R1234 B.n260 B.n104 71.676
R1235 B.n264 B.n105 71.676
R1236 B.n268 B.n106 71.676
R1237 B.n272 B.n107 71.676
R1238 B.n276 B.n108 71.676
R1239 B.n281 B.n109 71.676
R1240 B.n285 B.n110 71.676
R1241 B.n289 B.n111 71.676
R1242 B.n293 B.n112 71.676
R1243 B.n297 B.n113 71.676
R1244 B.n301 B.n114 71.676
R1245 B.n305 B.n115 71.676
R1246 B.n309 B.n116 71.676
R1247 B.n313 B.n117 71.676
R1248 B.n317 B.n118 71.676
R1249 B.n321 B.n119 71.676
R1250 B.n325 B.n120 71.676
R1251 B.n329 B.n121 71.676
R1252 B.n333 B.n122 71.676
R1253 B.n337 B.n123 71.676
R1254 B.n341 B.n124 71.676
R1255 B.n345 B.n125 71.676
R1256 B.n349 B.n126 71.676
R1257 B.n353 B.n127 71.676
R1258 B.n357 B.n128 71.676
R1259 B.n361 B.n129 71.676
R1260 B.n365 B.n130 71.676
R1261 B.n369 B.n131 71.676
R1262 B.n373 B.n132 71.676
R1263 B.n377 B.n133 71.676
R1264 B.n381 B.n134 71.676
R1265 B.n385 B.n135 71.676
R1266 B.n389 B.n136 71.676
R1267 B.n963 B.n137 71.676
R1268 B.n963 B.n962 71.676
R1269 B.n391 B.n136 71.676
R1270 B.n388 B.n135 71.676
R1271 B.n384 B.n134 71.676
R1272 B.n380 B.n133 71.676
R1273 B.n376 B.n132 71.676
R1274 B.n372 B.n131 71.676
R1275 B.n368 B.n130 71.676
R1276 B.n364 B.n129 71.676
R1277 B.n360 B.n128 71.676
R1278 B.n356 B.n127 71.676
R1279 B.n352 B.n126 71.676
R1280 B.n348 B.n125 71.676
R1281 B.n344 B.n124 71.676
R1282 B.n340 B.n123 71.676
R1283 B.n336 B.n122 71.676
R1284 B.n332 B.n121 71.676
R1285 B.n328 B.n120 71.676
R1286 B.n324 B.n119 71.676
R1287 B.n320 B.n118 71.676
R1288 B.n316 B.n117 71.676
R1289 B.n312 B.n116 71.676
R1290 B.n308 B.n115 71.676
R1291 B.n304 B.n114 71.676
R1292 B.n300 B.n113 71.676
R1293 B.n296 B.n112 71.676
R1294 B.n292 B.n111 71.676
R1295 B.n288 B.n110 71.676
R1296 B.n284 B.n109 71.676
R1297 B.n280 B.n108 71.676
R1298 B.n275 B.n107 71.676
R1299 B.n271 B.n106 71.676
R1300 B.n267 B.n105 71.676
R1301 B.n263 B.n104 71.676
R1302 B.n259 B.n103 71.676
R1303 B.n254 B.n102 71.676
R1304 B.n250 B.n101 71.676
R1305 B.n246 B.n100 71.676
R1306 B.n242 B.n99 71.676
R1307 B.n238 B.n98 71.676
R1308 B.n234 B.n97 71.676
R1309 B.n230 B.n96 71.676
R1310 B.n226 B.n95 71.676
R1311 B.n222 B.n94 71.676
R1312 B.n218 B.n93 71.676
R1313 B.n214 B.n92 71.676
R1314 B.n210 B.n91 71.676
R1315 B.n206 B.n90 71.676
R1316 B.n202 B.n89 71.676
R1317 B.n198 B.n88 71.676
R1318 B.n194 B.n87 71.676
R1319 B.n190 B.n86 71.676
R1320 B.n186 B.n85 71.676
R1321 B.n182 B.n84 71.676
R1322 B.n178 B.n83 71.676
R1323 B.n174 B.n82 71.676
R1324 B.n170 B.n81 71.676
R1325 B.n166 B.n80 71.676
R1326 B.n162 B.n79 71.676
R1327 B.n158 B.n78 71.676
R1328 B.n154 B.n77 71.676
R1329 B.n150 B.n76 71.676
R1330 B.n146 B.n75 71.676
R1331 B.n965 B.n74 71.676
R1332 B.n792 B.n470 71.676
R1333 B.n786 B.n471 71.676
R1334 B.n782 B.n472 71.676
R1335 B.n778 B.n473 71.676
R1336 B.n774 B.n474 71.676
R1337 B.n770 B.n475 71.676
R1338 B.n766 B.n476 71.676
R1339 B.n762 B.n477 71.676
R1340 B.n758 B.n478 71.676
R1341 B.n754 B.n479 71.676
R1342 B.n750 B.n480 71.676
R1343 B.n746 B.n481 71.676
R1344 B.n742 B.n482 71.676
R1345 B.n738 B.n483 71.676
R1346 B.n734 B.n484 71.676
R1347 B.n730 B.n485 71.676
R1348 B.n726 B.n486 71.676
R1349 B.n722 B.n487 71.676
R1350 B.n718 B.n488 71.676
R1351 B.n714 B.n489 71.676
R1352 B.n710 B.n490 71.676
R1353 B.n706 B.n491 71.676
R1354 B.n702 B.n492 71.676
R1355 B.n698 B.n493 71.676
R1356 B.n694 B.n494 71.676
R1357 B.n690 B.n495 71.676
R1358 B.n686 B.n496 71.676
R1359 B.n682 B.n497 71.676
R1360 B.n678 B.n498 71.676
R1361 B.n674 B.n499 71.676
R1362 B.n670 B.n500 71.676
R1363 B.n666 B.n501 71.676
R1364 B.n662 B.n502 71.676
R1365 B.n658 B.n503 71.676
R1366 B.n654 B.n504 71.676
R1367 B.n650 B.n505 71.676
R1368 B.n646 B.n506 71.676
R1369 B.n642 B.n507 71.676
R1370 B.n638 B.n508 71.676
R1371 B.n634 B.n509 71.676
R1372 B.n630 B.n510 71.676
R1373 B.n626 B.n511 71.676
R1374 B.n622 B.n512 71.676
R1375 B.n618 B.n513 71.676
R1376 B.n614 B.n514 71.676
R1377 B.n610 B.n515 71.676
R1378 B.n606 B.n516 71.676
R1379 B.n602 B.n517 71.676
R1380 B.n598 B.n518 71.676
R1381 B.n594 B.n519 71.676
R1382 B.n590 B.n520 71.676
R1383 B.n586 B.n521 71.676
R1384 B.n582 B.n522 71.676
R1385 B.n578 B.n523 71.676
R1386 B.n574 B.n524 71.676
R1387 B.n570 B.n525 71.676
R1388 B.n566 B.n526 71.676
R1389 B.n562 B.n527 71.676
R1390 B.n558 B.n528 71.676
R1391 B.n554 B.n529 71.676
R1392 B.n550 B.n530 71.676
R1393 B.n546 B.n531 71.676
R1394 B.n542 B.n532 71.676
R1395 B.n540 B.n539 59.5399
R1396 B.n537 B.n536 59.5399
R1397 B.n257 B.n142 59.5399
R1398 B.n278 B.n140 59.5399
R1399 B.n791 B.n467 58.1815
R1400 B.n964 B.n71 58.1815
R1401 B.n539 B.n538 33.9399
R1402 B.n536 B.n535 33.9399
R1403 B.n142 B.n141 33.9399
R1404 B.n140 B.n139 33.9399
R1405 B.n968 B.n967 32.3127
R1406 B.n961 B.n960 32.3127
R1407 B.n541 B.n465 32.3127
R1408 B.n795 B.n794 32.3127
R1409 B.n798 B.n467 32.1656
R1410 B.n798 B.n463 32.1656
R1411 B.n804 B.n463 32.1656
R1412 B.n804 B.n459 32.1656
R1413 B.n810 B.n459 32.1656
R1414 B.n816 B.n455 32.1656
R1415 B.n816 B.n451 32.1656
R1416 B.n822 B.n451 32.1656
R1417 B.n822 B.n447 32.1656
R1418 B.n828 B.n447 32.1656
R1419 B.n828 B.n442 32.1656
R1420 B.n834 B.n442 32.1656
R1421 B.n834 B.n443 32.1656
R1422 B.n840 B.n435 32.1656
R1423 B.n846 B.n435 32.1656
R1424 B.n846 B.n431 32.1656
R1425 B.n852 B.n431 32.1656
R1426 B.n858 B.n427 32.1656
R1427 B.n858 B.n423 32.1656
R1428 B.n865 B.n423 32.1656
R1429 B.n865 B.n864 32.1656
R1430 B.n871 B.n416 32.1656
R1431 B.n877 B.n416 32.1656
R1432 B.n877 B.n412 32.1656
R1433 B.n883 B.n412 32.1656
R1434 B.n889 B.n408 32.1656
R1435 B.n889 B.n403 32.1656
R1436 B.n895 B.n403 32.1656
R1437 B.n895 B.n404 32.1656
R1438 B.n902 B.n396 32.1656
R1439 B.n908 B.n396 32.1656
R1440 B.n908 B.n4 32.1656
R1441 B.n1045 B.n4 32.1656
R1442 B.n1045 B.n1044 32.1656
R1443 B.n1044 B.n1043 32.1656
R1444 B.n1043 B.n8 32.1656
R1445 B.n1037 B.n8 32.1656
R1446 B.n1036 B.n1035 32.1656
R1447 B.n1035 B.n15 32.1656
R1448 B.n1029 B.n15 32.1656
R1449 B.n1029 B.n1028 32.1656
R1450 B.n1027 B.n22 32.1656
R1451 B.n1021 B.n22 32.1656
R1452 B.n1021 B.n1020 32.1656
R1453 B.n1020 B.n1019 32.1656
R1454 B.n1013 B.n32 32.1656
R1455 B.n1013 B.n1012 32.1656
R1456 B.n1012 B.n1011 32.1656
R1457 B.n1011 B.n36 32.1656
R1458 B.n1005 B.n1004 32.1656
R1459 B.n1004 B.n1003 32.1656
R1460 B.n1003 B.n43 32.1656
R1461 B.n997 B.n43 32.1656
R1462 B.n996 B.n995 32.1656
R1463 B.n995 B.n50 32.1656
R1464 B.n989 B.n50 32.1656
R1465 B.n989 B.n988 32.1656
R1466 B.n988 B.n987 32.1656
R1467 B.n987 B.n57 32.1656
R1468 B.n981 B.n57 32.1656
R1469 B.n981 B.n980 32.1656
R1470 B.n979 B.n64 32.1656
R1471 B.n973 B.n64 32.1656
R1472 B.n973 B.n972 32.1656
R1473 B.n972 B.n971 32.1656
R1474 B.n971 B.n71 32.1656
R1475 B.n810 B.t11 28.3815
R1476 B.t15 B.n979 28.3815
R1477 B.n404 B.t1 26.4894
R1478 B.t5 B.n1036 26.4894
R1479 B.n840 B.t9 24.5974
R1480 B.n997 B.t4 24.5974
R1481 B.n883 B.t8 21.7593
R1482 B.t3 B.n1027 21.7593
R1483 B.t2 B.n427 19.8672
R1484 B.t6 B.n36 19.8672
R1485 B B.n1047 18.0485
R1486 B.n864 B.t7 17.0291
R1487 B.n32 B.t0 17.0291
R1488 B.n871 B.t7 15.137
R1489 B.n1019 B.t0 15.137
R1490 B.n852 B.t2 12.2989
R1491 B.n1005 B.t6 12.2989
R1492 B.n967 B.n73 10.6151
R1493 B.n144 B.n73 10.6151
R1494 B.n145 B.n144 10.6151
R1495 B.n148 B.n145 10.6151
R1496 B.n149 B.n148 10.6151
R1497 B.n152 B.n149 10.6151
R1498 B.n153 B.n152 10.6151
R1499 B.n156 B.n153 10.6151
R1500 B.n157 B.n156 10.6151
R1501 B.n160 B.n157 10.6151
R1502 B.n161 B.n160 10.6151
R1503 B.n164 B.n161 10.6151
R1504 B.n165 B.n164 10.6151
R1505 B.n168 B.n165 10.6151
R1506 B.n169 B.n168 10.6151
R1507 B.n172 B.n169 10.6151
R1508 B.n173 B.n172 10.6151
R1509 B.n176 B.n173 10.6151
R1510 B.n177 B.n176 10.6151
R1511 B.n180 B.n177 10.6151
R1512 B.n181 B.n180 10.6151
R1513 B.n184 B.n181 10.6151
R1514 B.n185 B.n184 10.6151
R1515 B.n188 B.n185 10.6151
R1516 B.n189 B.n188 10.6151
R1517 B.n192 B.n189 10.6151
R1518 B.n193 B.n192 10.6151
R1519 B.n196 B.n193 10.6151
R1520 B.n197 B.n196 10.6151
R1521 B.n200 B.n197 10.6151
R1522 B.n201 B.n200 10.6151
R1523 B.n204 B.n201 10.6151
R1524 B.n205 B.n204 10.6151
R1525 B.n208 B.n205 10.6151
R1526 B.n209 B.n208 10.6151
R1527 B.n212 B.n209 10.6151
R1528 B.n213 B.n212 10.6151
R1529 B.n216 B.n213 10.6151
R1530 B.n217 B.n216 10.6151
R1531 B.n220 B.n217 10.6151
R1532 B.n221 B.n220 10.6151
R1533 B.n224 B.n221 10.6151
R1534 B.n225 B.n224 10.6151
R1535 B.n228 B.n225 10.6151
R1536 B.n229 B.n228 10.6151
R1537 B.n232 B.n229 10.6151
R1538 B.n233 B.n232 10.6151
R1539 B.n236 B.n233 10.6151
R1540 B.n237 B.n236 10.6151
R1541 B.n240 B.n237 10.6151
R1542 B.n241 B.n240 10.6151
R1543 B.n244 B.n241 10.6151
R1544 B.n245 B.n244 10.6151
R1545 B.n248 B.n245 10.6151
R1546 B.n249 B.n248 10.6151
R1547 B.n252 B.n249 10.6151
R1548 B.n253 B.n252 10.6151
R1549 B.n256 B.n253 10.6151
R1550 B.n261 B.n258 10.6151
R1551 B.n262 B.n261 10.6151
R1552 B.n265 B.n262 10.6151
R1553 B.n266 B.n265 10.6151
R1554 B.n269 B.n266 10.6151
R1555 B.n270 B.n269 10.6151
R1556 B.n273 B.n270 10.6151
R1557 B.n274 B.n273 10.6151
R1558 B.n277 B.n274 10.6151
R1559 B.n282 B.n279 10.6151
R1560 B.n283 B.n282 10.6151
R1561 B.n286 B.n283 10.6151
R1562 B.n287 B.n286 10.6151
R1563 B.n290 B.n287 10.6151
R1564 B.n291 B.n290 10.6151
R1565 B.n294 B.n291 10.6151
R1566 B.n295 B.n294 10.6151
R1567 B.n298 B.n295 10.6151
R1568 B.n299 B.n298 10.6151
R1569 B.n302 B.n299 10.6151
R1570 B.n303 B.n302 10.6151
R1571 B.n306 B.n303 10.6151
R1572 B.n307 B.n306 10.6151
R1573 B.n310 B.n307 10.6151
R1574 B.n311 B.n310 10.6151
R1575 B.n314 B.n311 10.6151
R1576 B.n315 B.n314 10.6151
R1577 B.n318 B.n315 10.6151
R1578 B.n319 B.n318 10.6151
R1579 B.n322 B.n319 10.6151
R1580 B.n323 B.n322 10.6151
R1581 B.n326 B.n323 10.6151
R1582 B.n327 B.n326 10.6151
R1583 B.n330 B.n327 10.6151
R1584 B.n331 B.n330 10.6151
R1585 B.n334 B.n331 10.6151
R1586 B.n335 B.n334 10.6151
R1587 B.n338 B.n335 10.6151
R1588 B.n339 B.n338 10.6151
R1589 B.n342 B.n339 10.6151
R1590 B.n343 B.n342 10.6151
R1591 B.n346 B.n343 10.6151
R1592 B.n347 B.n346 10.6151
R1593 B.n350 B.n347 10.6151
R1594 B.n351 B.n350 10.6151
R1595 B.n354 B.n351 10.6151
R1596 B.n355 B.n354 10.6151
R1597 B.n358 B.n355 10.6151
R1598 B.n359 B.n358 10.6151
R1599 B.n362 B.n359 10.6151
R1600 B.n363 B.n362 10.6151
R1601 B.n366 B.n363 10.6151
R1602 B.n367 B.n366 10.6151
R1603 B.n370 B.n367 10.6151
R1604 B.n371 B.n370 10.6151
R1605 B.n374 B.n371 10.6151
R1606 B.n375 B.n374 10.6151
R1607 B.n378 B.n375 10.6151
R1608 B.n379 B.n378 10.6151
R1609 B.n382 B.n379 10.6151
R1610 B.n383 B.n382 10.6151
R1611 B.n386 B.n383 10.6151
R1612 B.n387 B.n386 10.6151
R1613 B.n390 B.n387 10.6151
R1614 B.n392 B.n390 10.6151
R1615 B.n393 B.n392 10.6151
R1616 B.n961 B.n393 10.6151
R1617 B.n800 B.n465 10.6151
R1618 B.n801 B.n800 10.6151
R1619 B.n802 B.n801 10.6151
R1620 B.n802 B.n457 10.6151
R1621 B.n812 B.n457 10.6151
R1622 B.n813 B.n812 10.6151
R1623 B.n814 B.n813 10.6151
R1624 B.n814 B.n449 10.6151
R1625 B.n824 B.n449 10.6151
R1626 B.n825 B.n824 10.6151
R1627 B.n826 B.n825 10.6151
R1628 B.n826 B.n440 10.6151
R1629 B.n836 B.n440 10.6151
R1630 B.n837 B.n836 10.6151
R1631 B.n838 B.n837 10.6151
R1632 B.n838 B.n433 10.6151
R1633 B.n848 B.n433 10.6151
R1634 B.n849 B.n848 10.6151
R1635 B.n850 B.n849 10.6151
R1636 B.n850 B.n425 10.6151
R1637 B.n860 B.n425 10.6151
R1638 B.n861 B.n860 10.6151
R1639 B.n862 B.n861 10.6151
R1640 B.n862 B.n418 10.6151
R1641 B.n873 B.n418 10.6151
R1642 B.n874 B.n873 10.6151
R1643 B.n875 B.n874 10.6151
R1644 B.n875 B.n410 10.6151
R1645 B.n885 B.n410 10.6151
R1646 B.n886 B.n885 10.6151
R1647 B.n887 B.n886 10.6151
R1648 B.n887 B.n401 10.6151
R1649 B.n897 B.n401 10.6151
R1650 B.n898 B.n897 10.6151
R1651 B.n900 B.n898 10.6151
R1652 B.n900 B.n899 10.6151
R1653 B.n899 B.n394 10.6151
R1654 B.n911 B.n394 10.6151
R1655 B.n912 B.n911 10.6151
R1656 B.n913 B.n912 10.6151
R1657 B.n914 B.n913 10.6151
R1658 B.n916 B.n914 10.6151
R1659 B.n917 B.n916 10.6151
R1660 B.n918 B.n917 10.6151
R1661 B.n919 B.n918 10.6151
R1662 B.n921 B.n919 10.6151
R1663 B.n922 B.n921 10.6151
R1664 B.n923 B.n922 10.6151
R1665 B.n924 B.n923 10.6151
R1666 B.n926 B.n924 10.6151
R1667 B.n927 B.n926 10.6151
R1668 B.n928 B.n927 10.6151
R1669 B.n929 B.n928 10.6151
R1670 B.n931 B.n929 10.6151
R1671 B.n932 B.n931 10.6151
R1672 B.n933 B.n932 10.6151
R1673 B.n934 B.n933 10.6151
R1674 B.n936 B.n934 10.6151
R1675 B.n937 B.n936 10.6151
R1676 B.n938 B.n937 10.6151
R1677 B.n939 B.n938 10.6151
R1678 B.n941 B.n939 10.6151
R1679 B.n942 B.n941 10.6151
R1680 B.n943 B.n942 10.6151
R1681 B.n944 B.n943 10.6151
R1682 B.n946 B.n944 10.6151
R1683 B.n947 B.n946 10.6151
R1684 B.n948 B.n947 10.6151
R1685 B.n949 B.n948 10.6151
R1686 B.n951 B.n949 10.6151
R1687 B.n952 B.n951 10.6151
R1688 B.n953 B.n952 10.6151
R1689 B.n954 B.n953 10.6151
R1690 B.n956 B.n954 10.6151
R1691 B.n957 B.n956 10.6151
R1692 B.n958 B.n957 10.6151
R1693 B.n959 B.n958 10.6151
R1694 B.n960 B.n959 10.6151
R1695 B.n794 B.n469 10.6151
R1696 B.n789 B.n469 10.6151
R1697 B.n789 B.n788 10.6151
R1698 B.n788 B.n787 10.6151
R1699 B.n787 B.n784 10.6151
R1700 B.n784 B.n783 10.6151
R1701 B.n783 B.n780 10.6151
R1702 B.n780 B.n779 10.6151
R1703 B.n779 B.n776 10.6151
R1704 B.n776 B.n775 10.6151
R1705 B.n775 B.n772 10.6151
R1706 B.n772 B.n771 10.6151
R1707 B.n771 B.n768 10.6151
R1708 B.n768 B.n767 10.6151
R1709 B.n767 B.n764 10.6151
R1710 B.n764 B.n763 10.6151
R1711 B.n763 B.n760 10.6151
R1712 B.n760 B.n759 10.6151
R1713 B.n759 B.n756 10.6151
R1714 B.n756 B.n755 10.6151
R1715 B.n755 B.n752 10.6151
R1716 B.n752 B.n751 10.6151
R1717 B.n751 B.n748 10.6151
R1718 B.n748 B.n747 10.6151
R1719 B.n747 B.n744 10.6151
R1720 B.n744 B.n743 10.6151
R1721 B.n743 B.n740 10.6151
R1722 B.n740 B.n739 10.6151
R1723 B.n739 B.n736 10.6151
R1724 B.n736 B.n735 10.6151
R1725 B.n735 B.n732 10.6151
R1726 B.n732 B.n731 10.6151
R1727 B.n731 B.n728 10.6151
R1728 B.n728 B.n727 10.6151
R1729 B.n727 B.n724 10.6151
R1730 B.n724 B.n723 10.6151
R1731 B.n723 B.n720 10.6151
R1732 B.n720 B.n719 10.6151
R1733 B.n719 B.n716 10.6151
R1734 B.n716 B.n715 10.6151
R1735 B.n715 B.n712 10.6151
R1736 B.n712 B.n711 10.6151
R1737 B.n711 B.n708 10.6151
R1738 B.n708 B.n707 10.6151
R1739 B.n707 B.n704 10.6151
R1740 B.n704 B.n703 10.6151
R1741 B.n703 B.n700 10.6151
R1742 B.n700 B.n699 10.6151
R1743 B.n699 B.n696 10.6151
R1744 B.n696 B.n695 10.6151
R1745 B.n695 B.n692 10.6151
R1746 B.n692 B.n691 10.6151
R1747 B.n691 B.n688 10.6151
R1748 B.n688 B.n687 10.6151
R1749 B.n687 B.n684 10.6151
R1750 B.n684 B.n683 10.6151
R1751 B.n683 B.n680 10.6151
R1752 B.n680 B.n679 10.6151
R1753 B.n676 B.n675 10.6151
R1754 B.n675 B.n672 10.6151
R1755 B.n672 B.n671 10.6151
R1756 B.n671 B.n668 10.6151
R1757 B.n668 B.n667 10.6151
R1758 B.n667 B.n664 10.6151
R1759 B.n664 B.n663 10.6151
R1760 B.n663 B.n660 10.6151
R1761 B.n660 B.n659 10.6151
R1762 B.n656 B.n655 10.6151
R1763 B.n655 B.n652 10.6151
R1764 B.n652 B.n651 10.6151
R1765 B.n651 B.n648 10.6151
R1766 B.n648 B.n647 10.6151
R1767 B.n647 B.n644 10.6151
R1768 B.n644 B.n643 10.6151
R1769 B.n643 B.n640 10.6151
R1770 B.n640 B.n639 10.6151
R1771 B.n639 B.n636 10.6151
R1772 B.n636 B.n635 10.6151
R1773 B.n635 B.n632 10.6151
R1774 B.n632 B.n631 10.6151
R1775 B.n631 B.n628 10.6151
R1776 B.n628 B.n627 10.6151
R1777 B.n627 B.n624 10.6151
R1778 B.n624 B.n623 10.6151
R1779 B.n623 B.n620 10.6151
R1780 B.n620 B.n619 10.6151
R1781 B.n619 B.n616 10.6151
R1782 B.n616 B.n615 10.6151
R1783 B.n615 B.n612 10.6151
R1784 B.n612 B.n611 10.6151
R1785 B.n611 B.n608 10.6151
R1786 B.n608 B.n607 10.6151
R1787 B.n607 B.n604 10.6151
R1788 B.n604 B.n603 10.6151
R1789 B.n603 B.n600 10.6151
R1790 B.n600 B.n599 10.6151
R1791 B.n599 B.n596 10.6151
R1792 B.n596 B.n595 10.6151
R1793 B.n595 B.n592 10.6151
R1794 B.n592 B.n591 10.6151
R1795 B.n591 B.n588 10.6151
R1796 B.n588 B.n587 10.6151
R1797 B.n587 B.n584 10.6151
R1798 B.n584 B.n583 10.6151
R1799 B.n583 B.n580 10.6151
R1800 B.n580 B.n579 10.6151
R1801 B.n579 B.n576 10.6151
R1802 B.n576 B.n575 10.6151
R1803 B.n575 B.n572 10.6151
R1804 B.n572 B.n571 10.6151
R1805 B.n571 B.n568 10.6151
R1806 B.n568 B.n567 10.6151
R1807 B.n567 B.n564 10.6151
R1808 B.n564 B.n563 10.6151
R1809 B.n563 B.n560 10.6151
R1810 B.n560 B.n559 10.6151
R1811 B.n559 B.n556 10.6151
R1812 B.n556 B.n555 10.6151
R1813 B.n555 B.n552 10.6151
R1814 B.n552 B.n551 10.6151
R1815 B.n551 B.n548 10.6151
R1816 B.n548 B.n547 10.6151
R1817 B.n547 B.n544 10.6151
R1818 B.n544 B.n543 10.6151
R1819 B.n543 B.n541 10.6151
R1820 B.n796 B.n795 10.6151
R1821 B.n796 B.n461 10.6151
R1822 B.n806 B.n461 10.6151
R1823 B.n807 B.n806 10.6151
R1824 B.n808 B.n807 10.6151
R1825 B.n808 B.n453 10.6151
R1826 B.n818 B.n453 10.6151
R1827 B.n819 B.n818 10.6151
R1828 B.n820 B.n819 10.6151
R1829 B.n820 B.n445 10.6151
R1830 B.n830 B.n445 10.6151
R1831 B.n831 B.n830 10.6151
R1832 B.n832 B.n831 10.6151
R1833 B.n832 B.n437 10.6151
R1834 B.n842 B.n437 10.6151
R1835 B.n843 B.n842 10.6151
R1836 B.n844 B.n843 10.6151
R1837 B.n844 B.n429 10.6151
R1838 B.n854 B.n429 10.6151
R1839 B.n855 B.n854 10.6151
R1840 B.n856 B.n855 10.6151
R1841 B.n856 B.n421 10.6151
R1842 B.n867 B.n421 10.6151
R1843 B.n868 B.n867 10.6151
R1844 B.n869 B.n868 10.6151
R1845 B.n869 B.n414 10.6151
R1846 B.n879 B.n414 10.6151
R1847 B.n880 B.n879 10.6151
R1848 B.n881 B.n880 10.6151
R1849 B.n881 B.n406 10.6151
R1850 B.n891 B.n406 10.6151
R1851 B.n892 B.n891 10.6151
R1852 B.n893 B.n892 10.6151
R1853 B.n893 B.n398 10.6151
R1854 B.n904 B.n398 10.6151
R1855 B.n905 B.n904 10.6151
R1856 B.n906 B.n905 10.6151
R1857 B.n906 B.n0 10.6151
R1858 B.n1041 B.n1 10.6151
R1859 B.n1041 B.n1040 10.6151
R1860 B.n1040 B.n1039 10.6151
R1861 B.n1039 B.n10 10.6151
R1862 B.n1033 B.n10 10.6151
R1863 B.n1033 B.n1032 10.6151
R1864 B.n1032 B.n1031 10.6151
R1865 B.n1031 B.n17 10.6151
R1866 B.n1025 B.n17 10.6151
R1867 B.n1025 B.n1024 10.6151
R1868 B.n1024 B.n1023 10.6151
R1869 B.n1023 B.n24 10.6151
R1870 B.n1017 B.n24 10.6151
R1871 B.n1017 B.n1016 10.6151
R1872 B.n1016 B.n1015 10.6151
R1873 B.n1015 B.n30 10.6151
R1874 B.n1009 B.n30 10.6151
R1875 B.n1009 B.n1008 10.6151
R1876 B.n1008 B.n1007 10.6151
R1877 B.n1007 B.n38 10.6151
R1878 B.n1001 B.n38 10.6151
R1879 B.n1001 B.n1000 10.6151
R1880 B.n1000 B.n999 10.6151
R1881 B.n999 B.n45 10.6151
R1882 B.n993 B.n45 10.6151
R1883 B.n993 B.n992 10.6151
R1884 B.n992 B.n991 10.6151
R1885 B.n991 B.n52 10.6151
R1886 B.n985 B.n52 10.6151
R1887 B.n985 B.n984 10.6151
R1888 B.n984 B.n983 10.6151
R1889 B.n983 B.n59 10.6151
R1890 B.n977 B.n59 10.6151
R1891 B.n977 B.n976 10.6151
R1892 B.n976 B.n975 10.6151
R1893 B.n975 B.n66 10.6151
R1894 B.n969 B.n66 10.6151
R1895 B.n969 B.n968 10.6151
R1896 B.t8 B.n408 10.4069
R1897 B.n1028 B.t3 10.4069
R1898 B.n257 B.n256 9.36635
R1899 B.n279 B.n278 9.36635
R1900 B.n679 B.n537 9.36635
R1901 B.n656 B.n540 9.36635
R1902 B.n443 B.t9 7.56876
R1903 B.t4 B.n996 7.56876
R1904 B.n902 B.t1 5.6767
R1905 B.n1037 B.t5 5.6767
R1906 B.t11 B.n455 3.78463
R1907 B.n980 B.t15 3.78463
R1908 B.n1047 B.n0 2.81026
R1909 B.n1047 B.n1 2.81026
R1910 B.n258 B.n257 1.24928
R1911 B.n278 B.n277 1.24928
R1912 B.n676 B.n537 1.24928
R1913 B.n659 B.n540 1.24928
R1914 VP.n14 VP.t8 340.659
R1915 VP.n50 VP.t1 305.154
R1916 VP.n5 VP.t4 305.154
R1917 VP.n7 VP.t2 305.154
R1918 VP.n43 VP.t0 305.154
R1919 VP.n56 VP.t9 305.154
R1920 VP.n13 VP.t7 305.154
R1921 VP.n25 VP.t3 305.154
R1922 VP.n31 VP.t5 305.154
R1923 VP.n18 VP.t6 305.154
R1924 VP.n33 VP.n7 173.596
R1925 VP.n57 VP.n56 173.596
R1926 VP.n32 VP.n31 173.596
R1927 VP.n16 VP.n15 161.3
R1928 VP.n17 VP.n12 161.3
R1929 VP.n20 VP.n19 161.3
R1930 VP.n21 VP.n11 161.3
R1931 VP.n23 VP.n22 161.3
R1932 VP.n24 VP.n10 161.3
R1933 VP.n26 VP.n25 161.3
R1934 VP.n27 VP.n9 161.3
R1935 VP.n29 VP.n28 161.3
R1936 VP.n30 VP.n8 161.3
R1937 VP.n55 VP.n0 161.3
R1938 VP.n54 VP.n53 161.3
R1939 VP.n52 VP.n1 161.3
R1940 VP.n51 VP.n50 161.3
R1941 VP.n49 VP.n2 161.3
R1942 VP.n48 VP.n47 161.3
R1943 VP.n46 VP.n3 161.3
R1944 VP.n45 VP.n44 161.3
R1945 VP.n42 VP.n4 161.3
R1946 VP.n41 VP.n40 161.3
R1947 VP.n39 VP.n5 161.3
R1948 VP.n38 VP.n37 161.3
R1949 VP.n36 VP.n6 161.3
R1950 VP.n35 VP.n34 161.3
R1951 VP.n37 VP.n36 52.6866
R1952 VP.n42 VP.n41 52.6866
R1953 VP.n49 VP.n48 52.6866
R1954 VP.n54 VP.n1 52.6866
R1955 VP.n29 VP.n9 52.6866
R1956 VP.n24 VP.n23 52.6866
R1957 VP.n17 VP.n16 52.6866
R1958 VP.n33 VP.n32 51.171
R1959 VP.n14 VP.n13 41.915
R1960 VP.n36 VP.n35 28.4674
R1961 VP.n44 VP.n42 28.4674
R1962 VP.n48 VP.n3 28.4674
R1963 VP.n55 VP.n54 28.4674
R1964 VP.n30 VP.n29 28.4674
R1965 VP.n23 VP.n11 28.4674
R1966 VP.n19 VP.n17 28.4674
R1967 VP.n37 VP.n5 24.5923
R1968 VP.n41 VP.n5 24.5923
R1969 VP.n50 VP.n49 24.5923
R1970 VP.n50 VP.n1 24.5923
R1971 VP.n25 VP.n24 24.5923
R1972 VP.n25 VP.n9 24.5923
R1973 VP.n16 VP.n13 24.5923
R1974 VP.n15 VP.n14 17.507
R1975 VP.n35 VP.n7 12.2964
R1976 VP.n44 VP.n43 12.2964
R1977 VP.n43 VP.n3 12.2964
R1978 VP.n56 VP.n55 12.2964
R1979 VP.n31 VP.n30 12.2964
R1980 VP.n19 VP.n18 12.2964
R1981 VP.n18 VP.n11 12.2964
R1982 VP.n15 VP.n12 0.189894
R1983 VP.n20 VP.n12 0.189894
R1984 VP.n21 VP.n20 0.189894
R1985 VP.n22 VP.n21 0.189894
R1986 VP.n22 VP.n10 0.189894
R1987 VP.n26 VP.n10 0.189894
R1988 VP.n27 VP.n26 0.189894
R1989 VP.n28 VP.n27 0.189894
R1990 VP.n28 VP.n8 0.189894
R1991 VP.n32 VP.n8 0.189894
R1992 VP.n34 VP.n33 0.189894
R1993 VP.n34 VP.n6 0.189894
R1994 VP.n38 VP.n6 0.189894
R1995 VP.n39 VP.n38 0.189894
R1996 VP.n40 VP.n39 0.189894
R1997 VP.n40 VP.n4 0.189894
R1998 VP.n45 VP.n4 0.189894
R1999 VP.n46 VP.n45 0.189894
R2000 VP.n47 VP.n46 0.189894
R2001 VP.n47 VP.n2 0.189894
R2002 VP.n51 VP.n2 0.189894
R2003 VP.n52 VP.n51 0.189894
R2004 VP.n53 VP.n52 0.189894
R2005 VP.n53 VP.n0 0.189894
R2006 VP.n57 VP.n0 0.189894
R2007 VP VP.n57 0.0516364
R2008 VDD1.n1 VDD1.t1 65.2132
R2009 VDD1.n3 VDD1.t7 65.213
R2010 VDD1.n5 VDD1.n4 63.6793
R2011 VDD1.n1 VDD1.n0 62.6034
R2012 VDD1.n7 VDD1.n6 62.6032
R2013 VDD1.n3 VDD1.n2 62.6032
R2014 VDD1.n7 VDD1.n5 47.7186
R2015 VDD1.n6 VDD1.t6 1.10172
R2016 VDD1.n6 VDD1.t4 1.10172
R2017 VDD1.n0 VDD1.t2 1.10172
R2018 VDD1.n0 VDD1.t3 1.10172
R2019 VDD1.n4 VDD1.t8 1.10172
R2020 VDD1.n4 VDD1.t0 1.10172
R2021 VDD1.n2 VDD1.t5 1.10172
R2022 VDD1.n2 VDD1.t9 1.10172
R2023 VDD1 VDD1.n7 1.07378
R2024 VDD1 VDD1.n1 0.435845
R2025 VDD1.n5 VDD1.n3 0.322309
C0 VDD1 VTAIL 14.886599f
C1 VN VTAIL 13.298201f
C2 VP VDD2 0.434189f
C3 VDD2 VDD1 1.40835f
C4 VN VDD2 13.3864f
C5 VP VDD1 13.6639f
C6 VDD2 VTAIL 14.9255f
C7 VN VP 7.76101f
C8 VN VDD1 0.150975f
C9 VP VTAIL 13.312799f
C10 VDD2 B 6.890961f
C11 VDD1 B 6.860606f
C12 VTAIL B 9.511141f
C13 VN B 13.22253f
C14 VP B 11.365468f
C15 VDD1.t1 B 3.75293f
C16 VDD1.t2 B 0.321269f
C17 VDD1.t3 B 0.321269f
C18 VDD1.n0 B 2.92851f
C19 VDD1.n1 B 0.684322f
C20 VDD1.t7 B 3.75293f
C21 VDD1.t5 B 0.321269f
C22 VDD1.t9 B 0.321269f
C23 VDD1.n2 B 2.92851f
C24 VDD1.n3 B 0.677684f
C25 VDD1.t8 B 0.321269f
C26 VDD1.t0 B 0.321269f
C27 VDD1.n4 B 2.93499f
C28 VDD1.n5 B 2.49107f
C29 VDD1.t6 B 0.321269f
C30 VDD1.t4 B 0.321269f
C31 VDD1.n6 B 2.9285f
C32 VDD1.n7 B 2.84048f
C33 VP.n0 B 0.030512f
C34 VP.t9 B 2.14269f
C35 VP.n1 B 0.054198f
C36 VP.n2 B 0.030512f
C37 VP.t1 B 2.14269f
C38 VP.n3 B 0.045809f
C39 VP.n4 B 0.030512f
C40 VP.t4 B 2.14269f
C41 VP.n5 B 0.784303f
C42 VP.n6 B 0.030512f
C43 VP.t2 B 2.14269f
C44 VP.n7 B 0.817052f
C45 VP.n8 B 0.030512f
C46 VP.t5 B 2.14269f
C47 VP.n9 B 0.054198f
C48 VP.n10 B 0.030512f
C49 VP.t3 B 2.14269f
C50 VP.n11 B 0.045809f
C51 VP.n12 B 0.030512f
C52 VP.t7 B 2.14269f
C53 VP.n13 B 0.825108f
C54 VP.t8 B 2.23331f
C55 VP.n14 B 0.820287f
C56 VP.n15 B 0.192321f
C57 VP.n16 B 0.054198f
C58 VP.n17 B 0.031315f
C59 VP.t6 B 2.14269f
C60 VP.n18 B 0.755654f
C61 VP.n19 B 0.045809f
C62 VP.n20 B 0.030512f
C63 VP.n21 B 0.030512f
C64 VP.n22 B 0.030512f
C65 VP.n23 B 0.031315f
C66 VP.n24 B 0.054198f
C67 VP.n25 B 0.784303f
C68 VP.n26 B 0.030512f
C69 VP.n27 B 0.030512f
C70 VP.n28 B 0.030512f
C71 VP.n29 B 0.031315f
C72 VP.n30 B 0.045809f
C73 VP.n31 B 0.817052f
C74 VP.n32 B 1.72188f
C75 VP.n33 B 1.74338f
C76 VP.n34 B 0.030512f
C77 VP.n35 B 0.045809f
C78 VP.n36 B 0.031315f
C79 VP.n37 B 0.054198f
C80 VP.n38 B 0.030512f
C81 VP.n39 B 0.030512f
C82 VP.n40 B 0.030512f
C83 VP.n41 B 0.054198f
C84 VP.n42 B 0.031315f
C85 VP.t0 B 2.14269f
C86 VP.n43 B 0.755654f
C87 VP.n44 B 0.045809f
C88 VP.n45 B 0.030512f
C89 VP.n46 B 0.030512f
C90 VP.n47 B 0.030512f
C91 VP.n48 B 0.031315f
C92 VP.n49 B 0.054198f
C93 VP.n50 B 0.784303f
C94 VP.n51 B 0.030512f
C95 VP.n52 B 0.030512f
C96 VP.n53 B 0.030512f
C97 VP.n54 B 0.031315f
C98 VP.n55 B 0.045809f
C99 VP.n56 B 0.817053f
C100 VP.n57 B 0.028326f
C101 VTAIL.t18 B 0.334491f
C102 VTAIL.t11 B 0.334491f
C103 VTAIL.n0 B 2.98035f
C104 VTAIL.n1 B 0.413395f
C105 VTAIL.t1 B 3.80928f
C106 VTAIL.n2 B 0.520914f
C107 VTAIL.t7 B 0.334491f
C108 VTAIL.t8 B 0.334491f
C109 VTAIL.n3 B 2.98035f
C110 VTAIL.n4 B 0.459171f
C111 VTAIL.t9 B 0.334491f
C112 VTAIL.t2 B 0.334491f
C113 VTAIL.n5 B 2.98035f
C114 VTAIL.n6 B 2.06919f
C115 VTAIL.t15 B 0.334491f
C116 VTAIL.t16 B 0.334491f
C117 VTAIL.n7 B 2.98036f
C118 VTAIL.n8 B 2.06918f
C119 VTAIL.t13 B 0.334491f
C120 VTAIL.t17 B 0.334491f
C121 VTAIL.n9 B 2.98036f
C122 VTAIL.n10 B 0.459167f
C123 VTAIL.t12 B 3.80928f
C124 VTAIL.n11 B 0.52091f
C125 VTAIL.t5 B 0.334491f
C126 VTAIL.t3 B 0.334491f
C127 VTAIL.n12 B 2.98036f
C128 VTAIL.n13 B 0.437587f
C129 VTAIL.t0 B 0.334491f
C130 VTAIL.t6 B 0.334491f
C131 VTAIL.n14 B 2.98036f
C132 VTAIL.n15 B 0.459167f
C133 VTAIL.t4 B 3.80928f
C134 VTAIL.n16 B 2.03807f
C135 VTAIL.t10 B 3.80928f
C136 VTAIL.n17 B 2.03807f
C137 VTAIL.t14 B 0.334491f
C138 VTAIL.t19 B 0.334491f
C139 VTAIL.n18 B 2.98035f
C140 VTAIL.n19 B 0.368927f
C141 VDD2.t0 B 3.72444f
C142 VDD2.t5 B 0.31883f
C143 VDD2.t2 B 0.31883f
C144 VDD2.n0 B 2.90628f
C145 VDD2.n1 B 0.67254f
C146 VDD2.t1 B 0.31883f
C147 VDD2.t4 B 0.31883f
C148 VDD2.n2 B 2.91271f
C149 VDD2.n3 B 2.38517f
C150 VDD2.t3 B 3.71606f
C151 VDD2.n4 B 2.80518f
C152 VDD2.t6 B 0.31883f
C153 VDD2.t9 B 0.31883f
C154 VDD2.n5 B 2.90628f
C155 VDD2.n6 B 0.325096f
C156 VDD2.t7 B 0.31883f
C157 VDD2.t8 B 0.31883f
C158 VDD2.n7 B 2.91268f
C159 VN.n0 B 0.030212f
C160 VN.t9 B 2.12161f
C161 VN.n1 B 0.053665f
C162 VN.n2 B 0.030212f
C163 VN.t0 B 2.12161f
C164 VN.n3 B 0.045358f
C165 VN.n4 B 0.030212f
C166 VN.t8 B 2.12161f
C167 VN.n5 B 0.816988f
C168 VN.t1 B 2.21133f
C169 VN.n6 B 0.812215f
C170 VN.n7 B 0.190428f
C171 VN.n8 B 0.053665f
C172 VN.n9 B 0.031007f
C173 VN.t5 B 2.12161f
C174 VN.n10 B 0.748218f
C175 VN.n11 B 0.045358f
C176 VN.n12 B 0.030212f
C177 VN.n13 B 0.030212f
C178 VN.n14 B 0.030212f
C179 VN.n15 B 0.031007f
C180 VN.n16 B 0.053665f
C181 VN.n17 B 0.776585f
C182 VN.n18 B 0.030212f
C183 VN.n19 B 0.030212f
C184 VN.n20 B 0.030212f
C185 VN.n21 B 0.031007f
C186 VN.n22 B 0.045358f
C187 VN.n23 B 0.809012f
C188 VN.n24 B 0.028047f
C189 VN.n25 B 0.030212f
C190 VN.t4 B 2.12161f
C191 VN.n26 B 0.053665f
C192 VN.n27 B 0.030212f
C193 VN.t3 B 2.12161f
C194 VN.n28 B 0.045358f
C195 VN.n29 B 0.030212f
C196 VN.t6 B 2.12161f
C197 VN.n30 B 0.748218f
C198 VN.t2 B 2.12161f
C199 VN.n31 B 0.816988f
C200 VN.t7 B 2.21133f
C201 VN.n32 B 0.812215f
C202 VN.n33 B 0.190428f
C203 VN.n34 B 0.053665f
C204 VN.n35 B 0.031007f
C205 VN.n36 B 0.045358f
C206 VN.n37 B 0.030212f
C207 VN.n38 B 0.030212f
C208 VN.n39 B 0.030212f
C209 VN.n40 B 0.031007f
C210 VN.n41 B 0.053665f
C211 VN.n42 B 0.776585f
C212 VN.n43 B 0.030212f
C213 VN.n44 B 0.030212f
C214 VN.n45 B 0.030212f
C215 VN.n46 B 0.031007f
C216 VN.n47 B 0.045358f
C217 VN.n48 B 0.809012f
C218 VN.n49 B 1.72456f
.ends

