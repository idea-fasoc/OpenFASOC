* NGSPICE file created from diff_pair_sample_0289.ext - technology: sky130A

.subckt diff_pair_sample_0289 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=4.1769 ps=22.2 w=10.71 l=3.63
X1 VDD1.t6 VP.t1 VTAIL.t15 B.t4 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=4.1769 ps=22.2 w=10.71 l=3.63
X2 VTAIL.t9 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=1.76715 ps=11.04 w=10.71 l=3.63
X3 VTAIL.t3 VN.t0 VDD2.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=4.1769 pd=22.2 as=1.76715 ps=11.04 w=10.71 l=3.63
X4 VDD1.t4 VP.t3 VTAIL.t11 B.t0 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=1.76715 ps=11.04 w=10.71 l=3.63
X5 VDD2.t6 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=1.76715 ps=11.04 w=10.71 l=3.63
X6 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.1769 pd=22.2 as=0 ps=0 w=10.71 l=3.63
X7 VDD2.t5 VN.t2 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=1.76715 ps=11.04 w=10.71 l=3.63
X8 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.1769 pd=22.2 as=0 ps=0 w=10.71 l=3.63
X9 VTAIL.t1 VN.t3 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1769 pd=22.2 as=1.76715 ps=11.04 w=10.71 l=3.63
X10 VTAIL.t10 VP.t4 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=4.1769 pd=22.2 as=1.76715 ps=11.04 w=10.71 l=3.63
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.1769 pd=22.2 as=0 ps=0 w=10.71 l=3.63
X12 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.1769 pd=22.2 as=0 ps=0 w=10.71 l=3.63
X13 VDD2.t3 VN.t4 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=4.1769 ps=22.2 w=10.71 l=3.63
X14 VDD2.t2 VN.t5 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=4.1769 ps=22.2 w=10.71 l=3.63
X15 VDD1.t2 VP.t5 VTAIL.t13 B.t2 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=1.76715 ps=11.04 w=10.71 l=3.63
X16 VTAIL.t5 VN.t6 VDD2.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=1.76715 ps=11.04 w=10.71 l=3.63
X17 VTAIL.t7 VN.t7 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=1.76715 ps=11.04 w=10.71 l=3.63
X18 VTAIL.t12 VP.t6 VDD1.t1 B.t7 sky130_fd_pr__nfet_01v8 ad=1.76715 pd=11.04 as=1.76715 ps=11.04 w=10.71 l=3.63
X19 VTAIL.t8 VP.t7 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.1769 pd=22.2 as=1.76715 ps=11.04 w=10.71 l=3.63
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n36 VP.n35 161.3
R8 VP.n37 VP.n17 161.3
R9 VP.n39 VP.n38 161.3
R10 VP.n40 VP.n16 161.3
R11 VP.n42 VP.n41 161.3
R12 VP.n43 VP.n15 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n14 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n89 VP.n88 161.3
R17 VP.n87 VP.n1 161.3
R18 VP.n86 VP.n85 161.3
R19 VP.n84 VP.n2 161.3
R20 VP.n83 VP.n82 161.3
R21 VP.n81 VP.n3 161.3
R22 VP.n80 VP.n79 161.3
R23 VP.n78 VP.n4 161.3
R24 VP.n77 VP.n76 161.3
R25 VP.n74 VP.n5 161.3
R26 VP.n73 VP.n72 161.3
R27 VP.n71 VP.n6 161.3
R28 VP.n70 VP.n69 161.3
R29 VP.n68 VP.n7 161.3
R30 VP.n67 VP.n66 161.3
R31 VP.n65 VP.n8 161.3
R32 VP.n64 VP.n63 161.3
R33 VP.n61 VP.n9 161.3
R34 VP.n60 VP.n59 161.3
R35 VP.n58 VP.n10 161.3
R36 VP.n57 VP.n56 161.3
R37 VP.n55 VP.n11 161.3
R38 VP.n54 VP.n53 161.3
R39 VP.n52 VP.n12 161.3
R40 VP.n23 VP.t7 104.386
R41 VP.n51 VP.n50 80.7699
R42 VP.n90 VP.n0 80.7699
R43 VP.n49 VP.n13 80.7699
R44 VP.n50 VP.t4 71.1055
R45 VP.n62 VP.t5 71.1055
R46 VP.n75 VP.t6 71.1055
R47 VP.n0 VP.t1 71.1055
R48 VP.n13 VP.t0 71.1055
R49 VP.n34 VP.t2 71.1055
R50 VP.n22 VP.t3 71.1055
R51 VP.n23 VP.n22 63.3269
R52 VP.n56 VP.n10 56.5193
R53 VP.n69 VP.n6 56.5193
R54 VP.n82 VP.n2 56.5193
R55 VP.n41 VP.n15 56.5193
R56 VP.n28 VP.n19 56.5193
R57 VP.n51 VP.n49 54.8478
R58 VP.n54 VP.n12 24.4675
R59 VP.n55 VP.n54 24.4675
R60 VP.n56 VP.n55 24.4675
R61 VP.n60 VP.n10 24.4675
R62 VP.n61 VP.n60 24.4675
R63 VP.n63 VP.n61 24.4675
R64 VP.n67 VP.n8 24.4675
R65 VP.n68 VP.n67 24.4675
R66 VP.n69 VP.n68 24.4675
R67 VP.n73 VP.n6 24.4675
R68 VP.n74 VP.n73 24.4675
R69 VP.n76 VP.n74 24.4675
R70 VP.n80 VP.n4 24.4675
R71 VP.n81 VP.n80 24.4675
R72 VP.n82 VP.n81 24.4675
R73 VP.n86 VP.n2 24.4675
R74 VP.n87 VP.n86 24.4675
R75 VP.n88 VP.n87 24.4675
R76 VP.n45 VP.n15 24.4675
R77 VP.n46 VP.n45 24.4675
R78 VP.n47 VP.n46 24.4675
R79 VP.n32 VP.n19 24.4675
R80 VP.n33 VP.n32 24.4675
R81 VP.n35 VP.n33 24.4675
R82 VP.n39 VP.n17 24.4675
R83 VP.n40 VP.n39 24.4675
R84 VP.n41 VP.n40 24.4675
R85 VP.n26 VP.n21 24.4675
R86 VP.n27 VP.n26 24.4675
R87 VP.n28 VP.n27 24.4675
R88 VP.n63 VP.n62 13.2127
R89 VP.n75 VP.n4 13.2127
R90 VP.n34 VP.n17 13.2127
R91 VP.n62 VP.n8 11.2553
R92 VP.n76 VP.n75 11.2553
R93 VP.n35 VP.n34 11.2553
R94 VP.n22 VP.n21 11.2553
R95 VP.n50 VP.n12 9.29796
R96 VP.n88 VP.n0 9.29796
R97 VP.n47 VP.n13 9.29796
R98 VP.n24 VP.n23 3.17991
R99 VP.n49 VP.n48 0.354971
R100 VP.n52 VP.n51 0.354971
R101 VP.n90 VP.n89 0.354971
R102 VP VP.n90 0.26696
R103 VP.n25 VP.n24 0.189894
R104 VP.n25 VP.n20 0.189894
R105 VP.n29 VP.n20 0.189894
R106 VP.n30 VP.n29 0.189894
R107 VP.n31 VP.n30 0.189894
R108 VP.n31 VP.n18 0.189894
R109 VP.n36 VP.n18 0.189894
R110 VP.n37 VP.n36 0.189894
R111 VP.n38 VP.n37 0.189894
R112 VP.n38 VP.n16 0.189894
R113 VP.n42 VP.n16 0.189894
R114 VP.n43 VP.n42 0.189894
R115 VP.n44 VP.n43 0.189894
R116 VP.n44 VP.n14 0.189894
R117 VP.n48 VP.n14 0.189894
R118 VP.n53 VP.n52 0.189894
R119 VP.n53 VP.n11 0.189894
R120 VP.n57 VP.n11 0.189894
R121 VP.n58 VP.n57 0.189894
R122 VP.n59 VP.n58 0.189894
R123 VP.n59 VP.n9 0.189894
R124 VP.n64 VP.n9 0.189894
R125 VP.n65 VP.n64 0.189894
R126 VP.n66 VP.n65 0.189894
R127 VP.n66 VP.n7 0.189894
R128 VP.n70 VP.n7 0.189894
R129 VP.n71 VP.n70 0.189894
R130 VP.n72 VP.n71 0.189894
R131 VP.n72 VP.n5 0.189894
R132 VP.n77 VP.n5 0.189894
R133 VP.n78 VP.n77 0.189894
R134 VP.n79 VP.n78 0.189894
R135 VP.n79 VP.n3 0.189894
R136 VP.n83 VP.n3 0.189894
R137 VP.n84 VP.n83 0.189894
R138 VP.n85 VP.n84 0.189894
R139 VP.n85 VP.n1 0.189894
R140 VP.n89 VP.n1 0.189894
R141 VTAIL.n466 VTAIL.n414 289.615
R142 VTAIL.n54 VTAIL.n2 289.615
R143 VTAIL.n112 VTAIL.n60 289.615
R144 VTAIL.n172 VTAIL.n120 289.615
R145 VTAIL.n408 VTAIL.n356 289.615
R146 VTAIL.n348 VTAIL.n296 289.615
R147 VTAIL.n290 VTAIL.n238 289.615
R148 VTAIL.n230 VTAIL.n178 289.615
R149 VTAIL.n433 VTAIL.n432 185
R150 VTAIL.n430 VTAIL.n429 185
R151 VTAIL.n439 VTAIL.n438 185
R152 VTAIL.n441 VTAIL.n440 185
R153 VTAIL.n426 VTAIL.n425 185
R154 VTAIL.n447 VTAIL.n446 185
R155 VTAIL.n450 VTAIL.n449 185
R156 VTAIL.n448 VTAIL.n422 185
R157 VTAIL.n455 VTAIL.n421 185
R158 VTAIL.n457 VTAIL.n456 185
R159 VTAIL.n459 VTAIL.n458 185
R160 VTAIL.n418 VTAIL.n417 185
R161 VTAIL.n465 VTAIL.n464 185
R162 VTAIL.n467 VTAIL.n466 185
R163 VTAIL.n21 VTAIL.n20 185
R164 VTAIL.n18 VTAIL.n17 185
R165 VTAIL.n27 VTAIL.n26 185
R166 VTAIL.n29 VTAIL.n28 185
R167 VTAIL.n14 VTAIL.n13 185
R168 VTAIL.n35 VTAIL.n34 185
R169 VTAIL.n38 VTAIL.n37 185
R170 VTAIL.n36 VTAIL.n10 185
R171 VTAIL.n43 VTAIL.n9 185
R172 VTAIL.n45 VTAIL.n44 185
R173 VTAIL.n47 VTAIL.n46 185
R174 VTAIL.n6 VTAIL.n5 185
R175 VTAIL.n53 VTAIL.n52 185
R176 VTAIL.n55 VTAIL.n54 185
R177 VTAIL.n79 VTAIL.n78 185
R178 VTAIL.n76 VTAIL.n75 185
R179 VTAIL.n85 VTAIL.n84 185
R180 VTAIL.n87 VTAIL.n86 185
R181 VTAIL.n72 VTAIL.n71 185
R182 VTAIL.n93 VTAIL.n92 185
R183 VTAIL.n96 VTAIL.n95 185
R184 VTAIL.n94 VTAIL.n68 185
R185 VTAIL.n101 VTAIL.n67 185
R186 VTAIL.n103 VTAIL.n102 185
R187 VTAIL.n105 VTAIL.n104 185
R188 VTAIL.n64 VTAIL.n63 185
R189 VTAIL.n111 VTAIL.n110 185
R190 VTAIL.n113 VTAIL.n112 185
R191 VTAIL.n139 VTAIL.n138 185
R192 VTAIL.n136 VTAIL.n135 185
R193 VTAIL.n145 VTAIL.n144 185
R194 VTAIL.n147 VTAIL.n146 185
R195 VTAIL.n132 VTAIL.n131 185
R196 VTAIL.n153 VTAIL.n152 185
R197 VTAIL.n156 VTAIL.n155 185
R198 VTAIL.n154 VTAIL.n128 185
R199 VTAIL.n161 VTAIL.n127 185
R200 VTAIL.n163 VTAIL.n162 185
R201 VTAIL.n165 VTAIL.n164 185
R202 VTAIL.n124 VTAIL.n123 185
R203 VTAIL.n171 VTAIL.n170 185
R204 VTAIL.n173 VTAIL.n172 185
R205 VTAIL.n409 VTAIL.n408 185
R206 VTAIL.n407 VTAIL.n406 185
R207 VTAIL.n360 VTAIL.n359 185
R208 VTAIL.n401 VTAIL.n400 185
R209 VTAIL.n399 VTAIL.n398 185
R210 VTAIL.n397 VTAIL.n363 185
R211 VTAIL.n367 VTAIL.n364 185
R212 VTAIL.n392 VTAIL.n391 185
R213 VTAIL.n390 VTAIL.n389 185
R214 VTAIL.n369 VTAIL.n368 185
R215 VTAIL.n384 VTAIL.n383 185
R216 VTAIL.n382 VTAIL.n381 185
R217 VTAIL.n373 VTAIL.n372 185
R218 VTAIL.n376 VTAIL.n375 185
R219 VTAIL.n349 VTAIL.n348 185
R220 VTAIL.n347 VTAIL.n346 185
R221 VTAIL.n300 VTAIL.n299 185
R222 VTAIL.n341 VTAIL.n340 185
R223 VTAIL.n339 VTAIL.n338 185
R224 VTAIL.n337 VTAIL.n303 185
R225 VTAIL.n307 VTAIL.n304 185
R226 VTAIL.n332 VTAIL.n331 185
R227 VTAIL.n330 VTAIL.n329 185
R228 VTAIL.n309 VTAIL.n308 185
R229 VTAIL.n324 VTAIL.n323 185
R230 VTAIL.n322 VTAIL.n321 185
R231 VTAIL.n313 VTAIL.n312 185
R232 VTAIL.n316 VTAIL.n315 185
R233 VTAIL.n291 VTAIL.n290 185
R234 VTAIL.n289 VTAIL.n288 185
R235 VTAIL.n242 VTAIL.n241 185
R236 VTAIL.n283 VTAIL.n282 185
R237 VTAIL.n281 VTAIL.n280 185
R238 VTAIL.n279 VTAIL.n245 185
R239 VTAIL.n249 VTAIL.n246 185
R240 VTAIL.n274 VTAIL.n273 185
R241 VTAIL.n272 VTAIL.n271 185
R242 VTAIL.n251 VTAIL.n250 185
R243 VTAIL.n266 VTAIL.n265 185
R244 VTAIL.n264 VTAIL.n263 185
R245 VTAIL.n255 VTAIL.n254 185
R246 VTAIL.n258 VTAIL.n257 185
R247 VTAIL.n231 VTAIL.n230 185
R248 VTAIL.n229 VTAIL.n228 185
R249 VTAIL.n182 VTAIL.n181 185
R250 VTAIL.n223 VTAIL.n222 185
R251 VTAIL.n221 VTAIL.n220 185
R252 VTAIL.n219 VTAIL.n185 185
R253 VTAIL.n189 VTAIL.n186 185
R254 VTAIL.n214 VTAIL.n213 185
R255 VTAIL.n212 VTAIL.n211 185
R256 VTAIL.n191 VTAIL.n190 185
R257 VTAIL.n206 VTAIL.n205 185
R258 VTAIL.n204 VTAIL.n203 185
R259 VTAIL.n195 VTAIL.n194 185
R260 VTAIL.n198 VTAIL.n197 185
R261 VTAIL.t6 VTAIL.n431 149.524
R262 VTAIL.t1 VTAIL.n19 149.524
R263 VTAIL.t15 VTAIL.n77 149.524
R264 VTAIL.t10 VTAIL.n137 149.524
R265 VTAIL.t14 VTAIL.n374 149.524
R266 VTAIL.t8 VTAIL.n314 149.524
R267 VTAIL.t4 VTAIL.n256 149.524
R268 VTAIL.t3 VTAIL.n196 149.524
R269 VTAIL.n432 VTAIL.n429 104.615
R270 VTAIL.n439 VTAIL.n429 104.615
R271 VTAIL.n440 VTAIL.n439 104.615
R272 VTAIL.n440 VTAIL.n425 104.615
R273 VTAIL.n447 VTAIL.n425 104.615
R274 VTAIL.n449 VTAIL.n447 104.615
R275 VTAIL.n449 VTAIL.n448 104.615
R276 VTAIL.n448 VTAIL.n421 104.615
R277 VTAIL.n457 VTAIL.n421 104.615
R278 VTAIL.n458 VTAIL.n457 104.615
R279 VTAIL.n458 VTAIL.n417 104.615
R280 VTAIL.n465 VTAIL.n417 104.615
R281 VTAIL.n466 VTAIL.n465 104.615
R282 VTAIL.n20 VTAIL.n17 104.615
R283 VTAIL.n27 VTAIL.n17 104.615
R284 VTAIL.n28 VTAIL.n27 104.615
R285 VTAIL.n28 VTAIL.n13 104.615
R286 VTAIL.n35 VTAIL.n13 104.615
R287 VTAIL.n37 VTAIL.n35 104.615
R288 VTAIL.n37 VTAIL.n36 104.615
R289 VTAIL.n36 VTAIL.n9 104.615
R290 VTAIL.n45 VTAIL.n9 104.615
R291 VTAIL.n46 VTAIL.n45 104.615
R292 VTAIL.n46 VTAIL.n5 104.615
R293 VTAIL.n53 VTAIL.n5 104.615
R294 VTAIL.n54 VTAIL.n53 104.615
R295 VTAIL.n78 VTAIL.n75 104.615
R296 VTAIL.n85 VTAIL.n75 104.615
R297 VTAIL.n86 VTAIL.n85 104.615
R298 VTAIL.n86 VTAIL.n71 104.615
R299 VTAIL.n93 VTAIL.n71 104.615
R300 VTAIL.n95 VTAIL.n93 104.615
R301 VTAIL.n95 VTAIL.n94 104.615
R302 VTAIL.n94 VTAIL.n67 104.615
R303 VTAIL.n103 VTAIL.n67 104.615
R304 VTAIL.n104 VTAIL.n103 104.615
R305 VTAIL.n104 VTAIL.n63 104.615
R306 VTAIL.n111 VTAIL.n63 104.615
R307 VTAIL.n112 VTAIL.n111 104.615
R308 VTAIL.n138 VTAIL.n135 104.615
R309 VTAIL.n145 VTAIL.n135 104.615
R310 VTAIL.n146 VTAIL.n145 104.615
R311 VTAIL.n146 VTAIL.n131 104.615
R312 VTAIL.n153 VTAIL.n131 104.615
R313 VTAIL.n155 VTAIL.n153 104.615
R314 VTAIL.n155 VTAIL.n154 104.615
R315 VTAIL.n154 VTAIL.n127 104.615
R316 VTAIL.n163 VTAIL.n127 104.615
R317 VTAIL.n164 VTAIL.n163 104.615
R318 VTAIL.n164 VTAIL.n123 104.615
R319 VTAIL.n171 VTAIL.n123 104.615
R320 VTAIL.n172 VTAIL.n171 104.615
R321 VTAIL.n408 VTAIL.n407 104.615
R322 VTAIL.n407 VTAIL.n359 104.615
R323 VTAIL.n400 VTAIL.n359 104.615
R324 VTAIL.n400 VTAIL.n399 104.615
R325 VTAIL.n399 VTAIL.n363 104.615
R326 VTAIL.n367 VTAIL.n363 104.615
R327 VTAIL.n391 VTAIL.n367 104.615
R328 VTAIL.n391 VTAIL.n390 104.615
R329 VTAIL.n390 VTAIL.n368 104.615
R330 VTAIL.n383 VTAIL.n368 104.615
R331 VTAIL.n383 VTAIL.n382 104.615
R332 VTAIL.n382 VTAIL.n372 104.615
R333 VTAIL.n375 VTAIL.n372 104.615
R334 VTAIL.n348 VTAIL.n347 104.615
R335 VTAIL.n347 VTAIL.n299 104.615
R336 VTAIL.n340 VTAIL.n299 104.615
R337 VTAIL.n340 VTAIL.n339 104.615
R338 VTAIL.n339 VTAIL.n303 104.615
R339 VTAIL.n307 VTAIL.n303 104.615
R340 VTAIL.n331 VTAIL.n307 104.615
R341 VTAIL.n331 VTAIL.n330 104.615
R342 VTAIL.n330 VTAIL.n308 104.615
R343 VTAIL.n323 VTAIL.n308 104.615
R344 VTAIL.n323 VTAIL.n322 104.615
R345 VTAIL.n322 VTAIL.n312 104.615
R346 VTAIL.n315 VTAIL.n312 104.615
R347 VTAIL.n290 VTAIL.n289 104.615
R348 VTAIL.n289 VTAIL.n241 104.615
R349 VTAIL.n282 VTAIL.n241 104.615
R350 VTAIL.n282 VTAIL.n281 104.615
R351 VTAIL.n281 VTAIL.n245 104.615
R352 VTAIL.n249 VTAIL.n245 104.615
R353 VTAIL.n273 VTAIL.n249 104.615
R354 VTAIL.n273 VTAIL.n272 104.615
R355 VTAIL.n272 VTAIL.n250 104.615
R356 VTAIL.n265 VTAIL.n250 104.615
R357 VTAIL.n265 VTAIL.n264 104.615
R358 VTAIL.n264 VTAIL.n254 104.615
R359 VTAIL.n257 VTAIL.n254 104.615
R360 VTAIL.n230 VTAIL.n229 104.615
R361 VTAIL.n229 VTAIL.n181 104.615
R362 VTAIL.n222 VTAIL.n181 104.615
R363 VTAIL.n222 VTAIL.n221 104.615
R364 VTAIL.n221 VTAIL.n185 104.615
R365 VTAIL.n189 VTAIL.n185 104.615
R366 VTAIL.n213 VTAIL.n189 104.615
R367 VTAIL.n213 VTAIL.n212 104.615
R368 VTAIL.n212 VTAIL.n190 104.615
R369 VTAIL.n205 VTAIL.n190 104.615
R370 VTAIL.n205 VTAIL.n204 104.615
R371 VTAIL.n204 VTAIL.n194 104.615
R372 VTAIL.n197 VTAIL.n194 104.615
R373 VTAIL.n432 VTAIL.t6 52.3082
R374 VTAIL.n20 VTAIL.t1 52.3082
R375 VTAIL.n78 VTAIL.t15 52.3082
R376 VTAIL.n138 VTAIL.t10 52.3082
R377 VTAIL.n375 VTAIL.t14 52.3082
R378 VTAIL.n315 VTAIL.t8 52.3082
R379 VTAIL.n257 VTAIL.t4 52.3082
R380 VTAIL.n197 VTAIL.t3 52.3082
R381 VTAIL.n355 VTAIL.n354 46.2433
R382 VTAIL.n237 VTAIL.n236 46.2433
R383 VTAIL.n1 VTAIL.n0 46.2431
R384 VTAIL.n119 VTAIL.n118 46.2431
R385 VTAIL.n471 VTAIL.n470 32.7672
R386 VTAIL.n59 VTAIL.n58 32.7672
R387 VTAIL.n117 VTAIL.n116 32.7672
R388 VTAIL.n177 VTAIL.n176 32.7672
R389 VTAIL.n413 VTAIL.n412 32.7672
R390 VTAIL.n353 VTAIL.n352 32.7672
R391 VTAIL.n295 VTAIL.n294 32.7672
R392 VTAIL.n235 VTAIL.n234 32.7672
R393 VTAIL.n471 VTAIL.n413 25.0134
R394 VTAIL.n235 VTAIL.n177 25.0134
R395 VTAIL.n456 VTAIL.n455 13.1884
R396 VTAIL.n44 VTAIL.n43 13.1884
R397 VTAIL.n102 VTAIL.n101 13.1884
R398 VTAIL.n162 VTAIL.n161 13.1884
R399 VTAIL.n398 VTAIL.n397 13.1884
R400 VTAIL.n338 VTAIL.n337 13.1884
R401 VTAIL.n280 VTAIL.n279 13.1884
R402 VTAIL.n220 VTAIL.n219 13.1884
R403 VTAIL.n454 VTAIL.n422 12.8005
R404 VTAIL.n459 VTAIL.n420 12.8005
R405 VTAIL.n42 VTAIL.n10 12.8005
R406 VTAIL.n47 VTAIL.n8 12.8005
R407 VTAIL.n100 VTAIL.n68 12.8005
R408 VTAIL.n105 VTAIL.n66 12.8005
R409 VTAIL.n160 VTAIL.n128 12.8005
R410 VTAIL.n165 VTAIL.n126 12.8005
R411 VTAIL.n401 VTAIL.n362 12.8005
R412 VTAIL.n396 VTAIL.n364 12.8005
R413 VTAIL.n341 VTAIL.n302 12.8005
R414 VTAIL.n336 VTAIL.n304 12.8005
R415 VTAIL.n283 VTAIL.n244 12.8005
R416 VTAIL.n278 VTAIL.n246 12.8005
R417 VTAIL.n223 VTAIL.n184 12.8005
R418 VTAIL.n218 VTAIL.n186 12.8005
R419 VTAIL.n451 VTAIL.n450 12.0247
R420 VTAIL.n460 VTAIL.n418 12.0247
R421 VTAIL.n39 VTAIL.n38 12.0247
R422 VTAIL.n48 VTAIL.n6 12.0247
R423 VTAIL.n97 VTAIL.n96 12.0247
R424 VTAIL.n106 VTAIL.n64 12.0247
R425 VTAIL.n157 VTAIL.n156 12.0247
R426 VTAIL.n166 VTAIL.n124 12.0247
R427 VTAIL.n402 VTAIL.n360 12.0247
R428 VTAIL.n393 VTAIL.n392 12.0247
R429 VTAIL.n342 VTAIL.n300 12.0247
R430 VTAIL.n333 VTAIL.n332 12.0247
R431 VTAIL.n284 VTAIL.n242 12.0247
R432 VTAIL.n275 VTAIL.n274 12.0247
R433 VTAIL.n224 VTAIL.n182 12.0247
R434 VTAIL.n215 VTAIL.n214 12.0247
R435 VTAIL.n446 VTAIL.n424 11.249
R436 VTAIL.n464 VTAIL.n463 11.249
R437 VTAIL.n34 VTAIL.n12 11.249
R438 VTAIL.n52 VTAIL.n51 11.249
R439 VTAIL.n92 VTAIL.n70 11.249
R440 VTAIL.n110 VTAIL.n109 11.249
R441 VTAIL.n152 VTAIL.n130 11.249
R442 VTAIL.n170 VTAIL.n169 11.249
R443 VTAIL.n406 VTAIL.n405 11.249
R444 VTAIL.n389 VTAIL.n366 11.249
R445 VTAIL.n346 VTAIL.n345 11.249
R446 VTAIL.n329 VTAIL.n306 11.249
R447 VTAIL.n288 VTAIL.n287 11.249
R448 VTAIL.n271 VTAIL.n248 11.249
R449 VTAIL.n228 VTAIL.n227 11.249
R450 VTAIL.n211 VTAIL.n188 11.249
R451 VTAIL.n445 VTAIL.n426 10.4732
R452 VTAIL.n467 VTAIL.n416 10.4732
R453 VTAIL.n33 VTAIL.n14 10.4732
R454 VTAIL.n55 VTAIL.n4 10.4732
R455 VTAIL.n91 VTAIL.n72 10.4732
R456 VTAIL.n113 VTAIL.n62 10.4732
R457 VTAIL.n151 VTAIL.n132 10.4732
R458 VTAIL.n173 VTAIL.n122 10.4732
R459 VTAIL.n409 VTAIL.n358 10.4732
R460 VTAIL.n388 VTAIL.n369 10.4732
R461 VTAIL.n349 VTAIL.n298 10.4732
R462 VTAIL.n328 VTAIL.n309 10.4732
R463 VTAIL.n291 VTAIL.n240 10.4732
R464 VTAIL.n270 VTAIL.n251 10.4732
R465 VTAIL.n231 VTAIL.n180 10.4732
R466 VTAIL.n210 VTAIL.n191 10.4732
R467 VTAIL.n433 VTAIL.n431 10.2747
R468 VTAIL.n21 VTAIL.n19 10.2747
R469 VTAIL.n79 VTAIL.n77 10.2747
R470 VTAIL.n139 VTAIL.n137 10.2747
R471 VTAIL.n376 VTAIL.n374 10.2747
R472 VTAIL.n316 VTAIL.n314 10.2747
R473 VTAIL.n258 VTAIL.n256 10.2747
R474 VTAIL.n198 VTAIL.n196 10.2747
R475 VTAIL.n442 VTAIL.n441 9.69747
R476 VTAIL.n468 VTAIL.n414 9.69747
R477 VTAIL.n30 VTAIL.n29 9.69747
R478 VTAIL.n56 VTAIL.n2 9.69747
R479 VTAIL.n88 VTAIL.n87 9.69747
R480 VTAIL.n114 VTAIL.n60 9.69747
R481 VTAIL.n148 VTAIL.n147 9.69747
R482 VTAIL.n174 VTAIL.n120 9.69747
R483 VTAIL.n410 VTAIL.n356 9.69747
R484 VTAIL.n385 VTAIL.n384 9.69747
R485 VTAIL.n350 VTAIL.n296 9.69747
R486 VTAIL.n325 VTAIL.n324 9.69747
R487 VTAIL.n292 VTAIL.n238 9.69747
R488 VTAIL.n267 VTAIL.n266 9.69747
R489 VTAIL.n232 VTAIL.n178 9.69747
R490 VTAIL.n207 VTAIL.n206 9.69747
R491 VTAIL.n470 VTAIL.n469 9.45567
R492 VTAIL.n58 VTAIL.n57 9.45567
R493 VTAIL.n116 VTAIL.n115 9.45567
R494 VTAIL.n176 VTAIL.n175 9.45567
R495 VTAIL.n412 VTAIL.n411 9.45567
R496 VTAIL.n352 VTAIL.n351 9.45567
R497 VTAIL.n294 VTAIL.n293 9.45567
R498 VTAIL.n234 VTAIL.n233 9.45567
R499 VTAIL.n469 VTAIL.n468 9.3005
R500 VTAIL.n416 VTAIL.n415 9.3005
R501 VTAIL.n463 VTAIL.n462 9.3005
R502 VTAIL.n461 VTAIL.n460 9.3005
R503 VTAIL.n420 VTAIL.n419 9.3005
R504 VTAIL.n435 VTAIL.n434 9.3005
R505 VTAIL.n437 VTAIL.n436 9.3005
R506 VTAIL.n428 VTAIL.n427 9.3005
R507 VTAIL.n443 VTAIL.n442 9.3005
R508 VTAIL.n445 VTAIL.n444 9.3005
R509 VTAIL.n424 VTAIL.n423 9.3005
R510 VTAIL.n452 VTAIL.n451 9.3005
R511 VTAIL.n454 VTAIL.n453 9.3005
R512 VTAIL.n57 VTAIL.n56 9.3005
R513 VTAIL.n4 VTAIL.n3 9.3005
R514 VTAIL.n51 VTAIL.n50 9.3005
R515 VTAIL.n49 VTAIL.n48 9.3005
R516 VTAIL.n8 VTAIL.n7 9.3005
R517 VTAIL.n23 VTAIL.n22 9.3005
R518 VTAIL.n25 VTAIL.n24 9.3005
R519 VTAIL.n16 VTAIL.n15 9.3005
R520 VTAIL.n31 VTAIL.n30 9.3005
R521 VTAIL.n33 VTAIL.n32 9.3005
R522 VTAIL.n12 VTAIL.n11 9.3005
R523 VTAIL.n40 VTAIL.n39 9.3005
R524 VTAIL.n42 VTAIL.n41 9.3005
R525 VTAIL.n115 VTAIL.n114 9.3005
R526 VTAIL.n62 VTAIL.n61 9.3005
R527 VTAIL.n109 VTAIL.n108 9.3005
R528 VTAIL.n107 VTAIL.n106 9.3005
R529 VTAIL.n66 VTAIL.n65 9.3005
R530 VTAIL.n81 VTAIL.n80 9.3005
R531 VTAIL.n83 VTAIL.n82 9.3005
R532 VTAIL.n74 VTAIL.n73 9.3005
R533 VTAIL.n89 VTAIL.n88 9.3005
R534 VTAIL.n91 VTAIL.n90 9.3005
R535 VTAIL.n70 VTAIL.n69 9.3005
R536 VTAIL.n98 VTAIL.n97 9.3005
R537 VTAIL.n100 VTAIL.n99 9.3005
R538 VTAIL.n175 VTAIL.n174 9.3005
R539 VTAIL.n122 VTAIL.n121 9.3005
R540 VTAIL.n169 VTAIL.n168 9.3005
R541 VTAIL.n167 VTAIL.n166 9.3005
R542 VTAIL.n126 VTAIL.n125 9.3005
R543 VTAIL.n141 VTAIL.n140 9.3005
R544 VTAIL.n143 VTAIL.n142 9.3005
R545 VTAIL.n134 VTAIL.n133 9.3005
R546 VTAIL.n149 VTAIL.n148 9.3005
R547 VTAIL.n151 VTAIL.n150 9.3005
R548 VTAIL.n130 VTAIL.n129 9.3005
R549 VTAIL.n158 VTAIL.n157 9.3005
R550 VTAIL.n160 VTAIL.n159 9.3005
R551 VTAIL.n378 VTAIL.n377 9.3005
R552 VTAIL.n380 VTAIL.n379 9.3005
R553 VTAIL.n371 VTAIL.n370 9.3005
R554 VTAIL.n386 VTAIL.n385 9.3005
R555 VTAIL.n388 VTAIL.n387 9.3005
R556 VTAIL.n366 VTAIL.n365 9.3005
R557 VTAIL.n394 VTAIL.n393 9.3005
R558 VTAIL.n396 VTAIL.n395 9.3005
R559 VTAIL.n411 VTAIL.n410 9.3005
R560 VTAIL.n358 VTAIL.n357 9.3005
R561 VTAIL.n405 VTAIL.n404 9.3005
R562 VTAIL.n403 VTAIL.n402 9.3005
R563 VTAIL.n362 VTAIL.n361 9.3005
R564 VTAIL.n318 VTAIL.n317 9.3005
R565 VTAIL.n320 VTAIL.n319 9.3005
R566 VTAIL.n311 VTAIL.n310 9.3005
R567 VTAIL.n326 VTAIL.n325 9.3005
R568 VTAIL.n328 VTAIL.n327 9.3005
R569 VTAIL.n306 VTAIL.n305 9.3005
R570 VTAIL.n334 VTAIL.n333 9.3005
R571 VTAIL.n336 VTAIL.n335 9.3005
R572 VTAIL.n351 VTAIL.n350 9.3005
R573 VTAIL.n298 VTAIL.n297 9.3005
R574 VTAIL.n345 VTAIL.n344 9.3005
R575 VTAIL.n343 VTAIL.n342 9.3005
R576 VTAIL.n302 VTAIL.n301 9.3005
R577 VTAIL.n260 VTAIL.n259 9.3005
R578 VTAIL.n262 VTAIL.n261 9.3005
R579 VTAIL.n253 VTAIL.n252 9.3005
R580 VTAIL.n268 VTAIL.n267 9.3005
R581 VTAIL.n270 VTAIL.n269 9.3005
R582 VTAIL.n248 VTAIL.n247 9.3005
R583 VTAIL.n276 VTAIL.n275 9.3005
R584 VTAIL.n278 VTAIL.n277 9.3005
R585 VTAIL.n293 VTAIL.n292 9.3005
R586 VTAIL.n240 VTAIL.n239 9.3005
R587 VTAIL.n287 VTAIL.n286 9.3005
R588 VTAIL.n285 VTAIL.n284 9.3005
R589 VTAIL.n244 VTAIL.n243 9.3005
R590 VTAIL.n200 VTAIL.n199 9.3005
R591 VTAIL.n202 VTAIL.n201 9.3005
R592 VTAIL.n193 VTAIL.n192 9.3005
R593 VTAIL.n208 VTAIL.n207 9.3005
R594 VTAIL.n210 VTAIL.n209 9.3005
R595 VTAIL.n188 VTAIL.n187 9.3005
R596 VTAIL.n216 VTAIL.n215 9.3005
R597 VTAIL.n218 VTAIL.n217 9.3005
R598 VTAIL.n233 VTAIL.n232 9.3005
R599 VTAIL.n180 VTAIL.n179 9.3005
R600 VTAIL.n227 VTAIL.n226 9.3005
R601 VTAIL.n225 VTAIL.n224 9.3005
R602 VTAIL.n184 VTAIL.n183 9.3005
R603 VTAIL.n438 VTAIL.n428 8.92171
R604 VTAIL.n26 VTAIL.n16 8.92171
R605 VTAIL.n84 VTAIL.n74 8.92171
R606 VTAIL.n144 VTAIL.n134 8.92171
R607 VTAIL.n381 VTAIL.n371 8.92171
R608 VTAIL.n321 VTAIL.n311 8.92171
R609 VTAIL.n263 VTAIL.n253 8.92171
R610 VTAIL.n203 VTAIL.n193 8.92171
R611 VTAIL.n437 VTAIL.n430 8.14595
R612 VTAIL.n25 VTAIL.n18 8.14595
R613 VTAIL.n83 VTAIL.n76 8.14595
R614 VTAIL.n143 VTAIL.n136 8.14595
R615 VTAIL.n380 VTAIL.n373 8.14595
R616 VTAIL.n320 VTAIL.n313 8.14595
R617 VTAIL.n262 VTAIL.n255 8.14595
R618 VTAIL.n202 VTAIL.n195 8.14595
R619 VTAIL.n434 VTAIL.n433 7.3702
R620 VTAIL.n22 VTAIL.n21 7.3702
R621 VTAIL.n80 VTAIL.n79 7.3702
R622 VTAIL.n140 VTAIL.n139 7.3702
R623 VTAIL.n377 VTAIL.n376 7.3702
R624 VTAIL.n317 VTAIL.n316 7.3702
R625 VTAIL.n259 VTAIL.n258 7.3702
R626 VTAIL.n199 VTAIL.n198 7.3702
R627 VTAIL.n434 VTAIL.n430 5.81868
R628 VTAIL.n22 VTAIL.n18 5.81868
R629 VTAIL.n80 VTAIL.n76 5.81868
R630 VTAIL.n140 VTAIL.n136 5.81868
R631 VTAIL.n377 VTAIL.n373 5.81868
R632 VTAIL.n317 VTAIL.n313 5.81868
R633 VTAIL.n259 VTAIL.n255 5.81868
R634 VTAIL.n199 VTAIL.n195 5.81868
R635 VTAIL.n438 VTAIL.n437 5.04292
R636 VTAIL.n26 VTAIL.n25 5.04292
R637 VTAIL.n84 VTAIL.n83 5.04292
R638 VTAIL.n144 VTAIL.n143 5.04292
R639 VTAIL.n381 VTAIL.n380 5.04292
R640 VTAIL.n321 VTAIL.n320 5.04292
R641 VTAIL.n263 VTAIL.n262 5.04292
R642 VTAIL.n203 VTAIL.n202 5.04292
R643 VTAIL.n441 VTAIL.n428 4.26717
R644 VTAIL.n470 VTAIL.n414 4.26717
R645 VTAIL.n29 VTAIL.n16 4.26717
R646 VTAIL.n58 VTAIL.n2 4.26717
R647 VTAIL.n87 VTAIL.n74 4.26717
R648 VTAIL.n116 VTAIL.n60 4.26717
R649 VTAIL.n147 VTAIL.n134 4.26717
R650 VTAIL.n176 VTAIL.n120 4.26717
R651 VTAIL.n412 VTAIL.n356 4.26717
R652 VTAIL.n384 VTAIL.n371 4.26717
R653 VTAIL.n352 VTAIL.n296 4.26717
R654 VTAIL.n324 VTAIL.n311 4.26717
R655 VTAIL.n294 VTAIL.n238 4.26717
R656 VTAIL.n266 VTAIL.n253 4.26717
R657 VTAIL.n234 VTAIL.n178 4.26717
R658 VTAIL.n206 VTAIL.n193 4.26717
R659 VTAIL.n442 VTAIL.n426 3.49141
R660 VTAIL.n468 VTAIL.n467 3.49141
R661 VTAIL.n30 VTAIL.n14 3.49141
R662 VTAIL.n56 VTAIL.n55 3.49141
R663 VTAIL.n88 VTAIL.n72 3.49141
R664 VTAIL.n114 VTAIL.n113 3.49141
R665 VTAIL.n148 VTAIL.n132 3.49141
R666 VTAIL.n174 VTAIL.n173 3.49141
R667 VTAIL.n410 VTAIL.n409 3.49141
R668 VTAIL.n385 VTAIL.n369 3.49141
R669 VTAIL.n350 VTAIL.n349 3.49141
R670 VTAIL.n325 VTAIL.n309 3.49141
R671 VTAIL.n292 VTAIL.n291 3.49141
R672 VTAIL.n267 VTAIL.n251 3.49141
R673 VTAIL.n232 VTAIL.n231 3.49141
R674 VTAIL.n207 VTAIL.n191 3.49141
R675 VTAIL.n237 VTAIL.n235 3.41429
R676 VTAIL.n295 VTAIL.n237 3.41429
R677 VTAIL.n355 VTAIL.n353 3.41429
R678 VTAIL.n413 VTAIL.n355 3.41429
R679 VTAIL.n177 VTAIL.n119 3.41429
R680 VTAIL.n119 VTAIL.n117 3.41429
R681 VTAIL.n59 VTAIL.n1 3.41429
R682 VTAIL VTAIL.n471 3.3561
R683 VTAIL.n435 VTAIL.n431 2.84303
R684 VTAIL.n23 VTAIL.n19 2.84303
R685 VTAIL.n81 VTAIL.n77 2.84303
R686 VTAIL.n141 VTAIL.n137 2.84303
R687 VTAIL.n378 VTAIL.n374 2.84303
R688 VTAIL.n318 VTAIL.n314 2.84303
R689 VTAIL.n260 VTAIL.n256 2.84303
R690 VTAIL.n200 VTAIL.n196 2.84303
R691 VTAIL.n446 VTAIL.n445 2.71565
R692 VTAIL.n464 VTAIL.n416 2.71565
R693 VTAIL.n34 VTAIL.n33 2.71565
R694 VTAIL.n52 VTAIL.n4 2.71565
R695 VTAIL.n92 VTAIL.n91 2.71565
R696 VTAIL.n110 VTAIL.n62 2.71565
R697 VTAIL.n152 VTAIL.n151 2.71565
R698 VTAIL.n170 VTAIL.n122 2.71565
R699 VTAIL.n406 VTAIL.n358 2.71565
R700 VTAIL.n389 VTAIL.n388 2.71565
R701 VTAIL.n346 VTAIL.n298 2.71565
R702 VTAIL.n329 VTAIL.n328 2.71565
R703 VTAIL.n288 VTAIL.n240 2.71565
R704 VTAIL.n271 VTAIL.n270 2.71565
R705 VTAIL.n228 VTAIL.n180 2.71565
R706 VTAIL.n211 VTAIL.n210 2.71565
R707 VTAIL.n450 VTAIL.n424 1.93989
R708 VTAIL.n463 VTAIL.n418 1.93989
R709 VTAIL.n38 VTAIL.n12 1.93989
R710 VTAIL.n51 VTAIL.n6 1.93989
R711 VTAIL.n96 VTAIL.n70 1.93989
R712 VTAIL.n109 VTAIL.n64 1.93989
R713 VTAIL.n156 VTAIL.n130 1.93989
R714 VTAIL.n169 VTAIL.n124 1.93989
R715 VTAIL.n405 VTAIL.n360 1.93989
R716 VTAIL.n392 VTAIL.n366 1.93989
R717 VTAIL.n345 VTAIL.n300 1.93989
R718 VTAIL.n332 VTAIL.n306 1.93989
R719 VTAIL.n287 VTAIL.n242 1.93989
R720 VTAIL.n274 VTAIL.n248 1.93989
R721 VTAIL.n227 VTAIL.n182 1.93989
R722 VTAIL.n214 VTAIL.n188 1.93989
R723 VTAIL.n0 VTAIL.t0 1.84924
R724 VTAIL.n0 VTAIL.t5 1.84924
R725 VTAIL.n118 VTAIL.t13 1.84924
R726 VTAIL.n118 VTAIL.t12 1.84924
R727 VTAIL.n354 VTAIL.t11 1.84924
R728 VTAIL.n354 VTAIL.t9 1.84924
R729 VTAIL.n236 VTAIL.t2 1.84924
R730 VTAIL.n236 VTAIL.t7 1.84924
R731 VTAIL.n451 VTAIL.n422 1.16414
R732 VTAIL.n460 VTAIL.n459 1.16414
R733 VTAIL.n39 VTAIL.n10 1.16414
R734 VTAIL.n48 VTAIL.n47 1.16414
R735 VTAIL.n97 VTAIL.n68 1.16414
R736 VTAIL.n106 VTAIL.n105 1.16414
R737 VTAIL.n157 VTAIL.n128 1.16414
R738 VTAIL.n166 VTAIL.n165 1.16414
R739 VTAIL.n402 VTAIL.n401 1.16414
R740 VTAIL.n393 VTAIL.n364 1.16414
R741 VTAIL.n342 VTAIL.n341 1.16414
R742 VTAIL.n333 VTAIL.n304 1.16414
R743 VTAIL.n284 VTAIL.n283 1.16414
R744 VTAIL.n275 VTAIL.n246 1.16414
R745 VTAIL.n224 VTAIL.n223 1.16414
R746 VTAIL.n215 VTAIL.n186 1.16414
R747 VTAIL.n353 VTAIL.n295 0.470328
R748 VTAIL.n117 VTAIL.n59 0.470328
R749 VTAIL.n455 VTAIL.n454 0.388379
R750 VTAIL.n456 VTAIL.n420 0.388379
R751 VTAIL.n43 VTAIL.n42 0.388379
R752 VTAIL.n44 VTAIL.n8 0.388379
R753 VTAIL.n101 VTAIL.n100 0.388379
R754 VTAIL.n102 VTAIL.n66 0.388379
R755 VTAIL.n161 VTAIL.n160 0.388379
R756 VTAIL.n162 VTAIL.n126 0.388379
R757 VTAIL.n398 VTAIL.n362 0.388379
R758 VTAIL.n397 VTAIL.n396 0.388379
R759 VTAIL.n338 VTAIL.n302 0.388379
R760 VTAIL.n337 VTAIL.n336 0.388379
R761 VTAIL.n280 VTAIL.n244 0.388379
R762 VTAIL.n279 VTAIL.n278 0.388379
R763 VTAIL.n220 VTAIL.n184 0.388379
R764 VTAIL.n219 VTAIL.n218 0.388379
R765 VTAIL.n436 VTAIL.n435 0.155672
R766 VTAIL.n436 VTAIL.n427 0.155672
R767 VTAIL.n443 VTAIL.n427 0.155672
R768 VTAIL.n444 VTAIL.n443 0.155672
R769 VTAIL.n444 VTAIL.n423 0.155672
R770 VTAIL.n452 VTAIL.n423 0.155672
R771 VTAIL.n453 VTAIL.n452 0.155672
R772 VTAIL.n453 VTAIL.n419 0.155672
R773 VTAIL.n461 VTAIL.n419 0.155672
R774 VTAIL.n462 VTAIL.n461 0.155672
R775 VTAIL.n462 VTAIL.n415 0.155672
R776 VTAIL.n469 VTAIL.n415 0.155672
R777 VTAIL.n24 VTAIL.n23 0.155672
R778 VTAIL.n24 VTAIL.n15 0.155672
R779 VTAIL.n31 VTAIL.n15 0.155672
R780 VTAIL.n32 VTAIL.n31 0.155672
R781 VTAIL.n32 VTAIL.n11 0.155672
R782 VTAIL.n40 VTAIL.n11 0.155672
R783 VTAIL.n41 VTAIL.n40 0.155672
R784 VTAIL.n41 VTAIL.n7 0.155672
R785 VTAIL.n49 VTAIL.n7 0.155672
R786 VTAIL.n50 VTAIL.n49 0.155672
R787 VTAIL.n50 VTAIL.n3 0.155672
R788 VTAIL.n57 VTAIL.n3 0.155672
R789 VTAIL.n82 VTAIL.n81 0.155672
R790 VTAIL.n82 VTAIL.n73 0.155672
R791 VTAIL.n89 VTAIL.n73 0.155672
R792 VTAIL.n90 VTAIL.n89 0.155672
R793 VTAIL.n90 VTAIL.n69 0.155672
R794 VTAIL.n98 VTAIL.n69 0.155672
R795 VTAIL.n99 VTAIL.n98 0.155672
R796 VTAIL.n99 VTAIL.n65 0.155672
R797 VTAIL.n107 VTAIL.n65 0.155672
R798 VTAIL.n108 VTAIL.n107 0.155672
R799 VTAIL.n108 VTAIL.n61 0.155672
R800 VTAIL.n115 VTAIL.n61 0.155672
R801 VTAIL.n142 VTAIL.n141 0.155672
R802 VTAIL.n142 VTAIL.n133 0.155672
R803 VTAIL.n149 VTAIL.n133 0.155672
R804 VTAIL.n150 VTAIL.n149 0.155672
R805 VTAIL.n150 VTAIL.n129 0.155672
R806 VTAIL.n158 VTAIL.n129 0.155672
R807 VTAIL.n159 VTAIL.n158 0.155672
R808 VTAIL.n159 VTAIL.n125 0.155672
R809 VTAIL.n167 VTAIL.n125 0.155672
R810 VTAIL.n168 VTAIL.n167 0.155672
R811 VTAIL.n168 VTAIL.n121 0.155672
R812 VTAIL.n175 VTAIL.n121 0.155672
R813 VTAIL.n411 VTAIL.n357 0.155672
R814 VTAIL.n404 VTAIL.n357 0.155672
R815 VTAIL.n404 VTAIL.n403 0.155672
R816 VTAIL.n403 VTAIL.n361 0.155672
R817 VTAIL.n395 VTAIL.n361 0.155672
R818 VTAIL.n395 VTAIL.n394 0.155672
R819 VTAIL.n394 VTAIL.n365 0.155672
R820 VTAIL.n387 VTAIL.n365 0.155672
R821 VTAIL.n387 VTAIL.n386 0.155672
R822 VTAIL.n386 VTAIL.n370 0.155672
R823 VTAIL.n379 VTAIL.n370 0.155672
R824 VTAIL.n379 VTAIL.n378 0.155672
R825 VTAIL.n351 VTAIL.n297 0.155672
R826 VTAIL.n344 VTAIL.n297 0.155672
R827 VTAIL.n344 VTAIL.n343 0.155672
R828 VTAIL.n343 VTAIL.n301 0.155672
R829 VTAIL.n335 VTAIL.n301 0.155672
R830 VTAIL.n335 VTAIL.n334 0.155672
R831 VTAIL.n334 VTAIL.n305 0.155672
R832 VTAIL.n327 VTAIL.n305 0.155672
R833 VTAIL.n327 VTAIL.n326 0.155672
R834 VTAIL.n326 VTAIL.n310 0.155672
R835 VTAIL.n319 VTAIL.n310 0.155672
R836 VTAIL.n319 VTAIL.n318 0.155672
R837 VTAIL.n293 VTAIL.n239 0.155672
R838 VTAIL.n286 VTAIL.n239 0.155672
R839 VTAIL.n286 VTAIL.n285 0.155672
R840 VTAIL.n285 VTAIL.n243 0.155672
R841 VTAIL.n277 VTAIL.n243 0.155672
R842 VTAIL.n277 VTAIL.n276 0.155672
R843 VTAIL.n276 VTAIL.n247 0.155672
R844 VTAIL.n269 VTAIL.n247 0.155672
R845 VTAIL.n269 VTAIL.n268 0.155672
R846 VTAIL.n268 VTAIL.n252 0.155672
R847 VTAIL.n261 VTAIL.n252 0.155672
R848 VTAIL.n261 VTAIL.n260 0.155672
R849 VTAIL.n233 VTAIL.n179 0.155672
R850 VTAIL.n226 VTAIL.n179 0.155672
R851 VTAIL.n226 VTAIL.n225 0.155672
R852 VTAIL.n225 VTAIL.n183 0.155672
R853 VTAIL.n217 VTAIL.n183 0.155672
R854 VTAIL.n217 VTAIL.n216 0.155672
R855 VTAIL.n216 VTAIL.n187 0.155672
R856 VTAIL.n209 VTAIL.n187 0.155672
R857 VTAIL.n209 VTAIL.n208 0.155672
R858 VTAIL.n208 VTAIL.n192 0.155672
R859 VTAIL.n201 VTAIL.n192 0.155672
R860 VTAIL.n201 VTAIL.n200 0.155672
R861 VTAIL VTAIL.n1 0.0586897
R862 VDD1 VDD1.n0 64.6872
R863 VDD1.n3 VDD1.n2 64.5735
R864 VDD1.n3 VDD1.n1 64.5735
R865 VDD1.n5 VDD1.n4 62.9219
R866 VDD1.n5 VDD1.n3 48.8931
R867 VDD1.n4 VDD1.t5 1.84924
R868 VDD1.n4 VDD1.t7 1.84924
R869 VDD1.n0 VDD1.t0 1.84924
R870 VDD1.n0 VDD1.t4 1.84924
R871 VDD1.n2 VDD1.t1 1.84924
R872 VDD1.n2 VDD1.t6 1.84924
R873 VDD1.n1 VDD1.t3 1.84924
R874 VDD1.n1 VDD1.t2 1.84924
R875 VDD1 VDD1.n5 1.64921
R876 B.n801 B.n800 585
R877 B.n801 B.n121 585
R878 B.n804 B.n803 585
R879 B.n805 B.n168 585
R880 B.n807 B.n806 585
R881 B.n809 B.n167 585
R882 B.n812 B.n811 585
R883 B.n813 B.n166 585
R884 B.n815 B.n814 585
R885 B.n817 B.n165 585
R886 B.n820 B.n819 585
R887 B.n821 B.n164 585
R888 B.n823 B.n822 585
R889 B.n825 B.n163 585
R890 B.n828 B.n827 585
R891 B.n829 B.n162 585
R892 B.n831 B.n830 585
R893 B.n833 B.n161 585
R894 B.n836 B.n835 585
R895 B.n837 B.n160 585
R896 B.n839 B.n838 585
R897 B.n841 B.n159 585
R898 B.n844 B.n843 585
R899 B.n845 B.n158 585
R900 B.n847 B.n846 585
R901 B.n849 B.n157 585
R902 B.n852 B.n851 585
R903 B.n853 B.n156 585
R904 B.n855 B.n854 585
R905 B.n857 B.n155 585
R906 B.n860 B.n859 585
R907 B.n861 B.n154 585
R908 B.n863 B.n862 585
R909 B.n865 B.n153 585
R910 B.n868 B.n867 585
R911 B.n869 B.n152 585
R912 B.n871 B.n870 585
R913 B.n873 B.n151 585
R914 B.n876 B.n875 585
R915 B.n878 B.n148 585
R916 B.n880 B.n879 585
R917 B.n882 B.n147 585
R918 B.n885 B.n884 585
R919 B.n886 B.n146 585
R920 B.n888 B.n887 585
R921 B.n890 B.n145 585
R922 B.n892 B.n891 585
R923 B.n894 B.n893 585
R924 B.n897 B.n896 585
R925 B.n898 B.n140 585
R926 B.n900 B.n899 585
R927 B.n902 B.n139 585
R928 B.n905 B.n904 585
R929 B.n906 B.n138 585
R930 B.n908 B.n907 585
R931 B.n910 B.n137 585
R932 B.n913 B.n912 585
R933 B.n914 B.n136 585
R934 B.n916 B.n915 585
R935 B.n918 B.n135 585
R936 B.n921 B.n920 585
R937 B.n922 B.n134 585
R938 B.n924 B.n923 585
R939 B.n926 B.n133 585
R940 B.n929 B.n928 585
R941 B.n930 B.n132 585
R942 B.n932 B.n931 585
R943 B.n934 B.n131 585
R944 B.n937 B.n936 585
R945 B.n938 B.n130 585
R946 B.n940 B.n939 585
R947 B.n942 B.n129 585
R948 B.n945 B.n944 585
R949 B.n946 B.n128 585
R950 B.n948 B.n947 585
R951 B.n950 B.n127 585
R952 B.n953 B.n952 585
R953 B.n954 B.n126 585
R954 B.n956 B.n955 585
R955 B.n958 B.n125 585
R956 B.n961 B.n960 585
R957 B.n962 B.n124 585
R958 B.n964 B.n963 585
R959 B.n966 B.n123 585
R960 B.n969 B.n968 585
R961 B.n970 B.n122 585
R962 B.n799 B.n120 585
R963 B.n973 B.n120 585
R964 B.n798 B.n119 585
R965 B.n974 B.n119 585
R966 B.n797 B.n118 585
R967 B.n975 B.n118 585
R968 B.n796 B.n795 585
R969 B.n795 B.n114 585
R970 B.n794 B.n113 585
R971 B.n981 B.n113 585
R972 B.n793 B.n112 585
R973 B.n982 B.n112 585
R974 B.n792 B.n111 585
R975 B.n983 B.n111 585
R976 B.n791 B.n790 585
R977 B.n790 B.n107 585
R978 B.n789 B.n106 585
R979 B.n989 B.n106 585
R980 B.n788 B.n105 585
R981 B.n990 B.n105 585
R982 B.n787 B.n104 585
R983 B.n991 B.n104 585
R984 B.n786 B.n785 585
R985 B.n785 B.n100 585
R986 B.n784 B.n99 585
R987 B.n997 B.n99 585
R988 B.n783 B.n98 585
R989 B.n998 B.n98 585
R990 B.n782 B.n97 585
R991 B.n999 B.n97 585
R992 B.n781 B.n780 585
R993 B.n780 B.n93 585
R994 B.n779 B.n92 585
R995 B.n1005 B.n92 585
R996 B.n778 B.n91 585
R997 B.n1006 B.n91 585
R998 B.n777 B.n90 585
R999 B.n1007 B.n90 585
R1000 B.n776 B.n775 585
R1001 B.n775 B.n86 585
R1002 B.n774 B.n85 585
R1003 B.n1013 B.n85 585
R1004 B.n773 B.n84 585
R1005 B.n1014 B.n84 585
R1006 B.n772 B.n83 585
R1007 B.n1015 B.n83 585
R1008 B.n771 B.n770 585
R1009 B.n770 B.n79 585
R1010 B.n769 B.n78 585
R1011 B.n1021 B.n78 585
R1012 B.n768 B.n77 585
R1013 B.n1022 B.n77 585
R1014 B.n767 B.n76 585
R1015 B.n1023 B.n76 585
R1016 B.n766 B.n765 585
R1017 B.n765 B.n72 585
R1018 B.n764 B.n71 585
R1019 B.n1029 B.n71 585
R1020 B.n763 B.n70 585
R1021 B.n1030 B.n70 585
R1022 B.n762 B.n69 585
R1023 B.n1031 B.n69 585
R1024 B.n761 B.n760 585
R1025 B.n760 B.n65 585
R1026 B.n759 B.n64 585
R1027 B.n1037 B.n64 585
R1028 B.n758 B.n63 585
R1029 B.n1038 B.n63 585
R1030 B.n757 B.n62 585
R1031 B.n1039 B.n62 585
R1032 B.n756 B.n755 585
R1033 B.n755 B.n61 585
R1034 B.n754 B.n57 585
R1035 B.n1045 B.n57 585
R1036 B.n753 B.n56 585
R1037 B.n1046 B.n56 585
R1038 B.n752 B.n55 585
R1039 B.n1047 B.n55 585
R1040 B.n751 B.n750 585
R1041 B.n750 B.n51 585
R1042 B.n749 B.n50 585
R1043 B.n1053 B.n50 585
R1044 B.n748 B.n49 585
R1045 B.n1054 B.n49 585
R1046 B.n747 B.n48 585
R1047 B.n1055 B.n48 585
R1048 B.n746 B.n745 585
R1049 B.n745 B.n44 585
R1050 B.n744 B.n43 585
R1051 B.n1061 B.n43 585
R1052 B.n743 B.n42 585
R1053 B.n1062 B.n42 585
R1054 B.n742 B.n41 585
R1055 B.n1063 B.n41 585
R1056 B.n741 B.n740 585
R1057 B.n740 B.n40 585
R1058 B.n739 B.n36 585
R1059 B.n1069 B.n36 585
R1060 B.n738 B.n35 585
R1061 B.n1070 B.n35 585
R1062 B.n737 B.n34 585
R1063 B.n1071 B.n34 585
R1064 B.n736 B.n735 585
R1065 B.n735 B.n30 585
R1066 B.n734 B.n29 585
R1067 B.n1077 B.n29 585
R1068 B.n733 B.n28 585
R1069 B.n1078 B.n28 585
R1070 B.n732 B.n27 585
R1071 B.n1079 B.n27 585
R1072 B.n731 B.n730 585
R1073 B.n730 B.n23 585
R1074 B.n729 B.n22 585
R1075 B.n1085 B.n22 585
R1076 B.n728 B.n21 585
R1077 B.n1086 B.n21 585
R1078 B.n727 B.n20 585
R1079 B.n1087 B.n20 585
R1080 B.n726 B.n725 585
R1081 B.n725 B.n19 585
R1082 B.n724 B.n15 585
R1083 B.n1093 B.n15 585
R1084 B.n723 B.n14 585
R1085 B.n1094 B.n14 585
R1086 B.n722 B.n13 585
R1087 B.n1095 B.n13 585
R1088 B.n721 B.n720 585
R1089 B.n720 B.n12 585
R1090 B.n719 B.n718 585
R1091 B.n719 B.n8 585
R1092 B.n717 B.n7 585
R1093 B.n1102 B.n7 585
R1094 B.n716 B.n6 585
R1095 B.n1103 B.n6 585
R1096 B.n715 B.n5 585
R1097 B.n1104 B.n5 585
R1098 B.n714 B.n713 585
R1099 B.n713 B.n4 585
R1100 B.n712 B.n169 585
R1101 B.n712 B.n711 585
R1102 B.n702 B.n170 585
R1103 B.n171 B.n170 585
R1104 B.n704 B.n703 585
R1105 B.n705 B.n704 585
R1106 B.n701 B.n176 585
R1107 B.n176 B.n175 585
R1108 B.n700 B.n699 585
R1109 B.n699 B.n698 585
R1110 B.n178 B.n177 585
R1111 B.n691 B.n178 585
R1112 B.n690 B.n689 585
R1113 B.n692 B.n690 585
R1114 B.n688 B.n183 585
R1115 B.n183 B.n182 585
R1116 B.n687 B.n686 585
R1117 B.n686 B.n685 585
R1118 B.n185 B.n184 585
R1119 B.n186 B.n185 585
R1120 B.n678 B.n677 585
R1121 B.n679 B.n678 585
R1122 B.n676 B.n191 585
R1123 B.n191 B.n190 585
R1124 B.n675 B.n674 585
R1125 B.n674 B.n673 585
R1126 B.n193 B.n192 585
R1127 B.n194 B.n193 585
R1128 B.n666 B.n665 585
R1129 B.n667 B.n666 585
R1130 B.n664 B.n199 585
R1131 B.n199 B.n198 585
R1132 B.n663 B.n662 585
R1133 B.n662 B.n661 585
R1134 B.n201 B.n200 585
R1135 B.n654 B.n201 585
R1136 B.n653 B.n652 585
R1137 B.n655 B.n653 585
R1138 B.n651 B.n206 585
R1139 B.n206 B.n205 585
R1140 B.n650 B.n649 585
R1141 B.n649 B.n648 585
R1142 B.n208 B.n207 585
R1143 B.n209 B.n208 585
R1144 B.n641 B.n640 585
R1145 B.n642 B.n641 585
R1146 B.n639 B.n214 585
R1147 B.n214 B.n213 585
R1148 B.n638 B.n637 585
R1149 B.n637 B.n636 585
R1150 B.n216 B.n215 585
R1151 B.n217 B.n216 585
R1152 B.n629 B.n628 585
R1153 B.n630 B.n629 585
R1154 B.n627 B.n222 585
R1155 B.n222 B.n221 585
R1156 B.n626 B.n625 585
R1157 B.n625 B.n624 585
R1158 B.n224 B.n223 585
R1159 B.n617 B.n224 585
R1160 B.n616 B.n615 585
R1161 B.n618 B.n616 585
R1162 B.n614 B.n229 585
R1163 B.n229 B.n228 585
R1164 B.n613 B.n612 585
R1165 B.n612 B.n611 585
R1166 B.n231 B.n230 585
R1167 B.n232 B.n231 585
R1168 B.n604 B.n603 585
R1169 B.n605 B.n604 585
R1170 B.n602 B.n237 585
R1171 B.n237 B.n236 585
R1172 B.n601 B.n600 585
R1173 B.n600 B.n599 585
R1174 B.n239 B.n238 585
R1175 B.n240 B.n239 585
R1176 B.n592 B.n591 585
R1177 B.n593 B.n592 585
R1178 B.n590 B.n245 585
R1179 B.n245 B.n244 585
R1180 B.n589 B.n588 585
R1181 B.n588 B.n587 585
R1182 B.n247 B.n246 585
R1183 B.n248 B.n247 585
R1184 B.n580 B.n579 585
R1185 B.n581 B.n580 585
R1186 B.n578 B.n253 585
R1187 B.n253 B.n252 585
R1188 B.n577 B.n576 585
R1189 B.n576 B.n575 585
R1190 B.n255 B.n254 585
R1191 B.n256 B.n255 585
R1192 B.n568 B.n567 585
R1193 B.n569 B.n568 585
R1194 B.n566 B.n261 585
R1195 B.n261 B.n260 585
R1196 B.n565 B.n564 585
R1197 B.n564 B.n563 585
R1198 B.n263 B.n262 585
R1199 B.n264 B.n263 585
R1200 B.n556 B.n555 585
R1201 B.n557 B.n556 585
R1202 B.n554 B.n269 585
R1203 B.n269 B.n268 585
R1204 B.n553 B.n552 585
R1205 B.n552 B.n551 585
R1206 B.n271 B.n270 585
R1207 B.n272 B.n271 585
R1208 B.n544 B.n543 585
R1209 B.n545 B.n544 585
R1210 B.n542 B.n276 585
R1211 B.n280 B.n276 585
R1212 B.n541 B.n540 585
R1213 B.n540 B.n539 585
R1214 B.n278 B.n277 585
R1215 B.n279 B.n278 585
R1216 B.n532 B.n531 585
R1217 B.n533 B.n532 585
R1218 B.n530 B.n285 585
R1219 B.n285 B.n284 585
R1220 B.n529 B.n528 585
R1221 B.n528 B.n527 585
R1222 B.n287 B.n286 585
R1223 B.n288 B.n287 585
R1224 B.n520 B.n519 585
R1225 B.n521 B.n520 585
R1226 B.n518 B.n293 585
R1227 B.n293 B.n292 585
R1228 B.n517 B.n516 585
R1229 B.n516 B.n515 585
R1230 B.n512 B.n297 585
R1231 B.n511 B.n510 585
R1232 B.n508 B.n298 585
R1233 B.n508 B.n296 585
R1234 B.n507 B.n506 585
R1235 B.n505 B.n504 585
R1236 B.n503 B.n300 585
R1237 B.n501 B.n500 585
R1238 B.n499 B.n301 585
R1239 B.n498 B.n497 585
R1240 B.n495 B.n302 585
R1241 B.n493 B.n492 585
R1242 B.n491 B.n303 585
R1243 B.n490 B.n489 585
R1244 B.n487 B.n304 585
R1245 B.n485 B.n484 585
R1246 B.n483 B.n305 585
R1247 B.n482 B.n481 585
R1248 B.n479 B.n306 585
R1249 B.n477 B.n476 585
R1250 B.n475 B.n307 585
R1251 B.n474 B.n473 585
R1252 B.n471 B.n308 585
R1253 B.n469 B.n468 585
R1254 B.n467 B.n309 585
R1255 B.n466 B.n465 585
R1256 B.n463 B.n310 585
R1257 B.n461 B.n460 585
R1258 B.n459 B.n311 585
R1259 B.n458 B.n457 585
R1260 B.n455 B.n312 585
R1261 B.n453 B.n452 585
R1262 B.n451 B.n313 585
R1263 B.n450 B.n449 585
R1264 B.n447 B.n314 585
R1265 B.n445 B.n444 585
R1266 B.n443 B.n315 585
R1267 B.n442 B.n441 585
R1268 B.n439 B.n316 585
R1269 B.n437 B.n436 585
R1270 B.n435 B.n317 585
R1271 B.n434 B.n433 585
R1272 B.n431 B.n321 585
R1273 B.n429 B.n428 585
R1274 B.n427 B.n322 585
R1275 B.n426 B.n425 585
R1276 B.n423 B.n323 585
R1277 B.n421 B.n420 585
R1278 B.n418 B.n324 585
R1279 B.n417 B.n416 585
R1280 B.n414 B.n327 585
R1281 B.n412 B.n411 585
R1282 B.n410 B.n328 585
R1283 B.n409 B.n408 585
R1284 B.n406 B.n329 585
R1285 B.n404 B.n403 585
R1286 B.n402 B.n330 585
R1287 B.n401 B.n400 585
R1288 B.n398 B.n331 585
R1289 B.n396 B.n395 585
R1290 B.n394 B.n332 585
R1291 B.n393 B.n392 585
R1292 B.n390 B.n333 585
R1293 B.n388 B.n387 585
R1294 B.n386 B.n334 585
R1295 B.n385 B.n384 585
R1296 B.n382 B.n335 585
R1297 B.n380 B.n379 585
R1298 B.n378 B.n336 585
R1299 B.n377 B.n376 585
R1300 B.n374 B.n337 585
R1301 B.n372 B.n371 585
R1302 B.n370 B.n338 585
R1303 B.n369 B.n368 585
R1304 B.n366 B.n339 585
R1305 B.n364 B.n363 585
R1306 B.n362 B.n340 585
R1307 B.n361 B.n360 585
R1308 B.n358 B.n341 585
R1309 B.n356 B.n355 585
R1310 B.n354 B.n342 585
R1311 B.n353 B.n352 585
R1312 B.n350 B.n343 585
R1313 B.n348 B.n347 585
R1314 B.n346 B.n345 585
R1315 B.n295 B.n294 585
R1316 B.n514 B.n513 585
R1317 B.n515 B.n514 585
R1318 B.n291 B.n290 585
R1319 B.n292 B.n291 585
R1320 B.n523 B.n522 585
R1321 B.n522 B.n521 585
R1322 B.n524 B.n289 585
R1323 B.n289 B.n288 585
R1324 B.n526 B.n525 585
R1325 B.n527 B.n526 585
R1326 B.n283 B.n282 585
R1327 B.n284 B.n283 585
R1328 B.n535 B.n534 585
R1329 B.n534 B.n533 585
R1330 B.n536 B.n281 585
R1331 B.n281 B.n279 585
R1332 B.n538 B.n537 585
R1333 B.n539 B.n538 585
R1334 B.n275 B.n274 585
R1335 B.n280 B.n275 585
R1336 B.n547 B.n546 585
R1337 B.n546 B.n545 585
R1338 B.n548 B.n273 585
R1339 B.n273 B.n272 585
R1340 B.n550 B.n549 585
R1341 B.n551 B.n550 585
R1342 B.n267 B.n266 585
R1343 B.n268 B.n267 585
R1344 B.n559 B.n558 585
R1345 B.n558 B.n557 585
R1346 B.n560 B.n265 585
R1347 B.n265 B.n264 585
R1348 B.n562 B.n561 585
R1349 B.n563 B.n562 585
R1350 B.n259 B.n258 585
R1351 B.n260 B.n259 585
R1352 B.n571 B.n570 585
R1353 B.n570 B.n569 585
R1354 B.n572 B.n257 585
R1355 B.n257 B.n256 585
R1356 B.n574 B.n573 585
R1357 B.n575 B.n574 585
R1358 B.n251 B.n250 585
R1359 B.n252 B.n251 585
R1360 B.n583 B.n582 585
R1361 B.n582 B.n581 585
R1362 B.n584 B.n249 585
R1363 B.n249 B.n248 585
R1364 B.n586 B.n585 585
R1365 B.n587 B.n586 585
R1366 B.n243 B.n242 585
R1367 B.n244 B.n243 585
R1368 B.n595 B.n594 585
R1369 B.n594 B.n593 585
R1370 B.n596 B.n241 585
R1371 B.n241 B.n240 585
R1372 B.n598 B.n597 585
R1373 B.n599 B.n598 585
R1374 B.n235 B.n234 585
R1375 B.n236 B.n235 585
R1376 B.n607 B.n606 585
R1377 B.n606 B.n605 585
R1378 B.n608 B.n233 585
R1379 B.n233 B.n232 585
R1380 B.n610 B.n609 585
R1381 B.n611 B.n610 585
R1382 B.n227 B.n226 585
R1383 B.n228 B.n227 585
R1384 B.n620 B.n619 585
R1385 B.n619 B.n618 585
R1386 B.n621 B.n225 585
R1387 B.n617 B.n225 585
R1388 B.n623 B.n622 585
R1389 B.n624 B.n623 585
R1390 B.n220 B.n219 585
R1391 B.n221 B.n220 585
R1392 B.n632 B.n631 585
R1393 B.n631 B.n630 585
R1394 B.n633 B.n218 585
R1395 B.n218 B.n217 585
R1396 B.n635 B.n634 585
R1397 B.n636 B.n635 585
R1398 B.n212 B.n211 585
R1399 B.n213 B.n212 585
R1400 B.n644 B.n643 585
R1401 B.n643 B.n642 585
R1402 B.n645 B.n210 585
R1403 B.n210 B.n209 585
R1404 B.n647 B.n646 585
R1405 B.n648 B.n647 585
R1406 B.n204 B.n203 585
R1407 B.n205 B.n204 585
R1408 B.n657 B.n656 585
R1409 B.n656 B.n655 585
R1410 B.n658 B.n202 585
R1411 B.n654 B.n202 585
R1412 B.n660 B.n659 585
R1413 B.n661 B.n660 585
R1414 B.n197 B.n196 585
R1415 B.n198 B.n197 585
R1416 B.n669 B.n668 585
R1417 B.n668 B.n667 585
R1418 B.n670 B.n195 585
R1419 B.n195 B.n194 585
R1420 B.n672 B.n671 585
R1421 B.n673 B.n672 585
R1422 B.n189 B.n188 585
R1423 B.n190 B.n189 585
R1424 B.n681 B.n680 585
R1425 B.n680 B.n679 585
R1426 B.n682 B.n187 585
R1427 B.n187 B.n186 585
R1428 B.n684 B.n683 585
R1429 B.n685 B.n684 585
R1430 B.n181 B.n180 585
R1431 B.n182 B.n181 585
R1432 B.n694 B.n693 585
R1433 B.n693 B.n692 585
R1434 B.n695 B.n179 585
R1435 B.n691 B.n179 585
R1436 B.n697 B.n696 585
R1437 B.n698 B.n697 585
R1438 B.n174 B.n173 585
R1439 B.n175 B.n174 585
R1440 B.n707 B.n706 585
R1441 B.n706 B.n705 585
R1442 B.n708 B.n172 585
R1443 B.n172 B.n171 585
R1444 B.n710 B.n709 585
R1445 B.n711 B.n710 585
R1446 B.n3 B.n0 585
R1447 B.n4 B.n3 585
R1448 B.n1101 B.n1 585
R1449 B.n1102 B.n1101 585
R1450 B.n1100 B.n1099 585
R1451 B.n1100 B.n8 585
R1452 B.n1098 B.n9 585
R1453 B.n12 B.n9 585
R1454 B.n1097 B.n1096 585
R1455 B.n1096 B.n1095 585
R1456 B.n11 B.n10 585
R1457 B.n1094 B.n11 585
R1458 B.n1092 B.n1091 585
R1459 B.n1093 B.n1092 585
R1460 B.n1090 B.n16 585
R1461 B.n19 B.n16 585
R1462 B.n1089 B.n1088 585
R1463 B.n1088 B.n1087 585
R1464 B.n18 B.n17 585
R1465 B.n1086 B.n18 585
R1466 B.n1084 B.n1083 585
R1467 B.n1085 B.n1084 585
R1468 B.n1082 B.n24 585
R1469 B.n24 B.n23 585
R1470 B.n1081 B.n1080 585
R1471 B.n1080 B.n1079 585
R1472 B.n26 B.n25 585
R1473 B.n1078 B.n26 585
R1474 B.n1076 B.n1075 585
R1475 B.n1077 B.n1076 585
R1476 B.n1074 B.n31 585
R1477 B.n31 B.n30 585
R1478 B.n1073 B.n1072 585
R1479 B.n1072 B.n1071 585
R1480 B.n33 B.n32 585
R1481 B.n1070 B.n33 585
R1482 B.n1068 B.n1067 585
R1483 B.n1069 B.n1068 585
R1484 B.n1066 B.n37 585
R1485 B.n40 B.n37 585
R1486 B.n1065 B.n1064 585
R1487 B.n1064 B.n1063 585
R1488 B.n39 B.n38 585
R1489 B.n1062 B.n39 585
R1490 B.n1060 B.n1059 585
R1491 B.n1061 B.n1060 585
R1492 B.n1058 B.n45 585
R1493 B.n45 B.n44 585
R1494 B.n1057 B.n1056 585
R1495 B.n1056 B.n1055 585
R1496 B.n47 B.n46 585
R1497 B.n1054 B.n47 585
R1498 B.n1052 B.n1051 585
R1499 B.n1053 B.n1052 585
R1500 B.n1050 B.n52 585
R1501 B.n52 B.n51 585
R1502 B.n1049 B.n1048 585
R1503 B.n1048 B.n1047 585
R1504 B.n54 B.n53 585
R1505 B.n1046 B.n54 585
R1506 B.n1044 B.n1043 585
R1507 B.n1045 B.n1044 585
R1508 B.n1042 B.n58 585
R1509 B.n61 B.n58 585
R1510 B.n1041 B.n1040 585
R1511 B.n1040 B.n1039 585
R1512 B.n60 B.n59 585
R1513 B.n1038 B.n60 585
R1514 B.n1036 B.n1035 585
R1515 B.n1037 B.n1036 585
R1516 B.n1034 B.n66 585
R1517 B.n66 B.n65 585
R1518 B.n1033 B.n1032 585
R1519 B.n1032 B.n1031 585
R1520 B.n68 B.n67 585
R1521 B.n1030 B.n68 585
R1522 B.n1028 B.n1027 585
R1523 B.n1029 B.n1028 585
R1524 B.n1026 B.n73 585
R1525 B.n73 B.n72 585
R1526 B.n1025 B.n1024 585
R1527 B.n1024 B.n1023 585
R1528 B.n75 B.n74 585
R1529 B.n1022 B.n75 585
R1530 B.n1020 B.n1019 585
R1531 B.n1021 B.n1020 585
R1532 B.n1018 B.n80 585
R1533 B.n80 B.n79 585
R1534 B.n1017 B.n1016 585
R1535 B.n1016 B.n1015 585
R1536 B.n82 B.n81 585
R1537 B.n1014 B.n82 585
R1538 B.n1012 B.n1011 585
R1539 B.n1013 B.n1012 585
R1540 B.n1010 B.n87 585
R1541 B.n87 B.n86 585
R1542 B.n1009 B.n1008 585
R1543 B.n1008 B.n1007 585
R1544 B.n89 B.n88 585
R1545 B.n1006 B.n89 585
R1546 B.n1004 B.n1003 585
R1547 B.n1005 B.n1004 585
R1548 B.n1002 B.n94 585
R1549 B.n94 B.n93 585
R1550 B.n1001 B.n1000 585
R1551 B.n1000 B.n999 585
R1552 B.n96 B.n95 585
R1553 B.n998 B.n96 585
R1554 B.n996 B.n995 585
R1555 B.n997 B.n996 585
R1556 B.n994 B.n101 585
R1557 B.n101 B.n100 585
R1558 B.n993 B.n992 585
R1559 B.n992 B.n991 585
R1560 B.n103 B.n102 585
R1561 B.n990 B.n103 585
R1562 B.n988 B.n987 585
R1563 B.n989 B.n988 585
R1564 B.n986 B.n108 585
R1565 B.n108 B.n107 585
R1566 B.n985 B.n984 585
R1567 B.n984 B.n983 585
R1568 B.n110 B.n109 585
R1569 B.n982 B.n110 585
R1570 B.n980 B.n979 585
R1571 B.n981 B.n980 585
R1572 B.n978 B.n115 585
R1573 B.n115 B.n114 585
R1574 B.n977 B.n976 585
R1575 B.n976 B.n975 585
R1576 B.n117 B.n116 585
R1577 B.n974 B.n117 585
R1578 B.n972 B.n971 585
R1579 B.n973 B.n972 585
R1580 B.n1105 B.n1104 585
R1581 B.n1103 B.n2 585
R1582 B.n972 B.n122 492.5
R1583 B.n801 B.n120 492.5
R1584 B.n516 B.n295 492.5
R1585 B.n514 B.n297 492.5
R1586 B.n149 B.t17 336.741
R1587 B.n325 B.t21 336.741
R1588 B.n141 B.t14 336.741
R1589 B.n318 B.t11 336.741
R1590 B.n141 B.t12 280.312
R1591 B.n149 B.t16 280.312
R1592 B.n325 B.t19 280.312
R1593 B.n318 B.t8 280.312
R1594 B.n150 B.t18 259.942
R1595 B.n326 B.t20 259.942
R1596 B.n142 B.t15 259.942
R1597 B.n319 B.t10 259.942
R1598 B.n802 B.n121 256.663
R1599 B.n808 B.n121 256.663
R1600 B.n810 B.n121 256.663
R1601 B.n816 B.n121 256.663
R1602 B.n818 B.n121 256.663
R1603 B.n824 B.n121 256.663
R1604 B.n826 B.n121 256.663
R1605 B.n832 B.n121 256.663
R1606 B.n834 B.n121 256.663
R1607 B.n840 B.n121 256.663
R1608 B.n842 B.n121 256.663
R1609 B.n848 B.n121 256.663
R1610 B.n850 B.n121 256.663
R1611 B.n856 B.n121 256.663
R1612 B.n858 B.n121 256.663
R1613 B.n864 B.n121 256.663
R1614 B.n866 B.n121 256.663
R1615 B.n872 B.n121 256.663
R1616 B.n874 B.n121 256.663
R1617 B.n881 B.n121 256.663
R1618 B.n883 B.n121 256.663
R1619 B.n889 B.n121 256.663
R1620 B.n144 B.n121 256.663
R1621 B.n895 B.n121 256.663
R1622 B.n901 B.n121 256.663
R1623 B.n903 B.n121 256.663
R1624 B.n909 B.n121 256.663
R1625 B.n911 B.n121 256.663
R1626 B.n917 B.n121 256.663
R1627 B.n919 B.n121 256.663
R1628 B.n925 B.n121 256.663
R1629 B.n927 B.n121 256.663
R1630 B.n933 B.n121 256.663
R1631 B.n935 B.n121 256.663
R1632 B.n941 B.n121 256.663
R1633 B.n943 B.n121 256.663
R1634 B.n949 B.n121 256.663
R1635 B.n951 B.n121 256.663
R1636 B.n957 B.n121 256.663
R1637 B.n959 B.n121 256.663
R1638 B.n965 B.n121 256.663
R1639 B.n967 B.n121 256.663
R1640 B.n509 B.n296 256.663
R1641 B.n299 B.n296 256.663
R1642 B.n502 B.n296 256.663
R1643 B.n496 B.n296 256.663
R1644 B.n494 B.n296 256.663
R1645 B.n488 B.n296 256.663
R1646 B.n486 B.n296 256.663
R1647 B.n480 B.n296 256.663
R1648 B.n478 B.n296 256.663
R1649 B.n472 B.n296 256.663
R1650 B.n470 B.n296 256.663
R1651 B.n464 B.n296 256.663
R1652 B.n462 B.n296 256.663
R1653 B.n456 B.n296 256.663
R1654 B.n454 B.n296 256.663
R1655 B.n448 B.n296 256.663
R1656 B.n446 B.n296 256.663
R1657 B.n440 B.n296 256.663
R1658 B.n438 B.n296 256.663
R1659 B.n432 B.n296 256.663
R1660 B.n430 B.n296 256.663
R1661 B.n424 B.n296 256.663
R1662 B.n422 B.n296 256.663
R1663 B.n415 B.n296 256.663
R1664 B.n413 B.n296 256.663
R1665 B.n407 B.n296 256.663
R1666 B.n405 B.n296 256.663
R1667 B.n399 B.n296 256.663
R1668 B.n397 B.n296 256.663
R1669 B.n391 B.n296 256.663
R1670 B.n389 B.n296 256.663
R1671 B.n383 B.n296 256.663
R1672 B.n381 B.n296 256.663
R1673 B.n375 B.n296 256.663
R1674 B.n373 B.n296 256.663
R1675 B.n367 B.n296 256.663
R1676 B.n365 B.n296 256.663
R1677 B.n359 B.n296 256.663
R1678 B.n357 B.n296 256.663
R1679 B.n351 B.n296 256.663
R1680 B.n349 B.n296 256.663
R1681 B.n344 B.n296 256.663
R1682 B.n1107 B.n1106 256.663
R1683 B.n968 B.n966 163.367
R1684 B.n964 B.n124 163.367
R1685 B.n960 B.n958 163.367
R1686 B.n956 B.n126 163.367
R1687 B.n952 B.n950 163.367
R1688 B.n948 B.n128 163.367
R1689 B.n944 B.n942 163.367
R1690 B.n940 B.n130 163.367
R1691 B.n936 B.n934 163.367
R1692 B.n932 B.n132 163.367
R1693 B.n928 B.n926 163.367
R1694 B.n924 B.n134 163.367
R1695 B.n920 B.n918 163.367
R1696 B.n916 B.n136 163.367
R1697 B.n912 B.n910 163.367
R1698 B.n908 B.n138 163.367
R1699 B.n904 B.n902 163.367
R1700 B.n900 B.n140 163.367
R1701 B.n896 B.n894 163.367
R1702 B.n891 B.n890 163.367
R1703 B.n888 B.n146 163.367
R1704 B.n884 B.n882 163.367
R1705 B.n880 B.n148 163.367
R1706 B.n875 B.n873 163.367
R1707 B.n871 B.n152 163.367
R1708 B.n867 B.n865 163.367
R1709 B.n863 B.n154 163.367
R1710 B.n859 B.n857 163.367
R1711 B.n855 B.n156 163.367
R1712 B.n851 B.n849 163.367
R1713 B.n847 B.n158 163.367
R1714 B.n843 B.n841 163.367
R1715 B.n839 B.n160 163.367
R1716 B.n835 B.n833 163.367
R1717 B.n831 B.n162 163.367
R1718 B.n827 B.n825 163.367
R1719 B.n823 B.n164 163.367
R1720 B.n819 B.n817 163.367
R1721 B.n815 B.n166 163.367
R1722 B.n811 B.n809 163.367
R1723 B.n807 B.n168 163.367
R1724 B.n803 B.n801 163.367
R1725 B.n516 B.n293 163.367
R1726 B.n520 B.n293 163.367
R1727 B.n520 B.n287 163.367
R1728 B.n528 B.n287 163.367
R1729 B.n528 B.n285 163.367
R1730 B.n532 B.n285 163.367
R1731 B.n532 B.n278 163.367
R1732 B.n540 B.n278 163.367
R1733 B.n540 B.n276 163.367
R1734 B.n544 B.n276 163.367
R1735 B.n544 B.n271 163.367
R1736 B.n552 B.n271 163.367
R1737 B.n552 B.n269 163.367
R1738 B.n556 B.n269 163.367
R1739 B.n556 B.n263 163.367
R1740 B.n564 B.n263 163.367
R1741 B.n564 B.n261 163.367
R1742 B.n568 B.n261 163.367
R1743 B.n568 B.n255 163.367
R1744 B.n576 B.n255 163.367
R1745 B.n576 B.n253 163.367
R1746 B.n580 B.n253 163.367
R1747 B.n580 B.n247 163.367
R1748 B.n588 B.n247 163.367
R1749 B.n588 B.n245 163.367
R1750 B.n592 B.n245 163.367
R1751 B.n592 B.n239 163.367
R1752 B.n600 B.n239 163.367
R1753 B.n600 B.n237 163.367
R1754 B.n604 B.n237 163.367
R1755 B.n604 B.n231 163.367
R1756 B.n612 B.n231 163.367
R1757 B.n612 B.n229 163.367
R1758 B.n616 B.n229 163.367
R1759 B.n616 B.n224 163.367
R1760 B.n625 B.n224 163.367
R1761 B.n625 B.n222 163.367
R1762 B.n629 B.n222 163.367
R1763 B.n629 B.n216 163.367
R1764 B.n637 B.n216 163.367
R1765 B.n637 B.n214 163.367
R1766 B.n641 B.n214 163.367
R1767 B.n641 B.n208 163.367
R1768 B.n649 B.n208 163.367
R1769 B.n649 B.n206 163.367
R1770 B.n653 B.n206 163.367
R1771 B.n653 B.n201 163.367
R1772 B.n662 B.n201 163.367
R1773 B.n662 B.n199 163.367
R1774 B.n666 B.n199 163.367
R1775 B.n666 B.n193 163.367
R1776 B.n674 B.n193 163.367
R1777 B.n674 B.n191 163.367
R1778 B.n678 B.n191 163.367
R1779 B.n678 B.n185 163.367
R1780 B.n686 B.n185 163.367
R1781 B.n686 B.n183 163.367
R1782 B.n690 B.n183 163.367
R1783 B.n690 B.n178 163.367
R1784 B.n699 B.n178 163.367
R1785 B.n699 B.n176 163.367
R1786 B.n704 B.n176 163.367
R1787 B.n704 B.n170 163.367
R1788 B.n712 B.n170 163.367
R1789 B.n713 B.n712 163.367
R1790 B.n713 B.n5 163.367
R1791 B.n6 B.n5 163.367
R1792 B.n7 B.n6 163.367
R1793 B.n719 B.n7 163.367
R1794 B.n720 B.n719 163.367
R1795 B.n720 B.n13 163.367
R1796 B.n14 B.n13 163.367
R1797 B.n15 B.n14 163.367
R1798 B.n725 B.n15 163.367
R1799 B.n725 B.n20 163.367
R1800 B.n21 B.n20 163.367
R1801 B.n22 B.n21 163.367
R1802 B.n730 B.n22 163.367
R1803 B.n730 B.n27 163.367
R1804 B.n28 B.n27 163.367
R1805 B.n29 B.n28 163.367
R1806 B.n735 B.n29 163.367
R1807 B.n735 B.n34 163.367
R1808 B.n35 B.n34 163.367
R1809 B.n36 B.n35 163.367
R1810 B.n740 B.n36 163.367
R1811 B.n740 B.n41 163.367
R1812 B.n42 B.n41 163.367
R1813 B.n43 B.n42 163.367
R1814 B.n745 B.n43 163.367
R1815 B.n745 B.n48 163.367
R1816 B.n49 B.n48 163.367
R1817 B.n50 B.n49 163.367
R1818 B.n750 B.n50 163.367
R1819 B.n750 B.n55 163.367
R1820 B.n56 B.n55 163.367
R1821 B.n57 B.n56 163.367
R1822 B.n755 B.n57 163.367
R1823 B.n755 B.n62 163.367
R1824 B.n63 B.n62 163.367
R1825 B.n64 B.n63 163.367
R1826 B.n760 B.n64 163.367
R1827 B.n760 B.n69 163.367
R1828 B.n70 B.n69 163.367
R1829 B.n71 B.n70 163.367
R1830 B.n765 B.n71 163.367
R1831 B.n765 B.n76 163.367
R1832 B.n77 B.n76 163.367
R1833 B.n78 B.n77 163.367
R1834 B.n770 B.n78 163.367
R1835 B.n770 B.n83 163.367
R1836 B.n84 B.n83 163.367
R1837 B.n85 B.n84 163.367
R1838 B.n775 B.n85 163.367
R1839 B.n775 B.n90 163.367
R1840 B.n91 B.n90 163.367
R1841 B.n92 B.n91 163.367
R1842 B.n780 B.n92 163.367
R1843 B.n780 B.n97 163.367
R1844 B.n98 B.n97 163.367
R1845 B.n99 B.n98 163.367
R1846 B.n785 B.n99 163.367
R1847 B.n785 B.n104 163.367
R1848 B.n105 B.n104 163.367
R1849 B.n106 B.n105 163.367
R1850 B.n790 B.n106 163.367
R1851 B.n790 B.n111 163.367
R1852 B.n112 B.n111 163.367
R1853 B.n113 B.n112 163.367
R1854 B.n795 B.n113 163.367
R1855 B.n795 B.n118 163.367
R1856 B.n119 B.n118 163.367
R1857 B.n120 B.n119 163.367
R1858 B.n510 B.n508 163.367
R1859 B.n508 B.n507 163.367
R1860 B.n504 B.n503 163.367
R1861 B.n501 B.n301 163.367
R1862 B.n497 B.n495 163.367
R1863 B.n493 B.n303 163.367
R1864 B.n489 B.n487 163.367
R1865 B.n485 B.n305 163.367
R1866 B.n481 B.n479 163.367
R1867 B.n477 B.n307 163.367
R1868 B.n473 B.n471 163.367
R1869 B.n469 B.n309 163.367
R1870 B.n465 B.n463 163.367
R1871 B.n461 B.n311 163.367
R1872 B.n457 B.n455 163.367
R1873 B.n453 B.n313 163.367
R1874 B.n449 B.n447 163.367
R1875 B.n445 B.n315 163.367
R1876 B.n441 B.n439 163.367
R1877 B.n437 B.n317 163.367
R1878 B.n433 B.n431 163.367
R1879 B.n429 B.n322 163.367
R1880 B.n425 B.n423 163.367
R1881 B.n421 B.n324 163.367
R1882 B.n416 B.n414 163.367
R1883 B.n412 B.n328 163.367
R1884 B.n408 B.n406 163.367
R1885 B.n404 B.n330 163.367
R1886 B.n400 B.n398 163.367
R1887 B.n396 B.n332 163.367
R1888 B.n392 B.n390 163.367
R1889 B.n388 B.n334 163.367
R1890 B.n384 B.n382 163.367
R1891 B.n380 B.n336 163.367
R1892 B.n376 B.n374 163.367
R1893 B.n372 B.n338 163.367
R1894 B.n368 B.n366 163.367
R1895 B.n364 B.n340 163.367
R1896 B.n360 B.n358 163.367
R1897 B.n356 B.n342 163.367
R1898 B.n352 B.n350 163.367
R1899 B.n348 B.n345 163.367
R1900 B.n514 B.n291 163.367
R1901 B.n522 B.n291 163.367
R1902 B.n522 B.n289 163.367
R1903 B.n526 B.n289 163.367
R1904 B.n526 B.n283 163.367
R1905 B.n534 B.n283 163.367
R1906 B.n534 B.n281 163.367
R1907 B.n538 B.n281 163.367
R1908 B.n538 B.n275 163.367
R1909 B.n546 B.n275 163.367
R1910 B.n546 B.n273 163.367
R1911 B.n550 B.n273 163.367
R1912 B.n550 B.n267 163.367
R1913 B.n558 B.n267 163.367
R1914 B.n558 B.n265 163.367
R1915 B.n562 B.n265 163.367
R1916 B.n562 B.n259 163.367
R1917 B.n570 B.n259 163.367
R1918 B.n570 B.n257 163.367
R1919 B.n574 B.n257 163.367
R1920 B.n574 B.n251 163.367
R1921 B.n582 B.n251 163.367
R1922 B.n582 B.n249 163.367
R1923 B.n586 B.n249 163.367
R1924 B.n586 B.n243 163.367
R1925 B.n594 B.n243 163.367
R1926 B.n594 B.n241 163.367
R1927 B.n598 B.n241 163.367
R1928 B.n598 B.n235 163.367
R1929 B.n606 B.n235 163.367
R1930 B.n606 B.n233 163.367
R1931 B.n610 B.n233 163.367
R1932 B.n610 B.n227 163.367
R1933 B.n619 B.n227 163.367
R1934 B.n619 B.n225 163.367
R1935 B.n623 B.n225 163.367
R1936 B.n623 B.n220 163.367
R1937 B.n631 B.n220 163.367
R1938 B.n631 B.n218 163.367
R1939 B.n635 B.n218 163.367
R1940 B.n635 B.n212 163.367
R1941 B.n643 B.n212 163.367
R1942 B.n643 B.n210 163.367
R1943 B.n647 B.n210 163.367
R1944 B.n647 B.n204 163.367
R1945 B.n656 B.n204 163.367
R1946 B.n656 B.n202 163.367
R1947 B.n660 B.n202 163.367
R1948 B.n660 B.n197 163.367
R1949 B.n668 B.n197 163.367
R1950 B.n668 B.n195 163.367
R1951 B.n672 B.n195 163.367
R1952 B.n672 B.n189 163.367
R1953 B.n680 B.n189 163.367
R1954 B.n680 B.n187 163.367
R1955 B.n684 B.n187 163.367
R1956 B.n684 B.n181 163.367
R1957 B.n693 B.n181 163.367
R1958 B.n693 B.n179 163.367
R1959 B.n697 B.n179 163.367
R1960 B.n697 B.n174 163.367
R1961 B.n706 B.n174 163.367
R1962 B.n706 B.n172 163.367
R1963 B.n710 B.n172 163.367
R1964 B.n710 B.n3 163.367
R1965 B.n1105 B.n3 163.367
R1966 B.n1101 B.n2 163.367
R1967 B.n1101 B.n1100 163.367
R1968 B.n1100 B.n9 163.367
R1969 B.n1096 B.n9 163.367
R1970 B.n1096 B.n11 163.367
R1971 B.n1092 B.n11 163.367
R1972 B.n1092 B.n16 163.367
R1973 B.n1088 B.n16 163.367
R1974 B.n1088 B.n18 163.367
R1975 B.n1084 B.n18 163.367
R1976 B.n1084 B.n24 163.367
R1977 B.n1080 B.n24 163.367
R1978 B.n1080 B.n26 163.367
R1979 B.n1076 B.n26 163.367
R1980 B.n1076 B.n31 163.367
R1981 B.n1072 B.n31 163.367
R1982 B.n1072 B.n33 163.367
R1983 B.n1068 B.n33 163.367
R1984 B.n1068 B.n37 163.367
R1985 B.n1064 B.n37 163.367
R1986 B.n1064 B.n39 163.367
R1987 B.n1060 B.n39 163.367
R1988 B.n1060 B.n45 163.367
R1989 B.n1056 B.n45 163.367
R1990 B.n1056 B.n47 163.367
R1991 B.n1052 B.n47 163.367
R1992 B.n1052 B.n52 163.367
R1993 B.n1048 B.n52 163.367
R1994 B.n1048 B.n54 163.367
R1995 B.n1044 B.n54 163.367
R1996 B.n1044 B.n58 163.367
R1997 B.n1040 B.n58 163.367
R1998 B.n1040 B.n60 163.367
R1999 B.n1036 B.n60 163.367
R2000 B.n1036 B.n66 163.367
R2001 B.n1032 B.n66 163.367
R2002 B.n1032 B.n68 163.367
R2003 B.n1028 B.n68 163.367
R2004 B.n1028 B.n73 163.367
R2005 B.n1024 B.n73 163.367
R2006 B.n1024 B.n75 163.367
R2007 B.n1020 B.n75 163.367
R2008 B.n1020 B.n80 163.367
R2009 B.n1016 B.n80 163.367
R2010 B.n1016 B.n82 163.367
R2011 B.n1012 B.n82 163.367
R2012 B.n1012 B.n87 163.367
R2013 B.n1008 B.n87 163.367
R2014 B.n1008 B.n89 163.367
R2015 B.n1004 B.n89 163.367
R2016 B.n1004 B.n94 163.367
R2017 B.n1000 B.n94 163.367
R2018 B.n1000 B.n96 163.367
R2019 B.n996 B.n96 163.367
R2020 B.n996 B.n101 163.367
R2021 B.n992 B.n101 163.367
R2022 B.n992 B.n103 163.367
R2023 B.n988 B.n103 163.367
R2024 B.n988 B.n108 163.367
R2025 B.n984 B.n108 163.367
R2026 B.n984 B.n110 163.367
R2027 B.n980 B.n110 163.367
R2028 B.n980 B.n115 163.367
R2029 B.n976 B.n115 163.367
R2030 B.n976 B.n117 163.367
R2031 B.n972 B.n117 163.367
R2032 B.n515 B.n296 77.7609
R2033 B.n973 B.n121 77.7609
R2034 B.n142 B.n141 76.8005
R2035 B.n150 B.n149 76.8005
R2036 B.n326 B.n325 76.8005
R2037 B.n319 B.n318 76.8005
R2038 B.n967 B.n122 71.676
R2039 B.n966 B.n965 71.676
R2040 B.n959 B.n124 71.676
R2041 B.n958 B.n957 71.676
R2042 B.n951 B.n126 71.676
R2043 B.n950 B.n949 71.676
R2044 B.n943 B.n128 71.676
R2045 B.n942 B.n941 71.676
R2046 B.n935 B.n130 71.676
R2047 B.n934 B.n933 71.676
R2048 B.n927 B.n132 71.676
R2049 B.n926 B.n925 71.676
R2050 B.n919 B.n134 71.676
R2051 B.n918 B.n917 71.676
R2052 B.n911 B.n136 71.676
R2053 B.n910 B.n909 71.676
R2054 B.n903 B.n138 71.676
R2055 B.n902 B.n901 71.676
R2056 B.n895 B.n140 71.676
R2057 B.n894 B.n144 71.676
R2058 B.n890 B.n889 71.676
R2059 B.n883 B.n146 71.676
R2060 B.n882 B.n881 71.676
R2061 B.n874 B.n148 71.676
R2062 B.n873 B.n872 71.676
R2063 B.n866 B.n152 71.676
R2064 B.n865 B.n864 71.676
R2065 B.n858 B.n154 71.676
R2066 B.n857 B.n856 71.676
R2067 B.n850 B.n156 71.676
R2068 B.n849 B.n848 71.676
R2069 B.n842 B.n158 71.676
R2070 B.n841 B.n840 71.676
R2071 B.n834 B.n160 71.676
R2072 B.n833 B.n832 71.676
R2073 B.n826 B.n162 71.676
R2074 B.n825 B.n824 71.676
R2075 B.n818 B.n164 71.676
R2076 B.n817 B.n816 71.676
R2077 B.n810 B.n166 71.676
R2078 B.n809 B.n808 71.676
R2079 B.n802 B.n168 71.676
R2080 B.n803 B.n802 71.676
R2081 B.n808 B.n807 71.676
R2082 B.n811 B.n810 71.676
R2083 B.n816 B.n815 71.676
R2084 B.n819 B.n818 71.676
R2085 B.n824 B.n823 71.676
R2086 B.n827 B.n826 71.676
R2087 B.n832 B.n831 71.676
R2088 B.n835 B.n834 71.676
R2089 B.n840 B.n839 71.676
R2090 B.n843 B.n842 71.676
R2091 B.n848 B.n847 71.676
R2092 B.n851 B.n850 71.676
R2093 B.n856 B.n855 71.676
R2094 B.n859 B.n858 71.676
R2095 B.n864 B.n863 71.676
R2096 B.n867 B.n866 71.676
R2097 B.n872 B.n871 71.676
R2098 B.n875 B.n874 71.676
R2099 B.n881 B.n880 71.676
R2100 B.n884 B.n883 71.676
R2101 B.n889 B.n888 71.676
R2102 B.n891 B.n144 71.676
R2103 B.n896 B.n895 71.676
R2104 B.n901 B.n900 71.676
R2105 B.n904 B.n903 71.676
R2106 B.n909 B.n908 71.676
R2107 B.n912 B.n911 71.676
R2108 B.n917 B.n916 71.676
R2109 B.n920 B.n919 71.676
R2110 B.n925 B.n924 71.676
R2111 B.n928 B.n927 71.676
R2112 B.n933 B.n932 71.676
R2113 B.n936 B.n935 71.676
R2114 B.n941 B.n940 71.676
R2115 B.n944 B.n943 71.676
R2116 B.n949 B.n948 71.676
R2117 B.n952 B.n951 71.676
R2118 B.n957 B.n956 71.676
R2119 B.n960 B.n959 71.676
R2120 B.n965 B.n964 71.676
R2121 B.n968 B.n967 71.676
R2122 B.n509 B.n297 71.676
R2123 B.n507 B.n299 71.676
R2124 B.n503 B.n502 71.676
R2125 B.n496 B.n301 71.676
R2126 B.n495 B.n494 71.676
R2127 B.n488 B.n303 71.676
R2128 B.n487 B.n486 71.676
R2129 B.n480 B.n305 71.676
R2130 B.n479 B.n478 71.676
R2131 B.n472 B.n307 71.676
R2132 B.n471 B.n470 71.676
R2133 B.n464 B.n309 71.676
R2134 B.n463 B.n462 71.676
R2135 B.n456 B.n311 71.676
R2136 B.n455 B.n454 71.676
R2137 B.n448 B.n313 71.676
R2138 B.n447 B.n446 71.676
R2139 B.n440 B.n315 71.676
R2140 B.n439 B.n438 71.676
R2141 B.n432 B.n317 71.676
R2142 B.n431 B.n430 71.676
R2143 B.n424 B.n322 71.676
R2144 B.n423 B.n422 71.676
R2145 B.n415 B.n324 71.676
R2146 B.n414 B.n413 71.676
R2147 B.n407 B.n328 71.676
R2148 B.n406 B.n405 71.676
R2149 B.n399 B.n330 71.676
R2150 B.n398 B.n397 71.676
R2151 B.n391 B.n332 71.676
R2152 B.n390 B.n389 71.676
R2153 B.n383 B.n334 71.676
R2154 B.n382 B.n381 71.676
R2155 B.n375 B.n336 71.676
R2156 B.n374 B.n373 71.676
R2157 B.n367 B.n338 71.676
R2158 B.n366 B.n365 71.676
R2159 B.n359 B.n340 71.676
R2160 B.n358 B.n357 71.676
R2161 B.n351 B.n342 71.676
R2162 B.n350 B.n349 71.676
R2163 B.n345 B.n344 71.676
R2164 B.n510 B.n509 71.676
R2165 B.n504 B.n299 71.676
R2166 B.n502 B.n501 71.676
R2167 B.n497 B.n496 71.676
R2168 B.n494 B.n493 71.676
R2169 B.n489 B.n488 71.676
R2170 B.n486 B.n485 71.676
R2171 B.n481 B.n480 71.676
R2172 B.n478 B.n477 71.676
R2173 B.n473 B.n472 71.676
R2174 B.n470 B.n469 71.676
R2175 B.n465 B.n464 71.676
R2176 B.n462 B.n461 71.676
R2177 B.n457 B.n456 71.676
R2178 B.n454 B.n453 71.676
R2179 B.n449 B.n448 71.676
R2180 B.n446 B.n445 71.676
R2181 B.n441 B.n440 71.676
R2182 B.n438 B.n437 71.676
R2183 B.n433 B.n432 71.676
R2184 B.n430 B.n429 71.676
R2185 B.n425 B.n424 71.676
R2186 B.n422 B.n421 71.676
R2187 B.n416 B.n415 71.676
R2188 B.n413 B.n412 71.676
R2189 B.n408 B.n407 71.676
R2190 B.n405 B.n404 71.676
R2191 B.n400 B.n399 71.676
R2192 B.n397 B.n396 71.676
R2193 B.n392 B.n391 71.676
R2194 B.n389 B.n388 71.676
R2195 B.n384 B.n383 71.676
R2196 B.n381 B.n380 71.676
R2197 B.n376 B.n375 71.676
R2198 B.n373 B.n372 71.676
R2199 B.n368 B.n367 71.676
R2200 B.n365 B.n364 71.676
R2201 B.n360 B.n359 71.676
R2202 B.n357 B.n356 71.676
R2203 B.n352 B.n351 71.676
R2204 B.n349 B.n348 71.676
R2205 B.n344 B.n295 71.676
R2206 B.n1106 B.n1105 71.676
R2207 B.n1106 B.n2 71.676
R2208 B.n143 B.n142 59.5399
R2209 B.n877 B.n150 59.5399
R2210 B.n419 B.n326 59.5399
R2211 B.n320 B.n319 59.5399
R2212 B.n515 B.n292 46.7944
R2213 B.n521 B.n292 46.7944
R2214 B.n521 B.n288 46.7944
R2215 B.n527 B.n288 46.7944
R2216 B.n527 B.n284 46.7944
R2217 B.n533 B.n284 46.7944
R2218 B.n533 B.n279 46.7944
R2219 B.n539 B.n279 46.7944
R2220 B.n539 B.n280 46.7944
R2221 B.n545 B.n272 46.7944
R2222 B.n551 B.n272 46.7944
R2223 B.n551 B.n268 46.7944
R2224 B.n557 B.n268 46.7944
R2225 B.n557 B.n264 46.7944
R2226 B.n563 B.n264 46.7944
R2227 B.n563 B.n260 46.7944
R2228 B.n569 B.n260 46.7944
R2229 B.n569 B.n256 46.7944
R2230 B.n575 B.n256 46.7944
R2231 B.n575 B.n252 46.7944
R2232 B.n581 B.n252 46.7944
R2233 B.n581 B.n248 46.7944
R2234 B.n587 B.n248 46.7944
R2235 B.n593 B.n244 46.7944
R2236 B.n593 B.n240 46.7944
R2237 B.n599 B.n240 46.7944
R2238 B.n599 B.n236 46.7944
R2239 B.n605 B.n236 46.7944
R2240 B.n605 B.n232 46.7944
R2241 B.n611 B.n232 46.7944
R2242 B.n611 B.n228 46.7944
R2243 B.n618 B.n228 46.7944
R2244 B.n618 B.n617 46.7944
R2245 B.n624 B.n221 46.7944
R2246 B.n630 B.n221 46.7944
R2247 B.n630 B.n217 46.7944
R2248 B.n636 B.n217 46.7944
R2249 B.n636 B.n213 46.7944
R2250 B.n642 B.n213 46.7944
R2251 B.n642 B.n209 46.7944
R2252 B.n648 B.n209 46.7944
R2253 B.n648 B.n205 46.7944
R2254 B.n655 B.n205 46.7944
R2255 B.n655 B.n654 46.7944
R2256 B.n661 B.n198 46.7944
R2257 B.n667 B.n198 46.7944
R2258 B.n667 B.n194 46.7944
R2259 B.n673 B.n194 46.7944
R2260 B.n673 B.n190 46.7944
R2261 B.n679 B.n190 46.7944
R2262 B.n679 B.n186 46.7944
R2263 B.n685 B.n186 46.7944
R2264 B.n685 B.n182 46.7944
R2265 B.n692 B.n182 46.7944
R2266 B.n692 B.n691 46.7944
R2267 B.n698 B.n175 46.7944
R2268 B.n705 B.n175 46.7944
R2269 B.n705 B.n171 46.7944
R2270 B.n711 B.n171 46.7944
R2271 B.n711 B.n4 46.7944
R2272 B.n1104 B.n4 46.7944
R2273 B.n1104 B.n1103 46.7944
R2274 B.n1103 B.n1102 46.7944
R2275 B.n1102 B.n8 46.7944
R2276 B.n12 B.n8 46.7944
R2277 B.n1095 B.n12 46.7944
R2278 B.n1095 B.n1094 46.7944
R2279 B.n1094 B.n1093 46.7944
R2280 B.n1087 B.n19 46.7944
R2281 B.n1087 B.n1086 46.7944
R2282 B.n1086 B.n1085 46.7944
R2283 B.n1085 B.n23 46.7944
R2284 B.n1079 B.n23 46.7944
R2285 B.n1079 B.n1078 46.7944
R2286 B.n1078 B.n1077 46.7944
R2287 B.n1077 B.n30 46.7944
R2288 B.n1071 B.n30 46.7944
R2289 B.n1071 B.n1070 46.7944
R2290 B.n1070 B.n1069 46.7944
R2291 B.n1063 B.n40 46.7944
R2292 B.n1063 B.n1062 46.7944
R2293 B.n1062 B.n1061 46.7944
R2294 B.n1061 B.n44 46.7944
R2295 B.n1055 B.n44 46.7944
R2296 B.n1055 B.n1054 46.7944
R2297 B.n1054 B.n1053 46.7944
R2298 B.n1053 B.n51 46.7944
R2299 B.n1047 B.n51 46.7944
R2300 B.n1047 B.n1046 46.7944
R2301 B.n1046 B.n1045 46.7944
R2302 B.n1039 B.n61 46.7944
R2303 B.n1039 B.n1038 46.7944
R2304 B.n1038 B.n1037 46.7944
R2305 B.n1037 B.n65 46.7944
R2306 B.n1031 B.n65 46.7944
R2307 B.n1031 B.n1030 46.7944
R2308 B.n1030 B.n1029 46.7944
R2309 B.n1029 B.n72 46.7944
R2310 B.n1023 B.n72 46.7944
R2311 B.n1023 B.n1022 46.7944
R2312 B.n1021 B.n79 46.7944
R2313 B.n1015 B.n79 46.7944
R2314 B.n1015 B.n1014 46.7944
R2315 B.n1014 B.n1013 46.7944
R2316 B.n1013 B.n86 46.7944
R2317 B.n1007 B.n86 46.7944
R2318 B.n1007 B.n1006 46.7944
R2319 B.n1006 B.n1005 46.7944
R2320 B.n1005 B.n93 46.7944
R2321 B.n999 B.n93 46.7944
R2322 B.n999 B.n998 46.7944
R2323 B.n998 B.n997 46.7944
R2324 B.n997 B.n100 46.7944
R2325 B.n991 B.n100 46.7944
R2326 B.n990 B.n989 46.7944
R2327 B.n989 B.n107 46.7944
R2328 B.n983 B.n107 46.7944
R2329 B.n983 B.n982 46.7944
R2330 B.n982 B.n981 46.7944
R2331 B.n981 B.n114 46.7944
R2332 B.n975 B.n114 46.7944
R2333 B.n975 B.n974 46.7944
R2334 B.n974 B.n973 46.7944
R2335 B.n698 B.t4 43.3536
R2336 B.n1093 B.t1 43.3536
R2337 B.t3 B.n244 40.6011
R2338 B.n1022 B.t6 40.6011
R2339 B.n617 B.t2 36.4722
R2340 B.n61 B.t5 36.4722
R2341 B.n545 B.t9 33.7196
R2342 B.n991 B.t13 33.7196
R2343 B.n513 B.n512 32.0005
R2344 B.n517 B.n294 32.0005
R2345 B.n800 B.n799 32.0005
R2346 B.n971 B.n970 32.0005
R2347 B.n661 B.t7 26.8382
R2348 B.n1069 B.t0 26.8382
R2349 B.n654 B.t7 19.9567
R2350 B.n40 B.t0 19.9567
R2351 B B.n1107 18.0485
R2352 B.n280 B.t9 13.0753
R2353 B.t13 B.n990 13.0753
R2354 B.n513 B.n290 10.6151
R2355 B.n523 B.n290 10.6151
R2356 B.n524 B.n523 10.6151
R2357 B.n525 B.n524 10.6151
R2358 B.n525 B.n282 10.6151
R2359 B.n535 B.n282 10.6151
R2360 B.n536 B.n535 10.6151
R2361 B.n537 B.n536 10.6151
R2362 B.n537 B.n274 10.6151
R2363 B.n547 B.n274 10.6151
R2364 B.n548 B.n547 10.6151
R2365 B.n549 B.n548 10.6151
R2366 B.n549 B.n266 10.6151
R2367 B.n559 B.n266 10.6151
R2368 B.n560 B.n559 10.6151
R2369 B.n561 B.n560 10.6151
R2370 B.n561 B.n258 10.6151
R2371 B.n571 B.n258 10.6151
R2372 B.n572 B.n571 10.6151
R2373 B.n573 B.n572 10.6151
R2374 B.n573 B.n250 10.6151
R2375 B.n583 B.n250 10.6151
R2376 B.n584 B.n583 10.6151
R2377 B.n585 B.n584 10.6151
R2378 B.n585 B.n242 10.6151
R2379 B.n595 B.n242 10.6151
R2380 B.n596 B.n595 10.6151
R2381 B.n597 B.n596 10.6151
R2382 B.n597 B.n234 10.6151
R2383 B.n607 B.n234 10.6151
R2384 B.n608 B.n607 10.6151
R2385 B.n609 B.n608 10.6151
R2386 B.n609 B.n226 10.6151
R2387 B.n620 B.n226 10.6151
R2388 B.n621 B.n620 10.6151
R2389 B.n622 B.n621 10.6151
R2390 B.n622 B.n219 10.6151
R2391 B.n632 B.n219 10.6151
R2392 B.n633 B.n632 10.6151
R2393 B.n634 B.n633 10.6151
R2394 B.n634 B.n211 10.6151
R2395 B.n644 B.n211 10.6151
R2396 B.n645 B.n644 10.6151
R2397 B.n646 B.n645 10.6151
R2398 B.n646 B.n203 10.6151
R2399 B.n657 B.n203 10.6151
R2400 B.n658 B.n657 10.6151
R2401 B.n659 B.n658 10.6151
R2402 B.n659 B.n196 10.6151
R2403 B.n669 B.n196 10.6151
R2404 B.n670 B.n669 10.6151
R2405 B.n671 B.n670 10.6151
R2406 B.n671 B.n188 10.6151
R2407 B.n681 B.n188 10.6151
R2408 B.n682 B.n681 10.6151
R2409 B.n683 B.n682 10.6151
R2410 B.n683 B.n180 10.6151
R2411 B.n694 B.n180 10.6151
R2412 B.n695 B.n694 10.6151
R2413 B.n696 B.n695 10.6151
R2414 B.n696 B.n173 10.6151
R2415 B.n707 B.n173 10.6151
R2416 B.n708 B.n707 10.6151
R2417 B.n709 B.n708 10.6151
R2418 B.n709 B.n0 10.6151
R2419 B.n512 B.n511 10.6151
R2420 B.n511 B.n298 10.6151
R2421 B.n506 B.n298 10.6151
R2422 B.n506 B.n505 10.6151
R2423 B.n505 B.n300 10.6151
R2424 B.n500 B.n300 10.6151
R2425 B.n500 B.n499 10.6151
R2426 B.n499 B.n498 10.6151
R2427 B.n498 B.n302 10.6151
R2428 B.n492 B.n302 10.6151
R2429 B.n492 B.n491 10.6151
R2430 B.n491 B.n490 10.6151
R2431 B.n490 B.n304 10.6151
R2432 B.n484 B.n304 10.6151
R2433 B.n484 B.n483 10.6151
R2434 B.n483 B.n482 10.6151
R2435 B.n482 B.n306 10.6151
R2436 B.n476 B.n306 10.6151
R2437 B.n476 B.n475 10.6151
R2438 B.n475 B.n474 10.6151
R2439 B.n474 B.n308 10.6151
R2440 B.n468 B.n308 10.6151
R2441 B.n468 B.n467 10.6151
R2442 B.n467 B.n466 10.6151
R2443 B.n466 B.n310 10.6151
R2444 B.n460 B.n310 10.6151
R2445 B.n460 B.n459 10.6151
R2446 B.n459 B.n458 10.6151
R2447 B.n458 B.n312 10.6151
R2448 B.n452 B.n312 10.6151
R2449 B.n452 B.n451 10.6151
R2450 B.n451 B.n450 10.6151
R2451 B.n450 B.n314 10.6151
R2452 B.n444 B.n314 10.6151
R2453 B.n444 B.n443 10.6151
R2454 B.n443 B.n442 10.6151
R2455 B.n442 B.n316 10.6151
R2456 B.n436 B.n435 10.6151
R2457 B.n435 B.n434 10.6151
R2458 B.n434 B.n321 10.6151
R2459 B.n428 B.n321 10.6151
R2460 B.n428 B.n427 10.6151
R2461 B.n427 B.n426 10.6151
R2462 B.n426 B.n323 10.6151
R2463 B.n420 B.n323 10.6151
R2464 B.n418 B.n417 10.6151
R2465 B.n417 B.n327 10.6151
R2466 B.n411 B.n327 10.6151
R2467 B.n411 B.n410 10.6151
R2468 B.n410 B.n409 10.6151
R2469 B.n409 B.n329 10.6151
R2470 B.n403 B.n329 10.6151
R2471 B.n403 B.n402 10.6151
R2472 B.n402 B.n401 10.6151
R2473 B.n401 B.n331 10.6151
R2474 B.n395 B.n331 10.6151
R2475 B.n395 B.n394 10.6151
R2476 B.n394 B.n393 10.6151
R2477 B.n393 B.n333 10.6151
R2478 B.n387 B.n333 10.6151
R2479 B.n387 B.n386 10.6151
R2480 B.n386 B.n385 10.6151
R2481 B.n385 B.n335 10.6151
R2482 B.n379 B.n335 10.6151
R2483 B.n379 B.n378 10.6151
R2484 B.n378 B.n377 10.6151
R2485 B.n377 B.n337 10.6151
R2486 B.n371 B.n337 10.6151
R2487 B.n371 B.n370 10.6151
R2488 B.n370 B.n369 10.6151
R2489 B.n369 B.n339 10.6151
R2490 B.n363 B.n339 10.6151
R2491 B.n363 B.n362 10.6151
R2492 B.n362 B.n361 10.6151
R2493 B.n361 B.n341 10.6151
R2494 B.n355 B.n341 10.6151
R2495 B.n355 B.n354 10.6151
R2496 B.n354 B.n353 10.6151
R2497 B.n353 B.n343 10.6151
R2498 B.n347 B.n343 10.6151
R2499 B.n347 B.n346 10.6151
R2500 B.n346 B.n294 10.6151
R2501 B.n518 B.n517 10.6151
R2502 B.n519 B.n518 10.6151
R2503 B.n519 B.n286 10.6151
R2504 B.n529 B.n286 10.6151
R2505 B.n530 B.n529 10.6151
R2506 B.n531 B.n530 10.6151
R2507 B.n531 B.n277 10.6151
R2508 B.n541 B.n277 10.6151
R2509 B.n542 B.n541 10.6151
R2510 B.n543 B.n542 10.6151
R2511 B.n543 B.n270 10.6151
R2512 B.n553 B.n270 10.6151
R2513 B.n554 B.n553 10.6151
R2514 B.n555 B.n554 10.6151
R2515 B.n555 B.n262 10.6151
R2516 B.n565 B.n262 10.6151
R2517 B.n566 B.n565 10.6151
R2518 B.n567 B.n566 10.6151
R2519 B.n567 B.n254 10.6151
R2520 B.n577 B.n254 10.6151
R2521 B.n578 B.n577 10.6151
R2522 B.n579 B.n578 10.6151
R2523 B.n579 B.n246 10.6151
R2524 B.n589 B.n246 10.6151
R2525 B.n590 B.n589 10.6151
R2526 B.n591 B.n590 10.6151
R2527 B.n591 B.n238 10.6151
R2528 B.n601 B.n238 10.6151
R2529 B.n602 B.n601 10.6151
R2530 B.n603 B.n602 10.6151
R2531 B.n603 B.n230 10.6151
R2532 B.n613 B.n230 10.6151
R2533 B.n614 B.n613 10.6151
R2534 B.n615 B.n614 10.6151
R2535 B.n615 B.n223 10.6151
R2536 B.n626 B.n223 10.6151
R2537 B.n627 B.n626 10.6151
R2538 B.n628 B.n627 10.6151
R2539 B.n628 B.n215 10.6151
R2540 B.n638 B.n215 10.6151
R2541 B.n639 B.n638 10.6151
R2542 B.n640 B.n639 10.6151
R2543 B.n640 B.n207 10.6151
R2544 B.n650 B.n207 10.6151
R2545 B.n651 B.n650 10.6151
R2546 B.n652 B.n651 10.6151
R2547 B.n652 B.n200 10.6151
R2548 B.n663 B.n200 10.6151
R2549 B.n664 B.n663 10.6151
R2550 B.n665 B.n664 10.6151
R2551 B.n665 B.n192 10.6151
R2552 B.n675 B.n192 10.6151
R2553 B.n676 B.n675 10.6151
R2554 B.n677 B.n676 10.6151
R2555 B.n677 B.n184 10.6151
R2556 B.n687 B.n184 10.6151
R2557 B.n688 B.n687 10.6151
R2558 B.n689 B.n688 10.6151
R2559 B.n689 B.n177 10.6151
R2560 B.n700 B.n177 10.6151
R2561 B.n701 B.n700 10.6151
R2562 B.n703 B.n701 10.6151
R2563 B.n703 B.n702 10.6151
R2564 B.n702 B.n169 10.6151
R2565 B.n714 B.n169 10.6151
R2566 B.n715 B.n714 10.6151
R2567 B.n716 B.n715 10.6151
R2568 B.n717 B.n716 10.6151
R2569 B.n718 B.n717 10.6151
R2570 B.n721 B.n718 10.6151
R2571 B.n722 B.n721 10.6151
R2572 B.n723 B.n722 10.6151
R2573 B.n724 B.n723 10.6151
R2574 B.n726 B.n724 10.6151
R2575 B.n727 B.n726 10.6151
R2576 B.n728 B.n727 10.6151
R2577 B.n729 B.n728 10.6151
R2578 B.n731 B.n729 10.6151
R2579 B.n732 B.n731 10.6151
R2580 B.n733 B.n732 10.6151
R2581 B.n734 B.n733 10.6151
R2582 B.n736 B.n734 10.6151
R2583 B.n737 B.n736 10.6151
R2584 B.n738 B.n737 10.6151
R2585 B.n739 B.n738 10.6151
R2586 B.n741 B.n739 10.6151
R2587 B.n742 B.n741 10.6151
R2588 B.n743 B.n742 10.6151
R2589 B.n744 B.n743 10.6151
R2590 B.n746 B.n744 10.6151
R2591 B.n747 B.n746 10.6151
R2592 B.n748 B.n747 10.6151
R2593 B.n749 B.n748 10.6151
R2594 B.n751 B.n749 10.6151
R2595 B.n752 B.n751 10.6151
R2596 B.n753 B.n752 10.6151
R2597 B.n754 B.n753 10.6151
R2598 B.n756 B.n754 10.6151
R2599 B.n757 B.n756 10.6151
R2600 B.n758 B.n757 10.6151
R2601 B.n759 B.n758 10.6151
R2602 B.n761 B.n759 10.6151
R2603 B.n762 B.n761 10.6151
R2604 B.n763 B.n762 10.6151
R2605 B.n764 B.n763 10.6151
R2606 B.n766 B.n764 10.6151
R2607 B.n767 B.n766 10.6151
R2608 B.n768 B.n767 10.6151
R2609 B.n769 B.n768 10.6151
R2610 B.n771 B.n769 10.6151
R2611 B.n772 B.n771 10.6151
R2612 B.n773 B.n772 10.6151
R2613 B.n774 B.n773 10.6151
R2614 B.n776 B.n774 10.6151
R2615 B.n777 B.n776 10.6151
R2616 B.n778 B.n777 10.6151
R2617 B.n779 B.n778 10.6151
R2618 B.n781 B.n779 10.6151
R2619 B.n782 B.n781 10.6151
R2620 B.n783 B.n782 10.6151
R2621 B.n784 B.n783 10.6151
R2622 B.n786 B.n784 10.6151
R2623 B.n787 B.n786 10.6151
R2624 B.n788 B.n787 10.6151
R2625 B.n789 B.n788 10.6151
R2626 B.n791 B.n789 10.6151
R2627 B.n792 B.n791 10.6151
R2628 B.n793 B.n792 10.6151
R2629 B.n794 B.n793 10.6151
R2630 B.n796 B.n794 10.6151
R2631 B.n797 B.n796 10.6151
R2632 B.n798 B.n797 10.6151
R2633 B.n799 B.n798 10.6151
R2634 B.n1099 B.n1 10.6151
R2635 B.n1099 B.n1098 10.6151
R2636 B.n1098 B.n1097 10.6151
R2637 B.n1097 B.n10 10.6151
R2638 B.n1091 B.n10 10.6151
R2639 B.n1091 B.n1090 10.6151
R2640 B.n1090 B.n1089 10.6151
R2641 B.n1089 B.n17 10.6151
R2642 B.n1083 B.n17 10.6151
R2643 B.n1083 B.n1082 10.6151
R2644 B.n1082 B.n1081 10.6151
R2645 B.n1081 B.n25 10.6151
R2646 B.n1075 B.n25 10.6151
R2647 B.n1075 B.n1074 10.6151
R2648 B.n1074 B.n1073 10.6151
R2649 B.n1073 B.n32 10.6151
R2650 B.n1067 B.n32 10.6151
R2651 B.n1067 B.n1066 10.6151
R2652 B.n1066 B.n1065 10.6151
R2653 B.n1065 B.n38 10.6151
R2654 B.n1059 B.n38 10.6151
R2655 B.n1059 B.n1058 10.6151
R2656 B.n1058 B.n1057 10.6151
R2657 B.n1057 B.n46 10.6151
R2658 B.n1051 B.n46 10.6151
R2659 B.n1051 B.n1050 10.6151
R2660 B.n1050 B.n1049 10.6151
R2661 B.n1049 B.n53 10.6151
R2662 B.n1043 B.n53 10.6151
R2663 B.n1043 B.n1042 10.6151
R2664 B.n1042 B.n1041 10.6151
R2665 B.n1041 B.n59 10.6151
R2666 B.n1035 B.n59 10.6151
R2667 B.n1035 B.n1034 10.6151
R2668 B.n1034 B.n1033 10.6151
R2669 B.n1033 B.n67 10.6151
R2670 B.n1027 B.n67 10.6151
R2671 B.n1027 B.n1026 10.6151
R2672 B.n1026 B.n1025 10.6151
R2673 B.n1025 B.n74 10.6151
R2674 B.n1019 B.n74 10.6151
R2675 B.n1019 B.n1018 10.6151
R2676 B.n1018 B.n1017 10.6151
R2677 B.n1017 B.n81 10.6151
R2678 B.n1011 B.n81 10.6151
R2679 B.n1011 B.n1010 10.6151
R2680 B.n1010 B.n1009 10.6151
R2681 B.n1009 B.n88 10.6151
R2682 B.n1003 B.n88 10.6151
R2683 B.n1003 B.n1002 10.6151
R2684 B.n1002 B.n1001 10.6151
R2685 B.n1001 B.n95 10.6151
R2686 B.n995 B.n95 10.6151
R2687 B.n995 B.n994 10.6151
R2688 B.n994 B.n993 10.6151
R2689 B.n993 B.n102 10.6151
R2690 B.n987 B.n102 10.6151
R2691 B.n987 B.n986 10.6151
R2692 B.n986 B.n985 10.6151
R2693 B.n985 B.n109 10.6151
R2694 B.n979 B.n109 10.6151
R2695 B.n979 B.n978 10.6151
R2696 B.n978 B.n977 10.6151
R2697 B.n977 B.n116 10.6151
R2698 B.n971 B.n116 10.6151
R2699 B.n970 B.n969 10.6151
R2700 B.n969 B.n123 10.6151
R2701 B.n963 B.n123 10.6151
R2702 B.n963 B.n962 10.6151
R2703 B.n962 B.n961 10.6151
R2704 B.n961 B.n125 10.6151
R2705 B.n955 B.n125 10.6151
R2706 B.n955 B.n954 10.6151
R2707 B.n954 B.n953 10.6151
R2708 B.n953 B.n127 10.6151
R2709 B.n947 B.n127 10.6151
R2710 B.n947 B.n946 10.6151
R2711 B.n946 B.n945 10.6151
R2712 B.n945 B.n129 10.6151
R2713 B.n939 B.n129 10.6151
R2714 B.n939 B.n938 10.6151
R2715 B.n938 B.n937 10.6151
R2716 B.n937 B.n131 10.6151
R2717 B.n931 B.n131 10.6151
R2718 B.n931 B.n930 10.6151
R2719 B.n930 B.n929 10.6151
R2720 B.n929 B.n133 10.6151
R2721 B.n923 B.n133 10.6151
R2722 B.n923 B.n922 10.6151
R2723 B.n922 B.n921 10.6151
R2724 B.n921 B.n135 10.6151
R2725 B.n915 B.n135 10.6151
R2726 B.n915 B.n914 10.6151
R2727 B.n914 B.n913 10.6151
R2728 B.n913 B.n137 10.6151
R2729 B.n907 B.n137 10.6151
R2730 B.n907 B.n906 10.6151
R2731 B.n906 B.n905 10.6151
R2732 B.n905 B.n139 10.6151
R2733 B.n899 B.n139 10.6151
R2734 B.n899 B.n898 10.6151
R2735 B.n898 B.n897 10.6151
R2736 B.n893 B.n892 10.6151
R2737 B.n892 B.n145 10.6151
R2738 B.n887 B.n145 10.6151
R2739 B.n887 B.n886 10.6151
R2740 B.n886 B.n885 10.6151
R2741 B.n885 B.n147 10.6151
R2742 B.n879 B.n147 10.6151
R2743 B.n879 B.n878 10.6151
R2744 B.n876 B.n151 10.6151
R2745 B.n870 B.n151 10.6151
R2746 B.n870 B.n869 10.6151
R2747 B.n869 B.n868 10.6151
R2748 B.n868 B.n153 10.6151
R2749 B.n862 B.n153 10.6151
R2750 B.n862 B.n861 10.6151
R2751 B.n861 B.n860 10.6151
R2752 B.n860 B.n155 10.6151
R2753 B.n854 B.n155 10.6151
R2754 B.n854 B.n853 10.6151
R2755 B.n853 B.n852 10.6151
R2756 B.n852 B.n157 10.6151
R2757 B.n846 B.n157 10.6151
R2758 B.n846 B.n845 10.6151
R2759 B.n845 B.n844 10.6151
R2760 B.n844 B.n159 10.6151
R2761 B.n838 B.n159 10.6151
R2762 B.n838 B.n837 10.6151
R2763 B.n837 B.n836 10.6151
R2764 B.n836 B.n161 10.6151
R2765 B.n830 B.n161 10.6151
R2766 B.n830 B.n829 10.6151
R2767 B.n829 B.n828 10.6151
R2768 B.n828 B.n163 10.6151
R2769 B.n822 B.n163 10.6151
R2770 B.n822 B.n821 10.6151
R2771 B.n821 B.n820 10.6151
R2772 B.n820 B.n165 10.6151
R2773 B.n814 B.n165 10.6151
R2774 B.n814 B.n813 10.6151
R2775 B.n813 B.n812 10.6151
R2776 B.n812 B.n167 10.6151
R2777 B.n806 B.n167 10.6151
R2778 B.n806 B.n805 10.6151
R2779 B.n805 B.n804 10.6151
R2780 B.n804 B.n800 10.6151
R2781 B.n624 B.t2 10.3227
R2782 B.n1045 B.t5 10.3227
R2783 B.n1107 B.n0 8.11757
R2784 B.n1107 B.n1 8.11757
R2785 B.n436 B.n320 6.5566
R2786 B.n420 B.n419 6.5566
R2787 B.n893 B.n143 6.5566
R2788 B.n878 B.n877 6.5566
R2789 B.n587 B.t3 6.19381
R2790 B.t6 B.n1021 6.19381
R2791 B.n320 B.n316 4.05904
R2792 B.n419 B.n418 4.05904
R2793 B.n897 B.n143 4.05904
R2794 B.n877 B.n876 4.05904
R2795 B.n691 B.t4 3.44123
R2796 B.n19 B.t1 3.44123
R2797 VN.n72 VN.n71 161.3
R2798 VN.n70 VN.n38 161.3
R2799 VN.n69 VN.n68 161.3
R2800 VN.n67 VN.n39 161.3
R2801 VN.n66 VN.n65 161.3
R2802 VN.n64 VN.n40 161.3
R2803 VN.n63 VN.n62 161.3
R2804 VN.n61 VN.n41 161.3
R2805 VN.n60 VN.n59 161.3
R2806 VN.n58 VN.n42 161.3
R2807 VN.n57 VN.n56 161.3
R2808 VN.n55 VN.n44 161.3
R2809 VN.n54 VN.n53 161.3
R2810 VN.n52 VN.n45 161.3
R2811 VN.n51 VN.n50 161.3
R2812 VN.n49 VN.n46 161.3
R2813 VN.n35 VN.n34 161.3
R2814 VN.n33 VN.n1 161.3
R2815 VN.n32 VN.n31 161.3
R2816 VN.n30 VN.n2 161.3
R2817 VN.n29 VN.n28 161.3
R2818 VN.n27 VN.n3 161.3
R2819 VN.n26 VN.n25 161.3
R2820 VN.n24 VN.n4 161.3
R2821 VN.n23 VN.n22 161.3
R2822 VN.n20 VN.n5 161.3
R2823 VN.n19 VN.n18 161.3
R2824 VN.n17 VN.n6 161.3
R2825 VN.n16 VN.n15 161.3
R2826 VN.n14 VN.n7 161.3
R2827 VN.n13 VN.n12 161.3
R2828 VN.n11 VN.n8 161.3
R2829 VN.n48 VN.t4 104.388
R2830 VN.n10 VN.t3 104.388
R2831 VN.n36 VN.n0 80.7699
R2832 VN.n73 VN.n37 80.7699
R2833 VN.n9 VN.t2 71.1055
R2834 VN.n21 VN.t6 71.1055
R2835 VN.n0 VN.t5 71.1055
R2836 VN.n47 VN.t7 71.1055
R2837 VN.n43 VN.t1 71.1055
R2838 VN.n37 VN.t0 71.1055
R2839 VN.n10 VN.n9 63.3268
R2840 VN.n48 VN.n47 63.3268
R2841 VN.n15 VN.n6 56.5193
R2842 VN.n28 VN.n2 56.5193
R2843 VN.n53 VN.n44 56.5193
R2844 VN.n65 VN.n39 56.5193
R2845 VN VN.n73 55.0132
R2846 VN.n13 VN.n8 24.4675
R2847 VN.n14 VN.n13 24.4675
R2848 VN.n15 VN.n14 24.4675
R2849 VN.n19 VN.n6 24.4675
R2850 VN.n20 VN.n19 24.4675
R2851 VN.n22 VN.n20 24.4675
R2852 VN.n26 VN.n4 24.4675
R2853 VN.n27 VN.n26 24.4675
R2854 VN.n28 VN.n27 24.4675
R2855 VN.n32 VN.n2 24.4675
R2856 VN.n33 VN.n32 24.4675
R2857 VN.n34 VN.n33 24.4675
R2858 VN.n53 VN.n52 24.4675
R2859 VN.n52 VN.n51 24.4675
R2860 VN.n51 VN.n46 24.4675
R2861 VN.n65 VN.n64 24.4675
R2862 VN.n64 VN.n63 24.4675
R2863 VN.n63 VN.n41 24.4675
R2864 VN.n59 VN.n58 24.4675
R2865 VN.n58 VN.n57 24.4675
R2866 VN.n57 VN.n44 24.4675
R2867 VN.n71 VN.n70 24.4675
R2868 VN.n70 VN.n69 24.4675
R2869 VN.n69 VN.n39 24.4675
R2870 VN.n21 VN.n4 13.2127
R2871 VN.n43 VN.n41 13.2127
R2872 VN.n9 VN.n8 11.2553
R2873 VN.n22 VN.n21 11.2553
R2874 VN.n47 VN.n46 11.2553
R2875 VN.n59 VN.n43 11.2553
R2876 VN.n34 VN.n0 9.29796
R2877 VN.n71 VN.n37 9.29796
R2878 VN.n49 VN.n48 3.17993
R2879 VN.n11 VN.n10 3.17993
R2880 VN.n73 VN.n72 0.354971
R2881 VN.n36 VN.n35 0.354971
R2882 VN VN.n36 0.26696
R2883 VN.n72 VN.n38 0.189894
R2884 VN.n68 VN.n38 0.189894
R2885 VN.n68 VN.n67 0.189894
R2886 VN.n67 VN.n66 0.189894
R2887 VN.n66 VN.n40 0.189894
R2888 VN.n62 VN.n40 0.189894
R2889 VN.n62 VN.n61 0.189894
R2890 VN.n61 VN.n60 0.189894
R2891 VN.n60 VN.n42 0.189894
R2892 VN.n56 VN.n42 0.189894
R2893 VN.n56 VN.n55 0.189894
R2894 VN.n55 VN.n54 0.189894
R2895 VN.n54 VN.n45 0.189894
R2896 VN.n50 VN.n45 0.189894
R2897 VN.n50 VN.n49 0.189894
R2898 VN.n12 VN.n11 0.189894
R2899 VN.n12 VN.n7 0.189894
R2900 VN.n16 VN.n7 0.189894
R2901 VN.n17 VN.n16 0.189894
R2902 VN.n18 VN.n17 0.189894
R2903 VN.n18 VN.n5 0.189894
R2904 VN.n23 VN.n5 0.189894
R2905 VN.n24 VN.n23 0.189894
R2906 VN.n25 VN.n24 0.189894
R2907 VN.n25 VN.n3 0.189894
R2908 VN.n29 VN.n3 0.189894
R2909 VN.n30 VN.n29 0.189894
R2910 VN.n31 VN.n30 0.189894
R2911 VN.n31 VN.n1 0.189894
R2912 VN.n35 VN.n1 0.189894
R2913 VDD2.n2 VDD2.n1 64.5735
R2914 VDD2.n2 VDD2.n0 64.5735
R2915 VDD2 VDD2.n5 64.5706
R2916 VDD2.n4 VDD2.n3 62.9221
R2917 VDD2.n4 VDD2.n2 48.3101
R2918 VDD2.n5 VDD2.t0 1.84924
R2919 VDD2.n5 VDD2.t3 1.84924
R2920 VDD2.n3 VDD2.t7 1.84924
R2921 VDD2.n3 VDD2.t6 1.84924
R2922 VDD2.n1 VDD2.t1 1.84924
R2923 VDD2.n1 VDD2.t2 1.84924
R2924 VDD2.n0 VDD2.t4 1.84924
R2925 VDD2.n0 VDD2.t5 1.84924
R2926 VDD2 VDD2.n4 1.76559
C0 VDD1 VDD2 2.31257f
C1 VDD2 VN 8.254709f
C2 VDD2 VTAIL 8.19853f
C3 VDD1 VN 0.153732f
C4 VDD1 VTAIL 8.13721f
C5 VN VTAIL 9.058701f
C6 VDD2 VP 0.629416f
C7 VDD1 VP 8.72848f
C8 VP VN 8.68282f
C9 VP VTAIL 9.072809f
C10 VDD2 B 6.3502f
C11 VDD1 B 6.89554f
C12 VTAIL B 10.40319f
C13 VN B 19.38489f
C14 VP B 18.045153f
C15 VDD2.t4 B 0.232488f
C16 VDD2.t5 B 0.232488f
C17 VDD2.n0 B 2.07477f
C18 VDD2.t1 B 0.232488f
C19 VDD2.t2 B 0.232488f
C20 VDD2.n1 B 2.07477f
C21 VDD2.n2 B 4.16442f
C22 VDD2.t7 B 0.232488f
C23 VDD2.t6 B 0.232488f
C24 VDD2.n3 B 2.05727f
C25 VDD2.n4 B 3.52548f
C26 VDD2.t0 B 0.232488f
C27 VDD2.t3 B 0.232488f
C28 VDD2.n5 B 2.07472f
C29 VN.t5 B 1.92718f
C30 VN.n0 B 0.751917f
C31 VN.n1 B 0.018257f
C32 VN.n2 B 0.028686f
C33 VN.n3 B 0.018257f
C34 VN.n4 B 0.026298f
C35 VN.n5 B 0.018257f
C36 VN.n6 B 0.026651f
C37 VN.n7 B 0.018257f
C38 VN.n8 B 0.024954f
C39 VN.t2 B 1.92718f
C40 VN.n9 B 0.742795f
C41 VN.t3 B 2.18842f
C42 VN.n10 B 0.703913f
C43 VN.n11 B 0.228665f
C44 VN.n12 B 0.018257f
C45 VN.n13 B 0.034026f
C46 VN.n14 B 0.034026f
C47 VN.n15 B 0.026651f
C48 VN.n16 B 0.018257f
C49 VN.n17 B 0.018257f
C50 VN.n18 B 0.018257f
C51 VN.n19 B 0.034026f
C52 VN.n20 B 0.034026f
C53 VN.t6 B 1.92718f
C54 VN.n21 B 0.679828f
C55 VN.n22 B 0.024954f
C56 VN.n23 B 0.018257f
C57 VN.n24 B 0.018257f
C58 VN.n25 B 0.018257f
C59 VN.n26 B 0.034026f
C60 VN.n27 B 0.034026f
C61 VN.n28 B 0.024616f
C62 VN.n29 B 0.018257f
C63 VN.n30 B 0.018257f
C64 VN.n31 B 0.018257f
C65 VN.n32 B 0.034026f
C66 VN.n33 B 0.034026f
C67 VN.n34 B 0.02361f
C68 VN.n35 B 0.029466f
C69 VN.n36 B 0.050629f
C70 VN.t0 B 1.92718f
C71 VN.n37 B 0.751917f
C72 VN.n38 B 0.018257f
C73 VN.n39 B 0.028686f
C74 VN.n40 B 0.018257f
C75 VN.n41 B 0.026298f
C76 VN.n42 B 0.018257f
C77 VN.t1 B 1.92718f
C78 VN.n43 B 0.679828f
C79 VN.n44 B 0.026651f
C80 VN.n45 B 0.018257f
C81 VN.n46 B 0.024954f
C82 VN.t4 B 2.18842f
C83 VN.t7 B 1.92718f
C84 VN.n47 B 0.742795f
C85 VN.n48 B 0.703913f
C86 VN.n49 B 0.228665f
C87 VN.n50 B 0.018257f
C88 VN.n51 B 0.034026f
C89 VN.n52 B 0.034026f
C90 VN.n53 B 0.026651f
C91 VN.n54 B 0.018257f
C92 VN.n55 B 0.018257f
C93 VN.n56 B 0.018257f
C94 VN.n57 B 0.034026f
C95 VN.n58 B 0.034026f
C96 VN.n59 B 0.024954f
C97 VN.n60 B 0.018257f
C98 VN.n61 B 0.018257f
C99 VN.n62 B 0.018257f
C100 VN.n63 B 0.034026f
C101 VN.n64 B 0.034026f
C102 VN.n65 B 0.024616f
C103 VN.n66 B 0.018257f
C104 VN.n67 B 0.018257f
C105 VN.n68 B 0.018257f
C106 VN.n69 B 0.034026f
C107 VN.n70 B 0.034026f
C108 VN.n71 B 0.02361f
C109 VN.n72 B 0.029466f
C110 VN.n73 B 1.19766f
C111 VDD1.t0 B 0.23493f
C112 VDD1.t4 B 0.23493f
C113 VDD1.n0 B 2.09802f
C114 VDD1.t3 B 0.23493f
C115 VDD1.t2 B 0.23493f
C116 VDD1.n1 B 2.09656f
C117 VDD1.t1 B 0.23493f
C118 VDD1.t6 B 0.23493f
C119 VDD1.n2 B 2.09656f
C120 VDD1.n3 B 4.26544f
C121 VDD1.t5 B 0.23493f
C122 VDD1.t7 B 0.23493f
C123 VDD1.n4 B 2.07887f
C124 VDD1.n5 B 3.59737f
C125 VTAIL.t0 B 0.178876f
C126 VTAIL.t5 B 0.178876f
C127 VTAIL.n0 B 1.52192f
C128 VTAIL.n1 B 0.441615f
C129 VTAIL.n2 B 0.028995f
C130 VTAIL.n3 B 0.021135f
C131 VTAIL.n4 B 0.011357f
C132 VTAIL.n5 B 0.026844f
C133 VTAIL.n6 B 0.012025f
C134 VTAIL.n7 B 0.021135f
C135 VTAIL.n8 B 0.011357f
C136 VTAIL.n9 B 0.026844f
C137 VTAIL.n10 B 0.012025f
C138 VTAIL.n11 B 0.021135f
C139 VTAIL.n12 B 0.011357f
C140 VTAIL.n13 B 0.026844f
C141 VTAIL.n14 B 0.012025f
C142 VTAIL.n15 B 0.021135f
C143 VTAIL.n16 B 0.011357f
C144 VTAIL.n17 B 0.026844f
C145 VTAIL.n18 B 0.012025f
C146 VTAIL.n19 B 0.141917f
C147 VTAIL.t1 B 0.045192f
C148 VTAIL.n20 B 0.020133f
C149 VTAIL.n21 B 0.018977f
C150 VTAIL.n22 B 0.011357f
C151 VTAIL.n23 B 0.944969f
C152 VTAIL.n24 B 0.021135f
C153 VTAIL.n25 B 0.011357f
C154 VTAIL.n26 B 0.012025f
C155 VTAIL.n27 B 0.026844f
C156 VTAIL.n28 B 0.026844f
C157 VTAIL.n29 B 0.012025f
C158 VTAIL.n30 B 0.011357f
C159 VTAIL.n31 B 0.021135f
C160 VTAIL.n32 B 0.021135f
C161 VTAIL.n33 B 0.011357f
C162 VTAIL.n34 B 0.012025f
C163 VTAIL.n35 B 0.026844f
C164 VTAIL.n36 B 0.026844f
C165 VTAIL.n37 B 0.026844f
C166 VTAIL.n38 B 0.012025f
C167 VTAIL.n39 B 0.011357f
C168 VTAIL.n40 B 0.021135f
C169 VTAIL.n41 B 0.021135f
C170 VTAIL.n42 B 0.011357f
C171 VTAIL.n43 B 0.011691f
C172 VTAIL.n44 B 0.011691f
C173 VTAIL.n45 B 0.026844f
C174 VTAIL.n46 B 0.026844f
C175 VTAIL.n47 B 0.012025f
C176 VTAIL.n48 B 0.011357f
C177 VTAIL.n49 B 0.021135f
C178 VTAIL.n50 B 0.021135f
C179 VTAIL.n51 B 0.011357f
C180 VTAIL.n52 B 0.012025f
C181 VTAIL.n53 B 0.026844f
C182 VTAIL.n54 B 0.056853f
C183 VTAIL.n55 B 0.012025f
C184 VTAIL.n56 B 0.011357f
C185 VTAIL.n57 B 0.04972f
C186 VTAIL.n58 B 0.031708f
C187 VTAIL.n59 B 0.283025f
C188 VTAIL.n60 B 0.028995f
C189 VTAIL.n61 B 0.021135f
C190 VTAIL.n62 B 0.011357f
C191 VTAIL.n63 B 0.026844f
C192 VTAIL.n64 B 0.012025f
C193 VTAIL.n65 B 0.021135f
C194 VTAIL.n66 B 0.011357f
C195 VTAIL.n67 B 0.026844f
C196 VTAIL.n68 B 0.012025f
C197 VTAIL.n69 B 0.021135f
C198 VTAIL.n70 B 0.011357f
C199 VTAIL.n71 B 0.026844f
C200 VTAIL.n72 B 0.012025f
C201 VTAIL.n73 B 0.021135f
C202 VTAIL.n74 B 0.011357f
C203 VTAIL.n75 B 0.026844f
C204 VTAIL.n76 B 0.012025f
C205 VTAIL.n77 B 0.141917f
C206 VTAIL.t15 B 0.045192f
C207 VTAIL.n78 B 0.020133f
C208 VTAIL.n79 B 0.018977f
C209 VTAIL.n80 B 0.011357f
C210 VTAIL.n81 B 0.944969f
C211 VTAIL.n82 B 0.021135f
C212 VTAIL.n83 B 0.011357f
C213 VTAIL.n84 B 0.012025f
C214 VTAIL.n85 B 0.026844f
C215 VTAIL.n86 B 0.026844f
C216 VTAIL.n87 B 0.012025f
C217 VTAIL.n88 B 0.011357f
C218 VTAIL.n89 B 0.021135f
C219 VTAIL.n90 B 0.021135f
C220 VTAIL.n91 B 0.011357f
C221 VTAIL.n92 B 0.012025f
C222 VTAIL.n93 B 0.026844f
C223 VTAIL.n94 B 0.026844f
C224 VTAIL.n95 B 0.026844f
C225 VTAIL.n96 B 0.012025f
C226 VTAIL.n97 B 0.011357f
C227 VTAIL.n98 B 0.021135f
C228 VTAIL.n99 B 0.021135f
C229 VTAIL.n100 B 0.011357f
C230 VTAIL.n101 B 0.011691f
C231 VTAIL.n102 B 0.011691f
C232 VTAIL.n103 B 0.026844f
C233 VTAIL.n104 B 0.026844f
C234 VTAIL.n105 B 0.012025f
C235 VTAIL.n106 B 0.011357f
C236 VTAIL.n107 B 0.021135f
C237 VTAIL.n108 B 0.021135f
C238 VTAIL.n109 B 0.011357f
C239 VTAIL.n110 B 0.012025f
C240 VTAIL.n111 B 0.026844f
C241 VTAIL.n112 B 0.056853f
C242 VTAIL.n113 B 0.012025f
C243 VTAIL.n114 B 0.011357f
C244 VTAIL.n115 B 0.04972f
C245 VTAIL.n116 B 0.031708f
C246 VTAIL.n117 B 0.283025f
C247 VTAIL.t13 B 0.178876f
C248 VTAIL.t12 B 0.178876f
C249 VTAIL.n118 B 1.52192f
C250 VTAIL.n119 B 0.67014f
C251 VTAIL.n120 B 0.028995f
C252 VTAIL.n121 B 0.021135f
C253 VTAIL.n122 B 0.011357f
C254 VTAIL.n123 B 0.026844f
C255 VTAIL.n124 B 0.012025f
C256 VTAIL.n125 B 0.021135f
C257 VTAIL.n126 B 0.011357f
C258 VTAIL.n127 B 0.026844f
C259 VTAIL.n128 B 0.012025f
C260 VTAIL.n129 B 0.021135f
C261 VTAIL.n130 B 0.011357f
C262 VTAIL.n131 B 0.026844f
C263 VTAIL.n132 B 0.012025f
C264 VTAIL.n133 B 0.021135f
C265 VTAIL.n134 B 0.011357f
C266 VTAIL.n135 B 0.026844f
C267 VTAIL.n136 B 0.012025f
C268 VTAIL.n137 B 0.141917f
C269 VTAIL.t10 B 0.045192f
C270 VTAIL.n138 B 0.020133f
C271 VTAIL.n139 B 0.018977f
C272 VTAIL.n140 B 0.011357f
C273 VTAIL.n141 B 0.944969f
C274 VTAIL.n142 B 0.021135f
C275 VTAIL.n143 B 0.011357f
C276 VTAIL.n144 B 0.012025f
C277 VTAIL.n145 B 0.026844f
C278 VTAIL.n146 B 0.026844f
C279 VTAIL.n147 B 0.012025f
C280 VTAIL.n148 B 0.011357f
C281 VTAIL.n149 B 0.021135f
C282 VTAIL.n150 B 0.021135f
C283 VTAIL.n151 B 0.011357f
C284 VTAIL.n152 B 0.012025f
C285 VTAIL.n153 B 0.026844f
C286 VTAIL.n154 B 0.026844f
C287 VTAIL.n155 B 0.026844f
C288 VTAIL.n156 B 0.012025f
C289 VTAIL.n157 B 0.011357f
C290 VTAIL.n158 B 0.021135f
C291 VTAIL.n159 B 0.021135f
C292 VTAIL.n160 B 0.011357f
C293 VTAIL.n161 B 0.011691f
C294 VTAIL.n162 B 0.011691f
C295 VTAIL.n163 B 0.026844f
C296 VTAIL.n164 B 0.026844f
C297 VTAIL.n165 B 0.012025f
C298 VTAIL.n166 B 0.011357f
C299 VTAIL.n167 B 0.021135f
C300 VTAIL.n168 B 0.021135f
C301 VTAIL.n169 B 0.011357f
C302 VTAIL.n170 B 0.012025f
C303 VTAIL.n171 B 0.026844f
C304 VTAIL.n172 B 0.056853f
C305 VTAIL.n173 B 0.012025f
C306 VTAIL.n174 B 0.011357f
C307 VTAIL.n175 B 0.04972f
C308 VTAIL.n176 B 0.031708f
C309 VTAIL.n177 B 1.39939f
C310 VTAIL.n178 B 0.028995f
C311 VTAIL.n179 B 0.021135f
C312 VTAIL.n180 B 0.011357f
C313 VTAIL.n181 B 0.026844f
C314 VTAIL.n182 B 0.012025f
C315 VTAIL.n183 B 0.021135f
C316 VTAIL.n184 B 0.011357f
C317 VTAIL.n185 B 0.026844f
C318 VTAIL.n186 B 0.012025f
C319 VTAIL.n187 B 0.021135f
C320 VTAIL.n188 B 0.011357f
C321 VTAIL.n189 B 0.026844f
C322 VTAIL.n190 B 0.026844f
C323 VTAIL.n191 B 0.012025f
C324 VTAIL.n192 B 0.021135f
C325 VTAIL.n193 B 0.011357f
C326 VTAIL.n194 B 0.026844f
C327 VTAIL.n195 B 0.012025f
C328 VTAIL.n196 B 0.141917f
C329 VTAIL.t3 B 0.045192f
C330 VTAIL.n197 B 0.020133f
C331 VTAIL.n198 B 0.018977f
C332 VTAIL.n199 B 0.011357f
C333 VTAIL.n200 B 0.944969f
C334 VTAIL.n201 B 0.021135f
C335 VTAIL.n202 B 0.011357f
C336 VTAIL.n203 B 0.012025f
C337 VTAIL.n204 B 0.026844f
C338 VTAIL.n205 B 0.026844f
C339 VTAIL.n206 B 0.012025f
C340 VTAIL.n207 B 0.011357f
C341 VTAIL.n208 B 0.021135f
C342 VTAIL.n209 B 0.021135f
C343 VTAIL.n210 B 0.011357f
C344 VTAIL.n211 B 0.012025f
C345 VTAIL.n212 B 0.026844f
C346 VTAIL.n213 B 0.026844f
C347 VTAIL.n214 B 0.012025f
C348 VTAIL.n215 B 0.011357f
C349 VTAIL.n216 B 0.021135f
C350 VTAIL.n217 B 0.021135f
C351 VTAIL.n218 B 0.011357f
C352 VTAIL.n219 B 0.011691f
C353 VTAIL.n220 B 0.011691f
C354 VTAIL.n221 B 0.026844f
C355 VTAIL.n222 B 0.026844f
C356 VTAIL.n223 B 0.012025f
C357 VTAIL.n224 B 0.011357f
C358 VTAIL.n225 B 0.021135f
C359 VTAIL.n226 B 0.021135f
C360 VTAIL.n227 B 0.011357f
C361 VTAIL.n228 B 0.012025f
C362 VTAIL.n229 B 0.026844f
C363 VTAIL.n230 B 0.056853f
C364 VTAIL.n231 B 0.012025f
C365 VTAIL.n232 B 0.011357f
C366 VTAIL.n233 B 0.04972f
C367 VTAIL.n234 B 0.031708f
C368 VTAIL.n235 B 1.39939f
C369 VTAIL.t2 B 0.178876f
C370 VTAIL.t7 B 0.178876f
C371 VTAIL.n236 B 1.52193f
C372 VTAIL.n237 B 0.670131f
C373 VTAIL.n238 B 0.028995f
C374 VTAIL.n239 B 0.021135f
C375 VTAIL.n240 B 0.011357f
C376 VTAIL.n241 B 0.026844f
C377 VTAIL.n242 B 0.012025f
C378 VTAIL.n243 B 0.021135f
C379 VTAIL.n244 B 0.011357f
C380 VTAIL.n245 B 0.026844f
C381 VTAIL.n246 B 0.012025f
C382 VTAIL.n247 B 0.021135f
C383 VTAIL.n248 B 0.011357f
C384 VTAIL.n249 B 0.026844f
C385 VTAIL.n250 B 0.026844f
C386 VTAIL.n251 B 0.012025f
C387 VTAIL.n252 B 0.021135f
C388 VTAIL.n253 B 0.011357f
C389 VTAIL.n254 B 0.026844f
C390 VTAIL.n255 B 0.012025f
C391 VTAIL.n256 B 0.141917f
C392 VTAIL.t4 B 0.045192f
C393 VTAIL.n257 B 0.020133f
C394 VTAIL.n258 B 0.018977f
C395 VTAIL.n259 B 0.011357f
C396 VTAIL.n260 B 0.944969f
C397 VTAIL.n261 B 0.021135f
C398 VTAIL.n262 B 0.011357f
C399 VTAIL.n263 B 0.012025f
C400 VTAIL.n264 B 0.026844f
C401 VTAIL.n265 B 0.026844f
C402 VTAIL.n266 B 0.012025f
C403 VTAIL.n267 B 0.011357f
C404 VTAIL.n268 B 0.021135f
C405 VTAIL.n269 B 0.021135f
C406 VTAIL.n270 B 0.011357f
C407 VTAIL.n271 B 0.012025f
C408 VTAIL.n272 B 0.026844f
C409 VTAIL.n273 B 0.026844f
C410 VTAIL.n274 B 0.012025f
C411 VTAIL.n275 B 0.011357f
C412 VTAIL.n276 B 0.021135f
C413 VTAIL.n277 B 0.021135f
C414 VTAIL.n278 B 0.011357f
C415 VTAIL.n279 B 0.011691f
C416 VTAIL.n280 B 0.011691f
C417 VTAIL.n281 B 0.026844f
C418 VTAIL.n282 B 0.026844f
C419 VTAIL.n283 B 0.012025f
C420 VTAIL.n284 B 0.011357f
C421 VTAIL.n285 B 0.021135f
C422 VTAIL.n286 B 0.021135f
C423 VTAIL.n287 B 0.011357f
C424 VTAIL.n288 B 0.012025f
C425 VTAIL.n289 B 0.026844f
C426 VTAIL.n290 B 0.056853f
C427 VTAIL.n291 B 0.012025f
C428 VTAIL.n292 B 0.011357f
C429 VTAIL.n293 B 0.04972f
C430 VTAIL.n294 B 0.031708f
C431 VTAIL.n295 B 0.283025f
C432 VTAIL.n296 B 0.028995f
C433 VTAIL.n297 B 0.021135f
C434 VTAIL.n298 B 0.011357f
C435 VTAIL.n299 B 0.026844f
C436 VTAIL.n300 B 0.012025f
C437 VTAIL.n301 B 0.021135f
C438 VTAIL.n302 B 0.011357f
C439 VTAIL.n303 B 0.026844f
C440 VTAIL.n304 B 0.012025f
C441 VTAIL.n305 B 0.021135f
C442 VTAIL.n306 B 0.011357f
C443 VTAIL.n307 B 0.026844f
C444 VTAIL.n308 B 0.026844f
C445 VTAIL.n309 B 0.012025f
C446 VTAIL.n310 B 0.021135f
C447 VTAIL.n311 B 0.011357f
C448 VTAIL.n312 B 0.026844f
C449 VTAIL.n313 B 0.012025f
C450 VTAIL.n314 B 0.141917f
C451 VTAIL.t8 B 0.045192f
C452 VTAIL.n315 B 0.020133f
C453 VTAIL.n316 B 0.018977f
C454 VTAIL.n317 B 0.011357f
C455 VTAIL.n318 B 0.944969f
C456 VTAIL.n319 B 0.021135f
C457 VTAIL.n320 B 0.011357f
C458 VTAIL.n321 B 0.012025f
C459 VTAIL.n322 B 0.026844f
C460 VTAIL.n323 B 0.026844f
C461 VTAIL.n324 B 0.012025f
C462 VTAIL.n325 B 0.011357f
C463 VTAIL.n326 B 0.021135f
C464 VTAIL.n327 B 0.021135f
C465 VTAIL.n328 B 0.011357f
C466 VTAIL.n329 B 0.012025f
C467 VTAIL.n330 B 0.026844f
C468 VTAIL.n331 B 0.026844f
C469 VTAIL.n332 B 0.012025f
C470 VTAIL.n333 B 0.011357f
C471 VTAIL.n334 B 0.021135f
C472 VTAIL.n335 B 0.021135f
C473 VTAIL.n336 B 0.011357f
C474 VTAIL.n337 B 0.011691f
C475 VTAIL.n338 B 0.011691f
C476 VTAIL.n339 B 0.026844f
C477 VTAIL.n340 B 0.026844f
C478 VTAIL.n341 B 0.012025f
C479 VTAIL.n342 B 0.011357f
C480 VTAIL.n343 B 0.021135f
C481 VTAIL.n344 B 0.021135f
C482 VTAIL.n345 B 0.011357f
C483 VTAIL.n346 B 0.012025f
C484 VTAIL.n347 B 0.026844f
C485 VTAIL.n348 B 0.056853f
C486 VTAIL.n349 B 0.012025f
C487 VTAIL.n350 B 0.011357f
C488 VTAIL.n351 B 0.04972f
C489 VTAIL.n352 B 0.031708f
C490 VTAIL.n353 B 0.283025f
C491 VTAIL.t11 B 0.178876f
C492 VTAIL.t9 B 0.178876f
C493 VTAIL.n354 B 1.52193f
C494 VTAIL.n355 B 0.670131f
C495 VTAIL.n356 B 0.028995f
C496 VTAIL.n357 B 0.021135f
C497 VTAIL.n358 B 0.011357f
C498 VTAIL.n359 B 0.026844f
C499 VTAIL.n360 B 0.012025f
C500 VTAIL.n361 B 0.021135f
C501 VTAIL.n362 B 0.011357f
C502 VTAIL.n363 B 0.026844f
C503 VTAIL.n364 B 0.012025f
C504 VTAIL.n365 B 0.021135f
C505 VTAIL.n366 B 0.011357f
C506 VTAIL.n367 B 0.026844f
C507 VTAIL.n368 B 0.026844f
C508 VTAIL.n369 B 0.012025f
C509 VTAIL.n370 B 0.021135f
C510 VTAIL.n371 B 0.011357f
C511 VTAIL.n372 B 0.026844f
C512 VTAIL.n373 B 0.012025f
C513 VTAIL.n374 B 0.141917f
C514 VTAIL.t14 B 0.045192f
C515 VTAIL.n375 B 0.020133f
C516 VTAIL.n376 B 0.018977f
C517 VTAIL.n377 B 0.011357f
C518 VTAIL.n378 B 0.944969f
C519 VTAIL.n379 B 0.021135f
C520 VTAIL.n380 B 0.011357f
C521 VTAIL.n381 B 0.012025f
C522 VTAIL.n382 B 0.026844f
C523 VTAIL.n383 B 0.026844f
C524 VTAIL.n384 B 0.012025f
C525 VTAIL.n385 B 0.011357f
C526 VTAIL.n386 B 0.021135f
C527 VTAIL.n387 B 0.021135f
C528 VTAIL.n388 B 0.011357f
C529 VTAIL.n389 B 0.012025f
C530 VTAIL.n390 B 0.026844f
C531 VTAIL.n391 B 0.026844f
C532 VTAIL.n392 B 0.012025f
C533 VTAIL.n393 B 0.011357f
C534 VTAIL.n394 B 0.021135f
C535 VTAIL.n395 B 0.021135f
C536 VTAIL.n396 B 0.011357f
C537 VTAIL.n397 B 0.011691f
C538 VTAIL.n398 B 0.011691f
C539 VTAIL.n399 B 0.026844f
C540 VTAIL.n400 B 0.026844f
C541 VTAIL.n401 B 0.012025f
C542 VTAIL.n402 B 0.011357f
C543 VTAIL.n403 B 0.021135f
C544 VTAIL.n404 B 0.021135f
C545 VTAIL.n405 B 0.011357f
C546 VTAIL.n406 B 0.012025f
C547 VTAIL.n407 B 0.026844f
C548 VTAIL.n408 B 0.056853f
C549 VTAIL.n409 B 0.012025f
C550 VTAIL.n410 B 0.011357f
C551 VTAIL.n411 B 0.04972f
C552 VTAIL.n412 B 0.031708f
C553 VTAIL.n413 B 1.39939f
C554 VTAIL.n414 B 0.028995f
C555 VTAIL.n415 B 0.021135f
C556 VTAIL.n416 B 0.011357f
C557 VTAIL.n417 B 0.026844f
C558 VTAIL.n418 B 0.012025f
C559 VTAIL.n419 B 0.021135f
C560 VTAIL.n420 B 0.011357f
C561 VTAIL.n421 B 0.026844f
C562 VTAIL.n422 B 0.012025f
C563 VTAIL.n423 B 0.021135f
C564 VTAIL.n424 B 0.011357f
C565 VTAIL.n425 B 0.026844f
C566 VTAIL.n426 B 0.012025f
C567 VTAIL.n427 B 0.021135f
C568 VTAIL.n428 B 0.011357f
C569 VTAIL.n429 B 0.026844f
C570 VTAIL.n430 B 0.012025f
C571 VTAIL.n431 B 0.141917f
C572 VTAIL.t6 B 0.045192f
C573 VTAIL.n432 B 0.020133f
C574 VTAIL.n433 B 0.018977f
C575 VTAIL.n434 B 0.011357f
C576 VTAIL.n435 B 0.944969f
C577 VTAIL.n436 B 0.021135f
C578 VTAIL.n437 B 0.011357f
C579 VTAIL.n438 B 0.012025f
C580 VTAIL.n439 B 0.026844f
C581 VTAIL.n440 B 0.026844f
C582 VTAIL.n441 B 0.012025f
C583 VTAIL.n442 B 0.011357f
C584 VTAIL.n443 B 0.021135f
C585 VTAIL.n444 B 0.021135f
C586 VTAIL.n445 B 0.011357f
C587 VTAIL.n446 B 0.012025f
C588 VTAIL.n447 B 0.026844f
C589 VTAIL.n448 B 0.026844f
C590 VTAIL.n449 B 0.026844f
C591 VTAIL.n450 B 0.012025f
C592 VTAIL.n451 B 0.011357f
C593 VTAIL.n452 B 0.021135f
C594 VTAIL.n453 B 0.021135f
C595 VTAIL.n454 B 0.011357f
C596 VTAIL.n455 B 0.011691f
C597 VTAIL.n456 B 0.011691f
C598 VTAIL.n457 B 0.026844f
C599 VTAIL.n458 B 0.026844f
C600 VTAIL.n459 B 0.012025f
C601 VTAIL.n460 B 0.011357f
C602 VTAIL.n461 B 0.021135f
C603 VTAIL.n462 B 0.021135f
C604 VTAIL.n463 B 0.011357f
C605 VTAIL.n464 B 0.012025f
C606 VTAIL.n465 B 0.026844f
C607 VTAIL.n466 B 0.056853f
C608 VTAIL.n467 B 0.012025f
C609 VTAIL.n468 B 0.011357f
C610 VTAIL.n469 B 0.04972f
C611 VTAIL.n470 B 0.031708f
C612 VTAIL.n471 B 1.39543f
C613 VP.t1 B 1.95864f
C614 VP.n0 B 0.764192f
C615 VP.n1 B 0.018554f
C616 VP.n2 B 0.029154f
C617 VP.n3 B 0.018554f
C618 VP.n4 B 0.026728f
C619 VP.n5 B 0.018554f
C620 VP.n6 B 0.027086f
C621 VP.n7 B 0.018554f
C622 VP.n8 B 0.025362f
C623 VP.n9 B 0.018554f
C624 VP.n10 B 0.025018f
C625 VP.n11 B 0.018554f
C626 VP.n12 B 0.023996f
C627 VP.t0 B 1.95864f
C628 VP.n13 B 0.764192f
C629 VP.n14 B 0.018554f
C630 VP.n15 B 0.029154f
C631 VP.n16 B 0.018554f
C632 VP.n17 B 0.026728f
C633 VP.n18 B 0.018554f
C634 VP.n19 B 0.027086f
C635 VP.n20 B 0.018554f
C636 VP.n21 B 0.025362f
C637 VP.t7 B 2.22415f
C638 VP.t3 B 1.95864f
C639 VP.n22 B 0.754921f
C640 VP.n23 B 0.715405f
C641 VP.n24 B 0.232398f
C642 VP.n25 B 0.018554f
C643 VP.n26 B 0.034581f
C644 VP.n27 B 0.034581f
C645 VP.n28 B 0.027086f
C646 VP.n29 B 0.018554f
C647 VP.n30 B 0.018554f
C648 VP.n31 B 0.018554f
C649 VP.n32 B 0.034581f
C650 VP.n33 B 0.034581f
C651 VP.t2 B 1.95864f
C652 VP.n34 B 0.690926f
C653 VP.n35 B 0.025362f
C654 VP.n36 B 0.018554f
C655 VP.n37 B 0.018554f
C656 VP.n38 B 0.018554f
C657 VP.n39 B 0.034581f
C658 VP.n40 B 0.034581f
C659 VP.n41 B 0.025018f
C660 VP.n42 B 0.018554f
C661 VP.n43 B 0.018554f
C662 VP.n44 B 0.018554f
C663 VP.n45 B 0.034581f
C664 VP.n46 B 0.034581f
C665 VP.n47 B 0.023996f
C666 VP.n48 B 0.029947f
C667 VP.n49 B 1.20986f
C668 VP.t4 B 1.95864f
C669 VP.n50 B 0.764192f
C670 VP.n51 B 1.22202f
C671 VP.n52 B 0.029947f
C672 VP.n53 B 0.018554f
C673 VP.n54 B 0.034581f
C674 VP.n55 B 0.034581f
C675 VP.n56 B 0.029154f
C676 VP.n57 B 0.018554f
C677 VP.n58 B 0.018554f
C678 VP.n59 B 0.018554f
C679 VP.n60 B 0.034581f
C680 VP.n61 B 0.034581f
C681 VP.t5 B 1.95864f
C682 VP.n62 B 0.690926f
C683 VP.n63 B 0.026728f
C684 VP.n64 B 0.018554f
C685 VP.n65 B 0.018554f
C686 VP.n66 B 0.018554f
C687 VP.n67 B 0.034581f
C688 VP.n68 B 0.034581f
C689 VP.n69 B 0.027086f
C690 VP.n70 B 0.018554f
C691 VP.n71 B 0.018554f
C692 VP.n72 B 0.018554f
C693 VP.n73 B 0.034581f
C694 VP.n74 B 0.034581f
C695 VP.t6 B 1.95864f
C696 VP.n75 B 0.690926f
C697 VP.n76 B 0.025362f
C698 VP.n77 B 0.018554f
C699 VP.n78 B 0.018554f
C700 VP.n79 B 0.018554f
C701 VP.n80 B 0.034581f
C702 VP.n81 B 0.034581f
C703 VP.n82 B 0.025018f
C704 VP.n83 B 0.018554f
C705 VP.n84 B 0.018554f
C706 VP.n85 B 0.018554f
C707 VP.n86 B 0.034581f
C708 VP.n87 B 0.034581f
C709 VP.n88 B 0.023996f
C710 VP.n89 B 0.029947f
C711 VP.n90 B 0.051456f
.ends

