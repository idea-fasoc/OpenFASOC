* NGSPICE file created from diff_pair_sample_1576.ext - technology: sky130A

.subckt diff_pair_sample_1576 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t0 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=3.5061 pd=18.76 as=1.48335 ps=9.32 w=8.99 l=1.66
X1 B.t11 B.t9 B.t10 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=3.5061 pd=18.76 as=0 ps=0 w=8.99 l=1.66
X2 VTAIL.t14 VP.t1 VDD1.t5 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=1.48335 ps=9.32 w=8.99 l=1.66
X3 VTAIL.t0 VN.t0 VDD2.t7 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=1.48335 ps=9.32 w=8.99 l=1.66
X4 VDD1.t6 VP.t2 VTAIL.t13 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=3.5061 ps=18.76 w=8.99 l=1.66
X5 VDD2.t6 VN.t1 VTAIL.t7 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=1.48335 ps=9.32 w=8.99 l=1.66
X6 VDD2.t5 VN.t2 VTAIL.t1 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=3.5061 ps=18.76 w=8.99 l=1.66
X7 VDD1.t3 VP.t3 VTAIL.t12 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=1.48335 ps=9.32 w=8.99 l=1.66
X8 VDD2.t4 VN.t3 VTAIL.t4 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=3.5061 ps=18.76 w=8.99 l=1.66
X9 B.t8 B.t6 B.t7 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=3.5061 pd=18.76 as=0 ps=0 w=8.99 l=1.66
X10 VTAIL.t6 VN.t4 VDD2.t3 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=3.5061 pd=18.76 as=1.48335 ps=9.32 w=8.99 l=1.66
X11 VDD1.t2 VP.t4 VTAIL.t11 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=1.48335 ps=9.32 w=8.99 l=1.66
X12 VTAIL.t10 VP.t5 VDD1.t1 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=3.5061 pd=18.76 as=1.48335 ps=9.32 w=8.99 l=1.66
X13 VDD2.t2 VN.t5 VTAIL.t2 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=1.48335 ps=9.32 w=8.99 l=1.66
X14 B.t5 B.t3 B.t4 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=3.5061 pd=18.76 as=0 ps=0 w=8.99 l=1.66
X15 VTAIL.t9 VP.t6 VDD1.t7 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=1.48335 ps=9.32 w=8.99 l=1.66
X16 VDD1.t4 VP.t7 VTAIL.t8 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=3.5061 ps=18.76 w=8.99 l=1.66
X17 VTAIL.t3 VN.t6 VDD2.t1 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=1.48335 pd=9.32 as=1.48335 ps=9.32 w=8.99 l=1.66
X18 VTAIL.t5 VN.t7 VDD2.t0 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=3.5061 pd=18.76 as=1.48335 ps=9.32 w=8.99 l=1.66
X19 B.t2 B.t0 B.t1 w_n2960_n2766# sky130_fd_pr__pfet_01v8 ad=3.5061 pd=18.76 as=0 ps=0 w=8.99 l=1.66
R0 VP.n11 VP.t0 162.631
R1 VP.n12 VP.n9 161.3
R2 VP.n14 VP.n13 161.3
R3 VP.n15 VP.n8 161.3
R4 VP.n18 VP.n17 161.3
R5 VP.n19 VP.n7 161.3
R6 VP.n21 VP.n20 161.3
R7 VP.n22 VP.n6 161.3
R8 VP.n44 VP.n0 161.3
R9 VP.n43 VP.n42 161.3
R10 VP.n41 VP.n1 161.3
R11 VP.n40 VP.n39 161.3
R12 VP.n37 VP.n2 161.3
R13 VP.n36 VP.n35 161.3
R14 VP.n34 VP.n3 161.3
R15 VP.n33 VP.n32 161.3
R16 VP.n30 VP.n4 161.3
R17 VP.n29 VP.n28 161.3
R18 VP.n27 VP.n5 161.3
R19 VP.n25 VP.t5 130.518
R20 VP.n31 VP.t4 130.518
R21 VP.n38 VP.t1 130.518
R22 VP.n45 VP.t7 130.518
R23 VP.n23 VP.t2 130.518
R24 VP.n16 VP.t6 130.518
R25 VP.n10 VP.t3 130.518
R26 VP.n26 VP.n25 87.0235
R27 VP.n46 VP.n45 87.0235
R28 VP.n24 VP.n23 87.0235
R29 VP.n11 VP.n10 44.9016
R30 VP.n26 VP.n24 44.2193
R31 VP.n30 VP.n29 41.4647
R32 VP.n43 VP.n1 41.4647
R33 VP.n21 VP.n7 41.4647
R34 VP.n36 VP.n3 40.4934
R35 VP.n37 VP.n36 40.4934
R36 VP.n15 VP.n14 40.4934
R37 VP.n14 VP.n9 40.4934
R38 VP.n29 VP.n5 39.5221
R39 VP.n44 VP.n43 39.5221
R40 VP.n22 VP.n21 39.5221
R41 VP.n32 VP.n30 24.4675
R42 VP.n39 VP.n1 24.4675
R43 VP.n17 VP.n7 24.4675
R44 VP.n31 VP.n3 24.2228
R45 VP.n38 VP.n37 24.2228
R46 VP.n16 VP.n15 24.2228
R47 VP.n10 VP.n9 24.2228
R48 VP.n25 VP.n5 23.7335
R49 VP.n45 VP.n44 23.7335
R50 VP.n23 VP.n22 23.7335
R51 VP.n12 VP.n11 12.6443
R52 VP.n24 VP.n6 0.278367
R53 VP.n27 VP.n26 0.278367
R54 VP.n46 VP.n0 0.278367
R55 VP.n32 VP.n31 0.24517
R56 VP.n39 VP.n38 0.24517
R57 VP.n17 VP.n16 0.24517
R58 VP.n13 VP.n12 0.189894
R59 VP.n13 VP.n8 0.189894
R60 VP.n18 VP.n8 0.189894
R61 VP.n19 VP.n18 0.189894
R62 VP.n20 VP.n19 0.189894
R63 VP.n20 VP.n6 0.189894
R64 VP.n28 VP.n27 0.189894
R65 VP.n28 VP.n4 0.189894
R66 VP.n33 VP.n4 0.189894
R67 VP.n34 VP.n33 0.189894
R68 VP.n35 VP.n34 0.189894
R69 VP.n35 VP.n2 0.189894
R70 VP.n40 VP.n2 0.189894
R71 VP.n41 VP.n40 0.189894
R72 VP.n42 VP.n41 0.189894
R73 VP.n42 VP.n0 0.189894
R74 VP VP.n46 0.153454
R75 VDD1 VDD1.n0 82.4548
R76 VDD1.n3 VDD1.n2 82.341
R77 VDD1.n3 VDD1.n1 82.341
R78 VDD1.n5 VDD1.n4 81.5387
R79 VDD1.n5 VDD1.n3 39.7681
R80 VDD1.n4 VDD1.t7 3.61618
R81 VDD1.n4 VDD1.t6 3.61618
R82 VDD1.n0 VDD1.t0 3.61618
R83 VDD1.n0 VDD1.t3 3.61618
R84 VDD1.n2 VDD1.t5 3.61618
R85 VDD1.n2 VDD1.t4 3.61618
R86 VDD1.n1 VDD1.t1 3.61618
R87 VDD1.n1 VDD1.t2 3.61618
R88 VDD1 VDD1.n5 0.800069
R89 VTAIL.n11 VTAIL.t15 68.4758
R90 VTAIL.n10 VTAIL.t1 68.4758
R91 VTAIL.n7 VTAIL.t5 68.4758
R92 VTAIL.n14 VTAIL.t13 68.4755
R93 VTAIL.n15 VTAIL.t4 68.4755
R94 VTAIL.n2 VTAIL.t6 68.4755
R95 VTAIL.n3 VTAIL.t8 68.4755
R96 VTAIL.n6 VTAIL.t10 68.4755
R97 VTAIL.n13 VTAIL.n12 64.8601
R98 VTAIL.n9 VTAIL.n8 64.8601
R99 VTAIL.n1 VTAIL.n0 64.8598
R100 VTAIL.n5 VTAIL.n4 64.8598
R101 VTAIL.n15 VTAIL.n14 21.8324
R102 VTAIL.n7 VTAIL.n6 21.8324
R103 VTAIL.n0 VTAIL.t2 3.61618
R104 VTAIL.n0 VTAIL.t0 3.61618
R105 VTAIL.n4 VTAIL.t11 3.61618
R106 VTAIL.n4 VTAIL.t14 3.61618
R107 VTAIL.n12 VTAIL.t12 3.61618
R108 VTAIL.n12 VTAIL.t9 3.61618
R109 VTAIL.n8 VTAIL.t7 3.61618
R110 VTAIL.n8 VTAIL.t3 3.61618
R111 VTAIL.n9 VTAIL.n7 1.71602
R112 VTAIL.n10 VTAIL.n9 1.71602
R113 VTAIL.n13 VTAIL.n11 1.71602
R114 VTAIL.n14 VTAIL.n13 1.71602
R115 VTAIL.n6 VTAIL.n5 1.71602
R116 VTAIL.n5 VTAIL.n3 1.71602
R117 VTAIL.n2 VTAIL.n1 1.71602
R118 VTAIL VTAIL.n15 1.65783
R119 VTAIL.n11 VTAIL.n10 0.470328
R120 VTAIL.n3 VTAIL.n2 0.470328
R121 VTAIL VTAIL.n1 0.0586897
R122 B.n327 B.n100 585
R123 B.n326 B.n325 585
R124 B.n324 B.n101 585
R125 B.n323 B.n322 585
R126 B.n321 B.n102 585
R127 B.n320 B.n319 585
R128 B.n318 B.n103 585
R129 B.n317 B.n316 585
R130 B.n315 B.n104 585
R131 B.n314 B.n313 585
R132 B.n312 B.n105 585
R133 B.n311 B.n310 585
R134 B.n309 B.n106 585
R135 B.n308 B.n307 585
R136 B.n306 B.n107 585
R137 B.n305 B.n304 585
R138 B.n303 B.n108 585
R139 B.n302 B.n301 585
R140 B.n300 B.n109 585
R141 B.n299 B.n298 585
R142 B.n297 B.n110 585
R143 B.n296 B.n295 585
R144 B.n294 B.n111 585
R145 B.n293 B.n292 585
R146 B.n291 B.n112 585
R147 B.n290 B.n289 585
R148 B.n288 B.n113 585
R149 B.n287 B.n286 585
R150 B.n285 B.n114 585
R151 B.n284 B.n283 585
R152 B.n282 B.n115 585
R153 B.n281 B.n280 585
R154 B.n279 B.n116 585
R155 B.n278 B.n277 585
R156 B.n273 B.n117 585
R157 B.n272 B.n271 585
R158 B.n270 B.n118 585
R159 B.n269 B.n268 585
R160 B.n267 B.n119 585
R161 B.n266 B.n265 585
R162 B.n264 B.n120 585
R163 B.n263 B.n262 585
R164 B.n260 B.n121 585
R165 B.n259 B.n258 585
R166 B.n257 B.n124 585
R167 B.n256 B.n255 585
R168 B.n254 B.n125 585
R169 B.n253 B.n252 585
R170 B.n251 B.n126 585
R171 B.n250 B.n249 585
R172 B.n248 B.n127 585
R173 B.n247 B.n246 585
R174 B.n245 B.n128 585
R175 B.n244 B.n243 585
R176 B.n242 B.n129 585
R177 B.n241 B.n240 585
R178 B.n239 B.n130 585
R179 B.n238 B.n237 585
R180 B.n236 B.n131 585
R181 B.n235 B.n234 585
R182 B.n233 B.n132 585
R183 B.n232 B.n231 585
R184 B.n230 B.n133 585
R185 B.n229 B.n228 585
R186 B.n227 B.n134 585
R187 B.n226 B.n225 585
R188 B.n224 B.n135 585
R189 B.n223 B.n222 585
R190 B.n221 B.n136 585
R191 B.n220 B.n219 585
R192 B.n218 B.n137 585
R193 B.n217 B.n216 585
R194 B.n215 B.n138 585
R195 B.n214 B.n213 585
R196 B.n212 B.n139 585
R197 B.n329 B.n328 585
R198 B.n330 B.n99 585
R199 B.n332 B.n331 585
R200 B.n333 B.n98 585
R201 B.n335 B.n334 585
R202 B.n336 B.n97 585
R203 B.n338 B.n337 585
R204 B.n339 B.n96 585
R205 B.n341 B.n340 585
R206 B.n342 B.n95 585
R207 B.n344 B.n343 585
R208 B.n345 B.n94 585
R209 B.n347 B.n346 585
R210 B.n348 B.n93 585
R211 B.n350 B.n349 585
R212 B.n351 B.n92 585
R213 B.n353 B.n352 585
R214 B.n354 B.n91 585
R215 B.n356 B.n355 585
R216 B.n357 B.n90 585
R217 B.n359 B.n358 585
R218 B.n360 B.n89 585
R219 B.n362 B.n361 585
R220 B.n363 B.n88 585
R221 B.n365 B.n364 585
R222 B.n366 B.n87 585
R223 B.n368 B.n367 585
R224 B.n369 B.n86 585
R225 B.n371 B.n370 585
R226 B.n372 B.n85 585
R227 B.n374 B.n373 585
R228 B.n375 B.n84 585
R229 B.n377 B.n376 585
R230 B.n378 B.n83 585
R231 B.n380 B.n379 585
R232 B.n381 B.n82 585
R233 B.n383 B.n382 585
R234 B.n384 B.n81 585
R235 B.n386 B.n385 585
R236 B.n387 B.n80 585
R237 B.n389 B.n388 585
R238 B.n390 B.n79 585
R239 B.n392 B.n391 585
R240 B.n393 B.n78 585
R241 B.n395 B.n394 585
R242 B.n396 B.n77 585
R243 B.n398 B.n397 585
R244 B.n399 B.n76 585
R245 B.n401 B.n400 585
R246 B.n402 B.n75 585
R247 B.n404 B.n403 585
R248 B.n405 B.n74 585
R249 B.n407 B.n406 585
R250 B.n408 B.n73 585
R251 B.n410 B.n409 585
R252 B.n411 B.n72 585
R253 B.n413 B.n412 585
R254 B.n414 B.n71 585
R255 B.n416 B.n415 585
R256 B.n417 B.n70 585
R257 B.n419 B.n418 585
R258 B.n420 B.n69 585
R259 B.n422 B.n421 585
R260 B.n423 B.n68 585
R261 B.n425 B.n424 585
R262 B.n426 B.n67 585
R263 B.n428 B.n427 585
R264 B.n429 B.n66 585
R265 B.n431 B.n430 585
R266 B.n432 B.n65 585
R267 B.n434 B.n433 585
R268 B.n435 B.n64 585
R269 B.n437 B.n436 585
R270 B.n438 B.n63 585
R271 B.n440 B.n439 585
R272 B.n441 B.n62 585
R273 B.n556 B.n555 585
R274 B.n554 B.n21 585
R275 B.n553 B.n552 585
R276 B.n551 B.n22 585
R277 B.n550 B.n549 585
R278 B.n548 B.n23 585
R279 B.n547 B.n546 585
R280 B.n545 B.n24 585
R281 B.n544 B.n543 585
R282 B.n542 B.n25 585
R283 B.n541 B.n540 585
R284 B.n539 B.n26 585
R285 B.n538 B.n537 585
R286 B.n536 B.n27 585
R287 B.n535 B.n534 585
R288 B.n533 B.n28 585
R289 B.n532 B.n531 585
R290 B.n530 B.n29 585
R291 B.n529 B.n528 585
R292 B.n527 B.n30 585
R293 B.n526 B.n525 585
R294 B.n524 B.n31 585
R295 B.n523 B.n522 585
R296 B.n521 B.n32 585
R297 B.n520 B.n519 585
R298 B.n518 B.n33 585
R299 B.n517 B.n516 585
R300 B.n515 B.n34 585
R301 B.n514 B.n513 585
R302 B.n512 B.n35 585
R303 B.n511 B.n510 585
R304 B.n509 B.n36 585
R305 B.n508 B.n507 585
R306 B.n505 B.n37 585
R307 B.n504 B.n503 585
R308 B.n502 B.n40 585
R309 B.n501 B.n500 585
R310 B.n499 B.n41 585
R311 B.n498 B.n497 585
R312 B.n496 B.n42 585
R313 B.n495 B.n494 585
R314 B.n493 B.n43 585
R315 B.n491 B.n490 585
R316 B.n489 B.n46 585
R317 B.n488 B.n487 585
R318 B.n486 B.n47 585
R319 B.n485 B.n484 585
R320 B.n483 B.n48 585
R321 B.n482 B.n481 585
R322 B.n480 B.n49 585
R323 B.n479 B.n478 585
R324 B.n477 B.n50 585
R325 B.n476 B.n475 585
R326 B.n474 B.n51 585
R327 B.n473 B.n472 585
R328 B.n471 B.n52 585
R329 B.n470 B.n469 585
R330 B.n468 B.n53 585
R331 B.n467 B.n466 585
R332 B.n465 B.n54 585
R333 B.n464 B.n463 585
R334 B.n462 B.n55 585
R335 B.n461 B.n460 585
R336 B.n459 B.n56 585
R337 B.n458 B.n457 585
R338 B.n456 B.n57 585
R339 B.n455 B.n454 585
R340 B.n453 B.n58 585
R341 B.n452 B.n451 585
R342 B.n450 B.n59 585
R343 B.n449 B.n448 585
R344 B.n447 B.n60 585
R345 B.n446 B.n445 585
R346 B.n444 B.n61 585
R347 B.n443 B.n442 585
R348 B.n557 B.n20 585
R349 B.n559 B.n558 585
R350 B.n560 B.n19 585
R351 B.n562 B.n561 585
R352 B.n563 B.n18 585
R353 B.n565 B.n564 585
R354 B.n566 B.n17 585
R355 B.n568 B.n567 585
R356 B.n569 B.n16 585
R357 B.n571 B.n570 585
R358 B.n572 B.n15 585
R359 B.n574 B.n573 585
R360 B.n575 B.n14 585
R361 B.n577 B.n576 585
R362 B.n578 B.n13 585
R363 B.n580 B.n579 585
R364 B.n581 B.n12 585
R365 B.n583 B.n582 585
R366 B.n584 B.n11 585
R367 B.n586 B.n585 585
R368 B.n587 B.n10 585
R369 B.n589 B.n588 585
R370 B.n590 B.n9 585
R371 B.n592 B.n591 585
R372 B.n593 B.n8 585
R373 B.n595 B.n594 585
R374 B.n596 B.n7 585
R375 B.n598 B.n597 585
R376 B.n599 B.n6 585
R377 B.n601 B.n600 585
R378 B.n602 B.n5 585
R379 B.n604 B.n603 585
R380 B.n605 B.n4 585
R381 B.n607 B.n606 585
R382 B.n608 B.n3 585
R383 B.n610 B.n609 585
R384 B.n611 B.n0 585
R385 B.n2 B.n1 585
R386 B.n158 B.n157 585
R387 B.n160 B.n159 585
R388 B.n161 B.n156 585
R389 B.n163 B.n162 585
R390 B.n164 B.n155 585
R391 B.n166 B.n165 585
R392 B.n167 B.n154 585
R393 B.n169 B.n168 585
R394 B.n170 B.n153 585
R395 B.n172 B.n171 585
R396 B.n173 B.n152 585
R397 B.n175 B.n174 585
R398 B.n176 B.n151 585
R399 B.n178 B.n177 585
R400 B.n179 B.n150 585
R401 B.n181 B.n180 585
R402 B.n182 B.n149 585
R403 B.n184 B.n183 585
R404 B.n185 B.n148 585
R405 B.n187 B.n186 585
R406 B.n188 B.n147 585
R407 B.n190 B.n189 585
R408 B.n191 B.n146 585
R409 B.n193 B.n192 585
R410 B.n194 B.n145 585
R411 B.n196 B.n195 585
R412 B.n197 B.n144 585
R413 B.n199 B.n198 585
R414 B.n200 B.n143 585
R415 B.n202 B.n201 585
R416 B.n203 B.n142 585
R417 B.n205 B.n204 585
R418 B.n206 B.n141 585
R419 B.n208 B.n207 585
R420 B.n209 B.n140 585
R421 B.n211 B.n210 585
R422 B.n210 B.n139 487.695
R423 B.n328 B.n327 487.695
R424 B.n442 B.n441 487.695
R425 B.n557 B.n556 487.695
R426 B.n122 B.t9 336.507
R427 B.n274 B.t6 336.507
R428 B.n44 B.t3 336.507
R429 B.n38 B.t0 336.507
R430 B.n613 B.n612 256.663
R431 B.n612 B.n611 235.042
R432 B.n612 B.n2 235.042
R433 B.n214 B.n139 163.367
R434 B.n215 B.n214 163.367
R435 B.n216 B.n215 163.367
R436 B.n216 B.n137 163.367
R437 B.n220 B.n137 163.367
R438 B.n221 B.n220 163.367
R439 B.n222 B.n221 163.367
R440 B.n222 B.n135 163.367
R441 B.n226 B.n135 163.367
R442 B.n227 B.n226 163.367
R443 B.n228 B.n227 163.367
R444 B.n228 B.n133 163.367
R445 B.n232 B.n133 163.367
R446 B.n233 B.n232 163.367
R447 B.n234 B.n233 163.367
R448 B.n234 B.n131 163.367
R449 B.n238 B.n131 163.367
R450 B.n239 B.n238 163.367
R451 B.n240 B.n239 163.367
R452 B.n240 B.n129 163.367
R453 B.n244 B.n129 163.367
R454 B.n245 B.n244 163.367
R455 B.n246 B.n245 163.367
R456 B.n246 B.n127 163.367
R457 B.n250 B.n127 163.367
R458 B.n251 B.n250 163.367
R459 B.n252 B.n251 163.367
R460 B.n252 B.n125 163.367
R461 B.n256 B.n125 163.367
R462 B.n257 B.n256 163.367
R463 B.n258 B.n257 163.367
R464 B.n258 B.n121 163.367
R465 B.n263 B.n121 163.367
R466 B.n264 B.n263 163.367
R467 B.n265 B.n264 163.367
R468 B.n265 B.n119 163.367
R469 B.n269 B.n119 163.367
R470 B.n270 B.n269 163.367
R471 B.n271 B.n270 163.367
R472 B.n271 B.n117 163.367
R473 B.n278 B.n117 163.367
R474 B.n279 B.n278 163.367
R475 B.n280 B.n279 163.367
R476 B.n280 B.n115 163.367
R477 B.n284 B.n115 163.367
R478 B.n285 B.n284 163.367
R479 B.n286 B.n285 163.367
R480 B.n286 B.n113 163.367
R481 B.n290 B.n113 163.367
R482 B.n291 B.n290 163.367
R483 B.n292 B.n291 163.367
R484 B.n292 B.n111 163.367
R485 B.n296 B.n111 163.367
R486 B.n297 B.n296 163.367
R487 B.n298 B.n297 163.367
R488 B.n298 B.n109 163.367
R489 B.n302 B.n109 163.367
R490 B.n303 B.n302 163.367
R491 B.n304 B.n303 163.367
R492 B.n304 B.n107 163.367
R493 B.n308 B.n107 163.367
R494 B.n309 B.n308 163.367
R495 B.n310 B.n309 163.367
R496 B.n310 B.n105 163.367
R497 B.n314 B.n105 163.367
R498 B.n315 B.n314 163.367
R499 B.n316 B.n315 163.367
R500 B.n316 B.n103 163.367
R501 B.n320 B.n103 163.367
R502 B.n321 B.n320 163.367
R503 B.n322 B.n321 163.367
R504 B.n322 B.n101 163.367
R505 B.n326 B.n101 163.367
R506 B.n327 B.n326 163.367
R507 B.n441 B.n440 163.367
R508 B.n440 B.n63 163.367
R509 B.n436 B.n63 163.367
R510 B.n436 B.n435 163.367
R511 B.n435 B.n434 163.367
R512 B.n434 B.n65 163.367
R513 B.n430 B.n65 163.367
R514 B.n430 B.n429 163.367
R515 B.n429 B.n428 163.367
R516 B.n428 B.n67 163.367
R517 B.n424 B.n67 163.367
R518 B.n424 B.n423 163.367
R519 B.n423 B.n422 163.367
R520 B.n422 B.n69 163.367
R521 B.n418 B.n69 163.367
R522 B.n418 B.n417 163.367
R523 B.n417 B.n416 163.367
R524 B.n416 B.n71 163.367
R525 B.n412 B.n71 163.367
R526 B.n412 B.n411 163.367
R527 B.n411 B.n410 163.367
R528 B.n410 B.n73 163.367
R529 B.n406 B.n73 163.367
R530 B.n406 B.n405 163.367
R531 B.n405 B.n404 163.367
R532 B.n404 B.n75 163.367
R533 B.n400 B.n75 163.367
R534 B.n400 B.n399 163.367
R535 B.n399 B.n398 163.367
R536 B.n398 B.n77 163.367
R537 B.n394 B.n77 163.367
R538 B.n394 B.n393 163.367
R539 B.n393 B.n392 163.367
R540 B.n392 B.n79 163.367
R541 B.n388 B.n79 163.367
R542 B.n388 B.n387 163.367
R543 B.n387 B.n386 163.367
R544 B.n386 B.n81 163.367
R545 B.n382 B.n81 163.367
R546 B.n382 B.n381 163.367
R547 B.n381 B.n380 163.367
R548 B.n380 B.n83 163.367
R549 B.n376 B.n83 163.367
R550 B.n376 B.n375 163.367
R551 B.n375 B.n374 163.367
R552 B.n374 B.n85 163.367
R553 B.n370 B.n85 163.367
R554 B.n370 B.n369 163.367
R555 B.n369 B.n368 163.367
R556 B.n368 B.n87 163.367
R557 B.n364 B.n87 163.367
R558 B.n364 B.n363 163.367
R559 B.n363 B.n362 163.367
R560 B.n362 B.n89 163.367
R561 B.n358 B.n89 163.367
R562 B.n358 B.n357 163.367
R563 B.n357 B.n356 163.367
R564 B.n356 B.n91 163.367
R565 B.n352 B.n91 163.367
R566 B.n352 B.n351 163.367
R567 B.n351 B.n350 163.367
R568 B.n350 B.n93 163.367
R569 B.n346 B.n93 163.367
R570 B.n346 B.n345 163.367
R571 B.n345 B.n344 163.367
R572 B.n344 B.n95 163.367
R573 B.n340 B.n95 163.367
R574 B.n340 B.n339 163.367
R575 B.n339 B.n338 163.367
R576 B.n338 B.n97 163.367
R577 B.n334 B.n97 163.367
R578 B.n334 B.n333 163.367
R579 B.n333 B.n332 163.367
R580 B.n332 B.n99 163.367
R581 B.n328 B.n99 163.367
R582 B.n556 B.n21 163.367
R583 B.n552 B.n21 163.367
R584 B.n552 B.n551 163.367
R585 B.n551 B.n550 163.367
R586 B.n550 B.n23 163.367
R587 B.n546 B.n23 163.367
R588 B.n546 B.n545 163.367
R589 B.n545 B.n544 163.367
R590 B.n544 B.n25 163.367
R591 B.n540 B.n25 163.367
R592 B.n540 B.n539 163.367
R593 B.n539 B.n538 163.367
R594 B.n538 B.n27 163.367
R595 B.n534 B.n27 163.367
R596 B.n534 B.n533 163.367
R597 B.n533 B.n532 163.367
R598 B.n532 B.n29 163.367
R599 B.n528 B.n29 163.367
R600 B.n528 B.n527 163.367
R601 B.n527 B.n526 163.367
R602 B.n526 B.n31 163.367
R603 B.n522 B.n31 163.367
R604 B.n522 B.n521 163.367
R605 B.n521 B.n520 163.367
R606 B.n520 B.n33 163.367
R607 B.n516 B.n33 163.367
R608 B.n516 B.n515 163.367
R609 B.n515 B.n514 163.367
R610 B.n514 B.n35 163.367
R611 B.n510 B.n35 163.367
R612 B.n510 B.n509 163.367
R613 B.n509 B.n508 163.367
R614 B.n508 B.n37 163.367
R615 B.n503 B.n37 163.367
R616 B.n503 B.n502 163.367
R617 B.n502 B.n501 163.367
R618 B.n501 B.n41 163.367
R619 B.n497 B.n41 163.367
R620 B.n497 B.n496 163.367
R621 B.n496 B.n495 163.367
R622 B.n495 B.n43 163.367
R623 B.n490 B.n43 163.367
R624 B.n490 B.n489 163.367
R625 B.n489 B.n488 163.367
R626 B.n488 B.n47 163.367
R627 B.n484 B.n47 163.367
R628 B.n484 B.n483 163.367
R629 B.n483 B.n482 163.367
R630 B.n482 B.n49 163.367
R631 B.n478 B.n49 163.367
R632 B.n478 B.n477 163.367
R633 B.n477 B.n476 163.367
R634 B.n476 B.n51 163.367
R635 B.n472 B.n51 163.367
R636 B.n472 B.n471 163.367
R637 B.n471 B.n470 163.367
R638 B.n470 B.n53 163.367
R639 B.n466 B.n53 163.367
R640 B.n466 B.n465 163.367
R641 B.n465 B.n464 163.367
R642 B.n464 B.n55 163.367
R643 B.n460 B.n55 163.367
R644 B.n460 B.n459 163.367
R645 B.n459 B.n458 163.367
R646 B.n458 B.n57 163.367
R647 B.n454 B.n57 163.367
R648 B.n454 B.n453 163.367
R649 B.n453 B.n452 163.367
R650 B.n452 B.n59 163.367
R651 B.n448 B.n59 163.367
R652 B.n448 B.n447 163.367
R653 B.n447 B.n446 163.367
R654 B.n446 B.n61 163.367
R655 B.n442 B.n61 163.367
R656 B.n558 B.n557 163.367
R657 B.n558 B.n19 163.367
R658 B.n562 B.n19 163.367
R659 B.n563 B.n562 163.367
R660 B.n564 B.n563 163.367
R661 B.n564 B.n17 163.367
R662 B.n568 B.n17 163.367
R663 B.n569 B.n568 163.367
R664 B.n570 B.n569 163.367
R665 B.n570 B.n15 163.367
R666 B.n574 B.n15 163.367
R667 B.n575 B.n574 163.367
R668 B.n576 B.n575 163.367
R669 B.n576 B.n13 163.367
R670 B.n580 B.n13 163.367
R671 B.n581 B.n580 163.367
R672 B.n582 B.n581 163.367
R673 B.n582 B.n11 163.367
R674 B.n586 B.n11 163.367
R675 B.n587 B.n586 163.367
R676 B.n588 B.n587 163.367
R677 B.n588 B.n9 163.367
R678 B.n592 B.n9 163.367
R679 B.n593 B.n592 163.367
R680 B.n594 B.n593 163.367
R681 B.n594 B.n7 163.367
R682 B.n598 B.n7 163.367
R683 B.n599 B.n598 163.367
R684 B.n600 B.n599 163.367
R685 B.n600 B.n5 163.367
R686 B.n604 B.n5 163.367
R687 B.n605 B.n604 163.367
R688 B.n606 B.n605 163.367
R689 B.n606 B.n3 163.367
R690 B.n610 B.n3 163.367
R691 B.n611 B.n610 163.367
R692 B.n157 B.n2 163.367
R693 B.n160 B.n157 163.367
R694 B.n161 B.n160 163.367
R695 B.n162 B.n161 163.367
R696 B.n162 B.n155 163.367
R697 B.n166 B.n155 163.367
R698 B.n167 B.n166 163.367
R699 B.n168 B.n167 163.367
R700 B.n168 B.n153 163.367
R701 B.n172 B.n153 163.367
R702 B.n173 B.n172 163.367
R703 B.n174 B.n173 163.367
R704 B.n174 B.n151 163.367
R705 B.n178 B.n151 163.367
R706 B.n179 B.n178 163.367
R707 B.n180 B.n179 163.367
R708 B.n180 B.n149 163.367
R709 B.n184 B.n149 163.367
R710 B.n185 B.n184 163.367
R711 B.n186 B.n185 163.367
R712 B.n186 B.n147 163.367
R713 B.n190 B.n147 163.367
R714 B.n191 B.n190 163.367
R715 B.n192 B.n191 163.367
R716 B.n192 B.n145 163.367
R717 B.n196 B.n145 163.367
R718 B.n197 B.n196 163.367
R719 B.n198 B.n197 163.367
R720 B.n198 B.n143 163.367
R721 B.n202 B.n143 163.367
R722 B.n203 B.n202 163.367
R723 B.n204 B.n203 163.367
R724 B.n204 B.n141 163.367
R725 B.n208 B.n141 163.367
R726 B.n209 B.n208 163.367
R727 B.n210 B.n209 163.367
R728 B.n274 B.t7 149.601
R729 B.n44 B.t5 149.601
R730 B.n122 B.t10 149.591
R731 B.n38 B.t2 149.591
R732 B.n275 B.t8 111.007
R733 B.n45 B.t4 111.007
R734 B.n123 B.t11 110.998
R735 B.n39 B.t1 110.998
R736 B.n261 B.n123 59.5399
R737 B.n276 B.n275 59.5399
R738 B.n492 B.n45 59.5399
R739 B.n506 B.n39 59.5399
R740 B.n123 B.n122 38.5944
R741 B.n275 B.n274 38.5944
R742 B.n45 B.n44 38.5944
R743 B.n39 B.n38 38.5944
R744 B.n555 B.n20 31.6883
R745 B.n443 B.n62 31.6883
R746 B.n329 B.n100 31.6883
R747 B.n212 B.n211 31.6883
R748 B B.n613 18.0485
R749 B.n559 B.n20 10.6151
R750 B.n560 B.n559 10.6151
R751 B.n561 B.n560 10.6151
R752 B.n561 B.n18 10.6151
R753 B.n565 B.n18 10.6151
R754 B.n566 B.n565 10.6151
R755 B.n567 B.n566 10.6151
R756 B.n567 B.n16 10.6151
R757 B.n571 B.n16 10.6151
R758 B.n572 B.n571 10.6151
R759 B.n573 B.n572 10.6151
R760 B.n573 B.n14 10.6151
R761 B.n577 B.n14 10.6151
R762 B.n578 B.n577 10.6151
R763 B.n579 B.n578 10.6151
R764 B.n579 B.n12 10.6151
R765 B.n583 B.n12 10.6151
R766 B.n584 B.n583 10.6151
R767 B.n585 B.n584 10.6151
R768 B.n585 B.n10 10.6151
R769 B.n589 B.n10 10.6151
R770 B.n590 B.n589 10.6151
R771 B.n591 B.n590 10.6151
R772 B.n591 B.n8 10.6151
R773 B.n595 B.n8 10.6151
R774 B.n596 B.n595 10.6151
R775 B.n597 B.n596 10.6151
R776 B.n597 B.n6 10.6151
R777 B.n601 B.n6 10.6151
R778 B.n602 B.n601 10.6151
R779 B.n603 B.n602 10.6151
R780 B.n603 B.n4 10.6151
R781 B.n607 B.n4 10.6151
R782 B.n608 B.n607 10.6151
R783 B.n609 B.n608 10.6151
R784 B.n609 B.n0 10.6151
R785 B.n555 B.n554 10.6151
R786 B.n554 B.n553 10.6151
R787 B.n553 B.n22 10.6151
R788 B.n549 B.n22 10.6151
R789 B.n549 B.n548 10.6151
R790 B.n548 B.n547 10.6151
R791 B.n547 B.n24 10.6151
R792 B.n543 B.n24 10.6151
R793 B.n543 B.n542 10.6151
R794 B.n542 B.n541 10.6151
R795 B.n541 B.n26 10.6151
R796 B.n537 B.n26 10.6151
R797 B.n537 B.n536 10.6151
R798 B.n536 B.n535 10.6151
R799 B.n535 B.n28 10.6151
R800 B.n531 B.n28 10.6151
R801 B.n531 B.n530 10.6151
R802 B.n530 B.n529 10.6151
R803 B.n529 B.n30 10.6151
R804 B.n525 B.n30 10.6151
R805 B.n525 B.n524 10.6151
R806 B.n524 B.n523 10.6151
R807 B.n523 B.n32 10.6151
R808 B.n519 B.n32 10.6151
R809 B.n519 B.n518 10.6151
R810 B.n518 B.n517 10.6151
R811 B.n517 B.n34 10.6151
R812 B.n513 B.n34 10.6151
R813 B.n513 B.n512 10.6151
R814 B.n512 B.n511 10.6151
R815 B.n511 B.n36 10.6151
R816 B.n507 B.n36 10.6151
R817 B.n505 B.n504 10.6151
R818 B.n504 B.n40 10.6151
R819 B.n500 B.n40 10.6151
R820 B.n500 B.n499 10.6151
R821 B.n499 B.n498 10.6151
R822 B.n498 B.n42 10.6151
R823 B.n494 B.n42 10.6151
R824 B.n494 B.n493 10.6151
R825 B.n491 B.n46 10.6151
R826 B.n487 B.n46 10.6151
R827 B.n487 B.n486 10.6151
R828 B.n486 B.n485 10.6151
R829 B.n485 B.n48 10.6151
R830 B.n481 B.n48 10.6151
R831 B.n481 B.n480 10.6151
R832 B.n480 B.n479 10.6151
R833 B.n479 B.n50 10.6151
R834 B.n475 B.n50 10.6151
R835 B.n475 B.n474 10.6151
R836 B.n474 B.n473 10.6151
R837 B.n473 B.n52 10.6151
R838 B.n469 B.n52 10.6151
R839 B.n469 B.n468 10.6151
R840 B.n468 B.n467 10.6151
R841 B.n467 B.n54 10.6151
R842 B.n463 B.n54 10.6151
R843 B.n463 B.n462 10.6151
R844 B.n462 B.n461 10.6151
R845 B.n461 B.n56 10.6151
R846 B.n457 B.n56 10.6151
R847 B.n457 B.n456 10.6151
R848 B.n456 B.n455 10.6151
R849 B.n455 B.n58 10.6151
R850 B.n451 B.n58 10.6151
R851 B.n451 B.n450 10.6151
R852 B.n450 B.n449 10.6151
R853 B.n449 B.n60 10.6151
R854 B.n445 B.n60 10.6151
R855 B.n445 B.n444 10.6151
R856 B.n444 B.n443 10.6151
R857 B.n439 B.n62 10.6151
R858 B.n439 B.n438 10.6151
R859 B.n438 B.n437 10.6151
R860 B.n437 B.n64 10.6151
R861 B.n433 B.n64 10.6151
R862 B.n433 B.n432 10.6151
R863 B.n432 B.n431 10.6151
R864 B.n431 B.n66 10.6151
R865 B.n427 B.n66 10.6151
R866 B.n427 B.n426 10.6151
R867 B.n426 B.n425 10.6151
R868 B.n425 B.n68 10.6151
R869 B.n421 B.n68 10.6151
R870 B.n421 B.n420 10.6151
R871 B.n420 B.n419 10.6151
R872 B.n419 B.n70 10.6151
R873 B.n415 B.n70 10.6151
R874 B.n415 B.n414 10.6151
R875 B.n414 B.n413 10.6151
R876 B.n413 B.n72 10.6151
R877 B.n409 B.n72 10.6151
R878 B.n409 B.n408 10.6151
R879 B.n408 B.n407 10.6151
R880 B.n407 B.n74 10.6151
R881 B.n403 B.n74 10.6151
R882 B.n403 B.n402 10.6151
R883 B.n402 B.n401 10.6151
R884 B.n401 B.n76 10.6151
R885 B.n397 B.n76 10.6151
R886 B.n397 B.n396 10.6151
R887 B.n396 B.n395 10.6151
R888 B.n395 B.n78 10.6151
R889 B.n391 B.n78 10.6151
R890 B.n391 B.n390 10.6151
R891 B.n390 B.n389 10.6151
R892 B.n389 B.n80 10.6151
R893 B.n385 B.n80 10.6151
R894 B.n385 B.n384 10.6151
R895 B.n384 B.n383 10.6151
R896 B.n383 B.n82 10.6151
R897 B.n379 B.n82 10.6151
R898 B.n379 B.n378 10.6151
R899 B.n378 B.n377 10.6151
R900 B.n377 B.n84 10.6151
R901 B.n373 B.n84 10.6151
R902 B.n373 B.n372 10.6151
R903 B.n372 B.n371 10.6151
R904 B.n371 B.n86 10.6151
R905 B.n367 B.n86 10.6151
R906 B.n367 B.n366 10.6151
R907 B.n366 B.n365 10.6151
R908 B.n365 B.n88 10.6151
R909 B.n361 B.n88 10.6151
R910 B.n361 B.n360 10.6151
R911 B.n360 B.n359 10.6151
R912 B.n359 B.n90 10.6151
R913 B.n355 B.n90 10.6151
R914 B.n355 B.n354 10.6151
R915 B.n354 B.n353 10.6151
R916 B.n353 B.n92 10.6151
R917 B.n349 B.n92 10.6151
R918 B.n349 B.n348 10.6151
R919 B.n348 B.n347 10.6151
R920 B.n347 B.n94 10.6151
R921 B.n343 B.n94 10.6151
R922 B.n343 B.n342 10.6151
R923 B.n342 B.n341 10.6151
R924 B.n341 B.n96 10.6151
R925 B.n337 B.n96 10.6151
R926 B.n337 B.n336 10.6151
R927 B.n336 B.n335 10.6151
R928 B.n335 B.n98 10.6151
R929 B.n331 B.n98 10.6151
R930 B.n331 B.n330 10.6151
R931 B.n330 B.n329 10.6151
R932 B.n158 B.n1 10.6151
R933 B.n159 B.n158 10.6151
R934 B.n159 B.n156 10.6151
R935 B.n163 B.n156 10.6151
R936 B.n164 B.n163 10.6151
R937 B.n165 B.n164 10.6151
R938 B.n165 B.n154 10.6151
R939 B.n169 B.n154 10.6151
R940 B.n170 B.n169 10.6151
R941 B.n171 B.n170 10.6151
R942 B.n171 B.n152 10.6151
R943 B.n175 B.n152 10.6151
R944 B.n176 B.n175 10.6151
R945 B.n177 B.n176 10.6151
R946 B.n177 B.n150 10.6151
R947 B.n181 B.n150 10.6151
R948 B.n182 B.n181 10.6151
R949 B.n183 B.n182 10.6151
R950 B.n183 B.n148 10.6151
R951 B.n187 B.n148 10.6151
R952 B.n188 B.n187 10.6151
R953 B.n189 B.n188 10.6151
R954 B.n189 B.n146 10.6151
R955 B.n193 B.n146 10.6151
R956 B.n194 B.n193 10.6151
R957 B.n195 B.n194 10.6151
R958 B.n195 B.n144 10.6151
R959 B.n199 B.n144 10.6151
R960 B.n200 B.n199 10.6151
R961 B.n201 B.n200 10.6151
R962 B.n201 B.n142 10.6151
R963 B.n205 B.n142 10.6151
R964 B.n206 B.n205 10.6151
R965 B.n207 B.n206 10.6151
R966 B.n207 B.n140 10.6151
R967 B.n211 B.n140 10.6151
R968 B.n213 B.n212 10.6151
R969 B.n213 B.n138 10.6151
R970 B.n217 B.n138 10.6151
R971 B.n218 B.n217 10.6151
R972 B.n219 B.n218 10.6151
R973 B.n219 B.n136 10.6151
R974 B.n223 B.n136 10.6151
R975 B.n224 B.n223 10.6151
R976 B.n225 B.n224 10.6151
R977 B.n225 B.n134 10.6151
R978 B.n229 B.n134 10.6151
R979 B.n230 B.n229 10.6151
R980 B.n231 B.n230 10.6151
R981 B.n231 B.n132 10.6151
R982 B.n235 B.n132 10.6151
R983 B.n236 B.n235 10.6151
R984 B.n237 B.n236 10.6151
R985 B.n237 B.n130 10.6151
R986 B.n241 B.n130 10.6151
R987 B.n242 B.n241 10.6151
R988 B.n243 B.n242 10.6151
R989 B.n243 B.n128 10.6151
R990 B.n247 B.n128 10.6151
R991 B.n248 B.n247 10.6151
R992 B.n249 B.n248 10.6151
R993 B.n249 B.n126 10.6151
R994 B.n253 B.n126 10.6151
R995 B.n254 B.n253 10.6151
R996 B.n255 B.n254 10.6151
R997 B.n255 B.n124 10.6151
R998 B.n259 B.n124 10.6151
R999 B.n260 B.n259 10.6151
R1000 B.n262 B.n120 10.6151
R1001 B.n266 B.n120 10.6151
R1002 B.n267 B.n266 10.6151
R1003 B.n268 B.n267 10.6151
R1004 B.n268 B.n118 10.6151
R1005 B.n272 B.n118 10.6151
R1006 B.n273 B.n272 10.6151
R1007 B.n277 B.n273 10.6151
R1008 B.n281 B.n116 10.6151
R1009 B.n282 B.n281 10.6151
R1010 B.n283 B.n282 10.6151
R1011 B.n283 B.n114 10.6151
R1012 B.n287 B.n114 10.6151
R1013 B.n288 B.n287 10.6151
R1014 B.n289 B.n288 10.6151
R1015 B.n289 B.n112 10.6151
R1016 B.n293 B.n112 10.6151
R1017 B.n294 B.n293 10.6151
R1018 B.n295 B.n294 10.6151
R1019 B.n295 B.n110 10.6151
R1020 B.n299 B.n110 10.6151
R1021 B.n300 B.n299 10.6151
R1022 B.n301 B.n300 10.6151
R1023 B.n301 B.n108 10.6151
R1024 B.n305 B.n108 10.6151
R1025 B.n306 B.n305 10.6151
R1026 B.n307 B.n306 10.6151
R1027 B.n307 B.n106 10.6151
R1028 B.n311 B.n106 10.6151
R1029 B.n312 B.n311 10.6151
R1030 B.n313 B.n312 10.6151
R1031 B.n313 B.n104 10.6151
R1032 B.n317 B.n104 10.6151
R1033 B.n318 B.n317 10.6151
R1034 B.n319 B.n318 10.6151
R1035 B.n319 B.n102 10.6151
R1036 B.n323 B.n102 10.6151
R1037 B.n324 B.n323 10.6151
R1038 B.n325 B.n324 10.6151
R1039 B.n325 B.n100 10.6151
R1040 B.n613 B.n0 8.11757
R1041 B.n613 B.n1 8.11757
R1042 B.n506 B.n505 6.5566
R1043 B.n493 B.n492 6.5566
R1044 B.n262 B.n261 6.5566
R1045 B.n277 B.n276 6.5566
R1046 B.n507 B.n506 4.05904
R1047 B.n492 B.n491 4.05904
R1048 B.n261 B.n260 4.05904
R1049 B.n276 B.n116 4.05904
R1050 VN.n5 VN.t4 162.631
R1051 VN.n24 VN.t2 162.631
R1052 VN.n35 VN.n19 161.3
R1053 VN.n34 VN.n33 161.3
R1054 VN.n32 VN.n20 161.3
R1055 VN.n31 VN.n30 161.3
R1056 VN.n28 VN.n21 161.3
R1057 VN.n27 VN.n26 161.3
R1058 VN.n25 VN.n22 161.3
R1059 VN.n16 VN.n0 161.3
R1060 VN.n15 VN.n14 161.3
R1061 VN.n13 VN.n1 161.3
R1062 VN.n12 VN.n11 161.3
R1063 VN.n9 VN.n2 161.3
R1064 VN.n8 VN.n7 161.3
R1065 VN.n6 VN.n3 161.3
R1066 VN.n4 VN.t5 130.518
R1067 VN.n10 VN.t0 130.518
R1068 VN.n17 VN.t3 130.518
R1069 VN.n23 VN.t6 130.518
R1070 VN.n29 VN.t1 130.518
R1071 VN.n36 VN.t7 130.518
R1072 VN.n18 VN.n17 87.0235
R1073 VN.n37 VN.n36 87.0235
R1074 VN.n5 VN.n4 44.9016
R1075 VN.n24 VN.n23 44.9016
R1076 VN VN.n37 44.4982
R1077 VN.n15 VN.n1 41.4647
R1078 VN.n34 VN.n20 41.4647
R1079 VN.n8 VN.n3 40.4934
R1080 VN.n9 VN.n8 40.4934
R1081 VN.n27 VN.n22 40.4934
R1082 VN.n28 VN.n27 40.4934
R1083 VN.n16 VN.n15 39.5221
R1084 VN.n35 VN.n34 39.5221
R1085 VN.n11 VN.n1 24.4675
R1086 VN.n30 VN.n20 24.4675
R1087 VN.n4 VN.n3 24.2228
R1088 VN.n10 VN.n9 24.2228
R1089 VN.n23 VN.n22 24.2228
R1090 VN.n29 VN.n28 24.2228
R1091 VN.n17 VN.n16 23.7335
R1092 VN.n36 VN.n35 23.7335
R1093 VN.n25 VN.n24 12.6443
R1094 VN.n6 VN.n5 12.6443
R1095 VN.n37 VN.n19 0.278367
R1096 VN.n18 VN.n0 0.278367
R1097 VN.n11 VN.n10 0.24517
R1098 VN.n30 VN.n29 0.24517
R1099 VN.n33 VN.n19 0.189894
R1100 VN.n33 VN.n32 0.189894
R1101 VN.n32 VN.n31 0.189894
R1102 VN.n31 VN.n21 0.189894
R1103 VN.n26 VN.n21 0.189894
R1104 VN.n26 VN.n25 0.189894
R1105 VN.n7 VN.n6 0.189894
R1106 VN.n7 VN.n2 0.189894
R1107 VN.n12 VN.n2 0.189894
R1108 VN.n13 VN.n12 0.189894
R1109 VN.n14 VN.n13 0.189894
R1110 VN.n14 VN.n0 0.189894
R1111 VN VN.n18 0.153454
R1112 VDD2.n2 VDD2.n1 82.341
R1113 VDD2.n2 VDD2.n0 82.341
R1114 VDD2 VDD2.n5 82.3383
R1115 VDD2.n4 VDD2.n3 81.5389
R1116 VDD2.n4 VDD2.n2 39.1851
R1117 VDD2.n5 VDD2.t1 3.61618
R1118 VDD2.n5 VDD2.t5 3.61618
R1119 VDD2.n3 VDD2.t0 3.61618
R1120 VDD2.n3 VDD2.t6 3.61618
R1121 VDD2.n1 VDD2.t7 3.61618
R1122 VDD2.n1 VDD2.t4 3.61618
R1123 VDD2.n0 VDD2.t3 3.61618
R1124 VDD2.n0 VDD2.t2 3.61618
R1125 VDD2 VDD2.n4 0.916448
C0 VTAIL VN 6.16672f
C1 B VP 1.60558f
C2 VDD2 VN 5.95825f
C3 VDD1 VN 0.149536f
C4 w_n2960_n2766# VP 6.10555f
C5 VTAIL B 3.579f
C6 B VDD2 1.34876f
C7 VTAIL w_n2960_n2766# 3.45121f
C8 B VDD1 1.28231f
C9 w_n2960_n2766# VDD2 1.63323f
C10 w_n2960_n2766# VDD1 1.55795f
C11 VTAIL VP 6.18083f
C12 B VN 0.971068f
C13 VDD2 VP 0.419153f
C14 w_n2960_n2766# VN 5.72405f
C15 VDD1 VP 6.22695f
C16 VTAIL VDD2 7.04042f
C17 VTAIL VDD1 6.99231f
C18 B w_n2960_n2766# 7.83192f
C19 VN VP 5.95995f
C20 VDD1 VDD2 1.28497f
C21 VDD2 VSUBS 1.451755f
C22 VDD1 VSUBS 1.931525f
C23 VTAIL VSUBS 1.0087f
C24 VN VSUBS 5.46525f
C25 VP VSUBS 2.519614f
C26 B VSUBS 3.699082f
C27 w_n2960_n2766# VSUBS 0.101339p
C28 VDD2.t3 VSUBS 0.176024f
C29 VDD2.t2 VSUBS 0.176024f
C30 VDD2.n0 VSUBS 1.31289f
C31 VDD2.t7 VSUBS 0.176024f
C32 VDD2.t4 VSUBS 0.176024f
C33 VDD2.n1 VSUBS 1.31289f
C34 VDD2.n2 VSUBS 2.97718f
C35 VDD2.t0 VSUBS 0.176024f
C36 VDD2.t6 VSUBS 0.176024f
C37 VDD2.n3 VSUBS 1.30663f
C38 VDD2.n4 VSUBS 2.59652f
C39 VDD2.t1 VSUBS 0.176024f
C40 VDD2.t5 VSUBS 0.176024f
C41 VDD2.n5 VSUBS 1.31286f
C42 VN.n0 VSUBS 0.05206f
C43 VN.t3 VSUBS 1.59022f
C44 VN.n1 VSUBS 0.07806f
C45 VN.n2 VSUBS 0.039487f
C46 VN.t0 VSUBS 1.59022f
C47 VN.n3 VSUBS 0.078116f
C48 VN.t4 VSUBS 1.74036f
C49 VN.t5 VSUBS 1.59022f
C50 VN.n4 VSUBS 0.689151f
C51 VN.n5 VSUBS 0.676838f
C52 VN.n6 VSUBS 0.28388f
C53 VN.n7 VSUBS 0.039487f
C54 VN.n8 VSUBS 0.031922f
C55 VN.n9 VSUBS 0.078116f
C56 VN.n10 VSUBS 0.586815f
C57 VN.n11 VSUBS 0.037622f
C58 VN.n12 VSUBS 0.039487f
C59 VN.n13 VSUBS 0.039487f
C60 VN.n14 VSUBS 0.039487f
C61 VN.n15 VSUBS 0.031973f
C62 VN.n16 VSUBS 0.077759f
C63 VN.n17 VSUBS 0.696336f
C64 VN.n18 VSUBS 0.041734f
C65 VN.n19 VSUBS 0.05206f
C66 VN.t7 VSUBS 1.59022f
C67 VN.n20 VSUBS 0.07806f
C68 VN.n21 VSUBS 0.039487f
C69 VN.t1 VSUBS 1.59022f
C70 VN.n22 VSUBS 0.078116f
C71 VN.t2 VSUBS 1.74036f
C72 VN.t6 VSUBS 1.59022f
C73 VN.n23 VSUBS 0.689151f
C74 VN.n24 VSUBS 0.676838f
C75 VN.n25 VSUBS 0.28388f
C76 VN.n26 VSUBS 0.039487f
C77 VN.n27 VSUBS 0.031922f
C78 VN.n28 VSUBS 0.078116f
C79 VN.n29 VSUBS 0.586815f
C80 VN.n30 VSUBS 0.037622f
C81 VN.n31 VSUBS 0.039487f
C82 VN.n32 VSUBS 0.039487f
C83 VN.n33 VSUBS 0.039487f
C84 VN.n34 VSUBS 0.031973f
C85 VN.n35 VSUBS 0.077759f
C86 VN.n36 VSUBS 0.696336f
C87 VN.n37 VSUBS 1.82076f
C88 B.n0 VSUBS 0.006847f
C89 B.n1 VSUBS 0.006847f
C90 B.n2 VSUBS 0.010127f
C91 B.n3 VSUBS 0.00776f
C92 B.n4 VSUBS 0.00776f
C93 B.n5 VSUBS 0.00776f
C94 B.n6 VSUBS 0.00776f
C95 B.n7 VSUBS 0.00776f
C96 B.n8 VSUBS 0.00776f
C97 B.n9 VSUBS 0.00776f
C98 B.n10 VSUBS 0.00776f
C99 B.n11 VSUBS 0.00776f
C100 B.n12 VSUBS 0.00776f
C101 B.n13 VSUBS 0.00776f
C102 B.n14 VSUBS 0.00776f
C103 B.n15 VSUBS 0.00776f
C104 B.n16 VSUBS 0.00776f
C105 B.n17 VSUBS 0.00776f
C106 B.n18 VSUBS 0.00776f
C107 B.n19 VSUBS 0.00776f
C108 B.n20 VSUBS 0.017492f
C109 B.n21 VSUBS 0.00776f
C110 B.n22 VSUBS 0.00776f
C111 B.n23 VSUBS 0.00776f
C112 B.n24 VSUBS 0.00776f
C113 B.n25 VSUBS 0.00776f
C114 B.n26 VSUBS 0.00776f
C115 B.n27 VSUBS 0.00776f
C116 B.n28 VSUBS 0.00776f
C117 B.n29 VSUBS 0.00776f
C118 B.n30 VSUBS 0.00776f
C119 B.n31 VSUBS 0.00776f
C120 B.n32 VSUBS 0.00776f
C121 B.n33 VSUBS 0.00776f
C122 B.n34 VSUBS 0.00776f
C123 B.n35 VSUBS 0.00776f
C124 B.n36 VSUBS 0.00776f
C125 B.n37 VSUBS 0.00776f
C126 B.t1 VSUBS 0.313202f
C127 B.t2 VSUBS 0.329689f
C128 B.t0 VSUBS 0.74378f
C129 B.n38 VSUBS 0.158773f
C130 B.n39 VSUBS 0.074975f
C131 B.n40 VSUBS 0.00776f
C132 B.n41 VSUBS 0.00776f
C133 B.n42 VSUBS 0.00776f
C134 B.n43 VSUBS 0.00776f
C135 B.t4 VSUBS 0.313198f
C136 B.t5 VSUBS 0.329686f
C137 B.t3 VSUBS 0.74378f
C138 B.n44 VSUBS 0.158777f
C139 B.n45 VSUBS 0.074978f
C140 B.n46 VSUBS 0.00776f
C141 B.n47 VSUBS 0.00776f
C142 B.n48 VSUBS 0.00776f
C143 B.n49 VSUBS 0.00776f
C144 B.n50 VSUBS 0.00776f
C145 B.n51 VSUBS 0.00776f
C146 B.n52 VSUBS 0.00776f
C147 B.n53 VSUBS 0.00776f
C148 B.n54 VSUBS 0.00776f
C149 B.n55 VSUBS 0.00776f
C150 B.n56 VSUBS 0.00776f
C151 B.n57 VSUBS 0.00776f
C152 B.n58 VSUBS 0.00776f
C153 B.n59 VSUBS 0.00776f
C154 B.n60 VSUBS 0.00776f
C155 B.n61 VSUBS 0.00776f
C156 B.n62 VSUBS 0.017492f
C157 B.n63 VSUBS 0.00776f
C158 B.n64 VSUBS 0.00776f
C159 B.n65 VSUBS 0.00776f
C160 B.n66 VSUBS 0.00776f
C161 B.n67 VSUBS 0.00776f
C162 B.n68 VSUBS 0.00776f
C163 B.n69 VSUBS 0.00776f
C164 B.n70 VSUBS 0.00776f
C165 B.n71 VSUBS 0.00776f
C166 B.n72 VSUBS 0.00776f
C167 B.n73 VSUBS 0.00776f
C168 B.n74 VSUBS 0.00776f
C169 B.n75 VSUBS 0.00776f
C170 B.n76 VSUBS 0.00776f
C171 B.n77 VSUBS 0.00776f
C172 B.n78 VSUBS 0.00776f
C173 B.n79 VSUBS 0.00776f
C174 B.n80 VSUBS 0.00776f
C175 B.n81 VSUBS 0.00776f
C176 B.n82 VSUBS 0.00776f
C177 B.n83 VSUBS 0.00776f
C178 B.n84 VSUBS 0.00776f
C179 B.n85 VSUBS 0.00776f
C180 B.n86 VSUBS 0.00776f
C181 B.n87 VSUBS 0.00776f
C182 B.n88 VSUBS 0.00776f
C183 B.n89 VSUBS 0.00776f
C184 B.n90 VSUBS 0.00776f
C185 B.n91 VSUBS 0.00776f
C186 B.n92 VSUBS 0.00776f
C187 B.n93 VSUBS 0.00776f
C188 B.n94 VSUBS 0.00776f
C189 B.n95 VSUBS 0.00776f
C190 B.n96 VSUBS 0.00776f
C191 B.n97 VSUBS 0.00776f
C192 B.n98 VSUBS 0.00776f
C193 B.n99 VSUBS 0.00776f
C194 B.n100 VSUBS 0.01717f
C195 B.n101 VSUBS 0.00776f
C196 B.n102 VSUBS 0.00776f
C197 B.n103 VSUBS 0.00776f
C198 B.n104 VSUBS 0.00776f
C199 B.n105 VSUBS 0.00776f
C200 B.n106 VSUBS 0.00776f
C201 B.n107 VSUBS 0.00776f
C202 B.n108 VSUBS 0.00776f
C203 B.n109 VSUBS 0.00776f
C204 B.n110 VSUBS 0.00776f
C205 B.n111 VSUBS 0.00776f
C206 B.n112 VSUBS 0.00776f
C207 B.n113 VSUBS 0.00776f
C208 B.n114 VSUBS 0.00776f
C209 B.n115 VSUBS 0.00776f
C210 B.n116 VSUBS 0.005364f
C211 B.n117 VSUBS 0.00776f
C212 B.n118 VSUBS 0.00776f
C213 B.n119 VSUBS 0.00776f
C214 B.n120 VSUBS 0.00776f
C215 B.n121 VSUBS 0.00776f
C216 B.t11 VSUBS 0.313202f
C217 B.t10 VSUBS 0.329689f
C218 B.t9 VSUBS 0.74378f
C219 B.n122 VSUBS 0.158773f
C220 B.n123 VSUBS 0.074975f
C221 B.n124 VSUBS 0.00776f
C222 B.n125 VSUBS 0.00776f
C223 B.n126 VSUBS 0.00776f
C224 B.n127 VSUBS 0.00776f
C225 B.n128 VSUBS 0.00776f
C226 B.n129 VSUBS 0.00776f
C227 B.n130 VSUBS 0.00776f
C228 B.n131 VSUBS 0.00776f
C229 B.n132 VSUBS 0.00776f
C230 B.n133 VSUBS 0.00776f
C231 B.n134 VSUBS 0.00776f
C232 B.n135 VSUBS 0.00776f
C233 B.n136 VSUBS 0.00776f
C234 B.n137 VSUBS 0.00776f
C235 B.n138 VSUBS 0.00776f
C236 B.n139 VSUBS 0.018115f
C237 B.n140 VSUBS 0.00776f
C238 B.n141 VSUBS 0.00776f
C239 B.n142 VSUBS 0.00776f
C240 B.n143 VSUBS 0.00776f
C241 B.n144 VSUBS 0.00776f
C242 B.n145 VSUBS 0.00776f
C243 B.n146 VSUBS 0.00776f
C244 B.n147 VSUBS 0.00776f
C245 B.n148 VSUBS 0.00776f
C246 B.n149 VSUBS 0.00776f
C247 B.n150 VSUBS 0.00776f
C248 B.n151 VSUBS 0.00776f
C249 B.n152 VSUBS 0.00776f
C250 B.n153 VSUBS 0.00776f
C251 B.n154 VSUBS 0.00776f
C252 B.n155 VSUBS 0.00776f
C253 B.n156 VSUBS 0.00776f
C254 B.n157 VSUBS 0.00776f
C255 B.n158 VSUBS 0.00776f
C256 B.n159 VSUBS 0.00776f
C257 B.n160 VSUBS 0.00776f
C258 B.n161 VSUBS 0.00776f
C259 B.n162 VSUBS 0.00776f
C260 B.n163 VSUBS 0.00776f
C261 B.n164 VSUBS 0.00776f
C262 B.n165 VSUBS 0.00776f
C263 B.n166 VSUBS 0.00776f
C264 B.n167 VSUBS 0.00776f
C265 B.n168 VSUBS 0.00776f
C266 B.n169 VSUBS 0.00776f
C267 B.n170 VSUBS 0.00776f
C268 B.n171 VSUBS 0.00776f
C269 B.n172 VSUBS 0.00776f
C270 B.n173 VSUBS 0.00776f
C271 B.n174 VSUBS 0.00776f
C272 B.n175 VSUBS 0.00776f
C273 B.n176 VSUBS 0.00776f
C274 B.n177 VSUBS 0.00776f
C275 B.n178 VSUBS 0.00776f
C276 B.n179 VSUBS 0.00776f
C277 B.n180 VSUBS 0.00776f
C278 B.n181 VSUBS 0.00776f
C279 B.n182 VSUBS 0.00776f
C280 B.n183 VSUBS 0.00776f
C281 B.n184 VSUBS 0.00776f
C282 B.n185 VSUBS 0.00776f
C283 B.n186 VSUBS 0.00776f
C284 B.n187 VSUBS 0.00776f
C285 B.n188 VSUBS 0.00776f
C286 B.n189 VSUBS 0.00776f
C287 B.n190 VSUBS 0.00776f
C288 B.n191 VSUBS 0.00776f
C289 B.n192 VSUBS 0.00776f
C290 B.n193 VSUBS 0.00776f
C291 B.n194 VSUBS 0.00776f
C292 B.n195 VSUBS 0.00776f
C293 B.n196 VSUBS 0.00776f
C294 B.n197 VSUBS 0.00776f
C295 B.n198 VSUBS 0.00776f
C296 B.n199 VSUBS 0.00776f
C297 B.n200 VSUBS 0.00776f
C298 B.n201 VSUBS 0.00776f
C299 B.n202 VSUBS 0.00776f
C300 B.n203 VSUBS 0.00776f
C301 B.n204 VSUBS 0.00776f
C302 B.n205 VSUBS 0.00776f
C303 B.n206 VSUBS 0.00776f
C304 B.n207 VSUBS 0.00776f
C305 B.n208 VSUBS 0.00776f
C306 B.n209 VSUBS 0.00776f
C307 B.n210 VSUBS 0.017492f
C308 B.n211 VSUBS 0.017492f
C309 B.n212 VSUBS 0.018115f
C310 B.n213 VSUBS 0.00776f
C311 B.n214 VSUBS 0.00776f
C312 B.n215 VSUBS 0.00776f
C313 B.n216 VSUBS 0.00776f
C314 B.n217 VSUBS 0.00776f
C315 B.n218 VSUBS 0.00776f
C316 B.n219 VSUBS 0.00776f
C317 B.n220 VSUBS 0.00776f
C318 B.n221 VSUBS 0.00776f
C319 B.n222 VSUBS 0.00776f
C320 B.n223 VSUBS 0.00776f
C321 B.n224 VSUBS 0.00776f
C322 B.n225 VSUBS 0.00776f
C323 B.n226 VSUBS 0.00776f
C324 B.n227 VSUBS 0.00776f
C325 B.n228 VSUBS 0.00776f
C326 B.n229 VSUBS 0.00776f
C327 B.n230 VSUBS 0.00776f
C328 B.n231 VSUBS 0.00776f
C329 B.n232 VSUBS 0.00776f
C330 B.n233 VSUBS 0.00776f
C331 B.n234 VSUBS 0.00776f
C332 B.n235 VSUBS 0.00776f
C333 B.n236 VSUBS 0.00776f
C334 B.n237 VSUBS 0.00776f
C335 B.n238 VSUBS 0.00776f
C336 B.n239 VSUBS 0.00776f
C337 B.n240 VSUBS 0.00776f
C338 B.n241 VSUBS 0.00776f
C339 B.n242 VSUBS 0.00776f
C340 B.n243 VSUBS 0.00776f
C341 B.n244 VSUBS 0.00776f
C342 B.n245 VSUBS 0.00776f
C343 B.n246 VSUBS 0.00776f
C344 B.n247 VSUBS 0.00776f
C345 B.n248 VSUBS 0.00776f
C346 B.n249 VSUBS 0.00776f
C347 B.n250 VSUBS 0.00776f
C348 B.n251 VSUBS 0.00776f
C349 B.n252 VSUBS 0.00776f
C350 B.n253 VSUBS 0.00776f
C351 B.n254 VSUBS 0.00776f
C352 B.n255 VSUBS 0.00776f
C353 B.n256 VSUBS 0.00776f
C354 B.n257 VSUBS 0.00776f
C355 B.n258 VSUBS 0.00776f
C356 B.n259 VSUBS 0.00776f
C357 B.n260 VSUBS 0.005364f
C358 B.n261 VSUBS 0.01798f
C359 B.n262 VSUBS 0.006277f
C360 B.n263 VSUBS 0.00776f
C361 B.n264 VSUBS 0.00776f
C362 B.n265 VSUBS 0.00776f
C363 B.n266 VSUBS 0.00776f
C364 B.n267 VSUBS 0.00776f
C365 B.n268 VSUBS 0.00776f
C366 B.n269 VSUBS 0.00776f
C367 B.n270 VSUBS 0.00776f
C368 B.n271 VSUBS 0.00776f
C369 B.n272 VSUBS 0.00776f
C370 B.n273 VSUBS 0.00776f
C371 B.t8 VSUBS 0.313198f
C372 B.t7 VSUBS 0.329686f
C373 B.t6 VSUBS 0.74378f
C374 B.n274 VSUBS 0.158777f
C375 B.n275 VSUBS 0.074978f
C376 B.n276 VSUBS 0.01798f
C377 B.n277 VSUBS 0.006277f
C378 B.n278 VSUBS 0.00776f
C379 B.n279 VSUBS 0.00776f
C380 B.n280 VSUBS 0.00776f
C381 B.n281 VSUBS 0.00776f
C382 B.n282 VSUBS 0.00776f
C383 B.n283 VSUBS 0.00776f
C384 B.n284 VSUBS 0.00776f
C385 B.n285 VSUBS 0.00776f
C386 B.n286 VSUBS 0.00776f
C387 B.n287 VSUBS 0.00776f
C388 B.n288 VSUBS 0.00776f
C389 B.n289 VSUBS 0.00776f
C390 B.n290 VSUBS 0.00776f
C391 B.n291 VSUBS 0.00776f
C392 B.n292 VSUBS 0.00776f
C393 B.n293 VSUBS 0.00776f
C394 B.n294 VSUBS 0.00776f
C395 B.n295 VSUBS 0.00776f
C396 B.n296 VSUBS 0.00776f
C397 B.n297 VSUBS 0.00776f
C398 B.n298 VSUBS 0.00776f
C399 B.n299 VSUBS 0.00776f
C400 B.n300 VSUBS 0.00776f
C401 B.n301 VSUBS 0.00776f
C402 B.n302 VSUBS 0.00776f
C403 B.n303 VSUBS 0.00776f
C404 B.n304 VSUBS 0.00776f
C405 B.n305 VSUBS 0.00776f
C406 B.n306 VSUBS 0.00776f
C407 B.n307 VSUBS 0.00776f
C408 B.n308 VSUBS 0.00776f
C409 B.n309 VSUBS 0.00776f
C410 B.n310 VSUBS 0.00776f
C411 B.n311 VSUBS 0.00776f
C412 B.n312 VSUBS 0.00776f
C413 B.n313 VSUBS 0.00776f
C414 B.n314 VSUBS 0.00776f
C415 B.n315 VSUBS 0.00776f
C416 B.n316 VSUBS 0.00776f
C417 B.n317 VSUBS 0.00776f
C418 B.n318 VSUBS 0.00776f
C419 B.n319 VSUBS 0.00776f
C420 B.n320 VSUBS 0.00776f
C421 B.n321 VSUBS 0.00776f
C422 B.n322 VSUBS 0.00776f
C423 B.n323 VSUBS 0.00776f
C424 B.n324 VSUBS 0.00776f
C425 B.n325 VSUBS 0.00776f
C426 B.n326 VSUBS 0.00776f
C427 B.n327 VSUBS 0.018115f
C428 B.n328 VSUBS 0.017492f
C429 B.n329 VSUBS 0.018437f
C430 B.n330 VSUBS 0.00776f
C431 B.n331 VSUBS 0.00776f
C432 B.n332 VSUBS 0.00776f
C433 B.n333 VSUBS 0.00776f
C434 B.n334 VSUBS 0.00776f
C435 B.n335 VSUBS 0.00776f
C436 B.n336 VSUBS 0.00776f
C437 B.n337 VSUBS 0.00776f
C438 B.n338 VSUBS 0.00776f
C439 B.n339 VSUBS 0.00776f
C440 B.n340 VSUBS 0.00776f
C441 B.n341 VSUBS 0.00776f
C442 B.n342 VSUBS 0.00776f
C443 B.n343 VSUBS 0.00776f
C444 B.n344 VSUBS 0.00776f
C445 B.n345 VSUBS 0.00776f
C446 B.n346 VSUBS 0.00776f
C447 B.n347 VSUBS 0.00776f
C448 B.n348 VSUBS 0.00776f
C449 B.n349 VSUBS 0.00776f
C450 B.n350 VSUBS 0.00776f
C451 B.n351 VSUBS 0.00776f
C452 B.n352 VSUBS 0.00776f
C453 B.n353 VSUBS 0.00776f
C454 B.n354 VSUBS 0.00776f
C455 B.n355 VSUBS 0.00776f
C456 B.n356 VSUBS 0.00776f
C457 B.n357 VSUBS 0.00776f
C458 B.n358 VSUBS 0.00776f
C459 B.n359 VSUBS 0.00776f
C460 B.n360 VSUBS 0.00776f
C461 B.n361 VSUBS 0.00776f
C462 B.n362 VSUBS 0.00776f
C463 B.n363 VSUBS 0.00776f
C464 B.n364 VSUBS 0.00776f
C465 B.n365 VSUBS 0.00776f
C466 B.n366 VSUBS 0.00776f
C467 B.n367 VSUBS 0.00776f
C468 B.n368 VSUBS 0.00776f
C469 B.n369 VSUBS 0.00776f
C470 B.n370 VSUBS 0.00776f
C471 B.n371 VSUBS 0.00776f
C472 B.n372 VSUBS 0.00776f
C473 B.n373 VSUBS 0.00776f
C474 B.n374 VSUBS 0.00776f
C475 B.n375 VSUBS 0.00776f
C476 B.n376 VSUBS 0.00776f
C477 B.n377 VSUBS 0.00776f
C478 B.n378 VSUBS 0.00776f
C479 B.n379 VSUBS 0.00776f
C480 B.n380 VSUBS 0.00776f
C481 B.n381 VSUBS 0.00776f
C482 B.n382 VSUBS 0.00776f
C483 B.n383 VSUBS 0.00776f
C484 B.n384 VSUBS 0.00776f
C485 B.n385 VSUBS 0.00776f
C486 B.n386 VSUBS 0.00776f
C487 B.n387 VSUBS 0.00776f
C488 B.n388 VSUBS 0.00776f
C489 B.n389 VSUBS 0.00776f
C490 B.n390 VSUBS 0.00776f
C491 B.n391 VSUBS 0.00776f
C492 B.n392 VSUBS 0.00776f
C493 B.n393 VSUBS 0.00776f
C494 B.n394 VSUBS 0.00776f
C495 B.n395 VSUBS 0.00776f
C496 B.n396 VSUBS 0.00776f
C497 B.n397 VSUBS 0.00776f
C498 B.n398 VSUBS 0.00776f
C499 B.n399 VSUBS 0.00776f
C500 B.n400 VSUBS 0.00776f
C501 B.n401 VSUBS 0.00776f
C502 B.n402 VSUBS 0.00776f
C503 B.n403 VSUBS 0.00776f
C504 B.n404 VSUBS 0.00776f
C505 B.n405 VSUBS 0.00776f
C506 B.n406 VSUBS 0.00776f
C507 B.n407 VSUBS 0.00776f
C508 B.n408 VSUBS 0.00776f
C509 B.n409 VSUBS 0.00776f
C510 B.n410 VSUBS 0.00776f
C511 B.n411 VSUBS 0.00776f
C512 B.n412 VSUBS 0.00776f
C513 B.n413 VSUBS 0.00776f
C514 B.n414 VSUBS 0.00776f
C515 B.n415 VSUBS 0.00776f
C516 B.n416 VSUBS 0.00776f
C517 B.n417 VSUBS 0.00776f
C518 B.n418 VSUBS 0.00776f
C519 B.n419 VSUBS 0.00776f
C520 B.n420 VSUBS 0.00776f
C521 B.n421 VSUBS 0.00776f
C522 B.n422 VSUBS 0.00776f
C523 B.n423 VSUBS 0.00776f
C524 B.n424 VSUBS 0.00776f
C525 B.n425 VSUBS 0.00776f
C526 B.n426 VSUBS 0.00776f
C527 B.n427 VSUBS 0.00776f
C528 B.n428 VSUBS 0.00776f
C529 B.n429 VSUBS 0.00776f
C530 B.n430 VSUBS 0.00776f
C531 B.n431 VSUBS 0.00776f
C532 B.n432 VSUBS 0.00776f
C533 B.n433 VSUBS 0.00776f
C534 B.n434 VSUBS 0.00776f
C535 B.n435 VSUBS 0.00776f
C536 B.n436 VSUBS 0.00776f
C537 B.n437 VSUBS 0.00776f
C538 B.n438 VSUBS 0.00776f
C539 B.n439 VSUBS 0.00776f
C540 B.n440 VSUBS 0.00776f
C541 B.n441 VSUBS 0.017492f
C542 B.n442 VSUBS 0.018115f
C543 B.n443 VSUBS 0.018115f
C544 B.n444 VSUBS 0.00776f
C545 B.n445 VSUBS 0.00776f
C546 B.n446 VSUBS 0.00776f
C547 B.n447 VSUBS 0.00776f
C548 B.n448 VSUBS 0.00776f
C549 B.n449 VSUBS 0.00776f
C550 B.n450 VSUBS 0.00776f
C551 B.n451 VSUBS 0.00776f
C552 B.n452 VSUBS 0.00776f
C553 B.n453 VSUBS 0.00776f
C554 B.n454 VSUBS 0.00776f
C555 B.n455 VSUBS 0.00776f
C556 B.n456 VSUBS 0.00776f
C557 B.n457 VSUBS 0.00776f
C558 B.n458 VSUBS 0.00776f
C559 B.n459 VSUBS 0.00776f
C560 B.n460 VSUBS 0.00776f
C561 B.n461 VSUBS 0.00776f
C562 B.n462 VSUBS 0.00776f
C563 B.n463 VSUBS 0.00776f
C564 B.n464 VSUBS 0.00776f
C565 B.n465 VSUBS 0.00776f
C566 B.n466 VSUBS 0.00776f
C567 B.n467 VSUBS 0.00776f
C568 B.n468 VSUBS 0.00776f
C569 B.n469 VSUBS 0.00776f
C570 B.n470 VSUBS 0.00776f
C571 B.n471 VSUBS 0.00776f
C572 B.n472 VSUBS 0.00776f
C573 B.n473 VSUBS 0.00776f
C574 B.n474 VSUBS 0.00776f
C575 B.n475 VSUBS 0.00776f
C576 B.n476 VSUBS 0.00776f
C577 B.n477 VSUBS 0.00776f
C578 B.n478 VSUBS 0.00776f
C579 B.n479 VSUBS 0.00776f
C580 B.n480 VSUBS 0.00776f
C581 B.n481 VSUBS 0.00776f
C582 B.n482 VSUBS 0.00776f
C583 B.n483 VSUBS 0.00776f
C584 B.n484 VSUBS 0.00776f
C585 B.n485 VSUBS 0.00776f
C586 B.n486 VSUBS 0.00776f
C587 B.n487 VSUBS 0.00776f
C588 B.n488 VSUBS 0.00776f
C589 B.n489 VSUBS 0.00776f
C590 B.n490 VSUBS 0.00776f
C591 B.n491 VSUBS 0.005364f
C592 B.n492 VSUBS 0.01798f
C593 B.n493 VSUBS 0.006277f
C594 B.n494 VSUBS 0.00776f
C595 B.n495 VSUBS 0.00776f
C596 B.n496 VSUBS 0.00776f
C597 B.n497 VSUBS 0.00776f
C598 B.n498 VSUBS 0.00776f
C599 B.n499 VSUBS 0.00776f
C600 B.n500 VSUBS 0.00776f
C601 B.n501 VSUBS 0.00776f
C602 B.n502 VSUBS 0.00776f
C603 B.n503 VSUBS 0.00776f
C604 B.n504 VSUBS 0.00776f
C605 B.n505 VSUBS 0.006277f
C606 B.n506 VSUBS 0.01798f
C607 B.n507 VSUBS 0.005364f
C608 B.n508 VSUBS 0.00776f
C609 B.n509 VSUBS 0.00776f
C610 B.n510 VSUBS 0.00776f
C611 B.n511 VSUBS 0.00776f
C612 B.n512 VSUBS 0.00776f
C613 B.n513 VSUBS 0.00776f
C614 B.n514 VSUBS 0.00776f
C615 B.n515 VSUBS 0.00776f
C616 B.n516 VSUBS 0.00776f
C617 B.n517 VSUBS 0.00776f
C618 B.n518 VSUBS 0.00776f
C619 B.n519 VSUBS 0.00776f
C620 B.n520 VSUBS 0.00776f
C621 B.n521 VSUBS 0.00776f
C622 B.n522 VSUBS 0.00776f
C623 B.n523 VSUBS 0.00776f
C624 B.n524 VSUBS 0.00776f
C625 B.n525 VSUBS 0.00776f
C626 B.n526 VSUBS 0.00776f
C627 B.n527 VSUBS 0.00776f
C628 B.n528 VSUBS 0.00776f
C629 B.n529 VSUBS 0.00776f
C630 B.n530 VSUBS 0.00776f
C631 B.n531 VSUBS 0.00776f
C632 B.n532 VSUBS 0.00776f
C633 B.n533 VSUBS 0.00776f
C634 B.n534 VSUBS 0.00776f
C635 B.n535 VSUBS 0.00776f
C636 B.n536 VSUBS 0.00776f
C637 B.n537 VSUBS 0.00776f
C638 B.n538 VSUBS 0.00776f
C639 B.n539 VSUBS 0.00776f
C640 B.n540 VSUBS 0.00776f
C641 B.n541 VSUBS 0.00776f
C642 B.n542 VSUBS 0.00776f
C643 B.n543 VSUBS 0.00776f
C644 B.n544 VSUBS 0.00776f
C645 B.n545 VSUBS 0.00776f
C646 B.n546 VSUBS 0.00776f
C647 B.n547 VSUBS 0.00776f
C648 B.n548 VSUBS 0.00776f
C649 B.n549 VSUBS 0.00776f
C650 B.n550 VSUBS 0.00776f
C651 B.n551 VSUBS 0.00776f
C652 B.n552 VSUBS 0.00776f
C653 B.n553 VSUBS 0.00776f
C654 B.n554 VSUBS 0.00776f
C655 B.n555 VSUBS 0.018115f
C656 B.n556 VSUBS 0.018115f
C657 B.n557 VSUBS 0.017492f
C658 B.n558 VSUBS 0.00776f
C659 B.n559 VSUBS 0.00776f
C660 B.n560 VSUBS 0.00776f
C661 B.n561 VSUBS 0.00776f
C662 B.n562 VSUBS 0.00776f
C663 B.n563 VSUBS 0.00776f
C664 B.n564 VSUBS 0.00776f
C665 B.n565 VSUBS 0.00776f
C666 B.n566 VSUBS 0.00776f
C667 B.n567 VSUBS 0.00776f
C668 B.n568 VSUBS 0.00776f
C669 B.n569 VSUBS 0.00776f
C670 B.n570 VSUBS 0.00776f
C671 B.n571 VSUBS 0.00776f
C672 B.n572 VSUBS 0.00776f
C673 B.n573 VSUBS 0.00776f
C674 B.n574 VSUBS 0.00776f
C675 B.n575 VSUBS 0.00776f
C676 B.n576 VSUBS 0.00776f
C677 B.n577 VSUBS 0.00776f
C678 B.n578 VSUBS 0.00776f
C679 B.n579 VSUBS 0.00776f
C680 B.n580 VSUBS 0.00776f
C681 B.n581 VSUBS 0.00776f
C682 B.n582 VSUBS 0.00776f
C683 B.n583 VSUBS 0.00776f
C684 B.n584 VSUBS 0.00776f
C685 B.n585 VSUBS 0.00776f
C686 B.n586 VSUBS 0.00776f
C687 B.n587 VSUBS 0.00776f
C688 B.n588 VSUBS 0.00776f
C689 B.n589 VSUBS 0.00776f
C690 B.n590 VSUBS 0.00776f
C691 B.n591 VSUBS 0.00776f
C692 B.n592 VSUBS 0.00776f
C693 B.n593 VSUBS 0.00776f
C694 B.n594 VSUBS 0.00776f
C695 B.n595 VSUBS 0.00776f
C696 B.n596 VSUBS 0.00776f
C697 B.n597 VSUBS 0.00776f
C698 B.n598 VSUBS 0.00776f
C699 B.n599 VSUBS 0.00776f
C700 B.n600 VSUBS 0.00776f
C701 B.n601 VSUBS 0.00776f
C702 B.n602 VSUBS 0.00776f
C703 B.n603 VSUBS 0.00776f
C704 B.n604 VSUBS 0.00776f
C705 B.n605 VSUBS 0.00776f
C706 B.n606 VSUBS 0.00776f
C707 B.n607 VSUBS 0.00776f
C708 B.n608 VSUBS 0.00776f
C709 B.n609 VSUBS 0.00776f
C710 B.n610 VSUBS 0.00776f
C711 B.n611 VSUBS 0.010127f
C712 B.n612 VSUBS 0.010788f
C713 B.n613 VSUBS 0.021453f
C714 VTAIL.t2 VSUBS 0.181941f
C715 VTAIL.t0 VSUBS 0.181941f
C716 VTAIL.n0 VSUBS 1.23716f
C717 VTAIL.n1 VSUBS 0.670762f
C718 VTAIL.t6 VSUBS 1.65145f
C719 VTAIL.n2 VSUBS 0.786651f
C720 VTAIL.t8 VSUBS 1.65145f
C721 VTAIL.n3 VSUBS 0.786651f
C722 VTAIL.t11 VSUBS 0.181941f
C723 VTAIL.t14 VSUBS 0.181941f
C724 VTAIL.n4 VSUBS 1.23716f
C725 VTAIL.n5 VSUBS 0.807529f
C726 VTAIL.t10 VSUBS 1.65145f
C727 VTAIL.n6 VSUBS 1.87689f
C728 VTAIL.t5 VSUBS 1.65145f
C729 VTAIL.n7 VSUBS 1.87688f
C730 VTAIL.t7 VSUBS 0.181941f
C731 VTAIL.t3 VSUBS 0.181941f
C732 VTAIL.n8 VSUBS 1.23717f
C733 VTAIL.n9 VSUBS 0.807524f
C734 VTAIL.t1 VSUBS 1.65145f
C735 VTAIL.n10 VSUBS 0.786646f
C736 VTAIL.t15 VSUBS 1.65145f
C737 VTAIL.n11 VSUBS 0.786646f
C738 VTAIL.t12 VSUBS 0.181941f
C739 VTAIL.t9 VSUBS 0.181941f
C740 VTAIL.n12 VSUBS 1.23717f
C741 VTAIL.n13 VSUBS 0.807524f
C742 VTAIL.t13 VSUBS 1.65144f
C743 VTAIL.n14 VSUBS 1.87689f
C744 VTAIL.t4 VSUBS 1.65145f
C745 VTAIL.n15 VSUBS 1.87208f
C746 VDD1.t0 VSUBS 0.177482f
C747 VDD1.t3 VSUBS 0.177482f
C748 VDD1.n0 VSUBS 1.32475f
C749 VDD1.t1 VSUBS 0.177482f
C750 VDD1.t2 VSUBS 0.177482f
C751 VDD1.n1 VSUBS 1.32377f
C752 VDD1.t5 VSUBS 0.177482f
C753 VDD1.t4 VSUBS 0.177482f
C754 VDD1.n2 VSUBS 1.32377f
C755 VDD1.n3 VSUBS 3.05458f
C756 VDD1.t7 VSUBS 0.177482f
C757 VDD1.t6 VSUBS 0.177482f
C758 VDD1.n4 VSUBS 1.31745f
C759 VDD1.n5 VSUBS 2.64822f
C760 VP.n0 VSUBS 0.053491f
C761 VP.t7 VSUBS 1.63394f
C762 VP.n1 VSUBS 0.080206f
C763 VP.n2 VSUBS 0.040573f
C764 VP.t1 VSUBS 1.63394f
C765 VP.n3 VSUBS 0.080263f
C766 VP.n4 VSUBS 0.040573f
C767 VP.n5 VSUBS 0.079897f
C768 VP.n6 VSUBS 0.053491f
C769 VP.t2 VSUBS 1.63394f
C770 VP.n7 VSUBS 0.080206f
C771 VP.n8 VSUBS 0.040573f
C772 VP.t6 VSUBS 1.63394f
C773 VP.n9 VSUBS 0.080263f
C774 VP.t0 VSUBS 1.7882f
C775 VP.t3 VSUBS 1.63394f
C776 VP.n10 VSUBS 0.708096f
C777 VP.n11 VSUBS 0.695445f
C778 VP.n12 VSUBS 0.291684f
C779 VP.n13 VSUBS 0.040573f
C780 VP.n14 VSUBS 0.032799f
C781 VP.n15 VSUBS 0.080263f
C782 VP.n16 VSUBS 0.602947f
C783 VP.n17 VSUBS 0.038656f
C784 VP.n18 VSUBS 0.040573f
C785 VP.n19 VSUBS 0.040573f
C786 VP.n20 VSUBS 0.040573f
C787 VP.n21 VSUBS 0.032852f
C788 VP.n22 VSUBS 0.079897f
C789 VP.n23 VSUBS 0.715479f
C790 VP.n24 VSUBS 1.84856f
C791 VP.t5 VSUBS 1.63394f
C792 VP.n25 VSUBS 0.715479f
C793 VP.n26 VSUBS 1.88154f
C794 VP.n27 VSUBS 0.053491f
C795 VP.n28 VSUBS 0.040573f
C796 VP.n29 VSUBS 0.032852f
C797 VP.n30 VSUBS 0.080206f
C798 VP.t4 VSUBS 1.63394f
C799 VP.n31 VSUBS 0.602947f
C800 VP.n32 VSUBS 0.038656f
C801 VP.n33 VSUBS 0.040573f
C802 VP.n34 VSUBS 0.040573f
C803 VP.n35 VSUBS 0.040573f
C804 VP.n36 VSUBS 0.032799f
C805 VP.n37 VSUBS 0.080263f
C806 VP.n38 VSUBS 0.602947f
C807 VP.n39 VSUBS 0.038656f
C808 VP.n40 VSUBS 0.040573f
C809 VP.n41 VSUBS 0.040573f
C810 VP.n42 VSUBS 0.040573f
C811 VP.n43 VSUBS 0.032852f
C812 VP.n44 VSUBS 0.079897f
C813 VP.n45 VSUBS 0.715479f
C814 VP.n46 VSUBS 0.042881f
.ends

